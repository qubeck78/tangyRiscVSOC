--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Wed Feb 14 11:10:49 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPADDSUB/data/FP_Add_Sub.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPADDSUB/data/FP_Add_Sub_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
Fkvy9Luzhz5U0QmYihEF0APEWVRqRpqaqFl/UDFn0meHh/NLt+klk8XBqyghCM5irpB3HYbgzK8B
kR5SREmw2XdhTEset7L4SBjY9idMoarm4M/ZNC8D6THHJ7idi/RieUJ/MJoRiPxokHzeQx8eCs6C
wrE5SJe0xcp/K01/zZK+5QYj1YCsknvEnTSJcGqev4ZSi1EOKI2h8UNRRDehc7T4AV6L0CcPd8dG
LYePRn4MWPPeG1NpOaHI/Fowpv51/xe9VoJ3hsuY1Ydwa86mwBY8HMGFLsV5+CmxtUdju0EvYjkJ
5LEqB+IFkbhQ5xgCtlgFinUdzQWyR+YXhSStmA==

`protect encoding=(enctype="base64", line_length=76, bytes=264896)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
aOmeRLQtlVjPF2Z0BRDo6Nso/O26j13YZIYhWF9jT4mAviy2BahPG5gor3oyhAExz71Rx8k7mOK/
ry4TzO4fuuB381e66tjO3mveVRehuKro5K0jDPwgMBqDAHTLPd7qn+JTGtKOl5PAh+aQTWoz9brd
47Rgi/c9t5BTi3Im81qiFJAWHX7+0fGKsol6A1xb44duc0yZWzIC552TNSb51UsTH4H6G9leK89S
5p0hgcTh2M509tJ0fVhc3VtXdpyy6/eZXUwHTiwTVljELLWVmE0c9xsaDp6D/rkmczV826WK7gCt
HefNFgjg4uCMchhZgtNjTwF1lsffBo8qt5AlE+g1/znwyPDMgwZhMo1RssbFlEtOQbnDRvXxztZ9
0dcDf0lJ3y/HOYgxGUyr6UkUnRgVDkos9Dmza2VtPRuYdde5m/fAG9HI2LH0w0M/FHf4dK//Hu44
2bkWYPfr4UQCFpk3d0Mdk+3dqM0GAIU6YUrfZ0OwJH1yjjXPbA/BDV3E+AUeilc3gd2dk+eibbx1
UC4nO/a6P0Y0UHpFOi1tyeo+Z/BXwmFvrf7llpthvd+uTsS/0S1K4Yl2u9g/EtA0nJQUwExBEfOM
1G68U/K3zhFLkqIbOsJaw+3AAQyRQQDOTVCyiMsnUqKGYkF7yU+sgElX6TP2Z8pvrEmQwjxKty+E
RxbnIizaFIKHruvPOUHAClR23vJ8TsNU5yER6Fcg/xd1F2Hb9ZrpxyqNWNVVa6hFVaIVJf7Rb8df
/Pw2HYkcKAor6WnDGNmJl5AVWMlkCxsbHyMApfKDnptPGeAEeIDnGjUOBE7fB9c2UE5uqsJDF2xu
1UJbParhagU5WhfVue4mdlKSA5XOufb+eiQnRpu5WEUK7kMfr45GzFPt5sYBYEK0WRPpnsIjGqYZ
zTaeYU/98EC04CDHAmsy0KXKUCCcp7QZz7h+8v92v2QclozclPFsxjcklTH2DksHdn0E8pT6I6Vq
u9Du6p7eHcao3HMlwy8Js+IBLxeQ7n0cU+/6P65tr00oRUhfU51IOSn9jlhqUqjk3nLILqDesiDs
kpuf4N3VQ6LwQlocvsVEx6yrFmTu6a1RQvWqOm8d456yTTOI9Crs2tBxoSbLXvJsh7iJ9jsaxZu3
/WVVJggkEyFjIc8fcpxlxUPzSl++z/ZdFn5Lq50StOoddg737qn7yEulmR5dLtQ9cndbtAYH2pP2
lMY7S3epCeE6LAZVLX2UjIwncvV1i0iQJpMpcsfYsWttpoQeRzWDyR8x/+7A/RGih0pt/4UtBgP0
eP8at1OqSvePjC0jPebQB0GXitWFOOrCAmC/vQ8JTuaCuKJq5+wE+l/zZzPsKi6o+Nd1Bse8fEnY
TXAWrVwHVlXlokV2hnjMiFPm9KbAiZFvnAeX+RJdv26wrw17pZEtXukf9VZ7+/zk4HErP5YubFPX
dR8Gk3N0da8yAUYqn+7iy8YxZL5nGXBAbYgn00ae7+A3Jt+w4v30Zo8OBpaBRnX8li9E6meyh+D1
FHHINTKLkdo3+BSpiV6ipkFf/Jwyix5Y0utRwRgvbtA2At1bo1rILqsWKqJ36mJNxm/4KQkGXA1k
WYeXlbkerejrVnF7pfwvVDrCeK7S0WgOAHXYKyfJaeiRhkNYPjJi4jnqqoAXv5ZURJ2rEwUNWiL/
A/5Fz1VeIdZglVFMwXopajBYskNqwMQ98CcJ5saQJZQ5nBxcD0ukPhQG3oUmShfWSnfNBfCaZLkr
vVtV0tr8kVUWofli3KerccyqxGMHPYB7LXL3F0lpQNDVJNyJejOrLgwsuWoy3zOE2jB1+H/B1yMe
pcveZBF3e+NblRO8MgBQXykSOWn5ZY2UUlFpj0tK5r6VVgizWNJc2ftfGoA2QfCMubu8tHFy6TGX
Bmns12hzlH1mddtNuvGTymmsvol3kqU8u2E8E49Wfh0GftdlB+vqPYFrpnQT85zVULH3jEHRSXIu
cB1yQ+BcI9DQJW5CkR1SqT+mYWad3ROsA3r3x5KykfZ2wRgzad39Ya809Y5kl0QD9us5uW0Q53xE
uIdk/4c25v1Y80zorlKSRmUMBGJr4LQBNzBcVqX7+7bvaPSSGhST1hSVL9add4yC28o/H2ckuQ6H
x/0ZHdS5i4muZfKExmCm9oHUGf+g0bs48UEGycFRrMZ/Mkd8Q9bQboFjC7IclzQNT6SQE5EhYj8s
weFZ4oVQv7g0YqlQe8nDHg9mjhr00/lquuZZRbviEydAeH6RrbyaDN4PwcG7x+w/yGoaJy2tuF67
Qm+kIsYJOoOb7EcMyiozLx+7MqjRIh3n0WvsBwC7U5z4hHvDZVexRLBWPjhvWC60jV/pgRrqQArt
XydgHQVaR0IiP+BUwjoUhJWDrf0WEWprWQ9jLebQRnY5EUhGM+IfJ1qgqvPVLknT5I2oFYos+uUW
gphSma6fJNC9AyGvnRPMYGo10sCrmx6O87hS1UW7t/kgP5SxOmpkZHbdV5t8RG/iUubEKgwklUxl
HK6LlHZcyspVNnx9ZCiEnRcwP1SXlbJV9vCk8p2me5PdIiN4RidkgPWgO40GL1eobUzAHVDi34kA
gLEojkNZsC7DOMbP8HeSFx8g80I6OrSMoTcsbCDScOE9ydmhgjqBF7sroLC4s7KL1l5VjXiyhegv
7lWPlKtIr1J+3u6gL7FxtFK22j2Hk+kzMIEBpsxN7PCKqDQWO3csPYJYi/p0QnG0Ro8BBAtXNUZO
qfoh2JDnfjkVz3Ev/NB0T5N7Y0tCUAyCNYnWZXOEqk98pmyk5n3ziaNxnZUY8tZNMHlN3MYCaelj
Gp8Bsr/BkYz23GfR0tSzp+RCECmuc8vWv5KSfsddB4eTRW2iPz69Q4wJ3Z80efPkCtbNiz7aJNDg
0wu4mNaIphG9OAgjSiXqF57q53Zgod/zMtNmpBUSbU4mxE5fUVu34T4VdZ6GUfgrsnyQ+DFQ+j2t
Duvh3PNTEqclhUKd5aS1Mk+qtKSMTZ9Ve7WxIU9Mhu3a2vTM0hbbAN1T9Q0Qi4vN3DgnwF+L08cR
CKG/dYyPot1pWW/osnyxRKPVqmdSXVowPtNhAkArhsKlTuhG6vtek6DvmrnPuHtCdv8AjcFbNjTq
6q8/WRAeT8ORK/TtPjXEYpUbdaI0HgKjKClqlUIs//FfndqIWd5498o8/7/IjKI625j+tEoyGhDZ
W2JqZ1icgEeZ/DJq1LtKVVDs1BQtSgcM4dRqfODclSyOukaF1X4LzeH52eJrck89B/8MD3ngO/Su
/SWGSARu44WtjhwYNU1kigS2XQJk0P4NhsomNenkigED/Y/iG/ozGaQH2Q6VqRRpCWpGGSA9SwFl
3ornjybaMdZWWDTjx9Y+PKEhmBWoBFHt8yj3PMcu3fK5Q/r8dN55x76SOtfKUZPK4JjUAOZZ4CmY
pjUwJaECP+8RdB/rGXL0Te5HKDeJL0zK12B96/3zLIcKqeJ9XLghRuI4x5LnBeiZHzap5rlGPDHV
iE6MDYaPMslsjTTjTxboxJxgKqVL62fQohGcmNKhHDYxt4CDsjBjj5ICwTmKaNjoGZO2qPAuP+pm
YXOXbVuVhJFum2Rr8W0Zt+UyECkWAmou+Fn9rXQhUhu+o384kd6uFOoW9n1KypltzpbH8YJgeBpG
USVGbnSIZ5bmQNMuxHh8fyEJGr4SqvG5ss+H1GKjgaG+LPIiQ2JwYt2KsV+SDeFm5NopsRFweLIO
ic7ImhdkCVo6DLazDXTJKfuRDZFOc2LFALtHriy0oPGWHMDk1IEs0j++u/UmHbOB41wk/cUY1rv1
HBYCwNhAacqCP3Zui8FKLOMryMQZZ3Z5cK5GhAsbHgPjK+R4qnu5O/vHmkSM/iS7itFr/XCUyaNI
P+J9rav4OHB1sSLo0xs/S2pIyjVcq8gYS1HFc+k0GxeoMVgqXDIRHT3BhTJanLIE7luaqYDGzCEF
xV+uC0Zk24YsylHRoQcP23Yqgp0WhS7wlgFFpQ5+QRWivo/lDV4OKE43epbf0uUjSqWKfQUMXWjN
QjLVOZCPRxekrwl6lVNbSdxqSeonZBlzmyeNThdfMtLznjCbYVi1OX2QVHYerBrpJ3T+GP5iV5Oz
NqfEEKO5+EuUxZphN4gSUYttA9YY5Ds7B3yapKhhaMwecKvg6DhA/XeTKSejuPRwkLRVe6f35joN
1I8NxKfcCnSH5tleReogkpIyGwGDiTu0iFRla/x686Pd5aIjWKFkJZK/oTIkU009Dj5fATfGL8eP
AlalUrpygaXtNCrN5G6knWEIclLdJRFbdmt+5xOjrBQDsyQfzrerksbDxnDMNtngnpsFoBQxDFZJ
oRgq90ZYj+qdfe/KA65SI9E/PzSzO/Kq2MTvUpbgGIRdk3llllw8rDYlcJi/V2m/1q1fXIc2h34h
PB0I5XNFUA0uTpsn7Qv+zUO5LO0HFOqhyA3W/QMUXG3+FG6tmQS7yrUy4ipbdpN4IlXxi2s5QyHq
GpxHNAbinB8Xn1lgYwn4IQ4EVswZbcP5FDJzQRZu6ZSTkpJS9pqkzNFQ0nEQCWT6H8pUpvns/yqz
+p+kDhr8WKsqF/Z5I1FQ4EL73kFK/ja3QUpU42STAwoaLSL5WrrWWm+Zat48jw0vFAq2wtvPSl9m
syy8fdRY7AeCQPP30mDetqqp5uYc/F5tuxwZfrtOt9vGZxJV5us7SFxukrunOjbk88ZOCoRKdmLj
NucoTBgCb4QI3nmEsm9jW2ncESCWMEabWwGDtO+A+4LC9+T8nwwiB4qtORG64Koe1UGxh3LlA4M7
mCWseD3IwVZdblRPAwYr/ulvPyGKvnLUdZuxrBASO4LdM/pPUn6D15kfW7UA9JqBHnmOo8COcuDn
3Ahd+ZbGX9ZqkMLNJyRGnOGJFwiekGb8ep5F/iWRH933GTPaJp9WwMeM4BJEGgq0OKmFbXJWRfPQ
9gJ/2uaf5bUJ9ZemhRr2guhCuVax7WwZzUj8IoGhi4U76NQ+TTwiYzWAMQpQmItITxD55C4WBQR9
RCc18euykkdt79gMFqPwoP4dC3l0qo2DL3Qc2HGXhSkS0ScesRILhR/5mF7AhszDxvYlNk9e/wDV
Ldd8rKw/GBf5d3/XdB7HDOHggu64iOtSn7ZKk44XwXEYdJbQji3XXwiBREmTatZtLFFkP4wavt72
jTCF+cOirXxyLvKV24diHK+moauPdgNsX3O+5djLfXmS5Plr2+MfWWmAgj7ukZ9rHHwcd/hNssH4
XUr2vL1JMg1rbmi8vk7691x2eVHvMqxA+1WaA+n3TorO9TnM2Ms0j4ZlN5xkcbKILZc5zK+bmj5p
yqQqzWE9QbZTlGuRsWUgVwM6/wFM7u52Sz47T0E1JwKt5xrSdDCzNWc7F2idvfghsqid/ADq8Rp+
Nvo6ovLbYZJMxVlwqrE8W4tzCn1RfXkqgF0lBpshPh2IalV+16wXmhoQIqzd7YpUS3KQget0uglt
0NKeAsUrW3AejbwGEIhdyTy5yo2qzhhJpD/XM7JhmxstSVUKwopV3lUJ6nvx7lG0/oIW2Kf7KvUo
kVhPsA3cL9grwx/2CN7q/yTV7gLJe7ZikE8fDSmu1af+X65K9NDMAVxRKsLtHFiaLcE96vswQVPv
P4mBLECuCaCIhKdNtUixEstfUhU9aOgw7a2WgT2oMan8B3iw3N2W3eb4v0UAlqTHSRnoin1kqZdK
5+d7/6ywSH0VeMSgaJwito1xHT1nGjpTcx5v89jOz2LNHtxM2efG+WHVTlnolCqdMDjWmp3si2ws
4XWUzwzLnQxPpA1lp60aE56N3TfkBWY24d0njydlh9L1QtIO783wXE2iJuFOkGn2IeEOp5mryr2W
erqIZ6PDTeRCFmZzIxv+nnLb32XNr4t1FyIotiisTAOP8YFChqH+o7S/oe2O1kAoVVcwzR/mpr17
1IKP1F72asllLy0Ugd7uTLw0K6fnYi1cR7k+GutotSIeICsyk472waJRhK6z43x3NT2CMdsCiYJz
wdIsy3jBxirLznsNzDKKSJXrSu7e8hYG48OZJCsHGtXGcR1f7ae+0BWHvsaT5XraqchUbwdoyKti
tFmvsqffeMTKOGnMD5HdH3AW7YqJOpW5wS0vAjIq5zQaQo8NFwAJjfagrxVb3eIAyqALMvvw5Ld7
GEuCEdswZMd2h/pb4ImfiEnlznzTvLKF/4+yqhcOuppsBrF7gg+kmf/y+lLjKCs8u2uUFw9o1JEo
yOy58Fm/GrsAo/dURNJEZWm9At/f/ejPwgC1ud1uBvqIs98tSRpbRxTPXZ+lhpEBK8lCPy7UhOfq
9/dBqyb8p3h1hOL0Co/PwuiLc4m/p/4LDZdlCeiW56Srciihm0xU/wxWKmxFetGh+K+o1I2HRqtr
BCVX4vKozJ35WS1hxgvXDtAUxNvAO3QbNJGwuQToPmL16bMGH/ui+HP409a0T27Vd086KTOaZDca
4GZEvzpQ90fuEP/a+GOnf2atuHfMCm2wstTN5p9PwyPCAAlvnn0R2Z/VV3wm1xr8fOaDwVS17bYa
u01xLdXNpqla8nNd9uz4VSOZE6u67opTIYDeuURTl6ddEC53aLfmlktlbsH85ijTHd4UkgDCgwVP
fvQFX7x128UoxIxWIW07u2L/Tiwsf+DXdFBr7RAvhkGZriLtI50s8FUE+Ux4r+V2wxmhTIvZCSaj
YaMxLpvxKRSyXO0dozPlxQ6V0+z9iNtrvtlLNyGN/tjq3U/h7an9gae6z7qCnpnW/0WB8IofyUHb
Y56K+4i5wIYgGb8VMxT86nUxOcmuNhJKZnbQVkJbZVK+6ylh8tCHOztBdOw+Uak54SPxMZGo8YxO
jpVXn15N4DiqWo6yVMYZPHnpAcCvcHbQ0LyhWe4sUDr8m46jk1xbhs7lohBfBI+YoNbjFCQfvCxx
eA+pX1gafVPKVYg+qU+keBz5n+pID9EFnG9qHzC6gbWWq+e0xIopkzKUQtZuTNhknDUxQyFMOUiF
gTqe6AC/Gy94gVQSVbU/LCT7mX3jcpnNK3/fOhRZKbe39xPu4rz6yweF3cjWcSE0gja81pk2y4NI
gT/nKcYRyT8wZOcMdUtbWmZ2XTQBbowZ+VW1e9MtGMWEhqWXgFYiDFaoYoc8Y0cAjKYAiKuTXdTk
Ab/i8FYStLJSYIE8992ZK41PcwXUhhyjKsn3d3smQKOEKXtGVdYN41MCNaBJeTp5AOH3hyxU0kGI
U5A2WtnMajfmamZ5fLENHAB/S+AzXkN1tQA3TCo9NPDQvuVanQdwcqANuMapcntWoCWoexQKun0m
uCedsTzx02qu2jnhme1Nd1dklAG0u5Ws9rHVtRpPVT0I1U7tnQz/CUp7v/bP1zotqfjmmh+v6T0S
byMhxZEn9T6ychfjCgNUDbgFpAJtzCHETdbqkFkfrivjI0HN+vUdmA6zfrMGCpgpmJWl1RidYrJH
b4BMnf90ekN5Q23SCJh2MpxXNUngvBxJjrQfpo6W65mDUfw9TLSAdIvmq6tViukamim6dCTaFuii
SQIvLhGGAuO8vM1LTRZTRG0xqgRuKXH3XQDl3/zfooe9NE/v+n2S23VfRjq2BUBWElw7hPW9e/ZX
ygLYNfN4591wuQ/4ISkAOx7gtpO24asjQ1aw7Ln5KXX7rIV/RafmsI85DQ1/kteuMTiA4TnvftNW
B8dAs05GaOMMvK14uVU9xAGdEPROLHIjgeJvxEwTBh36LkJm51mR4LeRwWm43Gg7LHHtYWKuY5Wu
IiGtPU6l5oicvoAuGUSmwbSQCBIt/b/Wqv0CLUbQVbFVX0VD++HFqcZ5mdfL4zbQzQxVds5zlmgA
O2V26dKjgDDoArhaJ9keZ6j1xGY8juGhnz/USvCut5LkXbb3Kblmab0lP+TarIS5viiZpKXSlIen
45bc9j3Uxi9nPIA3iAZB5YJUqbTsaVy9g+ZI8eTDw9Z/vDD/27N3ca5ABQQZfh0vJLC0brpj2IHf
M9vH79HLc5xDqPkIvmwDQipsqL1VNDvGvCKGIf1fPdtnG8y0Cp64uE87deuKkLJPSKof9F6eTxHE
xf0NG0ScSIuyCuIWh3IEpMLz51sRu9hw546qbnPkR5obKYhTNYIeNJ3YtVjiQlUZcbEcW+r+30PB
a0HpjE1HhujPJr91eSkkHS00lEIzTb4Mr+2Mce1F1bL4m3algaAljFgZmFWZMsLYHoT2JBLZp5ZK
a2k85Npemu/O1gFIeRRElHgJCIHaXVD1DUSTCvPl38/gQk57iNmF2tKQWgq66iRFwcNE+NAFCqST
GJmBNQID3hVrdb/9Ro+fl9anHwDI64UGgHg0+wH/Qp5ROb89SHaIVjAZejqyPIJ8vzyIqMJ6bzwA
/7AxQNlz7sfIDDw4DplIUZVwl1jP30XYt8wqmInn9vOAsJoU5rZWLKYX2NBZyCz2+uG3968TMk6X
P47vbbGIyPpfV7NHbkFJk4eZkwks/tqdfXtd+u59sciO19Sn26rCE2B9mLhkWk63Rbe2lX0lfUTF
l2YMPT0eAnV+4SsDa9YUp0lD5bwNgq4TPKDXaOzsuqLjPR8yQN9xthbe+dLMmNlehKNMc/CpXqtW
zcPL0wrQO4RiJQfXurLOm0W2MbmXfLX6HMVDSY/+IAFs7Avvj3lb2pD++aAytlLq+klE3sqGEfHL
0imUWFv5IBjVPudyhCUCJn6j3YpmRE5tsO5hLTJlUCeopxGvohrC+AtKFKEIDJ3gQq23kkqDfkKG
TQkwNzQrIyv6VBdmIm+XPP3bcPbD7l/5OePyLQsvqs1yOcmLsm9FfkvLYlgc6+pFwjq0J8IdxcOq
YqftmQjmEk46sz5ag7cKzcLwscV3+u/xVcbHxV4VeVy6cv0C0DKWcsqM+vkZNfE8Ib22PULCWDOy
qvPvZtBV9nPTgoxIqA1HP3KEn0WulbGIj059uQkLPhw+LlMmDA29ADmSiCmmJYofkekxcZ7Qx4Y1
2t8z4aVwmZD5yF/Le+HYnwotBs+Kb2AK4cOSNg49Ob94gb4+cMTPV17mck9FE+toKODSjbEEFHz0
Zf0C29yPU6US3oamuOqKg3Dm0y9ibGBwVOXTUs1VQJWabgeNgaXFi2m7MRnotk1ZGGstIO8UmU9w
/bY0Z0rQtz0JLS98ppMYnBX+UMCrDSLhps/eyxxq8+whcBVPj8ysIY15LnvQeg4NKg1de3Gq9Ski
CwUREqjGjoFk37JbNwHLjMXqUycefD6diARVpuTTkVVOqlrB/qLuXXYpN4etaaYuushwHyOB4rsw
eLTjpjKerITGMz4upVg68wTA1dvgfGsxEzW1vfN2L1F1c5Vn+zO0I2cpV1xkcr15/nH1iZu1bVm/
dA7OwsFkcQeYuAS81o7kOulGt1pnFd8AMRzLctkDi1PuJ9Bsv2/yGaOBU0Tw9HiVr6YyLhZHAy/3
okxjtzA/cSLPL4OIYOUTbVtCqfXYZWznSZhEqvz9AmUQ5tUheFhaChFCfqq0qiq9NBwZj5bz8mVE
/ncvGEC3Zf1LipeDJmETkENIb3//90lZgog0jPnsN7Twa0L37E0LcnbqfgkVeRVMOGXPOUlsKQLM
KwYDzLlNy32qLkcoQsS9FF3jlrUnHHpRLaw/+jVZpMtE1JxykNtRHItLJkeubEKzUs39vxKGmUAe
GjFwtLg2a6OhjTV5RvpBIiNgvkWDt/X5z/Au0IgflJPtHwayOHNxEkQJlEknQ0fnJlx3ixWli0xy
8INkg02muWbeMPtW8VUs4/5GjzakWtajfkr6ITvirAsnZ4gtgJkMrt70QQMhreYUQTGBmYl4Z1/w
wSlv/SzA1gVf+MXA4z6HhhWHp/V+3/5MHtEuWvgvUutjmmaNkDWPRSch+vjLW5b3ZJtlJV9jSQli
ITZFX6Z3QNyD4ewzQUTdkCtjm12NlYT9nDUZG9BEleZXFfkKLrc3B8ekrWvD/5eOEES1mKhY6P6O
dMG7qXKIRspOYxFtyeslG6R9KUTM7+3TiZwxKYu2993iW9PGY8Ks4dtHy1qYDlivixNbuIyM2yO4
+hjUZF4UrLBdV8gXCb4Co9Qn5JO+ki0X/npzyR8pHp7suGS+Rl/H+Ylcz1FBaHjb/XUyuAXifVx8
zMBu0rG/tPhj5us8DQrZhmTwnbIChqZwthswb/3vs5yNTHwCmzGImsz/9J8Eq54k3buspFxfgzoZ
xZ/9iKeptAHS7gdkZ35RAC3XuGlSF2gSKIvlyGtdJStcKJNuMV5pi8QdgQ+UE53PfIz9dc4Nj6qJ
y5If4VxhwHnw4xr8eiP/7QTOM/ELGRXd0yCNaenlRDaIKdOLBvRr7I34hHqBpHNkLCuDBP0G8LX/
tIB3BCSDZO1/z9HiIwwRUjyqRnmijUayGC2/Od5p7ty+1h0gxkjIxtJWHJO/Vn8OeiiDS1GrGmfV
2YSdjjnesX0nTd3Y2LeZGNsIa0D2EA36TZH99Y/Zu/YC72l0iTQIaDJmwYLesEv0kEUXy8jguFP4
bNuDTFqDPxRzLMgx2Bced+noWwnnnq8V1tjHacKzlgxmfC6QAbNvwG//CQH/b68MzpSfiFfZ4dn2
iA34HbpIHvBDRw67gz8CUHxBHx7Y1ZvV2Lh3Ta26KrMuSfHaY99VNjU5eLA3dNmBYwzod1BKTOYN
50siZBVG2za6SYYgrDSo0vfN0KsyH5yiah5ALDzz1yqYDA8ZIvRvP+f/awpVkO0lmStVaVDp6/dy
/BXjaqQDMoNsUpnz4SOYV59ZH8SBP8W3KwkMmiU18VukhGmdr9hQyNa+OTOIKFoKDzqIPjOkDSrd
AsOekJcnGd5f8FUZIVl2FmYJLI3JOTH7T0RFKlohUlLs0eaLvu3RiygyOzvznfmwtTjVt70WHWfD
piGy1ftPObXuI5fip3JdUSZKF3J8VAFB97jcwf56O01TSjZXTf2NVrOJiHOv9HDXMWRVc1asA54b
U5krpUM4XtLxoRUutCfCx4L1iFuDjjbFxJfb9P2oqYo6GfLBWXQkn0OHKVfc+57pnWc/faYKa4rB
d9cgI+CbBzI5KdO/jOyfLV/PeXkZFOBBbfP/KossZMSRB8mqsKMIeEsuWSShMUX9PwNwwRcDNu1o
Ef33/WvVgdI20Md6uQcl/W553u5m4gacCuo0a8I0kTANTZoj53MWcBMwVM7Nun49ipEK2Vm17eUN
OnED34cXbjFUVu9OlUSyIJCRTqN5CnA15cOLvOrszO6p6K8jhro6Gk3623ge+rS7SHXZYXqQpoEO
uP0DRrs7c1WkHUNLjjgWPtULQ3+VFbyXXTGOwKEw6TzMjzwKOLYgc/9DiEtOYi5R0j8VNhs3+TFA
tGd0BifGoZxlh5eGNNQuK5zzIr1tZ3bZxAUmon5jiQBcNR/RlwqrrAMKr4nHosImSy16UrGEFzJL
2RtW1nRUmcoPkwG4iKpdscWgsO5Dg0E3blZ718D0MDFdx8icU+WUrZ33AnyqP0W0kC4ynGVWGnCZ
wborPp2iJlclgvnIxbBg4ecVtOjQtSC0RR9Kwi9N97teqXaaIlJej7NpDK8F1pBs+5vPgLK65Fpl
gyAKV7tjQu8d2mxq+IN/W2V/u8HxyIFboLPnl9hE8nyTiefm8b7fUq2rqG2MELDyF2fOKJCPT1IY
CUqHZLvRWLcl0C9Bv5/3uVvCIUqcgI/ztU3P/a9tBo0aF8DL4jDXGpNYXqYPBrUlYQfbenyCQ78A
342ZBMMP/CckdjrMIu8yC0cMOs8GwyTFtN+iNanHW8XcHKNhr81/RGQwNDyE/KmkvwnzqLI5oR5E
OioDhB9RQRQCJ8StC1v3Cod/qqGAAYGhoc2MoTwMLcDXF8uRi28UgdpajX5v50vJ6AR8GOwj9JKv
b8cP58nuhltmlAMwFKe7vTydwAK7W4iwk9E1s4CZQ1LrB0XUxWpMNpZxekC8t/EOIXN8gZnKBDsK
oTmYiCuqxcPd+CKSzoBwHBpbRAYkvBGb5YUnwJ6mbuQPLlHqV3+e24IooA1uuJgbX9QsP0+hPP6O
hPxeIH3mY1SzyqrkKOyVMdb4laa/rzEGGM5zh/6qWZbGD5xIAxH0YI++O45QzGgFG/j4IPEeYq0W
HwuD5+6VZOsyhXKZTIw+adi9qXpzRiSW8UXzPfbniJbdQjPurxsS6r+foOEF/RJSeJRhnANGam6e
2ewGzvOpZ3QCuozf59evmEFgtlooD7VpFeNhbUvAI4Y4PyEDisw+J3pPG4IQIREDKJQChuv4/OZr
umjCMHnJD9nBVHpLHnjBZ9Ccl7ywyGknacVicQpVAwozkOjN2G6/DLXcmk7c5njw7sY7GqnRVaNR
Uk5Gb8nE0NNrt6ViTVd7CiiKfzYieSPjXUkLWA2a9r9uTKyTNAzAjOavDo7cQPpzLJ/uG8Uwy9NI
tONCnAGl63t4mfkk4Zn6tv7SGYTOdD+PMt6LtVMD2S5lP5zNUQveBjY156+a6HOAh7aTPFbe/cni
Sz8PF1308xweKgwGYCNYAa7H0ju/jPDYQEB0KBSBizioVG+93bp9tRTM084JL+ACPPPu5NUSTxRJ
fHxyK096b8IZYb/Oqg9Na8ac5FmZD6o1aiVSFnnI9Ws3KTcfeUsKeuXMqmDRRdBr14L50EBwIMaR
Vx88qqJCbdtthyFyxC1dpfph/GamvXjpaYewBIANPezqtUR7G3ioMBTuAU/ZGt/MBMVjz3heAAQR
jiWpPKycxXPiDPhbTXuxxJ/SPE5MlbOGlNYzRI8G2pzbLT6GZ7JXtJ543v2B/UVht6oelMQCVYrq
zBtQ+2YkssCDJ599KE6PdKyGXdxbW5Z49lu8N1IYxSZ3jGNODtUpBRYuNgK7PWpa/LlfcndVyUZ7
P2CHO9HgnHFFPbyV0medJF9K0hBY+pGZyGvRkOqcLJnLEO/bqISQkbdbVLv2k2T5BFmKnULkcGjD
36QaAZCp/T7Txa2UGb0QW6xmFUPIsMTQGHyWKxKMNvwB+E2wnERSx6/taP4NtK12NHe7LKSLn0Fa
j5uWSgDEdzDqwUX5UiMIR28ZtG7F8M/5Uyybn0eJ/u4yU5NmW456Dd2wPVIAr5pqaerBmv7bGTpy
RZGvDyFXICJC8rLUdAm0OIXCEIWrmfFbTYWVviubQ7oO5lt8pAmorWXRNaMEBnVw5QZwwLkb9Ccc
ZOwqllnDTddvkpNa2JRiiXWAO/B9SzsCPiqJo5OSXKcEBujX/J3YuXTZDk+02hJE1ozo4wCFRgmF
83XKTuvhGQW/NbcbEKE4qPV284ndNU9aB4jtdIwZkF7UnkJpp90mHUItgLQz2Poki+S/X0FP2+QN
4LcLR4tEbdYFtC6eCKmyvmfP4xlNCXisON7EBIW5Rh+Ku8TJMn2RmFxwcR7MonmovsQtzT7Gw9za
IKkcxoWwDA5gSUbQ/G2bgfiPnJYbFscldW0y285UcKpHlLszi50B8BisgfNspv5oY1ktJB+PS3Pu
U90R0hK5xHBsCFbborPgWL9Hp3fCpFSsPrmQi/tD4UngGF14DmW7F/YuAyvTTjHZUBF2OviEPTlz
DsoevxzAemtNUMP72CqkfDtOJIVt9OijUEBPP/lHhYWizmMfX4CMMSNC+rBjtApFG7D/YjwfGUIy
lTcrFyZn6jzrqs5ane0GOXTHp80axfyK9AqlhzRIOjuy7Ekwm8pNQTMelh35nINsVnnyCFPokeGA
5LFyn7KMaKfYsQmdhFM0aH5wR+ijxDaPPIJmfVfaccWvEvYxJL+UtXvSa3tg5K6TO+Y4XiFiWA7H
f/nyIwdxK7mRiEeXQT0giHhugje6A9zUIol3Tip+p7LtFkI/N6tGoq0kWIsUFBBtZSsbOAPtF6S7
CR1vlh2Mub+IY6O5HmFwpBg1G6iwWUvusEqCubiDbS8M3vHaoTlWsIw5pRr1t6cjKejgJTCrropI
x5R0fMYnrMoLx8lT0AdysFpnOyIdV3BRoqpCi9BFFcxfBklv5lKTmPB1HD/JaCwZUEM+dUceLNRY
vvTqbPeS2L8cAMbLo/Gj8Y8iwnVonWdTJX3bhM2CPr+a0WvpklHrjzdOCFJPPpSfOCgrn5TsQTlr
beGpTdneF7MeS+DUuaE+r1MkQ/3R4FeEZGveUg0FHFuGyEDmg9tAtWYfoQTZfoG6mc0sVVJXV8Wi
q/vpUmzfP/+sHW9ZU8Dm1EQJSONWSVuhUkWVPUg5vsQ05T/J3ii0AXNUA26dxCF2ET1LLua76MGS
d4Vag4AjQzMHG6y0YxHBwvQU3rrVMYMDA9O21TVyKOD4IHj97Gw8Y8WFu7lA5IKQ/Jom//cvErS6
vTnqacCDnwqyOu9Rktromn1rBycg/EIe4pZ+ENyARI9E7zrGJcjnr4RQ4mhpU9mxbeBxgtPZqnIb
lWzCWFVfuLYm+5itqy+xRI+THkIeETw0QAV3yaAL9SCRZckzebXQecE1bblxYY60NiyCYTw6AMWO
cIdJnIA890DLkbCXOj5pMHRxL6hWMS2K5yF3KcdaAHWLm6kQB3Af1oaWAk2sjL9oCppMR+0aOO0K
go+HPDFNdOZ6BK6Hks60bHP2rOMD2qmJVF9sIKGRuz8Wqz/npHMprm/6sK81Mi+8d49NWhDBfzt9
3pXHuKJGEOVa8NwhSEGu8G38+hdlPgy/Bd3xp8nm1GFR0+vAmZl0H+9s+1DBSt4nWLPgtpy3JoGC
7sOavyZSf8ch1+AurYL5z4wZxbbYxvYTN8WDSrCfxAINs4vW8vO2hib7zzTnxHx8seDla4XY8cIj
f5mUzXd4d1aV7M74rd9tscPeF2d7veMYBAmDsfFpzOTKS8/bCrmdcaRNaIuKwgjAi7W2it4Uuiz6
GCrEFfYiI4ViKaYUCzhfjBkKwb9hRlYODrv46gv3ZE6aUA1oNyWelccb3KllemfFfG2citOYUJ53
Z094h33sWDgkBG5mkuDYU3yIQAmkvS0XtHQ32/9bjnlxJER58h8ceSxu9yOiX8BLsW6UOpOovnMJ
NTUVXCYvMXYrLAHT5R8WiFGiNeH/buzusqpsfNCuA9RxFx+/daXptfrSTmmG31Ie8GCQYyR5F0Kd
7js7tjDQlZk4zwTLglqehTY5YEqo/DODpu9/Va9DHzXIbClWWWpM1AnvF/ZThE6L6OLw0QNa5X+I
OeO2WfXf9jdePF9UvcaGsE5NT67P3FS2UTr3FROEhtug5MfMvAwia/LOKXDBtbjJcOQnRVjhd1YQ
urXEVeSMbQ+qymENkYnt3RUgNgLivQ60XMaRD0m8HzcsPt/vWeVeP+Li3LSzw0jUqd6vIGeVZcZP
YoLA/oKhfgt5Hcq8AUca72cMa+aEMOiNjOqp44hzN+IYZK8+LrQgZvL7QjDMyD8f9R2Wa8NHeITr
t9J3DMUQmz8oq1HMJsI4V0vESVz/+figJec82q6zmrQSVR1kh7vGbFLxXBGgUp4frtQSe7FzI1mZ
nrh/NIaySUz2kLLFA+y4fgH7qZgZWkx8ttJoH9LtIMqgWBoOclbhM6fmMWUi1wM0fwtOvr09zPsa
lPBdM5wdule0kFgrOB+IpHezXzLlo6gLsuUv2CJGeRN3+ij3IMXvI6SsORbEjKsqL0SBo3LQgiJL
Fsq9Rc5zyu0gtMuUuv85jDpjr+pbAhORcZvDAAXRGT1EohlXoaje4yyJB3rgI8XQoVzS/kTwLwNX
UD5sGQeDRIdQuTemIJQQB2Jqjv7HttlOdg8vaYB/fqy2sIU0GJnzsP3jVQiOjum69giPkoBhpgLf
HEm6H7Za/rIeawFIaF9v6oIkcNicQ+CQ2yp4nMHVKW4D2xzYv0EsBHD91sh1LNkxDFX91cF9jhIB
rJySANFkVkmFu93BZY9sz9lVXqRYKgQlhjG//3QpBQLQ0Y7OVANuGHtitxg3cABMQ2ncJhuwrbYa
qS0aVPgba++AGM8MTPBQ4ry53o9BxP2PRxj6GbxOA3n7miU75+y1Kw4uIDJKvDxnauCB/ZG4+dPP
u1stGGEu1N/hNtWoUDuV/4ycY9V/RAHTwUiSm/8MVuLWnHPvIHqSaSOln81gI0Tp5LAmzpsxU+ye
VdDKke2dXyeesTsKz6LaNIgCQRqI2hKNpLMf0mbgl3r7fNqcEbk+qZJE7TGj5UqnfY2a1yc9wcfF
vASKRvx9SyqldtRSLBqKI/pZGmmz4ldz/nj7GkpFy4bvjoqe9Ufy6/HeP8Z2FVzXfLGT4gHUkZf6
+HR+DJgUxuvK3bGiqv4hkNIPn+cGm/Iycd2iFRIFPNKm+bR8c2bqcRlkB8mCqolaaCXz9As6W5B5
yvtS1dSxck1ILbbCtXwCSnXPSNQeybC/SOKHTj+RFgwEpqjsXHcL5CZ7jFVASIzJrH0VW9i8aG3I
Cc8TBHeBfs+Ik/cxPiMBkxavseLC4ovsiFyRdSzeKkNw2iuISBLojAHV25EIqgtLjVF4xP2iVJUb
V2lpMkTec2y4iXoS2nHiXNF7bOk9T/ZbFeJj42zFSL2hnWXiUXqrwuixqick8Kve/dMkepgW3ZmQ
ZPFsh8HuxVx4w7c1ETslkI/IKBko+hDb6k4vmPWX3Zypu7Qwc10S431mTt9ftCRn0JWTyEYmuWMq
2IHKBzmZOoPrq3JfrIX8C1/De+fLub8FFCPVwK3YZSkPW9miZ89hWK9IiBbyiNQmNUzfnIofU440
zHVuavWMS6xyZfb1lYX8/j4EqDmnnGtf2YJLV3eWL+riEg6zuTX8BGAzac8jrlTfo/+U2rIZCA7S
ifj8A/lwwPut7VOTlmeCLnxBbShKcsIyWzeKSjAqHYRRyO+fozq52Cdsst7SF1MSTPl3gDvwyEcC
ATTIQRoKBt97dh3RDy8F+OdOA6vmZwqiHxc1PFvkmsaQxYe5k/2nIkcaJvDnPHr+rdsdtfO4QXI/
x0b1d+p/8lL21kO6FjlIvFz993W7eVA8jWwC5HudL1N0AsH4kf2qalkdzgyc8YLk3udAW7+soTVO
oxDClv1gC6UVAxHn8BfHun488/DrxzK3JdHoxKAfssSy5PfX09Jby6RZlA6tLLg4psBTCWoeeMGv
dI3cKXHArvfuuEzO9AGMrSQmpFGtlJ3oD9T7y8Ttm7bOS7ud52WOtvb/kJS2yhv/riv0LL+sIY+i
nU58+Oqd04H9nG52shiXNkEoAha8tLTMhkGF+8GGMg9GsKKQ6s+hU43gByFh4Qpmrj51+1SZuGtJ
YRQVl63xi5sFjeQF48JrUENgTz6fqesVngcuh7m0pYCYn3ebdl/pNDb7nYf+dE0ksZ1zq28gXt7l
fQLW+lKDGZF6tufMPD4Eq0GVXgNMAMMjeiWGcNLlROiIBec+o9IEfKOwooUqxCF7fYXFnisjjf45
p/L3YvIEvprM7aHtBheJ0Kq1uxYCw4LbQgHqEuWZgl3ybqI2/nkfp+ONhcoMp+k5nITmO8ZeaVXB
76yUrsw6s/caAtX4PM5FIMLZQu4I+/DT2GixF90jkSSJKbpAZbfW+PgkDnr2dkUaGnocnz/3VE1z
cF1UX1jj+7kU+f6aXJDZlyhhHRN3L44/m+jvsJPqHFAsLRjE3xUSctB7GedAFWCr2iN3aV452O83
asZLPZhicTYcvZHB6bikFMDivXaUlcaRXTeaZdioZj3k+b+tm46sCjcXl/NfRRPgZKXUhW5+0CBq
HWqqu7azV7mnFYUrKB7qyLUZ3BAg1a8na55v+EOQ9RVGiYXSwZNKwJFoBLzrcw/SHG69okheBzGj
7sa1N7I+zUpP706/+QRzAZeqZyHRd9LDi6uz5M7l1UiNlrZg9DgWr1Z0s9u9Mm5yI31HXLIb1XvV
4GEIRfjaDlVFtqMUR8BPNTppat0M/d88UiXK4EF0F/SwOBQGxRwxtSkgBhlDUXC+QBS8JaW7cFhD
7j5XrUs6YA09goZnJfD3B21Zqca9ek7Jh8xmG74zAE/Y7QT/zozUlnDQhE+G/Tzk95pmeiFob67d
2bARjpbzxTfISW0krlZ2Ac+CNdRnuGmmyXUBvghQcXlNGlbTREvZwn8K3j96kQcoH2BJrlFeQwip
u4dcE0FdmFAc1oVv1RF+5oTS6uaQsEhvuSJtPdGgN8KIi4Ijv23XFKCqrpOjUUYbNSXtlp8rYOzH
e/1ta/YwTK4txjeLI97joooQGhSzr+bkEjEaSXWAi7fxAXk1lI3YIvWCuoKogjW+FcgDlrkL9vHL
1rkxNFTAPf5dN2NTAVcSJFdc81VLwZF3h8VR8JY/H7oeBnyQXU0VvLa8f38bVUAczpaMS+BBPdGp
dZBFb0FLvnb5hRC37XF9Lns/hyBWciY/4amalA25vjzwS3A3synxm7YmuN1wLOFhAUEBSKGzS2xN
88cls9A4qCg6axRXzmnwKzbF0jFpZjYsVpdoeOIbgG8lmDg/U3imWYnMjEbRTsUeqzZYCakBbkP3
3vWQYhWsLUhSbBIrdazpYzgqdC9CxaB4x61Z06vJkXfua0Vq2vmufbn1jlfQQTEEIfUpQrqBlykd
D9P2IOZtXJU6RU1KbjWcf5kb6caXHvxOHKTOOu7OmfQ7erPuLoWznpKde7yEfPRv862weeELAj8u
8TCQIr1GdGbBy37q+oxLTb0DzfLsBMdR+lLIDU3/626QAFvPfIHzzIx0Ij659NzUXhOvP7GwkvXb
LH/FEPYn1XZ+jzxCZiZgDAYSx+CVm+t5D+4HhMZTVQmANN2Jjr3tL4H1cq6lSi5ki/bNUO802Fv3
P+Ccam4ukohsJ0uo6GE307tDWge6JZbC8l4BfsQZY3FIxSqUaeNXlLQ+ERTKR9H9UWi06MlitmgZ
3QN1PpsXFat2Y4RRV7ekPkyb0R87ejpepIU3ng1nFTQt8jvg7upj3CVdsGf0FokO3tI5UR6LyEfD
Kno0EQ0JFpByM+X89SNmQIm6tRpefrgm0hlA8YXy5ZCyy7SQ4j0yw/cO5fuLtetSAsniq7cZTsbX
/ACAEFirLfPx6RL31CvH9VfFGFHjW7YYqezCCK2TSiTB2t00bXOveolxjYbWgTFtQ/Norv52JQVq
u9WSRIfHJCD8MPXngSh77DHio1AF++QB1ACGJq7AOyUspDCfOrHgvmt9m5c9nIVA+TEaJDZOFJlp
q9btcf/6yGqyFLEbAUT9v7uqrSsaQtoJMoLBl2ezIiJCTmXGv5fphui33K78nVpvfiHvNPWSS0cz
n3XypmxcyaJ5uptZiQZ49dhuiyopSJsjWVJAmetrk2+RR2NJovNyC0hx8Pz2zRjLVC/XNYp5ER3j
1KJjCKr9BpI+MJYb7laGhpmqRkJd3Ej/UHyXwl+DMZs9krDW0e7dq30283cvlUxxTuNNEKq2Ovg7
5mjHm1edaS2u+2X9qmJXfbqMaDK1h4TmZ8wYHc55OTSz91kl+Cf1Qdw2ZUTJKpQbRlb+fx5MWSVD
DrVSxHqDKsjTxJEkZzHNWo9eabogTvpmbQqzrNPwDYN5w7UFmbkBor9uy+izlMUcPawsWpvPc8Ts
sZXBz3VDnGl6xEZWnvhzQC7IHuI9KI1i7kDU8Z1d/t0sl6L9hVp5wu77U1mGhs0MljE8oQFdH45L
Ikue8djMfZZt6xuNW6gzCwR3UEsljo+Y60UyR8itQHGpy2G0ui7AsWvVd30ehulWYfzFis5K5E4u
ZgJ8+oNbqaYWTYJ1V1dRzmJymqQGkOJy5h/eF9V3T9kk6ISf23aTOoNskrPZbK9TvVA72oHxjtXd
h7TmQYBvzCcUPu4pEyEjrkStdRJd3HP8kN4ViChfJ4wWJ8TSfWkLzkcyWikA2RoBUIOddlDqJnyg
JnFc6qwMXmbj88mn8j0IU+hzNoYzAWXcPoF6PhagmC8Hg0rzQSCVedLkrYYjaeslC1ceDJfKrowI
9tQN+uutCXq0s+Zt5yD/tGR2Y9NSgxd6pitQKBotqgs426bNxBvRHtfFo3DYhyp7gxmOiIEipgMj
FfcGeoRi9UTc9K4VL7VhWdWZoe6dIDG/rzolki0DmfxTESZ3GFZY6eCX94ODmoAcOXIqfB2QvDgJ
ZE3tVcEcKwzfdbnGrVKKlh4Ka7nprNnHGITIH2muvoA8ZG/PfvZhiAvaMvRgHVqrrnJyu7qPhVNW
hk3fiwck1e0X/xwafiPS2o35GQWO7ySmjLqqwpdjBxLD9kMbLXcff1BRnKYPJqUz9NkykXs6DfXZ
7Xbil5L4ocBbTbmhTT53HCLLm3mJ7BcSWhCxdhE7/rlQjL2Q2wMZ7v2e+PKcUaOcB+sdsUyBq8ku
SWg2uaMmQtHhQmJPWGoxyWVpTGGNLJ4X7rLFG+XDDVC90scXhFrFHgRelGRE2MS9yUe6pHkXLq2x
2D3td7ynStolZeVfis8DJDDHBA/FpzzXZyzUeyH1N7Jov9yRMmLERoL+dQ1i7oa8LCg1ACGUl/PW
s9V0nMtiwk6P97KPJpa3gKgbNyGlF2QGGpEzLARinhAbma/fIy6MJvqqjeOa1F1GDuoVMN5rL1z3
4YVzIpH2EWLoLZ/yEB1C1UH1MHrckKzHrtBZHlxQPbtfMllY0yUOXQNIsdZmWiVU5SBTe5Atp48/
YCZj1gRNoG+H2Y/Jd/8n4j2vHyedxf2NdevhhLO7mmt/stvj795G4LWO20blBhX2yMjA8X2ZuAYb
0gRUO41883g8OOhh7xEooKy6Sb1iF1+it29Q+0GmWZk5OpUZMm79DpodN6yrXYAxM88jvqAW+1ti
p9UMVUTV8mv5jsXx72GETWWc2W67keMXGkMY5U71VvU5sgxbjXmIMcvGKZs7czvPvn3rTASGT28p
MHfSILa8+XrGOt5UZnM1ZDzmQ2ohcePm/+tGnqPz5lOa+BuQFANoO7Lp99PP2XIjkN0my7UApDKo
sdD8rwDx7o6H8U88Ndr39UI/aki9jvBLqqfVDP0gLCGngTj0g21AKbojoyfe3DSa2OkcU6ZStUI4
oNNg9LRgMgrX73beOg1oykuyMzU41BgjiW90ejTZThS6rPWAm6vS92IJ/HIRKDrvD10IBPkZ4B77
Sk09OOOvi8/1iuTsHHb0H6kqXCumjdzn1NPR0/C9ImjX0rpEgWShC7DrZHTPfxvDjQNMIL9vh8rC
qgv9Hy5vRsW38DUJ/PN/OJsFPkM0LCWvzQqpgR5yILoymxItg/J1UlO+CZm8xrmTPVBm4Xr7qFWx
Pxkqe6hJ53uJg7bqJz97DcpM6A77rcVubmaSSaLsp2R+eeL6Z6IR556eySTm4PMXS3yKAFsLPphH
iCZr6rLCeNGkawkiYy3pqsJVo0iIP+QHKyXEGWua8iDz0uEpT++zuiTFzTHERw7ZxuYtwdHIqJPJ
EJ09dDQaNkstICopFI5CLzhrGVlJZK1Sdnf1NvBRU5L+4mmBZrov2hU/EAFpwavGFl66Q4S6DPq7
KSseLkOSib0rgAdMHlZEAWEhEeM6HyTNRKQYhzNX+064Gmrz7NVMPAzAovuU/+br5I8eO54Dufl+
Hd/NGz2Y/JsdfJSrORgg3xQ03oEjdQZjKCMt+YKs7WMobilntHwajvmSMmx3aA5iv5GlU0ISdSCt
pVQ81iiN3xr0Pc4npmAN4dgqE2TKg2EWTb14Gu4n2v2wGSpdrPwwK7vyFOgutFVDm7hE+FuOCuX/
bGl223OviHH8NW0g6gUvtK2jifl1LH5iS+LBfWKQo2A9coqna1ZmW6SqGHYj4n3hmOv3KwkuRJ/m
KFE7Rt4ZkjFzOhqdSRvDFG1I69igC6apSJIA4prQYL10fFWCUNKyJl3xIa47iq6oPL66r5NFKaGj
jZeSC7e8Hw5ukNKzrs63UOPDVHlZ0uZMK2S5m/054uhGr5qdL8+ZUdjl1GltOBFOt3YiUifiaCBZ
TmNR8ldAgfTXJraRH4TI3US2kXl4A5sFZY50kC8GoRhkQLI7ZtW5YXczen3OQDdgNS2Lq3yxzEj2
j8Q6/NmpV+zM+rpeT8OU+HCGnPot/buBpPA0A6WOuheA60fpnLqrHdd9SvJln54UiYtZMc3TlmF5
1sk54OPHbwwYZeMEKJoI6mNEGVlSy/0pZDnxam8W4io6p2JAvZYbukPTksXm2Yq/vnLEdOOiNtkc
t2J8t2xpEShKEB2PpC025XiD+13yKewwTKR3p4V3FYBHFkKBgFfwDbgehcaVuUS+QpO3jucfGdpt
jXKStFLLE1A7VlFBerUfaHLkc9B1QkmD3EwZspyLRqdLLSMOcYr4DhqvDe0IBG4WnEY8Ld5G00Vw
o7lnRGDrq5Jp6aZed+U+JyPRCzsKa98Em3Iz9mlOONXo2/fho2JwrKOJtCMDUgvPHThkWgFWXIba
2+7o6VHlLqqlkUzWD6D47fJaoNlgL0qX9VcMt7DFqA81jRrlQT0YK3GZo4bmwqBZdGfQzqOcQru5
iQ7CMXveN+0A8PV+qti7p0RN97HKZpTVcT1VylQILo9E0T2hXnIuR1W3bIdiy0xJ9cjqP49rxEfr
dgMOxbqjlpxUJSosWkQNiVbZUfE6IjW3g91QMmJU5k6oBJFNPmQNXVI6Qm7liZ/Wh2XSeO/dnEkf
bkWjWdx8lz2TYvXiMpIEVIvN3HyZb/lT9bavbJqgksN2xbuZhY5b5cpcFVuzFd3E+YGY+fEgMc76
/WBuO1+wB8lZDle0kHpTCHcFSr3lvOp2Dkf8Kine2hZsKEd3lmfS43OzQOezugF7ZhuNLuQw4dVY
dZnGs9c96FuLBSMVmlO0yeF9qDLTrsb8FTTsKKYQnZmiphwpQMp4Yhla+CoZQZMji9VOEdKP3yYU
y2kTDoSMhrOIiTRx4YIeeN43MCj0ZVa11UTLiBTWpn3I55hJrEOerhXgkBObtpDq/0ehOlHhKfUy
nGgCIKIjnnLivNDxEXCjhainP8PcsAQDOidDz//p/EqvyaKM+XO1cM6zA4S0zjw0h9GPPcUUQKsO
+jnE+wQ2nULvLdWxFZUyhmA/nYjG+7SvqPyEmU26a7YKvIwUJUfe/zVzLtAfvDAASQQWfgfcYVBO
cM7UjMylfwVvPtIkG1GzZ1aCc54ssc4DstSbkdgECxtm4GwfDhsLqE4Ep5plduNRO12MVOJQ4X7o
wrrcz8JFqOhO7Q/cAdqxj6ZSsyZ2/bMPRMrB62hGMcNrzoqW8Sh5YKmZaPcUTWeNFPodL9bd8uKu
B1Y98gJf/3jr+aRzvmWb3Cshd6a9MzLPgorub8y9M/J8oZsXMUAomvl8Z6pQl/XNit0xIGG32th2
ZU+M6mibfGNYFV6xm30EqNt7JniUUOMsB0NR04cEQ2Wpdj5ri2h7B9HdWx1yE/aWlaXrsVQYbsJP
NUiKEtzpCVjnZYIdzbQ/A0az6FdO/pIHxQIpLyWKkbYtrO6EuyloLaTHQCHnEgZlYCvcrJUm5w7P
xjL8X8Fy5pkRivPNrkvh4iv/DUVRf98hde6w7oRtH6K1oD6Fut/JTXsqc/a1jetSZS1Bp5fVRKgm
yNQQBKMJDIYuSoWSkWHd8VsUmPUv6MIx001RTxyUIci4jH0o0/4B2RhvkTZzR4qal6V3OtTIAnqf
quGVVYmXTGQXC0zE2eWjWTB8B6BR5Pba5EvYk4i5syGGau/RyvbudfkxB7mqDYgchRc5M0ZPpybS
C/Hp3CFORi2jWlblcSVIxQhJsdufnVlRv1hS5Qpx8Y+8H2L8cwv0Aplw+B5DWmSlEtTSDhr8PEP/
vyKCPmChsMzhAiH14kNAawvBf5swJyQlmvyouzYLQYKetku4yY1ouc6/CK2QEBGQZ/zVnExvJCsm
xtpsJIU87oRiZDjTve66TVoN2K+bgVMpVpGBBAKJgzhsOZAVOrtMnf7bqcUDflj6WQOwxPIh34Ks
VNdNn6i1gcnNZET0fBU9vK7EpkkryQN12lJDP76Ce+Gl0JnsgR3RNf2GXvWLZ1wsG0XFjxwQysdT
tUNw2pDI+GtLt978ifQsQ9rF8fU5GrqGVPmNqSevnGS04Yj8f8opdjBGuvRuS4eqf8oEH2a1WLBt
tIEwuF+VRgKhnHFMRW3cccMluZGi2B/iFLbY7RtnSFujXM3gllWPgw0jyJd/wcbh1IUWYq2YLp9P
F1aSTRqI323sRBfHYzzMWmSgVEMdolfT32onO7Jdhe25T0nTTiFQQcRXk02eW5hTjqcXEa+wwaJ3
DQXaca/d/cF66LpYny2EYDWd3785U2bP3QD7k7O1ot7jB3bonXGp8/B1hoO4utZ/z66iSEzwypOA
M81ACd9Bla1AD3adgHLOtqCCsLwN6pftZWPQW7U58XIKx3iIbUkmdSz0ZrnBvAB1tkqbLsX/e2sB
LZ/HGd0zd8+S9meoeMY+MfKwz8IUSornjcVtj0+BxOaDRnbYwwx5+5+Gvl+kXNjgXFJSpHg1peLg
nTSX3zqJ7xOzgLdGFHCm97nczFYybECAqrTl9rW9jH3danjk17mA5Vx/9hZblqNIObiYRwKtqzi/
WlC16OV9wbD3EpXHXpwuZz+1hybcFY/TpC/tdFSb/fB5J1WtGCeHPgRNZoI1Zn+QInv+nKzj2p3Q
kCDG+3gIITvrTEIZxd0wqiw40hDcufC/4A0YOd/Goi4yxyc3Hv7uRRMWAv5lloMTnGyowbx82g35
x7Uj0sD7MenwByY/8Q+he6M5l8sPzO15vt9EbTRUtI0m8ENocgU5ovr0p+4UijZpIhJisUn9w4r9
Scu0JQURELEzPlmeqLO7cNlAt1fM3n2gCGdPsEcUWVB9u+sq9eb8NFOGM4gsYyuezloJXmpLLW1t
OJodVpJn0d9/6E1xNysJ504YGwURBX1APn6Nu5F1CGaLyaN07N60ua7QLzYWtolhri82yUd4I8dc
d4/nbfSpnD8yE3Kx7vDA2uAlCZemMIh+2Wlc43wQhZ39IaUotIKZIArwY1IjkPv9N8J8ofglv/ha
PvgBApU9S7VwIraiRxIuaGgR/5f69DzTBBOFXQ26sAEsUL0kZBdOjf32sYsOeNH0dCdf4dQjKbdH
/Qfo79HsAdSpYmYA+8W3VHRg1oN7zqXcAAcUCpsyxlHQaUthKPqPEOiX94Ed2t5ZVwWVG2nAD1mI
OKJQMPEIu6+hn0V7eWSvIS1HpdakGy53XwwwEeb0qM2H8fRSiiQlh39H14rxI8uOosvgYI4vxk75
+7Jr/bXf0nt13NBt3zKEnqcHLzz4yuQHItzNZG7Q2UdhfneT6b7tqQkvw8Gxz3ApsAMFVg3xwNf5
JlZ6M3ZpzyXZhnEYTU11cIZhHQIwcHjDsAwmAoMppkAvw78Bhjm3z1Kkk8oEN/8AcMuk4JWKuKk+
P50RCyUiYmGieNcqW2yVAcQKspr8iIYvt0uRncGvl2r1Rggkk/M0eYMMELnjYFQK0HjZKi99/Gre
jQ4h8ZLPfusuDXaLZUbJRSJFcyAKTVHFUHksKYNSuVpRFzILihobIJG0FehcEJ8c3OpExd3wHbV0
8+XHXnq8g2u2tNqOoSeyVDu1IbW57FIYV3wSIOnjxogtC0nSs7fER/QZer7X8pLR15dFL4j6JVFt
tzSHziiiw6hNVzr6qlRCKYPu0Tzgrq/h+Dp/itku4BnNSknzPccuRAfLfnmpZoZRkLqZ2mX3jzmZ
xqHy+aNyJ4m8YSeoasTsVyaWK9rG425QKNOvB3gC1w/yc9B8tquwKVQvS7jTLqyKX0K7Dpldwnsv
PK/RgfuYOHBSI2QvkFefhbKuJOy604+h+e9PEKB8QJrhEYybVYAu3pu6T4aI/WcQB8W4ifRkuFom
WJVv/uinkq5DZkvljnQ9nL1wGmNPKZM37YO3sYI7aSEQWr4+4ViWW74LnLerJM1rsgVIpcRgdQTA
bdBthxbPdhXHRwm7Sd2T8QGNHsQRtpn57p2bqksn+kJyxGotiGfHto3WY18S4gEiC+1loekVMC7o
Ujqqr3Z3Ckb0buR8hFmuBMpPrW3KWyixmKrzE5F4g7dqd6ej0nFu4quSAX8SWJPy6Mf24BlMFZKG
XAoE8hNQQyTCvf9wIjzMTMl0IiSqw4WV+iObuhOBREtLTCqrCDK3CM0RaPFbB6s3Ei/tmQsv2brA
RUKSKamLlSpFvlCljP65K5dMDGqosAfSvI0vlf3X+MLDrtf5Kb4ZdBP/4r/h35iJLFI4zbPHN63e
51enQlN5gmKpl3SYKKkShbiIaCo1vqmCWjmg6a1PUZ/Xb4GAuYmsbp6MV2cpb7jMBQcGMEJnLUtg
HUOSt0/b4otRvHF0RFvM/bEUXKQumcMMdKnKstEdipf7jbhpXCvKl4a8+lIBM+GrDjvLSvhgdNMO
2+rywQOGpFVT717D60+I5WlPTXwQwDvALIBcrpZ3QjhkzX2vVhQ1AzN/cqWTUrA23keGZsYJy7VE
QH6rlZQAojuegaUqVLdLY5gzV15cJXGPLtsztr83vJxtX0Tb6itcMuF/ybaYxPXfjypbjDE3A6EH
UpNeYTPFBGXu7dBKpj3obV1tGyfDFMctKt0QYyZeiJdeHw7nPaUOv8mA7a5dhAFqS1G8fepNpyfi
yS3U8ZDx6MFmIuqCdxDNUNKrPa0xZdqqrfk0zdK+oKw73wQ9/wS+6SoESlfgGJzAk1pvkQmM5jx4
9/ACRmh9ChM/A+Le/IifKGlfiHkQrBEziaZ61Ew3l1rFo/CG5s55fzaejoHKAVFLhIYsVaynWWnM
8WGQamb/VIZNfQomrGaHAMIbrCm+nsoxWnBGBDKlqFHDYA0wB6d32ymE5gxZh+cJET55QMJ58J+G
Gf+dnfbbt3JakhpgYHKn2xlJuAgcKoEfz4DuucZFABzOuBrswobhO11cy/G09/7n1kEr9TuysIym
vbs+CAg/c4LWODhpFkZkOuQ00dMRv9oW4lDlZtM0vtP8HhnWIC0Oa3M5H1fIEk2UDvGQvcIZFIx7
q/2jbgRayZmMRxtO+xGmhBwpKZKoQbs6HehP73HJ4JYw2/yaEpuD4IrUry+sBKNJMrymX/Kyny0A
/iAnfSY7GQ/II2r+unhPC8fyQQC+98mNM05XO2AsbdFLCtmqHt/3gRjy/A+58BwAw1psIDcgZ5aI
HKKMBywPQqmmYTgCau5kK4IXVn6GMe9CzLb09+TZh8pZ8fFhbi2S1W8uh63BKmeyj1LDXwjVTbq/
183pq0Xz8DdYkEM7M+dOZ/ClxEPbpd7ZuKN4eUPVaZhUom2t69HD4JQ7BQqMuT1Ofws/f+5OxgYV
yxkjK9nGgYpwNm5gQpOMHi0ETLPRKNm9tpZW9fB1l4VoJXYpTmaTJIIikW380/ghjIyUl12o8EJD
z4lNd3X5NUieCw4fH8iSvBkRZp2yqqljAESXIXEOFoScr6G1fHiQ4rnVmsawTmbKRd7FTsEsi9JN
OaCzWxi6fNed42gxEwpf9+BvNPw1ZOTzdFWXhMrHJM/2dTprAKAyreY05TseEBPjHGibjqei1Is+
CTmX0N7aUktCyOpsfOZI1z8qkR+cGwSzBE/aD8XOgzNOQQX6+fFAfqPgS1ibqKWr3alVzPksz32t
1tvifNitMRKjoTel3uHgInyePA3VyobAFiw0Eh8mSmwwfcZMM6sdswExiP4UdLJrI8qKIFwnFGGi
zE+A96XpGwvwB6MYC45YSB4qx8KYhWpyvX1qddl+4qCY0N7xByyb0Mr+8GFReS+Y2yumHLirO2gV
TWK+/cm9sI3odDp7UI1OYGA+kAsW7oYuxkcv8xx040xMeodkF0l7rqFf7auOvKWw6xZpYtMiwUxZ
iIWrbQ1sMVazIDKnENTQF8SwKns4hGghrLOndzxzxaJHViczUWkRKP4nrndJ/quRHvW/DMpyxmnx
5/NsCGPbS7aETkT6GWMhwlieCO6VYMjKerUOL5WP/LPpQS03QUu5494btPp9NE5BS6AJvVVIjqdo
FtTv0sdvULbrXNZuIXbW6zAZSTOcLB71DjWlQ6cJDGqDXYVX0K6yh0B4ZAfV3/h4Ap/DU1DD6bmP
JUohFLC7tR3yFMSS4YGcp2tMZ+4Ay5tFDBjqESYpiXkT3N9EUAZmGNVM2jdrB6e3SFtrUIYijmqG
bhfL1sOhg1w3wc59VY/h5CehcQKUhwR4kZMRWwdYGKtWJsijacBAkSz3BBDggC79AAgv3kjLVrDk
I952BryCIAdiJR430nzLjV/NTzvc+kVpf8/PzgyyaxXOHgziir/1+tzCcdfi5a9L9IbS7RQV0VSY
JZ80PpF5YCc/PyJ2xmF9/7iD4p7GQYL0rWyV8RBGU+lnG8pB4uAkV23iCjRU8YPGp9iYnAYEBd3c
qsXv3jUAAT5i7O5JItipLafiWEY0SsZRcVDrYfhN5f9SrxUq8qBrrOvPKBABDQ/18x+E2EB4yPb0
SFNjUTLqTW/7SKGEOHQd5/J8KoyhnQ7MVMzCWE37OuKBsiYTiQveW1xfQM1DVGLpWP0fi0I03UL0
uljL7pvdLFVMF1RP5zhnyO/JDyidjxa8ZTqbU9Vw/ldjBvzx+E7oyufEBPMeUNue/5OMvocHPoFX
HQyQNus0dAHQT443N8wcw+TYiphsDbuT/7d9iaPHQC68Fl+20+KTQTgJ9WZfYlDs2hRN/+QuxGDI
CyT2w77a7h/ivQUbVgHbWY/W7aMZoi49a6V9i9WkUXQbPZijshesszjiqpa9klpB4rSLwR5I48JL
53/3o4ollO55ahtk1f7cE1PNRT52YbD499hsq9ef58SJ3XztSAjn3Vp3RCy+MWuacm9vqlkupWoQ
nk1nZkQTTljK0I4aEMKJSHb/i/5ILIponxxJQp061QEcCPGAfwYx4csaH5BOp35pFuuJfFPTNhzn
qj3H75YaJ5UUHb62dsdPPY8YfYgFQg8dYtGPu0+y6qmMxjwG2qBq+rY1vTxjYiwN0ONYvO0vv2MM
unwzWy2kb3BfyaqJKWEXtOHI10rwhQAGLaSeBvkUSs9gsMSY/XfAIo0/pYvlP1D3WMhyw/uYvRMi
etzRQ1J4Qxp0ZxkCDhBjTE8hz3cBGJhdKrjy4Bi7kDl38IJ1xkEdjVB9USbDu9pAdShOAd/udPGp
8LLIF7da5GJ6zexYqcQ/e5n7wA7yQ44S2HZC+MKcHJT9b6XJ6+mBfswKu3k+OHetWgw4mXGvqYxG
ngMNypwd1Myc95/v0Xz6ZkCqN1auV7j9xbW7paizjaJNdGepEBhFpCwJRYdOE3ep9Rk8mrs1Eivr
r9BaVgQW5EisE3StrSwd/AXlKltmAvySci9E2A89erqAlq6DUxp4I8/fZUi4EO3mVj/0LV6UHuvQ
278HqpNqObkucmV2WRdpZDNr2X2BMYc4hul7vvsKBJNEOoRnwgZuDakpCKPk52qhHNBK7HX5jELm
rHvCNru+EPrvY+Bkig16OqNTkM9YdyU7q62AstgN+ZauDwIpcAJonEWp4IhHGhzmaIBUNC4PJ1SB
x1DrAe95jDuK62nR8PAdAJGuJu5kbMk6ztmGPSdMqyhyEFO8ALgUddkF2bMP0Z9hNle5HrW3qtOH
yBlpv+bZCku6TRRFhtZUMGG7Fr6aOufpzwHesybPTfJ3p53RSo2UxbqtqUD0cAVXOxNRkAjmrBvY
1+UOIor0Pq97Jazj3V5un4DF2+mqhRT80xBzvO1GqJCNowYelP6aJdMqgigw/HA/IXUlmH6wVvUd
V2P20Ja/FbQolmoFrBKLgIaOuoUcSt8En8L3k4hkJbvIKvoTYpbNfukeEPQpanQwS5DkCjaY2pKF
bokc/NvF1MfaPk+HqaivAYPmf4RgXWzTlfVk0j8Y1SI3BOMLTcb91M/023fWe3FM5gy2vcEseppt
e0AA9d97toty+9ALs/RwyoVD/2WAC/ZdUORVWw+mZfk6sHvpYKXet//5el7AO1NEhzHTQ3i+v9DN
JIAG/gcYUgkNdFO2EJO6LgbwsMukYn5dWKq/2aFaIn9uSU2m3Ild2CJcHRBOavuny8DSWtNmT7r6
wVaSJZ4ZTqUEp8aZCOE5OAUUum8/BEabTi8USOYqryAh0xR2FNEEAQGjZ2zsz1FTfe/vaaIDpTJx
XByheCV1EvkALfLqw3IRz0WFE4Rg994G8qDR5b3GbdicTVYEaXQbq/M72qGeigLcCogH42hbi2u3
p9AKZzqpHdMxGlJqPoI36wkmnA924PJyVXDX20yXSTbSH6eC7jWPlaBVP4AeUSzPgzZMeCeOAp9s
RaR58M0Jcga7w0Po2M5FiGNZ1tYNLKV/ppvhanlkT0YcvId6N9ywWXZtWzb+3tTqLznJI97djoNw
8l/P1h/RfelRmFhfd2YQqoht5V2nHH14G74anvibQ7Oksxea/uOt4gHQt6JQcIlc7NwL1yZPmrwj
+WN/1keKm883l/j7Hs4x/ZjcWr/4PZ5Gm96fxINCjw7I8dwG6EDA41UG8tshfYwMTMke409k5D+l
rKAPcLBed5AOnwzTU+Ac0ZqQMxDQvNvrdBHORglWxuknvkJL1BfLLuSGwdV771rJ+HD9z7FqLMr8
TYX/H7zrpiE9ygP1olM9MGZVSqQ9oFVyTQYdS60N2Easz9diNQQzgn+WEvw3DPcxF0ynQ46J9Jgs
zKVBQj8GfHvWO+InTM/dSa3gB3ZFe1BRMDV6CiiNcQa9m12LJlYzBWyk9UiUbbI4BNGWLUbPUe0J
2V3GBINYdZMUtD+lEE5tPSEgLFBpvkOsU5U817YToR564ze0FHoWYlaLC1pnfTRnnHXQXPHMjdpv
HeR7DIeGOAq2YzZrpTeFuindDJ4R9v7dZEiC+6vi4YZCxf3300zKbxb3RIF3fK1WQLIVqNWxLjBa
mVQUCFXXYpYlbW77e5N8kAk5mQNoIyMlQF6b1r13yMNHEHbijXXiSI2Al1zLdlpwItcg0j41gyxi
eX8yCXNmsB723sayafYFbV/yiogO36T+qteZBy0d1JLI+/SV+g3xUBg3nC1vyzUxhY2IpEs6+JZf
ZtK+GeEgHWRO8FVhzAcj1T6VtGQIk8N82pJAOdhfJGH4/9KqVPpcHIP27m3F89vVEp8GMbBrAmAg
zKh34IMgR7fe1hgkV39b/lvC5cb4j5xZpFlZoO0iqRDp5r8gyLPRZEJ/UO9CnLCMHzzxYejzxnOv
IZRkFcBJbh/inPfePw3IosgUoOw100GA+QF0KpyuUu1GZ6BbRYnsY7S365qmhzAMjOtEVO6evT6m
2r4nWV9AxoLoZsV36S3MrTFXr+J0fwEJFPJNkRi2SgOWWoXYq+d9pfr00bzpEO0Cr/BwnhGj3sv9
3y5ZttufKvH1WfuQraezJ+66sq37SHu6Ko0D9gOTBGv7zTrD6bm+rwYF5YxjprvIGhQ3eLVvv5bb
whArcn6AFR6X45y3tw+VsNk4Ds1DGl8jSWmIVH/Ob02HRwxyoIFUKZJt+JHdC0pA026t3sgye0ez
QPNTjE11y2L8qes18D8YU+2A0TmDZ95p6brV6z99cW8MdIsMT1/7lQznbYKr/6LOL96jaT2qgQtX
JaXkgtn4nmIgMJ/gvgBrNZ6qnnIyu88tJ7rcvd7AFf//nDvC4Y++cyzmTFADYj3o6xd6ybPskFjH
W0gbhWKq6qQstXcffiHlYUpjxWbRjYIvx8+H0saFTJEyzyKWqsh1YgsEX/jBRX0vwBToo+mYxjQ/
fQbGImTUiac2F93j9L2WLV4ikO6lrSw3BJOAKfgbRLDdzeGSkJJz6JvZL8b21Hw4yBdFeWl9DkCK
DcheBUJW14e3M2mTwGzCCYd94f2KdlA6MqhqjCz/CcmaAo5DwfWjSIMjZUU8szj6NI1iRwHKIpKs
1EmyFATVWPsbuZceXAc7efDqoNAbmd1gSlveaNkvP6fKeQ4XCkcv2tt+mQzEnbDKiDxoJ9oHFAHs
mCvSHUcQJ5hs0VlSf3A9wRI/zTk5P9TKXc42/sFFXZTdm+BW+XmjamX8FFyAztkg//eXtqr6F9xl
FE3228vUzb7yOzW8tBawVfv01la5EHWHYPSOlf57Gj6pPa3vRg4GlZhtiuOnay5juJ8WUI1t5moi
YTecEGbzbFeTyuuzAZWe0GFjJDFpbDUhu8i+oX45ApQs5wsm2pdv0uib7PAb3pSA6fIRaxcrm8nE
YPR0EjxDLyyUid/rL7qkELju+5l1R/4QJ7kJrvtTfLdFunYLIyUOpx/0f5whxEc/pZerlGPoOiDL
nSNLY+fEkFOMnqLaoOJ5GtxfrITcI7hz8FU/S5KaYlrrACYEhs/Y/TDP/7eyQHFEOkW+bOVZhBbB
qjkcp6DLEQ7n2TWIKppcIO2emHab+dSG75rCqNv4LNWshzZP0MN+p/SVOqcQ2ojsyXoUW6lTPzmY
HZC7Re0KeFv2jPn27ZFp0QAxeslcr9w3aG1hQA2aRpnE2w7tB374Xawe0HkqTnlGzPk7LPjLrEf2
aDm+9r/7qM3I30XTmsc3EYQkX22KUVHJFV1xDj5//dsCCNoIEeZQFpHaVQr6/iRUdgrZCiSP4Y8F
kchuxzoptk/r4okFtfbdQvK1cn24EdWaJlAglWKMRzCg0HcLJHq/QpCf+zH8g2HzXNCG2v0fT7M9
TIEuEqiYT0j0AtpTgUjCFkt3fxKXj6vBaIjrnW4ln0AvgwjgmutT7Dp/dj0Hepd9UTuUKk5aHJ0y
508T6ZWU80GDxbs8bwFTLolz3cvdO7d/L0iGYwUYxNfxxcJCRFcDCByfE4Bh/FYCZJ4YwF7tWhXl
rIauxLyDBsB0jSiq0Z52BlCfVBPUqTSe5p6zCbUgICRQfCH6Wm1ITOmJxSY4WPb83RMvZ7QXXp2B
5759wvOxmGJ/quC3H0oeg5FWukTyWU4Sgs1eD2izGeObiyzo9A3yBt8BwcPktCD9ZoMigjW1CXZ+
rm1QKHIS3OZq4/7RRPG+QaC0Xtb/l7htj+fiEaF6+5ppY+Kwi+QTxbt/sG+lHC0wo9FllnCogXdn
02RRwV3XPsOpkeMA7s3byhJpvc3wlBFwF6X4ENj4FwF9axDRu7VZvpySy95E5XeIToD8TvJf8k9y
navLacrF9U8pXZB4CSVeK3e9CjOUgegigQ2XerXDroYIF/m3fD77kFUOy3grv1tPrVFI/EmAHR1L
ctU2o3VhL+Yfg2RmAQs9YGGptkvUawgqh2mNG7f22RBP9+B280oVwe+GhzQHd9mRuLcqZ1O5/vfV
4O2uzJvZ06TjiMwyVyFSITQCPyud+hw29tYkW1tbdZwSxn4Zs4xJ0nCBLzRQ8EZ26MJhzX8vPQHR
f2huT6Pm/3C+Y/fGp0T7I0So1qOrrGA4ML12l7gW9XVurHUMGIk8a0ThR3PHQiJv0GTuSngGDqee
2GCWjy4ZB3kt8UiiIhZACC2GObdqAFfe98JUUthicwRM6g1TEg5XR5I108NiMLQUq8IGsdtDVczF
N6OiQhr7UzEoTd3IU0oZlDbMvFOGY+equoHNFw1WFyWzn2fUA3Gopbt3XVofl5G35wtCiFeuSJtm
iPKOvMrmiyWvOALpHuuxlKxbNinoCEJglrgCkp/704q2Wy23In8YujLgxYqSFrwlmA+sTBhwYZ/B
Z5ES0lYHPlVc6azkeKk/j9Ina4520Ntt4jyKTDhWN55EEAvVwAw/BCHGB7HGB+tjPf7Q+1MiW2wf
YRvdTAmCqE6M7D2EI9TSbKI+xzHLB5nWlS0PWKe/aeJ8EJlIIleRIYA1HEK2jMGuSeRvVk7oPqIx
yvTO/TowQVruE5d7XDdNXS00U/L2afMbFGP3WVlxQQj1kMZtlIJcdLWtNGtjvu/raQc/5vbUIgOy
80+iVXHJkt6KBd5wQw6rG+vA4YIpVuidzDa8mHjceBCCgfDBMI9gE20jdzGbrwAoClOpF7RuWkkp
hJF8g962sZEM4FeBUIiactJxn7AwZCuZDPpkgUIwcxzBYaZZI8+f/DWskurwR58znyMD41yO3YTZ
cGnj1/JJww3ufxxHJ9GIoJ93KFMmpA5n8V1+U9/c0BxxAzhhNKElDRrAt0hBvG0Rp1989JtkkzbN
6mUlNfhOjkrh9Zlu9mMp2JG9KRo+Vhgm5OzPH8v1IhOZ/PRswbBLVstrwBkvolqm01PsLVBUWnXI
tfHGKUtvAJTMMi360NYnrXP1c2NKGlSrzSclv8nY+Gy4o4QruuagtSMn2H51Yr0mwyyWQ2km/Nss
Np2+eqBzPTG5e6UCarNt9+MGh13GYtbWgc1RLoF7ZzeWXwVDivGN8/sf5/3uFdzyAhKL9EBTbqBC
6TWTIGSvaZO0PAllI7AqZx3TAOqKNB/Bncn3A/mlQN8m+juBF1bVf+kroidOiEDafIoAZI8Ctg90
uCYF4+Br15I0eIPpvQH6bHujqbTnlqpd1w6O7VVbUnafZhijcJ3HGbyYNRjUvvM+xeumerwxumKb
iK9NiDttuw8GIEuxS7I+g+N/Irl5OzIvcvIq1jMw3u6bZRUx+EVQRc8Y3N8NU94nP/GhB8g5MBL0
CDxlHzkdMrnwrnlPER1qRBmlTPWQBknebT2pF5h7VZWSevejO/6DAntbM0Y5O9iNXvGJ1W21rHll
NVUZRw/VwGN918UUqgz9+Y7H6wlm3CFhMiRwnKZovoJHNP+c8LnEwy5iL+iB63Lcbezh0/cXfijW
JmzKonFEchGJniDQ6tfrqDRAGzixOLgr2adfRg1hLOoDxuehHVfD5r0asUG7nH5KWwo+kttvK9IE
csXt8989qyX0xJQRR/1A0abj6PB/EdVm7isRQhJ15L7KUSBCZVWW9tGTiKGcT+NLWGVi5dZ5TRqn
D9aRnF3x1hUtRUho4TiCnEt3Pu/jbOpqxnnsjYDKyGeaARVNNDWpLbk8PbOZrY3PJ14KmUeEha0T
R7cC7t46faOVP3lqZUf/7vOEv80COxPAq/uTIuuQvFqArbGzM87KzVpVV/PuNB/boXGgHFU0YrbJ
hBAp+cNj7LC8b8bD99cFLd8zQztLfH29G/wpovqYr/XcETx76JmzFyohirDSGNsSY0sSHKXnDLBf
QdY9qypVkhb+7doX4JkCDKI9dlGLA8H24umkrJ+qUM9HiVSOizgl3+gAcII4kLHg2vVWKhiiIqbk
gqqZ+J06zdyoNi748Ulrfm3Lbh03oDYtZoR/MsPyi3RTOaIjpUjfsw/mIFmoBRvoCVpMJLSCLZqR
8S+Eut9KvDTUnp4IIR0jzvIE07MBqrp629zPeKxMZb9Gs+spRDSqloAHgLa2Gwo2sKdmaoDr2lKe
Zg2iVrUnWz6MWsgpGch7eA5tmZRR05ql6bBKAibVWZHtfhWMxg0lihxeexpKV6XpWmSwZODGZM4g
MoJcRinkRKP50sOMd+45GpkGiBIxp6O+8I2i2oY1wypl1EUUn6IFVd9qXbuJEDQGJ7g7Wx6XzcVT
VKRSLCkJV7PRiLBBrGE40qchTRZcwAAy/j9YvKW/GllFYygYl9XopngTWgcVzZUFcIX1IEApMfnd
FnPWTlBHvUStQbKM9Q1jVtGIssvLMHTX9Q3avKG0eNEh1D3M8fyOB+6+egpZerKuT+nnnnAfh0wj
sIUCz4ZFiL89zTskaXeOPxHZkd4TUCNUcJZUH5dzqWyr1EHzqF4wHWgPBehhxRn2E0VVrQQ5ZcoL
2W5QGBGXszkMtYjH6fvviKn15wMI/PMx/VynJ8N708Un91seH6hzggzyG4a2CqUDyRq+vVriLQLx
9mW6Rpydz8uqYXzVg5bzRb7nwuTbeQEQ1zV58dW5AhQnr/+EVeOxikhhqF5UTllYk6KXh6OdDo85
HfscDr8NC+R9eDhUgcTgZXnwDVqvXY+nU+qsxXzIZRZ5OmhTjiPL8FXv1gEp8I886tZvera0IY2M
d/w255WQ74sVbxoFYvNGP5PJIR7n08UCGuzOxFAfBkNAV1np2wkgbJmDFa+mfwajPrTd3dKaoDPC
A1bRQG/NX0rj6yUNLVKUKfkhr8aKzSeoi4EBtJg9xRBOyjKVBPLN008zWnnmSHHNxKn/a/u27YQA
PUHuhXQnar+d7Mu7OWEDI0IDXBIZHzSvus+vXkb3sUw73pkUKZAPWMric3rBtRn9YAJqJHBkzrlj
UH2nu8/GRYlRrOoKYX27+sk/BeBQPT/5bKAwhFQsHRIxHX6jOSZtWnRXSSClP3vTKdAp7sc2om3q
WSPMuiKb9fDypGcrT9kRcvjaB5PMlxRs9qQXU12YESoYie3jlf6NDfVKktsvZD/3OWMBt6tAnUUo
xfQ8uqr3qPLtN0ECRygoA+yXqQDEFM9P4B+wxY0nzDPiBn9+X1OyEfP0aHXhWB17Ag/pmEo7TVwu
EOa3xax97KsZzbrkPkjIFFqIK20vJvnGSd1na3fyI0fsVGN2g4GOmTNfGv124fOMLXHSQwm8y0Ic
fexPXNRebpdWoxVSFdJPMO6qUcmTJ7MzrhDpkAxYNq1wUaeXE2V+R+BYC3lseTsc2QGRLauppSOG
jYnQ1a7WYjv8rSPnGyCYXKXPt2JVIiatjMSkORAQxEQMB0gY1v2M0ZPCKzTo3ONwRLb4ZEoGpYU9
pLy6Z8nkOSy6eQeBdNq/2sHm0cfegUCiDFO2vum5cavxv1Si0TMjuGo1RnyLFyr/RUy/YO6QXKr9
CrE6IZoZ9HIWFXTcr85bzLkNJ2Lugt0ACv2VX58EHtoJ+KIh1P2hFFYT8Y5tjHVf5uN7GN4A+PyF
KCrs1zbMHz3/XHJDdmLKzKDWl1mS3aNwB0qFKgJ7wPReFe7tDlCsNShbLUICUJCpVbS19hk/iFHi
WKEkLBZ+WVc1RSakGhWu/+Poi5BfYJHYnyxdxsRWu9AL3zGYjwcfR0TLw5AffrqJGCKy0hqTt1Ub
CjdyYXdKGd8LmJrQDsQnIgp815d5gJaPCBgBFw1RmJJ5YnvgcKIUCKQjvkHk4m7YFqDr6MBFZ1g3
AIfX9mZznvCCLlb8yE6Y6mD86WxMVm88nthRUxQXwrZCVZKmd/P+YoUaMHOV8RYiLnnvQp85eI//
H3SF9fhtJw9HesfPfEaQ03Tgtk2VeRA2Sgm459/cvuM9TcFzykKS+bd2icOM/VBj41cPo1YVg6Z8
gmvljIYDcVhAYzq7hCyMdsC5iD4j2YCrxolXGg7JBQdPssLx3zyRF7/cADkqzIKk7+2gvkH0FfXT
dB0QGN0adS+XH+5ErdYJ88rwoR2PfKcDTpIe8acEWKp3NTl7z/7xYpjhMV8hOeAU3aLKWh3NEqlv
5RLSo264BdqFcKpZeyK2yWQlOHgQrt40wCvA2RLRZ6AwJbRnALMcC1uX0u10V9uXcVwMwxvqAqw6
glNYLonYMe2KmYHRZJmeLHzX27C3Yd58SWfO3Hn+k+OFnbWDbEkBJyGMK1DDDo2uTZ0czwaakLs6
ZxNVRy7gXBFfkNa7opaXEX/Rc3kUbVJGFb2TIFXPddaniu1V6dwetIwI6up7yjKznLU2aJGjFMO2
n36eccA+U3MEX7fXHIgY2728uTyHckpxeUjHPr1FToetPQYLW8Ysp/oKHqgMoSgcgKPIA8jXW008
lcbPxZ+cvd11aB1WAci6+gbFQ13g9YUinzB6KQj7tekaaf2j7Tv0dPmSRfqB7SoPBg2HcFAq8s5r
swucFTWNBVwclGrN8jl4afbYII4dXtFLJO6R1Oawd2MttMVT2n7hli33glraWzhx30OTso68MDoN
pfntsjC3vG/m0yW90Nih/2VkJd7WXoqaW+fvdZYSomAR+mPs0DEXAIcNT6Udn0xw+xwSfJtNuiva
qs++zekPgEen3nsR72Wlkk/DWA6EiReDCejT707oTv1YmjYOJjxI3MdeJC2LyIjv6Cl+WtJ97+6B
xVgPWyboNEkbNHVNYa80HX8UpV7UW5hxXcn63s+7AhMiR3Rzoxdxx4aSHMOAPXWsmWZ0vjjvnLFp
6TE28Xd2PDU418pKvSJaxU+QS74UDGTuMxXN49KMs3nNCfeHXIA+Ysz7KHcPTmJFuwu8ZCBHZP+a
Fub46zj5PZCChP/JkCtvdw7N/hy2F9JF4lZ/9AdkKa9Yx/EbkzUW8t8v4gtO2a8b2bAJMSBb/+/6
dRoqzIGRB9jchcjhaJC9pMrl6FzdOit5FxHF+fJsoyU6iS03WAHiZ7kDHWYYIDBwc+jP1Mx1KBqX
iJT1VhHkJCsqlOc73T0k5tFF6X+dzd9t5ZgAmsNwH8W2CoM8Vd+KbTPlT4Ba2FiHD8BoSAHqxaqZ
V8aENJ5uwkayGUsLGaOvqBnqIufzRd7LY8r6wfXBvLjokkSm2J8pGngujTjTCcKNlkbjEAhqKF5f
vegD0Z15hGdoQGT79aT39Xk0A23ZvhE3BRGn7gbXOOK7wgb4Qm3Odue+HWOi0dE+SLcv3z78br7O
U9vKBbOAa4ZxQy/oiGBIv7CtMMkAPtbXzinDjsfqvgSjsjarAh8V97nu8BbWLeeYoviGf6Xsc4XN
R+pExS/neQ2n5VfqnLJVT5TuJ/Ac9C6v8wp6+dEso/mAJmGHrYhwkHRHBItmRu2wopngDDcBaDL2
3VLwNkqbNjhuaKGO0hCPQAa6VrxNeu4D0KozeRORa7nLgMWDoHryau0Q8YsWiXYVPBkP14W+OiMM
+meViBLd1kEKu56vZBSFMCrqwIBh3NCi6nFvGUZrNlDdEFBU+flxyMMOr5ZEsFB34AghesWrA8n8
joO3aSIyNNum6HVlOgmqhnKpbZaBtrKJlmB1LcY/U1E+drGWw463j7sj6/n+n4yzKNnlpKlHMOwh
jBAmGoGTjjBiJnjm1oeywxiQYZ6UZdCM8WJqT66w4Ifn70R2eqgaCYPjACw9Z68DA2UKUoFuDmpc
FUGt0/eDqMrwrQCOphVvRouOxN1FoHoXYsjVmGfQrhDvBm9z5zIYe+6JF2MSCFpgKMS05CLF14jf
xOOZiGkLqra1ze3zL+ibwSc8c0fg/Gkmz8uHWCKBcInVJUTMe0GPuZLlL/gLAhOJfUuNDuA/BqCr
reFf34se0eIQ9rM+AGmP2qXNPvH8D79GMbJVKj9rhFER2XiG29ogqr1BzDHOXaMHKOpnQ/dIsYC4
FLhH4I0/QftieFZvfyrb0ekMYSQfS2DtnFdVFZ7iUbgXZuIDT6WtwEG1G3aeY4gfCVXeCq1tHvkI
xIOnkJVVhQSPznBVUTlNAZclWDMU4GJoWY66elC3UrPj+Z/Y0lbVNfDFIvXR1U7dBWApr96Ct2Cz
UjYIQ1tB+zrV5pncW9g+cwB6w03KxF2dEWk8Z1nj2Z7B6FKnsyJa1esl+p4OrdYqE1V5qR6FB90e
pxUasfcErz0DsT1YrEej+TYBtTgYwcErjYKH4IsZtA4fs9XlCFJlQBGwMShm+KQMwArdBITdGuy3
ryUHNq0VoY7P6f4OTy/oL9QIfiVIujoVSMcXs4hc9SlM8hZhHnr+KXC0uIt1m/h2nvu0JtARgCdJ
qEByW8TbPbvTAJqfuoeFBQwIsYhNP81YARfYon2IdwpOLTyBT5Af0O7KjZDeARe6Fqc0Wht7XvHA
D+dk321gk0haqaq6BMBydrCaZPamQbRjYxdzEonlbQPIDdc85cBjl4chK3/lDL/dRj5Bg7vDI66X
jaGsoSZnsMmBYJfE0LW7y1foIkiCyyqT5l8QRE8DVWJICYedxsa7pAtk/cZ5EHWjbahK0kkMQUMM
s3ExzCE0R7d0PogwH/Q07DbY5dP97qXY13c4G7yRwyZU1Gf+KR2JW0TTxshOrJVARhUcWEyrO/5z
f7qm1ZgrdAEa/vjiURJhBMhRUFom86yjGBjP6uAtOTyPJdlecWoO3K78Y7U7COYjeNDz8uv79zmi
QA6AJqlrv+50y3EN5PMHsXjWpTyoma6IRLN16KW68DE+vnNp6cf1Qbe+xcnkrtqKSDJ2BI9837oV
5MzsJuRBnn+VBWsKfb+GapOmVznJXL/H7ErbHsxw93CNRMmZPfOwNOGP6U231s6pvntoDkd4egA3
LzwdiOAChcERr5AOt6cJb0gM6KQNEpP/66OqnWC40e87BLyrSNksMq9aNFVViF9XeKOAjlA3Xdaj
nRaM1x07BGad8SdL69t5mhdolISJFOn4MooO9QhOCj4ea+EMztHrmd5mIaXQBffaL2zCnWI7kb3r
mkkZVH+yYD0iDWgw0Z5Riv5tyNL68gqzwxwks7IlYas3C+/GfRs4VWHqIsF+TIHfYVdmDcJjdAqS
cgCRugE2yZBS2LuR5nYFw0mBUYScqYG1ViS4WxDZimsd3hmc5CnZV4TCyUOw0aqOg+aN+nnMUdl2
t63zFKsrumgdIZv1fEL/Vma8lqHUNZs/MBOQQh5d+PSC4gTXRmfMW+Yv9/W7aJkIQww7cmQ1WdxO
//xPJM8oLR3MT0vJmcr5qiF7vpzyQv8lcdxPuXW8T+v6kAhz+WF8UbHoSyhb/tTuFKSsHHNbEheB
TV/Frj98x+agIQ9yFR7DhiIsPidHCdMDXysqDarnIvPqUenIi9ag5H7G/ENto1rw9uMGEqjVdocU
wrhp3p7uaFeiwW6Io1rz8ApxJcVKSGAwSRYbzU8bhnTL7x1OctUFzbpeQe0SVxNAFEVIT7XUobxN
Z0oEQebcZWjVwr2UQUr6NbvuGEMrahqEvnwznZM76hfN4ypF2MqDTHDrCrZUysMKMtCBU6zcd7rQ
n5SLohVmqyEu7WEeSV2Y82qkNaTRuaWlShiFhRGgSJrft7bS0djJR5HP7Vayr1vUA2+shrjz2Fxi
R4l98DzTE3Etdp41rlheLIC+RHqDlCUm5g++1oVM9C5VLvNX7POsFDkg0vEZcMrMJ/G3vcDhJPuJ
5oBy3ujDDRFbozCx7VYjzeY7W6DE/0+2zGzk+FzdRyntuWPWJMFzvW30CN34ZOWF9O8wf8/6/y+u
AS5XDR0pcHVtpv4LXFssWl8xIylhL/iDcOnJ+S9V9Qxwl/JbDq9b059TASPqfHJQTZgIrhO6rX5k
0BcLgEhdV7Zu+R/7yW33oy/KkzcaM866b4FVXeY85c717BaS1hSI+kB9w5cN9DaCZVJ5WHYQL6Cn
QdsZBkYltadtxnkD5B+1KmpBlm2/PGRiMcS7MGkk3si4rUWynuy61NnoHQHUW+ll5t1AWuvG+fLn
OatKYSpeI0NR0kG+U2qXpJ45PItv4voy79BiQTXZ+wqqvRXjDbW7o7XU+Nk0Xyg98ks86gPumAmx
UEjy07OTX0D71DXIKA3DIuY3VLfN88NJsmG3XP4Hh2B9BeI5UVbWIAEe9ky4Mxj1ll6xCw8hDMxN
4w5mD8W3jCNhyG+AoYvTH6cW2uMr6Q9XhtPLFP9dqGa2hmB48keDZaYpry26+4sIRO7MBnLdj9ks
qZ4fYSIknnMuw8o9Yr+RxiOVoMVMk+vxpnCQp+DG5ggvSyDpDolefQ1xCBf3q0d+dIJy6RHnyFqb
3wPq9LH8OVTDlUDdLzn1u5EFcF02bkpAwY1QRQwjbesHfBF9TYdXx+v9Wpwv0GnwT5wlf30g4sWC
PwWJTDibgzu+IqFe9JbFfC6eNsGMfRCqOiSip8vBk2X2GFhC6qcqPVhdcrYYNt6yMGxR8V97q4HW
ZNt3NTdm5q0E0cC6QXCWZCIdziZ+w4pQBMGIcylOPpKOE12CFdkevWWAUqd4VVstZg5JgBnPbhmK
YGiHigdGeE3YthPn0x2jI1h8vEFNKFzOJrfAKaFtIx7cGGha+ug/3GMUW6eRLWFwkgdHlSMU3hNj
/1Xbh6NB082dtDEkdbytzqV1VHlc1Vl1mnCld8cviIkC0nw5kkg4tisNuCOR/Q50tgQ+zZvM9q3f
AhPy8uJ8TOS/IZqH+OMEiOTUKTSMuBanu/ZsTSdutkf/rgVT24EjvytZUJ4hkaXEWY1nhu4MWchs
VT/1fKF6iFMc4UHSVfHYDQgb2WC47lBxA55ClxO+xNoYN/sm8jQXqZodJe4vM7Q9WgwDrEQfiRBA
DmzhQMIq4T+N53Mb4qhuQ323D+q9rDLG3/O43RvQ7T9lO0NEUTG4DUAMefvtnLsOsqxny9P4qHOw
HoKcywN9IM2pSXkGXeCQNP9yWMAvdQUFTFKeycgmhEKkvyai2UizkqUU/lTr9Fxxe6BW763QuWeh
xaIrv5OHAaenWikE8SOw706rviG7DbYnriKJ53kSKq+Vo7HptbDC41Ff5WRWZSRoc5jBAmyBd5M9
qHQp6MCUj0BlKpX60omv3olrC+ehZPxNDpFKUQihghvQWhHGoEnud1j1iexWwYwVyJBkhj0pPg5M
Vkx4POR3JCxOOuq4F3etncjCxN2b/VQtTAUw2BkFL+fQverrMH0zgyrRNHzstdjS0FPr98Xkej1x
8UHsQ0W54ot+1TVtx5+SrNWKAKCpi0BB/LAH5n1s6ae6PzvRGfrIdzVVF70Bv64PoszgYhKD/4pO
VyMeq08OS1tRAhrpC4ePtFSe5H5iWqh+KHmkKvlDP1HieCiXA27Kp4FxxBnBFLEuXmnyBD3iqCZ0
gMI1zSFMGD1LWDxiLi0W7SX8q8wHZPp4+UwJJN5mOghmn36VHWB+9lSdU9o9XDnxcZCzDTsfFE+K
XX20TwRM+9OrhK3DjF/Wiyrn4qb0EQ2WVjy4jswqM67Z+T9Zvhxs42QWUEiSqctHwc6q/BU5vQUs
hqEP0hI6STR48S3+nV6+yWkznJM1hneaZ7CsXyCdGCQ9SUg4hb4xOhK0eBQI7DqgChCLNk23AWUi
Fdw+Fyh5zCgISoy6pKagp42rcEhsYPOZwD8mqAVxuqLnuk+lvQHIYS+iK7JZt4mHPs+M7EFoqEW1
5p4qa/snKOg7c7zNBKv0Ij9rGFPgnYDI8M443q6AtEHBJB9QCFS+hpQIABcm/3IGHkh2nanBja2a
n2wR+33oxmaDy3mYf9edPj7MeEejLE+9ufbr+50qOld2JPimbFTyQ6TIXvzO7hBUKzxk3OnMu3U9
BYPcVwyw8QXIkN3qrp4OvITxoZEqDd/lrsK41ma600qzQwxZ1d+OToSfTuGsne6Kv6pmrNOOpQ58
w9bWGe619gIv6zFlyveHxVC95hQOP8CtbEiQ0226AuIuIBLPVPy49Ok3iROeE3oxPvIWVbRa5g8o
bWF9vQzhYXv8R3x4rwXk7BQ4fCz9AurJrBMpaOFQ0ZqhYg9v+qFnfZD94f7FtMc8ogQYE5KNaePQ
cttC4owFzCxCIcifAEIeogUnRv1LEg2cXdw9j6PI4/r7lMhfhuT+F4IRS/nqGLrmOcQoIt9DSuAS
pnO9VR5o4SIwSkmA1pWtWjMeRA6ZOV2QRV2Qn6LoH7YydrKHVPZ0cO5/lF3iJi4J3nZHuHbBWFuS
bjClystdao55KdaAyH/MjDypGmLXR03iYZX4/9DdVIT8hm4i/HV+l4nIFYkW2LytVnlU7RtF9m2f
MYE3s8ZGtBZorxzhrnLFPR6V6d4B7ZJy4bxZxwRja/tQXay4O7WTr0qIhK1IR9wcFpWu+kgz4wS+
KYj5j/BAKI0lY+OyecvLKjvtJfYUlnuGcwj7bD5V5lAHilNAx2NH98YN7e7ioCVOFPlp0ZjiuzuI
jORNx5KPk8t891GSiw+dTaCV6WnFwlGbyYe5T3cHvRkT3N5atRh8s275+CL1fLLss4G/h6J0pRKK
hWBRdVixCj27h+a61wC8kTXVrL83QzYKNeaBf6+3Cl/96FgL4wDyncqPGzrIH26sNouk2p6KwTw5
cHEUaiejuA0Qvt/3kNtnww9/i/eUgu1cEBmLFXW9ZFNFhdU6U4OsEwmCS95m33ETqv5XFRbad+5T
FiZaKatPf0WfAhMCuNFOQpbbq+xaD+G8aWyTJR3ymUup8KH82RIgDZO3QHYWha82n0oBafFokHwO
ZN8W+p8R0oirwU2lQI1Dnnit9deazTzmyAWzWRms/xBxFhapG5ACr0lU5jVFGn1TSIGfZguIM/mg
tGGyH7RUspBcOECJ/l7h1R5Q6MvFtGdghq3hvMAd8RQukTT8oim+NCLFdzI7xSDXMEr5DtXkkHPi
N81pHrU06cg/gK9NjNvOK30F5FE2CkuMH4ihkKmW4NYJ4UlI2jWp63hLzf8qSHGT5OD1Bq3Jm7o4
KFNILNDfgasBILddzsIHDmbHgsTF/ZMjlrY+w8KZkfro/R+yR8hv7nscuz3BTvvDwHrShFGe0a8T
nkLuhFAzBfIFx+RavxKK1WGgizTG8fjyQgo/E/RGDw35PJa+nZxbKwa9K8bPnn8KGKXl0HBsHRgc
8gUV+pMWuHlZucKng+eD7vQzahFychm2t/OYHdJRNMGb+9mEBTEh3awMAchGD3HVwCepbEtyflve
oHwux61hO4EOqavTqzH0D2/nvkacGmrfyjsKRrq+V0A2mqwroEZvFpfojRT2PjiGaI2tA4AvtZS2
891Vjzm8YqCdUj3a+yqAjDonpKtwBk8fT5a9ni8esq70OA8VyJ8yajdp4nXNLjz0ev8pqTpewcXG
EvcR57mT26XKtMf+bkT2C2Edma7VX1/xfQTbvEQnj0mYMwEUGAa9IDOJwxaoEeCnkWjWIx/H58wq
CGKl3t/EyfDkhxVTO4z+Mv4SN0nURuS/aYoe72qLiNe915MoyYryFZ6JkaQA0egI3PR4jcKythng
Z/4dea7ykvj+M0RJ3i81xE4Vpb6I1NQmFvesZB2cdtZML3Z11iKleV5N3z9UPzPSzl3Q0Dqj6HnB
cCu9xfWOrpuVs6Lk7tbJ/efTokmKmcfk0agDKCtV40xQ9rPmsJFPbaTDpRU3+8aLg+pKR+Vo2W8N
7QhAs6UqXeDQr75vM7hNLMXVA46LHlYoMLa7lgxO8CrGBtfhcCo8Iw3rTP18m3xIllr4kIRg0hwT
f+/BWL6w8lFn6nVCv6RqeR4ShzqiqruWjNvVpNhjfy9oDCjSvuQfrqMVnA/CGETczU408XE/241y
ELUCvsGiRgZDruA5ouWGKPz2itHvYmJF/NXbw6i05QqLBJgMQxeH70OKM/vdpNQ7B5zS5304E14q
oteG7W4Xm8A4beY4Ma/6+ewTSUzmrwxzP6FG/Xl6AgBWk5WuVROR00vnDNAZ2M/LEo412EFmQqsc
BgPe/Ya/fqsw0667pS3wKHUULJZ+Uxkowdwfax2soY0Oxom70sacDrHN6IrQmZyk2g0EdmDOnVXm
cNME4b12/uFI3oHJP+VhxQQyNolfqbrCf9C7M5Sob8EOtq7NdYLt1MLpzpQmQ867/u9HLkECbR46
6jjU3tnex/A9FbpGPBx/nfu1oEUimTINZaCLzhcbBt4Sii+FvVS+KhHdiFTJgUIuHoneDIh9+6mM
wqX1k+XNPVqCr8vAzn41bzBMyRjovD0g7byyHrkGXpBg6XGAEK9KOyMQeVa2Rjo4iYvmmLoHsXIn
MRUngQsO3kIaYmnHmsbLJdSee5uIBaQsXgpswrAc59d/BRfqwsPBEBGwNssdUkzmIEXKRb0TvKEV
IieXiB/XXSOq2qU+mk7Uie2IC9LJstbDO3OH9a5tLoR1BjauIOvGVzu6ewTU6dHs6XDDFlmnEQsk
SboIOaUYWsC+b51NInrjzzPw3393S4fo7Gu/F4cVxvQzCjl1k+urgmr2HL4P6y3Jrch5Uxa2R5ab
0mxzd7qT0nrBlkGllhG4W99T4D8d/kSHnn09H5G56e2CjC9MihvFbTHKgyA5chkrn949fUaPjmyw
mqkh9sM22EJdkBWJh61hs8prREr+WolpxB1rsZcfdyRcDPOfVMyInJDsShb6Ik3FtLGOjMGlofrU
kqp5tw4ZveIVYJWFV3Oo45YRpohlx8A8KXXDbMjLqr3xw/0cvRyEw28i8W3PplzP6DSGqGq3ERxJ
6A5U4RQ32hVBMtk7gddGyUXS+ewUGkKU95IL+2Ct5gX8AobjQ7/buvRc2jCC9Lef196J1nVNfDnz
P0R69sUr1EUoVBOrp8gq1HWHwGCIswceEIhTdCwf+Gsn3ydODzWu+aOcx/DZSoAoEBceB6hlO22S
LdgejDgyM1cmxZT4CmnWU5BkQplqKIKXIX0aC/h94QEQANyj/JC/u5W5Xsdr1EvhhRp6VpFg/EhL
frOoDqfsH76RmTNinlctEe33X01lCPOohwzA/lfDhkyc6y2t/Wy83TGRG+EgRwzCtbwW1wfR77gn
E2s48rU217XPoiAwipK3o3bW/yChjeo0B9nswNOv2WbC6k59FwJRgmzHLjgaC+aKZJ54SGdtcmxz
QNyHCOtl1W6eHg+se5V/DZZ6kl/kbQfODiT41tEGiQCX2D1wzTwh6VHSb3oKAg4vvA/lUyVSnPLC
OqwrORvmCOGoOfvsvW7Ii0Kr6deu3i2fNMDoZ//aqmTxXcm6+a9GM5MOmLGvJD+a2bazvY/Dagn0
hNDj3wBRx7Q56hDtW+092sbUgH2eXDvMVVIHNXLkVpAglXcDXu0rLMFltg/GEeU7GQYgzhj29IbZ
483xqHKU/j3OXk43ERRaIjN70LtbduhhNolpBqCxy9aDNQND/WRdTYgikk8T7oTlHYHuwMlzcFlY
UxZ6q18SPMC+Kv/QHdPgJqj9jL5+x6pP/n4GEXfvbYzyw5Fi8gQw4OeoMq6nv+lp8TO62DOI8T+Q
QTnmw37TqKIETilC45ZkuXZUBNHTnBJVKnNXbFXwFB4FTjG9mUUD6q+oizKb0wvfZo/hb0xL8EVS
V7xpenxMtIcl6FTo3zi5QsUb3L7Y1iNL/DF28V9I/Y+lumESLiIXkWSkyNp9/9gB965slxFN0zXK
/2frCHSfPDR6enJz8vM6i7fbeui2qqelts5gPbqWr8z8gvGlZfzevHFf92ANQqO5MnWPkAe2jXRk
Yh01WgMPQjcmWjQtjYDffTUTxPWxVoRxBKeDc1cDw2r2Mjcty/PutVyym7Diu7RY1/kIOX314tSk
wD/fYXiUffQ8ACyvaZDCgJJvjs48QtNkQn66vbKI/d+Wi/fYwDBBRUqCQTikgHx3c5DmXJgzJnfj
3ypISus5NDmueAgpLd5KjmPllPj3ewlBrewQGafuG4cM4Q64qRrKVhPn0bBKQ7r9Pic5/WuHRGUU
aKjGEOj4qK9CP5CZnyaHN4spyuoIz9Dz/Y0CpyjALCnkFrYNVv8WoTytvQZhVrZCZ089oxd1beCf
NbhbwD+DdC18tpIBa0AZcND24XDYkFv3hN2P/ERgZV0leBVox1rbuV9fGiOar/2sOiy/DRLXgTDa
t4hf8Y6TqDHWbhkFExi1h4nHOcfFMVoWWO+L5M8qQRbiiOQMcxDSmLMCKix5DqSO/NT6el3Tu/FU
pYyrx1Cr7KRXXPQwdIOU40lbCjTEh/+2LJ2b/cuvPcr1kQWFYmlSqkcI5flJJHdx0o5BMOeSk1mK
aR15nbHKDFfWeDTMa4wlhVPdRnnJU27LPJE8/nowur/awQX7m8TQ0pZzGmVlEdEFp4xhA9DNloq5
4L0ClUgcsLYGFAf4Ol5M5ypPaCLAo9Ml53TkxywPQ0mLnLe4wRoQQKPBMOQqmaBOFnKZ/T2U4laR
6DjARKIvPvBdywfC5J64yZS6OZ3qUUhpFwTn9CoCTVCRmsIVy2mVmRzQTyhQ4sQLAjxJTGMXoPEB
/lVrjBDJa5UeAyeWQ9oU8UYExRtivz83X96cNzMRWZOwpT9WItmm5N7p7na7e9YdvGx7mtug+PvM
8J5gIWSpV07wqy8xzBGzZlSLNe3OF86ibtXWfuCvjWdIvBl3Djk2sGiU2XbNvwTwCaogWx4CkOPi
SOyinBKfpXAJXtUa9qeoHeKs9fBK0dKD68ene/E3NfpnnoGsx6Jm/Heqh7+m2WLKeS/2kt65BIeq
bUTbjT+1WCZDrWufg149+bUnWCUch36EnxMUdt0CeKpLYBahA+Mst7V1v9gY++PAHv+1a8jtlJsy
0+TSPp2RFbB7W65szX3cMbsUpUBWH6DrwxNpEZ8HLAEIk6EUfeOaAVEeLRcjisrqN324CCUzq7nh
zMycdlop2mt5Vn9b88s+QwPbdbdW4WANiDs9LdSzEpeda9J27ddN92FHc0QboreqIlDQCjEnzyfe
AItscK8sC+TtRR79iEO2EhfEOVaaMMj0oStYO+XrBG9vJRwIV/JUXvSj5o+LDvaeYUvckhRSh6e7
SKxkMV7C4xyNjr/exklsgakeBdQJuBSj5Z4ppE338qxEXS5O8gp73n14QUulpTLZlXu7mzmTebgJ
iMeHBNe2az8FYW0r7RdEcEss2C4iENFk291oiG3MK+uRZZ/4HEjuvN9V4lBzU2twFJrBPTsPK86p
esgPJL4phPpPnffsNYAJoRHuDdCgDHMjxKgrjWsOu2GIeHBDxaqeDtfmHns5eC0sWfthukoDj2cQ
WPSq6QFQX+qi8xbleJ3P5T3A4DwjGIKqq5ZFY2Lqr9IBX4LNJ/FNSCFLlhz1xf+wyMvMJ0+aVzsE
vpbPPMKI5xv4D4rt/qgiMTM8Tkg5NgzTnGiy28Nqguic6GNRf2WeQrR93QidMAkmhG7JshzOtLeD
efiPdbOcVYypid1HoLd4Y3rry8PxIfP2LeXmxEbXOX/IjksXq5cjq+EyxMqDuxGPcQm5Q8J5Mirp
vlG5uUGvsQ5jZSJ0Rp2dug+lmKVIgpPyq0yXdkNVU6nQ1Ma/kSAMaOD6kjk4Pz9v4G6J3LpWvt+O
15l+7BWihpBld+5iINVSdTFqxUAPJxvCfc0b03oh4VHvRNjnrxcMaMENlv2xwM03IFozW+o/xe30
xzvOi0MdIXK9qAsdfKOGIOyn4KgmaECbBxdHo/G5yw0vWpVQrN0K+dzZkfWCgsEMK2InPZTTOvRE
Y4+/BCFRcHb8bJld5KXP8mRbcGLuvrWXfQMunGfnoJjo9O1EMJo1ocYJUc9EzHbub9H2GweM0SjU
wpfrti16lPQSDIXDz8dnJXuZb9UNUBZiGuUuMifKRRRekMCqoOZFPdd2rDD6/r+X4BrhhFW+O7Xy
TvCqlFWFOxk+HbWxT8oIDh5bET1FDQolqDG/bFJUmlyNafxkMxt2V5H8yjp60sao+Zyt+rSs+FXE
mGReTz8u+PuU+GZZWmgdTHk17w05n7wisDnKzp1t4QbW0vizuzrn0rDSPwfKiW3AoZsy35ZBlg6a
cEwxarFy+0V7Y5hSzH3n8wigBHcS9+vy1X2eTHohuejERsIxW4H2FAy2QnHRQh0wbMZKTwoAcqtJ
5Q2UjDb3aklKNl8/+WRFIb0A3fvqW7txvlYBoqQaeRJjAnXQfugROAvwE1awR/tCprje79VIQxJy
KRdCubJQxAsqKlHgBlTnFpyn+JoUO2TnsMgEH6S0ldvFBNVxK5UQBzcBlJursgJEuQQlhUmvZHYh
s8qk97olw5n+OR+k5UGvhHiwiINOPkvOJTOF78IygNmIjV0sRlHbLqyoAj/RT76uMMpay7KuyAJ0
g7gmEtx4AAZf7mfmzhBDskbqjZpoDMT3lXWFwt6Uoy/cfyB4daSoQfVMRUCERuPb0jg+bfG2P24Z
2vV/lnIFC5CQveH/ORbtMmvaWa8ykVZTZuIgx2rdBLbfRpJdh3MvXm5Ell7yDQpV6+HgBhOZvw6G
5opIldOkoN+oT40urh+KxIvfwd2J0hVT3fqcMV6E0V2f2uHwrPi6FVU6eP8M3FUQl4bpwtuYWxfp
15HPmsVbQuAH8mn4/43rU5JQRuR349dXyip0h73DfU/CCw27AGDgcc6b1U6oucFEwklNrZaPHRgR
SqUdif6iNatpstxOGc8MOBwKaY2Vw0sgmbDQLSpzaZThqs5ISPKkutoE0k6lrEpFm6bgJdObq1H5
gLcDXRHMbTc4ieJnKQzMqyyadnN0MhS3lwfEEivnMy0dH/jzptnAKC+U3IAtMUny5zdqq5qzIAmP
1R/9fJaUTMR0SiN+b+A6MlIjrgPJ0DbWp4LZgivA8ffS26AWnBUAyegWLoJHMoqHVNj8tEWmA3tF
ZaUJuFlc55BjF54tR5Oryaf9pGFaDsMgabDlbIK/ZwN+EoveWRiAeeOQGmzxjkbcD7JNah/6PDjR
mV0dVSW8aTA9YJ1c6TpaVOHcdLiFNB2a7FpZZkHT2LZpouVhpmEvpfdnC9kKVijuPN5sOLHHzQbO
E+fWr3nZ39ssqRT/Qtr83haL1RP4jvnw84CZbHFbQ97zXM+upvGK1dSKAs9Gt/ZuGgMk+bbNZ9bh
2hnboZs12V+FxKdHPpHKlsdoTjg9MJLRObHM4QuBfIUfAZnsP7OUGjsZJK8nEZSq+kcsl6viw/M/
Bex/nHL5ziDWeCdFJNB1h2X6axLsNjw4Oh2Ub7vur31ClCXMFnOQDNAzgxfrpQH0EAkVqS0UkF+G
2mnNBAdZC6oUKXgzr9bWkTr2s14+S1pNUwcdm6ehgZgWnR8XOTQGwGt0MgvEvsQeF/BYIwpo/6Im
6OQeZgRdAoYAw5SyVz4lV4fPgJxtrm6rbrwzdYggLEgFCh6jearowl/lP+Z94CLSYFQleSigc0vD
b9qkWVicNo5F9pMJS1rbV/PM3H6NoFZJqshJz9BbXA1fzLzMOqja+1RuMaocMdRzIm0MJ0xo34Pj
0tQlj0zWUf6e61SltEdGpi0V4BLrAqVcLYsPGdtHlCl1Ykau1oqr2PtL9Ie9sHl1RiJyvFh9X4Vd
Udaco2VGZ+AenoUTciOplImKskHnVqzMi8atZbP2c473yJspzn1d47R41Uc3Og3jfJbPCLPtCL3d
pwJw4MRrENMETXR7yaYASs0rm5iutjTu0WKv5ZWt72h/glZL3/vsERmrz7bDUjZSUodwK6ZzlCu2
bILQ5W1FtstzF/dkUmBgzdk3abDT2p2c+2nkB16bZQqxrBXma6CjdhJrwtzEa3fU/sx8129XrUb8
k3zMfg2Os/PkPdcftjmjjd2efXA2l5U31xlTRpSWSI4dtIIoAzWyRtLqMZJrjnCqxh2tUaskAyNF
zaBb5q5X8bSK3ofNSIcwIRXLiWkmQxql+MtSfShnbFOd4xNjt+hPjh9cpRfnPAtcEvlfDu6uIU8a
dNEDXVz+gPyqczZ92OKqzSa7HeknsBx9bKf6q2m1BJo1ENZ/t0sy5P/jrdxlxltPIdTNTVhy5kuv
1BXrEDtzVnLihOLsYExx0fYhVyKctL6VsORHpJxC0pQJ2QB/VWAZ2twewNsYxTbhsKtBItlb+cvD
CrRWwUluzE6hQ415zHU9nV6vBRdbP5yUOlNzKJu6RJeqLLMdZx6+gGZ/yfv2WnD2iRuygV7oPA8f
KZFP3qwWTs54O9PIrC/OTciP3k2L83NIMMB6pQ1fwo79mXat86F+i2cBS44+Sd+Y54jsanvaSv/Y
2vLt/3su3sV4uom6SpY8s6z/3cQjxl6LrUukmheGJC/lIwDnOMtSpzDJc7mXq5Z+MS7ZpfgoI1aa
9nvpTyNgoYLDaE/MFllBR93GWS02yNW1RJhnhK/uz3rdxz5iiICQuWaNCFansmHPm32WO1zlqB6l
8QCQNEfGv4NydWBTpjt1veSc3pat5HdKtgUjDr5O1MKWPqbTwZkBfdiOzMCFD4QA69BQtXOqNrPW
gGCMuPDtM7AZA/nNJSF1NW/lUH+8UM9eObMz3y6GbNP4b3Gpjq7uS3FJnHi6J1+byHmTCtrmfAus
zg5s+ZkYnBox3bcTkWH1VMC6H0Cn1Bg2yD0CkIkIUgfsoqBklCTtxuAI3QB20DhMAqz6wRDsfMVJ
s6L7U49aOFImdoylwNv76dwC6mAPiHk+DKpnu6dWhYVfcap+v+gY9rnjRtRRl/ikOjmcuqNL7vgJ
Dvz4wuwosb7qs+af/kkVgybFtt9UWXa6BeRn/WQTJpAA7Tut0Jk1Wa4dAxLWjRNcvKXlyCR+uSBG
OxunVVZP9gXIA+73H0bQe58nIJIiZ4XthmitneFaItvHklSvQfh/uw+YGG3ZSpIUx8iC6xLpYSeO
5eanDGMzgzv8fG5K9DCGKMmD+MAV5ebUJuV7yPGfYnDzwp9k5k/J2oPxFZS2SeRCiylDVy7aPJ/k
owJ6+MyqSWKFNY1Dk93pQUAgwfh/LehmhAs8w0ScGTwJhWb/9fBd8XSyv3Eiplfwmu1ake6KhhJC
gcREijr9Ain83jbS1aZbxlHdk/Srvl5TEX8EmTnFrtTOpZrsadWyoXzjhDIWmkFTHbFtzkYpi7NH
e36VQhH8Q35IFcvpqvj2TMWUPTrzyEmk/wSHJ1nTwa1AQGYpv90thG8D7I7XRrp56MIIdL9CqyPs
rPFJbmWToA2KQGUI2ESDoFZJ8HP9yS8tsZOIkN/KgM17QDPhP1cI0pnktwYmtNQtlIIGJMwB+dDt
SE02Kfmxn+GLKtLsbYlJ9CEHRMesVS4DiibSfSIddMBNQ/rJVVeQBJ7fFdeIEeBxN73dSouwQlJH
BdXPPWNQUYpxBFKsX7+1XsjqLHYhofHMm9QgA6DvdQmPBcj61vPtre3XletQI/IJeLotPDU4+pMe
nIlTDGJ3o/8llBOZHe2mdRmBlrlb17rOi9l52FiWZ2/uowCv+b+dxpVCM+ihITKxu6d0EIrRICJI
ZC7DGYnvxl0WU9ScoOA74YYDb8h/NBW9ZWrpkt1WOR6KoTyMz+Pldk/I1XaJcisSofJvZh+ZTLwp
HKHpL7c9PFBXBjZU6x/SDYePyA6gGGCQU9AGeWFeJQPqCTPqsqYUaPevN/cbNMvBtCB95uQdNN4i
1WJYE4OFO7qyYNFCsVTFBoEzdYnGtyuAn27bp29dhbm9PN81630l//CYVfxcfQydzX4/4mXnrgrn
jJ8fZ02hI2/FJAahdNANQveOdGpvu1XM066pu2KJf5CviKrkz1Xtybtbg58k93EQtSBoHOFVDxiy
9GpAUTCg3ntt/vGwgNgQPD4dv6oPdcqxkQ4Bfj0Wu8XnTilu8jpmXgjPeUvOxySZSOlmfu+532X0
In741GaI6L0w5K0lmdG+jKW0d49+NJI/8d/nxY9agFEhdrfKeRQMM6MEmQYcii5xjITHw3PTtUoV
a5R4FELGttYzz2Uid6V8LDszzXE427kj75vFihbkDgu44WfZu2Vy4oDcTSKvyyYg3gW5P733NFtD
KZe8zL6dRbAb6TCJXpPvElPUfy5HwAsokstngcMiUJtedqT4rrme4a0HfypbIrPOhgtp9FgtSFqF
G1UGhOq3cQm3m1rlMuBg8fBvRXwFcXe9gM/kvzRGZRp3sJhSsG68cgItyQrTCIhJ2f4WP67VsBoB
omXA7DFKyZpDXvCKyNRekI2UnuLF1pqJ898aD3tTkinK91oZ8tzQ4a+GkIbGC3z8j9Z725I4WjGV
GkduglWGti8lPMGb0YTx9/XDNUxo3hNqV42RZmhV7XVTxc+OJEFx+rBt2baENYMDRvmQa+J5qR9E
pftVkBJU5vlojEE6jB3TL2AnC22ai+y/5ERJxP453qWxt9DwiVTnLX+jIpxl+/pF/DEq7Gs3x4VW
Fd/d8w+dA6KaNam2mXy4KAGcmIEi8pBVML2ZtoDDT2s/yasqPon1YfoSN2CaGIg9KRFFsF5QIKxC
MrCsicpDxDhTjBdk0WOKOfXaEohFCS2wCuwHaqK6Te5Ft6qzmhQhkrVk/L3ceeJdNKZVzBBbfQey
TyNV7eV06kDpJ1xv1GC5vCh8Lth76CVPVXw3nZ66X4eHdocPJFHGmEdzVo4BZxKKL+vB5dC9h1pk
Px7XRy/S1/KAk1L9J8eTxfVaHnSjuSvPmjKcI2N8BHMaoT2wtnRiUPRp8YE2yoHj9ZwLxl/1bIYV
/8XYHy5Q3oPR4daxxSb0yEQERb4i17XVWaUQYU6ulci0J25UbBtM0jN2aJdyfvBiNjfTvS2ib60F
xI2gL0VzkJcxkcVGNRbxr3/ORwEYLX5+puH+S6lAwU/pkqiwlFuoV1s0dc2s/IaelvWm+lwvSQoq
0N3SAD4V5FAD6IeV7viEpxg72uoJI+LQ9KiZvpmpOICtlXoxqG5MK0JRiu3S26s2DCh/1IdUi0Og
42uIbeOJX1BU16zkkAUoN3NH3VDgH6GAZmXUMVADP6S6/vaemq812CB2pbNadJdjtg1I8FBCpFFw
SEyqjkqnWHNcCaN1rVdOvUZ5m/zpppJxg3nkE7SrkFvFicbRnrNNgdgOqwk29MNo7DtdtyIT47Kv
QT/2XC4DvllEyazmkXCK3GZmK71UGqXLJ8/0fBYXFG0M3KyeCkLUliCwHN+v9vgNJtKg0ew38c5m
XGE4DuaSs95AoZCOSR40EcDDeB4lJJcf94sHciAcgS33NzXFXTthXM/Km9HHjH1nEVg4PHGMe44w
kdZiaTkHsRy+Jl8isQf/U2geOV197e45/fGXq1x438QYdNoJgzB6yMZy5EWkLZE3dOsrMfyMgwbZ
+X3Ag0XG2C2yMzyPvzyTFad873kixjVQR208m9YKjrYvXWQy59bIyqujQwRN9+2Bd/PQVZQT46cE
lgTBdPyJt2T+jwR7A9QbzHjql//bRwqJ9FZ9K6a7MrpwEsbIzVatdD6xRz7oUq4ZMAvCdKulaIw4
/PFB/uPVQ2jndD5cOMaj3HYyY46fUsyWCcQUBpTnSomnem6N3SRf0JtiRiwFmVkGJg3fOPrldqkE
JmoeV/jFdXjV1tYvMODRTZajrBzns4ovTEb4E9TEdam3FDfFqcxMAWzZU3Xk5CVKrOvPk+w5L+Sr
U4W1AJ5/HjeMDNmDTEFsWw8T8/v3wuRzbATzenrXUgX6wEraE9y5OSnImFFDLkCHqycXqK5pY+UU
M5dgbbk+aQZpW6m3v6378LIouQp0B24+/eU11YpT+txG8HSJV31LxjLS3HPHpu8M/RcEmNXDT4uG
3ab0Pgf2HcgTaVl9YZvz189Pq2ovHJGPNsI26gv7fCWaf/U6dK5NJK08rIH2ryKL6PIpO2kEpIMM
XYN5f7KzuI2VbVcs9qL8KY3/LHkJ5KKrRUwJVtBuPByJsBUUmYv/FVamuMcpropJnZkKqlHxpUea
kPWCU+uCYMqVC0vcDUPss3A7GLvJ/k3F4jPq46knkv+YmNbFbudGsm9LM1jCwarHqCCKpZiR/cqh
b5q0enrVNfJykrl/DZO86WwtWfw/W4Kowl/S9vX+PJ7f3NjycFCQoxtlg0flOAimj/N9Fo0+C1N/
gkGuLMbU9yL3708mtP0OC2fasVtPGA+4u++xFlmWNHwFvoC1p4Pkort75IqvR89hnMKPqPwYSBmW
mClb5aY8fIa/eTDHogLSeqgLxDGq33rg6cbdgzEyDLF/d9HYZ0YcF62a8ycypL95pFkyKDfVlTf2
AZbv1pnsi/kgkYn0FxKhSBC9ajgdfATtBjILt35I5XcTwYdVbM/NP4ILTvrYtPxmi24EG/wj0Yh+
H2f5w04fXyWyWbEnokTrsgc41ezTEbwmu5pdw0u+mwsU29RBhUm6fJroWOFp9wCnXgvR8jiJKJe/
AKT7GJK4wiMthRijCKp0cBQTGdTt+JeXQ6gqMb8NWCZcyue/liylTAnhW9jXW3sZgUOQMRjcHp9E
OW28B+Eu39mvrx7gE7B2mSPf+2K4O7ykscSa9lk7OtHUQIWabrSk92cC35JABb6ctx/E9ISLz11t
uEgdmO/3YaGhQsU+seR5fE8QWN94utN+9ml82h8s3dXgmSik4q+wdrkxeZnGktZQN6hL+f1FlkGm
Zh+SeLarxRdlmaG4nR30zqPRRJ7VYZgjkcoaONCdxT6Cnf5OScNHoA7Znq04TkDvk1JHbMHKXeT1
0EKO/Q7vNhI9ZAXq0wxFQUnx/4wPe6kpXDLCjkk1DJXUUS8QM16aW+Apq6GVL/9G/2jubmQbadtx
jFwJMHLAlFgKTDiIfTK+sFfkQ+0a42BBj4z/jAIJ09e9wdocGupvsIOH2ljzyq3VRaZqezMHHrPF
Hino11aILpXZ63BVW+/ddPQSFbAEdm9398nFMY33Usq2PbAm3hybOlZjGgGO4+HbJbZlgcsbAlaR
SgELoJunx78WpDdqs86+uTuPMpOUMXJ5A1nAM9BHagn3fVJEPIZ07MA/6bPmTVMRxXbfvQLbmTo4
gcyCb1ociqXj/NMmLOV76bb6zIXycASp56K1+cmtHbH6DYIJZIuV1nV62WTNfIQK8bVR57aUW1kH
BMuqIadkoCC/JnfhoAHFlYkCQ+lhGTGPcOnXI7Vmm8kbPSV8fN848cA5Y5aw1a5cFZvZ/oe5GwFA
+OpUEozjjYmaDZY19ZRH2pj+f7ZW3wZ8HRxbxxK/DWQrTzR4f8c1O9PrEihHLj6fCUgLSQDPyg2B
BicFDeIf1+k0jJ4Oc4tiBH1sk+CdaEa+7Dx2ZMVvL7OrDssqM181VwqFnLMvAfr2q+1I6uEZgHoQ
dLYWEaswXSq7k25nPhZkMAIDbZ4Eq4dl6x4wVarWBf7VAaY47DgXtqne2d5ujLINM/khOx4ae4vF
+91qwYKO6fcekIQkioiZQxQbdNLoVd5ybEMRUgjkG9oA7zN0gWVXFBaJQxbIavGfOyVa1pTv1Z0q
BPoOjTIL/HTjlpXoAURCJEqzQV8gLjYTblgF6NwaMXdvHnY8UsM9vDEkw3YgHeFiIoxUEphJEXox
Owjihhwd7P3ZJPZWULnoBAz9DR7jNVLQJQFiKM1twCm2IP7tfsjwnlrIMBDZIT8386lWogYtYZIY
y3/GX2wpV2j8r4bthYyphL/5/LHPMMm/pkgU3uKUbElv/hCpiBZfKw5InIgC3NqcaBcKPam81eps
aeQX0CS+wtRcnCa1o8mvesI73BwkMDObLdF2ex0Y9AU3NBz98yPqUceQ//Y5PBFJJFO13Oq0r4Lc
hvZMm6XB5t0kRAVUN+dcFogpC1swkYBMsJZa2uPfHTpYmz7IK2iSw9iMntBY1XIZKxy5MiTuBAoD
JBQ72CJM5EGZi/oxnPIBGBVz2WOp5QdhRKdX/pmcJmnqTAOyzh+bf4XG4Ya4U+IjzzQZ3pyhJiBK
9KIEKnpHSedpH4zDJ4dkBfYtX2GAh3E1QPfRcyCIIAkkfUcFQm/vJyPxQ9RpaUFVhxHJFytYGDsv
J7Dh8jxoOLZdou/qSIwzQ29uoqRVl6+0j1O2wRTo7bLhgUB9Yw6rDrGGoe/z6WePXky243hiRuMw
RtwSGxwzn14zR54HIObH4IU8QAtj3piMF/Fskq0MyLVyeTzjXwj4IACPsfq10st/irFqlUTtYCL3
SV72Fv89N4No3MZzT+h8Mb/Nz/8r8BmtFWGjqZ4TQZ96krXiotSxUgjpZha3OCubWo1xnn/876oi
M/pQ08JamezQ2EBCOfwrWckyuS/d6h3yY31OW7ZEpU5ldClLJ6m4AVzJAHwtLlPvSpDT2Tv/Up2R
AEPJjQwiOEKh1oWHPZhXxnruWtS7dvg6zH0++ZPf1bunPocBSjHxmKo5kMrUhRKTDkVEhGlpeG3j
m1wYOG7mCAdtT6d8KkMW1Z5ai4YW1makGrzwihRfU/6rdLByCVlBz2i0eUFrKGYCd4xdZ6yYm6aQ
kdGFLVuaa13DiBtDYIGl2PhJaAJbcmmSKlBwB7iCLnSqLQxuMvC839S1/ektXs1qWz0uLv1SQIKI
tyIi7XF+CpMOZ4qSBT6EdDl8DIB4tMqi6xQjjAVzEvHezSz9B8CpSOW8D4b3IWvvyy+VyXsLKubP
wrXEr6+B44MOgOzpjPm2wG+Jo9LZpH3Onk4zHvB+ROeTRBTTfGAYHOBqYLemOvTGfn7zBB4FwSCO
Vge1kJAktyct2lOwab4vFjb3oaLWJ38GdgdnFqNNtz4macyjTjTavKpiCPaB35JhGeErVEfE/0tN
35+zZ5Y3e7dMP1M3rtuqHDnAmeF3wYS+rqa+sv1+o4zRkxFEpe39w7zfQ0xcIlVePZla6DmgCWOJ
pROC2AinFanITP7tKiRmzJBsvpzayzvRL2igIpa0sefGpcpILM3nJQ3yI7OzLywcxq654LeiydDC
PzVGA5w2kyBV9zexEnFPikTqz8KVLAeOjdXp59lD8E0bnENBXayE/J395XqAU3KAwpsmkka3L8kx
3dSIVg8FJQiL0voc5MWwBB/nGFQqi0wdgqXC9ZAolWf4KhyggJ5ZgFiUvwoS1/Zwpp+qNzvthXtK
5VcO5K9N0zdl6Yp+FlJMAU/IZBi1REmLy8JrtLNNqrWy/h2/KIUToNz/2CpBcbHEEbqAFQtSbNaO
/FwBSRMTfvI8TbfoXTdvRj3vqTIyQmRySGvtwnXeMYWlZIV6sgaK0ETYvfXzwkrc6WtPVakCWw81
WsuXaVB3IVz4ix1o18GCCu9uY+3DhdR4AV9MAj7MqEKRd9Al7AftA/wxTRt92kOaf1LomysD8BmC
M0rBtM+2moGrTNEnEB4NTbTKVxonNnqrHbF2pdRZfwvENgRjEf2EuDfyJIagEhE4T5gE4QAoCrVy
WrsB8fmwyIjneIHUgp9ogwN+FVjonyxEb/1KkcpH27wItxM01y/VgR8k2ARuA9mv3H1Apcr4GyKs
HeOTKywaTHnjhRx3vXGBCdZNVSSe0VoewSD6OAOABE1z6ffA8m7e88KW4x7aQNEbW8VtmGfskZgr
BcmqE2y/zPhqxvi7mHWu7eO2C1/ZwR2ISgHiG6nTvJY/RQZtM9b6l13/oeF2yc8yFVaAOEcR2pAe
2vPBMWBhTlXj3fvPB6m5oTfGgvmubkoTUBYn4wzhypxNXIZoJ+a+hDtFNDHthsmxruFNRqRqmI99
76WObnfZtIF0AvIy87ZVanR6+tVT57bj5jXGd0LS/eje9IBHF3QuRC3rkCuZBOE8NN5Si14RQVpU
XK3hhjpPGtto+4eEj6GCs/t5YAtMbVHqLZQL6SDKpd/DC+kU5V3Uqlf8zeE9rApzknxRz4kU/wh7
XV8ZM1YdbTvpgB1YKi4Ju0hq93xtc4zq0Qb4OrXAWJTxQZcCFmFoSuiSUit0C0hwd3PTcVLIzip1
o+4H9lp9Yn4rvzaUJ598B8YxAYVya9RVSQ/2YxBrn7LuQG2FSktt/PcBEIyXqMStNZvOWZ6v8dvf
5R6BYYjIfi3PJRZZYZmOnxzTQd9fL0lUNJsLXPJ9NwW6zEfsdLvFMq3OlAIz0Yjui2gfO9Chlb/i
ImcVk2A2VvW3QI27ii2tBjR9NXSdQI974Wua08Sb9ffS3tFGNvLVqi0AOeyBlM4ljjZCoxDHdLMJ
TkdODfYeFUGDPuwXBK7rLyCvzBfBCCRB076adtg1Cu17P57BcKkaVsi1oS7l9+h3B4J/9TUJ/kXg
A28AYFyLIrHsSuDRg+BNtUotpvaQ+fq2uVH9PZrW2gPHpcwsGw8b2m6H0RMPaYPJOas42EF+ZNT9
tJCwdm2CgtZS8dtFKdOgw47SSdzlcQtxzgvbfp9bG/Cr7NGUSrdy2CBC94xXNGBoUlHK7DPLqZiV
H8KsPf61lofG/dmmpgaLzPbkzSAdGFShi7t/Z51lLOoot/UUWVH1VggzLzF2S0V/oMZS+RaOQIh2
24sc2ygnKX2yT7p19R8l4fqgCL2AXMhq1CkjfNQ8UnLuZrXvqXkjGXaS5TH6O0AIGh/XzMhKfKym
4LXCKGIzCdLMj1PN48VW76CZKjygOsGnqwxtIXMmzQ2ghXPLrUgZOGb70lA+Aj2ynxnnq0Kve1bg
gJeJuPu062IIua1aCbtJzDiM8xW0IRdgMKmBvhFsi5N/ipRjLpDvG/dwiZQv+nEWf1F9wATQBeGb
GYrFEVrQFHg8FwnsnN/kPqR54LYrsEMK1EDSkiEEKT2dA9RaRzkYgY/h+eL2f4dek8DkkKJz7gVI
kDWHjp73GsAnzrhblXWN2v2WSLwj7pnxGc0BO1OTDjrpq4OMAhmhlil1OQ32R/aSwHB6vcdnuJM9
0sGppNumzUV3dKWLg0whPvdnQK6IPxEDZpxaOtmn/DT9n83rgUczOrdVheXUq6FXwLGt2HL8AJLt
oKzAn1hn5zXLIh7Ppn66i6NVf67CzRcmS47u4/Ha0TEsNqq0IVEpFnYyHV3jXureITSFwxTsypvO
av5o7pDqKABQUXFqggTZScsOgTemupY4Jfk/Ap/nje99b9tQ8OIx9aiuVFunowrsOnBS0ZwkSLKg
NdTvNeuh6hufrSD0MbcLw9VQp/E9KlKUG924aYg96Z5OkVCMmWIuQzq7umiUAyHDk0NqcG8AsVr/
UczhBbQkMiR69IWXwJ2XtymJ4UHz6u1cI3Z3lLem1nYK8zJRe2ErR+9Cxs4ckMQTsn6Rla3CfLOs
81pUPlTMJfII88oBNTqhyg3SFD4Ee5TWjVWGjRh7qe8N4r2B6pnf9gX82/GpkVhwyd4u+CGK9E1K
2o0EwYMb/GXVquMZ9mC4PguI/ZrTQdJrcwSOuJIViGFJnvKEtJv8v46V0BhPSu8LEPkwGBcPxi5Z
716dl+Ns8Hh3eXy0PQhhKRBdWPfx/rVXGOLoWnjXT/cQzTE6xL/pfATvOZTC2+UxEMxRWlcYzsgn
BNoplXiNiBV1KB0t+G5wReOKLaIQqQzSqqjFF7OCFRlsxo8C8vU7+vu4O+yKqC8Lmz1PghI8c5Im
7Zdp3FQIRAEsw72EGSZU8OkI0h8DSmL5pmlLiTke0dmjax33NxyBC+s7nwfuf0M6e1eyeMfizsv3
6hfxF7ZieGrmKwKH2ssbW0oUuq3K1d68gwMzDGGdj8xJZed+wkKIWG1Ek71BZglIkIZfoCvY/FSx
jGTZG5uM4Pc2IBjRh17+G3rGyx8DB5/p8BwaMmWWVuUSDFMSnYhr9vWMYUcPRtgpWBfYVDiO1PDW
ktXPHEroJwiJYQ2VlJFKceXf5Y1iIH2LJ4rhiylOp16dK/Jdv/mhDGIKOiajfTJqySZZa9OD9Aff
rx3zLbHqkvdNvVegYfOX+0MucrmEGnmNjT63rx/ndJAuSToakO+kzibxB5H6HcMhIQVGgqmxzBGl
+FgukgnPvpQCa6yrmKoE5F2q5DFpDK/pGELXoH2lhiR/poaY0WzoST+UmlTOmTrjJpsC0/pW79i7
BH8i5Eg9Y2r5wqeT6Js8gxkyjynvo3y+lxGJa4TTfdtLxw9B7mUQe8eoiRIX5pR560KvJCZQmmTE
1XhKlaSH6wjfvQSo9wgYhJYNbxlpnpVPdeNLMyaxl4OlKCtj+nL+NH3t7GORRLW5xt9fYal7zc5Q
+6xofukN24YiTYusrkx3EkyRDOPSp05mdd1oMou/TvlRBPkf+ukNKGAY2fIC7RkiubZImsonVufM
nOnSvcddHaiAtgVLvxHmhZ4foDq15AoA1Lc1rI5LCg/XZaYIStqDLkTuEdS4G7v+tQVaogVJ8qgH
nMSSqNZmaMhPpRTdD1w7riJPu3v4Sc8gmDC4x+riRLgf3bBwmGOUTNHblZpJ0pSF/ZJ4Uj6symNf
rw/IoDoRrIkD9zk7oFk8nVWZXrWWZfhiZuYGuhPhObhfjyq03K1ug7zCEeUlpxSWmBw0ZqJTNBgU
XwVtyrMeGiXt9UGz1aMCDBJX+5E2JW/UzH7bTAnm2o00a1QRuT3k+tL+MlL0AVkNPmbOEHPKWpJo
+RvfcFWG9+k+xS7AqAXAi9pZJUpMXmfu7f6OqXM0YDDGXcIDIbe0LF4LrKfSekPunmV4uzfwpfR2
Z+QYiSlnWjbHRZ+B0lrFGKgK89iKL2E0400Ww0/hjox6JwGRS9Bd+kzBdx0GMN+itONYsOceopAB
ZRTnZX9pOCnI4md5nXPsteO2lgfhPL2JuhS/5rlq68/lyr3rDeTbuSEBLfJ2LMuf9LVUYih6PPuX
8dl8VD1NinMaT2nfXHR9todX8Sx9xRM36ymB71ocfDAQCHLhvl0oM75j6y4SKD1PPlf3qzFZfueq
uie9nte0YuXuAALCORVWJLJNZMq28C4GDA2k2NwEeECnQ9kjaN/5/EQPj3WHkwAcguJpiePgGgXI
g9/4W4/kD0EObla7g7+v4nM5yLqDx3HH3XkYFcqJiaMDrao8A7prjzy8A1AGtBnME+G0ew6NSo47
LRo+Kz9GVK44pwUB9XalorrlPLd80Mt6ejTu0zcLutHgkVgBYNzAWfV1WVqfDHhXHxgMHSn0Je/K
/sRd+WXaqD0ojOpXrzt7a5+pFuKWxZ0BGqOcS02iuqAQWJaFJ7yP1PG8MGn7iAuri+zsTGTNJMV6
JDzTyKSJsngAvJuhctWR5WgrJ4RBDQwUKLEqxizJxszMmlXge28S6FL3FoM6EL2nF7GNMqnbXRv2
shUs0xDoV/lIxBq5IlYCLviylwwdQM2oi9ciK370U3ZP1blusUUey52ThJQgGMJnyn8zcYuLFZnw
FLWbKDWfBLb36zuScm+NtH8Lz1uPsGn3OOMbksFEUSqD7tuFDF8GSh0t4jQdQoyv9l6lcM8SSo+b
ixVJBfhlVhWvx6dnn8de/kUM5wSZahK1xsPjPK4UUBc9SUlUenuRnw2xpRbzdSY/9RTiKCqoBpqg
kXp/ulWkF+tNN37P9YTDJZ0Bp3Ls8g5eNgkHmc+Asxgv1hhjfUCKT13xbNhMBEUJSjgZdaXyyUNx
3AFftJl9TK/lM/WgHB4UmKFt55e9EqSD/MKF0k310lfxiIFDX+NcO5Jb2ynvmkYKALKu+ZJdAqCe
fzoPWLXjXaWhq2JXD4ZhoGlYY0fXghIxKDu4o50lUF0WOCNDcLR/y4pVP7NMfjEEnGCaM1f4xFau
8tSkcJ8NIXVDBAuW1zOuF0pAIRvRD4ISXODthNHBBmMO87w7is+724Ye/GClBLgxHjnW/KhnWvRe
VFxhE/ioI7pTdA22h5ccIEy6nxLs5XCmH84OcTidgY0qQYTsjIPOL2isc6yDEW6J/QLDUqBg7Ak9
hZ+z1bw3XePPAwKUpfDZNxACffZsKHX/6G7rFAdpQ/0KsYTvP7lTxco96Tqjc5hobf7zimpp17A8
FGoCN+KvAYcaVPADTfBdcPV4sWvWxp/ET9+4k+Tn45Eo1geXknk92pzDwLsF7bI4oM4RcmX7FjK6
BsQZYtofNXUO46VaRc33Ed66jQSj5RQFBx8GS+EmRxLibGvW015XLmzYOKgHuih59fw+J5uc0ma7
DSPlIkVD+RMsdCO572Ug7YdCO+DUKdZggWpKxwUn7ttoa3qDhjJi/FpvMIXdSusL+Vn5bws7Z/wg
2gsDHAaiLQOXwt7gioFaqWkA9DM7SqAoeY8BQbhA8zJT8E80pD49e4nnYPBwGGtLuUZ5U2ws7hBz
I4/J6l6Nca/RAq/vvF+c7XbXDMvp3B3xUE1zGVAZXDIoOx+QPb6jaqy5T1g3LoYfinOtjixa03tF
N72sYfUU6DlZBWXtr2g46TnqF/HhVKYLHa3dFDT6MndhZLExKiSl6QVRgYnS/YktrC8hECU2znwS
rjI/SCfxqVmBWJJfpeOgXc2SHgXL8l/ic+bOZFZ/bU1XvXBbIG+0XpQstrdi2U+ZBQBqLvFqsjBZ
j/TyyFrNMclXx702CkpwIBv2jm/7Y/KxHz8yqJ2D6Aj1lLuAfxvEauh9i+zeHqpSW3Vj/HFRDDsI
9OdRg2dLU5fBs96HIiHnN5mB6NmUJBtA0rOVFEAbauYBgMicpRA7HDqZWKqBgwzx8LiQaPM7lAEP
Eo0cm7tjpRYFJu+HgJfL2zSSR7dKCUuOQk2XvVi9tZrXnc6sw45TopU2Ljko/vLu7drT+cLPbyfD
xAO3mZPmDrwSpmoiZGT6fbm2eqSMwuMqM3qC0HP1IKOk9dQqB/KgGc8mhRaAB1biAmzZYCziqfum
2Jyam2X/XnCLdKA3qxmN7SUp0ff1zr0Imc5xPpwQq792YQz72fz2VSMqYTfVa9Fiaan4urFdx5rK
L2QoVYKu8IbbnwHTvIaXtTzrUdrd1BeCeut+QL52+1EqM5GXx+Zi4UaQ/bU9E5ZpOFcn+9X6ThU4
xRw3ieZWUCjw74COCBF0iBiKo8a9KUpzaVaXBzuyKN2s+wodWw8zllojtJ4R4AIdvV4r+2jP9OvT
wFXAMXqD8oUyoFeNHV40AgRgpARJoGoZMqsJv0up8yHQeZV5MN/5KxqUtvDzQdk985gABvTY1Xp5
ULhkvX2ktQy8lwROp7lPXVuZjTM2CT1Wstw2BEGj0SoC30KrEa7oGCM2Qy7RY9JPYkwmoVPARRvV
BKm9KkrdLNHTaGci0Q4lDpUm29w4pPNXXLeMnoC225hmr7nMIAHuUISzRhItusTdrn1Ms1fb7fKy
U+b4p0fbCDVh2gonYrZNB68iF8rtxuL+WMX7rTY69lF0DFa3UxlaCXkKNtp6tiR1hRQ1g3hFaw/8
KdXOTXZ5JXurKMLKk7S4xZvy8TKiq0AYRsnEpPUCU1yfKgf71dBpf9J+6Gp+IdLzb10rakwcl51E
YTFziDC+uO/PxZchJNjBEZJq7F9plQkUTjcy7cjMBKzRbHYfgU4gKv1IZH9fbTJrzy+YNdK70Kgh
M7trLxLuk1Wm+7OoiC3aQ5kbySptJ5KIxmYur2jgDgwLjsQluPAVnhBXs1H5+hA6b+C4xvwLUGA4
hLv2wUCCjD2/K3z6h6TrTa6pwxoRlEvaKhskznPwrDTFX6BAJK9V0N6YnQ1LdbDZeq5y9tynU8iE
7xRILuxaskn/tj/p1jHSpcy4WSnpG0Yx7oNrnklZxx5Lw4d3M2fPRBqiaRvtTlyCzHGfIqtvZ4bO
4js9jGrbPXqlZnEwsOoOAE3VZvvYj3TqDzxoyVwRpJffMxnydMnzj+WXmnkkIo8jHjWe8HvRtxg6
5gZk/26Vn08v9n8FjcBJfoLjZE9nzsgLtnw5Wn/Co0nCNf1C1CCPAhcSUE4zsDwup3KRsZVU8PHM
wAdU1irA0wrT3kBsz3XhD4wFoBGXvNXlTtECDaI+sVDumptemHyEAbVVrzJ9v/PjXrUGMD3GTZi5
R92B8Ywjy71rfhJn8D7mIlBBktLvSDA9v6G4oLZg+XnxX9lRh16N7isE+8pnU41J49WMtEeOrSo3
Dk4FJAi7lx+p6sRBWCqpVl1mVn7JtaEUWoXC6vCdii1X/wsSZmPbFpxqKRbtnG5hlzKsFY1eYfeK
VGtiKz96owkgsWsXxXsfG6n+RRsvqdokQq8QrAWU3R3FWU1b6JjsvI6mOg6IYST4+bGPGOSETiul
I5t3IDmD6EW/xriXh14SzYSGmBcwVyck1g/0KTabBElfP6u+LLHAqD2GR7S1kl+buYOyjKlvITj+
GcP+luegOk+PuMXeqjjUAQj0Ffwjv4qlPuWDxv5jHZ8TpCYpQrmtUzCnozL/TY1nWwDG29g590XL
UoCRfmMfZwX4eZgY3RLfV/0ME+PTcrCFNM5pkZjWmQwrn8dYSnhxrqC08gdu0Ip/JvnDyRGNeow4
YUxjrodv5RoKDdfG/xzohR88BesCRXhalYhQcTgv41n70PrDDdg2OPD8mObG9AnCM+Rr1j226x92
87Jl2lenT6qxfkD8JhhKv26EW283pn64P26Q753zyTo90djdo5AdpfClgf65hdbabc4htU3lT7AJ
DW/9S3SFUoTaXIOCkIuQMvXSJGcuXffd9HhNPL15dAX0f0tww6gcuMM8dzso0cGtvQxKW8faZQBt
Q9IdKFS4WK9kNASxDiwZdVvM40a85ANQSeJ7uYHhAgpOdZzMYsF4QyvWVvBxJS+jIAoZRrCT8IL3
4VitqS0ANb81iz1F7JVmp5/VCGET2IWErMZIRvEnJu/Mbxv3OsErgQ5IFCGCJFkhWNjGDqnkAbr0
L/fqzcM7J+bUgBxPrlOSOX5LMJu8Mf3sCK3V3sCakloIA1shWxE05FyUzDVe9Jo+BBfFnTHQ7z4b
s/tmK6g6A4MvIH6WBOmrUJZjTH+1hbp8neoeDnMbYeIq3W7eSNls4TGJTfBbyr3wM4uduRXP3ZrB
qZSyM6xMFb9jYiHMtOaoaCWx3VEQCLiHJVxdvJF+HEgXto/2VPN1Vn+exakf3UXmtGFpVXU+3R/K
tnfJEt9Mxu4eJVAdpMpcqtF6ddHtVX2w2kul4eIAE2u1T6sFyHMG42DJqqqEMX8sCj8cb1PYmDda
fFxDJpzQWoQGbrGj7TtPJ4Y6HdAXXTWX1eJTyBY6dkU5gbFWan1M/TgkOcgY59w8woqIi+WHyCbC
qQTlqGSGmSGSmnrb1EcNhx69gsHBMlfv0qJ5ml14K7U0ODVtAVSBdrg3c0L11QgdHcAQ5CA3+b1o
BHVXsO9fOOHLNgzutP0ZOFVvO6Nx9fwpp9dkYoOGHgczUCGKcZW2/VtqFvcRQ6RtRwlt/i9eUiVa
4soFVvEAX6fBvByKnCewvW87yeeYOgCNRSE2y4ZRO5cmdZrOAmg0+ZnpkxdAzGQ+qErcmrlb/JtM
8XSAGvbCvxWCUNHRifn9XlsQK6m3qBlJVFglL3Qk6CBQeCFZm4aVVt0EsKUf5M8dcZyfz7256YuU
UKpX1GYlv3VHpWmR2nvIyPK/uZ3AvduKfswbtFwSaMTLBNwU2rPaP2ZXSiljZWVEd6Q1P5q9TisD
wsuqBEBsmwOQkHCPFWCd3BSxL+ogAN5F5JNg0qWKjqRrDeqcxBVlFeCHrLqc0T/hjWCOc1yH4dax
xIcgWykPng0giJiopAUXc3fLmAR1gD2UFSF0oOi+SRSGXVSoef52kzPwwGEnFYtL9YjNjI1KhXd6
XJddvYZis1Tlp3lwfz+LK6ZgwuHk33pOVztecLrYPz35MYoZWgen0lq+8ag9VP1IMMhIjn169Dx1
sFyl1CSS2xdNntr9eEEKZqbidbINrj5YsH7P1MDcftEGmSSqzJgOQH99Swr6OFtK7UIGvdY1uaKg
RwIqR8oFy9oVYoYL3olaG3G4kVmgt/CZb3PGj6JcIsmV2x47q1LIncy2NCWLIlNGhL6j8jlomaRz
9hZKTHgwu0njwjtP/FcbMJxxhA2QF1Bo4yJp6CmXR2xcJD7iLswYHj7VXKx/ZxCnKHQYLiPp7eiv
Ye6LnJwyA0eNdelfC0wti+K2jAvi69tD15g1PeQgwoNk9GDf0vr9uu5oM76rZZKFECV/TF5cQ+hP
d8zhFGGnU8cWvbYI19QyJuNrrErivyBvt89zGnmO3YCO35mAhHWZ0B6x/QuzduZzJTdGv0mXcFxK
J1pjL+s7tEdmmHwMpZj/CzRaJhWhC3EmQvTGpy5AmyaGozl8wohVeFil0joQtOtbx8fLsNWXbb3C
PwyqCEj0836yNKwP+gHertX+9n8DS3szcFK7DUwHdQfcIUjdZRa6Xl+463GTxNYE6yjrVaBxE6f1
j8SDc7nubJqy+dJRIjuTWNEjYWs/UaYUYC5jcfCuI1NvG22LS+mcOCaEkNxWQdHwXBwa0dp8N10W
p9UkxQL8pImJSb0uONDiYVbAHBDK3SPDKIHfk+FK2AcUJ/qaUCvETsrJWyPQ74Cm8c5lVVxsPdiT
V4VEQE1J8w7CDjo501yQBuE/1+xnTp2lxAf2MvCfGd++RwuGkB/NLf+8uaIagCw8+DpRotejVGZo
dMF+feHqmCQ+f327r7LN9N2Lm6Qe9UJSmJn8xbD0TjqIrZ3sbpAtwMfhenSnTXGAnF0IDOCx7YS5
oj2hUvGfg+JGr/fUwGVBUcwjoH1RUuyijqLcjwhpTA57psPj2vQzJPGQn5PxlVMYw+JB0pnlGHfE
jo5lyaoIRKvnz/vtVJ/TuG2p2e3tjB6oXcS8Ge1ObfO2TQNzaVYRVVHIzCVqefEidk2dd3xcW4y7
94D9Qyl+8fqp8Pfa7rIrvF1QPmkpzg4Yv6suVHehcNDIkzytvm8W3y3Rbj2DPCa3zJ0fwAKPKcS4
hUf1bBoBFkfTdQJnl++VtFntfj5LyfPOfUWGkSLnb/+LAbsvCAfQ2z7E/j0lQyW9TSWyyw5ylb3W
KlrzWeWbdHkWVwg0GMPNi/98Zi3nlkDFn5Y2LmpMAHONBlW67Mr232qDOz7QPob5vXsg4tLPEiiO
4LOdlmZCPlgwOcUCZjVcMQPH0a3C27opzyZ79HkR1TCEHsQSWPQg32ercPvL1AecEgjwXn/WSgYT
buUUa6zi1T6cdKZ5f/zGsaVI4lSBQy+rR3fAT+PSK69to7Y6yQ7+YTISDVeoDOH0CD18o1sLp7aP
XkrKcyl+1nEyKIwkfuTeBGsmfPZhUsBTiy+E+cTMzIH7x6g6MfkqV1OpeMcJDKfNN7MlHBZXLcG9
U77JhC3S/S7H/JuyO7blkj4OYb6flc1MxfXXS3rFHjacDanWdzh1s4sIplqyAEzZO8bH4FzxIGgU
GUgQm0/eL7/iXhbP9fiQhZuhFALwOCwkE4WxrSDg9LLCX/bALWb//v3xfIviRs9uwL+A4Albvz8P
HfO01KTomLPtZUQCbHcXVHcFjkM0SkOw1LPLNbII24o06moVdjuEW4pqnvb5Sh2Cqk2R47C6O66x
Cu9FB6/lK4EBGLCmlbKkyAo0a7DLPB+POpsJg8o3SIGV/xYMz5N/Wd8MOK9oEV3Qxd/ioHzvyd12
RSWFmC9bEqT7ZUcTsbcCzuPRcWvLU3Pcu/ZH72pPtp0g1DhyO09D+W0rQycGF6zUrZRSgaK8dJkv
PW7OGa9Qf3makzmVHnsZ1rr95WatBMkj+SoWXSSIJkQTZPfAvJkUtv31TmnIvW8MOv8iUwxUWXVH
a5GIQFkEoMxW7KULyKWBRLw5Vjbb5T5TA07syowoEXdckEcr8HahuKLi3VgYZAvxTs+nMZBJIl96
52dn+hLUK6Xa3d1WlGJMqbf8+cKBxApjpARjuO2iDLM+j0iiU7+nM4hs7qKjLk9ZQiIvxfDAh72A
0uE33YKsPOzaOkXOOjh4+RKqmUghlE0i51tuLfFoFsB71qw/gmKFKe5/rEyWWl0DO71NQVAQ6axL
pdCRVPugOjVnPVRVkBuKUiZm/4JhtpX4Wgx3XtgRSeyZeZl0HjTP9GpLBdN2SBtoAe35e86ybzLM
Hd+dspKqXqa72D1ktdFWnJu76SxvnDEIdWcMUt/J7PAVncGmm8Kc/eYPqCM6qzmGvNEW611aYNrk
D4bZe8hfrdd02XEElsiT++nMw12c/1wfOuMf5Y9QkUwIk/x9A3FJ7B6e4TvADM6YJZBLQurdKlx+
PLFq4lem2Ag8YoT6Itcqk9vWjJN0ht15ij/26eTfBhz3jNGhZQT1oQstMYxoGmdjmHXm8EconMXe
rWWJr6dVvYWDYD1985NLP2z/pFiNY4zUkuM5HV+YLToL77ZCjkHw3VfxMEGgPyLUzrCRqAEgQrrx
wxB4OV2vZ3SNfRCzL3g1oDFtAXsnRhGMrQP+ywj+YcQOfbViBCTtDxjitE/fgiV20RQiTbleWE77
Pip6tsNdT/BTSLkbOG3Qgvv8tzlafc1Yx25P8fASyTknzdRPlFKoTkeycOBuWvGV/Zc1dydH7how
v6J1ZLDPfxcnvL8uFEPUpWoaNxYqYEbOEpHv1hQJolXlJHwY/OBm7hpmGqezq5Ku/iRZbGdJN3NT
SaGh9p+fcjoT/eK/swxkwIcztd2rHNNySc99q372CmdopZxFSKM3dCCgcTWEHdDO3tdQtwgCSp71
m44JH/r40GKR2WSPN2U125mo1Ftdi9SBdAEtCHC3/5i9QhvdQ7PG68T5gPvfKYD7V6rL1LGzruj/
qu6Mo3NeU9p2W5oW/bei8yi6ZwMeCfpDGIaSbB3gOc7HIGWcrRFilE7pnQbhfSCsysSHyHp6GsA8
8QkYt27iMd9jotVJxzPajAjvDIUPmMF+iiwGXn9x9Bwo10zAPdYJgqxBR+2LJalu21/JycAcGH5u
yMwVrsov9Vn9dZJzgBjlPtapWIu+hRfYhq1qjp91meuSQdQdyre+7v1fqJeB4TWBT3yy/uJpKybT
O8LrE23hGguUjRyok5lFov7/nSy7sx3zKVFpYzZ3Nu8HMu93xE8FBszmyM2aSN7HfTD9IePgxCyN
iufwl0npQ5Lrk3I4TrJi5ENaGyQxt3iwfpbw56TXRIvInZ3+RaHggpX5xTS2Al9hvscDRQNoAlcA
HVjaVG01jMc1uf0dOhlAMoA5zzcot5r8bhFZZvNuh6T8aQNSOelPOnbus/mAFVDzC+6XPfmezHgy
3kHHdfTvczC/YB1kwxB//LVBAlAsi1yq1cv1+NyRvrdJJi1iR77ZOXsXyOiCVsb52RPMGRVEiMXi
nNMA93iuGMwegdxAemknUsBowE9CMWwoIehkK8wluqQrxHSZlZn9QgjkO7eLXi41v4E+1UjgA0vG
Skg4ACx13ZA+ykVLjiVQwuoVMiwnlluemb2AoCUG8pUaOEiomIs0lXaTkQ/+949iBXVpfwCILwva
73BoW4/3IFXj7XD6o/lyx8ALzYJ5K00XJ1DMEQUpD8dtyyhA5BXkiUro+hD85tRKYusoYNayRnb0
VqZQBzn0vjmaZdniyLjQzp/jnU0qBbnUDoSNaAzz5RB97CGdIrLU/yQVcKn8DT5ic2D2O0I/xIQE
eINfWNXwJ7/0bwq4OYFJXLrqgL4Ir0EseCS/GC0olWV8fh0FxG08UJeLgTJgyDPDFc2LOlHvF5x2
VRRCQOi7omsRmrCAhQWksuRGSKKKsa0QV+MKVWLPmqG3TxNTkjhg9TUd9nGVjUPbBmeqXC8SroVU
zCxiZZWPhfKykPmaSBP0b8EAfit2aaq7viOCFVoW967ZN+qi9xwAj/X1hnmsTdpGiR4rpzkPBrWc
JjetMvDuftgiQ3uYuWp4NFn1kg1mv+nIumjuORfObe/e4ZZPMviDyLtsbEDllYfeM7xnVOaq8W3+
MJ/FuBaigwzpYQEC/Vg19/FFbfrUGWIhMnyPy3ePmpaIn12T5u4zRGbFQnPXpKstHE6N+Yk+hH7Y
K8mmXqFkez0jwCMSpDhBA6YI3GJ2yB5dw/P/dTiKEx3D3lTze0K5MLOHwoi131E8mB5tbrXse4cW
iljjg9JgZqc1PotsNMEBwHFF9Hu0/ZpBcE/gEwo5TsDN9j5upZEQlAazdCCajLREVYSWbaLQmKhf
o7FiENg/lbVa7iFfilR4dAshouy7eJjxewY/VwJZx+ZSCofKQCRPiVq3828/Hn3I1T9S9CmRN9vg
PgBKQknkA+J2n8+mxFE227xMO8M+/kdSE7AVyxUmGvUzsYO32NV73DUMvqlr3kj3rK+TP+iRnF3K
oPVIygHVkgvj5kkf7Ee9y6gTly83lH2SMltokg148M/yecEqIybgHVzTBHN0V/QJbRxdLUBAcxcz
rLpPDmMzLhHglHJmebarlyogrJxH/PEBpgMAeIgzbhoe/eVOiz2mR/pglNbB+Dky+jof6PpTHYyO
R/6A8ebBAHoVlgvgVLxj4Zht0QiVJCwexQs5y/tg4V91yOQsXdBbKFrDRzwzd7WMP8gLqoweAE+3
Eo+3tpCFJqP0cFTAvXeZfNTFL3AEpmt9eDd9EPZHlHOr3jP0mor2GWHX71+O7nH6REWskC2EgV/N
71CQ4zfN4wm1+8WezTXQ5sSsHhjVySZqD+aBWEWSDNdDmCusGlzC7KgRdhESBNzrEjX6JqJ1pTP8
5BEFZi3bhpXmTF67eiYykpeah5ogSOnnX/TcTplebjUuejHgBUbwqRCTkvAdpDjuYzVNXWqUWmaw
juFPwBfgXvWc32xuypTqVzO9HUcRlXTfesWO8VYiU0HuRC+TikYxY3ghvHRAJhcGaSqvI4T596Gw
f8RKciwOf/mpMqjjl2g7TRhuVwdS32Bz+zZVsohj1kqSdbIelkbPYrvuo78COsA8OErF3xLlHP/5
u4k8Ws3nY5pigIy5KjTlERWKe3nVUWd8bzL31VOBTTJJMsjWbIsF2zLEy/BbDeKRbVYrKiwLjYsi
R3tKosgqdO2wO9C8gm418WtJuLVMpnABROkF9abvQ5hNRTYyiKYkh/95JUrYup3xDe0jWGHPub0k
3BNuBGLRGBNWkZvZHt0jh3naCcLCenRYr93RhcUdVaTwuyqpqZ/PpSWSOloRmGZkAfZTR5JXvm8G
2JbEwDejnluxmw4XoGsxnkQwgMEvPXlUTyeqpzsZDIqzogeeQnCoHte5g2QIZs2slzIPFjBqkx9c
lO/Z5h/enXzDvsIXjQpQ/TumzVGb/0Np7QYfmHz8i/gPPDhJmYR4jak264b1LwnbTxPNTiMSwz/P
W5QO+kvCSgtPgg+KsMDQ/iJqbdSQGC2+5/4FqpQPthoL4Igp3bXkkypE7vBJ5nd/e/fwohQ3b1D2
wSHg5Ob0ALgOYmdtcZi7Ntry31eYQ5vqe5PMLO8WAB/ipfmGTaE9TSaNpDEuXBv3fgzJA3l/jdVo
pOivqgN8bErhVgPAgZofnqqcY/k/VRri77UrTOi5hJxN/+T2D5ZndJCN/MI8iEDX9eGX/UU8eTjv
6IBvwcJJ2c3QvVZQE2K+OnpqAGKAfyVhmUUhGLdJR427yX7Sx4Krc8EnggwuxV7MKcHKd8DPbhE9
ZX2kNag+wqCF5RwdM/F4v9zY8CE4vhR4zXCFUx6YlYvdSbOgWP++QJpAfWEci2zqPAC/O4wu1N5t
mo2d1q6aPbmYP4FOh7aRhvNdq/ZGNyor8E9jzJscJpv8c6ydr/C4TlB35+z9UZXZbyevFQA0geBc
nKGeeP+dzIBzjM8bGw6DWFd3w8Qfaq0qmYOsfPr4RiGCmSqnNHYA54wNfaVAuKk4oEHyNn4SvcUP
Q7CH4OqKxf+rD24K0hhCW3oIk6mywuK+Y5ZNew/rD1J7NmNw/T0B+RPZfQrstwHEoghEkAZKfEOF
5+xQsugmpnJPly70EH31KSd0x5VV77sOebSKzoaJZYHyfYq1P/UGS7tQuzp8pQ8vZv7OALqWJbUW
48WXr4RaQytBHvP5RivEva4DGITO1kM3PzsEaC23kzjCDLvbMXXRdjsly513xFX/7jCGJIAMbXW4
PhpgzO+bFPa1YDGqtxi8X7wqTNIRp9V5Vv8dvaV8UKiVatElg96aT7KUGoxJZcgVct1bQalLMzLO
koDrdWMIYGT0xt/fuuce8rMVpJg8h0vI6uMp+OkA4glykJEPBqxt6h0/h8sbRnWKfSYeaZfp9FT3
U27gH9HDY0C2qPj6+C0QjbGWMMIms/U2HCxUig1obiBq8ecT0qVS5uBr1/XEzN5FenV7DyFB86Uc
3FwRYYGWmQmGTlaV+aOSk3wDkQSW0W/qcnQYyvlQmraO1jl6gHWONe2RTVplm3r9eNWSacqazUuR
VwD8JHSzFR+CO7HFG6DPaIobUQUCM211u+o7o5DM/x3JEtKDYHkb1eyyqDGR0yU4iWqaY4fGBSO3
d03Do0sVavW/7BjXPB8CtId+NgAsSJMKtuXe+VmFySolFHr3Wv0UWXipE+JsgNarFdLCv5TusIDA
9V2BKl6SQvp7l3RSysnKYkuKb+bHreCn9E07NNYUMATcAzHQXYjUIgJTxh/6VLqXj8B6EN1Hs2IU
ZbruGNiDgkHxdO44fPKVkxevhLITybwfLSoYSoNUqpqBa6hgKTxh3t7kVcKSIACg33kWDn2c+yQX
Eydvdf9bs6bdl2xPLfWeRLLMmxRNMVwuJzx9Ix5ZF6cR3WJsvlTq7wb6KAIzzpZYCLLiXDKbmris
fJ2QOknjuyh5jZptgAb4hsQ1E9ggRY3lvrttXdsiRtc2/a3uCxCz8HcG3ztbLmO4MEoPn1ekK0io
/rOP9zus8+L8DHdIo/CzFUwKeqDLhaczylaTAsfUgKI8uu3BYstdFH/Yg/xGd8FrL6gosQ9zgcq/
X3eXCAk0A5l2Btj3Bk2jSLwTO9Bvcdso5iSVyk5rSLo7iwB8wgcv6BY8T0pK2Rp/ZyM8TjTDX6sq
ujiS7OENaZbluew6lNozHV/Ugf3X+DW7syZGy2A4ZUDtiyb5Ne516/StfWWuCpSAELowgn1eoPJv
63UUn9IlC4IJRQZOk0bdkPpaHuU8KzICLdvI8p5TBKWz881rscoPa3pvLxzpeF3e/66kCghDWhod
O3tfCARpQhtwSxRNDIvsBOfRhw9FogGmQuy/WGG2Kjg0Pwv7uPq/2bDugbPtu0Gswds4SHSn3FzN
NbvAuntwWLUmvotvpJcmN2j85q3wheS0kUBZSrCL6wgJ51dfpUa9MjZwM6+PJs/rnLpO+FsmjB7S
wFG7L3jYOkoEyIXFU2g/D6lXFJSu6kT6X0d4kxwoV/ESySZU6St1czObdYOtoan+TRmBK3I2EB//
HqXl4e0uaaelGCLoFq1A/5OmUPP3iobCJu3LUW2DdDgdiQ57nI1vjDbxq5LGU3Xz38u+TR9ZvvwL
jX7BtnxSlFjacp7AIZS6uj8BcQZRIhfBoj9apzPB86qdYzuM0SJE4Fj1+BUOr/P9ZV93nPbIbWGe
FpqNtSFe2apP9P8jxolojBF6GWjLI11/1YB6VPtnPSi7I9oOVD8jF0fN6NfiMKv7lmntyCD46BCE
KqdYitLUbYv4Vk4cnnKZJ9d8QpAvtZnx+Ngvg9wTsKrPolIN+o3lVqgr2ec1U6+BQtTpQdSm7AFD
YfGS+SkzIfOgFHgRYI3OdnLOuSbj2Agjm6FKM7ivvyE8pFmtkL4drlYdw3eijcgdPDAFulRSlEyI
bXTPPKmqMpIrn9/ihuG5/DjtKTR2P3w0C1BdMH2n3cY4Fk3WBplaaTEkfDC0CZStNLC66roLVJXQ
lhPHxHiLPfe3ziZFqXmYKPiOHkwbN+wxWVZs8PhNKTwJo4w8UIgTpcFdjFyJTFHdks+3km1Ebgfx
yQcn93eomXlAqae5EwpzSGGKqqxeGreveCwN04sAQUd1bhzeKr2TRbQ8m7ADJ2CRfemybdqsZZgl
uzuMj6qFxe3dAUtMUDX3jsYMojjQJkKjHKMXvC31DEJzCM852w3glZkCw33u+iIic/lS46wIY52G
71geq1wKReBCNqypKJK7ZBpmKuUOqagEccPtdSVWS/V5uGaavc31BwYPPyZi2S2vkWIWeNvH0mdk
g/fw5vQtPikabe+Bj+i+NMLv+h5rXAFXoouZ5Eqw58+aj83tN4QJaFKr3LfQU2VIGtJ1raqmf7HZ
/9bO1g6UcMVvWJoAgkdYe4xRqKADQeN0QEsR37v60qzBGMK9AfoqlpggvD61wICl79vavWFOplC0
MtdJl5CTYrblVQCcz4NIEN1VNQ1m+qkl1zZFdL/s0FQbAKLLUO/QqL/OmzErcMQY2d9tpWiMCkPo
yFMRDVwCry6+DRTyz11n29uwtU7z58wZL2J2Xpp96FAmNIcPUSDj5ikvQuXuhRDvifFYS0RvfpV3
tiTn8PgoscKDQGeGnUmFLZ+MR7MKlkAEVwBCNOSnXtp55ypmHBx4i0BkO3TUr2eC7gnhcf/T0+vT
MCo5Xe8EU2ELJbpnJUKFNtF8v3qlMmNoLDJODogiJQ3roWgIb4o0sKCmfTtdp1JockNZUVUKn8p1
j80V2+rYXcQrkfcvSc4+o9St/uaBdt9WGnXrNGe8hd1+9I+sgNbZ8SH/eMzopCANMFwmwWuyuXqf
rOZ+QdsA8LxwxvtyIN6uxyaLwyvjfMj/+5pNULZZ9vV1riQBFVli+EZxiMsgcbEjy4yAmneKZP66
s2P1zts6N7/H0HkUDVzDaKqFgf3e62NW8ka7mPr1k7/N/X0xZFTws59O2mwMUrebC2gxiPG+5jiy
CUY9a4hprI4BlY7R9BInukXt9y+C+pFu67vvtZH9/+O5snzhBt8w0zNZ3kyGrrDcVJpFpHfeCKL1
+NzeLqUouKVEzyLq1Qv6HkZmB1aqvS/Q+/Rme7FXUUT4SqpIqWnPqKiz4krdutWV/xJWC0lmj/q0
aDAIh4x0il0GZhAaNB6EgDj9G0SmaWB5ZR7ooidw4bWHLIF+7/D4LSPvrV/JY3rf5rA532bkHbq6
lRptZweI7ZAh95W9SaHr3sjX3uRzfTKwoOjX1BbnI74mKTlRt5iQghZYlpoJBG5icapQZ6ZQhxPe
N0vmdRLrZHRr09tPxLEozBVQ4wKyPAfI5Kn7y0cA1WfUgS4qkaJd0q5C9XqocJAp0BXargjfSzFA
SUhx0vIqT4+HHbwTX7H/GHo9Tz925tDVv6k2teOBtpHPL+3k73+MRpirfux5Xax1XWDmue0m0OKN
a9tKgcpknkvGsgWiOdgYRBUNlL8vAiHlJv0wq6+8wgZqnqxUZTY4rbl19+Su4KYGwEbtJZ6sLjYW
4oZXVdLSD5GVmg7UJm0mF2uhRaPgBQN/elUXa7Uy7CMIjGcQbb71vGttkYUz1QkL8i5MLfng6Exr
AgwVWZ3RGLW0RlR8GYMs2hsCRdah4FEl1EYAKpRWSo9Q1j+z5AU8l+6KJs4UQPpe0ZXvDjfJoN6x
jOJkDr8wi5wiMB0p20MXtNx2nqxvqWD58m/QEEsnO8/sOEwO/v+laV682ulRM8aM+2+R5UWMzMAO
mJu2IkNGiqWr83j7m4zMQ4cdtkAB0FMLKcXgr84Rds2xuRNYM8FsLZPyBcxulitaF3+CV8W0O5Do
BiNhqE0hL1waZvw2T+VDsqAcrbAteHtv4gc0Iu1VJpey3Ba/LuN4J0827yjJPwK+7AzjPJvQ/+a1
78CQAyxwLizEb5ng0cuRGOKrNslIpkV3R0/lALI3I4DwbNjnYtHzNdX5LXcBB0GwLp6zZ7VOudys
2AYmNXQfUXkiYWw4HDSaItvTFzXXakKmveCRs/8FTSsFRfIllLvBR54HIEKFbSe3+ByYsMRI2EDw
kWntdGIiGNmQtK89YMa+8pdI5bg5mCiXtSs4t/uMzwUxGMYoZQTZ2GFuykd+tKOYMx+KdP/Ofem+
FQ5CT4Lz/LJ3DR96auye5U19ECSGp6UnCyVHsTjmBL8LiieNHdPX9kMkU6V+wqmRm7dt8iT/J67d
yvsDQ0aG1YaK1+U0mAXqGImCph9Nsh3fG/KDAmX+SuHCBSAOSTD/3Pph3rO/4pr1iVGgXWg/Npix
Ig6vipELbfFXfKPLQwMWVbZAiShtxGA/PUE8NSZZP9a2RgE+wKHa2T7bzRe/njiTLF92BjM4weMt
y7qf+R9BM8yaxLPwagCotJyEFy7fRO/xPfkd5fn1twng5OPtsmFVuaWfsUmlkQnG5ak96SfzXzKU
H8AsgDjKjavSUa47YCBJuVk0Cn0bnptdwzkGWbWXq7Vays+fB43/DRyAxBcIEJO0I0Yn/KfZmNgR
eQs+l0ZhtFtHkVgP0lAaLqMrcE3V29p8kM3UO179SHqTs+6ihg1YT96gMcaTHUHuYiIBLEiX6ATK
SUx0AAk4ZLzyKdADg+NfvRUlBw4mai8bJSGPFTOntxCm0cLbuCdbg1oP+AjXN2SZ/RKy0KAr9QW2
fgUFSHoBkev669h6Hnikolw3sSKdI7322mlcez3gZFGJ+A/aBqw+b1O3JXUgpqDdFbrl2TKMssCp
2MMOvmW+2wETPhDDEEDfmzJjWftdfkhu5y/FOJqSWRsq5dnbbVAJh83/JOxL31bx21XosFfsj14v
VGAaq9fldx6/m0oMhAjAQffPn6oM7JxNtY+dOUZuJNnqGZU8pgP+ug51m8OZ7wXETB1jhxJXVhQe
nxdtuGocdQmQ2B3mQt9/7ei7XX9N0kdwUiumWyxh8ep7/V7reY55at21uTI658k/xPCKG+S16a/i
Fpb+bdi+LpSpeULrWFc8Ge/hMIbHP1Gzyc89dDe71KP2dn9VMgqMe9dhO+RCx33sxbvgSjOC1MLj
el8ECHlb0CM0Asgc/T/LMyVeh/q7sVMR0qHNtxbb0jcX+Up0LIHCX0LX0pbvKaattDD8rdbFuToI
iVE3dHCFT4kWNSLjgH6Qcx9qggFU76xkaMCCp+qBmKqa/x7R09qBaMeWULk+boC5xu96VGQpWtdd
ou2dY3G8TJrQMv6yU86cSFI41hdDEsJXq/H8jIgOehNoZhH40LFsUKNIo4OYzUgytZa4JIvDEyAB
jw7YuCOK61q9cOPc6pBCfwX31cKfsADXTTJn+QH+cgtLkXPiAsSQfyhQ/xyLEdLPBEYrZA1+sxVK
IyIt16FfIadKpHzepUSECqVMwuhLtkSST4x3kT7lg0HHf2IGwUT6tnJg/kTVWV1g9O4EtGtFovz4
dSRTy3hrTcsCWixtcA5EOny3ly6i7iJiGrSCAFeH52HTkFptCo7dY/v1BmgjXa1zQIBcgADuIcaU
FvovPBR3EZgDjoQnu7Na3uCGj4uHhkd85W8kJY1nVmMfkC+Gqw8DNamVA4Mlt05Tw3PFY7RIEAUD
7lovMcknDt3AuXj0TcQuXBlCQnrxsIq2WZkBl7fMAgeNTPxdVaIEgPLZLJ5Q1nhK+bpBvULBwrqC
aMbwt93+vUY6uIkLPC4PmAcQ32dyXmgFDulL7DQuEwUTupla5D213oDe9JFjYamdbEUQtCbJl5FF
SmTYeyqEoxxp7Qw2l1KW9dcwIQapJxTgvd/okKnHxejANtQquVzAJ7G3TM3W/CR8c7b18s4L/PYS
nU2C+bWzTMYLq0QQmHbZPkhlgMoufk9wxFKBTdC0VAW2I5qApTsm6B2uN7rUkchVjLFDKbl0lxb/
ZdjX2cId+MJtypWyYzK1Xiih+RCjpHiLJNvNV87MCsCjvIwsvcyj8DjPMx9JNYAFB7MPwcH67hcI
PyKMVLHrpKLl6/uvy17IA04LmS9LZ1TKstmpKkaq6fSBzMTEzC89yeyxAKQnE4dwNsxK7meAt+4r
ry2B74+awPnIFCIbMYPpZlW4mAcgN+WqhCvlBGW/g0BAlHuROP+gQNyljcjs+98gPRaAkmlcvSB2
2I1l4/ZW8EjqbgjO7/FdGv3Qy6SxxDc9efoAfe3QBP6quxwWQxnrM/YjTHxuDnw/nNMAl5e+lgsC
92ENgeMfW+uZ0ly6lorI62K7TiyjpjJnilwIpaGaTXt4lHZMMDUuGzNYv8lCNFs2NhAYhtRlnbGb
u6NJjpTaazoSN24kVUktelhoOU9fwztuRMf62zhDW3891+7Zz1Ua25q1XHfe9lGy75C1ATDGkfll
Z72fYyvCs+caaZN5JaaSjJUAeu8+s3vNVs8WL6bUyVHJ7dLqhtLUPRK0KaHi6aLqMmRZnxtx0S26
S/59sP30Nbt2MbzWW2t5ZXS0oMyWSwQQ5HEuoW7dsX3wS8wXm5kPPJGSd3CwY/zXpfpz2wxpe6Go
lJzuziwlALNsIZ5QicjaOsP+YrQToJxporTWIJSXCVawJYfF1b2d9a4O7ciLbiDsseodEC3rynMZ
tFctzjS8y309BNWLExVxygnO2rqUSu1eshIj+M+sBJ3WWq9t+7Ddwhy5tgBP4o9CqMVfOytrUwfC
UhYXOT2IhA6dlMIMqSmcBbwMQW5Ul9S/mApz/PFlAj+JEm0k3mPL8SKZsdNvS5JU2PShqwpGEhZi
3pvVwR8kCTtIbw4YqLsn90vpnyXWwF5wpMgU63ADo6xdwziJdgZttTUnkTPbzDhSN4s3CVE3Usuu
nM1mHeCssoVPv69x6J1qFS9dzvXAKc3ZtFzfz5PiNyhl/jAuCW2dj+ybXZXqMQYs694j8FxkTLMK
sYNqabD3JczJ+oUOBKTD4SK1PUQHwvbg74McjIkqHtwf0sJ46132BMqWHcZ78VEkyPVbeeMWcyJJ
y/H2jrzNx3u232PpvPXut8tyw97qVxXxubco3vTZ57XMncQrsT5RtlZ251ST16C4r27Qu/1wguIY
wCNrS3J+WJvEkcVACPVRtOm9BNRXwFWZQazivIV3CitpyOzl2OVYBOhaNpya6RGWAf+t8GLbXLND
Lv3q6PbJVGLrygkiyZIL/NFgirFN7IMdJEUue96oAhjmScWgEzba0IASERL1+ajtKc6wEcUA021O
rz7Uz8KS1hXocCHmWllYbz/iPgp2ZONFLC65rLsWeP1UqlgWdfMNjKfFQLJWqXQi/Y2rritgGui4
Ozk5MF4WzQza63NQBN9GDZbFcBWEObaXr5x7tlqAp7FIZ5nVXPjBEtpd9S9XxkO16a6gQ+6BjbhK
rR+vbBTq7M2XhD8U2B5h2pU+CSIzw6qgqxsZ+o3mjNVrwld5RronNHVKe31Mq7HEbGD7stj9kpDO
qePW5Ar76b4q+5Yrq97ngV1vd/SqiVhT9vqmP0wyfy1zV6H6Z0gFI4tQF/16uSHaET9+sPY9uz0N
FVeOFBiHIJVCGIctxT9MXaRK23uZFByu3GgLIaawHkDeaKk/SWDPD1Wv3VWYTqY4vSuFilOzsOhL
PRG9OglPMfKoT0IHVpB6o/uGDAb0QvgvkRvS2wj740VSE+BwzRuJmihdeBaGniwMBuMvs2ZsUHsf
M6tUlK93NCDibC5KSCuG84hyvQ5PAxXmHUaAhXK0/d88xZpXJYOlUCsw3Q24hjTcaI9bQvp1Szbf
6jHJonBQkL/goWPOly7cYchNWCC5OK6t1Uy9FBTPk8soNQQzxoR6eCqBGqBU7bh6ICo5q930RlGn
dl38QC4gQRNKirQF8ZoXiLxAkSGjSY0GUfWPBz8fD1j88SK28fTRHHJhXUDTPguRE3FbwIznS6VU
pP6GbxVVqncw+pobBjWCgUSvr1wsmGe2FtKJ9QQc30HIuSmI72G1EuI8QdlTWw2RGFf2ibpZLHM8
9ugjCYT0BHyp2lshg5VkY7tphtuFNwET3JdbbVnxpo4ms9FFWdYSRlYPT2OgPCB7ehx2N1qN/r0v
8cbAWVBv0dx5SwAHf6TncGZ/dV6OXJdl2wJmmYqwx7P4qT1a/437GlSLQk4RqT5ReyUrCG0K/g8z
Q8WD8qO8q1//oC+U+/Rykyl/3qPf0T27hrnWmorHmCcpppTWs7jOX0LHak1yk9LekkmOhY+UkDFm
O8/tphlcvatMe9IaQXjOVPrjqoWdGTJlqMkTrl+8AKq6KZmReOHskdgjLWU+GVMpX592NoCt9Xp0
4go173EqCDALzLI1J+W+0xWIkih6B8GJAFUtccWWpaebt6z9heq0limcYca6uQ+yi243o8QGDvQP
NaHHFYnEGH2fhZc8Yx4akZ+7stHNAwXFULR+oT9NT0OnZykmNfipj+RYQzkSUOvaLAI3cX/o7mIT
cxnJeztSQfjqBWkSj/tmZfWL5Z75q5yChG8XnAVXREAESdeqipYfe4vvgmYvAkrpqjB/QncbAn9U
lTgYMh/Fvae39Ivmwmrz7/j2AjbnSmDIHjKQlIfBVgDigv4fvmvi6wWsp6OjMd5JzsbIpFQ7lNSo
6ljEfsaYpwBAmTTmTV66qi4PKFv6kv//zQCfXdqGA9pHsDQJ+GRqGkeUzXZRcbvtHNRKA6oHx253
swFHzDMwhAQ4X+AMyCDMN2fLJGrnsQkC7wj5tjzYMlns0jH+hxXvOsCUrLwoZDWv1ecnXrDVvhi2
KrHab3+uDoUrPzPsfZWoyJY01P5L31X8LdIsPwUy1W4nCuqRhCtkccLF6/JUOSe80Yp4GR7im2kP
3DI21OeSCwcZAGiNOwVFr+dT7dCrery00+9OH0BuuWXizm7ebgh3qOMMmkVr6WFdA78vLhMcRfz3
on1Ogai3VMercivnq96esIr8B2Sq/Cst5AiDrp2VC2/e0725GB0gfPhv2dyQIxkoOiClGKDEyv4o
0kLeBkAaMA+5cyAoNgn83WOVW308ukU3lTnDvh4uQHEL/vbafDwqxseAhV+LCJ1O5vGuNjuQVTeo
S1jeKK19CzIDejSMwRRKfh1+Qjc2WPDw2zw6yFmgvYK5rgmJDfku9G0fM056uYP5TmMSk4/Wd7mQ
o1a48rL0WrLc/PurHTatpaNHSeYQHvL9GR5DFanC7h9SvH0uXeD8As8zBS/1WpRKFhtRfIeEO/tt
oRsc10/hfRKGtGROnXxOmAr7BR9eTPIBhhcM5tuMrYI9j9vFJ5IGswSYTFUlaofSbiiKuxufQ7O0
Op6GlgBE+JepyQYFm2ET846lvoA/1iZY4ILy01nz3x6eaUf91FiVlM3Vpfqq2kDKpz+gAV36VQ6v
OfywhfLju8/+lhXQH7Q+n1htPs6ZYSshDZJhI52BW7aytCs97ApnlsS9GOjHWzNvkU65SWm25B9b
uMsyNXY+4emlwyoEFXtS8UJ47LRIOnpvksNBov4nLFOv5/RvIvwVCAUg1funHM67vTBuK9bfK5j/
xZEN2JplPPWMYd8ilp45vWhqw6SocLwBr0Qo73oZhaZ/sczsw/WyXHyqMbxvR4YVzFrdld5KdIa5
wj72gdWXRXDohKfpT60XXpKSy3+EwqpjexFLQh2RMezidi8DeG1lqckgUBVTGE9apl7ISNSUZqOE
kMHDr31kQUZVzGCwTJvyjpvk1i7pCAkcfLFDJ1HAPBONoXEGssFML21l6dkeqh2Jc9T4z+t3+KT1
zI8969KEaYc7AAv4dbznR9Q5er9zq+RWhLHLsrIyzukB5ufDOxG9Utpo/gsk9JR4LhsYKsQdAraY
QBwbHO4zSAniAtT2c+NypDd01Kcc/O2uM+pOU4OGFoAfOBRoj/CJSDu3V+bGZ2XVdyJ5OJn1XH3+
L/QoByPetRt7WWjSnyL9JxtLhd17POhvZ75hP/qa7TAk6fRdbOVQqYex+SB9PgWxM6z+/6hiThcV
ogFkVvdSZ2m/G9RuJALMvXwNLhDkdFu+hAkNd+mt7eMVrmCjhwrjP06ib276dTjrjE1FDnd2n4hb
sDEGlwtudOiYZdx6WhnXZ+wbG8hr78V3u3m0JQ4OyR61Y9Xfl+K69QRbA/ltXTCPauo0Qz1VUnRg
2pzxGNJRQrapbn/fIgODE68PKF++dhM1HdrN5/7pGM/74NAOqOayApJ64ijmC0qg68VZDVULGhzx
V4wEDCcPn+KLuiKfOZhaVRCE1v27g8iNxYsUrUya3ToP1tns55stFmAYPvlPvbTi4DfMcYr732jj
q4AlVKbvNJ3bE5M3sfp2Lckj6Pbysc/I9kDpr1vBGIg/rw/ZJMwqIkWZCATTrKnVUFV1Le2iDtql
abWeHP1LMeGjS5xDF1uTO6py35qZeShAtOq7floX1UXQSHIL5T0bNlk5UsnaAtXqLOlevjRwUAol
YwwOU/4a7YLMJRcr97DNX7cRgEDJbyExZd4d1c+AhVc5hstM8SCD6qN8MJOACRPhAyA4utikNGHC
1w9u3wUguK27Hq0lq0xZKTyMs435NmY96VZpB89uSkDkdb02o0pnI7BfqywGTwg4ySWFF9OkxQ7a
B5cE968w0SQZsoEcP3b8cvJejLkVN63mhfp1pIyXYKmwzVGJkeO8kPbBLRcA5w6HnzA6awL7NDaw
0rYrF2Ga2J8255Bd+go25XfNyIg6fDB2nHYIRK/F07UqHJ1xor4O3ZIyG1wTKf6pqN8Qhk/DKEKA
w6zOMU00CtIf10+37Lt+wV8d+10DD354AN3P9aL5+cvXhEa7nFXvaO31oMmF0NgkcmsMF6BD9m62
bCs3m2es/0yqejdWlhHoewHwzNwUcLvBVkWqMYsQnUznjACWF6NaYa1Eff3NgpTRNTgJg1ADecJv
7dp1pBkkqKCwGk/8f0zisv7FLpn41/n27Ui30VZ7W+P53nF3ZZ9XcNkOus4apOEYkyx46fjnoNyJ
ZE0U1KEF+A+WB3YbIpl+LcRxDOrj/089uzThMYWVEXqDGMkpmAx8M3B0sos5Zp6yqTflZYZneDIv
FDiKNMTdVAe2q2auOufhRYEdQq9mfbV7/6eXAH2R8W1bghhlHg8uBnVZf+d9NqsM6j2SDxYX4WFH
Pb0y9CKNiYi3yb8Jkb1rSsfpUPkzXHnj6S2IY+uHVY/Ttg+gnOk5QDFF7zY5Pxu/x+kcbSudLeC2
2kYEHy0ocTuvgCkjzoIIUZ8tjwsepOUSyEYvG9xEu1uUAa7RS/X+rsaUvw2jz0YWGmb6A3piQmme
wQF+XqdkftSngKiiwJ7SpSaZYCGCvCuFdUaeWvuLPhFwFZtsQczFYV3DhRlJ00Z11XYmYm/rSm95
qXuWcOEowrh/j/M14wMcH4Z8vXqvgIgUB5WAMqSJoFwgE1z4U3Ctii1By5CI/pz4zHHJNosi7lp9
orleclSaxpMegJnX4kjOqAe7bEjvwtShIPuJSHTkRSORDK/wG3c8G/+ojnYFKkbV5Ad6dXSd051o
1Pt1feNzi/4dj5IusHlaimI1VBo2mvCigjj5pmOmHcfF6sX9r/G1aWUF/od+UJE3tmb+8iCKalHz
mH7AHf9OQqUSJzsLRXfb8b4Gcx+o1LuqHDAnUl9HIWR1aSC4Q/h5/cv47dXCcSQflN2Ee73n05IP
HJA2MM9+vM2fO6Xyrg2DOBMaflbFH2N8tv0hNStF0CZXN0NvkmW3vyddm9By88GiMPoDaARGFYvJ
7BOdDZwoDoRU6EKMwJ0OPR9c1/Pygn1/LtiPjIoBytOU7cq6oHx9FD3VSrkFJ00am/BV45IKULnx
imtHeSogsqMj+OjHpPMMeO3k9Zn6fX9enlTmuGXHdq8Af4RW6F0727je6O1yVU+ypVRJA9KZpyTM
T96ioZ5Q+x0zTBLlTpD3O/UxEU7BUg/kHJ1r66UC+j5dcyJI7K+b9wxlQqjBacHBQf/wdxs2REYC
y9p1Z5TxTUi0QS3NAuAsf1im9nVLUgvu79Hgz2YehpFnlEjIX4volCl0DWRDADcYu9EzkD1gmdPL
0VkojttNfgiyaqUWRKkC05mvNxHE/BnhmE8LOYncMJa6mYBAR8P2cNe9GgHxYDzFSQh1jW0w9eJi
tKgTt7wGMJazRyifFHtlxSdY3gan//f4MZGL2sMw8yA43TQN0WofF2/Fch1/IqY+vO4VFOfKU9Gj
dqFaPGDYjVXnyCP0EApjLuyq7Y+tfeLOgl4Cnki50b6T3uRdwDcWKW7ZqLGnL8BBrG5+WSPed8WM
StOrNL1k/ZAjxgkvW/OmZPtqKaOc0Cbygbl5i/PRgMLhLktXTGXjvb4h3AqypzcxJFa3sfdJkNmw
PFD47UP4ltypKpivcsNrERa6Ce77teIp3XpGlYB03KD+wtuwuFiTvt66QAhwX++xNMQW5VyVXW5p
A4sej2TAyHJnYcukedn1hqqRvBra1aIt9vb/GmN8XPUUW4FK0QP2g1FOeDQfWfg7rCIRhw2/C13Q
GbZoRyAP+1bAxjt8zeMPmvtil81l5L0z7irVhYSOAhV9TvBrTlbul9KPBERSdDbn+fD9q/kU7SnH
gVeT2+p0YKA1WJZAOWvFQC2mklKwT+xzEhIDQLDbGodOp7KG2EgKAu1XToIbbHSShWUjPXRr8rCQ
MdvY6i9fxcGEpyXgEhRrXtcKfgODQqAiIm436TAKDSiFmRiIEIxiozoce1tbGBtYjO/VX4++Pp16
LVVcCf0sm8ja2X9hIE+/8Vk+bTx49qCTPpnIxqrDPEKulDTYUzawW/9+PPil/usCO/2H6DX/FNRk
g2B/+q3MscQRnhTYJrs4jOhyV+HivohKaTLO5QUsjFHsmpUmOdAra4PdlGhkH+KElC0fTfiO253t
/fbnVmi58G/kgsylKvDfWIRuRj5l/QvA3zvBMRrtNQFxJn9Cckp4ReS1D0JUdEO7+M2jF9FiwsAs
a/WgmqK3b0+oW77qgVHWbgwWmTdqj9pKQC4pOigPod4OLih/tuI0eW8pq7t7GZ4CLLjisVvCGWjL
dFhc+SzxE7FO57+JdGFEJTrDfLVMVGQqoak6cVHb2pvGPYPb4Hrwnz0c0nC/YrkdaEn4Mizg6VC7
Ka+XadhVtOBVjZcbGa0rheMAn3UWYmog27AVH1eeSes/MqOsF7aMH9/jE/G3gUZsgI2LvpekvVI7
nXKnNn5ZbfKNZzvjeKzWNGPd7ZH0QKYrfjkC4h203CgAbexSlC2G+mMFybgxiROIJL34Wu3HwF0t
F9mpEM80ccx/IrGRl5zeY3fwksTbZAVxUGHgc1zxLiKRgWIYt2a/vWMOc5l4dOhlAlXwBg97DKl3
L5udtM/+6ksheKz1rC/kUlGftw4hchCrfaO+tfwoyCA7b4PRiBlmexOJXLqNqD50Hkmo8My33toK
9sBeamceQSuAHGh6+Adlx5vhCBdjvqG3nNMqqbzfCjIhm9TsaR7R/BWyfiZ/BXVuYaqa4gee+jH6
+6xw/VlD51Sa7wSNjs3vTenFRTlUs3Bqw9cK9sbTY32wbERIcHuYfdS7xGuppBkRvkPLVEx8flHO
cS29HxpLSg/yIIj23MW45H0XCnFxk/7Ak7PeWdnuN+BGzEjbirgGjQtnGWSeOpmz6c93PZB1kuoP
mrjc7mCsj9u7E5SGBs2mEYm+WPj5Beej7lhloYtiBLZHNsQVJsOkG97D62DUgTJ2AdZThd82Kog2
5pfw0lTgrc9plkws81IN3Ip74N++uL2rx4DvF4vNldhMmWo5U7w+DIHfJ4Q/7ZXCYc2+DmLp9PLH
Cw5B6s8BOfHVQeNW3e6jc8J3xRvqI68l06Qpcbv1eGsUzufOvr+8ryLkC8XkdhsBSnnixtdoQjnM
GwHAf1U97ZfPBA/1a2PGLdLQGYJapVGFc/JwutWTs+fMhuaOY4n/ScXfsq17fP6T2rbKPG3ZYLa4
bc+kGvjpyDf+eepdlu348B472hnoPIjF7l01rPefR6dm/e7AFSEJagkDkLC0PbFx2sZmub7rygG5
dfr3BR6riOPzWRPg3DbCXD2fN3hjYbRHQPZoTA4upLlBWo2w9Xy3WrjCs/qClY+LsawKuUl3Ctlm
b0Vejbyw4xXJa16hTd95OIZrU0eaGJzq/40ddR+4yiYu6NGKHyIFqiO+A+s+KdqlpP40q/Y1FxK3
OpulfylVPvMUwClZszKR+R2vJ5nJ/6UOzhUyE/Lc1IP55aYH3NjS6VoOXamX7VcNVoby8feHMleG
miYjst3a76qH/RZcC4wxG8c8ssFa/JX4IxURymGxSItrQfAfmdcKKEb94ftysnL3NEKnEH8BkkIl
rYlpU69Ksms1iYCAczkS26e3L6KW6cLF90Bou9fWymabt8QucVt7hr5CAnv0Jm7j3yhmpj0ybkiE
6xJrT+bH0mOphWO+lnZHmE1mEzrZt35SrxwEX6YUUZNgah45kKPOzBZu8fs2Si0l2/UnnnnUK8HK
a98H0L4uXtvKie1lxFwkZK0o0gkbRuY3pWLi/CvzvAhPyeCXTBPDpESPvFd+R90tah2CleesS2bh
dZkSDcTrHuGKbZ7jOl8x5MoLV9GU+MTn3JYoRtUB/XswawaIRd2ksAVW3ptO4p0Z8kbLo6wwgyXU
UAgWLRljRcN7XHKAPHboQ6CjXWWzc2OjZYk68dZjJOnz5faSmp2LyDXWQQkseXuvl7W0g/6NparG
VF8pa98mn0IyS9/y7X/lnmjbriDTJCnOUoQ3szYRZmNZG60mYB3rwAQ12SYfb7k7hpOOfclwBcFu
YEtkQE3W9IAmFsGV2mtiLICXLCMusB9vNhPfpOr0ZaS8zNuryo3jCZdXYXr93buR1kRqX4NRBHPu
9P+vxGpQlOb3cbYae4MeHxKqBe3hm06i2g2L6byihktoTUMQgmZC45JGyNkgBYVg/nm2yqR4ppMX
+fsZPnYL9Xf7ALiJNseVT1lcICRO/ClO0ZNNLCEJeqfJ0+4uV7DHRCuEvIRfisWjWxOJXKIFboDR
zxPlyzRRX/fiDbaTW6UieNxMunT4k/oCG8S5qUF7I3NbCHzwEbQ8az7VMtyMGxTBfSMSaPSVAuAT
meuLFl/WZyFp5sJ1BzFLhmNsHbDGG5cDc6zq/cEahUGRuDHAtlpClIkFyKEpeNyIaLsyoiI6rMUd
j7jysom6vs9a9nGscdbhed08UzsTdvB7B2k0zFZzcB7rMlwH9wpoudWFsQva/LkM07ykY25X9dZ3
uPZYemrgqb+TXIHdhbvAWqYvgsnXDlsV5bB4EnJstLjoxS7BF6Pf4e5UCTko78xk2dxE4ey/8AHe
yLKtsx6yI7OYQ5MG839K31qwpzgMqmp85+KsPL/upgoXjKs7+2ZfAxnXRFlDuTiwPDCAegzwDQZg
XhmiwNNl/zL05sS3PKJoxUYLCUsx8zKYMpjGpZ4O9qEwKMtAY/Dc47740F92tsd2VAMSFQURj36s
cPdai5Re3ke6PqroZeRzim8wJ1c6X1m61fqrAcaTPH6Z81smiev/GxXtwUlkaxz9TrG6cK8UqfkS
oShC50lEw4a5mIRwvKlqNX+boXWO01NTD7bD+ah08ON9UxaSp2kNakzj/4togYW+Qb/bPOpJZreM
FrdT+CR0qJa9/nXExasHkuf/VlcOjupX/Q8cX91Mxi/iPChlaV3Q5+muGdc73+unsFxBpBWJB7qB
rYpuRf09DxNn+8Sdb8HlY/WoZjhu2SZ+2vh5LhZYr86d307UOjs7U/gCJ85+G1+4/W5//r9ubD2E
4pt08N/7nwdW/JyHaGoZ7JxPIUlPI7t+Y1bo7OOhCRlfyKP4WR0PZmQRXAkzAliVoqIAQ8v1i/4D
4UqGuOYdj012aRB0rXAhBk1xnoruOhBgviqCSeDH+/p9VSdzI/u+69G7BHEiVmqAHNzFlrUlfqDl
pADGhc1Q+FiMWjAekkHeZ3xirQroi8bq4JOTi3SOqm7AjheT8xoZpVzrdZXb+lYXEgetWg8LR20R
XTEcc+jgdLcnV2vVVKkE8FRWXqSyuDb4usUq0KGqGNdkv2An8jDRJ8e+9su0YN2HCmD/+cMbYFAG
bKQ0FBWOLlEjJYhViOuM9Hv/69f8MxiDzyqKheHOYWynpKSnD03CSkvCoOkHy83aOXCp2+2w32rz
yFDPuPTYj9MH8xyJyV7SIipmKfKlAWnfUXTo95t0aZBUmjvKLA7hiCMPCIbWJGbTUYqlOf0XOI/a
H1ZwObuOzBMWktzYvu3D2Q+uyjJe4asM6uuFOReG6aJ1UG3Uz58E8ehkkEo7TkjwS02Jnb59k/4g
2pZKMhewr3FM8Twy+xq/VU5Zw+6dqUS5daeV4h7qEyI/kIY9u3hLYROyFT1wJ2wYZO/QEHIvj/A3
4dkpEyQ9snfKQKwnmTqa0drF7QhrzNESqXn8sp6tfqQg2ip18i7vXt0RgoZH01hFtQpGNISlV4iY
sl7zfrc93oGmc9OfJd1ajzqqjgm3pm18vepn5wA0skd1fF6uYJSQi9OopPQwMkdRpdqosHVHbOTf
Cg16a05agVrcEOz717zshdUU+drqmz1Bxrr8kqwsN7DAqzg++TjJlpwaqQfos9Vqm4ZhX4oS6pLb
PDdiwsKQkK5rN4tcD78vELIEBF9dPoPmd/Gokcb5eSW2kj88lKpeU/AsYcB50JBUItOHVuTM+a/f
1OkSzr8MZwpSiPMibo2V7vSHKm8GpN01hXnDttGsA/ROHyjP1WTKixoXr+8BP+4D8MkXpXuFDix3
qPM2FMdYGOveEVE2b6ZeeFZvi6cJ0vilSL0UtY0ODAkOpGAl+F9qPTARSvHu7DZPwuJyDZ5tt6+M
A2Dg0SyR/ujOtGToJrS0oLQBehW5/ZSSDVhmjBzAuLU6r52Qkg65kdsbE1j9F24SyNjbhaJedxWC
mwkOSZzpuHZwFjcalXSO5paS/6nalpUsFA8NUtDmUEpXrh+Qgg4VHvKkrr4FntRrUYM/cvD7KHpr
YyRl9VUQVanWKCi9nGXw/URslsv2xeic2sgRXjzztXO5gl8t8MtdftmxbMhclZskMhsjr7i2nW0Z
2Yd1BcNfMAWPzcDqUaDB+uBKw1KmvFtuHODBXsOVb83r2ogFL8YBSi/AQS5hNxeH3IKHPAjELk6A
6Q55BbCdgIlUzJ2l1c1JTCT9d5obHKaybLbd29B2+7svb/reAWOPQruXqdH8EfG7IrCT17U8iC+w
2+C5jF01QSZSBi/fYIFHw+OqvazVRKjaB/RkYz+n02HPKp0UtMIUuA/i05yNkReb4CjK5lMQa76B
JEZSNcxwtLpCFXNBtyQyW7XPbUbdQeVAh/fKcsMK0Pwo8mm7OGInJtJD86PXRb6Updq5QPMfU5IH
EWzWwP+aWc0erMxH3pqYyZnI/5YBrtZYJyZ4eZQHhz2mhYJW1o5EYVxWUhjiY5fU/aAVi0GvCL8e
BpmbnmMRxY0GGMYRtGFlqizYXwt2vPAAZHlSxWQgV59I78+8G1zHFMNd/Pu6/WK0lfTy/h43KTim
a4SEWOUDUkALkqch3Mb5W9h0/XGRgiSNsbeCc9VOtotmV72ThvOGIY0KHpzxTL80wxudrMsrS7Ft
UZrifFBgY2qLCEoy6NkigsZac4t1YOGg7jyk4k7wYizhHzN+Ib2zNqoHKlSvW8T2UDC61+50eJGO
Vyf6DsSYgcyL/gm8CTXqgHnvKGLHJ22bjg2U4jm4ZWlyqtoqK0YIOshnUTnEajexKcQQ9RctA3fg
NhdUBAKOiza7HEa+g4be+NgDtTz73/J9ceiScIx9XDryCcBEX/LT4pzkgR+UzjymZGCbfMVKMd56
awj6xDpT9V1RqT5SHzfrm8se1/hZWd5uBQMNjJvFKL3TJ5L4E8AoRLPmhIOFu6jNa/XpEK4iD2lX
jWyustHMU3WX2Ug1hVGTB9Cbbyy0GBLwJleaBluILu5YQy/nvebeQvPntDDKbJVhtnUtRoOcgSMu
1elSO+6lV4W/WQA3YvEetT4sO/071Hwx5TJb+6K52eDOs9UppC0GzWM2pHWeUooS8nboczCuokHN
qfyg0tQR7A9A5CJqGvxC+zJPoT2Z4D+AHHs3uJQ8lyxiwcl7lT4wFMx4JYx6P+05smbhpa8+GMU1
KNZ+yKFSxfINCbVoT9mLn3Kw0ZPBs7TemnNC17Rh8GK/jRUmbZW6+Bx2Zahq9Q+Jz2QS3wvEMimL
rh87UtxmNHw7zcrYvTWWO9tIcTNWysIJF2JOvs5m6XsHo9crUkILbC9IMVmyzvx2Z974Pd0HWHvB
JH/vV4Vt5jn6INEZkUrMpB53UWamR8W5oXG3MDgtV3iHj1wagXsq3GA3imA70S5xrYXD1SIrazmm
JaRPVY3QnipGkmjeCQpy94ICMTD/G+bNTetyfL3NtCG278L8H1Dn6BgkhRvz8ah1uqbmNjMZ8p/l
1j1xBoWLG4XyFnIfjuclxJLtmBPirrhjnff9cHSi5u2j+RUe9wWZfdmrjJILzMlmzXiD8L/zB57R
4t3coSj+GEF1NYbeFZsjxyzc86Yumu19+Sk7V7F2UJMl3wcR//YIzPAjPGfEWw1NzyXxEajWQBt6
zH+7QeY2AzZV1l9UAGW1oeH83gInbDXr2enQz27Yvc7NnrGWBsH1KRYI26K7JwovgbS+yQbkfXQR
QhChc998XZLi1qudqnl4uB0YuUy/SjeLxMcxtcirs1u5ZbLwib10Bma0LcG9a+r2S0vuu3p/dzoO
a7NzDaysIhmw5yTZEMI7/vT8RXr8c/2Pk9JryN5CDq2IuiC2aZf6DgvGMzrReAj1XYPTY9EFqe+/
l3JdzTMXcRylhc1G8mGZSGBtc7pHq019WAgmt+AtWy2TDRvfPqcRUnnezDvuxUD05FdzDsYAjCfe
Ryx+IlEAiaE4RIMlj1fOkQaOvvAMDlLtDn+JF2Is+xqxd09J+zQxVW2OjzZYpmdkIuIeOUl/2oma
p83t0vbfKCPBJP58dVgegI+RgFIv9H6MKPjRQplo3oTpNE1vNA6JhyWTZe6/b53z0EkAHOEPYrSK
WPOW1GU73Ta+YwHJf4yxBJTdQhX0H3bcb2NJW7E0W4BWCnq9tXIoPKqYWCcsMJ7CCWCAnF6JIW4i
6V0Ib5zPIDg3egD4BcVRAzGpTSwUX9/4mz/viIrgtMksMLHXUr7XrD9hoC3AayIT1nrXTxnNET70
A/nq3mTEgQt2ul20CLNBQi8KoJhVCi5kSfw5j0yNL+VmY3CYRbdsMixAuT45giwRY8/nk9J4nIaT
M7DheUfJ58r8DDP5YYlTDDLI+SVS7U9NiRk+r+mxPdsQsfW7qyNjvPmDd8Pn7H2mce5StKExNVM7
Ficy1fzB6JBjXZTMVD6+yUsuDoNT9vUxr2fOzuVSe7rartB1V2ExHShUbGoyVmlMnvKyU7DtTwXc
Lu40K3A0//Kycyph7ZAhFjVyzmg0VTEqEgxqq0hSHJh+ecfIAxFvEpDUV+q0nsMYOrsm9hozzSYs
mC2Z+RwVY/cExuw69OxR61V8nToAaSw6T7dhA4+BM1/211T/v12n3EBRKQlBIatFMohvDJ87qR8X
YeVTr3A1veo6i7eox1rXuXIAawjXDtgTDZ5DyssQpjTlNaNq0ZYaPmJoEzce8qXG734o/fL6Zzbu
FfZaVps9I9QTzEGd4Lch5IyHYBGqvXZm+oymRwejrvuM3IYIgwTDhQV8QquqAx7iH2uVQbErJHkz
K9cnChA10qwjf+cxgJ4rNsW+9j1sP7wwPtU0mhuGIR5Y3+xrE+CEipLDMT9QpTOdCjkeAdCX3Xd0
9Wm0kvRmnSk4RSMLUo793QVz+zk0JoAK90j7gdXn3GcrShhuRzTjQ/lSmDSKPN8jQhqTgdEKYpxC
++p5+Ozk8Flr8zcgKwc33e9Yll2ma0I4ZEc7Nw5gr8yLu3GEBvHJtTDOJUOXaGrZBIQDJQNPBU0k
U2lVwg29cxC5d9UZnaUyzQAWT0IUuHFRj4c9O5KfzVjfHSLAFGhEY35oKfAUYLwEDgXSG7jonqy8
Q9pQzr8NCN/z+qpJBxArlkTtoZegAQueewON00noAf6SkwohQ+iqeHj0GLzEtfDF9tu1fOB0hkWT
OJUEXi9gdvpmoXefIAu7Xrm2HnuDTvJzSiTyQ+eMh2A/etNQgsMRymCR7/IllE74jnN9NaaSFVhX
MWqfS8y/vr180FQqNI0enCwRlaJYQAHdQXhHQyVR8jmIAnAz9W3TxkchntTx0UZygPbWttEHmn9g
5QoPPB4E85pxwTPCNzw0Ckkc2yKD536LBVy5+Oozp9pYrgzajDsXXM6Ts6sMHv1qGxz46CWaTTaZ
prVy59pfsdAwEVe1SzdZNVjhhgcxMqXxoMhlpVOHb1y1SuyEzenP1qY+DOI93jygJ0UE6VHm9rHO
VztIdSNspkAy18V5ofoj+iLl6LkQp2hPtYdgi/mGkQwI40iys/zQnjTUg80pCF3dbCc1c4NTlTsH
6YQb3CGfLHoVv0Cqn31hFZ5ZbF/D59N/8fN0VchAf484aNOigWv9nSLuC1/t14Z93sPqGUljeS1z
PYgR28lGrvZW9RUCG8Zppl+dqLDCfzq0MiEfA7bBDU6gs3v0mpWUk/jHYgFgakGJ7wAjSkmhkJqC
1U6iZD1eYVyOEop+ur18gu9NTcPfzd8PsrDBJAbixRxCmXpN6eP5bwUt9gC/9ECeOTCUvTyCnzJW
cYdFopUuwblcG4TwFVV6t3neZG1IZhy0iDVfEo2YE8TRROzpzhIgAyKwxLOy1bYB+UbLbVSzhgRR
Z6Oj6e/Zy6IBrmzqg7FEpfyD9M9WvKgZEO+Qug70uKGolAoQ6SM1TrIqRWuEISPqO99xBHyQJFvW
ALLiLpZ8PaXDoH4OqId0YZQQMI+Nq4p/UOV+KUwh1MH3K/QCg8yJKvjJd4eH98cJ4EWPSgKlKXNx
K18eDK3N2GVb0aEFV3p8i2kVlb+LjqUcl/UE4o/GxGqyqvsnsB3mXiRxmLxGB/eGqKEK3NYsah56
rycKQ0g6uKVFyI8u24vNVaVWGKozIvmlId4gEfheUAE1vgYZtZHQSqeH9aLzZJ2a232lRYoi3chY
bCR4/ko/uW19ebBuIJLXMMRVcK/gSLde0DrUvVA9R7kKJIMWdkHfJY1FfEFYDelF8m3L1kpOyAej
JI8RvPhdfMKGxhrc7YfifMFGkgQqXXQe0SMJqzXjEbPRPvKfabM26jqirorMuRXZn78LvIalJURB
UZjzdlnZ4hifbl5jOVC9VlnrrmOiBwlEyUxEmcsfeaRSPKvB+LwABLkg1yp1d831+LZKCLhoJ1aq
Nod0JX6j5Gikhil//YtbwPg88RUGYf3IW7IhGpkhaZRoviy9+jmuUBWODoGiVb7iqn6lwYUhPz28
BF1j5hNKR5PN/b8xOzZb2QsbpEgvkRrWtSvEaUWpQU4Gnm3s1zOtvqnCd6RiRFpbdMHOvVDJFTPp
OTT3H9FnvFloUIqYhGw3K6P+dxOwbO06I2IsYM7LEgNBtRwHfFoEa8nnYFU8MBMj2ESJr7X6ohoi
UPghLcoWd93imP9dt4BCZHSZD7E+iSWFaOwNSh/cdn0V1QbCH41NYZCKmfGE53crx/gm7aVYKved
bAOawgUWp7dJouieQ5i52XMkqFuJ8FSVJZ5H08IGoXrjJsHv/xMuPEPP0GZqnua+sMBLb6VQ6HcL
GskkflRyYhDW5Ykwas+ssBCRjd3fJL1gxIITc3AUQNT3R9Ndj0OKlUCTzz57eJyQMZW5j/mYqDat
4kb1wwiQHq531MoGBFIy8Z5T7eczsGdO5VqQNsPp8gAvQPQsECJt1/GwKCcw5q6OzFDm6VngipGs
bKMX5xIcQTyNG2PDrUuv5RYbC0bMFmM9qqEOHCc+2Oa2wh1VwrkCPFxnDB6nnasZET7aLOYlWJMd
dxcJZSweJ21XJAtukDDhG+BSk2KaP++FRHA0c595DDoPpFW1q9x0TCVSPos1wVMVzlzkJtwugvUA
WVbiNUouS1JYIMbVSMUuFICtD8OO1zl2elqPfthDg1P4Xoi4kgsIOOb+9dz9IfMA0eoIgHdNXeTO
kyMoa6WupdP7N4V1LtBCfv85r7FvEfVUxaXVQp1kPIAxK6OEMSVtpwKblUDHS/ynaq/G7izKS0sD
T5mrxg3H9ISYj1l+DiJ0oHWcYPGd2axtzA9Fl4A7U9EPIr3kINj1cj1GrD3yYBCvfpheEu5jj7tm
l66Ll0SGUr3knK1H9Pvo9jAkvt4x1ED+TE+dRJBunau0st4iPUiJyxwNI4VfBlxjlpQ+SrEGccM0
ZPmnA18Nn7b9Tot+x7dmnvJszTkM7IWX0G/ChXMvmjwTHRosgSvCt6YywSL72terNYlIdQD1iVgk
55fc61GshsUqUl0l47rv0E9ryOP1kx6BBhsyci/bcE+etFVfiHRfRJW4eowI0KhtWKdTHqiJowf8
qxjO8RtCUK+uxLGZj0TbbRuaQVqNIKFF2J7T3zgnL4yPML9e9W5JzHTluS1A7xiSE7wodxVPjiNO
yvQ6CV5Rn4jMjWAW9Ip02iobLqPfwQZ1Xd03o+UJDvayIiALfy2oiJgAosBYi3xuBNe9CrNVSmAq
JntuOWDoZyyUp7u4wdsU1azCR0CBZ1sEljNoKr8EAZBHrXNv7PFtWYVHHvE/Uuwr5HLDI0onkmOM
cKKvbvevM0ID5PBqqi/LPXMaeWb4MPeKmC7Zk6GQJODG+IulmXBioVfXmeWWXfaFEqWyG/QzscNp
G6XI9o0op/4LSB+cQBESF/yrtWDh+AeJfohGSPlGvR38wqukDB5ywpr52Go+5O2qxDdF2Hj/ZXjb
T7zZHZR1B1j7LG1frugTtyhYoBSvLFEDFXBsdcMjCiDR8/I56YMeQ1IciyznU+S1iGzVYF+LxW83
QdZVpeh6C9+YIDKfDFmQrlJ90tEMVnKY1Y+j7YgtU4DtUh49sdiBeH4ZO+Yn7HO25XUq/xS2MaVu
ldFSI7TJB43TrXfIxqrBslF9uEAn6J9fyYL82BiiGOw/gcDddXYCaphEz98YwESQmDIkLN74xfCS
AeD+h/6t9p4qdK0sM8FBu/yL3xIlVUOtu8F4aLHE/lP80tcXotA0sJMPaUKbvuZJviBxl5+5oFBA
HB3LPCoc/ZDDw+9mbMJj37F0RoQjKax2K1oMyl+tcQ+D7u+DXiaM7UK2BPzdVa/wLYTCO9w9UjRU
xdpHsZ/OJV5EboSjv70KeYflbF5nq2QESniS12JTInXhzN1f5Kt38L6gPBlapG+f0bBsLXzuwgU2
2XAt9IErcEWFwAB+TV+hvvG1d13CBwOk4KhxXn91fhgka+NtkgpT/gdRMxD3eOTJDEoWDojFEyyG
HIcVppQkm2yurkwvInChJ0+99UxISIWKIoU6oPhKmOdZIGlvzo0E3TSU14WNZyc6iex8MIuohMoL
jftXJY7luMe3Sms9qzSDC5/Tu0Ds5D+XVEUMQaH42Jaei5Qn/hru2S6lzyXJppgvjEe3dIgEq/7W
SsHMp+mM2VcGzKU81xge1V6+dSgMcdIALN6qagwTQnskf6eQdAwQFPy/R6/izwexKls67CwXXtjJ
EgLrRkus27fWAVuO3tAln4OarswOfd4ORHfPx6/R9Ln/xdx6R2UtmdMV6loXjiPPd/vzehmi0nAq
Jq+9U8R1wYhXSa3hI3Pk0Qk/8wXCYxXDiwpp0vBx3yn7acuxObrWejn9hbRMt+7GAxVcPk1i/vHr
yc9ICkux5DNnWFtq+1+TiEZKYreMLHOYQhGIsMVDaBb8nBDu8WD1Cy0WfWzKVEf3WA7YDE2L51Tn
WQnMuEXvMNxfQ0KWS3ACW5lCUGl1mBRG0SOhPjwt69J2CjNttVGo8HSxWolTesFoJnt7nnRDu8hP
tKiE3NmqmKVA9XXqJp+5xltmjN3SCxXSj8ENZA8p3SqRtOZ0l5j06gPBkrsRXZpAbaWzlEvUbf0T
IxnUeDnOpO7hZEUsGUEWC77Ca4f9jZTc8fBM6hsC7L1RW8Yhq37N3yzjWBx+t9AkpBvPSs27pnN3
Z/kntZneOexbvyVl2pj5dlCHGDeaKU/EgnEDZXv6v0xB1RTr4q5vhUir2DNvN9d9x90fIz5hSX6m
gjGOw3DimR93o4aueh5+lI9SJXhiBEg447fpg+XTJ+jo+52lBSa46clKLxRY0w9/Gzp5FzjikK9l
NcJO09Lbl3+xLyDqS/qFANOgSzHaV3TJVH/4LjFXrlmRhp/J09a2hy0t3aUNUjillHzD0433V2cB
8+Ozdjcp89+/mFhIhDDmFRYxXAJOZeaxSzF8w9EJTDpmKWQCxOGDpFkNAGHL7qrf8SwAMrH0zfDb
y94DKX9Z9MxdODo6mY5PGVTaNQDXflHVRWAlYYPXCOwUOeLxVwT3oaNllxggywMan9zSwtzQ8/fK
ejWGRqt0IjwHZlxuNZU//fp/1v+2AlU6mvNbt1XYrnbLOXgWXuY3X8SLbx3hpyGULfd/4xrsibSB
gQ023GXz65pNo7p45M+PeoLW99lg7/TpkVusYE5Ci9pdX+aLtuM8mlUMziyY5CfiANwYgTQ7SSJ/
YYdLt1YnkwjeIGLPSp8rlaDKgI6enqAESqcUBcQNRHleWcpCCjPDlOMdYNseWEN/FcmvGrQsuApi
j6DTJis0QVmjcgX2Ya9th36nK3mYjWl/U9wEuEtqMybfNVYymU4vTVpS5uUYgT/c3XLwayHyakg1
1IGbdEVsvlzXe+ieP8FCJMrMLTYmg0/n/ybKoGjgKu4oPjZjSVQL8WvFVIX9vKg+N+FZpaiDa5s9
Y2YNwV800LOr9HArPRuZJhw5LGjDpZ4c2wZhfrcVXtsqO3VPBCkcbj986KyQuU1B0JIUJfNZxDuD
Fu3xYpuCTwKFqTg2HfKHFVjSRXryGxPoWsUbDMQECUtxBltMzEZmzldz2amd9TyJG0L6PjdsBvn6
ZtRQxy9VD88lUJX0sqONCjXofCT95jCx1zdSxDiwiyklFjmsicyp0PuMFzzeSa/OeplCAlOxHajT
q9BbDSsKurlF/4opJ0FuvjxX0FSKTasvI8DS6aCZ7hBqGOgaacCS1tlQcPAxlN36NwM8HyFAbuo2
sLkkn7ITj4CNlfaM1hgFhgs48/j6aXiaSnIeVVc7Tz2JGHxaWL5HJuesEx0yTOUFS38eIZ4R9DOw
bn1CpTJixEY6eVC/u5fAbAsUx2RUKltOlI+618rh5zunE3dibTzPbL65CUAGx07YrpQccFc5Adkp
isN7I2sQjwA5Q0EmmLQosFHHdU+/Y/pLKkle8v7MP1R++VwF6QfxU/1OAppYDHqNYXy18x5jsbc/
dPeQU0J1AwOhem5waBPuonid8ZXps2xH7CVijt0gJVag1AaOfmodeRJVC5FtE02N0iOFjF9KM9VQ
fr0nwLDpHByWuoMVLnlsovk0Q6xRJqBJbhBOYvZem0t3yS3nkHKvwgc5N5lUVSUYFmEcM/nBD5fH
xxuDlN+NoHkyWib+NznPO+H4wcOWfi4deA/j7Uk0x81u8HISfTwIZ/z/BSFr8qXljswBCZj/8unI
NeCnLAhrUHLYSsl9tCErS8Hqqz9I8IlsdCS0D59at4kp4Rl48oVK/eZwPAz8j8yUHIh07Sf1RlB3
HL5qCtd1NqVW8o9MA0iYa9pHg0pfuQGTIqudLuKebk5QDrTiow5RDnZarsgYR/HIgXmahLin29bL
N47Tx0g1YIVHzqxWM/tT4x4PXvsrVjMIObqAGoWVYoN6Jf6ehf8JS9cZI3Bc8xYvw3xpoKDm5X1P
7qTKy09Ngs+czbbfGhGHQXYJrDM8dbKnKAjXFSs6Ie2SF7+uythp6qMxuT8Hh+yIlWmNal6nyOnI
T5Wrh5ZGnBd0yLyfkzCkyoxMoelAsejL/a8tmzpUpMfIMvUZMaLjcj+HUlGaQLrjdag+iBK0D8xF
1gZ5ugYHWNlrb01/9SKr/AqdFiAGZssHS1RSYgBdGHepHbG1UPEBQplnfQvnLz3Jc2bsC+eIdz38
A74CK+/Qfla2c1cyR+DCNy9gkG7MkysP+71eyhPmg8R0MqQC1cN0FPDIBpFa+FKtYGOgcWZ8HxTM
aImpgQuvXpCLLSZtIUfpsm0IYApOasF0x0g3cVP3o1iKG6X0cHNOSRvSc3giNIBIwC23ZfeXJGWA
H7U4v4KRRMKvrn8PTStNGO95WuS6m2EogYryjrKctoCOlBxEXZHYAUzSaUkCZcyfNuELQitRV9qw
J16FBf+mn/zXYS55oRhlAZn0WHigUsFUlGAh/tiSclLyIS9aMbmziolc+MDPa7aFUDmPfGWrURvH
ChSsh2VYdBC0u+qQR3zBjiIeCl/U75fbfuA471tnQYMNITUydm12Hl337/wikjLeyfa3Oo3RGLGr
smzqbKIQManyi2E3XZXEEtD425Z2y925E3/Ft9QRrFMJun1mJ4jwqhb0gpRd/rAWySW+sSgRoP8r
3tR4clD4bF3SPYZN0ynP5XK1xDdN8zkdcztmdztX0VMbQHUlp/kB/OLaXFgUERvKA+rMwnNq5to8
BFLYGkURiM1t7IHmXKwkooSiB32qGw71Nv35/fFWEBA6sMjluP+zf1CS5O/w6gJGldMKAh9nG6w9
YVkTLtC3MG8odIWeSdsqjwxrmiD/UmUz9RoVIMH4KdUqLgzjp44tYuPjWH1CSkyw9zTrvDWGITt2
btFkLUKwkrS+lsEq49j2OJLIp6Yb9Taf20nWDMVZx4Debu5adc8xh4JKv7Xbfp6EVurFupxQ02Hu
zItM2nm+nFms5zUnzugDB3+Mx3zURPWw3L+jqBPMhi1oErNwGgNvkj+wz/s49UfPV0OWGDni1JUC
MrG5+uoLaA+cIpVWe4r11Ji/B8to9EHOpr3sNy+DR97ayv59tOtKE9HmtSoJfdzOFJA23IrddTCE
1Cai2SnACzlGkLMmLhdgjGHvLhmDToIhCiGKn+9uAy5y93nHqdA8D1bEaMAV1QEmnUhnWXtfzUkS
skJ0Gv8ZAddF4mKGUcUNfLpSqByMd54MBifZGN1qQ3OEF0NJ/Y/PinmRUzWkvjX27hKejv3hfXNU
I5jRYwOcHQXUPKImDwU8+G6nHctd+rMkpt0Vj0PW/yYSaqVqti/ngk4nCIavzsehhu2mSqLACO2H
5tEQ4f+5FVYZnsRBGBYGo6edxvoZwcebIxg+Tzs8RzscuSIFoEmaU8Rkv1kjsnIoisVAJmkNQBIN
UmO91kZ6k++UlO0Jx/Eh0V2lS2zJxNsTms7F1AHRgm51fCtVUjMoKQK2zH+mOtXZErLGNdinX5y9
n561rxjTORpxoqIFxqKbtw6wJNo8zd8z7/CQn2jkMf3nfXQGJrAHhqui52prVVptxuwYAkK3dz94
omiYicWUDmYtsMi+oH09ZgRzAm2HBXKN296tA5n6rtctuHPTYJM6CzhIoGHPrLeWqWWJJvT9Rjkh
UjFH1QaF4qgB3WxSiYAdL/q9qUQE/G3rnziwNWvLCJOVvBBC8aYylRd1J4W2KJzVEQQ+sIXkMIZA
fwW0UH9h1423EvvnoYjgL6r42iqQLXKV3sNufXUyHDl3w3gR76DRE0sVaTN+BSgvJfxe9cYbXZZz
4rHx7D6a+SUvneih2VErqcgK03UuHHz/st/NCtTL+bUf3j4AjcM/kDsUahMuLo54lAKLTRUVENSN
rm2YcQM2e4lNyz+DeOh1juYJuoCJ5Jtb1a5DjzS39UJ81az4yr3pYUZmFvuv2YB2XLJ69hy9AsAl
N1JGmsKwCeX5szMKhJNxr/vpkY3/7S5ExspftzKr4lmkIMlUnouCEoUGzMjpQ8zXoQoEB+EmdGal
2kep7zrRcYulR5mEv6tW+QrNxBOs35NC2oPpuqwvZhfE7sbNXwvCt6iCIJnF1a0USOVwglBIcoxw
q8Geeuy4YIMi4O7/WHk0/VrgwLyEsO3DDtdFC/qvmQz7tgPIllt0XUcPFfV/P0FB11il6J68wn2S
T1Dpigej+rRoUfesobNoQNCYwc6a82GtiYT3sOVcKRH0HLd3KFKhwQUc5lBX1ZOkVgkeXpf6raEs
o2YZPWsFF24DQLAh5Wj7wLe5nfHQgUdmsnUYZ714t+BHHuA8JUBCOf9mDJtctN2KLdDUGKszzqkP
o3IEpCwVAeFg5dVu5w06BSh7Ge8bszYoGhjjPlcu8sUAm1ufHFzgsK5inGNvcgIikd+a+HLG0duJ
sSYABP0ARvO/2pdUBi7yix/C5TIoAczaLxSKJYe2OHWE9sp2MwVrFLZnSwNVUkuBRPECFCHWrPD4
LBQkd4SJ+2LDNjIdgre/L4AJu9bIM/J7EkMNTNVV7D0QbzQsULIkdYaBG0qsX+tZGfAZgEM4t8pc
oz2vbdSstELq54Csolw/xcsp+l7vT1JzVUVEG+MO5OtKlykcMwzhC5PHj45i17Bv5T/3TxV9nqim
kyu+wEENCy/kPJDKFv5yzRZ7E86CLxiDCM7czG56QGmEUPXhxEcx6wc8vO2ppnzNkj5DhF3dbYuR
Y3scLgZb29fFk6wck48XIc4CkNL5trL6iFy2LySQMPSpn6wmxAl6RospAxHdOPNOtVzc0odyxetf
3OoQ+EQ3ZwvwQEPH+htQo7VsJ9TNU7vgHp7wEE2xXEG9tpZrOwQgOolQF0dxrKkKJxcUemOiYbSA
qAXMlmKtBmqyMrjx0te0RcKrv8qF4woiO4TxJEKBWdC3r/Tq4azcdjYkrGU5mhu1fI6BbPDNKrdW
IMmm8naNUIsy1b9UsVcsaHQfwWUO5aYrq/ZZ9p3UOQ71arIde4oGgTT0LYZe7pFY4qwO+W/HoZTB
a5FJSPSF72hGSa/IxdQy+rvgyxn03DM4J6+zEv310IJzgnhj/8njdMIfmmVhPdNH/Lq6Pqzxam57
QRWXiKPOOSjGvIjvJI1C+tEwAM/4QOSCgkFRxbhz0poIL7tQyHQUHuUEEnJQxcZoux0fSxkpHIh/
5+56OLtTo/+fBL5u3+3uzQlXL+0B2DmZaEtWysqurxyTbtATzwl+6f5oTZfjvAWXFlE1i/HMUq2B
uOfQ8JiP+k0j4bw2O+dUGmslUUME/5ikbIrbIaoqyzRiItGKgm/gBEHmmDb2EuWk2Qm5M5nV3zJy
PN+6luUdljttxWh7p3rfWztIX0Whmjh5amWzy0h1+kcjM8sXAifQv8SKZjQFSskWFfEyO53Lp2K+
3Fx87hcOQlf05A9g1hGyVoid+vWurVd8CssmwB6CaZk9HplqOENroE6LNl7P/RkdfkUjvjar2pYD
JeWIxAdrk64QYImFL775nXONjNJFVOAdsBSdmforeyRF8ads47K7wTPpzDRamMu29vnCC3tKb+/g
E3a+N2EKMtBgRjt74vGJfHVZmXYzaK/OT/W3jOugeUvOzjWTLX0DNDp0oLmcLaL7ds4pkFCBALKn
gkgBsOrt73frAdBw/6uHv/8m5UHbymGHyNEheD4ozeGQxfke8lr0ue6s4N0UeY/SG+miJRobAJLb
5SdGhKvvoU5Lj7/wn92w3v4zo4BMyULYeVe9ck2LTNL+tmjfynJcIpcPgZIZqNIEvysZ6fQ++uTa
A4y18eM3tXl4hHK+WUvhSYIWYNVPid54y8yBCD+JB8W3D1/2oy8ZtFnMRLESGw61DJkhDZBILlHE
QKVfJLO+z0wOFN/km/fyxHx2KWEirOK3dtop4o1HSEYL1XDubeK+k1XXFDS4c5OJn6XssMzEyWzB
vYWOUMjFAj9gc+8xvisAaVQQTS8mafX0sQ/1KVN4ACAIfSNQs/CIpP7VXrgzFwpyp6rbT0mds1+u
s/Hb5jVo+Yqc+BkvJo7Ry+oPZEPSow1IlBaGSXQnno0OyQxGDOrnzn3u+BbvGcMRTvqCQK6HKyfm
1wzFizt3hcrFv45ybHz6lbsgDxUn2ZoNU5A0AXY49muKXobslbZ3HntJv+Gk1YDQLnPKPADuTVbp
ADOesYH7zN+dJxKk70YQKrcUOt1QmwLqojQgaPTHBCJpGRa0yS6v9Wi4aqkeY5vLwleyRIc1AlXW
v0mLTQu3Tzvti3zn4eR9IC8LJ5EC851RTpxE1thxmfL2ju5YfzTPhngLdSjjZu8DAcpZwBWZBYwa
dUV6YxKNvuYEI06x45/4pR7arZj24GUyRwyuigOjA4CyJaKWaGgvNRehiDlGqKxIo6pwC66hjYBe
VqJGvRERjs17PJa7F21yRmXoAIZigOMGoLb8HsL0VLDoCTDwWkNj6IpZhxjuTSfmAHKadL9PfJPD
U4s5ipBJuCc/5qciN9W/KXgucs2X+KIvdidYY6Bv44JJoxh7U3dw1bqMSK0gaOiOiFQF6fE/Kcxo
lU9C/CLgawJEUkXtGE9L9V5qODqMEC0TZ50423mdSz5/1YXYs6qHDqgZrWBZCAfEoEsfJ0Ee7EzY
PJpFYt1yqJ6IRtU+3rYnI7IExjRvNHr4n/hqs07DHVmx5uVz6Z4nTiiJqRWW8lRK03csOPJwqiVk
1k6osnKxocd4CQHoXD5c2tGqfhZg1duxQtzvO3hsjZrw20HxnDxEUYIkrKGs61/yVQoY0PiRHhcg
OTHZFsgdCouA8TK3nPpR1mwNnYaF5YmA1Gz5dwMDxCAfcrwu/lEykNoZtTH07qDIPtxOLOtWhxNH
2utFs986xZG1UMBMMlti/QdNR3WYwuQCFxhQbQYIVNSGdzAZ3c5b7PqJc7emtLu7ky30FrBydJ+H
NGEzxIwY4J2LEsIk55uiWqxv+eIyDMXio/gq+ZsrUsvpM9ZX8yCNdJJqH11HfyEzCxYEJ1dt6S/4
hi/B+pTJwEd6G13sTSf6UjNNRokle2wO8IaQiZuQPDFOCU8QIISrA6JYd++avzOL3zUbnjq4xnSB
pIF6xfgpCki9Xj7SmDSV2sngT1H6zfbo8XjSAkouOVtGx8F8PbOzzbp9hR5ZPnMTONSXlx6Zg5tZ
cObY3zay+rBBiZTWybAzH0WP+Cij9PkzKhwAGsAjvXSSLkZrRKHfQVbOGJGy6FcQa7YgMMS8W59o
xLyOW+bEPheTuSO92Tu6voG+Ngy2lSs/st/+yhldhKNvWypqZZ1IBE33DcvUAed+Ouucar/hNSn5
rGng03qaypt0DKTPml5lbL3vTdzjuwzrpD7zCd5tW+behWlwT2iUxxGSdTt+mB4eT2tnD7SgAKXm
95EjGmWdEpeazOgHkYeakjepKGuZ2Ms8otqdzG0GOEcMGssF8r2SFFPLujDEC8YCSA69/mXlsHiV
WpDEUndjtDQanORppe50ZpRpUwE1BVW7LNx0zkUH1uyG/sZ6jCWnLFKf5Zg7Q/QHlczxac99veDV
H2O+ctrV5OtifEFfgaPByD2NeouwjZRddetAg0vRTMLZn+sAkG4rpkCq/MFYKG/k9Uu+zhFZUQkN
ClQfRnYK1kSYCtJ1dtJeolnIXQ7YUSyo4eFLenBrzmHiAyvRpVD79WpEZOUJNHT9IU+6iCoD74l9
AVLcec5bz1mg7+El58jAXpCpdeYnzjR1Md4EOpUDcmEfi4cOIj3NQuRWyot6p5VfdNjKyGAjl3rw
jx6zKhETaNfW8DO+NZqYwKaic0lPabXGNmfC0thUNKB1IcXhLByWcMKD9OSj6EyCq7muscMqGycB
hJJTXcQG3I1vsUnygFp0oiS6zhc2iel9wNJaNFu1Ttc3RfxpXh3PKW3cQ28gW0f5ludQRd+d+XhP
SvdmYcJNxUhpnkl8L1qX+UDUEuYmQtG5ww/RzqQUp++0lYxBf/CJVVEQKYcQMrNoz0Gad/983ZVF
bTVDcv33bhmlRRv3Lk1yce5DoZANFYvi/re/Uy15wsQCLoMBBLWzpBKMy3CouHk6YDVrSVy2lqsI
f340NcTXTeSG8epS6qSVCI/mLgWsKY56vDJJBC+WDNXNJITtMOCopMWTo6omDW0C83RnpA0yuCfV
fciEsiP7YGkR04fn/1ny0uUl6pQNq7vBmlyhr1m9T8zFpU2yVzTqlr1cc7wf+5jRHzmZ9jgPkrFR
tIInVudsd5tOteWJOsQWqDrqyTeaA10rtArwuj199Rr+SoVNNHNCFEhj5j/jl9tgknuZXrBiMTkR
pgyKZ3BgG0VkCDervY815NV6x1Fp/v3yvp9Dv1emYDOtPr/lESMgJP+ri6APK/Vw1V31S8/S4ror
sbSPTLmi4303O8tL9tTw17a1kVxQekfLNZSbNz9xxMZHkKPbVTEDdoeK/5L0Pdm+23UAS12nxnXW
r0wvxLlB2LRxG5tWoSYjXKAlf3ajudJw8oYahVQjW8Ue/mF1pHzuhljBQVhWquliyued2fJLqWZ3
jF3dLmjjrsUF9iOr6Ol3YYbWtYbOyh9xzouTDpY/7525/3mPgRCnQApVVEjlDiHZDpVmvSRVELsW
OlLW9xYVjtpeSpz3viaPO0XTjhXXqJeomw4jfEPpIpr3Cz7iNEnuaHkA38sMhydV4+w3SsjVLD9Q
VFaPz22Bo1tcHKrWs20DXyPowxeQfA6u4Up0Q3E3CY8q/atlcpPAd9TSXV63c9bBfob6svcFf1V1
dzzto03UpTFHqQzhst3c+VS7AFRmHhih74FVyKGBtRxnprb3L600kTItPzaUU9xWpYhvjZGpwyYE
/bWPoIZuJWb7mCfnsE445cjVLhKiLBx5Szx8cWuwEApkvx1kBItrWLuLyVFKK1UKzprNNCMQepFF
oSl+ap+MDN8VSz1WGOMBehm1TNUWiSphHX/dcb8CmUTI46ulTPKCncrHORwitE2AxotVL+tHNGIX
0DwXNKV46Gs9St+IZG9sT0rL7IZvQYRbF/ta49eULd1/G/clIVDhbe/QM0OjkPEekMWEAg3H063Z
IeQFr5bCw7J560J8bq2hCDbm/Uco9QoYZI0K4lgl+q5frMKFBPspcZ4KeQq/s3GSaz3uPi1W4zgF
DbGFbC3esh+nttn2ZegQzT8e3pdor2vC8sI73z9xrzkz77Pp514jUcdhoVUCJb8sPEfhbAeAbDAw
yH2nwOXkOG04EUKuULry45tMdVr28e99ePiorvy0TSB1qPrmhKsGbIPZG6yZD+JKkVRYdOEOpPTz
IYDb2Db8tJ/EedCKXur9zrbtu/FkfuoZQjBbwjvJjQy9j1Wq/y574qHvSEmx4aOLfKBANjvi1TNL
IH1wlQzIyJ+d8IO4Lqgon1GstEFQ7+6H0+69Ys3gxgu5sx9f7r0EWeTWjRLmQi5pZ4YYlB2Y+QAu
8Gvdj8cST5sS0eS522cQMtOZE7pnVMvP+IiQ/+MZVN0pM8HzFEyxpIaqWS6M45zYEwaCcrzLyKeq
nh2l2yAgA7J/oQBdBJHu4mh5r/p9Nl2MGMG90YH10ha/1eUjwM67WIUeM5gOCBDEJqsXaSafjTDc
WmiPlwkBsq0vsVyQMTJRoHAkGJatjykG+CbePyYzs/fUkYdyoz5r/710RAArkWFYEyi5RsXx+tHn
TpNItHJtf4TnELBz6el/nGm5AxR3WV8OhSwG0pYcyEC5X+etolBqrdm25EDwq3TOdr1Ndlvc1kYT
73fm469bnHdBLmgf/+LWnqAKltvSyzgjGFSkLUPhjs6h4zR469M7s55Bx8MfVP9WlBnwMYV54p8E
Vc9c5VSyN4fIrqby/LS9YZuH5YntEdry6fo+nnQnvhpMB20FlEsed2CQGe5ltsdNNvLiWF5bEuNS
6UoI1EYW40uPsxmW86uRLAXmd9OHVeOgos7V/QfDUmYRgkeGgSCngnsO+GUha0y4D+9X7zTaTNLN
KwVGrbJf/R+Fa/XKr4Pcszqw2B1bfaHxlV5LTVQoMrPSmN23wjSgQRBB00mlXNHn2CX7zxukmJ5v
QZRSzLdVSbhwYnHff95LNk00GS5I7gH3ygLPK7OhyUssFedHCm6+8net/p4sNA/3sLc5c8BmE29J
VVpZOhCNrUHCIGeNdvaOED7Ldjeh4sQaS2TTj89CHfUJRCFKlwsUpLYUSZmO0j4SdEEgC1OVec62
f/bXO7BFr+eU4/L4OUjiubipfDnMv+dKNPfd8QpMu9N4Hdbm5mIIHKj6XHMUtleDAf/cXpI8B2/s
iWUiq8XO+2ol9bzcnIvvZNm83I+zA6eVs6FQvmeSva9FhY14R0CJTLcxi8Mijrl5He+ftupE1yyI
mPNdYOSSootKuS6wHIxb8enJbmdC7GgmBdKzLmtPYdu70CbtfNR9UQYLc7a1fAbMjxUpmBoDBJfR
LbLCMMb87cAZvVzHMNfbI29TF6KqS1DV8E18luw+3bhYkvlgTwyHc+/o9mJFq+UKQar1w7L2QXb5
29se/92uNObfmlGjcsdpVLDhMuPRMc9XP2FAnJ5RvpE6XIUdGs5WYK0oQ3fMjFpcbsw7KZ+iJEgp
93LdEdU9JTT3ngpWtYFihiopVXin5ZZkjHYuyN9x81AQfKusgq6l+MkpyZu/RgEBzH8YfWbpO/RD
fu9KxvSupta8C4/vg9/CcLX09dL/NL+5U3iNDaVxoMs1h9PJuPh63JPutq1fxdFyMF96sVgnFsHh
cGaqVYOlNWRkrvagYKMnCei+toBNxK6iIFbYNfUrU1bsdDvNCib1sbE6JwG40IPEF/3Fo4ppOH3x
RNtPm4iwhRAFqejhIwi8za6VGeJ7Q3HbSb94ZQ7W8GNLK3wv9I1C++3eUNg0rghzfAnM+J3h07L1
a+1EHlL5a10V9UPSSfP2qPyUZPTPWSHl3UoUqOqAMBF7fTRzzg+rQjjLhtWP2Ya/m032QSr/rFqE
p0EvtyKbtsOFYX4F0rehniEZmEt5LJIgLnNG71YS5gsG6WTHyw+xGGQzHwcqXd+MjgURxO8cztOQ
VQZR6CjBwi8OE/kVqjRw5v+ervSg6XPkF2t1FWW3cjwS1grpNaosBZrzti8aZTtENop71Fha0spF
PDPDkzM0+n8TEfssCuRyYWdcadBm3eYxqNS8gRpVpu3eqOEy2erckEE3oksn6ZtImBPDyG8blFGW
7zW7eYDo+jpT3WTpFgFy0rMAZCTFDlMtHj/pj3gEUdleEwk9dajLLIUE4DuAxZByWGrWbjRadYrF
bdSDbd2PZxAacKF4Q0QZzWaVKNJb1hxmYvmlT6r7OwAPqqviUQYlrVEBsWNR/lYWC8ZmyJCj/UBg
lAvqdzvM9hz2KATn/NLrKg6lhoclEOFcepvauMCejFN/cl81/XO1sH8VCqXlhCGnvmn8G4I6fXLG
33npv9yb8naO7mMyhjio3SS6wyANqRKgnQFAV60dv4S1mHpDWkTnN43gEPnn9eTUMGcOChM+qLi3
+Cj6wcqIzjzoY6wPozPhKeSaOxrilZGz9fEONvm7V6LcWhxzE5EDZRZ65yIBkYr0wItu2mJgBc2Y
ESvROVvcpqUoQut99aIR6Lki1Ygc+hLHa9tDTj14Cr900BLaL/zMDrwNtu9hRBAwF8AXpJcetOhK
8glynePwmiTmXxxCOWkQfKDNAHm9xnRZ6AOgRBDu7Qe3Y7FJgrdjjVuRjlLzK9hO3gs/gsD/X8Ub
gR+ZU8x3MAPPKXkI4r4YM3cFlqKycQ9iqb+hVMIyeKqREF/broibv+jnEmn70sHsn2sFDak7ukHC
6WjTZvvWspS+LSL0Row3LcIITPdsuUt2oy4iihoyo6vlVKQ9BwFgBnxwRPuC9KxOCnWrSVEaOWkT
qM0Ah6zpFgds7un+LArcTiYFoT/hBhqktvnXyn3LipFgYgWfTanjZSeo9OyIxY6EglCXn8A2Yl1u
gexqlU8Jnf3W077ZasJBqQjuOC+HhmlpW/u+dsRp+hPROh47ZH6ujEpthTXAYjRVOZd0wbEkwyNo
EhqCpejYzGSG4eJYxkcLQ78PAlSPaYbB3Z1pbVMfw78zSvXPbwjO7tUhLUvOBACdzk3iEfOZ6ekU
tptlJTZM6Avul2KZ1D2hQaMfZof1LxdktO1hhMpDqD0l/IWoV9GXFBgNUD/yeRxfesYBGH3elowY
10Ig0K0aYNjmH8eVNlRld1/OrNLSYbxUne7xoueBt0JdUFPJ+NoaqNiI0xa/cExFKjEwyf+eJ8pY
Yo4u0hZQflIUZYj3fwWM4aET06NKccUq/tX2V2TepUZdytAMuffyH66SGVFuWgbQP2ieYZtTU+T8
DRf4MpF2bKkDN35MTuG/611hWqHdfRRVPt5QDiIFyVc6I+1t4cX/jHhogrGgMOonZrfw5qiwe1x9
6TPSNa1kUKPHgHZDp94G6dNUtjCpdIJW+0q3EXGLsp/2wVRVxhl02axxZ+MEh/TMyyg+198CwWpr
zMkZZ6yoU2sRl5I9iZfhBN0ZxgCbJ3R58+wKz/0NtWKlu/pFAB8afIOw8Rg3zb7hEaVTGs/GTRZ8
bIMF1YLllUCvGUlCSEs0DPIRHJesslp2Y7qCxMbOBhtcg3Cg/VPiAHroF4L1XcN+Ps3eVangrW2C
X4y3camYOVJ0pyc1jSxBTdIrYNP714A5YOfnieqtzV4xX27JCcE5uBZtxO6gwsdYLr7Xscwqn7g4
CpQdPd+uuzSCz7vlUSPit8S/oaIvrvRzfTRyVmgBJsObJoUkwEK9Z9H2dZ7tU2uywNlW+crvVJcY
umqvs+NgHg3fbWzZbq72o4SwuVTZKgCVWfBI1q3SRDCoMC7rjrsofvZ310vtu8Z9hHtiG0Y9yfJw
YaMNj4Aoedblqo9PQ/6zH8PT/6rAEc9LshMIMk0wOMNDMCjatfOkoAilYx9QYxk8QV/moZOorBhG
C67CfAuQ0b8fJvFaPDqiZHFPcFj+n7v1yZuVvNlo456ng1xILHY/QmB+wKXc5yMag4S6++oY8zAD
u4rGROMuebtWyAOS4LCRiTknVqVEmR9YaY0SyZ7T09P5s8sLeAabImPz0AhZntzcKM9lqKpMaF5t
8BFijCYsVHFvfsKAzXS/5RzzgMYo9rbyicJLye29zeaE4lNEeOPXCsjF4mQKg37MM0k7pQmf7t9d
wzeEt/4afuEv9LxU4q3hjLjfVEnxa6D/tWAdjzRATJfNtp8dx5d6nLMGhMmp1elou8cibn8IVBYf
KWN43Aiq2XPpb1ZteNPUVrmFMX28Xo28uFZpuaushr6t18DrN3+O1KbX5Xr5OoET0vI69/SzqFvb
eU4JT4UdOp1Pqw+dTV/d/HfyvWfVhlXQUCcRYu35+1uZAzHenRbDCNroXGdMSVjn343pX2vZ3zGY
sV0+2BJa3TLZw5Bb34GTGPMT6NSMuh0weiCUv3uHvwYAt72oJJUyHkalOnSgX67X2CdBFkQwAaxe
s8viLl05fwce8AlyjF84RE5wKmmvHpIar49fv9fB2lp93kRDC2atA+bfe+SPKX3juzNOEXFXiHzQ
q5bm5WP5Ne8PD0DEv+X5SZ15+LsLP4CqV3pfQJ58esc/FhqIZRwgrCXjw6Btv91uXOYK6HpVW2l+
B4hWDYDXBQzCnfB+NcBseoQAFn2ZBHCKF+nouvA0Th4QkToEXjOBb8aDqgQVK/0Fv6tRsgC2B6Vn
rodpwWH01AzQSOBtnh68K6a14jbfQN5rIzYnKWBd+vQKcn0OfXAIzxB0N60fk1qxegMe9DdLMsXq
qiKmIQIL1sz9ztqC+WoXxHLKI21Y5KF8f0cyJrD6IipU6UF2CbNEe5oADknHQcOM42tH1ZPsRZo1
ItGL7DYkLSVuXlP2thFPIyf3Efp+KUSxKDEOlLXitskOU+Izh0G0wSmr4WQjBl83oXnk+mdBpiqb
DXyzgyCFrqeQi4ckIAQ4VIAkkjE1VRIyysia36BZFufgHL1JOm3iFR3a0mOyWa7kqgsge0OjaTXo
gsBBQwRzmQIJnbYssbSwruHx6nT/FXUXSGXxbTPgcPyFTJfmrLmk4lZnHnjNd+baYe2poDLXDxrg
XBGj9n0Wa6PqYUJeTpPjzeaL+tyNO/bmdc7VQ/Y+3+TQoUmllD3Y0zIfP8MnegEiLf8zhE5RQBjn
zAdWQKJuFCH71ARRJGCMTdpqgW8WZH651Vthln5igZ0zqv74bYOmJLBwBmVpFYJUm+6wNox/mD/j
YikkjA5cranGkVg6+S2kSg85heSGDyyg2NVB28gACofMiXVle2Hesm9sNivEPMnHjDFnrciLLtCf
baP7/lO4HImHgAS8lLgHvHatzktdaMIRwQEdz6jVwxIAqlUbnA6IZWjEXilWCfY1Cka22Q8TSINL
7oy+qCcljM1OYQlDvZAeXI05Y9MTvKngsH1D5NU6Aopc1zwPcue7CEfYmHlHFB1B3ioeJnZAD5vP
2dwpeWAHqZT89QU63N5/gN6Eo8G9hHP8SDb8bLspWZzqHOS4pZA29l9jIDqdwmECn3FxJYkB7XxP
bRO5wsY4tVdbwIjWtF4+1UIV+g0zZtxFP/ZebZ6VBQHWU4dIL2RKu7SQ1647B+rUJxVVmptSELW/
YvwtmJgRgpFpGepipb36J+yeyIFoZwkiHwHq7ICciU9ULRAoKfecqZ7ruxEfMLVNepNiao+k9xQ7
gXauuUiy7sFeoUcmZaU3N4upZKqM4x22/av7u9B7K3b45tNlhiqYqEHcoBOprqn0HfjoEicGf0CQ
r6ZIyDjnD5lL/P0Q+MqFy4EP1+kNwg1+bY4JEOGz0W30VbPqyb+imcRZk58hFUB0q0d+/pUDAPmF
q78wmadVyJXqUUYPztJ325GAC87ZnLA9oNXauSWNJstIDcSua7Krla+4WKsZY79/1pZ1H/yW/PFk
687bj8LFPTB85lPHHQbhv885/8kGwNpgAr7+6IsWqWQC3hDnB2QZjIkrtQ2HGvDHlzN/5c427DAC
RxD+x9Bw+KHJsCUoYOOf3oQFxd1x+ODFkk+s/tQwFJFNZmLkzkgGz3sQ1ErSgU/2wdwWAZEJDJlq
zh2L8YfyDcHcePTR4Q3GXtrHzbq5OAPFG+vh4a2aOLO1P47xD+9HG2BzsDkBJVuXTxidtdPIXj8r
I0E7WDyz8+rWgSXtkf+AksROo0uTHdm1PyR2nehJbOSgZ1wqii2TboZ45gaYUlBgIeljDLwJMNT5
OAH4pI5L1sRJqR7IKXHKmE1onpWDbRb3R8rRaryH0JwJkWRYBVx67kVbuOzFlgWkwAtNj97mnRSQ
OpNlY89SKlucZdpzSi/mww7WUSr19Eg2iodXCh3z8XTCh3af0mQ8Et337K+C2J+0Jdrb0a+/3jFh
gLqlP//XTGSemLfABLI7UA0WmC+gmHUUs+kY2l2yHhZoW1hJ9/hzGquk0Q9sURnSvn56PXCTmMjm
r0EA+4IXwo5IDj+167P0H/RfvcFah3DcuWWBgnNy2zjQ3kpATo1HTwpZPfoIg0Dh8VmW0D1CAMVC
SawfanaRUSzlzV8XK3uoBh+NADX4nJdKUJfEbpL51jCahMZLjiqeBgAvv2MQSp+TKbhoSLEC9ZK5
iLqWzhXFD7ESbyq3uoojL7TCmrE84c2cinvPMdx30gUcMgp1szDSebhkhvz0eKe35kUVLDJNjPm+
0EdGmlvUElULD87pDMWifI5k1gaCN3pN3oJf30XGpHjWRgO0IskuUn3uuc3SfyAoGMf0DyY5TMvR
GgknJaZoxLojDQ25kC5AXS5HBQJrXDlJCyQicEQhfE2P2PiP+r6fqSv/l5L5sTmZkypKszTEkvCR
Y0aSBDMgO6wHpk185+J08EP6nWbiDIlZNN01sG4Pc9RdPjjIcAvHUB3DZ9NLJT6tYcKtGqTIQVOu
5nzhkgYPX5pRQBrI+UMhG+vtnDVkjZSu1SdQBem1rtD3Y1mBeYxlAzDPw+ARj4lDosH8vDW+5O+V
s7kBYGu13JsvoOrqNqMNcMk5JywlacMoDQnCBlo570ams5V5Zldwwz7LZ3/4NklrWRfpJbAmWIFu
KnsOxFvj3aZfErbkNWG6pqV8KkKstJk8vYsJVlKbw8pP1NvHvBYrCpYlpU8bPZUbxctN3hUz59WY
eIQNsfu98gfr8ZogXJ0ADqSg4ejLYs66x2LjDKuf06MZ75TcS9GI8OAiiliTwPRPs7B/BKOtVyWY
j9YgS4lO/I7z9o62ASeBESM8wCTBgMXNVY+IxD5Er5of/BOWd+PdF/UGoykw5eeRtAvcYx4X3bAA
itOiPtn3j73sZOOvkIIFQEPMDDN0KkwMNI8a1XXhSyj1BSst6tAWtODiYBJGhXkSP0Y1cNxxvSfW
pphu3XeLrO5R36EzI8bWEOsvoIZRO/0uQdXh9VQW/N2KiC0j1dS3KO1REA6glKzb7MoPWGiKAVGg
ocsGxmRjrNlkEQO9m5taStnodXeFxqZj+JodX9+jegIX5XdrzKQ9ZKsKpdg7f7M9cVLqGsPOL5wO
9gHlhIHRX8EDfDbDYJ0FFo5zFZBcNGLGF9xHZjZKsmcqXb9Nk4eBoD7Cb9XJAULgwFw6isoUJlVF
IGMsaE+c94m4BJPTGknTgEq/L5GtVrUPsy8SxwdJq28pDsLigveWhEp5W5ci06ejwZv4nvyT5UQz
ehr0bGsyrg9TmqElMOuh+skVLBR4sc3/7568O8lFNfMtIzambNUd5oV1voz95GmXbYuj63mh0s1X
Sbiacxl9mUReZ7AybVbXGhbL7SdBh6v9EC9kN/REVPVCxuKI04LAgu0Q/6FhFziiVbCqPVU7xkyq
XynDhZCZc4cC/H09kMDuqgQTtiIFJnRk39zV9SomlcN+cOlUw7WyenxT8f504ibjoDwem7z6NFCd
qRvHS0WptaGHvmC33I9pxj3hg8fIj6WTlMqMR7rNM1Jh0XQcT4SiJ14x82KRSa6NHDIcZcu35E5t
9ajjFcWj8lbHCgzL6Fsw6OHpGuPjzZWad4I10yVjErShb9Mmusl+CLjzZ5CEQaT0r4FYl+6i7I9q
saCCeRsuGte5ruRICwRBoVRGljQGS/qYJHOvesRUJF+pmexjDe/zijKKi8PQXUAx+AYavwaEGuUz
damrR3vfQl3U4t0TQ33PWcYhLHDIGPCXegPqisfb/KyETxRkJgtsVjZ6JxMOdy9/pzjhS0x9Y9Th
HU6MU9TJknoAlleDqIYmbtmF0mnSM3o96vzCCGbncB31YDcJIWWTvfATrzkCPPAITaWPiLyfljVi
7s1c3I5zt584Vi8s3xRLogXwM08tJYkd5FxXN3DB2NgzAFZh4cyYgyHmnd0takgJ3hhXlvQXinwC
BxWit5ozc11Ni9l5IsWWxveh+gGJgVLhZ/EZBni3/RKsUb43lp3sqYd81GvLaRutWEhzLResoccj
hsozaGADl87x0TnSCv7R0NA+9a52HEAZoRVvsQhUpOX6qXtAiIzsjDyle124hM+1ckTkh25wTzAO
JwD8mJESBB/hEeG61brJJsHelBVRTx9KuGTZqfLa2wJuw7hwYaua2hUtf4c/KRtMg4x0wqaao0lL
LZQ0Sv3mYUJeCXBq2DilFeNIZmNL8d0ATgZc8UEv8aUPhVYH2809qRP9XAaN+AKdVPqL35jpsCsJ
3f6ES56onue8p+Ni4h7mhEu8Xl0o8+a+FMGB/avAWuszmsgIUNYgCMYR4fMEbMIoomeeJiCVCuW5
09xbflNw2EkkxMbziWcxxv8YnJbRWHyRy5ogjyN5If4oTCHL1663ZjdwNrbZxfsBlH/KUWEIR3Gr
E3X8UEKGaeu2/iq3X81lvNLb9iw05dyiqKg3YIc1W5PRjxTsZURMuK2m66KAVZqfVIDLwNCTfrly
7anUP2eR0XWhS47iva1K3uH6ltC4MRPB4oxIq8HONdha1kYsrX7V07FI6nHB/lTEuX3Qfj4U26S+
cZlrw9BfhYMyKPsAKIdSqs7ZzNtc49i6w/OE5f5IaUB2P3Rb7ICwIbXVTHI6bqLWeDyfKC47P/ST
Aqvuxm37pq9Gz2J2mb9svZhH5IiTq767bcqUbkQOIQ16OZ7dhtUfsFVsoX/uaXMxilhyHjPhvhj6
hVZzHnV9BfQJKjOn8k5jA8itOcbSD0QZpUIB26TvbMzPNdUBDsMsihrmo6jJvzoxyN45K4MsaEaE
Br9XdJPuS2dRdWrVwBY4eV/svZJU4MtyaP65gMc7fXUgoGOZuT+lR+Qzz97WXo+t5JAFQ+WJUj2X
oFaTQDmoCzGRFKQw+i8NwpOrmjtPy1d6Hd7F73eqJPya+AoaPANrm+ohFWsm8oQqUkUVvHhW/f0s
Uek5Ls1mJqkkP5cCJWRx8xhM9HbrAwpARuk/7s92nnWcUTAJALpd5u6CWuUzDCPdI9zUDStVNLPl
XOKCOUiecWetKRsDohi6LIZ3RpXmLyrtenRIbjJvTjhWnsu9l9PDVnQSoQ2izkjDenmS2WKjeaG4
X6kegrt0mbUsW8nxWj2VRyRK0HGzUs8YdNbaD/6uh6L2Qfnh+8bAL1Yg/GktLozd++sc3KbtudaH
z+VO3YsA6n+MG6d4fWjrbAJTp5RO4pOcHY1jlzoSq1PUEblOv1mSOuIdhi/8AD70BRUHMo+VL6bt
Hx9XlfDK6LpSDzwmBmm0PSfNbN17pr22UoJwhSpKjc/Zcp+tHatbuhocrf1Ce+1tkkmDJe9hP0PZ
NdtY913P/as5ZxO4XOUrEBX3felkpuH/JlyvGnACBty2v1KJbGrTMAtyXpX6DZ3wInmF2trKLm+L
jqyPBHdfKB9rJhGD4jk/TGS7pkj5rQdopfksrku3qUiNwE4gCWnhwVx5Bx/CVqS/S5nmKC9c5dfN
WX/8a/DpUbCtWbQKGd9ny9h35COH7TrU+E/AlrWjxQIHjE1WDZ/snDf88fIaEJKrDE+VwP4lzOgv
nHUWeBVmWGPeMnUun3767iXJY0IZ88cJZNrUAPUE3WojJwmZ7KLX41r7tYhiNDum8ByoMEWs2eKB
KiEFSY5PaPBAnI55UOEIslngd9nROpfkiNqJqk/+8G5IlK/Vjgzjk0pEa6mFe1rLPgnhK4U/PHe7
oPs+Fz9xHPI47Ge6pquFK6utpE1lGnyJZMUsXiD1Tt+GVTVZ5m4kSGXOyPNNoy6gHSIPvnE0h3SU
MY5LTa6DINFD4dpne+WSTsT8YJCDE004ZzwPmOkhbZTv2F0xhL/R7pWHitKOs+Gm3DAKX7ONyDzD
FbveRPYdGWfAWfYI2gyQLQpS9V5IBQ8RPfQEtz9F1b4w+59sArKwCd2nZWncRnp8skdHnmMVD3dF
clxEoLPgAcClI7WKDxJDQPF7YbPtDMCxmqqKGz0xuM1PBMuAwi2FDqkjmfKShldon0o/4C2Y5sYq
gzb+zi8udDJdHHNyu5BVjq7Ob0v423F0qz6Et0ZuoVQjnEhye0e6vET7jEzyCd9DAR9pgYhPfbev
b+FeNrXddsT2rk5GsKMutZSB/ulex12rSIsyIO2N/CCMFVsrLaUhrv36d2Y9H2Kbjp8ZlzI6lBPC
zZ+JTUfd2l4KbMr8s6LOinw9CTZR7Z/SkykQ+bdTwMxvekOgL8nfCRSTGeys792rikyaTTQP3Ipv
xDxEHZ0rRtpMNuceaeObZ18i6qAbbOjExvTGdepKkpF69Y2fXkV/TnfXHlDGMOlLFtcJL0wfpGVq
jnZi4fCtg5FFYBXnMsWsjzmZRQOEbbeXz8PPyYdzflQO1PaHG4eJ3q+zihzIPReCDbSRttiEg2QK
7nTQsczBpO5QVIb1rubtUdFknIsUGNcg8pMTLiNHIthhm0wgH2j4QZC0PJbYR903rMNH51XLy7Mk
xntVCTP/ah2PvlJCZaZQI831COe06d8zD9Fn+LMDiBWMesxIze9Td0mt4KVa3Q1b5Y+Db6Tpz+eg
YmhusjW2Z4au2ICZwBNtk7ysBwYIt3DMApF4hSeUDSoClCgodf6qN2RT9wXp87yFWeComCJV80PB
6uJk8/GMdFG02+Gfb+kytXXLFF8eKGELl9laHMeT05DgYctk4UrzG/ev6rlc0G4jsYtONPpTCpcz
eCqxvU0SQ2LZUBkGOqZSavYbVEgSpdTozxJ830ppOHeE3BqAvJvjjcEVV8oF6fgLmV75sGHuzd6K
D8Fmoxc0KF8vXzXIapB4Np5z9V16ZxtNsJLj7WD9FmYLYUyPSBuLmPfKB2ZZWOxMlVi7De6rSDw8
WN55xz7tSoOFpDuz8NFq/6Mtw+iQ35YRiK0f9zopTxiIvkdA5HMETfJ0Pl5E6TrvVsJVdAaNEuKh
q6YXAtT3Fjk/Y4Lk2nBCVswu3tnpzpqxG7QWr6npxjzvq83MbYgIiboitnpImhUnCntjKExBAT5K
He2nULV9XBpnmPqVCnrIuxES2BKHwIxMRsBhbYT8qplaJCVScDLNpZJt1j7EAf1/31SIICd8fsZa
QrIg6t9F9IlK7TDjvQ2GWNvu0edH6RVbekEsmRMiwI+axMwn7fBVybTAUO8aFhnM0C/3C2+AmC12
f62kCp6Vu2oieGVzevZ8wHjfo8CoYAmuHxFptV3QZSvtKOHofQpr4MoTZXCtabAuINQy+WoKZS15
1rsMUgQF3MtAm3XvIixLAP8yDHwz9vapaz2POV7EP/1Wq1BWbDwTzOYo5j/irX6X8YG5HF+sVy2a
ZNhdYxy1kq3p9SbBxX2okLC/upjw4tAemJ2a/LyX4JlkbyNKDwT3HB4RnUMkcnCPkHgncY3JNXV1
sGFC2D0e0fJrswJ6qp2Dq6EJFVf+W3I3G4fEy5NHeQdFdc9jqn9YuRlYOzahP86ELO6opiK5L6Ba
OlJ66SfzvyYybI8xETgyzsgOS+17mASyuaGW5Q456760vX5WTIeWaOzAhRmM3Nyqh/QZWmxUgaoI
Neojk/5TRQXBW0leXZUIDgnd8uAz8fRvPu/xRXKQO/lgyYNKReJ+Pcsqg1wQ/W61mM4Ucko1Z2rP
3YkhRYCB5DX4TfFtI7eaRT/EtsoxSGhPv1D7dgrOAcjDXKtuGyphn1za6/UIarq3GrZ9qEjubi+n
LnjlZdV8zGdko8LsOnuMsa5pwJwH2cVYp0sysDVmAUv7L0AiMdFiozSWhE0AXscAyBXXnCwn5DJa
MAmSJJvu7E/8KZBCCizZl1rEt/CjUIpKSnAVcdGcd06J2IBWdd4YZ7OjGATyF6OBqwvx+FDxqSuK
EsnnjfPJC5dMVLymzud++rhAxo+JvDpyFUoytLGw4UnmQ46LXe2xVgvX3rio2q34oHYckWkxWaGX
4gWcrGRSSAymy4DYIQF/z3vVE1nLj9sqNyWLfAFyPAV0mjELKSkQGxEKm5jgE6O+UxvXpLiQPwiZ
T7QAnslbj33+OjE//HWmeMOG7vxiyHHxjMp207ZjLHLdRfJBB/Zwct9pIHIax/mJXwgsX/VIeiYs
QnpqK92bZEGucXGqeHimbRv1UZo2T0mBhTc5nvegSiEPjStxwkog5Qb2fRIOSSIMQ41Cv9ogEgkj
PXD2O0RIDS6z7cZq4A6Pf9cRG5SJMyC/EhOueywydoBuAETTQspbAbvUaTOVG7X5FCT5GgsiHxFP
TjZeIHRfIuC0Va0mAngzPWP0ofBs6sEmgH+yexo0P97cY1naLyNvqmr8RF9HSyxw9QLfwhIZtWw6
OIYb4Ty66oWXcBnmQgFRDm6HE7bqe6sKY7Gb4dXK7nvtsEUH1ZsC/ELEDcM8oB0xqcmQZzhtuH2C
6O71YLy1nGQOlwla+4fypc6eomHwekeInSE2pFlGpEwvnDNAYosMcy9y2hIQZ0JwwKP//WvffcjV
jDcJKPMhJLDBCqZT7cx8hBxDOVXirivyp1jRs6H2ZFXBVKJg/uXHd7Y5htiLrowGBNSA+JbzbCTC
45qWWJACetyw3HzFmorZhsUPiWk71xih3dWLZ0wb5JJ9dBtDFvbNZ9tNvAPRV/sQCO9LZbHf25yC
3WsDJNRP3oXy+hC+gDGBM4nsBwMUHkrPdFONv8wy4FrspVSstqJeocZL34oLgELjzBhm19amCNXM
iPpS956hZOY/a9aTEz95U8nFPaH9d3RH07V+Yy9zuZxIAsADYgffOfFKd9kV3IKCfcpyvGRiva+h
J+x9BQK5iqbQ3rooz3Ji67bVEZnvdZiGzUDfmxStwyUALbGoSTUoYv3DTv+Afzo372OtpYM1IWXA
xtLbK+LmGXBQOqx8rs+NhFNdEQs7SDb3V2QsMd7j3k7o8/uvwZE/mT0ZKGHLZi66f5OGfm21zoDA
lxfN3dG1/PA6vyTEoCLD4a4h8cYLqq4ovvifTWVNg2TjDoFwDIGe9y4JMdp9MqbF9n4R+1c0mPqp
YIqAuYkXmpigwPar75gtermw0Cgt3hgk4oURF4rOhIHk/TYZ6pc25sANY8RzhjA+VZqbMBlHL2C6
at7oEoWulOy05vICFtWvyZqthYO9SPG+78ig6FNKFetId89LbaTZeXKbrOFqHe9/QqjVGFF6+8sW
aQg0RUCvHCLml9yaYTI27GiSmQ+J55P5rdiIrJRYQ6PvRJS8BNxbPZURi7yxzS/IVXotaqWVLgs2
0kMmlUA47rEBlStlhLpPGw4EFNJ2SxOvtw1z3oFCt3VNZbjDD6ikPuUvjtBFk6rliW4fcz+ogr0j
Db4Nus5/OsL/Lp/aYLwoUpJHcWPazAes9sxGpe03n20uRxgR9lQyi50m5XwiBC70k//x1Ztmc1GS
resrJvZPqwJMAUWD1QQGZgGH+g//ESRUYvBfBgfF8f55XZ1xZuH/c2QqDgQWW2geFVBupoM4Tady
QLUATGHJ0kulkEaobND8Xo/9zN+Z+DMNDTqwvkcmHuwTvc+WRBHn3Yr+1f4EIgVya1mzpUOk7L7r
dL9VorkQz7K2pr5TAsgWrVR1y4qeh1MOanAIa5i5qbz2N8VbKEAJCt2QxG60ogRwA7Oio+lo9koT
cPBkj8gGetcI84cx72g7jyBIOAoVQnXCNrH2i73eVuHv0YUBr6aHMTYd5GpjgdQtIMK9MmkClC6J
CTmv4KL3KDt4b+lZxJKioNkwHgFqvw4OYxmzFMO8U9ONMyuwrcXfKukHZnPa/d3eQm6jUG954Poe
THdxjaNiMzGrmvgy8TyuYfV7bozcg+TtqAZigBIOQlnHqIzzKPU2PvKbiqh2lCEnuZ81RLEZOPR2
hNqgNiYuxxRUVAK7aSsq/3bprzHAc53Zk2M+B4RTxgNVvhGH4ceP5dV7i1YmR3IZxTtMxKR3jpkW
DGYkGF37nAj87+AzJfMMiIysiNa45+3Q48cn0ildDux1gk4GgKhgXOzh55xMK3OLiiDKHtF9+0Lu
QvERAnm6f+hxKF88LOGsvwyA4ME80q30jNKPawutO8qa2F7jhAX3wHsmz0F4J+kPAafvqZoAu6dI
KcBMnt5oyBM9Fqa0x5joaxpqq+f9wcaHNjRnqJWijGipgMuJRHuH1GwBqKi2o82zczQh4cujGBhz
U6vH2n8RfU7lC2L0KeJTLlqmDmWczwLBBfwbcR/uTUSTdhs6A008P6MtjcH9F86tqu6spcGQjQHj
5pffhPcDz3urT2PCfKinug+RSwaIXEG2udQkuwvu22eryxeCKTflezMchSA4u0ZQdoZeYWOsABcD
Ef0pTU+aa5kTfJZWN7H/hrcPuU2Sh4aasNobtox31ZTw0MnsQ6wAuPpUlUKlQffM1J35hKn+xuGg
YyRn+DQhNOAywZsEZabOsG2J5h+OcqA9f78P+P7aVtrcb3DQW0e9IFwS2jy98RG4ONPkhG3TVLAu
FpqBYuB6u/M+lKACm3pCz5d2EV1maDFjF5fbnNUB5u3i2B+2KRbk9AIvrPVdR5k/DbzdBFWAZ3AA
7Eo6WEMOIIBkSOvMQ9i13Pm7CDaaF1eS/4AQFeuLqQPN13fl0RE1T+v8OJUz6z7kRFBd2atf/Q9n
cHpOb6MddV0TVcQlnjh3qUGAx/Fuedc9p+tfv5M3TtO+kzz3XlWIPTRJa/+fRVLYGbFHPPHhQiJ4
P3U0Yt9QUzthxSWOM1HRmK2hevppbqFssOzVcfKchTUlM1dAuN9mGFx/40GifjwJpaTNSy3+GakF
BUFpdd9NeTGAdgdbWRhErxD81aghwTHwldch7sMps4mXmwzF7O7FQcOpP3Jdk/y16AoL2XPkD0dr
CTRBXUV8ilV3u/MPjeVhtY3/Ztb3Dd4NihRRFFOIqTLAfDyeMqKBdsWRVo7vR5LcYOJM6gmyMi19
sXv7Sl8bU8hsmCDXAtTdFt23d2mQzszbvUGzjGrqkWuV+UNhR9pjt0Bdr4nrJBAT8dnNKbJM3Br8
4aa2aDVLCnNYJ3Le0jnfy5vel/LvpEgLbc/u0kA8+cHwKTvPOqF9vJPzPSKM06QTz801QSDANZDu
l49ggxRNBwC7txkw87XckGZ9fn+fu20gZOhV0tYwKToD11RAlUP1utkwFSt6X9miAl8kzm8v6zuS
tEkGh6+DAYuw/HiaH7g8INQjqWisQytqQJEQIZ134Oo+42WeN4YXoB6KwPUsc12PJi6P/QgmoAHw
h4+zvl+aikrrrmnfhG6kyEfn4Yhx2Eiwm7rzMFfpuF4e5kYnSEVpAf4euY8ClWqxolzcIX5tN/6L
Fx6vt7VQczvFgmxwr7wTlOHA9nK5dQyqlLy0exuaC5CimT19dVg63gBU3B/xLAXN7nwEUl9F+Zpx
Nuo13KfeTm35EGToSTb3wDwGCSwYiPlvhKUXMrIel7c+WQALfG13DiVzoMhv+NlMfLzTgE99KILZ
AIAOk+2+dsaL2pwOB/3FyPN2BVfvBbL1Sw4bfqnWaczs2QKJs8tMT18N2BPHS5JZZw3rueVQ4jPW
c2Lrlus7nmjnhPt3STEqsThiWF5yZc9232zSJ+YAA0gSHEh7YyetBv8RIHLYSDLgZIbFits7q5HK
sLYxM5G2NFcNpjKhg54o8lk91BLzKK6gL+I8Q6X4/gd3ajwpxGIBALc9v5bHKuLd1vQU6SIX/gb7
QQxChHZwXo8WzmDjVEKq3FGsVXgfrowYyaADEhcuowAS29rwpTipjpNo1httWDQQDpySZ0ZTljZc
9MOCYhnJAhhT57aIUYVw0Hrm6uhQNnh0dzTyDFgBz7xE9rujlzSyvmDo3J40GBRhgqsxNtQOfrFl
LeCX1jsiMGfDx2I5RhRhftHMzDGdoylnPBHbVB4uZAlAuj6F3Fh9d8tGa870yNgfmGHSLmht+cos
WpxVUqXwN/Cg8q+rYvbpoRU0fU8NDwXOyaX0tjOtpxHmz9OsCYibGqKZjBRB2WfXOMUjvBM3fChV
ejDVBenpAwGJRiWdPyo2Y2RIM++Jqk2iCO06mLrJ5b2r0amHS0b6jbtuhavwH7s5dqPpvifU/XGP
KAibA+4bsgC2UtQIbb4LGgYtD8ruPb0RaBlCcYkRzb6ydUU+aqxgdjAvcbCi4r1RoF3TG0awVlBs
myGzR7on8o5MBKDlBxHchmGyPUkK0HxUI62VDd4LGkx7wYP9lcm0BXvBefTpzniHhm13JTuvObg0
GPkW4mGNktFJpPmNSmagl/RLRYgJWSsApubbBByuUAFaGxCw22IwQNdwT599ENG50KBMWBZ8vBdH
4ZkM5CwkUvXcNMqzzrvNEPEuMsArCMlPXsmVO2wEDfi4/G0zTQYefGL8EhXpLGuVLa9zf7aYN2l3
U7q414Qr7y63XmckP38TE1GS31R7o7D+a1ZcLLkxUDC4Ul6yTlvyjLOdUvQuto8x0dinsVJiq26i
8v4yp8/0bSadNBcI8JMz+NgCEH/J+QTRyoLVEIOy7zXiYR0IL36gXpvy7c+1NzLCookP8lAd1+Pr
cnafNRP1jp5BwbYz0Npj3tsIGbCwGO2dirGTWz5RPLn/VqE/veL3iBpuPfwTeqekoF+ArmlNzdMM
7Z2uxJp7vGwMfieGnGacP8XOPUzdmxpBKBL55NXOqklU+SPj+2aZ4MYZxU1SUxISp+dlQQkEWZoU
mvNxWT7pffMQ6zQoHSniceJWXGL70Kjt4WQeQ04dS+VXw80XxiGBfxt2j8HXOTXUo+TkUt1OsdqD
h/K25Au5Ux2f2OqV23is/3/1mQRgAuqMzWE7xHsJuHS/HKS14spbfwAVamQKYOWZ29tbZhYy6CM6
yhc1sD+iYgQycpS/QNMYsU/uqJDU+sH1EZD5doUqXAK+yIiZF9isHuC8GQSbqq10p/Xur7UtzPN6
d71zbODeUMOd99lWCWJ7SJoDMacfWCwPfuz0QjaTuHx072rYbjyEzobDZ+9HUpoJN7/PvR8SQAeT
PoJ2bVD01rsX2F1ry0WoFtjQnl+WSGHP5KjnpI4T4pq40uADJnMtBztUims8xQG4KmBEJmjq4q8s
TEMg1EkOEHC38EtszQy/9GEM5geGj4imznjgvHcYuXLrheIcq14S4iYjNl5kyjU1kN5XXEaAUpyC
7KB9+dIlASWU/J6oN0u+qayhqSEb7Db8nCTSwz8hv2rzGis/q9WSdAK+BSsVgBSMojGFbpe4Cx07
ZcV0q3OBSSu3DlK+LTQrsOj/Qohhj5D1zUhCnxDfO+dlejJGAFSAwHXGYfJUzSNQPF0BGMoAUqT/
j75VRk2FFldoGD2rMRCO/l3HyCo7kyncSP9mcXzeOxc5xgpADqFsYGWQDDppi47VTt7XdLcdjd0g
2kebGpcJLfzjcNFPoL1/e9D86Cb3l3nI98ehm/cYqIokEcNu97uaPDggQDcDgaYoueEsLUWbNE14
QLDTW4ZxYkmKBqICm7w8VcHBzehFYYYArkj0Q9cIKKvlp71VMQ7XbmsKi8H+1E3tIL9iT5LnvbFb
n1aIc/X/4cctSFD1/sohO6MXpkP10KWXCiPNLX51j3CFcgkm4eSz8CgOsu+3BQGZdSuMxoXDukHj
8yndm3XbrY9HqXOY2gDBCq1E/VUT2AH2pMZIJrIScsR5ipTD5Gq1DLs69vM5dX/jMuG/v9Vz4JuO
CI1XGcpz+CDkPvvxHs6Hrn4qBB0BRdrSBfLnZ1rUS3vs1iKaJTeXn2U2SGvhadczhz2yO2TWRDkx
HLNOA7pJz3s4MoZPoRKuNpxnNIUI1pkjHcRFQvdEWZrlkq99qep3c4JW6F98mZtX3ZXqpu6yldWe
/vF4vHcCwqFjHcSY6slKfTs2j5FsKU76/F1SUH5QZ1nsyJ4VsYms9NNUAxRvhFVynOo5lFxHp4mz
8RcqlE7EDGuGKoxG404tdOGEclY/IQgxOJem8EAb/RITpEG/MzyQiFkcdb3+FWFeEkRoatJTcKIM
aYB8yACDTND8EpImBbx4DZ2KE7w5yKI5+HFk/vMIir+N4FEPs+MlJRnM8XL0t9YcCdQlKxlrKYuF
lgiZ476fY39t2piPec2n63/emb718dZ+0NvOXpT23IlTPcllW5yHcRhO4AKiijI3JY0BKFG/VGMV
V9A8xs1r0ssN/euGjYW+SFCPLMtOQYP4YhyZcDGL2P1BvQz4oAKgNsUglVBjRVR+gH+f276LWgsW
4uiN/001gnxHdE1FS55cxXg5jCwPviRKYSZ71WL1v6l4gy3+WZ+X7LFSfiNqci2D71pcPjG41aVB
l8RknhEfYjWSfLSprDpj6UD7osCHBGWHVEEDOcQ3Ek+RSFDosOtkVycTdDtyhhSYe1JrK/TaCSf/
qu0dnI4bVd5HLEImzL5WMu9qkhmVu3UAPmVTuW3VtLW1ydut9ItPXFf6DUFme3f9QgC/Gz/aY3PC
O3AI8g008G7B+s1Wx8plDnIyY8ZOXEntqI0VwYWcIsFM90G5XC2MwodFhEHA0hky8QvEVjv9PXpZ
i2qr6B2IsiMNUB3oSdFWi0t3HVq2hcJgdTvIa8CTyb75fokVicZ6bOVMAePWEICDFDIl2VEoadMi
/zA7q3SW1xQVTwU98tBeAqbytJIwCv8tL+yKLXGHWTutHl+sxXwbRqP02QW3CyiCW2fsnGVybg9w
S2WQ/6eFGkBFu415ZUUipappq29Np5J2ytywHNpcCoee1hqHiovZo/CiBIRFvn4wUmEWRKcZQkZs
XOpH1SiA5nlBtbr2rR22T7MVpceInKrsMRHk2Rrq54O21c7bz+GN8WyKbjfpCt1gE/zitsOUHL7K
TikqTeALpnXVy+xp1H9raJeStR9kH01WGWIBC0iZaFm8p7o47rD+xOZGkKt6gp27fuAQr6/L7EEo
/uB2hlYuMn7ynUeKoytJwfBe+WiBYmDtjVi1LTTcDEpXghe5V70Cxr2EOuWO4vQAwBzVB656zAIC
RgxwsSlUbNgC17LuEKz+5ldtybKO4GGC7OPDjyHTyB8PgjbidLQkmvipkp0Fh/SkhlUTNzvSf8mO
o+CJmiJpsTreH9MTd7vKxaKYWeK2SOqUilu7eiFwg35fW99jfG7QIZ2M+o4OEq3Vc49CEWEb+CeT
DTYKHEfpgIe5Dx6D43J/Qltrz4uQtaoPuKtn076jnonxvMjtUxiWNFpuQeV2AuNyKUpfDWZ/kHbk
fLe13PI9POBvg4oLJ/D1nqG3bLSp7a1OA60qB3z49UBouaF5785L/mCohOeaG7t0BHm9aoi2AchZ
NvHZPOZ6dxXU5eibE0Xff2JPF3F/wRCX/oaasZ63QevGIuSx/S6lTlnyLCZ+81qdVeUguJr/bRcc
qoHD2x/luyiVxZRKa803PTr93A9KYgLUy7wn/1q6XZd9PwnlghErr32QgpNadJPv/quRKKw3rLp8
21+hu08nTqYuHItDsqpa2vwFxnvtIgshJUSNpmMPWf3H3EoagQ/WTbbMpkCf5be4GU1hlnMR2i9a
jDInS9evUcji6EEWoP2eNrCFyZWWH1IvwHFZPEqKJp85DEs0Mk9lDsvj3BkdbGZYfcDn1QIqqhxX
8PbmLmb2t2SNW0J7JiJy7Q/pswWFZk6x4NnMKiJwhSJZIo2BVx5GGQiMHYLxi3MIMu0LecGA5ckQ
6xqKma1frQHr354LcEk8aOTvOAKTK3CZbJ1nnYiPbAGjUFyrSVGGLKABa34sgDfrC6wb4Xk1/0U9
pMFsVKuSM80Uh+CQt7uLvMwfBISNNfCQ+3mkqiVEF/+QO8pA73blv/6rrxN+14gzq8iL+X93AFJN
Zutrq7vLqEi2OpauBB4QiyziqSjFgi2LFn7bLFMbaW9eqGNYX+GcxiW3dZSyw99Fl6UzKIvx/lOl
7N+my5WgJnEjA0s3vasg8iY72JOTdiQoWMDIA0N5OXBNCBSuQx+C1ZWAx/HcRDC/aBTK1RIhA6Ol
1aj8fChNSnvdpmSem09B7h5L0cS1LuehyBE1Y/lF/fb57mL0KRfWnvwoRlL9wpAmuDXpzyCudiKH
7rRfn9C1YQHX+9P4dVk9ttYCNklHlb+9Lb951uCcBnY0BAQT4plTfdyBr98RZOVof5/Tr8j+ko79
noTaP/BycgzI1dUc0cam6dZhI8jbAZ1yWBitXAyUabX+uqmw4otHfVjJFmbNQHXT1IN5vsfP8BXP
LxRDlbFuZH1uGfsHZurSYP7qyvnmvs9oUM9fd6SBVuu/51ArlxiMduOGT9chezYXCmX70MzhXvlU
RYk7ECDF6Hzeak8uV4/uYuAYslhZ9vdyu0yp1p9wp1VQeEYmE5b9rg1HTxv0YTlVmL9EQfuipKxc
KzbJRcWM1u+FOIC2l5LFmQs60Cp8ctWvewmaQj8D5bL7OR+JjffGFYuER2DvNN0XLsQDABiuagdy
lyk5UozSP4wCcimvYP0tl17YrXD45CTWDQkq5yRFtFV3Gw9sO5FbU9l8ZXskd4UlQJui+YjY8BkO
kpKR9hqf5ZnHPq/weNFIJAlttvJOvGyJOJ3f/HcFAcpo9rB7z4ExWkohc7YrT+qeFtmPON95zCkG
efuiU0dXoVSbHP+GQtkI8YwUurZLiNblW12VPkKSM0y48Gf82eu+VxVwXwETNaOMMdOKswo68QhN
uMtQmh+8ToEkWRLzKGwyaPbLiRjpBkdS4P5lJOXIX2CAl4nA2pTTkOY/OBr0qa4YqjQvkknoDA+O
GMkaktXG8uzEWvI6Vo9ivvJZyUMxZu2ZLh/E0yw2OzQLrrFcxiPVgJK2OLqzr/qj/3H/A60qVQt9
iLyEvRrMW0PFKqst+vIEXlD+FUeG3B/tPcv0TnEWYF8i7y0AXZ1gwFnmDyA5yh5qMMLQXFt1xClB
4/9vsDsq/wnS7y5oMtfhn6c92oGXvuJ9vtqOKA9ucguqhdGzHPTs8ktAgDSrN0HCJvVMJ4ffdqtR
3TEmuzUz8d7SJ0+2i4B08nIw2b8hXxjpo1MM85371YG+YR75XMxOttXSmJpfhBt3XlIwPhjYsub9
wuqd9tJgBdfhPUPHrtIF4i0Yp9aHkdRRc/agoIOhpM4e/9TRmnCuUhektytSh0A7GPLwlUy0USXv
b64oRzvZwnCOufBYuNWWqgMDowrj4RAlpqTaWkTOj051q9B+8iszhzBjs0iJJZlA2U638eiuZLwT
JiHfohXwRDSX8pqYr4jPeZqlYolJUPsarc9OkIXGMCha78D24SMVIFkIVgZsRJ5KP8HBqfPe4/yW
SYvzPhubSaMHscXLYksflKgtX8mn/uON/S8EssPxN5Z/36z9HN86ALkuvA0HKbomtKlArk8FEBjt
mvnUYH3zNJKxLcn4NOrmaLtSz9CgJxcYPrquo6biVacyseyrprWBPpmgiTpvEzSYFPQytdBl/icf
qGtZDGhREylO2KdLDDUwqlhOv5RjPMq7xzg+PS6S2+iIpnOPfvMSRV/u5WVPzRMJnQjkMvbhGPJi
UNRWXuEjVtp5BoMhTplzaaPitO2HFtKXp/B0DWh6VdBk5KHxx/PgmI5ewAUzYoPTgGGMIcWq0KM/
8t8O6OvNzfir+iw0Hi+oSSEYRVWQfef3NCLDbCatCGPEPUzXVgiF2PVdA1NNNK1ZEiODupWaVE9a
DkSikzl7fNojLE++VAg+a5UBLu6nbWtloLOtRnqzxgRQDEk9i+FIfWXPCwMxIk6J36tONApr6QRX
fkukixGVTKL3ciajRz7YiDE/4vTFZxoZxPKZl/1AyBZaFRY2orEKVZlafzApm8vEWkXCMe3zta/e
fXnRIM9Z6kTtb//Z1EA/PGnMyQrHs/tEuq8jH3OHbh1TvSAiANkD7BerbL/Vnke8VmZrWYn/9jI9
RjtPtkSTUahU7sjtvIOaEVx6bGfeRUIN4486p/fKOSM3EHmPicE0A6urk4yYMnOBcL7QIWBe0Ufr
vdI1PXn6L4LFzaQIufYQ3n4Q3/QynrzpTrAlxHEp03czCJh1K9ZL4dpskT1YkJKcarTjkaHlUfHp
rguLi7ZYeCXPP9sf9w0Kmhf9rlVztoHAE9E+rqy+xwj7bBnPdWFOJxYIKEduzpz8+AKkEYSP0amd
tzypmP38YriMoEcKK7EG9jq0Hu/BppCI/jew2/Rl5F1ft/H8UNP3wFXF4p1MRD7kjo5oM2eqgXpd
uYskwqi6sAifBOoiGKNjGhNmN1e5srsEObabc8/vN3SGsJxnVi9jbnsSUq/BSE2kdxiQuHBSe0Vz
NsEpFLVG/oO1/eSyFQDLuUeR9SK57qXXXTTOB0I372/Sf+VEkgAoWL+MGi4Ah7sKypALnOAzZ5jF
m0UluJTrMX7VORw7BU126pnguePpzTFEtN+SFERy7MtHhM2FzjQBxvok2SEbf/7hzI+v86mzLrBp
nwZD4hrC7d/z2QtxB5Uw15SwDr8nWs8+HnDnE3ljKkNsO4I8Gaj1zbpPDjbLCGyNmILKdmTb5LAm
e3ziDz+R0WMn9n2aQWcWaFBv6sd1qhYEmbirQaBPkHbp9KOIJt+fCtt2bNvhYOs7YReNLEVb6+of
ersBTF+NrPV60gJGviRmUxzjFP5eZ6cu1RBdWuUhD/2NvUUmV94xcVtqPb81dHfOqPS51Do8O/ti
o47Qu1+wLszRdukYLixPOk1bisCwCooT0jypfQJNjU5u4bx00ORYHbB51pGAMtjaV0B9NYPPPkA3
5+F1TstVoAH/ZCpP1r5ZJzV7g6C1eTqUousdMf62wgqYJbvgaQl+GG6ikItjs0zhYTRrc//3oiu4
JHnINOysdHjuX5GoPGHltBBDhF4xzhSFYJsvSfTIDrNhVyDgXyt1O6VQ3KB0P7DB7UQqwjM2UE6U
8R0LXetBaULuHCQN/4AWaMkhOEntFGDUxF0k1eUXaj5h8hdwJzQmYlwlA/Ob86XdJ8JZooPXq3jV
6a4Z3FjurJVwH9EeepqYIZo/lMWtLMax7GsKe+ZdAPED2hiCyv7ZjCskQAlfjB2wOMHE+C5B9rA8
EQWVaUdT4xxUhDbtK8M1oAb+WLx3l2gZ0c91SK9nT1sXF96ClICO/DzWsDtR8a/syEUQQ60jfBTw
ysoFvqtJBb6+pk0bAO+iOeegpYGUI9GPx4xUN9ALgQUr9K9LtB5MexJHYevZJpA12t8er2sD4EKp
vHKUtRJoO4lhzeMuLzdEe0l1Zgx9lrue1LEoOxIQ/gjqQCQQtvJTmFhJ3X12AXqP5NEN+PJFXmJJ
m1iA2//poFn47GkPS2SLlKZnqJqI1GydtiNxtaSkKsnK2ocQknuuQq7H8NpXNJOs7lUx/LJe2572
OdZNZh3u4pa9NJu8u/dNfMeoB6z2bXM3v8jskHf7YRLTxqAImQH4mrjwR31tJQFCHl0j3ZmOPOKh
m4Ox3jctH/S/XWUp6X3Dz+XLmyMfx0Q6xLcOIQXmsS9DNDqc9FItS1DrQGF8BEVE8J9rGAIultFG
LuXEwACVfEVHa++1Ib0qDzsMBGVXQK6czmTpFlasxDa+yLyHcjfD3DbLa59isrfDuOu3kxByrAFY
ud6+YjT73qWELvkitwEfNIaaaPj42c69fu2bs2G/5FqVR2zzQWLCQXLesVJCvo3TfsHEZ0RjwUme
Ubaxr/GOwQPrAVt+fNQlA+Q7TXAL3DqKhaWtJ2nWJXzWozKJt8gtI36O0SXx3q8FL+GHG3VSr8ts
DRAKypUzvuhjNGOUqddypX/7GmmFy1KqRNBHF7AEGX5HGB1l+w3whOJAnBXBhewfKjlKENSBVmif
5bBB9TA5sh7ViP4CEMz6OrTWjY5jIElRdvw7X6EEyQMJ6orfoqZW2dACib3643dMTr0J6XlmlBXI
DRv66rd5FXB+UBa+81wAp8TsndkueNqXheAw4ciMkZala6RG7q0+GPN1alVogQoC7gELtKHs5WhV
cI7uD3aFSsxSDArSFGgpu/WpUJwY2XsYcEXFu1Y+kOOWRtsURWNJgDfrXjtlJxLbBWPpPvDDcARu
m8b5XAy3HneXJtIi4zHUQr87yO3lw35dUc4HCVsbb4XGt5Yqeb4EpWfpP/4Zcpa2v7pV7pPF25IJ
YwsEwpAwTpV7imqQZxZz46s5A5+MbtvBUZu5j7biUxJkVu/YPU8bpzRfPLCX+ryOAb0GasH7wc2F
8S+yu1umcbpQY/DLWeIBsXyJJ4LZWSF3z4arfago1kEfCAupXZF/XFfPNeRM5AEUpKqtKBHfZoFG
hTuMfpGtRG0BnUbBz6xbTbd9lSHPF5KeM66Q+psVQjhcSjcofgwsfnc7kI8M+tHa+c11/RBQmTyr
Zm0TtGBJ1xPCPAq4IZ/Ox851qi6yFohi0NBhAyRhsZSj4yu/PKARzI/S9odw4iMTkLPHcf+hPr81
SNjfXzao0Ez7DiZcthm58uThuEaW+AGiVMWV5TGVBJJOG9z7p8faPtkKtsAPMeovvEv9Tg7EZ+bb
wD5dt9ZlnHwRkg0MxhjT8ZFW3gBfPgwxq6PFDP4tzMQtaDbb1IBOl9GLaNOuhTdVp8jVzTa6u+jc
l6Q4rEgvuuET0V4wZzrszz+H2icB47LteSPMRTIvdLNE1Rtiu1PY+OgTgyYH70VTQ1dkJZt8Jvyg
wgnz6QaGqyzihqUFlco74i3axWFQM8uh7MWly5ewogawz5CCG7cfvMLDlx9PsQsdRNK/MiJrQWQN
/f82vJ/zjPCUZwdhAX1Yto014lxam1C+5/tNSGjtCWFn756nnmdVblYUH8JQ2XUCgSuQ3U3PZpgL
LmKxflhv8pBQDL6CEgn72IXioOfOgE944qdMHrxV1GSD13RET6bO0OdhGrqD6j+gCmpu7oqGSeAI
6XcfvTuJY0XPKkvttRkiowK0ddTrv8Staz1kLs/UHBH/4KIw5iFk/Jj+5aTUlu3NYUFsGC60C+zo
/JYLZGemTjzABc811NCUtQjYUJnahkdRj17CxJ/u8TrfwgYdT1+HiHak8mUDjENxyrRAvLGlKmzw
oEWQXGCim2hrqhwAYQt5B4j0T/YgyUvSjpt0i3jCNZoaXtMEmqXYSQbw3IXkowuEFTYVa4/PmDRo
7gB9ksdsBnaXpUoa3nEjBYKiX7WOswa8DkshBwkjc4b+6KzIAprNFoyBJaQjqV5yzz3GP7/kiBoR
XEdIteCQu5abDmW9IgV6rQ2LxfdF7V/OGZNIpalX7fzuTLyHqyRg1gfxSpxaZ92/YFhiplsTnMWY
qnUyS1UDtX63Ty9dqYeTHGUHCEeJE+LnTu2Y2VYWJOsqRJUDWqJiRjAGZUtsurovc+8vA0eDwi0N
lBSgtQLbLQ8hTt8EX68P52zJEqoBWVxrtJfr6KryDKA5f+zu1+WCeZuu1f2DfzC54km+XN1PZ6g6
6F/AEeeEM1rt/aDJBeOVgh+zBJKbNMh35uffVokjkRYIocaXvhi7Ufa8S9Gdtm5kIpGTsFShtCnO
VTzPFVb+FldZq+rateKFKJA/4Q7AvFgS/ZCw13d5VTuLnQ7RsWd39gwn0IFOz340h9vk0C9yRc5C
7McKHkf2wsEtGyRz373VsmPv44xGWEC53wYztNpFBumELUWaaweOQa8SYjgspxWngDz0YMwkmZ12
hBctLW1lLj5R3pWyocLUDw3ViqL424E6wvlSbttP5psXWlS9N9uvBom+1yXiknKQxIwOTnNZ9xKe
Boqdt6h40QcQbn08TJGZfeSweANWnSODV7KuO8ZWcbsoyPPwId2D6m6KZNagDhqI/7ipG01hRlPp
UdeP4llYqSZTiahxxwk6SXNn+M08TUTwWtm1l3F+RA9rT0fIZSdedZB9ljO/e893wUWBlytGy9wG
veyXQIF/SSxUmN09lb20EIVskqINAmvjWvzLVYpPv3MZIShuDTYN19MSwGVZ0dDtTzA13urbK7l+
GNAxvHDz0wAA0+8gUEAEft1RsIWK1YnCFQm7qAic5TomggaVIokI2x0bkC6G8vlDgpgmFskHKWkO
iEX0DqE6m/wWp3IKpfrJrpZxyrll3WRVPNWRoBoCqKIiA7IUUy4o196xkDuhnIDoHe465t/mP0+F
rpdrbclpHaUKGt7pz25Tv4yBue9sakkUqAkmpxonBDU8WqoRVE3z6EUFr5oC9djBwEOEmf+tmgEn
Ri8ajSBkmT6OiQ95jeI+IPqF84LaPnbYa1cZ5b8k44wLuISy6zhg0USxFC97BKPJaAP65N3FeXVr
4dyT8t1QjrOvD/em1b7f0pf9Ulh7x8NnX2uqDHCPrLLJdJkXt22xs8VO7gF8z3KX6d66GuouRhk9
rGOsUv/RTVyd1GQ4HdVIwUpct9Gj87D1y3FRKNAn4LYdM43Ko/nUtlEvL2E5Mv/q92KfrVKG1Tac
ojqX4nuUk06JLwostgVelPqjWRqpLL1E/Uynda7znKLEs5dGMRDRJapYnaFM+RajxyuPfunfVQ4w
CxYpqRH9TGR6ZcDI+e5Pfr83x2s5bkGdU4DHPk1S6bquTAT41AsrWIDc6pH9DMNMB0Km9C3u51Oa
KhMvFIDgszA1jDScsE6NwzPu2E1FF/r0ysTEAuF4ByJLKYE1vXN8pCg9Z0LKYSdcC4su/2/1WRGq
Ie4quXb8tcQlf8vNfYjFDH5Qvt5QtEZZp7zgchfArYBKSNR2cEBqzwew3Qmzl55w7zdBuAfIUMnE
vnl+hsgoBAmqQjBuP/48m0MTBxDrbDcmQtHWirN5VdcfDl8dqAlK3D9hoj64VzbzhLwwfYG96GS8
kOFHhnXNC+9GIto3s4ZbTab9jgk8Tz83FkffzqLq782gI65ZQcaOgcH9Bonw9zpKyEHgVbecP50v
iBbpUfE45YsM6p7EWQu1eV/FrCQlw0Q/r4rlIiQPfWMSC7YZT5BbG8rmaeSqWbnRf+YRy0HT/KH/
B0s33EE4Tp29LkCTR6XJcBfCydE8LMkGy600I4n4M5lfY9as6pazlkYyDbXmJjpugpE60KMrM2Je
5bZWTnAqPM+dd0+VxyVbsHLrVwv5dAkMG+KQZRqi6lCE7KkgUR+Mu8Vv4yH+KhgYAYta3Q10cK9M
HVceZKQ/nuOD7ZZ+QIbpbh8Uxi0+mqmi8VQdEmDYkOkoUex79fk7GC/i77ZZBNmz7dSExJGFIkzz
UHdGX5i9VYrCX7L0D8T1NVKsfds/P0XAfM0GwZfRFvlz0J/8jrg304OS0rU889OZA79xmFBBxhZ9
AE37wCco91RU1XazAme5TIy4X/M+NWDYDcgjiiWDIG/AtrIvF0Xl7eU2ziFumf90iix24qI7awZm
EDoDxFrY6/2er8X92fBmUI/SUhNSHQNJXqD/xNLcElXTPlEsrbBTR+hDAWAlxITtNVZbY9EAPy5p
E+Y0PTnmNyeeWbzDAbZQg9mEbi9B1tW/U2XCDfzZKYmublipZJ2p2mjdV0T9/kAedXixnVBqCgIT
peSvhIuq6XZBHD3BxHu/A6afAExMK1ISPP9Ig8pqo4zsKsWsANvXuJl/cUc+eWPBizyw38SAe2GP
clRuKS9b3FzhkatLBpGDsiyuQwHnP0NriBthVC24geL9r/n3ek1yso9B/iddjo6YE4CWgiIa2emQ
DC+pfXnbaeCw2gmBw/8bGIkcc4ItQ+KaUwE+JvBHIUOAZSVTuzTAzQ/yUIV1TEQUIW0+F/YCE9LF
VBv7Be4FC8/XC7jvVc0LNzOBxCbObPqYCSbgNauRiN+iKQSFRuc1MYdzF2ZtHlSWIM3ePd+CNMZ+
NsUQm41LIqKCA6v69QylSNvxMadrdjSR+QSflNOc4HbuQe5weVhfoUu6/kuDDN75BfCOqjSgyvaY
N5tPVJk/mE7i6HDGRrTKFd9YFJKFUeaQxL4tCV3gFPE7EjQc/uaTNDMyU7o8BLopjhsEIwxdj39P
noMXe8TFxGu68hnEvO/ZKjWsQVLSB5TLE/QIW+3CDhejgdWGa+hO2aHX2zx7ufjzzIaLfZmtC4eo
FX879DkKPZoZillK9B2X36epuGTn+vxgwSAWQIIwayOk43ALhe4zBs6eJ8difpbi4RB4rXtT/8bJ
zYS+RtHIx5RgbhvOjrdmoAyS928bgrTP1VzmmgzzKfQZQx2jn7EcE44zogTVRm6fJH1L5WfX7UAQ
MGqlS8Wcrds9vbEvgoOd9aG9KaNF2XNq4Rvp3vGXCyxaxncAvgkKLARueWXmzbgh9FpZ8VU1Ul7B
im70/VD4bUox1VyIQXtb+DxKK7VqHI227Ni9piS3jMpZBbj55ciki0mahrUTEZ9QVWD0EQIs6kvh
0RGWgixHn+JIMJyVWHl4GeKPjT5zgNSKCYg6kckZymcQmRxuGUFe63NmiNVjYyTl8opUOnkKddgt
ouR4L8h/pMvqOl3jIxJod2pBoZxx1eVuco9ugYMzEUuL3gnexajpbbAPCTIuA1CDLtpHtdv03iSA
Xt/VnioSO90EfHxm0HNU0fnAs8GWRkW3pQCurOiMchrhsPjgk+Xi0dUwGf2UFUfLIDw19d+veW6R
w0eD9kgi+4IybX/xMCuhLBxkMHyqT442hZUg+K+ud04rmWBaWMqlEpy9xUNbZs0BuMLTRv4Ua/Tl
4Bpkk4Di1ZI2Wkwvz7HjzgH9dcal4UgFZIhkKVwsQbtsBemCUzfosxEKcBo42pBY3KNrJjuBQbPM
ROrOc9jhuCUk03RSxmZ9Qe1jhicCDQSzEZtZXyLDAiycZNe7udVrrc3qMcDTMTykitFaxwBz60Wv
KlpnJCuxYp6TXnUT8UUtYLLxNmlVR9Rrqgqr5ZUAiwvENZCGjW35p74sz7vBNNkU9XpO4zvMWHyn
v5L+Z6mLfws7cEcVTV/ktxPMYdfY8d6b6Ciunjv40K991HX8d9/LzXiLJF+IRzmkTFHUNRnlAT7r
OlkHWzTRYlWaIgUIHAggt58v0tsUWL7kgEtxo1vrrojciA1+R1Sc/b6ikXoPnJY3Qn4iL9KNK+CN
uDjDcKaxxk6UQNbX7UCNRLKP25uXJeM8Eh4n4jXrfI1u5gPYrvRM3g7zE7zQHp76PrtypwrpUQ2e
KKh8efpVv12rhOl3FlwdooqfgLubQxTOOoyCG1UIKooE1g7FQIBBa4PtRuFcuVOIFMRnZFTPBXHr
n5/btU8cJ3Z1dSqWJMB38Qu1a2eOMolVlTLodjAhLo4IHllMlstU04UELUzB5fexVisH8/f6hk5N
Fv0k62VC8T0wL8zuQvPIt0NXMSaDb4XmRMATtfQ8Bf4BCLnLb1W2/sc7ZvAF1pFFJta52xN7EsaD
APzLKBblWrRqcO8P4GMs/umZK9OiPLaahScqiSCjQZ3e/b47plnPinla2XeiolX+isiJLxmAadFv
ry2V77Za2BBqRzsqi6GsEPkcj54mmXjH1fG7uexMuOzueoUN6J2tzKpV4gdnsJrX6sZlPPLCRvPD
LQWncAVQxpFU7jOAUwxxhXYGr4WkJ0VzoTZUvIcESLCgxSwbSk5kCqT6lE4krQDWxC3tiTWDI+oM
RdWqy++ZgU7s2fMMML3sq895YiPvAszcYVkAWyjQkPirO2bqJvRLSZ1kSR9iRcFQEW1JGt/L0z4x
IEHNoZbcaeY/cQrOnyG9i0bHCySRCq0dbwgKCNGGRhnsDhsJ3ISkLkFZ1QZSqqH44b6KIZGC5SQE
RDeJJrt2XUdVnxM5vKtNg2jGSG5rGPLaGSoLQiBzrMK3iM6DuzreuBRePbw8NPvfIoB4MdmWbB1z
tbVcF7zJnBiiAKvd317Kn0LZkHEBGisAsl2oR9B9ix8cVqOYuC/TPBR++RIGeuWDaVYw7T9yE/3f
SAcGZrhSp01DLewSEzXCkxrlP/S/XtdwYW//6k7Y/vJVrffSeClpuKDL2Nt60LzafXfWSM4TNjz1
9UckZiu/6ZVLJNqKt98cxuSKVN5RQRRoWeB9wqPdk4DA9B1bU0r6Qx36gyCjmkmE5+tqUGj0TQ5v
pgWLduwyKUfgnJqaw8BOXOmYfC+4s4oQ/1XKhgZtOjLLr8PGJ5qX6+RY/B6ZdpQWTAi3gQ/i4zu5
qC4YVy5uBCP0SP4EkJFQRiOx0K5FGXAhAmXX8xCMoftVWCXKVSUO+EZqDKEH4ppBsIQ7nhSIG+he
jghJAvG6F12cQ3ReN+Fxpd4/d35sQ2269yfCzfHVcElL54tH2QsPwOSop9XiirLkrAdBEU09x5IL
ZcgqtKKdIgzrZoqXPxzZcoJ8KQawHMk/ImHJpLwmAuNLQlAmvCAXPpdYN/LE5kuzVnxw6p4DWYWg
LEro6v0uoo87cDJGylxDMf299qvYsZ+KscRx1VvU4Boaq0z8s4SuL/hYaACP6gogwoirnsy7B6Ku
B2IH/XiaZvCOFraBSvO35Qrv0KUvc5VRm72ErbmqyMaJA5hN15LzmtBgexQJ6ClcH3nFdCuRMHUB
IJGPPc0rBDdQGjLY9mVpiDR0l4guVNcdYBE6WGTY1HurHeCdJArOpwNTmjExt/zETl0eejXQZHAp
kfQnu4JENqzrSsuuSRND++ISwSipCZvCTENH4glRR1I3Vb1voQkMopKJH2bRUS92ZTCCpc2MbFzN
lyIGm9R4tO3t4xMPOFPqNvdkk5orGIMkn3d5VTQrDm8CE/WCxBT/viDE5KOZL7GxqAPAEQyNl4RV
npPkW7swp9hPRkCrBQPWA+tRbY6qTyVY++jnFABnCv8+vb6rPTYefmBLwT9GuYDr9NcbdnKrienE
jf3VB0CZiQRHzbygc680KtKIIUP91pQ7PE5Ok487sRaWgWOU4cZWOke6Ofq3z1vTQAkLH9H3at/g
gadhvR3tsL6C6tItp7Mh9l/quDz3KGLhH3iM78x9dVaWpAOGIeBnX0fZja0TXeLfm0flt4WivqBQ
g1brINnpvRWDAgr8nhHoPKtvs5LDzxIOkoMsBdDG1K5FSqtu/Qx+XO//0X62ITgioxeu40gYN9oC
rEHFm+ekvfkAIKhIqxvG8Zqk/TP6D6gJtUxsEWt7khnV0aCQ1qXIqHat+VptahN9GLl4f2tPm5Tu
ubyMIEENzcbREgHhb7XXAB+xQrAqyGxARUJnacoE3lgnBHlP0nLtvD1hF63ObhWPA2MkzHbCR7/8
QH3Gqz2tTykekwB0fjWdWUrmk8rcKSrk57/R4GGrLBQcVooH0FKcX1Z8oKi4oYp7gyB6zeN2/s8+
8xCzJ/spt/A+pf1b+6FG/bl17N8/kspgtxpI+kSwv2EA4AtHkIPhu3HBEGYETQaMxOvYTYayCLnO
iiWZH0YAu3SQ6vRsJH+iVAB2mRBeqOVQegp32fX1pRghGPcCUl8Yjbb0EGIHwwtHWOU2CaxnvgbT
hRIs74USaKBaqO6DSi09LGgOWkO7ullo1jq9KNKkDIjsuOuY4+2+MJ49v/Q1jNlT8JkLq20Liirr
JzCucW9mJ83ndQnE0AIm9ltMbJlI20FWmUZxneQ6R2Jz1VLCRam3KtBfBO2F/fAohekJmYBL03IP
iuwhJPmAY9f6CgmJ6wp4SjDlielOCvIXPL/Bu2OIbG/K3g3mX43Za2WRZ7DeDG6IahVv/p1oMEiZ
8pKaC5z6H7JahhqCYkpYWMMhS5KrSPs+co1sPzHNSCWFMdEj+zRymeeK1yQUctww9FTD6Wt4YEdS
so7Br8z5DzqvE//3V1EoKAMnpHMFSOkDB2cZ8feuU7lhNfKfrhn7uL+RQtzCnXAR9ea2+DuuoTPo
sYeDysmC3OrLrdaercAGskgSxdEYIPuwVotnA9szINgSfBX8aMoDiwdpxM5/P+qsa4CBGPFgBHmb
VstQ3ZEA0dHUQWaLqqYdV/juju0YCwx3K35SwMhI/bIgNkVgy04yPjc/SFGpnTOLzlm/r6aAWEEH
/134z1RPCN61VpwPKhiCdlcpwbgslkRu4JR95cSEOJXZl/4G2Su1RPcbdQv5Ds4HHy/ZVYrH2524
woeGtioH6hFLU1W0P0QgFZetqzoBWHHFmXy/SqEBqTOo4N8z2eptc4P2dRizlqa2b/nfGVB1QQGB
q9y5bRqS0qS3lZT7F5VxB+oP1T3gUXD5228hNm0Lie9mrjwQ10i4uvR+cvaCX0Z2TtfhS/8dgIzR
cTcF/MHV9KrW4LMDzmqzQqfEhkcJBrpq3Ut4JnSdX/uri4lUXInacoddE9kyfb9n02RCUqpl57uD
9JL3etZMfa3gTglS5GI7HqRIJ8sDtVMGjHabZF5/DhaYZDcLyitd5QRGDTS1+dyEBTHd0wPGJt2u
63Qr/BrnaeMo0sTGVF1+7jLP0cZ1kAy6ggb8+ckGraJlHcQ/+hnsJb2/39cGRvDur1dYfN0lhDn6
rrNJAR02rK4SL6en6BGYwtL5VLX7Flh1gA/m5VOl32FjTwkd5TzdjGogulozgOCuKaNj9NCny4vT
wpDMH7h00QLhkTTkXBoAtikPz+w0ySo/6dR2ISVSbGM65a+DV5ReobAfcvDe3uCQBNAQDrriVzbN
4PKrpJH63QWd4IJkXg0AU23Rn76varbJtVvFLqR7yk0Y4xr3AHsScVVOhqplMqpIGunB+udz/dKB
ciFOcr6r/ehOrIqw/Scxyv2em89VHw7lI0kU5VIpNjwHlNjuXateKzo4ewlnahP0Nnu9rw0FnP/J
hpNXtyL8MijdNUH5tZL737IMxLZFLkLCzmjIYaYSRTs8wZcfJypT3yVf6uiO4MsE1zEziXsmVycP
x/kp+ph9x/S2wM43gY7qqO/784qiJzz87fw64A1S+Fbc8RZ0Kunl1FVvV4lJhVh5X2MF/XQR52pP
z4Fu0myPqonKsrbo45p7A2WxWm5qtdtJ2JNLSGXh5U5nGEoUeLxZFLWM2cKZTtKgWHKdOJ820amG
iIJjOZwb+i/c++Z2oKynmUBEAu4GE9d6bDcDs0RYrsQXJZVOD8EBsremxOYvOQmGwuphkXQBQSQt
SFLW5hGJ3D6VDLVB5y98BFTHQ5P5q34d0fU+c+psgL01BoN4p7R9PboaJVyqVfDmEMBNcrh5vcOF
g74ujgh7BrhZpI6U3xo/J2qeGGWwhwTxQjiyPXqeYJjMdiTuJ0fmuAfrVL0kbODm5qzAxGq5jGxk
KHuMHr5UGtKvb7NJF0hSsq1ryag6P4mVYNhX248pkYu1qZ50RcfunI2iBjYrOBCelsMVrNDK8+1o
oLRTLxVoMpDgSf7suWhV4FE+hDm1mmc0mFzRRZJ7iiHZWAuCw3e4Vu3DLlWMjgBBHW1TUDSOy39y
NytYtsZ/ey2dYatULl5L2/fHHTe2afOGDvM7UuQ2mfZC3cRMeskuP6JcmoknHDoEYK/JwGYZWJ53
rC756FuTKK4p8BVwbeEds43ExRTNeZ/LhdGX5yVsoTFgXri68PG9t+m+fx2yXJz4ngE+OQfcN3RH
0WsJbWPcZQX9CWtbIErJoy/hkMShVzzIOYOlzlW6clCmNuKDS+Sg3pbG6GDXxZHCVAT+Uq59tawS
ePStUqE6hWt3CP1PSOsnsOpzdungoA2sEGwWvVg+QKMKRZDzFlmAfC7N377PvW7yWjFeULpr2XC1
MK69l7qURZc+TniiRsByLsNb8oukot2lRZHP0Qj0wbJ9UEcgOmRgFTgGqUkaPXro02zHYbUI4HeF
1CSKuKDjX+uYugmrcn74LYVp8UJt/FJqfYJOCZfD72UkOb56KpROe3Hh9M1TwTAkBXXbcUVf/Xna
8KjtL/p1XLajIn+jNBMmvFryBy3wOe/ychbShXXcQrLk/I472y+N2VJpx+jMTjWygQBA0b5j2Joj
UP3UNe2POw5BtDh2vnfZ+MhyeEnDMGw+byFBJELfVebeFLuXDnq5FA6ORY+2mo56go/YEKGDHc5M
ij5DiMdnpgJi98G20PvyAg7JQ3HEKjOeXZ/D2S7RPxD22t0dKLm2R3YwMuPt1pcg21hOcQW2+qa2
LDqyikNKUVA3x6tSHXexq5rSww8WWJKvyr5e3Xg+JyOrdXSjbNWPgdctHeOxzp/iW96gdObRNSUm
kadfDO6nKrMBAuujiD96jNu5rB5ms7EcU/F5NtniuGtXu5irl2BcHqv1NmnCne9ClbXgI1xHz4Wa
I/s0NeoPuxPyHrG6gv7FeX6JjS2161Dz8915gaXsepYucaNuiDxX1Cb9/p/7sIszq9RvAZbmJbn7
qwMmi6rB1NHofSlxD/6x5iXByCWCwMwx7QvFuIc+Fa7WFPSFbIdLL8Qf1ynw8yHKw5r1l+ZcCetT
N7gbyk7Ud3KZ6N57m9kAU15wN8GsFbWYxle8LE0yfi5qwMSuq8IjTxAZeq3exlmwcU2SA+ewOzRw
Ack7AWmoH3MHV7mUVK5wJinOY+hzURMzWkRL3LN5gfQ4gdCPIiwihjuxJccqGuzl72sw4N5NkUyt
yH0vAgGLsh8ieRKSDvXDy1gUBb4AAubKcJjyxTDe7aGc5C84OKVYS7wBrChjLd8GZv3Lzh3exg9j
wbO4/C2zeW2Tvo4WeJ2d/zLRCXujaa6pg/47OejFB+ce9/ECqOhdGVR0L0OYQ8oU7FnaR+gCQBnF
coCYj4GmAkLDZ5RR9CaTExmWT179R77k+7OpxYMUcxZLSkH88skGQZKfqta5VgZeP6KVaJUdRTUg
spDrB+f+6gA5ddObnAzqGJ2X+GIqk+c4M23vmCKQY8hxvGdDXXRD3MnOWSFnPE2NimOUog6sIWSI
i1nzd/ZkMCFUTYnWDIIM3yB27qM0TCDE8Y03HxZweFfIAFN5nKL5eh+CpwwYq0AUCFamrMyN41dk
slc0jU2DPMMprAw6STZtudfFHTbkcg13bMZ+gydLG0ekW7TwndE15QYJw2KNRr9OvnXooIYxspQk
30FkV1bqmbErnyaMqAhAgWhwsmnBS+bCjFqK70mZr+Z0hMPLOIY7NFsLMatupDxFh055/8A4ajBS
dv00YjOUIu1XmXp0gqLGAo2S1NbAd7ySq096t1xDXjpju3GTezijaL2imJXTvSV5sxLcds2O00c4
sqCNNRuWtmcDFtfjsX/kzlsJ3hDJkcvYIvRH3kGgxjDBAgSVOb03XutZxSfnAXfP6LBNhsKToMVF
6FQlSX4Cf0IaZJVP8f+sa87ZgXYuidM+yCy9hCDoKXi83WQnyxXMkjvKbVHe93vtWUkWOjSbYJ/R
u1DH7ICe2lnqkeeEXs1Je7XF0S4jmvRYsVNMI0HJuc7DLD5ydGNpn6TRfkc0Gy8E5zvXXh0KAkWF
jSHI9wHp511qIiEqF9mL6gI6ZjmjQLE1BixyDufKbc/Ovm9EG2MbNqy0loVgVQPZthBGp6pUeQVF
YNpqiOC6YGGHNTC2S/0fY+CELbGaMMHZHrR7wR5pP9osHSpMFvToFKcX7ngQN7UAfEd1Yv9Hr62m
96lwJYwslCNivvpfmDEzCV7esDRXbBcylA0RDtNAnASaU12Aar10srn8jRpJAL+NNo58Q9+LX0YW
h9UtcLfzozt2ct35cimwmLoAtqCQxPZnv2ZWL3V6haSTJkw3OlqJo6/wSDle7gQI6KFtnMVtSDkP
1sH7EufimWenJD//SLkFNF3gkgvdKOXVtvhYsSS7jmBvBMe79ijFKO5yzHEIJLzz3tyWFCe1dMDt
kSsGXtoddQkqR8rUhi/NM/H5itLY8OSXi9rwmtHbesTPzbuxOn2loZBRrFNB7/xL9uzVzRhqOeI9
7vRASLWktuNZ+v83FQES4ScdzBpx2stj2SrMBrAUwLPN3LG5DFl6n5uYcF1hlGX00ONXQqUcof0g
S0md16QRbEVcmUa3yjCQySi6NB7PX5zwyJYux49ANXKGHticryFJvrqd3L4Owh00bhL8rgBY03zf
dErtTJariEwyC0ddw2ktLib4LYuH4EfIWjWVjKvrlVTUHuHEO8n5HlkPoPMoQM2mzaw394A5Na/p
abOnX0w0ZspG+hdChdBOP8mOrRj7hxVP/Hntd/B+oE7IUBpF7SMu1amHM3zfyCJABTb3iBnRdUXW
TIAYURUlGa6yAYpDxDqv0yVBzgAkRERsecz80QA9rK8idAA/0GZ2a+t/Y+bKGAfJIgpWoiv9dydR
EeBvaovkqSks2pL28L93y/wjMFBwfh6q/oY6zo1re7r1k9kuwqNW6xRiVedUV9ejy0LPTnIHOh6H
vjrobiYCtzqhYvR5+53aaZ1Zo03qwh9WrUTKPHt4JwH7wverGRtRTIRRDP0f8i+MZiXdbgPBs249
MUoZEu4/jA7Dt2P849zr3JfK+FOBySoXYefux5eEPp1C5BuAwUzglCFMBf8d0OU8ur2U8MsqDa5T
Ppb1astO96eOKNtPHBDAyvq3PSiaOGf5s+cMITHNGYd+eVVvBeGLc2kCSA1KVgVBbHkTAYtkQLKk
Z37QsB6BZbNWvRNpdsV2r+tu3VqNakOxCh29zGe/fxluPZyU37ccUnxQuHYsO9lSglXY5QbRBjgD
ddCG5DymZcNxhQ3SaLjmevBZTsauoH3gEva/YMhGTFefnmTIOFxxDQaXIH9mWXRW3+1bJrhQQK4A
N3qowu62vUc2cbEyiMhC3B0xwHf16pTALK5s/NofnY1Hu2TbebUYxNIfpjbNIaNhjWHkKksF0wT7
ZF6tDuvtTIkujKR+ZkT2gAa1I33N8OQTV9hyhX1eaS4/EiC38SwAWVDHSW42k9nf1y9lf3C9xc7T
Mb5Ru88EV+pKKreSftELg2QUxyzKQMGaWP6GrebDGNlTUZ/YI5IvyCBNN6+w3s6YLyvmJUZQg0ox
QxwtrwEw+WS2jZcc/4UxQi+SVoCXG6sV8LT4deYCJSYImCBhKr07S4uQVxZijpmAYvFQ0D6PiVfe
OsRqF8Yl8dnC1a11LYwzF8/Qur2gcopf7luiNphz0wBRVDs9lrkhjdnLZARXFJjVU0PHoOYtDMzb
W9zMrOsusVG3hxn4Z7rb0CayEptM7ikMv1TD64BntYeRY1fqXkaVRq5+d0BzYQULB0P7CPbQ5+I9
Glwq5f2k0fQ7gVb/+Xn/N65FZQNR0+v3y2BOg5iTui5mGOilm2czkdn3cazmGHXKUA0ACsSBmBKN
CAAqFD4EXWjJDT15/cE783klPHmHngFULATLedmXzIuRL0nL1ydabAr0P/FoBH74/rD/dzbrrgbk
syzWqbpyukIY54dkPVCIZ1MLkIjf8rZW4NPce3wi2l5pN58hPrcCey6rJ4+xda8JmgH8DLzpUvwK
sk1JrVApzM9p9qoaP9kvWMgbEqFy71gH/AHJcqHpgyLab4xso3Pc6Qx15xgJe7g7+2HwhR6qKtpN
ADPVHIeITfCGy83f3DMPDjNNDFSUmrmIhYMRP0+0mUKkynAM/oRZFI83vBLIMDMlroZJqZ3KOrF3
ZMHz6OB6gs3nNljvKN2BlIbAx+5VdWSv4G+z+A0xKWOWcr17Vu+/hJpgIhpzJTKU6hHmYd07rg1r
0VY7h5qOxQlV4J9XIGEYjMAsrgFJETTpuiv4sFPO7/a+CH/+h8KHAuAC8g8OrN96lXe9TrH8rlxg
UXkvVZ6F3xTAdo1T9xwzaipF/drwrvtm384+PKKuNlE/d0Q79XjZY5AhO5X5X/jAYxiJSKWF1SjG
NZnwxbsnKXeJbp+lFTtmmzU+E2NafbvCXQTA+n9RsWSvsplMUI+qvu6F+Y/8Zg1jUTyFKRc7eLQZ
LdZYONcQGoxnPkVLqYweZkrlhFxjLQyagU0CR2SQ1mtMviI70cZ5B47teoGtS7HwCX3WRcErU7m1
xemRocoU0RfKiMRnJMh+0QpLCBB5MZudc27PAuL/wuaFOmHowNXt6ju32jiJDXpB/2n+nMkTD9Ik
IrbdLz7iS326OpfXsPZtV5cJklVMNr7XKFQCURg+rmQEGdyLzYcffEQdUFUpBkY41n6H5QRl5YYs
KPc9CUbVwF9f4Ue5hTU/m48cJ2UCG0fjBs6gTYjJqfnptGrjb7pjY8ojunlY7MiwTAgOegipPrZQ
hMWYbRF30nFSc+qE4aQWJpKWsKgcot2giNlqTtWIaUO7Hi85mMt4roo8d8RA1xisHkuykRiYdUye
ntu3Rp/sak3QZL2AQm201j3864ijsKfDPtcHIzGI9fqUGew6qBSJSm49FrDVYXD3jQWL+sZd29hV
oufQzENOz118qXfgDA8t3CLxz4rKY/3xSRGItX5h6kS/WWHbr9+TQ3imo34ISweEwsY7uc+GpVG6
pn/QHIrthaAC/OofLXJTm3qhZpVCz1ttrAAgeIyHvfAWXSaKiNCyC4rdvUdD4/Oz5TgyLaOaEoRK
Fq69bzYHAQ0AOj7MXOXTLihiMIO9zpi/AXFWY+bUVeKS4yHrz5KTI9gztgNkqMjDIEeE1txitPl6
zQllgK/OEU22fGuDevTSnnmBzrddQzX76KF2UdGqfdMkfrYE5L6EbwagcZghaEmIzYSRQqCT9UWo
ikzlRR6GVGndINF9yXIhPKYDAK/ICpnDTccpbBlCpwRf0Bdvx3G5H8Dn8KWNcX3fY3BpHwPV6InQ
hwVo0X/efqoAW0gc8AldngR8KCSmG5JYZOwsWkGSlYs1lXzUPT03ohyETCBy2AzebuMy+kLDR4B2
9x/NHhkPCBC014sdAR1+yZ3nzgMO1KGEEPKTR9xlkBOhwdUIJEmZedqcdPfRNtNXj6QJd5+24d4H
y2uGV+q6cZXcfZWcc2sGh9/0ZrEzPeLYFKVhrIKWrk5K0DuD2SNMXRanFLWlsO5eU4u+P3SjD6V4
o8+6cbnht78i1GJaS4JYKMgE4K3OasdpPBzvzKgCTWo1Gy5ReDEVB0rYz5KH2LoIxlr+wCjEIkKV
RAVHU5mluYStifvZ+Jv0yXVLkNVRPONG/EuSfNEYs4hjxc7AlG0oHygiidxpcncVRFN8oqPj6Evc
pUjeq8ixngRBcUOOcJjASv/lZJhqdyTWGYJ2MKTD9eIKp3D7h4uPRCfFmBlyinpmDDPXCCVhgAJR
3PgBGYYzcmDlFdYJZHPdMTNDkOAcytXE6XSoHGDd815v+P5SSn5rvopxY5eYjQ1bR9H7XJ0KFchW
jESvlEHgdOGyN2mSAETMpS9hf2rYg5IkyNx4V8r/4DLvRWPUJcGvYilOp9fHhDgPm/Pn9ZwZFJ82
50RhI2RYo1SYfAR4wPR6pkPjXmbsa8SYqQnm+jX0DEjn+TxXXs7Vi5EHA2Ya7AopabBK2hpcfVzP
Jy/wPv2jfoiKH32KyH7nIQwbacUlXIIO+ffVoF1FBbDAeFMSR16nGmmWNuumOw7qjUSNq/ttQNeg
0eM77X66sVgnzHn1SinyZItzqbxVLbw14zH6ESFaj3xxdb9T5Wmkyiq7MLBSIJXgDkpUy3Zk6H7t
vGT14Kl16FazD8ABqv2p3QPNJhnwhMshAOoKLUVA2F1WkfSTSrAZGZ+QR2BQw/cjin4bP5LBu4GR
d3U+o0+Gj8m4waBg/UrNx+khpf9u3nGTCQro5njnwDzYOZpqDl0zDKkyZNXora31t3Fj1Sz+Mj01
5w7YhqJntUdJQpWFpJgwcbauxsWQBAFbUr0gDELSIN1zO/YUPpe9+QUvkoODuHQ7mxhtniYVkv10
RJqi/WIQxIzJ3fSnO9SDJeZ/yIQ6woVSXN8EG3JLNxIla8nfhwbLpdcLL1VvupIOllTCJh9X97LR
LHJGSE4EHxxRBHhAynpWqt+lCOXOyhY1/oa9iLKXJbBLkM+VE5kVIOGeivYx9wiAs27EwnyFfP4O
qR9b7fXW/wAd4F17Oc5FmtoUCAAxI241cGR/MX9lI+rUnPmNO/odnAQcEo8cIYe6QyTD+LXYNEQa
xA0FqheFbYe7yQLDgrt6DpsFailOFcldyYEixAodhuG2WMfizfs20FU38vTvYt62+mVWQe87B9nr
YtefNBQflYq1JIQo0ygUmwYi31hTkEm6U+7CT+6aA9WTE3YNXnmJMmM80PFP/tu/ZVS69JWeeYCq
86mUXt160W5UQwDaOjZeao9PisJvq88qBLqXbRaCL2DaSsng5hx4xTKQZMB9+tLg9WIjz0kwKwLP
4Rg/+QpHiKWE9i6krCRCzNWqYYye2Fe52/a8zvNSyVAEdysH75m84Hunw+0UdzAP3Hbgqn8ucPxN
cW9xYz/tn5jGInp3AkCDRzkrtk5j9L4FeFRD0/llSyGGC6fNiNYCvauffZmmKG0Qw6O4ZmmInpY9
W9iLPL74EsI0HZQfp//MSW33en86M5hByt0SK72h4JKMbdYV/TelWb5Y6yfqTve3MR7U7fpk4QYQ
CM4ZkNfeNi+gsHdquAwDHON2wGBIQ0p1MBI5yxeb27lHgnWiu6AKlXnLpUKvt5XuQsKPbDrANKSG
hKbokhCUY8lCmavXU5flvLYKoa3aK1fumJ0UoVS2irvhZTZILfERLNVzXNDg09EkvwfY5qfuMshE
mKjfDgko+zLIiZRMzirYLDzr/QxNI+5nJSwOL/u72mMpeixIAB1EMnlnYfjNiYXGjRMJumyyg5tq
U7pV3n9T1VYDqcPFTinhD0X92aH8M1yRinlw7rYJrY0n90+ddbdqPFbY6JthlGuquOnAwCcJ5DHU
jLCJD8oiqkJ1wwDvB4nb2DV8j6kgddb0urerz3GHYuYFCVo6hOdvUlNDekeQ66qtEQ6hp5FaepRr
zY2ooLlCCxe3P7xn+LJQ36tBVau694KDCAJT2qK6kJZRFP7gsjbRBeyFiU61WkS/0nu874OnzZQG
YFZbZ6uMPDfA9ZXcl/EQd1lIIZ0OgJuDpq45AFTfifrAAJxvF3N9eSyHuvcoFheaWGRcdExfeb3P
2ivJx1Nx300/c0VrtsRpYVtxVccSfwNZXRwRR8/einVkd1Dtz73EFvFBizmx8wz3TcXQlkr/h7ru
E5bJMbY+ss8LgiZqE6Qp+0AYV8cU/jWxjprqInoaBydNHOQkzAjLQMub2KAQDZ94tfhF78P6GfVq
qeKVTEkdLIN7q+tYdq2mhY7UlU0V16APOv6LBw3uWS7uifFcKIfY1i651lSTjI6E0gCTYNkhbR3K
txNIdyDLXs8yM5zFBjX0X4kO7qDJjXi9krquN/3p7njJ/Nxgkw4h+j12bFScHlJ5Zn8TIyMjZZvG
iYBi93E7KnO4pT2qZxzPPIbdcelH1GNk/vsDKGjz78UVRe2WG6YVgXXmqUaAcJWMgePVqhHyUVry
4RaqXqk04xqhfNb4DL0wg/Z1nftxseuWR5RRqx0gsEYyp7Z9DOQVpYm2wSfkcl7+UDGeukso/VWA
X3MKq2qeanT6Y4+mvOe+xypWbwuxGpz0wNrlcQzX8vdhI3Ox8ere1QWcjvT8dAINsvUmcFXnBJoe
cZ3CanulZSzZgmCEPjZxtuEE8CzYvb1qxKAPNr3XTvrFy+xImuFi4W2k3sR2mvFjLljX5GigNHUL
m6fSQxzSXugqCzhAWyIYsP7RhjYe3MLaZGMpXSkP/IkCcod7kN4xZBE8G8Kut0E7+8+9XIRKAcib
2poSK/9I0h1BARESbvHM8AkgbnilxtRFASBHQ8ceL+0XBczqXQxTfM+DelyXbVmrW1WNJ4CqNXDc
TbwPF3r4m8ablD2p7RKGqP3L31I3yfWXxRTmFnXmthkQ+IKS9i4C1B28gdJyeWRykCV8svSUZQsA
Ucf2yjSPCxiB45KQXlWnllA394qxZI+Tw6uuxyYwlK5+SnefccukdKU8lhyCOgolOp+/r4FvSP8k
yL6RHRDAkYo2q76TzsC6Pavf7nT9boTPVbJcg5CHapYhh6yjW5o9fsH33Wz6yF7jhCfqQrwTuYC8
GUy55N4rpbnzBjbuelqXXxBLuJ8MzXthTGVZpXB5j6GxMGfW6HTRMLz6wtkLTJP2b/LTvTR7S8Pz
tI+vLTcbD8PIH11tLUKFPoi1NdAH03YVeH+Z0xO4plL95o7H5iMDg3PXjUGxqqYKRCA+B32kuIfV
0lk6HsP2EtcgiFjWsnz8xGlw3tlfjgUtXUCSx+JQWjadEaf8hYsqlB7OpK79yxLDiPAbjQ8RbNPm
xwlEWmg1ctfLRWH4i+ezSqGKZXII2qqrlKtAdLS1LuJSt1urJRgIgmXfzONRKG11ZhHwI5PtQ6ls
iONRJWeS4/wA6f6GWgaJ7oO5e9bjWuwP7SmnaLZYFkVL4nTRKU7YoavcyQ61Bw68x8MtnOA6BYBn
AtA1gev+DdkzhAzgeh85Fr5yXFzFMZk+/nYu40PuPRFWcpiG3/52c5wBogst9ail0smFuZhXW7nr
ymu6HD2q34ZV4g8mw+LSVU2qJ4HXj8vRSjAfVpkBIVXY4OeJpbVsD4OPVrv19V6+pcWBptUn4ACY
1ETtBr9Py5ZfxxNOz2eBhSPVFImK4UB7g0FxWUuXYlxCW1t7C7oapmSmYbDMh8fbotYSzOc8traZ
8SI2MfLYDszrb/zTyeo1w1Ucpt+tZFwlluk3M7GpGER8amEjQ91cy/StNvDppD/g80BWfziVF+ls
uHpNwmTGQ9ZxGz7hgh+xPA5iU8sBI5Um2/eeUzbabrbmHR2JvHQgT9a6arcu50fWTswNJNvhJ7iK
z2L6ThqK15eao68YLRCgfHD/kEO+xefSHmg99xQXG01xK/FUgz76ewtuAdU53jYMTTO34sPUb4HM
C+5MQfua9g1ABrba29JcZtCqvyhlzIwZB3evIhaFmeEJ5WVeirdsRM/vHba7NABYUrm8/IHJWOKV
PyTBOrJJzX0xaDizTGduSlBWReXya5tIYw7eBJox9BbbbinAuQAR/sPB3JGLedk3a2SxCB+CsxH9
kdIj9tvrUVw8BAugbP+TCtR1i8cXoancw7YDLOQSzDXVqo4Hl3Nb+l8B7KoYP3vBaRIpRcQROtwN
eLk2VgW50wOjKpiRyDJCiuwVYpIy3eWZnxZEBVLcjlg3dhg7nLicQkXwm3uIwIM/lgAgjHWOOUiH
nKATe0en0bmVYQt2454ZONBGWrOMhW9iDKFSP94g0ywZghoimb6XH3pQJEVLhQsaytrm7j+BL8vP
IbH5uxzh0aCx8wIWIVt8rIuHfmOEMewmP8QPlJeQJr2Szq62C0+dtE8VxwFlrxCEDTW87w1L6gfd
tCV/DzcGGBdloKrK8Ngr0/lfzKQs+VnyiNz9vReG9KUpKE7fM/QwJ9sZgtkJU79yDNBjw+KXTOS4
CWoDQz8k5WllPxR8JFICd2fiQgvuncDgtdr3bc/75DdF3TVrbBZFIs+ON5PLDljRO8aiAli67omq
tgwoxzsTs8ts1rMwEwzesBj9U2hro6helxCljMzRv+mlDa4XPE1FcLJCD+GDhJKL3JZJCpHSH57H
DvNsp3XlsiPxuRR+Ygqnt3EgIXcKZ9w+vowJ9FfiTnWy9UOjWkbWE3alN/+W4Lf6UoASMNlZa1Gu
DTVi+zTgJQ44pDgdLNC33BP8+XPyt5A6De7tvyIh0AmBq2etaxg+jwFX5Z6/f7mAfizUWdPtwp4k
nvrYsACJevlOiR24/2la1NqKNgrn+83PyDcrnNM9vvUrObvFYZ88HCEOBcLsvIg1Kyd4TxOJN0lD
QZm3hTxC0E88UstHpxjv7rH+xrRNEimsOrX7OOB4GDNkEa5o4geRUW7IKZYqEWhmvIL8rsD0PN52
A8aiywgwOKZh0FimtBn6lY2n0MTmHmh2JtFgK/wzh1kKWbGILsNK9eYkDFU8m86ty7qOcLQmY8gl
O8ptQAtVjJ5N7W4wGzaFixZuVHVsBMp8hO29SvYbUXYBPTTm4LYY1i/vfefbI7g/KbhZ202dZCKH
IqQ2wj0+PzoZC+fXxOaCGIWF5gJP36qDWKVx8h+RFzQBbqXRosUbDOztBaMGrBaAZ6x4yTDX7B0v
bwS6hLDXTAhAb440Jr93ziikE1OsjBmZsP5aNx2kHIGSUmXfDIXWAN0d3kKE+14VrvL+IAZEQgLy
1e1eYkARo/xyZB2984KeJNaPfD02W6w3WF3J9o1XYg3Ik/X/5d6cWGXIN5LRhGISkUuE0hTCXlNf
4wPNVwo0tYAAmCysockkA9LoKZ1ycOI+LYGV4WGzMdUWPsiusWFPo1BWODUl6lXao0X/NTgrIugi
R/4AcCwd9KlHj15oJaWLkTMlRDo53rxq5PqVmXpfZhRzB+/G+j/YZsqm7Rf3TbvjgnqePISVx37y
K6ZEMfemHOKLrhq6yHujPVzcXhQUBl5IAkr0x7aKYTujTKPQ5waltHiZIppvCoo5T6AeIF3YcecI
JHdnbK/GeniEa4aFzDfRxCG/eHRfFB/kjzVL0fedCrpO9fiaUJC3snVqAzEFISNewocn0Y0zvKj8
/Rw/Lpu5Rm/arPFL8t31K7ZltuAovwvHsX7CU7gkqNSebRK8Yw3nTGeHg4sIfauVuSEAnS8VDoBV
TupLgO7UQD9wBXZ5xNuEYf/UEtLDpajiljsxyY+qpbjEiae3gv/sU09ANoSXnGCgrI+QAywfki5Z
pi8WUjyNu1ymu+LvUSklZLRoc9KwL0Ri3U1VcneacXzTKseKuwgpnUeTK5FcxieHFMR3C0rzJ3Ik
d8tGe50YuuEeufDWEKd+NlKeoDFhimgVY/W0beP2EZ3ZPKv4Ymq4Qug2ivrxLaw3tcWD4GTwjz2g
jl+g86ViBFyQhgM+dUED4Hj3a9/DB9haKtLDVNGmWVobKdASJKqMWIBJCJ+GTRG66+Modb8Khzyo
TURN7HB22l91LVosKAz6s401rvnh0+irAJKTIXjdnQGBcOh9fS6Y3Z4+e+mTgKtTEkKGqhJcHeaq
cfDP3vOrAZV0Ra9SXVZ4AzHQpr8ghLD0G7Bd0aCSLJA2jvZeYjrN1XEdgqqZyftOum/c8r/iOLwb
DfEYPtIPyYVSHnLGcOeO40BUbu3besyIgcbpgqjTr2CMGbZeBRT7SMfVm4NhDhgNh5kzVyiy31PW
hxarjRmwX/Gj9QjvXitNWD6c5t7nWTshJXIpvtPtz97AlMZfxtVDQKBmwE01cLrPtQeGqAKvjLlB
OjHOO6agwHFLc2Ng00MJWoro3FEHZg9qeLJU+JCXkHW3fjllQN3wfsltx8GS3h/P23WXhjTT5W4S
lRNJBMqjLawxKgUIPyv7PVondIrGBwxC7g60LcpyGY6IwEd3nICiU1/W9WcRLp1AgIS/3jtc0lxf
kZ+2KPeGMVhKly1gnQLqmDxnhAPDiWGsWTMbKz3uOW+GmiPtNg35dqEnvVpeR8jgNbh2NgARlsjj
LfP2nViyXuRBhuNuEQJNwnOw+gbRFwQ9XKLMn8uOfXSdvOzcBH1CQT7Dv8FHUvwsCNhYX1ovDSER
eFYNjdVWYAwhVo7IR5KSOYilSoVxMqZnp9dxy+sloHIo+4KMfA7OhPewSlzyTt0PPg43QzlBOT9N
jH8dYeSP6Y+qcXRye39GcQGkyYuRX5w10d/+4ZedYzDGH/yO6NcBK2kYvIIS/Br5Tn45f+hiMDg9
YQ5fCaoypkcQyUtmyMZBPmYeCgGkhWS45Ys855JjzQ9dbeijvCwLy3HQ2fwopZ1GRgvGMwMt+sFF
ztqCK67C4cPG13Iu3fFB5JGhpGPdxxcNgPJc9AZZ8yXgxYjHx5EnnHKySXhIZxRxsRvCkfHM6A9P
lHRxqxPJGNa+CIN1fr7gEquUpDysliYDasEHKhX+sLm1V+ZLfoJguPHB6cmfj5HebPsUyhQlGxqq
+/Aw/2U3A5FlRAjCoJbtjUbYKhol6gvBKUQwGmmSXLtzmeqMabBlCr4rtllX1RhD8h7mKqNFYtWX
bDgpFmnZf+Hv4wU3wt5wB2m5yigCykT3Ion2L1FmDP58Hnr5h5KQGWaawWWYbxPNZsihO4bOrxkh
uFXLoQUMrtGTx54P5sYfxSOMncsahnHvuxQwI2osVfrXknYTwmtKugeZAzTiJf/4tjjNYtq+a7KU
AmnXot0YNbPk4f/MuUHblV1GIPgYSfnEmsiVPFRtnvuTSuBjfAIov8CXPcc3+JRtWVmvAQEoy5W4
8wUDXEy8yMwF4JThDousXP44mc9hYfyQT6Nzxuc/fOuq3IjeGDw3dsWip3/OFED1ysG4LfBpuZly
svBdE8GjXau7EZW50iZM3Asq5J9g91uqf7X0A0r7xV1jJiaQlSGY7M1Ij4HNz7KwqSWFMj1pd4r2
RFmzCTf/vApnvj8C7Vm6I7IKXuw9v6SKQ0xc6i1sjCBpn42RdqGm5pAIE0vwaoogOUqhHAyVvdfA
+USGVCg/lGQklrgrS4m7sfF5Ej1H3fplp9W0C2AzDr8cD6Evrya++pFXPAkb+M19yYvm+x6Zs765
8ego+oyv9cd5L0dXIjUNpyDD8GqdAD5sHote25aHdu16S7NP+r5bV4SReDNNWIy27VD09AT6fBaR
RZKhcrgRjccGsNxRefHuXdzu6op0t8NeLGXdkOhm5LoWvOp4/xvU2AcgjJuETmYUipSixQ96nt7K
2ajGNIYMbsxaecSBLIs5ida1D7jIuY2yvLFw7rXlA9NNgij4igmB+qhkmM4WTkJgAtDsTBbQXAgV
/ovNUCLwoCQHM28pOq4i5YLaPWdQC7o9gIuAINPGQY9ZbsscgMP4HXi+XGBAltIgMYRS3rvLhSqC
oOfDx3FJ6gf18Xr4tID9U5z358Iq9ZSQWoLNi+VDKVjlP6OoqhI4vHQwmTctSaZKTJlFilLTr9Jt
5oKr4F1G0Km4uMXzwr72ayh9XRMPhjnn8DggWBMZ4lvmZKqbQovZ46qfUhBMTE3mPK8omqjaA8Ss
Zc4cx/y7ttAaG51RvaRxYnhrodpOaYSb6Q7NGgit6UexxZb/Y9ey1b6+FWzU9PpkS8ksf2GZLaTb
gXrRO20Z3rjJ8ob9sQlwsv0ToH7zmdHh3ACHbw0fyZTwvvGhgS82nbK6DN+MdswQDoGWRkyEL7Ek
DPW8LCyBDJmYqyIGdk70mVNUWqqkX8zOCnINYcLTNxItILbsSuiyHs49n+EXU6CLOamM3sySeuyr
5o6cN3MIuUbl7tsVVG7fSFwQv8kRbS108MEDttcIoQOWJQCaeDn1ptOKiifusNv0gEstoyzTkC9K
vU42ku+/+5eDqr0CAAXEfcQ1yPBJ2nzRyg7w5v5dpSKGQ7EgmN7+kzNSLbyTs9msIVv7TN8AfB8f
t/iw7aLxhL6MekANxn9+GLUUOHrbu8SzHrR3F5ECzjXaUmta449UUaiIznVG+lcEtLZMbgV+gv+4
z66v9TFjMmntJ05ryuKIbMTedM9ft1S3nRQkEhQY/u10cY5fLv8sDzJlXAizZBW1rBJYQZkwoFhs
+L9O7IQYuM4hVUueGmKfMqhNYB7bexnjbdpPNhTYJCu6BDPh2KZ/b6WVkUaTsL9f51Z/tXhgyi9u
JcuFam2i+hoggBQW974fgL51tf+UD1TVqDUkIOXwjhmMPFRhz/FpW14amwtMQgnXNgAZLnyDnDkp
nVGk/E4OkBTcjmnhXoG3Gp3GsIUqNgOtaW6O5afoUIEaO85BeRB3Mnw8kXaHRDIKNMkF4eJ66QBQ
TJ3tbps2s0RAq19VEla6Uwzwvb5r3oV60xRfIvvYKHXUV4foAez/nqT1hKPE0Ieb6gZHZ8Pdiqms
rApgxdOCye/sS2v5XpOV+110wEMqiiuCwe4tcHC+AOb3qO5JgnqEtPiT3m6v2kCt2jaMQzRWa7ML
DgorkYPDZEN5xJ2iAtYOR+s5nmqgGegM9babMSppb/uymrrGjIjySHziuN+GRBMepE19uVlqu9lx
4RPGmFxM7p6EjYevuq3c1qBQXlaGcK8IZm3lUn2Rodc1Lkd06esxcqTe5eEcn5QjxVBnls2gaT/k
gkO3FYI8gyQEqyMJ9IGBD0M2om1HNJUYDL9dmfwO2/oEjEPtJjq1USFBjdNc8duZBqYfXSZhrOZC
5tfpBewIIGKcWioQsw4E/6zHZXrJNMdKG4/nNiuxW+NvqsFWih+9wDhyIVMlbHeylRPkHh1vZ3js
Xt1CXd56wPi6ngYRgwTYxhQryhLeroEq5ECoOzelB6ZXXAOfoal0x/od+avgf/qvdNf2cs+P8rG+
2u1+jLYLyu7Are7t5gemsT4QeCmgTLDB+vT0go4UPBo5rKSLvES2jFc5IfvUE3Hbr5YN8ZMl+5Cx
fM87yxukpZP6G1VPgEn1uBQis/xLC9FneiYDYBUtvnvxMfLKqVXucYKXy4g5oOVyqvYojC5/k5pC
hJbimdA3WI45As/E290ogKZWMGnDJG9nUls/jBh+IC8Ae/W2o5mcXmrrsAzWg9osSxHA+wqxqfTR
PRVh1M83nUHk4xsuWbSTlOceijFwQce5RKAkcC5R5Ofb8oU5hqvagbgtsDIQLppy+hRfM2Re+YCp
ziZwdPT68m1bs//E8VmtpvUhHPAbGIwuK4mZ1uQi5/yZJBn9qeL8cmiTniqDTUNixjK9wclKwlKg
LeD/l905tzpTwku+9nRXp2prk8kbuT/fRPdYxiaM6UTig9yGvwcngM3JoYAB6/t15PFg8jg92bQq
rgeKYr6CDRTX3XKfjZgFv+INsa72s5PyrrkHKOoNz1ExXRtRThYZPFJCA5ha/xh4adwDvId2WXDc
6H2KTHCtnILBvK0ZnAVXrvrG7pKS42EHYFqCzh0SutgmHXIkfVcFO9JRqdJQYPDNVlZ4nIaCnc0T
JNIX5dXAor44uTVCPYAlES1apC21TTk2UfkF/16qiK/lcWxLysSkjONyOoc1udIeYFDHEvc1V5Te
35C06og5xQaNJTS4pCQH9duQMT+LKzh5HE9r4kk+SdbUDau1mGhVPb6C1HkRnE39cCw70qupa5la
0F2NlyanajrqPP25XYNF1dt9kgj9TsKxIsHlw45hvZPhCIpEvrhVCrK13BO13BWgLbx5pHL2Vdr8
IJ07mXJrsChEC0+aUobP/3dGkkpd7xd0R2e8MLLWeBiZRmD93EqoDHkcm4CkGG/WcnL2BreYRDmz
zHs3S1S0czKykQo4gWbSyTMUmIiUSqGGGnHVLA7hdraiCyR34v5dHDSSgbESnw87NSAb6vx4iuc0
hY5Ybb13cG6Ud6SCiWVDiBSup1lCVS6CCxKGWoTQjLmBjBiKDxsbaxeDOcKSTPGmcdapnGJXv76p
56EMiVz2iuvz8NQ1Bf9mEN0Awzm0571FEEp5B98MS5mA/6l3yh8yb7PIoo1/v54H2vaTlTS7+1lf
8fjeegnO5bQUyozrQXoLGXpRx9eD9BVYFhK4C92ruAfqgVZff61CdjsBVV8s+q1a0h7Jqpa4o7MM
KVnoLsTkndMFOGzEFalGtAtL5TcjpTS2i0PVuLJ+f2eJdtHY1kSchGdFQPI8tyfd0e71N5IceOVo
ikfCFolQUR/qr+gkY0edpKCQEfy2Ec1EdkAXD8UPkIw5ZvRXvqUfzrLYFAa+SBg0tcTkMStItYT+
r8PIwRm0wBvQt38/qxfxWpr+RUU9oN4RGT5T8em9yhogrSxWRgK/9qYq1P336X2/b1bGQfWFoYfz
s2T6NIlPIZvlk6umDylFeElzrydDQYbvk4hgGsJqtEPtL0DkZmuhFaI7Oy87BxSXk1GzbtnnbRzs
w78PeNKGVppHzNvDeufcT8N2NMq9iThkr2zIecED+CmsmMYsdWqsPfu3866XdL1QcO7+ciT+Pl+1
FJm5jaJvNrfOaFtwWGXX6fjdFnQLVHZbVKgR23BRdmWfG3oVwr0pl7jDdUb1EoH55pAu+jMZitCM
oMDRvWcK3z3XzCDKd8eewyhzs0fHkdSF3wzJ5FNirTUpmfhiHqsfQA5osFfinKVYE9HMKq6RaZbc
A/c0SAQHYKq/EpXD3ZN5ktvtIEN7FejeloDwjH0uoXY67lKlwQ+KjcaVaTUrg30jQJIusNPeja6c
R4Dy7NwKzn31x3E0nz52vzIne175Fkt/VMbMe/75j5fy0q4ZsSnaox3IVcB0oADOAcSHRjwPGAyJ
EIbbzvXVziqblNpu+NyEB3HtepMTlbbnNL0awFrFlWucQ2DuHHNdklnLN7n/3xE6BoSCT9nsx9Qi
yeE194lNr03bYUgMdTJcLobwP9ypUu4BY5GQLgPPs0+8RMwNf4H8cxDMs6T/vnPCkaPqyUt6NWS4
BivS9C7pXnZ8qMK3S1Gc+6UYpP4VdNABmSbDVfYMPU/zEnngEzh/Joh0AAEqUutIFrPY0wTmuGPf
3g65jjbdSIWvzvIYfbh5aVmsyJm6qgLPV6fP1jdWmx6ihlclvHsMjKW+g/eSzB+dgTK1YIyKJuUx
DXmzqp9hw8C50ptm7HH1IIAQwQwU8kPYXUV2+vI4de5YfgGdRWqMFnUGYvhDrJgB0n9jArcvHjkE
IDvjF22tC+x85v4LQW909h1KFA6ebGdVEUSBXHdZT132SkDZ+tYFMurKRea2YX9/uKbEGOdEggaS
vWT9KXJFrUmvwZIx60Lp8JQRmKMiTLMGW/QnNjmADHqDIZU1318pOwuj4Rvphzd11hW9nmjHnsqh
Xf0Nee0vKtcRc56oOrIMMH1Qnhn6/ONfVa9VA7q4bLnH+oP321SbpdbAQEkgVUQ94tAtypp8hh/e
tCt4yxFwvuP96JO5Y2c9OZd3pySYWPPiEcjXJFWdVGIVhwDlwS5GOBb6pPzVGiQSDcs1Jb3Bltya
vxzIOUaZKYBwY9r8CpXSXarSHhtKdTjBpZnbenkrt998c/dFKbAZLhksBET9/3OEC0eU3rX7u4id
Hmm7Hbe08PLpIGPE2zC1K1W61LjwBXmJER6XUPEXDXjcybdmHNnMklF5byb9cE6hzHcLMehwT0sO
s2YaISqjZeAbTL9iqgFCUxyDxvOnocKABC6EVMsOCWDl4n3oWpYJ1/J/XbLQDRcY8c6isLwvK1B6
tfogF/BqaSlqttW4EgStz3BSvsYYS1ijenXn92BvtNMoARWEQ4TL2d+2pi5iZnoAmXsXnI5AnkGC
U4sWNxoH6+OKNiBga5qOesiBiVmDdetsG3jbSSJO6Hj9ObL9wE6G2PHiEXi3cE51H/iI/194b7Ow
UdfiEJOKSvAe/ridp9UpfQ4usSDj6bkD4cu+wymtFKXrpAOtO3FIzaC/epfe1469jghsZ/7I2gPr
bFAbOdEU50hyUb7fUGP+P5ZcHSObXIOW+r1VgrdwlkBbaPle/rYswGXUtUbBDHSd7yKWuojqVZW/
3TKparFsyzzn39wvnLmoKfRyx5Kym0mzWpwiW8CAAMvn67kbYjfuTqd34AR0OF+taJGLl0GsFCqg
ITj1K//mwF1qaR+VHUUGve3WlOfAjbitlztLU4XA22EbCvKgEbIdkELcslo14NlEgux0ZR5wKaIQ
Yoo0JjI1Ggrvmq0jyxossKHSPUUCcl5SBk5jPSd+wJIah3XoIMhVsNQXNUGxmnskvOdtvCp0H6AU
rrS+xIT0xtRKAaAmxRK9Xu6ZjBK49/6xrQoD+tyU21USPSu5kDLIDWbc5+GNI7uj3htfFEJxfdYb
r5s8lgPwB9ij0N7txiNYxNGj61Wrift1LR6TYUmsQ5yv7RXtJhLwNTEAqG3P6jueBHwYvKbb+Wva
mZZ94Or0VwrYueP6JID8LRNCI+aTpab28CDvutqu9TSXIKGlExDQKBhbakehyPjikGuoz5P03+ad
eGgdStkE1BUXHME0OUdhxNd5hCela9GRgEgfxeXqs6mSpJpIBf91MOGt+nNNKoxANPCuzCA97Jt+
CQCtPvHW/VHyNimEyWPCBXZhkjY5JPkol5AHVoWtm445V5WHUO6eQGA3jzYf6iftmyTPvanelgEo
TtmHbF3CW9KI4/aFRNiijnYRrn3l8Bkmwh10Y1I1DZq1ZWychlDE0i4arubkHTe1nq8W1e8GePj2
rXw0mU7rMjkatPRtopaZ39A84r0wX453njoBGocUW9IfkE7OaIMR/TWcUvmVDcY2Z2RsGkRHE0/2
QKFJjY31Px3POPsHKZGTygfuEaNlvHjojq2fSpT2nzL/mrpQDOpmCgpqjsxIdH9j889k5eQh42qu
/Z4pLBOeI+n3U+//6N3XoVQWLYEA4msmE5ZdFr9gNxyg2SFbsqz05WPzBkwtnPvmppNDWqQRMFhR
5L20unMl31+fRYmdR456kvyRzNBm3ClXgzh+w6wPgPi6yr8QoTN7+JVv6+ReNkkr+U9dX8+Y6rq3
iaq+qNBS6Ny1HtYq7DfwPh/eY1JgNKb8FiyyfJ/K24/bjIVPaGO5mQ/LLS3oityEDnnrlxk9JEs8
eNNw5jIqYBLVdKqsKpKm9WxofhJ8MI+xK6kXE/sDOMaSxG6HdKRj6q5RCY3HB/zDUohQNvflnx6O
cLdwN7ByRf979Cfz2BWOuF3wJZ+pN55DxfC18wnmjf98Y5oKQ/O6MPsVKFGabNBP9+6khQo8P2bw
3wEvYyV5hB73eEpzEzZSD4MEwEaPON4512g1+bHp8LTEqkq8oN4LXdW7+ymEYMmwi/1s3hszFGCe
sm/bg11IId8m0FJt06T2y5DoibwUkhAF3GVzBLHnCGYoEB1codhW1umEsQaTYLshoLTOyeJ3zKUP
4bByRaF/1PeGaQA44a6KuhMkhhuwO16J1OHSj09aj/DTLkNOnQKfw/8gEhkUIMih2HMgkcSjIkwR
5lut7XX4UJT7ilaxN5wTgo5TNiDHyECfDMovZe/22N9Z1lACznqxCaVlM5l/OwTgoJALTO8zPueV
V/8Q0wJT8LcT5MyWXViugK58j5owMIuayhQ6i6AE3rMsamVDZZGH9OL5f19E3pHkoX5/KEYRGNfV
TjittGq/VquJm4cBnNyuWEFX+4dzO5gNAAUmYq6CbNXrHf5TuxAxBalj0rZfuehp/Q0LnIlxRRti
sfqjg+55v15XIA4u14Vhr8XZqmbnQCS6J0OmX5wVnf6Yfvw6UaqsrdJSg+5Rh0btT6Di93f36j21
ZytgrJNvL0qH2NziD9EmCeiIkA3zOLX4WzpZgvckHNHzQHyRAetBbSyeq50ffVBA2jfSneBLKm67
F6UHgA3VPo8/GYBANwtEE0Z0++ieHjr9MFfBrCd1EzmZZl3GOXvCD3NxUuNUpKJHqkY6T1bmPlkT
TpVkpY0XsePNmOZKkhJegk7GNW+NJHakKBU5iOy2Lp7xIwnwc4WotDsevT+1ES383zPBt0cSQQDZ
FfKmD7jJCOGHn0mhcr25ggn7AhkKNZCx0Bb5pNerL2Qzp1frnmqmNkgiLHgQJQsv+Erk7HS+fUmP
XGm3o6AKCVaBejFD7IXo308UZnptIL55SX2hBAmZ/F1MvSpfDZpaFjebJPMtP6s81aLzw2hdTp1l
FwQXOtQVGiepPCaYezZMOVFnh8sg+rbX2C3lc8EH5teMKI7RQp+uln0+PVT4MLAeAINppXKS/3GG
7pO+JT4wUIJkezhYsU3C2sJPP/5FO5Cr0nD5OZkLuS5+skz5JRZR68Jze08LKKTAxSLCpVpp0LxZ
5J8xB3kWMSRbnuu41NvxkhegyUteCbW3Cy3IRKovpL+FXK2q2okTWCLAlCZJCQ0oARize01RoXSD
d+Io56DzD7X6+j3QMtogFKUH8vZQbnopotomv2PGIMTnHCS8J7JIRoUILDOrudebRqjtoflCnfpW
snRKsaUg2/0yR+fPsYuV0WVbluCiScdoOT/3pweL/WTSIm425Iz0+Wa13T6Bn5TPXA/L+phZZ5vP
VcgkrnULpuLmh/XEHMhWkjpNvGQM/PyTV5pmKaATbfX5awSiLRSvmID2veNqcc95ptbJ0YAlGhaS
y9L7mevVMM0M1rDmeV4ksDchJ3MMGhmR0noPguyVX2CG3ZgPksOIHovi3ZUI6jl+hrZMfqbA7kIN
hB/YB/kBnMIy4/1t8+WtC6xX/vqY88Ibjz2kgEdccxvnLm1vHC8ANnje2fspr2xo11GOX5+5fVka
ay0G0a5iRhku4jRHXo/hq2slYme3Kw1/ORSjDJeA6MvH/d/rjaq8+LXy+Thoi3yDZIw5jUUtbi8J
jnTu5H8U0Qn5sIJgprgToNynQIUUatobre/KFMx3JZyQADrg9Ztr0sSFans+ncM0gaB0ORifgM8H
Hej3b3pqW4Owzr13wm0fUQkJfdtVYu0KJjd4nSFQoyDDj/IbfB96Ymw0p7D95LDhVq6Os64d5zYu
2leX+hH18wDyH8EXi2gXp3dw6/U/ZVOgb9th1etqPV1xdsdn8XztqkaLIsrxrbZgrrAdx2VIxHFq
C+CO65m9AMZADxIeXGKbsGsKfN/QTAVmEmpVH/08AEWsxrPkzWVo5GFXMrwayXS4EWnpIsIAEDEP
2s5KFHc79pX7WAMJqA1NsOyCs4F5U1o/n4giz8yPCab3uX8GzqlNWgy1bRjYH6noGxw32Hd3eQmm
5EoWaDSPB4GpQJdl/EGC2eSR5BzEtH49YsUjHN42pabJKBOEf5BQrKexgS4Te829FA9l5P19iW22
/6zxN0Ko9+Tl7p5UnEn/LBnkpo69NKrOdAx2ysbwhlC/3IOUA+YfMPOxK4vkRgfUC5uHJ2Q0gUJ0
Gv77MHUUsBBXFW7k6kQfLNzg/Wc/7lmHPSY1b1eR3P+dJm5MyluGXTrNelNl/pd9NZY6WEtDLlTw
hMOr+4UENCj+JZjR2Mjd2EM+IERpjHSGrijywmBYyf9r3HNgTci/0n3BH8/i0NHPvbIFyAmJS1tq
1JTc94nuZ5/x2lXRVLSBMMv7aQHuAkZHsldjM0sEjuQRtUAdWug3dtwTUErznpW3/M0BZFX/TiwK
18D3pz6Z/BUfNGWiyFp0E9KFaogX3o4S//MPiKv9J3b/SLTa7RlhPk2UeaVmsiKhzTDuFb/I/T5d
Hvous45u0zqfGgNMkRDkoQeo0P2cXOwB3AwO4OQ8AgtZ7jNBC+xDn+ZEUfEzWXBYtychwItxjHy0
xjJSyWbwRPqrNq2OZmcif1UfADuxyvwc+ZDJJPxcjF4a0VVkvSFf/idoxiR5Nk0c/tzwq0J9SX88
oJdmFtnGdR05XjyC+EAZGdYXkPusAB3nfjFM/3RajKqYORFLZQP7bCADjEPXENN7BEVPbfJCOhPB
bPn9ER/Jc40vgnxlgoeYZqGpLxB/H6lvLX1fsm+Bm5hkQCXjlbGU7IPjg0NttVJZZmjnOV4kmTGL
EfEH8zKIDD8fq87v8TslQfZ2/kAobWTk9xwfQbFFgHHvbFOaDKVaMCrwD/s0IU+JlsyaVUIs8qIr
cMmaAbCY8s3XYXDkfF8iJLJWT6ei/zbE3n2NWKPIDk8lQuFkiJj0C+O0CRXhias4uCiFjJvpJRMU
KtZQzWYmiiOFtaqm3yicLdsiIaysWKU4DRUgSISWkGGY4S7a+JeHb7BqwsW6AbLciZLfFpAgrmFx
LsOURAv9FNjoE/Qv3LFp36BSzPm8X5gkYmnava7eF3mYs4Vj+ifLEipupHIzxYkG8pUX7U18bq9Z
kR+pxUKnHFdA7oXE0UHD4UGFMiBRFjx4Tw3k2EdaNJlMRj9Q0YwVNbBq4PnzOX/PWKVqRKVpF6IP
uwHYKHqXYTcmiPNO61ZQBjuEgExzbLC8Nll4JCN1OcPUEvMQ+jSP6u33wT+Pd3LwmTXI2lE+gw3X
71DReOe/T/Cc9Gg94FWc0T4QeCMAxCp+gHaCEsSrrXtAF1mk0QTtnWCXmw+X0kNrH37NWM39UQ8p
V+MIjhpuH0Xpd09ZGpCnSCtPdjY41AeisF6Tn1iaJxurNXROmCp9ySKZ3SHWeR3oOUJKcr2fCh6i
kvs7oVKDVCC0zXOzZYhtFVfaKyoPaxMdAoQLidY+z6etmY4trqLF0NrO6fkiWbv4WxeneuqBR1/k
mZK+lB7uvTUf5BdEJMXeYlMhD4ulm4pXz+GotRpnosI0I/ncbInQXsQpmvkaOg3UAwV6+W0koMRV
xE92JWn45DL2/bmFlivkCaWa3jYwiiQq27jQ13GKbvmIt6pjG81XnrKjmXsy2P0XshCrfSwf2Ozd
ZFEmP6IhX3uweRk4tYDcXoQVxD9K/AZB4swJTJE3/oCS6rAGeGR+L/swXggI8GF+Pm/Ww7mXf+pd
6X+aXvHRupLoVBTrp/tN9J8uLPJyENQ/Qs5tdanduhJA/FAFLP+u5+BPpgvNj9GFUCa/twEDDoar
84/9JoV9rrNiVH4HOfm+1PaUw8xMVvVVqKWYXLb9NN40MdUA3tkqptfag8K9Kb1aDHZWtHMP9OCo
hRnWXWoi0Fpdf8EGWhsB4R5BORSsObP+n7Sstif1lHmLHjBIqr5JeWVcFaXY56gOcMba14Fcd5KU
KuZQedbcyQJ/Regs9xPCPcFYoV6qQIkumGB5x5n79TWyo2YwXROKVOkJbLu021Ln7HpXgqE5MJGD
j2zy5SFAuMfWKMDo3LRxT3SiyOWlICdWAVjJYXEkQCxsRlHODALOIMehJediza4zTokg4XhqNN/E
HLFtZA9gszRiGdmuBQhvo1DTegv8oYQvnii8Yx+ffSlGxGCMiuXAsgoBQ9LEsSvAYHnX+/U2coQF
nEIkfWDo7mO5cw9FPwbSQG3VboSWCeXK5yzqK/G8uJsdtD5GrJ1IUsFwe8jCt2C9dL7x5eOpNGiK
ya5WTVeHEIKKwz7P6INbiuiidGP4m/rz3yPR6A4lU3isFAmsTNkPe83zA6vjLYLFWnvQGmXyKULa
dP9PGXbGTgCcK7vefObkx0D36duXoNmuqO/phXm2/QFR0Wi/XRzja4HcH5MFQxaDUlMsmQoqtT1s
P7FCN8U3k3/KS/yyDUE1qO8tfmbzBrIOO+huAXCYRgKOSx8cxWTWlzZc4keTtahfX3jsUJ7+NPNP
fJaNi5HTnbQ+Lx0UGegrJI7jt2PtnLXViKcChsTgvdHr+/a0Jk/w32RcoERYhTRAzTlVnttMp/WY
y15va4fqZZX2ArL2opB+uPUFQRG5isBD/orHah0I8/mRV1iLC36WgiBpO/CChb2Qtt1SrVFlc5Eb
lQp6y+QPWiYEDdU2+tDC0ZZaO13/9hiqJm/vfbiC39s4m3xvsXEWm24yPtrJkXEsAUUcIesZeJ0M
gq2rbxAggmjtuiOOr3yT5zkDwfp4QTV7rxogXIOlibjI2A+ou6jxk7SuWwl5JzFI/hLLbBFtSgGq
YstLbmAV38uLVoh+/ARRjK9FWGCD2PUIctRwAz63V7LFzMw/islN4goEno2H2obFRyCd8CK3GSqk
ORTHfE4RdRDxrgWV/Y5SrHV4Y1R7sMx8xJwUZV26bRFoaYyRJ9FziZWm5N+ZZ6othOK/0nE7oXRI
Xx0FrfARSRNlasQel/GiB8Sjjh4RvhJ9Mm9Xo/VJKoF739q22yWD2MS5b8KkrQ5GwQ5AR5f63OzJ
mWNzrbICd2PBrJm9+fg9k1jEmpqqXHf8VW0Ygk753viqjhRqoo7VX3BrgQ68n3cpJRcQlhlgIn0+
1G4OPOeuoopmAW1Zduq6YuUK2m5pDfePAE3jpO4v5qZc2oR9JAhFKsCQ4dOmEdUX1A7j5cS9MsSn
tk1eeRud1vBG6Lmmn2FX/+8N0PdgeI9Ad78BPC3dMuRGhucfuqc9z9CcG3pMqmdmBEasYshnIxQY
7ij6FBxMoej4KksU/ySD/Muq7TcHL44//GA1+5NbGtz/cr6pjxgl8oTKCc3WLwIJ8VW3RL8UkQVW
K6mWWNgMBhEpeaZRYbEKpVH7lEqjVfk5eTilvfDPREeSURjn76H5OS+zKJZAGUYo2iDh0xTQw7SK
if9PXWu369wco40X3WeH6L/ijdcwJOrlN48NIUBPkGlaKhA7qbPCCfIh7zxi0c5EIhPJBzFqApGb
0sDNseianmxtyUJuH27wX2QvzaUQinG9FkxrsVeeyj9RJQ8hI8dgSdgdu52tI039Bo0u0qzqywgz
MRYI5Hy9/GHyYOgSD6fcMMaQP3iJQ+5XLchc4fGGnImDwWhweNw5WLL5v9dtYfsNjZ+hCE3RW41R
DfSNzc/6QYZUT6yngz96cmQrlQttEztVVJQ0/A94SYsdgEcdnuaIW8W0WRv++OAMD0O5vGDdXeCt
K8yneWvSLttYOWxwqRESOuLXPkO3tWxdDILTKvqyDqUkwpE/GqoadCETpQjBHV/bp3ThP9guPdQc
OkzpCEc8Dkr1KvbN+RIJbbJSnGsPucwDzyT1lSz9szM31IMmIM4sqzwwz0mmPxkttiIvnKtpuBPr
sSG3JS33Um0PnbVEZkuv4irPf5V02M5arlgTRXjlG6QRSpLn1IxHxxtZ+HpnrkX4PLKGNA4HpsAF
XXdZtmdfE0JmUtk41KLpwNOOlwuBnC1/aZh/le1usYguf5PFjk6McBm4msP53Fv12udRRyQjQUlW
8OH9OnTV9zmAeqwJ89klyF1vue8H+bAdRoVnbioDqUPAjFrvkdNeXr9ERTQ4oO72kz8QKbnF9Hgt
+EBiqS04gwsrmLHByhhoisu2RWOI7CUBK3Izop90wa3RsKCzYQ05dsFNoG/jc+CqqqSbTUA4NldJ
r2LATcBiM4gDnRVbw4zjCRlXIZQSI6Wz3oIAJv72dTxguXYS9M+/bX8dKOsOLGF2acJE9RbJBhFO
qWoQaqin2LqCELyoCz7QpVQHnO27BLSBZOPzmTSiA3m6u85qwawKKDZMs9+eXjCIe1N9XpM6DghM
S4W3/OkKe1zHnn6RdG4fPddDRO/I1mnjLO3iAz7s/6RhW7lmKRikT+c6FMhvAdA/vcwGFp4J+tcJ
Mb6KglLnF0BwGHCMfPh0TfbYCWLENm/gA+nNw8HtsJsdXJMmILbsVLipPOPyhbq05OCegMGOkEiL
0zk5HwuCOZ0+4KyGqFyskmtwvHy67oL3c37sN0NE/aZMwRI183gF1y0IA7eHUP2Y+fJkxqAaK/wN
wznho7Qyh9BSvonKgbhObsqvvzINRnat5PwR0OaNnuc0Z6nfVGrJ5jzUywS4Drb3G5ET5eYAWufv
GIUjimpxmed60TcS8rSJeAJS/a4sJW4cvsUKpTos5x7fX2wVWOVls7XdTp/XrSSsjqeA+NV5jwMP
yNFxmYTMvmzFulbdDdP5+uMhZ1VSe0dqH4XIbOapfpCR1+0Cuhn37/daqaaw8JRz8nHhN6DZASmY
wHWMNAIptF3uP6W0Ia6kp1Za/R5vohRhHrjQ6SS/3UhCEYgibxnY0ORIuBXX8VeE87dswGpkm7hv
XGlRo9VQOukaQC5zUW5dxQh9JSi3tzv7JxEsqmdIunFFj1RmL3jqLpk/WGFfywFbpog0RGPRitWN
cL4s4s7RFPMeXzDWI9Wxg8WobiYh+m3j5ymIA/LanF/TLkOOG2i1W6vSP4Odjot18vKAyJ3evp4b
q7891p66MYEHxNHKy8CrffYZoM8ukLzYYljSfhyM63oRPzpz+pNYzD88f/FQQoASo/LXAbWo8VH9
+ic89O49ifN1E3Bjk2f6jgJ/3sBhvA6GrCrzcHBHe6eqXxcIk+B6Qb8iFdaJ+zf/4Y9kqIMIF9hR
BHysebfnTYTcE/heZtEMq6Kx1WvaX/UXRRA++GHiphP++1mIhIFYtiTPtxXJ8zRtSFDkwMRiuv0/
BnZ9cLoAVgFz+mnmcaZZ6NB7xMQWG1PvbU2t67hA7X+UxqDqzcBUX/6xI3RFhzIX9yEC0O+SXUyq
ZZ62gze1x16WJJlpi3y2ff8oum3pF5P2KeXUHQEfQzX+wgIf0T0oHKDFVxqPOiBUwt8egbKvqIPd
zGohsjym+lTNFHk4HlAfySawLrPKvsXsM85GqLVssgfnuR+zbhJUCfChgp67/tZFIaRi6wDlq1si
7lQXfGAKLm6xqMBL0rS6R/rBllNWem3Zeo9oM1BG/1PQO8nP571nKpXAC0Ea4nBoGxKbe5ke5Yjr
Djzu2fLOndUO+AiKhJEeEEhgW4eE3GOF4OnyWVQqgJXaqbwctoNeKs8jM5gy3iQJDCWhhHD+LQsm
TaPcI+kVlVD/Pt+G7REIqDa6WP8rgOOkwD0R8+PrC6VntngS3U8W6NoAMv8scF/g+lhjpYvFVT6C
VElySyELu0+iHYxyv4iEpKLUVRdmanKR6I/X2x7OLPQslfuXhwal4r+Tc5RqrSSFNetUtvnCEkWm
G1iUj+ATiJlyLyDMOFi8ux+H6JZdhKJcWBuTf/nPNAZ0x7DA8GFQrRCOQiJS2gtKgB3tAw3xrdhK
UgLQWwg6ZiQqeEGrPLfu4EuTcWznTvhwIpypp/QT5qRY1lrd44rFpjazktY9gjMmbzjE1B38bn0Z
UbuDCDCvbjCUFL3JY2pHKkc1agsBkcek3gMu1LYKWIXeF0+qhDJq2InfhQUHizUphtUbjK28t1NZ
vqCrkdIWynbdxbSKBWQBZGVYbeXlyNioqjcTdAG2r6I4fxt6xTRwD8SrrBubzaANi95LXCkZSO+Z
T3+DHQaWmaTkCcdXmJCrqJhiK2uI0wlAO441wawjGCdmc0Y6eiRTgAXMbYkIM5mgrxZxVe+X/z54
XY+CeCo4H9pjJB9z1T4xcZy0noN1oFp4ISHi/79Y9JSKtBjMTSyUhIRDdu3mpbjJHavBze8rdK0T
FIgZcImVKhmEgjcZ0xFxPXWeV5coLen8mf7JCQXCNzKXEWtUe1xbwV+RMDRBLofTRDJ86AqGUala
+Zw8tl2Usc5LIJVp7eC36fyyqcT9XzTqbOCrHr54nVb2w5lpVzBizE5i8n2wRnP2CygztpTgfCH8
2jtyV621G+RvfPj+d3+hfMy01kUCDPYOlVqB4MT5YDoaDlgiF9abErHA8S7tvLrUDslPbeHxoset
xEht3I+z3HieBQKmA+AKczg8qy/yTYH2j3e+NinW3v3EaxrMIVF+CBBszYBevQd1/txYHRxaiUOi
R/2XdyUwtlaHaNnRGw+lA+94KdU1NlBSdKhgwi4zhgHmJ5hBSHOePm47U0qFEUTgX2kHofjpJaRe
dz6lLAzfGZ1W3xJJhVQBiI2Q8nkFjr7hEV/hJU+H2nL6jacmfdC/RWddl4LXb+0yaRxbXIuKHxBR
RMzFiQHIEhu+KZ9cmlVXa5k7AUveYYs7YmtlGyQgNtv+4++I9W7GFySd69Rz6BobXx14sOb4SaZr
9JV0ki8sMHQB8ByGQhvNhVrB0OFOEREt1/dbGwcESHTYEIO0/keeI7a9nBiHKFNNjzvQ/gbLgt+D
ZRHf/w7EkN8NQ9IIJtPPDEpRi8g6mnBj4BuoatvtwjnugjeLOP7tMnBHUYkdiA0pcNDFZ3uHBb18
gRqnI48V4K8r+mg/Xu3MzuwI2o0eXVopOleXhWfz+2Lmra0+W6UgTULCf9RVa4n9Pe2FYXXWbM/A
LMVTa3Bo7GYxeNGBPC2nyD+vIgIR+w8CDNlAfPmrZAO1G97AQ/bKSVvli+zFtU1uD7326pIsC4D7
EucBooC0SOGPAiN8T0rDk4QDrdyHJ6b6l2R6GGifT4vVauQllVdfw124SP2dg6Yi05LMpIXgyFSi
yUJx9EmpqBc/UNp4RCZ59RYD0Wfr27iJM9LpTSZQo9BkX9zWz9ETK91SR5Mas84z85Kun/lmemGi
R4RDdKoBpMUSQ2VuWy1/hBmLB4yhSST3MdTV8hyEBAV8xJeEDg3ecG8UKA8PDlWrq8emKt8Szv1l
WqPNUJVl6CUocDR2SBckIyma8ZKxpEkiOEDjYxchDovx86ueNXT64IaIqTETk8gpsEzyYs7m+xnA
8VSImDEF3UnOkhBsLp94nSiCcmNGRQg6W6g90taL4DrRp8bP+IdtcTBxFWqAgsjJJY+QMX3wAMmz
dTrrCpz/9eMIJE+Rv5feCUUWwhZSWnqQc9GffcWv1KRaiMmdggyXdaCCVqMnYQzggCRSV8/5SD7B
GrbBqkM8+KZPVBQ+1mDiinRMwoQSIlMVnIgemfDI4Jf0FQbwFWl/kvufhsvubsGUqc7DKuCwKu/R
yp2lJ8tkBj238jDlk1hao0Cry/qD1s05jMIoQMYezV28EenHQh/XpEtHnbm9gpDBOriILQFgWjhb
9CBaDrYfPbPIOnKWpzGXaV1TjoeN7gMMpUeSDfxknOQlonrq+wm1uQO4ygG+T6Zla32p2yFQZP4z
3MJmQgZlxO02H//bdxDaNI5DRuxDD229xBTvbr3RGnf6fh/rgNWSexF5bJgS6+41eVywyvcj4fyJ
eDLxYyFEH6BuH0Tjkgs0yH5nt/qcDRrVkOU2vaPfJrJVgRHG2hmPoPXI4HkC/KvvL3NpKcmH2MZn
LAy5iTQVfBhNAEuJ83eanfPGDew3ryPEK0X7hHsvGM/VFoHhJq1Zw6DLKgE6X3JxohCHUOsSnM4F
Vg2mK54ccmhJNyIibCDmgWUzAPt49VpD4fX3yf5XBMor3flN4lu4zMndVZFzmdYHPhK/61i2gM+9
if/ut1/7A/xDQ8T2svqS9BF2oZlWZLWSnhTUJQdAm8OLk+clYmmmkWnSsKJF/RM/+H2Ok3Q/LR+/
SA9j1GKIKVSrBRYb4aw8z5TA14DSxy2KlOVCJLmNDRn8zancYPPp3X/EQFP362ZEtrL51AKQYCTo
MsPXKB2BRow7cBHUyzmDMFEUjrOtANb3AbksUT8Z6SK8eiaXTocevrlp+EdtgoGGhZF/GRz1BazP
em/LULobRpyJRC2E9zcqbJVTIJz9z7P/csrb/ZCEE3Yhh1bTYSzOunIYAnaXneSZAnndtmtIKyiH
e8QLp2tLolFrWS5ER4n3ASYLpoLRZlMqUBCnt7sGCZxOL6RBs86sTU9oseffwKOhJZrBvDeYG6qi
tR26ZUXwxJT4veluku37keRAQiRDY/Chletp+n3nCYTJfsz82M+RwS1V51+0FD9FLVn9zv0I+B4y
Q70IqZLyR8kexp/N+7XFXQxXTprLjHRnOhq3CyH9p4VlFlzjh3uoQBFqWV8gXl+25WGjp7lYpf6G
D1NmAU1e+6gr5rw+ELLmSTKqu+P/JOgqAjIIuPGylXLsaNl0wULUCPGX0BlLWVRIiwYOfXuvuAc+
fOXEDjo0X6AN3UVYTC3E2RD73Eh0BdtSyH7rnJeiZJZ/SHw28tqjJCICxYGAd+3v3Gd2bYMe2lRN
0EVMdeEFQVA5BGenuC2R/8GytdcoiOsVWx7aW04GssxnquiDX/hZG0/nmzQb/FsoH1ihpsX0u0Am
vX78Rhaob1Yq91YSr3OONA2QSRwOYBpdv4qilMnSAgNrqaLAGJaY18DUZn5CT9O3a0Q4cmhUvJAr
mpBLzDIq0qQSGcQorT4QlZQyfSBYjfSFEHtImFyQ9qvkVpcRUK6EtrbwcDWGUwLPh6W7FW8Mu1cx
Oa7PnOflp1KQfB4N0ECAPQOwBo8V21GfvqYEzFSqDQo7uXFNs58BmOoBWXQ9t9yuVY4Fr6qzUxi1
5sy6YiaMN23GviYqCxrPQhL44uz/Fzgbiec1CpImc/PVgLVCfULGRAc+owk0Uz34pNR04Qfqblyd
rQ7XmGwy1hAekeq8L5njuJnUI0s3QuipQzqYP5wZq1/I8wLosHpvlroyY5YTXl85ZZJD7FSORwTz
opgASf/rdDZWJqTuZbiJK81L0PlsAVQ6LcFANgVeDYeFMEPQlHGzCvkZqQHSGD9KDqgq9gMOgCdD
46eYHJVfr8Ipd8Wdrp9wB77tKEa7RN/c+MA5Um6XjQsZFG2CJCrCUbzZGu9vz+vajqb8pHK15tVb
fR+K0Sub6YbyaXzXSu/ZBjPQnOZ4KsdfP1k0HFsoczYHFt1wQaM6pYSR3vjzdeIZIL4edH7d1H1d
fJR7okWDlUTlfCbtdwaJyQU4rg82W3iUu2EB/sv1Oq4z/HJhZ6itieVxoV9/d8KfSdnaZHq6AsuO
/ub86LyJorD4fcDBibbxLBMoBCFGhEM2CfcE/w7G8h/l77baTymjuobpfrrUvQ2MeDglFDX2jdqM
aDwxjsMDaopAJQuHentF7PdXQWyMj5D/PkYUEFoDIGBhkqX2Av6zaVdF2d8Ij+S70bRdoqeLE6WR
bHjfd9xTxBNRUjetuDO3i+MqiEKpI58njqrHwHcpMEkPDxfWLsl18SalzxJwrZ6F6KzuNj0t4loN
Zsi77pK6hMX1M+eurTEb+pFLe589/eHf1OxWXALdhLnOTN2XZCGQOQfoti977xhR1hi9LESQ8Xpp
QSv3BGqgVgo4dWKxC52NbK6JpbJhp3Q76zw9oaXiOClYctFbtJ5doezZDa/PK1s4TSfpmXvlAYj9
hnUaCZ4FPw1X9cuNYRBAaOGFV7L6KwdhL/TMcjJpFYxti2+TTnNWDCHNMHVrW/IqLlb/TCwLGmVz
X8/Jbih5CxzjM9LbUICObsce0DAgnmir2jJx1ob84Uavhp+aQYYY7J5sycTJx3xXKddO62BMkVUS
sWkTqNqJ1OGZlR1Px+SMvxt53pqYJSUDU0XCBvAgZVkM7q+117AUrzj5kqL3vkeNOKPP6dhFf00B
S2JDSsiU/ZxYz7AbCkbe0d+akiYj74aLRFJvLYaOsRmiyyg7T2GKoyz5g0emJxoU1lnYCsJmt6sg
kWvRt/6ao3De8pdSZ6BRgEsM1zDg3QG0Wr7x+kcNjeYSUJxEoR8DrHwJ+11xFRrGv7ShicoYGETV
jUKmD4vu6zglGRJq4ZbYxW+0kkOtXxEAsBkgF0URckzKqrZ+HrZnUzcOCpRJcVDU4jpSVE7kRDFS
h0rN6NgCgTSaCFbgZlbSfdZxqGO3GaFFtSafYrLACpHAe0OogXmJN2l1xrFIjk7mDueTP9UYY1cq
fuRtSNE4HmYWUqxoLqyS4kZqSWzwN8swoM6g08BnOPh7aL8EzfH1YI+VUPeDKlCvZdUrKCeNawGO
6NuXY4V0bAvPJb/+ZmV3r89UWkJOm9Icm1qYHfE5z6j8Jguxv5uWZ5xOXXnWHSXuztODjbSeI7D5
A+hlAy1nXHA+Mp2Bpkaqsxzpciriar/3d67zh65sT6kuQb7fZL77TVIyBW/001CB0F8oTrNB1je1
CEKeiBVIyBi/wtu1aPtJx+zBbV36Hso2DBsOB9rudr4YLTu163eddthQjZm1yAs9ou5NlStcmNWt
LCGbXCPpQz4G3maN0H7ikIhI8ORPj3UEN8CHKAKn3BP+WzFkjolfupbrslXxH2Ioj+IJhILmXq/T
UX5bVm8LIccsZCgLHc4CLfcc5psSu6iTj1MIkLpW+hsRzZktvzb9Jd0mRK2Fm12jRQZTvY9PkSol
Xqkyikp6EKOAfSeD7FOUzwIHmJFiEGrN3jSskMk0KMr3Ma8bijMfev8ykpq+jEyUeExVx3npSvCx
k6jvogVrFyDWS+8y/BjWf8A8nOKDoRh6QuSTnSpAjaMaTMou5WeyZhFNOKSKSVluRwMWBAi98YDD
xFS432OITtsL8je8Vbh6mOUxhx97YGlNpTtVVbPBi8imxEu9x9VSQLl3QTpuFRVsl5CoIlpghAOn
VMTvfbeUlV3f0tL0J2nxpFcQFmmbbFK3QDdMzihgSZivl5WAf9xGdJ9ErwHxbaaQOlHOXoMcR8km
CsKx6BDPudrEECQwSEvIYQnNsjVcJSVp1u+xuM129HJDbqqnngCTZFP89ksWgygaxTvJwUeO8sFE
kr0J4aDCZir1uDKEtJzEkncp64DgV57BD99g7qai/ldZg414CyR/BetQ8T04EJFSgKhCUncxfgKW
iBZCcrnK/8gjG2soMnW1kic8H+4C83+yxoas4P0s52DhdNIAoRML5Gne8zi0DuNBcyZaFzagsAGU
S7GG9aXSaPdZATIYykrukiu3fC99kMs01iLXu3ajOnTCevLrEbysB3KXsZVMGSPplwrsA7bnfoUJ
rmF4IDlj/nUwgc6I/+tf/LbNFp8rasjqpwqTtx9Ca8yjVTxjrXALLOUC0PymTkMBYG0b7HAScJm1
z0G1EU3vzczdWnBkIaA7fqEQHvruItVeX9NKEBQ5xNog1NfWnW7uVClFo6l+7DW1lH2Fd8hRKQoc
82Slg7KL3xeGiZ04+cgcWUL2MUxAvyRmL6BiGtKiSCgHQZ2Aao33X1W1EtTHxx/O0cYTZCx2vJd0
Zee+G14o1Mkz2H2MdsovhjvSJcx/Jq3QFVMc8dsrPq7gvc/u+oawFSrsByN+L37cF/BX+b16H5VN
KlqIOp6ezROT2WpEmUCslwQUP0jI/bFJlCQEynfBlSg0TUaYSFwnC+JNTPKhrFoE+USs4Jcn12Nq
7fY9ju6CpdHpWw7pbBxe8/ui3WWnDftLb2tL+q66ZuHpXeFzbPte5uRMiF8du1SfX+6UgFl6oRxK
/0fdmT+nRMVYVMKCAlttOObduvZAyFbpsgzD39BXlEoYG/cpDHyRwZoL/xa9G6glGN6L0KSUqUo4
NUx9w9QpC5ifoIb9gyCednrL/ojR9W/1YTeP7JNPCVFcZSGKEnhu19/7IZrDOHSRBn0ZUkX7pebe
DPa+A4RftULomFBRxUhcO3G4DL/NSu6WX4is9aFUwWp8KKVGw9SDSWfCjdAAPUxojZcDILlBBG0G
KYBv+6p9enldYsnv+Y05GqztAesnoan3U5LRteRKmXq6KtBVUjjRilAcMlRun9vmh8kbjLYXL2wl
TEDUenC6JSJNkl4mUEO3/59BBT3DFuRefQfNl/Adyv+FriKPdv/j02BU2+gkMNmsaBzzylJ7MYZs
9d3w/LYk4oPpaOPI/+nXfz1LFi7Jgh7xZB4U2PBwqF/UJjbgRYk/tv06MmlKOXCgg9VkRU5K7s7h
PbP2NUAT4v3fPLdBwV3LebCMZi3uuaNbWBtsyeIft/SvazvbF25gHVF+YlRPSZW9K1LCtJ9Wc7bp
MKvUI7Vg/0bCBoSmlpW9ZZWd2yElnYSLLLOesQqK2uQ827rCFgAAGELVh31EjXpG/25cJG4dTbG3
0SmzrCwKgVCNiTGyCPgLio8+jd3xO9Cb+iR8k1Zt5xjjv1RCdP0k6OrB6hu+0tc+p3IvKFBybQVh
9BRa5Q7bcwUwByKzl4oktrlzpS4u5hfY+pJdvzHyeasBo+vAEFZl7Pr7v1v9M01KLR/LQo8X0RoV
grHgQNO3uj2K6+b8LtI19G89bvxeuyD6gAwSCW1HgEoRJwkv6YeftZATLJRRFqnX1AxiEpklZQRI
SBw8t0E6VtADQhOcu0QPFbw7t1ANd/4avtt2ffYr+fLCiI+Bqr7z2FTsb5aL8v30am3S8uvw+vU7
BFCu8DUR9tz2/9JLvDZDlHFIxGPWWDU28URULP0csv8aTZ2gG8AKFz7595Sr4IrZQdHgkdteHCr+
I+PFjrRHKOyGczry3vU3G5Ongc0F1fh+q96YmxbOTQzHs7IrAgzZTfGNlhLYhkB4f05RCMLJqlF9
lF/XR468GHl/DMjtwwrWY1DvTWZzHdxFk/Vz5AMTFJfImYM5CMiuyl6VdkLTSOysHz6Y8xH9EVdS
HB40rhZJrckHjalNpYI+Y4Vw3CiYgKcmX9s9XGy7oA2ljqTEUgqRlqKMsmDdIQbNpN76ILpn+k6i
Ycw2s9efdLor30166mRPZ71tGFg/KtTzwzaNcs7Y7J4umaO6in2LuIK6Cz9QMdQnINce9dKwfMQp
1z5InjGEWR7EAP9iwDa8zvWknL9MhPmV/7rbtXQlJ9OBdL3MfqjoJ3W2Gy2Z/iZjiS2uDIHfEixt
lS7s997T9AccwqkgZfHxuLrkpf3wwCLj4eBFOD3+uOSWS2iN2IoHXk1oBhp1phL0dxlyn50MUmx7
vnt86t/nyWOLmgxda/RUEA/u3DON/dgPvKSZzQW9a4QYP3rmJ2x2iJhhqeASU0ajTgrVF3wl44Ti
pBHP2O1fHQ8+hYgZ9kX5+hkAREyy8uwQ5wWcEEH7cOG6p7ZV9/v6jg6GUCZBwPYnE61hlVvQakLo
usxKBuKx74itFPIeb8HYy4i3L+L5sKL1SYUjx6WF/QHTRU8zrkXcgDodoEp+F56HqCAwrM27G/hg
FN4XxqysZISMdM4KEsfLrJshcuQ7ryVY0q7TPyWfC8/ur6LsJtluFiRz3d9JRHHjqQKEI0xVZLn+
W25CSV0JsOwE1kidW5yBsXdFAwTaEkFolNI0Z5ODVDKUfK+XylhMFkj2W2iuExGkQOf5+eRAG7gG
RrkkU5OZg/5d0CIKMAS3fAw3hrXJhvgFxZEFaKM5C4tfnruKjXVprc0TGdkasDN8jgB6ays6jaxH
XuX05selRLvkeCSmB13lQ7jCa0hmtVxxXliZpPVGvWQtsPYDw0wlF4/07ES/0Lr4H6ZnT6nFMCkp
8waiJO1xBLHKCjc6yxo125bTV0pcBID2+SEPvP3QgSwhLKDwJO7zgTj0TNhO5SkZRIF8CBnZRMWj
/isg6HIIjtlC6M7MQ632zj4RCIrpXEkWRxQEoKJZSKQ6lvYU9goXavEK9+u1neN6Itb4rAypipt/
xyKaWabWVaFvqZp3uB54oFDT5Lnfg3ncMEDfmm0zHeTnZY5fJghh4cOS3LNa7r7IKyUX4+OoWDO4
ShE1mpnHn13Vc6gOZHGd966L7K6oNcKAZ21pq1hRMFJTU5bU+7DQg6CQ0zVATXX3l6PGOPb5bvdw
E+D6iBP/cxPhIu8z9NYFAJKFFMxzXPi9xBf7r5FUBbgwGosKIniev9aelWGJgVmnGFjPlsPF5gDH
nZiOZPgxndXimNH7qrLurJ/OLLDzUIi34R/RdQ8ut1crD77GVtYSsTswyDZfIdiO9TFO722Pg4FY
4M3VhIHMuCWq0wAh1LgUzjaQpLcOUaeUfmNf2Q2kal5RVxE0fLy8YBxn9HDSv6tYi8y/go2GkJW/
wOASIZ8IuY8gIuRvWsWB7D0l0UH+3IQhxTZjbZmZuyK8AIAyD4X2Y7+N7HXigbiMcmJebDbOLHPn
NS+LJ98Y5isAkNwchI162LfpObHpbbf73XYSW3wTSkqlPeqF3VYgI/FdH4hKi3uy4yZjQG6tw54S
DYVhg6vSZ9SkkD7fvX0mH+YYTDqD9WiiBjbYiF47uIkorRjwt0GdRxZkw72y9n3joYzuG99l4I4R
D4/HovBSJPsnV47W+j8MvGevrVRbKOeAXIu3Q0ujT5baA3bKniuV/mPgBpYsq+bxGljalugtaS/r
IkdWS5TtDZwGumWVu0r04WWg2ENEjFQthY4axjh5t2m3S9Pxkxlh0a0dRSjIwoeDVe4MQNYSURzO
CKm1dfrYidqnwPw+yBW4oKglEJt+Dc7WC4GFKI643EKnlMpe48FKNMNsU1r4VmmGdyWIFnBcVtSU
r3lpcTugCPuKNM9YYfbZ60p+uJLsylvY2bj8fQfwAhESsk8eQAKpJBGM8WBZc/bRIXmq8iTw2l6W
F9FzjYDgXxt4d5oYe1qG6QrqSqeutF7tGVSdpfEh2M1QGzd3m+7y5opAf9L37/lm5f+t5TMBH/4W
T03U6bX/pSUVChRW89YG/CgQ29yfhKjRmshppF5012M13mU4raYl/Fj0jUqFcRzckv7Xh6n0p6aO
uhi2RgeHVdZP3UUxQNV47v5EfJVuZVtbNaBSFcZ+SXNXUkp00yWUrmabp87ivSspuPzCv5IZWU77
dlz3/2bCc1U5KIAk2XX6SJt2GETas4f1U7r3Cw6ob04BQHIWhP9JW42zmd/NOGBN/ZdGoMeAWBBh
Lj6eTnyH1eHQ3vsV8u8u6dHuRM1PnJAfC0rio3p1hY64uLQFslkm8D5+Y1snYJJcSUNoprQoTvx2
NGBKSe1Ab4nO9Y9LSXMC/UupSuA0Nbi8SoPMDdiD3+vx0OhWrdz+guJHi76xrSQ6IvOprIPuQYDw
N2HMjOAwKywkYbCixbAZ8BrSuB63/BTBRE5wHrhNyH5XTxPDrIx1JA0b+0VkG4I5zCSgu2Zj5o5+
8TXk2Iz7HBRRX8DGTs/P+O8QZ4vCzqe8fZ8YW/AQ6J6mrATAzXgZHs+6+pGhClo3Syb3yZ4YFqAn
yAAWXtPY3PRsjqVWNpAo/t3cZJ+crugAu/WqrviyBOQkY4j5cKNznGN9wKTts89C37rNan/kIRCE
fEsoBuP1NCu9HvfMM+qmh0c+lmUUelI67hgtE7ymnoPy7wsnd/UYfnh0AcUWHxLGn+gT68z7qJ8O
tsogQJImZhEbgB/cZZisJHwMuTN2jtd/lDCvx3i+4wKL69TpmxcScFSYJyslUkliS2JoWFXN4bVo
muEZebQmeKc1Y1eVH8zF5f6ta0xuHTdiFca4iPCqxTu0Y5YemsyHYKf+UaGpDv6y1SChZVq1KE0T
GOjC3LDC7WQ1QWmuaGC36ASjrI39vCzpiWRgEosUhO4oUb1VvIiS4jQbU8949N1oksFv1+wolzbc
ekPoez9R4/oaz0N8CiQMH4gYCEDvlWNuvnSbIuZ1w/RtdZu5TelYNPfPk5d3+HSaS5MnuX5xA4Kt
85pkwNIB5F1BAxqbjz70hepPTjmBMOxaODcZRG17HAMULKpkDSUZg51niNFR36CAsCjORYxfyoxj
QQhCwSts1lBjhiAIJqJwRbEKU/Xlm1mHAyVj8bS8LXu7hbqpTGXgNIjnKRkgnjk9M6dB47TJWrER
oWaAldiNYWZfLWEK3Ex2yuv6MCwUFdXjCB5eK10xa0wMIGFGFZwjbLMSXcxClMU6Iow70oaMDm59
1NP7RP+QiSgv2NYYMmDzlaSQqUHDMn9CSMRaRJyr8aKKxYYhDC34vfjdLJX7vbIlLTEMpYA6n6SV
ai/gyoZucW57/JbN9i4zxVkVcogR0V6RuIyuQppLShrtv3+jz/CcecDOUdWXVYeajafuvy6TE+wz
zc0n+ischYU5UUUldYu+eDLpQ23FpwtKObT4teE9J3cfhZBgsmQqVinTlBnYX3em+izF4f3dn1OT
gYuoXQ8YjkO0gtuOl8RwuH3IU/mjJzfWHHrX8RCm0ot969PoqHZ9U7HpDPLYBkOrCSLaw0HNDGTF
npCMAPSbzESjyCTx3X4im9G1JVQ+5YzW0Cn3VD6BGGdz19UEOq/7lY0YuAppUfSeBc3NAto4HBn+
gKLWU2pNXBsn+uznT5r5/QaiU+gmp/m4AXhoHZkfSQpsJZKY6eyTt8ZeOH/ORrW/q14kyqTc0DCH
Drf8fNklXnjm1Q4Uzzk9LQLX+oKqqk55SAJ1LGPoqrzzG9s2tRa/CHrVlSsVHXS1og14hCQEYJs2
amsK6uVfMtVfSlU2LRgratXznQ2CBfmlNRWHXbcowlagIWgyR0PxwiBKOQq5pts8J5fuZPJNrYU2
sW/BSv4hgV+o1wYzGOo62b2bYOwQarWl45FoEnfv4hXxKKDnHQu1Sjyov3BPBK/qchikEWHO4zU5
+WiqlyrXFNuWGDMn/Dn58Q0ER0gytHUwkj0Ex8QOGVdQRwX06o89+Zlf5KoOoK1ZBFiPeQ676N6h
UcVIuQBFQL0pKVYD/4zg0yLTVlbj6fvRtvCiNo+tMJXMmTt2FPCHwOPZDhc9RlZEajAGF08F2/m2
1eYybMDZVfNyx47mmFXqh0ELqk5yZi40qdoDBx6/iOQ8X7SwyguYWK/ekPCg4ELt1cVtf+v1tQAd
i7wLRUE7i7m39XLk+bLLo9uCUMJiNFH36GakidSmBD1TdZqGGegpEgK6q6Nm7p75n1OBlfl5xErC
2+LlW+QspH5Yrh/Lar6YSKte9a7hLRK0kKNEOOy5ObtKYrjBJzAo0kB6CviO6ToYCqLkGKYYNrHs
vGwTrd890S7RMoDqEDa7pY4nIP+4nBmXPhUzb1/bJYnGuLi0Q3mdqyt7j084KtVRh3whWZfGzxEG
fTt7UotrgqgIj1X5LF0vmyVuNbvwp9VTtyPP8sXrVyFeBa++4Un2T3E37INqonMESQgN3XI3XnzB
+idrchr8E4317n+AszZgHiiz14DTxxyYaKaXMLnD65lrOCQBsmFySVUQbuQn4CiTSUWhe/nIMvSG
qrMeTzehEqc+EJqAJz3LsR1w+CSMHezCQQRD3sxai236L4r6OawmLt3jCGr6XaRoT/FWeReAY5UY
4VtZRqe45KJ7pKgpfh+CEcX/37F/UVS/6kwIKiLL+B0PY5MvI9ySIqJWu6zf04/3gA5nHtLniH//
oTFVxZwT/ZHzeKFEqE8XbMdH70RILidIZ0r+XnJnyeQxq7SOC+VGsDwbsMbfzFQ0VYjdIj9s+LmG
ohovu49btNet2QRAY+GgLaYIc/yxrB3vIp2Lz9gQPk6nbPt1QLhOZ9fsFZhGd407yomao7uENCW/
Toi5ktBQHnOTN+Q1v2fX+uLSK2kyl7MS2xkmwJ9R06iydbZZzosptZXtma3/XmqprVYCfKlaLjbt
Rt7dvglp70YndgZt6ERNT6yGh1UVfvXPg83hxQQlK2YSY6EptrgajfAv90wD3+XiffdzAGkrX59a
9dq7sk6cC5a+5PbxVxyoOuFsUzY6+QQkbURwZ6tUqmGzAeaTTFm3we36rVVZpP7FsmdjfQ5la712
yuFmX7j2HE0d30RmWDJGegPklYIlTDj6d24HmwQKBqAN+0VG4uL5TRGZ+XA4JquXfeUQ4haXyhAr
5eLfITEiyRCNiKdtCPoGLjEgF+TwRXvoJ7mfsniHYYPfG0cW1InlzmjSrXPxiraFTQX9Ns7s9o7a
QvginkXtoqskSByjWj0SAKJYhSbC6YrMKsILPTU5EY0unGiNffEQR1Ew+K3SiJXzDlts48RYCUzE
Lw1YgLbAiIFfuWKq2ptGRycU8uCd5lBTWjSFzubc+Brc5GZm5QX6LJfYnHASH95B1XCldakh8t9a
bfsHFxerwM6Cz95+ybfXcgMqjUKNcs4WysYFPOZtHXXmfBEMjTBOo3KcffpVD2Aiw3ko+eAn2PJo
ZdMiMiztV1wS3MaiD8zeBbvPZcLTu+Q1l6oUeUhsIqvi0JsObGKOCat5XjcrzoeIXD/X9AzQagq1
Xg8CT/uupLO1IWtQg5u9WyjRqFUQb2WqY/8PZBjV4H2ZGdVf63cDu2WRoK8oF49YjBOpROgW6sWN
nHzNPNbV9EnpiV/KjylJwNd2u0yMSxsMXMtQWF2YF7C/dt25vYiz2I7Wre0qkP3QFXuCUFeiuP+F
UMfmkY5d0AGVRJBrfZqzKsLv/9C44VAvpBh4SyXiVWscuppv0Ig6wYLoCrAMeFB/5cJC4hvL0vpu
JxvBmxqwAFsbeX4keF98sqLb4L2RyrBXmgQ00pUIZdHjZ96WS8ysioGjrbJaIZZtClPu5qf3GaGv
ISxcUPTsNQq0wqOIVauWZildZw0S1/AB0SUkzPEojIe2HqySgNVRoq8wAjzTokMisSvXL98JaJf9
YQLHivQwKlOWsGxExoNvRjFnDf9vl6kogW+qhyjz737DGEn96ayzGplCui7bNXQbf9DiQvTw0z0v
FVk6JzBcNTakk76zux8GgGDLVxAEXHuYIsQJw6Bay0BiCGV6Kjr/UkFaB5lJX8RoXyXoJBe4v0Mp
CqO0UcXemtAq2Eg0tX9dtJ9lyjkznpKC4lDyAODDVP0TqkOQcXgZHURQhONYM9FcCSM3p4SnB2Rn
5HzS+SJszUr/w5oY9u2y1cDHwlYpc0M4T9qvexb6bB/C03DyKYmI/41ADz+b1IlIRR5la/IaO2uI
Hr9lLsrJfgGNI904mlcouhYoigFzRvaJ2pZlSOzu1TNurFIB6+McNgJ036OhND4LAxwsNDBPSK5L
41zUlvc8oHP+Usa1bB/LKDgF/BwXeeVbJPjDf+q+TSvU2QBNitKJw2YC29xSPYdz8V5TM34bDTyZ
LmE1en/J4KFngDt6MSlgigPzpeRhv4y839sZTf+Ud92qFEfk5Xa1wc3S8BxkaBzQTnf1hFbbPqi6
ZL1gHL+CElulwfdGOkcANWUMoNpSPuLs7J1P3AaxV/77Tolcxney0DrRk4/ps99WYt+JYPS8AluZ
HAFJ7E0VE4HHxF36X/kKWlsCccTvwuUTaFmr+AW56zx9nSAgCXGMoyFaorvrgH875Pckc7Cr+lSM
u5sRGLqflKS9IKcqbzd9NgahKVXjfYkJXoKhu3e/xbYwllyPErIF720bIrJh8i/P6FmSogRuwvSY
bnXBLsDDR2eGFfWelAps//cGosJnRSrVsbaljEq2SQWzfwslACPDQYe/8rVijbKLIqMaCyt/Z2XQ
Er9QYEJtZ5FsvUbUI0CoXJGmTNqOS8/YISDldWdR7i18+e1A+3GaTEjjxm4Cmpuf0+Z/FO4+XOdc
FAkx7SGleYeaIP5xNUBlltbd5TJLruP+9MzFXx9W+nqswMtzb+UnW67RBEQvHzOrJ6nmgrmeN42a
dwPKnDxC/Xg7eU0Nb+dFvoWU2/B+CB94KgC0OtQvp96YUY/cynMyNWWG9QlzYBsGZwq0A3RT3aj3
pg59/UuLmCsK8jogb2iI63UXli6FYp8b3u8N5UYSrvPyehb1RTgujFqTMkca0msZuOCoVmUgC4NV
989QQCwlFADhUyg72V6hvG6Nh2y9P+NP8GjtxLJe695FG38g0LydY6kgGzxkNtWhVVJswWQ9DN0S
+zM/SwyWT/JIuuCVIz5vu1n3qYUE6LMmEEAkHmEmWCSnATLktoQwwatZGlmn1ZSDx1N7LlWTicPT
PC49j5v0Ss2x2cnCMTVJ5n4zHs2AqIjx+JdF7fVrZnsmNc4lTWkaua8jJF7foc3azM+9klbxa5r8
KHdi1G/cWTcmD3NNFoZB52bvWxmYN+jM4WgJwBA7qq7Otlqf2+j/jZql176Ynqa/W/9ltCXfkPNC
dteJy6aTR+9VSBiRZMptSDVrUKQ8EiUVYfYfNJE6KUK1aqTd0w7jhZk5jJBlogtlayiDtSdrdv6t
c9v/ds6CY0JZX71YpvjNZTpgYKLRzXVD5qAEeR/ZDQL4LtuUSjDG3L/v+BGS1RvTQR0/D0kLGpb6
+4jo3dm1u9HFqbdIq82iHp7ThwRdjeI3PubFcW+OBLMUp9ki2rD70Ux1Bh+91xa9G2V7iY/IXJi6
05L1jCq4BmeBdwFso6Wvow9rM7T/5+Moq5VgrO+NkOm6+pnew4/HbwL2Kaa8Yrpye4QHL9Ed6GQD
BMrX+1Oko5uI3HUgrw7wbeiTz+IfDniVXkieMcjo0LjPH5R4DU2zsIDGSrDxpizuwgwNR6udkyiA
zKjeVuwz0PsksHskJN272kt0XdQ2k3Hj7PmkAjySRTpHm7WDYSpPrEyR42FI1pIpXyk/VXJLb+m3
W63yl0pZ3BVDsDmRbv+1REuFcgxUowdBiVXHD8v/0vGOyP59BLUZrbWU/AloPKzf9sDsD0b2o2VH
eX3gBlVo+LPW/vXUfgjK+BgT6JmJ1f8wtTY088oIsV0G1t+JXLk0ngrzodZfLgAPeTlFimuBazBr
oa0zG9v8rOAt/6qs8RrXjfsUVVQXX7TnbinxParFcngLRoQO9+tqeKORQC0zID8QIPrUTQ+vXDSz
e3DFs4noYGjpLikQJA99dWvc/Ee2538BLjWpxuPtQ5TNAo2shYQCQUMGH3bno6j0LubhkxGJNqQZ
crOV13snTfOHoDg2vcFuvqXkCVm9ZgtNNe/b7tg5Ga5pCmgoKEDQ2LXij+UKuaTsRdCyh/rwVD29
07TJdTULw0DPFWwMHW5MQHqUxgXpxOeHWDfg3VLlKRXz/z6pzKRoqyHcfJYUDPCRyZuQiGeSfcr+
pevKEMa9YBOnaPfGqsrrVSfA8Hd2/zqQR0ze/nIiDIsc+VV/dATXyIXLCylvNlRjhWxOCQN4qthh
uOjQgxxxxobD+Dm+OtwHnoNqrvAqg0ISp7dCW1gnYeN7Ak3q1WeQpkm2zWTqN700azUnb1SEEG7c
RYpFgoPtG7e62qiOUB65AfPewpgVonwO5FapOTBclErFk9Oe6dQlbpAsCYTOxTD8DnRKOz7EC7VP
Gaw91EwB6N9k2gNMgcCweiGR4IqiE0QALIHTrrMftqkXNyNbAlX/UIbynB9CncbZRc4ood2/iPAs
GbtGvp5w4nZQzcUsgae0fhbaURfzcYj8l5jrOCJ0vmROoAxPkdtE3lP5LVYAQCcXxVs3u5AJCKTd
hNpVSwb9/xN+NVb8UKgpe41+onv3xmx3egvrPfc1Nmq22w1h57IP8kaEy3vGTVYiYnGBAAOtdX5b
Iu+uxHQ0Iq6SdX1Iak9sIOIPERo/hAfmdlDa0cmI5uSrigSdwStfvDJ1z/IgFE78UcLcjNxSBHiV
hIfBdsmGDGQOMXagwiGz1PKF99yuqjRU8xe9bkv1fGgWnUY4MLf67mOa8XpdA3BSQvL4UgkdiYzs
Dt52mDU97IqaickbDeF7vWKZIpjNKX3m4JoU41q2KPI3sCVJI6fFAmGfRkuflBI1Rq00jmNyOysi
MVfDZJPckDVa3m4AHE99yUf1QI/Bw9B97Lg8ibDl4YG4z8UcniLyV+IFbviXGm+QiPnZBWvnc1k+
0ANhpHOdcJ9h4wwfz4L7PjvRmJbQqdQStlfjp/TeGklQpTaiNydJoz1mLo3VGZl8VzAYpnBhgG1B
bHqsJBtxugt4pbMd4KJSgGWk74uUFFv0ZFl4YSSuFoaBwIrqE6G/TG5SrYeIoYfNRrReNpr+xINS
bomMti6bXcvspBHCS/BtHob6SPh6EgZJFoSMaKD4W+/t9SeKXp2CQzzdWe6k+CRMG0O6tD8RAgSu
3gcKtD9PrD+vay/aRJIf1h8l1BtHSunRyzo2SWd+yuCH2HeenIKL7qqzVliAe2Urw9oaDX91sWVU
jpUFqvLOyUVD4P7bKVLW4Tqq11tumEe0sP08vvAoNK+VjqB3GC96tdQKRJbNkgfhDwDpTtTGRZe2
ZoZJE+hJOzAYNvPItD4BH596yd2wxPOF6jtrY0tsFhnWJ5MRuxHCXVEiHDM5IvEvuvn4lfh9U2yT
dPKXGwpOQAeDGwD0yx/Stwln7tcC8BjpzKpvXqDPDBWNMyOWSnMP8b8UEY88tdaQfLRGCqQf2Poj
YvUiNvhZhIFsH41fZ4409LLxDcOc32YM+IsVWzf0kdREjdR/V/o3KM+SclKvpbhBtkFXjqpyIW6z
vZve5vaYL8WAAxjFRguHOV02LQOOZywHBommF65dBh76K3ag12Mkv6qQjRf0g/jWkp/9WZyJG90j
SFM/ZjDOAnFHuW70YiuK9mprSpbVQMZHczU2CDlviyj4+f2C4RSnokx+vZwYAS13z4j1LXEYDjmm
X1BhmgZyYw9hF7V1pxWO4eUKFI800t0vvCLeoRqytDh00cD2kVygFHiu++7SxV9iWRSSl4663CWj
A1lpTTQcleygsvqK/npXEstzEC9R1YJor/c3xjHer6zSxL3eUPsHPY0sVFk9XTglpU8pOokpUoAQ
iptCCXLkcpsWu8V61eExhYBDXYeQPdYIL7wY32vC7ddHsBSUclevZWFONICDuFitD+Dghc5Kpp4R
A80YNdtl937LRnk1g8a0t9NQ7XMne7mm7oT2r/D4pq0RWAz2Is62sejKmK20gIZINbpmX2Fo3v7P
cfC/+z++ZTfwhKDy2c9TJjB91KgHdhxia/j1IzQsBimIDOzQXSv62Y3q1n0idOPS/TD1UQb0dExw
feqCOLwgjAnuQP8iEP0hqD3iixAEpzcAHlcDRqYDkXiIizN0zmQ2ieOCr0NLikkE50QP1zuODPWH
+UiVcaU8FQ3A+qsMlgDjBukPdPCxYeeK1AyNobKG4cS+a6DHHKnef25UbTrvZZVrAHsImwnOCJF2
L20jiajYidMa9ffyBnWb/yN+v7YzczpkG9/76CQXHoWhzsQp/3g6/F+HpKIavu7tDjm31PKjRPim
qxJdEQmH/mg/UZ3BGJqfoZfR1dWzSSS4IXMm8DCpKFSnItEP1uNO2Rnw2Ld/zuOe3RfNrQpD963T
NGFvfTeFRIyLhJ5z9Pt/jTskTsHSVIhJvZYMRZ50eFgsLoYq5EbDO+PicOcDqMCCS54hcqXqUidi
+Im/chmvkYwc03wcjwlHATej7Vo6zAUTXQ05cmScHEdtvWqFXorEwUOqZBzdaUl2vu4AUqdiJ3lF
dACFXHjxj0mUe+YzPRoQhu4SZt5prjox+I0Sa+uM/D+/15zak281DnC89zCUsIxMjd2ntlPc7m0d
g3kCY9XQ1A+vLZD4Xeoewstr5I0hzu5/Od/qilXQYRNSNuiZ9QzY5+CugTiSykJ9xAUGT5yVVQRr
m77AfdBEli1lIVSnezuYGi1Pf0MrTnchH4568E8r2wSNfsOSxzaE5UjZAvqf7cHmCktKFsW62ink
4EkSYXj4K1i+iWDICa2Wh4YG1WQFfcbnSxoV5q8iynbHTwwHXqHVgKx40loe9CwQBJGPoRG3I6JR
uF4x3adkqVs3rgIX9b2zaSVZvcsgutv/xDguFFLPOcxTO/MJVOMEXPp79V7KsMzttYi7xQx2LEYu
7zqoZAptlnEI/+jVOZWDGWS0rlWvbso8u/9liD8MhFc3IBEhwx9BfvmEg8O/Kutas+QSxE1bZ58U
d6CV0CPpo1Ym+KKk8ROv0iqmHuupfJgNVjbx2ofcuhufpuwCuULRiAj1bzMrZ4uWCl6Ov4LW3MDk
z0DfLKkThbJC3d2974sw0tN5Pr0lun1zA3y59twm2XqZFlD6aW6qRUyS+a+XSn+WVOtqAWxHBdZ4
/IFmsF+IU7PA6eH/rUfK1vwqzZZpqx8QQ+GsjoXx5KB/VyFMI30Tk741eoTWYGUimUxkyJJR85/6
exj0jwnKEiPEzw/aUhg4a3Ys4dKz4CJdkMFFI8qvJZRjWZ/kzAM+hKA0IFxcY2sWkNT7wVyi11FQ
PhtXM3s44iN2gK6HScGdjKasXH1V+fshKG/Asc4hA/TBKseZGt9fBCrljX7eynL+yB+q0bOHQHKa
n/enDCm0I5GoOisN/z+sxyDvPjvmRTGjGwRcPYIN66Y9FAJMgyRFVwXSb3C4P3s2m3rb7Fk3TYUN
IgmEDm8IEgBbGTJClXJMkIaiRZfEoml4m7ys13ZqnEW+rPXYkX3Z64VzNFHFSS+mS/q2LuzYWuTn
6D/XTcmewm6TV0hmF2/rK/7T3uJ1gl+cikKC7VEFzAwJAvIQEcnEWxyaVgyd/SOnlgSEDdOxHsyf
XnfPc6/70Zx239mHlcYhrcNUX0Sq6UeLTy9xn8uXkFO1MdlB5ngwe6FL2bzWQDZ50tTB5DmmFL7I
9GwfNUoVFeprMdN7HK3UoOuTWVp+oxvfuNkyo8kJqRUg9ECBTtzzeSNFiN7mMmp+9mVz+/2CCX4N
fmHtTvhUPHlAJ/Kg5IqGAoAtqraHbNzYB4QgNKI8wgSxTwghQ1cBULupsmsoPECoJKiwLtgFIYl1
w0eNxdtL5LG7JylwzVteoOYWxxHDEVlEzDnTOeochl1ZfeqJ3CLQgolJig37NJe/Hfl4drWjNtU7
r0cEPk+lCKKejroA/PQm8fzVLEt+0vW3r49KlC730VLJo8KU+9Dsq897D2dIPnO7U+T+ifxDAx5Q
hHyAjnU9c7Bh6Li0jtIcGiH7t618gtKC20I1gLTsgba59+8HaZw15in7VvBAmG8LZqYPcXhkWBba
uiEknmI42vMTHqWmB/eW5llnxlhM4CvBXnCVJ2gc9VACXUFS367vcWswZWexuVQPbuYIkeUoDUA7
z89LyqcLEca0v2t42HMg1jKFa/KgZmkFNVDzDU+QE9ypRH30Bf0yHeXYKWGA/o58TpQh6JAPjhPP
foBe0BmyOYeSeFXaMiU7+eTXG7LI/hnNOrhcJvEbKTFQSYATIBVrRkb9ewniyxOHgXsHAZBTM0uE
omSgzvUnEOvugZ8PEO35tnIUpLKfg9Qzi41kgt/stlcEv72BAL5pn/NCoOtNmJXjco4mmyJ9tPuJ
wYWWQzJm9v2xVaaVD6cu2M70V2yzOepb1Wqjr4w+K0AJDsYtUZl69MG6FJyXOcXzR2npbdiazd1c
FB9QFaMUZv8xjuioGgE5mMtOL/L9Pnl60JCwHT/hT9j4G59RwwsUlkwTM2BCMlCEdHISzz3PYlWc
D8119oqT430Nxc/QQlFue0RXJceLhlwCWmKOCptw3vXX+Wux2Zfh3Hq26DYPv+L7UFA4LzCxi6VH
6Sagl7G8qw2URi2qKifMum6m/lUN47M16GxmOUztKeEN+c65UNmemGqAMQ+kyMwX3v0igKivN/aG
8cEvOgXkvmD0AXoIuXwILQjfR9f1cFyp0HcxIwsRKS4Ti9U69dytTvKy6whg8WTlRoiIs1WyhTgX
m1Se4ztEzYRiJF6Aylhk7f/gp9fWIuZVRwx5k0Po/KNctqqrrLvK/5XTRXC6gm/3ek31bXVtHD/8
3jgRfL9cT0/VPJzJXBGsnv5Gh6cTgsbeMgnODMULFsoFpnbqxVzKf7IjoHT0cvSb+amVBLzP+FHr
NR8qodSnp2RVuXjcAl0IQvipGvJeUDWvpsgVyxuvEH55MnqoGbryh0pduAcmIAgV4E4l79k6N1V6
ceU6/M0k1oFIfiO8Sk+nGkmSvZwE7KMu2TKBR8d7zTKF7RQ3xna6oHY/fRMndxU9HQ67K2p1Xdzr
/mD8xpeWqqV0hLcMW2nkXDfSUi5ISWUdVTJ9oLlV14JvX2dCCoM97u3bmzqNvVcjjDu3c0yNG4aK
aKsyohdNkpyEYfV4f5CHrZ0K3K8skFkVnhk9efSZbb7UTwgJJGigIc2JYISgV8PPeeE/XbNmhNu3
5VDlIK0IXDF9TcSVeSjSsammDXt2HLGub444+dlBF7j3m2RQQmQ3q4jsQr84KFvFEuyfT20n6hO2
3pWbey+yWhxEtfVr0IUwhsDgWpDwKnAy/ebyvR8Pr2AJ1A+hAGDshPVGMi3P7q91rEueCWubcdz7
IOcVfVQa1zVZ1GwKE2+Cr+zwLq9rvwHiRV/1aN5HsAbdEuUJZn5P1xMLKRlpXTz5ay2xEL8CO/PJ
prlBoj8cdu6b37MUldtAgWW1pqFCciHmKsE2VuUH5X0cgKrhs0lmsOLxyF83bUv+53P0H3CAH17A
rUVAU/7l9G6SeQbOjMfJ6Kj29L+IoZkaaa8YLifCCTtavEh+WiNTznDyjQJ+dRPrc9vzvjUNrs6V
iMGeUON9Jqi0v4Dq+8uYq7JdD9ekjMCg++jj3n9YDEOF9nKl5yjql552sD1iFvW7nyoeDIV08Ig6
xXhMaJzb7uUjKxrlD9/4qyzG522HSM+BGqvVCfQaXX2fWRDtntzUgfk74xYwk+XHpUlXJUfx4xJD
p07y2BexMzbwUwtG1b86bRDYu3qtqKMJ9HsipVuORHmREQU2qL0TkiM+UxzSRV/t3XJ6Ag0B/+OK
qlKBEuTi5YSNeV3UPzwckFirop8Z+x+fAseI8DDl7rQv/8SMpx/Xqv+Gqgn9iykYlpR6NAZOPzmL
mzshiiq/alvBoSQ8bDkoE8BWDix56mQsZbK7eqOzlaH4JIRqfLwDqN+wJvamKOarjqjvMrqSdCBR
g4BqWBIFED4Kr3QIoP18ovNaRrfo4VWic/iSudfeiVD9duh1BlvAuMHh5hqSKkdxv/90pTclLLTE
NJgRaR9JTT824NlibbXfTlDP8dqK6Tj674Xf5vmSfjcKPYAuR24iQ+XI3BcT4xX+fz0sjz9iHcqS
PyLTw64i+9J/qIkjr9zBFMIGA9q9akSwBo2KJMGFB0AQ7X1eQAQ72DMR6rJDzvaH4vo/LxEjrEEq
6IotedTsg/AGnmw0EmnyFcvvVNAaMRb/MueTI1vNF4069NoEuAYu4DALLBfibJ0LdGktiB2o1BXc
B4hzgcSsqoFQSimBSMVzZhbd2MTz/ZA4it2Rx/Cdg9fvOH++5XJ6pyRl85giwTXwUaEWgb/oCTK1
jziA6bK2UTgb+C4InTlzJ7jNwyi9RdfcxOSs4gTFq+ZzvsDLE4Px8Iz92QlrJUTq1Gplo25gDq4i
OK612XDIYTRyXeyDR+iJZYdamLp93Xbtat4KWuuSFoOdC4QRaZic4r71UoRIg91BHxeSECcdG/cF
BhN0E0SgVavVcUzuvgWl5LNMKy4GPmyBWtzu+CsooXiGCZd68vSh5MMqQpwnXbdqfMVRme+5Z6ED
15OjpkIADjVTtU0RCeW3qRxG0Nr6JainXPv6to/HRwoK7pHUlo7UdrEwMSPsakjpRq/V9h39QrAG
tRRra/WcvqFDRUVjnDe+I7levTcZeH2EJml1unAT1/ZrUgc79b4Vmp9Z1N61eo0/kNz7qIjHykgq
gxsyD6F5SQWLTqgv+juffgaaiaVFz90p6O6B30drtOUwT/KvdOb9gTXzMCyMGHFWJLtzTJzKgOJq
WylJg9LnKBKSSj7o1wrAPAeCE05hvSRSGWoDGy9yUC3ck8MGYj2a4ZXWSpSD8reKLn/FHwkQwp6M
OMHenkkJ9KD0z0dCBE0mgRdQ2cCWMWSM+22bO+AhjWgNbwECtVVh8c3zEo0UGdISo80DJGerOXlE
G5jc2A+d6fRDYdMZxVlUWq0ivnORHxiU3zsK+I78LXH43hJiF/xh5dAPFYlUfTTz30cXjdpyrSzs
AUnb9Hw5LdghL76thZY4ASC6bJxoBmK1B8BPtDJr76Vts2PpREseTWC2NQhUP6VCmZJqqKffsh2N
B/xcnBHRpiO/C4usFbl4KbCzXEbLCx8NIahXhOgBKIItZBWTj+eZbYnrklgtH3vJPPvakDl5++td
fwQPP5b30B2IaipwauZ2dpbXXopo7qtMkjfuByfn3qV2hXfwGRdNkIknZZXgm08ZGQaEhxF7JCT4
iKngLYrkCALStsjxxcWPMYyg0jxY+ITmRBzOoxlHr8aySe0hMibzXSUdhccBHLgRwDhJ51JhaB4z
Mpn41JXiwQoM8PHV43XDodvUK8m0iHTKbirIbjm3xLwCJbKsWSn4Tth2NkNzpKceF94QKTcKxqcq
RYSGe8m0TcsUglkArl+Rw/EB0Qb5qLjMMMT+ZPRlbFI7qOu0AE4iqfB4LIeZSMbZcinsBpUtld+9
P/nS1UC5MPgPL63JVE6p7VfydsGpW0wUZwMv9IjctoSKBmRAvAoMm7LpF3r6oSQFgVJh2p9aBc4s
7wCxI5R5uPFDrn9ValrpHm0wksDMGSV34cQVrz+lxfZRrPr98jocm9g5VCxePLd8+r/ssG7b8Arb
pMc9oSpNvQkGUwomwcv4qQQRziiX1ibiGdoHy7q83MxLUwgfDAQKFyjsR7RBKE445y/ehMIB/ClK
jYSya7DCSC4iNv3SOPXu5aMK8lhYj9GEAh+oFynpZ41VxUyEpHuhZhN5kMyMyMKukkk5pw71bLzN
Dckxg8trjqZPM9f9psgS2Pnrz4o4G0FaS6cPDcLDwINYKGo45SP0xMfH/BnSQ+c3N1PviJv14/8Y
W4uwNUevDceobObE2MjmScVikF5TfW4OHMWqj3WujByxovvH0+abVVx3XzUZbgAgZ5fGakDG0+0W
JBymArOmSbKB0KtewjWD755qvVK3bAmXuZM/ySc7G0FG4dvBbeWXiH/Mwk+aILbB6Sh0N2OKBH9h
zGU20CaPvZY6iCyJIyavX723UTmjzFjv/Boviuh7ajxCUMGrNmN+wvSVm7IwM0VY/NA7mn44crSm
PhWvJECLS5V2Sg15KslwSqx1P80wDaLkx17Gg30JlB8ZXefeAHZ75ZEkbKKT/awkpd7C0TKQ6jeM
ISWEJPiAHWZL3p3r0pFPFpE2yenpfqkuJJHdsYfowYpjnSZF5w0E08IvWY0EaG11DqPPO1YtIcnp
Rb23tnL4YD34PLdZAhS/tCEyUCfI9z9h24+TT/gQG+Prh7PuFfBbm4XLYD1sRnEHbueQaePn5oo0
Ih5e6+MH11B014X6XP5IYE0jM819UCQfgQBDA4pj/g2fkv4eXfjXI4ovZlaDl7XmdQeULyHdA3F8
UCfzUXBUps31UKlRtejrLBcsgrsgEcj6Fo2lwMsNTwgdcchlG1SKbv74FTAHALzUzUOe+Z2lkINX
ud37tFawbBH/PH5GSBOdCDKpU4qXmEv38PCVpEvFwL+BrTepfezgEQWj7fUad/uBBoevqk9hrC4Q
kxgLnSBeyITniMOOOIYNAPznWuv6MDl5rluadOoEKhuibvYa3iyjrBWf5cizFY5eFoLH/6Bqdegx
W4vZErtkmyN6lcbS/8IkluUIIo2w72LaNBiBN+xNkFvMiCHbPWnru5xe805ISbiTfVzvz1wpYKRC
IRLXtgqipcfVOWBZYkUO0gHlPsYU9fnziKiAL52EUZ9PxH2VvzPpU0+mLJGURWnbV242FHZGkiKp
BOLx61XBbHQ+tGPGPYyl46xYUYNKIf6dYFowlKRQ00Sq4ZQGS99gGcP6ozV3N6PrgSMSs8OspWSd
YHfPNvVFzhF8Rej2kZWDs3Kj0DbRjJbVW2AjhFkXmx5h+pKxTqgqcLD1Xz0wk08vsKeI1F3Z7uV4
Wh2+V0gYMaOfbpqhppfqhTyDZM1SrYs9Lht4/nRcVstcfGoKkJEQh7qS3J6wCtJnUILG9qsiJLiK
j7RzhW0wnacfi58DSk0APYMHkLPFsL/DcjguA5L92eaYx8n3bhNPrQA2ZGkFGkkfIdMj05F70FHh
/tbVkeLz3K/YRGiHT5ekP0n/Qqp8T3stCCzERcA9oz2JYoiH1+haUsGa+5vlZI29Q7iyHC9ve9i8
C5DKCkBsbVXrFQxc7g4N/zHcXztGgZKPFg0O/6Gp7AgqiVlfG0ACBXu5NUa1B9HaCD5CQRngQLeZ
5r/iv7F3p4DYdtfhRm/V9oRhjaLWKBrZTZLU5IXW3zgly5K5g+HnmpeyM5aSjEWJJqOf1J5Wz/bx
HB2/QP2T5SGfqVFtIOSq1MA7yuikMaOFOZjCmQbtDSsd5Q7WpMs1Qb7BczUdfi3GaXwXhh4ZnpV2
1wwq7fHVtSZybSzpSGPWcD/+v+0K9zSKGPZGPDW2Ixh9d0win22pi1mTP8I+iorFl81+jew38VM4
kabpycyau30r5CGuIHJSvweUHLl1E8MpsJybLPOcOoD50UP0tDz6WQvQBQkPjzo1gocU6Cpgn8Mz
18cwEXLi/GR6cTHJr/xkDrUgLdAq+kwzdkUpFaob30xpw8bSj5a5rngD4BI5QpoAdHLI12q7CYSS
9s5KaIUOiKOc7f60OtZGBU271uhs5VLYkwzKoixcEJY8hEmiGaABnqVX3JcqmyETjePcqi+x4tNB
iGXB5FZMOvULb+DQGaHiSzx6vNP2x2pp3ycofoNbt5dIAW9TnHiEh4RBeH+3owBmaV3LaG5wIKqf
1YmVwG5BWio4rvVzMGZu6Yy2CxhUW4q6Txxf/rL2DGdrtAHwMbAlDjBc6kp21vQQvo91Txz2j1QZ
rGhsdt2X5TA4E7vABLCFlfIoCgTG9KDm53Jb3ff3yVPE/Q6kS+nO560X68c5T0byoogHWcfe7oIz
exbTTWjRzW9mKHhGF2adLSZAOdvJp6he8Xb0Y9wiiXiKkkb3p6xosBQPSceDlnKNOHX6URtBVo2K
++FaPbCuDY/6fr7JbyP91t4JWemxC25Lus/21HILUP97Dr5shNQnPybEmjKQJ6zuDi+EVbUaMgSS
ZEnjORNgVt8AqMXAaYXD4Z5xs9lO5gBw0Xyn8zbeBXemJTCaTx2xsURuvj3Q9JY7rgmh1GSbiVQa
iGto9NiLjwmYBlWOJkT05pr6/hss1PhavtkKnNDd960leJVEuhqpJgSvLLeUNkqxovWTdU22jTEe
4bO0VkKEAML1LpPxx79R50NmDFw+0NC87/ukpaWhte9FKM6CcY5kd61dZNWsrPfIh0ggiQZ0V45P
5Wa3toRdLJMxTM3xXAYItYS089U3zp16rBxJAcgliYfR1QfwK3nbmva+BmV+O/M4gx6u8D/EfWeD
FDmbOf0hM4JdEobfJAFJ6475TV+clexcFAIp3VCpQ4WjZX9HAWU3M6TFSyZ5BXfuJu9cq3MI2s/d
sZgqeQWjpfh99DMm2NoZs4sWR5nrWfcuiy/uJk3OkesK0WQyBximh8ZN8/YSCnqD+rJvHhS5+Q1K
KTo/lYXbm7CNxuCyNP/L/7Q64zOvOjzh4sFy1TH1wpSbcUrHdAjMIxFdNqWk6YSVb4jUuQPfsxod
YR0w3DQHE0XTZRIUN5b8I5mnRCFBrtki9O5H+hR19ttpqvW17zrV3hBaxMJN+dv3oH89IVAztiDF
XMuEwuF++wn/zJVXFL+lisn9GUDGto2L3RN775m954/ATtLtbtQlrzC+Oc26GSFJ12VOyRTO7go5
DBTnZwxDsi6qmUWwqScyxAnRYEexf7NhKXhktV4KGuwOGKod52qVIcUtzwLxoVOPNf1e9kwDu4RC
DWeHi9/ItPLVpqJPoxKskXNiiJb3jtZRkdIKy2FgySaCA29IXZjOlGoZf8j3FutZK/z2jNk0XHgW
CZaXcl2R2sRkGN/8hRRn9eFpqBgoO1wDxeBEi9KvJhlF88xErGQgygCV3lMS6jd9DX4a2cP2NtrT
z9Coe8HSFKblEmG3133Y2a3rnn/JTdhgqSigEUp9ftlmYowOONVEmW2KD1kbLbwvF8a3xcnAFbXA
tqb95GOUeXs/pdDRA+IcGB30wDw4lR6zkNS4+lndge8AvvaT03Zvg8O/6UUjYmzxebkelm8dbphP
K2dL/C+od75z0MZbNzlr43bJJz+eRf5K9ZBDhSuSVClDFX1CE9uActTSZHgWu9eAsvU4/WcT6D0O
AMOx9iDehhOXTkt7Zu8vKAaeVgqYsC8hTsIaRJNRHOmkuSYO/yU3v9C0R//C61TC/uq4I16t+94b
CDB+4hfN4uYAWRiygy8dr3tsZcd8393Jbphuyi8qBF+fZRAp0t258p/j/jeGAaALd5YLWQFg5Ivu
HFM+UqGyFERr3OZOejeYPCgVbbUEQ/h1vv2kLskktW1c/o4gmdilqbN5Y4/Cnrlc5NDrJrpkoyVZ
rAd3VojWvpKvhoJVol/uuP6f8uwtwI0Vzo9EPDqJExhUJSw2M6Nd/4EsuXMd/BXd690TKbX0R9mc
rL2B5B9nd8nmQI0iln/VPxxnm7jr7XHgOsm/sx4lKKWZK5cPBeaQAPthufNM3oFwgFI9TlNorF8k
3R7jX9KI28gXzbA8natTIbUqeBLRyY5Qe8Heu+U+xA9bq7iPTNrzeSpf6mhmzp3Z+IkcBob3J1rD
sSYZY4buMkLguF6YM1Kd723VfCU4uY59/FHE5hYWZvL+lkelRCYPNRfSAgBmWBwXHE8yfeeQ1yV3
wYhf2oxSLXl5tg6QmKC/46EjjgUbLZ43qE4s78H+xj0gx8tNy3OyOefiPDjqCDkb2FiTe/Ki/q24
TZGDZnBCfrTwXHYbhTL2EAvU6dczp8eAxNOKnImwAw2QDG9kqFy+VVfJaXd7zgUODN63Sq8G81N0
SkyRt+UoTxSkqh2CuqjdfR668TQ4tuPcX2Eb1l0gkKbyIrXhwe/WQIJX1MDuGqMmnsz2KGG6buhA
bCm8qvVUR0Qn0Wmtm83sMITNHRYSrZaXnbQdmfIuEJCfHy7WKULh3YGL+7KF5FQtWjCNmTNLt9CJ
b+mjYnoPalYFAs0tR6yy6qjT1ScCs6gaD9Nhr7DXnEzvsCuX8QdgDKb+sOKyLHNTKd2MpMesPFZ0
OJEwWEH22TBt3gKhOGNojpEDXSWC7mvjcqXU5EJw9nPks0VsMfRaha8Mf5ohjOQOXj4vYXczIlTP
fAYbljX0MBsImLNUKAiTBonNZwUNnX6MZfCA59FmScVImsSuWT1C7vsMQS7ogAHaPZlyERMmSTMe
vc4jtOkae/q9PjVM28O2ASsyDYeeFt9pdbIEkGLj0WdvJ5Wrk3q6RGGYEpPzk/k+Y+jHCE2v1YTC
ztjmy+pGX/vNvzqYOjHyUQlEGeEQD/Mi3YIvbUM12LDETilHNUcLDDlA00vXEzrzhhVV1DvH7mfW
mwHYv+JT/dsyI1HPt4X+gGFq5aVKSmqoBYIIOmjVC0Xb9gWl8n4yylYbZCIFsRrrxvO9evHGA/B5
NvmGmfzKX/Hgk5Il20li+9Ph8W20GkWc0raHTyFsstVQmXGuVFKNrYiqH0C1f0c08wmATkjsqg04
NHFdv+RyBEepllwbF5BlTV7COLYOfhBYcvEUVrpruJFIHxg3BA1SJMDskNLjoEE8QX1/iHFMHzxk
3TJ/VgukICQI2EF/OhaIIpZVO0egqNBA0y+olSbxAgJPVeW9Qk4TrgHk5IcLkKkvP5mguicnZS8y
GK5pZENDd684cXXwt1aWXyVfpY3NI9C9BHCvTOAGiLsP8g8WVuSmFK6V2C+5+LSDPXQ2MEkbKMDa
2lKCmneqzuIgoEQZSZnkn8LfErGkrFE+zG+XdJVnk+URdh4EFa48Tr8YQMFyya+OqZFfUK5OOVCZ
BlBD5ghECLYY4v8NB7yYyCxcwVmG55UuEpAWJUKveHzvE0EBYRgPgrT84H/40102aipM2NuBPx2v
gXD9VyC94kpiq9jB3HqkroUsl8IzMwUtYgGd+bO1Ud0nqMl20esKPqC33QtfEC2XU0rYzBtevWL+
VZWyVLBDaOC5XJV9OQheZtaHK3SOnoIxhPsuuaZhwDHS/JIKGbCJCZwy0jXqn9xht812jUeA+CRK
Osm4nZ0+h+1lBjjqFCT68jm6ppfMf8Bx+hC96NfkteO0QMe82Eq94ZkTJ2AlxDGMLddcSHS9PjC3
MJCwy6der5eLlf8iKfnMeLH4dK/LpdcMOBI1ELvkQ6Qml/MIP1khruY7F3JzHM9J6jppOjxMW1uI
Q6TuH4PF0bNYEgrbUmlH4n/JLhw91b9DyBwaGc8Gc5OISY06J8T0uguFmrCyAD1xK+H5RSuNp7fM
FVE7q/a2ReURwnj4VXmd1Eic8Ce8fwgJyL259aDZ7PRF2SarMSJnhiPsa6GXC1nylVSdQzUFEHOZ
rbCuurcuqjjGHHMQd7pFP/4EzjmjNQhXoAtnx2me4j0ip3Ye7IVndB77IJbhtnkd8E7OYGf092+g
wCSYqmjofwIUIz7ZWDgLCA4roFbJSgDUVUeFq0xBtltDh43jEheBJMj+ZInuutu0cLz6uqACjtT0
uGoAMl6Lj6Io5+rygCxFyZVM+n5K4Nv8Cf5WHoCRxAodA3jpjkvZclg/dEGnt/ueUr6lUnVdzzb6
Vi9jHWl7uDRdTyDIDJLpt3d2mWBNBkJKGe+7CTskYtAHyOzJregog9Ocjp/I2KdfDPPCy80HwEwa
/fv5UidKGzayuEB+zqwzlVmYMSADSVPh/GkVmxx1JiTad8aDIsJBRVFpvasJSy3UMEm3R41k/kst
8j3M7jgJKKCkPKU/lJ1M/Cf+IHQlT0cqFE5jhw3XJ13SEPrLC4qWZzmhnwE1/pg0pwL1V1ntk+u5
79dDLtBw9gm5OqhHQGZrN7OGwqagi6OGELQDJfV9NQzOfQa3fAEijCe+ZYQ9bwxLjdPvXc7QwC1j
kBykRwNQ83XbbQ1XMD+Xi+dDFRjV1CcoGONa8xK3i/HWts3nCK1iQczZwstJb0Mh5KDUhxmW3Zmw
DwR8ZJh4ALw69lB5qF8qYzTMgmrfmd+AQ8WxCQsOipPMIaUInjBA+2GG+hmb2Njlu5C/Nxv9yma1
BrHnSg1U5nU28Nt1eY+mtP07b+KT6mYkWW7QG6k1oZ8kEqjDEFyhBZhAPsrizQJYOO4v4RGDEVZj
pBYwbrkfF/IHqfIhLnehiduTJWqFjriwQoGxFcDP+D9wCze8jCcqW4B1GMK5gXKNQ+ZUQMYGDRWk
e0fnV5B70xv/Sx7u+HCnKzrlZ1dlZA+Wdy+3qZZzTSNHC2nxHmO4/VElITrsmMg819hhuxqgU/1L
4evUtFZxz3KXbTlqNeiUrP+lxpTOF2r8WOyw40yT/yl0Gr33KHiTpfushXORlrCyiYaq8fwaZ+sZ
hi1OwEVZS164Sl/G1ptNr3zn215k2UtUy58/az5BRBKb9QzZr5Izg/p7TszjyZz5j4ElwLu8r7Ma
M9cbLspIV6bJoyL7Cn63sfuFrY/kLLI7NMn1dbsEbuDyajtdNSshHsswJ6MDNnrQQPy5jhTyL2Kt
pjTlQ9eBsO/eAT0R+dJWVW/mx8Tq63eJZlAhEwXkJSPSg8hv61b990j/Fa59L0hSYjWOshV7SiHe
Zv8+SCrsdEkIry8LUjYVEWCM6p7xX7g40iX8X0JcFhIIeEj7rtspzQCb1O7puNKorrVyZfrakkzy
xKbqT1A1gKAcFaaEw/H4FaBhXg94NTIjPAdlA6yegYQsavt5YiRlq8glJexOPz3fnyKlEzdDwaQW
yo1FwlfzGU+TZ2nkRw89r5u0Z9ThKGTLc3fjOjfJ0REJAzpBL7qweoPcVgK5bQoEG6/FwlzY7zuM
7N+jOZdaSDty6Bn3mf21xRLlKOhMUs9ROZW2rI8bnniTh/Nwq3d0w5KdTKxaIDiweI6lqQncB21v
ylEflkpydQFhO/h1RIJH5kMvkgdyF4obH843YaKzBbXRBcIPsyn5GT7bsYnZVhckO64tiE7XA6i8
yORM6Q0KXqPwhlNSMN+Ja9ASM1OtZbIKiWUUyX3BdaAwBNE/Y/pV7sA2iMd2W5J8CZEgLDosi1az
XaVFKS6C1X6YPXVEzjAZPLxk9rSWuRzPJSD6VmsGLhPLERQUcPV3wLApusXkWcM+B2CsSt8yX798
9upBLXP87CJHuDYmvh43JOYwO6nnKXewCtM60WZN7m5KldlFKJFcQB/AeezN7FTZAXn6v0W9l7NZ
FsTMUHaduIMZx1R/MyHJDHVfjSsPCgSCMxKP6qb23qs9vioS41EHZku5NpCz4L3/odkC5pNrDgds
YvhrLbNImcih64HI5L9yHSiZgYuaZgJ55LkkLKwyltGbz6Rdf2Jsm/ZZr49tkGGwg6FHsERMCUpU
zNnVSgN2D4cBhGqRDLaYvKj34jFKRTlif/pn+ZHvlrVc0OsP/cQW+44ATy73guIoOMFnjqR5ji65
/297ObGZrv70o9w27pYNyvdCCQHhBCWR2hVeNpFb0BzQJpfbiMta6X7cYN9KRTA3IC1TaJbgXYI+
hGldhPQ3zpj9OdmB39NnNmERAsdwtRITcBv9EQwHCUoUbV57jfM14JoBHIB7unX7C8BpZwjFIjQm
W8W0e0PayciivSNaJoIVuRJBRMP+4v2AkvoEOcRiHDhziBdcmJdW9V1muy7gtssol8i7jfy1RsSh
jELNtuf5g+yfr6AS1cyQxlITRK5kb8eMCXpx3X3tG9nBieauZBx2mSxz34xO3hrsDbUTxQtB0u3l
vMjHW5YANdcuQ6EEcT2LIkegOBAvnsRCiYXZ3RPc5QVBCCGDRiZLgAkVHdQp2TqLKzLfmHl1TieZ
rx43SF+jGchZlK7I73bN5JW91O2/vBM9n4HvndbBmQGFHy1zcQCbGCaTgc+unQXvpxgW0nfjnSud
KmepqqNDNIbMTs1hyaEAlgrYU5vOnNSFeWWasmR3Ce2ckPKR6c82NaRKRDh2CtpQPUtOhf7Q0Dsm
uawsAd3SuuIibWN8TzsppSv6OuI+6Rv/8SVO7ackGJLWWf6mto97LZMv5xPSvXBEW9xqCe9b2g97
XC8gz/9oCT+fgZ7jqRNIBxzpNpvWq4YR11WPDJsgVzHnW6JVIt8IIlVYSie0KXjZIZGJOwZH7rqt
hhDJRqkxTDsihsBj7oOjiIqJcGKEFhettOrIxa3s7zSjeSqdvnhtei5EPi0vnzRWuru9SlOoqY1Q
B/Hux8YtkUCYNxs3C6rqObSzQyGQwbIwUxYGbBPGojwEUGEHADx4MWWmabjzMowlz5wUtZn6BuvQ
Rf8jmeefXflCR5RZFyCX/GdJuz1TyLka4L1XFvy9ms2kT58Djdn05vf7VH89TzzeoNWfORrn8SkV
Afd3zNi9kMxSMsxqoGLVaJHNX+3cJmeKSF+S15wkrfIqKVjA1YEwppJwhm2sovcg9IUnZkRye6fF
WBhizUVT1xmGtkiZ9Kd0O0MMd5XLlj5C6qFj8VWB2bxapvkiz+/6eIZF8ygXgDzmJLq199MYxWWO
mdQvaUeNEfLxga+MPLFx5sEMJDjR0Udtny4jhK2VAojARLKsxjGSZiXYaKNVjLIsWEucSd5XTBFV
TnJTld8MURnsKqL3AZme9Ckgx749K6Vi2xl+k99q+TumzH37V3LbPmI7y7EKrPQeSjs1wk0gdYLg
mUwZm2WCIIO+kXU+8BtRxE7smPBiqhWerD0tcaFkhywhNBQC5lvSkvNXypNV8DnVH1WWpPJUi8Rd
gyuAT0LAfli0SLP+GhFkm0/3Mh3A3eoydH5efcgCupoysOM4M1Gz0YbuzxfdEYREWNCXHw3KR8EG
o+mOJZmCzVrNM2tDpoggQend1zI+KFsAkrQX3lU6cRJkT8oQpetdIbkTolpEkISSUjD5VORVtfyq
m0GAAiqKlp2nH/BZnDK1lDkvCQxQzEbVx80tbY41p6MF1E8RNFsySrOI5gA8IVCFz3VWSZ013eF0
kbib/MaTJonLMmKWjS1OyP6s2ETPPPrP/yViWKVZZ8BJmA81l2eZR1yiVIF9eEekJeoCaFpJbTqD
VMr7YzoF57MAmrwwdmstH9qd1nrWJmyl+grpoQ1gMG47tTN9aEvmKEedylvWwLWuW3io+8hxgmqt
xsVioeZarOKqfCCRrMNAJoDmcr1RlNuku59IaAxLxKTHbbNFqiDNntLhZiT22EeO5ggx/xjW3cbt
KAcOPIj7ZKjMndiy/CGlFXBazggUtXZJzckCoBHoX0/inPMaaaf3KNqEnOTDhqUKEo6X501z522D
xFCTaUYAAdB7X5YeB1+Gb85FQ9lsUU2/1RKEPCl7jpSJldghK2RaKBK2RPlZHlt+Hw+NkGim1aX3
WLfXD+hJNULwEvm4rrzVw6Gkq2vf3QOajVdA3TZwsFNvvf/vY1eAM8B10/ygWPmYJfgPXLEw2ZnU
7VCT6XZXWpIinSYFYs+UA2guPw19EcaMq8EnrrjjPyHn9dG/Rj6f5/Q4zLcx49H7Gc7drWJnR3sX
527RATT6JwHV3B+CCMKm4iyM+4nQdL+qI191lbpPOWJBNLL8c1BmNF8dfXJlrkOl8nvD89xZK4Dv
PxOtpyflFjnW+8Za4q3g4518rvSNmo6JG7koH+1viqIcWgjyJ6uq0K7MnMoPGH/QW1TKpNwOTSB7
pRVOEBdjaBAA3zhUltAvizssqVpXBEE8qXnkQ0hEnMYvv3quW1q/O781nOhQMtocWH32A4DKEbj2
9vjMMZNwqfb+p+q2ZdgPFl5WU0VU6JcUVQzuCIv9u2OpV3dO2DbZkMMwDjd/mmhVmEMQZOTKWZFk
7ehBsUHC/OVq0qdX8048xgPLzK7m/wBPg6dI1WcHJJbgo6JO/hUZNwuJ8mudFd6hR1fzucwc1ImH
kMEnU3rxq1BB2I5PrxaxPwfA+DCWRfFr/qDrIbQ4SMQrU68KHB9uAhztGVdMVXniSuU4AIDVVn7f
9YvcwlSizxQ9YQY9lGvm7dCBj7AeUV9aZfkms+1J5v3UNYiAUUguOYZaOPGRgst1ZTCw1KnpTIzJ
mEkILDKAviduPAn/164E+/9voS0y1QkELMtApiMzLDAnpHA8WkYoYhss7If+NOxNb7V5zJVE5nxB
PUNmTJOApOFDwXZXDxrE3kItkmhsVGOoJd4cTd1v1gR7J2x92+JVnLupAX2e7G9skBRoKwduk1Ue
6qXRCQseIWPec0qZvfQ26gNAadNEfyIXkQHfMQMsxSvv7qboWfcZnffGMixv4mCF9yD4Mtmw8z/P
n3p2mlHH01RLu16KN8ZQQkz5PrTBgE++DhvNMmPOb3j390Nw9+UteWgDvvptkWF8CC548Chl/111
fxAi1/+lL9wFMGZ6AlZWdbr9lT7cfAT46dkl/O3aV1GDIBmIpq0U2WNTVYoj5v8Ld8HOXdNl0xV0
Y6oa6f7nu6YNuqRzwD28u7OC5eKzXUlkuof/KhHxxFK+ndghZABz4vhgq3gUJhvBgEmY51PnnIeN
b1ZuU026RvG3+KIk7lBvO95zEioSQS2g8YAqno2PQfPzOO9yN3gcjjjB3lKKh0bubupfXZK+lEpL
nkYhIv5pQZuB6vafhiLHJcr5WNJZ/qxZTGPdi1rAT/dWCrwhQY99p8H4+8NQg4r6hjKkoFsQpkvw
pCfyM/pB1MxDq6l7CAW+S7L7J8fmxxnQncSKfTHVYGUXhKkodL/qmxY+xyQ0JwwS0iSSnmwDEb7o
t+cZ2vobfIUHI6XV1aebi2ef+Z8AF4Q9YmXF4tPpbBc1tntXorY73OujRFfbH43iVbcPi8QWr7aK
ZRty7Y3TVvg849K1VuBbxrX+1pBd4loNzr+AzflBr/s3pdP4jnlHy0I0yKUJ5ng6Vr4VqzD27r0k
k9e4hufRI1Cpic6LD49dfiqfH5Mt2vezZOHx9QGJjebXkns5jMkjEqRDDLyR/RbyDq3wy6GB6gGu
jV62nE74rbS8n7xhafD6kVDYu3vhVCwlmFcF2amWdfoXFT6J2pg3DJEh1U61tm04duYMWRwsoP2V
VMsl2F+fyoUQ52tTP4f/Lf46UWmN/sBaZvTFW1gty3du3oFiBzfiXSre6VtFfNtje711FtCoxXWu
hSPuTD2FvW+FZF8xqARB813/amp4HPCvV6KomC1LYvgslHbumPqREyZLYWuvpl77ctEA2jPM9FWG
XuQmC9EFnNn1eDycse4LJ7NZmf0Xwh3V8qAEcQZqtdulnQwwNi9wyRB+1VwU8j8dHU4hJktxvWz2
bMnNtexsmcY5+ZYezK6A1wwS6ie8+nbTewzx2bWhVMYp/RV36H+6cy73qNgo7PtM1bsUWIpLvdHv
6cZ4WTH5fNq/NA0a7m5iDeTeVSdIDUdmYgO6rEblqIi3zOOfx29pblPeDMn8pcUJBRk5cYXMLQOo
M0mVUT9ldd63f9oi5NqkohQGXJ5r2kDm9zVHXbek3jZDrYbGHiGkNqxK0x6CQS7329pgXrcSCaH3
tjiklRd5fKmSfpoEZRiPSlIkvaHH1CqDGySViKGxpFd8HoFg1DdPhQjHK+X8KrBwZ9WsCE+aPRmx
HpWmHBAnkcUCMLPc4eGfC+pSjsx5TftfZxy47KON4rAnIxHjeY/QX+XeRlflZAQQcRzBOWwQKO9q
vQ4D3HGktLyLxrwgEGvOVlADaFMOEN0ZWV2KxVkYsySjrG+hUCRk8JDm6moeVnN/GF05F5lYvxEo
VN3RBkJ2XzTptZ6phe8xsl/DoUGZHg7k2TosV0ABU8dq3gpdtT/ZUgRoCvqyiGLnpH2gty+Ec7KG
yecSMEJcJcPircJZGRU393FW+W5bDLGp0+gFdrNK9kEhmImd4JWVgd6TBkvXflAvi/qerVgulAfg
Pu2K3BFIb1SLiDMM5T0FBcNcJEA4vCQ33F/avpuAUI69qCW0QLUIL4WWoGzMYwa92fb8jre3rkFI
ZI0bAy68qYwjpx9r0sACX1on5TUWyLoew8i2HVegBDHar9aLHK01/TzWlg+XjaKs8GJ9K7BaykZY
ko0pedi3NfAYseIKkC8ambFGb4cGpG5NzbhrZnF+PGllqg11w3n+UjEk+W7+fnbr5N5/i6V3dGbK
kqmAFO78rRtRy/3Z5qShzIAHRvRRjrOtPOnwUUjjbuwY8vLeEzTzoZYuava7FgpcnaJZjhJPtvnZ
sA0beTvg/E0YTD+cgcXV/HXP7PZhf/nqOsLxH6A1jFoj24DcqM5TTpoG7M7b4HygekRAFZY6B/Fn
IbeNuPKqW0rmr0EfJEIn47zjJNUk3TEbN1ISeCHHSJitMWvxo9vmUn1EE98WjDh9HyQ8jKIDzvyf
/8yeMPXX2fVZuOBcoIcZS49jxFkbpKx+riEJ7dDJPRJeHnGbqp7/9d9W+sJw51U0kaCuOfF97vik
3khfovCKs3b2omyq6gOx0is9wiglwWsblQ7E1uu1m5L2fVtuaDBecCkmMoRDD952iq9xSpgn2dxh
UPNQFU4JvbsA7j8VtaamLo+EvGG3LDuxpcujrZ6t/SurNoyv2t3vvgkuZOIkmkIzpiiy4RroaYel
jMNGy5fJp65Pk/xNuhgAYohA887LyroUvSN8xCX94TDiZzLYT6/dSZ4yJduglnCh5kooQKMrpqdi
RMlQhVQ2OVkpEzVky4y2cPnVev/A4gaM8GGjaU0LogdcfVIj3adEmPFGkg12VTRuwXKA90++mwCL
b44wewdc3ZtweVQZWOf+zjyW/TrUss4JZQo3jJmab7ycusAwWyZ1QcJQM2dNnfvX1ldLSepDbQfB
7Tby7XBbyYVRdec8yU5iwB7FH/KA9llyxomzIIfZqqK1uYfvGLXfyAK9nBqWg4NU6r28yqFSm9FD
fokwQsFuxZBuUs3XfXWfVAqVjXODBkYcfpZNzh4pRsMpM4MqMElJyLQSX2NT03965EXRipHlUtGM
75HQ39qywN9wUihSLHmGcSgiUKLZA+csQNyZVXEahjiMA45zsEjIt3YTlxHeP35uDV7+dUL58Kz3
k3sPu57FMclutKx3abJJu+hZWwle3oUfQuYkTceN2aS/VYSPMhiTtomJOmR58Xk8QL+chjgJvxRq
LQu4GROyfMz1tv9mAkq6J/MlwqCKoVIDKHuRdKwqUbFXrALfDJwsk7dSrTUPJnpTR8n7MsFyPSrr
ET4E8RFgPcsDlbbnCzpiLo7TUBI6WCA6rmWWzi2niHBYC+7G1WV3y5nrw3B+zHsdR9YUztwcqljb
QFXMj0A4CsJmvarbTuuNoNwq1w5VXQK623K5e/+Frrmc8ynOBj2GJosinPjoE9mJAWBOHFoFzsan
PsDOZhpnwV5VsZIwgccg/1+aUnXCzoKdaWMmmy5qpbqefKjPfsJPkY+5sGITZN92grTpZhJwC2kY
knbhfAdtnRZCukcwCQA3f93+N1oBuQDg+adT5Qm1IUm2QwMmIZd44qbizFkJiXF7gKNy5M05VK/T
RqMWaVTdJYQt1icWlTwsWbETyWYAoYg47e087rPppC0r72YCMEgmFQ0B7lVtJrLePl1pGNb36jFW
wz7OPR8Y/8GIQgrv2UNu+Sv4wdqY1/y3URem6rklALbMBJD0tqw5X6LM+WmzSFYDn8wptg79YCTi
WrKpTO0Z4qmXIF913CegzlAbQ+xD47ukRevTqFpffyut1Ll2nxFBoqtuHUAn8+WATw96BC6F4RAG
a+oKTUoW4HVfcpCrgzxvX5cQ+iXCgegAwQqi+a4sneQN8/8NuE/9/Y0r+KLt2wWylQIAfGgQU2ZE
7AyQ15DlooAPpOSHuoCCAClXe8Os8GdysVSxSYoxOjas37ZWuAz4kNB/2GiTLBlQMfsL6CD3ulU+
t6tUZXbTmAvPGr7wQZRYk04oQ40DntS//wE33LfthlX4AWzx9N1OVeCFYzoK+0E4gG8TD9OAwKM6
3EWqOPRkhZC51KxODxsyXIcskqcqA0a5ooySJntSteevNE/1ERnPvOP1UV2mklwX/c6kgDF2YrWO
v38FOagqnDd0eHgRF967IYNjxUbBZlfYRTKiSS9GYPKea+P3w1m1v9I/WjJT+p0SV2fYFSoCKv+Y
BYQRDEKv+ZXWTohjbW1kfI+BSQE+ISXNtSBRpW2WUFIKU61+jxrU2NUYBVWAre7xfdLSxS4q2KZR
8/25lOh5wcABmObGuGPvUVyTqlei066e8wJStdjkUFTYxKIz/NakHww9TR2NnreFXDWIUGv2e0E9
tryq/KmohxFzhpiA9iFp/Dn2J9/Ty+/b3Lwm0MIxcqGIqbKj5aAyoM6xfIpxA9KqxTYaeE24bmrV
8MW5cvOrsaCvEvfN9roRTJKFbQky7bDjLsQpCx43/lRHDzX7D+ZmzHS5UYB0PWsvznnFCuPT+wBG
jWmoOAFTi3+ymAXN24ktDjVJMwzTOJKEayPpWh2drxrFToUCP2emv4sAOeYG4B1N6AKd5pULDiYz
Krvx/wMH5o6k1k18vK5p6VaCIoa4YdNCnGLV1/HPUqvp4CgCKum/FJW68VD3ZL6FwksuAJbqQS2Q
2jQiIkpV6D8tJzOEmdgBapOK2WWsr/yZ16f2tO+KhtNKiiyS/i3v1mgqeeXolBtyRlK8SJAYTOmX
eWUoNYeNhN6nOmjetLnmQtsEPT6BJbmf1OI+MGOTBh/+n7JaY3k+ruTjD5dx56Zk5KbXqCQMixrY
I6cIT3CmoB9QzqEruRCP26YdO13zsXdx9BlrtHfTJgVW+N+E/CyRN4iS+u9F4uv//X6x2jWNP+r+
HGZ/6z3Ex2Sj9ijSPr66DjWAN4u6SaGtKK5CoAZ/sP2LwAOyaUWhkk807aiLwP189UazVb69sjup
LGkFlVUEHkCdV+R4dwlzarQXwj6AgfoDTfzwmbpfPDeNQWmRoDtAWzYo0uBarY9TnBij2LGxMdEJ
4StxZ8luq/bAmBeEDC/TO/WAIUkv9WnRQ0mRPxUtJesPUhmxoWO4Mi2sNUa1M6axRZPTXM4TvUHD
NNra2+INaRl4cWjPjhZAhcCbjZwjA6lfFllo5BsJMqsoTWL3PeynzjUVDvcYgy5aE4EaOqFfWgII
Q5yo+BUtf6RiIrw2aTzq2CMz0W8eqn1DqUXn1aYyMzeSNisa/5+EaS9vp8/3OpohoPvQVFmfalw1
b2cXqaMCZ4M2Fm8foBeCrHmzQRZRONb69qEvThqrawTcegoR+chlAXiwF9Wf6PBkXXWVJ4LAER3A
XeowJBbJxpyc8GEJZXWpTJl27KN/q3+fPaP9uHFF9ldJsTauPyiYIImAHO8AQlV2FuG6kIBNltIv
/F7SeC9LUgwI6roavOhui8vbyQxWrlt9Ru5/QfpAFihpPKTELeY40XYlDP1p3ZBJYusX00cH4oU9
co/jGZSqc5xfVNa3SSOQrjrihuQwpQ9ELvOktviLaLBr+w2IHO3VvgIfTzH8kVOIouvMml8sAt0E
R6L5yHrfNcmht+lFkzOIjFZyjPJUA8lFze90PSaB/QlwXmdcim3T+pGLazkOx+ycFC/Zoowy8Yzf
K1bWWRabVLeofoiBqqky65mA52Fv3nNT/FuiGJwp0vRt00nxYIKB+hW7+gPkZWRyboeUMonpDigS
35tbOvFJ89ZX3oMJ6MVLZ+ZEDAmwzXYKkcSoe/pbVIm7bEyRePTS+9JFE0ubBGn/5EOnQb+GgTol
QqAl09Ps69FrF7Crk7V/+zYSGkmFgglxB7dbxjfEqmeMmLhxzN1krhca8/WYOevj8dMJrj+7w4Nt
DcC83vTeR3vx+/se+YYqKRTRiNRasJ2x7UWJAjovS5Mse8B28trnLSo2TgX/kwpBfA7YeM5BMlks
CoVHegqQS9TpmItNmPj8hNVLE8JGit8d1SMcC40mRcF6l4qYjHx03RQ7rsfuUPjXvZKsHjsVJ9hD
9mzSwAkt8iZDFHsz/lbgecq2cY5fkShKAYmOb98Swcj78oibzNLx9BVrYR/3Kqo8jwNUFUq5hD+q
bnZkOyAJ0DvtX5JLkHipnyfxfQZ3yAX0o9HeQ39JO8JknNA11DTh1WnmA8GguoyJVQCjcqDDfHHk
JMsxBFE3DOgt6ZdGKUEl076lnYD841+pbsF8DNfYSMp3dOd3swiT+C5afFuDRMG0Y8Op61vRNHLu
409W7e7isr7F+kH2ahADYrrgSDwGcy+F/RdWJhBj79zCwVo5Zcn9RNYZg1cIn1knKgGhgMpN66Pn
ArveaVAEhc3tofTMd1Ge/CMZlakuOegJbG1wEglEqPCmSJ+PMYzeGiJ81IO2Ch47cH9QQ6/oXnon
0kdBA2iC8aL9sDszlmOlJ62yFAHJ3FeKbarrhpAll9nzHebjzbyaMI9t7NEbh5OSQ1HDRvIO/vrW
6WLUvSaYJM0mNZz4Bu3yW9rvWa5xyHOmx/eA/2htDjuJ813G/CFt/ohLgjCtIUMF76Yfan5Iqh/x
sv/kdSOWJc3G4jH8yJ/7J8xzO/lWXox69OQanJXEJc2MTgkiJVZf3vwGHjt8HKeod/nFLDaXnyFN
jFymAfk6ZB8zwZNOYMUDwWHvM0vnesXcDvohU2qL3yG2pQ0IK+rGht9f2dLjQ+zbPblyxhVQXPK3
1ivmF9kqh+Zlil2UwotHAMAX8X6hDGzzELrXhQ6Jo36tc3eEpiwWTbQjvDJ/BhHM1L5W0+iguhIJ
kj2xwURQWGbmdGkU9rlionINqyj479kQAK4Ccs9buxRmwiRycPdW3sZme5kgyo+2YAbs8g7rfNnP
iuyGrUzSfllMewnQ1LesTMU9PM8xMImuHYXSc9OmlkA5mhYslnFR4aj7MCwZcDF3xUGUhyUu2O8k
CqQPkoyGMKGwkDN4hnapfiVmiT0GW3nKrzlSm6+kLXU+ofGRChOuFMwbXR7ybpzndrliGoIkQg6Y
D0dN3kGP/gkLaUolPoXU6hMUUMiL/N9pot3EQqI0dHhEqK8O2tCfsRNyq8pBcZsMfn3xOhtwg9Vk
qSM5IQst/A1+R+jzE1nIy2FZqkGPscCnW4/u8wUbZR6Y6n2zTZ0q+QOcjXriZMPlTg4l7m66L3bK
uvcWli/OJu1ZuHEHi7I2zWXbqmTqLpdtzwOXgE3F1Oz53T1McnjQNJLZ7xTVjF2rRZ2uMmc8b+eO
/FiF61HX4mBH7aBZriiZcskzuZRyW/AHB9ZqqhwCNZL/AA0rckt7eKD3H3LqUUrW/bjs0oGbUrdg
3b4oQ6Lcd+15xvi1dObGDwgYKTKe7egNYUUNt50Q59Pc2khHj/4FS3yLVgecYmNrd6ugGe6K4wS6
hVHA2pQzboL0/g28yr8IKfFYzvoNuOKFalh1vbUWhqsqbkjzftzkHaMCc5XuRr3U4kJr5dfU66I1
DHMdmEdOKO0usd2UGckCGSW3/dLKLlIR/c7aU0yo/72tinz/taBD9hwlg71AiLTGwPZNX8qpAhLu
nnaqlzKjhjVPZ+tXthVeJdLyzF5sTOS8tNiSHCa7jit6egRxOCJB60J4FIzLRBY2Qpu+VJnVbqtq
yWt6HikiRr9PeoKxERgwXOki2DBkxQU9GzVfal2Mn+xsoYggC+7u8gw4qyRYi5qc3Jb1ujG+PEg0
zPUROVzAJrPiIEMRUFO8wH+pe7n5Fr7F2dGpphyQSPSJq7/iusPoqaY8EX9Psu1LREOOWoXSNbOK
pqUxkugnXmBRXfmi++aRB60OkyrEtlXE6ltdk4r0ArIR/5C1DI3ec7DuH/B1huBle6FYZAjXABZ/
0C53zEB4PEHsiTzXmc+NkUhGYo4ksMzXTyFEvDtLswvTx0JtZSXZwaMMD9bjsZnyibn0Vi0bOVE/
9mZ+dBSRYNV8h9ZpdCHhUmClo9cHYXiZRXVtf9WVgQg34f+EZvAX0ZzG6AQkJhXIlSCjbUu/wB0a
wLH22pUrdIqmw2JszvjBiKIBzFHwxKi4uE4KaZSRs60ImN3NWZ5UmwDnrADl9n8wqbyGjy5Sp4kI
hRx81euAq/wyn+7eMo8BvOdGxv0BlAEbSGKp/Q7bWyWGuc6j8QNiQnRUQ3G+7YnGIvwOo9GjxJy2
FG3UGTRiRSFtJGh9Osr8PA4faJ+cYvb/Lg5c/XpVrt6/g+ELM2pox5skdIuvfQPSwU+oZbQZDdRz
UDr0pYF3cLpqvmbvkY3GLrN3+x1OmRrf6uadwFRabsXX0YKGkA9THDdud9rylDlF26Cv9MokZdEy
ILGBrCssVjatAZFOduRs5kXr/MlQrK6SYWCgQ/lkQbFJnjstEZ7ap+n+hwPAhBzZz7O/xPUQycDx
tla+N67/LbqFgiSeuiP/gz3ie6Ob64SRBQqQLdGwHlLZpPJYVqlho98T9z9jL2ZV3KjKFuBhkwHp
L23fbwnVJvZg7g4ubf21o6MGxJ+t1thHGPuLXJFQsdmAvitO9FShNxwzTmsE9T80zsh6ymnLo2W5
IzfR64A8jfL0BnWSjSUw4E/jNLbPOBScs99RnTiR/mcJfSmaYS7cmzvE8hii5ECW2/l2NfAcK8xv
V0EWGDPQsscURDYtwdEChgQwVcDI7Ehh+EDw4XzZX3lUMw9FMCSCUFrAnHNRjlOZLtcVJ9hPfNSv
y1KTlLkEE4K+GOVx0ui0Y6aa/gJ7lb7TzeWuKwd2SRy2gxZxhJoYsFxLGcGbjwlv8ivscTU5i2DV
3KQeGiFHI7OKp2MrG5p2YGzqtfyxohNMG5RE03ZOzqe7up7ifsDt696Dp77Ih2SNHo2ORK8BtNmn
st/xBtULbak+xelvXBBUH4guLP4TSpFsU/AdFPyhH/REEUn0mMnJTCwGrlUjUpPhf4SygIuQwmKl
BMFnGta24TRaUMfSzJcFusGZ0P+NtgWVrC1eNlYu+2P+V0Tr3GNnq/6pygBkdHOZJ911HKVlvdo/
jOzMSUJ0RdGIDzfX5OvVs0z501TJO95JgrU5/96ILy26sL1ItVE45tCCiu+98WqzeuLnFdD8dHj4
Jp7r1CSI9RshkDX38YUnsHXYR8aEGo4jcn/FZ8GeTG3ag0ehuvaTxCXjmMft8+AnmVsgaaBmIy1X
x6U9e1hcg4S7Zjqjgin8R/UZilnmr8iRlGfPY4dHYNZnZcQGcFyFd+EQjsHYun/dMs+T6reJKzfv
+LDJT4O/v00J+c94AYM9UWDV7NLx5hSuBgUVEvAYb7WrjaZc2FixZKtosi+g1AlUSoLnEUyUjbCh
eZVo5MKc2N/VUcBGM9faYron4dA1JC9wCsEURdR2ZHpiI/4W3lZnOwI4MsoSuNdCXZpM5GY3Xpd9
2SvtdW+nzkb+A1cOfFnHYv3kGovU4hyWS3TsZfSeTt62XgtLXeTdi9wy3F20I5HS0OlvkWlrQvZw
oKsGh/efn2yXnFVevWXMui91V4Mt8t5IvuaBPk6fvAV5Y56zPh42S9Sd3+ngkBYPjO4vp334DRz1
9Jkb+3QMwEfi3P0dGAG+xI7r1hHrTfjueiBqFX9pQ5wEBUX2m6MDYusnv3JtMu8bJCkUgQxSiwcS
HipU9uZIvrUMOVdA+QDXD8blZzjIySgQmZkMaRZs7LQRZMvI1Nd+uE3U64w5FsKwwCSzxF1SLHju
/+ihdCFIATB1x9ZpASN/6SE+UQ72qrIBTXy1/64qnQdu1KLGYJbcd4pIv8XsnYvEmoAbzC9hc0co
3pfFyM3bqprHAY+OKugg6ANjwvAdHODbyLpP02yTfEDKPB4m6Av7WnTXuigOFdONEbNANX1/tz+C
yK5KLSCM4JKaozx718SOOKURBNEucNQpJ8FTvQehYAlHnyAavJM6jRAyMSzmEZdBXtLgfYIEL2rv
kGqDdsxCRBKUHMjMpAc+t6TswqU6wvxXXNbwiUeI5cKewdiJnchu/na1f3Y++m4c/k7NgB02VtWW
WU2AxP8svEgoDn9EbwQjAzhR9WTaNiIqflDmMLi4bPxZ4Mxl37DWimYqdi6fmseYOnIOm1PM+sQH
Tjmf+JE9AlbrCOUMO9RpC0RTaZHQG10GKDmQVBEm8sa9TStpQv35lhPaVt0Nl1pGBwW0NxBvvEY+
e3a3lsU3fKjJzy8oLgOKvzpS6Lfiz6puu/sFfQO+908kIAP+trCHU2J4heKHEQ7/5JremlT9aTu8
3OqVfLeXU0hkQTA2i/jQtnFlAQjES7Q8v2wfXtMdlepPLcwPtZqCDgEhI4UJwQoJ7edDxw7ob0f1
6O59doVcudZkiQgpPlGtqbPSXPNOhALWzZGsB6vo3g71MmImdABdkR6WHTmeXUHln9bwYfxmF7Ad
3+s9foV+cdN9QhQ2oJILxWLZM2lIvp9Z5haenYGaJytpkDXYbhqJdm0dhtCOu5p9ge5y4EKCawt+
2GM77t8PZ2XC7Fanjy3b+N44fEe24W1dElI98TGOXs1z16cE/DvUP6ix8aZjRtPTkbSkrEFKG083
zZ37SPLog3mzPuW5JytVBfyNkr9CRm4Pq0oANQuEDZ5frgSwt3P/5eP8+7gQ8Qplchs3soqS5cVh
LT443F1xtbh/VOFFu3/VE28ArSf3QsW5z2U+QIfgLz4SoZDHvMAjibzbm55148lvNeV/8ZPxSK4p
fQ9OqjR7sufrvHlNiBNgvrx3qYl/K0bRFVfmdEIEvEfyvhxcLy8ypAYV9QFxwfgRu4AKKf5to/+E
ls3Vlyil2Mn6XVb9NKTR79ZC40ZBrmcO8SUdj74sOOILcOGupO0CU+WOLT+2Qq+xKeJ3va4ImAG1
nqa2aExOOn1zor59tbQyuflGLZphCtm8xM0LUxbtIyUzFMj70mfPpwEwMRzzprR5qNw6ythQ+XVG
jS93itUAAz/3ahQcpd6Y7xDLrqLP9G1pri/PfnPzhFqvgSTOG0X0uJF44ZoR0KwP06iCN90K4C4h
B7a2MvWqCTEeiNFvNNhxn3Z5S1W1bqpH/T3KaFW5KJpBOpylFLmSfVZ9DdctMKUusPyYmUwaEAc4
uzqhDnEuqquLLKfe0+hsHRqNkRsl1clNQaouLFXsDUerpEvYFcHM+IWqBxJvCuxK8omcuaUZBtaZ
0+fvtPfgFEDB7W8wFRKk+eay1ZSaqHthQYru0wFQPG3ZUt9ugTGs335sxQqml+1IXIFZ9VYo1yIN
XoteuUK8bZYQpRYxeygEp7V6sRkeuiaTr3x4ljQw9nnvNdtVDSnq3arp41hMqGkn822XDaLTyKFx
Ps4Gg85SvNq0lDRAvKVEZZsxFAEv1yUg+VOxgw1XKbjo4DEm2sLctpMp67XAn3siwubySvNEoK/k
jnYdYAkN1ZhNsDyjfVwKGby613aRBMXOhoCQXqFEKicL7Jt/38cfuAkSf1UaeLC+NRlzZ8PNSR6c
jBwZJGwaM35pHDrdphVPMiMNlw8QZEXljPt+Mpn0c6ItZOCrzQZB4rQWKR6vqjJlsYrYJSAlg54n
9FRStVLSqfeerXmduYi9v+PKGM+GqvSHDJkNmj5SE0flUCSBksx1gjJqefVWXxDx+ZLDB+0ubyAm
4wWgMz4W1mzpOAnJAx8SnIl0NLQNrSkqq6twgu+unVsVmUyoPpVTzUVnOX8BxNDUlpQiGlvdYDtV
bUZpwwWCDJml3Gkv1ggv9wi76bUTGB9pPyYg0C4k3JBFMXvHT1aWvkP2uBrLnmQ7X3p8v7Pxwcwc
Z6bkhjYRS/g5tLSwro9iAfoambPw+f6Vupf0+1gbkXtGfWeaUmC54zOuBX4epQZlpJQsrbPc6Rhu
5cjFVA80z3Uve5WB7bPTzGQqQqrorDq8is5Z2BYyEsTYr4LI+Dq/0ey6v7EkMcAlfoIQoEBxXj1y
HSVKHk+Pqe9jhy7p3grZg0QOpxv9f+vXvFWDo1t+EQmXd5kjci8os/+lN70gTkrm3bkG4WN+dkg8
WbCEqCE9rw40X4Pau9T0ctz7BKnK0VLiXTSGkedXmnHEbKprb2/N95yz21jHN6JJ0JoYO2WE7pR3
V3Ny1ivxSzayWqAN1b9Dnh1rPPXlrNeJ0V6qxOpKU0klu7bd1t3vQRsB1N/0n8CzZeyRvolD5GT3
FxbhWySsLssux0+8CQazBL02UQOpcxzjeIwoToJlBPrSnfMTO6S93oVX+a1RoeBjEbhl0R1xAMOD
q3YrlSjlRUe7AN5uHz8MoRq2SkIPmQ12o/IQxWWcpgubi/jO5izThVKuLnez7LnOCdP37oTcTMSG
xCdNVQu8pTXZ3iMgQ6Uv9kNsbsiEhVZcDMFNVf34LMRGjy+RM4XbNj028e4WmdjFpFdG8+dNSelP
EZcxNYERRQ855zm6zB0g3HbfZBRtvRKi9cDUI/04DiJD7u8vpy33CBjpFziMPPa8PRkBp9zyypOl
Axm8PGukyuvuV1DUt56vnPte/GZeP9jvbQsu5/1Cs9eYuLMPqeuRad1N+V3H/KKFBy90MWfU5+U9
Q1zgXd+Zx0pMG/j/UJAO9P8fCwuGhNzJ+cwvZIqI4vuVXKGA762oTQpzFbpO9/ueq+txPA1twC04
BTI/rvsl5AenqXWbVLxK7G0oKDT1q5mAhgaBL22eaungoQB6GXAfIt6paOjGnfXgVOP2YLUVJlaN
LKNPVQJ33PMEio+TOa0KTt7S9dWPXbwPL5JXTy9jdFpP4qTqmdA13xFyjHkCNZl0DxLXaRvCGMp0
TucYrNArerR0R3E2zJV/bXoTMkujQKz9ziqqGYwDceRM6DUAEHz2nQZ5mErgjUYFpANOreMkYBEd
fByGSQF72+c65BGBjbOT5O/cdYMGtEPSlgaf5j9ptJCwFsYH+LFDsvTbyvFST3GKVcCG8XX1qCq3
44pCxNkbIScnUMwcO+vWFwxDwJb6aPREsWcUqthgsUkoY3he9msqfCyQMvVM8mieabC6OYeZP8gn
7mTTD0O4DDgr5Zuj98AvHIYnrZvo8AC6mL2zoXgZZ5V416RL4q0OL5mHw/XUAnZ4Rb/3vgcLH4hH
AjSMed0C4mlAu9KEXKwNcWysW+JodehcVP1HCCgVGlLFsxA8fonAI1BVOuUAy4i6lDQ4FUHZ6QVv
2/aGmI9ZqLy49ZqbZyYOOBk2zG90KCg4Ry25FsWpwJ0Ly/iIRgTD4F9UIwQotaAKcPUM0ulJCWCM
nzZnM5JXMON1MG7v2aoKBX68EA+zRnkjo7hdog9Gu6//oNJLMaQcSxWP94cvcPEWtp47co52MwCW
ZIqScQ7a42fzF5feQZxR9NuqC74U2DA/NGBu5Ko1lLzjIzDRL7ZXbEnsA+vWMs/G5eefZnG+YlEx
H67She08cY8dkRkj+J0S7oe6a7GWOTmofO/h7Hubnzg/tWD5+Jg0cDMmypV4Z+DG1btDg5z36G5U
7eCPvdKtCl+aY0HDPISuEC2xxQoCC0Dy2tvKnBHzDolvBaNLvQXd5/z7OQI4uNYMTXC7ndbLoBXD
n8geo9XdtV0Lxu62T36Hhu6BtAl7Zh+qKGY5fz11yhyoeWKPumPUgb7ugBnY99yXuO8jqu/NLlsC
dfqnWerzD+JqzDd6XGOMmJYCLwyl/7Hqdja/3LNPxR1j6bbHuQgzXOCzqiKpb/nfW/PSBvzTAbCT
9yxE+RygCC4J9xny12pY035Z2pMsGbf2+WkWK7OdlL1bk2HXCtW3ycUcqvLUZn330GkQ40tYQWTU
nltTYmsA4YA/RGQxPEp0RfM1rbktqEPcrn0Uz/uWXgL4dvqVRsmpFuuQvYqyxkn+UTJgrVOBHAJn
peHtFwDpqUBAX6Xg0molKKEy+UUApEamo8a+VR4bg9NwzdFbecEUF6a9RRmhzPWsyA2mpbwazRoy
i7o74TPit2dG33F2ssD0Pwg+KJ3muCXdDe0SpBv+f0oIrQyXLdtEVMAiCgVwF9v54tjQdBba85uc
3qLtc5EgLY3nGq0cKV/JOVuLnW3JyVWFdccDTTJcKnurUS38obvOchWaEofxuSl08WO0kIMxTy8L
KA5UoMLxo0x1qu2v4wxuwKQRWgHA+W5SwTlrZftwjL2nN/M9F9AFCc02rqKjoQcdbCl09S2+WP0Z
KugnhZpenmGon5fMzAhqCtkLLCbqJ6IpZlTIuG5M+Mnsgya9iYF+BGyJCyWRAAxNAkli70i8R9ef
gKUjLDL0IWQmwkm1txMdTCKf+0aLGvBb23DlWdujM3yQpKGQFzwk1XkxNP3HIcuWB73QYOhVNpTb
811hW/p+kYpt0dbSO+pw7DF1tMMd0F/Oq9yJv7313v29aAg0Xe0J5M2tlosue6KcjGGhWjUAjeiZ
ERr+ZFVI4ctkP6+cQEwu+vDSHWZJjYGJQt35ky5D3TMs1hgGGzGAMQrLSHSTSQhXG6e1cet8qpRa
Ockv6iXD8HHJ8E0yczZ18D5/kqx0R/X2DZfp0VEtw/5BsZ3XPMpxLpo7bnTgCHVu4JbpcIVycXFe
WplA9Uoa1IOsdtEXqW/yB6syTc5rMoe7uqwsTwV6xnFnQSm77moAw74gFiHm4H0HzyZWBaO35UpU
4h18xEWSKzpQb0XDb4ZxCG3F8kW4/ADa2wt09aCcdCoOWxGrqQ/E/d4JeeWOexhqT3uM9iIS73KL
w7mczQq+H6G66yomTj/WK4cLqAuZ02szvH5qj5Saj8KDaUL6fHB2QztKb8xVfPJnCljvKUmqYepO
u01iGOUxKUm8exKKnGpjSoU18CHPe0lMVL4zux4SfDnmlKciOMtGMAa+UhRmGAeS2tnjP6HRUe8l
FIGB+tgcbOZUREBwY84tgji10Ju7Ribkdp9+9quF+fxhvv0m/3m1lmvUW+mUDu11jVb2WrweTzGL
PDTQdqw2T5Uha/CaYUsb/fYmsW6AHUX/HSvzGIIjCPpg36FPVULb9cYD53DEk7IBiesbrNaIYPRs
Y2tNZchFJM4kFfGIuGP2dT0Y9u/QcAXSaQT7CyS0XC/MuFym76E/zcCdVeZobqdXLW5Ohi1RG/Ee
X+mVNMnuau4fUsxLaRWU9Zb/rZRNjEPBv6aRUofdmuXzUIVEMwL4/OgEXRy5p+kxvQvWCV1vcIDO
DL5O1OV40dl1A5l3CXWoBBIfdAftGr7uSwA3avIfzVBvOe8fA8vV0zcoMRjzuBm9Ksv9f5c7HYq/
83PyKgaP/nhWZ9HIqCo+m+3SrzvbofVcEDKx0O/UlFV48MeZsppYlrQYcvOQjEJ4jj4XAru9/vVH
+yP89rqtL61llNjMicahtdxwdV8IAfdG6dd9M+MzfwmlUxwndnrXIulZ0DKWOHvJ/n2I26iyZchf
XtywqbXUDf3k0DbpeSXcQWJyZANoAvXZWASfbdATiF0LDILtASNNokqKwlzby8kbd4Ma5fRaGHLo
vnx0EtzCgL4JrfTS+ikR56Q3sUguPZWuwjl1vfkFZ/BdSgWx5f2Fz4BKE4XMKTiG3rW1C2gszNoQ
vhTuUg97Y3gKnZqNqH6QmGh0NEcDazoAQgKa1gv58lpD4PIDb48Ra65LzMPGYn0Bx6hZ24KzLjOL
+/tKI//GgkAY5vRmBalUNXsagVZx8HWdySTa+01dU7EX6/8ZwjY2/AWARDReoXB5YWoWTUYFMywz
MlQzHW4cwPgf0ZsNcaxyP6Ka6NTwraeVBrBbt/z83sykM7WlzHkmR2r9G/6V0SR9pzzCLLHVCVo0
NGQBSIwaqdhkMitCwAhM0/FcVPT1ePme70CsqY7QPbtez39ycKsKbgH/90WCqOzb6SM30v/dV3Bh
S/Hot83m7oD8gspHpvtyB4QmAw3mfWK9LSI8AV9kUVB6ALTtvOLSZtmCKLSGs+bfPDwgI1DL/d8s
UUxViToKhibORSa+WCi2Mq2WnGt1lv5l597cT939T6dDrs7TaOPmDfQ2uG9PQX7uElbxueLleGrU
yIFKELgpel8KePkyUq3cdhNBbae11zmWBocav7NOKzbv9JmDnQwvyrXupL/cVAc1MWItzHd3Fmbk
NyDInVXHYsnExTnnslIWqiEtmdpLBhNrx4HRuYx2Fyr/pLhTCYwgPSv6YaPrN90uHH5zHUSlwlzu
BML9QTg66TGNGE6sTwUobXAPByFoHgRl83UX73Ux5stR0kDY3sC/vP5uxQk4fGYL38bkM7jnAAV1
oTiDRHVV5O531sL2GJbKHHlobjJOg6NVeUOUhbtkT64h6O/tTjxv+hePQMJNLGZT9S7JzXOyj8TZ
P+Dwprb39hcHTIwgJ5/DJATev8XjvOQaAU8yxGNARvLdmfRsOIYqk1Ka/el5NhuV0+EFYhaNqpoR
aUG5+jjOqP4OqW4meMjdQzV15pxBiuDNtT6wxR4EZK6JuZJvmg3JCloBfD48yaovXiB8/+CyJDz0
RJG93Ya2ZjzB7sTpaEPQs8yW1dipD9N6pmMNuDYr6+KssQLvecoh4YuVEHN2bPa4rxULRck91LCU
5g3mLIabV5BcTdBjgWQhZY9sY7O5XR6Zg4j0temOqOQAMWUDvhigT2RFpYZfnPNPz3UA21LrQ7Z0
H6zSY7dPGZH4po+3gwE+Ywx+nbEo5CEqxRO4rIbzkC5TPwla6K6TTrnQKu8AR07enVSsjLghIQK6
MVi9CwHTkl23mZ9QfP1n8MVKpq2KFPbglPjw/W9lEShAtpg1tBACQFoBXBq0q/D1Ibez34sM9/Q6
GQckL2n87lAzUh/cQtYIlDhaz/FnCFa6A6bnV5VKFsjQaj93yM8oXHmgN7NDBkKVXvNHBgbH+5gg
DV5dV1i8ABrpui4wEEMvSyPorVOu6deCnFSOQRe1fFZTkSMKPZF6LTMq0uqtXfYMJHQlyW+AEtW9
DKDF1lOz4xDRLnUoNYZR6V05XNbHlvSs0+4T3TAGg4hYgjFHyY+g37w0ap/9bNDaSfDTwH9NKrBR
BFozJYD06ngLwgk6nLsZaA7pKeRAg5vIfjEMDbAp8kkORTKVSdX6bNGLohAAuVNBZHkJAWlCUiyG
CEVm7wziji+iV1cnWuRgWLppGCDxzWITcQz5oF6TKoGLRI995diEU8ceKcR10/C7CXFgTW4HVeYA
H+jFllXRnarbF+vKF6vZkMcE/JrF8p++VLey5L6Ydh/ik7RkQueYIsizIVE0MmtwcVnx1U4tESjf
qWcAxm/xFKrD+JodVYAR1NaotEfxTI7qCdtW9jbv+KzCW/m+JhNLymtGHXTQh1gHp15bRPa+7DQz
NCkeIplHpvs5/m1LTFGczzvGBIHyCc99muxdBM4oTb4qtELlr7FW3MqbNdSI1f2bSTF3a7cLV+/Q
6tVy3HuDMrqaXPR3vgNPYRqhHQ89N2RsOEcu3nk/btY3T2HhMYkhGzgvKvve5FOrIIQAV1ojfvOe
TyfbzssrVMQXoSQaOIQc4TiZAmdmyW9+I7UfckzfMkfdORiI8siS5NGvRTN6cfm9E/O9ztWVODHU
EsdBl2zfOX7gRgOyt3iNd+Q/oYr/vDP9JEtZD7KzdGAuhwcpT+L/lntpiYOT9GVN0TjkIn7x/BNK
loPxN7Qb9f44rUbTy3gwLv9vb4Op/yURukJpiwXPtjfBRopiGZqY5bpzp5uf+T/jQ56H5NgW4FeN
Jg6yg6fiHczTDyTmMABwlDl0nGWVSG6+5Xw+/AxxH8B+0prnzXi/A209VgoxvleaKiXFs6VJuOmP
vPvtUoMkHMS3lMvK10hdEn2FlNzmBqv/Vb2sBo9vBEjx9BTuNOWWfaAMoXvoJO/SDdI5rxESGZ/M
0q5kMivNjoyqSydt5e/+GnWV7B5B+e1scF/d7iQLd3rXdBf7gAvCH1MnqgeMRNUdCDnuMjEs4wsP
sm9V9tXIzksDIOn1+H8C6XU+9vO16AqdkNGZ/wzRJjE7r2F8xLYcX1dDWL3yUaXWMmo8VXi9qKCp
QjvKu25PESP17h7xt+tipaLb100sZv4NK4px1X9dfxx8wG4Gpi3j4tAqkauXB6m3t+g+3FP7+2Yr
B45FVJGPI0/wtjb36pGsGDBZ7E1qozv+d++Kb6l1H34kswYcmCNhgeowgAoLyRTvm3X6bLPbPAye
WN1jPakzUkzSbZxu0bXcswsljyxY82y8Xwjuzq18ocybWOFRNyMmtBT/tDO5IuWp980S/p5K8fB7
3AVAhSLNTPr7Otth2WDbEHjt+vOnPMbfo3U926SI0HXra7L0rExHwRgGsdsHtN5Yq/kbda8nRdbc
WPNFNjVHA2oFtZGnJCJgQkaU9J0m7SJYjJD3oA56ELE1N2yujLCyD3hwATw/SSmo72NGBSM0YTVu
00/epMo5MyWTQEvdrw2Uyn+BOFpuERPxlNhqWKedSWw7Zv3HhUIBTEhsqSBvDA/vQfwe9xgLrhF4
DtbNQq/SWtRNtlqu1eXi8C0118kBxt0NfDCYi+9sPXwRlpvewQ61vu0W/XF6hGSJH/oA5kHEC8qA
55Z72foRr4PJhmcimjNpArkQu+nP597q+Y1rYv1NQRwTLnyj6kECBbFhuA5DJbd9lPOC0ydNZEdQ
Bzm8CPRAVR7rSBi66Pmk2KquKhSiCTVT6mr+rEzjKb69Hqh1eWAs6UArbxAIokhUKsura5Encxf2
/ISZvdyS3sZkqirwErn6TKj7g5cKjAv3dcs9vOb9VK0jd9M8PE4Ppkc+f2fAdFJhJ7OBQmBuoZyZ
UbIPHvYtIpNon7RjZV4ULLOr4JbDhRcHB2KOXaXQ6yRcd6GkLDRLXgXimekRrUzdgPDLraYhUnvB
c4xvEHW1FKWxjIfYNA/qE68GrXlu+u2KUiLbIATn7ek1SBTq+Ipferkh6CQT4+csb59LAEqGo7K3
4/eq5rigDHdvPUQzAq0rhChOsbj9MeYLRzoKIypEd4TWfi+xJI8yZ0Rq/MjFV2s2q7pW25MSu0bj
zRUmWjQRTgKF2OavmSgImyK2kqvzF3X97WvasBaSYLOum71GTALpp9aIhUd2WcymeP+vzjqCJ7mD
KZnen9Lb75J8VNKTISd07NY0OPhqh+fx6Y83XO1wOPvtUFH+ZPNU5s1Q2glnAUqlLUvM7Y7M3SYt
YvH95Zq+iKTgVzk9PBME+dSIuNQHfSjuPb1ST4IynLffLEYrmR/I5pq72bGPqtN2KAprbM5CQLq4
Z6OREVQNSXyKGce/tU5WDxnQYaoQsNeL8xIRW/ow+BzgS0+TccrTjT8xemFly/jEpr6JFBfRuaPV
u/fHXzyJzf0x7QhxV9euaKbnLlDU5S3RR5YSNDrMfR7K7G7t9ZPjow8tjWan0UaX4QGN4iAAr8zi
c0/KhVJ9lIICcNfx+ZhgyHeXLpsKVc29WAt5NBhTmkiC0WvQj6742UFJlljS/KFy/bJXKQTMEhe1
/N8zYdj4Pq716BCLhn7NcLrNRtkGadh8QYq8Espb7HtoRhoacmdxZZ2NCY69dEe16+BXuu4k4ijI
9nfDM4WGCG+PXvj+Q/t0XWEon4IbmAg4sKFVoZGqXP0+CYTUOgfvxz/UWNFbyLlEM6KG4TVwD2Ov
P4Bka2sC7LHFF9F9c8IifsmJSB/WJQm51ltekgEemEJAV2nwcLrjLhaH5/CEj4PO98tgFqnWh4GZ
KjZtRus1J+qPHVCN3n6v0H2zwgR7MDWDAxIU0IWFCyFdKDXEKmsWcWplmPY5OpHROlsxaLnuquRH
+UhFjW2nkoacbsLBA5WAbK3BlqjuLNfWwNH/vZxluQgpc7vwe7AdB5frWApi5hqvEMDDEY3AEZrD
ATLSVXEVryULVMprQarrYeFQbgF0M1F8fLLaVaPMk+FCiHvUA/Gn0FOOBg4tbkU2HZwnF5clnzWV
wCosFONHutui66wjFEsygwGm+hY/6bUBEtEshoqliWUpSOqheHeQSWBMjATXyx5zFhVDxqkS2hRp
jV5uUFdb63W/RGuuCfHa9pMSBhyHUNjMUwLJk29Ajf1A0P5ptLmhI0fE0czy1yPDRfWBW5jgVxwj
t0XxBd0lgQEJhm3pqY2IOhCW3qHl9r8oJeEL0tOA7HWT7vA7erJaUxRZkjLp4fdZP6IB/QU7Ojk8
bVO1iPAzog2yG43OXBuSUabwl1NEWExi//t2PMUUajGs/CXnx/9xrAHpjHvsX3Sx9zl5NQElPJWK
CsXEv5BWD1mJWWssTA1nxHJZMg3xPmTY15piZzFuIzqtVCVBW0ajytGPdTZnCv45D4aIikkUy9wq
OiJ0R0EvteX8Wb1Djq38t8oJuCWjiW7lwUu9lZbLcg8ehk9/IUcn/lvZqEuIka9vVzQaYS60zZzn
BbmyQRqovShMtpitRUgsWF1ysFiuGlQ60o3flPmGUaNgaHOyeHxkf0PWvwgKdlQjul6YYkxuZ2Yc
mzNPrF2s7sR6ZmP9PRTKkTbTjGMR5V+zFjRnouD6+CuW/mZg5PKm1XXyy2tDGbXl/RoynJo1kNOE
Hji5K5EVCKVFE2F330bJC5X7GV2i+X2m8iyDmdcP/63wWA4mASO2ZIUV5WHzh9tCt9KN8aR13sKT
M7P7UiPdJtAfxIP6EaG973MKAJ0FCmEicZFQ65YRYh6LfIMzMbXaSD6kh8Q4FXOSbg5lwcHdygYw
Aj4u34sR+eeo7tsecfkoMgU95HSpANzVqEfRxpqFCuFHmZj0n3UuQpZlQpDfGRcVpYl3xNByxDCs
GMKdNIoYMdcIx2S8LNjW0Fm7oxVDATMogt6ublqh5RapqrEX3Rnb132esSvn8b2HC3L54UbGPupr
iVNEDMkRnKz1AyMY+myI00VOIQauJkzPHpJ43DhlQc3EdCgKCOYHmE6UtjlqmPBak+aJcW7gkQ3D
R18AGEpCiUsU7d1gqdfrJFDH+n0BnL2GT9U4YGY8NhFdMu1Qxb4EqqToMy3C9Ccwn2x/EUcGpTHE
iNv6l1OzRUJwF/zQ6yCvchSLHymH+fUjheza2fgLYbaA0mtNgXaCMSm74c2gOTXukAeRDU5HrJ/D
ACfeokrpu/zCdk+8+Tztfw0fD/8O0LCXWU1eDTR0SLAJ0bY2gKC7C7A8qRkD+9nwRQvWsrzUnniJ
X7/dfZQDu12TyTAkmh686b+pIOWildGgaJ56kdZhhFtm+KDbIViVSKuLlSqLbnhr3NNl4NuFOyZY
2C56FDTsa9ePlzSoXwAFBgVV0oTC+NPlX7SFR0FAw+K02CfjKPjSiessWkHd2bvG+oWElHAM3BJy
YN2PltnkfM772MmP3l3eVe9uPLkgHMdZALiGNEnWg9ChtGkiRp7ShfE5XnEIy59Mn7V5ISJjEDq/
J8xVNM6JymdSQFWsDdvyPXrcGQSj8SJp1iW88BORj8TVj8xcDPBLTwV9Wk96pBItTBULEzdEbVg5
MlkSV2b2bQTD6kbSd0AxGlLWa+92z+GhOO4tovsolMFa5e6fsk9iky76KaG5U9SgzX9B8WMRhL/7
DBEopyk27UoqomUJFOr3wK/nM9J2aVOnNh85AedGB7ZhK1lw/d6Gd53fPhNjjQNO76/qFKZ4omRK
CMhG1Ov59Ev+hr3OnxxdMRm/wT3p/wMopD86UwECo4mOGvkphzQUN2mIy5lHMDuMqqO7b2Q/vn2F
W7TDd5qdrDj9LRw06uUth9SPcWR9ot2efus8ffgqaZI3J9HRTpQFJ3RJJkdioom8+DYEdeYEmzky
jwZOFMlxpOoZ4cJGNSdNNc+2Wugno2RW71do4SSEygBPyz7cB6bFmz5vSKJRZI/umjdD2zq3sVSd
W62XiGTFIjM8xOzzeXsqmT+jnkgkQIZpiAToF0IUtG9so1C+9OOzpqrjLsuredw/2avzB2fjvpul
BEvX703Rxv3vwchD09HcuLGY5c2BgxFE2kKl8kd33vrfURkIQa/ndn4BQ+wwTz6vvpWdg5XCjXHI
yKwypVozfKVX+nFvbvq+By6RC+V2I4TvsggGfqp6WqpVfOuF3ZF09Lj4fhcP9q08qqwzG5AUpJHE
B2HxblACE8Jje39awjFXU5c8404aPU89rDDW18tVcZgxnzEF5MDwlpFvyL0e1NaF2d/EcMP3AhS0
MC7t+cyWmMHP1L4IIkvmxNPBGi5kFnIn6s1XBxrOK8PXIso0e8BQcX1tx3Dvr8Xv79tty/d+MsFX
SreNe0hcklsShOh8/ICgTGu4VZ1SnsNaqOmhGVCJM2ETmf2I7p4afWyOYkUfeb0S4KsDIxuSUaep
XdDxVE9OdsPb94N4ZIHFmBjr4OCc1tQ+j1A3NSKBqK4dQLrccahx8f21plEa9dj3xelFFqt2NAFU
o3eYN63s+OlmGBT5kEy5afCKrS9yh3J4+h6JwqS5t3MuHYBPl9a6DbJyrl0k3lGNOFN911ocNAZE
WJtFC/VvAHwDWQ/TxTVVqA1QUQp6ObeGyPt9EKNcgaAqnbDsdnFYwiScwLBNzxja1FcqQbJEjp7P
LCMBdiyA4HnuDd0LU20jXe2aGtcy0r5SKelWC2jhy6F53IDW9JFQQf/+dBPKfBxp4nBPb4sVzqg9
lzy/T6utknFwUVqz45IJlrDlHjY1iDXnvC6MoPjf87ooZro6LPW0XsOD7lja+SynCF/3OW07V/CE
8mcInfDiH+PBcAQed8U8/G9Kd5NwMm8TnKCw6GOR24GPnS4wXnCXwqDFjCGsGY1E8OtcuLeL8ncH
awF5yTAci5+4tmudVLet6SqPAnSU+iQQwLyH01d6dHd/iEx4HII39cY9v3piRKEUceuTlfwtV/3C
kJytjD8mWnfzxdRPvAXwZgSRs5kAGok8vQm8Qcg6mAlfPkIFDc5vObdFeCicCaQXCI9j1qkTmnhQ
eVxF0w3WCfhTZOKffQxqYnknmqyCS7s/gFS5Dh1SaHpZXzUxzVeO+oYYUTwjdMlk/98+u4ikqvAG
pYAjGpOMQSQm7VFonfnw6lL/4ddmQ1zeocIryjiYeeT5voLOMY83Q9L9FUWkZ69PM6Qa6GJAQI9/
xwAQeIYsngfcpOElwr9IeCu+YcAC9ZfBbyLy98YghPB1fjg7OzPAZVmaGwzmD1TQiBu81cPVN/Ti
Jf47rnl3Hfj+ukpXL1itjMCq7M361baZor9AHoYf1hwxteQY9oilCxT8SVRN1jdNfjaiGRl2qX18
ONtPod6b5AuUPnNRzka7ycn1LEyCPfnBtdAVlzMyeel6Btpzt1W8V0IZfo+at+/FAeEvqMapz24V
6mg4iAWia6Hq98ZCcQzglbbkj2X2Ad11BcpkOknZdsb9mHh8iydFcnRBlnREO+U1zt8iWew+A12b
zQ5GOBOvO+jKWzDTHNCT05tficYMyreW3+IrufWoD85A2XqkE6IosgBGmegyztndpitwgB0SjABP
FJ7AWPliD6ro/9m+5zGv2xh2I5JMgV5fWicsHGjY2osof1rjR059lAnt/mWrpJzkZ8oBuzh/6ia8
twWIJIuhs8hCD0e61wWHo47kX0pywq6u7zMFwL7APwnnpj+WTA6dO0/2M3sUIJk6xf3hO/2wZEBw
glHyIEnR9N7GUkRNtLS6RZi2fh2jmBAFkUobEIH4d8A7CPPj/kItgSjfzLOjwbKcbZJyjyicapcx
y6wV3NKbd/hwVwI9K9pmcfe9SSG1KLwPxOSg01KnQBSKz+V796+QriFNHAy2cLA4FREZkWVN1YvN
ETGVCgCMU6Z9RDFutrjh4YFmzlAmwSEvDL8JqUh+BuYu7btqKUq2Z+3T5PfbzjDIb4NJYv5yZEGT
XjuJtbk4g/z9Hi8GwAqvkX/cthEQqM8RwwsuTDZ7lSv1lQH3/hMOLXyGY2zJJc2q7y4OZde2QXOJ
SiW71tRadpKAVrs4JcEtNBqZDXqCMD2fkgvhFD4+4p9cidjuQzQyYb5UY1/7JzhVsoLIKfDLxRAI
qLwt/wiqSPuxXkFHHa1Vu2VWNNAOQzi1Z5PElaAgjTqyS9FqMPoFBxD8y8FKDuRfK6TN3qDHt18e
X/ilyJxZOA326am73wBcdXNaP0JOrG2r4sopN6rhpC6NWYSE2YgzkuQb/YDvBfF5D1ECAOf5bgrO
NShNkei3levCwB/b4ipyqEQCUKCO1u1v3asQTYblZ8FA/VhTqcR1I5HxmIpLM39kUzG0nVhwavFZ
v/Vqkp27GTtKmEa5F2FhNmfObDBVkY3u3XRdLxt5LY36I24R/SJbrBew5+Q4tDlRG+sKvvQ61Udo
8B+RpazclhHTMdDrRt23FSbPQZ0recyYl55WTaZsNh5sSXr9z6zaPF2hE0fUhF5OVtp9gvhylYgY
RObXSNZdEHObzcc7uAEJQNnsEgv1Pj37MiTZIry8vHUWiC/4IW1ssecMlon/ym2XvdIRWsxPO273
KG+Mm50MCoX4COZg4uqOm/wvOK9wW+2AszQqGgxpDRsLFzE87Urtzc2IeOmx0WnPYXwuTu366ls2
oljg+5L8fNwbJJmpZWSxIhXB05iX0QVVzNzP6ISqi2k/OQCTgHfG8Wk+aQo+RuC7xSw84+RHHc62
p0ygDoHd6/AS6mhJW3Z6Q+aMlXNOqG+GuREH8B/WmaPRv8aEyoJZZDcSXDut/3XixFl6+fFaPk8D
it+hiChx0NLeSZjISyu2ZdBzVEt37JTp9Mo0WYYR0GnsCuypNMBUV+kEb5Ygj3ta46s5TjXtCX09
fHGAqx3S6cnW1yar6kfX4WhhP3wDeQRau6t2V/K/r/WuxebW7FvF9vsdp76YbkDVuGhOekq9Yo3w
U2ySANBRCqe2TD+gv0ObMY3nCx96VS+m9Dz1kLAKYtSRxMKPIPiZvNp2ZskE7q2nYqS+B7EFkUfm
0ZGFvxesAb+Dsl45alFl4loOkON41lYyREWY4aY5bjtPOM8kLI4B27prsE9xYXLAORwkco/lXaIj
xOW7yZpVsc7NFZbQKw+puuBEO18V1piW9YiGugmek28oRIb7Vwr7V2TQlluHKBQHFzRXKk276rx1
EEtb0rDk6dOIHO5AoNDus64TJxSl7RdBsz+ZwwzTyRd/Rmmat3HjqgwUwlMS93CQ443xe4B3Iien
A4CdA42l98//WXYXB+Sp34ioWWSwhiF09SmSLHRd4oY8PsJhp15XNw49sjZFn4Kcbhv+Cm8DfCB8
tjTrMpxJahi7D3XwG5PEciLUqIGwNB4LNe7Q/TJTyVx+IaXeBGbk3p8HfRpbq9A0YHZmLBhXW6fg
NKvxzQjOoumXIve+TaRbJtqSakGM01zr13HIjVyukYPMJNwjD4ELUV7nRGHuVyhm7UWbSn0iH4bW
V73OMg5Bcr34Lye83kaBFANhAfX/E1nWSsf1Z3YmX4w4d4a4H8C+fYvvkc7wvradAWcrfHvxZ8kl
FWTVHxvQzKgodwsAkgkXXV37qVWR0KYOlalIaX0McbSDGbhvvXAcIuHYyVWwJeCyc2a7O1fkl6C9
LC3KUBJyEKKSOXj6SyKD1VrT+H1nB+OytPEyCPfmi+/x/rVHcnt/vFtH9LYUqZ0ljN+YP5DuOv/O
wfQn32DtH6Gku6vgmFxaHXSoUE1Obk53tLpa2KXIcHmmeMs48qDFifRU5ZmWcTodFMwB9kwksPo2
SBXsvsZ66ig/b/1aXHuAhNSC5kMxW36fBPaT53K7zyZ8qHjSZHZeNMHdBr1X+8KO+yDQD5YyV6+Z
YzIziWL0RqwiVxHg95uJtNSk7hh40skDWZvfLFWfeRRMRdZSYhjqYP20pzOo8fz3bHrZA1i/F6iS
0qb+z7z15bLufwk5Xy1FDAt/q6SUYhqxHL86zXh9yvT3Xb8YIgBZQwvIz5bZkp8jWwvnc5SsaSaH
vYS7bBcSSJ+x9oE12LDaY6GM9LNdvaF8oyF7IkxPz2o/K8DdnmuFCxGhO21ckGM1WMG25sIivZL6
wwflV8oFDPaZkJX0pG/Tdtx72h+YyDt0bTHinf4nI/gnSXEQJZpmvf+/6UA1PifUSOfQfPtHZqkv
i/GvD7wyoBfWelK9IlVYDYvZXbHfAx+SsuSL2eeSSu6/0y4bhRf2h9CMdmVvQjicBtVfk/xSb9qB
mXA3aNN/h5fP+FEN1eJFkBvU9SKDbIbmbTi7pYpOpq3+xTArcuyYJSKLX1IJv298ROFL9IYciCME
0prMIgdXQdDEla2cTdOidkm9USwdyLXUus7Ny92U8zNE45kRDA3wpa7+hbxx42btE4z50kAUYnLk
WcX9yuKN1AQtWdqdB3RBS9wexnrBeDNJoxStts9iUV/Szk8wFh7ybJm349VVEjhU2GKqYpDn6gaG
IIjGhZLouxBZebzNLUuStOLbQHWbPExV3h28yPfCy/CS/OtNI1j4cKjII9zfSl01kO0rnKhq78sh
2eCcMEf6q2FPJ/C+leUyV6X2ja9eZe9NtTDDOcbOSiuzOJiZhiyZkF+A5KTlkTTubcOLw3ZujRob
AH+lNoldemSBFDOvhTKVz+qxNw6Ju/UzakaRxfEh74+MlLrlXrylYKSFBgzAYYyogX7syBkIG0eN
+JqISpfd/uSBqKebVI21Md2bX0+/6cFQIvDPk5XOwp3P7wsqmY54hDvaVOcgrY29I8inmqwCK3Ix
pODOqQjnzDsl3gyzK7sy9Fuyzu51PbdH/T9rP+vBnkKjaQD5wqUobR8sft8IhifYBn3hc3PO7DT9
UGTYe6Q68733gnD4HPbKhHLQcWs4wTWiTF50pBGukt5eecy52DK/W0WCB/axkn1SgRxRPbzYrY31
D4a8WbBw7qRDgGh0ODAL7+aKjo48vjyMTbFEMWFQI+a7OsgdX6Gy0ra4DcaJbZI5rp+SwrvmEDf8
lP3DIV5SKlImzusIFxVqU40OeIZhlG1ocFYCfsHp4dO4P4xAxK6mdvMFer/Vw16Hk449ZlEuoY3N
5d7vvdvXgENLh6melYx76VtB6mY40fB9Va2IFtPFkTgLcsVqiKZUQaiQeeSidnGArNqBok+v3LPz
hdszZ2wshNeHbz7GoMYIdLl6+d93Q2hcmiqDMw+1xckyVv86ydPGaYYGH1tYsaCcqd8RqBAa24u6
+EvKNVXlLOjYB3lPskzvS2tVSeZZQUKDcqqKJDFJUHvww5rJ/y8plyNYapXCAIqPcfUn7soXybRq
/HdHPglNCUmZScGrzLEd9762Hw/F0nyoOfiIJdDQLvPS1ATY7PiGFiG2AB/Rfs2Pl0IWECFgzczW
FkK2in8+CwJbe8JHFQltpVGMgnR+bf9ApKkY6e7RO/hhGrAl9baJjXBgaTzkC9VxlXyB/4rl2oc+
LTudSc2xubjhUf0iZ1lbNAlLlW3iRUPEyxVVzXiqyZ8KMJUR6fVw864K6eAqndWoBJOsd89i2oeP
dJTi6LCUSonlIhpeLQWhv3vWOQWrPhB8OPwayHiTzVodE4XzAs/PAPiExA9Mf5Ez1LvOLVPLJIO1
Epv9vokAPk5VPY+B2qzVIytFLZ2OCgWZ+OTRxfKLSGmwf5bu40Q2RnTKgrZe1E0IItWbnjWYlzHz
oGBjka1a5I6X0DzCQsjthUlLIfqcQm21Ld/muP8Ouems1p25Gs/NYt+lW0yDs/eNX0AyUdnFClvJ
IijMkFeyqR+nKT92HeS39LidK+oa1B2LS6L1/VwoEGasai3FLrX7YKpX/hAOGAZRLb2g+lwEprkZ
gbVcITQQJUZXGnDG4NkFgsstvoTsOtSQ0lj8ivXmiG+DQdlHuodiAdRa6ph0Pm0BTDwwUUSY6HTA
qnqilTnFetc5a8UXNB+gkTqtFjmNehzhRHcbEX/tMWQGwwG1JWkE7sA9cA2Fvxmlv5cB0Tn4f7wq
FmhBxVwno3MBa6NJZlAj/OPRcaWHkjeGybP32LaWOR/JHE4GQuIihMFYEEpWTlVMDnJiWdQSPPRQ
X5AE0b6trGVoW7sjHs1jfgSsRWkXE523VFUw0Xh61w8O2kOsqJ5yo6aDn6xRYOTuDSIdWB+581bc
oLYUWz7kCqbX2bDrH4i5faGid/R0eU7F/Sn9bCru9JNV9efE2QKNOS7Q5alnCCXOzFhcp8izAk3m
wPWwWIZKXeIe5oF2bckEOEsiiK7jveoEIB1aDB38fNnkCETox8UvKW9kxTvBY+Gr+2/okNcLC6/U
Zvx7vgWFnDtiKxxO4oA+wgfVMP/1a3tEguUXGibULIrjVu38sjZvZ8KOa5mRob+hIX4ZyAsBLxTz
Qk8zQaslNSM3G6/zzbKXczR44bRqtcaO3c/d123nuu4dLxwKDNOqvpJuSq91rgZgOiqzeAGUGOA5
79o+PDFvb0iP5nRRlpTkiTH8vVHLQopAOepsfMFg+xSygz+c7OUcVUSLXHkNGV4/PjoxG4li2FET
Bx24mB1BT7uK8Ow86f/kGJr8weVtVyEsgAhlsR1mGZplmqEcVCp/dylW9cdzr48JE+1/vp9icrU7
qGdq5/BfNEB6VfVCmi9TKtb3DTaPROLP2h7NCajBBGb9n0S6aWO7HeICG84pUDUcITKvuKgcIeME
EPHeuPow6a/rJeQ/nJ+f4XFh5WCawpn3UFepMj5PsejARL/HADz8qK5IvfDecrvVnrxD/Puj+FhC
MrjSIX5FAe7Ya1ZxsiC9+qHKGBH/LHV1x4YLLPYoTL5QSotxHfaHL5F4RrRF2AEU4nHo0GjLQGsX
CsTU4S70jjCxKDqrKwwRXSkMschwSdfiIGXWSzfk+QGs7/d6mIw73Yvyaf2dvQSAaWGGAQdlDcKk
u8wgz8DOLuBOGRVMzwQoaCkcso769c9pwa3azbQIlTuHb/i+2Zkwvzspbx/MUhf8HACbkdZdxkT2
EsboXPEz7i18IipEcRgGm1VuJAWgTPefv8PxR78DPzDW6CyxOuwwhdIMki3Qxj0AkGc8eU9vXNr7
rKdVSUApPfInzCj36qFKLRjjMtLq37BTXgnuXVJErYcxao7KxAar1PZS8JlGcHwU8V9cw2wLpD6x
7RRD1fNyCynUHENZmi998r7rvVyCzqO9vvAVMFt28ZXdiRYZKDm52yyPDFHjr3X1Su8T8e2clW3+
U+YVFVkAA6VCcw8IH1nB+FCBqhA7Epmb/V+P6eTWno7mCdunQdd2/WflkRHTF7pJQEy2WiNqnI3S
rWeXCDSajhD9U9yuKF0bU4H1FQHCUrmIegUdw1jfSqRdNBCWkb9Oj215hWj9jGgNXuZAU3+jtWHC
CFWj1GmKf6rB/v4AaN62wvakoq0d9//OogAfgcKxQlorIaZKmmVNLz2EQczD09PVB5wIkek/fXlT
Q0sL2Cmm8Ply7qMEUqqyuav4hQ2DPTTw7YHC+VKAgi6uMmwL/kRyRSxx0A6idQCjIMZ3c6ZtrTPk
BBR1ptckQI7f2O7wCdWUg9+E5l49tQkJytCa74Af1ChebrUYdpdi+5n6CuGQup5FpBnoZjKmEZ5p
Dry827k7k+pvrY09kpVGi1i8N7Mfp+J6sUveJnfO9+sdZ4ycI6q0KvZCWqC26VqToKR8WamrO7jD
RVlDlz/5SLCHBEYdoKI7x1Ip/nV3X08UkkSGwyB2wlIdNmC3PwN1qjpqRvVO4CQO9YDSY3/077m8
KjcoaGeN2+9KBrMB6dql5UK5cK0wz1Kf6llGHRDSjtfUbAsMGib26HPS0JoOG35xUERGA0/QSbNe
csxtk/4M03z5G1And6BJ+PFfMrY6wtz8CIg9p5IGfZSesXmGiUzthQu+po6wi1r0vNcRqiRFSDn3
GzLr9y+1M/l0I71VIdOYvxwNj0tfYdEBaUG8yO+oAUHOlS6AwiwTAIIJlnzHO3+BnxnQZeVv7pVW
m95aiX/IsZzyKm9dIhayMnqj7GUnzqJ7l00zJy8L7iOwbyo9EriYxpczdBLZ7WfJKWBfTeF7ZSUg
3gxNe4yTc16OPX+hSuKj1B4+WxIjPGqmusneUyywepsXQz8TXhkaCDrwz3uu8wUA8PopYBIeqXYu
vf2UlKTqkVXzh/fmR9Eq5JS0YXGNExuPv4qzG8ojYwRDQZgPcmF8oMG3MQYJgyddJ32gAYpOtRh4
r4MM6HWmq/48d2OFiAG4NrzzgoldIjDCHVcSGjBUMit2WBOoIBzRk1APYuN8wpdBDE3uPb0cWmlz
3S88RowrUiXnb+MZFdZQY9lW1VDUHiVp3avLWYCi7UJrB+6mEFknkHBvSYN0xul7BxcTnnLL7msC
Kmu8kjpuPRE+l9+Eb17t/YkKRAQaR/mC6ElTZiW4fuhsz1dwlJdJ6IZxjrqjZ7zwyAqHylJD+GDk
ZBUTSDpyZRUL+8r1l8+ft3rTTjEbrd9pX8dDzduL9FDWE7IbmkcCWexbr1L/p8w0rDndKikPlqHT
O62GaAGlppayWDFgzZKpqdoiua1eT7nK3Z5WEdBDHxhxC5W7mGFftwB+cvKu8bIn1aN0scWrz3n3
pxENHF1A7yrAdJZiDmERsuK/18sJLfBwAwjgk9I0ip/zWZhNmnkVwfg1G3PC1FGwZqasUvrQPXwA
Iinl7MRIv7biv/Hm3CA5wDNdqprXnVtERWcc+43H8I7zoGvHJyaWVZ9PeEK+A4toKdrPVsyqKLSI
x2/fINW3aSAPOlQq5SbfrIyQvW/2r6WG3FVYdR/EG7evN9H6iGTT/nk9TPtUeDsoyX4pjr5kGblo
1wQGrwo1gxukHOuh/SaZ+v2EMXu2BHaTm7y+fe/6b69UgfKbnbF75g/kakhrykw+4Uaf5GfInfMR
dV0zKs2wQzwsQBhOxWIXlq/FZ9yxqZ9nAjVHlQq9w1fRCc+gKEi3F45PhEaqzyLwBFjbxZR4taXz
kR/3aFTa8gSViDbJPEDV6n3q2TTRzCZZadD7o/0arZ5lbEFVWxYKptSuudBeWDhXlbabfVKnGnJb
glIGwinZnzCTfPJleSk+CoFMJo+I0w1Fvt93wfVnOyEXxvbFk9iEoN+qK0PbrgJYdELurebFHOTv
DBJpEaZPhWvVRLvlwGf5n3eoYJX30mBtKvF1b8rsrSbWhCe1YqLRH3j3dorc0Oz7I49XsyAnB2a7
jom08jW0uYowx6uxlxslrAT19ie2mF5sAMTH8j6zpfAYymUroutGY0IugCi9OGE4xaq+IhYw5WTu
9GpRcl/EuuGNKADMk2vnPZH7rcsKfmwaMndOH4rFPL5PUEsy797FR2czGd10odWQ3GUey2j28+ds
uzocWOkZnkq6l9XL8w3qgJoXZZ5r8WTahguTe1RAD0Ub6+x3c2YITk+EPx44wL562YBjyDiEKy5l
qqnslBqovT4WwB+kHUZMDk7FOa51EoVw+qoagFI92xWv5JaQN5cQ/HzhrVCAT1s1/B6zo/PKU0dy
02LSxRQjIFB+adoPwDC9mG8Dow0cJ2/qnzBSGIbxVntdFpsqhY76k8YYUZPcrWObOACXd05Qcc3w
tU5LxVtOhTeYvESdAuCI1Nioth7vbkmdrAJyuYcDc8hPO+2fcZ/MKB2EgG/DZmrf8dqXMJxF2q4K
+gL2M6soo3yENDfpRdMgsFxye6OhkaG8b0ynKxaeQjzG5OJsMXSbWrWZTPkX4rkOuh+xuzk+75hH
xP3GLweG09kqq5FhbGk6waBC3BRfKesXutWqwlspsouGrqZa1kLpoCg0npmZrqksnn6LTRkK9B8/
MPE1l9bl+gO7PwNLLT9BbNa6lT+S3Pb09C52DUs2R/D+9VLqzyEBpVWsVEEcmt324JaSkdlxJPL6
McV+NTaH+1ZmAeBku94i0VOpfQwSxiOlpJIxgqQICSHDu70oQqnRjpvOYKT3Fu87pLlvJlJDPG37
iCdXCPOpmCTvxG96tMCJJH9L6xI8u7VASUuwejYN1DhVRNwZyykCU5alhynlHjg7bz/ISL/eSi7u
RW1PIdJi1lybOcTeyyvigzACJNRCLLjA7qKHCWj6q7nMWb0z9jpRH0IMO+7EABcF+PdF5Grj/vY6
osN1oVUsba/dZEyWdnua1ln/3XctaEtQcbXXICVBDy880ezhhn4H1RywXetrKl1KGRbTqkbNnb1A
P/9t3LzBNDXP/mZ0AD/sHWfFv6omNh7ywSVpXSYEade23Ux9sPpwRrKctiZ+jWSDpcKNErrHeewz
rYt5WBXaZqfn9vQRmeKe/48B6PZtSHgxbtViugd8n2PJx6Up6mGmGtqCe2z+7Rv2Wdo6IpZ6Zsxp
D2QfQABkpwz+iRS8kzYja6fp9SxpTqkMvybl//QzK7xZN4K1A17w5Mi2K1/ZdqL1+NJh+ossgy4Y
cD5DUdC1F+hBBxU2JydEMhXXdGrLSnU/njsI3NOzgoTEze+MLM2QwpX3h+oBaCeDSLFDDGBAv3DY
Z3dWP+niFodpstNHexXYsn0Uy23b/qaeNv/SJ8pD90G2o5Kd7ctTsX3+Oz8sJOihtA7Pw6d/wXfD
yZdd5kYhLftNV1WSV0vPXPlBMaNCkgkrOHS93HVp4qh/T8ypdf7GeZQxjNPq8cXC1ni1PBryBo19
TgUiXF1J4Nq0L5Ocy8sLQ7KJPLd3SdskRJoCxVU01xsLvI2y3zGoU0DLoz4r7yztMZqYgHmhGV2E
gSc/p1Kt/aGkA7jcNzi40i9bhhlZt4yL+IKBC+mcgkc/YlYCwWZT8sTwMROucDjjCpUj04PwFI5d
cqguPR4W62uBTW325OFjzsaLn66Rbx/INHJSkzLDkhc04I/YikWvc8GvKa3le86kaNMVaTqCDpLz
I8DkKyQWe6IXfSNQDDQyyKdM1R0V+AvITZkfU+NPqtP9MMJgPU4Vj4H23RZw7o8nb+sqPeoHO+og
tmLB2hUq5Cp577V9fiUMQewhCKX9y/Nw5Yr1SzjgyjkyU247xaYFCgUDz2filCh72Z85j+2lmo1o
9DSEglF3BHP1LGBm6twIJit+BXnXu8Yw15cyDhd12ujkRZIOjahHn9pInpnIAI2hqryq+s4sJ9+W
ZowiL0eZnssogTNQnMwUmY2WdLNC5wMwb8Ye+4jXceftpuT3FZh4ZtRgxdwwk3ZvaQ/vVobkFXJf
y3gzV2d06YUuUDioI8s+ojZ2Et20ZbVVch+wr0U98dPASR5h9FvXX2zD11H9RVCTLTevxYxrRGHi
fWaxavMs/1qjgxMtt5f/Mk0QbCgvNv10QFxBBwhXDU4HQz04O9M2KUTRIjuvryjHWwcnowyYAvrO
VamCSaSON4X94pgEpo7JcnklHFn4NuZpxsM9aa6Vb649OkjeelPp07RrhX4gForE8VQAhXf8raec
86KJScNkxNqUGy66lXz9Xtg36aLOklsKAnu6uHHkGjfMYlccQ6s+PMCS300sFedFZGeF5EeaRNhF
pEEebgIJB52smjNqMW/bY7ZmTJv1EOAA8ppJ3iXBo+gJjSN4VGz4C1IWiNzvxf3DfgkWxOjZipyG
2wAr2OBPx7a/miq+i3MSKrBmeQUG7Bp2R5HquRF76PK+3e/WUEU6bUFBVonwjTa9eZ1GjiRoCa9c
5Md61ixJku3Ll4gd+ANWdUT3TMqNPAJliHI8H7Cn5NB0sFoD/pz0byinSSFS+VNL6ZWbz+JcSTVo
IOqtOXWSqJZlJkedO1Zy/eQY7BO2Cn/mNIp0/quvSd3B1mJ0QITgqA6mJdBcxFuf0bsRJX+UNOOg
TPUALKhStFjTZoZyUCLyxIugNRYFC0bvUWRHsdnqfc31DtDd/n+nsiSYYn1EKLkoMIPYKISwDXGg
+c3CtlkNaaLDTR2kt2yj7Ak0lCSJY6cz+ipTSDGRPMFIxNUdgzEDBQYFjOyd8VOOxiT3vS7xN2Uv
mhwClsFi3BaHhnCiTo7eNnNywiO5QOadHC9wga3XCUmhyWwsUtVtz8EgMW89TufnQfUMFT1+wT3X
v8Xhaz6Q2/dXuOfuFXps4/6pXgAyfIkGP53jodrr6H79q0aew3/KlUhW8Nko97koxbC0r6kFum31
YUsHVPu6ENu0Kz5bN173zergiep0jPWQk+jdehp6vwXlijimvbEKjm0Z8R8lJOYYtmMzE5Q6cDF5
sky9eaOEJlWQfbNV27XD4ekqqj8mvblqNKCtj0/waDUqFo22J6p1UZV/OXFQgAwUEKBbzafi+dFT
ryKobs88Q2VWuxNHZFCTlKLPNulOpqnw2QapG//n1gEUQ41ZfEFixmSB0JHd/Mfg6STwq0wnj/Aq
xSXdeYW/VTyF3Bg40jkfj4Dl++EQNgRlIGutApu99D+OKaI1WIqKNbis9QOFaLehTiMf+Gv5S0EP
Kx1rN1E2x2kL5Q+J6z4iSV94uX03gUHsUQEzOgn1axbnCaGhfudaFiGH9/sJ3QL8mLATGnC5a2xy
5ZY3v9LQh4K9b5o/YhUDIn7KRDAg78qmiKFMWN9QJHgUq6+A+kCy6AOiSeYSaqmW6o5PCpO/R782
ZLRRP+pCVSZaZACYi+NjJOI9azIc7qzoi03zI8x2Q2vDIvKJU1ZlUj7WJ2C/iprZ7SCUxybCk2n7
IuTZzDudkLRmJJ19UJN5m5DQtWRIkIQGDIY9YJmQ/TIXzIoPVnw8ygI7/cj2iOQGAxplNzvh/jBs
VM7IMdFxoEE8pZZidKVmHI+9Cq1PAU3yXYquFZ+ti1OlYxW7mPtjgxsnNSaSjzz9v971gCYvrSOf
eo0GuEZYoh8NsU1H6FbWKixJW3s2ojrSrCtTNeV1f6V4gqRg3/5oyqIe7fShQWNhnYpmb+vsBpcJ
16motJvRBCPZUYxqb2WyN+/UAc0S2myNqLrXKw+USyz3eG9UcOmkSmYYrlZtv3V/BCp0T2yrEOo7
pECNvspf12mQruPktl+jcSbK2sBd3AXnGkoagTZuz9dhDzt+pj/zCf+sdLAQTdtY48iOm+/kcaQZ
XcPDSzQ0NXDWItfFQ8waih9+rj7wpVMjUhoJxzy2dOCy5YZFqBOh99gPWRU2qCL7+DuzWA+6clAd
QO78rtMh4PEPjVkQB5MF9k/okGauSDKmIvjEDW0u/KZZNF9xUQlE1pYYjKp1MjHwMEXkoZoWOJPW
1jl2q0o1my5PmEf9pYZK9XMWjN0hqyxrtskzqx2H1k4u4SUPVXYdAU5d1vmpBjQz0So3vosp0pcH
k3pYZqJB0dxGkG5sVpEHTLNdS4Fk09mhHdUMVhM4bsiKOdhrNA7kOnwG35P8VXnxm1HZxSfV3EOZ
krqHTUVTGYMH6aHPn0RCchO+TljGOOaklgbxOXM05atriOkgIl9cSCvYE4fsqT/AdzK0IFZpijH3
+woBmWaxPQh3YOMudu1PsXfmzRyTsAtCQLUcs3FTabjOxjQRU+cgBWRW2U0r69AVVW21BWPOUdDc
DWyU2mXgSTDCbyk1HMRlpGSj5qDnSnhZa52vf1vzsPqsXlntRHUwZ6Zx9bjAa4AYKi8SMEd8Py4W
1dedoPrWq1+BWwol38gh5HBQas6fOOO9ECx6QctE3jqbP1nno6qaVxw9KsChoT8yaSYRh8nY9NLY
Om2UzPsN8dd1M/OgRbuLWLRngTd0fus7qbkvlpWZ6GLkGMh5wL5c9lVnkg5PAouGZqVA6CTtvfn5
XoTvnMwOCHHYK+1hErOufYdMVH1slh7nhghg39BQeC9o3sP5G/Kcbw/q5vnjjYZvbq4YWMseRGzr
M/b1KumZkMz3OGDIP0YapYZzysQdTB5eNBoRSN61lMsm3LT5OLz2kElAvTYjI10N+j2AbERMHsla
ikmnpyCHH6cesW/tEAR5zlORnE0SYj0uNq1PkMbJy2BKryFtRcpz/dSPZSbQGxuNWBK+5fFT1Q0L
DT44sCIdteyBqrY8MCeRLEhYgpMXacQlqx35t1xF3BftHzgGUil4oSvWeWmC0Ppwa5l6fMRcCn0S
Y4znJ3+2FsEuWR5lkrlkiU7EjnkbvIRBrFPZFJAs1mvC01d9Da5fK2elvFN2bd5JmHVm3TP9yCYJ
vXw8OMKuP1ixjyDghpQy8E7loklfa8RIggC0mPTc7nBSPTJjreMWbIbbmClOmp3Lx1DcJ2HpSFmH
1CZR+FEpPfL/81fRP1iDWKdC9RkgHkjCEPbFhbyC7Jgo9pfeeOJehtb6/Np6e2P82VEYN5mVyKUF
079kUO3RteyyGULjs93OIlvg03s7/eQnsT+SEwXYnRFBMPv8vD+2vPbzB5Uq33RbmL4mowzH8fMP
QRpGlR4Yj3hWbt16C+z0chG0LvnTHFlBXpVv4pq0Ag053unGcytp9/PQ4vkkJ1cKi1idU0o/odBz
WbTo84u60Y7Tlq2tERgSSs+mqmJ/TOfzP8oZUhn9Gaf5L1oAs0X3ccGtiS91xzMPSXZ2JXonhevd
n83+QvxgNdZ3OJcWtcR6gZ8qVp8E3l0ZpiB89Rl0lAYv4Oh+znVPWe9he09LbMhAehok0m5fY9Gn
fMTQsWpi1lyxwkuIS0UKZzfKtwhojFUR5WCYh2z1+69xA9UPk8EaaDtFQnNNf4xJnmhMUCNPi7XW
3ZO/38KWrE4igDLDRtcnd9IU1uDMPx3V3qtxPzd6tDBKwQG2K8T7uBAfpm2pfcEOjNjYWW/Oj38c
m//FdVnop8aLc4GPTj86Nif4u+s6T5J70bz+/sRlqSC8KcmugYBp2qRAJSnaoeK5/s6mmFJBkHhx
Hay8zSeOooGx1OteAOFBmWF3pkB4ZI3otsfSyLpRZ2mWqkDGYRJzEbVvTrquVAv/GxwXtvBzb0du
+0y7XYQ6weIKEjJyixnD2rCMla8mxQJ2Fcw5ecvADX+gzKyiBj99u4/z+ziNOEWtiJ29co4+jKIO
9LIe106iEvIaHru8xksOrjnaiJICnegUGWZw30ZXjMkcRL6TtXtrzY6rIgF+z57yxA2bhCbtkwf/
UeFNgcs2IfwMf4YMln0pW1KYr2Nn/l7veG95igUdnik2OZOpF2MsPBMdpUn00iEMPFYjIk/szyzh
c10wakbDBwQEIQCLyEClZqa4zBkdJE+siFCn+D+nx/mgZlMKfNxc1qVNR4Ov5rAouL81Bu6jY+E6
rkKppBYy4xO3sdc8AVXqR4rNxA5c/JGhvR9dCcUIkYG0LBePfgTp5T57087E62d9fSCUiBql2Cdr
9uNPe4Gcg32Z0OiMa7O6N9eDMLVKOXx8bXKRhFEo9CIXIDCjJNPIbBi+DOa6fyxfw7AMafP6fyru
fiAiW8XKDu3xpEUsqgVZdmVcDyM4O9s6LBhDaYfvlMfP4kesv30vbp1cKFIVbci1hmatFLRugA6O
D2nmE9PQPsX0a9pT/lh/omuqKsFdbe3TgSRnzW3zm2oXjPjzmzj39I66r6CBMfJ/KxPmazLwKZ0R
RX8Vc5eTnjYfUlGeydkRDcGghZoAcSf9s5LI/ge/YHVC4i6FSZ1Rm2PnwM3PAxCDZfSwBHakz7ws
J5+eGkYl9DrYM5rxqcGm+OpAWEqaoNgBi4vzYjUEyFMGB0goTpUzwXsnOavtR/Qa56YAxjefOCgh
I8ocEelbebA0j4S7okU5ieQug+Q11Q9Uu15NC69pWWooiprvGIfWXbWun7YjX4kHp2unuNo7eqSu
Y2FwItv4q60ypyaliCkWcvZSs1FX06aOaV92wnbt0N4R+txu/UHKTB7ZpNeUCq3YXrd1zKaEUKht
IiUzTFq6RI8adRQ9EdMU3VEfqMdnafIZ7g8+7HsHjMpE6Zb4hHxbw/s4F+qGFbJCe7365en/yU48
IQW/hc3ntZ3hMVIBMvG+lMVCjPyNgmLkEv+q81geL7pmBmwUkB7BHOHbAOf/dSjIFjlUrzU1V11J
WiL26ld2dFGSI+bpB9rykg8iYzEy8A/T1XJ4AbEak06Y9awr9oMMRYQWSvVbYqqVz2D3Cqe2024s
NWbOTOg5tRHqP1ifXOEjsRCXVye/VfTYMK5FWkohH4+u8t5WAvlcAfKUZxr+56KYyG1hnwFcNzXM
qpjw9l8csRGkOB1nDqngdrbZoGClvk+qr8zLk66zXC2fKlYOFPpORQbOnwI1JY0BIBS2dp72k+05
tSHvHTKxCDPFD3DNSlps/ZwAalJjPhqK+L6jc9LRxxqpob1y+PdvvScyt8AuAqyTvO1d8fRo9IeS
myjGMtsLAnB3UcHzb70xFA62xXSPT+09S93qTfdnpU+8YZ0ikcndyH4+tNuI+NX9ijrarG70yOs4
KeNyhzMYX385qKuhkY8roWVUdsv9+W6VXaUIadTUiMAID3uaJ0TJTRABnNIFReV1aKCxqdb1Ps1Z
MqDu1v4rAgdcyrTMCgdCic3iLZ18rQeLloEjFzjf+3lXbHlZeP758JdKBcmG6Q+7ogYU6f6TeyHZ
yFdvwM8PdQQ7KuGX9INojSD5p+t9nSql+0933Qw8+EOMjaqQvx4t4rZxyC7zdnYTbVOnaDPFKJE0
VlKd/eSIWwSxdSaVhbXOU+dyPNnaP38AyQXBgrtmg1cs7ge3zzsE2+fLbvJya1LIcPIllGCk3FCP
nWG6eJzEqeThUN+gaEs7G8H3Uect2aX/Ul6cYiLbmYUMSNrhJoktX338EKjHG0lkfZxUePNo9zuw
8/7/v525FLYps+TywGXaGiL7PK89QiqNxeSfnUfcSmJ/XNXOIcMEwej6YqQgSAZ0vZFnI3ath/+E
GXESaG3u/+MZLQGY6zelquhwgg+sVfpx15suKNjNtktKaB8W2kpoLhZE8mAtiJ217BwLW9QYVPo0
qJCMVa3S0Ht2Piat9ktWD//sd/x63ibmFLzHUW5laQyrJZP5sgYsKT+wRSn9IQkFUp9i0hMMiqsn
VM3qmo5y/YPEpQ4xuicUa8VkhOYKWvNqN6nSxTRox7Ex9/fChiOczrvbqmmVhwI1ENHV6kM8Q4Am
GWeXSYaFpnC5L9tjAutyMGQtfxfsMa9pupbsH4tZkcDw1EeM9a8atEfQVmi5YWB9W7aJx1yT+i5P
QvZbixHQ7ho6tI4m2/tVBrvyNO6l6BOdDBrNrznqEhfpqViIxZe6F7MLQtcHK/gW6nMCdfMbvcsn
TXuSfcSDjuFh1o8pV8+IeunPmKrkm5mAQpzTTMpy9maN9rUWXgVvm+4ekvhHMlnYZPYtQT1uQCt7
FP11VYL9KTB6QX0+lfXnZ3WkvFotMQK4I+C5jjpKarpCj0nQb88RldI+LT9sbDZviqYVSf+1P1XW
ysKgUb0nPkJpXSLzFIaSP0GGo+6SNf36tILIm90ju6E96mQ/ia6r7WcNOI+jl05gMpniUVbmCpNJ
QU7tgKg0m/4wheiFrqku9U7FXsWek90zAU2/ed8N4SqCIO572mfusqrvIKGhxnM/T5Pry5QGdef8
9BpjQQxq2AMSYk2OK7j/FSfgeoZWSYJYIW7SuLqkv4hOyATYgXlp+ubrbQafhlHRoznolkhHjOac
hguWFS5RSFKW6CUJIeb8oDnI/lBW6Tu+meWhGB/lAvZg8E7zTA2gNpo6EuU3dykfFvqO6nqw/T0F
SpPu2VfvCbhzQKxHl4wr36YGHgkDhjVglbJcGbZdUvvjDg17x8IjETb4u5ZiXDv/Qjlf4dHhb4Ok
QfrPeEQ/dkrP/HOo/U6wndQL7NfZWUzwPlU7Z4B92MV5CZzpSm1xmsse+C9VEFhgeMOpOmtWf/D0
yKwYniLk5/7L35kdog5j5d/beUHRPJJvV+F197U7wru8w1H0fTM9DqWJqXv/S/d0HdNJv9RHqY3W
W/f0podcZL+2N9QsF+rpI5Mbidt2p7e0r2S9LhZe7SEpJUSf8nfqNG24WLTqduPrRTV1EqTaMn5O
1aTmAFXgraoVl5bGCMlsC7gGDm6w5QP0kFw0zyq37eSQLnk3SSaT6jEwURTvEZi78R8HT/1PyUiE
FEV6OdyT6VptR1uZ3nquTcGuWUODFp84STEaJhjOPV2GOUojYJheZ8wHFktNug/RBqqPzOqy/BOq
dHZtWw53ltUEjBuVBrmSKZDOMtFrPB/uXEye+wEsDf8NCLj1z51FYWuxcQDwjHjJiYmIPyOT5NVA
Fk7mrRGVWB67Tn9LrKN7/6V/1VxwzwpXCqzvR0wvM2KOYCMpuefdh+fX9/dnEvuSOV7S2sFOKO/d
CjZfvxvooXgsiEADFIY8ExxqysE5axnu5uuX3UAcbpoq/JAaTlZaI0SYQK8vgczRZLhCVt7Xc21q
OxUd+ERTlHKw+QDEqXH7ie+ISXFl2isLLl+7NYwpKH3jpeGeFHfRHmht9vQsH46xvdtJ9dvp7gXB
ON3zWwnJUaVW0c9Y12Fggs5PPPxCrQ/++7rFlnispzkeaFTuT7f/A0MKLC6lmYKjgLxuIx0s6wzL
WgoUz69XheY9J7J8faXEqFviiWbXqtlYrLa4NQeGpvzkvUnyqLil+Uc3YxhNO8UzsaoC+DuGEgqA
EwukxgNpC/TCA78mucIO0tBO8Hci8HXzUmVmoiZgCYCWlwQpJM2MV64qCb3KtRQVZGEdFnRMI08q
I6TrkrZidpLCwHcaVe/5rido9SzQRHNElXgQNsuhpjmrqxCBLcZf5pNn1xeu4xkipsRUrUTgRbDo
sXvqeaLq3Xi3Ub+aJgpiqlEQImlCQ8NhxfP3oiU9BFqKHz7XpFSNzrhbDmc6MXgb3dqz8pJt/evE
+aR2Ms0b+b2Xn5zRCRX5JY4D2N9WrhBO7mjETYD5dTqbPA3XlepdmjDFLMlDDpx7yWPgP3KDGks/
yDknvHXU1daX8QlNqBrD/rt9CHSGVmR7RSmNwHiV51HXpO+N6rrnTuHY/FKghxhrjHEUdxtyR4Hx
KsjHX3dyN67AaK44HAP30pCgXHJFJqG7Tjc5BvdEHlw8SFKsXrsomc6k1U1W5YuQ5KNY4xRVzUh3
8fbpR71IfuANd/cl9rTcWq7xYJylY2L1Yj+VkuenI2ze3C7X1+ay22E3yMD4iZiPwulyZK3tfP7c
PuQ7WtJWRDTb2FSn6TjkmFWfyg3P18TiF4c+Z00XxTGnS7KteWdl9LT39S1rrFx8WRzP3UEOTaGa
9onJgZi/0quiZFu35m2Zk17vn5SSo0NvvInowi5eSPGKUAe0APps92Q0LMzKyQOQuoVD0UMjfImy
+m62R1NSFMEwTCgsN+Wa1vkeZm3Q2c33FBYGi2QB/2Nmk1NPHMeOFpFKUzf1hOR4f/37YgeW6Ytq
WNU7hi9zkSxfKzY431EntYrMNLfvoTAEDiZ0Ze87T+Eh/legf2jVyVyvdZFdxRQ7dcHsC3vY9Gaj
xPPkGiVygbsxmVf9If6FntXfVKI2W7jJ/HtiNHhVEYixZ5zEf1pdMeb7S9U4WrVuLP8KVE6Zqop2
0LxYhR1n1sw8GDL6Wd0lp+l/wVsmTX8MVCScWzLnfnqfdVVlTC9Yfr72xhYXQ14c5X1UKbL7db6D
oWTmGDkrGfT+J7kEf5MMFn2oQKA08PYS7Jw+F6a/kR5bFymGZoYtAODNwxl6QOU6wCxQ6Gp6lxBE
ME2Oe5TeFI18ZUS6QzWN2JKHfMpLU9kC+xLLwKkYbmkz65J/JrcaJZ+xedLQxaJy0Vyj9uZNJcXJ
X4KLEP4hPuffTQsY5Aa/nkc/izka7SR3Rk7wqVgpgDKGxFn5B49E+DhQDJpN1Q8YGfu0bI8I9ws9
Lm9feyKao1ZPlEoj1THwLhbhNgZ08t1IAXHuoKKo0sJzvOn2++B4J3MBy/z15n++RkhS11UCKKS+
UE0bryf+csG4QAvSyeSjYb2eutVelOwLaDI0I4nqiU5TlcojpgRo4TxchHyWoORWMAR0Vz2KI9ni
qsLAgnU/zFL4Q2gnfUPktzS0LAN2Yh/k5NQv74NxdI3Ayb5vN0Q/ta0jRuuM3H6M+xqsPo0Ieezn
1cXiNqaaI0O45YIzk8QFXlfoMdo8I9rTzdFPDx9h5wQCh4hX927KtIvXbKe+DidTihD2JdCsCziM
u51dwbIqDRFLsmyONeqS85KXDzJelrEN3mBn6X8AndHswdzor1ixI65M/jxh2Fj28TitQ20GZl7r
X+vP+idIU2RlbqVl1cS3c1bKeh6av3xnkI/yOZRtGMP4fc2B3QSG7tg8XszfnCKlEeaIPuOYypKj
Dt9ZTnMe6WYV+Yf5Lqi7tdFt9+KY0rFMSaJCjXVATXXi76FUGrdMil+mPeIdBLhl83sPdJ+h6Y2/
pimxP28VADr2OsqgXDj5eek/F1NtL3sbfQv9oNwKtswBFJkKwH3u6Kvp0CC3CUcvYZiqirSHnUFH
CtbHL06IOC5cCa2kFHl62MKVfU/YByxAiIf/jMf1rSRSfvDPFmMwxezIu38LxWByr7GqFVdRIwik
QDLZSLpfB88+5MLO+zI/6hgIViDcxqVhdDDz61p9kZcVOBoJMPGhmsRjKSbEnaR6XMciapCJnA3p
8NpvYxjlRvn3p/fbfE9aa19eRlEEZYT2ZLBzKKYix2C4ZezZl82GCl8FmebUJZ/O4z8SVK4uTO31
8EoryKFEthDdd4xwg+Z+XAPMLJG89POwwWTbL9WuVtxHzfZkqmUtxfVLhdEVfQEAmXFo1mdjTRW4
z33xQmG6BqHpB8fZ5nsHkAsfJmzzy5LWLeAoncCe6yxFKPZkLVB+OeKZLBPCpbRJySW1m4nAOy1U
PQFx4YQKQOuzkScrYKl0rCNjFnahouYgl1W7VcwVYnAfa2x2aVrFSqodp/mORNH8aUFTm//k0hTU
ss6VDs4R8ZgeatxewBjZJg2Ku2VJCaO46vs1zy4ITcb68AKygaC2suQP546xFZDUxLuOnzR8L2x0
TURvNZ5PQKvC+PwN7oD//020UD/iX0wTaBLCqUVGSR/NcgOcp9U2Yp1q9A98NPGNglB8LoOj/aBx
oWxR9tHU4tCs9t/roOIlzP7ABp+Rt35I/0pWCLzhUSNB6wYzU4Uas6j3c5ZifBf1AqOtPuFMU3tK
rTypK9MhfZ+pDjzZvgEabrVxBrX5kZ3qo+dYH15ZMG6Nk9vqwbgNmHPEZv7PPSmqcQlA3MO9vHQd
JgNUxP6PfyYXCY5kxfTOCQT6OadNTDgODAzLGp8ICi5KFBGHpKbADzdKayF6n2mWiewPqaswH1K1
YT1c+FURRbAjTtt+oHAAeaCAXwmlmvtWQGjrrgW2C60bCdhw9ktFOAY3pHHUmGXWwlV4Q0Slkqvf
mxWYdtwpFLUxh33fJsRofD6YGsGGwAmL86QTFc6i4E+DlbjXC82hrq44FXr9lyAWPPzwwMkIseaQ
XYg0U07DOVwIu2p2Um3Aa7oxyThzVgh86yROJ198B8gcs/1m8uYBz1QoqtYCTBCrwlcvyhyPYkg3
ctqjsiq1b4E2TEXPbjuWGONSt9Vhh8jNp0r9+lnEigv1TjLaooG9NUpyZ3R0jRfn7Uvb1c37g7kE
Q8oyGiKzJW30bfz299fPvCOqf6SpGlEoU+dmmyScpooX+Y6aoC/sVl8i3GUvr25tPymL+HJVKSbP
GCOeMvsZK8RYnttRxjpPNt7qKlAd9gpLyUyvzfzw3pM/H20iu1HrW27Qjy2KA9Di4mn3uPr/H4Fw
SZ3ZF7jGDxxy/LWyzHKS9T1rfIZO4SLSTsi+ZqxbKYbiEyMjsfZO4uNa0quAv3hOa5WuUqVcw52I
ul+kBoOuelp2u8fiBgE11NgbwDgW4l2Vwh2gQB9keQhgcDWehg2+ASu+20vtW4i6Zqp8ASYiItYB
FNQ819zaQY/5zF5t1g7jNdvFEKdAVcX0ybKpTZAeo3NxmWBwqNyh7wZVQtprBlqFAH6nVh3wcebG
jHDlWG4aIzCdwPM9UjWEVHQlj6foiFuWREuAt75Cg7EZQ6/zPuV9ECV4gzdnMiPB7YBEVcyviQD/
AL6LH0+Cp6ihvgQ1MvkpHE0IDEujqsk5JutPGPRlr7/1GGlwBSG6vNjoEWyXsiJwr9wrL2rrn2nf
8aYOGO6+9wKXcQABpmxQ25TPDbmYT8fxUidCqy4CViMF6m70olUM7MP0Qtcml7IM4aVKOWflMEZN
p0zxC6qe7oQsOoT40o53RL//sUTf4lK0dF36v/UvJaKEmmkvM22tTFpR7Tv+kf5Zcdb725uB1QIj
MqrLas5X/D8utijcAjka/XADUAWHiCx1TdfcForsxoiEyhN1B/hfKcvI4eR4Qj/+NzD4OeoWZMn1
nOc10l9AL4mJLvoPVj3gh5PbcTUNfpBviRDFlcmV6L7O0WBI7S4emjM/CCU5TAUR2BXAiYEV1WU1
dqUaLE74iG2WQ6CmqdjPxK5Y55+mhSMIokW7WriWw7cmdQIJwvUi5bAMVbCRR/zZaF5TUzbRhHBk
95KUdDO+hyHWFHG/RcnX2rMcZOjb62RQDQmpa+V+FylzcbWoAPyZbZaTaGSxqlpFIGni6JbIAD9/
3/eiECVsNFFUdRVdRrNpv4czcDqIR8G0oI2+GKqDVPlcBhXSU6NGCM0MIdyiMJTNJFMMV6AGbQom
UQgSPo3jVVJXv3Yjt3A0dZh8S6+b5fpdtDfjRs1QyDaJG1L/n/nB467pDBg5+cjmMVNRxQc1NEeN
w++nLm7EX3HwFoZZr2IWLSzFUf+9IsDvsdwtpnKBTE9uF7yYWWWjJJzl25fVnqzSh+aGHHQCZZpK
qRYTooiMwX/GZvZkhWtq/vN9WHYQREqLym9dZSYxvHA7/5/aNbFGBbFHoRYPZ9QNt/juNYL1smqO
LVpTm9Ddpo4X5Fqdwf6AhIi/SSEEGmP9cAa+vAoC/eNDpkkMPl3ma+vPpDjZVvSgM8xb6jo09MHQ
VU81BqZ22iUwBPm0G+N3yVHR03pT1sdb54KqsInwl3kkvxErLzRmPe2Zx2e9opMMkkUY0vL/Rf0y
CXKRA1KL/CVHbyk/UnIweuxKeZENpuL4EosGbWS0UzFCpr3RnRMmRJ+8HvgmOPXhH4fNgM/VN5k4
5RP8zF/OdXVxKq9ImcJ0Z12o60KRJVkv0yoKnpgJ18X6VDmklHr+GW3bXvM2CGjY/K08HosYsy5j
TJMatVQOKyELdJ7NDiDqp+UPbQg3ehHqIojwwbP3xWdO2y4i/KUPAaWBhs6FbuSrxIsOEgtSyvpF
DMxAb9sLzn8JDf2IXf2HeHzdy6XuGXZj1UxNAeyJ2fgPzzaCBXnK7v9/Jl9uDzGcsNzgGMoYJju2
444mlSf9oTYlJsRc5wuPYOOJq5/yC3vEmRuGAqKu+dBfvkSF4DY4CiiiVzBfhubAoGMLhsfrKv4w
B5IwCgHbNIp1pXV8XVfqrKuFgdmAESzJ6KED9eGksDytZB2pAqb8F8AL1B9jdEHPZ/0/a+DHfKDB
6/S1H2SJaIHlIWXCcQtLRUFkU3tKlOnzJlS5uWjnJJzUflYLOX8fgITJc7lPOn8GnG51BmKeQJUx
/jZkHZBThBQ+z0kFfM5X3Uy5zkiZ3EphahIqpIf4vJ+e36z6ZF2LlcI+c65vDW2ViRafmxJ/AJtZ
atqvdJ6Wv+uIexnYEsXoGpfsPls9lN5jU9q2CPT5CIlN+vaC2kYfeXdMpv5jYZgre3GfgV5eeuaC
G+gwin8NJ4G5FbrTDV2CcUM1wjx1ucUsWiehSYl8cyARLnh/TNeyykJihu4GvcsiAzCUWLGvBEJ6
+aWToWnD7P/E+2GCE3TjDFAXgQZV21ulwxQMoeBw/Y30bI63CzIottjCpjZkbz+7E4kARXhMLWol
C+VML8DTkHHA7K2YbYJYqIke5Bd+F0zwfOExSPM1tsR2Gpvn1Xyg9fGnaUxLHcoiMpf+7ngQsCBj
wz2z3QknmUcWPczjBjqY1QtsKJ2B0hCF4az9BZ1Qtj2Aod9sV2dKgyqYG1c5lYCqXBTWWj4A0CDs
EJ9Ro92d8L5ivehlC8c/lxDSBl/rep9CtL4t6NzsfMZC7NEnDkK+hbfOwNXh+JHHbSVmJZFdLYYm
U2QHqWNwp0Jbk50tOj6WRzmwAJcWXOQY4rRb49efS2hhN9xebpv1M8COn/KbU8jIHWYyGDRkJ/iE
eScYXI9oWaT0pb43vrQY7OpCciXjzW1BxJ2SqxUj59+hsbi1UpOi7uVNK/SUvK4iuhgACvhAeyRm
lNSi+5fifOcQtbOPDQ73vtDS+QcpwJ+8xesI1ZgP3O+R3C6neW4SqB23cfBWuNPRA8b/ElHw5DLl
EwFgJbvnakufht8nW74s9O4zppzDXNJ6V7bUUyUdYILODthLfEnNHB23GTGf/DbpQeijVTbdBZpY
pmyriJclsLtlH+H06aaUDwfgNpgn5WNMHeIK+nJffcjAjNp/IyinbmJOIRvG12HElGE4tzTenI7p
xAoBn3uYsHj+tJ2ha0+MoIKIb8gfPcdOm8qLpewN+l/eBp9KSEEFzOClPbcAqFx3K8pAXM+q87ys
oa8PMwAywrU5kBCRANgwGISaaQTA0o1osc88rYNTelAgzYReCJ0ChmnuCzvux3t/qXh0WI2Sd5IW
NtW9Dko84PPEdXNkh6KIGLpwtyDlY1pdRmPnWr03hwqH1hmYljPn5Bg02EN0LD+euVw2H9a+7pdl
fPd4wlHeX8QNDcW2qggn6r/MYUI+WLv86b9wbQ2GQo++Ntj/faPzfhpjXBuUJlQ0qbP3qC+UOT8K
DwdxDTnRY+XNUh3/q6lN2rJ4ZsbngoYahMBK3HUn+XrH51VoawYdthXQZl84+tVD/xezBEePuSTl
oL/lBP3FUs6DBZ0JcALXsqeX4o3jtZslk4AE7oB8+u311e8cvd9RO/xbah51TTaomcugTU0YdZlr
NlAWNYthg+r74gHU7SqhHFU8KbCT6pTI/fjphYSDHMysrTg+Vgtb/TXHXw9jAMz5gI7OZIOv0pq+
lqGOT+u2aejNm9p+0Ztu3kXeeGj8IGmWBmHmdGNXvqwZExwsQVjxjRPcjbEOc8gFthqKrdOXYUTD
9jhRCUA753zYXr+GdhsbV7iM+XQjy67i61dbk2ROsaxmiCHR1ZXozyjNkCT7jK9mAYyoPcZE0MBb
73hDOH1MpqC2zLjnKnXej8N5Hhm2m6SR5vbjLIzqEN2CTfaaBFc2ZlAGzlpl0J/fzaiPbtK+tzcL
s6wUl7uYBPQqqCp/NGKnL0OWUyIckOjD3JrspKVY/00PGWY47Rtxb9681BAoNnfy2/nKOygX7YoE
ePazZkX6/508hSl90iL4vI7+uPxSpuez69lUQPMjoHasRXFN6tDIrDL/R/fDGJ40DLd1Io+L5H/3
UdEXhur28sfJ+IhyZ/+1nfF14/SBeoMk8l6l+d7/cM+13hcbEtCSsjR3ghjGhXr+W2IkE9g6r4d3
vPwVpYA/A0Gaf+K90L7nOLTH95urHvBzJJqgJZ2vVqwDQYa20nR5vxbgTwKiQo0BAjeKwk/R5wsS
TElee0UA0vdYzlo/7bJldj7Rh2jyB4vLyStkjm6VCNvVMGvTI4sXhol2yvzPgjvk8jGNlmlC2f/B
N99DqBYzObyvBN9ahW5clIOgZAPinLkUrSCokqK9KyeDD38VQv3D8lm3XyR1FdXLtyh9p6I8339p
uNFsxu7nfF4azs9GAPI4+bgLiiqPkIFZtXHqeFgi+QNWuBVitP4hhVV9D75512D8r1rJwUJNPou5
TN6CXGSLVtqr2mPf3MPV7KxLccg84tcplyDEfqSpH5I8IxgvbOjqJIwQasGeeTpN8dMAFrwIxfkv
BDL4syOJh8NbVqJaXDdEM5sXKY8+swf4AnqdVuvc2AhENddCwGCLMlVebiCw4sI4hLXGOiXLHlBr
bgIloaizq7bwlES9umWDZrXf2CWlKkx9wfMfaxTsTNVy6WtIVGlf8RqzJ9/RBKnvddzHP5PDWtOE
QgOislO30oEhaLAK2YZH2F/kK71XkeIiWXth1zT+BnRP2Brt7tp0dDp534xKBdcBi14+uUVMtrI1
bBKEE6UzdYm5ycRbBFlL4whwxPNfTrNoJ3JHgReRoXwjtrxWB5T1KcRc5WqZOI43hMdQmShekRvS
fKHCwE9pReLdnLJTsrzQmAtOiEvjprGpjnAAmB0FFW07WfNFquQMWNg+NMPmcacv31Xw1FiAJ1zm
VTffPXVfnzlXyBYQLcrvwruDgnUuq2s6xB1ZSumLYQP2Vu8f0lD7l9BKqr06NtqQN2Gj/A8g7Kei
ImkxmBawgxHWFJnLxHY361LsV1OkleLqcIdJi2iN9IZ91VbyRlAOkTGbH7+K6989g9R028ID0FKD
HWngVqNFalVhqe6FoxnWqqAHobcc+LSVDkwcGtEn8Xzt7w8nyn3JQzggzrL8ZQrjgyqYgaQfP8oG
7zS2KroUnxloV1wMawWLtXxR05cGYiXclZQ04vqxjMf2JT7mWCXO+R583MDBtiYxSXZV0+glZuPi
0ddAESrS+63RTzkHOkS2/rmQaibY1GNqaDG4U+yF315BV+bFhBiBxZeWzNCi+nJlVTTlU/EJMRoP
wDokX+Jm3lgnxS2L47imdLSekpIa7dOL/yX1AhMXsTfCZ/cfmoXBzKIdIh60B2t8hLS6WkQWkfFb
EUs9F/YRIO4E8v5a7m0Z62ZzLYdCjn8flVnO3Vtrc+ps60KMAXZ2G3TXArNjatfxR8s7dDcUGfwN
EA1/VZi3r8AHn+GvsReaF7r/0KaOURD1Exkq1ww6xSjAPH1lklZ1CobP/Ku3RQyPKpg24BYwdTtI
T3kXJX1CTKvvPrrOEH7aWOWp+XEKIEw0S+Luf9EGbo4rjG/ZSHYZ22p695E5DDD9XpLj6WgaewrH
EHd9wWiL/ZERXG0xVPrbYuTT2nktjJsUXI7c8uVLR4XDA8ZdBVpPsYKKhLCnBUg3BoDKg0EQ/alH
OorUyoT7uh+ynWcVPmiexnfhf47sVFN14BuFziwRCKtgopQDyEyJ/XDW6EB26orUYCF4p6u6I69w
VKQW6G7y9q4pSISeKPZ/uviobN6VS31yPHelQFO7cY5k9p+MRSaaKiLiOTJMFSZ0/ozgb062R/6B
i2edi3NymZH6xlHNPEjCLYVpMAih/wtGjYxKjTtgTMFP5vd+efqD1e1vllJ0cnMpeABUZCVOVL2Q
KPKRwksKWSx51lHh0Q5drrLfzOWOu1Fwg9M7SPNjJoEvm1AXckOx0FkXZc0nbtIAzIiIMwTTp0vc
51rGZWD07yr5CjLJjd01gPBHyfB6W1rDzw7D2Z8/4X9yI0BzYejmV7x2TiN1qzL+vTH+55uv7pJK
nehkQ7oEnv8ZhBWm7rfhav2z2wGwKoV+vA2bAThzHUIOtlB4YzyhgzroWqI0gMC6K/9RdeXmMxg0
5pf/78aylN851Okgd/jFDjgiq4VFtaxjTg7dw59HDI7i5jaqCwrRfcABaiKDs/Uk6reIywMeM/K5
fVZ5YtatftBrlBLlNGY6KFhErXO7wYA1bROm+9qsCev1pP84zyGXzxfNioLM2LqGRohN1hB8xt0m
+/6Q+TlcmHSX3G1m1430qLLBnwEXLMhA5NLe6K1X9PeXXEUODN7kOCxbDpO904uZ2vlXWMfA1z4A
yCe+atIBdAXEvYbkYmqnG1VNQ105zTcN+VIyWtYFIq89EEc+WhADiX6nrGjO97R1UHtD7GfVzggY
c0U/8a2i/88QX2le1K8dPn/6hh+bhvkggdAbipqrAxKRFFmcpNc2aGMRcxs7VBRTu5hFVtuOpzUy
/vfzJSeSiuDX5A4XbsZWdUW+yyHsborY/uRNd2AgtMTIYzYdysCo94DnqbGQVRDK/LYu29SOZerh
Z5GF7ZWBWJzOUKYJcf25hPk0Rwn0xwEMDbVYYXgDtWsBKn4mwrE8ucyVTq2W6hP+sToRadkkRS8W
jKRFLkm1dLrLtmWPxHwJJ4E7fZlhtNPSgq4M0PFhpSQGAg9dFZzFvM/FA84oYTYrNHjvb6UPtvk+
0oGxl0tHYJ2uvzRtPzTZkbPJC2N4JjDkikFE34fyIf/ZDKCJADBBdjgKs9nJKqLBfVzI/qIEnRlO
avAqkpLequOV0ck05/aCBx8EDd4mhzclgOneR5BQeqsOehHnqWNi0oBaNQvMyO1Vz37kvPVYK7wR
FrqZC8BwDYWPiF4v6u1CG07NQ9BoW/WSZFyO+7I21hG7PAacEPVgonI7kth7g+qxNWqYjo17YqCw
otkn+nPGySiM0cAH3f8GbY74ZJao14KNaSpg+4LDd1eBrvrkwXdd7EWLQbRTp60Y5EGzkMGgzuRK
RLyWjqueqnN30z62kASs3MeqYm/lv/TR8aRDmwQhTDBE9L9oy1xH4jzzANP2JIvQ7DHQ0N0JRaZ1
PgglMPhv2gowzDXDph+UpbV0pADogqL3U6vKOq3mSk5S4KK23m5UR9HxJifnwMsaQuAmXMBE+Vel
atsybGhXTuYKheyNVsXYkirEC1WY+QVdkvmAg8+lwrViukOg0UX24jJDGFtQ/xzI2owYNNyKR6te
lJTzeLlV54Ggp/3OcV+od5jBankONExn6Y3ZyAr72KuHNL9Iwvzt0i2g4P2CS6nsoKnLfLSNMYy/
xzBSdTmV3GD1/hVFaNXO88oo0005ScNO68p8JRBs4oS5OI6g8DIr9Tac9/sOEqS5AsQvV+U/F92s
p6DK7jxOe3psNkL0CcPNRYnO6keBazWXBwaQPRtJ+9WNTIzhCW51DNGp4oVGZ0pfK1utve3LFcR7
cWySitnn/LJQ065ivxmYhSlsoco1TnQQ86J2FuTHaN3M6FAesQLq8zfIHtj8rzGknM5A52iTmN1m
s9s+KjKPhCMLFyZiN6H8+3JppCJ7wd/LMSLH79WE0MQ4VFPqZxSGudq8JaqnqYI2aaDsgMmbVLqp
4LS+v+9DAHMQ51oiqlL1ycljuHFyAROuGTKnu6nSoytnMp9v1JuhfnnVkzyZpdeJkBNb/ZffcNOc
G9pVfM44Zu6jx/W7LkmtzpWF8hRlTXvGWiWub/rDbb3QsGeURaVk13cAqxoI9K8MkC/JZNe3FdN1
Mm0BfWpr7oGn2hNJTr9wcC2RphipwDnjx85SYDoFEmwqHP/A5BwnQWPXW0x1z/bD5NyimIADX8gH
SWoserimCLR4pOrBP4rg0Nfw/ZBsYITROBTieK8Xc0icbpsFIbIBkbngz6UEnhcHSlqP6drH+FVS
0yy8CfNrygEmTehFKnmuM+qnc/AAZHk3lPliSgPR5GjmelaL10xc9h3RytPaa5Z3nhJQgHbukCtq
ZFkEDvv7fUwCuPd+hG2yOOl0NYiD8dCSVx/VwTCshNJ7U/NfdWF0VXUng0rP6H5ukKyOlO4l/+SP
eCC3CFKqCBh95eNtHR6Zc7K+wDnJVyjQBmgPfO6ttQn4F/8ZPY4rQ4FBzouxVQm14x3u0I3/Wvpw
xd50a8zk72v15cMBZo219hGSoPGMgVYZpl7AniJHdgZXnsvF/gl2ToCS4tUc94N6C2NSMM6pIrDH
iRay92GDM3pu2W7r8aUOAB7I8tZ490USVQAgIvVYrdniH+gdX1aPjIxT3dEJXnkjaMASgpJcfVml
+0C4beb2W0k1+9+O8p+MWdB1VddxKaNQqslAPqM9FrVAh3O/0PXKMvOuc6+dXo1vAzpME8ggY8TF
kZs1hTogDHZY1dnoijgS/hUlXVVouAdtkBOdQeDZ9RZwo/i/M1B+YBC390cF1mznJiDo04AtOaQl
UcvEh+1TehsgQMWP15nWdKZkxnK6gyQp4Cc2SVyKm8k0tUHZcSC6MCHc54Pa1bKhIdapib3VVbsf
d/5pg5pktR78j15LP81UB+PbENXn9RQ8BVENjkxwrX7CYAF4MCSSuyfpmEE4Q/ylJ78+3c5fgqIa
dUABDwmFGu/I5+OKNFvPiHSrR0+nVcP5zRCiIdQaxCpGr03DoE8hGY1GNnT+LJUrh1DT55oG4IpS
/OMIWES8iI4+sgzT3cj73633qWAU0T0BsqpK53HoGs1//Wjns98UIFXl7Kf8XAzX2mTCAYypo6mq
OtcLlbfPDV/n7naqBqoxqva8i+PltxGGXZ6MRuNSy8OQzX0BjudPXk+G2NhbeYTScnW3W8fZ6pmy
LhdL2TBuS2yxdZTDVEvsnrnQ3MQutounQok8LLdPfKxLVJEFzyjyrZY3qFgbAuuIPCbRaCeNvyAY
2vmOyTGxvKFq/hxgm9Sge5Cwq5aM62OFvrbTPuDpm6Axhj1dKlJ/y6FtR5q+oi6PGHZwtxwAm6+F
IF0B1EjtiKc8IPijhp49xr/mx0JN+MMe9c/mbyiqfeQ/rkNsT1F53nm3LPrweSPAO3wZh2R2m6u0
y/6008/pi4TsZKplxr92Cloby87XIrZv5yKmp9n6pXI16BC0lG3SExn9ngb2wHgwn781pWHKIS0P
0+1hZg93MkMlz2vrQU95IB5vFY8AQXsGM/jucmASiGZb1iyx+xLCxyxQlYW5g9Woat/X9/vbzFIO
SbnG56LlCkefnCSHPCekVV5nFgkWi9tZRGffoa9/drX6L5Iy9LMukt29zaesp0n7o8dWap5+OgH+
kA9than1I+eOhbCuJ5ULqeXUjVSeIpw/wcjAQATRv0wi3o6zyW9qPJpunPiJkg/jkYHIe8UqzK26
Xpj0SPK75KfteemlBUPGMjM04JuC1XkbVwI4hWCoByArHC4zJpSv9FtMPJRg6h4E3FzsIFxCqSwW
h9T+XDCVVl65IEK6LycOXYqsxOKSkvSimcTRmdMvRS/KJPx/n8xXvGtrPJ3dNjHY6l7yAf7bjaYD
Mq7bV1ExTX9UzS3EcQ4/dR8uk22BoFG7GX1PrCsSBL8Kutbhu58BeoIti5irVQJmO0NS6cdYLXJR
3ew1yeiApaSaZvsPQvIvuWwW3RorOgCUvHuuJ0MhtRLSYW1UY245HWITkOQUFBPEAlMKoVfgOQp+
ct48ZjobrmCQlp3r6bsqYbXb287DTipAKKrQ8kbrgoey3lqnW79DfvnMG1jMtNN+U05DVGsmNzK/
+oTkRwcyC1G6Hy4B9n3MF7+tBXWf5sdmZ+fCAP2MxBnkC2Ind4xzSPJQ9FPT1blsy2CPUxQ2XOaD
XZcBwjYbtSrULHNgIDptYEGMNWAk7tDhkNj63VqiWrMlWqFuXWyQB1FgRqotuSyTgUCGfwWdSIxM
RFJ/TQQYftTrvX7e/93jVHcJUOrKChqTY+tUiTKTofI3mOGbWWfvpOGLw8O1lZ1g1UZCvKPM49eu
Tyj8psHUVFniURuxxG7wU479z2eUFqfeLWLpasjhRagI0wTM7q+1RitAHkYzRO2h7bKwkvzDSw9O
8Agew1W2zllDKmez9eKNLoUAWAgS45nRGgQkCyvV2EJmo/sM4XbyiOOJv3LJRQcmR8EokjiE97Qh
Xp3CslffVA0wL/ftCPqk6qoshY+NS5J30boVNVYe7egnXzM7FpLTjK0NxV4MJ5eS2X+p6lqpl92r
hC+fubPy39LG+nkuhvLUhiJnqQ+h9/Pg7Otumy6YBya6DWrRPfySHDpAXiE6FKNtAQ7pv1gVSFjt
HNZVSEGMt7CgoQpcQScMgeDWQIYZ8mmIk9tt0OlMFtG4fMdrwl+mdLCyiV4OI36n10TnoJImE/Gv
66q3dKhN6gMjXvlpnLDeOZRCMy4Xh2nVb1t8kDHlm12nI3LzJQ1EBIpxEWqre81UrjGPqEe09NKy
Yhqd0aANsSefB1geBjbNaJrs03gFnEyDHTjt+/ccjAOlqnYgrfhJ/wD4bO7R1t9vpqXh5QzX3BAe
TKBJlbDNVsQSWqOVKdY2QhQX4SDKduG4reeV0rOJ4ifPaCOVjvcLwGwUrA1nHn45XwIUvDiDtR3W
NRAaeiGBw+x6ehMdXYQsyaLSIlMc7/ngreCQNlUKhY0wRAVQAEQvwC5v+5H3LzzIqr2d6cmxp5+f
V7N9VwoOdMvGiryC2RiLVDaBlvIj+JZG+03itoWaqC6/28nbbWY8blC+uh1KC/MIDXwKtbOqPbmm
nPa3mUB40n9n6fibLhr9qNldIeuE0xoy2b5uveN+L4koZ3wRYpoY5tsMlnfzzTzSKJvYqaQpT6BI
B/xd2P5u1pjiFLJ9eOz/oV6frS3EINBr7y7LfLNjcFjk4A+YuKyhzmwaka+vobCKLqdlTcYONS3P
g9M6BqGdoZfWHprGqex6dy9kQPU9iO3wohXfbX7DpeX98lo9nuNcswO9qeY+g9yM4S77pHDlCf2g
jaksYie6T+HD4yQduOlEWyaUcfKaYWvqE2NPjtKTJhQzYguf8ngcAEHWi3ohX6PJ1FK5/b0oXF1O
tUeJQ04Po2eTTfRhb19VPAqLrD2ux9P+C2VoDgdzcSeJ/oA1snJQuzrBAVXSu8oinbZJt3PKr9sM
v8QjFDJbfJmbig86LT2V0XpgzDuAO2GEUsZsNM8jhfLCxDuho80Hn8YRVIc8KYeDHAVxw1ZrVR9x
xbRX7Zd93+SyPUciVHJRXQc9hqbD7X4GYHQNiT3xrRmoH1Jdtq+UXh6fURpBE5P/9XDKre8uBuzU
3319owBG1K/8Iww+Z01jR4+ARdAoDygaY5OPiPfxs+goLfCDYQvxHvTQsRm1NOwUW9cbkwCLSYLr
hrxPHUx9TlCfsMzHHjUQByNktAbGSHncl5F0ioBW7MUn/ID6TqZsUFB4wExW+eB2ELjQUrezr7Bk
Lg+0zfCkKU9itCocK4WpE1XgGif2CftFnpdDcXvqrHJ/hvDMgWN3OAlGIqcKTlkSG8cGAv6MQyXR
8g4O/NhWbGzCqp0+J8oFqjF/ymEDdykA2D91VrUtqyVYC3jL9quOhX6VDe9Cd9iUHTKWR+v4YPKd
Vd5garktmF1FP64BQamGBIdPZ1XItfn5if04AhDWSVAr5/vkj0VygA/MlRLbJbzWpS1CKtADIha4
NNgFmE/e5A6wO+aJGtsnOqf0mOuTYUnXeWubBb+U/KxMe4qF6yLQqA7usrIWhhslBTIF5dMzxjg0
uRWyqFjCokJcKrKhHj4krimnXiBS5qgex514bJdeS1CS2Ambt7r3dAypWRMwBR9DIjMxm9LH8nGh
6KtxZm0Yg67NeSRwsEL8HS9yCMEHXX11lmsZ2NJEOU5EyySxly4AQFsWPbeyioGb622NIMR6xYXa
N67TYcNmLoLsMMGrH/UaLIojJL1BosxsNR9OqTpSmAivzUzRL4xYfoaNQ0Hq9rChiNcJmDdrAk6z
2ziot2pLlEPeJNkDpKNhEpZU37DDvjOf77LTVpZPnF7NKpMgLUHQm7qDoS27CP+hBbJw6Et8m9ib
BMougNzBWpITN1M7c3tsQbgvM1ITUq6zDjxH08RwodokwDvCZjGDEkm3Y7ObSzsMPNCpIYYH3tjX
DvNrkQwMXGO1nMt5OLPP1dSnmOBxkQW9d267+UcX8PblOhCpwF0cXHhM+u6f4qA/9tMb5LHxXPql
+QNvxdq5vhU3JwLQZXsQmDdnO/TuCKo8UDEvupOvuhf9zFxfXOMyTD26DRf9XNfgrX1FI2B/KN78
tg/chd1INZmhMaOQF/XyEpgZDxx6p4Tx/D1IXRCOMgYUicrq3ydNOIy5jj2tnWZXyACKYkIrNKOJ
iOLx3IhI5kwaMjKxD54X1oygNY3A78jZbFdLknSreHbhnsKEO3pUYMuWf9VGsEHqdd+/YMH7xHzM
d1i0JRbqypKC+C2RJ0UBPrYOapg5EC8Wsmzrr59MGCqy+tn+uU/npREYgDTyPwWJxh5420mEN9rz
Vh20lu/zkMQ2JHCFh+ehlVNgWz7OKKFIwt+kA3b0xuZbGNmHeVLmDU3sKOsiI4QwOxvugUmbsVKx
tESNv1YO2l8yUBgBljsHgflR0Ob+1WWcJcrVQ4z+wp4nUvWghSbmzZLOV1jNWH+s9uOJJUQY/UhV
/A6VbZq67ZZo84cCFV+IDx25l37UOz9fortCvPcezSYBTRy417KL6OmRGq5qw8/n14SunlBgUwI4
ojLKpHuIql6kRXTETl65E5NIywNqiBI6PwpDyKztlQW8YfC3kYYY0kutjCB5MKOoB3cAyZx5dp47
Ljk7go1EhHclYkJY3yHyURz4lMzceRY8m+I7sjmWfY72Zt1awbaBz7AMXDh+hGJCIErp01O76nkp
T0TVsj5XHTrj7ifpeiaW6vy5I2EZttyhrleshaaI7YvnIajwowekGZYP9Ri6cGvCj2TcqrRqt75O
NaReEzFUgzUZSOaQ4KgOyJ9toqzY8NL3T+IkeEzPNjWvcRuVcc85hLLJEgnL+xLXwahtuxT2Q9i+
agYnpMZYEyvBz+2RYoBa7IerIdHxSMoIjprTRsNrNS23T4KVguWAbOfD078EYb5Ug3a1Yu6CV4XS
Qx20IglWognNxTU4p6CQGBY9db5Ki9P99sa4IgPmqanYELGsTNUQuQOHFsAxMYqTIVRS52CEhB1U
PdocyqnR0SWfTqjCnuWHU2TTfNUiMevCWimgtVMpRirwKrFCF92l9spm7j8foma/8wCG4MP/KvZw
QpQi9P2+iry4jImcld+2gatB/qoy5yFmwmUMLlRrFcofFlBo91tCA31HqFDBIbXIVK2H3Z/YYznB
O/W5AL/sR3dyKG+greosa3TzemeqzLxA5LQmIHaSmVqIeb0re1EnORcti5XZARz1CK8uWcf/yZ0o
uCZYElU98ZYbb/SxPqAg6/OReoDIJLIEFwisQ/hlVqh9KW3XnoA3GCc+W3twe8SJpfKdds6rd98U
nIPAWqIhv9/R0CmSoLft3uIzjgg448iEimu1UHl+YQBbzBLLAULaqxhw0ZPIY0vCa7Nu1qxMC/IR
52kIqXtngYEOu67/rvt04LyJtv0EuF+KdWOvMUxWYnp4as9HOVc9RDvMJJOaoZ+IY7SpfGQavOL5
X7SpGi+5g6txVZK+IqHaY4/f/5H1m1Q1dnPX9WTVUN3ER7p/G6OQORHNPUYoCW980G7m/cihm9xy
1t6W9yR4v7ZjnzxrL0t52gqXl4dtflZKT6lvxsXmCoLXSatMbDhnhNBRA5X6iMML3ZNlXYeMxYuD
EmExtHC+ZMZ9Nj9iwJ96spoZnO5D2UKmJ7DqyhNyLQe5pLC+n4dPNo1OWLOlG2vgZ8/YECKW+ixi
tZj9b/kUPh4CXziStdwWFYp0A3kPH5tj2QrXLvqHFOZDjpVR5hKc1fndDpWtpIJfD38wbl0GTcNi
xbLPbeeK29zTKBDNbOYCwXhlQ7nHlCaIHQsXL0gS99dSP8q/rXeI3xTlrX57Pksiv+L4oahXJP6k
NBtANmg6/wGpZLCoKzPGLN0VbJxrLnTW/WwVtX6X2OGZBuPAn8hP3ovE9Yi4vIIVh9mMejB773aA
e5EGMsNsL6QLtCrXVTIwXsiXHjuBJptsDmnP4jkYtuLqaGvYkBGJ9ip4M122npUxFCI1Cgo5XjoQ
0zVLS5XuoxTmZ/zGTyOX7ZFTCHzA7WPCLt50l2RY2tGSG98Rd1EzSfAYi1wzIcn1olKiVeQ/DiUx
6o651ZFsu/s58t3wuiinbu/WgRLj075PXwxbn4gIM0tiG17M7F+YImeGCmnxsWSXDYhuV8GsMwmK
FJbtiXWNWTQi8TxDi4m3vAhF1c5Y16oV/f//55t2tShQw5puJExParEaERFQUAZnxCUaNLk5SXJt
QykZu5ys6It/nKXEaZ57tE4gt2naGhd01OZU9ECC3FRq3YiA9Rs3tC2cBkyO6FQCm7KCRj3cOzap
yHGbm3p4TuxV2ceL7g6Kbqom70dpn2YitOv1/vgd8iUcQ00wGZnOnCOaesdmFP1c8BFRKD5X6YeJ
Bkmd0bowKxtRRmp8U6Qc/k1vQ7jKhE4Rn5TMYZR7SupH2h2mTFLgteZ2/FkUUZ81z2Rkm6icW34E
Mr3hflbfzDaiiKSwsf2VcBkjxoiCnF0q7aPmvqrZYX9dgelYltlPWukla+tusQ1ajUOjcK55orhZ
WHXeS2lkQEyKZgWzPQjuSmeaczE10s/gU7m/QGZtuD5aVwbm1Ozvr2Zwy4ha+KFWB4qxUlGXEu6f
n7DA8evH1Ig/sw1/GGEE/S18kEgdVLbjhgrIYlrdKOw5TjahkxcdvyX5BGqwch8TjKwbxfO+ImxJ
MSrL3tzQRff7ANYLyvhHGjYNwqZB6lPnr6oxEh/9LdUSyvnLtEa5g4Tfdq7GGFi+/COH8aiAod13
fen/FGZAUDBozC5W+YNVRCXgAvggbiBbaS7tRUTp6efu4kr8sV08B3pWwYlRekJl5ysX1lisyiiq
CRUeln6c3AvwEgof6rlJGnQwaW2gLygX6Tkbk/oDWJ+4OSgI4jtAF3upybBCzeAKFCtFxAqTWI2L
GX16CHBL+dYGJF7ro/wdsaD1Mv19TSsvag5RX0hC5z7puRAWJm2rytAHWcMb73aWbIrg4T8hPiQM
z4ju4gQSBbSW0QZMR6qil/PAvOGGWYX93v1ug93ie1H7zNB2bjnJ7vR1/IGeVxbSUb179am4pa1+
eNC64q0PFS4oOIrWOI+Riq2OdC0gPwU0nCQDChJUQfP5oyjIqUg/yLTzR0wkW4vl5dDgzi5kExzf
78aeUDW/cGti8irG+mw5bpL18NOxsr2uz8ZgUULNqDY+cVrQ+PYyN+2htPFVmua92zQuqRjohAyh
nnCDyvEmRvDOW0BmtNTM8u/n02J+bGJ1ao/o3ymsPsVqqhAXtw/eydvQis9mQGNBcVUcraHEPCYS
UJJKJiUNdvQfgrbjVnkkFwev3vWIeh+ooduqdTp4745D3IepDfddbVzrsaQrlIH4CzXsFRCKEDxy
L6OJbcGSmX8k14mRJas1srZFOOhFdtA2dLi1dL1QFSwF9FvXOeHo+u5R55pn0Vq5rZuByH6tu8Zb
5sAJtVWhuXMZZnzPWY/VjlfeTxO1+tSr835p2XYZFnRk9aHvKR+yeUiXAHMy+5lLES6OdupYO09R
M718qOWZvXGlLNbW6q3dtkhg1VNJeGGLtfDA7mhLujmuigWoZnNOZqggeD6yh9r3V3FJ3c9vXoTS
hmbJDaKcVnraObRQR9D/D49Cu89DpjU1zis04IUQ5h+WuT9FsaeKfJckLd/mwN/KWjSxf+6w2bTI
go9x/piF0cazaRBUKJYFxWlSaYwoJ8BjN+w4H7Ut7ZazBdad4PRrVRgcGutLGbIDy+MAv/++RCyU
k/p9RoIz64meM/AAzhBof2pcYsCDZYn+cEAXXN9f6l99sT9t8Eztv/WRczHUTcLxxGiSQtY6DC+V
XYl5/NKG5ASTYXiSQD6T5EuHZChl7DUZ837ETZGoNSHHRf6kEIWKNgMUwP8yFr2dV7mCyXjrLdYD
2xf1+pc1HCnV1BkCbeysLqFWsIgv1OYOGBafFf1cQ9EIxGYTpy7q7NoCQT9LVjq3E16qRudfJ78r
CsAEpApNBeoqOS6uhMLv/jwJVvhzB0gUqcTCIIbp/2KSgi6Y5lFXItTlHmfsTk2FlZKltU+9u8R5
CDYcn7+Q+KSfmzw5A/wZwWa7Oh3qiLozlWw0cNJUOv70HFV2RR4KBy4J77D9bw2nLk/o5c+qk8Kp
BE4lLX54nCyWE8xFLWIrYKvWdprXyjBxoeaI4L5ujBRkBnwBsuFqtc87tzAWG5x2bZAx4VMm7SqS
jxsDskezzwZzFYtQs7ttCgcyy81VmFzi8YaWll7IrSp3ujLWUYdFkvAmuEkpj0lADe7lSwKnTEqv
j0JelFmO5VTrazeP9RYn44k/Z86H0eljLkJMJEiayyyQ2smM97shNk2snSbJgYOPmSXwWz5Uq5Uh
XuNbXw4riwcRAMHn4Z0wSyp7sHqznUxFi1PJ9O0efml3ISsEQMJi8brU1yHmt53x9xKqnwrRpZnk
lNs9eH5TYAsJreIZ8nHuW+LFJoq1QMofcsM8D5hRGKfJPrsgRG3bTDJttIl36/WPLVABeflgf3+w
52gxI2xDIu2NmrviW33AePRyBl6JCNyBiN5TmGLfurfPV3AclofdrJB3L4gWTajf3x4I77j+cDMz
QJZoDhxWhTpwrV3zyH1lFDr/hzF4bmw1HgZfbdhcoCe01DLidBTny9GSTUElMRIXkCd9KYa0q+eO
mfT33uQojro9exeBC4tY+isKgRihFHWb6aSCdGrZoRJsW5HFtLxtE/LrI+FwQ2JtUgjNBfSvFgM3
c27MtGDO4BcOVF8RjJbp02OFHqyDx+btuedTscqmnHHlIwOrC2d2MAIga0/LcPC3UIIJLMQiZTq+
n7ArlgpzwbBb7+QKQ/TowCz+iZJkzNPY6SKU7OjLZjsaLyXVILUj43iNQ0XnT1ZNtNlkyHQ/JmYB
cTeLN1gXT/no07aaNUv1tQhvexvlBmxDNmjhVVW8iHCk9kW7mcN+18oeGVjh8nVDBjXkrJpEATZU
F6+qrAcEQbccoTMvnd9lVUjee2fsPDIj0JH7m/YRAMPVrMU3zcbFyKYQLzzBSbryaH8cbWtKH9Jy
iz1i0wHJ5aGzFv11qm3MtV1TsZ4U+0Pq12GGkaaT1y5vg8W4IIc5lXzJIDvASgIqIVvDPY2ZiCFI
25zGE4Covt91FQiL8/MxnsusPsf7QDF+YUrm2wUgvmelAubIm9KxU8T2AOiAUrE8feCV5HIICVgY
vHUeCKvq+qRM8iW0G1NOH+GMpA1xx3kDkGAa9FAm30RQWPa08vdCOs9FvF60CCWOM1PR1YV/hsB9
8mNpj2zMzmUK8HfPE6qynfavoRNcQ8C1qrsFoBmb2BBi5++KRFdffiufv2JOWia3hdS/1xrTkN5W
T3E7YNLed4sXPbQ1UU5HiZoAE95oHxYDAg5wCgpI/97qX3Y2OfAge8pCf9YpBFLkf+NBhvlvwAcS
pN7MPXeq7JVqpR3PjNWS2Qtu5+RNQVBKiwVqup2VAmbG7aZPGNKQcCZ+a18z8q7dDBQ74otDAnvF
dqHNHL64o3KI7HBoOTTQ6UnSQzrqnOr4JDxZVSORwVRZbSwn0zx6Sf92TP/ENivh9mteVQ/LkKp3
Y5E8yq+1Jwc9N4CNhXfEhkLPeELaG5digvUVJvSzccQykr/RdTLC3gt6RYMmpevvMBRQmJU4fXNs
dBZ/AsXIT4HNqaT1COyIatj4DV6lGj+2EJkU0l/t0kdhtO5XU3n4EEcvI6klHfHkw1HrM3FFIbJr
tjyPpgR7s9fXX0z8G7zB6iwog96mZOAPB57UNVxSlh7A4U3nnDNEx8AghBxXHDFYWSkXl78XPySu
9cYOD7psfMExvZg55Wgtwi1Ew0xOLlKtJD/neN/sZI+boHviVuYoHNs5rQIst6YsCdWN66UtDqcg
hTaWC+SsI11EUZfzklf1oGqe+zZ8OJdtYTKzh6kiwNsnZtqRdlcDQ5BOI8OoYkWP0yOwKzMI2abR
/rj7Rc817HqzvFz7SAk+zYNiE7AiIGmGP04vv4q42kUS6btRJtGE7MeEWFW6UT2uIdhMjX4Iu9+y
Tb0NC0EAZ+jopX3rqurava4LaVK5PpQ1sIvoYFMrVI5hvIeOS/K7eDXSGYNXgNhMLFjDc/vcdguE
Vmg3ydfsg4baecFjeBHyt02pAWKWfuARQChe9okSEBqHwgDNWUhxJt2saIKJKbfGeSG4f8IEwQr8
3SjgpLuweMH2cDA22osLc79J+2T46n03HJwZ90a6UPiUr1WYrtITbWByeoF4UvpRfKmimUhD2PPv
GSQUgSkZMRYICgbk285zr9t4Tptd9YXkNzPfdOtD3x9ltn748QxckXFK2of7uV6zU2I7xTHUq+W3
85wi8EcLg+XxQjLI5sZsbgu3lSQCwrRlbqCW4xP2lkJzuQ4bRSrBXMqiI6+Mh99oeiGjgKuNepGL
dPnXNc9UzhPjmkxWGUwwbuCD4z+VooOjHi6QilVt+x8is0F2Rm1ntSTolCJaiOweGelg6yVwfpD6
OnmelV8Y9Lff2rCUnVD/r7dAvvICbCxKOWTlJJOdkcvorJNpO+oU1upwUWGeSseIXi1sdNOwwi0P
HAt/e8D/WnalHhGBIzOuA+Bagz5AmB3dPZiEc2fI/cZQtoooXXr+4aKbrBWIYQsXD1jIp1TTpu9/
RJuso6nY4feC+Prwd/oCXuow3Jer4X1/p8/qQj/nJo5oPnxN+RtEosjhEuKPdpeIkqkYle26EKZX
ZLg1y9sOwcwiKH7E2D93oTRf1YfJ0qqvckUA1FvLLs+IWQNR5aEPhD5DYJiadq0EoEiqWrJfrlkB
ipnGKemz7PZzaRVU/6/UzN2NOlfdim5fjgDY7lzk4tZfWwoU+XKFvB+XAM3ryJbOMimtH+ANq6Z+
oUJKJfPq3bSNprOuagwI5OE+eRea8bIlMbUOZjnac1X1wZSEeUgmhkYXh7FcA0RifiMpZh/+bI2y
THcQubqJgbt/yUvxX93nEbubAYNVRuyB54aAVe/xrqHIRUwwJCMnna+pTTyU8mDX5nLAV+LJwBb+
KnKDOV86VsnCMW+c75KlIaTC4JSZ71DcsWlZBHjhlrmYYASloCdBSd2GRihUADz9V4sy4WVrtQu/
uiPZ782jgiUo5SjbgR3Dq/Jk8VwggQK4b58M/7bJyqX2M+DCoTcXVJ4bdP9/9N/3NFOSyMdm13JX
zWo0nS5hZ695wgnKxVs4fn4K5KHYjkzGCKmcH/nKA/+uDkOCl53vgFZuqn9bpLJWXubdG2Tx8lLv
prEadFhQqtFixAKxP59fsFmoVB9Z1f/X6QmOMl36n9X7Werryll7FX72iFPrbkZGQNWvNsQQ2q2o
pBo6FwCOHCKKcVjHTS/72yAzpP/+hROeJK7v6MK5Pve1uJdmeQ5VTBZh1PWIY94/oY/7DwWw5tdt
EHO1b/tffGu8JiMLR7iWQRwbpz6fPRUgadpPFg/+v61c4Ve5WKVAWSOZRCwkCFqH4W+8McGQyJbi
bx5lkX5i4gz7y/rZPV0Wk6J7tHyZV30PGBKgIZHKTdmnSpU02iFF4L7F0B22dG/076DOiaCMj/1X
sUUVLnmnG65lmgR/ghbp/MKl2V76ioaWPbNecgHrInYuvYKnK9L4MtaF7cT4a2jSQX5nuTZULR3j
1bo+OpEGn6SJL6UkF3qu9r5+pNvf8U3F8Vzq+uKwUOcHkTRW07sIUnuxO2WG7D2HVga2ETmufP7G
BTGrsx13lPX9IvFr5O5CO+m4MRJsE9oSan5q0Kh71kiTPCXeuomh9e/2Oz4RZkHY438OrpR52jvx
WLhvmppAvOmD5cdKtrEDRGSjOs2JJJqYie964Jg9EqNLTOjTFFm8xQLvLzohdSdChLo9jnKsbLXT
H21AIRKmqXzxX2csOcNwuY6OlnrtluDQO5V6W4a+qJSF7/4HcbkAipFDoFns0xVEKkdTXShR65OS
po1O/eRCMalNbPsxg4Lvto2h5vJLMp7Lf+Iu8kJvLS0ugX26J4IE/KMizSTtSoichHlD2YDMm3Af
S8QQP2HYgTfUcjYcv/+IpcK/SBV+mDFgc3L5Fp4IIL/1K1IYvUyth0X4MBAhc0ykshf/p9Ecbrk3
J59JZ2K0QKrKuG9gx5sXEhN87Jn/RjZEfh6Gw7QppG4I4MTtnVgjuLPEIf9QWcxAQ0APOs6h/A9Q
FFlknTHeKMe1R/k+dJJofSF+2SFnm5AL5dvZ/DkeH9JDcL8gkk7FezCaDGpIUC2rKh6se1G7GFId
rs0ZmlIHQuIz8tysLIniDPufYANwHePlBoAlfmbHjtkUj2z3DuyIJL4zD4DzHYxQlZoeXEKKMj20
40xvxfx1WnjR3eOrrHGK5PV1179p7Vuqx6laeFLjq9u+8OJg0/HUnvqr0mXS9mFh9kC/YQUKPc8d
A+svBhoJSY/myx/vZ8fv3K1taTAAwLje1HTQSTwgPfZB680PYO5B2t8vA/x4Nuov/MnALwUPpmoB
3Px3YcrgsylSPuL7DanAgQemHbBj/aQVw7AZ22vJI8KgGLWAQQhD8I+pw8YRQjuhQ2VtUgrHNa/b
DXCqepY2EyKPw7AllSUBEmVtboa76Ti5NnU2Yqq8SuFyYaZDA4NynYjZoWRid1DloVlxsVex4OwF
fjptmWwCoAzGA/lgeyfX9c9RetqpYz3wIn5k90BNlr+twnscOizPKWUBrSJJE4q68tsVOGSWp9i+
fJ6DWMiV5O0xAu9bkf3L1lY+0f5COUiv/kzEBO+FcJ6fVetgKzZZYM4LxHCdLTCUz5Thsqi6BqTV
IcQPLwMixVJymGjO1gYsDqvTsBQibDsq4O/AwSosyS1NE5HvubF+IbAK/sMVGDY3cwkIitRnMpLq
pOm6AybAQk4FQiwlz5oqmxG5klUGIy3asophnp9w959uXTQYF8gMEHaX3kqmYWU1E2Z9pjpUl808
Ee9yNH9TsDYMu6Z80OZNggJzASU6+wy1SVwTT/+uphTvSx1ZJhTtggF+h5gKX5XTOBd5gxXvpPj8
XztPuFMc0oYkddqQ2d5Jpqb5/JTVUIzDlZ/wreNTdP/SWzfAvg7Rob4R/AB+Nww6osc4KRsLFUwS
l3EIZL9AbXZ0TXfWCCh9sLaxAm2rfxBZE3gPReZMNd5ny93CV+BnIkJ0Ah5s6xEm+QrBgGKcO2yO
e6Mkt3z3YbHqCMGRdYyKgD6kH/PjAVKNfZo47M2vI1e3meaP4OKBW/Ulq/38+gb5qVCYGnfetaeL
gTt4faK3hwNeiT5utAyQMrylfUy7uZ6L9M+Z6F4a+bHsMVQR9amT6T5dS5j/bQXtt4OxYtwlOMTT
TiOIruYFxH/GEtnyaAUaBKj0XJp6uN8BIffRFLxjyMUzoz+2w0DPve5bIDVnS6UtRKltimuNbfK0
VtR3YpCvibwoN/QxwxqksFjTD4mm3Ihrduwbkpo7p+njy7RHF5i/O6nG+7jt63ZM68+ARcAX+BFb
q0TQS95YBuXZGB9fXbvYBiva9y/6CKxEOI99vofWChs+CxKJa8wnAvF+ORNEAyRY0PZ0skZfCUSO
7PaXmdo9XISD5bL6GvbP3vSIcmwHLKjSUtBzjvUn4fI+mRrxkD6/6wGWmAOZFyFyPF8aV38sy+Uv
B3uoQArfPw+yR10rn0DtMt8P6E3sR+6/mz8YrLJlO/LD9nvWwD7nwm513PDnFHMi5NH/6EMK1Wuz
yBvdm3DpaA0+Sql6gn0ej6Judr/4q8Cbau9kBfRci6kaNQwueW75ksqKlm6E6Rw9svVf1XvhUMYt
Hxb3N7DBSLEw4eZ+kJ2NEwzAVYj7mSvMVEBBMG5aH3iQ6y4ECIB3nZ4QZL1fR//ESScX0TxgM9aV
Wk4bV5MvsvdXujcgZshBysELlaWdFQHXZvqQiB6iCaPrr+25Wui7b1r0z+TkAxAPRw8yJeeEh3KZ
tIy0XLvkHSmlI39C+Kzgmq6TbS/eTDdFPUgFOROy4CW9Uh/U3kwUwr45YkOfyJBYkA2Ka6VABKmE
9ftKsbFHibA65Ljm9W+9d1goGEqRMq3LrgalUH//da2l68zSy6IL44DjhE0JVEcY3F/Oo0KrSg+d
i2EZF6iJmw1SSBW/M1W9Urlly5zl5Z7JdpGx6DDbopLxCVenXJ7RG/LPqp28T4cNhUL/tkJ2AHHj
6O6BN7z4J1xxPEE4tA2cpoRlgmbLdPpgTzMX6LuKU1EUaxG7IYYss93hZUMgkad6JU72aLk4ErDB
9g9Rgnx9oVxoMYH1hgXp2z9xASb4DnyINAVTuUSmshCpV8qHfVTiq26CM2H5+o3ESxEo/wPwol9V
qaWu/3S74hM9+zyssiug/UjWD5fOEFP97DDyDoWfaL2C+0bPD9MD8PqtuQFVF+ex0fXFfSK1qMSX
kWZQwAnsxvbKVWmWH4HBr9AHelBw9dKS38XUhXhKvkjbw4XVMq4M0cA+R1t6VYWpGRoL1hpn6aGJ
bM8pwOf1dLqRdqIg3xYwehroPhMJbF6FLcnqUjwUnCu1+cxn2EWranToeiisCxGNe68a/xRnTmjx
TQ+G85v6MDhxnm03ySTYY/AzNzrdTdkLL9ZNdAHQrMWh4i7brkl3Y8mLovg9+gpygNpx+NoK2WDP
uTulY1lwGTVUhn7G558SoQulfaU5v9usiZENq1nTecmpGRDfdjRRkvJQcUThx1w91tQxX6UP4vCt
O74pxnjzx/Mj9ZX2QfKmDoKKt7RGmP8l8P4Hu4Wqq5HXuqsio2T128aqIpDlbUMZEgZ9evpAdwx3
IUHYqlE4NqEzFxQfySZXAhwSgSqKu40JE1SZBaJXmkXf9M2IaljpXWh216KoaGv41fD4GxxhJ7aJ
O1giwe66/sv8hX1H+qH7A5JZde5GOZSXdv6lDdpSfyyMNleGGHBuPbkesU8h06+o7DBjI5iV7tcd
qZFgOf3jjVV+6XNMI1FmAvTtzc7PQ/1JQLxpLbZaysiH3EOzo2yWMtqOZkvkKtwhBm+ioXg+isOo
BqRzugC8gwzG1368YyojnGVxA/O4pla4bvN5V9KHnTM0px9RbdYoiKc98GRg9YEK+osV2OsTzZuz
Oo7pm4nFI21Ae8bqWMy26JbR9DhXAX0UOPPxj26qDg23AYrSXvo9tBU2NpsLbFIeeQYkMavEV/YH
wZZkehgG90MmfybeleYt1Uq/0pCIEIRua7Bq3AfOMbc3CvteqBnDRf2gdq/1w6w5luxqB2l+EgSt
WmGeWSsDVI3tCdyNyLmz0+pTyeueiWRX90BwobzmJAOTIHxSE2WuHwJ9E9ydDzfBJ/aGUZlh18d5
4EZSjN8vs2Purpd+S+PTgq3Czd3k6fGptn1rrlSPcTvrlADusoPXs+CMOFvZDxSLqJGHy3rs9EW0
MV/Y3f1XRP59qMCLO+T5FfY9hZK8Si5DjwhFMeWaUBvyoEiMuFPdrarvP4jP5iIQZ788H5Jjl1uJ
fyxNt60pZdSjao7yGtTDa5ml7jXgVt4O3q6AUbVzbuMNPjX+uKJheCqMgDG1Guix2jUmb3a137KH
C8Jm/Py/PTmqaG/sAIlkzPnJQB5oEoFVE47+GQm9pBPf9uMRinUv4rwHmZv6j2QNdJ4BgGT3IUY/
wv78+/H6vrkY5utWS1PBM3seve8f1/QVRUykOE526/Rsd72PqfBRmaEqGsZY/6gBZJZfiky8MQJo
G1V2Din2mibJOicMyDvciKYSV2QSynhRiUM/XxXW3Vmu1zL/aUrdt3lIC7A01V92ACyZcSRZX0tF
/GI0EzAbm6c98UzUBGdArfo924T57zygg3kR1PnOJ5D0jlMefamkJK5gHCZu47cOq0JBP+CoSRes
8Q1+mMsdaYAi8J49a0uTkX4+t4VLl1PWB4v+JPIbH3UrP4vP4vCW9vzzKFTXbKAgM9qeais8lXpj
W4lr+3vbN6ev7NxH1FcWCZXMpYzKs0ZN0RqMpM+k68yX+n/JSoq1DfnCiADLHDp4GJQmfhWhkHjx
h0R0RwcgWjXc0rPIb/XqNicJdns5lYKNJR9NjcDM1hxBI+jKCmd2o2We7kLTz4i6H9LOS12jvfJ7
CKBMRC4Flh2TYHrtlMYTtLCO14ZgPqEMagAKtLu8eKu4TEHo9SOsTl4Pj7HttZe+xjp6tpl8DLSY
tTVMVjx2zXNP5kJmKn8jH48k3ebSv+yW3o7IiXlAoYlxzfo4s2RILFtMHyUt33IeyvBx7LC7kAvC
zCn7f5vbyuw+CBaUca9QCRy5G1Mif82qveRVHMHLHW68IhjY2lMpYJMDyup53PvaL9y8mgaEpF9B
gghvbRtRyrOlKAyduv9pAhbpWvTRzsqto4uMbXenQlSSB3jMdjjmDROD8R1kvYDbo1naTjxxZaj4
sp8hhlYdzHT2E8PxgjOuuTTmVIDN1N15Be5tO99jg5QKnJ61p866addvHAIrAF9EhIR9raCpmAqf
f+BYQd6V8+CS1K0tvqk+UEK4fIzsN7OxPMVFyQ5ogo5TutFTETIscjGcKI5gPayCOBgCsamBLy0q
eF9UGdEN6vtPBF4Hp3joa3kCk3BTt4nelb3rrX9wd/GKAlwMNQ5D4hlnYiKIsN3Up5jdVge/Vkp9
P0IeYAx1jK9V7LcTNyNMAdmdzYmEnCd8JICpq3xAQ3z7P2a6S65epBJEU+v/ubnLVvPvwd7naEV5
mqSebXgeaGJXSB5B7Sp5nd3wdTdOdL9KcQGn7bxNOH7C5OYyJRCoxFwNvzCOUElc1+ZBBm3pPOai
X9WXK45nxeoUk6V0ACwsPiqFtfQS1w+shPpqv1wtqaajIcIm5WUA2wEiqP4Xrze0ffGuYDF6qbJJ
bOG5CMitPdiTBdKSiYVxqc0AEdSb/SDWGJGaTj1mO09zDFmjNIUzX2NK8JV1wP2dpaMKunkWVOYH
vN9Nn/BrfRa6HqpBO0Wo7RAu+MKliX/ZFKJG3hsbBuUsjudaM3s8aXzKK7ZfcBRh9G3zo7nlFjAc
yQtdcqEST17E3m+gqJXkXAQhCW5lSib1u5+P26VT/mChMF6lNL44Me4JhP0bkrvzS6UkDwa0fKJ2
jP+M/VBEE26Qm9NjUxOEdT4HKw1w67eTa4QqwIsL8xE83hpFdzvV2PpKkTD4uggliSVAgL14b8PE
Mo4l668v8kQTo9eKHTn1qc2BkEi/3N4UW2mjXLCqUTtyEB/uffQr97DjVDtRmuD6VaoJVFGu+d2/
4DFGSkr5zNluQLgI4ExF+mMnzu+VYKRAPQwYEoPbKBj3WyWO+o6Z7hPi+6jk6htZT3RrmjJnOHie
2tnhIO5dHCE7JM1wbUe9D6z9oeErfijVKFUZEHKKClSaYPQUXvDx/YCkUDQMw9gpPWLWJFK5dEYZ
Snc7l+Kyr9OXjSMN7wupbMqpPwrc0PqsGEzEZ/g2ceWjlGx2bl/kEkChLgL56LPyzJmD9FW9LZ2a
+WuC035Dd62ipJyENS8TdTimAZ4YgHtwLZ/Jj7DM0zDRhtudUOwKduL3OlFrxRoKfUjPNIPpjesj
o6Pox/p4JhFRpK9hG0bnpL9N/W2Ka3BysVebBgJQRomrZt2M7L+6kccYRm4gGVWZTE+U5cpadUn0
/UuI14rnxohhW8yD0HDRF7GIefPzIw/wLstWRkhHL3UYXsn5xVAZA/jJE3qGuPMdMJbFYRmoOKYT
rWrGGY0znnqYpjuYkxUfeFyiKbalfPbT5qHyzdnrAWHRtsIafUoHyEHutqgCYUpX/d/gV6z8j+/f
CaHfvrqf2MuNRrSJJj80YaZ9ilfn3ODYIERcgzLzLEZ+d1KVZr6x48FEWpPBpY1gDQQe8s/6pAJJ
fwyz6Pam+Tb4eGcVqDmeHxe8D/UmEZZN1umpbIqed6lOsOt48wViXKt3LDJopZsN6dhaYb/JAn3M
KkFCWUXCGL3hnxeVSAEeJdWH9N0ptY7k63xlsMVr/nMeHy8J75D2Y1sovrpx+Ad3x/P/mHZSc+k7
OHqq7N9ip2O3DUTsKXTWXmH0qm2AzSiATtwCwStc8+8zPZPehQC9kPRU3laq2MK/QCak1MyFmMZb
fRT7g+ZNVcRZ7GKbE4D/cMxp0PH1LvBAMYjfP79qJRz8XTGSWlqjK29QQtwRM4WC/IMu5mZrpdOB
5QTCFDDfPK9tbWSmDC8ggDIKRt5kC5pE9SKSVWFhgR8di3hlsPC1bAWAc0/tZgEKV3HHnukYFRJ5
HiShYWLVu63oer5VF7+283l1lTRw8CrBc5blxD4H56p70a4oBII1k4dMPMuUKGfI+b05a3yxdAds
5zrYtbXh0ZzVEKplN27XhFpwFpvCxkkjDA6rg6hyhzeZ+sYINqOkADTJn+QE475cllm3CW57H6s/
/f1orK3yQ8mr06DQl4lSpme7hP3GabaTgPP2uwLYHZt29XolB2A+GwsD/bSkOTYvG3vHxd21aTZQ
ihB1AgqRUeBuYDui2FTMLgaocplKL+LjsSndUm2PeZ3F2OKAPhhj8to8WffjhCRzc72nbDMPwfvw
3Id2X6MQFoY3MG/32evDUqfnjmCACp1ZzGce1oFfYAQ3zCzfrJl7dKijlGpDX7oggenUIsIRVjf0
4TkvZ7qoxOeR4qFX2SHXte8TdIqbcJ/L44y2VUTspxvqthQT2DwlOiHx7ZvPtCPwVMvx0Yj9ctRe
1UyYhazTVRkoabWplD+HG60wbqpSQY74jUBrDrv34tYbAir7Zbs1GUSuO7cRtG9dvSnMSeMXWAhk
DGI1TD/q5pZ+91Qx78dmya5p+bt4QKjshEHy9wmow7f3/aGqExgaEBYm6GEbk///XcvVfrj5Fu5q
bD6LeqBAnk/AUNw6H4HTb6d8F65aEMB9upUFK5YwQMQAyigiWpMrHp8UhZ6r2RjyBw5QpcCX0vFq
U3vz2UrvgxNHJL0vaBp+Cn3b4EZjLWHHUGJ7W3DW17HfNXw1FPoNIus7ukpWve80WPAnEKgjISew
i5xY6uIQlb1tT54Bav5VptzLAv8tkPzWYycrOof4othoI7Qd2jsFl1bCKRGIfUc6YvDeHtJ91Tra
T3Zh/hFRYD3Sp0pRJtojCU6WGMNG8ygmvdQCsVNYukdCpIVCXQUEwtYqQvgHwsb1BjlgWPdk1oAi
2nfi/NDbJSkmgNrRjBQtznrlszE8SDqQv9/HfbGlBVAdW753jLVrlco9hsNT7A2E2K/gG8nqBoLH
v1UZOiQFQD1cpGJPH0zgLPUh73otHQrhTrkipVRBUDp1j+10ZsXsMjfu1iEHEqM6HPVUUDJceA/F
/9gy3YlQdQHrxYNtboMND72gpOuy7RYUt/lBqKkCfsLLzMXfF3S88pOGaMEEWVk0ukDtvS/Fe6tR
O0qgiKMgia7qbpa2PKMPlKy8DS1KpxeMe74vKUtRJtkOBWm2vpLyk78adF0q29icNTQxHUMuUJ4M
LXUaZJFwA0LcbQp04xB5KvMbbbT3tX99TCzrBcyc+QfMTRB6HDRgdP1XUmupNISpAOda7/Yq3n2L
zq1yTdE1w/ZJis+gAyblWw1SbeGXrGmkFjex4F56cejxd8skeb9T2JPzT5Nqgf43srC2MsDquXLO
eqEfBJe08qfOa0SoL55t8L56k9Pp6wM1ve/cvTZKp6d8vTym0vf7XycALjiUqIOMVYxzK9jIRpFy
nGUsDWGkUWSxhX6M1gDNkRNEh1lA0Ci5mKSgrnkUXOsIrBpX1N70yO3KQTB+qBrCkP+9RSNurlpk
9pm/yqwWgEIs0ghJHTe0IYCruuU5Hoaim+C+sYgfP7YjH3/kB8M9ycY/PsFEPzDPQyhVEBIV4zpE
02bW/rD6ezGORpQGBxsp4xiuTiU8KJa6sJNtutB/aOqxmVoc3PYFaceClAKa+tdc7hsA21d3X0aw
NMWQ/FapHsDCKH6YL44ggVCzynEBo1hFYQnwt+45fW+BGCR47n1wjOjgAar/AheHXS4tH91SH7G3
9gERRoD7xFZsw+KvTeKU+ndwtjk7yAp41CwGjLbg67nwX6XYcmjlfUP36T2ffdBp8Ak0vJ06WKhS
ILqkjYCZA0/dr4zid07sj6Auw6Ubi+EIqy8qoThFlsZ61FZKvfcpwVIr1TT71puVH2i87B5ZSt0f
pXo38iyCb8Q4IZf6hUOIe4eL1s2sY3ELFl5g8zQYJLKT9Y3/n49tXsoEArNXG2ikTmU1oSbkVju0
RVGlG5/49KSu6/hErMGJmqUVYn8YokVR2ShxqghUXcdF8ss8MRyrEgRzffHc3x1CqZrQAqrSs7S5
6o5nOKogNHd3SqzK98557QAL+dxljRkXooUhUyXRUsoscxDtwhQAxaDYrW8Pr0kHmqocxFMSbKML
n2Q+briRzAPPtx7WSGFPF0O8AjLAtJ395v2MRp+1ziBIGbib0PA31ZRn3dLVjhxL6KIeMCJOU9bT
xjGICJZpidvZiuJ35bD95U/H6DglJ5TUqxwjpSX1zpz+qGPZfbSL7CooKLl/yC1NWAE84CoGVVxT
ld7wC3Rg0dBaRYk4R2j4iakMUl1ugno++Nc1sH37MGgsM9+1KdGfL0Mdniy8SxBgSWyj++t4VccB
5aQRY1CQJFjCXMs9aqNpzIhhRXyycWLP0aChsmRAtBAYBZSd/ndirjxpnoRzc4nLPhbIJDUi05Nb
WVUvBoiBmH0dQYQvNEgJAx/bCamzPkXw7JIUVL88mERlIoSYsS82ZPfaUaiBUwTL9LR/1qRBzYJK
gCL1IS5d5+pQtpPq/YTtsH7EKsfQHxtgBtc0YbvDkGd9VEh32yoW2+pW0+qwn5vzrqYwt+AY4Ltb
bojWBa4TdckUor5vRm4mrHK8U+X99kfaQh7sS9JrT3HiPiZ3/Npcl+mMPmzCqDRAzbTuqtqyuT/n
zNGQ5o/dAxm25sH5nZeHhESOQtsGVeU4Fkh5j5kMtmiH9SerM9KuZd+gTs57MtEPHyMpCIYtaN/O
k+bVLBdeQM3UIlGbbkqq3w5nerKXFbupczfYr5g8OkK09zBOZvPpFwYWSrJiSLdU3/Vb74iz5+BA
pRZWqCawnWFBMa0nMMY5gDHMZ4xoCkcrcbBvoxZxEbGU/QHKFQpGW3x3q2a1KdqV6gAzgX8DOn0K
OckZnoUhxf9MfxifRCemqEKk1zlqXL3c19CovIvF1U9ub8fnTFFgn52CTBlULOHa8IGswgtWbt2Z
tqbB1KLkS90HgcgGjS+WVA8lquF4Pxr7TSdK7oCeAtH+ZjDK425h0Sfh9CEx8TfFT6hQrwJHE5Ur
jQvjma0Y0K5rotJqv+8mvyRLxlZrtX+ItRUXt8KgntHi8vb2WKrQx5Wp2RzizBk09+CpEHnFV0KB
0pRz5tKvAo8E8fVhst9XCk7PVuEI67UdsRLu0nyQHNwsiN/rWbwTmjun08FQRG1RxD75AJrxcCOZ
RnKsjW8Qlw0RxPvJk2+NL9MUhX5rDJZDXoEGFKh310998vPd3ddv9lfrTuH6ra0MK9Md9k/4dB3y
C0W+KrAf+2l8C96xeQ92utPR2l/D072vBT6VwEFbpyIY76w9RBY7Iq6wZRkWVwui5+OC6VDcvyMO
o5I2uPn8oFZGmFhS7xQPGSABmWqyPIIOtoEg1V9vB5HgFsVK+/XW27EpDmVMXPKtF1FDAn3xsz77
OdevglLcBbgzkYkFc9NE5HbZ+BGPtLl/ihbvqRhuBvzjkmB1JFUKOuuV2Wa6iTo87rgmJhGG1R6j
c/VkhKYPQ8P6COAT6SrSiSlNoM4qHQMGGNPw0ABFdlBAEryxzMGDV1K/I4rIiDdCmUQ0Ecx2HYBM
NQ2sba0yCZDTVcfVjmgAtuG5bxsjcb+DvUFhUiN76mY9oR0FPjP8o0MYyCiK8oqN9BVUthfEhGyV
F0olEEZvzAjhMNfTbPbNPESoMjMMeD7xgO8feyKQ4V68j8pTRf+ThPwfD8VtJFDSMAxHCxCHdE1F
0QV7WY2/HdmUeq3gjsQYxq4LSqMRZBYcPnDryZiF3JgY+tQdmktjXoKDsb9jjl5e6yFx7cOLnAWB
q42eMkDmHrSvCQqeP/YlFfEba8EbU7DyOA9K39vL0PIM575fGERb8vkMQjEYCmKfePnFMePPYq6A
DD8d4QvCi33GjQQcHEcAbok06/ls+Ma+21worfuZPm2xu+16KKxihW7MIJGzyXToipEU9LsM+LD8
cBUh3NOOHiGTWJvuev5/mrSEAYh7q4m3HTpzczpjW5r0Gpmm79A1+EMdggUi+FKtZyIYECaIfcrQ
CaMz2mZB+mKt3g9n9/gYGr+KVzGkGJgD3brq9f3sL9pLbXkZ1HZfX+bKhfzEVY/UzBWZidfqtVsF
OvmiOQ/LJU2Bey2hFqyUyyMd5/UIN2L2MHjqU9TakeL/iD9saIFXF0++X6VMV8kwGPBkMiWZr3xC
IXR2nT4TtPM6M7/HsrgSbgLKe7D8H1s1bshEN10NJueG2wilzByM/LsQb+9OYuzuQNwlNXDc9yNp
v9TtFooo+1WIZifmOOZgBTJR3BHsXWvj7vuHeNVaenmfJQSRkWfMYRl3jxXKXGI9ytoRONtSvigY
LMi6bMYefDuVdwI7fHpX+VUfcl7oTj7amxgJIOi+cfeOZn7im1570yLXoLI5MZbU1BeY2gF4q0kk
PIXu+TqBTAZF9+W4+lezLuKDxN1cLXdVuPZaRGUn0y8oBo7EA6RVblHWDpRk9DS8tLzOq4usfNkx
cI8d1qbmKTKSClIjVZQufAmLXu1iOvTpr61MQBg/OqaUv5gAOBUkVozfQXki49FwV/Nw5rGsc0uE
e+z9uL6o8ZYS85dUzyQfm9H0UTkogctLT2jjX6VA0WbPN9xlBXKuu6Fa8jSCPnqOK7JnIJdiNVdR
1LGQ552T13f5jC7b3U5cV8qrZYxov0qUkqUOpkangu2IqC/9uF0v/Um1HKf3cra3NELNyyfqJHP3
78+LFXI9wozaJtgIYN447DHzmu1P7OcwiVh1qtWfbHaFG8605QHAkCuj4q+HDVUxZNlDGRHPa2ky
xWYfcjvVBHqEKEULBJtWhsmd42FUNpUH5QvsbmG0KSR+RFu4H8pQ5FFqXJRZ8gCAmiPg+63f3hti
HVRDVGdEXPX/NW9+jPC811pP/dhhm5R9tnZRbds7n39pjv/uBoE78wlcjTcPvI7hL4UqrMV2W8TV
vpEnd/i+R8sls06cmSJ5ueKa9/iqYt02R/H/UGqKiRc9OzYq3pDMB83VE6LgI+A2EAvur0rm75JL
wLXb7H3d5UY42mfwLO2nXT88tLE+dSyM1tfpFI5YNxeoh2ZP0KUciExiYhu57JghnuzKmkFpRBRo
cOZebzWRjqWXY7FG2WuiDQpuUg7EFYtn5sMLffspOa0KC9GW1/f9GAhCPdIp1oO1LVtgMMCzs74i
9YJLmhWQabBN4EySNwhRYubCsG1WbUrQX1cqqNYGzXmGCvLonk+yXK42vRAyTff9xqzzpZw+ixla
RA+cv+IUtQllX8zC8YWzXu7HcUhrYoJH0xO8pkKAKITOSP62wFKo/3t1wicbbBXCWugARSKVh7E0
sedNBToSaxRGZEfYDUYEUxbWWBFEnUJUPnuN5pYXgwUeuIyYV1GHKuXIjsowUwq5dkoVJS2a3/yx
svgUOnC8O3PtwE23Rc17+fmPcme8RbRqonw/nqzwlsylTHV3zlJopARlyOT7alMmtIo+/mH2hlw+
0ntMoRFA+y3qB1oyf3B5g8TE4Kpd6BmoM0gDkDmIkpba8dBara84xmKRmuko3uJqGwTg98nCYp/H
zDQz/10x1RhS+sWX04wDWFM7PE/QKrWaEkaELPyPmPFb4RNiBgpX+5inFqVzGIMiHtcIYHSBE/WR
/ysdeE3PiTfh4o2O3AGh0FsBZSgjNAC7cWmfXewHYBojxKbCiREonQouX9SRAq1JpL6CQ98kBhk1
YtGC2yLx1lGdI28O0XUZogXhbDLx5Rr38mBgLFY8SK/TdjRXrXHK7ke0mIldFOBD89EL8BLu4HCn
SnsEXbY/5Kos+K472USvtjnD4wnm8qy0go5LXvV/FueCeR2ukgVeNK5b/nCB+2mqahFHBac5EkOn
dl0z0TjBqGcGQwrLJwXcGhaI9waqVT+TPagst4ox1JRkQ83XhGx1i9m5sWV0XKR4lEL5pAq7oF/M
2lxTLDTqUCuwbpxSy/7K/huuDHgwUhT3Iyj06LTXfmfEk/inuPGWDqSXbueRi7+60AGWsnlXDEy1
iaWyGBNsvlVyLnODV7b/YwoxbiyGpR/PUGyWKhwzr+0AadHwZmKCRUr2xA8D0cz9YAT73D3kpjbc
jwpNmu8sv9OBCXb/CYJS0g+s9MErR1K9zYU88wxmwOl9bv8eAkcD2bzQJNJu9sx9/e+4xoVaGebR
+M40Eos1wHamvmA8G6vmrJI8EwWvHMPSB53fCM5MiL3NDvSyvkQjRDS6W19HVy+FoaSr6azCH83M
/HfL73zti4JdGFJIEXQKLj2D1TxCvAqa4APj1ob0nCM4mWEVpDkcXzGcGSbNqjmsZP335ZHd8ZRe
jlPVIom1cUsDRt8+kwe6kZR1skCqrbksfZz9WRkN3xYRDCZQCXKYIzFinOT35p5KAnz0tYAk20Ix
r3xn/6KxtwcNn/jns5Mu9UWc6B+HDcO3ZEIO3cyS1elMT6mTs/qXOzlkCWUQiymQhe5RIDXNMtoF
BgxQA+xf4wX6BCfSEDXtLyFinRr7HtGjUa+5o6NZTSwAI4hs/bXTB6Q+hvO2sOZDDtdqSZ7eduuR
h+SHCcCB+9InHoDXrbcYWEzvIJSLY3ZzDZ03afNkCBWgzVEOcWm98x8nF7LaigQL/NK5uZGjkbpb
nl8EmsY+5gWmtiVx3V6b28SI0h+5lu4/uPkrbfNeIJ1pc2rApl24wN00s6kJZh9wiXbIVE4THRi4
9qu/7pWjC3plcAxl6NMZIUoSfA/eFFf2dUtPCMZvS6ekowH+/Y+gkKCgitegeBDtxDf9lC9L2uzQ
9IX5z5dt1YMROJ+UPtVRx9wZd4JZrDkl30TyEwyLWU4Dzv/X3dpD2tX5rlOW9nvT2/vFW2+v89mm
d5c6nKUr7Vl2c+3g7fiQG7b8zMxbO6fDKM/G8KomoOcOODjhx8vyq+Dyauika7/013RQhpZAluPj
54S+XCj9j5nb5bd8ogQJfNtQyGS4WeazSdxPabsKp8MZ2k/819eGtW1YHhsWvseut3XN4Pqag9g9
zumtHcePcWxedbfK6BKp0LpmXhhdfZqYdBNx8hO2lXcVXWs9ikWvPlrDl4ixWgvS1VTCavoCK2NC
VsLH9n/o8oVycKJyfKQKL03bpVVkNz+Qm5OEf1VAVp/VSu+KzRdAvat5buJuAhtBnfmc3x5LtloI
IMZo0tnBvu5/hx6/pNg5XMf7B2LK6DZr6Vlb+jc7+4Y50+my0zb7Uq3ImLmo7FeXF8eKJGEmlzzD
U3voq63D5cTN75k/PBEtyhB+l8Z9O31LS3OxHybgtVwuNaHj/9g4iR2uERLJW20IIafd7i42bbO+
fyzEQ6q6OtTgd9h0pWg29E1REoP2ZrgD7YYqWjDY55L9EtMr4UTrUw7vuyclmAgxB0FAFNc4Bocb
aBrwKMZ773b1XvKTuLsH2LoxCJe9rWEsM+qjcAsGN62Erf2CvsydPPIVN5q8VHRt6SgZtd/NWU/A
C3Jv64+Wt7mJe5IrnOd5y+0yR6d2yp7SZSe4vhtAFkOaS+9wbQJ71ZdsN6YFYgZf6J2b0p18a+7q
TabvxXWwAzKHc/uhKfC7VlIsX1GZ7PbSM4TFcpCCumJGr2Q/FNciP+uuG0tgZ+S/7MdAPT6SWSQq
Gz6SW00QvMoylFl9GYT8rWSiu7nkeR2MlFau/whLToO8PRRAU2jv4VHLLWWe1pCJztgFNpyLkJOk
EC7XYFOEAdYDlIP0SUdd3x+TdpBT4KPb4RA6eXWfpQ2BkjcXrmqh4evgraqP0IpMxOPJ+8hNuAb6
TScpycxTmf2ZqbhjUiwBXvX/QZpaDFS521tK07N2KHzVjacnUs1wMFiZTWNSrQ9o/4WxHpU/EqiI
fE5tYzj7tJnxF5F1h3M0q9DUT/PFq9R3tqFlUNreeglxbI0vNieU5rViPrKegB68kjbR/YYc/z8t
6E0wORkG3P43PDR6EwAsx78AcjiUFLvBcQ6YcgQ51GVYW8MXYnuIsyuOm+xC3AFNwcunjfnMGvWi
fYEB/IWctaDjQZX/fGXdY7AGc40QFlnoTsgzcXbk9pYMKfxvDByk8PCjXhnRb7IGcVS6lH8VHin2
28iZyzfPA8kslbZkCftryq2Uaspf9YIa0l8STI7xloxnqrxrx0d9uB1nsfoOLCztbU+uAJQJecKl
pxw2bBwoRZQOdKGiQ2LpllbOPVA1/WnMNlFf5EJaJMZvGWaMJAkBtEnMURyLxldLStrfZ7h36bnu
vrnVbFvsD22Ck8BkC9znEY1mQWbBhbp0TiEb7h+p+rJr1pE04RWx3ESw6ffFpzjwBOr0RXLjsePQ
OChBiAqFxKazwii04IIH2MdaJz4UUiLXMbAFZJ8WjSNHgDQ2+Weatk33oljGVc2n3aWjwmALU/bC
nzq+eO8QN0CjSfN+vIlxKQQunWlW2ryJz97XWwb8EAQ1qfpFrDaDj/jtiVhYbzNbO32bXrZPzZnx
+u6YWgidmOYuopYWPcqLwpMBE6qRzOrVbWfgFSOPVi9eVLlVROsbvkMjtVaPfyGgYef4RRv512TM
TAvF0ZBEVOomB6Qlhi8ZNcXZx7z+AClKkCftdXDlzY9l6rNqLgJzn6zToTr+FUjGYeQfEAm7/ZHA
XQo0QqCKNMfQ89o20Wa1KZ4mCGhR3MF/Ny0+fKgKPxxsOLFBA9CRYHWVDFEuQ/epm6HSI+jFxcaN
iSmXaFJHxsPRJHnJWOVRuHiuiQw3e4eNPjRV7mDVz0rjZjko5u26f1a0dlXsgA+BRf3HbkHci39v
c59UDGvHApMyZPWWToJXAbjC/3gPMmzamViLVK6XgReLKXGSprquTqXiSnV6St+tyVu/rleihl8R
tdFtNWGF+gCgknwN5fulHgKhrkl2zSe6rLxgKyYsiYyFLRn2aouhYp00FAXaMxlPZfJs9e0utfhW
p+Vy5XiVy2+osNcXya4xekDA7Paukk4Rc74Jt+amPsQlQjNUJEuI8L25YIkqoAISTqESCBYqgHTM
J5MxdsTx9IUDfpZrBma3ydlhoAUcDwAD8906Y1Ieo9lbdnKHI5b6s3BK+k4Gdh95TkWHON1G3xhT
QYcZN7yViyFXnlDIELXfvBDfKlCLiPvJfbNUgaFfkvjvV/IusAEkr8+6zGQ+KeirVwZYDh+vZEFA
D1Lg7ptMgrrliodLy6XD8UkX2Cv0TtwR0DPoH03s5nMqfNSJkLN/XZ/FMUoPlBkOOMyXE27DqJ1H
LN5qx0DxCEP8O/4q0ydOdOTo3WJ8mnzFgdcGNE4ciJ6AterSvKn8b8j8acP52oLRA30TABQ10W02
oSpN7l6agjJjI+aHidfUWRgpHki3U8KaugtY7UABfRC6lIA6EZlWAIiErmN/MUI8J39KEuiTHZCA
LgmMVp1zU4akq/9nyFwF2xxD3LWETvcoNA4RvdW54mnGYJKXgRB/PzGJ60AP4t2LNk51E3NXvUsb
avhIyjx5i9okR0hLx8mNLnJ/lpe6phJ6mjo5NoWsKCNhFbtVfJJ5vzZVDUoU7fDh6LYHKmp+uGVs
dp84D4vusVFwG/AkaBhzTXuxoO0ApQZBSylsp3L7fG1bQ8S+Ziu7N2CVUrM2y2WUF/Z2ijExOCOF
mvEY+l6z4/qfyWv86nT6DdYHgiGg9CfHxp0eZ1ZBeVn1DlbLUWoZllQ27zpdu8/nkTEjSIkuKrcg
qJjazJv/UGp5qHDHvywWwzyEbtf6DlCm2VWxtJevVOD0dr5mmYpBqKp6pY9hKoURLbFcdpaswBRM
FZj3mw8dQveSzlRM47MW4zyXBRpVhvRHHak7aJ6ILx0IKPl/HeLiluSn5K2Ytnz00qkf3v0RE9pE
Z2wHuHH/bpbA+ic/qQ6Pt49IhU5L42gg+aEOdfeaPEWin476A8SHBrwePOcZfX3i1nAA76yqD80M
bB6oPMHaHNQZaMZwWOnddVFe3MrZriK10vTR6mIwhljQgAn6oaiS24WWqlARhBnsRXQ3fIXS4qPA
37k+9cAezLnii9R2XCD5ZEvzbYOP4IIAYwKoF1BU3YJMGuJZqOQ9LQMuT154KtHa/6f2Qd+GyTjj
rJgAxwQRfZjCznGAkIJRY/g2Z87yK35MGgWmo2QTqg75r8nC6eFirGILVGdfSwqlDo5BblezwHzm
HWDuyRWnO1Lgsm0gMX6a/SG7rpz5ccW0j3eX3RtZKI+5wgONC7hYt4/tyY9nb/ebAlr5cWYeZylj
V5kUYznGUghyO823rpa39n0RfFzrTccvgvMGA8h7+FtJlWznw5r7equrfyz2iPY3ufbB4rNxDsaU
t7M3HPkiEtFy07RIN4EI4kDmzRsoKqqbN1AGNM+EneyEVjkRfrNoMrJjwl57zgkpEqSWJLjOmh32
WX6PeGwH2PmALYsWqLvOMWK8sQ94iaQBFxPxhiDDDZ1wwM5I5tAQN1Rxezz987wVZreQd5HT65BV
gs9IDZPOvuEGH6gegBTgXRWlWXt4BNw6PTRTexDE7VUOsHO3MqfsEolpiUV8n3wUbJQbo0+Mk6r7
RIPAGB1iVoSYysipgSgwJfY8VUm6V8L339AOHrGvNohTToju5A4N5HMfgkIczUFWqWlTbkDsEGd6
znktgNfBM0ecLfDPZe29puCwNBMrpMuS1CDeSx3oH65L8/d4g1+RkQYkgdlzFZNJ/bv6DMDZ8gh4
8jbh345FNc2Z0OJOLHseQCZm6jDJfLDbJ/Zc9CjozmA94hSHCE9xiZxxGNP2cM3UDiubgjkDYBs8
pMOpd+tayZbI14ob/LEMk2HtTGZR0HSiG0MBQY1sf3OU1mg55x7wWrhmvU3McGSo09J2B7ADIQmQ
Cp8y9OmemAgVy83p70rZ+sP9sIo8QI1lbyBYcMHwg9s0ZW2+v+DBZTuN2ezTMX5IrUL//8i7PwI9
JvYTmYjaHw7UCCsAmoPOfREVbOI+a9qexyWSc8vruY5mDiJM1OlU/N/+i57uh953YSybC4TMQBLJ
MyCVhAt9CCNEn5qkPY+QwA/2IfJOH/wSJgI2D9w3tjQnrxFR0oQN6l1fwoBbObtinVDFHDFiG5oY
Yt6lv47vxykERxgYfuXph4XHekhMUca3sCPywNSEZMsMSdr0TZbHftDHYiJpLWcznkHdoV6a6s6E
c2s3hV6VRf3ibdYIJKbaDpUdse/Ihlsrl3GaIj0gDrp7GZ7ZUR2Llj0uc3hMmNBrZ+tcrH1igupV
jjILYPyIU6ID7SkmCron8zqARuPt8+qv9u0dgXWvK8SFQZ0ZWB7oOO9V7yn+g4PhPRHcMlVy/0cI
FrDIc+8WgWg7L62hyP1VYSeqnUbBcCxuDuw2Zks4GcVH2fruouOyRs/RxHT8BBWn+n9weREmMcA6
gtSp924m6jPeOYa/OoLDazTNVmTctJ+bPwCLhc/jCpDxvWCRl0t6WJNWmTtMttw4vED4Yx6QKRzU
4JiXdb76QN0jHaLIbwP75VOEGDirVRq4Dd5Gg9GsuxXhlnLAAsjia0O/q7b2ufH1RkcIe1+RMHaG
7rCSWEJy3geVKgUitydH1flIDBNc2HjGWPXMuNtPbqPDlEbFx7gR1OPAXynQPHc5d+KlT/zm4QOH
/dOnXdGx1xEIIFaUD8Ci8gXyrttphJGYNvaYb3imskjX3x2AuAl7Rj7YLmINwfi8m/GmMDMHoF1N
vWhXEGMQCN5YrveqGsAVYnDuZWiKFpXsE5o2RZpaYs7PRSlXXkeqE2QT8fl6nMa1fbqF/C+qMpWO
uooBcny9vIMvs9Ymnjn0NROpRbNnkAM2UJISVko/iHKINAOAzzl3/VYpzSqoPYERrquPQtPDI1Mt
q/CS6hEIt+OZJ16r3jUAq5V8VyfdydFNnhsGmCQRtUpMnYovR6hRsYqis41Q8PxFnk3sGBz0WAKv
fixDBSbyvpQKtHc89btTL/fDEozmaLm6D2Wen0IKdZAHq3EuUoUzbf0/EI7P0ZKqwzZ1Hefvz+MV
wzOefJ1n6MDOoonbUsAozHqf1Bc1Q8swq6VPB+zQy/pxF4O9a1+OepWKnT7k7MM90JlSBsGA9iZM
dIN/ICy7TRHuPEJjACZYG/izVDoMWTPfy4GNnKtlJSJVGPbCUPuMupP5jb2FZ6itb13t/g7NTQtd
VQkw+j8oMEDYrxjmnKEsVSLQo1311OFqQuFXyyhBPoO1qucJMG3+RZu2Au0w3wR4w/5nkqNTut5o
f6Z4korWGJqjn5LzbXHtxeo9o4GDQ+mGXDq8OTYTbVuwh94P8C2qaamv3wnK8jDpeX1LrRWUubTj
bXZgIGJDhwjrzZi6i32csdGldU53pq2VdHdFr97Hr1+QQr0gRVcMVOLUFp4B/y5JJrRZvJtLi54h
el0E6Y9YxNOG2JVPweIp/FTY4/EYozqR9wWWFeXQN5T0fIWrOxggGBka+2xi3htLfpGns+AXcLqw
8+xdr7wSJe7nYS2vzaQ8kpm3tZx6Gc0yywGzMA4gZk+/RsYWqHTQFctpSj0qrb00wx/YIJiKCpe6
zJ3QzXwWiDYBjOwx/fbi3jZOx2sp8GZr/Gn9REmbqS1BHboP74yk9j/Sw8gUrnML9A/ftQFiyKCT
joXUul9Qjvkxyid1UjVdhsFTSKKpWkRLOxv1In0TbTTDl3mg2rBoQimnLT/HzjX5bCnhJKJVA0rt
mmFx9Lb7UdP+cOst1gzwyHEhCexje0+B3IDg2sBnL8d/MAEkC8PLrIG1d2qiRP1OyIil0jxLwKWc
KHRzGO83zpX4gqwv15R72KUgFZfXpvWc6iv1eurzlvT13Hs/4n2gityHfn8XI190xrBclHl2z5DB
JCSENpa6pDAqWpUGT95i0QNtsQ19pjOr8FTsZiwSH75eaXKzjgzU3YG7WnXlIZmGdCBw+g1VyNu5
6zHmrXvBGFLVxFVwp2YUGQJ4BAL17yN69q6nQMZTr3F2NSbopjurrrKRq3d7tsRSLVmXdJB4M86z
U1fapeuz+I7XqrJGimu0mNpznUyv5CM45+FcWrsStKA1Rgxs3eRSYuzNZibfAJ1+ZOAPk1uxsicd
VgfEI1RY4eY8rYgFFqj3HlciM2fmqERCTqVb6Y2NY5ikvsFHfY9pSO+Vk+8LMGFlAMMv3nbF1NJi
2QNkN3Q100/SFt0o84vAm/APwMXHe/q/+WxqPRMsJkShMsaoGaa4YJppXv3uP1oD/fnYFmYgq1OY
tM+Z0r4BGb8MsKbb1uysyKuraMRqDFCFIDq8jKuxqK5xzXPkXejZIhLY8BNpHueTV99QcvDCHlNa
VHyozcGc5jaFEWgGVtU9VT+k4sUvpJhfKCCWwy2YO1FYNrtJ3f2Pb97Hhhd9toxyTDG4X4cU77k7
GX6ULTDbMQXIe1JwVnigREPYXUhUWOggBGRP337HxbRdhoffnAklp/IwFHPnSz4Tl8kWIKmquEsl
8ZL/5COwdsKZpj+LIw+RO0tFBlDiiWa+TYsdXMWI9JAx9m9K9ebFnr1wImuoYO2jYU3VjyqcEnP9
tIYOkW+FNECioizCnJ0zleGXuJvxHTjBzdOY+mL/0K2Ys8nKf0jOR4/TvDqzykBxjxCnlEbcI+8B
sEVNQ8PK7FFE7T2ivpNOqjLuRBXUdqBcmh37L3MSvEGmb5XskRTH3EotT54GvN3lpp5VrAI+vqrS
JIPzP+0W+9QRyRRsdzzbANw4tKJHfIQVCZrzer/ujFX+wio+Lf0jLtgSsaOP2uw8hlfu+TbIVM6S
ZXzEM/qzdOLknZNKfCXdKkowOZJ0D9623KlOXJJi3VW58sT+I5L3L7VgLgZnhGlQQq3uFcBFoJKo
mPxRB366hbPrjHnTXLVzLhlEW9qEWY2kIMMJnY95kXLyhPd9rPDa+Afom1azYEC8TbU81UDTXFmo
q7n9st/y6ARe6fOpuvbfafg/Lr3XDBtVobk0HmB0V3u00l8hrQTdpJnEjYWdGI8VjZiNfJUUdPh2
ffzphqesYIgdj9/mohSPwgFj4i0LJOPv++Y8JdEXEgmjXJuuBgOAT5QSBYAhkv1xttxeOubjHqmW
7i5d/s/wPUQcevZQA6xKVX/zlXLAzuMmh4kTFQh5ohs7Ei+Sre8JvDffTZ9w8nQv12MpH4DzbD3C
KXJ3+YOUm8WBOOqCs8fyzc7FeiMk84ECxuMYHA8EcPIfiFKVaG8yhapq6rAS0gSJs75HdBgRVVQ8
i8yQ/c8hxk06EWppwc0XhA4y/QozJuLUZzQwzSvdO2e6vxKBujGYgEHVyUqjjVIxhWgu+bFljEHC
9cWPQbgXDoRcwFfhq+K69E2VBPw2569PtdobnwLSqKsI21VMjAoLCi57eY5qHQAtSSnTHDxP7h4f
NgNN4go9Pwlk15bGdvigrPjGrXknOvl1LL9cAEUtvAtt/ogbs8VGSdKLJPOqT31oH3aPkwrN7UwF
CMWDuwI9inBRijHDkTf987nJZBy6eP7Vfw05v3rIpamg73b45PmI3SkK9yYg+YKA1ksVipJMk4gA
vYBa4C7X9/OjXyDlNWqrt/Qm9LiFmIHt0bBbxg4Ko0u5cp6Gh+v4JrnPDoEj72YQBzdgvZ4jxs6N
YUUMk52Y0l+plXjTOwR+Z7iVcB1DTStuPP+OXd/qeQbI1IXq0YGbhiTGM27w7pnLeK9bywaAeGir
pKilBQ9mdKP9OI9BNK5B3Kz9TOu5e95dmK5fWmTSXrVmRqbnHnvHybrE5hIEjB2/mEmXGLsel09t
SbFRvWnwr3GJ2p3AS7NERzQ1P5/keIXJzM65tKyVVMEIFWISu4cw1mSKLS/jpb9Bej4f/+tb1Eh1
XpKnC5p5vbF4C8Ao74i4Vls7fyKv2MDouzHMPWhO2fYyyZpB/7KGrz3d/V0gISiAToivNR5Wq9jJ
GhLEQGlKJlNiM1J58jB2Vve00tmTH/rWm7Ii5J9bKQ/eAZ1m1sG+S1YRY3nkbADusrv56EAUqvXl
poCksfdDSCXyUBLghOJk2+vojJNjWzLoDRnu7PsRdZFc37cIXlRj718qgixAQdynUMBlS1B2yhE4
t77+Di0BdSck00ue8aT0QLap//QqW/stPEPzZ+aQTiJvW0jAbplJbH8qtFEOqwIXvK4kv7sRXAuS
TGRl3d9yTyKsyqXukGrGgx4sJv+XDpI0kvpLro9Hh3qTeybc+ecqygs7tPwjANNvA3HiVzPf+7Bv
JxQlHk/Fh/D09LhU4jiXuT3iAQ5518G0RMs3ap7Sw/02QTmWMNhHMNM0jcJDnZ/exKLkowoHh9xS
9fhOmimlmwEQz3xkp6yMToUJ9u1EEy/AeNr0PaiSlndiflty8Fa6ivQKkdq3tmycbWCgQdptbyt2
sKh0vsg56Q3Bp6U6GG1QZnplbWMycioPbKyqv2DS8dixQ2sLTVB0EgLIBL7TCgAp01KTDPEL7zkw
V4beTO/+z7zivi8vyegPSb/J/0iZtM4fKTHdyrwPUjQenhHNWfj3sdSgEGnSNOmatHcEOpeWWg3X
NsaghO0zPV0HmDtAV7xES2Ol78ZLKAz53dXI1qLrai4MFHtb0U3vzvBtMdommsMh4g4L/4dWG0MX
MEtam+Vqah63IHKJZDQ2NZnrPaLLoleNKiphPnYchu92m42S7J6KVkmb4aMmTE6EoL8Iu50AoqRo
HYD5XON0gpkM1vwcZHMiwJEDg2wzmlV2rkacnyAy1fyYplfCuKtZ9Z1H4m00P30K6eDymLnzlWxr
JCJ3rzb/9Y9yh43XOykyneLz+n/Ay+2rtaNFXWZlEX5eHlhxS9Dk7+pMZg+yLdOgPfRFiqP0sObK
ohM6OtljJBIljpfzVWZGVNBkvhKzG0ZvyrPCGMlumxOR2LHosO2Cbo5QYfzNEJ96elbQGwBME2O2
hCDJb7OiBZxf9VUF7cfvE8pwzwDmdcHxfBc1RLLGnOZ8joUCwxL4npCbPSnyumsP/UJa2lI78rlF
W7f1k3/iySlaxWJkHg7/+s428Q27K+w3qCxvpoMX/9C2aUc4u6xUtJ4MKCSTPJs+IXyVFDmhagP6
oBrlThIYVq7sjZdRN5BbhOxWJ6CcYQol5gqTBFm0huvRxAPk6aAd3n8DqTWaa/95I87g+vP06Ki0
M/fdSVUgRyaj52G3Dr+CMpy6XHl0aCcFpEn4qn5JLUE6M3j6wgaBXjIUoEey6v45oVtjJTOanHTj
cH5Zr0ZHzlJ2Zt562OpNza6TuNCyIHY1pR6zzrBa9tiiIqIWSioUtjBfh0lrcdT0sAQrEyjyYvmL
NmVVV3a5lbRcSIhZtjr2pRYL0VofoaOCm1LHFAhgVL8IOO8n16IBp2QwEaKACAU+3Uqie6UIy6jv
WY5oyPqSG6FjmFHvCrvdNXafNSiHAII9T830tQYA7AMOk/TxShDfTUEWUFrjKqfi+7hwIZHI6tcS
7p6MDvnsLINlZgl6A6VtUnStbslI/3WIw4ojDh0tteVl0sQCJ6eYT7NtCsUUz05Nx7c77Wg68iI8
QRkA0RnKpYG/8Gv/l6IdvBKvyEsBQWqX3r6LdMO9zmOxs88LrBBFWJydwhiL2YYfF2iYOqPZC6aE
3U+BR4dOBFvOxVn5oSRVcHCyt7RYvXQnE6xJCQ/o+kVQ1fxheu0mGFah85zud2pd+dJWEQsqFKZp
sKTz7IMsJlS5N3aP3ZEKDoY1IB31Svs32JIqMlMb3af7kpEJczDc6oTQ763ojUiVtEXKuJEqc6fG
BOXZboEWQnMXYNaXx6mUOHZ4VmjtxbnrfcXsLcG+F7XLyDtqXftXIBK1CreQM575O3NeZ9rW9tDX
4OT8kZMEaQyNrjoROKB4Jc/FrwN+IxjoUQ5Q/B5SRgINMCon2Ysu8ykKCxS08EJjAQ7v4JXpUTHE
bfcC7GHPvPG/Ukv7cskHY9gyzsftHKqm7kqUTKIHRx7jR+siaZwxsSmGDOeGRRyxW4fDaRX7B8nh
j+pbMxkcp9Tazjmgjxy8EfUlkwqBWltO3B5u5mGFlwMw0gFGMTavwC9VSLCYOeZZ2l5FiNob8Ngq
nZqYnk3jXShWi0CF4S/C85lXUegfsfX4lk+8pRD3xAXjZu7G/UMuHJPrLdY04LHEStCE1Bz8P48Y
UegKzN5lB02UHeXgreYR2aNiV7EEuQOI+/euY5ns/Smp89CEAhtC+BlhyT6vmIuvokVwBAq9rCm9
ek2dliwkkNfnCl+ddPeatbJw9SWVufRCCVQsR4ybAu/7zGBdUqYZP+ADHGUsc4iSafy5b1qhkUcP
nXa618bO55KAoSwB0+g9wUuU4ESWSTAvX+4COIG8S9Iz/0LgSiK0TcpWLDlsZ7x3osbz0+YXaO1E
m5OMDtVHUILp1jo+T44XrcOgKNa7Z+UdBMYocLjdi/BmfO3/eyAKysbV0yZSiu997aYqogkdSZMI
34th8yt/X2uMvGqNqmMG/DQ49b75CPQT+bN1oCjRzLkaR9HK0zlgdDuc5djyfQHHrkr9ttPVHg+r
i5b4gndyWTVvwvk0DrcWtISseqkrTk9AR/DrHaueB+DH0NZQvwKIL5NKiL+ug/Bi5Iwln7tU80Gb
rXBe6bwsXRwkjQxKb7j/pttNCwqGiDQGQ+sLGiU3zzu1fNW4xnR0WuERq0WQy7ZXW1jN1bnqZ8nB
D4XTQOny6/e9oMdAqqRKAj7v3519j0hHQrrHmj46X+hnoKWQoCpsSo6P42NZQSTu+pHXhXQuUOSv
GpHxXsmDQ2G7dTMjbJ2jVmf/udT/OfjB78azdrHliNRu0Qk5s7w6EzTBXFBNpNxM/FE+gEz6z60a
0G2xwY2IoYf+G5my1CwZ6iAk1u+LScV9edFWfXeAcfWByjudYhSmqUBydOax1RhC4KfBrYRmS6CB
05cVTq7jOrc0pmVP+Shrpc1GOE/xpn6dw5nMV6KDDX1rPqEAKwLbsKx2e5MLCXsOka/tdgIhIUn3
GGDhoWguTahyw5x10JDYxJvcUfNVv7GgDYdx08GqTRz60OAN6Yr0ghUS9geIYvEMWqFepjay8Edb
6nEza/wNthel+HW5NoF250aa/uDp50ZLXnUcDTRgUsBg2BcSF+cHyF+TOgmVvSyKzjGPkwP42cuX
pyKFBcVqRkpqfDQdXrmhlw+SwYPozmOgVrL2dra5JGlHegh1wyBwehmtEl1TFRiTNBPiYDodwB0N
M3/ggPqU58b7qeWA9w8a5vtNaOv+UmHJsDrvT5P/tY+0m5yHjls2iXGhcP5K+IYOjjhJGwuJPAjp
b/ggOSjwexg8+polRW5OlQNRyBenerTpCUGOqFx7r5JH/fn8toDeJJ93XGj2MOqI/ZXHOi6Q+qaJ
L/Lmw21Is7x2fMKuOmSZn4YhTVaV2m6OCSE2eY0oBcsxmLgVvAtCB3tm98sJv4Y19maajxVU2m71
U3IwVaa8EX2cAx8rRUlOIgop9FzztY5QOXEJhHmopV1djgolPHaMT1shwky3hZGLzOikm4w+dvYb
SZHQMvTWmYmas8RghDIW6nDA2vh09QnIul61bTqUfv58yhm3AJYtvHM76uP9DStydUsyMMgnXHUM
R3XdRnwhWyom6XcV7Kw2eMW3V5M6fMGjpAGNgfd43zNcb4yU2ptq6LsdnB9AkBxmFQA7NJnbX1Yg
GujFRHCVZdczZfpjmDnn6/wd6gO5Jc+9yhRkkCZjjxBSJJLxQoevia3Y+B6nzgEJQMMKVv8CPJz9
hVxLFnKaY9lOa/nq8IsFxAz/BNYJXcygwqgwXxOX8nSdIKT0eZDleSNm5mcJnSIlQEuPISlG9dAN
S12Z4+KwtCMsjd57xZznP4kqbkx5Yec865/mtQ+mEEBg8ZwkFH+Tbg3PInOZD0B1nxeZKziVAErV
F+VkSRpTGs7rKiKhJ3b8Ee8oz7jJHpaRurchDOqDbpRl2U/XAeKGJ6mACFt0WmNwD41gQUnfe9b+
kSSwngELvCf3HfkG0q0xMHDnqVkoyj9voR1YUG/QcJEl7r5pAEPD5xTTQshRD3sfsNzk7OslP0fp
PnUhbJGx9yX0sAlttYiWkiEkvL/ili5TlJBPrvG0DB45jRSyUxIpUIVhqIaSrtfCyspzBx2+n+Jr
9lxV04CjaG+VzwalejJjSgnwmzqQWAnd82UiHNLdXzedOWvPU95G2P4WHUM6bFpTVgxO27qhsS4J
5+qc+i0moLm+zeJFSURJQcBqytwgdJBsQtheMPzjisdhfaOVtY6VPASrXv01Ix6W6JSVWdMi/ZjG
nvAkv0OlaT7qnueTRDvAUd3MJ99JuMGl4mwrCnmee+QCw0jeqHWCutwBNlFmWlYTs49pOAfagw9Y
2C526XUdyqc+0ABJKUvrTxNh/JZRzOVfAwyituPeIwJOAamCneMXySV1gtyvqH8RdzumPj28DeLA
pPEc2fBODpksSUmkpapZ8xWOdmZ7kvfuPo0c7pdTC2NBMj8UIJZAzXEPMcChuLDIeplZ/7Z9ecuh
0J92HjuOwEoG0L/JnHuTx9lIYuYpX84MmTo4LmAgGlo3lliS8AdhNrX/ZnVXqBSniQJU6HI8bNWn
HfoXIZpG0t/vGBM6GcIRDYuZSeu0kPaEaJdc1E9NtvtTGL9xrPwXKl5O0kFaaqJd2ArvKRJM2V6U
f2wYkoCWHbiP02XZvr+pFWiHqO50oPG3mBfRMNmqqvgCTLVzz4mNaI3gmm9rZUteMBFB91zB/l3j
WX/zVK+L3GvaXVkCp7H4g0zoEqRjKaaHtemvi0sU7q0cwc4rQA1+3ua7vUCinaST7uIvvmHaE08E
RmNZkXsdf4qTblribDVTUilK7nqHFQY5wbwgsQZczx9yuEbmCA614vmu+/c0eqiEZdXb+6YLcRU6
DMpWhJgKss5RL7cjJjC7k/eO8C7Ab8+B5TrV/qnScDTAEIQCXODJ2Gv15Ofu2X8suH16Z4FoIAx4
0IxGUoQhOVriNrnt7E2GsC1l7gknB+qjgCMyhmi4WQeWhrYTy5GgA20dEk+8BTLPzTqrZ9z6cmfT
YRYPRyLkOmKzcHeLzP+VRPqzY3U0cFW8u8o0LnmEFFEQtE7MG6t6UERz9utHA00z96SJ/LGKPcOp
b8dBfnnvY8nKIwEISOYQQDwB74sXrpDKn9JYUV5Yn9cMxhqbJR4yXd3B40Xjy6wJhziy2CeFVCcx
p+H3FkKLHlpXdQKyQs03JmSRbYghsBEdgYPsCG1M6dqoeRg0UHXJcWCGKpEUPqJD9SBb1LXlt7gD
u6gaLAxPMGeDAfrXn9jhnl5vPuj9aQeJ9XwVUBQ9t2LRROGK4rkgfd+QvqYTFywY7RFVjf37jQF2
aoYQfqJTF+0+5qltm2LIE/38Z3qY6NTVslOHgqv0NjOJHvF4OTX4DJInchkRIHn8arImLni4Gwr8
uslKDLNNNMsAoqTeqmuOIggBNtglbK1B2Y5dgC24CQAUHle+BeOXCRedys6k4eQV/kHx2/vfIBG5
mrGqcyh6ybrblXWcntfATJ9M/X+pC4JCAB4szKGJn3Py9+m4nCPBGIPrCRFGiDXVuDxPnuOfYh0F
6QQnHBSVL7ztTlrspNkh7tmYTr4pBC9OpMxd9ZR6NWEB9mNiup8bU8fVSEGfZX696yBQcV2UxQPF
66BpMdHbeFzaDoDr0Zwt60pfJcU4opLrk29NvL9sAPaXkqiu9YP/aFzWvudq4THtTzZSYuXNttzl
+5WqxfGS+Hc8TzH+cSjt5Q9AtTG6jkMqa9yGWSlrDXfZ5e9xiaNiW8cs8ZHq4UUxSwhV10UvIIgv
FShBaaipw5e60Ofxqff2P7t1mh9jWTAvhd7lGwkPSVfDWF1D+AqMLzKSbNjHvX1pYVS7xHxzH+AL
qNt/JpKJbr/lfi0c1rbALxTsxPrQTwLhYKD2iBjmFt2kV+2cTOrLMjiMkPiT5HIWfjG9Z0c2qtP/
vZYsKUfriMTPVPvlDj8DMxLBwbcD1Hhebw51LEYHf8UB81z2uiaNXIVNMCO2/e+aAIn6Nux1ju7C
kqfdWuP8ejpT4MXOPdcwD55UvfdpjFeBn1ehhBWm95IxbH7aNiQNQBtHCuJbCdVOcwPmgQy7crSK
pIUuR2y5z4Y00HanH1x8x9F34xNstS74KlZe0cQCwTPPHWzUEqHePu2ZJlFyFmWXx92Mjsvw1LY8
dUQwWPxGew5evPjKQ+FdXN0H/tK2Mz4gQ2BVDGnIq0dwv1l6q4bZulAqMfCcPr++4xcbiO5hm7Gh
2kmkM8IngZMgiRr04mN0FBJUnfOPaqXsYU9LT31owXEyyOw0ZUuWl1Spofk9RDfNXVYRam4gsPcZ
iLMaHoGbOqQ1RdhVDd4syYkgQZoUb2jtKbsXf+E/2R21hbu0Z/Yp6HPhIIYg5/hDiRMrGhkwdgOE
y5cfSPTuh7VwJaUjtjuFWCZcaAEWTbrgPi68b4TddRnnG0zqcBKvevYwMPI96HKP/8b5WE9JNScy
mrTG0lFDoFfkewpAUQW69nmnB529BnZlzZDKGuiQVZ4UJt4YVQiUfc0CUwYZ3TbfAw1DEJkAh5C7
pWXC02ETWiYf1GpmtUYEYyswMbfkOZ9Y++DY5HOsupwqG2aGdEPBGQBNN3baQzFp8UKiUL3CGdGg
kw0eLWOL6JPREWStczyQQf42y7RclMLA/S+4IPvn3obogtUbu0hSUe+9GAkwnr030r5Z/OVhtZVz
yMSaQb5D2dHtD4mLuvN7ryEtJG2jK913whwPmgNLVlqINZ/G/VmugqdjtEf7oVSaOIqX21x65cNr
oKTXzrPI28TpwlqabRDNIzeDhUaIN4EE6qirbDfWykQon14ERB9Eh3OETfefw65A5MdUKOSiD77N
lsqSKXwzElBeejnLwuzjDgl1HDqVrQcgmpLLhKkMIrSmMvyZkg/yOuwlcXw2hLRJQ87bqw5zZ77K
lKdxdXGYCLE6C/zikZTIVkKBX/4b4Yy7t/93fVmpS7UNbK/KXvUFZBikvBAnAVCosJwtlLffjOxj
1EKXGOL2JP00L5d66TOu29WszpeleCrHcSuEhDS+4tnNNWRhmDCSWQ0VM8t+gsDtsPk2lq8o4Cbz
WvRXCyqtY8V7Qc0nO6jAFwbDeopgRspAu2NxHa4Qj+5p8JJ3ZM1CEqM+Lsryf2HaEqkkdiAt7fqY
0rph86fzkv1XfXRCOHvH0NvoccT2eRMuMMVeg1YNm+/7aGutjumT+BnlfQuGldEL3IQSyuta8e55
W7LUjTpRN4SdnsKKB9O/6Ks/sn6n5EI/sG5FMBVkbtONnO0v7e5vJwLcWZc34seM9+gnXHMscerD
EQ1sVSdSTBAW9g4TjLuDXxdzQDfQQEuCzIB/po0QyQaD4Gi50aAUgGOtC/oMf8I7Ha3xZGZBCCYp
pxlCzcam4FdBVhP34Fp5XVnwlPogYw8SctGjHDKtsZg9ZbanrKntfzfPAtz5zz/JSi4HyKsiVkCN
PbviCmVF0EWtYDpnpSBm3LjfV3GkKr8qN464pwD6lrnTiFdlZQn4WTzGlSs5CXIjZXMHrJCV5MKN
cUdLIux7wbJHi6W+GU91KVj34/PCCnYCQ4dr02jWj9hbVw7E00UV3e2WSsM2sN4FiNowZo9EYFjs
9BqgqtMbzNur/pp+18UslY99LXZnGb+6KpKvrCCM2v0vXzQrJg0K8vO5sUGRB7YtRh5lfhkNeA/7
nvMEvcPoReBj4lG97bdHnytwMTN4aVLjdv/WI9lNuBH+Qlu82IL2WojfuxD4O7IGuIQUh4hFym7A
jzM6DkhjZxJoeZivryBuSJ+pgTZKDeWaRyp1B3FhwIZjcpBbO4X5CNDwSqxzRr/EMkQ6rS19iQkZ
DjlwGSOPR9pHXMgwuJIr8TdhDx0NasB515IyYOQfVSx7s+15SdGymgz+kixx1lOfZ3NaN4Rc+fHx
B1BAYM7fQHCfjxf9Rd0D+ljFIbpCB8z1NPPC7uepCONEo2Dt6SiGQSizKmippFK/ApsRJDr7w2mU
VWiphchYjCZBsMaQBupbqgkwHtkH7rH4N3YIsrEX4ebcD/p4vI5jPpb8HahjIRLgJdSa5iSWZkDb
WdJAbZVV4dd5YwZ6nDERZaYoi+acEW0HpewcVmTQIIRSPaYpqMAJv9J+5a8G+x3fA8Qgy6I/CkJ/
o497qFtFQcUnJv0C8OUhCbW/uTAsubfBTM89MODF6+9s2srOQK0hI/P3KZSb1Tpj0IHgJCSXM7ND
MhyUYqhC4H8/CNdplMY4LGUB0iIIUKZtpYPiadZGv0EtqBZcpSCtZy1AwRcIh/uFxQpwgzK652Ds
YgQ/l8KHd88NfZyUSVlbjjNrYN5dBIfdwgKpQ7fKH3pasI0qvNq46BcN7SEUjnlRPNYjQl0Tz2UK
jePFPWi+LoQHbH0DEOa7ocSGD015erpjnUHtcl/EA8HHVYhI2Kw/KLGLEwMiB8wTZslhMQXQbb8Q
tYVvtAN5VsvRB80XpCg38WbqrUxbFo2ROX9SaWOz9iuUcaOzlxjmYdOujm/FRdUFTF5fQvvnqVoy
Q3nNZhdERIHu14iEPJd1uY+kt8RWK6YP6U7//scVgK/kHjHEpSUxSW0wnBWGbEmSZ/yiQvXhCbCZ
48pVsEZfjrca0arSCJMkrmb8kDU/XKrJ3YWAKmAtTMsWL/Q0ihibOT34nR2zETN3Wqfz9IjY6YnY
4ytuMh/7Whj1czm/sOZsOCk+OSQw9J9SXZFFl9OpaQSsgfFztXhvFJiaislFRKAs13RReOJD08L7
TNHE2Xl+6xcR5Gk1HJfVfYXUmOWSRehMOn1SfALI3wBnqkDl7A6WS6ok8KNGJwRa/tRxV2giq4Nr
jX/5JLlhJ8n+Lyt2cNxoZdBpn3fbOJX7IFZyo8F7XspU0+8e2FwDgmtahaYuD+r2RMiGdD6qqjet
321Av5VfeaeZuFixjubM0/jQIjURJVsYX+BX+JKIcasa/AY2/WCIy9XLNJ+HMhCc1m0fbG3/uaaX
CwnZfmnMf9YUsWnh21Bnghzxf9qr7+NGYPYtY64kKiUcThCtGlHXqbL8UE4/4kkIGm2P/JM++eKI
1TQuQ5oGLu0s+GqYGNaSOMrKBPymyb4mZQUpaTULhZTEzMYc4VPDft8+yRRNpsQuUakqxvv9I6jz
tqDumD7/vpNiCXYBkH4ixniLpP+LI5RRl6Vdffi3dCC/+f5ODh1tCVM72yAlc2RoV+pYaFe1P+d5
kkyDVfKXQxZZNRgQobJZFpjBjU0iZtY0FWruIzX+wMDlK+auMaJHOT0hkatLzxu5w0ytlYrYMAav
WmgFrGav3VANzKrApY+hATZKfDl/0d8MDw0/wHChyeTW0JI8eJZFfRasRqdJjvGwmMSgAaOwiWXx
ElfMw/+9sIvLiTlYep9k5CSIw0ei5BieWS+atsYX/HRpv+UDJa/n/3Pl6g6uWTyvA8tVoGptxb07
sRhQ3jjbkHQuqXutlVXGFyZg0PhhQ0rQ+Q8337QI6R/1/RklqHKN6314KFMa2AC0AnLBcC3ZI8om
aEMPh8GjMR7dn4LZdJgDTntFI2/0HuGPy6JSOHKd8ZIL45tm5odvLW7Y4MHy5BJntRRvQ7UW5xj8
z2aw2/8lsMQUA/CEvhTRvrsL75mp+r22YHXkEsSejXUCAPgka1w607Oom2JgXgfzld9qVkPf0Eyx
SjvaCMmO1LMoLhIIZ8NZJJdskeLpdlKWS3omhm5h7BeX7PsI7h13VUH0MpjxabICK3Puk6hy//ed
HYEEsykokKAC0wGZLbi/0pQL48V5mmanh5Hcxe1pASzbE6iVwbjttm8Lfpt9BDMUpF6OGGkVZoX7
vHN8nTDGF0+p3O3jZHubjh38Hi46kUN1Tqsfa8Zdn3gCH+S+p1Sn+x8M3okBIkptS+LLHA/dgMg+
+WHospI6YyLLzUEbL54jpHFhTR2+vQYhedrKVRcoOjcVI757reegmneklJo06I32Kcp544CXaAm0
r/afIYYCRzaKg8NaGN0EtdTptfO8um5Km4njLb1fvNBKqikdUGu6byYdoAHfg3uDY2mSDOE980dF
68Fa0Uq6JQrtNuQZ5vZDaKch3Q9bi3PBC+xng8N/kM9jsV52rITCvJZZEkw1Z9K9OkSdNHQWY3Ri
7x9fv0YZSqHRfzMD6XtUvjhjDl+vP+WDWxOfQ1r0K71OYgCoOwNiQWhcsOiqUnejQlwL7ljtLkVf
eCv5WIw/p55vqeeelvzvjmIp9fH3pOs65P2MrCFpYjNKQcrO26eFYIsAQ/WAWlH5hOHYdiYMs2cy
4PnbxTjNzNJ4OafxFGw2R3RfCpCcFqrsavGiaNMB5MwUhnRELhC0VuOfmulxTMp4wnfFXzbKanV4
L7wqWWu5J6++32d9aFBZbwX6EsCqtZB7ULnuzb/j3nTkhwtaHlo7Goz5XnnNQS1YodxzLvX9qFd/
PrOHTZ181vBlhrgJxWFAR4f3Hy06QrxhWrvQtKn4h4G9Frr2b2mn1n6NcJHRKSWDcDgQGi/KRG0K
YWWaAe5JT4xKzWwRT+R24hmSsWn73kZHz2BosfS8M5A2jWOiFcAdRkB+/9S45v7Lxdjs1IiGUawV
V0GN+yVfQLkA67vdrKgL7AzPaMi8xIEl6bk1Zz9L9bWjFGL9pVhIvHWuIiX6RruYcWPD3lOr8BX+
WJD1hjthv0aGa1D9yt6XV2jzFszuVLTXwNP8W91/Gn8GzXFDaZD6V3anH00FBJg8KlA5YEPypZU1
aMUAsPpcjZQpqpzgUzFiXh/28Q8FSN3ziwQjUQg2fz72EVjF554hAm52nlVxEgld7ixPy1nd/kk0
z5vgF/V1VKC8hlwbiUcHfS5k/IfsBh+xgbyMHdOnR+4yeb8wL73+sOF62Kig637Ez4mcAU0G11Md
LDoWG65RcCEsv9Pk/tg8nTEI/yX2hFw29eSrzlGPjvxAi3TsHrlFQ4aagj5YHOHQ77dKXgxUmOpR
skYy1O56JiOfmX5hlfaQ/O1BWb9/Sc6kDp7STNN0c5KXK5rA9XkplplyJTGKFy83tg+wVpniNVDX
MR9dNU4GpvnCnXYgC19CgtTbdW1lOVU+4rNJamlDCCUIOSi/i27R1PuztTdQmqUNwjYnJRzBBKCd
QNoWBVwN6cUVxd5DvnIYgmHnAnJh+I1Tuv3Z47nZU01p5t/mqGRQtE/W5fq7zZ/TdzfvR+RZm4D/
madNM94dOkypwLTP4hlPzfLQXbw7cOGfbTJLLAaAb8cOW6LhwkfloEzROYJxLWJCKhzX4tZqGmhG
7r07JjH5IZBPHgdOajFbFbZmyUbtgHVtehGjmqkq523Ba7/sF7/rxiSA3PSrs1rWLALSk4MFjvag
TC9b+TQQxhLHpvgusiyuMzY0L4PBjJP5XTXMt486sjUMi1CTaE5EctqyOGQTExXM9hG1kRhZx0cC
srJowYdUKqC7BasNwuJ90+x2fXK1YGP6SI7SJuVGgYFZMNc1UDAZDkZdZNbEUOILuP2SAx4wrHU4
PhtCMOD9vvN03963NbXOw/rZ2XpEvXtw+aJwftAzRNEmpphOdkt07rQlXfoZKQeN92b01L262MdX
gHo8FQlQa0w/0y5mR7dEQIJZBuoSXujCpGtk9vIUff6Y1NEdztoK13CE7Kz9zGOmCZo7vBKgn0kS
4RTmee5hrMnG/+5Grq0/PRPqD9vGTnIgh7tFCyZ7a91pR2Ko5XFp0UcSNuUQuruybkmwx2ZXVzAs
Gpb4q3b/axc074yIIV35ouUl4NRA5nmU4vxn0x3IkyiHhQd74wMeicbQP82VlB5buiXjVRrnRVXw
HMt5lbMPYhRjuxtjgDb+q5+GD3/YnrsXm0NxVNX58aekJsuxieWh3l2umXK3k0Az0yIybkpjoHXA
WbNV9PtdqpQ0T0CnG0xtKTkHV98q8oNVA5HdlCE8RHYk7BrbGRy4osYaQ0DNODGY+a0Rmybtdq9A
V2snfmXY2OTm/6uThrrOpHnQgJ4vrfYVMLgqk1Pq5nezdY0xLrO2RrjEaKvqmA2EhR72oJ/LlSl/
0rdfe8eUffZwAGZBSqEIri79akgitn0D5HwNYdBzidiAO0BTlmGf98UHceeRtMEmSQu9Hc+ROVAJ
olbVKBFsWPMSaxU6IYtBmZUtz85pMZvmpJqFvrE5/366CSNChwn0jmtmFNXLk4K4cPwXKDtDLWJA
9Kq1krD1XmpdS/UYAqtg6eDfKWWUyOVHVhrxN3ivOz16jlFjpR90/1mlPqTSPv+tdXkBdHAiuH5y
vN5noHpJNzngHtp/ef6yikLLqm5GzdVEVgDazdTBeHW0q4HYSNRDtlJCVgCMdH2t0ma/XJ5gKmor
OEfDgM95lqUVjmtcvxDg2Kcq/yu6dAL0I9rnUnQZC5lIvXrTEiaXdBLrwSk2XzDZvjk4jbsWRZ3C
wmL0+E09U5VmVP5koE6NkIiKUFaXItdkD0Fz7iXKYwGwCaZ6uN4ZHLgLKapsoMqrgzu8BLaIuREE
aJZUylv16D2QDh7D0yxte+LtPuVRvExIizdsC923a8rmWWpZWGqEKdt8QZwWAV0/Ru4v7Zc9n0Zk
vf69B4Egkw4o4vDXUPG0LHsVVQaseuNi7zjmDBgym0rs5kCIKlLbwX6G/rQMGaa0LYKhTqcckgW8
6RyKqCISJOQZXfaPD5O6iqtsxZIHu+jHfXowR1VE3ErwLmlpR0vLUdWiGQyYIj/u3Bfb9qSK3a4r
VlnXyRExMvAXqIReMiiwPCBhJEfe6YdqARfAI0+DaR5o7aGQXngxKL4xyYEDXSTnIHFs1otGe41/
V/m5DJDEKLtPq19idy4UrV6hixp0ayMButCs9bxgCv9u2/jXtLsG2wIBeZgd9BwM6uI2aQ39eLCZ
Kw2b5HMoVKrzVzVJApixojGAYtegJs+SfUoAoXAlJds2gktRXsIgGIcCkk0ezndPA8vTujKtB0yx
BTcvHcK0BZl4SqLJeAUa8vaOlM0iVS0WFI13I/YucZXS0rKsUKbsjvFpWovzDVSmQTYGtHqMheo3
gEIrTzs7fbbrZHZwWg30bLaaA81zc+NLraLuYGoWTgf9rztRhEWW/435qdBvvBK9TdPI0eW3pTxG
+v2MgjID9avcum7gLMfU/jsMorWH0ZkSi7mZp+ag/pNODj04y/vDwAeCNRIgXpmNc89vB/TVi0LF
74zagv7Z4y+MmPixFpEbz1agq0nVziGKa85K3CAGj4HLNuZ6r+og2iUaHvPr7XQclrNePdm8NycX
L0i2S0XtNuLGRl3apYujD+4LNtfMYx9+6Vv1f0w5FmdXIGjyTQ3xvLdCbBqtbwZsHFL9M8Zw2ulT
J2XvO9yrSvvFTelCeocpZZB72V6/pddf/KsMGRbmux0aORCeWaCkGZYkooDn78MvZeIwLr8ApfEs
DK8IoooEC+AVmFjMro3gacZetFME7HlHR/a1zW5x5DQWEuRaooYU8EaqE+oDhY889KdSVMHJC8RZ
vWlmxY4HyzZqgaaUC2+oz4wWgi4s4hXy3pkFO8V0MXrm8+w1oWctpMJb7DMiX+A8PXFdDM/HnY+c
7a+48Kl/WaVZe1g4cg6XzPaL46MVN2aETJPfPi5p3EJvgV5XvefTrjQ54vXlSZgw291fJ1ilGeYp
3UbdWbKU/B2TyOfxVqRrDwMU7cYs5fVfwgJ3lI8XhXnU8MdESc527RzkWR3J39JrRdqn66w3kXBs
Ia8ysu9XKYWqBMKCH1L7zRNL+RJ5fbjL47wTueRqp+RUyfS++rbKvzU8fNARE/84nTp61uJCPFjD
y6xVelUJRq5Gf3KNxChz9MKPYuKyd0Oxr0oAudgC6TOxuy2ssEHwPic2gBzWkXMyNmxYUCFhKu8b
qSjBHYsvyTEO4Dh9s1e24IFQOgQ22x1+f+/oaO5bHESjuDBkHSumu7RXB8YutD514UG3CfXpd023
l6tFGF1jkyHqmrErRsWI4mzQXprNdJAIg4F9Kvk/F3M3sd3YHeYTrfpv5cdaw2etGzs0em2BuiAB
M+51Miu8goHY8W0TiozImaWfNxwNvyTHt2HncOWGYwFMhZ0xDp5YWBPPP++vpq8o9Ra7EwTb7RFV
OI2gd2xkBRkpZck4ZJbD/LqkL7raaYm/Lf/XzCQKFPMjOri1EQFJCWAnhZPCS/Umk+yF0Ek1gv1X
DUzj51BFCrykOXH6Xi1O1hq4SCTtwhU6jdPAFXDtZJw+ILK+2TUI2IIUukt7Q1X74oNLQiMnMovK
SGlbFiUKiA7i1bP667G+rB/FhMKAZQqJNAPUSL5ddo+e+5634n0n4rREUXyE4hY6bb1Hh0ssneGp
zdtOf2jgrKv7WQoil06Qgj52ZGI/ra3IHR4IZg3owVuuzpk9kn7GixvJGJ7yONmPGdgOXZBWCHG/
Yv5vXRKwN3k0OlsnTVMgIoaOHuwn6bAVn63WDufwxCunPdfB6J4RkJHaFJljPk4ZCZVpfp1LFsva
HrmEIziyxPB8x67hNIRGIUDYU94Ce5J36WGKaz984cYEobBTsYOUpl8u0dUmH3qrimpmotwKKzXU
rMHGpDOozST3Xu4sfrW8M6Yqmw1tAOuGKFH8OWYfL5T0LhhxQFBQC2KA0eWGTgyyTIFutImARQvF
Ymk7IUgVUY6JWKC7I1pQDT+TiojsGSyu50DoMXj4tx2Tkv1PgcXmlqfua/gHpyTYHdn9dcqc6zWi
YMnRFKisPoiySsyfY/NFZxcHOXQvi6a22azk+raq/xhaXrChXdChDnUouEE6X1uXICMowL6LcDVb
iPlHxQ30uCyYK4C9fjSIKmScGfixKHDyHsG4xfDHyPeQq6X55CAGAseZhdRhmVfs0s5jxiShFzgt
SMeuRk+r5rSiCpNigSTC8vYcKnfNzur2L5GrRINgRrIH+aRmrFwIwOK3YVdG40KHkdB9vQcLzjU5
6ldth7fXWmVOXsZ5UG3JQzez5GIZFtitunUP0wq2mmGQ3MhGH3zIEAb9plK2pTAzeLaDYB6R6s78
mOdunMxD9SITiramj1XhJyZlLdtZSs/BEcdHlUrxiRKu+Eim3f0MrCzJKx40LwotVfJeCZl6dhJ7
u3qbgs4XPz5s/bjTcq4R3nBUyB64gycZKz0ZNHb4nCAnfVrej8zH9HPr0s8CgX7LTfbmWfmhsknz
RMq69oQJhiHIInSHwKI/Tj7yuXDTz3EMrAfFiF6dR2+NwkawDnMBKKHFWXI0yhrHAaZsJlMWpSkL
poCLAvnZ6XQHpEQsT81eHKLOFu9EhCC7mJzqjBVLoGHlZpS7bn+98Huwam3WV7bVGhOTJJHuwCgb
9Cd0ktlA7wf0Q04+wT6GIQYdeQOU3AEq8QCgO7A9UOsZ1dc6RJ5pSR7z/pd0Nepor6Ha/lbE+FzO
h5nJGmcvPTDBtXFXXxLYL6vgEAp6jJk18jQp3D+jYAolhV2cPwGWMkTSWn9qIihF25CEMM7naQe+
Ty29d1fqbRYYbRzdluc9aTxxbGO+TjCPLq+jVyViVK+fS/whlaZLBslT+LGDNkE7zhuTuiIkoBaY
dm38pNwmdAD7lhyC1KIayexZSZOIYOGKGaAEXroGhBG704ym1eK3g0E0xqQKEIxYFkTEGLixANpD
FPVfnC9nFHf7DQzWdhsOplvUXNP1u6jMOtc+4HPPVJ4QM5tzKW9p6d2Wl9LackeRjDHSKkkRYkrs
b8e9hzNQjNDKpqE+4SLtSr5Fx60A3P13fdDnjFXPQRz25BpQKFLKB/ktVi6sKViKMjzxnGCLCyyr
M7wMPrlBy+0RBlr36nFjKbQwTHC3e1CbySMI56+krUCl3Jegp1Z9JK6O4bK4ZJj/dSUIv7s+TZUd
/DuoIb9EeqdYezLoXOpwwwPvzDwExFeVp4Kio8YpjE/ahZVniPw0p1pXJur2y04U1rVz+Oz6HKQ4
0nUSFrmSRPDmBWQnwOQ1UZfh2f7SxA9M9Q9+5ageiG3MHXLMhZwBlSuy+2zCOdKeyeJ3k5vhp2ZJ
8H4iU0JFdItmttyjE4sXReXdl8vIFCMCZdsHUVmqxkJYlvbGIl3MqXRyo+nCq79BBgAbqaQ8vHsF
JQztFKjkG1+ODCtpDSy2D/7Avo5J46yODL8jbqQvb6jQoeZWUwyFq8E3DXbFYIbw0L/zJjZMnxRo
M7WsLuVb57wM2HUBDOaUwgZAwNeTdwoy9APdTvn2HdKeYLFs+r8hCyj3ontmfkBXdMuXLWI98EVZ
CpMr+ciV2ROjZZCh7lOYWwYE08ml2s8LV5hkW3y19vsVD5xP4AjNYw+pqaXzog9jHqi6YsKGlmlV
1VZpH3EROlPd4bzQNilXjuFgD62JTSzSPjP/PPnuiY4jpPJqLezyq4dt25hoDa28IkVjn3aBPfQD
GGSoHQcdPxhuUpN95t+CavGCYxdkKR0dor5Oi8Upv6Q+Mdf9MVanEwEGNW9uqTC5Eq2iqO5lGrZP
BNN/VdgC4IFwnzEgY770z9vDuZzicn5VNVmwi8nWD8KOD6QR7SP07UTZ2SFb3rD12r9JlubFoG15
4pPPgH+b24z01rOQM7EVGc1SJdyoVlKzR+Bd4yh31DEPkoos6lmwD22FjC/jwg1uywKb35ClFwO9
4cgCqVGEE1A+qlSSRFrwCY9lSerWswlUDsF2k+ryfjbGwoO/Iory4XKNhSZ9GzHBXBYByqVonwKy
TkUMg4MPFmD4RJ05c9ZJcqlqza13bIMot+Maruq6u1o/Ty1MB7mI3gd1e4CckU8LGXdsPj8BviNd
u5M6/oJesLDmiISKRgQtlNFVeTkleRbksozpMvT4guyQLoX7li2HawyoKXZuNCDv+7/8YsO1Hvx9
bp1go/v3cveXQHfgBRgfDeLMb9ubd4knc+LsvK1xs3Kt8TGh6bOAJ/vB4KdbBQLP3TbuPOR7yduk
V9AX74WWfm4wPPucgFm27oAc0qKoDeePvCS7BHiQv+kGpo7RwCgHkavq1Jm0fNrXgP67bR42av/+
QQ3wHg+GSj+lCAhhUbAzUwimWkwJikO6g0OgoKMINKHy6G3YP38TrPqOjAQzor3F3cpJrVYmA+YB
QmPA40Wd+45AcVWn/Rauy65UewxCp4WF4x76cQAiEGar0rF7/lCNnjB3ljr6LZFhgUJ9V3PYVZ1M
nggRFQ5Yd4Qws/QJGDIrLZg9xtOIxgT6yrAnsyW4/bt/5ulps7NNlh1DQXVIrDSX33VCbhUigVG7
6g2WiE5KQ9mcLe+K3j9RfwuoHdSstXplmf4XlMN82RQq9j5RdNlrYGMnOPYdv32XCAYn2NqvLwwO
RuJEnnojLu8hyy33z0xxUfNUjlTZlEJz7RPKoTT8lD6V4AJhWhjxpwEWwGyXuJ+Nju1A1rlro3Cl
3b+VsQMNJXXKucD5fjqJjuHIltTp3aixHGJe3txGMgYR9o0/8+zV5kqqjuUU8FSRLNhYJLpr87MJ
qE2u4gVclOggfCVMH+DS7+gWJsBxNyfvmFT+MQzCmE7JzBVrZbdY98srJlu8MnQOrnZ3pycL5s8A
1iuqtYlXTNRB0wJNzuXwcLoNX1f7eYWGm0ExJWkH9H4ezBJ4HG9AmyqlmEjWLWy4ys4dkM7KyDOp
q5p4LKNfHRvalgOVp4HTLa4EOJ6TcQ7GTZcF6xlTO3vMl+k7YarBc36RVd0Hm9/bqCvUqx/BaaVK
et7CiUYAtAk69Ky4UFjvz8ixN+8s4/OkYNelAJQ5Nx8rVdzl9fjW8bZiG0RNnjYxiZYqQRO/7dmw
0d1sDGJN9VFuXbllR95FedFbTdVpBNubYOsja/TlzfV2oe02ctA94sxLPQn+jPJPwUeK69sAyI4i
M5PQ9/FQYysPZomzJJRiB3ESUCCm6wq1H63VpiDd/ALV1Phx9U3Ae4Y/opIaI+GHHoD/HjW4wpDB
lOTkDZ01NdZ9HQ4nQhEyo9IucihK0LdJR6cPuXzDFdxqXzD53Y8ZkYpIW0da97RsoZYof4EHPjsr
r4obDh96RsbmFkoGgBFLc06oKEcKjCeQVb4Oykh3SRqmaN0xfqXOGn+T9HfP1ihuDnqMMkVRCijr
qvCwkzOsrVrCsnsAoCa/BBO248o1s4RChHz1uq9Q3AmGv/FU4DI2y2aBGcbAn7xCfl3czCARY0It
/H7B79hLI3ufKeTtnHbroCBh1i1AfTeivNKtK/LANJ1jpJh0gC/2HWxD90xJ0YbDn+kpgn/z6d7Z
qOQn117E7abH0DyR7BxAIE6LJeGVvRf3/tPJvfPB/0eL6WkbKjHcguf+X2D9VpVdkJU2J9kNOeKf
L5BZr+ntjMYcZiIbB+MCQZMH1VVJQk+MRIHTRcStoo/tcdHsNakkWwKNyApSvs+hgjtOSKvq9xY9
Oqpods4IatwYvXjIGNvDSEQ0Guo9OmqwcqvQnKJ8UunaXFRHjXcPyTlqeQTY+6dMydE0Io3D1z9W
66vr+w7kF+AJ6W/z9BnXRQfRgkEslF+jeNd7qOuFH8F26L41HKb2f/Z25w9v3CjDN13O/DZqJP8N
n60uJEUWDtIFhEmXf70L0rGfCtrJJh302ITrL89Z8pi6RhJJkbZCYAOS/bjjuqPPP6TEDVS/rlQy
AD2tYxKZA7VVWzlVTLRRtY5R6l4KtVXkInwhZHBMwZ1DMFb4+s7P2dvb6zxW+c9mQ7jrM9Xy2zTG
AiwGCRF/dZfNHfr2MrBRqY8QvN18KpV3oNwL0WVmSaBoilQv+phpD+LWMMrrJyc+ULH0coU4n0pE
FoLdB70tg1U9qY2fym3QOY+It2g6h+DubuphUwOtOCYejSu7XSxnAuaeSac1NJtBXhEovoSQKBNM
s4nF/Vgo2ayqE390bTCZf7Q7IrE72WjjbXIY+qFynTRSKnoskDNoy64mcvK9boSIOE22hDk5zpGy
x4F3IjjlPEX7RoawsB43GM/CEDBBGv7Cg311lUsqyKOSuDwUC36vW2yuOjktuH654n1o/+9pj2AL
r/COUdz8TpbNNVgEHV6ww7c3wi/akMmvDfC5C2/De+4z7NDKdjua0T4quoXjZCKSdMogWMvEmo82
eDLGmLTfz9JpTl53Kso2YqnNUGm7F8xl7ITT2hy+Mj+dkWMughRaZxcKqvCvE0TKJPuTsIUpnBkx
23fNjr/4TvZVrct6AM9fgsQanINvP+dJzd1/psWY7O2GHj4u+kqSAVxlMFzVruxdAtUrRLvhjfbX
B4kP0COtrFrp8bpzZW6h7dQ48kA1GXFDUJcd0SlorUkRTUQNNAKVAktOxM7SD+WIqqkZojApR5SC
Ykiz0WtLjuzvRxWehTXsGHhEXafuzGxEaNAmksItIjjWFp/B8lA2ueYZ5ReaiAatBk5NI0vS2pQf
R3lpk2T7CcnmYqUSLAWfbk4H+rifiOCpkScoCHI+yQZpbgSKfyaa7EIgSoyJBpskOmanWuoMNH9Q
jSYOZBwWbuNw5pWtZK8IVQfUKyBGeC2xLlhsw2qMSmAXfquY+lHopQdcJHErRVtNNGLwuOsC3nf1
xfOYQy6qloApdGJhVfAP0DtlBaCKnMB+oTBmksWdFc2gUKYtzLStrKe/G3eG0S+H2DFTH8sMFo3q
K+F+lGUcUyDbrlUrCd7owGe2/cviyEUyUhq8QS9Va/Jxss/PdGWTJz/8KZT9RyxBQ68ybDLMMEt1
ZP69Fo2maByZo6EkFjKG2NlxNb9njMuby2d0f/8MXAgqlzddthMbgCAGg6jFCeFs7A9VTHrq6iHa
V0K0LfxP8q+/89tOcqkdtAGfO4IB/p7O54dmw96PBqB5HE8b+Z4yWjCgcqBQhYKuxGA65ofbU/AH
u9vlZKQ1S6dTvUowt6y86Av/EnITYccyPy7lunogNSSbwGRFxw5Jl3uIYiKBJghWHS4zWlid1qkf
tpFoP8AKwMUHnUPkGJrpeowz5qZgQxREitgQkOeLlxFXRao3oZbIMde2RgKsk8F3W/WvcNoQZejt
KAD7ye+Fqu8FmGdLSpTAdGjquOoHQFJaxIvcgC3aqs4ndI7icDDyJs0lyBMa9pXgwCol9sJ8/vbF
LpUwRWO7nLCkfvvAYeGvuYoLvcXYtnds40yZPm3oRlFeK5s69pWG8xjCZi6UJyLKbY0UVNlhHd0J
t++SCidmixVJzyAxbNC4E1Z8ESMKwGX/3H3l80TQmatLDi2vafL5P/w6H2ufcvrQMSOpVWvTocdd
sv4//MmDQldGBukP8+exxhTFu4kG/d0qPJaAUTcHUv8Yi3SDCJJo+9geOlT/8FqguBtGRTkrShy4
bMP+gVAgwj2u8DPmYQ997Irdjm1sOqJ4LGE0WCOOhYJDD28Uv2zq//2PkUcFdocSF6SsWMWnTFpb
WY2VkD3nyVGmn1Yd+Unmb4diV5B2C67mLmW9AkYdB7smcIzUYLeNUVb63UoCGyo9dm+EebILjimV
lTAIxa27ivWr+HGEX2XzRxQujEpHzo1Hv2XiHL0j3TKadowHledp0Wjg0lEiBJK47VvTwiXEGNr1
fwGHymauuZHDV3XKOre6ncnrvcv1yYIOIfI+ZJbm63uBt6KHuggPZ2Z0lx5x7hrKNmh1Tk7lv++w
sqB2u/a7avil3dIoeG5YuNy1O3U24j6yGTJVUdT8jbkSH+WNDn6VVBdrerNlxsjQaZAxeHUSCqAU
CsRwy5zFmn/neYQZx1VuWqVPSbY9qonmuJhWRHrikySuLG8JVBfMbxX8VC8OgYA+I0vQDaRMrU3B
PDIJKtEhm4/4qd3dyLZzYSIzwm2iKesHwcP62I4e2Wtn2YfGbD/M8EuDgdeQaKWr4YLs8m3MuQSz
qW8x7Fjshmz+WBWRy8P0ThBwiqI7ll+G5L6a+SKm9goWnI32qmoJK2e1YeFPcYRm0i0sbwXjGr/N
iwvTRY/0jkhY414BB9gIM8+iUbEoUhDGsD1v0HH5VyHOvLdKxlMVrmFDNGBq+Q+9rqtyhVQqLwFC
esHqIDUwLyHzvwZ+5moupPtPOEUY0nKcCj1Dwqbu9CXpDHAzumMTP2j+ai24qwqcuJ/HSr8pbCer
0xFDv3oabF2jmbyhpWvlaCJTjYgwoy+WmZBaS1QZNwHSF0PmbNbjiECqnotFVHC65ab5lH9EwtRg
SrUWZHpI7fqtb42QkFmsM/WoJMb3LRBpAXY8sIILd4lraJ/LvPOKbHP0tN/JA6mTXeP2jUH97iUI
APgPy4XNGMS5Maz1kUi6FpiAii6MAdaibYjIksYjqs2ztHfB6Ep1HDLPJpkBQt0vEts5C37x0mQ+
uj4hA5t5m/jSVJrS8G3m74SReISutQpkj7lTR7zXokBQJNjiFw8O1cYu5r4fGRRCFj/WXpLOk8ml
/ysV0nWGDgrUJFgCjuYr0ioSsVpkyge6EvK/w7rLF0UFnNHTcBUSH/9e2//VssQZMau5o+TBK6q1
vmXbtjU/C8yR7S3vhiNYy66EybJYkborZOmQQeRZx4+5HntGWEHAxO3Lh9kn6dIzkVNQSVTc6zHC
wMSjo4r6gq3OZjVrFrDPRqXo/j/jwFGBbhRm0WBElUnOzg16CxvDyKGwrMNhwPdFqANKDW7ZPOta
4rEC2KDMC/oBmwKKVIFyqf5njiehNdKUGeKrUfuRL4EFXilTWBvG+/EzZTc1GginnGwG7HK94su+
da0CsJSRJK3RS3EUqanCQImTl0k8HACmaT/IAA1kUPhdTIK1+8OePyL1lOFrEoZMaN8asc0TV8JR
pd1CeqBbFaQZt8Q5d+VPY4rGnTc1JuBco2hFOlpRFNNBu1AMWEmC82EwZirgbFFVEbKXXH/0SaRI
7sRcn2tAv9tgRixfKEVVly0Mpch6SPs0Hm+qYLEAZ0K/ptEwnU6OE+XvHiD8LEeBjCu1FRbBWLQd
yhsh1oTK80uA8sMnB65R74cqXKAoFwLCcjZm4gC8BbQ9l7Rodh+4mXd83y9M1yUnETCybYTuCAgl
co7eIzplJ0hrb/hK8rx7Y6LOxm32HctJbE4ILvJWIFrnNzWi/SRzWcl57atPKm2mu4pLL/PIbv6X
XhCLo4mVuF7AetTCX19WCIgVawKcnoXCf47XCuD7ppkoGLW3DpJdtmpuBHyBvYneEJpVl1Kycopg
Ra4/3b4qbDEmxouH4WrbdxvTFrWquJsWfCqV+SAkJBxIOSfM8N/VyRMavOADvvvln0vcFS5ts/sd
cGt/sphFn63/LxTSI0wlcfvABjDPDXDBPJsvsmstOY6prRJ6ik1acu9gC6Qmmwxreta3Lvp4QaOp
bkvbVqvhLYoG1Tdur3/bPY3jTjwZjTVs2kBQhYgd0P9AALp/HDg+Rc6YzC8KALg18SjAzRBsLRzU
me8MQsuxHIHY/KspqcJffLSpUPz3G8DWdeRmVw9mkZSzt7PE6YfTFvRyu70x2OgsES9zZ6hQA8PT
Cakf2G/mb/tssYEUkjIWXeqWB0qr3NDouQzuZfAMUzGn6LCCRA0IngA+L2TiI0TniutAqvvxXxQ4
4+0gU6l/W/GevmoJWqeXopbqKrmRD1FFv3DCrsM0lsBoLA2MT89Sy+VGcSggfHLxARp+Hq6iGE6q
FXO7Yf9heqvL30cmoDCkNo45YTfMPsW//Dw5HGw5HxbaxeSoyq3dNA21JFmAl8rz5zuPamsUbdPd
eYEJTMzFG3q9Wg8u17RJgm2RJuJM2Ystui5SLDP77m1MbDLe9THfqa2Uj1cpPnby3gsN3vVlyw1l
MUnsfZ/T7/8F4VV1PbAiO9hsSXSboxSDPvdP0olCK6oNYxDjgIWFQw2zOVxkmeFdUs0z0EcMX/yj
LMuCP1aOJ/hfir9SLSSHm6VBYKQ5WUvc986R7eYzB9hD95IKc65eg9x+Y6F7oGa9pILEjq30+NWY
g6zBCjz3xKJ+zDwayuweMbMNLPeUjASlVvPvCL/mwXn/WHRQjahO0yiyXbcRdow1fjKzLj6wumPx
jahOrpuSgegpivMlKVkHdV7G/nQv1whsuaMMrZXTvxdMmejgjhjFPT5zRyFE8jRjie93Em4m2XSe
yBTGrkaqat8hRihcgm+WqTmd8QIg+H9LHOPW1E99Bwil3uG8ah5hAcjLLMTukk+expLUc+GHd/1H
qtysqyyoate+XZqLH1LyqQ9B3S+elOoi9+luNn0rg9gAQCuw5b/CWQRZ9HUF9XlhJBl5gLIn6q4S
vxDxXUYXdT2ebpmDWcTr4N/wJ2tXMPoMwOB9RFurmCTLxzOWs+lW97BaHhLrKjlsg5F1Ksk0BzJE
ewYXNgEc5ho5WzoDpfdo/i5ZLITg4uklA52v1qjXG7seSN2VHnM6lVIRaY//RIP+VlERB1dkMTP5
1pQ9IRWaL4ypo9XQVgJXGjSpbmNWnSX9P8YbT/VMujIKB9Y6NxIgd9Tpqy7cVWlfDymZi395xoZM
dDbPU3BuO3kkiOuQyCWfFwtrFNuwcXs5cPzJJxTBrsDF2G8FkDZRYtiL34DJ7bZ6Bpdq06DuNObY
cK0+saQF7euZtKj2XSX1sRmN5iY0F6Avo3GxW9s1g4DkApAmrfE7jc2LziqX2TPuIBXDMVVXZvX1
jWqZlvHHYDa6k2XxbOs4+Qroy32tIHSOlesNz0B33rDYbrm8yAUxXqJUTMhAgnALZhESIoyreIqK
1ftgrAFWd0bco/n8/4EVhs8RFaX/ieWBsKLhZnb38UZIMYT18nRcCZ1mD9cNBOA7gbs2eKEvZK+1
apAOC1ZY62Mf6sE3wmFp5/25ctShkJutVd0JVgLJs0k7I81GMSQKxwpHiwI9VdkFVrpCm1J1+x39
JbMhmrFQ9zNBHoCSYFejggY2eHlndwGdq5LC1yE4Qkx4xvVVE3JBHF5jyaLkc7Jdimsu4h0g2nVU
2Nf7Ge/aRd08eNBPed7JSk3CAZvt/GG2AnnNfeDJa9n7Qv7AiR8KQUguZHO+A508d7ozzcvarR6z
5WWU8sLH9Y3hJoouvcisDzhmMM+BI5m3Ha+ihjdrD4brJfyyiJTZE+jheczPQZq6CCoV1VwAyMZt
li/7R9uxhPjszqdIajUWKtxxIMvOwV+9ZFPpbwiSNLbQGntfTglJpzvaSylA/TuSazY9L/zbpgdB
0KO0jXRPGHlspoxP+7K5MEFSl1+529uVpQkoop+0eYiknVW8BLwCFcq4n6P11Mb8v/W0fGgJMcLl
ge2TztjYxe0hXFpN4Ll4ixkkypi0eLZrqsomm5nrQBWFxsZBY225JxX3X+L5cVdHtJ0db3I9fLTk
lIrm1+Sb1DrNxxnqAspEPKP+dd19pvdJt9eTOFtphOUSMCEGKEZ0zHv5ELlnXQ4+6R4O7SxB6w/P
B40PZoyCsyr2yzKqIasLFOSYxJUkQRo1qZtviLxbWg5Ebi3cc1QCDtPagEhDUF346hbaKipTqf63
sy9A9932QiV1V+cYi5HHl4MjQemtbSNolzOCmwsfhgRF6dX2ElTfjtRlg/ET8bsaGYCAO37zSl7G
gqHcUzyNnJr1qMs8ieHjLk/RwSB22iNUlAXk57wDaJGQ/7dhCaP81TbWi5aXWHyokWib5BtSbzm6
+5iIkhVdwzL19rO+SYiBZWjqU8O4vlWoUsxfIMM7t1Ky/psismxcI0/GEac4B/7AJM+7+XywiETD
LI8WEvyBH4mJPuwJe+I+CGCA6N89yvt7D4m0ylpzeRHIM5Xo+Ld2Bt0BkQ/c9jUgAZHAuZf6gDwd
F/9SuejWHAJYiTbSzxwUBoEuJJHKmD+sJ9w8psmY7WkR8ab43ffpiA26E2BtlmxdSSWQ9y8z+pG8
KinOwFnzno9z588f7qftQ1iP0za+sgIFGBJqnGpmg8N0/zpnK6X0LXGciopR8iCxgeYsqiWtbB1H
IDQ0xSfrddvBWa/9pZpAtLp0WFAzoq3bW1H5IGQlQAMw1OvpxVec8reWI9TGRcQba9dm4z6LGLGG
KzXLnD0KwHHYtL3HyAmsnFo9ltBSRYufjLqstwP5JjJeoZc7wDSkyNgxIIakKypo2nvYr6HfPYpF
88FimfCU68UkLIebW8vRimsena4Gao492tm9RvHZf68vNTosmOXPbbvY8/9MEoRD0Fe8ixe5Ux06
uodsfDfICvC/MQGKaLXPzVd92EYHxbn6YcB86SRCFFpXAaxr1td8nr3wvKM9obERIHgQfn+jIDte
cFKN1C0Xmlph1gfRABJZvkmiYlTLNVCnbilXwO4vTaNnQk6M6B+nwmb6N3rtazRU+c25MrqKAqVW
oYbcoxgcuFgszUw4xfix+HlsZ0DnrrF2y7G/O4lZ+y+rid9MTKxwX26l9ev8uty29Mk2I+iVVwC6
5gJP034S1OkSWVOeZoIClJJsYUjy/Fcp9qI3JNqYrWbhonFzAhlwbtr59Y+vQ+3IDUYKJ34I5DMH
LuSaZ+/vb7tB9+PWW2s9LCXK98jhViRkvbJx5d6ixxRBevzI1jEWPVY2nYcGe6J2o2zUbjmEAbRd
gsJrA2kM7hxBIeHRlojXHrIQL9E8GMF6sSlI0IJB+MfM1o4Uz1jGDuAhLPXK0LOCVQae0vWZTG95
m9fJIdXmeAoxFIfptAj07yKKCwmPGHA4sXBDo6geftI6X7ckUNrtCIRSx38M/ZgqIwfiJCZxjlGq
SR1voEg6s0G0CCqAQXfu/ncVDPRPbKGCMZlOduObCj5QD4ryBgjvPAIgYCa6zE9CHNiHt4eO4u6P
RFLpUNY6QPrDXfOuKkTUllBtGAAPM4sWsypuPIfrE9nV28mjbJSRxX+td5B+s0na1rhiKSr+uVYR
7k4/AjaBl3H8XfS3+pdQx9dTrv3lDAAQX/Fai1s2oFalfWCohxoG0V9+4xcRnRsnRFmbOg0dpW6a
qNjgN16/HxotJgmAQFcPpoIavsZbF+ELBZK7scuNHSQfAkXe3o4rwbdh4dIEqox/VrVGWttNi4fZ
KE8gNM3rMfDeb5CzJt6wu2N/hpxqc+wcLmKFypCWceT5t7ltcz4aiviF70zThrB+e1Sy6ZGs0mMG
2b314tgr7iJFQfXo2wSzcWDvbaX0RpmzmZ9lylm8e+91Av5NJehLrzjrd9LfNTVezo/eHKLPC8Jz
TYaeeXfps95jfu6fdecwNMoeCtgaDc92TBRcPJQTP1PjX0XYIkRlVdr6jk9V8MHIhTgkqoolCHs/
fLDDw1N+jFSBeDWH7PPRsJm5FIuu0UbxMlDqhu8AtFE2rodzz/xbTBzSy+iykXouacotqwozKL67
pbqprzU0pux84fiQ4yOOby6/Ll2YuSCN0OfnzPxzOQHSVU5e2LyhSVzccYFFA1vMAJOgN8WIW7aR
wpxLUg6gseera49squUBNxpTaSClW45eBGPAoXY3nQaFtvPM3Mhni4Z7+/+XQSKE5ZhPBYWh6Yj4
E5qD+dTSmpdTXChKsFCIZIHR0DKUYknUVydUnlyS4xh0WfKQI7LIZQV96waLYUhd3fpg8ATvbang
JVLXhKnrhxLz1nyzlwwvan9vKGC7HAd/6XBxYokEPy+gbsvXXqAu21sjtyZ8ZfE72wr3LROzHA4B
VpbxfqdsK+xxoo9zSULRGYuGUi3Oz3Gw2Hd8LHHfGbhbtcdZ5QGOjic7jlkk2hZlshw9kBO4hPfW
DVqaa06PJpGEEoAaqSLnr8iDg1WwXeff+CEw6jRwx5t8jpA/VQINWIIo9GcAqvWVnTHjf8iQRc8I
HRdWrNEu7BOG4HAtsMi865AFA7WJeLNqsTVNQDutLRRWGtG/82I2EMKT6if0fLelURNF0xeZcNpb
GgG0MDzQyJxxCPyz1y18SkGuEZOxiV5MuJoVtE1IgCuKM1RTE71MmekIWyIJNTtfbA7fkDIl48Fi
f0qwoxswsYELFsHlawhXiPRuNdN/rNlnv19+zwblpnGJ3akwAXFfs1uhFzT7HhRfYvAht+peLedu
E1HL8cu7D9ViploRENtddeimUlhWPMYgVfovAhbGmC33GRDZVd/9PWeRa704Pa/jIcNe+5EqKR+9
7D2jmhfCx7lqXCqpFVJJKQ/eV5sDW/7HZT0sB0OB9dybX59ViNqbRt0/Bt2bcV0dMeFX1jpe21we
tAehzkXSCMbahECDWQ8OGPrx4eucyX2Arn9gqvSn5IC9ytSwpbjnOpsiIqiDQyA+XUgApsfqae9+
O+HKEL5PrwnuAoWDYoCCDQKBPidygi6n0qpLZNNF0vqZjfYbPCTwM1P+3sAZn3BihjOQL5DGmWOF
iAMK1NkyQtFLw/B9JJS9lK28/lRX7q2pkEtSS7JRmGzqQRx7HmAtSKptz4tTcnMQsBBh6kEnonak
+vxKn61eC2AzwCYoY7BL9CAbiBnIQTqN8nhtzJY2cwSav+KSGUBztSZnLImTOlvxgprwg0fJWujR
SaeW2/3jPeFbOtfb8WOKMif2TKyNPZmMA4anmPF4R1c6+TNzB4VS0ZachyCEJwUeelu0RVgY+b4A
f84PqxSARExMfBriCikAam288B2mUymW7fO+F5Q7PVshGPKJ39lGFqtHu8ER7bRbZSEpxG/PY7jg
P190unQ3s0Vb1nJ5b3QKZyWCKjLoaHG72eGXKEuYQ/FgS4CTpMKUL4h5nL9PcG6qJQdawToAaA34
0QFQDc6QVxhfQo9iYhsLfJA1Tj6DbOKlYh23nckJPMvmw5EZ93SeURPo2zXQ26UcoVW0G+Sgkdho
0rfiJFXmtbOEjEzWlIGinET5xpDXdc7MMqQqhk1PVBd7e3rPWcEFFlnzEYsgp8RW2ZKt1l1p8/vB
W5MyB8sM1mmiCk3Xxj1dXYvx6y5kljBX1Qx3D/LhVZO6MA1EZspWevxB2xI7MQ511K7/ZebQuXr3
sV0Cfs8w+3cV1YWjMfkxY1To+pc8X6pT2NMWz+R77t0CvTzeyCqpCgnnf8QyBMQQJW+VGqLyspeF
2/wyDXVWj5KSnfSWqFPMVs2LJ5H7nNQ7uRB5GPW6+ZYOYoJzCt1wXrnmsHFenIK5adgRbiNoD7g6
l7Pm4HePZp5wINeadWWBoRY7G//yOOkeriHr7k6rzLnez7qTyJ0IL1bPKSnI4863i7qemGN88b2y
uFcBJoy8T5Q0y7Ji5Rn0ACWJBpFqmkk7vpiLM3O+3k34ShIUn2Nc9qbouyOQ1FTzJmZb4OHbjJI6
O+L5t0UpGUwqCSeHFQ87iGUp+VFb+owBmt4ICuzDM5ByRDyDiUshCHOrJuqiqA4K1hwKhj0ymSNU
2hh4CwtEBU4AnsX8jb2FttsUCisxPR8GFz+jBQhAdJmSKFQ84JiYNZTKHeHXZTE6v4mZkwdy8EAB
DvRb/zuTR1Gz9fhRGhyII9i5HeMTGm6r+ZECquulXHfsbUr/6+GzqnyXRpKsAWlJQnS750OKPojC
ypwJH0v+Boe7GJvHpWbGodH4jco9TFgnxVe0atSpxST8S/gzvmM4m+krRs8kFldh4T2KRAehIW5j
nEk4PWoEj4h/hHxRept7D8IjZWxLCMo2N3Obn4LnM8iMYFGBVC/KV8E/0/XXIT+drAtXHT60oS2M
afKTTT8HSkouEwsNsOW2aQ9Kf8nLsIsQMSSwleB72mGG3WOGLlhnaMINPQ0hKfcsBtfvCc0OQHa3
+m/FD72v1JSZ+qtkvM1LoXE2XGoYySVfZWovY0kDwwHo9SAI+e8DA+6uE9Xy59RC+nVaRC/VY5/b
UgKPtZEAfFjjghvFAbFxs/+DDeOuvlF1aSlXbz9Aegk43Q6QuYgpythbDWYLnKs0SXwJTLrP5Vd1
/OcD7lkCMUIUcKYyCQDlgNiu8PCeh35GgsnnGNaGz5OCxsHzYsKma/W36OEbmxVMXOTpZLxih7FL
EfB03qU5Pax7lyY2q4JiXwMrucg4Z9hwt4SRz4z22C0/Qt6M7JHOKmrh4Na/TfjwZU46OPbcnjuQ
JegOnwW6gXUFO44QBM/gEgSB1cxekZWhAHmrHuc5l6kdJ8f7SOKg14u4DXibvp5UAQFSppaGrBUg
N0puUsaijqENd72SuSwJTB7Uf8X/9LZNTlwqdOi/7cO4sT0uGYdxhlxsHd+/kpzeEfduR4P8NavW
JaMX9aWoERBrJj/09M0GRoKDrCENX3KUax8p7yYJgDv8XxJd2tgoup9Ms83Q5qz+0jKqAPNY9140
QTk2iyRh/mJvm6fIjd5ZYydYCNy6ij1/wkWYEtQh1av4SgURGzuMmyWMk1eveZ+Bu1i3afTq7VSC
DcnX9h5jdwEbOjgjY2u8sXzT74l+gcX6grmF0FvOzW8fLMI2bX4K7p9DyqbFp0zKF+EttNsPMNdL
8wc9BUg7vP2uA/WjQS7pwJIsGsexphxRMF6P/F2bXC/vq3u91ARJibxFV9yQkHPDt3b8H/OisZjD
01IoQqQR9iv8PHSczdYeE9WTBdHe3LfYgW9wyPkATWwgIeoGj46oU4Rs/jI3eA5/OoK1HtVjAfV8
D7ol0WANAwlmiqyglY8777gngjyfkcgPQ9a/IWmb/KTzujvnbjUbLT9EnLy7ypCgDrJxWTXaux8F
huCM4Zjg1CpzPjnrLc9N0bNOGUGDGieoSbD52yKeIKsevABY5xBikg3UPu3Q3qKEODY29SKvB48Z
7HrwPJqeC+jnHb+0hMs/5P9sJpI9Te+OPQGW4oRmNKqv66B/tvXOVIOFPY/osnsOMjSqXRIDCtks
HWp+DLZuMO2+BZBNXBGaxhrPKwWrCat8sbxCcMgo9NbCslDstQkAl/B1IXrN/xphfMoEjpIHMEYk
Z0HXTA8zK18gfqdpPNpmdSF4DO9qobLfR29eCBXRMlTE72rFwE9UqG6TwmAZD9senb9DRiNzsrh9
3QwUCJwMZ+Kw0NEjbDjmWCxgld81LihwKsEF/nIFiAcQSvxaId8Fhq8y6AYSm8LqkhIX7D9hBelr
HjhP6MPPqmUFX4B6HS2YYowk+D3uY6OQJMhi/m+Jfg5uOdRnkCom/tzsBd0oM5txbHKX/m5AIGf6
ta0jZKGePE0Rkuu/t7JyVpgrG3UNrTYnjdqzB+9PEReCkyMgiTVdQRpIkeOZQHiAtyAOLNPlgMBY
3BiTLHXvYtogeQ5fnxWOL2Jkfu4/NkKKDo1Z2Z/iud9X5LMfl+PksJZonCWMwNW8b5PkuDvlS5Aa
aQyMniqenJOsJhG6GljLtPsx2D9GJvpR/Wnxfdd/0t+2MhHbAkpFLjkf4STOkzx+ARwCPA8JxaS+
Nu/pQ1XKHiK5mpKaFgqaTqyKPPefJJkREr94trmPDuK3DP8Q5X8rfNhHHCzua5Vzqjo961+zqHWd
7zJH0uNZ45mrJ0gd7CDV8YiL1+JMBj0GnVmMtP0j3/b2JwS7v+kyQlKpqnoQr5OteTxSekdEE0n3
RBfxBXQIWahCCRB1mOjBcsxKEV24mZWa1lC5vBspnaFSqQIyOgVe5zxtWkD0rIm45yTLATVh5bqa
5TVqlaHQtNSV+MtOBtTEKT0lcXsga2qc1Z/QXPlVagT58bo6tMjg2tOBIn8fIAlYpue4cOCvkb+F
7t7yoMQawV7U/LblHWeEn7aW6b1+Cp9KAQIpQemSztvWDJVKQj+zdxAbn4jaTxVPOc5aXFv0dUFQ
tevckO3Ga+GzDjLEIc8Iv1/yji+4pIF3qW1IQsYpGqjGA2A5sAajZo6IOA2++cp63pmX+Z38f+Sk
hIFJEXtw6gyWgDlsXJY+k2CfLBfbozsNtLFpTncU09NJETzmPGgvj2k7t+nwnwXNsq6OhU8qwFol
jjsKhUlSojS1wIELgW3wBlQoCv0TsOmxSFS8YDxwJzoIdCrLxT/BZLeZYK4mR8um9MOJxxJ16IG3
4AzbJgvcVYSgiZtHr/KhT0A4pz1mdPr3sYf/Nuyy7mZMaxnhUK6hdvpFYoHOM9TvcqdE/h0POtRt
L0g5DE21uF0vrkx9GuVpXH6SII/hhuSxfOCL1GUu26Uv52L+Qesqgo0BE8EbKm0IOb8VLqmM2Nt+
7bbGGkhynyi4yxruIh22PyYVtSCIKsEL44t9pk4TzkaO5ozWS4l90FLHn5uVN2wXJNWj69QRBOx5
2mxq9dC6y1+vT/P09a78EpxsDLRhMDYcibG5jkRIhNsmP/qZsG+milJe2eLUUnYNSNdNICqzH/gC
e0XJ98k2CgmbZbm0G/rNEUXRYtIocxcIzZ3gWdpH04FGbvWevRFY1UOUdfegnG1wfRe322gXwVwG
ZAZbcA2Rajdwxwc1JEpOv6sDMysOVxJ0bqp57/msCmYsVOfLb+yq0oO0z/y3aF8csGcQxNNRhkgw
/JeDxMe5OvbePgm9FViQ7TkyaTf2++5/24pAMQq/vPmTELKE/PG45BL797/jXTBeF+wlyIt9STJD
JBo1hsoX0Uou/h/co7NmwZkLcq3wrjY36te4ZbowwaMJu6nHx8OeVSrnlMCHELBpOIAHI6WOVOF1
XMsNrzw23NseSJfunJo5cheSs443Ky3WZwTi5/Hm1WYWlCR6r+/OG5gYPzgriESBVsEgKRSrB6xg
CUO/NctGebwHKemw9hlJTRvo5F096T0H+R/wJjoMCkge7PjodfnwaFhtuuNi3jppErv/QfklnE6O
Vh6EEvm/hNZmGcZjnT4QROtjHulsvibgo8o6tc4ZOjVpUdyAskzTCWEa/Wm7msn47koOppnzITHi
2VBXFsfvPJ1MdLjOZmVIE7TSKLxgq+6Ed4Sq/u4d4cHBUZtAI8i9JPIfkWlnaashXEg/whEMn4Oh
/6cOOCUkjyrzX4RIX2KLMuZHYbCDTZar7KH1lB6ouxcffW41TGrAkqVbquBHKGoTyfTUrf61JF18
ZkiL/OFQeYnn6SaQjcalKAuhsvrDeiS7TKB99v1LY3shE4aphE7xqhcXbaN1oE8Z8csk9xNGQjdi
fZbf5aJNz28D9aey6Jpf+hsuMih0vsoT5/U9ZXazAOsW1+QsmaULkAsKmSQpTduyJRBQ5X/z9Cx3
1J/BmfOG/+phnCm1RPVQfi9i3ni1XPpsTemP4hLt+vbWx4o0Je1D0I2yGWRZo3gKn1RUGSpn2Z1D
ckeXD9JXPuM/fc4vy+z4VFWvTvwqcMCqWDJ1xaG/GyCOyw4UXA6HkXxNfL/KDGvRQXsKG0KTdEVr
luiETIw0nzxeH8ef7F+DlTf2R5jU6LfLybfxQnDU0wWUhSWk0pSnoeR9wG8YNb44FX3k9UETCzQI
EzsP0U42r+Mj07fTVPu9KI/gaACv5mvUbvnBfeWoeLum3tU2du6Dya0Q8B1j8RbA7wIEetaC09ex
MjASccx/bFbGb+alfaPgZP5M30vwo+G1q/wgtwV1Ed2y0NBTAUniZkhL35I5X2HTSvKBill0U2CH
CytKPBlN/EXycoxnljfxIvqekzsTv5Vp1wCn15Zc7BSoX1e5Z7iYJx2sTiHIEuMJx3w50+JVDMeA
V43cKMgx1+AAIMOfgc1vSflf9P0F/jn6pzN0sR9/PAVOG0isioYiO6f1sJH71Q/IErQEmRqInO0R
q0GYlG//n7JkIL33tiaT6+PjiBBgKBHJe/+eZazm54gpCaObMB7xqbYILQUWLw+EGb9Ctl8rJdde
I5rF8NO5WwZdnDoJ0QVkrB0iA9dSINKk4A/JmqEpdW3NShALX+jhzn6IRl2SonDrrRopg61rADUh
RuJ7Vu/XauRwwZZ8qVx+iOnNsHHPIxhDqTaXQKDy50QV1VOCiT1VYnp/Pw+Aa+qYtBSeS/U1jnYL
+kBNibAbj+E2J3V6bVBZyB9RcUjD06cZroYQo0DQJpOyVfeX5Vo07pyR1fpId8oTSQYvASLZho1S
N+drWAh+eAJkMuvrK2lUhInLPH4oY6D3lb7mhLrUAyKC06XnsuJ2q9hy76FNiI+UQuJ0iLYTON8E
qlwc9+Dz+0rz9cEaYtzX6ehhmrlwV4icFSfxZl/sRsBeW6o2EAkOPFWClxpMQLpwnKporQ7wJaoO
oqiMA5U7/gNE6jYuVVNVX2ueD6yL6l27O/AT7KPS0/yzUNhU3t+I03Pm5p46V10fvzh1RV/J7l07
jAnBS28j+6nQ+PyxP4lT5pFDekk7jjV2JvOOCGdDJ5G6r12vGlfWbFwO9rXZCbQJTwOaI2Evi8Yk
PlKRYQdDaVZYX4H1QzAnqW8YvbcVDnjIqJa1SbZsdF0sGVe5ILU0at09qsprOm7CpQn1u7irfWjW
O3JHvbdqaVjK/NPTlEgq9PoQwBo3P1LJ/rIzVfNtoCiSx3j2jah2Vr6qmg6Y+hi5ZsC4ghm1IrT4
Hw8JoPlXa2yrlSPcMHg6ODipNJfiLHg+JgPwFrK5Zayl8pgFX2oUZeXFgB9PLYDD51PYX0ISyC9Q
VmwVEHwwti906nrw9OoRyzj+4xhJ4N1L+lsozDl9/hmPkc/vglhCRpHuXJOzYtqSgBZZeLVYxc3+
GENkeDv/So6jSor0xpdlgmcDKqFWFRL8aviV6XY6WtrcU+kss2AhB7hQ/CQOx6HUCB+89/igC2Aj
lr/IYV558HFVW1FgSlzo14D7/1XOfW+ecYjOTIS2Qu0nJQa8sAtG4xpHtCIm2gltMkzxrJRroxq6
wN35aWZYg7IfSJPkPeQu9k/KF4SSUg5EfoH+DGOJS8NQcZNzqP/5Ibigdm5hGrrWLiLkvfDN3XLG
apfEA72S5Z4z48tghEx2u2TRWFQj/7Q+ZsGPNUqRExGqzKt6Y4nKeXeQipH3G8chT6G9zK2hBUjj
LbiV9kHP/IlDQATnNu4CgieAucBglYoXqpgGwdF2PClU/4pgxv3jynysLqFdSdn7pDJovvRdHENS
nVhkHXHVaPzaKkm8YnF3rDXDyfmCT7WI7/CtoY6ZwFwSYL7mG8dEqegNzBlrxA9NyHIvA97NQMUi
l0xr5hgtDgFev/336ZV0ORQiOUSmzDnrftq4l//yfPiPPuT/641spfv82tlttKsZLQPt5+oJQqYm
UDaCUD2zl8XbYkYVoGWMNGJLVaR4etNZCoPe4alC+BvoqRmycVDwIDQK8oMB4ToLObiFDyk7oWKS
4ZPQwPDib5mTssTE44N+zJcaixLF+QM8RNF4s1tlERujkdzv2jmQbTA8Ur8BbVlOTB4uPStwGWba
5asFtkQy9o9wgN+xu7/I8NCSGzAQuN2TvsAtDOPmzUG4vJWPg3L58+dIBQdKYe+iN0mQEHtxbZg9
BgChpVQAM6poTO1H7VEUBn5mgSwDAvoObiIrhPJbYu3lOg710Xnnj8tJ1Ee7mDSaHwJ7NffTrLfx
Jmr5ZQJZ4qW20DbCm9/ZjOVmKESOM4ue3KhQF+zc/nBikn3IHfl5ZBCnPnFMVNzbjcPzajyblj2c
q6v+ACuBF8jrjYyJXrNDzAZhflom94OyPAZPC7zJPGVQv+VpwBub8x3AoB+UApqBIsLj7QRA+2UN
NrSwDUswT+I6+s2pk72utHsSSDpJy8bO6jWCRql6WvSMt/uhvCgCgq+xkBpwBVwch4KG/PVaVK4W
sCX426n0gX/+nRajBTv6XxLBfK7EN4ymNUo/Q5hvcOCMoP8tJu2pgKbFCNWnqv4tkTkBfN1YcHUy
VAyJ6TlADYOGGNPDAr2v8xCXYzI3UPWRpAr4lkk/Ddo/GMpSUuxPnpnGBlhLnP0kNXsVkU7I7rUj
dWINAfI0zhhV5TG1pt0OM9jl2vJJbWe9XE5o6di3KThjRVal+6NazeYdmB8dUMLijpCXsr5cGckx
YurFAk7N5VuVgcMesojUl/15xgxatjKzP+kvpg0cEqqI1C11q3Si6ZZi/kZRUMw1bhe6dxtmREU4
LXNtO45/VNjNZV923N1KTuOKcSXuWJChI3kQnYJo8Xkm+5+G+bebDn4yDZD+cSUvMFJCVz6u33mw
4thxqi+5pJ4aIwkb4BKEnbz2emdeFPC2UodU7YoEdxzXn++65X+6R2YsNN6LFroZCFs098/9dg0p
unO7DYGuiWDsSHpU88PUfGbQvpDsQX3ze/E7rfutNVyWb/++8nwK2NlI2Te9EBDFh93pUco9Cma8
CzVzilWQkYTDGo1zy/Fljsawxem8Rli+wtzq+oZvqnCJ0GmlULCURhOpdY8nMB4qFflMXVrTmuBd
cj9T6RySI8LSh/HmF9nD5VB5etYAutCsRWPCr+mWDCtqBo4rRI9OFrdM91HJVcG6sktKCOjsj9Sn
C7ZZIdFF3kAPikKH4n/tvROSLW0A5zDfuXqSjRJd+sbbLn+mHFRiYqA8vuXmLHiPUsOiVVROp4K6
Mv9STZg7jmrB2z6mG32husZoS0Pi0vXWojLvmDvvfmHeQt4t5Cnz4xzHDoJOAhUzuqnwn3FUBZ7s
K6ARd9HH6wqxM7AoafbK5fTUNatfiizPKY1DvM3fAeNtoY8A2JmLh51qSxX9x67K+7Sxxx7Wd6Y9
Jl/B9vUm0T/9hzVKlQZ7dvotx83qvkXyZV1XwREKDMMIMQNvVwWHEUcNIrhWgpst8ygj6rJj0fbI
DCmhaSfL0mbqmzIHyEw4a4ub6cjfBa9s64V2yGSKwbYWp/DAEeK9spqtyrmBy2/nxYTPOBiyATlV
xg7pHR55haOjRS+4zQ8cmGZRHYDHQd622PrUQnkIX86WvTHFAKqQ6k52rBpCDJ9GxJowSRXE/wcB
aELd3IBwGUmKUT7NLMA65Gg404s944zyRdVodZvIznoRmv9P4mMHiDoIUURFn0pgfKKqwcOD9smN
s9PTxVTWsRN2cnVy3Apej/hPCYFdKzAT7/fOWxf7VdXJHa/YP/sOydLoeQXIHgMdQfxc6cuVeOR9
h21vyV2t38pXi+sO4MUA0Abg1ew6pB4oW7txDTTLvEnKAEEm82XEIKgenJpMkNrv6JKfPhPB42dg
1JKy7VVvYjqLnTRwdOBpy5apHi9HUyQUCEc7xMWzsJyUiunua+86YLhFXc70Shdx3RZsSvEH9PSK
L5fW5B9bpHLbbOX9jAe4PWSwIyMBHxlQe3HWOkguqcXna2tzxW7Kd9t6lclShq+L7wpq7OQG9DWx
qjywM/8JwXMUg0UkJ5lsQlJWuRMFJZouwJnhr8zX+b1en+rCzmRHKnWNZg67+IDoFRCk14T0sqe9
UbUiSFqJn1smYnOO3tj66QeLYIz8uBlZbm26SF0ZyyRwL0iGfaFHfbFBnc1KDmsCOcEzAWyXZpkx
+0vSL6EN+4qZhBX6S/uGnMFdyNCCk1Ig7vSeyMu9wgFF1xj5cQzXD4LRNhdcZdaO/OLBTSK8bBcQ
TdUfXFJbUY7o/wV5NQKOqYzsNw0wWj73nt81f0kTkT51nv+P1a3L7E/tgEgwWI7G7yQJLZvwTDe7
xgTZbXLXX4yETrPdGweXLbbkbeQloBIeKUMk+Va5VWleqGgsaX+laiVe4Lc/nrK+R6/pw+h2MvjH
JrMi2EjQkx+bPCkApf1P6lY347UQh7VGnRCb7RVeH9YV6CzoNYCG2rHZWzQvSutW4KMCXAG8Ou2C
2B1oZl1eLdN5v2OI7qq+kOwS9P5s0AZGX4u6M6b8MYrlpjwdRJObms8ZfA4dYeGL54SHkVSaDS4M
u8eOaAtdlKWI95hku/ZFEvK/h3fMvfADZrUcl45kIrR82J8BsJsplYAqy2In8b/5AJNHSO+R+K1t
+bxx5i6JE5kOKgVN04nP4szUjT5q/7N4ydeURsgFwKlURUNpqQcStELaX8ecafycGepKA/Y8Q7x3
z/1vLo7dXxFTghGMWvaJ4Ftu28WOT4GZRapN2Xytk/Nt4wtNnFWF4KNk8XNnJnJ6N3024euoBgSe
SyGaIqnFEMugCXFWi4/V+SSlHz5l3kx8diUrnddNtVPI6oCMz7GlRr5H0b760Hw1rLeZys8GeVea
JG2FrjqlvJ1FDhNhSIZ+gjtMKLr30Uu50xv0rftaSxZ6Uc0GwY4sw5D3hHTdW4rCBBP3V3AWFg/a
4A4bh2co3Z/NdQMEj9reuWn10U7KRcCYxRvBI9sKvoUX1CNnnTDXqXmZl+Cg3EleXYYGSiD0RDZz
eaE3yVZfUCr59vurdXrqyVvqT9aLduQVgvtrNStZMmZ3xFiHWaQ2raXMuVnTe5MoXWEsKtvJt8n/
LSU3Ue95nPeC/ChPHSotVYaycImugeL5xMFR6Qg1MV+XJUHN36Nflh5pQ+OCcJcLOMhRDj8qLKHl
TJvBCR5mwEUQZzXZbESHpTuZTRTvrysrdV3wYDfvByOExxTIrAdNFbbYVNXdnsmJXpvoTk6WQ9Z9
DFPxo0+oirkkyF5UMj0j4OP9TH04ogNW//5pcp6ZSqrc03SP+i8SvQjJ34Py0U7WUGsoPgR7q7zl
DtAQ6f/EWYn7772joNIru7bazsEc4PCgyvqaMqK+8n03jstbPN8Kv7FWH8mhwqJbhdlYHa6gyRZO
1QBFo6HCrLxWDRp4ShOPtb0CMMP2E2G6yfXFlQgjLQ+T0Iiezfi1cUcuKKpTuaeadH6K8v6LD3Hc
VwYbAHmBXSgkDGIeuLomu1g33Qb18xkgx5HEldgviLvXv8VxScTVWDIZ7jjMh/sVnu/yb1hfz9XF
SrD07tIWlvmJD2D5xKyN4DSD9h9Tj5WFUNzILyUhz/PxY/m8G4/1eY7r7iwT5DqvZfj4Rv2teXfF
9QETZvzU2RERhmrj7bDCnlWSXQQJWGMfvWGTNXgYhKlsE2YNkV2bN/ZbivR/FPkbNeTu8moL2BzS
Jw/8d9JeYM+pAkcsG60wsibI8EH8f24D8N2DolqdihTc+mNjOhU5O1AcwOGViGz5x1B93XGCzwVC
rQbXgYxj0graQhyqr4Bxo6Ll76/1ZxTBavjBRqlxtVaiENxHJHqPRLONtgoTIkVENe8TPy2h7WOL
Vzi0eMHbsiPm/2iFKeUQ8xYyppegM4y71Dskd61ENgn/A7dG04y/NkAg/TNGe2lqs79X7x5tH0aF
Qfht6/tdophBkFrxdl329ej7TeB0WoHbenauiZCdWQEz+uNAswKYTaNV5iTucSfh7HMfGnzDM/Wi
EdjKJpEa/0/hLUknnWNoLh1YZ/wk4e/KYRHJ5gq+du04TDRKAK8mgYYzxAMxvR9H0J9DrkN3mAn5
N1o5w77Yto1sw1IwpeggzMZxAOSQLJv7vetM6zt2RAq+qtQUfX3Ptk1PAuDO6Qb/uiRdELUTPmeF
y6MuifE2jkSjLuGlYWo/BuEpHUWkDuq1had++M9ZKvvKMQ1ugXXBPjot3G2DpZwcT1Lm4Io/GqNo
/O0YdWSJF8eijzzBx7Qg5PFajx0jlJdFgG1Q5OxCqvJxFhKjSJm1mtnQ5NRYQWA1JuzEFjLTNR/e
sA9acs20QwA7oKdnqtgyd1k70X9u5zfn7LK+V/nIqGzio19z4MA8dbfkC5LxJCpCBiQslqTJGW7C
3DLunbjZcCadk7Xq4svh2TEufgfxogzSDNOwLyGxbEZ6Ni48cCP7Ebmj61D9g2kfurmhOEZEXORN
AP88gFtm2wyOLabW64crpFPIjAkzPVkKBXWNzuh/xDxv/8ib7aUYpwW1QYEe8a1+6nRLBcyfyY0O
6WpssdZywc5L7LWhxxYoOoonlZWcIBZ8vusPCw5Ep8Fr2EapYz5rR+Ba6cnZtwd5xJKvP3dr/ob3
84RLmTbQqK4WOXRCyCFQWJgtFH18kFae/X4Zer7GngQYYV11Keh/zmRiaoTtcXpg9FIEIlxhjAFh
n81rmffc/8fNqeqDA72JjN6UT17NONH3knvkEBR+KIfRRl0i9PdwT+rsv+29RktS/F3kfnR8qdvI
lRXbiakCN5jR1q8hgTR2Lfr25jgaXZBSI339eNEE5DbR9zmyWA6UpG0c2QcMzPZzX/NrYROec6l/
KJwsIK7jq1U7Lg7X+OkmiSAjGJmy6GZfKLyjdiolKiHS7VpAObT4jPxWCVqdOegjEiBfqIuUyL2w
ERc8J2CIz/jA372x0IvKFh/yuOTuC6Rq7rlAaIAbXv16NMJWzmKOry3nvcxLIL+ecUxVJI4h90SZ
pu/NWiEQugL89afPjOKUGHcbGBdNqdu2FE1H9sHpdgZEafUiiSzw9EY3r9FGcSf2G2WqfgJucbKT
CHUXcAeDg5U8wMRa/UQAheoY++sWm6wSH5ITflpoXtPR39Xh4XFUbpAC09wATe1ofB0wZnj0Swia
wCaoKghMP0WgFqLjydhf7vuFjvbPQ73kNfG+IXEpKufZntYeHCjAVfdzakomnDHhqcw1Zj1boMV5
Lb1skn0IgCGQdzLAMYSO3QNXKuFve93/Xuyp4JS5XtOgtiW1r/KHBDJ2fibRXGCMH2EKGKmn0IZq
MF3U0DG5ROYMuX+ZefxxbOHZsCNlQCGpddQY5VNxhsiD7GVZ3CA/AC+57Sjv3jhmtzzIVFoSEOCa
S90uPjlyw7YtDKQ4+EdqFs+kOeHzQ5xA3aizP2424xJV6qOMhj4QiHfo4JY7nCYvzzwHNF7QcArY
OfXCni6cJTpjzvzrS/Pv5q8KVd5SrXaZEcmzFydrQNsHRDqp+2tteHqjqZx455ZOzSiNb//rSko3
FyTLyXCNH5dt017BZPeIiUssZdAwmf7sWv3BtNGqZ7y8GOh4um9RRpvZZVn2+FVNTbms4sZNBjQB
thiK/JceJ/PEhuGNEDmjosouwi39G9+4YgA1RY/g2jT3cbacbLwn26yI+9Tdh10vjDAgEzuWPSuo
U2xOjA9dnM0XP3mdOZKWfdAGFlpaRGSdweXhVDsbLE7RE5DI+aOkygeNzYCZL2KV+as7fwU2polf
gP6H4fr//2yIkBABKGJ0zqAVW6f0eMVyz5KbTQ3Ga2DNaw6RGrWDMgNN/OJYulPbMngCXfj93c1C
ebdnQkbvwT2xLO3sRTeSvJLi1Rl5RIg+ack2mo/oEL2CoFi2bACkk2BIuiUq5lm11n40DHxrF5op
Kbp9GqbdSYCVdIwwH/KYlfttWAwEsdtk+L4djROV3rcoIlKU+ePcSlOM3nucoO8vrWJSIBrpmNI7
BzKligTpbb1nYc4c9j3nQLq71Nt/jbpiNnrQjPX0uST12p0GUmiyR9WcNablMZ/iSVj8kM4zgpJB
E6UDjpjaXGMAGEWls0+zIUFMjUqljJGvYBJapj4HMqv1cDsJ1Rh/9nM/842hxw/i63rasyf33Noe
RwWXIKcHqqGojzE6inMyCNwVDwuw1ObTT+O8eAqMVux3CDGYcFTVP/P4q0IcgzrdQekGD5x0NuXr
BWLy9/VMw+LrMaP/aMHkkCv2clmrazXv0gFR7fFlCOP3OGsopOHrtoikGeDfkGa1EgpGYGJrYLGh
U4nR2X5CSY6mcqzP1iV4/ajMkb6v/5Oj7xdVpTpRna8vAEgXapiTDUkOsiHEW+UPv4FimmCFgo8B
yZFGy4KpE2XHY+wgLyiy9NXlB9uMYQL0EILp88fMQ5t0mrbvMjst+sjHat4EnsRbZYfN14WN6YnH
Z5Uy1Znr2Juze+TlNdzonFaC95ePPdVFZIwj/C1N2kjRWOUFzN6Q+soPNQ//CPsMInl8nT1MhWOM
zUzP0DHcbzWBN9w8gmaNByTpKSICMXpoOumJjOizjgAYwEO4DW5QOUh+7H1AoNCHoPbsQEJqlR1z
LkYLfQLgccysDXVIIbXB/WJudYo4mhoPTDin+lRYxWt+ImkV9KtJhxYxKJ4L848ZVloXsuNdDAzV
9H0CA8vmAqzutimf41vim1labYRs/drNDQK09ITSJQSrEMP2GwufuCeMfC/Z7OdplNbDWDtuaOPC
RhYBegzjuUo94Tj4K4ypqurvLMxXSq/uehWExxtAcGh5wqzb0i7q1fhIVjCsvTp9lmxozHGAFL4F
sTKIm4vgvICC1Rg5Y2HsHV765JwoNjExL58W4rWbysZ4gzGbWuMWE7/GZ6kNj2Nldi/Q4d+hPMRU
vreF2ZpQMrfDp4y4QqiO8oZyavgtNCdSdvcFYmkhTC/5td13tmkfwERdawjlRGjebYjabLez5Pwl
iDwo9t+xn1uzYajLQKo7BDiDY/5oxnpG/P+Ox18zo4FfV80nvxyLffr/1JF5fhB01tFNxL+xpplD
Sf04GG4ogvqVi6EEveeD8SeaYeuoLO6sSHxzTaI+PiDbHzcGO7MPjRmnf5H8Z4f5SmxfHX0LF4zO
TGvktumIAv6pVFsyEPkcZbDSjlZEaPDd2EsOw7bwMVNKEBtstWCugK90jWchRbZnqLOmIuNQphgJ
zLvPZE7aOPZFcpz4+ue/aMkZ6Cu0Rr1UEEVeFnWHhZS+Qx7rCXt98VWzFFfY3ahNX/nZgXpeVJR9
UCeAS3/MkYJpnzyqv7M29+ipkGxnFOyd5+iv5zjPsqy4hT/kdVeVX0B+aqgxtwqGGm6RqP2hO5fF
xTfyY7mED4UM9PlzfgsQPMo3mpUL+TJdCcbxOXZz62zXU54VIkWd21tDbxL09TUPV2Ts2EQvgeql
5T6vf/OemHgutce7kR9mYnwnU2i/HT78QGdmlnrg5SdDMTwJZg4ar0jypR7MSPcVJsuke5yyWjlQ
J4hCzOrmpYRj7LsacmhQH5EQQwn0+Ex6u8TdOkvCSFjaeTSVkfhp+i/+vrMM307O2hknxFbRuKpQ
BhF+VNStuRunReJQyQoRfkhCxH3FM5oeSIjluBoVONecL1wM+0tKOQvav36kqwLWCKr4xb590B87
E3NAb33g02VN0mZle7crvn5gKVJHv3RwYn1Uw2Xh2cNBFOmN03Eauo9qxNkmWjsN8mmjIwlBs+Wz
BUfHWkicVYMwD5Flqhf4qOQWPZsFJhPCMdX0Kimvg8ZJscJKEoKyHHW24T5pki0832NwPzY/ah9D
VWW6k0XLiH0PwwtXgimsVCtWWYspYFWkelhGg4rUmM5e4ZqqHiHuvF+1IfIssAhxpZb9cIcWywBN
TFyb0MerIl970v1phP7AnRjGCm7nq7QPmqciWiMe8XIKTDHi00+Aee5QnHRIljGBJbTsDhhszY29
OeLG021lVrgEVq0DzxDICUgaxIOme8NinpJLpIvkTP4cizB06zmPmiCT0UzQEGyGn8k3b/yxUDJP
NCBArDw+xzZqZEDD9mAv8tgcpM+YhyKbarV1GQtUjPGgC+zUX2jgSA+2PgXH8ERrc6ujpPo2mrKn
Q1sIPlWqi0KOImGG8oOYsmj/IkBgK7uoENo0HI6iB/RWo4vhyC86onmAt2Vz6+6dcBGvF5TCRTgu
eKavpDF8IsBTVzj5VhSrQH5Eoeutl/wSfJSl05vlRWJX134OGXemPFvc7IV7teyTDJxa2Kc6CC5/
qRQzpOwILG+lLtnfYJVefP8bxBrkuqPTZK3DUXiqNlN13TcSDMnxer3kL6RDcVi+oZSSft+IQBPb
SmRuAkEprG2EsFHiFl/XZidbmIALG1Yzp+gAWC7C1ffrZk/ItlvB0AAVNi/T4QqI+jx409s3raPB
+YuY53m7U2HULOYwi9hetF62T698twnHnKr/Qs75+A7runPJsaRoMrLRGas+mxUy8MlT/lZulDUt
0bd14h58WVJKHKUye3tSanRTxFUZ42cuFaxtFiKE4EK4ehW5gWvVdo/HdIKC+su0eU/CH6hfdVyX
SCAMrZUzsUEsiTbddz+ZPlCmlBaD5YsRaQsjAgkl1aA+vXAOG+kwLLfaOuIkuwtakTpXzgY4Jn+/
C2Xe39UAuNlh0HImIstWUOUamN2tikyIMNiPt6tEuUoCnXJI6dII6nKwhL8XlJqekLBP+Szso8wS
W4hASxui4HEr0aTeub7eGr2F2j4eG+/VD2/IUfy+P1zt/IBvL1/Cswu8TZZYwmwEHP5S9bgaFV3j
pYKSBptij1Onjb3loRmHFAHGFH3aqqoYAYfIycGOoEdky6ndFJW477piAy2npl45hooraajXE3Hz
SDZPnj8bhfopB8T8WarrP1LxWpGKvACF9tPe6ZlpNzpIyOLiSgEJEagJSyk4rS8tQ8oeeBUUDxpG
zUjXvvO7z65UwfCy+566sW89+8+0JBE6Oxakq5iqNIKPeqXY/NQfaF4Ihd7T18j1Bx6r1PU4/Wwx
E1K1UApa5icr5y4EOtMliR45i8ZNZ2eXn/S7uiGzsK34Svi8jUN4aTcRIONBgaFpQIyTXiwpYsTY
HN+Y5VrwmjvgSG+rbObYlvJARvqCYfIg7EHOZncpV4/G2D/G5rZ5qXaYwxFdd3ec4M3X+Ed00hGC
AKjMZAQR35UxOQGxGe6v2pgWtUAK0HDnD5LN9ytJFHiHO7x4l1nMreO5vpVtkpeSV7CYkUJHv3QI
S4ShpiA4234Fy3uW2dZArVWiuPLNJAsvbXFAiGgHqOgqRQuCC1cNNaK092kxaqvzwo5PvseTp4tR
vCafygH125iG8efjMtfxqiym0YNY2bWVw1/lZQcQweJ23jIsTBbyuTDV0Ckdx+TbucaWSD9Ax2yM
62uakQE8NeCKgl//8P4s8RtNWpafgdYyq9D9pUNmpEAOoAmgi6NxbivFd20SUBSP7dy0wI7RnYxs
uYTvNdD3p00cY84+1pTj5ZF6tKlcOH2r0ziO6PcRiHI0rKFY2uf2HqwAoRuOI98mtZIFW528/29Z
6psDF87lJPQ7SaNL914OuO7LMFQMEvvWv5Y8AyKWKfG7zk2w3mMyImAzwggbvh5gAUcg2bf2djbD
fnqm8R0tptRZd/dnJneLrntCZp5oTZLYvXY4/CkPntDJZHA6yJIfjbF4tCfHo/WFS7qVEUfe27y5
zWZIlrUvFM8jO9I7gFz+jQSYXsjuOdg3h67BIIlKlN0kzfr2613tHrjjpR42WgVPgFKvuAV3d/VO
l/Mb0tuLZSI7BKDRjhkJx2jT8hYhxxx0fC9P16dtuiJf4EWIrz9UPQot8RKSQ08jMn/ijovALxpY
3hVbF75oqGuLYYYXr8jXqnEYs7IPQa+0YV92q+wRJVWbRX/StTpZvhjSSawDFHSzCTYDY2cBQ2b1
o2TTA3jXeBEMbhO2ObnQd55hWauK+duwlrZHXJXr/e4T3mBcz81CQPVnluosyvecNSLmvr93D5AA
7ZKDbJ474r8aTJXnCEXd5SgvPMOKR1Co22/TmuDuc4rrij3Z73D89wudjmB7HZq2jeHKkoHNorLK
oUmPz3Kh1Ki5B9sh9ecF5ubMWcm/d4qeDE6al5JE1DHaUHvskgKSn/NuVwRzN/qprajnxLjc329r
hITneAMAktN4JlVAQULy6dBI7Z3cVSGGkQcHbkA4lsjx9vvm2Fn7FuWuC89X3+Dv0Rj5rY5TK8XW
Zg2cyk3poqHdXVqOpT82i7omQ1Gv4vXsJsXS83b2638ZEDxKQuU2GkPjTyZtPZ+/ZHzR5EhvU4Ic
soixz3Q1ubr9jT3aYHWfMhxMXZzDNkQCF+a7WJ3x2aUUs/4rVn8NMhEdKGiQiAkhUUoZ0jGngF0f
dUIUZm8O495cSVoqlssnLYa783cgzVdS+jz31yzed+6Sia6Rp37F+kIg2Lcjz1jvx46w3TNY5mF1
3mZYffYz40ei6/Rz1sEKrU9pgTFrcrN/ZB4JrLRb+c3S82fZZsFfGxClW0ewqkIop35/VBw1tVZJ
zDykgk0FV9zassg0N4RUJ0ROx0LpYcdozPaTlkPqhs54mG7NxbvHSP8UnZNon/CWIv2gMF6iqmKN
0QnVHouM72RZGyMx7O0rV320ZCvWxfkpGZ+k9u20GVLCL3L0lBME1YrFnQIOsIlDnZ0poAtfmx9A
+79QSzGrUVTdT92lldZzey+N8Wzchpf7aWVEGArw7e1kXwVJL6uaoq0prwlXll6C/jLZiWc2DWUm
gVDFkVoqyncMmh00wMRl9DXp6K3XA+EnjXOGllF6LSy1x9li9fjuFs096cBINzWRhxCJ/UEgYi+I
/nVFb2qEYYKJFSebM2ZkQKbrMcEz4RffdDJ9EEMPZ+hIXfTRs9lprWeuoGr7aulAcOkAkE3XLcuq
QFzdb5dsobLsMOWhC3oNtwNRAqmY+vi2tG7HSA9VAk41iU0ATLDojqtSM+OoTvaHKLyks7YggTh1
Pf1RNRv/6c5PzpjJhWqAgTTNJMG0Ok7RfQHhw9NToX0NYEf/dVvIu73mYL18t8s5mQuTf5uC6FQt
WkTPNdHpcte26Ij6h5fdFxq8EiePK+y9CzA4HL9ZsjWP5F0cJjPZ0oF7Eg/35u2QRH5/4ogdglu5
WoXHFh54SELJr1JDhAr2w3Tt7DPzBa9MrvgesSf3XRB28xssMGbwLekeqRFs/N2PhZoxsE0F8YZx
wSxv9uGkyH+kExyZJevd7mS+8GYOLCuqJkqZGHxIwd7Enq+HVKSFyJvrkgf8L18Jof395QlA9JmS
q1+P9F/tydGEIUkgt9+H8RRMV3p+pz6Cm7Ro4WpjU9lnRZ4DBxEJvfx4gZU+9nLOS0YKsBpdRD2G
zO3E4hyhMVKsfNgNTvXVD3n/8ty8lt7SKv/oId1gV6bHPvRFboP8a+gOD1ILqJX2Q14AP5xSB1tj
6216YAMJbdIV0DuExCSfFr9qPOkULyPqr+Q3cR+np2Nw5/5DuVTkHmt5BDFyYmflnRpxtiZ3Q6o9
zZm/nzyhw54+SYYuCCXJI7XHT9/5c3WVJVcru0oj3+FTmk1LUufTM2sMuQhNEdZmhiAeANmowY+l
5NE4DSOdTu/E1f33J9TTPx7i+uppxdyzIc8d2o7EZksau8h67NUzSJb9P5PzSiqZ9F0U5HIP84R0
Iaac0IYbBn2BJTavgA+vwWR5hJsfhq9puqIgRlPXRLEuTbWeKYASaa0DsQpCAfh1IpHyXbgj1Kpr
5Ax1/hI4DLiC7a7piUyZwe6ZajkdkFlYakjFCY6NW1nXq13YF0YH7MHMByKYwUoHHZsmPQluE1Qh
hh2t1H9drVuinWkp+JOyNRtqRHFgv6CD6gt1e6tkdDLtzwFT8pbfP9Df89FaEaTeS+hC2HjL9w+H
5953Dx+miKLt+8aH6DJTnlIZkv4OZ5N/AFy7NT9SPdzFeujz/5d2uJe0QD2qp47Iv7cT4o4sFeTw
X/kdMMHv9zykHgj1dmPMoeuyhRvvEJ+zKSgDHa2gfuW3eR3bEjZSIzLl8T+/s06G9My9zyDTVm5x
tSVx25ZXrhew2GOQUZK8i8tbG5kQjeT18L2D/p1s7wwwoQwNoYpch9qPiR+6kiL+24FT2AXFNJmT
BmdVBZe0OkeV44UxHLuBRyhjxHJM/9GQD7Mr1XtC9wiJ7CYoGu9LMmsdjjmmdwDIn3rvP9apPQUG
9ugzs/YiX9WGt6rzMtKIRXvHM87ECEkO3etiucE1KIFBU31ZMqpFK2ML+Wmr9lH1le1WxLN3Oxdf
o4lRDLnz9nDFxaIc5S1/EeMlokl/atE2DYFvzBOzFqlyRvtX4385jePSwEMdnWuCC1y4vn5q+4kC
dfDz1t57806zBpcKc9h0LmRse8MrYus3LdzWNCvdSfRE0i0KWtMz1sdQNa0tT2Srsm3QPzNiwvA0
4HuaTLv2s1/sxcLJAtlcaxSBiUAerQVOuzmtsMo/m0oKM+g1Yk+L+xCMUDlLbwrQoP80+dcMApvv
+IDRb/1PV0uFXCa77x5LBxzcvnX9Xf6ZH7lbX2AajAofE43/zJUEXQXXWjjLyeMSvoCF8DS9cV5x
VACjU6qqh5LB409oAxiIPFTXpHfgQnk5bQ3euGQAGhY7bwI8Y4WiBvBmk3GCirQtgANtSyoEfNBG
bWzA4UGCHF/SN/VHWU5eekOj1JuovAb60RuUkT5r9vZ+NV8YPf/LsFjcmue6YRoaugVmBNIlEJGp
1jsvmCR9EK44evqNblRyxq/FeTvS+090ji7xu0sQBgYA68D+WiH5MGTNHJrq1jAaG4YeqD2ggxaB
2yS6AtujHh7kmtrN/P1umzPGoRQckfCT/dR5CMIdePF4GGKNsmUvTmLirUwI09CH8zW7p2PAmke/
WZ6AFbQTI9x7PaW5+NDBPLRA9HbFRbhKO/hvEdCx6M+talfDK3FHy8DpfzvLm3RpUYr7oFQf4M9L
y2UAg5THr1wdf83kpIhMRvF5ZonFe9OJ0F6xCZ1ClIlPrGezYjrfNpX1TFXbxdjOm7jK/FCcU7FD
EmFVS9nB5+la0y5X1M8JpgNxfibtCPBV4Hd6aPdyVYf5KZLbU9uWphYPcT53KDcAW2ZwbM+C6Jcv
bFvDouGkrnN6f/5fArHgcOKvjKA3IFzeBt7hwssUnBLxacuxoAAgN7ezokmTLkMrIyihp+lhp4jv
B+iNsVXS/txesCl2Wyx4IR32Llgfm9i58d1QfQ0+nWxKrxL4gYttEgBLDCE5Q6gxPjDxlbHt3qkR
FZZ4fAsdG37A9GjJf6wBo0LvFj90VIufqiD3/0GRu6PpXY8gVpVTDcwAnCdTnURgbU19Q51EKK6b
dpXC/8i6WSpc73S9NQSLDpGibmzMzVek5KTgB4yVMBUSqCm5a9Oc20zicRKbfBmIRDjMnpaQTeRr
uzwCnTc++IJLQR0NVTWmL4oR7n8jfNnKEJ9k59z801iC9v2wSIsuLgKq1m49w2HEL3SenJVbD1Zc
8HoInCp/keI0Y9+qwyKTRy7y/0ebW8sz0PFOZr3Ad5oPQa4viubvFFcT0FZ6LjmOawnaJpcsBCqR
uaaLd/fAdA8eoauo1/CbJU/LHCnWCkIduJI+o7bn/I4SYy2FiC5vH739Lj6P5MVVyRspRoDnemCh
sgZZXDlxOxloJt3IElwk/XPPEnOb1sJftx9S6zS/kEAlNPeI3qKInm9sPpVGL/NX91z/XJsoiS1+
QSTiZnKc5nzrnaGP0E9HVkh9711XAv4pJKc7LB/a3pN16KsCLaaBXmpqSHwecoNmZklGIOYxJO0k
xXQ461Ccl8uWoIwt0JcDtaSYl1RbGu+pWVGZlid5TzV8CfcVyx9O6MrpD3cpfo56p4lFB7Ewsyuy
+Ki6q/X8bQGyoTHrkUsaFgbjnTXS3+A0QMUdx8cSc8qljJiNJNC7SgMR9qcqQg7Eskz4Yg9UPiqa
412QLlQY0RRRF/kaOSL28b2Pq3ds86EKeS3nweSLSl+6eVX/A5ay4i/TFIb2gVXXQz9G0A/6RWr8
GD6T7B0Dez3+CZ6eSvyrYba+6lHXSAsfpzXbAt3aCOv3aRN9WFsus6ZqXtavLCx3jXnSRPxPLxSo
+cI78/4mMfZyqH8MQ49gJWkOn3uE5msF5NcTmilduTptmefe95ccl9ATSlXg/mFlkiPeR+a3o60R
pegvraeN8c18IZwTC0ZEgH0T5MZeXO/txl+C2F489HpUBTBtLl2MblY76dfV/F2XabvqMPdg4SKe
4t44jVjlerIPJqDLntGmhqze+QjoYuQ4JE9C4fthb171OV2XpNSzjUuEs1nKeZaYLpvk6iC6wUP7
sOF5se2N0dVz2BExsiwvIYGJCb8zGVZwiXDVN54CDZf/55/V/+qsvXoukH+m16B7tt8HG1dubBlx
zD6kGMq/CjODP0PoTR+SZHXYFJSIxJb7dZnaISWX6wg1D1Q8Puf4/JuwowhSVB6tOduHQerqoMQu
ZzbeoqCpbeae4Xm1CTuNn4509SAqEuXldUe4WBy/zYPmMj7vVIfIQ1vIlbe3ouGBCZAGODc94pvO
q5/OCAVYN+rEkDnrOYomoqObk/PgTgQ5MG2RIA1iZ+/ScOTvqSZdSwjZJmCDvge5qy31ZZ/Dvxjr
Qb3ABNtIGEGfMgd+vrgGrxUXiCd3KuHCQNHcIXTVncZZkVaJmnMMa0Rzw0NkCLfWWT6xLFZQ1X2/
oa1RAQYLSiut/i/xi/+vofr23Q6+kO7xHdpjqHZnm7zmzZemZFK7gCA+q6U++BEfjeUJYupEZzf3
FYou5RO7v0vuksErAo+hGFwbwyeL7gA+6CtfDMNFr076S7NWEVCj8nklJfd5m8wf/NIiYXbNCOAQ
gmdgWF8nO9iJBnl1Fam/rgirQZZhJmBCh1ctrSizVdlLhNHMdypD81dHttJJLw1+sFGi4sNu4+bD
TfFS8COAkdx2r9Hb9zG5Z4HiewmXRXm0TNxiAjsW5b/lJc8egInbTEU873tAo+stzuvxBl2k+Sco
FsiLKKPJbJhaV4vkb/YfHbPVyxcKnWVlmeRV8muwMopPCFIWH8KWpwsuUTEpcwRQyYJEzZ+Q3Kjp
gKWEBR9LPe/GZPnVEcEgtDaPXcUZUB4+qn79do/0JHsziS/D5/aA38cZdxQsCumGlZDuVRaE2IYv
vjccrjcf54psGmUf0E1wkNdR5j0b6KC+Q0bG0ONmHoSpaf0CqjlUDBOpLh/Vbo0t4d3pnuvvapZk
hNkIKdKso1LyWLKWNzRZeN0rdCbUuR5SeC+vaxK6PsAToDGMmqey3KM7UcTnC9CnAd6qX2WjDJxG
6Ap/VD78RYj1mvg7eWHnbQUQPYnyA0ZHv+RaxHyl6R4zMOyrIWa1JJ5l3NFnZ5zVGH77b0+HNB3D
F81ss9Qgm29nNF5Y1NfrkqMAZrHeYMwaaS14OUsQ3YrDjZ+5MiqFLQOVASckBeEdDv4j0dM7XtdG
6S4OaTSFQBYn4sp4L0gIJD234kRaaZ7hMediI9c2Vu2BaGDDZpoa1dIF+rhBcystKsHvxkGFczcI
+z57bMfXpvbnikl+NSDNLoAnu5KFi0PrrW0fKmDzWi3SJtuY5KPsCybX5GYQDYhhAvNWpHq9cSxh
imlMzlZMyH6wgSuKoESLhlPdBeyIDfA2DFZBueVLFnl20iNxt7abdCSYFfx8Y3U3BSuNQ6vX+6iV
xm0DI3AIqGBIbyiDa+lVqshJErZ/6/+2B7uHQFj9NAJMvY/vcSohwehCcsRorzbaOc1GwV8LL80L
K5uNWDvo9F/BgTkVMQ/tfhVt+0ZrPkGq72J5QcfZCqAs3VNB18rDQLmflZ0l0GuKV9FVl3LYbnuK
TyG8Mckd5a6QLGMpMzbTxqI7A8Qs1NG4YZuE2aQyi7gQrzFRkzPzCq77nq+y+vBtaEbPRUS7R35E
W4DVgtGft4/R3UaRGyc7s040RXtekH3CnRt6UfI8lO8gEYusagkg734iJcShGVDXZbkWzgLkkJdS
k3+Lk9OQl0Sx7Qw15YfA7RynziIKnCEnQPqX7QzGATfWMIt/r1B7fZx3SnmqjVD5eiKo8r10Jd/v
6K9gkKXYRP2os5J9+JSVwRsFkSZTROeAEF/3Xi7Qf2dfx16uRfVgKuaYkMuN7Oz2E+JbboX6bfDj
a8YlVSl6QaGoHQ2J91Aye621hIOEoFip+NGV78GH1nrBKgZYSpehNBihw1lq+w8OyXoAPIL85Rz/
BYDdbblcpXD5bffs5O25jrnJPVcXv3RFGgaQyn+qy16Ib5S61DxecBy/nno4Mo6QV1ijtxpVPXJW
pFYVwh1ScZqc/DnkNEBiISnkc5d56zHE3202IQFnUbZTnV4T4cIihv2zn7YdzT1d6epQx4K395/O
X26l4XXbwY4IPBhQHYs8/Oier/hMZ3TB+tDzGu3TSWh4n0hCeg6jSJdOgCMYajnA1tSMGY0UfZpC
CoYyC9Ix7UKWlq3yP8itP8+VjHD+wBBsJisbGy35Q/1xKj4lXhIyMqQ9kB4cOdn4NJMCBUyQIwbn
RrJ/0h2tt5RPTYw1nCIgPVXTWforAphU7IL2WnJ1pwzZZHhOJmbIWGCn0Z14tjRz831zKWhj9PJG
AN7spEzsGSLmd1Glsj0a1Udo3eIhMQ2udtRBfu6eLMFmoVIWmqDXZT70s2iPDuQk62y0wCyIg9ma
o+WRW4Nk9HWKQlo17PMmszxNob3VPSZETpKsHxH6FW/d8fxL1ePK+e8SQPI3/7hPCyjfx7QD2AKl
RrhA5yu6pSukNQGei9xCL27AP3LGNyzu+doGr3HBfGOfMaggmfbhEUPN1fgrvRoIVyAYHWh7BtEw
F7nh3nhVe8uSfbvo1/66wFtk2TovmXFK2SIJvZSh56sljPsbvCT/5QQ56Wh3jSXWYcbODW9vx/AB
gYvyCkKK11Jo5+TQXWpuDBF1T50XAXiJBYBxw44kHRM6Q6hBnDVhWDMOKF4pn8SZgXjv0I0RZQpU
5Kaq9S77/3Iho+TNMZEfg3EQp2rEaBKmt6pBn5hn5ZixUHW9Ztwbc515GLvClOmcJ4YDcnb74e4b
A/KJVt4nKNmoP62qx8Qm2liFKs0C4VZKMjfGB8ksMlIeVRsdUZwrP5XQYT4IBz8fTuqrCyNhIe7Z
EhwznzGhHZ+4KVLxPkW99CgV2p4/MeldBOHt7VYj1ZRk8hGm7b/swl09Xf7+UJssKjJvcFuoGXFe
IjptLVm/2wjC5I35h6z0IxyGfgyqR6ZThPuAAZWMaPqrW0BsJ6IzPfszuaJ6U5EenOXKJEU4S7cL
Ux5zzRzZWxh2ORSPGR5OrFTC1xutEdCshKMuziI/8Wih/YZ+vD2zje72LIng/A9TYoUlPjCdLY/A
Zyy7+idG4DZb9Fuy4KaUpF3Q8gIOLfGx5ZgN+8h6YXA7huoHiD+/Htf0Wwx2FX65Zt9HSsOzOzvA
fnXW96AYMXAMTs3s7N3AELf8Z6NLxHHqAcNGWbEJ0tVR+ehcs/wyhP9vEK1Jp1WMoa8HA2P/Vgc3
zmkBVpJdOXTpXaktCDh/o0ccTSJ6xhmp2ImoKZgwIJUq1lQ+DQoY1NhS7RTnd4LVlZ2XyjtSMd8u
mrzVnkoIL07plzIIAb1ccdi9MBPqNcuX3KrYHiXwtNMpmTWgxPvAAzbrkeduqVnU8EjrBLZqpb41
uV8Ms/oS09VIVBo+6k3JgTvJyb58aItry55K3m+L5sS9jwHV2vBPoV0CinhyNTxNptXo7WdgfToz
mftYFYQM8WWbE/YOpVst0YbIj/f699kmKuIgiTzNtzxvAKO8yI4ejZiL00J2OXeZiCrAJA0VEBPc
BklR7tqcp0/MvKeLnYaedNyabSPncU2+vhdl3pVFd+YEa1sGNZSMowyGB8sFeNt1mzVi+sVmZ5Ar
B4++JgiTPOfdFzPKg3iPVXf7tclmUZSrwdSHTciizLRIlR9tv2rMbRPEFqSYz2CMr/YFfpsvVGi+
/v8fUwhrpiAgRiQUGuvzRUvLx2sfwPB/h0Z8JduNcrIgTp+TiU74RCK9I+HjrIehd4EWq0Avxqx0
3/zp0b0XC/baztW2OlrVqBuapyC6mjzRFj+oBGaIWfDURvo96cgIZlO6AJwLKIW+7GIKUjGxYqV9
6oNjQ1yAZ/3Zbsxj1DXaQqIHAXcKh3/i2BPwqOdUF+Q438JvaQtSwOpJCDlcVkliewB+Yne0gE8C
y1YK09NDPvqH8ME7px+1245M2BfTsbord52aZKo4VPDsOARNC9pb4NKJNAmvEKcz5pgDUg1pMzOt
EIn8EM7TcD+0DSRLBy7c0QsX3BkvzQCa01btXw0H4Eh8ZUUsVo9ZKRc9cJBa2TkM2coNfJLiVf2w
xaUw1jtN49fuyPw30aIIlMxzFUMiCGvQ4IgOtJ/Tzy4Ly4ujxIntOr0zI8jM2+JdIBVklZMuEm8z
MWP3EaF4k9ryhzXIpvY1qs4VwK+j8c+WJ9+fqp06KazJHE0j0uGzbL612q2Brz8bcalzTJmc2XDX
54eInHtIIUa8i5m3DjziuVkOjQgJU/4SnpueBIz1aiH0bmS2HL7v/Eg77q3CcUZrTst37ghxSjPv
RE2YFd4tiFa3bL0P5taoOKJG/1YDBHojk80W4DZju6mAry+0o4tNsAg9cFOrtUjteSU++TSx5YVK
mgly7rvfJVv2ylkmK4EV1sMW9Sc5prAvfyT+rIXpG0xREGIAILosrZk3CTKEqp+pGBEoHRAU+PTm
qawN7dKPIoeFDw4Af95qdksuPCqhnyOVfvT1gxKVAi53BFdh89cUbD7Mf2t0CTmPmPVlanK4ZkFF
TSxRbaA+6KAZcwJNdZJYn2J/iB/PPn9vI+HX8Dh2Z2Wi+1oZzpFjG8Nxqwf2qbenxKE56POQBH38
ItqC16yP85E4rych/iBLiTQ6HY+p7EeQitraqiQgo+XiCoW2djkM61vUqvz3cEHlL15sY2b1KyUI
w70UT8llrQFjitl8qUEZ/tE7Kbd3mbFX78q0e4TZqq5OkIAp/QOQkCKuPh15nYXtwwATkFs1hePS
zySS3/Ya+s5OwSiNKFndmp0+87syZo8E55QqZjM4dJXoDr52hW1FGe5FwLDxYEG6leBHlMsmXkbQ
q9hU88++QElpbHcq1wkubzNQtBpNpPa/QweQ5VA/2vKyEL/Qr376BzW5wzsm2lkwJVcvFbG866ko
YLZ28K67MC9+kE7Ef4GuskYf+yeBb7WADg7039uUqDEGLg/AAsM3ZLcngBt4pLJNnVc4CYc7Lbdc
NcQqiEAf6OYGF9ALCYLaZHnHB9UkMYEWDIyww/bIZ5z3hHScKFjrv9PALA4jBQutV9NDhN0TRWpc
ICfmjtbeNl69b2BltUloBi2apLZ0n1ppHuFEGUrWq9QCk1rBJB9aNuIhCb4Zsc8i12dE9OEHIj/l
VnNenT/QeM9vhvn6ujKDx0qCjW+c2FWf5SvLq4x2tTylVbBBWio76a5PspY9+huZX69u9ya+Zr7G
NjSnAQm54w9c2BkkM5d1RwE9BS5PgoTi1RoIEoMYUdDuzqGJXOuwmaOOVTFRySJiWQIWnhpc1Fmk
TDaYUfUbxcN/ur7brYWb38l2ALhXopI//pGjgPX/7r00cnbtLj9fOJBvn9hlwG9d456V/vHYGD/G
xfviJLV6Zw8T7F0IaMMeYym4S/n2Aq15IgrhHVZSnu4o0f7aEacxxpjv0Guftj5Hjvb7QKp/gcGj
4sSmmgzvSTP08CL1XiZx03D7jjGGFhJOP+FOFchnsw64wRtj7/zbufc82s5cY2cLfmM4V+GvFQC5
zwdiLiU3V/+HxpjmLpp10VAwC/wQ/Z7qr4uj1ZbEPNnVcbZjwstLMeT2spyvj6ZvM581ahDFrY93
rXOM4RfdFrSHn0cFBPBDorPT9yVgFlxz6YUy6IuK9++jyTR3p7ItY+/UnT+pfPoH8JmDp8riTu7a
iQB8dK9Sq+8o5eh9gN5nrSH0Z7Qac1Mfo/GkcFw+dhbedVy6wgldaWBEooI04SLkoskaDw9F+OVe
6Or/mHHUgz1jr+CB0lTw7rejQ3sMQe7uD2LJZbu1bfl0GHx1Nq0WXE5jfkWDNn3ARb0MsUFz9kuT
BDL961TD2vRQkrdXPRxi10RrIqhRS+FlW0CXhdGCS6VrfLlTuD4ixr0n2Geb+WtqJ2B8XgIjxM6v
zhsnAsrmM3XuMXMDhXL6/ja9CZiGOlj6JVF79drv/8KujvZ0icVpziFLdnzCn5UXiB9Mk+MS5Hc+
XjSjWkAmKjfk4PyQTQpyGvq0/1IPLl+B/p+BiYLuCUF1zeBbotJcWstckXChKFMpyvWjejtPohWI
JA97RAD1iA3eIJS235JWbQpOJKh6GSn2C6YKA1xE3Myh+P4eE0hvaMIhpPGu3yMWO9vwIWHMcfYn
CDrytwOIOkUvuOXdoK/nmGmR1kt1r6vpn/rHGT2zTaTBwPr4u4mmviBxS9vfxVegqrgqVcQPabvB
KiY+VpqznTH9RDQq/doTbwNg9TgQD2THO/3+cXU2j8UrmLFyAyJ86AWIbLTG/SGpBes/CoSoUJQf
w2GvJA99Be1KhHAsB59z4jkMwMUDGBXywpHbs7FIDQo/BLq5f6jks3TF1rYdtlkOxi5c+HVE/AH2
mCjyj9WB5Xl5gONNspapwszpzIQewL9eMlGhTvXT3ob0MFqeUPPDsbnl7H0clrMtvk3ECf+A6R2A
b+F5+UTCQrJ13k5Zw0cIcIRcVR5bTZMenrH195IQpFGqzH+OdjTxwcVxjFXAnSm0LmZXr/4Mb4E0
pwbU9LHfHOe17SAtLtO2xktEqLIKpm6b9gsb0hW5GbHZCp0AF8IRpzLP3K5iElMuPMGx1kd2RfGU
0qthgMUrzjGJOnCoiH9+VDTZqhL+G7illjGuRQ34bmdA7n3mx6KyeuAZ7vz+vH1QjT58BMmmi4DP
WC20DWG+FlB+WGn3bHhtl2FLwoqsBNfclZGnQYVOdEsqxWaryldOfGckYvztJ9zDpGe/od5rYZZb
w1hJOob8PMHa7+16cIgKbNEEBcYYYeOm4wMCMNuj/lmjDARcgF1kls7p0xF/cjiiFcmiCjMQPq+a
C40n4ZLO14xpktJ8fRFmkgTFrJU8/jEW5y0j9Vi4FwEVRoY72tUGXufDGINH90n5EMOsaXVGi/P1
auQWqow5GaLvn6yXXORHYBCIzpOZ8c2FaE6eBVq4w5qQBDMQb3N/jR4gK4HJ134sWsGmWR0/8q7K
RGIaroi9VJqE97aoLTRwyqPCrEKhzEWIcuVy66rg1vI06aJ2tltJ5j/snCfcxpN/7RgCU3+A6Q/i
dFsM0jFbtSLIlnF8Ceg0zY+lEbblQa7FWLjLEm6tp4cRpHolHcj19g6VHwHBCo0tUBnqyum+HI7F
3KskHy6PXp+iV/gDpccWFcqlgn1WVbcXQbzUWLTvkeW0Gp67weol7gVic0gVF3boyESryTsXK8uG
sLi/gkIKj+RaI6oEuXaNYH3ExOiU2KPS/jDfvKVglIpXUB1rd/s7c9KVbMu5fLMTfzha/d1b2bZU
u20jnnz1IpDOLdJ1XYENGVdT9/NWNKWLDrzw1AhB7Rax/rgiarJf6FmGyH6Qr9Hn68F/yfEUcgOl
yPHT4CvYIg3nM9pUgrRZ5+rUjyQYZsw5CTCYdHuONwG2Y0Zog3/gdIzr4tFBwTNRhBTrRh6Ce8BU
BQyWOx/78wAOmrxsz2XwJOLy10ZLiFwMWx1XSNP7VrgVd9RlrYS4IjpuuZ45iNKBMuP0bUJ8jTwo
ip5zzAIbtL/B0eLHiM4XoJiq/wSxJvOmpJOmEEvXKumziU0gbHmk3DDUwvIZMqiblXOwt2WBgr+l
V2x3143idbfH7uaXukitG3uxifFpzwywGhpS5nnjlAxyoSpMdZWXTQh4xT0J2EPDKFubk3ij5dSB
n+owMtFsBrLRJjPoOkzHlKMbXSu1PPtjLLfz5B10qLlCf80s7M5wL2u/fEe3TMmv4wuVLziEs+og
dK2ioI7E8FQs7PBgDRmM31o4yqngQx3Zq2vLDTQ08asy3/5FQiWf5n2TF4Ovop/5fGgptkDzOpTo
moDy2EpaiT6d92mIUosjgaS4TqdsySw3kQsga0NdJLsr29jDRMorwggn3xdYYASBvzeRdeSeE7i9
hIaMEaNWiUxG++slPbLuU1iJq6mAGwAHNejOoC52v3UPDOTXRy4HOG8FJhl12BCC56O4SMZUb3OQ
q9yp4u1sxm8PRr6zPKQHPUTPkuUtQ+2E2u759UrJGxpEVGHUAufSVyrG1EIgtIowshtNf1VNpB3N
ifS1JPgTLa4uHVI7He8++plhXHEJRpA2STvzbXcTzPSNBw/59OVzDAylRJsLpTBLmr6RCAS+eKdJ
n9awZHFCIFN+bdqLg8uy0ZQdRqp42gt4PQNVtunf2npRmucfvQpH45bpLO9Ip80c+yxxJyrXDtK1
PkeD5JprPDglDC8SBTJDbmgkYWGJNqAopDjeMlxVxf6JqKW6mTaFgn/j0d64ZZQi+kIAE1W4sVL9
ipzKSzehYMbdObnyxAf97ZRJ3oRTZXibbQInBV5EDQWluVTb1wjxIjNuBXXCII0YxMxX/90EZiDl
YLxokG9LkvvdjHa67IAZmegLKOcDpTFz4hrd0MjtpIEiUpr4QSlxntLibh73Zvr0AB4UcuE0NjHk
vWcA7FiDDf2eSXCGxK/R5dOTvJyKg646JGmLn6QwE3YAKCnnZt5N4cGsVY5qVnHArFYZcNRkov09
E9K0lJ99rVOjNzDEoMFKhEpBt95BpXHzYQoINrMmje7ktRhs1Yfxx5y40VKeWrgxNciisccXQ3Pa
8lH7YeNaVFsvs0qtDigssK6YHO/qRIJDuyX7HoC2KhJvuFcnJAbWq7IsqwkEXB8Nz/pBjZwDOAQN
QPokQN1CBmMXM72ZUMrVmkvXC3DDg6uAjRMRtRsYA01hVNcN/LQqXcMvytVDI54TN2/pLG+Uy50U
VClQLZP3P2z830/bLXhidK+FeexLjJI/sqSS5RLZXyYE4sBHQjeGmZeuMCBbo9UgyltvKCNbcJ0g
RCpFH100v0nqVVOHR4a8AtdnW6kxBPvn4Q70yfdC3Ig8dNIDlWlknhpMQJHUOVLun6c5meI9EMzY
NdJURmttVj8hIcTrtoG3f4hH5ITYY40XGBEQJ2etRCtZG1cs6zHvba60cU6NhC4ieNnnh1xPjPyR
CtWdtxRFhkNmwldg27TRTgVCPxZ6slhMuLI+VMYbcURQ4ZDTY+pE4wvMlWFBuWOwzL4kylXPoONZ
lUzei6qb5ukAWY1Jl0qXnW7YNPznDMaYej+p8sfAXAClLg/ID9QCcBNyv1f4ps2LnN1JNK/ztkdY
1rsIJCPotVn+k6vBb9bAT80tQaxTawrQxul3tBaVRHf3NupbIgETBDv49v7pcE6kd+q3pIOiLVtv
SQ2WWS1YLNC2mm5DZ/ZmJ6PPFTtDAbHWVh1VILWWa/nG1UWNcTGpRVphLM+Bvo+Y4dEF4paw8nPs
KKvahJOMeju54dk2ww0kXiVSR6E30CUMLWw+EcGhEUtO2pjjFZ+Nm5jUrdFM76Rqg/YShpZd5BFs
6OQb3O8Wi1Xf60v0yTc8Q0Pa2pHuvYYTWxND51LZ7NPiPAPOYjVM71dU+sgSxYTK7eVA1i6u711/
H8ao3Wvp5TLkIF9xxP2/EtFgw+McglvIIqliySCO72tqQkPUFhvRMXP7vRPgOXbkXkO5R18+SWfc
Py3kGgSY+pyTbLI9ODwUbDbbqFSjFobNrsUEg54Qkdd1vVsvXip1IUB918gkJYm4ucaN/ZD5gKVF
obfICqwg+RrOV6grvFjo+/j33BNWrGbUdDB57TaPz6lZQOVP2yNvDlJHBk4tzQtAER9MRikCCI6A
rea/VxCwMnWbjekWpH9BT4fMTb+dbngbNvCpZKC5MGNyquBGfuqoCP3j+VFLx8NAtdXkOHCP8hYB
qeMWg6IrXwoLQbsPFnHQhVJndfsuXVTPbD1eCH8CmFx5Jc5Pw/hHwawckgA6MOYbb4a+M5MQwFNU
68GJKHFE7PmmTvteFWfJGWYbzyYDe/mo5V0onogAZSXiarH/1mJCd3ecaGWEOy1uIvqwv45OMRrc
MqEE9lu+JXfGEasuo0DhZOllbkxVpkR8EJgvgaOZ6phL7maXKvisza+0avSUU+l2eRZxM2A1ayM+
P11ph4AEWKPcdJ/2L+d9+A/QqJ8fhaHHnkHL644rrGZaRqNuGGKNf6PVqlheDbYLzjJuLUi47epz
3i/gKf4+uZpI+WnzV7U/d8SgLpKGR2ISisZTG7GlU6qPPorElFOaa5bXCef7C+9n39kAbgrg6nrm
A5GR8EjOHyFW1DoBFBJcMeOTwLLYsTba3n+Z0SKyXMkcsz937UfiHCroGRP4LQhf3W3dkaHt5vx7
bk1vdbd78DSZEPgow0hEaQ326CFyfe59af1pCKMeZHVDX/n6Oqi+yrzi1gNdN/+ZsbUZT0O4rlhU
8Maq2+QvSiSBthilxO3bPcWpQVRyulzaajTy2iLimrMirqgAOXV3iG2DzP2Ou3xglvGpQAPjQ4bs
Dpwhhi1EO9zalidFEZzdO4wffsLxTapzf+P7EqvPZL9PrRZyibF68wTNcu5M2kTXuHAJPM82VgLD
vxZnGlNeFlSgZDUn31Z/a3dMJ0lAVMvTvKj9LdfUM08mGBmwt7ItL0COBTu+jHy4K2rWQDOSSpN0
gQUOZtO1zHxn+Mv9eeOdcTkddqiZDAXfBRquBlajeWOeuyV1WlHNfqGyBuatPrFI3vR4qU8J89hk
sT9mDHU0Vw6Xzn7KrljsHojjCg6IJbTKyIY2JnMpWKbRPb934fQm0X7hsIj6HNkbmBgOt1M3SEiW
Qz8FZI35xYZ03wEvHH+TqYsYpPmFL8EDHxI/ojb4mdSNF/n7ZQLNOflAhsAO9D3W6oaZUzHGZBXi
zDNrP6exb5cOUaJ23i85ESG6KGU4WVv2Bq6GuJ/gRU8hZH4qCxaG7gdZcPmDDQpUYwQ/qc7Vi3L2
jQxkRuh1JV0QHaP5ABvngwV5RH/FTwSegtCDGUogGPyWtat9nIdySP9Keqr5gFQeh0NOTwOxhadE
Mx6Wwcw95Mdh5GJ957ObiVyOfHVD0Y0tKx/yRNRJYqSxz7ipy/yKjc31HxgNnz9KU1SkH4LVtUnk
+TZJHgoh71tpdnZSd+z/+CbUPUAK0rE3tgP7+NlX3FDujJSCYVVoxieh0IveUckSBrowukarXbC8
4NgrcLSYzHH78AXWGNCCSZ1zKkcLskD88oixNdQqDOHsDFs8JnGceur5x07oSbRJDIA9CibsXMOC
j3WoIARF4j+YfweDrz9rCRSNfbgFcDBIsx/IK0YrP+x/mq/j4nKkwg6/grcGZIxG9Lh0p9QfbQUP
zL0yDjkbNKIDKcqCtO2aUoY9IosTjK3LEhXOtVEx66a+9BDFj6ValzAoo1WvwrxyTjLgO+xuDgim
SQKiScX6CHxputiySVVR5u/bGjLKEG4e/Ddcowv+WtwN/yxaVfB+0I0WLFwkPm8m6OvB5Brzz9ob
YFkcV2GDmXlJpN4ip57+f17WiHxFqkF99+KQULWwDDgN6hSTA5hrGe4ciHG5LJ6nycRUBfkqQ6+U
hvydnASeqAn72s8+KHD/mHwgcF2hJuHI0pGgiDkIk+T9olyV1pTKTEE5seKJobYRw6HIhCt+IhKF
OB7IlJhef9rbI4Fme0ZAGVFyu95CgjyjQDXGsHdxP/7IVta2wHcIFowQTtr+dafVUkMif/rMZcHH
wLURXBWRwy2gX7NBW7/q+KlFGBTYVekSNhhLmZO22v41aIyfxDJtLjmlqx48wXHvs+eEcjFvkugm
yIHX2C7L+NHc/lV8nsowK5i5O7PCsaAv9D4PSqh/e9fWH5lKJUplMPmlk21QFPeqoxxibyDiYU7a
Ls9/seM9zTiXmz/k6DeGhAc+URTmmaWrliPTzN7sW+KkMDre6ZEXqPLopJshiq+9k9rJNM4SXd0C
rLlhpoFwvkfOL7beSIJsxpNH1/Vh/fb7eN8ZvbcHmzEsVMRGVUVt6M+3kY0RQFHFdkf9NDgbE3GN
CwHqT80wRDH0SNaioSg3CjlU1Jja2IFMnNZ45cpdaGPxQ4g2KBcWr04GRJ8CFFGmC9Jka8kJ7M7f
h1ukiWOftr7Y9ctljia4SglT4fvWypjZREMFQLzcEUCz1yk1NsZvMuKF18U7bzg+YTiimVvVo1V7
P30epTxF3VavA33MQgtVdsOEPPzyzWu4Xy4x5Ym6JBSXRjA7D/8TaxK9gIjsSZuB9b+h3Quptk+C
ZFCOdbxPRaw8idmKfP5dn6dW7gmtCKKLkyjCei5BHFlT+zO1Fq/d2/00WnTYCLwq+Ni2ovcMojJ+
l0kO3MfXA5XfUuHhTw7aTfPSBkZR3cJaRWxoLwPJMcl0Ol5dM6m8lBXbi+xWv7bD32NiC2pFV7q+
U2Z6JMJooqSmlNPzCvygjT2OazrsPwl0gDkTX6tgwIjmBhsiq5gUi4Z4Alw//apixgiAuR6anfpk
dC025Y7Y5Kz5j6z1xDLBz81CKJqaL+R7+53hXd/RwN3D+sW/gpHNM24iGDFotETDOpFd2vt4JBhp
TrFk07dr3h0J3rkHiQoSfZgbVLHyTRIIkUln1mZ5j5yIma7T7Cf1eC4vF1zwRedSlAmDkP8EYhO8
DhlBaJ+MRCGqkTDzJRz59b/+AlFZsVCQ4u9C3+EDdlAONHU02E/JH0mQhHKN5FCwPsT1zoMoSA1k
AlWbc8jM4lptSRh6NvaCkYH31BKx7N5QbIM0dQB3I32AP4tF7rvc4HzsaQToRIJSpDj2njG9tzKW
EYUeFU8C1P4fMr3w4m5GxfAazK/QMEX2X6TTuxmA67DEZiXOuoI4WQbfCab9r2aybSAJC4Lk3Mt9
SAERWJFjNXGpcJpTvGfJK3/1KtmFtcizxAHsML/pBOWGuT6j0UqX8TT/D6lnCSkMt3qWN3vYcrnF
rrzhjo4XmRnUdh76bneSJdPjoo+rjGOrYCzurPifobo7BHXPgKdaKW58XAlsIbDhz1IOjV9/d016
A1cNpj1WUb/L+6PGk21xinCNqXDiMr3H9zYAqCkiz8bj3U73N3+sH/y25jwQXJmKMSJFK0b/HJYp
zxv+JqooqctE0fWDDbqyeO4S4YaVDjO2xLMtxM3vfQO3CUb2pEKDbi7GTxWfc1Kjs7Nfrx//KZAa
yXVP5EsmyU/WEkVsMjHBqKJndhoU3cnboN6NhD+F8DFewcZVbW4cayIPz+GKtodp7bx4cJ8/FBpG
8aZOUNDPkUel7NLwd32oQjmVlzGVCLdGMCaCir6Y3kXlhr/jNBTLlTBE+Vf3dQYiiUpws9b8jX+P
wG6BqwbyJ+o6JdrfnefwSmtDBms2tdaUoZG0TCweP7u0CuQIbIdgWZTPcbDjvxpE+Sy9inwkty0b
rav3Qu7aG4Qwi7w+iy8JxbcYfdIwkaebMhT6rsp9eq4GoBMNGSfFasAHut0Hrn/xwEkgbX2OFe12
2sbPYzX/43enE43t8Qiaq1CpXHq5N1YEWthbTJIcC7qlaMqk0HxNMMyaRKFvhXv2rNYGJ4XVqUbn
G+hWx1yauQfit1V8OPA0EY7ESmjb9n0vwijod99iApZ2R/xBGbi0bITygxc78nX5+NCSQOk15aS8
LFl4YImfyH+IJnIdReLvGUTYDmUFFbJ46DqBAdBYPZ7dwwgs0Yo2zOEg/7f+KqQcJLJXUxPqL+5t
WadZ9y6N5oh/tJCXhb2KfzmGedi570v3tgAxEXois56lgRvuYUET77nhyAen3KDQ9JWiWMLHWcCP
S76uifUlzxMrtQw+BrirOGA0GDYwE/PQ9Rjf/J+7jYhuGBv3j/k13bmIJLxj3GBM33Xayr0EYY5d
7l157MPQGNV1+r+HrEkct3t3A2Lz/B5T3DGn5nlV4jTx1pc0hP/ysZi9HhP5mn5wrGhnyfbzSkL4
2XKN2eplWe86J/08RkWpYv8kVw31rwGl1KphxBoDJ98/YKHshLsQUNunDUDS1i4uwPOuBphiBLtx
sW+lvTZJptBP5PGYUFBeZi3hsxLTqGhqjc04q4UzCa2f8bs2IlwglYaTnqYhVRK7MQKbKCOa3/3Y
t6Sosw1/lUr1bcmnk5Z1UzpwbCBjQKK0N3ffxVyU0IVCdjKxYa8D5qa0trPudDTUbYPyOu4k8ZEA
JC+fTDvs6evuDtcvGkzU7DXW3olk/xPYJoyODhCRspJ7dsD3wN0RdojRZugujcRlnd451kcWwJOe
OwV5QTAP1DnITTL170Sw4Ka2LZUaBDBx5Kq8HF+sN3lYI1QpI9OXma2+0L+OU5O0SmElwA4p+Dvg
Yr0q7NWrsR1d0VUl+tg+wM7UW9K4lk3JkmeyXEvl7FEpF0yvP63to/f34bJ2dCY5fRKbd0W9sv5A
IJ1FKF7Zykb31UqLBLvJggLJgl3xoacfkRPftQnVu53iQIOa0jkAtel/aHwSKZKQ+mtBf5b3scaC
flecPgMJyKv1RpMTslH1vjmEptY0CZ2Jz0axXSOrV8HEOBzDXjRRMRFjLu0ea7Vb+Np6DDVyuQ3L
UGeiCxFf4XmTQ+RySMVK1Ii5tD0UKt3oTcbxv00CpgRQ3NCD9bT75mjLSBQwyeS0ne0721gWSqTz
y9opAtcQ3TLruzzn7KIoAZQsuRjzBesPIKJHOqhEyZXL/5luwUUla7tTFEcZNISKgB7GYkzl3xqF
XZ+E6v+30dATzNqfGw7PuVadJZ+R4ely7a7AX6xAUuUKg0/5VTJdQew/fCjrkPd/+ACDJW052XIy
xt731azXNTlikAo8jWRpT2W1M1uxemI2rn/uXoDUGsC56oorPw4/9mx7UFeuBG9IC+Fdy0awVIqd
IqV3ySmw93AM84N1p1VnFulvvpvsel8V1is/2PvmvbOmNKEg12NL8+0ysYFiubZlOyR79BR/x/Mi
L+jugrF0IF4rcYlxUsSbB/xjk/+KyeLui8sJZ8ZdLC/E6B3FD4pXrf3UXThpgu7qYMwB7v4S3OxN
7vunKeq4OwjR51I9humU/jgKlvOa3E8JYwh8hKJlobR+f4U5m1BPKPFnYhi5FuMe8Vm3v3hkKqeV
nVxeE518Cnx0tBLK74xRK9MIZUk1+OnT1O+ZNlWzhEHqnUQVYJo9bk6Bxulg6fETo9zOJo9Juwl4
YJPGEN9ymrGFIF+49HNh/nKxyeCoGZDVd4XbTe98LAovRS0sM2LQ1gYrDOqBK70d8Xn7VHB5xekW
Q1ISfU5cWefbSvs5NCkwRaN9G4ZY2pMYiNgKbCFi5WBdPkXpQEeZsAts8dyl/pV4+wy9Aq8C+VV/
CeqsamDZPY5JKqoC5ORI1TkkXaFf3X9Cop5rhtkw1MUFOYzT5iHdIYSPH93nHKn/qMMkjaoDmLUZ
c3xyQ/mVWWgonqcvBqwXD6U4gGgZhmOx34oJLohhyse5v3FOPwPtdVY/XhX4ZwqUvxBsjctuw7CT
NDUhmmLLuF1OK3yMUJsm0nn9J0JoV118N0eDOX0KH60WAmagBkUNa6avcEyf5/f7WFHvK0t0/G0o
JRkjwfWAHAkq7DKXwW5iNWOPP1w+HAQgmciCbYKICdgt4G6Pd18AThe9VitQHiv2XOFWWybhrrQU
aynaQB7vtlJDjsuXg+vQKO1cP6Cx/oOKrYmtlzcXwF8h1TqxOSKv0KRZeBd3ZDaSIulj07hP8tKL
iDAoiT3HftuPRxnYvensG8k1noX90NaSnaXNXHii9BdRYVACVYfZU+4zGJBxNW3uhXMlBU38df76
Ppo6X/jaLi9axBWphTz3/xrJX+m6+3b5nBmef+dW0IGG+tJt+fitcjxM4YC6irpXSPs87bQMwhOa
uC96/+vXOCDw2XgzcyXYtbwsmEyVpf+OMyq4m0xiPUPZD2kbCLn4C6XdWB8Uz4nwurWGtSJiL70V
zw+LbNzO91ob5INZznpNFZeIGR2A+zvEV0sNjXNbyHR1w6wrxpCL4Xj0t8itJW7dnggg28UqJtPJ
epDM3aSLZj1qq0Jmay2hBoOh+mdaRm48NkSmRvRmhRZzoNpbA5hpnymXdkCRsVDnmpqoWZk32XAe
U+2/DCnVFMJMy7zZixW+ml5YkyTuWWJ3hO6m+b58I2ox3ZEy1Nvqhp0+ejTsy/wUCQCyLMEgtjlu
bvz/sp7Dk4P6fRaSDuYKMKde4DQH0XMzycbkFib7+AoWeFr/LgsTg2r/HV1cDl+H+MN6CJcENNjw
Se437Mn3IDGoULN2LLypPXu5i0Ac5SR9OLAQ5KsyJS3fkwuyvNHYN5y26njGGMykqaSAoP+YH5kj
aPxTLo5t+Vm26CDH0TlaEMAMC9dhcueoypqLuYqIG4efXJSHLkR8p0aix//B093a081HfuxGC8Zw
mQxSOzzxGXaHy/sgy6B+F6rsA9hMY1gKF0MkiYC2/duf1jTn2Ri6O79oapt/Dqbhmi6R9mcM7YHK
sDCrW94GEhbTNK5ooSFrwKyXZeMevjc0OPf5pFQFZJ0rDjvxCy+V9psUDvvKu9A9vWFXocW/t/oF
GUsYj6lWyzH1uzXasuV6p1J1uu7ptECO75wdsxH/eSCyLg1b9iQSOGwHDckMeJFF1dLGOe4esQL9
e2UPdNnHANVFf8ApJLLjZc36ZCwDmY9janyvZtHJxddxikC1bb9lAkN8iPplS+uc4AOaBZHEqAg2
Gq2LF+dtw0uyUfxOgw+X670bJE6Xy5Jbd9j04AFCHxL1kUileLfZgmdQW5fg0UaOvrC3Q8u5CjAy
Tb3o5vR9RVBPHWcgNd1z6QSbxpyUg0/e+RyJE7Nnr7zt0TrIh9Ii+m6AZdFlUT85Da+Llq1T5kRj
fcWd038pgqzgIcKVEMkzgVQQQmY+2u0bWjl10ME1N/Xd0QAG2cjfZkJPNDIL1lmFZrM8GgZhJApB
NdPt4y/IPT2spRcZhuqEU742Yws0D+yYeTrGfyhosRN2AGsbYJTUr5wb1oHntK2xiojQzr+xhigK
NvBsLnfaUnwMF6QlKzMWkDJpg8LITsTQaj5g86pQtveyY/u1LWyRONd1I5h9IMwKQUl3YOXu3YKh
epPujypCeCIjDJeqpi1EPjXvQEyXhCqTaNxMwJjJOHQO0fkpCXOY73QxDTjfuhZGdegX47/5WUtn
p/xzdsgTSYiP4Sum+dxunSeV8MtmGuDUqHCmyX4LqMBv2u2L+ixCc4WTLAtaA5qLWyh1vjyaeHEK
tc50JMEsMq+4jOiBpdCNYPj65WdzvVAOaKiEZ5lFcynoG1NWtWNu8k0yDeMn84CN2dvMVnc2j9VF
iutIsFvQFNO5JiygCFN3oK5PL2x0c6WDw2BOOP7VdtH96vv9As9JhkE5/fFt6Uz0RsPYl51Gk9PD
SozPLf67nDYZyEgExfs1lM24eovxkB+vGwDP9YD5uVEK8SCWLHuzb5sai8JZnehwEaa++QYUP+R/
qklmu/3+7lg/drxWrHA578lqQqJ3Ykr20sqHEEH6QpoRjAZVA3s41T6g94Ljod87jQcNZuIba3q/
gSlQIBas9qhSQHd7QDOZKGDoQSurAdWQPczt1+9G/H5V3exUnRLy/JzGg10wK2hKndsUIQBs5JwN
V0i4JE+1UlT3gm/3aDbFLTYJD8bHVOhvzAR1q43t4PuVtpMAyAEnLSqqTp45UZ7s209x9DDIoimP
X0un2eb3lMuRDqzoVirHCJOkNeUX8GtE/i0VOiLNa/fxKvzRSt85uxtCp2g9tUkkBTfNMy2nZoIH
AY5BJmkKQu/VQZYRS1lQo+Xzprf0EWFqPbNeMezJALMv3Y/BCnSQh0b0lKU8ip3yXtioVCDf+Cni
veN9eJnV0hSNtaESOO6c+RhrKUjnh/BbP8M2Vlz65fLuhplrYR8MkPL9QaFC73Z0Xeled1Lf1VJU
I57hdGISqLE0Q855dLFvhHfZwhW+OX2KeWtuGfrCufK09hcBv5oaVA7Xov2uufnKvsSCwMdtCnAS
3CnhmRTe5+Ysg2lnXEQGhtDiLvfXptlVE1QtjXb9VRaQsEZypYbv8OIK7Hd0lZXwbkkOuuegg4B7
Byi2f7cXgxJ3yEB2eK/XaZcFVrqPLduJnc/u4BLHb8hd3KztYaiL9tolywff+9x6qONP6Sjd1Iva
H3z9vKzX/U0SdQB/k+3SizbC201MmKl0mR+v5JOZBx2N3olcQlzEC+T44KagIZk+8h/7UTHvAuoH
8Ot7kY8gHwXGEnX93EKziUMT2NP0T8XM7EvhjisP4mT3eq0MY46lv1Ts0kduAtYRmYqxps5K8nOk
qoe0rsUd8msWnsSTMpVRvxvrzsVi8TukpsZM+u7y9tdxExHrLkE4hXBLcyGLosbbTixn2uHq3X/q
+FAreKyVM3c7oupbd/TqSoOeW/P0/0oUuI9ZVocxZN846dYyVL5jIcTr1jbfhxl+gV4/CpB9bmCV
DjYJ2VJ1yCba+SyCJPL/Nm1/+uFNxObm3765qg7WughhLN+gCifzvXsucoEoxisZ+OrAwVjpdbv1
Rrzg2eZW8nFxkDVLNyx3gHPJYAY4X7c847XyB8KPR74N2HP5L+kpJBSMOFmnVfHYOD4kctUiZX2K
zIANaLcxR63EskP19eBbUp21cKM1DKxfMPikE8ow9yLeLcyWiXqesbuTEsVSalF+Ge8eWKc8qHUn
e6YItOkvyl1G3s8Qe1zWcWobd2uNdJTNl5KDIYWd76s3/1rOl6bEGS9xGUqsy8nBb/vCuZrNMRgk
iz3cw0QHP53wwjLxuxZrV6OU70WW3wBc07cfu9KEuXusRV5S5HUubOUghNI2oW3OoKdJTq9Apkza
CopgOyiC/JFZng3lbg4vgQcC5y2ckM0wIZq2Y42WddZn3gk04NWJdyoM6walW4cfTDES5YAP73gl
YV9smQQiLuNQk8x2GYHlbb1lFL38HEjMbai29owxJXeZlY4XsFN4TMuYcWD+WUnNLIw4sLXSk3Qc
yRf1TllG6F8oAWLluEPMdH0v2aEG41T/zGPgcRny6m0cSOwvxoMOQe9s7Q/oXLuzyuULagkxN0lf
r7YOs96xDLAYPLroqn+fpRqXGCgw2rG/SHP1uSA1HH9W6j7Pwb/FemKvjGcRjR/Kv1L8/olf8Yd/
Z/8GniINrmJ9WgTAFHDhj2254F8byYWz7ITYlFjc6wbTYNtZV0khLcYICE88TsNvUDOJ4hTKhsSO
FEeOA4kzecBPFg8Jq0TMvN7EUksUb/s2L+fpN1oaTtKs3d7T/s3TywbjxbmhkI328mMRNQLH5tb5
txklHj4X2q9qondbPixJy686e9GovzIcj+IbKOQby96eRlaKONdgTtAUzcvWDZQKjRkgGkgmaezP
u9XA3N/Is5/tHqTZKQ77rpxIf2CUK2Muqc0diGpN2PucZT9/Ewh7GSjx6FIWUPpv2rO0Rq733eVl
fIgE6dMFJK89KXi5Lq4dw2qd0dcVRaDdd+bxvZB3vPULBqWu/eWBZZRMvGgHlVPoPCs9j+TL7blS
7HJszqv8XIMVisO1B9sRoT3aKD9Re7e4OhzfhmlDXp9UV2v4knCtY9eJyHUwg6d/G3YDNxZqgb8+
cRfDhy9PBNPH9DkhMDohP+KERB53ecwouqDHoZ2mRcqXcTXWdhg+9PntiGSWMAdmBQ33jeDlrx+M
oU5JTs4T+QkWRfsz04tmURh1xu09hk3fZJiCNqPwmP+4G/BJz99pNBVpHS/bn96+L3lz1m0VIxbn
kPUVWlmY7Hohs7WdnkBXd44rKZyYrfxOTYLqenIwhM5Biz+sWsK+ddz305IqHUvVZv5MspBdXZr4
YnUscHyfb3ecc5Sm9bnWdrYXGIIFlLIxjfGwxhzoniSzxJZkk1R7Scn4ayOhECUuEK0NkUXR+HpH
pFu4sleHwuBTE2BUl242wYQ5DRArCzpBXI1Vv8QEidcP02TrnuY938BREG2KjN87vXvvLc7vilxA
VMIQRpFDhWXEqI54hG7sCsqyQx9ZoXyH+Q9LJi6N99d0T3cCjt/Z9pwk0zmJ4w3t++SaeA9i2tO8
2PJTMiimNeSfy/tZ27PLxw/kHVSli5kocDS5PiZeXNMsbbgtbcO+kMkjQ5hCB8Nf5bbWsHbIdyvJ
pZJ6PhFHwfku0qv8gTvCjtYQ1DImHP10ikklV0hLeIDGj6avdSP9aWkjehKkMusfhvhAwVTk4X7L
pDGBJ4n/fZngimfbm+NzQP7FcOjOWPqYZuLJwETc5ZC6zZ2cYw0QVnYTrbvJsaQAEF/CvExFhA4v
2TE2gZOSlyoq5OgmUHyvzil63mMEaxL1FbHWpTcfaUxyjmVQAgoUuuh1Np/X13d3r1/X8DCfPJSy
hSHCbFzX4CxhyFB7bMKMa6R3gilZWTPX+nLsJ9i24kUBlqJuAk/ipaQTmaqxdQ7yiX0l8pNbGFw9
5zziF/qBElOlzazNM6ZhV75F7KxoMvfFaiEJjIa9RniiAMijjnx/T5dvJcJ9aVoIrgReud8vSXM/
HYiU8eBWhUN8by22kh7QjaJ+CWzUdGEillH6bvH4szHR4ai6m+aIcu62aOWynV8vIDcQpAdK8/+u
xUv1T7kwlS33e/GuBIwyxd2+vLuf6yU+qFjfmtCgTs3eRt+2JHjmsjbIRWP6hHb6smusQRW1nrpo
VwEVpX7ExUXIJ7tJXIRFs3cKF0AtaFxHBZDlcG8UAmZ5nP+6o+Tqq9ZT5MqAbCv4VLLQKC+TI9j9
bSrcFo8RkuwgTRE+L+UJVmc3kn3AJ4HEEm1wdWtINf5y+8evzmTdRMbK3CK8qQERWEwQekfnWush
MtpCwjhuuNAucGT7KcIgceFw3MiCaIyDdHgdwbjoXD4wDyn1i8P/Jt3PttKQgzGR9NyqLc4qnosA
go1/gUJ2KoFLRySzWgOZ4h6bwdccpIR50PHZ/4qWZDEI+bfz5RQtb/Q6g4jRpCZC7RpjQ51tNXv1
tKJbfIlosC6nJ6aF0i4YH2qhIFfy59XAE5FBZTtx7gnfNw5FhwkAR+wEGQZsP1LNYz4GzDVh5tFs
lgWtFyN17Di7TLAgPApYpoxVkqCBGacRDCmVfcw1XhfP4g4X0DLeq2f7lMTlEtp10vuVAz/zwPu+
QMM8wfCFRMiepCJyVvJ0kmwCSk1Egi8PxMSDuON4KQWzYnt4e9bzSfWaLQ60tRGIuVG/oNJHe5Mc
MhfbAfuXpGvtqVAlmDORZIyXbsaGp9Yv+WUTs8l15oWfV+/IQc+FKyRC+OF643aBBPahMX+KEdVL
TSeNUN0FR4fo5hAMLVLRP3keeU5FZfddvhW9xyq8ENz65WFeDZOJd5ZxVU2JsOutEoI+koFKxE+Z
hU5/35rYq7C1JNjt2MqIOga2ZR8B3q1yLfrdCEXre19mEm6tvbfA8lHXBe9fVHfdC8v+mUUzQ3fV
sRCz5lQ2duegUfg/WWwyA2Hig0L4uBMotbJus5fJhb5LfQpc5OZI5oBZ/+KUBezjCvbVzQVtYVHE
+ehM8kMb6j6Mry1KXWbyNkGFoqpT1I8JO3OJqB/3gmqijDRP5tPIvqpXtFPZtCebcZ/ZzeMJn1rS
6IUjF4EdAu580l5IePU2LKIDS07aa3wiZqIbZyKL+S4ByyjQdNdbql8lYMCvHkcdh9osU96sucSu
B5Qdmk14PiTLBjrWAgtXNhXJk0EAQl0BfFA5vSMgQ/MaaEcfuzFJLVkag4uaAxjG7bVHh8vQJuld
E/+SzRS+jfAf+O62FlFGJgA4DZrMOaWrGXtVwn8zZUqeunnaEYArK7z62w845XgQU0s61CgRY9cL
E/uw+U7ThN/qkN89tgzdmjTDf4z5/wLI84OCiGlHwU8HJ+OprPlUSxxY8Lq5U118Z5+ryScczDQo
Lr2TtJkvA3XnJSfSdD0S3NwYRnFMQYoNBJcGxq2nL39DCSPnw/APqRpfX1If5QMSzHo8qg6Fn4K8
e8dd7Ys8PgUXfXxz0n10/Emx70MfcWxY00XEtVetSpzicHg2Zo8asRTI7vW+C0QXIfAJLxVdL198
hkZN2kCNTUo9TCWZYHCRCkEuqJhfmnhZNQ9GvXNehMHqHpPO/R83CIODmHQTOzvLP7u/KjcqYvPm
flMPF+mtdz7/szR6zJfxV+jmL9C+8p1gbjxX/khYhVsXHiZBPqvEa0dzy4BHA7sRqkIqVciAT61a
sFx7SiIOMpXI3Ju4Q2wWLbC/qIhKTXVki+jto6vE8i7oTN6eayzeq5hXa+GuaPTMTcaWPxKtoM4a
gZXf9xQuXy43Drc8dyEH6IBnFdbIemKdt1hFZrxJWx6QzPHP1SQCIxNPDuHx2BXvq0tDF/T1KQMs
W7Gw0o00efEiFu+hJWDPfb45y9KC/f+x6twgyTD8JoB+1+r3TadjYksJkCqAev6obdalOHV9kEdN
Moh99wROC76rLG3Ajzb7xzZihceggBjkZl9Ziw+nDx2qH3f3fDWAidzdfVi9rZpA3Y3UupFsaYme
ixCBekgq0KCdzzSB31PfacbQGdgvrV29O/MCWQuX0pNrnZrhchj5Wu79h/BwWfgMHnr60aYT9zI1
P28/eQnr6TSRYrEWSzz2nomrT/HPV77R7RKsN1a580qGsHPuIN3FV0RA7zsvX2wmId+WYxqFeA7w
3t9Gl4VbPZGxHjpdyJAFdTM=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity fpSub is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  data_a :  in std_logic_vector(31 downto 0);
  data_b :  in std_logic_vector(31 downto 0);
  result :  out std_logic_vector(31 downto 0));
end fpSub;
architecture beh of fpSub is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \(FP_Add_Sub)/(fpSub)\
port(
  clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  rstn: in std_logic;
  data_a : in std_logic_vector(31 downto 0);
  data_b : in std_logic_vector(31 downto 0);
  result : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
FP_Add_Sub_inst: \(FP_Add_Sub)/(fpSub)\
port map(
  clk => clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  rstn => rstn,
  data_a(31 downto 0) => data_a(31 downto 0),
  data_b(31 downto 0) => data_b(31 downto 0),
  result(31 downto 0) => result(31 downto 0));
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Tue Feb 13 23:02:14 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/Integer_Division/data/integer_division_wrap.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/Integer_Division/data/integer_division.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
mHE/yqjCvkR6He/FA/QH1mwV9JKb2VlbMBkHvcetqccfAuzVeGF5FZ7oqIApy0cpX3TDA+BierYD
U4la9hh1dOmPZ3fdDQMwi6hEuOXjjVlFqpokIvKSVNsfmmsOgizPax6nfh3WVNxg4j2gHxX91RR9
GOOgKSiQuGHINmfZ2U79y0DCCwJjAlhhf79mg9Opzc0HOwqxYUf9ox4Dvf8fYv2+uVIXkoSeSkft
bMq/pKu8RtbRN+Fq41n/6pErBBzuJQfjuT//tNXX95Dtw198cYNplcpHDMtZCU18lXVqQiUVBXW9
2XqxaM/WkjWl7S4aeZxwkiAJeoe3hZfiIqvRAw==

`protect encoding=(enctype="base64", line_length=76, bytes=491616)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
xZD+dEAIGdVGtB35j/wct45ZyiezCi4BTXg0pKHpdxlbGSc7CzzVeuXIMypx95ycxe8gjni4PEc6
mtzLP/MbxtwIJY0TWv5tu7mNuPY0mlARBP8p6H8ksY4X/2Idg8FTV+y7BrApPDnb1RjRGuiDHw2s
AZ8QWw/WDVZ7ZdRMjsRGDoCjI8nKe4T9ZiWfUlBrEkMqPnPoVF2cz5iusr7ohDy+xXIvJ4y6/Qgm
NDye5lF1z1BnQWAfKwLBUYbkHcCZ47bb4TAM2xSKbfXmq30d5z7kET4EpWd2dnNrSfhTneMlK+M8
36SoGX+jDA9tjL6wCQ6l0wk1yrSo3722mTFZF0q5lqByWxom/UBzea/oY7Ne0h7gtkdve7Uv7LW5
3UunxXPmQOuHrGtKnjni8gzDAs1Bu/kl2IRlFzNsw0IdzahiwOMfYzO+aqDZDxwtxh8jnPZVY+r4
SwC6ghEbVtVbngD3v9Np3sFrn5oykdX8Xd/Wg2XSO9+erSToaQG49JkbiBp5kMx38Q+MSrUponQF
YMAukvekY/5PZ4g3dNvL5VHjZm956GNQF8r9p8H6zyYWxXx2rzzLe/Z0ecuvvggzFodhhwnZDq3n
S8asIOC6RK5JoHBjYG9naHuLLYWb2foFRDarq81/EMfwwtJQ6j4sZfhw03W+dJznd6v5NLlBmYNX
SDSDY3AsRzdKCvdeJ+I4pfC7K5d77RaBcVPv0tOvWI+l5kBel8qUroTnznaznLYi+dA8C9eg/NGd
W650at3gAqqa0L4hqlK2IA69orCekWWk6Puh9WbnonHNqZJnSxjkmYFie9ImQyiullg7xV5+S6CS
MzvmGyNPZ4FQLFIyY+8ub7KSe/XyMsP0aoP6mTLTIU6p/UetpHm/qweg79Xsb4+sQnQ6+Red4HXs
kXupvvTgQmYXDlrum7OAsmVReQcqgobfuxpKRUVrXdSSLzQ3lhgLGISGkLtPkeLqOnKuOLPEvcXW
4R5ca25SEMcYNvFUeb4xqdbvXhUYHWOORyV51O7Du2OVz/uXA3VwyzNWNuYa36fzvSnEEOMObU61
vu/0ad+Va/tuq1hnZnyjMq0RylwOa+Fz57CgKlVDvqNLh9KkSlVb/MZI+OTHlR1l8J+FuTfuU7ao
/VOnLvLgVO+8iIuAXoloWqvaAWkeOhAPKKH2mGXH5ty5tJdwE2ZNQZHKkdsy1oJEZ2khyo7TNwZz
IgF8Ntyer/fBbtAhHUFRnTBn51ju9e9dJ30XlZ1M2xOLtATjTv1SRPUUVXmTvaLMTFK+cHu81xSC
iD13D3tvV5kqpRr37JbHWRQkN1r6q1TfnlNoGCU+Lsy3+pxRPT5o17Vm2e+mjanPqa7JGdT5zvv1
RJmCxeK9iQipkJmFtWAY84JEzhg6tzvJ8XNvYkZGPFSO2gLDqM9/tzGDGgZhkdfzj3XDg6xlAoVl
tfa8tTnXVt+L3pq0JKW5x+80AVJmP4Fs7hUAkdewZwF5MvUdaD2wdYyPxU5AoUEzsYVsc/X8Az5a
Co5zeARPsnyhqJhLDvumC9dsdDREtpC1/FQ7Cq1Xd3LVoCwBEryYOEtpgek4ScLXFL3K3K+S+mo0
2CMaslegUWC12UtbTqS5kR/8iZOLxR5E/a39ZMMnH2QyayfjmEJ9BSFfSGsG1btHdgkt+BuobYWJ
ygdndWNjQXiLUyLOj+gXAh9ljgaLtx5rZyUaCczu+34GcIvsSv34sEy63lGEL/8VVpxAytWRNWiR
8FlKPu/YjPT7/gQBxOaOVb2WFGjPI6hAxfK22sje5CnVPknKsSn2QB8pYcHM+S962chsfXFz34bn
I6dKXoUbDD5eUNWedzJ+AlkgTVSXNC/Ba0sYtcF4rqOIQ9vEhrJu8XxTB3v0YdLz6Z/KLeBzJXdE
mdZSoKJdrJ3qB5/H7V9PL6gwjTeFq6mJtSBSwRfS5lBcrVEvGRXLFv+W7eRPYf3bi7sWTgnU+MjR
AkOtzfbnBv5dyWrKczW3+RFqc3oZ2IFLcAHaPMSt+Ill3Df5dooSnzmwAvraiM6nJsH6ZZ5vNAJ4
gbNT0jWsTBxLxCG3luG1x0mRnRzfVy4c6uUt6G+SB7N9naY5jIH4fnhWjWGtnhB34V9EDoLTzaFa
+70ZvD9ZcO8BJj45JFLmzIe/ArBRokxfMZYbx/HUjVTn9zv0CqlMKgIwLVHCCGmMqzLzCDDT4lNp
tPgh3YFycpSGzED00D77zF3oV+DV5MydYCC92ZpC0zX7UWczvdVsGPtzZ1/aquCQpjJ5yh3U61aD
aIDdEt3RLMfDg0tp/4nBaUuMdqA8U5YNM7/43hNHThlQW2zG2IqTeSENgdYggJ0x5He7h4+xQNjl
rcWOyL0kXfyFkrPrnAegB/9ikydNDMf+W00rWzDZeN2/ClE2Mnruaq6mfq+6UOFSSsk86SIEEZVO
D5J10Bb+y4dkhbNRhcClYWzhbe92pedIpn2aC5oi0MrcJxOA5WLj/3/ibfG0ddpK2uR177ggnLh1
vRYnRXbmkTO6Y3GxdrQmuTa1p9chXromWRlEJQ+D5+Qwq3/SH9SKS4DQ9zPQP28JWrKsK+T5odpx
2gUsxdLHKANoD/+xhvzCOz3BnSZzKpPU1C9MRpbOS4yCOKvPLu45T8OFG9/HwM41csMzpjHkCrJx
CvCiWceftoitmDtoEZh2N7j2HPujf7Yz163UUdXLm3BKSpc6BdIKwJl4S3Ej0PFYwHKymyk3jnxH
uLzDfLGw4GwCgJoif07llS3ED+hUdjFsF3ECwfiig2MHtHwjlHe/yeLcid7wyZVUxr5EGcbC9TXs
Z6poVt1yKd555QTiP9COWe8TWw7bcx1eA3BZOoqODmWtW81/T+bOWlE+W0Lcpp2Hg121JOVYdbT8
S5nORKCnCOSj+NrbXITNJT6hDzXIlbencVDvuOEUqgXHaRn+CAl0z6vGZW7J2QxTyna1drgw4TjB
T1h4mi0Zk9vOPVI2y3VCe9yEqXBqqROWnLhBYDR54DnMI8bDhdcLLkStXjHGGWOoeukjmkSWANOR
brojYAMLMd+IbAVd6iDZeA//u8KLNBBLms0L8bmybacJGuTCVWCwJsGDZEFaL9wOSpnMP/AnfqWp
deK+brckdVs05eEP34nuiogXNtNTNjPUQxA6qD55KA9zWrfUKrbnPJLKNGxp1+YrJfYMKy4bK6eH
O9KlvnOxDwbgueTQ0eJx02EXMPrhXahmVr9B3xXzvm0a3iU9zmsK/ETGJWWBJowacyBcvMg972Vw
FGpFhRKb1jhETq08cHuoZ13RhWdh4+0GbRnkF2u+a0RkZvKIq88woDC4L8fsKxA0J0YCgEhayqTE
7oziLORaiqtxKKhF84KWtXxXC3u4c0WAwdMQAmDD9Yml9JnwoOJRMvfnlQw/1idW2XvUEiBH9/IU
USKuhtDe+oOZhL1KiWFdzc0PWzMRy1/XynDUbGk4kTd4mN882yT6wJBd+zk3uxRPYqhBkTSxN8L4
wv8YmvvAIuw0+5uKTATOqqygiPn2e4zK//0REMwCcb+f00Mc7tNxStPhmdwwh9YBlOzNr6crCZa7
HTx6hIzQBMP/4nAmwlK45jJ1Wp+HxojsCZutJQo/UhftURxruNORQSEQozwpwT6OrqFLfJPGlPST
Bw4Lt5UaEXwweMkn32y1Dl/lVLLbwSLzwnSO7km+GlwPuLkYdDurPLEySRvBslXb3eiGX6GxvSbW
Z0eNK5EOsjAifKINXKGMr/0G9fJFzvNw01Lw4FNjpGBS/4YoEwUGki78dp0SVVgQ4tBEHLAMBaDo
dyHDefmIOjBTbDEEh+04QX9ypwMmscKJbX8Wy3N0r7KEly/qQpZRgfeRwQ7f2n5KqAq7OCd+sr/p
CRnn5ml/dioCXGQOtuFK4E6RE5FrHMLglKAmFv/VQnTowey82Uq0zOgiZhthLAHCbdvGkStP0zcx
uHGnXlLSBWeni8Z5rkI2VTEw3atB/j0yxWS9A7YdFVXId+/LzFNMcNZEjqxChBfK4vTr3V11Ek/0
0nnR6HPUa2fNQvxa9hhtBgxTPXs60yqWZDjr+LCw9Mw68bXkyuHUgzMdo9bTOwKv05LB3yXF1S/V
wVVLdVhlxUh+SRoQqccLbyk7UJKcNzBzonuMCswaArZSqwih6nH279Sv1qGVKXsOjgZ+XBs3bmxv
2K5CxkCz9VDAj2yy8/a2IHiTyQ7I7d00q/m2roElO8e6sl3Wa1j1y+ySVr2AGyqvigw+f0CJxiEZ
Gh32c4o88cALV6l+eLCVPT/Wfn8z7SPeeAu1QS5Jxz6ER+FVherSawUzZ72grHgI5HH2CNb0AiJl
5lHCY+++dR81yHZdZMlNrDkruHfZk3+8iF3nUibBHosgg79Y9lEJdKQzJjeqhQxfsud7DVZqhthj
XLFsir8bseMZ21oNz81XJlmfgMwsgraUlMsHWdr75CKVQaixWYD9u+DqHClt9dMz5qt9H85aBLR2
ulifHQFmFn4/diBwLuUQBYq/vd2eUyW4bVnieo/2ms0k3cEl9VH0/fdBk6oTUjCaA1WZUzEGlg2g
F5KOzLanp445J0Szw9Fd6V2n4znW30YE+MVtO0DSf6hLs6oWqz3sKMeV+X+SHl7zsK190k552BD5
lqt+XnEVKxdxTCFelZfxYNUZmqLIfQf3IEOKf0UD2L2B9Wv9hb25oN+HwT3Xj44mM3wvOR7M/lHS
Hg+1xIRJKogqtFTWifYY46NECsO+Bc5sN8ikAgW6n67dkWDZqTH09z+LZUo//dSv2CcxVpW6YN8m
P6EQw7xIuyzN3QBf6VTYi8Uxc+Yk9r71spC8FCvpRMiMpWPUB0PCWkAdVpY0x+gMrNQXe06iz8hJ
YAFfo1jafHUko3u35L8OQQ2bitfrj23f7Tckx/Nb5uKsgxkU0IMRuYCcUnksU7GHej5+2XT9HMxx
OS7Qz5AkoMCPfM2VB+pn5+66nShiDW1dgu5ugtzEdBgpi8xckJ6r9uiBBZf5SUujQ2RNWRH9p96p
apYIktvFjyXuoIuCP3/6Rn0gcO+UG39xbdJdUI3TnedFsf3Lx90pVXRlUez86QeUKtSHRYF7my76
BCm261sDUtysiWRc1PqxmqcajB+IiG6mYxMK+HOXiMMrqMF9dZAjGQhY2UILJA39MEglKhNgkc2j
QBqRzOkjz9WCa/+nkHXxkbcdaz+LiM2B41zfcm5G489yhiqtdqmzmwApxqMZlAx3Sexkfn1/DcC8
syLOI/yA0DwWUDTjr22ACD/wH96dC/i+TpHu2qT6hb8VLQGAiU0sLT3h5C7eJSxtS/FWOYyiYB0Q
bQdUGI9sXRdolnoUBtG/T/Nx1uiQRH6GJS65VZqlP4LAo7tvvjW42X+aooiwY0aby1cKFa5cddD5
6iuf7iVWAekgjSPE7E1c4c45gdmgByP8m2OHYCxd6iksPycP5glkRQRRGzSsUA06US9NHfk+gSDA
anDJFoVcssUPrzqycfkJvpU5CW/EgG5VqUk1V0wT+Ydb9vqhIQS60sB53kayU+a8JAog/b3beRsD
b1oxItF79nt9BZtUE9zoKW467wnyJFzuj68FbXEvPP+wcF1hjUHiCb6lN2Rmt8U3NJ/e7Luq81G2
/H3cCEGb7ICWBNLunafNSQG65Gc0lKZCzrePUlUB+Tbow6w977bMN9hNkoncUmMF2oxincXt/rQ2
9W+L5XTq73VYr/ow7Crn15TY7RurlImzQZUp1o/97GRsxHBNvQR7oTpEz6l3pbiMZOWDWfBJr3ll
5OXpPgnpb+dY+jAjLH9NLjWLy5c/L4OzR7SD75Ico8sWRlYCz+BpJDDE9XSzu45VpkDpUUPLu18B
Uci7Yedw4d+iKqkcIXrX4YNEPC5pRJHC2gItmhMxnEousLh1Ok1+6ykA1/sVyywalZkQB8uF33iO
yjU1IQEwX+HgHzzNCmztPEXMzs+syCUsTz/ImK5KxRJJCymQP62R2GN0or0D5zslO5kdWa+LnLaL
Ay2EW8VH/6wmKSYPaXrtoSb6EarcqlP5ghTl+Wf5JXBVxVvsV58r/0HpHobqRk3pDBBKO1tu6pwT
Nb5wunqAEVNpH2lf5FwD9dHcFzgnzM6Wfa4ZeIooGAfsW32AsWHNEyYuwp+JP3/5EcIYOSfDXurV
VDNiQRIWHT82TYsjkFj08rbfyOKj9815ASle2uPP24VoX7eZvUWFPzuPhLIferZaSd4zfqfcXnmq
bxrJWX0hQBvXAJ8MgosCqr/XjxUHGHJemimAa34D6GWKB9Wnu2uftT8Ddf2tHIUHgNUzRq4G4kPn
ErITCZxlnt1ccloqW6fAazbFBE9yBaiN7oU3eiQSvuLHW4GVlg/3LZcID/ihHC3xa/GANsXI+5wA
HUPax5YqP4G21nq7Uo7MZDQKyrGO7Y0kEquhz9Gy/vOFOZaLvEvBesDbwdpX8frDjhIIqCnu2PmD
dyMx+TCarUGPNmAqXlqmI1n+m7JthQjokRsyy0rT5hiuoCori1JHEcRjlx4nDYIJ+9aETZEBNpo5
4Ny/n+cNm7D1+R5OKBBWOPBESY49Z54gzFpBXKQP5lyMQbMueD+sYOjgZY8cCPCnLQw4k6++fU0s
z06TxClPLS4asKknq2b5OtEzIc0iDEgrF5cBYwhAF75obI0o5X0K1YUilqXRyIeLIkCDV8QFgsLX
HVv9ZWjc3kQaV7qNOE0CaaBxH3P23oK5MjJXVpVhrxtzKndS+x8YGZ+gxuBpUsvMlxHc/cY1QplL
y6Kyp6rCLL6VZGX8iGWVCwufZMKKCnNTsoIQZBiiomvM/bPU2Y0lgVSbh6ja5U+hbAgcbgE9uu0g
+Qy6nyO77fR4ArwxYv4XpZZDVhimfFQU68AIiiBjtNpwFOwAUwqLcc++xVTJ7eDQ7w+jfwvrM/ug
HyyX8MZuXOup/6G7HWPVlmcN6zccOT6b/b9P+3nwAxnjZbDbIos3VFTh608QpBeRPrRRUFrVfGsT
skKXqO155olcrUKLFz6a97cN8A+gK8tWumJdiK8qr7zXHWt78DDRSjI4pPMk8/oH5u/hzu0LrNtW
odKsDpZuz0YzCCDb8mw7LAABuv7O/VimOrXyOvKyhIEmQkWvDHejudVn5KKgKbHxpafr8/Bx/6ia
1GxghLA35dux5KBOqxnvAQHehPdC5j6wOs243TGHpzIf7DKzWEzJtEtpnKvAPKk1MGC4ncCec2GA
FrmM2fozhoQUiWmm5wNY78nI4feC+g5f8ABEpbi+SIdAMdB4fKvp90hNpc3Z1+5ys0FFDZgb366g
FYdQ3RwnvkwJq8rBFuBBbbHzFRtrf0CMS24LD+lwLBWtrVoe2GH0EbM3r3NPyP6d8ZmmRiHjIxLp
rQQu0o7OxyKRgACAmi3H/b0LDqdan+USm1JH9aN0y1WNdDlUbPIEQaG/D0i1IioJrDwe/+CuXrmX
H++4zdEL6hXshPNse/M4mpLsU3aJ4HQn9Qd4Ji+2SDa/oalZmU8v89iobxVNHbN+dnWp1/5dHnFb
bxW2IgACBNw9NplvptsdjFnloYEIakhOFgDVnb2sMCM8LxzvgYLzBUtdXetHIboGg0W2pNYnJrgb
NrrJu0uQuWLxlOSjYh5O+AdcVtUTPgELG65JA+tDhqPTaeDeRaDXGaNLONr7n40gy85m5IWZ5EFW
UjckfWWBSB5+dWUQ6qQBpYBr8NYLjGiAZab7a3XuSvJ6Q3bHZ5nJJ3tWGHq9MtUUGhJV/ZzU25GK
D7jIrpU5o0la8+sv1WZUni9iIWjB7AcYRyyeikBwzK1PKo4XYDiPIdAGvKdR8blNG+56ieHAoJ7U
wjJ5l6SZlJvlpymjONP2Bq3YjR6i0j8Nawuf3JDibH50MAPpHszdYAM1GgWc4Iq69L5/5jEEVsH2
X4MsJSMHWuS32n++58YTYF8VjLtFX22j35HFsfTegHY+rOAB4hT4oNyV9SaRZynx7nKSvF1oJHBM
d7CggK+ujEJf+a2miUKbsegfGgccnW5SYqP/yYlG1x1FajiyGHcnLU/wl95AzAwsD/3BueUa+fes
7+5KA2u3HenmYJTA7RGo+IAysfnBgcHmdqGqAi1euQnODNs+aw/PmMS8A3UmobWphzysR2V4WfX8
b8Rb7ma8Dt4LfnijIhJWWgSG5C6O0c8WFOmMxzX4VP8mF1kraMZEOXtst3y/wtvioKcIrTUFLOSL
aCy6ljM0cFM3+VQp37PAk+o4L9GYo5tbPeLZBl2vkmrxvQNxNSrlNCYZ0DkkSlT8N+R7YKMPsiQY
Q5k79sHm4g3h+cdfz32qkmMdJI9Ea7LXJpcAmrrrdpkvhX99yq7wiGq260rr0PRc7f0Oo+ofpvtQ
dWuzruUjkksKJNkSPsIJmWCcCbKW2qJn5AYUXIirUAdIf0Xteblr9Prpj1A8KleEvmf3LcVRbr/v
mpsiI2LoE9pNQmwjcYnPqQcSfFiU+Hbeu0fpcyPaNzNDfxPT+g/rlIO/9K6Nkd5eI3sJ+rSO4OHs
sRGQ2pNWrizlWA2Up30n/C68AIQWcRn4vxEIWrqhXjlZyQJFX9hE9PWWX4VGlBGzvlLgE1l74QbG
cynL+WKqiWOpM9zKc4pdaYA3IUbQYGeNQ7K1vtUkyiZQKwR6KL1Q6J+lVk3tmMnlBDDonlzc/Y2B
9V60Q1/KJubr+1u8fpwFmmi06+1LHrB+FJUyNjETltl+JYNSLuXVLK0dtO6ZGT5J16QZH6W0llX6
SDPhaINiWHVNUZ0ZDOrLZuUWZxnToDpwUDkHRbPPBJC96jsOWlBLHbAGR3rLTXxQE/eYaMJlJhDf
8Sco/dWvLTGIJUIg7ztmTBMqAhL/S75YadcxI1c3ImRo7iSpgBl2KK1+IuonzKS/EqsoOTkD0ca9
b1UVmZHnDI410Mbs5B+Qj4PHuP88hABM3aS1lCFxhfUeOHSo69OEWMBwG3kK3xw0EObF0IQB6IPj
MOIvQR2E4o9XrIfQrbTVGQNRzoEROQHUQoiCSAqnzNmV9UjXpJQ4jIkkqdcCxH2uECBAVeZbyIVK
gHcM12cm5w0r3Kt55gX4J80xYOqArEDBtcGXgqp9NM32utzDiMbf7Ik7RNZC6wBFzDhktIGT05/X
/qXne2s4FdBSPpbDbJv6HHRCMqowQZwS93LP2tSrPSXueIRyj5scEMi7TFIuFNZksxtHl/mnFDSy
jrFZ037gxnr8gQ2gPabfCo034x7UML+UXDz2prAuz9ZbeopArYXwHPZKQF88UhBIsS1McWjgTHFR
56QDO06HdYDhn+vVEIBJUkNCnizNyOG4povpESfl5fXArtT6z487w6Q01rMcD+IbcmlPAzxU824R
0HEenUoB2g0ax53Mzig1EuJyFILVwpRZKF9s5n9AkUJKyFY8YuaOpgbGcrGgDkTrRmeODSsO26h0
VQuGKHyzeLHq4SymtNXmpTHvzPw7aoHfA1SYz6kH3esUImomeRZnDHPlwQZ9Qx0qUq1vbmV1/ggh
Rs5G3M2mn00EyM0OqBjJiElwC67cr5HkmGL4SqMOQEsUctBH0WXwIhwPJMielLFaVFyo3rbmNwaP
XvcHX8dumlRmyubsYYbCfiJ6gSJa2XQ3elJ/6QKUbPmzr7jqRyBobNWoYT8quijCoAoTmbguyrPH
6rHLqpMrkb9dJYdPeQPFZOk2yM7ftyupLnzi8EaUEZl3ZHUZajswxeMlB5L4s52JFzp0GSSnrDrS
kwau4nCtbLInEpKiHqvaly5AIsGCVhz2O5UAV8BxtDZt7yEo6wEgkZpVcjv76F2NjxXCX41wXrWw
u/O9WYb5znwUES5wl+xkOe18D+bX9NAZ4mPgy+3a1xO595c+z+IXdWtWXguc3vBhCto0mF0BVLrm
26GnGOdoGyNoGqiKoGCJNwyQZBJjL/fqOwXlAtG730oObsXnybqUQRajuoc5vVEF3Wxy4h6dGtd8
ca11vTYLSFYZ23Y10WBnFj1ij+8tUPE8jFilF/HRKRVDODPZ0SgAciACNxcK++IIWhN4USQreBep
lH5pGGb7BA+LcqUUE2w6KxNlGBmymUj69uAj//CUDekySqifFB0CoKTnfG+B6nlzJO5IuvZiJZeR
HnSSHyB++mjrv3gQsA1A/0SkOrh4sNCjc5ErOSx2QQCX2y+C6Yi11m3lAcxQxj8alsTWhgtpOcP2
Pv6/mbPr58UBDmxl9dKW7h/WxfuDoz6BfGOjjUsryV5NCJX9Wzp7QUqyH9hd8Kw1Ufnb/oio/HMs
6jxRKk2Qp/DCjB8a6TUSHSSyg2UrA2sKVytTBzx38kZpxHqiwYSqznfw51+B45JLRbgX5mYpw+sS
YMYDIdweXJvBkbJQ4mBukUblWtUbGc4zzyUuvZmjmSeambNO+MhW4g8THHHm9K4ZEYHM3c4g5co+
EhvmTkW0yNZI8gPkYmStIbgJ1gtbDnZy7C4CkHlJwtD9oVjzwaF0bzt4ALJ7sx2ACXEAADSH1tDN
IjgjCujw8LPe45H6E4EZDqiPeIFQQW98d3Nmzl24AAuEoMsx89Eiujuknb493vOBAkvzPQiMulUV
RGDVdlxsfz2bAKZqdGrcPwqK6eBaonGsn5nvUOUj5sAQ8ND1GSlYZemIUj70IgbJlhGbB7LdW5OD
R1rykZ1kQ4ZUmrt3lSxkyMmxuK7sa0y3PWtpJovV5GA1qjB9BBAOPcrISNjELcZ5cnqPShtYmQar
nNPDzyrRuGP73KvMcvwHIfauX4jivYttAGJ5Ft9v3Urhxh/GAzHcdeRtHT7+h4QxPiWEy4HCXKi+
lnLe3xqVpS/7CJUqCH7qmuhJ5i1trWXvzN9aMqmpEfS/UTL7ZIOTCCi1+ih6P4H17rNdB4pK58xm
5E1cD/YdDyWcy3/rKQTwesCjnKbAOm3lD/t6XQ1CbyrhsJSBC7UsEgzwlMqVB3BFssp/EtevcAL1
10I+SAS2yg0VYQXA+W5BifRlO6XFTSfXVkJuI30c45JngPnoC4CVWYwUQI5gM5/GUB+KSScejljB
QbkTP3R8jUvSe8Yb6B0Yka7ltiATjYFAYu5oDB4mSrdVdMzpUR5Ot3nF4rydrck0muA/fPidYFov
CeqdzftgLwQrwUnbhvWhwXcMsFwWRF9UaQLH0WFhaj6NFSFu80zVo0R6M7ccH/BngI/4zTdxGyvz
UUujFEmBpmx3fxagUdECdBekDXtMInrfh4sWod0/jOxdMFb0z6UY4Ndldc3hUBAyQ8Us/5zOeDyQ
Qba3Wz3FyhsE8CO5gpjmnrNWZulSnigyJbPhsguKDvXOec1DEPy4gGSP3pFJEhuu1Q4gdxxdjC+s
24hkV7Trc21WLU9r0dEAFBFC5UHU6N5mTkp5I1g9/jkqDXSFfvhkRrMLI6vT8k8jKU6KOCaPxlOH
2MaguPOhmlNhXX2TMFxTs/cLL6uN/d1xpQnMpJaEQeJSc55CGP0Uaw+206QWxC8Zln1Xlq0+oKF1
P8+IH60VabElVLjoOeOYpMRo6Mr4J/0rtrf0bsyvIKjQVuiSETkVlNVGs5Yy34mCSEDDoOwMRv/T
LTPV5yRGIPuui8ZuiX3X0UnEpPBB4G53hvTDjcgz8z8zZRPpQbGy8QE6e3/hT+7qLKpEkWwMDFqR
8Q7SgX5com+ywfIJIf5RkIBurhk5I9LPi/OfV0XMe0yd9W3YZQUXue5sXYyPNrB4OuxrlxrbpKnQ
6f3Fs2t/0idiG+wrbw9RpVJkMxcR75izNzBGpnGV+t8tYDMP/XtAbloJyjsRZe1IP4Rp85+OnTtT
fvuj2mbNat+/6K5YTwWt7Ak0C7g1vRN1qfk0ZDFcWqbtkh8eFzs0L/8zdWLUakTDg5f73YepHxJW
vl/oTxmlBVOhWDARpUOc/HDe+PU+EyS73Le9x/VJZ6b1xOz1zJfBGGiARAJ8n5oZ0b0+a/rbYuQQ
A0H7l6/XCPp3aaCQHP9+lyw/7o7vFL0rTECLFlSYv8rIjmCL676fSlX/DOgzynLs3SXEAwo0/R1r
rP9YvefuA5PDt+8otKoC6aEJUom5jaAYYTYWjgHmu5Ak3RtNQxZqUVIHeHKN95RYHEDC+v1mlsWY
agvUOzT17ARO95zvRnNm0M6lHYXR6kYhSaQgOEKCSQpuNj1xIvdIfKovN45wc+8cjaw9+g9BBZfR
S4pk/adEkg26NZBMbBUb3NRn5+pK47zvlMSlw/Kd0zDIXTra6sKfU+hPFcscb4sHWaRfNlTAuXJp
Ymf80MYxuy7hfJKsgLhU5DAs8VZvz2R7kLFReUD3XwfMF/hi2zDzqRzLGAKxSwFCFEvy8Gmnq14l
6dXht9Z0dI3LRDnHQiURvpqPw3k8HqQKixWyiFIDrytFuTZKgCD7ZN/FzTKfA2XvXApZHmMh3Wdf
EH27airJGX/36NSL+8kMNzyoLVlNwvJL1lPO/75v2LZbUxCRPSWwXMBEL+0OPPGKplVYwfgUSSk4
oPcWM1TmbVLb/r5fOC6fsxr4TGj5SD6G+zwnsU2k3B8NUVkaXqSzcmHR3UkVP3w4DQGUWU6tLc0f
WBh94fNSk2QVUDJb1cBzymovUlHVlQ5Lau2E0iQ0uWeYJqeeHlOF894ZU+2F5PGiuIA1Mb2XrpLw
QgTQqa7a/IAeDxA9h2a52V/gwy8IhtkmyEqI93yJ+M2QJLYkD3tI+hdmZQJCPtJNaZFBHkP/10Fe
/OZICfK1szCkDhY/fyxnMpfR0Pd0QQqxFucI5TVV/nWbfuZAYqssvZCnUdLzXm5JXn5iD5s7/sA6
xL0p43Az8tKQ+3YQh6L3ks/9W7haMvzo6UkzjPeEl+R+ZdnUeP7AZ0fbCsHiM9tnGLxUVrchjGqo
hkB5mSXUp4Le66Jkl94mM137aj/UojzBlWE97H8pZV+YhHhZxCNAMSqjliklzAxLZ13TiBRE8hWy
PWkPQZZN93hI3R6VBU7mUe4ZbqdLfvDJRzv/J59bpyrlD8Ggur1QOlWQj9CdH3kMcOduyY822mM1
EBYQtu7q2/j9yks04NsSFBuVYWiqggX1niyeWoNUoLx11C9zGJYWIDRwV3o0QivF/L/oXeGNzNOG
GtSbZZQ9aaVM1Yn98JlAQigw8U6q4aro0hcjiIoHnFO8snvB4NvDKffxIfDGBUNgBF/E1oUIekeO
lYztqhTEIfTq8R9wEoOVWo7ONOUNZGEG+DMsOxkXcRjwMu6hTs/U5HP0HHdnPAQ02AiGT5yGjKTT
3l3cdUMFMZfrmboFsAZsEMOmujIgezkdf+V5Bk7XeRMOYEuD457/GYNE38lDEcHo56a8/y+yx+35
8CDJcym85OnBD3lchQFiLw0UHduoaj69kvnwuL4EKpx+HI2cJwAQv5PXCYfJ/ntWn/1vvBfcjV5i
KeP/GtqFn78m2R7nS81HZn1JxsG9c/HlZJINKfuhFOEmOTMufXkjJw2Afz/qg5lX7gkb8LRMLllN
aYQePiAW9l751Fkn0krdCpOuD+AvHAq0ktT18rSeb4ip+mQZGDbKwsEf6T+QaardMIPY3HtSUBEz
mVXR6D1Qv80oeUrPe94h9dyfOtfxY4XW5SKPTfobegL73tdNvJXbHKpMMteIXQCCoTYeZOeC6S31
qxX6e10MccjHBybpXsYtrTXoH6EytcrTOlJNFjOmkJNwOp7nLD3fHFRizU/YbtNg/jIMgUizWdeI
OtF8meb5nPrE6x3mMrz/qOAYvasT+G+SfF9vSolaYQSRXPaS7ejGWfH5tUr4PjiJieZV/eytv96p
iZ7QzE34Pw6ah1FRKOMPy6LtHVBcjowx6LqYN1MptgkRD8Mbdu4PxIt3qIrDygl8gqjmrPvvfJQv
sE3FYRRHfgaJNinussK97u2VJW4QfGXQsWnZT9NsQ2Lh9rxk5BToKSRBseKn41W0uVMugpT97CZ3
WJE7+xd1NJviSwRruQJvakYoSVkyjCxJkFS35evmE409wxWSmCRuAU/W/oN8UW3MPVDeZWOQna/1
mtS1QNApigfWEWtL04/IkblnE/ep7HiONeRMG2NJLoPgpPjjGD+Pd3ovbWLYGf/GSFWlMk4PbsFD
E3rQT8s9HcNTnTobTWZ/wXzvrb2CLxFqB2Su4BMDBqPVODUXro+SVObKiB4kAwn2nO0X6aH+fGGJ
oaLDPtxSdtYdQDgH8CaPLolpjLwuxqKLeTULRKD0T648D+tHbWe2VuPhDm2nUc7h7qVV+6s22IOo
lyVPUIWPJNSH2mNpmEoOm48OFYUJ1/PRYDO+YPXZVveR7AEc0kV2LkmRZEmO9q5z127fpu3e2R+Q
XTjf+yAcZk7Q7fixSGnK8sEIVJBkSI7TcynbYoP36sEd3c1SoN9mtnJKkzVMdNbQ7i6s6wCvNkVu
di2ktEpFw6vV5A4gD5v1rE7B4xDFF8PHWhAP/FQL2gtH7Vp1bZgtP5/iv4yh1Gt0B8tuI/Gj2OI3
gzrZ3/mUe758GPcMxia83rRJp09HG5gNMwUfOBqbGGse3FszQpfkHHEsoSZu8xxOjY4PYHMVNnI2
L6fL1XbrcvtbO6xEfCDvglFlnpOQDZ4GYKatH/R6ZCHySmW7x7NXT/oqCNQVGtuj0OwJBEG2dH5d
+Z22WNh0OQo8kl4P2h36aCQfKDzV3Th5hdOtXYbxI38AAF6C9u6rMBhIXe1zP2CapBFVDmb/W5Zo
O1nHd/tmZwKXi5YA/4SvD4cZhJ2cAeOXzXZlzBx/IjCRBFH/TkIFoeLO7dgDZ5HjEJDjjKxwP8C4
D/1xn/va6U34naRrtPNyu8m/77lxTley2sfe1u4r8Qw0Kn2YPsOTAHn8X4i3kcHk3YAaQBUXaFj7
AllJPVpI7+h4KyOlPomUcZ5GGZNJo5DB/4Mz2JkK1RJEO8GbgcOV4QtwPh/dW+gaPwiUbkZGcwkw
33mRAJy/N8FjMI4qR1+cjxColdlwNUDgMpzdqqymHJKAS08HZc8lfivIBFNzKtBsuWkVZ9AxfWgr
RW/Aa4XKbRvda4LnmR+8/AlF8y6JcDxv36vXjlQvOaTc2ksnppX4k7pca//JQvTMsVVvZcZiX7/v
0Wa3OaGiQcM5KQhabmH4MjtgwVYz0G1OvXeUO+ku8WaqXiVNjfUt00lFCBC1KEFsfJx+xkKNyVUh
8QugX9yH3iQQqA7AkvX8ZUd6e/1jK3WenZtXPZUBuweQ/4dSEsBBg9ESwlNSlurS26d5yswazM1R
sbw2ny3LcmeB2OF/D8sT3u0RCoT4MJ+PWcqkxj4l588S42Z4u0i53V3ydSJ02fgMRNmflCqAgjS1
EC5LGLtZ4Nje04oLJjCoSIjctf+IWZiA7Zv7EMnKx6zrTnkedeCcONc4It/HeuBhFDXvsW3HIwFD
lXjCUpyRnCfadkkOvoMDpjwKAhhomyvZNknHM+mrD4Y4sVo90Y80lulslgptg9EXBXDw3EMg3Uc4
feNsadrV1e8LkalhB301dLSL/Q2HA6G3LpbH/63En+SffLCt3Oyy0UQ7jgHhf8jAJekNKuTZTYXm
KNjw1UcvpusERjimA4DR2YdUJIuDQK+MxQIDLpl0X/F+LhQVomTs8SCrVlhXR2BfalSsYHqbG4ip
X8lS7GBzlAVrIKZ/WeKM8Kq4VwT8Y5PQeYvUNCuZVkTFyOIpqlcgS/QDw7/ZXyxCj4kT6hjD/Ver
G+XbEFacKOq6cWd90ESaeHy/teUt2Cq6VBPL2/rFQKMgfjByQ2Rw2fFE+mymiacSoWkdDbQW9S5W
4AfTOIWOjEXSRCRS1HAqJBEJoBHzQEWRasg+0EvSYbf9hrxQhfAEwaQUL+hWV3aF9s5G9wKQoJoX
xZFOksGKyJd3jtZzKzxZSOCFrSx/sLcYo7xsOPu1u1qfHDHBiVXV28UprlTXQ1r9upoeoMqd3J2T
Xc6zMRFZAiZUvXfVkHnzcVxvkOU2DLUkRQjY7sig7ZnuFa4vV3B6inoP54/tgyzPWL6EkKISyHrE
G5yDN5EtIrmWluJzjaIl/MskHhLTWYMxveCFxlDUNtP9xmq4mCuOHdKx9uGxrOhJyuYOx0Y4CAc6
oajdyzj36a2tLHd6vDcbikeKtHQPuedYV+zuy4oNL7NCNcoDv1OmaWukCVo2i5RBFGTDMOstUfBp
lluxICY8vcVp5MrT07d6/NgTcFUkQfupNMBNZPQu0Xo41jA5ibw2CLQeKWOBCMAWuUP+V10T4n/x
y7gu/NH+2hQOBnN09w9F+DvvvJPRjgV6Ha81bbEV6MCytfg9eCqIaN+AHzDIc/eW6yU/BaFkR/7M
uHOhDWWB6ncFDkvN/Xy/VQrAKD1R/rRJO1QXWWy/nlStxBMEbd8Trsa8zgGScu+qPbNXrVkvokI1
c+jerdKH0hD811FugX/3cKKbKO5ijKEoQWqPYbFUWKhnkv+WSWbQ0LiS+9Ek5KOc7/zD1RKbNPaN
X5Qom/puhb3OWktOi3Y/WlKVyO87uvy6UVY2U65MLz18hZyZFdAhTMixJnwf2Wx90tDOuXxuWmmQ
FDzMQ1ypbrfh6knE9qAk7NgloH3YKu1zwDpAgr82CtprZTVRUA+0ofPeIPLN/MFjw1M2p0sDdDb8
wVMPPrKQHaLPZiMYo9sxKBF8FCUjrBQzICGFzgbZjiPNxEyJcX+ZZMUSj52L4udS9T/gcA6dVqt6
4YHsHudH34wjkJuSx0HKNXATV/83wDsnwTYwqUD5xj+QaWgPIHeoDmyY+rYwXbM0tW8rP126m7HS
et7WqnhQNj6/a30y+iHY3Xso99d3LVL8A+Xqj5wvYv/udYlX3uuSAbX89U2rSOjCp1LAlLLOqiNl
n/gB0r3D2vgZUoTAKt0BPYPq+eyCadQNJK6QuOYfHX0yAcKJS/Vz6H2oUv5ywBt7pRAboZOTwYje
DxIN4YTNBuQUFwfN8uanWm5evELWybq+OIggjex86wPSUgrZ81xgfuK5bt2uQYOeiMkc4VdNclEd
KBz9G00p14CXhj0GTKR66FtR5DNLOhWES9ljANw+tYcBV1NHtWJOvhStHXOTMpGk+zsQGA/m3k3Q
EUVYd9W1FHISV1dD806VsUt6b8UGVKNmvO4c1mbQY4wN0Ens9vmq/RyzCSTTKzsdJHlz5bwSaMvM
a/psRKQZS0w2pq2S3q34ccjgaF6z33xTw8FhOaVxwr+PH43VJ92o7FhdehfidODXR3kcO95tnthI
N1pKFOZyBq97zVBTZ1k7MJUve2Qwxjh5pm7VlJdSOohc0/vKN9GxYITmlo8h4c2rF36xe5E8mWbO
pdYVsO1TMLqqc0M8td+kOhEeRObyy1V/+QLAN6ZszYTJRRaLoRl7IWHxB0ZFq5o0OrmVjMuJ3/cj
UhjeksFGX15tAuDige3aQB+4aCrqqltRqwJEcbKidJeNwbSjB60Wbcuxs/NbHO3eUNinIrPFAhNa
3VihPNA+Z9VYB/wYbJq5aKp3Jd3NHjglYunESQc8qEiGIIfQ2PvKRL2uJ+TNhJzV7A+yHEvPMhKt
EHRXZZFwOPD1I/mJRKy/V4Lf4R/t9yBv+frzAPpl6WgB6jJoiDhmfeBcaUvHk8DDrWIeSt1A6B7p
heY9z/RfqyHbW0rJo2TgGpFl4YjrTvK4kJY5IyIBOJDxFZqwXpJfrUDa+4pWf3YlOQ2pgaCMwm0F
3BlsRAPZ8VKE0B2/1v6yOhu1u8v58CZSdZ7ueTms9S5vOaGiKLQ8QPSsfxHoXx8AKqwK4GveyZ38
E09XIc5EnWhCM31U2X+Z9wpNvgkdY/77YFTAoFr28qzxb8DX0h0bG8y6Ts1fhBb/YwHI/KRI2hWv
G3aiyjKJhFOtbfZIAN+KhpuYTe5u1nYOwXc++YJNCafpex+XWD+ldTN/K4PmpzFM5xYw2c5Zk/hg
Kz7rhonGG18HMpTik6tzjPW1qv3lUiQC5D2HobfJcs6i7O/107tNIRu//hrg1pAmzxDRJ18TyX80
B1CBzSgG8QdW+CfV4dRBWl36FqEe0mpcM6JHxCJ15i80iyH4hkEDEPiTK6+x1GwBhMSdtr/9YSfn
g0TAha8aTaHpxlv0apbwbYXRv1tYa7UojFURDGoVdX1xPC9FN/NuF/AbOuv7P/qohh/bJNNhbCSY
zbMwOSrV5grN6SwKKMNCiiLzQKiYaGl0AmYDjmrbWpIezcCeCizBoQcYsEa+fJOMoBEVOjXglfHM
6Fxmzy9iy2+8bqvZIhipWyz+YlhwjE0VVdqjBGwTBgTMCFuDYuRj14WDcdDIYoXNEviwir1TpfOj
5nj27AVqurVrDtSwWvwiaLZp73o5yqN6xqRP+dHAqYj2RX721+JDopGvxxU3JCue++xhSknKYBNn
na9zb0gdLa7rEZcYk/4bST0W7/lK/tzUJ1M4HOLAocUBiLVVhGw7JDq88fZ7nmsll9z+vVkryF2e
V4ya56aG1jj1jXQ5kA2ytcFf2hzC2FqMQwUQ0Pn+WAMrSf9obbl6vPyrWosXcJ2nBR1cH8EFy1YA
BHg3MvPezWjLwcfx5C3mWjfyPquQPfYWyep6/S4mQP84PAJYn7ue/fEJz8EREddJ+d7hCUps7r+W
4EC4FvqjG0ZIe8Fl1QAbYIcjCM++lFluMCPtzUEG/5v0zctJTT8RMxmk0jCbUh73EZol95hwNQYk
jRacxTqdfMrYAnL4aPbfkR5ZOMM/TRqOrZsqThh2OUq+r1x6b/iP++hPdwJBqBewjkY15X+c9p5t
DQTdemguo/uiQbUpwxDrBTFUYUG7rl0cHSeP+JefZsZZAblh5JboL2oSFXns+Ycjq3+PRc7wm+k1
8oVpL3p7ZjSoLnEsxxOtHPQSd3tjLbpjmqU3GaiyqYqbvw+3EONxpQfX8u4u5B+ruU3B7sbHS6d2
H0AUH5L3PuMmh1qS8sJqMjj+1HjtqZdurDVs9aJb0W/NIcT22uoueOl2+ifzBUuf3Bz5GBchXPVn
QbSHs/0pRUpOGVzXxYpRpwsyqTqsHTlNpkgdBDJLf+0qHnGY66AMuO5hrwiUSRL0BYhlUxM8/CXA
2g4DSxKX5OjWr1Q7gCggnCV+VOJ6gASkdmQKIO7dQyiVDvBWk2ha2aWhDktD1cmeePakjsk60WSA
PXe+aIah+MAhRYlvLpxxBe1EcvzJ8fhFvnjDoIXDwzRe9QjXDNXcpVbOQPjhhK6LbcE0ZOotNRaO
WqLwovQEcoqnC2Bi6o/WB6U6qhM5+u1q7FJEtglwmKvTHVcZFFyXpJ75VkB2wmXIyVAilVrH6l4w
mewUl0aw+CcbFJDd3h3FOsg1tuSMsrT6uTXcLsGhxvBQLUXBYyWjSXJ9z2siFY0dzLnPeXduRxl0
7HQB3WF5sZHA8SwGQr+Kg4bZdrT78YAMJtSggvxWx+DMh9oo3cmYMvO5PUf9DK7SaGs1rvVqhMt+
mjpiRHVqZvBgFheUIBzOWHbPFAcyspS7fmmfYgcZLSqJHdUfwc0qm5G71+ZiubxEneTUL/ZUItXA
DxYs3cCxDJ1RITyL85E7iHT4xPYR+teMIVYBwLzlCuODiuUMk7FSKBWnXepFK6KYqRuIlD+QpVc4
I5SDomqPQvt+aJoGEH12QmEwSYN3SPAdbrSjmAJfUbBZT3TXGAUvaNZVUZvxE/mGvKTFeXnawUNl
6PqI8tjZsJypM3FQr9NBOnv+IqC24zDY3ujxWX821KyKnnj17dqLeeqZqR3IGnuVC/DdU/yGRNzR
m3HmL+uTh16GeLCNvbXHG/X90g8X/0OBitGbDprL6fGcnSbqNgZG35zEsJAYoYObrfTh7Rz6QfpL
CmB7kEB5X4ypdxOGwKgWJ5XDC2REUJcG8ZyO8x8bAU535bsEdjGkf1qpv3/ffREQFdvKIub7fl25
FJXGPJHV0Np55dmOpHdXALqwAyahw/kUxM3JFnwmKzW/PtWCbCNpaK1S+w4q+M6u1vFmBgLpKpN9
P8KpKdbGqAAyCnpOk5O12VKVmmab8WukvEsniAhP+IQlo4jLQ1NdFtnJhpXejafWKjY3rcLulUSp
/5/8lInxzbZ2W+b9sotwFWoo0XPYgAsAYuucBZJI6n5GPZe9xjnFA7WDCBG2oXGYQKHnOvhQ5eyU
ewuv6vrWdvKrA3KQfVzEmH7i7ffCIwBkY6+4kleb5t+AiTARI/PsVgdjqJAU6bL+nQQ0EExhLkWy
p7Y2L83blwiNwj+HhoSKmoHHsUIQpNlNmzxrR/SEiIwBdGgyix+J5cW2FH0htRQkCgZuVSw2DIzK
hc8NQvnx+OG9LjaocXCumHLgl+VO5SLS6engzRoidFIIF1dB3d4yjEL9nt/f/8wcnOY4Hr/a8h6m
YEOhbXNgzWpgEmy0t/nvrRn/dfsiIT6RADQ2ZGpRVdxKSPJYbL+WfaEpRAtySQQoWm2odvkkdOT2
kdsSptPuV3nPE5Keg12mJ3xvWIVFt7rHdCF12Z9JPKMGcTDxNa6/sMTPnccPtsbHdEbD1wbu5pRA
rE9nHAklQxTxV5grKLp3iofqiAgJZdW80+kI9tmbdAqrERBrmPgSno028iNPjiAZ+NNDnG5UzhBZ
0TEY19ghIGUeKB4ixkbd8kHSvMWX57oQ2zLlk2XLXzUFPORVbNEslt3wO8XK+FIX+2f3wWVBNHqz
/WhKrdJChl8z1AjAt8831IfnjRgNBNi6c+FXaWafXopAZqExGI4xxRyQTgl70eD4o6/sZNyof4Pb
s03jdgbugqh4GrROG3G+tIckE0HLpWDy/ENs+ywOkgwLSjEhCr4h2GpoElDOUCXM7GF7PHVx3YXS
+vQbiszV33r9fTK/nAxRN1JEMSs4Ifmc0wOlqcDrZq3/U96JzXQilGB/w2mFwrzu5mrvqxty6U7y
/2b+UuKLYlGU0KeTNaaulyCoWjAK8uxYI1G57JqJjubrhAsocA2xKiX+pzR+6I22tbJovZ/H1ZVw
q+UJ2Za3842M9VTdhUdyv3beeNOcFew/aujzObJDQnW6s1NLO29p4jzkBOF7k+Y/K+UTM2ZVF0ik
yOOft0EeKkNp8F2RNaMeqEtYFxvot0J4X/V0zZsO3M+Vykksej73/B2biyvTPjl6RaXJhu6z/UrS
hOw3cgmT+iafh7wnyLVVIZ0nKnz4pBGLtHRkwH7Px2uqFqkOqqozh0QHpN0DRcpLIRBSI+61HntB
/1LRIftbRzdYMI9dvxvyIW3KBKnsfae0vszibVLHpr6GmTti03pYokSNXOg6OhYdMbGjq+Y0xIsA
vm9+WwzgW9FOtPvTZYWPza4rxiFsczpTuglXoXD9lQ8+If8nkYkWq8es9kTOX8BfORPw/qAqKe2V
JrvgS4ssulOLV0IptWuJXAOgxrZeMfSOQhfbKtHnCvCjTpzKiTLy0CSczuFIpsSHv5AYQVebo4Xq
WSTc3stCWbORbNZd/WXk1XyxxgtcNj79XBEvMf31YZDLokQ1WtXZIXN0i/Xm8BRnT2U/yxizP4Ve
ErNhfQ8jnYQVCudMs10wFpYbVXaXPUIQxVerL2dPhTQSEc7xrrkFIJCWH+lHDEdkmw1JSCzWpoLY
lOpxAaVO/sbCKGS41hqpiEXY4Ty36Fw4AM0yJw9F3nLXmL6OR4AiQXH42jils+I+PdG8EB8yEyeb
yLpOPAYPQJcnj2tvPvNx6jPuoNLGB4TDOjC5/crh3A0TNlVXY+SiBaSNuoLs7MRZ2fFMzsa+6jaE
k5NwiLZNlFtEsqgRjUnMc9EbrezEnLa/B47UvXyeU29ogV3uQoWizsk4hzN817Floj0jdOe1aXLD
YPERmYWqq8loJtnhsN239pAC3mQqZowFLM8BU7lKFcy6neuY6FtLaqZUaBKjvTYObKJWcOe53t1f
Kka/amqebRp88SZxjBZbOK8W0iHHYXX65BR600eho1VdyyQh7CY3ETRoj7mzAwZ44K3CDBKTnZt/
yhD7Nd/7ArPNAWqpLK1R/Eoxj3thvL4pQoAd1SINuVZnFJodZ1Tj6nC9FTsnBiU/RG/6oUZD7a9h
VDmZp8Ugnt7X+TgOCe5W1PZnTNM1DPI+xiWHQDkjxEp3NpLg501+JlT7UnVmWi6zmDlauoezfj6q
5CXadDUJuE0oVVPIwHeJCmcrJZq3QVoaKgSbfg5XIFcGrBIlyQuwH0t8WhKN6wMyACQuENqH4OEF
BePCQC2wYHzQfR5Xse/9vvdRRsvEVCX3FVnf/EqjroP2ynFkM3pPAbMmsH3N0kCG8CzSyKYKb4Qu
5GnIaEAPNt78oTLbfYG/kVcAMyaEoYdU9dAPDaBjW1dVFWyklqfO5dJFcbEYEKEiSiz/pGiI6339
H8zAdkxxGWboOiCQXnaenVBH/VaAWjDSHxY4Kq40+bG3VMZgNNSTXA9umXfGoUuUWUaOYEg9DNZR
FOi0ealNtR+TFecUhS1lDDzld0cNnREd9xZXeLLZUsBClpBtB7ujtQIJd6i2xf+7JJj6VtFxrzTl
QuCV4/iwRYrD2FSejKVNjMxQ3GWxdcb2ZQIlyw6W6tV2kYGZW9IHT4vWxRmoluthQuC9bVqBhmcd
3Gs2nrYd45bbBPAUHuAixTNyJq+MxHsJoYGdeou/ZUQaaea5iHsU4w3IIY4Qu3I3Jy8UkV+4ZgFp
KT/OAj8rH+h3Zx1ULLdBYZF+nxaq3E3T0YZjET1iumdRsX/GVWoYj5r/Mq05KVpGutBDmuEULfcx
9wHvUbb52U+DZIA7FK9ZST2a9vUZ1jVwe48buZECpVEADw76i5ub8/jmA7wAJwmNJisBnCKNNSBP
XVg8ss5KKycj7q37Nd56gtt1ud8a/PWhP354GUJzDgIOdRdxYQ6v8a1NMPSaoO7p5jDDEC0Nkx5F
0MPd/AtWYyN+iUVQwgk9eR4con2w9L5SyH1V8n7H3DI6CzmVhmYv0Kh+75jFZQAfNjbeVT5PTIy+
9/tFTzbxGfxDf9joY5GmJDsAIht/MWzmdvc3rBR1lAN3IOJp2b86k2KdfD0ucHIggVTewkg1sohr
B8BwxiggxAPhi36uZuPyiq3wKaw/XZKP418iUoPHN2kN8nDHcyWmcIcD1UaStv5xUhyNjWRQ4tN+
KClCFEZiOKTly8kiHeHxhaYX9D3cfkd7RqxvhQb0Iza4qO634UD3muOqHCak3RLdkQh4uoJzeFk9
4TdE2UBhXqafMRSpBd0eMuWWQEaAC7FEOQ/iXB25/oKlSEK5z+lcWG1CNqVsMAZwgVuxjL6TrGfb
897OrtOwfSdFUeD6Gbusf8E5RYYAxF9Hj+n50sHCq6BziKvLMkHDBduM2AOPPuHEVuoMHpY2ymCr
+KAx41RBq7pb3OV5XjMvFVQijzFxnz0OvJwy0bCjT8Mvj6GnGSjsCe9Jm7gntt1m5f3et2VteUou
ooeY4pzIYMntn/EzlD/fsnmX1XquZvuF4rCadN/ccRCnhPCpz7lUXaqhAFQuCe27O5M50rjLItVS
jOOJNl/Ngimn6urLYr1bLxlZ8mpv79qWOLGp73yq/4DfkSrF4/7Za6IfMj+87cGJkPu1P/Lh2QxT
PGx25wMINPFapsYKeEWPprxyGhoCBy01Qo1SjXkX3O0wK1OW8q9UXdNFxrDNxn3Ejo2ugJcdH95G
GXRpqbDuKPbCJhbsdyokN9e7+KxIt0N7JCbHeSY+AQwod3gLzzl/iX1ZdN/lWkYytkIp7jqj5gVm
wA8bX1g9YzQBmtjBMwOB0iep/gi0mhB2vAVy5dwXDeauenWRf1I7ldaF5rmxT/lPzI8kfIga/YOU
5BoBN3VJaG7rFzQP1Qm3eyENn5sIg0xejma/f6sNC+S1h3SsGhXZM+E8OmxUZHfI0MSjEJ35ZRWF
2EP+ZuEmN800XfGobfjT/CS0QgFb12kKMxVyrQG/naCCNUXTRzSapINw+8gLEEnD3x8Z6wJtzEUW
rT3H0uZSGp67gszcniL2qk99DovQ0QpqgMIcs4ahjpYUBImiT60UvNL+pAXT/e+o7C8HEFx/6fan
1efUjD3hxMVL9eUpPfxv8NKiwuOMGNqsiTZs1/wMUX7CsjD5VrgJ9ktveGL08WrI62PzMI6CjrFy
9j+fIxkUwSU0yDsVRS5THuXUQIZ2K0oR9fO4scZWFCeTfsn6mC2fAx57U1C+W3y4ikYLAnHq9nUc
J0SH3NS6YAcS2WrKJbDP7zLf2DA6cg0EOzvVemIkCEWk+hFaLENX7pYJVci2hV99bcNakjo6PSUa
+Oc+iUbBgD8TmwprMbyXqjQg+XuYqlqsQBNaRc0aanWdXoqmuc7qvp5gc7QRm6w1fU9jI1lD1y4F
WLnCCbq83uAM13NioQ9aIoad02iTSoqluomGGG4YqZ+Jp0CSC7fjwduBaHVBNb7OnN/NTeDJ0rhy
DxZ7SGCEZan0LtoB7gIAw+MPQCKZUlQjerg5vHN7PGDqIlFA1A0MKRMJtfM6s5ThMZB8US81HVgi
wnkhjaaYXGLsMLoFKq2IAWwO3+Vrhi+CoF8CWtoDjwCiu5EEJ5PmPJBU5HkP3xyV602uec/SBrQe
6MQsDTXJRCu/qnuIfRG5p1FGeNqe8cAM7VW9tEjbIvfz2zPQImmL7X3Pv/6xhgGsX+q8o7yM/7s0
0Fx37vc9okYJq4ZAexG/4bOyqQA3nd1GGqFl4KH/8HGcR3goBwr/h/ChxL/wgz8tqgPm2AKyCXF4
m+GtkOEw5dR8q/FgFyyC6MYG4+COIpc6UhH6HYP2S5V7vwJv1CwJcSwnhdqgeAThLxuaJVhmzgG2
JUGEunNuVjocyk9lymA+NPIo836kuVUjNoXAr55nmsTJ2HG8dcXdoCD9gXatdPSc95CrmvrpPMC4
fXzH33YqhosEQklIrbLFYTIiQowTpD/ETF9fZkES9flSfAgDPUpZ/jhWbIuqb8vn34cV5DimprXw
tE62uH2MCtn9SbfWj+Q3K1erNSrNC9nxprFaC0lOBLz6cA1fsWeITSOyQ/ILg+POUDcnzftrlCO7
A6knp8juHS+Th2x2FldiUlAgoMMK/RtgjsmxWYNvYtHZ7xfrCoD2NmyeOP47iJFdj5RuaVdIqepq
XumIor6NQbkSpMFGxtyUYMhPcWraAlYD8WggUduEYjzAhEfjZp+qvQhEE1lrovYqOBgZav7NbZAg
84a6Tg/KCdLsicMTw/Xw9mKckRb0plMO7Ihd9jc1RXjxCNj9SI6FkkzfNfXySwKhS1wZI2QB42wq
IcJ0G7Hl/MQ3oWt9l2ygk2eA1uEaqgz+0yFIaUI0+aUENexDc0iSWX+1nXVjhP4CvdtOlE/nbPqu
6ns8H5uXs4JiCKbJbNsZchwVxgNyuQVg/hzxtV5GcahC7pqLU4xW7GSCj0tAXu03wX6dCn5Gy1iD
WIjOTwXK2r8rvzDIJTMtZCFlqr8E4sAVPLvR8NbTx7bPCTxJupfJkVoJxp7IYhmXbJRjJYMl6ToX
NoB8sROJw61MJZRastzaWX6LPHyQqSsEE9zi+U+bnz2GKAcIX0gDYFv9HWbcuX2Mvan3AHd9bl4K
plBUvOhW97dH4pUBvwujr0u8VR9kInfUWVO1wfn778JotR00UMMy89gVUw6rKzXI1iGhAWq/ZJ45
7NipNlUQrAVHnuSsvDa3Fz8nuU4kpGLKVOQ0hixu11g8MOfBd1WOv0DA6hHQCKtHLKj0vsSBVmSb
rnLdU7pi8frl3heT+M+UN21QorRs3tsetbDfBG6yfsb5gq6XYoYH/ZHYWpKW+9oKlDBd+5KNCWNC
PIMn4LTycDs2k1aEo5XTsFSoQv0G5riu2SXCWHxp7r4EJqdNWqNymusyLsYHPpbGSLvtXj3WWxUj
CM/2xx8gNRH4V0h3iGVP0ZeG7U2OYO7v6mJRk1AU8e3TN8vk9QzkmUDC9LIq0gWD4lgLhrYbGhdh
gAfa8Uac5W60QGpl/5LkROu3WZR95rXXP657/XEYihKNpCHiXS1PMF/sc65foO+ZUoY5H5+at46r
DdWVCYMU//8I92+LaHKeXf7lbfmoZmcdCgVqKV6+kAL+I1/JYSrQMPUEBargQqL52KKGug7oDveg
NDUzBCEXNLhgWP6mjXEFqK1StEZDnq4aJOM02RM8L9yeXYw/DbcwqENorusWym/siLQUMeaEuCm0
QcOOyUoyFU2fNZ0dhmHoxHAnzV2b689VSW1UffY2zcZYqeZULw2s1FdIHWngIm8wwyrHF8J28ZYo
2RMnM2XQTg0rAexa/8oh4oVnhCIELDVs+yPwW3131Wh0/kIYmhDWcV+7U+daxckKCMbUfjqLQGdr
pRfg7z6U8jGpUCX85y80Et6x7eTMB9NBjireZUyAXJYi9fO6rWh98y7luQl1DLSL/ch+RRV/XXRg
jpxg9pnW591JppN1hGmILGkBVTLN7WSzPsaMMzr3gHOc2qhBBy55jzXwoWbaF2RKvZPAr2WeMI/0
K9bVNGWiQ8/IxRRR1SRYOZuXSSUUQmHay4/JPhTNCztKNgWekbuQEp9DkdJBFEMOaZr+cNv+PEDW
JVkcUVe4kifebKaFky1nvBXLAq87oa6OdFiG8lGK+KbAvGz7fn/6+KvVrgWjWiz8gDbLN3OqsmCS
uwIHRnQJ5TDYkI0UEo9YZ3Zmo5MIBhABams3tkOrJsjfOUSiTGwQsm1vZoHerS2uaF5iiJiSCKan
5j/VEgBPCrJGCgMS5AwM8kmqw+8tRfq3TK/BCZyoSz710MvQ5O2hxb9Ap/CT+QO3+o3o1OGjeb6i
uZLVZmNuJoD6Mh7x3MK6G3ly0hC0P4nuL18Vi2mfgJ0p3Xt0QsHdwa2rMAGBOvXSIE78iuKoESKL
OO+Z46McKrUInIvaqgmEsDigMsiHpq8SyAT7PEeIG/1y1f4GY+FVBodFob5CdXYb1b8rSmIL0OxL
+qPvcDShjhapihCPDBoUYHOxFcj87tmLEaZ0ui2euK/uX3donZAGchKA3R9DN8jKcLn6sdFLtp3h
Mjy1J+8b6QgTw1WM5QvA52esbg6V3lxMdHd9x7dHeLtzQMHJ0L+KRmGjCptQFB/eOREeGXr2rvHL
dZhoOtc1mmAGPJ9S+AGdgW0rBdwj/ywp9UVrAbIk/A045bSwXKx4g8CGLjtFrJeoCSYbN2QrXUNC
gAvEnApj1b8RLSH1TXDq3Ky2ckW+tWl21nj4dCfzmoiP3qi+H7nr1my7ag067rMxjz1dnjJl/+EZ
o8WETnEbHFfOgJXfUmtEeMiI0CYUp0QN9ZdeZChQlB99F9O0gd6lby4/GHBAQ5oYZJJ3M8InZFe6
tHO7R3KCT63w9fE0OPMm884OFz/vcF/8BU+sVd86euaxhvknlVr+grf6DQDWoyxnMG7TlKfPVWYS
+6njtwa2aL9DYnptol7VnEaUYYb8HRnzMrHQK1By1ewi8cloEXnVLC+uhVjIfdpZt/NFlL8mXUmO
pTDyddASzbTFXh8xLXG1G2jH5THy+Atvk3qf2TWL4RyLyzrL7CEZUSMQ5/TMXEA/JrQGY3yGiXne
zTeersQAes2r0vxjBjIWbUh7tvXNsewjoP/FESrWGonbqb+AfLIhIr/WvcD94pIhkkXDR10cX8iH
WinYvk3NKhEjXdbUYQCCmz2/p38rJoS0PJIZFkEwAxL8LP6Es8R+yeOwEMy12vW+dTwayoFsdZXS
F3yIMlWSkzphuJpNjRYUvOr+1kIalhM8SbZSd8W3Q57xSxGErbh/l94SMk+QTx+3SaIK3gV7I5mg
iz+FXXtM1uYtQBnUCnVfRWY0RlORsSgudikRTFc4A0SVrj+DLNQlfpZLs0EacdPeQh3lIEGXIYF3
pORolv/PCBTVZba1+N/dp75X5nOBx3gP1ZjUBbm3NC44EPpsl+vdQcb+KLw5rXVgSou2RXOWmP4U
ACYl3TFf5bIP0Cf8NFXNkbSVyOHW+iX5GLW2L+GGt0S5lDKWM9fOsU8goZRF0nAdlsxnKVMw+xCZ
plpJXTyoc4/L3mO9sUu8VXwbLMixeBwWevHAL4VOGo6ey2zu25oELQAMVCuEbN8SGlPeFIjxHyIn
EfIH9o6jZZ8iTJhTy9lXu6FozIrPCRpjJHivqElD0HuLFOpnHYyE6ax11i82vUKU6lGhL/dlizHb
fXBKo+s9aRR620NUPrG08lIWfTum/VL5ifH77nFX4NDCDaF7wd+YSoKrAeJ2mLnu9Hio8/Gbgm3s
KJvM9jnG3XBMzM6Btuai0LbjoQrk9Hba9Pvhahkht4M2y/V3yXkCQOoy0VIA94KdlORvTlAR4mkJ
AsKkhKtMjOM2iz/3vct9z1et1r1i1f2xArrMwW52MNVtRryLunj7ZDVe7iCbV05mrqniLEh8oo78
/KEZD8kcwYCvNwEG3w3qyDYDYI1ralhvpD8m4nibDDi4ofBHys22aF8ZAG2T2vYXWiZgrSfRFfVU
NQuw+xZBkt+15VHqQJOwtLcKQ1hWf4EASI05ek0B6YHLqNWSdNpJ41SDgp6AnnY7kjuqgXHEoKAY
IPN1wRNW7MpG5dcpKQ72/ym7D7LWf5ey2eFsPQ0Nx3DPfL1G+hYEcRR8oBy/CyP3bYPsPX3119Ku
BGNahS023w2Pg6lp1nYI0tf7SnaIHJl0GYCEy3lOjBErWDz09zpjhTlEmVuPOfXUauq6aZUVoTv0
pqUIqp7agdBRPYb86cvrja4w2Vnx4iBC1sWx7l0QNVc5ZPi0crmXQjH28vVcAS46I7Mfvqu1mcQ/
/kan2MK52MywnzwcHFo1yVeIzGaUZJ4FwFTCs7sNSJjk77hTl69kb1Beqyu5dIsU1y7OTZHRxJX9
L+koI+7dT6EzeDTfsJA2TZd1iv3FOgGXpoOibmG1hD6qeYqG2/2Mcyz2XVCP4UJnlu3CEzGl21If
2Uj9fsKoBjI3XUwAXvY5Ec7v6NBjFTaYrsyaZDYf/diAV/h75/M3jFjfU1Md2QLlndJOrz4HyEHT
hf43KcjP4/N9UOS+K+mv/a7Ky4yVizfgucK3ESwN3MIaw12oAblCjqk9ej36AwocAdiAKVGrBmWe
y6EdOGFAlNNNQTRtPY8xfmsgYV5lbfUjk67TZT8IszOpWSCP/lO3eQJA8sSS3kMJ24e0iPVZXEt8
5zLjmfZdGcdmYJKZfB3mbB+VQf0mbdSEYLf6kJ/ctF32td6HZqnHbukyxSFvBPKFapHyKpCKQjK/
Bc78ukYcggdtddjJ4zQiOZlsSTL/ovLAuPd8b8sYyUeSNyLnroU6+6a1QqhK9MPpX1syBDfTtcj5
IJ9x/Jy1FInwfy55wbb7fDyu/x8DXvfhZEKxqgW/KixAsiILQ8pAvRkT2II5qsnW6Aba9FeU74PK
zAXBxKq405iLHaNIqSC9dioMBWn3lyOcmMxxGlFZYDQN/7J8k8aIoUdwayKqNKkh64TRigPXftpg
PejUdbYvAUMdtSLa/uxJ3wvRyixlUShMfwc8a4G+FxaTziED1E9RxWpBhmmYjIK2eVBXr5/kK8tO
jDntLouNxaRuxfXdVqG2/BZ+tMRnAO4f3w+mmB0SLFQz4Sm91fmD2A8ei+lh/InAZtxvX1iIS5tJ
Y1mSwXQ4ZnYUBlcUUS37KAOHc1qY2l/P6r+pltmOQIhQfwI310ctBZy+O6acyt0lSxKxgycFb6hP
/+1xqnJYrYP74ngmEDddZMe1rusmBXd1QhWMCfSSR8ZU4ZbXHRYzfmIs7u+laxJfdFhERH5yRGwZ
afm8BOywfJqwdrDeN+/0hjq6o/n9mXzOoGbbwhFiN1Y5jx6iPme/GKjH+auGUxYVIokfyKP25sMe
mw1OABvktHUkzBpIQhdcWOBnoz26M3KEx2BpaZwVFGv/bEgEVIRW7LyDwvIAx19ASy0WGk/C3/WD
luw8nL42i+uOT4px+ryNmWLp/hIi6hTv5EGc5mFv7XRMxANCG/zAmJTvTf8scbSRP0vgXjVWAMEo
2zxLRtNUklZFUJlkOjZkiB6SqDqOjFx6U2hNlbEaIyprlwGcaIWmha8Cr+FSU0iMU+xNoTp4T3PD
CQgeVnPSE/pGqaDfcVtTyNP3v1lWQ0DFtl3j9Iz4NkuG956xzBXU575eWAbGnlgY1fwJDfpHcPFA
FtmfrT+i1cnO0iU/Lb8FZn+NHkJPGjwCbccIUGLYEuTwJwBD9UnOOHT6aZNPOFgq78iDAInLeCJC
HX8em8v3TZ4J+3Pwdln+3IF8jUsiReXVXJb/cwV0nb1Ki81Ua43rIn75tzQJas11EiyLm2p/mZcg
YZas6nXr26jiRVCMToJyTKQZJKQJ0J39gf996lJXVQ6GddPD4u/q97lFFAYp/ZFmJnkFNpIqIdiE
NTNTkc6luL9TU4L3OUFnKsT0lIGhIJ0krNPCo2Wr5khB//Mgvxw7NnHDYLtAcND7hDWOYjMWXq+g
Ofs9rv/mLqZ9FIoJ/hBcA/xq8QYOM9bqd/voVA+k30Xkd74S9N22HW7dIN5LRWd/cEKEyY5/QE2v
Idr+jDPz9NY02PrQM3STsm1Zxo1XXQXDmdI12bKZnXIzNtHslHCXFCl+69e3wpxNacX8z7lUCDcM
DDqIpPHf8BAni/UqALy3DTc7xcgVILqCXfv1J7AP7QIq6G3zgQZLQ3OaU5KVorvek8uTT7aMuQwE
hr8ndv1UcIvmCmla5xPHG4XCOwNkdITE8n4RgxW9tI739mGv0QWCwHYES8ZbkYIq6IYi4f8HfDcc
qiuKWErRAO1aXaN/5GdDZmPFtj+CGBRoOCGHgp5/ZXPA5it8y/JikP1SwNJWWmidI202qaxFMTC3
OW5AMNi5pkgiBs0/DfV6XjzHGPNigSAQbHhQtqvB7RWe6iCc7XKeB5bKt19pP9zXCiLUnIG74nT0
Cq3uzhEziGOOb08la+TfHzBlJIzbbOeOHnRb7EhMi5MAUkiC45SMXATqDmwXjETs9HBY+/+pbk5Q
VJz3mZzmzT7us4Oj2LA3rCy8DwincjFfDUefN++AWlW2BDrBV9zoomEr5GzhRfBcTFzdGTSiGklD
PSJevO/WsHetaBsWqnX7wUfo9Mqyx8vHcY4ZpXvGTn8h+nxmK7prILjfRIzZySI/5p+dO196OEEu
pP5KvN8YABnLjBZ4LMPVtBYiuf4370MMK1I1qHkxDYQoIsRLwT2CpzO6SCaE4OiR2DQdm1JOlrIi
Ijl5mTf1zrw1B9J+AitYcyxy5U5EhWEikru5+YEiNTUcuxJuLp/F/vJ0YvGo2PEhep+uKZwmr4u3
pDl9GBr4CDSfy9+80JC+MB8xQ3lPatR/xMVC0lcZqpB6pNex3OamYS6o3jj3mJORWdzVOaaSVEQx
Lurw3xXWs/5dxNxzcHGgf6qzWZC5UE6L+JyQVnfN+vf+kWAZ0SpPIZu2+c557eilQKze/esiLrYh
qpmgqFJkmrEgcesvsCoJmIvnf1SDfFVRh7dG/UnObLMsipzQ9rd2iwdkJWLfezIj4QHNv1AAAlIi
4Bzu9HjjZrHwjKSBdOn9lCJazBsHgN4hl2WYThwSXghX/mc658GNAtU4k3OYvOz0JBQaFY0sbl03
eYzDN349wZFdq6vxaYtTK5QR1+OwXvzcchNT9Vpx9uRVorh9ddOYltGAZ49ig+WGwZvB4jktro8z
W8W6K8vSCvyJ9mPWJaL4PInkrkjm4q9WXKpi/ChnRruAwdUv6fTYUGUlrq+iV7+xw/aHxMraG91S
+ZF9iu4fhH5oWgz/UWlFWkDfLudc/lsMrLRyPviCpLSPSEyjklSs0yRbZUTMc9dEXUdJSuU9zN1N
R28JpfNS+haRHmcoVN4gAhqxndjpgwF7BMUxLWP+LvmpRNOA0GuNe7E0BOisYsfmaJ7QKC91v37V
EgLv8m9q3nIDOeTvWkQYNQ1ezNXLJzjIexRBhj5b+BAG1paq5VC8XScYRriIfg6hFj81GeT7eQUM
JLPiMYOLvbpwxWUPwPtvq/tNru6xRzxY+3Wzy7CglQKmyIqHGRIp6uYJEaZnrpeDPjfFEuLCghog
wkmUn5nlrK6Ic5yEy1JTMNaDhausFtTDDx3jro9Fx0/AlduKDy6ZTmfjHTfYB3iuZwPR57q74l1c
v4oW2hEV08565hq8RvcXKtUK6UiBBfgsmtdKbTDA4WdPOkobX3qS3RPix2mEmFqW5j7ZmLPUJ/y3
DeuuRxizSRCCW8/CqHx6f0KwAfsaUzika/PX6Qem6I2VVnzn5GQ8DDBRgrACghpLIlBtrnnc/YO6
FYv0oQveSppUkVeS56K1yGZ2oc9cB2it3V4Hdz2Elxnq7qGhxAIc/O9X4hQD9sHwAmEw4mKVyJ8g
vLuqGBpM9tJC34NW/1njrguxrQIHkObeeeLYOk+p1bnZdfLtWsidbOz+SyZLPnzJziRdAIwulKdB
VqaeA+ZK4miX2/eQPa73muzDOzDOYAL766Pv7M8+N5a6iqDrl6jWQbsekkaLgd3A2Cipi35Q2i2k
q6S/irxXpMitSS4cZ8b/j2duohy0PDnoZy+4mVJru6gqwKg9RqUpQmMD7w3U2bxuETTr7L11aZ4l
Vwo2DIvrcRyzJDMmJSSvE5R/Yp/2Lu5R0G2JV4AMUcQ12qWfpxeJq0K7mWXtsBW5AWNSkxCpJ2q3
XqwudxRCBbfHeScmI1mUqZZLfr0XZ5rviWyXQx3b7QfAztRyY5/NxDlaqSQ+6mUWllK5cnx4BpA9
uGgltVjg8vO9WrtfLwN9EOV7uILEdoKqF2CcY0ClAOG7NJXEzBoxmEao2Fk7Z8KhASMGLHP1B6N/
43MSmDN1BZP0IvtszYNHGFeQwaLVjy9JJGj4kUlIO10qzIwOw710NGRWZn2/xXZ0xGHnCSgsYSHA
29/Zam09wZxWCmVocut8jkM0qkcjLJ5QKC2QimARD8QzsihhxcmvHckghVnxflGxxELf931rePw7
Vq9p2cNXxIkv2echmcG7Syv5hOPMQSAR21G7mbjZtceo5nNC6vhtEXrWRuGKLUecfPVtUlhA7nmZ
EulWWDz+rC7dnXirUWwOj6endh2FXMnl5eC7HRg7Rb1upDNe6LPd7XKm0XGahFIOtwrTI//ZH37D
rA+wCwV1hpPIKcHkWiN+uwP1GkOggTEZ15oZf0RayVsjCvgHBm44e3zvRAxI1R/FQgzGMDiwf38V
u+WNKurN8XNrMfCyU8RaQzOg6uqkUQMF59v9tV2JWQae/PcKxwpNuqJA5YlW8J7NG5623FCDejnX
YTCMa+pgs63NH8GqMCD65hXTJzA966uW14ReGb8k2iL6/TFbEB2deTVu3xpe/320aBB6tRbY4VTx
rDR+3Mv4JZGNuRuErod4DQnTJQx21LrWHN8O70UFrvH5nIEvMhImKX8X/aEPm1siC6sXwiHlUWct
vvjdceowiTQIW3QwPy+H5EDDzX6ntwGIbkLwPxYJU629vnZ7UmKz83aEvqb3f4ycofEcn+3guTQB
7c/0K4Oi1YQTckdQXwkqy6VVRyUE6zAEI0g9tV9ikQgfrLDpGynqInc6U+qNhqha24cXjufGSMdK
pRGduNSaiuvXHGFWJ/zDrFecrRY/IM1Thu0EnBIshYB7fFCAe4j09k4ui6zuA5MkndY83SXasPuR
jeF/060Ztnd13+bda2kkAD1cVEVd5acYVFTRggogk6FFb0+WBbcpqkinjCYjXx82Suv8KzUMD+Jh
u5AG9d1Odi2caqCOSJvoSoGMhK6CWzXteU6X+aTvTLo4mwd9y/4IHnnaMMlhYcroNjXEEOGE0npk
G53fsD4BDi6kDsd+UsPV3G1DwLoWZFZgglDjZRx035zAhEQdd68DWpDIoFJzerzo8YO+hhf1c7YJ
mtl0MPO/UPEza87IAGZcu48Siy+U7RjqKneR2d2uh+bf0e7OoFjQbjc6waIIgEoMYN2hzi5nBegN
2GWBciExWY5FSFMTHMw1ALf1cK/uj3XEM2en0IDQSe61tPCZacludYATaoCMGtqI1Q0HXjr8xVW+
Ea9RPaFZ5Ubxob7UAxTtca2+NhW0JOjB7l+ia40lsW2upSqFK7ndiJszsD2jqyx8ds2T3N4tr5gu
cT8erRbtb5Wv0PJDA6FLJh8s8Bezhl0luNSkXDXraFEXNOS7MaSJ9vLhzBVhV2MurCWX+RpaqHri
PKRaq9g+mcFUafSRt96kyMj4ScR+659jdHRriFh8lK9/R/cxJoy9RjNu6jAFh8FCF27QlR5FX0cO
MzwxBEYUypTSqC+iWMiBzPWZtDquDJI30rIpZXrTAFwvosmoUxlOJqkUqIb5ARApyyWQIWOVcfqc
KRdZkY8qcfv4YJPhP9gn/UabNxO20zYDR3ujztp2TT887kMUbbJmWXv6C1qpSexDx3magIn/5xwm
zeebaOnwROJFjggsPb/5mzNQzBJE/QQYtk4CFX9ea02ph7LPjoVfcfXNN748EkWugwEEuXD8uTcW
OmF8LGhU5BODkMob3lEGJedUt7Feuw7PBChdp+sYoIHZlIVKe1CUY/7Z7A/RtRGPSYNFoPJXfR7H
XkygTvp3+ZhwwoCAAtTRWnUR3aCpuV3uKZ5BxGYtYH+bi4WGmrgj87sKKdh3QAO04iUrLp3RUexl
9pUHWI1+u5NdTOjDzhJJM2dYfviSStS47CQjVc3ABFWfQ+2UL6sMRXKSK8awZxl2Fkd1HuFB2q/D
OCrbPFGNMRWmgiwMXEbD6fi19uMDbYG4mqO522gJtvUjUsLzM29QZ4ZtYJJRvLIvzK8qui6Lqgug
TG+668r51o+LTT6voFGvaqGGREziYOR1JcBJigIQDZimMsW/bDWqymVPuxs/CQn9JUxSflf4OhX5
3vz8P6XnA5sFeeW8R5jO77j1DabBBttYw6JL4aNCtrc9Sza8G8ueXKaPcT1/r9E4RegCkOC4nx+I
uejlZ+hDeZBmZkDRFslE5jyNdhzwgz9vp8Q6l7+D938DYjguXwYwO/bHyErbp/c3BHMCxGK45FNq
eKJYV24NmFw5f33hDvGJf+sX16YX7qWrqTh22hi8HkOBXf/iGy6rL0sabgnO54k3g3UZBsKc5E4W
Fg75wqNsmUFxcpE3XkhrCirjDYT2lcbYYC56yICfiIg5mKkFF8PtzW9VmosY68W96nvsbzDwqUHN
EBefA31osp+5l8/tn7zvJeZ/SphmSHuMXmWpzGkruEK3F1a3kXpAFuIjPg1Vyo3Q/N3iWykZLC3U
YbzwAC7Y0StjI09AI6Yj9eK8Jdce+g5ndqrSCQg1pBzv8yBZuK8Qp7kMjnjbTgPciWTsDFERoY3I
uJOf+tPo6TvguZANev3sFv7z0MXdV2YbUm6OOurcn8a/9FFki7fu0IoD9fIAYE7gZ8xMZO7ADL6V
NqM+J9d3v/Lx5yc6YnOG+e7QwAVc32vJA3YMzPXRO4CqGg+44NrjhFHbp3ocytxGj4EzZausT6wP
fl6K0r8v99oGZKfHD0AS7aw5IYMC0aVdEjNzHYsy+DH2gpnWe3TXWME4l70bRYNbpERFWzDfUR+0
JlyL36zfBbuu82ynv9Y5ffUq7kr369Jz5gOWe3Xh+7/vMrd2zoSv67WKQfsPY6H/EVCFkQtw0zpW
t1Vrr5t36SEnZDJZdZSYWUmHyUYqs7Pmdik+hyvCkIqZlY3rhRg6IZgW4EzVpYEEQBuMpRrQOKjs
whw7cJc+s5gcsy5odVu1N3e3m3fY7FGmMNBkq600bym7IHhn81860KzPZf2d3HtMkeV7c7fA3KT9
1dnd8VYbjQTtLos2rpI75pDZO3aIpcWOKUAEe+Vd3GSDlkv/NfmYEPA/fqjVo6VCGEv6iny4r1Df
dXjxytu72g50vCGNpkxuldWXDS9SHcaCE1zQfj97SvceJ3YX7fn/TfH7pEh1m4KXN0KnTQdMya4E
6V/vPc6bJ9NphdtipafbaRWGItqCez5qvGi0d5fl3ZEw0y6SFvX3ApR05be6CKftUvpwy5Oxs7HF
2EqZuWpXVMg4pXq7jH82OEMFhXvWfFiekOoHMy/8GoOo2Cmndyyq4qGWKHaMWfY5mbNuFfm+wCiB
afDPxnCLLn2eMsOaI4+ozC4Il+B9A6DYvYNpwPNfHKrqCrQMWk3od4MrEi9cnTe70hVXmOuLfe+p
RN59P8LPeF7O//pVv12VMdhg+panhUHfQM1BdsUQ5g8GY7IEG3/55xilmgqhYSJfP7MlRtVOrNcg
WlNJafP7KUwtHTQVQWYFuNTwCIeHvZ81uBdA9L4u/nhtqoUbEsrky99ZIyXEZLPHmZY8YEM2qLRT
HHxTLTDzBNMabvHzA/ynXbvW9Rwvh17wBD/G8aLDe7xFHzDkQd1S+WtTLfu0Iy2Dy8qc7tL3QSql
ZVZLRNy13riNxqrd7Q526ZnTNCHA4XE4nDlho1eLOU+8fLhTYGKDugp74RmVMOTt+8pMo2WjPGww
5ahmMcCYUiPON5/qwYYLu6emh3Lvl00Jli+V26tvH9fIXoyGuyKGx+2A+d08xXHdZe6tNe9b8N0z
uK/NuWQMvlrEjJg26UdfvVnxt2rSpZq86wUbC5pYsa5rT273OhCWvUPtiuWT+LhKvFn6H7bE0t6D
aKuOOxbtlvc6vBkxqqRX54P4n7FhVrmaaENyvkR0v1p/U+rZL7atPKasJ8AAtJe9nzy/iBO7CNnw
5VDh7jdi7YqenxprufAkdBdhyCAOXTJOGqaNPV8d46QVkzv1EYPRXFnb33rAOGZDrhIni0gEg0UG
muC2s1cc3Z7bEysZ0VNpbGEAAbVIBmOpjYdB0025XFBs28/Gdm0FIjSas2fYbY+ZXZpPz2Hl2CAS
8b8TxNMgNQUv377yKmUTrSMMMwmPEmZPi9XWPl5t/uoR/Di/b2kRT5emkZRxsHVzL9WL3yzyUGVY
GydNzmAIKEjs8Lqxe0z0qu/6zcHGQYSqmg0xni5D6WEk5l3P4vdlbNaDY/U+w+x1PvKOXOn4xsno
7rwx+O1tQ5o2MWk9Y/Ke6MAl77EJ6t7IdUhH5H8WwUG12Mzn1JIk4BYbY6rOIIgqJ2hvdflxaKVJ
82cGO5J65ciFMFj3yRmDJPpbwlvJ3v0If0Nt9Qm0RIw12V/Sf3K2T8LBoMYjHoa/nt5EeZz2eGDA
t9VNbllfpMF0wsk240HQmmytiRl9Z6Sfuol4nrVWNa4Ce0hWPhrLabeIttK8O/OYT5H+9xH1fL9l
OnA2lgNLTxM8SKIHFD6KIL/m4OcHCZchPD6kpacwkynt9wuwlwKZlUIPfa2WVoxbohstC6vxs2kx
9gxD4hMdn+Kdd5rGefZ0F8xGIeZRu2jjv/ikwVabQxuFKSZn9+p6CghXzlSgw6BnfMLzfsZvL/20
LuK7+2BqSBpe6mfiNjv75Ivo5a6l4VXjKpU3l53DEjrCToWbFCmlO94+Qo7TRITHCnViRK3SbGQG
wIw80jx9DbXtBWQWskTbQLKQTkmWJwpMsGxWK9E5sx1tHI96wnebFcZ/Wu80QYwUn3zmn/4GXiRJ
d+FeAqXsXT1yDLD7wzQLmsQyTm8GjgIqRhrtRYzU+cgNSqcCMtoyA2UnX1x+BKu6lQiH/E6uYDjk
RdNXQC+SD11pFAtUa6GljEmlEvNIRZbTouhk9KMYi7W/if7jqvq2dbA1yi80Sb1Zk7LXoeouvcNj
cwpv/DTlioTW2gYfwMccDFjpjkVkrvviNRPcjgV+JRIKDngN0n0se8Flr3Fpn0GfEH3RH+F+LS1Z
arAq6R+T4gZDYlVpchlbeB9ZY+ZjaG5Jsww2y8W9MNInI3Lr60jB2CO8vC+wawoROdHjlVp0urvn
lXfkQd18Z3eJtcwRUCAyvcwDNPqYFVX61C6Kluob6vhGMIL8ZT6VfFQuLzn746IP0leiLiQYz3PC
cZzGgwPo0m63TlDIQSQthOGH3maUpIwQbTOzqDL/ITLHUSl23jL3JEuyQknhZy66INSIZciWT6QS
V8gLujQgoXO4KRc5PfXG3eAofexcKKo98zhi8A5cvxH2zEkC464OZcUPmuW/FuHbNQTHPoJHtX6k
1LmmOoPSNTnF8YB6LiVk+kc3Tf0HvVD/gR7LQZdJQPoi3aOVeGrbLxF9tqy+QynFkpaT0pyK/48W
PjOme36RxhtrcT1h9PqvCJA0lkBw2gK+9SYY348hbAkVqCJWd0b13w8Epp2aX8psSI4xm6/oHRPn
jqE5XfXKyZxyGo/npn/oyXwsOReRAAyrNvG8h+rYjLsnQcj9Ja08GqaLhnjaeD8gSx3HabuadnJ4
b6+8jBC6GELOZcJbs4tbRQSdHt1PRCcse4wAJFFnUdFLBjt9snYB7vCsbTosve37xKYJar+X/CU2
dI+s65anTh1+/99TCnQMAlbL/yYBve9UyrCA49XJcsikpfs1IinrcA7AEcqDqpeYH5R1wyHVpHXg
Ap/wQQtCOICoMKbTJM4NidjuQYLqQbXe24DPq8WTV4mzogQ3nKqAkkcCxkO6rFefUpHcp+clsMsX
MZS7HaWzuH9alLSMYIY4lGSr6hZAHT5qFSgLF5pAc7J4fCZXrGILIx6R1Y7YJTftUgbem/Imgn5P
267AHBCdPWWtLCDRUJlWeZyV5qkqWpwW2wx4x2Oq/N5oHq4Q3tNq3TtxvjtxZy9Op4/NThlZMbc9
6/ysrNXw9zQIpmnQDySJ8S16hyvniSc11drCV+Vt1P6JV5bvJCxUz3OLrB27RM7fei+fT+i0Zquz
zEZcOll2HRMe4lut6dzdqQwKCdm4UlotXjwTKNbZvKLHjMF0MapBZOTthCbjIAcA7ZV9UXE2ZZbA
Z7+NxL4UuF32TKfeKthJFwkp9EETnKwlGJui52zzYKHYzwfApqgCEdnoJDfzS97Rilrk4dGtEzxa
3cN5DsoeliGwcjW/PuM95PJBqSgU2kVfN2MAWyB+XH9vf3fO3/QkBrpVDusPUK4MTB95o0TnR2LC
GWj0pcJYtleL6qxwY7Bof2hSvFmhsGcqe/6+mMOQiF5QKzKwN4xfIN/sN2oF+ECKkWbV7smIGHp4
Yrv1vKiQQkiBLWQpXcDLTH5cLW7jLoDhNdVTnIUOxAcRLKxDJboGqUMXXV8zA1t4G2s5v5TZN0E8
iSa/B4eEFr6LlUcb+NIE6Vz4Xn+p9iAhA4761htQJnibwxsTzbFOhv/T/PA5nWKfbb40xPI+DAUr
6WYiibeLHQsqABN70quIKpwPIpxD6O3B0C66mQiIm6VF6H+7BsAaNSHuxcZDmxKoe6TE5VJSkIS+
DTywA0vpP4fRcc1skZZLkW64m+dbI+r/gItd8NC5TW2WDike25PQaNIuRHUdjPeoz1KoqxSPAvgb
F+Kul4+TvXwj5/w0syHwdoUsDpBNBWYMaFjCMBlwwlNZKluMS8h+y5gmJPV9asdbn7+kSa7bpAsb
HYaC31GddJ7FdROcGPqbqXyB2Jom+RdFJ62d8QKXTHTGgQlNZC1qg+IprMF+P6nMonbV+eDsBNux
FEzL285FwgLUakGx/OMAJu4b08lIThdAaI05MlzD6+SDmqydM0GBWHVtLk2096QehHBlgkF0dUE3
/9XsgIPFYRQXJJEHHBxO08F3pEm5lJpIwz/skmbNpoW/3d77BvuD0UyIxo39CBVkC+mF8eIadJ/f
jVG+F+aGXaM4mkC2sg/QzFebHlZ3LJfsg3DDcZwkhG5H7YCe2a4XT511NnLYabjy63/kux1ua1BO
9ek0wOlTC8jHecvt0cxmLDVvn7YBUeFDzhhBNbbV7gVKASVyIqgZ/sO6mwMxkpFZq9zqzmOZETdc
Qa1WtvTpvsypLDkan3YL6iYg8Zr4Dk4lvN7spz5TM0OztDmlTrGW7pdPUdNfnKddvQv6+cEdFy8X
uwVzQUcnPjGAljmamr5GmqlP/yRG0Jw2RE7AY6jRj5wWOWasidjaNxBUL6443hqL8s62doGonOlh
3+tUU24tXrhXJnmmSYbhqaa/d6T5Tp8dXsgURSzm7rDH0tcYIh6KaO0aaGqxVnDGCR93xzx0f9zP
ib2W5Y2HtfXmlHlS9cdlaDU8RA9CgVJCWjE/beSPsHMFLgKMxrTjhe4viqPywdXkG+YWJCz6aduV
Hs6tvHbm/PLsg8hGpfDKqE7jpNT8Yu1fK9Sv5KfIlcbTfpPM03OCEhkWo1dGZI7356rXNPAXwDkG
nj3ZD8H/Irh5Y+Q2IwXC4VfMNtgqrYeyXdrqZl7kdcfWorMI8EJ/1R8sXlVEZn36ZQwr4JhNRRHo
QwLs+DgVDicVf+eEy9sfS1Xof9qYKWX9oBNVRflUhlnrObNQjXYkKB6O45j1N3OOXqwYrK31DehK
ebkD0gZkQBVXmSE1sGiLnkto7J7FpyBWrkEmA3xx7mfBmTGZyZngYPThWN5AQlG8AlffgV0J8/X1
X7SiJe5kPGjjV9YV5N4PZEiJLfFJ0oEMx+W2oiOQe6Cz8xFQMdYnWRraOiSRLY8qs9qsIfVGq4kt
7RTesn7qf/H9I2+E2HNdqSMMAipqdl60Uvpv3ck35j39AfQ0zR0OJkyowizoEwXFvILaKvGEQhET
+0e4XXbgW729+Onujy85auWJ0dDB18i8Ppp8MoIqHNvJAUu+RTmwHEvi4sMulYzJk/d9uGocIOx8
IOteIF6zrubcRHhPslZ1EsJb14wVYMhJx1PehsiKOCUTfnV0hMiRyZP9pJgb9NTuMyigG4H3lbgl
OHKN9vbeNwleSg8GmuD3ery65OzY+59qwAamVZvEJ4mvoH3MMQBp9Oia6qKQr+Wuxw9MQ1zCrpjd
Q9aSdSbeLZhQeewam5ZFO/UMBwEWveer7FaI/jp8ldcR26MXYo0hTYPGBbk0S+iKSwoOb+Auk0r9
GDGahaNtBFx1A9rWbfuIPV/JH5igN3z3CleC6COeAfV3Ghjmrbf5koqWpsOHEb5EX5/c/tTsl2qD
LLTew7y1irguDeScx6lzvxab2h+o0K4Dd+iaUU+zyBg+zRphWA3g9S+n6S2gwhGLc7r7Y2kignYV
5LieU/MQfiKzZaV05vP9SLDQn/E3H6nTs8+BQpqjL1Wu6ypeNM1d97dHbav/UMoYN78e9ZsVWHSK
U4VjUjmE5J4DcWAv29S/A335YZHpfu46UU0CIalKgTVJ0dpiIExjO1Tt7d7NoXNsxMPzMhx95Ut2
YiVdJ3UJi35GVaJ7qbAAUKa7e5CrhRPY1UzQk7Oa01sMh3Hyr/7lVD9dUNy90nzjOl5tUw+A5hHx
Crj3l4hhtsJJcOi/atda1x0vYEwgJz2Hu3i1hEbk2Rv1kGJ2a+frX6trAeww9fPHOsVQksLqmrtl
j5+NPOiUgUOQ6R45htYj+qHsR3y1eFuBdLK5307619kU23NVEmGQZVqrfPdQCdD/kWj8eZOrZnTC
mwjjU0Ej/mOIPWCxWucKqpoyaA1YCAvFK2EK9o+dO1sCav/XX3t1ezFvKFDIqXg9WJ28I2Sf9Ah2
pHJpTywaBR2im4hXDUKbmihcyQsITRtnzAaOjo5N+bBo3Trn7ReUTW1XBpudvtAN1NHMvjD0QTsD
GgPjEL6z2wVDC0KbwbAh4xlTbghsyluKhRNZ0/GjpMbdv6RiwMAVyLXtQWIP8RaoQXkNSZQdOYjh
hN4hzLokZhVY+xVlV1IV/bOjiWle+isvzafSruBTx6GXYuXw50ilgVWfBDc/SpqLfn8OYut+uc5b
He2FZXBJ+Q5y73O8yw6VQUJWpdse9h8qATQoo3A7G+/hwpni+II9mXjy345m1oD8dLqFsk2EMu0N
5S9Im+EExyL4jEqSLWSmPZZl/gdKHf2FIA4S/trcH8BLKRj1SfCuRGJW2/TCYAOK27oDpOukGrfs
kaTTnshryk/nLGgj5759ul9Jd03zMhrOKMYrbBAsvjqELBB0NTLUw/BsJXCxqT3y0kO5yBF+EpuA
U4OdCoPkKvf4rklZQ16CjrwD9rh0YIiy+1CEz3nYY0DKM7vWsHcxnHbDM8gOdeKIRnIhaKnaOEIE
toLCdkvKfpcVzNLIPXFc/RpBP8uTN3GVbN1S3PvVtNxYm+wu6aX0+vc56U99eOGwUKhFVg2xMlbI
9ozZJUh56EHipY69dABxpSqgiJMiFYEwPyh6q8RR2VPr/bZmGfs4nJMJVR+gsqLYW1l5wMmGeCO0
z/07wLSnw2WW6DHQaHAs95rGMyMni4cj1UPeGtcwUXUo57ATm2GCumCmTk6DCVKtP585lSC4kgVd
Q4JESLiGbti3j+YMqKNjRVSUiOx5cSfCxdMdqZdNZv6wVNE96R81ORZgw9zVqf6mIYBq+tQ8aDWP
4duihyT2ZEj3fxVo8OK5uJCuGeo81jGP07bQ+9w3cKVvzhgjO59HHE2ua78pMGhdWSDP1WmwNBST
W4t12bJARxDVVrcrKXOtNxYJ2l44jrT8yN0JYIjjXu1w9B6TuNaTa8gE/3nmib5HXfYuMFSVm8fY
Mgm8fGBCo+xOl1DGejcVTi4b3DDIEHhmUaWhGP8GDU4X5Op66y0AVg3A+0d27RGULq+orYh1XLzk
PxZPK0EY7ccwFUWJpbctpat7GWXO79BLhzP7/7nFj0aEQwT0OjZUt1B+uUuLtJUyGagye6uwPVIu
T3QQwSysf+Ftz7ly7CFd2K34GKCqBDJspXE+EQehwniQ4wa2DIgHMQyGPVaXJy/+JsNh+rAC5JZP
8eBsinPeuhr9IAcuD6lq2YmaRClny+JQL1EMi4uSseh3c/LEh8GcVi37lKWW3o5Nq0hTZteDtB+P
TyK4MJeGBhM2z+4XA5aJZv1CU2i8RmbC/6mKOCw1nkXf6OikaLuVCArBf2iQnsDyLJF0S1yo9dPw
68uWqHwBcxyDi3BJpGgNK6rarZwW2oterR3CVi/aGmFaSU9SYzOLE5eICdsdh/+OC68xF/ccPpCh
SMEWahMPlBlyJVAMYA9csJHvIWusqBJ2tlbYM3Y+fyJAriiTos5zl7P+ibkQNdewhAtTjEHPndBK
1hePw0EBYNJ70hS3V1BUAA8XZYFE8CGT1alPTjErlIklHIUXNpnCvqPfLvh4nVUorjH06s5ewdrE
Yc/H9agNrWQ66m8p9tn32rDfywI+R7pQqc7AC8bBNx7Exab106cAnqCH/2drW8RXykW+91Dd3+eC
3SQ7VtMJjhs96D4cfq+iyyROChM739S0oZKrvAJZzumLuGN/OtDfIqX6ZDdjoLvMoYx7ElcRkXme
8v73+D+ZcRVaEomRUMXdWUE/Fb5lbN8Vw2JDnLE2xvrWEqqrmS5qMCbO0JWsIeTwZxCj1RrvvBvM
QM9PP8QYGygVMyuHgQKPJQA+D/3yV5Jtu+pOH1uW7vC1l5pn3+0uqjvgvq86b0//hEoKhwNhFUCJ
no37N94+a54kK26c3aEifd1U5oYcfHng3pGFgNfF+CgkhAaEdCopbyLCMvUnb4WSbjcxi2D6Cj3E
+zOz3Rvu+tGi4vEgrGl3zPC0J+D8tzFTZr175zL+m2xKbWXIR40VDF5I1Z+Mb96Wyjgh/s77dMr3
VfGZcRjSe0hgW4rxi7dIOx4orb//kPsKbAvynrewfhHk0+XXuqMwD+FS2K7/AERFRXdLoub74djg
I5vSRrVWih2FPUngLAHaO1Gha+sJb/Kp6UK/mH52ZqZ1bUda1x2bWYRZWXHRLDQQ6aAIv75FAvaY
cqN1S0YXM/04IAmMkysNvvEeojCdzaAsC1sdJPzgJ9jEWRsEabkGAcuGCl/UZ3VNpLrBaG+dn7mS
1HSO0UQPT7yRPk6rLLrd4M9+KAfLU/jVmHxs0lqDnzbFksskyk1zRmln/Ue7rQPtFDcbkwr4oweB
K+PTyxPCxPxc3Z3ZYd+/R1lICaLlbUVUSS1fmcXp9B+hD4YEHIiyUc19pkuuJtPwA+Mj3e0flk8g
qn+Juq5stzqV97g34sV4sKD4U4D1qgw5wB1PEBAhP75UqgrI106qvxd7ZkCJuDGhcRC5HSUbyQuG
TbeP9EXBiyRLeWT5fWvgNrxjVK/OFE2w6+eqLBhjGSPls2lmyv2nor6HV4Zklq9IA8oSPX2gMrnK
J6IGQP9lc9pYJr21liODARbbMdAgRS05LncT/NbLFNPai1bxdKsOHmLwaYPbizLfRBSahu1dDhYe
mBVfSKR/L4S5I2G3jBMRpvBhuI+zXtvaR+1txRV5HIKuQCt1QeoG2RmORCQevq46KG0MwKIqAis8
nqJBcyftDXH4ILeeQiSLTwxR+H5zLDUflgHm1gB5n2PuRimetvTeHAfmcD3PXy4YiIfCcaTQal3q
IAeQe6iYtjn66DgoEXFQNmGjwdV8rUqcLWUHmezdCTqWmS9uXqDN0LD6XVQT+lftVwRlGonyrZwg
iqOlm7d340ItBcEFG7A9Tbxii6bbWXrRZQqIdf6TNV5UYHdrCKQ+f7HzYmi8XXA+KeqiPpsvNFGy
gOTgpnnmYF2Pa/QGoYhM5j0zP8SZzODMbHYyhO4Tyyw5R5txVrro7BMq/zN+I7c4it/1uq3rbTzK
UH7q8PpzH5g379oDGcvYfSNDUw6wAU0eoQ1JhTFLSQFdvAdKLgp3imJqictdSKiZ5rp+lPSpdfn4
+eRgav0M6xhxNr7Ky4Y/B1rKKbw/4qPdvnpU853uE+Lemp/fosnIW5NJmlEN5VsZ2Eg0zZpyWC8j
FHpp0l963A43L8Gwbxudsf5FgrPAeJIIsn6sS+y/DrZcb2ILIVfgrWmj1w6hCpqFV8jcDlU28QAE
Y7p2+G439Rcjcc3fq+SANInU76L+WL/Lj/Y/7cdwIFP8D6uxu+Ws7yZXScKDel5UwtGIuGi3Z4WB
nTdWE55e1rMDhsWosJWj8E3DN0xoqFTJ/vF2UsF5c3sAFPwDz0BYfyKJ1VvfsW4ArlvL9OSGLWsS
lEKtmm18opnLKx8eVZ8ippBnT59ge5MvBog+4+Zk3MzhSgg3MM2B72fOPttRxrQAxT/6f/jgeKfv
OfiX1DtxjWMP8VOzoI+e3R+czZJYwnt6XIfyNAErzsZ05FGhkme2e00XT6n7y1X5lMRSlbosgHJe
9F68mq86nIJvcJ2x3i83xwzePu701dRn+IHBHebrfkYM8pfHSzGcsT0rOoerdl8lQLCAfy/qQ/w8
iojaCFbt1zvQe4QwIC9SdmZruczzJdyfsCNOhCi5Kx+jeB19tYDmPcEnYWPPdYeBS5dewaFuvnRs
rbcOeMoZFySrycev+xODbwQsKZ+ekQ3UJnpN0sOKdtAMVOvlhgOZQuz92lnwCEQHOEuvJO/Eysls
wQBI3MbgSXK1ie9rZpSbIUUGXiBpzvDywGvuQdEntZCoGeB95A82wzqD/cwEq3q+Ll++IGKiSond
KXeYt846XxTG1/0cGAXpyNeWr0Sk7Cj3XVqxCpF9lOuVEmHRoMr7H7g/Xaqk2UfE35Unw7QRT4gy
pIJtI8kbTa7THf4n1GDnFiUONlHLn8H6jpOw7AKlecGhYURMmP0VcMHqPt7Sj0GxJCYVV/oaAgHW
kwZe36JldpQgzSvnu6ZxhPVZoLHKm7WnEJBuQGl1/ztzXMnmyrlB6dZVIpWyrVocmmBe4NNJrXVi
VJcCkGBMHuOnl9oAkSdni9zElePLc4H9OqZQ6Q7Up4zDg6h4J1NYcUWUPM3d+Djhb2ZVtj/G1hUc
KZFKU+F80whWrpefDTF78sPfr9ScErO4b9vHuiR64ixi/anLL5itVY29zqzbOXZ+nhEQ8UWyRDBd
Di8CP1gIbVSHnnPiWeKSPPU6bEdoqQma7LwaBAIyzDAtCZO3RIpcF74VQ6I1INL3Fd+JrXX33mGa
qJknePW0NkCh4CORRsLY8WZldJGdDxZGNipDArxs19IGw6SG5lkzKeZSbeiyfPVcpzlv/D22ECvu
AIQ4e7jmQv9DJgpCBEp053cAiis1ximfT5EY71SPCaGw0sQTyFXwDwfCm1O3aKr6rmhwt0Lw5QFU
cNmmhUV0sXDYrgkKeCHpj8bZI8aywUwp5a7z5A+6LS/X2dcDDhbr7+cjrET6v0avLKtNzI9wBw8T
aQImsFbrKUi5FRNKbsP3YlYxhJZqHv8bRF4iF8jucCKVNl/Z9XsSMVn9nGNrUssf5/1yjJqMibWf
kdBaTmKbWB/amqzmtybNU/bD3BmhtjVxRYz8McFvjr/efp0bj+yjA4sWgbA63BxFBAez7F/RpOlC
SmgS9moo6OuqORCa4upneAyh2zK+MvTIn1sf1ZKOtR79LYswtIz7od9ePWc6zofgigToMv8/bWsS
Z2iD1A85ZTkE+msgKA5+feuwkBpGuT5ehxQ1/kOIzNKr/pzGeJabaEbdmuCru8W8UinAi4HkuFqd
2CFjGguIqX+RHd5Z9SiDwRPya6ujHx3NVIqn1zelwGOLVKGJh3Hi8e4OPeZfNX2wPVwfNwDsSPJY
N5B5jPq/dJO1mExL2v4RiIWCFeHkk4OgSq7ifYIcm6yYVlywdnjFFiI2MN92mTFOvphZQwYzQfe6
jYX8la8rPP2PZQ0BwpAssB5LEkPSyfTS+7RMRk2D2R4o9a/P85s01OqW/L5tNfmg8L23GtWeHarW
jUI5N27aFZcw1XRdz0XOa64WR1pfFhJU3ipe6UZztau8d9iGRyp7baR45TTwxvinCrBsjU/n+62K
yOAumiOunmJCEYhILe0f1OzUuxodsLE+U7P4rxkwvfE7qSsz8kJWorcY0oUp0VAkG/34tubxvup0
JRBK0SsxxRCBSNfABN81DVl0mt+NKYr4RlHjbXw7D1QkpfPRPz1BlvzWSWD7fCHjfVwJbz+4XymF
T4Gsb8iY/fGWzHwvweqDjOsY475cuC9LGjDELGGsejMxueEkpMJRm5om0yQKCI21Mu+HF3y/aVdq
mvE+5lRbbCbszVa56SaxKRYg6SxnGy4DhxbJVByq8mbd9QxSbVFgFsWKxC0Wo5/mZlNMHuH11FU4
DWqV+eu1/bZT9+GR9IXvQ1edRvqn+c7Qg250iUwQWe/6mNQfXKwg46BnRsmhvYgxwuPaZ73xvZ7S
znTa2SOlXvq2MAACGODFJTh7+0fv7c/Xpdobxtz79+KgxPl26Le3sbJG/9zNR6vuKz8+oX/KShM6
4iDaKYvZIiXshFH+M7kjyIFzS0ViU2kQMjqe56bke/+KyIQ2Pc+JFAEc3zzMvJjfAQlQByc06Csn
Y6OV6JJhn1vP8I8pe1qBMVSHfMqqjWItoU0fdYupBn1bbmhzR/eFXO/corVrENTUbA/Mg1qS0vOj
ds+Jhuw7jyEDF7SModu/pjoK4PcbjbB5uun8zX3nXmbYAahA9zpHLtgL386OUsg6dWWceZyfIP6C
VIADfhW8cwyB1yl9r9FySNiH0tOejpCkJ8SnldkXRR96LHyGRDAtx2Qjo8fNATulGfBlt1XKBh+y
03OYPDxUTkuaLwXVKJfbgs6fhSMUxRz4eGz3b/MzB2FN69dSVQx/EuMrhX2z1U7ylrTAgoCgmqYw
1+K5DBcW3GtKo1FoLRj/B9uUjsI3Eu9ojsBZQGUcvW/xdkI8MihGkOyA3GJaGEmINNwd5k3R+GfR
7ME5eR3yCgot6eZabkgyeRAyGFs8ucQeMtCy2fiM5slDHJt/iZwQGPCi+HbUySeg3LdvR0Hh9u/W
5JcSGV/sKokrRLAy7azUv4z88apxXXTOtKvvYhSoffX+ZWISvcVksufKU1DTiMKXFRTT4UeDrcfz
COkq5dNGHYB+biVBeyOY+Jr4V7rWtabnHg83aN7wZ111IHIFzvn0JV9QhfujOetM0CegqlpoPqc2
K5Qrd/MtO/D4IMD6M1l44B3IVBZC2xZ6dmEjfu08IstUEzCNudFvNPhHfgCO/B7vcoNAVtSDjJbP
QTip7fO13d0/nm4SEla93+dunwHRDdt6iwEKPw/hxgJUvv7BQ+nVC+hoJZtcd3s8IM/WhL5ELORU
3CgrFMPHdTkDzF5aB5hY/mlKUobrOuqvl8M7LmoJiry64i9hgHBwfAZpFYyZlY46aT5TfJoY/buj
sD5YouOrO3MdDcOIRWeuUg49AnFse8Om9ahR2ilvBKqoduQltPCuVdGY6/ebumAgrm64aCkSsZw0
x14Da7LofxH8QI5cYzRkt6BwXQX8uFZuMPe73qaIO7IFVp1fM2aL+xtHy9lnim8um232WhcHe6Ff
jVLAuRN928XK8dQkVCbvJWEFFd0mxkvGPfpKU17BaDxDFOJswyZSGbcNUwWw2JwcRo0jeRH3B9Yc
CINyl6icxN19gTlcMJxV1VzanpRmaQ0A2dvuvdTechmrLau6D/sYuTWbZrTFvCxgp3TbjebS5DEu
k8ENauIx8kzC3M9dYreIi7TfEFQxqHx/FvmLLZzks8zouxKqUiDcM/ZizQoYLPh0EQ3i2DmojiKL
xpa/2qQO6GhoMXMfI7sGCVoqTPkOSAj/GDeRp4wawDK+884Eba3j96g2rq33Xiz+tv8+QQm8zEOZ
ti0CFXfeYHC+CIBh8pY6U6+S5WPGr/WJLYkOcf3KeRo+8ntPAmhv29XaZ1McTiEK14AMxZ4jrKr7
z6RKzcfKJxQ4KEeB3VQnrpPXxjAv3+il9JAzVGesbug2OEzFEpfvZVT5NPJchlUGMN9NWXoSgXiN
DEYUGEWGy9roe2uSJAxno/4SLv+8zO5v/O0saNvg8DWpiDQpjV3l/G3n2q4+1iE0pfuwjteXmsGQ
uPZGxMo0ledjw3TL91glEWXKhOYA7IbtivkjRtl/w7dPZN9DHfs5w3JxZG6guMX8MscKQUsLfEeD
wAVWx0yHanZzFGraYVqRpCgp7pqo8G2MBcg9m/ZqzGJNyuH9qEzKa4mFnaze6m/wsNTjbwmpDryg
1FUJP1roJ42kPImFX9byIEDP/l5KBMSoug8Z8fY6pVntvHXaBsUfXp5JOlokYOA+HIUiPeCBiOqb
D1e8jHvt5q1Qmfwl1gKj8yPHUrIfydK0O6xso6ri0H60O2i51g4awv5/H5rDG/OlausitV5kklI8
RkdGtnQlI4Bg+SxLcy6Sz9kMz03Cd+JXOBOZijimbN4Ez0qfvB6qvpwClNrsbvWK5mjXJjWqvCoz
NOL33sI7MjFQvQfHHM3e9wernecEVfnNariBCoUTnn8BWQkuS+JxwFwzAMUZM3pcPt4S1UItx99l
qkeDu0wfnBzx1lAdg4RWWJxRa/T9alf/ZlOfu9yde4qXGTFI5tTFJfq/ONfdC/towNWGkiwAdC1m
HSkzMKFkh7BPXA8ykxQtxMgL26Ivzbw9pu/ukHxpDKKRzbgb5l9yEKE1UzZurHjYbdGe2RVfb1+8
KBFFgE8z1RISMQ4hX3PNkRwlHlxFTSVeJgXurSzfpjr0KMxHNyHG0y21VcFw2dsIO7RPqjDNQ0+6
UQpHDdqrpiPAu+wEuONbgWPnECUt+2reAPB2eQI8ax6yMI0Yp47H5Rnquag9XZCLKI+p/tKRyNUO
SaJ0xXTF3bBnFBq+KoFi+AJCf1+CfLJ4lnP+8sGIzSfkC/jDpSTVwO6v4exy4wmRT93vB3GCbRDg
ZJwzi4llgNpXdBlkwVN1IKyEbc7ghXMhJ4f5M4QDzZSadXBu8ePSwk6smud07Jj5GWh0oSpEzTSH
D/xswVUKqYW616+WIItFn4GMRqtzq5oG6IF93eGsFSZsroHb1jfffkaYznZsUC/OREaokuv+giMZ
tmBSJOl86OBhplbSAd7vdnMUU23XAwkeZybn7Qc578Fd9mtg6qUNhGiLyTdB9gvLw3Il6Uk/CwFK
4ZqK5AC6GOJFu6lX7h1ftw5ofQME4q0uXnw64uP5DVyqF6NhnWmeoUnFGy4q8nJwTcAN/1aG9uC6
PsC+90ml86SQi31Gl39jZ0rAeNOGuoBrbmx9R+sMcROqHbzi0lml88GbSLTFB8qoDsa2gQ1f6CNS
wJ0J1SztluAFok79Njb4BQrpDCiLIe8K9yLNFNCgc+mOZ30Hp0weFiq4keb0sAWJTzp73Tflb7W1
5LZ4ymDo/ny3Z88bvSECf9AafseIHdcHrqh36QVphFFYZ/DxBq8rj/zgsvWZu1tA1zylCtbBJdtB
Wb357CaL5z477a5bJCbU2NMpZak/dCZuePgB1qr3wg3uz2O4rqalF9DBuP9yzYSjm3KN8758yUAx
E5jfQkCAiyBVjlyuAV2qLHSA8Rp11J3zxTlJFgQ6JVQA301ipGDwXuNxm1EUKyDC3z32IK13oneC
B010zd0ac1BjEqZbJdP8xG39DYCobOILvBoPd0YD00MGBlxHmoUJQYIhLMUilR0Xzql4p05ZvNGK
MfxUA20Jo54qfNmvuBkOR8JhbdnQPMHZzjVBtOBke3irYiLi/er9FjjE91DgUK315bfRt/xzrr37
fmEgTj1DCzFLd85MFQTKXi+ow3RgNVJvZvg1lpm7HaLTSV8RJz6ZOsRr+GMXuCOFBMN+6L1NdQRP
A6bUu07EcJglYf4kSguH2EuZw9Fhb6vLrZxqzdEqbFX6iX3uYexAuIiBGsZKUYbLEcHYcCol4KFl
cmuUzwM/SeoFI6w+BZj9P0XW4uXU7gj7QJgZsC20cjaetY4NFbrapZ9ekI0zmuBfofwmil5txAiG
ucrsh0JClUEwjtazTf2LSQrdQ4+jzekcudnFx37RQoYnCf8uQan3h035aR4g1D8NXWeUHiDDwrok
4enD6EnUoRRglyuntZd3CXfLBVe00MNtvO8KoFj6tBpm0zf/sZXZ5nUyJ3pfvXJr3Ih4U8NlOdZT
PoBkcE92cLs32DuKz4tsJbr+wxAjw3lzFpjW7F2w8b0F/zAH1Se1GAchs10CnUOaEBZwavmXLo0k
EAjiXeN21wwjwOwcFK6wX5E7mud+t0lQSQfKA7Mxb/X9iiWABwvGQ/MBNd8/ICqQi+p+mh7RhAxn
HC8njXne/t58lZVsA94ghWJ9yTpHBX9nIiEJdn88L5eEbgTgAI6NwaVIXWuQDrI0cz9k64XSY7sY
o4D8hnLDixkwuz7zrVrfj7HspTs4Uz1NBUWS6tmLxmx2IQVazaxhN6n7dqkUNKJRs4x6HFF8eMQ2
WiR6ivUHjQHb3VtuaDyeM+TZI/SLXPdyzckMOBwmXdkx71ObuAMJo1P7grlcGT7oxORmYhQumR2a
r5pWliAunvt1TMgmZKF2dbCe5psHY5BsqUZHiRCNBDCIPc3hgq1qLKrvLeoDljj1andTgVSPxLds
hDxW7kscaydjtVEThmrY4De0a1+eW5zImsICMQedcyZ5qOB/aaV6Y0uc1v+1qLWsj0GuZfOMPq5g
3fNtj04RJvNVKzCR5bMgJ658FK5+VI1hdgQADp2pFddjtA/s7VjbXVenUYsS8XQ1uEEhsD60A3i/
2pf0VSXH9hzvq/NWzLnVVUYHpzFIoBZm5CXPw27chBjm+6Us8Ntr3WJnDtlz7VBS1Bj3znNWu57g
NfTnXdgA/c/8VOzmh/vZutuj3KgKyGE5h8F/sjoxXiTfvpqWE3mDyWwk98PSFt83MQ0yhjLT6cWa
EG7mbU8WD10Ri5iecBda0x4Jzo3ulrpGl3Id/NDdQ7LGsQ8Jg83qp9VRpojL4b5T/5LqsGnSX547
lvyVKQJ0NAmZhXr4rJUs9KDBg70OIJQGTfHod+DwRBdqrXzjtc1//gjPCr394QkXtmzRd+ZcWPIC
vZTTmxyJRevaaA3jUGRtqNK0QndRCngtyTmIGiD2WbCrZcfQiGUdzMTdkCSafF5y9e1ku2xmLkRa
pSqY7Q14ZbYr1lUQNxoTRfbE9fXa+QEIGiNWntd5yHW6HBWRJjZIYz5Lt74M+ZzUCjeDizbduTjf
38hgCpKBAFzowYAtugBoGZOUsbumqp8zHMAQRbR+8dy4jyFRUXDCMILyJyU8T+V6yTKZ97wzLWvr
QC76MQ5obyfLawUsmYmNxLA35sTaCTLk3Hm6W1TKQlcKHI5rqEd3E0LIXT5KzhB3RNfqPXvA3quU
z6kc9sw/5TDlJYgrYWI+4fK1j3NDEZayem1aKNFHuokB722Vw7R6+SyBBLBp+OJRMztBp0Ki+Rlc
4If06pOvNnNmCV4hdjN6mjtCOdgUrIo73gXKVh5pc6CRKpuGJ/MxXrRZTFrHsmX7TC8dpxfijT+s
XPsg6cmI4Vw3RI2Xs43mHto+mHPBVA7bn090VYNth/LxsvCh4p/TFxzNvAtWfMw2rRs0qQMr+42V
L9+NNL5Ux9GIHXdvXdwxDM1qhcSYDhD4IoGXNrVWLUSkZ5omD+ek5PW4fvnbAJEPsEY6+5HCkK1z
/6D3h3Sv9IFeODshQ7+aF5onbQXkswNHTMDGJnxQJF2ZbcRtCzSsR21OzaGH//o1Zbppqy7zeEAq
NAXjsafj3hFxNvva2q62dW3ZS8FDHgTbafLHpRGQKrvT46q7mPVH7FJ2daQrn2PAbVbNFy/7Iay4
aVQr3e6+LYUpdltJEzdHvOd9U3nWBfjpaHSbtWFpczFliapYFvavquQ88aPnls0Me33HdjWzz/ME
EY61N+5FOzHFA+aP7RRgpMqXrpEIHjCkGggD91NujcFxPcBkGGSUn6KdiEbgixxs1TH2AE2fE5T+
O6Ok273QvE8J7K0QlFpRlPR1JouFu4UXZ2rJ0Y1aV2yEI8NgH62gNpnzpXhMlFeNfo6gtV7SjH+x
84McK1oMRcg1XKa6l4kQ36CVOm7+gQjhlX0foSkmrDdWZ0qSvvw/IJc8HB83HBdBKCX01Obnp9Kc
ddCLxG6gjGk92baSHYeCO3j/HpYyptxPHOZGPfX8ZWmuBzUHuxeMjR/xKSkQ4iJg4BxIsShL+PfZ
8M1KiuljectHCYTZ3m4yE4LG64f467SxRSrx81DLXvzf586u0Y9JQkrZX8VQ8/yW518mfwwl/n1J
+ORXUYDb+SRrhPgMcLD9I6r4hqHVOw7oBVqNrlHwQiBZD0x/bWNYYJTYb8OeuzF8dHAJXjSHaJ38
6G0EeCZmfvkSl8gOOAPzj27td5/zCgbi/RHwn+rlt3LV7hEQ5uQxL98HTLLfO7JZM3b7FRhm6yCS
USGKvLakkSgrpUF2c8BpU7V9HVqNTQXs2+8NjNgXPcOnUkppvK2LKwwNbbxeZE4FBv9QFbXn9jHg
kwUblXg3oXlTm54YivUoSOqUqlD6XTqYkg98Gt9ry2FbM9zSon6/+n7ZfjgZv8szmemMFxAoIg0z
3ggvv2pOadtVW14owF1uyfHi2RNBigEfbBJZpVqDuOjctVsYMdDSOoFSKvgdRME4npKcu4KKeURG
TUTIvEQlXCwBOTSzLjDdinRqODiRA1Drj7ab352seo9KRuDHWAgfFnm0ojXjfBLXgEIOREfJGxZw
VfpaIWzEL9+dxZCS0WWDzzZx507oBhyuN2g7I4uhUc7ATcdBkIJgnFt0NgWEwSiaIT/lE+uhSMAh
bM5B3gPxhb7+fLuyvXPxdbdCa643Nr51eJ+NZZ+lCALtsvi5HwwngRxWK9PDzjv7y8rgEx1LZHsJ
8BQf0lb58Omq5YsBuNESdSZ+lwsd79i9ZyQm+sO+5F+IjmDm/J2Is4Zsu3dJgnpeLm7RChSg/D4w
vLKLZt52sw83SoPPxYrTJhgzciQuoMqBCOnpGCB04lEfojJF/4d4EzOd28LJTFJ/NBsHnvTCY1h0
e76jXcn+aODZtzTMMR7dBtwIkJazRg+SaVW6YomPYB3PP2oC34wn1nU+lZMtpGdNHwfSudpkP8YJ
m3vZC/WfEe2w0xhwEohTUt/FoO0KR9xDcQ5tQnWXM9VOCkXOvNMXLYqPAyJhSKbtG1tOD7rqo62Z
6MVb3FqTTLF3NfqwWeixjc+bNL6ifu/6fAUdohm1P7zKz92Z5S0LlUthsmPALLB5H6EbjcFg1/bg
VcM1QV3jO5CPLx/QAFtXnJPPTbqst4Rm7FRYhLivkWN1Uhv3DupkcnSJRz24c9O8uJjfwCjSei9R
wlD3ithge/eSpDBzoFXrkrjV/jeURNlx94E6B9pm/hNXgQyiS8CdFCwVouGDrvdIqSMWSvZOdyIg
e5Kx0G/LSvkhXl55ao3YuGu6UaH9PYsolOeCsc7RX7eBu4it5D0HuqK6Vn8rTqX4s/cGFoXav6nM
ZmylFBcwNZQl5mEwBG2sT/7udxxEGFNqLYrqwbDWq3Yd64FYYTMye17EWuWGzdt9o0OmeWOFru8N
my5WHhiw0CAIAovoq5JpQ/4CLxxDCYenqgbnYXdKQYVhEbGZpBZyxeAYIvrb9ZiWNbZqszIcCF2F
atw0B0On2kR2ftX6l6cgxNK3F0D9NmLOdXdnIfmvD3ZiMJlES7xiRU1zCwjt9QbCANQV47s+cOMz
fQKwfIxmvmIwy9lGPJvJLTGgjVv9iVR8TO4xNwdkxgZ0ayycXT1ufR6c91/MshdoTadJRz6j457K
LOEKSI/eJcnjmfN0ulvOpdduS6LQ7m4CB5VBGIajNiuwdqelJ/L6D+9CKgKCQzh5BJsmMbx4sdCw
i2Xa940hUjJdGvIgaMEAB3+Sg5PzNWxO+Jz+Rv+Nxy5rD5B6EoXoP/RsrlAueYT1KCo7TFoOhXH+
UYvXbB0M6oJiv27SiTsyUEGI/gwpmTKDampWSM3Zv76RZ265W/89GKgsKWLYA/H4Z6hTvIxIcQZ1
LQVqqQ8zNbtNZrXY7krFJqwAv9aM3mPQJ7rRFvND8eFJ5goUl/ceij0PuMLcsiHDpnPqq9Ja9jNp
SC1i20WD2UAm+vEgCCDAVAuUYqJf0a6IjVhb3SEfcoZnR+3IzLeSC7s/tN92rhY+TT86j4wX4JQz
/Pj3eW9TmLkoUQUo+UQBQDX2orL9utDKZdhi6fo11eTg5huvtkFY6UmoEHEp3qa6SGhc0uRlWWCO
5Hl5chbJmOxJ2Thq0CMyGYR5871mCLz+6ciVJCTW8FScw64oL3eo8OunZfESxiPj/OBfRuedGBg8
n+zrrX7GkFerFK/3bW0mEZxpQ0YzgvZX+YtG+GBGQnVBNc4Nz/2bI86VXuFtKULS7F8KfvD1XRaO
YxCKiJz+l+/4H9GBU1y76QnPIA51MCSy5BGnpWeBqpX2aI9/3I66I3v8Kufv8y0OoPXNqOQxBQTY
Ru0aODjMOG3O5sqhZCpcyc7UB3lzs9pTeIxDAelztY8Eo/nx+Bv5CIvZTjKLVADGwtf7SCTzPWMr
W8dNiQ3JFbAncUjjeMY0zZmM5m9z8AeSkTpht3CM6Z/OYzFbn20XDndK4ffUDx2N5Av3T7Px1cpi
+2aPnCApy34S5yKbfaqf7Pv4TSAbEVtbfw5ZpxSnQKlseCkI+5hgpejEE5Zr9/om6+3dpFwUSjpq
k1c0/zGrG1TtXu1CsbeYmVyVAcD4SU/XakVOTOxsGT0t+N2fy1yi0VJwIJwkGzc4whUcPXZUUYAT
ZuSZ1tZ3oanvcEBt8EIe2LlCmdZ81dOmukGxhsPOSSIy3dgxaJxfbttf9tTlDdedFzkLRonCnA+B
YfX4dt254Mk9G9rGTjJKiv9khumrS3cDdrEUTmthoDXdjSUbyim68qbOqD5OpnEDFOzIcIIAElvY
UljOosUXtyaWTQoB/3Jo3tDdSpx7Cr+xG5KFkdPOXao9V5BQjdlXhAhQ6Z6WTy2yuZrSO//l5D5t
DAfDg86SvxNweFkJHFPKdxLM6SxVnneLmzYii2UnFNFMhGTBHpsHYM+/L7K5wvd5FRU6f8k/vdIb
VX0Hu4rKz8Wqpk9Gu8uTKkiMvUmmR/KPmM8taq7oKisEmq5gWuBhC+2SYyZPDtnNfvjYUu380pK5
bL5HwJ0fjUdaNUA1cHe675Z3FCwEmHSlDMfcOpv+VsOBpaF7GMfCrfWg/f1a//tgPVAnR0ekTcNu
5jsduUBXcvFI+TaxM6tvj2Co3nWLtL1r70TOXy06q53E347t/Ty1T7YL8J0Lk4d6YWd5OjEFn3j+
76fB0scfoxK2iAwJaDxqEx5TVZn+I+30xjpxytYPoUPdz4nGE5TjnyD1xS62277sNaEAfjAyrtLr
gKSQumVFSGhCew2i7qT6fmAq3K/z4kgqB9xrPd8Sj9ZdAWX1CaMhbfdC/un/8R1JYKmpl+gaaPeP
/BCoujJxyX4Tfkx+9ribqVoSJ6C82X44LVV0qx//UA3FqPntRcqgVwBiq/kSzj896kIS3ff2ecpz
AQyyo6Y3hRvRsOjIEJVk6zQnujN4P+m6bHtWiGGv3ICnTXLw5QwHE732zq1rSO3K8tFlnGyH6jmh
qAyxKsKImYFdOzy2tCeUM0BlxAynDu9wytb5o3nrro3nm2r/HHlj0zUGyH267NWuEUuaMMKE9tJM
KL9zRq/P87cDKyUIMpmZz9llh1+J23SylRfZxYdDvyz/htRW9SLtSf8Syxw3INOIOkAx+5UG6ubB
BX1wTH8cZZi6hH/aFmmYnpDSViXay0dcPwoBjUATrr2EMvvd2oElxY3ZesRI42UMrC6bTSOHBV5l
oBM+O6IdUVvXZpjR0jUWpFirnFEihTHp6DHVEs9pVF/QZyiMYq3aKdUOtJpQToyunsILLlXPF5di
P530DXpVTv2xlzQp7uqfS44szcwygIR5FYnq3rMRZlKwPixtxHhDCq68S071i0u6GsV24+uyKO3D
gB3JUtyrMNVJwMg5zdnxPgWn6u6QSVPhfmFBkhcJvAddiqHg6+KUfkZsFrTHNf9MsBKIbbaON8bh
dBNkxg+qakXlZ2kueknlmLaF6VDf/vHklj6/yraHFDyVnZSj+VRiZsDgNKYGbCeGIoKd0TkJYJeA
cBtBFx25WEBdtkjF9l3a3klPKFFTMHL1fkyAbZFevbOOLC02Khvp81unYo2Kp9Kvm3A3OVFWaGfK
1xiPxah5HABUowkoJDx+GIlwMzO/fQaQjym6LltNCwKnmvSX3U7L7ixYhRKX5HmMnOVjPQOm5pES
Tzr8rI4SxhpzISLaLEotqEZwTzJNJ9sr8XmdiGiEEkopF2rqwwgLhSSQ7pFOjQxTjsf/+BDsdjMI
1tJk1T/XgtbT8At1qupP8c4nuFk7VvjmvRysKC98HKTH8NpIH7u3UIxkiBMFL6JAqNtVdOAUcu5O
Uv74o9XpOXddMWaF82GPJ3hgMKD+6bU2kketiDj20QbSRrtU5MSShuSATURkK95zjr47I8G+PB4W
g5XD2skktsbs/svjcZTgXE4fNYz21Qu6rvkS+J8PkI6ePXXJ5EQTK61zTXSfYp7WIDbaPYKHs3lJ
CJ0hg3Auvc59rHIk8ZkexX7zpgo8h+cCllmO4mNBzyf9wUui1h9Wzk912IlP2Wfw2FRHKTrufxef
FG1fK4EXiD4NKyk62867SjgFu2nvusQf7hAJe631x/HI9dk+e9NRB2CsqzzDCf5F221Y/IqI5TnT
IBDXWEklnT6kwFZoYpBu2+hVY2+dCfzFt0YRZr49U43vQPo8PAnLofuxlqgxqdqkEuZZbFph44xm
sJZ7JLEYdV8Eh4HNzogmgNh+TPCC3w4BklisDkPlWYfCygUZlBHcfjyRzZIe8odRy/HbOdhzwwDy
v97T3Hu8wz5ycabUjdxUa6Iycm6bT6hz7Ijta4iXv2OaeTWvNTVJIRf4CFY8/lgSppex8Uoxlzmj
wHP4klbatIdK/BXGTq+jOura4J8pUIAkHozrCRbxCMy3/eSQThTmFJjMcbYXD+q5AiCAkR427uhC
qbkBJS6p1iFSroGDHftCTfFPmfb9mmI527h/XjT+GdZgwqP/cEVeqAkWOAp6H6KBRneKL326ALle
iLvdSYW9jtjSuCsAYuQjOu5BXVvI6Rfj//KrVjyWSo4Dgg0rfHfShJduyva9S3fKxnQh2itkL9/Z
Gu1p7XLdDDCSp66tNDVsTjuel7/WKIwT+/djnExlCth2/mX/Wnp/DV3Jk2ycu0j5dEwhBVbphsq9
lCjcPtdHKSMcVXndFjJf4NS63qCCojedWgxPUIitMnYHnh5VeySGyJLUQluhE8OenForFc+pLqWi
AXsNxzMBE2jmkfVZmYRgzsM4OD7gy3794tOOYuGiRFdJGVsM+K8awB3usl17sHIQXiNdfUx7fnwA
LzOUR7RNBluGrE1xit0+Iu8E59mXHKEaVg1yXg3+TzhgQC8+496OakAMGfiL6ZLMbkMtQE4gdF1E
76LH7OnRQQlPatIFjBk0mUGu/Lz5qWnn1y03nSfocZdat/dIuI1sBxlh8HeQebmDNaabdWWkYm1O
I24Yewdy642Vjkzj8dcQz/uymfDeDe2T7Z01Cld2aXnfrflJlgsJUPdF/IWx3JauS4a8DovNZ+93
zjfet6LXfJW9XfevSloY3GHG1zO6RueHJv6ELhN8u0aGsd8Seiodd7VfBernRHS38HdCFCj8RIxK
loLZQmyTWJLGfwL8KeEOsUruiNiuvBSKXgTtJ272vMYMbPzWv0OgKttkQk/Hj9WmR+ykn66HWUmz
jELhQkWxqGt/0ywM3WZSy9IS23HD+FV13+As+XchnSx3LVkxdkcyS1T4jPJDKEnIazs6zidM8BN5
RNtaw6ZRDuxUEZeJRM3UK2vBCKF4a0NDv+eJclI/OBIaD+XIawGfVN/u+k0KiBGUiYbONoyK/pQw
/WlIQ3flERy6lWxd79N9u5eveJhYBxIJMG1Ez6DDuWRSK4jDmzpPxZaY0v4Ybf1r2EVsoKx5qFNV
y+p72v3HHnNElngSOAtvhcJ09+Ldnm2UkZ+jytzsmys5cPSXvrVVGIaqK4V8OeEzPumS4pUtKyPP
Zs/EXDuEDCAk9nym2nzlnTcTB26jSTw7mRQQZv1Lmqw4QaZsnE2fGymXwWrgAF/fjtmSpYCXrVHE
ss53vdFxNOeK4tCwGqpklJJ7q5N1WbLXjh7UTxKWei+qXVrH9x7eS2NTebnTi2+oG1Qv72maLiMk
wljmldRWGok5+d9jI2Qf3+9m7TRUem4C5QdQBbaHXMEQ1xS7V1HdM/m+BDhcrz6+v9nnnJJBj+Dn
DKt+uK1nCCrjVC07mLnbM06zlGbcJq8uMaezWYyAcZx4uYeFKYfq/C7J0bBj3ld8IH0dDfjRb1nD
9bnoaOYSUcbwrkDnCLeCoZ5AimEaKiC8umvUEcF737rFupaWV3eIs2sK4Bn0Lqp1ccA5Do8EcDO1
azF4yA0rcj08ZLxmAo5juwa4HsOqDFVSgavjA0WNqSQuL3W/0Q6ye6SU5dj3ypgcR8FvUSH5bwZW
xxAC6SR+s1v1KUwqJckzPe8JWmMpdAxWTES0WdxCkCciH3aNMRAvfDvFIL/iNmHiCOFM8Ee3GWoi
Uj3X2i2eqWaTpfTh49Agkm+jl0uyou7qZDFQPOOKae8izpVRPqe/FaKU0xxUbsUeb6uVtBT451UT
GBKKCT8KEW6T4DmnUyZdtkNIqxmXSfwoOXNBCTEEFvy2O3GvAFcNxUCPUJPS2tjn8HRo2mAgOlAh
pGsnU2GJHZbLdTCIOBfpKylsFgcGCYyGF+sbPDU9RRXXi7RyZIeSz7dNd4uh8v/sS9x2yNjfoRGx
es81fE4CLGMthvA42xxWI12c3+dDMMk8sUM2rn3/hDC28y6SwUc86ke45RPxirNetsGnJ2ID7a8p
JrRFqWHQZzEpdtrpqfl1rYB+QXmfQAYTvF3dil18peafkZovQsuV/xez9yBq91h7bXIdPctonqoo
MKcqkqrbosr/EQeonsrbBikJbXAEL/7uRfNGFbfQaZTibtp/jcLw0JDkGtzHS4GvSV4Ei+BnaZM7
4IMi/ul+w9TqEnXP9+PFI+Hv7QMhiHxrNOW6OUHAIa/PVXFbvC4q3TG6piJRfBX+73YjLDmI7Am+
bQ7Ot71mDhxTRKyTCvqvSOAC9X+C5wssKnYuGJLiGmV4T3qoqBL/6cBC5gL0kKxgYCjxx/NePGAp
GRn7kndW+WaaL4Jky+sPwTSIM7DQGrn89FPQHOkTCzxb0PO34XOWZUYMYlKRVatYkn6EADsfabcN
H0KbLd8o0RTV+2yvpZkfNFwbLizB689s0aPtMes7o7pGhvk3fLHOJJSynm4pdSlZ2hEhRctq37Nm
GBMtENhR8exjjXfYn5i/9fmnkPo99508IrzBbpOjJh8yQDP69ZZjwIU2ypiQlzmOLAgR+t8QLRXK
S4oeZsH75pHPkgcwYiFC0lk8Zp2O79yitDPjSfvYTICu2gH2zww1U1j+bvX8YU4l9p/AUDR8qfEC
Zc7fU4uGsRKXZl9/SJR8FHa3W5BYjVnY3DWdUbpZknAvQXqHNpEeAJf+8o2Ca0szLdqApGY4H5z1
ROW8iwZ8fMU5foVMLi6TflchJJoh4wcfTwDT8JZ0c4EkVSrhoQc4i3FwoAPp6xtkXPEAkNnTxLnz
2GKMpFZ3+PvoZaARxlXQzpljAKp4vwhWiTBnPkd5Sd95SMR9UschFKhbqYSLOSe4W8qvY6R09eTf
jIYQeb2JbkA99DyxJe078vU0Xs8rtXgzuSb8gtc15qpmKouD7OgEw72R5qbK//qbysutJ/nue7gn
G5+zId2fnQtEgCCF7wkE8WqoFdhAuO5KU2YqUtFblENxq8Kf2zWOMQR5zrYLwou1LAAEI07ioGqo
/BrRKw7S/1tUEgFMhkltVpkT2yC886hLnudrnJWaI4C2nUk9pQbCHb1Q2zN+9chwdVPQnKZtS9Nq
oi3ePChHDYl5P77AyPs9twcieXX99UbFIKqA162UYMHgX1oLhcEqu5dFdQq6bVfikzXvccNnJQd3
VRtSRXqpFjX4zgYxXUl2gs2SEMjxmO0Zzp8LrOn8QdB6GfAxjMOsSmYGNlsyOiTys/o6j8/NfjLy
Sz4eK8DGB+k7H9d/EPpDp70bCwzeb1yZuHa1HQ/DYlWjTjmSWgUpkJjOYxoV2x2ADyryfVm91x1z
oIdSiC0rIwlFulkKDEe0/yNFYbM4u0t7zhWRB1r6JJeRukCrQXd02i1erRLwlse8isL62gAIYOZk
GQyJvlrHGPIXxOPTPLgEbkdgogmD3gOoGLYEx/fy2DHfFB6K6SKFsc0khaHY4VqXeZfdIQAVHZIa
46jeGbt2ndYRl5eQQ+wcqYEBdONvpVujMk/PKQ1NFi0Ew+LboyBQUQ1QeOCleKMYulxo5ltq5t4w
etKnRW5tZ3TZK4AblxNxAXZ83epzr0yrrAvD2++vbilKBLkd+CEuDgwZUp5Tl90udEQc0tGH6lRl
ghazYQsdHjI9/mHK/QLLQY0b8TLIWVgcxGgb8p+w6m1grQH2ZP90aRgPEjg+8zZQi6LydSgg7TMS
yp5uTQGjS05FWaPAto8ekKeNVXrOD0LgTfy4gFn/tUJPaO0ASEXm2O0XxLcbUrHrof6DEqgZI7mJ
ZeQv3Bei9EjeeX5Bx6yLo2/RmqiKjLkK99O3Um8HPFUDVG1VJcuvNINIuUJ773wTZWYCYICzlXAB
q2nWb7lkNJPXwiY1ACkMSn0OlIboF1YxFC3I4hKqPjgG4gsxTTOSvLKj7vSrkAASxB6fZpj0I5U0
haD1FKXzm5+fqB2KH1Hwm4OXG2VBXc3e/I0IBeHfvwiJaiiuVqhpQpXd3n+bVdoyp0y/uDLRoQTA
KWWumzAQfgh5yHBGE0lmeN6ZBsoA8PPQRI2tF5pWF5YoNFGjsG1t+JWeWfvVS2E7IErxmYEfTJdr
2lo3N+naFgo4jjirt/kCXuYuFvUwIHrta70nXDH0MyN3vaBrunPKok1WCcifCw+nYT+/AHHOTNJr
TojxpYSSt5MzFLr9mQS8fJOXN0dWoQ47QND8EdKvfvjExzHwFm2ldXYjGWbWX7oaTYkHkX1AFFqn
qHVMILAPgWzpZ42dFYXtuGVM4EaFPIrhfHCTjJXpDWSKT52i9R+57+t1fhfOPNQmCoyk0r4ueDea
/kxmddQF9iSINvOKlOZxVVVopSVV+CY3eAjSatewH1tK1g2aVltr7moV3ALVmjYw1m67+OkZTIPv
TAdnjebPOZkFqJRCRo4CDzavQXoCNRnRcDc5CRGBeF/Pvdtc4dTdSp6BZFha/DZb6gXC7cPGddC0
r228bl2IR3Gt8YJBAJvX0V6v56FOnh9UsEKVO1T6/N+Sw+/lDnxMq5dCQNu5RickYMDoCYjTRzWH
jSn/YX0NjiGnGexhhrOs/u/HkFHOBCFOUM0trPDVwVdXZIhtYMloNFwrF15b/iJd2eYsxK94bybQ
dH/4/JOacy/b8NJdVBirK8vcziK+RkFyOt1LnRLTMCzbB/Ym5MCrZzZ2Yi1yRa103afqU8QEqtdj
XL0eZuBSmOOO6lDzLkFrHoxvVHSZyO0rMy9O5vUWHnNtBUQaBB0E9gc5APa7r0YcDXnybzhLFJAS
OpkuTbDSJNhtwG1OPQsDNcQDTcy0oYHAsXN4ZcmQslocl95mk2nA6V5RKJQhHWu1m2iIj8xGZh7j
9kArnG+fnvweJ31isA4bxODMrLW7/Am922bN+5EXmeCAFchrrlz2yurwKYhzqRcRHCHGLIZ+43U2
F5/4rnSdwtfxXEBuom27Q3NPPiLtSFbtogafcFt0sye1esQWqiXQBlm86k03UtO5a09n3iIRHp4e
JSkVi3Lv7M3Ml4tQ5ibd4OfCAholvl91rCbVyzVgX6KNhiO3WuNgJ0NyrbJEd0efJI7tkAVrAsQ5
/saiQ3X4kaNLFznb2F5FW30IglWG8GcrevZm0p1Us+dT7vMDT0ELGMppklgLlMfS05gxEq0FpViM
JhrITh9TSR7cWQ/a9R5o10KU+w8XIghS95GRzCGIVQVfWbmF3URVxURO2t+lDfXr2W9i2q3d6SVF
IxWnGDd6INz0ALmVJTQT1f/Y2SYysZKWo9Nl5DUJAuc2S+GLwKCZrcf92pDWW0vkohhdfruU1GgK
OaBPHorF53RMya3a/TrWtnqCZ0qtl+nEO8/DwbNWfGgWCKMLGNzWFAL/dqp0EAOcW5ttUsD6W5nY
u8oOgcJRgMowV7TWvUz5WuI9ROHfk9VZ5StUmgndLL4hRRK0UBYhFbLY5pFg+2CcbbKTNoLsB/eg
v2yyBtdYgYIlbtI0lEjC+CPNL+vU0JfWXR7/P4GYnKBDi6MgDoEYrwydy4vzyPE83YypJvHMCapk
T61tLPUg3+EALyeJugWFd0AufF7fVVfQLmkqC6Zby7DU8rCkSUNOa7xqRlHKD5PPZA2IMrExLb0r
07rlNfIb141hvYLgJqgtLsDFhMbMJemFNkNj5hPDwxb49+JHEdGInRBgNCQKmI2LMblGt+fWQBhr
SDs3cCkJcYAD6cLvb3TXtbfSillOkcrXqu8tW7H5cVOY5+UvTo+65QJb7Utu0JNAuYrZ1yR+hk7E
SqmcvYp/hLqFAMk4uDOquWM96DHtlAqjvkMlN64WXXaUujHp/V+XslGGxgx06xb2w6EmH0Cf9+lH
Cs8/o4hDnwiz3Rslut2TW3pYGkMBDkVMo++IBEqxfPc35pyTdJp5lKDRmgIVEA9hybpjYwY7vZHX
iC7qElT0B6Yx3SjkNCVpzJeQj/VLiJyRVPcMbouSCzdTaEUGLNw45z126qeKvutPPn2irnclCL60
cDDfJ8W4TGVxtFLPOBmiwqHuGqOMpfdfLI1hKDOyG3SeYCcFAxbZM+yrimJyQSlCvxH7tXaahUr4
iqwf67Fz80wLO1BbuhaoQgiis40NJWyNkcdR77/GTUXT6XPD4NfGmvh5UuTdCMWAcA+198b8+09K
d5tBnOkGKDQyBUcr0IRnQWY+kF6R7n25yIl0GAzAAXeOiLc6rt34744OgxHDHRji3Jsvv3C+EfpJ
h3mwCtBrDXAQhLB9cuLLgWqwi1uDWtt3VvRSl7kXVUNoDrrEGrM64GiDH/aFIrAUBvWy0csza7HS
i5r81DRxRUZOu3optx7iFzaY8Y/dzgxYxFh+o+yEue+J717MnZ0ZjD/Cod8+1Uy1pfgWsWgqBKcv
QL8lK1ApaQYDJ4poTVw/+Iw6nz4tF6Efg23Yq+5xCP18R8J+nJSr4f/xlj/NwqVzBVjXj9rgX2CM
fCiNbnTiSQBvGUxTJvBNCh1jtskScYm+viHZN9Q2TgFDLUzqpOHjKgmt6huU1tWlXgjMyfdN7kl6
qgqf89hv9NZuRenW/6r2jtwoA+yvlo3460N+K6Y5WSDKjp5tsFK7qG2B2LqIxSV1WgUklCULgcb8
en7/xKl9IqDzLCE4SDA++Hw4m0hW6uLcFDpWV6Emp3w1ZPfMPk8sxaVEifpxXLLf58oP8XWELUcK
Eb8Jo9nh7lXidkdDYr0QiXYQ8MNGxa1bDRGqO3J0Mb/65zLO1xpSarqGr1GZ7gbCbbBN7rVnAgHB
pc8OvZRBf7uH02YmNdLzMlF0+0LVsrS2/AVTNp8OfnaXH0FeJBi/FyZ6Os8M0fSDHZwy+LNoABiC
78HNc2GFGaas8tEjcpapO/g/96cm3YIcGSmwGUl0eg5gjPhq2xU7YPckGhlUlqMHpFEb+KW0nXg6
skAd7y4i7YiVoKJS0RFsLFZyrkt+Z7exNVh5EcAP6iP46lrQryRTaccRScYsXD15LX5Cwwuvp0vO
J6ooNbGfdUWJv3jFHvV/qM48YuF0QRYINtkQG9SyCQqTigzPrFPcvqoVi8RWRVPDkAmyPN1yub/n
PmMJOMOayZij1Xg41mVXdhDXdAvvqzzq6HphIyvhMW4skI4BypbJJYuGsMvtXKilXz+0RDX62OCd
dTEzw6/J4GzrJix5X/gpZCirh0O91TkcdsBAZ9hqotF9CyZM1UNpbfZopaGKNhjzw11tMiFez5WF
dIeUtB/Ihx4isby+w5/orDfXfxBlf6MZC/X+h5UGg1crO7h9MnsHcR4LjXVTSKtDggktw3/oNFWu
xuHZdgs+jbKQUEtI8T3GRUZRX0gHOExPZEXG5n2ugdVd8qiq7BJcpDrKVD52XdTPyCxqu63+E0nd
v2gTIw73LHVFMrwyFgcJLrjrTy9D7H8+F3t3PGv1OVuFKmGiWHXCXPWkjQ1XYxXoylmz7sWY6Z7c
wAqRYOYWWv3lps9Wf1OBa9UVAa48YwRitvXlvpBOwd1b8xUskug9DIk6uqiLNJHsFk9mpGbl2DEp
pFgshd4bJJSjeP6oLSeNLwKlo1iOlBGk6ocAIicbScByHrQOoJbLKonU1+AZCR4hAQVX/bZ9Qu76
svVwitirWqi+xMMXgLFDLfxprpKg83MEF2JXmTBuBz3Q8HqKqtcula/A9TmhFlaTZzDt8WMZjeNv
Togvzr+BQD7tPX3EB+J2uZ1rGy8iy63F8uA581r+yjR2O4EPHj/QGd/Oyvicflp1PMqi2Pgskot3
t6aumxtrtFs6ALyqcsdZvYG5JD9DW3EXKpFaKIv6DwqcQjPCdtkdJrF+3QwoG1sKR6Bw4OpV4YOk
OKzHhOqODNj69HCsxfXR+uDvt8dkLXcHGC782ltFTyccM65wrTYS3V1b5agJI1JfpZfiLb4fVb3S
+rEBc9ztngXHTjMdSLL50VQQ6vYoZAc7Z/m8Un1xVN/53F53/d3/kitMnlMn9kW3epZgaNCKczmu
7hV3GUVC3JPzarlKBbwfTqqIkOm/xzu/tG5deYkntQNH+O383ZYPtL2dvND62IwOxCtfz++k4U/r
45ipXUMEA2GQ7VaLR7YbDVgYs9QoMics9K2kkYzlpAyDcGaBGkFlFQp3iiU/U+Dgmfe5PRsTZjOM
vEzMn52OOyBrC4RVohcJNHwB11fi2NgI9+nF5vr9Aa6VDBKsucjSzrvgbuE8Du+WFrs4CNOH6qLd
T80TplUM8I/I8PKlNCHrs9OCWOtUlrjErF98a8eyNILgxCqjmdTwlWGyruQ3u/+fRdHfarudXJT2
BJS35LVjBy4swZOdyiaRoe5kNmbWQYOZGdpxANG/xqnOOfKG4FhXNUAkhLnp7y//tWSZ3qb6svcQ
+JDXQTosP9/VkwShMD7bAs2Zhe7QUM2DPDEHWwSfqwVPDa0wBz5bDJpFFiwhHW/VZCAWOxsqMtDQ
E+FCYYE7vrNPkTQWVovUmU8MPT5QX5B6TBWR11ur4TsU59JJ12+ETh1Yh7aWN/LiQ7jwxGZw3drN
QBHefXV8b+REWhDiYHzCe6opekTQBzouvl90jBo1hbOrRkF1AlcordsfjPn4xw1NNeoL1ztlbJnL
0G0JS2+u7i68SoUO8bh+6SJfKWMWxgCUfswfrL1BnRShW7GQFZYpAmFnKLQ4eEvTkRNiyWzHHZ07
nVHJ3ASiDd+H+lVmrrodh/iIiw7tPlR5J7cfZb4XZzlGMJoKXef7tusTHUZNH9Erb7/9k0U4cPYT
3R9XNgmuxTBiA/kok43eEVTe3el8ESbEn+zHGXqFG2HddG2/IzKTaCR8NtfLO1FWHwo8byIRTMQm
AH+vB3fDX49lhgzoyfg+Y93Y2IUTuL/i7CuiXh/VsvPMpYaJgmnBnbcuXR+dOxV++7Jyt3yhGhFS
JXbmnTI42Ib+UF/+4h9/UrNqsVLCdYWDoSNBn+RnirAu84JPIjN+eDzVQeDQyzjYHMaboY64qhOB
/I+Lxu1spAa6xeWtP3vrPN7f2k1iaBVslaJh81zPwSdMFuoR10Xc36EC5yZb1IBh8/peVlpv33Al
hVWoHqDDAgfzIUY1+iaKJtFu41zZEWIwV7yXhs3ESaDNI1WslXY6rjyGgxA3M1tiedAt4PzvFz0n
mJIY4XP5SFvgfJV49JGpxjTWtZyDnqEx8Xl43BUWmNOF00kQzQuqgerzq/nM+8ndvXScsOadLYfo
O+HIiW8swVgs14n7YAz6I2rsux+b8Cm0HVkWRFWAy2Q1SLkgLceX67jHTELabuFN4v1wXvJiNvOB
gbEjQy05AeYZevBPVgj6WNNwlw2htqc/PegLW79a3ceUsHABSI7tBi67voW8Cw0Me9JE9DeTWzBV
Im5dk2pdvDET+fjWfk7qxQtOOuLQnag/U2LFDCHBjHCmsxiLmGN3gOEAlY7IcmfPHrQe5e9N8+vM
dfi8/BGqJyXLxa9Qva92H9LCNA9n756BD41X0cih+ZxbHe/NBRPrWtNb+LiM4LPLV9xaFuVMi1t1
yaf2JC2unDY+E7TN9Fzfg47RAoWHaLcUpEGPqGuEOoXGNPyfTxdlC1PmNkHzZ5WdqwZZp3CqUboK
R20a09yBzFHVRtokjB/rwcQu63pnxIoFxe0jlA6+zr5IcZc3ztuk+tLjTdcOogQaU690CyyP3pZh
46AHkfsuiGdxOTYCPoE5Beq0B6F9ZqZGEKMiHnrgTJVXKnhPImfOkszS0r5I24wFw591hCL8xdv6
KkOWACAdjMXzm9uRr2GWziXs8cXHwDk3WyEBysmmoDDjAES101PeoK1ZpWBVvyhz5gmtaIP0fJn5
ux9xSx+Bb0ihu6kLYem6Usr/Sbw9+fFiUebu8WtcBP8uNLhki7pYx2hNd+BZx4yWV0Ysn7vUilQA
6rfgP8+F40TyZm7/4mKoYDMLW/wUkI7Yq1sPfxAzTWLu2Jkp5Yrlf4sOqYvibWPjOz9fTEQh3DZm
tRLmK4S1zCH5eYnGIDqv6sn97cUlBfc0bTt+bh9T/iELc38r3M8WdLNCL0OFHqME0TdGrf5Ldz18
wgqLuIuel4BckddIQGQE1Vb4FNS6iM7FoFzQ0Btb4TUMxt2Uj8PUw8LYINOJfANEVtMk3J/LsqmE
+wzsolCFfnB48ad85mKVZsxBnrEYJ58/F4oEep1mjEFDzkjopXaoH7r7by6QO8BS6naFdFr4MJlV
cxOfMIKkQIy/CQ1aZhb8DVpwaBLdzXLZZ4XQ8vRUrErFB76l58zupaXT3FtH5XT/slMhFZNbZGGb
NdCBbHdBR9ENVQJLFkIzqXABuv0EF0EyDgOJ3cKMSXEHdao6K1qNMUDvs7ZSmJdm0AFipcA05hYy
gLuGnbJiIUtDNXTqZG7QscYlbD8Ebz2Tb2c3nSblCv1RAgoL6qeI1nBcaXNCWnlYARJtNTc8OEHw
5kNEYegW6tk6ivXCyDpny7rnRmVoaE/Ful5U4S3AchsCnLgVqmVZ1Cfsg+OqHB4v0YDpPILk82pn
0U8QUrnHsESmslqtGFGJIfBrypNSX7x9cyWif6lMTzj7mpSAa632V3neBQcQCDorRHv8TelTYiAX
ABmAELE5VQMiUKbdh7fzVCJx6o5uLJtm9Dtw9LpzefwKjiFD+s5eU3ao5l1FVGM0CUwPjuc43PBn
EazZjhtB81DTvD+AWZ6XnD9Ww3dCeTUM4qSYilu1E5TYERV9g+ttJFmkC6PMD0opC9dWIOsSwzJk
+r3lum0XqJqe6/QdRTQd7llDri8SM+puX7wQ9QqrGUwSHcDOHTSt471QKQeo5VsFWpSsUDNhVA2K
V9W0TIb5b+wvk+6Mh/Vs8Dcmaaeuj96D//PsPeY0iszO8f5kAcXXw3Hz/OQBk14YCv/1AGb9zBdR
Vcb2j79G3I48U1+DFPdP0dVqdj1GYLZ+Rsoias+Z9hH3hrameANgo3qB5FBoTieseHz51ogsCPcy
WODXMJy0XQYHoMwyQ3TLffOiAL73oX1Ou0VLMKVxeI6yQbfxIp0MqQDerShoVj3gY9DR9ftiqIWn
ihL4b18Ycc4CHNmfBcIUeBTB5OAG8yaTa6cezk3HgdHITW/Gr60dpVqYnnu69fUuORwkIIghLHJ8
bpOdaVk5RKYRnmjgeFCizO4mxDKgWVbKHWpj0c0yopsLLsWpJpl77IxF6rw+XqV2xQOllCKvTSa5
CZfZTNHlFjMl/vb/OGEd89k4hpDHiT+Tvnafr7+qnj4aSTUsuN+zvVFZBs5z3Ix/Fh6yF3qxYr03
MSDh77YU7MLGC/qKiLn7ICvNRUBRFv/p+IWTZSu7dOFaRYWM3yWUbQGnkjRjqxogNqbZRX/rLk6R
DFjVdAuQYxKD6eyKIYvki+Kvgw76/YKOlmrvJo/CqeJMOpfX0SKn/QLzdtuSXiZpt0ra3jTsEXsr
qGGcg7LxdndfwKxo3UqRd3iTUJxe7aSDZix6InyAqY6ZAierDsdA4ZvDVST3FO/8yqR/po3ta6y1
H2sIVEr5A5UC0i0I/YZLgi7WnXAZ8JwUSvdKEqibn9ssAceAB2yvNZuUlb/K5FGS+rQ1YznlP91o
eE3jgHGndqb68+YuGvoaej/RN5K6UN3Nkdl3QF05HKzx+RZPLcXKeyu9ZFPBTH1JhGqTwb1+UHsZ
ZixPaX+gMmkqUX9lywm/M9HeQLQuIf7MBssUgyupve8V7rvWvPy+ze8fhDw2dgEj/wksp0SomWmb
ErpVzrrTRdBYC4yp39twMioG3/XpJ54KjXuI5FJAcuE4rLhmXFbWRFAvjsrRR9nCQ1vktYefNuaR
Yev8aahUK4LW1OkAuburX62CEPWEJSn2ZVFOQoGzDp9FXkGBq/UzeDx4kZpZtSOUkqUmr9gO2qoo
QoTCvVROug0qju/u5MRh0tK3hUArSU3ys2CceCHmtJlHDVzVvY6DvdpEVH72v6Cn9OP9+9CUMdH6
7WqRo3bxyahGfmotlosne2NwEkSeQ4xiySxVIuruyWiEgsQ/pTk5qHgnGFEq8yESmwcIC1uwnU69
IRm7jYR5VfsZJCQJS/5zJnyeAJ8RK6vBuJzPLOLSg0NnbzCZGvLLzjpSDNbzVB9pWWi6GRv6quIl
5SUSAC5Ck/zA9t793nzr+qZQre8NcNiCee49Ak5TAwaEyYyLjAoCODKpZ/hif0fY3MTxs+qHxNmT
5tXDoLi6qKX0iOrtqs5u48L3hIgKzcah6cJT2B+Cit89OE5BU8YgVZN31cye5yBuN48I5nY/wzv3
d3gs3Yj/A9Hb6BhrmX7cwQy8je8zkIzVZVFc8EUdRiXWLnC8DO1C0KN0f1kzFHupj7FvB5daE608
iDo5EV7ytzz9PXS6grOVUxqjGkckovtExdpFTGs5U5lt40RJ1clwOqBkv2fXvSkQ2V2BfXq16yAX
L/LrD2UnB7iGHCnYCxKV8uuBGS3TUtkfBUH25QhUaBxkvAvdF0y+MIjPvxMrK27pq5NFyr8DGAGP
tTTZ9Gei8X07IIbgdEebYdGx7vttYeeBpl/0hTIud6njhWIV31aH2LXB2LTyaGjw/liqQ192ZBba
M8Y69O/6wFQIOk+kVAWO86cIW7O+rU3Oplz3TGFZX7kwl04Qqsd11jx1LYXJAoP05POBfrFhpN7y
lzx8onPbSswd4knSxoSGbR/ZCAQtV7QtO3MxzQuaEKad45DBU5+bI/XXJ0jH5Pyq8X5ZhoIVcopr
vBs97rbY0ltiLH0iXCLFAz6S3Jklb+OV9VbxeLtmXC4d7nk2kUOKe1eFL8lVpGEKbANOn0N26slp
HSl84QpYwQPKLNdZCPuYvdZC+LPv32MvqiZIxawrXjsEboL1ZfvwEVrD8zI4VaYqmEbmcYNLmdpH
xE4vuBW5CRh8Wiw5RTEyKl0Dt87nIHCMEzna5Ko+vzigMb23c3qtNWirX9iO/Y6rOe8JPE4GsEeR
ee7lXRwVcZWI9mD33Lech4XbH2ucIYTwnLvRhBUSu3BjXWGlbfD7bgkqEwGADpzEJuCyXvWP1v/j
dQt8S/l2vb6Q+bVRzIyECNgvHipyH78CowOVKeiZ4Syk7hurfTJRB83UiFS/YYCeOaSqr+zDofM9
e2SHWEAKJBn0m8gruDXYf4TGIJc4jQCMV4jPZHv3HTqSOc5N9d2NDMTCs44UQ23PojaqTMwZjKuC
jA2X5JaXcTR4hK5CKZ+yeKH4u7mVrIdI/qdC4/YpNcYktDZsGH58tA+Oc1+og3OvSq0AAoxyiawA
mX+YpOvQdrHgAebHnqr5wswXBTMZaJGlPpZdEyapDu4SH3M+wFwYBzvvo1UGg5iikxiXKWXnr9n0
vtJrcN2THbS6SNeUdw5rBVRG83bZ2KlKGQfnvZ7j7RxQo7LpWczDWM3Zu7vjzXI6bDmJDsDLEVdL
aMIWhoXvagAjnav5lZYuzfWFOkipKpIt9OVTIfEikv4DzAskgluiMmDwO0AFAdGuNkoq55OZGr71
bN5WH2M28wqAEic2X1TxatMwFBd6N5NzAcdqi3N+J6RNRtXGTJ1IqnHvIGW9QejoEzUOc0YAf5ro
J0gTvGvwE4BMqfMD5f+n2sXvKz+boY54CoCV72CkA6wf15K2hX166dU7O0/Zx8JyeCq6n8in+Dtn
y17BkMSpVjRB5GWXytgSCt9dV1kUjclFHufRSn77zF66gGXm7Kvi/RaVHULHt7X+snl0fbYRHzOl
/+r6bgJ/RNsUqxBfM3R6djHmdRax5E1ZA2gRJanSKauMvWCsdvV5wc5AOcnNNzHrvs/31nLVJkoW
8vR2tXmRGhWybt9el4sBlQqNPjyTBQW90FT0epU0vDO3aG4u7aspuZDHQj9+bboMvs3d2Teb5hqi
irWIJotdt+DtCX5XXqZyczP8cwl86H3Osvr1ujooDXINeKlMymwRgvxHR/fSn+0lwS7Skuo4xDLC
wNTvS/8L4IoyFzfcQ8PsEnlgUNqoe7IMSTW7PxLkgZw6PugFxdh/iEH7Ebrao+PMkfPA9mfu9yVy
eYTrchlsTCz1oFf52Kh/xum7nWPUZYfIOb6B2TKBEY5BCvbiZCShjSlxC4j54Yt6vMw2ehgz3F1f
KSkUG7kyhgw+8jKyzoYU0R10fE7mpL08DCBI1ojBGpL0+4WVjYBIlnGwqPXHdg1zL8Et6kYiur9p
elAqPHENogbgoMX0fOpQASzTem6oBG/KP+lnWCMNa46U5rey7RN7EdTtnMlotljHke5fXgEZR97H
eKRt924iGWgu1d5yc08YWZO23yBsJOD6T+JnHAKMC3LuiZxRJklryujafECC+wVE3KuZui1jXExA
xDSh3vSP1f6q7LiQWymP60/GhJrK+IdZLGJo0wsLI43Otes3cq4l6eNc4CdVlc64INE80T3aEMUY
wrJVEQlRg4iFLmSgzAhaxHVo1HrtQPa39OYJoQfUvR+d6d+F3P80NPdDBa/xA2NzV+Va9GTt5lzJ
pRIOHj1+Gb8lnB0+DL23QMmAcwHx+0wdegvxq8xXhTB/YtYISHS6zvZkdxnb/k9+IUEuF6iryUFd
0w+dY5KhjH7I0CnPmKqZJwOhdiVwF9xcYaMH5XlMujmqZ+FA5JWQVtf0TmiPN27juSv7jbNt2yct
6wFdWSuH6p859eXYS7gUTBWrTyLwyvN1nfp7LZVzed8bKecibWibUuo+2POVf3jDizN8yQu1f3Fs
Pim8yguNHTXtp9L5Wlou8PPagEUmsmf9Bvtfs5ib2qo40xiQnsHULBrZ+8H2QhhmRJmH2wfDSDg+
HGWmbyyVOWn9erbBkKfIzsJewhr/ZuFscL/IsnCvNsHkX7uqphC5+lhmBk1PV7SbjiL2G4f7w1Cv
6xGC0tpdMlb7IRTzqhkwHrRC0EOMu6yqtEzDiss9o+jjijO6y6Q/ECOvxD9lE5/ZUaHDcoZUTZ/p
jtM6VxDxbBRtfnYmYeETOcmLriu+jUQ8ULA+W5uHxJa7MEC++rhhARaJnyaB3z/9wlsV9QGrZAkx
oYgREYGCm59qT4hMcPfWmGheS5mDj8OVDdPxYRrK72cmjmWNvGwnBXYa1ifJIfuNtBgq8WY1NRTX
Q9hWj/TPQUpv4d7bXmRCmHd1k339d6jzUfseE1n4ig63SB6D9T0EQNgS3mT1U+waduyj2Ds9ZB89
odBaB1Rxa4P83UItzJKz//SlDcCW9W1To4N2kAYV5dQ0RMRgPFO0nPJ03cGltJ8v125u4a7QyApe
VDPjhhZjvFnsFuWV6vI97mTfwH9KZ0Xie1Yo3QIcRoW7pBSfSgmaiAGUZDOLVhVp/5e4/xcu8AFl
9lb3duC78HnOdkC8UHmZtaQi0EaUrksZDRWTQG9PnIX0yYmDW8I5fGteTPTvFwczLWzzNYAm9BYx
jafdXymReyClmTwiMRBqiI/nuA4irpisN0pmgZjk8sIOJKAWA28L8URUbTNBfFJzYrD0lwNs+Ga6
ew09iRCgCRg9FaQYRfSHIWXoJCxXJ8lOtKDx36famKE2mANZz2k0xIOsIYDh3n6egkJR7BgWMr4T
DyVin+0WR1G2uTUgallMGfkNO55QTO2cOhcCgLtRUFXJkV6y3cdjuPCXWsyXzGITxvYBz9/5a+rS
eyJ9bVaoCC5iBkVqoFsduEOnf81+wQK9hRALALoBTPsoyShKUlP/Z7J/XGeSqEwkv9NJIb5TEgzx
cg/lg39vj/M6EMOnCZB/q5frFnQ3CMVlBGRgOtY6BQmTpFz93mJGah+j7mgCP0cm1AJ9q1+ot7la
DQL5w79HkKw/KK2ZEVKpTpQFeJa5acP/OnHVBDMlX2I4oSZGQlDJ5UHqQNGeu4QNuZTv6ThQnDtX
Yy9tNH/GPsvVkUOMdJaPgc9yfXlrUiXwQBNDLoEPgOABja2EwrW+z+W89DKSaX8p7hgoDVi7YPD9
8ufizlGKyGguR+ZPgUXdqoWh+ele784CrNGE5e3CotzswYW6lcNfxotSiel4G9oxwMkLjf8Xf04W
rKfKqLAYeMSx34o60vItp7Ps1rSSKBk3XOoGCrp2dnCVj63ICb95ejeHT2GnwhL8zJRQaR0mUrzU
xGCZthQDzuoBzeRG3mtY4SptRL63zJZ33sNhywcZm995aQYZKDHvgscI+LjBWVuMvKqtmuWlTamc
FjG4eUjwMER7riLiPdLEX82+ej8yNfU2A0xWgUA+5t9U0dski3uKcetDO2MGUihdOsMh9hhfrbUt
JvsQPkC39czBpGULtSWUC09NtxqcS7w2QIcej0TUsdw9JRN132J+71gMf6sLGGIxVST1OtULxBAL
2Gc4XRxNcOy3Wrg0wQ/ZUvBUjE85pZ7eFOGlPsU1B2jAJT2xXqY5tyd4utUA2HlCzVVKPADaocvA
y/mCtEQVQvdBOh2n5T2Y7GaVWeO3wmdvTn+j1IELAiLcNulkE7XfoaFzbl3OVlt3Dp44cf52O9/8
uP6YcsgY0SFDMeisCAFxbYR98oeuWWzuGm0tr3vf3spsGDZ7G7POr2RpSzRU4P0SwW4fnkd093Nk
Zzwve57rpVver2+KFdl70w4me+b6rcIkym4iDu9IpxJtYnO9QCPMrKwX3PwDeynBWsKMqYY5/jFg
e8Z/TSgGh0z65JJYr77lGb4RSzOL8804LHl3DTpWG5nAINx8svMLby+6PrINFCmXzH/PWL1vkGjn
i5m59MznFuFSDjrSRjZ5MtqNTNu43fB46amtKzNLsMjzQCfN5Kxk/zv624n3+EzWmjgXwU9d0L6R
4pwVr5zDPPYDFpIB5oWk9E5ItvvuJZki0a35BQ3RgP6AMlsEC1pjusyzynaz3t8aBcfaz/1FnRdB
m1fFljeakl+8IIHCoqfKsZS/15CaAoxFkJkISefkkZC+fzGt0tVeCIkJ92+oU1Fu9xkISj6LVy9/
8OJuboQcriLBV9EAxL9lFbBCqXmRYwiI2GxeepevEeIGaqgCLVsQqTMcsyf2KkhrkEdnLpq2inwP
CfjvawA7pjclIv4QG2qcMxvGPxRSGMaNR9SxRYld4/JLIxiJ3SjWmGKngYDh2kRbT3r3OcZt1PGL
38PSwHSkak+md9jIoDV8nen+yeyJvmFPlOZcZG4lUfSI/ayQqEyFp1Kkcw2ZN9BDdOuiLwEXAF6R
5GTz/celNrmyPy64H51BqEZCOxFosbQEkZYEihE52+erFma9q8TwDwnrPocM9+98zNLe92wO+fpz
sohXzQ8ppZRw1G/w+7XIDbE9VS9ytQSQJbuuHv0Uf40ELFwrPYf5oNbxQzBuHsdpkuvGfIEAEFIO
sj6oNCPoFA6f242S/jl5RG8+9guftD4CJFxyBBymEy/Ad62U3DbyDbvZH/kz/j50TJ6+3FNQbnUX
Fd6f58S5UjPP/j8eItipsE/P5nGv8Bf2wM2qz0rwaCX9CTJeAfDug7ym/RdrBCoSpvgMoaefM5bp
8L4ahxEQOL4pXbOcPpBt+yLx/TtlJELvt92AgdhgmE4lGdRizZhyV49UTeg4CvXHtClBuQO2E1/Y
nXLZp6/EUEjuyIpcbNw8x5b9NQccM2HKKbHpNJzUHDmIlCuCgLuFYGxUopdMvC6AuDG9iMXE4khn
1FmH9mm34VvhyVxOSU71emXb/h5GFLv7EU6V9LOV9yDIx/TBGhFVIkIf6hgRLMUnoGmEmY5wPlIF
8vyNzXk/wp+iYmSUTKIpxL4iHEAYS20yZmOvaaJIMwfZHpNPC+Kt6kZiUTdw2izsljdqxMUvMZGR
yeGNvqK/9B5u5H8h1NniWQcNsU8gO0wLOZoccjGr6QeQM5Yf7zcWKEkucoz7iI7tSTNmVG8eYFAd
nxEGP+3MI3NeWNTXiLN/wk1BOKDXAIUkj1Sn38hBBiwXaz4Lx0F1ofDHxZ/OB9/dPbHayuA+Yhse
9yGVuaDfWPpfNTNy0stF089dMymB+xvQhvVXGSofbZfZXhTYGQ3uOiohM5Q+GWc/N928TsYwSLzC
cu9m50VLeth4juVPjzUBPNWVwm90w2zorbtsBOiaigad3yv7c86dqct1BjJpoy6XCAvhRMSi2xqd
+6WtuKjnVWil2m19Hf3InlyigZBu/ci7zCcvsPFsLQ4VeOhVZOsluyIXa+QiC0f7Epy7N8PVFmxF
JHy/0Fm4kuLsdDABfJObqHC2zHbUfbG55Sa4FoN9o5clPBuUg56hoPC90CLAK5Z6dO9HYPUTyfE+
Z+c1bWHcfGP9Lx5qzQUnGu2jooTu8w7dkc2DNoSwcHquOX31F46mDhDtR3gzzF0hcowtYqtCF0Vk
bz5tMNudE0vDuDcaKengAo6vM4obGQYOjljSUP994HGQ28CzF7/AgeKkMvj14ouO2wJHGOD9E6mU
PV8+uyN7Q4Qr7tqQwhDJtNewBDGbzI4iijMKwxkClb3Ew5uIUMVOEf34uKL3O7bdl+wVvOLmeUeM
sxTD5WXIsFzjUhxXJSpEErRu9YwHU4t6gwURm4fYfDIpj0pJNwNHMjXhEPaJ0iuOGdHKsJlKLZQX
5D2sAsQc4GgxozLHF+K11DmCKbcaNbIn3FyukyI684ryx/0Lv/MN760Y8yLOYQfYDm5FP6AzejXr
CiYrpxNXivV4WHdLwYd26ciFnihukHBQ2nDPOLuYhhslieuKKkUCdpKhghyYycJRZwOw69TvHhxv
XWY8cmQK5onpjqniicId5MffHC+bWJWzZFwKEWvlDpTdnXXKjIu3o6s5XlBX9qRCe7bEWMAdaEoC
cchvZ9M0WLZ8WTOQUBPhfgBG18TiQpOEO01k2/hcODpNbh0UYNbNVVehtzDivorIJxkQBL7sjLkk
TZZw7eFlUMX0B1CbwHYM+ACgUXNCy+TgBfxSgqT3oqB50G4MhZGDSWQbN25diqOV+wujFYApY7yQ
fks+ozLP/qoKqWOgbz9zr+yWC6uD2Td0308EBOMEr9G3GE710peZS32hKlVaQ/Uu4F+whISW2oUH
D/TKNFWrBSoOrQLJ3zlVKrTxeRPtNaelziNAyNQZmQpXPMra9yP6Ydu8+438WhdfylDn+k5qV2b1
Yg/00Ob0RpWJPkn0//lglaVk3+extlqugJU0/zNiVRMzRuvsLq/pcIUuszaKyVzVczJZcOw8ian2
kvsTgZST3TCdJMSv5uDhFgBAaYKpSTJZnhEyaamyEYq33eLB4T0pxVJ8YYCeJWlsfGTxGYRuthp+
P/RWgaKb4G1AH0wY1V3R/qsiF+tWqG2MNdM/C/n3+pc8EOgYOCmfQrAZf5j9a0cUw21n80EmJrq0
S9s78W1d1w+KF944N1aHlZUKI5lG4u1K2Tzb9oGAB2Epk6hny04lDlBeQ37BEUjpXZPtCBLRtcqF
AAHMwkWww1MV8L0750WrYaG5ZIyq/S6N/KJEL8QKhC1CiUCewg3GbKaVexSFWWYaDjd/3sYU91gr
fGcxJa9xF8vdnvYhF7CG8nZJlIDDmsSOWEPHoPUtOu3egR7LD0EMgeNAL3q57aFU3igr+3v5aUGS
MfasaIfK8zpVZr5qII8EnhQTyGssEwom5kpqfzH5KJAshzJC8/4UWnxXPXSRie1PY9gIkXEUdJB/
+zvfm6+5TQp/T6zv3//eVygoxMQcJbj/5uQSKmuU4CJzBtDFFHVlJ6O8WAieUoySlUrzs0HFPl93
2ztMC6hqN05ihNQ4CkeLPoFExrLtVnPdWqhkB5WKzN4J+tNshoPEWBCrGz0PMibpsyV6vQTihEEy
l0IHD9xs1L3PRSLE7OzA/jF+rAgVP9xpV+2E+TrmO1N+OCwpH0xhn/uESIEaAs0Um0y0wDKNgPRp
8F13yjAkDYbFLSio7ZuJ+rSP7PociA2KTiTlM3QiIh/FWz4tshGIe4BRhWyZJC4j+g/9JtU7Ae3r
U3BY0fP1H+bCastns0a4URjIm5bQ5fHixq0qUbx8ElZCazKDUk/qlUzXNQgwbsFJT5RD2jFAkSrk
14UJ0i/zgEYgwNtOAyjNWN//GPASVqEXfGQgNdRQB1JuZRcgFh/hgf3i7fCsMruDN6vvmDJQqnjN
v5/gfNR5QbaiMJIsDFSvJvlGLv/lEXI+RwLxes1csGJ77H0CWmNe+BjIWTVbuEW0lbZ/lgPgkcnh
gChWpyxwfdCyDjngVaw94yOUbbyxxSO379CRdKdCem0CgePQsIWZTikyh2MHsZ048rLh9WKP6qnn
Y0x9YbMmmYDUnj8qjyu+35YaJA1kgAsJ4hHwTZeALBmx9yJww8EUxrkaXObnHI58FcB8ZvcYhlcG
GIHOuYnbvt94117jyLI2gzwLfhoQcHthz5N6731MDEyRKl2tgK+vsOXQNSuGTh/T0RF0yyT9MWgB
IQTwUnny8bOkRjoBS5LiS6HhRGo67TT6COIvnwO5P2C8qePrvnSk345IXg8dzeCv4NFX4LdQpfHt
PNGb+EsLpRWpWeNJneOcsvWCMqB9388TbjEkL5tULSyr6MawYcDiJZUq8ZsnHd0r3II2HwS5td0D
Wd7vMoWT2+d39uZ/sLgxGE1XOxZj4TIzdHD6cY0h7d9kW175tOvJXk6AyqiLbjlOK575DUBBnze3
WjvwLwqrEnyWWLPrQO3/SBQbFYTaasQnP9yMSmoHdO752jjpxZFngmevNB7xB9sADeiAy7/QqQtv
agWfRnkvI792gffW7V5Cua4ohyxOwg4nmdhvRwZaQfYpbWwzw3DyMIEy+3749oiisJ5YGhOs8CF9
8rsaRdWrPLbou+wnV9gvA9exd3KDUcEuYkbDaoimm1n7VlE6FiFzhIry/MGb7C8FNALyDUChVLmt
yFCyPurFsNFm4USWwilpATsZaymwnXy7vOXMiI/6eX/msLvy8gxUbdGQ4OOllyAdLNYCt2dpeNO/
WnPjSP2uiWWtkKNNfOTPvA3BkDinjg6fPV22diHRsxQ7rTqvb3EzWF4CUGO4bE5+qouiFZ9dYDGQ
A7UD373aoclmk/RNbIkRwdJgY2uVuWFMw/uBr1QLnsPv828YTLykPyj2WKRJ62oBt4DK0Wf+pV29
j0yXXGPKNPjND+UHlEjMCYPdxWKlR0ZTWLCyxGbvr8ycixkkBJkLA7M4oBEPRWyc6I0GFI230niu
jQL/Uy+4f+Xp0neuZcXHtRFIcY65+1ZJWH2gQEune9tHjBW8O55rJRQGOtyk9yK9TVPhiwVNEdjW
iQmO56yLEbXbnoLw3Eo/YEWl/rhi78uriWGvyeKQjZBPGe2ZhChWgFRD12eePzJGXLKBUSxa8pGi
vVbE/NDIwaLSanoPqDXdqPbGpv1WaiM4wlDITo7t+TTdDMKwsmlhYbDspEcFT0hrTeJ4J4HWLFkR
PmW54CYbDMxKYg1jm5CkyQAqCtoBRpRt6ADB5aIcqtos/pD7YfTZ3Mp6BI9KqCnTPXuHyin9NJny
pcZG7Ne2HQ4zLZyHICF85nhcYzAU34OeXDomVmEArKHSJycae8QshgA0ukciFPtGjXnLcxfRT6dT
b2yC2Py6UXZtEUO8UvLgUPpFouO89LpHrA5tPl8LVsL9sFrnTcahbMOTEOq+b/BtXaZ7jT0dk7ii
G3DLnCL8Z2GVbf7Pw9+ZsJxoiv9NRLeYhp1WNIw+tS25y2TJ04Zx34N840Eg7rg9t2zGFSPrJ3Ro
2+S0+qnNHwFPCoqGAk65uoQxQ0uk1GzPxdl/HCp2pqJA4RSkvgL84SkX5mr1xwLNdTXXglwIFf6h
02fwqDz1lbX8gPferjrhWeL9TbH5wxiBpxvScbwcD1CaIqaByoOvTMwtZritKjXehVSaONWxdfZI
ge2AUI4j1T7hvRCp/z7QWoCGbTZQLJk8zgFnUlA7YlRxhPqntH9beNQcBnE9r4Y/mJHheNG6Apn+
PMRuwmE5vf17GlY93TIte883qzhqaiIQfqkZNuHkMPSXr/lsRfSf/FxD5zG5igWulA/k9VZA+T4g
0WJ+QCjBYsBhnLWjT/Q4wkIr8CQd5TTxCrTVM0NRD2AJgv8Gg9GuAwIGAW+6iutpqCk69KymxeKU
KE2WqFuEoBm8TMFOf+JQI5ph1T5od0bb9xi8oP+A3AvHoUtUuhtDXblUYmJiRav+CQ/T7CwJZGL+
vda8rOQ2NsHvKU08UVltszawLnun7IIGC4JdSJgfaoQjHuA3+nr5gBwIq88ubOGT234WHMASeBtz
aGDp8B/HaDhaKoFg+Y4FRxqGPQ7sH6IpV7JfoLT2+5CNRrNdhvtTAw1T26IbMIyLBPBKxbKLUhso
7/ClSDV9H3454ACz1/AGEW2qYMjFMO/ED5D42dlbuF1kg28p7bPPRPKrbRQa9ZV7h+so6FUicnOp
+Z7Go89oandrUcwJBrlyi24usgLZUMpToS8xnOVLzl9S4jRtXbBcKCiosr4neoFQWE/6DOTuvDm/
9QaUf1NQ2aMJqe80spCuS6clN/c8gbKVWH/5Eumf5DtIXRwjdx3hK2TdXGz6V2spcJVM5AmJGT4P
HX7xAVgHbwrx4v9EQ8rrgXWQ2LLRTUkNmk1wqb4r4dc/lj+IjA/AlrPenyaZNRE4YU8ReoxlJOgO
1LcVCbBQaLYdYcV6RzDIzLTzMjJjLS3bfRmdAnbmAJVY3wyIXAiM0gfhviqk7B0yBIadz2FK0o0Y
mES5PiyXChwyPOsxHgxUPs2r5aMPKvgS9SbG6e6bTUe6Yz4Kp9j+qIFjvXqz8P1A/Mdj0JeMmxwR
JPVZdMr1dl+LSZeX3e8NVUwu+wVX6bWXLZ2+asZBX5K59/XTnLnwNapzPlKez/x4QA8u5zZHhdnp
jy5ECMxYfHQ7O3hrwanO99r4lLEr9pDZr+CLUuWZmHCnWNcSatP+AnUuTPSf60AY8wAvMuveJflo
RX8cfOFf9xFKzJ7Am50oIQI6mJ/cd9GZW1WQzvHpALBZ1PJxCNOoYnq/grVBkzyO1qGO+sgksEsC
mcmzhI+M19uTZUheoT7tqZPaj6391HaFOdpLDakxNgFRnawuMBXtgQgx4QD+8ifb2EIDteAluUO8
JN3H7jaLNMslbSz20yT/aluBtORfH6ufpJ5J/Qce0As2Svbppkc3sfqVS+r1FIcSbP6RxBXTy3re
RUGdulpuLWH8e65hqfQRY0ZnkN8wVNeNWFpPTNdxaUKcyOBsjWlev4ysHPe6bYeW0d9mGZOoDuFu
RXdgf5qr6bADwkBS8oCD4fGNDa/h37rTl+VvINfiCVor+OHYpPYwxBd68VrCxfgb0ZBIFarzIRKi
n1gUUdy4dKk0Sq4mtqI/j22x6eNdX2LcU4n0raByim/G8DYq5k/YOKWbVGl6aSBF30MAGLiWM6Ut
ZOM7KlDCqDWKralBA1FvLjJ7VgBWT5w7Ij4cOj/KXcn/50Y1p+su9XIOB1HrTPoqU+x3l6RTMTWa
kTeTlnaXCFgIHtEFUqONn7qq4YrXPIzZ/qZVWp2Fzi9p4CSHblYlGPqpCxN1g4Z9jrD2M2pO6ac/
1A+N27gN1Blr23CD9g/A0Ebnw+pm6Uf1l+7WP6arePDNBVp7PfeYE99J2AT6G+HbHBbYRvIfZLr0
sm5/qfSr9Iusg2Ygq1UlffoRjjmyNhpXBjScX9h1uE9x1vC1cAGYYjdCNWpgxpASxeHgpHmE+D1J
K959RJCmoWQSr6UcwxSHHG3/WMRl04baJpt9MUzIfuHd1P2CDnxLvQNvCIU7am+ad0rnbOMtb5pS
2DfdQZuKdMO/ka3/k2crhyY9XQIbPvTFBjp1T0tVUDQ2fL89Xi7MKCyTNlmuepBTw/6t1kpffg5n
PGjPnZ7xy5WV1QJ8VnD+z+syhbd6s4La4CnjoVAE3HCWM7zLQAnlFqWXymrtqCYRLmGQFlv+hv8g
XtQdf+xxGVFMAcz6YEADw35jNKkj0musPkxCs52/8/MfM4+495JvOpukO43wUmEFpjgb/ELr5t1A
AhoWc7qL+RaUTMfiDWSKBCCD3xbULw5l42BdD+KUzuUcFiRZ9cXxhMQ1hEMlASvall3/yIJ636sE
fKLdmj1uC1S2EjUh7dxiyKTcWEfNj8I9echV376S6UFyknwmIV/zbFzyocIgFKUV3e5po3Yp1a+h
VpqYsagfRlcudJIcQSQwMqp1VpvpJ/ElsYhLWmhGMevqHhtc//erqPUUmFb4sBgPAsEp0iWU5JZX
tMe+4CPVIYFMH35ySCoRziWokKDZu2G8rVWfwWpdQl7whPKHHGK8tOmyRgBUQWMAh/tHmqBSHZuD
8zrz21q3zXi+FM7T5+QgJR9uKsZqjEUQJfqVxv7Yq8b1QTw/DrxmAmr5GVnwsiUZpwmxFEm+tN1y
uzLMzuplQQ1KZwAZjYhJuPPtqnu0Hk6fgZRvIJSuW20XwLxIFkuqR251+4yBAtgOGJNu7vUa0ijX
kGYimfsujNVMDj0fNof0VIaUY7KITLotiv2UoubXbSf+otILy1LsUJ893yui5r2J4hxoq85w3Bx5
deB/4F8VUJuFIxZP7+OjlQAFQgmBYCTPEIcx+BRln15sovwA3YT34Z0TvxmsHWPluO9AOl/5vzSM
Bjc+NmCXjXDSLPJjvBXJtbZFYLyeJqOc03NpLuI4XFG/1ozD2wjSHqpNg1HyNcw1jAsQ2Ou4M5qG
oQDZFxTzOC1Vm1Hi5oXTuIOC92210MZuKVHzR0cjlagn/d/IJl7SsPq6+th9KJlefrUtin3aShBS
CSjTnYz986+7rzDDGhAV9kPXxvtfhmDV6vOArPjFXONBuM6fSF+Jh8Fo0UCk9r13WSi8cGFD3fs9
dx1HRVTavupr6042qy7DfhCMkKhAX7yjmQH5K4J4v2xJYpm1/kuYA/3HVDs/tjGLDXzTpVE0cn9X
hyLodhjpOp2KmfMgcu+euOmfvAqKJ+Mp7h03eLP+qBdZNHpCCHvpvsuIhJmd+5CKMo1yWJGOirEB
X1W4TKfJ1WD9uGnrAnNDRIPZhI7l3LdSzkuWAUjbtW4/A3CAc3Z6OnjcD1xw5MsEnm9zHaw0KfKy
Q+UjfqWMZg5ac33jGO4ztFmAYr0jbGtlL6FwPDkRHjjHfejQLJRjACFpVWuyS7ruggqj8rmz9u1D
fjr8xOSwMWVfqTdFdzVk4D0b3ak8CsMuJBDd8BXZfDePAbDxGV/UtVKhWwPSga5dLVHxCo9y+CDZ
LNIuVJSPbn4+RysE6vpIagS1gS5e9HYLR73lYfhzXWIk9w/3DICwpDvmh1rVJmfc7Rzlk54lMRQN
owtoaKlCtgFrn9TWgcKedRU1dyyxwNmBzs+QG9uq9/SZAfvSNaivIRQ3j2li7NJkDs1Eyhij5gl5
Vhp7D17SUl6APGdHKrE99gcL4GD5smeVFYDWT1smPyBAsh8DVINU30RCx2hZFmrii+ubLBkcZyHJ
wvLW5H6TgDfhwrv44/ge8fO5bZjHBdXJvQbjCot+Offb6lYtoD0IufnQqlWY7DlwC2bfNfFvtecV
oWprXbS69RB4pbJyy7+1QRyPAUcJ1DkFEr21t01EoMl/dswR1RqhMOTi3tYCa9kWzRLJ1OnFuFu4
Edn0MDuQeWG1tLf5CjO5n724GtUN4RzIbR6eySryKeDsmEh+TyHbl46DiPyING8T64trBspsJh3J
MWws33z+HrnYbKnJeeDR/JxVI95jXeFf2R72XrHlNAiRFQObpGZhXmAQwp/hJABIiwc05cNjmS29
t1WBRtLko9ikjG9Lg+MshUf+ghqgJa5PELuwmzaU2hX+m9sHw7+9QwBzcGlK1EzNdIsRDsfPKf25
m5heaTX+77asWld5BdPb7+cLF0YjEZZ6D+rNPkq+E8bWd9Lc3AenCp5iia3sOwojkAbNq3ZtuUuS
QYSLwaRXa2ozoBGMub9nGfyMTG0pnPPAX6dzzGqeg8DVME2Od3SJqyAnQ2kwUD8Rfz2r3XfMHWop
L1FrxyUuAQ68IOL1TbJlRZTOkI9aa7UM04eg2YYT+sYV13cb78Qwq1ABvdR/HzxSPKQAfJGzid0r
lZm0iOrQ9O/AlntpWpc5leDE7UbDMAMfOuSijyZ50S6hAp5Juch/AoO/ZauKzQiivjdl1IciXm7W
vKsJ6MmSy6dWBkEZ7vJoSqppNzVzB60lt182v9rgrN4KBrg7MPZlzdtVGLAVecdO9xnwM6D6LGR5
xbdAla/qRbN2uNJK0pBuCX6ba1CZ2eLBuja9lJQoHHzj+KOsivSlJoWDtdP6ZdeERI+Uw5qvFc+E
yw+Bb1ajNv+tJFQlSzFp2Eh164sKXxVjFm8TbNGzcwFWQDhkGlW3Y9Y/oaoSTqWYqG+ak8hcrjFf
RaEYc8wVoXZMCsRRPXIPRpgE1N4urapY7oWHT7297F7YUm48aR7usclb1dYsPmCWIUSIFyHq3YsA
wuYsLjIvCsI5XBfNrt7TRnydWNIISp9CajbWBpP17okdyc0cxk/HJbg/C2i9yOG2Xg45AYiW5n1w
mLfdZ9GoTRz1LL5rhKRt2K+vtsQhXJnU548R+JORJBKsmWuDubihfWdYRKsw7EivA2bIfviDhvz1
KSmRcdPmDPvc3R7XOJTI0pABj1UtyT1Pe82A2bnPp9ehFbxykCa3HxwIVZ9HJ0rV/U6irG43GeL1
v0ZPLjgoYnpMaRKRCpdT2INCdDGYpCKGkb/qA/pQLi8fhcD3jd6C+2+FMPW6RvxhcDh+imHoJw8R
kTZ/jppn1ZyBC4e9r8eIZS5suoRvzlqBgQB4oxryaLuGJ11ssGXTDhhe1X3IwScBKOYpmr942Y/2
mEUBFa1YGuZhU+BW0JsIoNSF17psLHoXyOYCKPBa2R61/qjp3r0G6pxd3sKu2FQdaVAvdFcXJ7nu
1q2pnX17B9IrT7mqolkFxuOnE8zIA+3TwoxmNy7aKakjosQVg3TJuRnp3F9gM3eX0soT8WMmSF1p
kgzpwXyNG2HwLra3TK31FyR8MCC+PlZUbMQY6HEVOf/UeR1gW6gPybsk3YBtv2zq00zfSOwm+Vqe
Tm4W+2lJCv9GsM6A9Ai6chx212Qh++a/TmNOoN1qTfevk/ylYoOuHoy/PWC/NPLwuXTqwDsUlBF/
z24yGX2IcxODRue1TYDSbHirRQe/WNdy4JSW8klc+TL8/toeOLEItOm5fFpjix8YQtrugx8N3C6P
yuWUFFIpQPj9S7Z7rD6t7KSA6h1dx+NrX1aeriEyFtFNXW2has5ldWiVtzR0+GVVD0om6A+W253h
/1s6Q8+S9Rp+E1slkjo2h8VmtvfxgisGkPMXeD0u7lv81XqmbMIl3O4oyjS1UUNRGh0M0q+Fip3R
p4Ksr0XWuVnbaatz1BhLti148aOBgHOhgWT8vKWFDHttcXmOHJBcto4PthlD23E28EApaHc/5D3o
ekRp9EWQG1mFGc+9FaKcvF4pegLXcZtwlz9AAs8T2Q7GZ+5t13sfaHWzyLW6LnkhS3jAkGSfX/KC
4rifbKgQtf0LhIsldy6PZonmzQGefDO787Nzcjw1/0L05B34MRGiO0ZuBWVhVa0nhy1KACxS0E6r
/1JJ1AL6HiH758b18PYc1+mVPCGMEsK8t/FbTNq5/qOSfbd4Cct/cmO3kW+JgaFAmQL3I44iOIhH
cXPAz8vTwvlcUlb1JTva5k2vw5IItmI72xcR1bt8c53nApYpp30CEaMpdDAuA8FCi0mFLDnJ9cAx
D6w8eqdTQ6vIImDCsv2UWEENmPFvyM7cUwKC2gRmp4gfSq8gL8ddnQGMsIfxhYbMurE8t3Hf6X6s
+F2LWh37UTID7nJZ7+cWfzrhsC+Bekwi0PBUzk64y8pC8yoORLxQhVw8KJFLV98/F+dTa08yBNbq
DE4CXh5tuHcUlrZC+Dm7vBtyeUldD5gu1ZL5uSYNGgATanEJSDEISneSlwrRa37Qs4e/T2fFyPeS
kBRfrnoSiNVAjE0HjwXFzsBlPrvEM8C0/xlLr2ko17fy02DHVewq0sIgtMZ+DhE0NmHr+VExA3sa
CKmN1Ljbw2CCqaNIlUuZ5P4Pw7SiWLoactg37miSfVeNBqr/qGZEc0NW69EYLPFkhqcHRjyyDmyU
N0Q9xdRkDyRumfWEkWDm5e/qijVLJGRnnQKr5f+l3tIyZLyrprkrAMJn6pQsM1SiGi6KbbRG5081
yv27iJufeVhl9D/kmvncGiPpjVcU13V9GOSGXvu03xAc+lqxg0dqKm32llU+TkLsthsNJJ9YtC/L
evZ/Tfbfba3RNAGE/z95r4CoWUO6LFDrenkOxhyWQNgtJKndiGar7tHsOWL8I2h+dnPAOMPVAKV5
KxID1JKJR+ve27Uyx2FBLW/f6CZoVvE3+v/gS8AhXZ6ZKiEKZUm97eL8NZCnWMKARjQ5/AXbvxDP
EaPL7clkiVd9nBXkakO97KL5fXn7Q37TMFb3EhIcUnOTH3E+F/mS+DpZAoU4ePbnu1bVaU7hG8Fe
ghsmoBDaSWRGEcB9d8bCmT9t8s4DiIHjb56Hl6d9PA/qeylAcmbxH7KBTeG6W7w1clIOQVovzjGp
fddp+GMXWct9rHM5tyFw1G7yePSDA6AX6Dfc7stn9H4jSDEsJBJTggQf9Hs9bK/s/zf43UXOygBh
c3mPEFX0or/vBjA8w5Mah2x47g6pk2u0dByBRYNcsNwks4I1vRq3H0Xoq8jFpIzHSXHT8epi8yP3
oJLnP2MnXSpSWr8a4XkuQdLNR26NECx2QCb4gSmj28JkzsFfsFLaMpfD57dlAlA0iXGuyI6AFQUx
lsTn4Bd6GzIUFPplxRBBpvu5pxNhdpVMTdPHkO0/CT1yQaslDHhVTt5IUNEzBXFNW7O2tSEAeMwq
pqpjtZnD24gYRO72zwGFzIU7ENZs5fzMVpkSafzKnF+IjfNwG5yBTzI48ssJtI7n0yIpD4QHDH3D
4wjq+1CwG7EvXMjX6y6IccWgn+5om04YurinrX4csFUEZWuZkD6PTraARLHTsPlj/oluyimzPdsw
HIZIRWCxy6nzJZvYWNK009txMzTkjdr0Q4pF8008ieTQW5XvtsHaW3oFEnlCOozEOdmwz7BamAQo
tRTdipw1qBmW1YH0A1qXXCnDCdbUUap812+9OAhd4cRGz8jcVCFZSLyHh8zfI/73ngw5XxrA3a1K
o/vQd19tK+/ogw6fzu9s4DWP52Ax0+LX61PCE3tMizji8H7HzbuJGYDx+SIGm7OPHzT4Sc6sURbX
ZYs0WKcIOx5iylPPx4+bQi55g5nlmeGIWmy680ZysAmsFKf9hevy4kr4zFJ6hkaf65Rldppt7J1c
0W3QKKyYT3EZJ8llbOulpJcGC+FEtKZVq2gCCwCEcbsjYB8KfYobkaMCjMurKJ59nwibWW/ghGXp
CZyETucUS/OBdWg5KN3mlk46SrByt47P21TF/Vz11fqqAlGQfKraKyQ9qW+PJBhTdhx5lOmgiSTI
tS5Mym/A2cYrZMJNgr2DJx0otWGbTerHVJHqhAzdwYjdoOuyPqdYVoWLZxmnvh3hj1tdLVE83HN/
pcqSjBto4l2P6iYIlE9ntLQU5hxhY11OmA/Cy8NwWfHiprqYAGBFwEH2Lq7KMQEclHivBhfl9Lbt
gOwf9D6D/EaPmlRyQGx/535SJQPAI5808wQtTdd8uq9W5xLfIfQkYpNwIquTJnG9HIPFX4xmqii7
QnknJDlP47I9k9Nzi5stwDMmmLCCh7eGd1NI6IMsKw/6obW7SgEW795miSMuYFm2NOvnbSOq6x13
Jm7LTgA0GVMFPzbnowLr9G8wr9q6vcaqpYbFZdDHFd61bvT6igWzsPqreTDDkKAZPH8p37hBO5gN
e1SoQg3GRwymrLkWf1JIuuZPJ0sVAWxmlJvSfTIPQNVjNXvNgQqwraO0T5ez3y3D8sq5F8CodW6X
yPDwwpEqZdB9naKlVxSXZB1q6hOeICM5K26uahwb0iLjHpIsYGb0xwE3v8IshJG8sNVm5kapFPxW
EypCWQ/5q8TNbLG71at/eNE3DsHlHaWaFIOsh6047iRpIyCS53uLgId49sAqh/xBaTT9dDCfauRa
kM9pYFZZ9+OLV59oD6yhg/5x8RKOi9r56Vd4yJZCIW9ncCkmNedYRnLmPbxruT1vWD1z3JeJlR6y
XGi2rBsBjZCF2moE9EpjYCzov7LmJeNlYQs/R5UyBXSdSWsNvkngys1q78955bvoUnSV1LSJJS/u
CC1HNLYpg9oeU4NKlvDZt1JwtcoxYyQViQX5VmDZ8IAmCFY2wdR0pX4N2HGFZSduBiNeCXA2+zLN
VQYRDQ7sSjwnIdXBUmnsw/8UDel1WCt11wEAutX73kyrMnH1cN/ZJh1vnH6QGS/+0wX1woQk5k9W
byCGDHWh0OlC3Yae3/Uh5U+bWKfyTrDAvVwenXi52R/U8G1m4OiMQJ8kn/wvcNKAeQRxFHoTRiCs
hDclMGMNWP1zZXYEm4UDoEPBNt2iwVPwy65gk3w0XTdqFjOvXTjocusslr9pdVJJAuPMow8t+UYY
+blH4jzwRGzRp8IVRz3B5WH2h/8ewtCQ8/+JvPcYTXrV1Shsdfrx9wo4En5DdoAh6byXRyytxT4C
ekAiit42q2xYP7k0HosRSr47P0Sl9WWj81+xcjTIEJn0QAKP5ocdENOXw1VR+nvqDYzqxWtLldB/
MV/3+93aw3gKy3MJkQ13KAZ1OWod/8vpwillR3nazvrSbhv2dn33b6KAiegRVejGasgqp8+7PFuH
W7hVVfSLv14+gUxnrLP9Y+Wxbpaga2CoOTE9dRfWRYRK9cr1Yi9JRQaGqh2K+toWASfL6gATsG4+
+0cn7DIG28aOQV6MI6MfYHYVO+xLthJ+C1VeHcIB4y8xA8+qvomDLm78GcD6DgaBjJoAlPU08mpW
Z8mryrCer12FG0Q5/NRhxGrlKo8as7B36f67zgoCv0iitRGnPJ+P5/2/Y6mbxH7fXoFNkr705hjJ
fAz7EnZE7BtAITvR01yDzyePgwoDYY3RQZF48JQYOly9t7qstR0JEAffSThCbFwWfEzFYGZ92J1J
Ar/j/5+RAdf5q9+1W0wfrg5HTG7EVGwXTmj+H5CDZdh+A9hu2ECDLz9treYMHHi5nozfKXb8tAsy
fuiiL9iOOKPwb65LXGuzbAEyGNRZFbfRoAA1MFiR9NHb0oxBAfMjNgI8OwqxfitgBPuzJQMA2vXW
mWbwf0bP616ZbS6Nz5HD3ykCM9Gfi7BEeUxPbNkYOAVSSHsm7kdXvWvA8ohXfYC5rgkJive1le4x
9U3RrWSmfnhwWv853stVGX+USh0RzF7c0LbFDFf+9pLhaTXo3v7uH5b+SQIyjPJpD1XuiWHfZ87x
g7Zi9n+3mCyauNWf9UfBD0Tj5D68hKCZSw8H39Y9Y/kc7XRoEA3dhK6jciBF3+4mRi1sCxNX7uBi
tj+Gf/ANNMKYd+Vg7I5jMI6zzC3DAGVtQu8c3pGBd7AnPzABvlknWe52gQ8NL7NXtL+DIpOM4xBz
+hWqG38Sz61pOek1shRctcGhfxmGInF5IBJeh/Qt8DqMjlhmM23QYvjp/9rQkIs/MAd21V1lGGnU
feGBs5c/XAfrqdnhO8ey3XKPUQXAyMIfSw1Hr2fW1AqPXAsxQN26QYCrmW2YTO1g3Nl8V+HMHDb0
DZDWc4fnAlAduHc15Q0MxNDgM48lwbyEHviFn4bd6ntCav0XaiIgN1JsWaXe28kseCh5/nuQym87
8xc0LTMwWiWl9meVh2jCNLHD3IPp/ChQSEpqy0+1ki0/+waUVhmF4ze99iIvIfFkt35bpEEqKXAZ
Ti30ZmqG7LrLhITWcvzv+cy242UOqSy+cIZyMSqVbq5q6KpCdxn2DLPszuFpthN2i3gkb1ODngjv
y5tj4kdcH0rsfObRX/PQSVw2rhkhC+CfTCbP2ep5kZrlSsOqD5e932lpZqtKJPXbBNWOgyuitGk0
oJtlE3rJxWBo+Sqb95Vp5HhOuil0z0jti22FdUEI+HTxoVUzG6ua6dtXE7oEaS5jnLTCL8osmNwd
ok5pl9wzCssyso3NDnUgL7j2TEYT4HHzkE6wFaAU79fIzKNRS92IKSLoMAWvKSNafgWPykDz5j5+
xnr4HggQIuu/1A4EZsIHgMPCWBynfiT2LlbGaf/Aq3T8q0HXOPz9FSKC+tBJbZu/pcJ+287HwWCs
lc3cQorgp1Ugzp2/pqDsDzlnac+fkwtvInWPZ0UHTpRlOf/LqceHrk4HDVvOt4fRRZJBUKOUdrzP
3GC9g3ejAGBkAVUFC1tkL2dW+NUNP79Jwc/fdqRVSQMfo/TmwJ0N/63g2fVxr+w4hxQr8RYMMB/R
c7JGo9uXoFlqRnvPhqPPYiCV949p2h98Gj0c68wvL0YqVa/KH3gzJV+FAX4tHNieDWafP/pGUS+u
xFmJBwEKtBNz0KMgfSiL5NP58XeXYqWEwJF59xFqoAAYnV17AvxEx7NPPxn8kWyiY6PWu/o1UGXZ
Bf+mpG0EG+K/TmnIckDIRjw11Hn1LhvIR1YoYaTieeTbETM0XYX3u1clH13zSl3/u1jsQ7AUdypp
M8SLL6oSHdftoeXPeTFAnKdR99Kn4X3gMAxALN6XquQX8xBNQ6HtAhOozKIKaFaRntAiJhTwHOnv
yzaaSQxOn0b+m2Gt3hPqxh8OK6KO3Iit8mWrv4WYcwgMWGPm1ssGClovpRCOAsYczm8WMkfUv1V6
iPojENQXT7JYDOy0cHgJZMS4cRGBy2c6BA2hHhf1alZ1KrTzkzPsf10krY6tU9KV62q8D9EN4LfW
GPVcDyTw+iYG4FMv0vQ0whLrSyVCQEK7qxFrRz3Uaen54ejWQ0LOsz/Ys+adKv+/5yhDILBrXlXq
H4IeJP12s52vHWi7kbJMkS1xKv3BzdgingMeRh7kie2tic7rvqwmhEMjlQgebRYqhNp9tV6ymBt+
buwAWbgm1jnkQorjONr49g8+YCtqmUMw7Anx+aKRRRtHIzRWqf3KxxhbPetggFgM/T+iTEnI22AS
52NOGGzHTMhn2HHQD/iRyeWwyQsAXbgyU2qhGX/H/YPKAjwfnmNWbnHnAUAsxvABimbXbGH40gPU
rQJQc+ckyV5j9dnbcJIaJ4W8smof9YF1Le2BAnfZaQ+nuntPBlxaOfZrhpxKpfj9b+zDSlT9Ka0r
cdEok27cPvSQDdwfNgWEdxcZbgNiMUz7Ytz0Wvj7a/YQkkvVXeQOktmMajIDJWu34lxhQ8a/Gccy
jNESUoJfEJw5S50WiQfCnJRVKXWLRYSJfvvY8XvgsqX7lITCwRmhdlmvvsyda/dxVfQYEe+gqVKG
Nj9VWtog5QU7b6VceGwa0VssmcTt8NDNDTWKVlbykjElWJXdYXb93oJ3Rl3IIz3P5q4VIvmV/1lr
LMrW/pBrYAvZtWEfTrAK0QHNwJfeVkh9JfKjvPcUZEJO86vwIBQFnUKmCAO3XkhL2fTardY6kOSC
dgMpehIEJSyL7K2xSgGe10dxBaUsBrSXzA0scJSpEFtU1UXQe+Mp4NSebN4QH/JpEBNEaqd1jmHb
O1jYbbNiORpYPKEksSwP4kqpQlCZZTJp8SPv5IRiKmjSyzCVXapSz7YrubIuP0jzfNZtbTlOi7mW
AqfIgX8/geBU7LfhIX2VLdgz4wxEaIgVuVnboEDZ7rC2Fx7HjAdnOWUOoFeqIeKRzoopbceYVvY9
B80z5rt/qDBigVuvdKxXMd7XQtcel1qN8ODJbsLIaE2a77ZuO4KxZ9nAORE50l7zCyoB5SJ7nkzQ
K/D6ynHRywJqhN5zd7ILyt7DH7cT5K4rkpG6sCM3b9nclAOBIp8oXyztM67tiWL31rZb+pPuqb7h
AtykzzQjg0N+j4bRWUua/UEP8fgjjQF4n1LJwUXhc3AFB3v/ypy42yNbeVJuUuEExQu3cCDYEt7I
U2Te8VakZ2pesxige831LUnlFhvaQjuDtBIt8Zklq2Rd6C5NYODaHvMGGaTdmhI4jNLn8Hp91nlZ
YohRGdMgKgtHASS+wYwXTPro9FOt07GuFaX5C8oROit/nsa5ae4KM4ar0n4YNViNgzQe2LjD016E
uHN5h0DAHRV+FvuFeriSVpBwWGO3Rpqn7jz4yCWXeGZt3FyQXBrq6d0Dt1lnuXsXjLRPiMtadpHN
yQg0PlFx2KivzjZhrSUckbxc3sTPGJEMOx1/0c6ks2DXVtffOwgxD247nXaIINFHnV6SvSRCvizk
gEG7xLxLoENpxhgp5mHiDcDLEBjboP5UeRyBOiDjdBGW9cf+95hZW9ubIjpefzdqLl/0FmCyS4EF
a6rHWORV7JrOjyyZ/oFZZdcD1NUHtMX/cXptdNSf+nTT8M85j6cB3+fXTiTjURrk6tQ5YH6D42nM
QX0K501ev45uP4+/r6VQHJ9Nfwkd1baYjFSytFg+rm2jioG/4CJ4TwMge3RtYywoHMPORPq8zNyw
ODsgxlfvT1eyyvzYRY3k9z6SQIRLEt9Fsqs8+RhOM35FusHFANoyfkK2yjtaBKEswu2CwoDyQfxJ
H1NkClwpxmbfppn3JqdD9OKhIrgglWmLtejw10//pjNcFOGhT5y+9rMOEDGPzzfv4yV3YXwkk6QD
mg3GyVfJZuiXW2NmVeo01ZDICchu5ti1Hrjy9X1C3tStQpeJ/u5CdFf9AhXuvs/HRHTAJCqGVq72
+6nsQt9w1LS1ii31kqvqA2Sf3J5lWpzh4+r8ptO6fprp0xIsOWQrRAoJ3ncX73+udAlJKuZbmMKd
eyoxp+HaxvHd49NgWEBwz+RaeZAg8pdWfmMkd4S1l6H5Y7WnCKZzy+RVS5Htrh22Gn4ZZDN24ASV
PEU3MaIdbjIjIIMf/+MjHpsjV2refAuPWm+Y0+UOjLhbh3yV8Idrievz3J3hsx1AQq9LfAXc4oth
IJUjKL76obX1BjOR1TvoSfNYeHxy1+qJb7U51J1wCnkKzrr7WHFnIlUKqYAsQ8Ax2zmjjiXZByon
uaDlsCfbu2TUC5R8/FwtWoMvYZ4d9P4wVMg0Txx11KvpiRjTA+zBqhR4QWvxLHXRMR6qUCOKOL+H
/UIdJZh7/JlexzxtN1PIhxznGbU39tzZonrtEkiPutefK/BvswGQ9pLiVwyX4IIw/PTbV6xEDnH7
0eITwcqs3xlJuX3O+hdeOAlv0ySv4Bjp/oCHx5NKptrIRbK0BS/bO/5x9Dw+WdKwwhBgdsHstgDe
qanUZq93D2ili6g5Ck9/wVi+JZkzr6+B/A8scUHVF9bU1V2M4x6tNfvJYKVSdjFdBiM8RbyLm4bj
095cGAx7HfwH6mNH4Yfr0K2s8KYatB7n+7qNXRyMCacHBnqMs7leTEfXyc+MCs1Hrp9xL+sICstT
wJ3qPpdRzxqEGlc2d/FtqwVNZQNUO7cyI7203oKS5CwtMuDhvh0pBKDuoQMYE4//8pE20xA5/lCd
+bkexduK9FmpKyJuGWyjhhLpha727nngDiYmk5D2g6Q10lv2LbjLKnyGJL/S/MaXoPDdbUB0jPLA
u1iErEGkuMugZhJJhDaMIObohJJr7lqnLRFA3kMOxhGe+WUy6yrVT1AYszxAC7vVB+FQUy0bG7BF
dYZ8eobilGIMKl80JgCikyiUwhokZoYZn26B1MoJ2MfaMjr0shE9tvff2Ho2pbTh1FJHcD/kerFC
FefJJ6fUoleNytBdfpVqxRFTIJW0QO8FPDqMhZEtgaAeVx6Qf40Vu7ZSsJkyvx0QUNp0GLD4ZWrX
VuBhCXTH0z6JzPoasMkukbx7ylDJ+ndMC263aXzuDM6E1A0zyE+1erLFD2GL/d70Te0+sw5w0LLe
kGI5HHW04VfBthvErlfSaMA+XuDzJRgENDnzqdnfezFRuL++knJ5BEL+maNy47fJhFjwneQWvjFi
e0ulolwq2TbGs8bMDRvUEOjxbSl1f7pYMByBzqMwzU+tqpaAMVGOocIsHdP70tPWZvXE8iNI/lmD
/IMsKu8SJeagP9QSmfwcZGELej5VnVSxZ6AW0TUc4C2GVlnsOXz4w8vzSzEyvyK/IfQTIYMTT19W
f8m3bNMNXPj8RFXUAUs1qTKtwVfZO1yDswckQ891u8vpCzgIp634OkcFCJzu+Tz2scnl3Y5NGnlc
QT9bxvh8hCkyZVbhc8cH3i7ri73idh1PY6pPxT1pRuZfRqvlVgCkSxEMGgLu8wjBhSuZse18pDlI
cGZ1GAmRR29gPjTOFA6p3yAqNaVf2cg5sLqDWDTrzWTXR5MbbLVU2a19VV94A5fzH3o9nNES6GId
skFRiGzi7FSjXuRZIqUTBniRjp/RKXgnRTAYK+s9JuWHTT/q0iUudLtz9UIuephkYzyOx2xQLbCE
zyXw1OM9DAGahTmw2FTd14bECDRk6EBQI+krF+UBZSaotMm+37wgm4Q+bdKDza4mhiUg9se03QUM
2P9/JGAHxEVfNeD3nRJOBCE13GkBYnAqYWVcKia9WWY/ZMhAzDeJmhWkJqHzzB/r3VypYSnXb1LB
qxR8nPOlzP1IJR9Wl9XH5/DIoCh0GEtIv+PGNulSycYQCRxdIyXvQ3VrIbBicdt+FWNuuIo5z+Q6
k+8Dcd6VOoPpTNwYvy8OFnUvT3sUsTaHz1AFd4W9+b6x7oH1Bmae+SyTq0lEhS8US8uUwfc1Suvc
EQAVDAJk2YGm7FpKWE7fKzpgflYolmt/AMON3a/YJsgu3aStD4kI74q7OzNPo2XytXc9oJVAimNM
Gf7de47Y1iNLW0rU8kXQUffQwOoZvdLzAKxlc4HkTIfcAyYsvemEgRHxhtKaRWRxgrMX4XfQ21OO
XJFE76Dt0pvb/8hrDWQDUUOInq5WIgnYIRQp9k6HOL5Kn6tLaEnj3Hp99xIehLTCH+t0iGqVdwM2
Rgpqj1G8fsZB0ZIQY5Iq9rNJeQk176AEwJ9fHbVfzojr5MeGrxYxBzbV4Gp+usPwna9bfJDYQToI
pgQwArtNA3w8XhuEpwTOGSRkWnXlqZlvuOfpaSrjtzqgmaUiBOICEwTX29Fs6X2IEcvNA7/dX8n5
tJ9vHwaSWafhScFzJrpWtHmvoD0W3yZfdWucJj5qBt8fyilnYMXruuhLp+ob3gAH3AfCOwktMX9q
RJ4advBnq25Wqoy2+hLDtsiecL2Cwk8J/YNwr3pGNvxTY5q/ViTpl0eBP/E5Gj0kg+xSNa1gHi2h
7+imTV9qQXkZNXyaAOMQodtSTCRuARNVHM4DshhOHcfKKuEt8+82CMokp7wpKsgaiyofi9pNFky/
+Z1xA8JfRf/mS9yZ0PpgNRUW7sUTJ7XpJRonpih0AHSkkUI9r03kl6hHEDeeQZ6Iz3Hl7Dl4vi70
jMoaIPWjcENZh08rx2UuyfzHpT3bETyhN6BlDHxW/EvNGrHUdoT0L2ZKjFt47GgF3SQ94Gk33GRO
nkle9FoeDxzU3yiiHAs7FaPZVkrhZxGxii9/hyvXyLSRpJarwserJAshsElTeS9H05c5TJfedeqM
wJunMGyPvZSasIrKXrFy7meNjZfKX8VaQhrNaRW2YI/7qTjY3v8HVxWLkKuoqt7CMQo2CoYm2Pk2
23ZsJ+A5wVP1KBtgI/B+KGKdJblPPpb1nJclCrItvnoFzRwWQxttb6AmEqMKawVooVQyCSQOeFrn
UUkPH6Qj3XU0ZLKedCuHPRGEr1ViPUII51oepBst1Dazgc3thYBMDsBhrUYdzEB4A0o19vYY+ka5
NYIenkdqlYBG2Nfh/7Zxyo8m9K8MRgo4jO57APwsaLGQb4yuYmCAo1EDAObSKsx0dcRmxhQ+1cvI
PunOylzBQy2KWsz68CE6I9L+2zYcTWvLqRNRUt0ScUXhqfWq5jELuGfdi5I3YYp54S8k7tBGE2n/
Or9xx/zpJ5kKNDJ6T7k4E2rvtuRfPNFE1E5yYZbqpTJgYLPh3QhaPnvx5Mcg70NweUXvkPO9dNb3
zdqEHfVdKTfwx6/1lcO+y/0m/iBmoVDkywM8NkFhxR/3fEojHk8mdML8oRrSd6vKJfeTq4oxUVNt
aSW3UOlJTSH6Db391lgFaoNun9OTsfpG5GOXD36yYR9C0+BzrzDiQWBnEf5ONtebQHgjA7h6Jk9m
wuk5fvazxs5wVDmG2SYnlk0nAF/QxRRxJHXzH2FRq91rq085x1GbzHLUPgw6nZsNTjOu5XyI4Mz2
hC1jW14Ah6AUxwih7HmjdwYWAbK/94d33h/fiFQTsH5VNUdLmXViOp+/I67KUqfEKPD4qU8PfI74
lncvuQ6qm4KubIB10Pci6q109YKfyvpDzHdq+xxY1YRWYZpnU9Uuhv2T8tQMBUbWZzPVr8MKYNlM
Z0xe74zD84Ej0bSebyMvFuMEfYgMRVc4t3GDdaD2I3F+zuhhOR57juW+9PPurrz9dGr95XRqJmqn
pp1QiPZYi+ebVLAobHt4niM2c2nlC7zlrLmkhryAq+WV+kL2efa8QL9BsNI3t2RFIFyQJW8wpEEl
SDvmgck8amiW7ZgHV9MFfc9joYkdo+Cvo05QT6rboyPBOBZ/5WPQ9jOA08DYSB2jKrgC6lQ8KKk6
NzKtKOxEa3VKLvyJED7s/EwRKt3n5/nyvRQaoACXwdsFeSJCqOG57VufqA45v3WgMsmIIqOtMdc+
qW12y5HDoR6jcAWhyUrKiYR6DjP98Y5VZ2RfFFXix3BEohsSA6itZah1j3Q+buxcL6GBcT/Z7Zd2
HQRn+4ukQ9rSwYsbhfsE1JehZtoziDMpek/KVwr/eYtDQ9Y7T69R0YXzqZ52TgU9u6nztqzAlUtX
j55TL7fs3xpAbhHqP1U3nOgWny2jStZ4cNM4d8YIAFP2d11UPyld31ktuaskhWIO8DadRB4gAErX
fqOhd83p4UV9r67DH+1B6lVltIjFQe9JfeinGF3zSXRcXJuVbDb4OmCiaMjPVxcdMpP+hl4yAPaU
cxuUO3euzTJYhHJHL4ZMqmAxGSe5eII/pSKjdLIUS52th5mxNa/INizw7sU5HIicE6YXcRtiKEUO
aP9xCcSlDEcMd7uXUQQt/JFpabsTRTS3pXAtK7zDBO6HsKqOrOZTHF7jlkI5vpE1ctnqGTA+fTfR
UuhfhzjAoyvTaQX9N5pJnEwEsuFpZkQF6aLbQkMhudboWOfY/i7poqhbR1arZ9YNfOOE82kzhoiD
1ewOGZUxlPMLUEBCpP/Wf9YMQV/G/0sv94b3R7aBfR/p6QiDKDWFjGbJroLKU1S4fyUbNRNLxtQG
XSk6p8PUF/vWqec+BahKhlXXQV9QH2FWKSUHeRZsJFoGlB56l0VJd0bOSZRswF1HqcuQP/zUMSK0
w4uRU31cOcCR73USjoTbHuypXpzNYmuxK9uBW++aoQ9V7y046Uqny1NDNQvK6LFeXCro61FbFccm
yn01EaBNlKxKrHkNC5YuU9/v2DD6i/S0YLjN0LlVHk0IyM0n3DXjYWJWtOUni16mN7tocF7Chcoa
QG9ZKbDW+JhOjbeK60mWsXtmKOIghv7QSu6NSaKYScnIiRJbjt2dtFcj0SdOFsukOYoOMFpMACZm
37oLWK1SYkSthpmMrTcEnssRSsEwhfdMvZdY3K/fLqrPdgsqAxtyRLJPNjYPQSWh83U+HiAOi1Tw
iyN9YarADY6lNjWXoLsz7kTct0zU5VkmLGXG24U8eqgR/M+Q51kjD52II5P5T+J1CFadncvgkgbd
abUofCXMBwm0lBzgJhgSKLv09U3nfkr8dC+orR09nU+Z2cRnLPOb/uIBcJBPGYTEzYubJPA5mEUR
OlMm4E1gv67wCVKbhUJQPkUHjj82zOLmqzsQZ/gyvq7E4Lt2lha3+3zbHnN9R+2VJ4hOMXTNnUiY
24hQ1OrbVw9AwJQdc160lZ4tVXO/xYFBbLIy7KIw6oyO0beuuoRycEU5KFO1X/OXMAop0bzG5Mfz
LsbSFBCNCUhbXd1nUJqqgZcQB5Mx3WStSHMG0KsYy0MuO88DHVSeXQ8r5UVotueUwm0CLB0BbYPr
NAE0BtGINOVEE9Cj+KDATx473z9EeMJj6C1D9eglVAJK+YZPY+3Qgr1fbtcncA5cS6jHH52lUVCp
iQRVun6w3aRBSPb7qKcIBJDDNHEp31dkVN4TbmsM8OZyIihPaki3CL6zc3SdCCK4Joal7ll09wN5
dLb8Ac9ntGH+0k3ezMCTUf+RntTjmcn34L31/SAqJ3Fi+6n0yWnpmI7CBwFIBbgcvCY2k1/hgQJl
GupdDd77YdT8/ZdEJpRbRuxSmVcNwUDnZud3W1N1MHXudpMOZeL6fHmbHLYzQO35eDKbSz9FW/Cx
9XeuGu2kIjgIasK9nEqF3MibyFIY1kgmOc2WHCARE9u8K/2hqSRsh5jUOL8I7h2TyFztcXdJR08w
96MpLwNOr1dALd2vSMLUsAwcwoMdi701XggtWAhdU19lbv6yr+bJ1UiIVIQfbwqC1NoQEHlnXL8Y
o+3+aVKrsmJ9578oKa1jXrnsybnna44gnHQj+albUtpJz37EOIes12LRNz7tU00BFBW5DfKrWMw6
lkCGMhGUjgbgAMuWXYIIk00ewY+EHamvgsgy3EsI7l5C+x5p2a6n3NT4SZuAiVUxiGNhoFpF7bj8
x1OpsZA+/liJdOgs2jjfKGvACzoANHl7VfOpRMLh851tL1O4dE5RpT7vtdvl72on/bIpIIAFmK+a
yKSuL57Yj6neCMbnbQ56ljiG+uEqbE7vst9QtJlM5KfWVIKnqrdsFOFPyJhX9+p0nj4xZqeBOiFT
XTyhbG5L83KTesYuVN5p1AW0nd/kBR8QAnB0MRElFfrEwv7lMZPA+pfBCaGvNsjd1ouSdQTlbm2S
UdXkP1MrS75DGNJfG2+AfB5voW1/AArsdM5jjQZOqUhj1ns51SjDqOID6Uk6bWoULgpVO0SOi9dS
OSV0wlb6F83NEV1oYSrkeXKgrriAxSxO+ON9vzB9ItGvPWUK78a7psuqgxjBUGdxHsCV2C9Raswx
cPgSK0+knRR5gzT4Lg6763mGFMwfpwbSZeRrj46U855olZ744h8xuc3yF4SsCCMcKA+uu3mocNQM
f5kbwWgQLAyAAQUzMI1pCzd3grqlRJ1djFid39K0lG+GIRkw6jPwTbWCA+w4UlLdoL04ckb+W5mJ
bgfuhOZVysnq2/ELoz0QKeygYRVR+WIOF2AQjhTUePL/5z4wxUqQbse1r0/uzer3M2mw4E+R8aS8
e0bQCNS2OLcXxp/JlHDWAjJCaCcKU8upNiSfRPc9/sJgU921VyEbTWhsV3QJjEYW/Vh/QVPacj9V
FKK64Z1SulmzqdEfuZOWAPJ8isBw/gVBV9C2FsqBaVr+eqAJYM1ZXX8KuA8U//nSm3L7GPYaHzct
nbKh1VvdOVLmy7s8lH4lbCEaSfdEjVueMizz3T/H43nv/r80ASognGY/WyhIGPSbjR+X/cztxGCT
UnFgiXXxS/rM7M4stFMI0b6qtTGwl0VZPaBYUwcdvRTh+3v5sILZKIg7+3GZZKEQoA88Q7Vcqpt4
YiEoGetrcp9LQqsk0i4ZJMiZWHZQIwoZxUNR2v0mbHiXT1A8ewVcyq0Z+JVSWCvqoZa97y6ljzl9
atrxrta/IU3bIoJeaVksvWSeUAZle93mfU2XgSHb99jbb6uQSY/UvBeGRLsk4A2mNYDgM9+GmpEa
F9jMAax1S7w8C4EXr6NK91XU5Be52/4XTjJcaGOqrAd20b65RAWv3P9rBEbQUppzKAgYwoOX++W0
WziBMNs9c8pkZC7Mgs1LYxkV/+GYl3vhwXYzngkBtlpG8jiLg0R5xdXOnN5opC8FKhHOh3Nc83y+
tx4ZpPaos0JtCCCi8eRYjn0n5zfncZ9fqTLTZ0bOG1rLm2DC9q15HMULigb7K6e554BEcgt5sYtT
rNmlNLNuhkYQvsrTh4INPUA8yTKxV8aN7fkoqbboWa3kV+f1IF8AEVmj5Ur6cZrAuQ9lNE5JEoCI
GLFa9s8XLWgOGSoL1n7pY7+/qzDd7LHVONAFO5I2vOT2sFZhX6jkORMtQf84h5SHYsygRrO9oZ3F
VijjyKRpSlx04J/5ISuk4/J9jiHTS4SJ7rjSW/nII3s3jE8aRv6PnIWiH2q8s5iTw8IyHrHFcHnS
CyuReCDgOZPUUHASCDBDZ88CJ/1Mz3AGeaf3O84eADnQo2vo6OiW6+o4+KAzI+t8wp25EiNfMOXK
fRGlVUMRPhqv+twZLqmGWRp5Tkk85456FetqLLpTX1l/ukSb4gn/jmhGMNRopXvZNTseuGBIdns1
XpBvF5Vh6DffkpC3gAAnBkxhWdRR0o2b49buoRt1Ycu4FKQWo4t/q/L2KJyrgigBigECuo24vNN9
b9DbG99qMb+WZN3eIrCVKIR75imRwNBmm+f6LTmC2CoF9Gu/ep2Tc4459OWoQ5DK777kBlPFhjQR
RtFSXVpFn1kDGCPuDL7Rzp1WnaxIWrXcxDeas9MljESGqwVisOg/VGLpJuUKa9ZwuH/rOjDTdAaP
xJeljiw8QHw0OMKXCsK6TSh+TlwdhzBuEqoG+YtsvmG8AdJLpwhLlsRas6NGtpZJbGS4glrDeTkS
OlolwEkGuhk1jfQ6tVlAf6kOlyd/JTZoz9h7CNvJvAHVmDQNb47dmIeFvuXe0v3aKYkyBvoMzRYD
MkjV/misZ/+ZSnEqHVg9jiuOlOHF4rWV004X4P+klGWF+85w0j84jUA0uOEhmj7WgkWf/h1wiMyx
JCeaTB3BTeTnDdjDZCAkjc0fg7e98DggxQkKeM22SWNbrvH/zFnd1q6ATQW6XOxpxI6IR7JiI0vt
o+giZLpGhSrT4edh50LXhR99czQZDIp5nwozqeS5AIE/QHlxC36/qAss+tYu8Uu2vFsblKwp4QU6
5fZE8i3tIOvtM2zizat3+4HBgqbggDUc5K8Ih4NDieb5JOPbEU80fozmu+sbw8OqyLlA5jDj950o
BHjW5rll3YQKAnh2UyCBYQkwz3cp3wASGo3DXE3qWgvccpNLmAFU2YGXdbkzENAE0NZFjVB+Z1Xv
5A3MC6BMrNypM5OX7d9q/Het1hghLJIn5mD2179sqOkdIV5NW+n76v124lPIhJYRUOEejl8Rq9zW
HYG+Nnu4Tv2q/usBbCFyOi5ukQla58xjlac1fPdxZbJBrvcfOgdtPfOWeF3pNlTqx1ZuWTMpKXJb
1IBkQa28cuLduZ44i32OYH3GITycKpso4mr/DZ0hCllWjbuQjYbYyd8+ERudkNQ7e44YaX4ZyNhN
KFV0QXdbZly9yx5Lyqf6WKBja88MlZaDP4+3tHzXlJpzG0UO+tKIeJ6DXteUEnClWQrWlWi24y3r
sMscGPStATtqn2dxSm4Ip4yb591Sy+TW1p6S4SkvIPQwULu6fLEDeNP3JyxRP2ds3nG++wX2f2Ib
WGc/DFRxHnfr25sG1NG940INapPPoHImqshFRvMQzWce5EvwxNYjy9fufz5amveROlFktdy/eeQC
HJfo2t4UAjhsIdAWj8Apd+1+pqZMVkJLN3Rpy1FtA9do6OlAKNeRi92FJfnywA623uz+GdX+14FX
K2u33YpsLui4zWmbZJ1lkGOfoGgejC14rpi4ydr8vnZVH5WA53Dn2l1UZmc8r+odV+P7qDnDFGXb
oyzE8M6g9x6BlefyQi/kmNHWegiqUYs+/y9ppkx1zfd9UjDyuv0R2dg8GkANSCZHeoqOy9Brn9f/
jZioqfOsKjh9pKnADh1cSiBHwGn5piGSN/kToZ3RhngWB8tkeo6L+XCi/ilbmFFMvLSBPceaUB1l
fDChs0xhKFsTAl+OTmObex5LE2vLCATTaW+trdoJbLabm+D6iUwdg0sqtXG65zvWEYSrl1cAOA0r
8oF8L14/w/PfXr1swZHt7eB0lMUB1aOaTo7K7qA36hTDkhazA0hiSN2Uz+uSOW6MMKQ2G3OqOXQN
mpgy27WRUiTw8KvditVDTR/XoFDTr2tQqI24ay211WFxLkaSk9cY0Nw4Cc7VRTh0xcdwvBDZtvqc
T64pcmmOtBKXqaT+OQtE+vkDlCRJDP/Zdp2w9bou7tike/ZgEoElPLRumgO7GnXR308wjr+CSc4Z
m/dfxI1IzmqTqfk+Wf3sCx92y6C6lauycoZPI2flwHeejgkttFUs+4Z+HHlSb9b6IvovNiRCv/KY
0IpAIeOTCjQmxr7ULH6zbdMpvbR4t2sWxRzBbI6Idnee1K1Svd57WxgH5Jw2yub8eqWvRcpip10P
wAXDVZIGVzgo6qE5ZoPURzVnjVv8sCI0bi6wdwmEEhpM7MfBRnt996JkP4qJdRE0TUIleenHMrWm
ZAyT9zHfp/5JqZJ92WaqOF4wSTZZWShX50nBky+NRw2xVKhvQfPcrqSXYNbIv5M1DzQsj4bE7Zn4
5G3DWBJ5e9wm4gbnFsXp56zZQ4ErFlNUyoP1zkYfYAW3qu7G5zIfXX0ZiT9PSunoEkKrDYMplPO2
9cE+QGsj/z7645se2vsIb8S1qfTMwmBy8XTmzmhi6vlNgNIJr9DiufrYjR/5dabkyRJnOZ8KTgl+
7rLoa31DqVwAW602VFfsvK43WMc7+DPT9e2Uf7OlYTR8k+wyV5IVQBtMV85Ggc3MvgvRCaJajuA7
kKeIFdbEP46emkk5NcIjryGGzXwmWGC7Ipbjuut9rEk+LsJYRJJklZBfTOCKDliKUsDGccOmY/qL
WJZbo7P8zu49bl7xMShyUaE2vWT59Ucntqjn4dnFR7pZSpKOsvyXE0kxw2mvMOvOF+b8nTPS8MaI
z+MF3AfbrfdrXv3dYn3yD+bB2Ve1cDtwsNhxZDGKtANF7k7U7oFvp9fvq/VKnkhVREg/C5XNu5Dp
xBjZheoE58iLtsusaU66Ffdgk86aPC7vOx+BYU3OTuW1pqlIRyGbQCagcoW8h46YEA4nW+1D2M2g
ZeVheUc6YywwCXMq1Mrd4LNAEZSt4+wHLTMK+NWsbt4Vfhz9ZZmYBaW/bD4uzITrOs8/zwzf8UyU
BpcjR20Os00tmhLf+iayB6sI7/xIINDmq/QoVN2wMWzKew2AB11pEj/mZC5RMB/lxVcR6vULPLXq
AxDI0Cp863nB1FAvCU4NF+HMIHnKInaVvKkr8XdaZklM3GfuURgJOdsPagMIwv48ev9NFROITOKB
zbqYwB6rRpoSjnULY61U+BsnSEWxbowIfwcMTU9Lz97vZsjvrRGtpi14I6nxLmrrf1/HvUyPrgEs
TVSsGxATrVpI/Gw0H5dcz6/exhz+rrN+PbqjdIJFXruLogPdKikrmnnDFG9kwu58mzQnLZFV3VIi
adtxXdjFiwAE2yBvv6WGaxJY0kL+8gxV+eCFoNOLfoN+JGE/C/4gkygzJs4enKfQQdCYT0vOjLGm
dvJeOfWL1XajJu6uKrGsev//xzHojrMJw54XS8e7+sqAJ0+uC5gFc7GDfUvndVPWj6FykOeGYMh3
xKoqBdkbpANO2KofoE25eLbNnCJdnEW7WGQtEd/YIwe3MxQhD9mI7BxTkWrTlMEDJtkDoXAN19Ou
8nHyz4V3xNsWQ7BAavq0aCPArJ+tm74T9k5w6M22FQYYb0iqHhAE2890tHHiUd5MOQk5g8bqKpN4
cOCxaJjuJlTrKl2mbsINX0iR+rbBINLR7Teh6jpiEUiDAUmyRm49Twbbulo2dCGBfKCc/UGyonn1
p8stCuRBT+qSQQcnCaZPokwiibo3LgVlm5zebc8fnQgSS1IDd3dLtoUcI8awLx09PCTpX2d3uhDD
b/Y8q/e5wQbYxbpJBmSmYQ2P2oqgqc4Ps4lno5TJ7scI+6nEo7QDaxlSSU/mHH8Nfg59FCzkxefW
o6nTDOV+v6wNo5H1dJThWVbbGsqnisbyN0ZZ9E/gzuwdkoseYQ/LR69R//Dkj5K/rkBi+Hbngjx4
C2nNVerN+MeSZ7b8PCc9mdGzXNaF0sdBSSwHX9aa7m4L1JR0PdF20+Ft4fhBp2/crmQJmtUr/Cce
UoncG0LR2vVhfEtW6KmYWEDvs9OKRkQmHp0XqNoctyOD+Yy1wPNi3k2JclM3VDjkkRLe6kDoeRlx
p974DyGazBDqVZRJx5MfH+tCNlLuTUZfsju23rWhclDY7+zr6fNO+3OT0N+VeqSvnlsEXgXjmAAf
mtFppegV0jpnCFBbgLxS6HjHtva5YFu7neUJn8qBO4YD1JFctg4DNfPmU4c68mO7tMAzPg0gnCmL
O4DVhZJogTg4ftQIbSK3jZDFylcRVibyHzHAezprKrj/eLK9RbfBJkpqNju6yJB1CE933i+bw+Vy
rP43XfIo1olEscLMawk7p36GwT8vyWuSdRLT+leYj8uKr/1SM+00c1ck9kkKxHk5fqiHSuv0Y+hO
9aPAg2krGtCCMggeI2UcV41eneYqkaStM3a0xHQ/VZpgvhvcAy3RBZbKwuNIeKsJW9JNN9krYjNk
SF3FAv7gsi2u4Gz/B7HFwwSd1+bwUXUvv71/wV/C4vT3t8jZnycENQlrwXTF0i+Vb/5fYWYQb5qf
Zharx5QuiIfkqiTF0Kngo5lihQnDsQuzkarwdJdkvFbSoD2A2ccSneGsDYjb9o53ofO9914z3UKu
ZeIRd6n7iOjlslcoFdU6nUOPUd3i5D3WkK+tOJgDWYJeXw0+AGWPpBkZ8Ht/t9mFNfCFFuNV84uA
hGO7OwxkUW7TblbJf5DDZpYcHBaLhiAatq+t6JBPwBMY8brdp+LHFnFq9uF3UB4OwB0F9mHzR0gN
p12uz7z6dNj8H+NRZ1XznUKJyVUj1u93l1ZDATYjQXeeD6o96Kp64Jqu+GZjarpgPWeqDBuUHPkz
9jkIY8Ftr7wpys8RW9BaQv4RNMo9wnYc9sONFzpcZ8Y2sKYPSTgJwz6sIxKF08c7D1BvdtAjTk6S
e0JtMKVaM4hfWpwDztww1ogGnO6cl5SW3A8CV2uG9XkJ/LzTek5Hzt4YW5VI3u0arzw2J/NPSoba
jIQbSJGVtwe9Z1bWATXxBXw9mEYImzzkKxY1dS2ZRpQ7lRXmd04Bu3Dix4gOoWa5lfcJ4D5Lr/E4
XrgrH4gq+XQ6BKc+GwpQJuh+bNVlIh/0gD2Lq0Q69h/e5/z4JL9n7uQCn1CVbGTjE1oIaJp046Ab
kdYK6eHZsvE+H5azfS7gEA1rM81OTplxPwJQmYVstJFBT6O8ojsBFuOG5NpXgs1qVnXA7rFNEC5s
7F357gtq/HwB9U5elxu8SfTE1Saugr8WamyJIF8QyU21tl9EO4r79aLvna54GR20BaM0uRALL3hY
XtQhXgTCfKdCi3ZdAaADiRGe27RhZrgtjfA1+/ACxKwtlSJ3zYHmX1gFGq3sln38l/ybma/oNN9e
skWDuAM3NB27qY7uvdiaP+S2PAIyCbuJxetEWVsrGl50VJNn1UXcTZVQsKHcLJEEvEGQADOAwVWI
irKPovkXtW19caf6W574YUaqz5OWCPZ0DWNN3JzMe5vdXvaft6HVAF+n8WwJ0oKYb6Gyaj2vyUvq
iTEWtmDnUbzqsxiBSaf8R4VPMQp29n/zHNomm+IFfJJDqO9VjDsRPOP+Fol9GYegIH4D4IvbAAcS
jbL14C8sO2R15gJXLOmJSfzn4Ht+5Pt+3wSlfK85Nueygf7Y0a3SENzJqxY2cd921oAhrOgzeKCQ
XU781q76VZX078/kKg2NiKwPCAN0MIFdYqwfJocBOXgVXPiSMJ5RD3RbGXgrPVF+z9Gd7XVuBtTf
1bUJgsiKAE3Gw3BTA4aQA9QBgSGuSB5duCLjbV8bOXPytq3seFERDDlUXXj69mciU/cHTWgOjNLE
Z3LGnfCLzfYhtKijDppQI/CHzhtli7+nTk7vg16qcvGD9L0z7BudCtMzMosAlHcl9/VU+rq5RkR5
P5z0DA1aLwh/Qsd81NeT1GVgbVZ9fAlPpuciv6w7HKFYeikl9zQ/BjFGLQb3ypWN5MSHQMn7n1WG
qo5CbZUxoUwn8U40LzwF4OZlgJkzLzdeJpdREZXddN+k9ko3nBLFrBq2Y5x9Pg85SWjMZAqCx7Ol
GBsCt7mWAWzYX8AL332dYunS0c7D0SOzZI7tlJPRWpIg2jYm/hzc+N36wJlMfEh3YDOjoyEM+h6L
roDK0KSYrBx0yQ9QKXNBD2ZoQS3Y+diaQvDj5pLAlxrJJER96GVduiAEtO0q7MvOsizc++iZw/Fv
ZFEqNEPlTUhe8FNmldpo5yaY6HwtSTWsnz2gGiAmWld4hAAokmHZ2xrEAZQYmElec+sBaaJYmMMx
tiwbB/l+ai9s+etXLMfWzy6usTRSVgtdfkvIXZ/vXl6sLocfTo5C28kuyC6lUzk4rF1lU5cvsiZ1
KSHm8TPYwYIBDpYU1ZJfMm8lgttVE+fIpcJ5D/FVaF3I1J0hvUHSy0QeFbyfWUB6dxoSHv3nEaU3
dzrqvAIYJrhJ90wu5K5E9lxspnz7uME0XDLKE43xP9x17Rz/jAjCR+hcOb7NaK82DnYRKxdYln0b
gnvNsP5If9hY9ZsZqttKpeqHeZxoUR1FS1Q3niDUfpsZ6u4GfOLis4hhivpvie4RZgA20fIaEdom
+y/h/3PrNcS6MJGP0eQbeOiGNkQfdXJuB4MWXOu5RkHU59cggZ2TowAY8ZUaoaUdho5QerpMVLm4
SJF8EPmF9LBtbW8gI6T6M7GZZRSBatqMA7oF6dtEpjwcQQFUFUJbt6R6iadnGCDfI8EvnCUnOoYx
igQmMPicEDqYn8sgxC+VSZrIFPSvXyiTDDbXCC15G9E3If4eOZQLaOKIqV1zDvgQJU6XazyYebSc
yrwMF8uc3RG065mo/eE55bNRXR9lpmFtvgeCXfIDQ82nLHg2m4sury3NKMKb5HKDwVrKAHtT05vg
BsRyvG9kgDtzOiuGsZcS4VVWFPSZWeqeFFQEE9hXWkJRq50b6zLL6bgH3oY7Ktx0UfiHBMabq/yU
hrBJyNTL+pJorsBG57NMttX9NknNe32wkRRulqQxmukVpv/FlTVPcYjj/7fWwvFkqlz7q4HElb8k
Sz5QvFnvdIw9jCNazXzHHIMHXYEgjI5tSzZp/09njJDKEBGpDIGev2XEa4nxW+xuNKBzNQ2OXDwU
TCHzz4853JssaOZOlk1VyQ3BvxABgDXbQIXH0LoO2fbziLujIs9ovclPMOzFNO9UTgdtdQI3DiRV
odtUKtq9lNmOSydZbPsKOhE0kg0svhCkbE6fK5z3zNx0C/zvnET/JwKW+KF6g/PmxjzECRWnpP8o
8ja946gqsg1aZd3X7sq7MlUc0PVxzJ38eQqdgfb0W/OyIgRMcmeHXH+woOT7SR8i8bqsrILygidj
sI+Otjt3cuvASSckBZ45QTg2aV0PPMqn7LDPw2vHbpcBnhrRzUDue3IF9H+Iev7bX61ij+x9uU/5
nj4fwX7JcdXxtBPrl830a6w60pXqGamJhENLEwSq9MlpHiDh36O2suswO29rmVqLdxsRNyafOysG
VuNNaWpJd7fmlvOYcuX8CvQp7I/fLn5A7bPQKgImpR2qmsv+dACkM1M8BcO4gTaopwZtMpdWbWRe
TfvQ3qCQ85u9OL5dfSSphTyALNV4LiMJVyG8BpTKjhQL02H4Ngk6eRv3ZUqRGj7AujBJ8NRvAH4s
NqyKz8NMwlpTaHWX3tcNghxTOXIA4OGM+LcxTT4UxyLmG4ybz2tUDEMg4UYb7HzUAfrAWu0/5K65
nQHgjz/SD8RXmaSLy1j9KBf6B4Hdj30zbUtKEYx/ERNQE2uchFNNEICJBsOVVbn6DbtiLCiCnu8P
U9o+ne1PmvAg6c/4p9fXmd7wC2akbzt/xTnRlO+criLsGU7oZ9XdAOCzivq3+6UvXj92Ji+3+DBx
nFZYJpV8wLftiBiamUkhhv2jP62EIxgsJ+FmnbicOENRiYNG6W1SnxEMf8jZKii1hpMhcduzQkhg
19TyOcbiwFf8LSsH9VpTGpI9BX0gq8vqOuFw77ljMXKp0IRKVyFxJNw+uEy9MHmowZ5rT3jDwdFD
NXfb1SuI2CPuGM3E/m3bi+7V3NUgSEF0nKr0x1bXh3NOGjCaAS40sNozD/V+VkcamMxr9phudSHv
npaY1BIR/HS3odOv0lBoP1Lms3SE0tY+9Pum0MyhkCAbxY0gXtAtpzEsJl7RrewINK3cwSUJZA9m
ydVW8V1TpJDRQJ3xjvAduQpGVPpIVLefu/W3zn1zMQB8pUcvvZUfIaov38BqFYKQoCi/g6Eam87A
FlDoYHrcjq1bchGlQmTeZT6EpgGE8D6Jzo7Ig7NPhpB+CNaLmiAYp8lOQRqtPz6sBiRXctqC2wqb
AnKW3onCb+M2WVtvysALJ6WxV4gdLspvAMAo9CA63Bh8pPT5WWwAxiax1haWhkQmeaUlu3AIuw+3
rg1j7ESkAhLRHrFugyWbR+AH28D9I93ozh9UMiO0jSK24Kf79UWvTWrz5r9DdHrge2cYtamrQFV/
DlIQbkB48nEpoII3y6OMG6z8RW26DI+0fQw5yugY7nKWG3govqeKEznn5DiXecMvjUcHjYUSW7Ws
ahQGRxZt9nS6sbu/6HdeVTGKwqDIP4NO13QNDsaC3qeS4BenMIubgKEfTJbtYAhq9y7VYT2jZQz1
3pCFsc1tdq6g64g0HLOwGKMYFRJVV5LLmIs2uyvh6vO7LLSDxp1aKAP5y4s8Hs3iip510qvybmgO
8BXGwIC6iQn4dVS9qtEoO6gmFBYM2XBiWaZ0VG77uhmljxquanHrk19UUq0ZuT5UMtwk7JvXIPeK
iUwc7JRQB7aVigXvkNVgDkwwffihyi8NojPKcqHFYGAE9D4x7u2U7MGaznJB+QzJv7Lp7h+pp28Y
KNwrYj+IduHdaOCZ4HofgQaD/MvJc7x9HSYFihu3MxZG49jbJvBG8mOPW8qctf32oeL5XGwNyWuf
DODoGkIx+h5dfaav9p9x8Ag7LMQnVO5e5Rd4zrptGE0nDcMguoyWa/Dsc8sXPEZBWJFSqeOj7EiA
zUEu7NpRmp13SLRF+64082GB7k2Rfrj9W5+CCNL/+L9Gj72MgrhuEPs+m/REn4iC6fJP2ZZlV1vA
l37SbdzdQ7KrOxCrJh2tcnFr94W8WuqdIr3rmYLtfLFFGWAuTBClfDqAVYAdKT/F6Asgq17IWEex
M2p6FhBgJlT//pvuk3WHViMxjWTbebZc2k5N5W5XcrDVfeh1JJZdKtdqyIEcWBeV1bIyYh1UE7w/
RBZw1ali4iC2GZMHG+/Xf/e6g7yMWdmpChtZTvowa605l1XpsUfVPJfwzWLnc91nQCtaf2LwHBJG
HpFpIjCGmt8uolOkYrruukjxOzdVbDXIzlQt23j+LaIr4wL3mZxKUTS6weM65tjn2oWu6/SALDpv
8wOH5ma4bsUrfONPglyMbFWKHJ0HPw5APUtjEeJ3jNSVKdxYyWs/nKwDyOuNNjBd6t5jZqJ2omm0
/oAxGeYnhUuJ86VqIJESkORtAzKR8POOHI5AqyOL115K88eR4gziNM3E+Gk4mkozqCAF4Oug3qWr
wTtzRdYpgtLJc7ZYy4oB22ybAwVpuGzh9dx0k7EVlTVw+Z+oL8oxYxv5UIOXSItXJTf1Dcj3J3DV
wnLARmgQYRnUJho+qfQwziarX3DPii3RHJbz7UFSqtdoXO2aIn31tZT+KDaKoPsfiiXiigvsbP3u
W+loDF9d6QkfDDPaPoWZjRyyENmlbpStzecWmJ68s+fd8BLu7sByQQv8OscK6MaTjYyzIYbZ04iT
6n08SiTb6QAaFDc8qr6e0prbPG4/D6FreE2Xski+njWenXeQWxCft8/8UdsU3CsuGJBgaoOoXBSy
/BL0W1FmGgJhxfstviW3p8fbec2ZeidxUDxgu7pqW29t/C6D/QmQjroDwVnCHa9S4rM3JwhLjbNk
VFaNe2fQJZ6OGMetT6X27ud1g2NBitsHFFPPezGwHona8J80sejvScsQg1HGUJoWFeI7n91gzR6O
4YV+T6mT9G9iWiWef1m0s/Wohi7ZIryuDPuJn7ZTLAhQwFEqzYUAo5qE+HXt/8oPKMweFF2yfE4f
QwOIG7csjbeRFNGnhdyzFAlw+t5/IEI1UMq5JT+1WFngTfVEJwOcbFpRwo7gsAS5Cwydnq7ncTd8
ZZ2PGes55J50dYp0Rruv9MXOjTtxv3MMlZTWc//eAI+piVsD+PDZlH1V3jYocXO3/Kdpu5ZQvLK2
+2RJ4bUNqAgDwARZqCehWcMkFtnv4Xtcl+MjzSfUapZSEVeqxi4UpUzhEy+OzdEkSBCMFwq0ffeX
+ztJyd6zwVBAFhSAlOcZhWSiVi8vI1/8G7yf4cvS5LZuAM7eUiLdmIDIwZWD7+dd2Y8xuEbY4JvF
bbRMQApeNEvVISQpiF91avWfLke5N9OchJE50blXIjP+cI5S0rKKKUuUuqbyfv9G7LF3R4Lw2T1F
Fd9Of/mEIiW7Y6IZCO/bGYOjn/DgSyW6ynhJlZYzHCfmaXjaWyZYZYSu4MMbtv0WhjlQHkL4fNAZ
DAc9OjFxDv9WQzy3jcvnASCYWVp8lrMUBESlUbLQHB7DQYsSaTjsGW1zA6FqVg/8+nvb5NUcMefb
4WwMPHUbS/aWd45XEBkJ2ZzY9GlPsBFaGBb+PLAA/+P4ZYfwrPkSZxhQBeIkzFPB/moKhT9eDI29
+XiP5TWQKrdEm7atVrC4PTR7eBIfQzVOwYUlhAsEqE1JmZrvGqquqG9p7qqk98EaBscI3xLnXeDT
kflOYh5F671Jtxh1GeGMelos1i5faldv/LDzqkpmCqlZvYm8mFgepPS//fmC4uQ7EHZTtfJhBojs
MVvnfHfn8bkcBFE2tB2TTA+lAAswKFQPqPnJFYtrdApRT2ZB5GSJIWTx4s/rbG1Phe17T3TM9kmu
mM1h1jlFE+DuG9lGFmnPDiT73GzgDIsexT+r3Zu46WCiJGrTrMuVmqc5BOhpPGY8xRJOAv/BkVEM
mfwI7T4nnP/EVm5+sSHl+fuLYmI5CAfeXjYFrOG6B//dbfpucLAPygAGp+Dv5cjoApLHp8iV+xsi
k64Vfifp+XWeL0TD1d2toc4mXilh1i9BO79xJca9xj0An7mOKAL2RW9jVFRUmCgtiEvgE6hi63Wc
PawtslJ1sGqYtN35Oa56DKlK9qnBoxZRg5xtTKNoNXFeKWI5m4VpMxsXnKlzbsGMs7c93b0JTsOS
YrywDZFdwmWkWk9H0c5kR4YwkWl81fQo7oTKUIXzNlcGYp7DqF0aTnATWV3oplp6vHPgzxl4TNIK
ePYlUbcn/VQduzAsnl11TsfSLQc4vG9Iky/eH8ePrdWwQw20S2udGQaHd1umN5TQNNzK6zfNVVwA
UG7aP7HjM6vWk5CLQCyjvmJCpVjUHOP0lYxsm3z468l71EYdnRD4RDIvIb7mfe2AAcSYVWjYbZEH
CtLisY6ajSI1UEGSKxvVFDXxcTg7wpzCyKJS3uV+E0Zt1Snv5VHIUyE19l4RM9cba9Qywo6FgMKZ
0lvuNs2iZG/BALUWMmDNRLrpVYCR9DEKDtiQJmeWrURjjHJUr/qR174bwVcm5Lhtv6IlPtw4yWk+
ywWHb2F9lfPeZemm8NktJ74pYhLG8Il15nlsEz2JwBpQHX9NtMNX7FCboe9SfD91NhhksBgaI3oU
AQ6L1WFvOUSEHAqRB/qAT94RpLuiDUoW1CcAUzULV86+XQ39kIl7qxoerj/4Q7CvLEgtYZNJGy8W
wWeHQjIMxo8h9ns+oxhvLiqx/E7hrMs2YSo2czb3j7dnFZ5afJyY3KBwIVradSQUGxsqagoeraw8
HTVwS343ljNH5Q/6nf4ZZIStZG5rFiRC/vGmYwU8Nd/ERRbNWv18jgn7d+8HFipMeOMmklNS9vUK
S/qe2s1cts4mkM7j53FL8iJ8ZfXXVrY7rFMZpr3w8bodu1VZzU75pE5sEQRh2rNZJXuiy9RoRu+/
n46GPNtNarigb8iULd4pYhJkBcPqOeqDtBYp70XYgfqby9eupUuy5b7yq8i6OJsfsNeux001/5p2
hoa73J79hg5Tei4QA/4sw8fsI8QJ4jorXfhO5v0fqHF29nLrQweZyalD8ZMIWcPYW4wcLTL1Hd9k
1V5ITaUDndQ9KPN4dASYMvwN7qWPFwUPYmS1G53MFfBaJeOVK5w069KvEl7uuYKW+3wWd5whQQV4
AsWfyp7LzpwBku/xWQ7e7vwk2BY1FgPEn5x4NYCa/FzNyFWb6u6aos8Ulm2uyBuJ2DrUnGQAA23r
mGulNGj0wEJ5MuQq4RXvjsQRb/b5wZp8eAQ+dfVbtU5OP8RMfDnykstNuAyM0+dhUrX6dXqH/h2W
6n+iW4sPc3+OXiGa2kcHRzuKhdLC1w63qJGhvpJVkaysowIXW7X5usjzAdCxO2KbrBhpy5eAFcjK
yJZWwXLFm1KdmsXEVfRLzrA3jMDkjhcflH48+lQZuwst8x+iu0+lrDm8jjJ8XYEYxlfeYsxDCbTG
9nyzVMfHcIzN9ZlXkma7N/Ugu0iqZZNZ9wnagDs9kRVgWJ5EJYhHwVMqlf0OmJhgkW8HttRPUqGn
rJ1sPlhLgJ/fT4bQ9ArSak5jQd17Mcim2zwKuaqB6+s17LDdJTJc6CxCE3yXutdGHBNnACi02Lw6
roNfBATfI7JcbTrOgOVi6I/Y95NjABOHqSR11auexZ3SECAm7yqNW7voeOtTkea2GUq7LIu2FT47
P3kGrBZ3p2uO70LDdViNH5CdRI4QRSg/rRLIkhW22IP3ZMkVvgq7B24vfpiSzqhmxgVfgWvILF5T
rnqhwBtGy4y4matzSaU+KhYs5Vu8jsbUrb1GbUeZUDas0PN7GyQBhNsiPpi5MlAxWizT4k+mauuL
YKnIJB+p99+fACRn9twneSuw0cOlK9crVbmHs3nPJksn1dbp0VnQhTwKS5YhZypQbkJa3vjRWBN6
JnKXvl+VozjOazj+D6LMOZMgunc/4rp05/4GKo7RnHgPSfpW9xkhdCHUHrr7g+ijJJRw6yko5VUz
wH/VloNogyBIXWc1VQ8P1w3XmMDOwwEhQMTinnF8sY1tDEa/+AXTJuyTg+HseFG9Ro7/a8cJdHI8
TG+WhRfZ3Ctt4oOgxizZFn7Rp2lPeXmrMzCuYiD5zZhX2+Op4IUfdVZg0n857aykHck/kgqtqQiD
kz0IOQw/c8kXQ56to8ukpvSABs8Ekiojr2dwjZzc48kuOlh8ippMlwJzjyhlHOc9xoBw1uSixIWv
zj/2S8eWdL0+zysJTyoY+R0WraX1Rv6IluF/oi5xSdPl7fVwAc9ZdTKf43KUa4xFiark/iUHepzY
KMTMt7FH2yfB8Odi26q0fyW9KjJlhnXU9bxNuTuGGWWOe78sOWV89mP8XcQ4HwcyPUUrQ0d+SM0T
1uptS5TiLi1Um0jRCGZ5OHjLGUiINJaRxFHnwhPzx6+HwNRaLf5vytirRWzfuYt5ipaSENKDWAZT
cmLgwwjCGz5BaZruuMG9DyXFN1L7KP2hR71pwIw4L9muwCC9XY+1dpYgfrudEuMDSt29okNKw0E4
FVq4IKO+zV+WgAlphpN40bVJU3kk0UU8GSpBhyVbQnfpo/oSeh4G0zSeWFA5eTw7T+Zv26U3MTV3
mkMaSNkucXNZiDE0ApPHhO/MskPsFVEsta1P1wt7eattAuXw1Wa4y8JtmFeoIZfcoMe8Csixf4iP
CwCefWr/G3iwitLv54YlZQb66C2iSniKaGM58raJ/zTOYEWDwBj2Rnyuy02R9VfrPK9EkNeFgEoO
WYP74kotT/sA/V/DKK8J+kZ6CHCu8LYlA4J4UP3mjQu6oXS+hbwVAiqZRo1J7Cuco+vT0vPgWx9A
rQRGP2l8Bg3vroVxku9oMCW4xTbLr6sdEQrJ8UqKrfy75TlgUX89kQmiGoPhYEZuYQtxS9Ohg2p7
dR0DdL7xQUSivc1FmTENS8p2QkM49NRQgoX0tdlkChe0X8dHnjI3Z9KoZAT6R4V5+BBX7S7xTRKH
14WgHvGFea6U3BVYNHzUR+SUXFJqo00aAlXOfyC4+Z1lzEkXMSKjvrCTTFGvQdt+vCNk33jek5NV
LEbYvy4yg+jkbibOTp9AhGLl/vYhRfAolMyzypvGu/1vTBgn9mKmtEsoKgk3GEn5IN8AfDvvk1mQ
Y/8VMOJxCFOTxPtlUloBW5SCf3aF7VAlsik59JhrB2NZEbRpDgLG52KSidFhb2HflXGcugAVzQhX
24eGClNzbG0wKCIrLSaPXnDNLHmgwnVEYKksUX3ufHH920AtewzFut9ZVu+kfHNlsfI1VEXSNH38
J3Fsph3MFFj9FwjU61leJqPiEf8ru0Nr6rPVEXmdJb3VeuujaFZOh41psyz6l1SRpNgsF8gyJhRj
86rGlw82XD6Kock4gz5Z3rg+DqP6R5f4qayNguolu4I6UoNadjujVIiCQ+j1fwvNaZrqY626EKOv
7mizGwYK2qwaqmS5SatLaN6aPBQBQVZUCNthyPPSgMlqsqtVpfDNQ0iBPGp2DWG41BTquEcLVtdb
FSUPRRacJhe2l4CvFimP6U9f5hMwH6dfdmKtoqp6Vk5DrxPOK9n/3R+GV23a1K79z8VXiKFlpE4T
SlRLOM2t5DwpN0CsgErAFqgZ0uFdS3cfxUwmSANmfoJ7aGINYL2JfaIiq2QUBSzMNMTEYGuuXvSI
/D8hlW7vfV3sYXGPJdeKypgp2ozfKnjRtJ+Xb2vXggnsWckXt4WyN0ARVyipooS+1u/Jmu4FKOkP
zCxZDM9mwi6gohyMbOrvqbs7skT30xHcBm3xcqseZdL7h0iNMqUrTJuFSw5GmFj4CgDb4eHzP1KE
DeAbBTD7NyDR3bFZBzeOlj/+DdfNrg/0i9oyEmk4KW2LibaQ8wS70lzBx9qtV+3ylSgrT1Sn4LXb
sMptd8DwlSZ1ua6w7jMLhak3hA/GZWKTEhOUKu7F8lp+/0TLdAtiVLvY+zya/TFpXwj/r3EQG5AJ
hSi6zjBeUrqp3Q7Ou4P67Itin72iH4ujN0NH7d7dqYcX6REXprwJ+Zn5eXMw3tSuqOQcZ0YFNicG
kVFEDZx36CEzt8bTApq9W9MxhuvL0TsFZaXDpvJek/Xe2q5+2JXFjnsQERnfHKvaPuZXMp9MKm+g
9HIOSfJHDdMKHGBEnlIBlZbhe7Qh47iNRAlbHg9CFpZo1UYc0n3ZGKLOHZNmsh3kLb+EORT/sBSy
G82+uVVa6qjp2A/C1+2bYIlLtuNHgu5rzcojQ6VKC4rJ0/w1cBtr0Uy/ZPKOC3i/bPGYfO9snr4a
uFJ2dGukw/i4fHs0lWKX5KFMOvZPfJlXZhQ3Qx+qeJyXzvjnH/pbK3r+mSBjMo/8jEHQlodLQ2OJ
s7PEWQzPIeO0KsaXHStmKa66QhM1pls+B2eD7mzZIgnfzCEKc+gw1jSCzfnyRtkT9eeyVpeSSf0L
2ZR0jKAaDZmvzOSotCJNfIY0dnqnZsueegfCPmYevzbuavESBAoz3EGSfxVVbOYbzwJ3vJ7ALu4d
jIu92caZilB/j1AUf1VUtI3+s62Ve3HSKo0sIrd++M4aJkSOS9mtIg/g9iou8aP8ikeMo5nBxUPd
A+Zi/L0g4NNFomfEEsrwtlMo0389NUuQwy0miR9lbMoNR1Zr6ugwjN10L/XQzvo57jgN566V+s1w
cK5eMWBRtBKsdXsJ8BVLjeExz5afOJJnKhZW8cHPX5gk1I88tYQHBz10u1GhkQZx/HBH4GAk7htn
5XAdY1sKWl6RlYtXOfiTnpsyqAtx0dM9xX7/rmTlzkQ4u8l2r/9qux5NGwAv0dV3CpgyJEgidUkO
zlGaKQ3//njMTb0H6KefIRYqZXXLlyplyuspL3gaBtRnJrDSWdrUADkYT/Y/BISGAZrNkIWBPXzi
2zeUypMTnQGvQrrVfxcTx3J09Ie/oBOnaFxx0ZEYLs8aOOVzGaElubKZg0dm9isiZxzuEEUrKA5u
ruJt12nBFy89TfCKmT8xjga3iwPblXt9hSortOB1PfGY0tt7VnZA9IhmYECAe95DQK+U4Xk5qpO0
QVySXG55nGorqJqwbmd5Nnbh0yM8DZQv5XcppeuFBUK3xo2EhP6WEsNEh3rpKwkpjKu3h/9e5lHe
zLXMR/Ai3IAf7RxDPnj5QIpxN+T1fuGb8aVvEIx/vKXg4R5p/8mKaVlSLefg4htVq31gefg4JwSi
1spZ+TaUV/CcSV0r1i3pC6qZMj3fD4i1lhXY5DzGDh4Wj1KUUjR9wtnFhIjYGPytQQpapICVJpGZ
/dqOvEgC+lGDVKWZkOAuJE7R2K9hq9Uea74W3wXamOzaPsMU1NGW7DEKLblWJR6Gal2ahDdqX1PA
B5DqOhaBpja/LHEKni0cO6b1SXKVGe+0JILAbSbzztRTsgatLBQXlztbCw0U+Oy9bLsxIVpRYns1
8CwM6gy1yp1icafI6DX8iGkHRvhXZvKPv/2PD/GzWDnLQYoG2TWEVagw+mu9aIm5b+JR5v59a0Ok
MF4hCVKhzO0o5fixLr5PVpvADKRAMbfHTpbnEBhk7xzoAaVEJ90q2pqGxCirIvWYAmArXoyMzc5F
OXBjBNyL0x7IQqPZVRFY7ZlNePZ8Ya09/5NvKK6U+hLJsT5u7Y1Dk0c1HwyGCfy60uIbiDYb29Fx
6HEgQV+PRexuCB6X+1Fywr5q+h5fi7jVSdprBnEASwo7414Q9GM0CcVlw2NDGw4gLKPajLEBeWv9
NTxY34UCG0I4DEiFVP8jQ/TqQDLmNqrwy5KY2EVxa79zjoRTd82XosAH1OF2R2Auc7I+ur89Owd7
LVBUWJjedvNNVoB7e7YhpyE5QCIfhR7/aeL1PSiDpUH+0He3Nwh0jc+vF/1VpiT/Jc5SzohpI5AD
snmCcfSijhRGrQlGcAg3km73/aKSFTwjCzotU91vFWuyd0k9h+3V/Nf2Z1xplyPUYBZD8viWr7lY
1tiLqt9JmUBGI0UXUbp0VKmPGuJvdIMffzAP6QlfmehDvdZqUXYn8a2ykFNYRzIWrNYkbE47hyRk
Fgfoj0mrSSJjvYVW/js5Gn5k4HRVuQ4yn3JUuou6OsodYxTy9TdApuhxL6TK8J+9bOeG0rKZMwNB
lPaDPqGfgtQmsYER2hnEiCJvjaHGshSeIZxKBD4pmDZIPfVFJgKuXuG/sEUUe5rHHYDGd7s17dow
Kv5CoomJ+kY1xXc+veZCZMp1yKbFcSIqLq7hri64gca1xvWnFUz4Jg30QWHYcz5OejmsiB2ghqga
O2785E1L/xK2syRWatCuQbZcFWdTy8w4Lsl1ouGCM8qVZV6nD3uNE2N7IHTYPeNz3AKd3Poct+oX
zxVIChmvKoW9SDsLXJWEFaaKNaZiuOImPj5gr2Z0UrfDgGGKEDP2CHBHWAsdC95rwexHLMUsF00k
GnxjU4V6ZppWAIsCLlpaT0c7dT3znerZ23MrmKzSjc5yG+JccyNkilQ3PGlUZVRE836j+wrqJmnO
rxF8rTLnHFq4NUTAmQH8XRK2DjFRgowm3XNRgoZ9Kx4y5dgfMPE4qnVVV/GZ7vigd4fHTbM+mOsj
VvWWZFCLZc3We9R5BhnNPwenrvxA6KQcWOqhlScXw/6aTMHJaBVwOwTYdHKXaT13zPkCQpw0qZ2+
wm6pb45bhoUqKxkt5nywheA/tViuXnVgz2qCdRv5tQn7WF79+2ZALTzg5YZ2OUEavSawpsICzHlk
VbY8rIGa9qoGhbhXt/pWkmK3oClFbieS55SXvooS7WuV+b2ESWTlBiwhX0aOAvM5930Ie3nh1035
05XOgbWtrAWqGeA9YCxfdQaw0c+GWzjaIwzHFf76PBEgAfFGZBccTmIFrhNtq2dX2EOxvRDr9kIM
VTObOOG1fBJ9l69rWbQ75JNLfcZ03wcSd1G7DlAQBe7r6rmFsaf1oerR+Lakz+2qI49cAMULE6iB
DTOignUv18MiEYaqbtkxba+QDkRnGxPLpvvaxjGShFDaNBm86cvZHe7Ofb2pj16Y2Iw70Ai4hVSy
8lyuTxa0UZaFKL1u+Em7CT/o4f96Y7h/nvDYRxffK1LHA2gY4h+p4KYsYjgxQe0zB1DVQovvEUoD
Hg3d80OXDCM7olCtNC80fzvqIVyh5j9VIsqlbGuWd0wVStY/myvOms4o5nBbRhY6NNv0Augru20d
TJ6LgD4DPHyAZRCFeIOjcyCJE4zTbYSocHzGQZP7S45lt6kW4IVg1ODHhiZtdM63xcMZA+15LUD+
8qHhVGmP25XwzxLkcys7AQ5YeMO+4cmGKah46y23Z7IfgK7lT4Jaq78Lo1PHmt07NVVlqBLcJrUY
UD/Z8x6ExPiCbqje/SovCdhO3BD27Iwya60hrLnlMghcFt5ErHD52UxQ0C5HCkKV/9RKNugKlP6l
wde+JMtnbSBOjwiEW/9QqdXhd7WvKaoDZS238cZkgonrpcxxwR13udAYhh7s/HO7c/fFdQaIVk4f
BdD2rgDjJpNWx/bG3x7ow6q6W1pjwUnr5OMVUR5ZV7kPi9Mvc7nMAeVkopAeqQdCkaCvGpTMPF+D
Z43YyBLz5Z9OlBnVuZ4xs3F0UPKgrqWb1wHqCe/nLKdH7HUxu5d2LwPdApIREM7IuxLq0/Z4Ci2k
CIb+ze4vBX4ZVIyaV2Jz0sYihVKYiMfYhsmgyJW45b1KnTzW6EXHp8lFZ3knYS+PgKZIdqdnhAwe
/YuWnp3gJX+z8DizudJbtZH5Gtw5zkLgPqNUZg/GeLAaMXt/8MkpfLNDXJ7dSomWFtsujkz+ikUs
aD93KU+r25KQmX1Hs7NlGLWqmhvpf8TfE9ytY6f6YkHlI5mq7FezIBbrCRxX7AGEMpxIHxWxEJY+
dIMxiGsIAKVIpekNROtVRKn67jbj38iy4ezBd8eOMtJ4DFpshQgQiMTX6DLbS2qypNmYMxogF9W6
7IGMn7YlA4ZYmOBf885xxcwPzVg5w3SZXD0P1KAAZ1kCqVP8JDm1dd0Vsz3LlCrJF7ZL3+YV5qRs
ryBRsEhVH1hH3dIFPxfwsygToEUzyPInj8AQCKOM7rQ11BuQGeIerfQVogIQb7AMn3rFQwauWxGc
6/IhV7tg4w0CzeE0QfPc+PQywR/bFaiU0aGBQw1VKhdZF1xy7oZj3ghBmaiObdispdl+A4p0F9Es
zUnE3UXqyNJ2X9mBw3W2YcB/OrCdVc10BW09ObbSiov32O+OqAhbi33pr+ckJD20TqyTvMPobdKo
UwNYkKLgsa/ixH9L1A59jM32We1es4yjiJ+LoOsw+ZbKSAoyiDeYIqB/MiMl2PL+0LYy6lBdJmJb
/sNEikzTn3tCZgCMNatABdd5NT2e72HM4oX+pwFYEUHkzrq2q9viLeveH9Z55PRDyK4D1QolzX3a
zqzK2uss/xgvnZGlchpLFbw8fYJElvSV/cvI7tl/B3iFRrAE38dDEmkfZI8LPpjwVwWCNu2OXRLP
K2yM2c5HnmLR8wS/i6QoX5vUPJH/v6V+MQxweRqVPHHTQY3meWE1ZZH7fOFjEnUbRMixOOEpwDCz
m/8DuPb69O68bnOcspLycBDCvBqZq3iTJh0q4IhXQduB4kR3nAR7f8uTPnhpKAce35UbSHi06IVf
xqgFIdGpv5wIBR4gcxC0n2ocmbQ5mRMsGCs78qVSucmwFz+rllPBQSvjbfaFBrOLP6MOOgKsNgjk
N/QTGxfC2poPmkFeqRmifE4zmz2Gpu3TDOxu3P6dGrG8w54Sx6pdOz/EMd8FzHBZUuUf1KfuYV/n
Uf8SRMoXEM7/nq/uMBzFDrJV3K1rVfuRIg9fn3GlCvGk7r2eOlV5DO1sZ5l3Q4hCR2klB7ykcchn
6yF9FCgG6owEpKy2WZsg2ldAgsRrR3UfkdMkpVubVkfqLG5On7M8dF7tdwXE0CHA4LesC+Q4IMcb
z1X0lmQSS5JTKnbQgH/ZTiUhYeN/+nakm3vIgJYfZqMX+OruNf2omjJuOU8EukKIaBIapsbinOpI
DODAKI4vMqcRl3JPWSWSnHcGOdCpqlfFHKwH0g+NTGQvVO1S0Hj/TSrIOhqkWdcyS8rHnAFThRkv
4enZoueRCs3nCFzF982L+PMuKztRl6luoAiX/6tbeeJaaKygipsFdB/Fi2+agDML4QqV0oL5y63b
JlqMc4cNVEmKSo0xMVBMLFO+oKLte8ZfAJ4O9ZGYkq3KzQoTEB8dlvlwQep7GPY9W0/qXWvoJ/9W
3dOMFLDSnMsMW1t+5IgPiFca5he7leQtwZT8BjESuwUwj7PPS4JKafvQpiSZsYU89ziJx6udrYs2
WflAP3Wx3gx5/tKMIs2xMBpUPd6EdJpC1Tus8PrjxkQpWgXi6XiF/dWmV3E2b1edv+XIlQsgHEK8
PSxtftg1Q4ji4D7A7/VsLXHw3yYQG5sekq8iDt4uwIL//y+Z9pf19unNHjfgqfZmyDLzredCSRv6
i7PgfxqeNDzGLdwjfCf3cvyl66JRZhzFE6zR60s1QVI5q0FtK8H1pk8BOesjRlYNJwTkgX5l1XJe
YWvTkRKGofv7L7KkdOliU1uVATM+HOuA2zqmF67sno41klSrY/TLw7AGq+wKF7KmifwkTYIckw8M
vs6u7HFRlAl2RqnKay85v8/IRVWaH+AGpoqXsfFwdTqolFZJdC2JEoRU5Hur4zakWlWlENP9EIyw
x77S3r6Q+lZJGVIlxONw10SG9qwQVCHohZx6JHextXdtoeJiXEZJftxXY2SGGzsl+qCNfUe1KzjP
28jJl49myyp5i706W4ZfepicqRhLIuO4rvkpwKHX/VOXfVfGsk+dXrktJrApOEj1iLP1ppWXYzit
YwuBKpBXov4h2D+HbXwHYUTwL+PQsx+HnyKLqL2kmd5YR0ax3GDRM+kUKYD/qM8TlMcmw+x4iZYm
+90yhR9IX14YD7mEptLd2liAyb2zSr+ngEu+gdWhJexl7I1+xlI+cr+jyDh8qLqgr5zrpf3mStqN
wfcEPEjIDCj8inm6X6swRijcwn1rEKIlwu56MQaC7gHn8pUHUQXdT5DQBs2fr0qufAX9Z0+8Tupc
KuuiyS2ycQFAB2BAiMtCxmu2nttbKC0zLa2l2hrzE/JGk2hrCPyg+fGqXGXFPpo9Nb1dThZICZX3
RkevdS7KveHaxwM/AXUBS2ThrxOh4aSvkFShA/3ZCyLBtJKSAs8IVVKQ+o1oMMn47U5Wijk5ujeT
KffXVgDlqF8fMGksr3NgYYw1bo8ForRtWBy8gl+YL12qxG5r4f9aRlqm3CKM+1ukIB2RoKJvk2t8
5+RqEd2lTYPKxXwJYEhGgXJR9ZoL6U6ma2MhnybX+SMOW1Gbhb8LGnlR9o5LMHnqUlKnE8biKmwl
kvNa+j7HGRcF0pwl+mCKXjqDXCi7esr9W0572uhsSrwMCB4MBMH4t++F0XFsArAO8qsZGFMHCvrp
drSDy2hDo0iLGtrrNKqZ2TjcuGfdl/d7ZU5h44JLx1FrLXTTMOPNZcXJwkzs9Frrd0gtHWT+997L
G7UjqMhlfVdzf6g1SPKBCUE4TLu3CAkPnSB1DVsgvuvAhoK9f0holrv61F7Cgc7eweqwEgobwGDk
gwY9rMsAVqo3uyMdMtmaTz6H5jl6cGuXBkS+g3aynqyGrKfORetT/V3+UYQr+O7d8hdks40wKuJj
nQQOIMEy21tHyJUnBsJyldGDQBfT4dMiiJ+N8qz4xzkM13GK9iSkQgBBWZGyHaMi/k4+X+KxomUA
u86OISETO+HHe69FCd0EPvat8OS23VkGg5DehiAeKjCpZ3MMap4bKMqKdkBYqnPIuxT7/RW9ONvW
L3jhHcLwWbQSy4A6koCGaPccxYaoq7+LJoZEyqDmDqUaCo03PwwYccfBDL3RmHaJ8X2+5MQFKCyE
xccbHCWMdYedviyk3xpDMULI3O2Etw0Bu7W1v4sBdC+wVSuApvbvDYyqQSUyYjIZe3LXocYdKNy1
Da9Yj4suV+sqwjd89+taOrzG+pJ9vUX/K9On3QAIw+puGYNwthtLJHWnzPnaTxV0Ggacg/YgOetm
Y+ccVPjP5hPrOHv2fgjArG8pwrzQPDvB63cZqZYO/JDzV194EiNNFD1xnc/kFD1YAxRs96AAuNx7
/KrrycLIqXfMJ2rT8NHl9cs6eiLEIbfKcdPwoc++bz2Ksrq1MrcVwbqM/EVxljYCJEyPxL+sTqM3
fcpb2i8eZvPyHUEx9AjwzM6GTXoZTTKPumVzaoKTVH6DR7/QUmRPXJvPx74Lsw7M3WCNu/d5PQ7d
hMsa6dLiBKccKPOOcRmH3RFi79BB89VnFnKBJptj+N+XM4hkMVmAw0i0ajxg48F7durIsirPW4FJ
hpHtSjWoUdWWlpuhyisa7qzaDcdkGSrTnC1fd0VucWKnyt1p8Opa39Q/tX1SYL+VqAsOyzNYOOc8
Sv3Ief0QhxZCxdJ6pqm2epWsY5uXkkIKT7nuVCZJHo/b+JlAcq19IgvxWMWREABeXr5NcVMNQZDU
J/gFIwbukxj/u0xPQaOfmRW2q5BlNmR6v0qL/FRjsNC7JIpwF4LHuOawcTC9J23q4O9MiH5BGsBN
bEkWBZn1OuAA5WdGelV/4TDyuToHaLM6NAuMjSN39iWfk93aBQwqlG+wx4bFEBJp6JVoMR/q6XmH
V324j1FgO66QzHctk09HjrW6O84ncDUn87MZE+Qe0ifHEeDsBUQ3/FnE4jdHrqkX3D8X1pgs7vZj
UAr1YrfS7CCrNr0QBdwwnxs+Ef6YRNxNZXiaZsf6nrYglnHdQloMEvcu6tB4jXRE0jk6B2B2TnU8
WnV0NsJr0nyVqAsWvkFMlleqMRCsfEOSy+mnzzSO3Unx2GRu5UH00em5Ea15YQo0ZvnQGWEFoGgu
alr7R2ZWvLTtmNw10AUNSpLsD9GKsUb9fJwC95E9IOexkC3+sPpxdUAhpfsy6vR7YCEfzw4tV3G4
k5cYC3MuSxvQhoPYzSLaFzGPRjnESWb5z9lmrHs0Vi3RzvtMAUuUHsOp92hE4CxbaAn+3uva/hKa
OF2fkeu+zmwgEhLC9b+P2GE7VoSWyE67L5UB5xJsW7IPoY/RF8tF82Pe6lOWeqfvBDOCPYiDa9wh
Roj8LRIa40gr4l84s5ttkw4+a1Pwd4UsuhIjiBL5CJPMEg7yZ77Te4ywa6Onfu5U4/AWGEw8rauM
C9f8FM1/dii/OVUbCdESGVzwcUYx5c8zhuf6mNOxKsPGdpBF45lXubwTRpBSadPCRL0zTp6hsOGC
oIvVrmK+Tj3rLmGzZdoEPkSw6U/24NDQ2AaO3FfASt6gOSRO7jCDcRy9Isj9ZzzhFIQmQGV9SvEk
qOksgeqtIMz3kFr2yWEtGZs39Bpo2VnHXpx9ACazW8WzUTN5KxRYb0yeel8wF3j6AM4hOMwdfXDz
2izh7tnWfSIclGSJ3eeSKBMgdJ+NGq5YYvdWwOt8UWVm6X/SHK4qv1pL9snBQrP0IylklxRi7BnU
Jw0krbvpSr5CCJbmT852ODxoRNWZThNMAGLq/fZvD1JJlujIFPWiozookDZF9IfKI0lqmPZxco4G
WbCJoF5ZDb+Z+6l4NZRduCV7cf5EoNwK6ADJubFZ3kMvbqAgUCK0uM7MAjipw4fNQ4Y+NnWR++74
StADTNVAZyTFQ2rSNtthpPsR3B8juzR0DARnMecqSDsxH9rthMeKVOawy5L9Y4Y2G9JlHpGQiZm1
qU0Tno/Ehx/d8XMwHsOvAIcc8vBYZvjkV+tsEgchFPS223ik2kpQh4LcfLvn8IXnxtsg/B+rwqCN
EF5VZ+9RK+1xHj+P7c0Rq1dsraR/z4CGoDj5OyZsF25yRrUKBnloYKvbzeggJlO6hSdKBrRcvKQy
r9Pj/XL0sAZWg6rfiCp4oUiwvT8gmaFJeScH5FhEt6plGMIzPOvJ6iLetoUSKLWZlyOWcgWqFuqE
iDQnhiH3RBk9iQF0hqaxUkV/UzojsW15lTOIgpKGrZP5tTZs0GaLNtrv0UXasUA56O69v8R+sWnj
9g8CPuSK6cWS7plwL2dlR+YZY/bvYdG7pnF3VjsKYZ5KzxEzmAdJkWeaBegYJGHJI4kVKVVs6W9S
SIUeTKtlkFb9fgeKAm2IBJJ9hIpAs7ORfcI5YK+1yxEIn1DJnaNnm7vSYV+/UruQ9ZKSibKGTM61
85zFIEf7IPZc8a8lt1fv99RkeyLYQiDrvUZcp88vsW4eMePe/0ytbYkcmTR/J2WDFP1Gij5B6i1T
1YgGkLrw6YIFDmXhBtNxFfm+wmv5GP5b+QRVCWzxaqbvZdmLqehS67ncd7le3ydjTfkodQWj8sA3
Y44EagBjERbLftVkv3+I7M0xTLpKoAXEWJ1GXNA8Kww6+LFi/R6da+tjq8seS1asqYGHLRcP3CCZ
zGihLD/wm7d9FZPsUKkwtmkysWYvPxpPxoA5pk0/D/3qWY/YqiRzdxp9lQaDLSaldxwv7qWWe40q
pmZH1H7FxcFTCl0qCBvaeut+3TpS955+O8u25Act4IJU1I26eTyHNyqBaull87b8Arjxmcgtgp4M
/hLxC07bQDCAQXkwZ3FKbLLriNe86mra5rhUPVYlTswMQAqWFaBUz+GJ7x/AeK31iiSHKarRY2Pu
NE3grIbC/XX44B5SB8JOFlCRkQeAJds5WWaHOS0YlfTUG+noGa1EG0GELaLfPe+rvNat1U29+0n7
ZBYalyNEQRMOzn6dpLICbLvMSfzFU/f//ZdJ7U/OFpcLTd0Hyn7nbQPlNlkra+Ye6tvZoG4mqnI2
Fe6vFGKX0s0BcMSLyyOT0GbHIi9LLYnJ+zL822NMcjJOmsDqtJvUYu/rAoqNxBzr5OxzgbR1cxMO
SBJ3nQQy2Gy+3JJvQpAj20n09r7j1T6GqBoUqRPo5YzjawAd1RBvgDSG96B2K7KFDAuQx1Etp3Pw
L0U30+TYqOnRhUVY/Np7dPOQasC7DXqHRze9pyVoVFzDocdKOhXe60QIpoi9ey9RoPuTzD56dWVp
xYx3cysQGKtuoidofTr+DY47jrC+1YKuxvb1qahe8ag1rJLJkOF1utj0hwXFxB9Uq36/q+QI7yi8
nlL7S4v+0yjA36t/uE6sM+PovsOlnihpWzo1MOrDnSEU5kBca1ClowkmHnXYvHf3DOkT9coA9yLJ
4VFzAlGKEqmUfQVAGrbxuCDdM4zMeI3LEkh56Mk84//3wJePZ6rKrA114C81fY4bv3eDtWKtiSea
dde2vF28Q6SAwrxKqj8DOzVGLX2YmkAFde/rKI6xiE2kGHSmfDzgOGPZdtkGUye8YUN5nOVdQLaN
f8SoG3lcuYYn2Z2Ja2KxA0N2sEbkXextJMQPkJ+hiUphJBxV207bfgLsIyJ1B+fhuyPjL7hPvGD2
Sv2BS/tEfMYIiJjpvrnjoA+kZYSfuCh1UzFdclQ0IRri+G6eocROZqy4HhWOuQbU8x/ikT/xn/Sb
CkDz4F2MzmYVnFj9hoRxYWBMWor10Wv+nFcQUM26VWBj4L/J0fx3fpr0Zy6ooEMr/Hi2/ZuH41Pm
FTYcuO5+4lRFH/So7Re2GJuxp4319DaQqeHv+3dfBOp2JRgEEBdp9zdsT0FuKeU3l9P7rW1jPwl+
XYgEuX6kE5RQ/rJuNpNqlh43s8i8vWtFKbLpfrxzWJCUz/D4oUeoMf0+enejMWJu2bijldwh3aHp
RHJ/ickwaYjEudNM8dLvGQQfvI68yZsNG/NR4g6j1hpv9DAjdhtF2ia5jM90DvUdI35506qs1ugQ
sZK4NpVPtd1EscKplJKYUS7M2uhOOdhubarqACWsU60KjSg1eAthOrrmF08v3c/I/EuJQhcdwNLz
vWb8JWtdqevyb83JPn+Q0meHbb8hJbwH2QYqp338P7rps0pZZHl/IcwJbHq+uw8JqNIVQwW3zP4A
DQs4VNRiqJ5pNfkxV8XhJDkGbIgL+EVCaN7VJa8zsCWp9vGtmQNAPvwaPlvqAAleRv0UnTE/EJOm
9kQcv00WgbxKyjR4LyA1QpK5sovaYC0tJy4i6lTKfkD2G2m99fchzDd2K3idbYhQS3nL8D+F0Wsb
dik9E8nSnTm3nzE4lS48yFmTRgpR23ql55qUGGafCS5Xk6Ni4aoWf41q4/WvLYVu9FymSUMDQGJV
1wS1RQvLc1JwCu/ocQJVwPZQfGYNCL6OL8h0iXs4F3y8XCWIa7SrN66GJhCaE3+PNjLSWgvCmZ9R
C3cjHSoZcrhrTBxOHfWPHFw2i9FiMSfnPvmBod/Mqz7Va0bk+ukaDfXF9OUM/Lo5Lw9v+psVWlr+
EWujCExXrqKHxyRqRGecG8rZbV4URxCmpeYKh6sao6kSisp8lPuWbqDLwMx0x1Uuq8QEslSunqJw
ZJlR7YvRQoAuDJbbFGE2SAf9R3ktO93zoegHjYVwq3XKRpXgNRQABgyiRNUrxGngpa+PfUHRGt5O
VHkPmnvq1uxXCJF6KGYoX/Rr5o+KMYkWZzUNFTeYaqrRmKJaZSBRG2HAKKw0ofP6i3HlUX5551sR
LUJqjWpKP7634aSDHPHsqUoVkhHOYIly1mzZwRvJb3N/6Td4kIdJwe8/h/xqnCFTgPF+TYeueK15
IrhK58lp4YTcU2M05smklWeYNNfknIM8gj1+IcXRalS8mNSUgP7NRtLN7boDA7PIsUSctfLx5Yfv
/JV5yo89OsIiRqO3EQhvqQ7tk2jS/aAY8PoxFxsA3a5rgHtoXSlDKSRS+AycGr72bcDgwkpIpgBK
8OsXbp+JDuvrbguPxIJi5IQ+LNG914vShAU0jcP+hBkOMyeLfVM17olHE5adngjFbWJ6jWqMMeOe
zZPoacmDSwMAtl49JLCjPg+PLx49Pp+vBKEoX6HaW2MV2IpbbBC9my2v39DZ/tsrXw4oCE+oPlzJ
EJST/0VfYGBr/ICChzSSwD2aPCbYNV8oS/eew6q99a0PRA6rolJbkvBWv36Zq/f4Z8O7isAN3m24
s5xUpNuMHRwJNM5Pa5ywhyk0Hu3HCtB6PznH4POUTwcQ/x/oOu7bvB2q8NNGuvTQpuC4QCPzS5XR
bLBnWXJO3S+hZIBmwXRNq+ohUH1SQqbO8xrvOB7OW9TFi7UT4AG86XoA4sUCHMw2eZQthKuiAj2z
7g1NPl/3aP1QqNNRnf0ovRZLzxnok8J8HGNFTAOJZwG/1gm8DYFCpqungpp5512EvcuB112F1mTB
28Be2HTBWMIQSJA4yNvCvdJcSLt0h0tnquVLh8Z30NUqYSMzsU57jhsSFbehT3P6fmKDTWvcnGW1
/NxIuZuszni4dWrm384oiVf4ssA2fkefKdA8AXrV11kiCcvDsv+VNsWZelqa+zDLd0TDBzF9jSva
8NGGREXkjK1umLJBogM8BN04Hw0rqlWs7wEVzCXBzTUvO/qErmYmJNfTQ4rMYthKI9Vu/Py9LG1u
nDmSUTy3JOqaKHcVk/0T3T3AfyT09FKQB3XEoTVt93Q2Yy0WI6T9On6jGHsxsuBC79a5zfIywCIk
nLsq08iNqTI/VVOxCZ0YJmJyMvhdya9BL51zLp9g3HKu7SnaVq3zB0VjVjMD6fpBF4myQpm5N4fm
kta31snxOP4Il5RZfXYyKjJyQ7n7brp4tfqBM8k7DZeRm4SwXRc5SMlt1IZiOO61YA0VvGFs4OSG
AHyhbGDmYgXm2E5VjyD96pAThRmG20Vop57HgRjugL1C8XXtVXRJ7xkb3PKzqDs+6U+QfeLQmLXp
gZtulj19cB3KnqCkUYSqRPU0taEq7TFlUn/QXe9wp8TrG7iHAX8LGqbM0wlQH9zjmGRADhMl2R/j
tphm2cPJUY7UnDTKeJStu/2hqqW/XtqNvda1gInLzuYQK8SUhOQefTyJFB2Q4P9ITFDuaGJaAgjK
eF/M4R03+C1m5UsIMQeb0rjqfoAl6/cYjD/ApzwsHHhUak1pyTY4T4YSbAuSkw5ieI6l5xqA2oAd
XyZjTrRF3+tbhaGv1oCH6xjDk8hEh9QX6hxRdlEWCi6aCHtqB3W0+ZpVjdxZJTeGjDQUxKwZ79hN
LFcao0hfQ0HnbqXmfEFJui+8klpXSmoMZx7Tg19ED1PPTlQx5krAvg80v9m9Clxv7230v7OMM6Dn
gwUQeFC5Cqz7ACD5RjmaH4gUKYV0+aHL4QQNpAjih4byRmQs17nLZ6ZvuH1bd9Fn72g03I3ASb5e
ns9O3SoNBQ9KurZpXiHjMnUDu/w7mCtBrHRBjOxbVYG4Dr8n6jjPGq4mdK3g1aI9DD+lChBiBwTk
sM031vSp7ijFuuWYU54QdUvvHYTUrs/ThCjwRSZooNQQ5WJwCWHpIuSTeuaVNgHtFiwgGYPrdGhS
bZ07aP+heCm/sIeloXX/nhr0GCFKKTAi7x14dAmxzDyQ6EXrzHfUao0lsmUiUgyjKxuC4Yowf/tZ
jpKRU4uKzZigPQ2GpvsGZ/8Jbt/wuZhCCrQMZF2WRuR0udJgvnOAlJ4+cjGGiUgRaAdfUVL71kOh
aYV7SqKLGpaOBmfcCGSw6pEXK7NslsyqJtGZUaxj6sWSzToWb6rm2VtFigJSg3xVkVDSotHNfQ8A
F5VomNevo9fNvNfypeg1igV/Qz9ebXMglnmxVhpr/A7u1qSLK6dcXuVjGZmeKNGNGZpEPLxrby87
d4xvvl1Mp4hWebkdx0OvYBR3BdWnurtztri7bQ3h1Ip95mbJ43sEHewgJDwjde++WE8fHK3H2FVH
WqvDA159n/T+s18TLzhl+dF1i/tD8NSgH0xxOQszy6xokaiA6ziw2Pq57UsdjxggyMjrwQp4apx6
abA6GGScNfFhG5FP34vya218KckdbDhKf3+k2y78RYy8cDoeyqKDCNZNy7YkEMbcFeT9goTIzEn9
H69T1IBrPNiTf4Lld6zff2Mgymjp+V/92LXOyA2QaNzZx5v9pvvQCcRpOqBXfjepdErr7zMDRyTv
gzJ8pRC7j9mQP0U04IAFxQb2wYp2WiMYzS5c7yjnoXZJWWON05KMtbu7tKu7hRKR/ijNufhM/C9k
mKtHmsJaw9DCgIu6G9jCEQiIAC0LOfqEZ4geQM0JXc0b0ssUjGkDprPlsLeFZOSCl8Mt18XQO//6
PfcE2zYNDtiazmh2SHT46H9DK1GPjHxGIZZXyAtPHCzKWZZJGtgj3207ZNfMc1tqS+Gvr8WiaTzR
yaGW3EQradKd7kJkb6IwhUKqgvHmXJAyQt7ye98ULHukW2JKpK76vfG9W/VcV61aczWpOIw6DRoG
fmoT1YF+fvWYQX08JSrWkHxiS6KnJO7T1E6t1ZKxUsBKOBFN7KIlJBJT2x490tMC4puclq40bkJ7
1c7yxOQxwGJZJkDjYABbfdYsAHRSfi4FGBlSyIW2Mhvd6g5XswHPODByoQ7JN+m09Sy5mXLKxZb6
xxlnX0apPhJfv2TF6n5otWBsjuMtNGlmCIvvQLJBN3gG6tgPrSQEdLghe6iM0JrRHKovUGW8qYRM
XY39wy4p8ma3zq0En+tEyyEMS/nAS/JhirGf04ZrqUHL6gsSfOA6aXCTKww7Ux+podKmx09JuulA
9b8kQhbTKD3JDGIoYjk1dlOLe3WImD6nCyJp5Ihtzh79KRQ4t1RRKmdpa6X4/xmcTGOPcZnU3D5z
1sLkMR4UfmHb8VwdfU9jn9iiVwK3nTh3VKePZgeDE8jm+w8/ZL8O38yKxhgbbd+jBQr6yPdOP6B8
AqiSfR0/cphcgdZT3+xL+hOySwRvExIyfRe4QC9/7iBkLEOU4gpWAO50XNVZqK1r0j/DF5QWv9zt
wDyZkUjvvBeZ0i8mCQVNwSEN0FeJVzTkzJevn0B/ztRfEwfD4Z7pJqnSs1lz9P3suwUQy/HW+GcQ
E2euMBOdxRWjqAWhwWPnGyVbGAUsnhr+jnS0O93nZSae54o/I6l2T84dYhvYUafUAEVnMF7bmrkg
Rd2+YhhXePKxJXHMxgm0JZW+wXfb6CDq7XT3cozIHjK7ClXvudGnTNayyOESAWUVZiDU4rdeDW5o
RwT5Zxr2jdOLx+te2Z1J2wl3KvsZLjGgR3FaJNOtGdVWy9AzTCd8N06LgP8wBdcZzePIeBOxHMb+
mgvKcFURn8Ax/w1Nk4W0DR0w0pHCUNAdvR58CYgDNfInO6iMqc/FWN3+EmKpffmpjss7EEKdoau2
Ejd5EfV966ENOgByNTswA+ODNLmulWzJ5jYdARqkVYN1IJbaOWiwd6smrI/w9WX5+BS8ucsCXqOt
adqiUEs5eBt85ZNvj9S20sA21sy060b0ypDpJFQywFSWRqrKGZLEWdtvQfsWp9L0xD2Kp1QhMM6h
0dEaKTNoVdcDosMelcGlY0zCBlIsiwpcyOhdlmX3xNp4iH5sIF8AxVsJa5w+JRAjl8DwiocepdaP
3WKj1U60B5pZ6jX9Rjbi3qOnDGo/hxDGLo1f/IRUjYP1oP5BYDcBiFhpMT8wX2TjeZfooZCJt+mx
+EUTchzyXMiDBVJoyetOIP/AnyO7gUCWyL0tBqYNX296Sf0fzlUEPgEydeNnS9pRdrRkwcwTmrk7
ptn/d9XaGIRF5Vn+0YCS2aZCYAannslvtdco4Tz5JpubVXEuoxFLd4az72G/VAhlcDq4WGJQHRMo
SDeJ3RaRjfeqR2OAJQyRdLlpooGq6BtwGkEALAGOXMYB1VB/9pMjw5vyAVgAS9zMERJfdV4/o+OZ
pnJgml/wLggeYAmTH208g6BoozZn2qXbFoVq8KaQLSKbo+PmR7fXAikLll3QLSIui6ub8DRIFE25
pLMA53WqNWL6mIlO9abE9G7tN7IUWYuLr52PabFD3kaHArBaQkSA/W8DX8fbwNWdIbGmzd2muzJj
DUKydlKJhhhP+lAehBuq0NHakQOyx4CQxT8Tqauitw662qv0viTHhXUWNRrb2vcHCw2uHug96jwB
IziiiyfMgPZvkv21rqq7fHa7e03Df1DV77OBYyCZ+/lJy1B3D38zJ+x2TwZVKfzP4ZY6VSPwIDfG
73MHwSucJ4i3dEvE58hvxeq1NAQFRTtkTqDDKWsr756lbCwwkJsXtFEJeFUn9riggXFVRF9gL4aC
Ln5Dh5RTDu0a6xRiN+TYraT+VXMJz23m9JjW0t+TMSLCbLrNw9Vb9fr6jzyLpzsc56wVA6y40NBb
nt+XeubmZoPIGEJraY6QyEnGFhtXA0o8DD6pLgW646sMB3uf/1/3JTesqgytwISTYMCRXDNvVV8z
ddjJo9V8FZjkGQb7qVQohFlQjQne+Ls4J4Nhlhl+xG0C5kub7PoYKFu+w4ZXhV4XN5GWYsVaBgK8
MNrrsewi33mAknvTaeS+OasM7ecs8s+4HlKhfPtyZ1AjETKGq8YpqDVAU5gAS3gX0bLp8B/kpGvt
B7yJF9fp1eVY0cMerI5+aHsRKkNWLSA/TF1+DAOlMSvZRj0hmIqgm3ycZIw3mYjsm+PSKohWP7YM
FBu9QaikbeEj/kXgemJd8Tl7rjDrkKmkuJCVNKBv3rRzpERn/TjvsJ4QKUCBTsZZ+KRj03FcZyAF
0IucfOZg4oHVrBEgPliJsMijrb0g2pBQ5wYlh0yl9Co39RClL7OU1g/TcyfZvzTeycjAApUb+wFV
z0lJ3BzkAFdRAaQf5QJNUCaulOD9iBIDj31rOmsiDNL29Xxp/0LG0UvkeDcqgF3sB1CH9QeSmYDR
i1SepheUojXLiv0ttP5Jtaivt+Tgyc31Djg9yQKB+cte2Ko7HhGuf9UTbq7FSdyZv59LcOQ32DK9
vHFL5feRHyM0ljU77GtR76cwI697XhD/xBlKRWRJC4fGhwlz0RktsYjThM+xTWbpalJKOv1k/G5v
DkS+5Q+t9TOMsAu7Xmdw3LU87kn+Z9CtMkYKOaBPncKPkflHHGs/3P+WBb2klCEH/kgh8KhpbuI+
qR/w2ZUwHiIpwGSwXrXFuUEgKk034UJLuMScNoN97kwSFGHmtIxvAK2WW2SkUl4cawBoq2geWXp5
Y9ZKw+Lo/hs9VdjyJqaowOryyS1zLDBjdOGre/vpBzU/6/goKBq2U0W7o/2doei0GgdtjdFb2gHo
cWf7zJ1K/D8Pdjwi8rGa2uryG6p5135ESid052PKSzfqKBTbj7IDaYmdysYX8MMhNIJXveJzqyqS
Uw8d/h6HbnRmbGwM1g1kL6RJHX2m28oShf9t5hWPPKlaMQ3XvuK7lrxiNWokqfqXOYybxPPVI1Sa
2Eal7FmIbb2VyKU4WL2ifdrA/7jQssIdYW8iApqo/jIlHX9mpvBzRpAmPc9LeMk2x7Df4gtCCGZx
1g6ka6Frt+XoJ6BII2JIk6djUT8FsjqoFmmGUNOpCzgO7uBKbLRUDarA1iQlrIytex+Z4Gah1igl
4RYuWIhiYyELA8hCMoN2FkT/0wqBesdzeaRC3XrNsrwaGIRyeOGB4rCLpWjI7M+w0bLKn3VLavcJ
DnpZjlb79XEakGSBfT69ShEs35t9/WvtaTmMjmOTL8NnbJVAe1wEFJDATBvqyWqaiqi6dmISFpa2
gC+oVsXqvwJzIJcHMQdclKwf1kSG1eBNFoxG7/GzP1Qpk5vFHA7r7qz3HLDX322KSdc/nbSnm+tU
Jmy9L0S8NtUMut4qaNjebE3Zefv/4ndBGINvqfrrUEaex6nt+tzVw09DMV0gCzyI2YU9c2gAXlEu
1aKClTUJBQuHi4XsVJkB5uOlncs+5jUgzb9h++F85/Qs1sxdsIZ9N7+U2RgeXs+iXyeQMhivRgI/
hHokSak2vxPuixUL62EdOp1FAnCOX2JSAPWJzNJ8IiMYGFbrJrGWeR4er2XI2eVbeM49aqCfDAHt
i05FcVraddALbv3eZwWm0Sv7C84l+P3Y/ASij6Hr8xTwAVmmAo86iwL+TV9zFYLmuYa3LXMnkRaA
zlvk0UC2hAoNuq7afOcsDjmdiKiTdjG0uukp1usqMH82xr+MLgzuApy0Su56w6UPWpgHmd5yaF/W
VHlTrEXP2r0w8NFPCdwwZaUrlQYojEoYl9cAzdq1zTSRFPM4nyCLuK+GdEUQkLmG8el2atdFF7xK
ipENFRFrMdIHwyES2FKRgmu/YmoiiQaWUqwfkrt6ByBLl5pouVr+zmxcp4RfzqzqCFycXhb1g2e8
run1o9X0PFYu5Abu1ROxAsZFnwOTXvr7D8UZFgFwPN261tTvdYqe3o7fuo/FaZDcQHH8e9j7XkQc
OyDD7st9R3XU6CRvkpwAB5+Z9ZRah1E4BiD8CQ2+X76Du0vTbcLOy3AEUvR4IdwGn8/YwAQg4EYr
QbnFlvyP77t7M4c9XL1lqYmRZBH0IJlhNmWEmhnl9nOenPqQGSouB8Bf7QaRyYZOXSO1ZX3viWwk
rg4VExo/84AeNCBFff4g4T4dZcDg5G/6d0srWmRjFy6J31FlD9JojX1CE8WfuMPhzilD/ff6Lk2u
Iauk6YHo4uIDQIaEuwQdazy7G/O0od6RFF004tKHYHKNiAmZjU5Sp7hDcqXe+YM8muCa39S4s0+d
eziqf/HoS2AY0f9uX77lhXiGgSQScxic+9E/8xnEVgivoS2+QJX54h81CRF3oaBLTqi41A5EX9I1
7mIVrVgEm0D+r2ffTLhHfcFZ2s60wDgneVAVdWORmszNO1yHH4th7XmDujzAYS2szPwRSIAn2J4L
WkivaXA3WvkgNqxCUzkkGUS7vcgGb2zILYkVkzU9M9zLtYh+yEvcJ5YZb7udSmCcDGSzDO1BWq0k
WTsBau+LXMD4s5PjM7qfiHTNTwwMChU4IlX+00g5KywUaAxsif/asCW7x/o4adDIbqbSAwPg/4Xj
vhIYS89Hjy2bS0dg5dntif/baTjD87kSWF/3oJXq13zHO8xpCJ9Dl5MDOOKn3C8CobJ08SNGQe8F
No0Z2CfBUZJRnJbVyMFbkJbIvbjN7AEXARY2cwV8phMrZp9huGy8w2ohs9GxPPg6gYxFXAqeZRvw
t5MBgOabumdAW58Y0AsG4J+0UzzEmKRYmIPvXOhZz6fxeDBjnGcU5G7ak83JxDnt+LK0rDn2/Nfx
TCXZQuDqegHM2IIAfDIm7wRht22j3HYfB/tGvsK80/BLVgUUJGEphK0oAozZU3iY9TkgX48qloey
TSA6uDux61JoR7cP88zaIIzT1tr+7bY/wqAQtG/Y2JrxhmmIliFLKV/+rlCbiQnC9hILGGF5SBeV
VA5T62/xIXzdGIGygxQIwzK3MIdbAicSvpPOa8imyCoZ5J2+yaspRuY3OMVSrMPphaGHLU/sCcmf
GdZqPsbBnire6HfyXIdnXdNVhcKMGpwCOUf7RJt45fJoDeWpOyrQixbCw+GBgzplqa+1ok/DS/GM
2BigYrFgcYI3FB57/+9lUWMUsAhaBgjDmbu8lU1vOIqKeikJzP0Hx6ixmi/ZSzLvYfKue4zWCAuH
Vl5aUvLtaXzwbfR0AQiA2RLUtxnif7YkT1CAJkO4UnsMc9nFxG7ivDQXC+id4fmtiSYWWXzD4bhY
154fltwI2vULcFtOq92UWQ2pIy6804oLBO96Ytl/va55OGwFPZW4BGGurCGKCl98bM0ACWxiQayG
Wl0tF2TIT0l1DzGXhrGUEKyVJlphQ2yj3RBLBHnEhH9yxxmsrR2QcH+Ri+n5jOKwsl+CXauodfYJ
rYiu76/fF8i83d/YdWPc3JCyaulHP5P0agJ7/+JljKmfT1IAHG5raFGmDYg+x/Ka1YixQwySXYq7
jGxPtvk6mE4emeFLcqSUVFdQANhVphb2iLfclGVVMefHBoGwIDHQXe6hvlARbbfVx1+1jJiNel/i
Ozr7Uut2v8oUqWERbpiZmbaZsijaKiIm9HFef2V9sdfdQleNG1cm0ZkfJK8ZWA0BRv+8UWuzOZnm
dDdtCemKjT2Gino8MjuO0tQlorz5c0/kpWjngOqrLmVhKMRpQyjzNUNfEm7I6b/frGfnoTFCW3LX
+0sOZgkRS08j6r6rKpYaTHhE5tmDVZk9ZVUwrJZGu8GMOWAJtH+haQhvm4CoA9BkuQehnv6NTnJN
oFiNM/5ruEy/U0KHGEhgHk8hFhJho6DCYUYUTCeU1HfmV0+1QJBq0XHqCYXeK9lbRHjT4mPcnXio
mZM1QtRkuTLZERja8BRMTxUNyXFdOh0TOOMaHlLAeGIxfjbnvWtkRUf5IhxJ3j3Ag897MX66IDai
3c8zwIt80C+gY/clZIO7BADVHU3ECJrNou9cyP0twHOVsdPsupHu6fDtZ8rw2Mn9ZNsLJWQrcBF9
ufBG43XxB3qsVUl9gjZGuq+QwSYStKZXWDadi9iLSd51HJQst6LiJuZTLXq5Ch3luVlz35v/7oyd
FmbIHRNT52IuAKH6GW7enThwP+kLxkgDgT4NKRXThMNIvfoYjNrg7kuULUS62RhCOl/TXUiBBK3r
d2CDv1mbrlAvcdXIYB/poJAmbyXj9KQoJf8TAhNuuZzdyj8XhtawqgtOfXscTwXSMTKGHgRGlcnJ
MKHud0SX9NsyqLDe+bf5YqzXyxZ+U37/lppsP3wgPpYH3GOIQiEmPz4cuQri7CKXer/De0UcmVdk
8kmGaWc5uEbt6CfzMsaSIcaDflzVDhvSCHbcDE9qhaBpOlFIXA9de7QRYKJZW0BmF+QEEobqOsp9
Szmxazz2ThHgV7Yk7TjMElFIT3qYQiXQJA3845PGYc677B3Cg0Es+Od6QiNLCncubi0rY0M6fWO7
Ysib6/buyrbosFRE8PGhyomOgCSFWlBLpPYxomrup2LySN9KMGoH7En3NvwcPXyZc4vOjugdLTYW
LqY6gmGXx1F0oDHpe0xvRmlSNr6dDZ2eDmJbQK571mUXLvkC1FdgXEGrON90Yx0o4YS67Eahk+4f
r8lLmkEKsQSiyaLLTupKnvXP2+uYkhyUSh0iCSQ6sBCfkQP36KWOdQR/weriMktRLtgOOnlearJQ
9Ffc3cKO1pW2hcl1g0KKqDEJ3OrniN5Ms4tGLIluiarZrmFZOVh7Jyi0YLxSQe7HFoOHz/rJim6A
WRDCUSyytVWU/YEgbHE7Mx4tNKRwO6VPHp2rNzM6o9X8ZSOyA5bnK5hV4oj3o6OJeTuQJkbSXBID
EVYJXlfMh01GaUddq9MZJIVtCMEhws6NDUfskbgb6V6CLOABqNk2y3kMhfyeer1obG+mJVRGP2Z+
BM4NNIKrEkG5njjtlocYgIFuCh5qwQj2stNmoBsVPk8nQ5+cCpnjRPrdWxW6mskKr/jZLr2Gp9uM
A7WghIbAWNouJ1i9OXUis6fgSVf55GZ9bS/EwYX1eD4SUXDEqUxiC8i6HUh3WPX9XIa+AJDxY+SN
JWWXlSGIxlRv+inZ71tyPfykEEZ94JzJQcY5TZ//5pj/ACX5D1eqX5atrXwoqaXP9BVR24OHFMJM
soytQvjd19mWPQXAtIpQaS9EHgswnMfAiu5ot3yfa1U2osDUXgIr236UnlZv5/vaR79/cer4OU/I
uCx7/8Gg6aMkW1pg10/j4RhiczUDNaHE8vjzktYtc0hh5dZAgE7c6uUYdzrUmTKgurDnBnFWoOKf
0a2ZCHfIRvNvoTgnVfrFN7eiWa3PVag3VAKe7/i4ZO6sKKv1+g6LhkKB9vEtBKj0mdIDxT83Hezr
2+1kFFz6iAPSr9eGyoDxgeh3TINzStdasCTfJ48EA/y7Xxlh4woISWnu1iWW3t24ZQWyZw4y3moR
o+cpM48ZllreebuOGPdU9/moHtGHCmpsQHv+pVlU+63MNXRWucDApoKRLLlHVXK+USxLP3aJoGH2
Oy4QY8jn89ER+xF4cAyr/O+ym9QAUvAq3mZM6wWVZO+1qGdIeZPmUhkYy+BFZ9CVzQvtLljwEk2H
1OVTdzypGX43/lT16E1+VtSNIdbyADcNcMxc5u/Sucvyq1SbgdCnIBiKJGHzRqiEu3weDwCBhP3v
mfYbQ8CKUEz4UI3kDIjHBrW7hGHnf7puqWYtMhu9kymDAWDiQROza3FQ1VWI6ibxnUG/0Zxyg20Q
P/75zKpiJ8rVt6DyEvYsXI1XyEc6bOZh2t6fCdHEz0CC4FnfoDAvXgjT6vCRDUURKRHuI5Xg5/l6
LzLJB4M8AXcvyqq72eyfp2/nU36mXjjKVAk2os4glsy5qz9dib7Lnp/GWVeGDRKigp6HNd7gX0wX
DP4oXFCbTFNJQDxx+KINvW9tli2VaZBAZZHeBsExbYo5/po/fEE0x1ZLGAP6zBb+NuR2aW772EbP
0/bN3JUAFq/PNzf8YA9yAgap8Y7DmJizkYLgXCog+a3OseY/xKk1UVAXwtnip00b3xdGR+wgc+Sw
repIb9q9Xm1VBYj5w7plnPKk5B/b6GsOKBXuR56CWtV52V4PG3nB2vMdb1T0Wz3tm9b//QmBX7x4
nUwqVhPOC0MXjcwuXrOjoSAL8YZnx97c1bsQTl9IRiRy9m5h6CzcEhDgYiocK3g9J48p6nK56sve
hBJ5I2yvlaAd9KuxEescHKZLh2bnTKGH41hRhbdnvXKJuCiYhhWDF93jW6s0uJveOj9zYg8dWCWq
9TrYTUTtOeTVJzqHx4Xh+nm3tBImN0wlE1M168eeNylCCtRw4pucbknDq9vL2DjLa/ivsn4vyis/
Fmac9V0YJZITP2aRtBHZna4omwj16auF0Yjb9iPDHQG8yi/yKS9zdt3o1mOZuiHBJu0KWAIcaa04
4mFegSDidAkN1rZymzGSH0hoRV34N1oOhBCjsZX/ofSN8ynhEVC7/DXO9wMryylYcIcp1eRYMpUZ
zcBC22oV3jgKKoMtr3O4eW48SMMNN0HDTNKPEfjDOD1QlBvGQ1NaLLFlfXH0mP67CCoJmpkoc6uS
JmRo46N7dVsfTeGxlsgstbCDmM8dYVByiNqi/sPqzNXW9dBQym7dhMzsqTWpPauRgTmffmbsbqcs
9b/lvMq2Kxsha0XmHR0F0JlnOeqoBA7aNFpGD99osDaRN9puSolsLTQsAoyhUuJMw0nvZXExRp1X
P4BiK+Dns1fUUaJd2ibxyh+Ubeh+D+pizO/27edYo9JCfjG4QnkPdMfe97sjk07fxO7PGPxSaBzi
srL6MYZ+BFUd/kUJ3nOVnpvm/pAQRy8L6ws88HLjumfYqn7IwUAKhUUA+TBPa8zcx9M+ruwbKu9O
JHzp53mux6IYWYHI0wDdcJtzk8gEAgO57yp8/QAWiMwiMJJPL6BsXrKtpPUl9lcRx4wg4x/+N10m
zW/DRU2I0IpzjAtq5jiUUaHwT7DvSOz09gF7/TTFu9HoKouEYZs7gEE+7o9sL90FwukTbWl0wNhw
zJcGWaTz2F0L1ichhTFsdW84q5+bEbqibb3UqmDR5nvCL/UaW5O+o4/RskoWyhGx/k7owWG50DaT
qGzNQv3ffk42YwQehCIR4R8+L4oEtkmSOuvHeiJhuJo6Wt4Lbf5jkDmYwbLzqLnMxpjtk1Smhbgh
G65MViPkm54OYa7YQXS8QSIOf1KvNgwkD49CBJDQ0SN4kSjEQK0YXlfuK2lfGWLzubU63/sRonVC
FNHX8H3Vtm+vBfVL5FzAs5UJhb6icSy62pwifhsXx2sRPtaKHcqxlCAXvz8hg4bhDFloJav4eeOY
z20oNXoiVwlwaj5bzrkwWrcT1vTVN8b1cPTYrpLk8Vf8e0mOX7J6wA8qpzV2+iOzQGZjZq7Au7pF
6iknebbuFAz5aEivvowhA29JmxhWj3v2t1SLBcYm539YisnaprvfOcqaQVIj47SAEjTHXvPcUDwz
gP8BRNLB2qPuuWRzHf3xb6TiO6KOrSCEXcLHvoELMqhXBfR+MEUgwSpcgGBK0Il1PPQE8AMeiOXN
7rzD8bG8FV8J6F0d35Q1mpArsGPHumagBWSO0Yf11oH60L3xSWGOi/Y0/uNS+6owSEyuSWobvABl
zwiDZnLApraRGjBoPTNIwZSlKw+UfdtdoEuHid+s1QWpQ7C/Ukicb2mTLURZifuBZedJ+Av7OTOf
8QmYAVlBn85AvDZEOa2uu3fJsylu/WndCyvE8r6m5+vIcFWlco2NfwT1mv8c/ysBXcovy/Rtj6tB
9Dbr4iRm1VzhY2iDuD2vz0gQ820LIEo+AvPG5v++GUCbSjo6Jey53AtrBipXc+jOE/IXLlfhhcTT
aKbOV8DFU+1cABG3KMKbHQPDfEFH/CmX+npZzNyTZaUAVfQZ4lWX2YuY6izKFevFAMIMvY7/xdgp
4vMPDYCD3SE7XLeuo4HBK5djgxYBLgshdu8YeTqzwYSERcyAo+mT/jGNBvRLDeHjvDKy+HcPiG6h
5PH3QFbFD+uI/8Y4vYVp1gVz3i5Cz4Fcueb0jFLux7gp8zsNhNrO2eKw2a5qMLAwwWRjF9ie9xMN
gSdqzt4Sz0BWjfp8QpZgpyWUlajqazbxiqHD9i62I/W8taFomA+3OL4pTwZRKMYDVsIe+ZlaLRmq
DhzGgnm1o5g3/IXbP5/x3PIpLIa/iwlqyo2feWm5FB5VN5ful3htdcP3rTLoE4vRTVNOKBpVBvjQ
dl7C7xGChgRr5doZioDf73Inz9e7mN7xEGRZmu63pSWkjYqOTGeZ9P+fyOsmeLPYDGHBStHQr8Ma
7i/72dtcMC+K//jJWRw9k+eJhNIXywTd5Xl3t9+V5djfUEEA7eV3HAo9MWqTapBYBQS9Zsl74NQr
Oz8TKBJCA9moJcILsFru0SEvxNjYNls+JyeKjDx+3hELtAMYPTrvBon/2dkgnNX1iRVN010dFc+A
9pQVhon+m7UqIxhCl+S6f2nj9r6yyjrLcUABDFDPQHOu/OpHM5zV2vth6HylVcJ5d/aEozFEIcxy
YAK4ACXkeuDIysLkbcQOKlIALNjSRep8u2PUG9LRxkiUmEHDbaZKp36PJvIhqORJQew2PJz6a7u7
zNPk3d2UDWTnn6vkUJSe0r6rVoNZfOGhFfkJBTYNjnZ80cOeCG5RKC8uEoXZmJUaCfGaoTetCuWl
q2JdWenyPcPLLQRFGBAIJHm97G+1+GwaIVZk8g9dYGtySP9KNLgRxdafChFMZu0sc6QXhfo9rd6R
oO4/17U45IW5hpLiieVQde9O01z9Zfyj+k3L95S/1qiczNfxkjIZii6qwVE07fqUkbfOk9BVJPIn
OD65JUfhDzRQiKkNUEisK1GAi34Z/Kb7azAhviI+57po2J3VRmfvQmEZ+LC7FHQeG3ZI3rthPPZa
5vil+tQQskl2/IJg+oqGte5RUkFlyW44/v2C22eAlhISQlYUapYAN66F9DCbr+u4n7hAiYfNa+2V
uVyKseqDQTSBBX6L7hI8cD/IjQ+imkw2eQeFYLGLDJ4Jr3ZqG74+nR9oCPWg0+3cO2cpmBlgL240
01n5+YkYNbWsDVLgaPWqe1NGKzsFoXYpsVIP2hRuMIQvTohyccYq/AtY3mbyCfQnS3+fSKVZ3fRe
xs7GHXM0DTWPVVrLJgVNmOBZaKsUS0ml8mqHG6zwN+cv7pkZv7m2DxHD8f7hza8eBQG94C6b4ozO
23DIuZf7itlUFjN0yJMWG4N8qk5pcIJZbbF3nQRyEmHLaM8eYqjyDLkf1PUavbyWMmqwLlBri8JM
cf9UsKlOCH2pd0vKLtP98eRv68RXCIG1t1ABh71fgIauD6mEjAART6fZfDxonFndTbtOmNy/hiaf
iMvd9PzOqR9aCZx8LKEeDjGxu/Ht7KyG4ZUCvs1uTvlerSDc19e+H806T4mb1gNELgsmOjwSQwq4
M/8zfDSXvjWUKhwEOhqgxKwR/4zAtz63KweNLzbT28nRAWjCo7imgfKh3gU7n66i0DXW2UaYbvAN
1bobv+74F6bJlYROb8jRLN8GEhSgoleMj6M/eg8fMHGiAVZXHBPUw5M/L64u/vaWW9hNlbjFKlNu
AVSesyZ+YjxZYgYnsXfl0FjacRUilsPqYmdxcIxP6LNZFNW0Gs/89huAurQTjybSAUdHEdM1kjWK
GyrK6eh07hFqEziqDicB/bSXqnAKi+Aj0i8eRjhAC/hCPsbzF6jePjPAliG9PiGrVHr2hnmXAL0T
WiU8ZwHPahbn+XmDLlIYNkHwU7ORSNBX1uWAQFKZ6j7VFPKCV+BLkQmMdVA5ZAPdM1nqG/al5zsf
YbxhRTwkRuVJc8UN4Zaz0z+jcY3qXiGYLC7UoZjCXvA1Ziq/vnfcCMSC6xoLOrIeN3sQUC41ogfC
0tDGKfQ34utP98DrZMy6GJGwICVTktX5MlG8FgQZdgxFmPEJs3C3iCcfFZE/Az1phBv8qeugms0t
ML2p164yj1/RKfPWmJ1IgLIJgNzhP8CwmUh6v9RnCINmbmbc/mX8213HzcG3s5G1706ZASc7OutZ
QbDquRfZHsyfOFj+LRutDIb74tFaMI4V8u3Jf81se+abXpBxiJh8zSgKwgDYJ79cbjRdWM6NJm2k
PhymKfeJKLcjRa3VKtRiXvFE9X7EDiOyWd9TiUfuHxEwwZbNBW1voeZeQVOu3fR7z2B0XqvfffKe
yQosPYVRKCcYrnTGr5qey7YLzEBHSP71p9FClfuPPJndrH4Qg3ABSsGOahePD8IWbK1dbctyxI0i
btfTgyMq3AcarggwP4L3LTBfEnYFG/j3IxPEnH+vedYGbWYVAL168LMrBsf9C9lrLz0I7nI04ZXR
AvXe0ICScQS9/PgzAO7J1gjBsnHhkA6sY+53rHLSuLGeZ2F6z3tPFrCiOe2hnoDb+qF53/VLAiSn
mCLOCZQQ9hBkZVIE62pJDnUGTF4/zEcKEOthAImm/o2gRQWquezm9JVUO73ZThZRU3PBT1VAeoAa
rIlPurh/KS+ZnB8gnrnGHgJ+5NOd/mflgv1aCobciv8dCQVpBZl/eyMKR9VDTLHMf+3sINgBnUz8
NVp82mZEGQg/7ZUGyiQQYZvxUfeklN8dd2BdzYDEEvMJI2utVTCir+y8iRBUEfhbdr7rrb0pHy08
qkqDHAO8PrY1HjzsIXJIj594finJVbte+7ygkMljI3J0QIegGfTldbT1QDmBa5tP7kZMBxn8OzNR
ALzx3BhD3Eh9vxZyzp0xsU/fb6iGvfqX8IGvfelPGhAesMPtGPPgcEqz1iWjLiWCibNxgWahqo/B
PPYpGxs2tQz/wGpyjLF3Z2naFBx81MN6AANdWdxMfZtNPNkJUXJMhgNi1ikHurH1ASaNezvI5y6Q
ku7Yojyf7l21xkxYcyI/KjDKxMEb+rbRVIlI3b/k+JGCc5fW0tIumapSVqyakGS68Y1gKxZmGBgx
qUlqQvYz3rGK7pcpIJCH94yODbBFRuwn2O/Cfze4yYbKcFWIqKuLSiC1EgflNPCXPOgj356ESyo9
AQ8RQM8il6MBitM5WioTtUMq8+t4fNPiN8mYaeh8JrA6bho7t9WZ6W6dAIBR+YCb19WODs/vyKlN
BsUKg/vGUtWalsWIf4Kg2/6slLnZYid7Yt7G/72xhoRzxdphd6hM7TLeg9cJmZjQH3nfYYTdl2UB
fvOeo36jYKJy3BD+emT5fcyXVN+QYdAA59XRWsdyrEIN/AHOknKLG7hkQ/iCkj6odw+catby6uXv
UK5gwPTZ8eYz+jkvQxOARvngxtqa2jHXvc5rNSrCxjrPYs9T1u1tLoi240nPtNBcKZ0aRifXuuXo
A7XxPApdcmppUW4cwXVnhiiM5VTCTWDsgXCE30sMaQlcXgfLnyXYkF+ZU1QZPAcBJznsrJY4O6xM
HBA0kMbHqI7hvhpMbxJ8xt87VrDXzhQiu4Ssi/6XmjY7ZwiYcOD+FRcEy975IjfxXGEAZNByFPrW
kBYacFLKDrm7w5WE4nhYd5wt+qa0dAEWCE1J0xFwH3ttQ7uV/5wjcBJqj0dAUn5xCuuc88g+NbIr
SY9GEe6quUiyV+b2RB9tJzOe49KkYOS+TsGHiegUFAWEZCVzs+aHd+bCSg68OSRryBuLNLl50laI
QQlYoT95buy82I7UAd3JnX6hxEQo3z3djCyL3hMmK5q1+r9xkcSydW3wKtvycNc+iDHe9IEd5fOL
jq4YtouNWl7quA+IEZLPkxWyr0j0hISUCIVUcskXa2jNoN6IYEB83ZgQEXSavaG+xko+v9kl7ZwE
pcV8R3dCvw6KHF0RZTrTSz3H+er23o/c70VzFcUh3CNQKfM1e0J4URoUN0IrHBnSFougcTArThSB
i3ql4GBidNuSTZ9Pt5xECkrDqew0QWhKnhqwq8fULDhzd1hHmJnnSI7A05QsAdMTeNUgVWd5jShm
GxHO3vspFzY2paPSBf8EUce0PyPb28K2mzwXaAFxOGy60t5mJowKecwp0NkD7zbJM2sBXInERN5i
WO7xjer0VgdU8BCv1SVKiyburoyjibOw+wOzlyuZF7YlB1KH0/n7C1Ff36l9g7YzjUNPdy11wnGx
69brnVPC1wHQf+OIbrnA760/ggXMajz2tVdfxOYJ0z84PvSOqP8KuPmgDNNz2QimxEAzqvNJL3zf
MpO14JN5yJhkt6KrszQDFj8JNBJO1MFn6rdncPEii+ytkPvrjhfKili9UomBgCClmGdj6m6qZv7k
2OV9kZLA9HuJvJVU2QRiWXJ8cJ5YMF3z42ev06TCbIVrd8cFcAfPfh8Y6iUmjBZ12Nc2UrNXVT48
moCpDFqs0atEZ66uKLNUBUv3a5nBrac0cKabuvTk9ZYTUxbJlBBnAfSrvyrIEffV6zYbmCZRcrwD
LImsZbMYq1WwRwUwignvem1BSUT9Yw/nMGwW1DHFQZvoDEPY1MAiVafbwPgSs9MKxpDXLQfymGdR
4Q8al04cu+1rG6VcVLpssElI70rJLTP4OmbIAwseHRCZtB7htx/zZZ8yONqKFIuyynKwr6So4ZB3
5loEiMymjhOtARZahipF887WGuIMxxP2lnvWGJLSA3u4yi0H2Om9kB424pW6coqFii1WSdtaJ/gy
iDqDMyX9d2AxfRcCdA7fqMUbUuudsvokzKQyAdLwPH71cF5wEJAA6powi7ZJkt0+yEYuoQM5PUdX
m2h8gbwR8KZo+ZnBCEjueWQCQbcNGh9r9msKM5ShvqEeMKxwKUjLPwk+MnWHhFb+rguiavJucePv
ESaHPnaZufzpp/oxR9xX8WebWa+Zyq9kDMZS6NURgUhIC1yftfuvOCUvra8uxFb3OrirKtXDQW8y
54OC8BtA84cToYYJNA+nyZ0BuNh3RVPNZutNf2VizFC8pHFGCH9XEfu6jf1PftT3hfCW5E8wNSYh
fKoFnpWG81kirR5u2ZuiKz5IZCF6J04OkZRco0y7Q0sHW3K7cPWtfuIk+n+VeTybh3IcOVWe9Ad0
gmetOECIYnXTKQI8jcpjCYTpHpS04ArEQ0FyGWowv79oGD9jzvXy8oBq9W7UqDlpvmW76hCIZkby
EggrzH1n+Hsqselx8JeRHjbjq7SbcaEfsnXnm8ntxWvhhDK1jOvR7z+jZmn/5krZkJyDmXMzNnr7
ZhdhVU4c0HNc4Ng8iqAY9SUeV6zfr+N7ReP7WbCJoAQEoJYANf/HMCq4a1eZP/AhU+8ZO9XCuC7H
tbQpoilWANc/So+DXJksL1dpPrOU5t+imTZ+NDUqpmIgq9ojZJc9NjjzAgj8I7bvynUDP+lqzmv0
WxwbapUmAO0TEMPIxPERZDDIkuxiKp+imHR1JiYxL30ruo00lby462gE/fcj2j19emd0aPxkN7bw
mZD7vY8ennuWQAfYAtI3MV0vTamOh0dvJDPFvCs+nibAzLpkdfzScDW5ldLZSZB8Xg9jfgWbZsDi
6+krcT9xUUBk9eibKa6DZ7tQpFbGhj4rW7dFh1ECJywwcGyO1jpdqLqHf+Cm+zXzyGcp2U5jSdKS
3ogKMj9Ws28uXTN7Ou0WhY5SNUKzf25hEt3aK1vp4074MpR/aoQS9FW+ve+W/4zo2VAM1hh5fpzR
ZPxUF8NHz9U4PlL3rqCrACb3+DN8BcjhwU/9NPSJGSbMeyNPMKCjkstYy/Bz5dIl3kt8sEirZz7x
8GySQmfUi0BAHaUmd2uM6klbiW6uC3mfKuD189qal76C3PdSZeiFQJDS/dAvMytFnFeAu0Yd8Szr
Lsw2B3/Yj5cmQUALCM+nS460sE8MI37XmvrjP5s4pGRXsnJb6uQwCb/0MIhLi+/yEYj4bXWR/FjI
Uect+2SC5TFeu7qw51E5ChhRnWxo7oauzagArbVjsdcLQ+5gZ0qzzMHvrvBvoEG9mX9+Ew/yz+dg
WzVDPc/Jf5hHTQTlTV7JB2rejEVIXw+JyruH35KiQw9+znNmA8OAOMc47uQsDfQpphsyubQ4rVMn
psBw/X1E8gQu+GNMPnbIwVumcShuaEFxHS7Gqe6ZGhAaQNT9NV4J8zSUfTtRRVq6hNxVOw59zgNM
AVn4GgD84fiJgGk1J457F3gp5OnfV5SadstSbvFT34KmYySrmLD/qjglMWUzRwngkLWpSvj+n+Sl
uHEN99cQxFciePWjtWoP8ZaCJN0LNd4a9aAjbbp7bYPYk94JTLX9Kdd3JI5yw6aTKMFhdVUh6wXY
tLLi5txAC+oftnzfOXMcAJEjhwkQwiqHcjCTdLC7edOWIQWOM2mSJT9X17DTGGWcBtKXes+27cFj
lBm25C7dYMxhjr9CwFnCci/+QLL0BTc2iBkqUNaaxSHrK7J1a+iMImZfdVy66gUtWV6naRT9w3H1
ZsXsBNNirncdvA0TOypHE8tWOQbC1FxU0IF+KtSQIeeLj4nIUB0w6BCza+tgK0VVvIVTKsSb3H0W
2zXzqvqZceGkCLch0Pl+88a4tGQh5VJ6FJlOcLSoDw0gKy6WOHo5Vj9OD1bDI9zPMilqZJKesJay
OWtzok+gSZXYG2P1bvXrQjnmEZC5QNiqcJJKAlgiOc87sIDdNK7QOfgh0V3/AW4SezyNNBdVjpXP
DV88KPJuZ1SWvaJ53BmFB+Q0uy1e+XHNL48/WMyKlPyjLZyO9GmEG5EZlErYjhkva7oLly7CujXw
hi+KCsuLGaX7ppVDLvLsP44eiqWRQ8YU+S4i4jGaeAGi+C6/KgP9wYV6jfM3TeSnBE/dvk+K2vrj
biaF7081YA/jpsffNaR041/uqobbNF8m1RZOQxU9ZYa8ZLA+Ob+XiM3ay4Wvy0uEGczzmDr8JsRS
hs+DI4lIq0BbuUMYD0UK5wrsyolKCWEuOFC7T2mbD7aEKdUtyNNy31dW56soiiNxi1os8y3U7/O0
oVbf1rkMWGq0o354cDt9aGFqpWqJqi7Q623wJeoDozE8Gnq8uuyIXQQpRW0EkmkFOTgMg4CxmxTc
9jAOyWwW+VV9olVY+qY9xjZ5aFLKL2980eU7t3CuLFrG2oY/WnAT2YZTpDsMzU04Q7TaCFSn8jN4
dhGo0Zi+BFNCB0ddXfQxSJiLCmkEsD8/T7J4SdI3YMCkFYUI4LwT3YR1F5O+HsEeFMtQTeMKqlOa
ZpcjC9xCgW7PVTdo4wYFcovFRTjzXQocUWdowYJVdnkd423YAx3BiUtX7HwliUbfuCkOpARaKxpc
gBdgYhtcgLaztHDU/xSOrU6OJj0lT0P49SdX9T4CfsSHmlBTlM7G9tb9AgCcYPqgJgVoUiZY7X6W
p5e51++AwrONnkVc+GvNSBmpCuqoHABprffz5JLdZ04J9n0FFJZFVnLssdoK+PuZqSqip5G3qCNe
dDKxOI9FY90+i+upsgfOTa0McyKgdHxjpc6kSng1stM44Q0O4l3H7O/ErSIf+3cRKbrTU4UvWwYf
VXIdp+4jyGJwskCa54d5lmjGZLhnFueLzQ+7Xp+8ddibGAfuglNcBNehEDniCBjKc/v8sFmg7M9x
UMxBON9opjnjRTmGp6to1iLynbxPDft2QDUMWdtYzFMc3zOtXTQxVErVSJZ898u2kh9jY0cRSHE0
B4moK92XPpNmrfxVF4jcEj4GyXoHE1mjgoQlC3q6bPQYDpJp3jx9+QXFBiTiHVlEvuLA//ycmLUA
fFheARR+nbaJH7JC1hQ1ezfhjvxhm84Qs3qJpwTEa1N4NOzFuXADHw7TScFwA2f6OCKT15emuYI3
BD4wE3ibR1wDS+CtVSXbJC51k3xo4nbTSFBBBjdeE5wVE+NmYtiGEQuDz20NGij/DyVrWlXjoF73
O4Q8VA2AZWBbqnTfuFcKALBkV9rZih03xHSJuMEITfQbYi4QcJe5/x0ji755gM0yMLXItz7ytHiX
m2M9VaCHVD2D5IiD9XmRkOTS7ZbiYEq3/mjABODM1yekMu+44u6JaY7HEb4ElTOGLGhwXcjcMoL5
Tvc2vlZPei8onJ4/y/ZrLoqU+0+m9013nuvyFrhaKOozi7YwPTgGhH48c4SiBKgS5ri3BHysDFdj
p1YdS+cCkrvDDTPDX5Ve+k0N/Cmetbe2e/JBNuR2JUsqz7lzsxLWaCF8sgkUZJsQfLufSOv1RxWW
g2TZLpr/VpL7m3ADAM7oPkQAFNv8QFUgg7/GzdW1MmkqDD0NvnmkBLaUx4K1pLytY0HfjYl6JXt1
EavdneoNNRRq+WOmRb7A1kB4lSLcQLgz3R0eFcn3YWl88HOERuJxjEk/JoZQY5W3aRIzKMjUHoq4
SJnrcq8Z8CCI3UWG1r1rFU5q1g2RnzvRNS7nxdbTyB2TeEt2tabHaoAl0b5okm02I/wznk4Mgw0+
qLyYSujIQ21orgOU6ccbJOzIFFhXNzlwx9bB7112XMD4mEW9i7Z504PW4SqXBc99rEHKsokvdPka
jU+6bWOuA0XHiDMPQ5AtucVFfRUb0GgJCKL8bT85n11omTCAWQxMZ38EpTJEwIgWV5WslBgkeWuz
fKBfU6qRqU5yLXzlucWhwpEYplIMiJ0/2JpTUOgwl1d9kNsfgxulWB612YYbsItGj6+lg1z8I1Fv
MbyEJQXGkF1SeaVrWoY9dKHcXmRE5qADGq0lGUnFe8Bsr/w8+AZcaYYhWSr8B3rMpRdlsGoeLQKD
67/65Ygv0RXOAFeDuBGn4DyBFUjps3eAmlt/94wreFFx9/YDf1qmWftcrBWdYifWC6nqgsxV6VCG
VT/EmE+EDuAC22/3BaiHe3awaeIbjIFABIVHc3uXetY1NfcoQC+wCGW/+WIOjVkJVlXGZzTWPrmL
FZgo1B/Lb+/5dm1Xm3npU1Y2mRxxgKQY63qVAwyhkfsRXQ84NesG1SVVrw2H0uEzfrB3+DfGJJmb
ZWv4SGbriS6GfTZXAphUmsVn4Kwtwjzcp8ZWr1CqLNYv/GnnANRvQEGPT3OooqUitCe2RyDwAU29
Rdo6UbdSj9LFUx2zrt0u2Y4Sca4ffaq1gkrpyN0lwpc/ioX6sAGiVAXKMb/FfLUvL8EwCNh85LF7
RXb3QjHU5+ean4TMfFTgRbirxxIxbwd1ot4AEtJ34N5O+6vwStO8OvZKsnXgyfmm/GQKFwL9rTmR
Nt4+afMwgCSdnvb/wrPWdwhigkE/HxDz5m/XRXvZL1yLPBRgHUlZ9lw4Oc1uZNeB78VF96YUSo/a
DYULtFfvaVAQfX+zDsAUhIihiyeZYhfIHphVHoOK6OmImSaL1HTG5J8Ia83tbH6ZCz2gN0LAFeMd
ZJM5K8LrnnmZZrZhJV+7ig4DZXcm3TDn/cGOm660g1xhttAri+63YS2WQ6Yk3FxH+8dFgB86lUEq
zonUrtlK840KcMjW7AjWdiYcmd9sUySr3fIgyChM4m0Xj79KhuzyZH5chd4Yc9k94ZbfkI7JLdQI
QsE9fbD4g2lvlzbZbYWEvh6iGoIxuA6Kqj8RSHoX9Eg+WD3jj+lHLQgZpk0eNl4SLusIR6PyAuUV
97BP49SApCLlBPB/o6MC1+Wgu4fRp6eXC6R5iBneR+8HuAbiiih9ILWo4cQ7RT9Xtis6uMCisUaO
uzW4BFnYRvA8Azn/d92bPLzPuF9HqNtWtTFOIPPB35Qx/YG1Vw1IukOfjUHJYE+8MfqTi5UsjX8L
MpT8mqX+oItKgaarcFFkXn5+J973R9Ya+bgR8Pqsf5/arG9R3gCqgCeeVZ6rbUF1gGe+cU0GtXhj
XEOFtY8t+QXOZkAE2zXh6DXOinqjp0J1ANQ+a+sHmqo8Zw/XrLhtg29+FcK7UHS6y4Fro4EJf/VS
y/d0fje2M6cZU9v2V/VTKQOHs1JxI3XjsPQcYDkgTkIR+bkwzMEIGDNTPIxfJN357HswOgmmkbYj
rSDjxCxkC551qF/Rjp/UQRHdg9yFkHq/S6J06CFPcXggbJbJigVwMPsvGfEWYWLZTTCDDjV3EuhQ
qSncyVsAHyvLHs6/RwGCMpJrs4mQjdPom+PowWy4rV+hOb77urCtkFbiVhHsV+2gesW99EG0tQtV
70OARLt5iEomgN0hLRZAeRJkFcZloaLzdWs7FnWcJCODGp0K06I1CjYex6IB0UCNy4cjr0f9Xp/8
qnHTVhRNIE8zlJuOysDUU1mn27DQNYpWatdybBZqpDBwC2kD4U3L8YLYMwooCBHKzIO54pB7Lvz6
DxV+hQc3Z6608Sct4rPqqueQR8P0eb1p00kEunb9vbBAo4XIKEXbkXvAizQL/wjU4dSEi3BH4YbY
9WB5VXrLelvq35o4wQMXZmT19cQE79VL6w3mo6CA1y9Dhc10e4jg+QsOEkERAWxI3ATIf471Na11
34znAiouWcTFSMMt/4R3ZCGDv4OeFje1uaXvZlV3sQGcmUVUvVgY1ZhBDNUCwl+J9HXokzDP+hwa
D3a/6j+wWHqEg9BLDWOYfOkmn2FznB3yVXTyITK4YdnqNyMfRz/HYHRJKs1w//aBEH42O0kcq1Zj
/GbbfH7IzGf1xt3g46G++sx+q1vc52L11gGh2QAV1WOaVYj7N7x99xwy9ppBFkw+LG90vCLoR7ge
tk66aq7wPXdD2J4iCtd5ctZiaZ07Ez7eYxZLmHV9D5khhOO1aASxLy/smv+YCqNoK+ugj5yqNvNN
TthZct02VRLTt46ygeWrumSFwaw6qwdayUUBS0QfniAugtak0oAdVPqx3/37nF2ku2Ac/AgDjGRg
daGCrAF64VE0ZUw2NPtjnBLNdCNcF9J/gc8wRJl5BQyWgp9+3ga+W3IsB/Zf6i50dd/Al7H34u0Y
JTWexdMhOfUEz29cDCg9bth0Uc/TzJ2N6D3P7IPmCcqMeQv71aJ7KmGSBcNUjTGC77GEzAeGc1F7
BHDKtbxOGsfR6t6IwSW9RzfmEHDYb/Y8OSCyA/+/mihy8XwD0I0AQVTgg3t8CihJuN6mwILJ5l23
bBe71KTDDZD/NUcRVNLB29zMjmbcQc9+v2BhFHhNrygl96NEjRrq1xuU8kICCn0D085YPp/MTI4Y
hw2/5WVFzt0Lgt2sc8NiO6sVefzIJsl4A/fP32H4YgrAFP4X2Yx77K0wk7baV0My3Un6DBrx+7cd
UnaaG5i7yO9HFAxIett7y+LMGFYiMvb7auymmO2pGbYDQUZ7awbvqHPgjh8IaS0qWi0c7CyDZg83
UKk+ilE/cfdRnKCjEH9dXZFhM4uze+c6oNAaFre6GgZl1kaKBRlLcjJSNzEoI91GKDloZrBB95Br
Iyabw2JepdYW6/jPNbssXwI5oSdrRJUukbEyhFTHnbXtU78Dfo9r/1FLcFAYsqnhB/xt7KoJalp8
l5FVA2h0qrKHq9G2DV7hcFPSnTt4JSg4fXpfxkG148zhWgdLkEtcK/XYokwX/Rpe5KizFO8Ht1cH
ZEd8sJTCCqy2rwMsXGPTBXpxHNXD+wtMC7VJKD5usPKfDCeFC2tdgP+XzRk+XjuN6tj/nMaX6S+s
I81vZvKhXGDrPcM2pyZj2S2z3BkLt4EySt94ovRXBIUz8DgTzH602yqy4f35KAx3v49wAWyyVj+E
kmI4NkuCRUtIc73K5gj43KwfNm6RDqaRxYS5ZXzHw4+/LjorA33fOcJC7UCxhvu/Q7r8AZwzESff
DYUA7ZNzrA9UwlOk8HXPqYgEQMcGnBa41qyxLJiFGoMcKhJm9SK6SGNBzVokwooX3Jp6uNC+iuhk
n2RxhQcLMb3aWGz9PSPovRIG2eflJ6a8Yr5OEr58wxlxTFXLi5Hi+Fv5tQ0n6UAwB1b2vgzxf3zU
WVuligCdcawLD3NYCsxdq6APf6HEGu/P+nVk7Ba6wseVJYKU9RYLbUxwITe7dCRYNsCE5ZEyBX6W
jX2yrUGMeKSNSgy+fEVgk0joeY9QaW9EYg/NePV+D4RWqB6jygIM/Nj3db3WMZJFYqJMh5VxQmAm
Me7iXmZEUTEkwO9/61P3MZ/siRHgiWw8UU2+Kf61ywNp6az3ZwmqLHmO25ELhGxtaJkA1isRPrFQ
F4WXF8vND1Td/Cpw7h5PGQ9gQV+ra9A2msUKCABlC0X/mK+fpWk0JvQ3Vo6UXkR7ERRdD9vgbQ0G
FZq6aYZhk9Lw5P8k4cBtMokCJRBRNAqc/J7QteCdeuDkHoNqKFawyuH6+2z8cIZCEqlqirbtcFs3
MIYN3+EXER7G5zqbEVnyL3w7iAkUlUb9LZTRXR1SUT0V1uS8rOqhu7TadmUzyyk3QnCQBJ29Z6G0
fF8nV5Pd9WpoAUsNOUKeOUcfMeSCheENOrjG87aJGB8RIOB2GiE4FOAKxS9KYPPvfLhDc2P3f0AX
iz+j+h4uhXZq2g6gv4nAHjeZe/4eKvvFFisx7foHtK5y/588MJWEE++GlWxWMToBS+0DG+4gIL9C
6ncGozPd17f2R/5v52HdXSqiwQg6KoL/OZtt0JDiCzWLhQkyS//G/OaWYFgt/YA1//hevXftrgn0
WRnSQrkZRD+Od7V3KmsMCsRNG15s7UfH/LZiP8Bg/AJ5pBg4TGCA7UtasqSkH6Vra62TvBkOVG3x
RLXtYE3ye9xT0dMG/ruaEVxDo4bsn+8FtPG2hBtviHyJ4zqYFq/yv/munHIcXKfrVTWbNnL+O93Z
VYMxPnkn4ionAoZgE2oDA552fTYgSYbGWXcUYHnU2xHPJIiqRuoAiBppDWWblLOtoJrYM8TUfgwG
Ca1yMpeLaTumh8vRxlzMcLqJNzp1bm1CtWPI9GPBjOVC3f7ReW2nkh6LNrcqBViEf4REWOEdo6r0
+Ywu23KQjjG5hP7mG09WhRVgiM/mpYngVHvfVziMlkYmNFoxjO6bs+GDwrciDmFkJkJKswwAcsvE
F9Dg5Q64jUySqyzPfOq/7bmjGbXi2Px5JB8awtE57Lpl+CjpLQGTEWgtZuOMtYI5vynQPc8/BIZS
pb91bozrh9FKbigNBMHn/fFFEhreudqvMHQj5fcjFZuAxdkMYGYw+jJEwndTOJbSehNA2wHvp+Zi
TWirNWvSqPOxO0yA3DR887W3o9PK9suO5V4DNEpVmNQFNScUJJJA6gLXzxke1Ob+4iUZUUa5dDoD
bylaiEKTkzRSa+n5cXRgPT3yzB7tq3hxv3zY8nHafcnWuSIAohN4Sq+jhPddfcXcx468btfmpooB
10NthhEoiyIB7V5kg0nVjqHXd7ZF849L7J8n62kkFHpy047aSfB+2oCSbA6r08dOiNVuYJxom5Gf
ApP8RMDv/2F1TPzafDAWy7alfNKIhqYPfUOdwQlgUAzehMt6C0xs81YwZ+/CfYaB3/7oOww6sWht
GmJ4wj14FjKrY1pqwMiv4s1dHxsRiDtgPai8kfz+3o+MD3n4EO8Rfj8jRlKaDod/m505bY6qHS5B
2UQqL2q+HW2jRL8/Y1z2t5RvDu6fUJoQafSUMoipRKj3nR67750RpHEunFBRv0d53RiUxB/qxid3
zIeQ1dDeXfOUT/W9i+uB87+kOqWRGl28+L28PEibxVllme1taioR7Jet2e5UGF98vsjYdR1BnKZS
5hHeCCVU3QTuVXoLr9eflvx+vaYNfTYb77yS9wOv0ZacilmOPHgFvK4nvjkZWNbnkajFCa7l1KA9
Ru6P2Gn/OaZY8+UBeFt+evJR94ytsRrA/8mGPo4jLWlNVXN2BuynutEFoRHLHZ9yuHO9gnm8VEgW
NSSdqVk5USaF8lPWr48J7JyFiRpo3HA7+Lc1e8J8VseCEhO4AVXxgoFxCgigEN6UEvPWZnk9w+6V
ImFDDwao/0PBJ7ig8MY+NBOjrLflftUEGhlOro95ZzXFTOccLjLQH4QQsEu+Tz5nXqrg05OftHKt
uStOtOBfi4ddzjYu500E3czqBH68l2r6EutTdbgHeKU/P0PCYyFHhM2O4Z3Xg03rPha1eLbPT7X7
Yuw+x+sk/JubFueSRvwgw9yHO0Ntbnav/Yh5Has9DmMDm9Zk64J/4jD92IxoWxcDxLhioM4gNV/D
lcmJHZz2ADicfIRZ0Zo+zksdEkR/XPbgh3QzEIi8bpsp9D8JpIOAp+RX+Pd4wqefbX7AiW2BuuwY
lZukdExXQ52OcE6CHnRjG0W1Ua3ghwtdAhpqaxC6HJUjqd00Np6h5M2FCOjf0YGxHJ9zy10TH+Z3
zGyHxEta7vuaTzpR3/OMiQiI7erBcPvK1gpBv7bTzIV9uB6sKw/ZXDJrxuMJgmgtakwx7917m8Mr
DrX7u7U/2if888HEL6sxIdb67216ucQjiX5MoavaYibvx7JMcm17cSJ538/QdQjUuiQdaHo0gy5+
AhaYVaxs2BUVBhnmNhzH8Lrxkf+8rKhMr8qx4BYqvpwzLyRIsenSq9mtO4/GkWeb1ksfjxvviSSJ
yTVXPLYXkM3Fgvn8Ol9TFHpwCh2jOWQCnmh3apegOsYv3owt120LvRg/8gEaNcZeDmaPqItQj8xR
ynXVdHFhS+nuVtGLNsHpkksVLoWLPmjAaM2cbgFR+ZBYlSgZkub4QG4t7ERmKGXkxDLnv71lKxik
Yhq0my/I75Jfe87Ha6nAGbVL5MBCa5Cxgt0bpptrCforEhvspVoZ8F7MJiBqh3Tj1481yaX4864j
EabRuRz6/Q2XuYe6ElU2ApvNhrAwSyayE52SugYO2IDa5dKhaVX1MS5hA/eWMIMVTlBuoPm6/gJR
WSZp1UDxnt+5gD3pFuTJrvCkYaAGth9aF0oE4rvm2ii+/sVR70BKW5C3l1IPEPwUway3JzLOKagC
QlCsVuVNAx3XIb5dvGyDZLXXG9u7/wL5NQxBpfZwZvXmxQC+88QSY7XJNnjkBuHSYqHxIs+uRBY3
mXZdBqCdgOEHwHUKVt8rxm4cSYnKY9ORz1TGpEwwZtFDgtjd8ory5CSWHJ9IvXnFVjqopO5lbpGm
5G/Nt3F8UH3tI0uBG4nS+ohnhuijDl2Kbiq4nsbgNGEwcsJSFanHmminuP2yfuWZ+EApSB93pYlD
0ZP+6OB1IR+5ACu37oCdP1VPiOm56/tR7vgvTn3oKMejQRFVq+hE0d0vzn/cGFpezxAsa+IZUPK9
prfG4p8Ya/2yVGY5O3m1IlXyZ1oE/jtKg413HGfWX9B+7TUEQ3JgsOy2ZhfNhoLM2eeM7EODL1hF
/TMskHEhJqcoKE+g3Wmy78oi8sVAQbE8tOZkJqShyL44pKPtAvYXPJsaoR6smb8QlhrCOIjrgbSS
vxvrGYHoPS1i4de7KdegIL+BmIyb5I+vctflzHjmLcNMIo0qEHaMiZigWZ6Ap9p75okKI3mB7pHB
xtgNtJAsVgMwezYziCLsGfXiBoYnV8boG1GktLhPXg58EDxSvwftW/lPsJ//OL9M/XxI2Qfwws9Q
oQuzg5qz5aOhLrpuoN/C1ZAFhoobXcAfJvslX4MDZ/GiBEEeqh2SI6Je1I0WCROkBo2CLh253IdA
/NAxiIuZCxqa/rzzeiYETLGKK1lYiORgTQeUmntvXE+nQLpjW/2u83n3ZN9NuVyu2dO1/ag5LrqI
7BU4HSRU+bhiMciIwOXn8EnuQs/r2uwkbidkZtjIayq9Var3NdWbhiMpPm6vQX2dBeAsD2wO8wux
VmEabtFD84Uyq2YLCwaeOWSYEzGrLYLN4PRBGjLNZ94r25Aoky5BUTFVfRcUkkZ71UpD2guFCLnC
GIvToYS0O85UT6EKBKC6QEeB92LsL5ayz/dr+lR3pp1kZAQ159mmfvrlybn4dCLzftDOBrTYslCj
hXbDuW7UNFoYVPqFO3iPsqwQD2dfIo7mZjuLOYH8Jo0Z6w8M7HL6FCNkYjqfwl17n0W47Kx+Td18
KxZQE8XqjY5wPfFZylxGHPGH1QMTZUGqiTY/dj+ye5Ag1//AT3B4Eodyu5Wl/5JxcghpQJ4qagCs
yNCPDxBa68QWqBJEdUVDo8PlEPLEU+HDKaTJ4DdMCuDC2JoepafwTGYUE76GUFTvXGB/NxZhbZnZ
p4Oiys10DpIWPKqlOjtjRPfWDtikmmg2bKJ7+ofj/FNlL/efoQ9hEd47zitRd0Iwtgr0f6QGQUSD
L+CM8t1Ur18OphcAdJ/p/mSTwml7OJGPIGP52n1EhwVyd1dnCPIWTAsXY7QyobZT+Fl1a9EQGQSt
864zgcZIQ2dKO1Rz9MbI6QMw4vCoL7U5gKL6rW6yM/YoV5fE5DmrE8+hMPP9PImzgRivkNj2DcDh
YAlvSeMBHRPF/9Gyxj9w1MNEH7xwM0E8LVwhsrgekqNbXupsUhYDKVeTHhVZyJs3F4qiU6WmzERL
oYcx03xxn1QZ2H3cgzEpBWjTQi7V192oGKFBQnjgRAd/mnf3bHqEqZDFYaWurH5dptoBQc3Qc95u
vCanv/VCKzS75LyuuoHYrXEVeLSpjVja+riHt+Rj7IWlPQ9ADzGgE3jGalFZVQQ3NDxHSxRMmKRY
IcNTREnIZsh4F6Ul+/w2N/Jy5f9kCc7YWpWD+RWhVy/Ah9KgqfzcUUCn0pY48tzzR1EucW0Ms8Gx
JashIzZNAkWVWI1HuRZ/MY1AIXC2skZLp4iTN++4bt2fSfKU4NteUUkKa3r8eQdP2EfyDaWkUouj
z/n+/wfYp1nBHrxd2kN4QfZhM8H1RDqubwkCEkra1qboBj9rdfdMt9hNsfR8jArPfj8epU4WodM+
aG6mkItI0KSdH9VRxO0Oqy3S8zigV7hJSVyfMuDBa/5WWs9W6fOLbK7YwMEKc6qzPyFfEmdEdAwm
iSNP4bIiJEDiiqMG9WyugaG/3ASj4KvP5TOpICsXu1WMRjdC2e3lxQBIoNS4tKW3ym1fYanFosz3
Gs//3N9XIq7aaarhTDhyT0outfwpFvBwJdXsxFCMnBu8PyrWEaQ4jQU/I+PRJks3Q6Q7pQ23BMZI
94+S/23l0ZEXWGS3zE9rHlqGt5dQsD5kgxFd00q23qjc1oPbX6WbJ/CrMxpq13hOVnhKxtYBe7MV
uetzv5/JBvUQIlAeePbveslnS/owtousV9QjQcw1zPJuPTY6LNNoAHLMNhW4UPtE0l7nOp4iHuce
+h1sa+SmtroKzeUMKxnDZa06B1fvv5HE92AYUC3zfJCYiFrR5kkHsIGUti31nKboaYuzwW6rMo5U
dmG5pPChin3fdup4b6wagyhEcfUJrvFOik+gbSZwTslNxHPu4L2hqJq2KaSnFOE0L2Pj+4UZGOTV
2zAJ1n2KXWJoiNP/PDNgzJZVEsoigcAMcnw0Fos4UPtgFFvGuWQT1scMQqbDBVK+fSST6zJYoG34
NUrbv7JDuPxTavTwZCzU/u8Heb7XMDacCAmVqSfKXdK0mJ34vzwTjIcZiKB6AEaNjCmcdK4PfHYE
CkY9ggou9Ml4qo/GEkL6ZAuPtkh7HXYmpNuYu9kExrU0HA6f7rOsh/uxHNtUWyIkjswEVYG21XN/
RpJYEWiVxrkiG8izVt2pf5FBWSo92XWYBbOQ+iIE7H3OGVql7Wb6bFS0hF7k3iXKuRHU5ohwuL68
NsQ8lipUxKMAnb3pJfgzY6ikHOKD8IcW2N4gDqXrKiSAgoJLpkvzWJx+sWsbWJO4KwENyct+VBW0
HwnmbvO2mixjwvkL3B1TxedN/EVvEF7d/rzl0V2HWNRQdZ8Vu6JsudsunC8L6YMRxqFnjeBE8HTk
+A2yKFInIBAgpUx8tGssBD9wpS0UuG5zEi9P2trdVy/uE0jVMNgS7ya9oso0Vz65TXODRC4epP7T
a0ECtMjnRnDeTbf8QsuPE7xvozBj5FyoE92DeuPt4dHRSt2Z49K77lBamVu7sAU5T6kEgNowihAQ
VHxH9MqSBzaPMCG8vmuYj/1RxNyRwJMK5ML9DH1oAWOjeekiDCrPrRXgKXGTiWcijWprucH++m8h
Tzbe9ifUJELoASLUmfue6Mfja+ro/unriFtgcEBqHDrynJ01EKybeYYLu8z0/is8w6Z425pzRl+l
65D2PH5ZGqeWbGEW6NlZPw/+3A3HzYhDvqptuyEDMYKFjcO0ODqZI77w3dsIQLUiE6mAKV6thaNx
VL5s4JidOZB2VhAuqZCMr0CanVLyPLRYpfr1cyw73vOmcr3fYVojTGiCdn8vdj0Mq4Na6l2nWNz3
VZiWKr2YDrdZsr+k9oDNcucS49n3LVF9WmlynDVfmh+c9hgR3Tb9ANiQlC85qCzNdutj+bC7yVQk
GrPcM2YA6eTxY9mCdZyuAVsvv7qs9A3KWc9o5MOEt2mva2a1nZ2jdHM4naw8JeoG0PzJjSkeV3/0
tw4MHYT4F8lhpmDScxwN80VGH14fIXY31vYibT+ql27u8/AyjmCGlnxIDpg9uTPMtfLJxf3Pat2t
w3dvYXHWLUD1ei9sVVcQuwbyARf5Btpa4qW+Seu5CwLQ6z4f0fkQxtpHG7RjX3eURxjRIY6+MwOB
c8aSNp9jbRAJCvNiAgCWV3M8IEjFe2r+ZGmAm0IqfImstFjXqhImmFWMUkMWQCW32UGXT/teiZIN
QMK1Vfh/DZ4DJ3Kso5E1k3iquvAuT3SzzgmmDXL8EHW0fJKp3RUf1ZHQzb5KZ/bsXf5b7m5b8Z6q
++vU7W+wG5N+kmaWLIJBGH4wk3gGbIsEAhmo8Qr+HCtcs/3w1auPoqklnhoHBrT39z9NEQ/3r2GQ
zJPG/khUbwk7RXtdjm40ft8EFilPAnkYhVpNyD4wK9uyfDsyL+PjmJQrUFAeUs6XMvbQRUs1OrN0
LOv5jAbIMgH0CFXE8gjmbxARdR4FBqKb0grkdzcxg+AjXkO9fBq+XVTOTaobQQDLEQ6/T1Vb40Ad
e2KwD0XqfLQd3TTNhrckxYu2Ui/CZsiow31DOJ+sH+tFLaMo/r3QKabBgPNFDx3uwe/UOFYdCCMf
6yy4QmFcQHxqJCjo2gL4Ku1ULRGEgdxIbIYmlesNchUIlWQ7EtWJbz76/Pui3cFW4jMyz7o5k+JJ
l7VKI41MHw2ybSdwMJ6C13h5iCIsb/MZ4nuS5aXM8kwp8Zs3lVbzmhezmhmeRIM735x5uyOFN/je
8S/FnlkaBP9sx30mquy+8iZRW1bguYza/QzRB1LKNV+fMbcH5gLku69nVnlsVR5zopgyqBQjmrMF
WAVQElXi97rqGEGyXOOqdP2xIt5cFGm4FENG6g/q8cv1mBlRBCyLxkAq0MVxdyVxtGsU0LNI5nlQ
Co6hpw7Ck4WAicZDXUVBMrikg0EWwTJ4k00Rtcrl+biImJwapHJx+pgewy08eIU17U3e8glSSQoG
b9hr6x44EoROeCAUlqOsG2VxXuK0GLE14bJNBmlErd5cgshez/IFItJBRekqcMkXyWnArxZ1lk0D
xf8nUZ5RHds2tAl9bzckSQvNTe4T3x7a/efH04tJ5D+cD3RSQqBbJoIJVlbTfVooVQbYjpDfekaA
/CfA6xwLXApDszuUpOAWwz9A3Hid3zW6eMSuR238SdvUBdaV8DSqp58H5Djd0Onq4rHZAgs+lF9m
poYx6kQ+7IRrEmM3M9K4ZYdKIr1ekp4wkC8/Yux4tqIA9xMuD8/6kTmN/L285PSKw6eh+eHU0Cej
SD2demfeh6XLVz2AVGmy4n8AX+j9AIiM5f28Q4yIx1Q1VypfzfIA059VlCCwB+KWE+As+jTTyPPk
MSLxqjCewZf8WTVwiG9K+mhz77toG2KdSrYd8I88pFh7jYEouyrHuuFnsUESek/pYUyL/z4/FqIg
tY9HcFCGwCOe1nogxklwcL1/DY+6VoFWQbUdBqLQqeCMe46ZF3ytE3ELuaZjCs3OVOzYmtiklFIw
TNKZBjzZoMugYR05mIHEYA8WKCGaWnS95qdb54MZE90tXRj12sMQlC4lZXvxqj2W1S1XD82DrUdt
pA4KWnlVluBPhpJZto9c1WzceZbkWVDiVgcraS6AWOA3EAHTWhRHijNK2i6BuJSgXTptqGSJ+cqB
iGJdDBj98qlKRxg7S42AJvqvWuAwY4iSEgtuaORGsFNlD7VT5pp0JD+v2WLnMmd0nzHHguSda9GC
RI/2VjZNAiqDxZ4HJrp5bopc0ZJArvVVIo4WwGfG8v8yANudOcOUOdPhGebUsqczM27v5+uXtqrg
cdtqLGIiSUwfGRODzim97oNsOgIcrwUYteCcrq8YMLVlC/+eVpm1Agl9prc4jcVgDBd69cdcWN5n
Wzhi6ZPBAtU8f9YZIA3J0DSWbzNhbnP6+BmDIHhADWX0C7eu5mRIiRtcuvZgmOELln5EMnF4x1ff
ZbQtr3GrqNVh/pB3bUBAA0Te4pcIeq2VbomKybRtxtcmgVNDuMDRRGvUudbKYYprc7BbhvQFljcT
3w+mvx4wAlI3zNIwU58hF84UFeVyL4+SgiUlGH/lG/vPvtpf42mYQgCaL5kdHrlpnaOKqK6WxQBa
VNb0h9FYzfEBUCI7vEZEa5RL7ZWmLebZwrO0Zq6u4D/BiA30xeS/te633G89lwe9M/IMziMjLMlA
coDbzT/tYMM3oMqyPjQaOeifsGpPRIu3OM92CFAVu/+mu5TxuWBqbbW6eYttlQpNRSwpPS6IQq5I
MGu2ufOruCxzrW8gIGIIiSzNvFfNFIg7qKM7sR4G/tlKA1vxkuecaVMSYcMxgWa71D4S43iLr4Kz
osEdLw4ioxm7BqwkVRLxV0bEuJuHiugU9FBO2vJS5dWRGSaZziUJDY1fBRVcBpWX1/+bkvN4eojq
S/vd6qDEJM4JUcv8u61EPtnNq8U8BuZFOj0XpwB26zrjy+bamNC1TGVBIFCtDPYWJBT8Nj48yZI8
Y3jhQ4x7GvhePtue+3hgMme920DBj+Xjq1EMLHz4l0E8/tbll11SkYM0UnuAytSk0t7yL3Cjr9Os
7rCGQh0F7KLxZPfHthUvIjvyAmvkW53Bt/OWs5MGUBfpVmt98aB0JEnbaImjve9dKbh8Te3WRhEQ
/gQwKTpz7x0xrqY4Z0FEDZ8Inq55d71xLiRPb5BCVdbnIgf7OLsq3h38IYNtf+1eX29MiaR7+jNr
QhNnbdaEhSy/+5FuJAZZCgEWLD3akiFXuiFRoUbDdiU6EjsEkThch4gpoiK8CMBOImpCsDSQ35x9
swOuNSxi5rgLDypyqbjOSxqBS1v2yxPz1vHClXF9h4aiIOGOg0SNRwdJwIQWJjQbkIIS6VcZWxsx
stAdP+ThKLWZOEHpjbMMRtwyO3aOF0//3MlFmqbbLJGPZRuww78MvJTEjyDJuKIh0HI2WhQEh8Zw
jOL9JuoCfAfxjFWjYMAbDHKGp1KVgh3Wfj+uHYUuRq4vvOIY7ZKp8iyRf/l0vjW2wQgckXeG5I7N
ng5Tj5zJ/SamqD8te36rBoRaexpYAxFOF53tcvAyQvd/Fk2MywVsPmN+DyYOTr2KckOruciy0JBU
/XU5jOxZ2PuL204XSXvNNKg6O94W2Tos+dt8JD1lv6ETzsXjTyIJ9qBdMFBDhJI+Joemsyh78VHm
skBIN6j18MdjSjqrvA8gIVPWm+CNd4C+Og1qJ6jszdKkCxyyTnry7xXW6v02ByySLrH9Ph0GncZc
UY5AXaIZslkpdQCY55Vt/RBPoBxey+2K3yJzIylTgHGB/FGOHSe2Wp9fatMy6n/+VHB8hk5+holO
tDIYK9LpLxkJykvK37f2Lxb1g/5G0LmEZfFbQSUCxoaqnXRQLUEEAu4N3r2OCTmD+i0lPQ4ufAVB
M8XkyuViNOFIZ78BqFVYYPjZkVMJEpMIGthxArLNxlmf+I61jGXmcAxoKShHvPfBgn2QylTNF/Au
fYNhmogWgyICTLIdxqnO5pZXEHngmhv2mNgnPzVi6r9iwty7odhmMbCI2R1SSJhRGsGVul7flgdZ
dAl+q7MrThoGlUrmengTwztN1ocj3u7IsFohPCoOd6nOVyEjVQDk9eCrkYMK3oyECw2HjymX8C/w
++5/hZAppJ02a2IJ1dhQF/KmiOyJhb3nF/6sC5/j8o7nkw+zRHjOh9PcjRjFLHPOI4FhJbYYKsgr
IPzKUl5FHZk34MNdF0bhDHDKQuCcpVZA8GeQeBpMsdCG81f7k8wAf5EskBCe4SODZDfSi7derRrm
j1Qte/kZtmnvKp5lVFTj/2GlqyIxCZp+Ua4t99NtLbbv9tk8rJ0oHYu1YVkiKsQDUlx9F5dFp9SS
ohVb2Lb0GXbi6h0Ki8RG8XOAeFbq5d5b1rONfMVUFmSfZcyWbhIpYY7OAQE8HsMnYOM6LhRqBmUA
kJfHaci3Hyf/6/JXQTLNReu0yylgqxYmN2ZolxzyE1/lZOKtbtqOM27gBXq+OIcncuCg6sSOicQB
te6S7WXCmED9Bgm22jh93uw62n6OlQfzVrDtF23BVaIu3bz5IbTGsCnauFr7Qgq/dmksQAhE7AQe
XWvnJue0s+nUj3b9If4qL9YrI73lxp22aplHCBqOx7n30N3aPk9iya5yzjj+DrB6fCk8buBHkea1
CHGoboaAY/x4ZmRTfp0dQi+rjZ7A5b87RJiv/YrrAD4dIGUt2cV/Xkl0CkZPAYMSERlmP7o2YDo2
xabljrs/Nt6HHke+UTzCZ2IrK1lHccdo3WegcsAfhq6lTUlCpoVI75qQcHmwkzBYJ6xZaRO+bVqY
GxOCq0H2oltb+bRJUvMrCpWcv7ApV7Miox7oR5LxziHdrikjuaMO4v8O9r47eenpifdT1YwFoJDA
8ES4uJYGCUk3wwz98f0Uuz9UBZpan9NL4pO+KXLJD9fWgbPqiXMsAOhIo6j+vJGdVaSR8JX2GZDq
qXIXpwJu9+RJEPyIG/jJ589rik0VmEmsfbDscmudjTwPt2UbTiBOnlQ1864RmWYT32ACFoGmBWtu
DPHMS2ZlH1gBkadaycCJEcQHJ8cVUtG/6C2vDbzK62uswi6EDj5ZVre7Bk0+/rRlXp6N+RD2XUeM
egxO/TtjN28EkDX01+2w7fdYOwvplxSvnTxfro2gnqJObrSctqsWJQ74k8DfDZtcZEffvygFUswb
7gnU8VBvVcDYTrC2cTzJl+CnhTOVNwCs4Jsy9oSbLrEHPtIPbCJGAL6Kjowt6epVjWrB7FwDQbgk
VSj/SZML4TjUZvUcCSv1PcxNgR3k2M1UcgDrv5IWMJyFnWr7FaXXfHE+kVfljxzIOsm13U4E9vsq
O9CuAdaPVXQYS/ip6MCDK5shPuxBtzZip7TBEPZNkwJ58DT1fxsVZn99So9nCdRg6Gkc5NZJALA7
HNV0b+bLLoFa44EqcFmz0z5RUJm1jR0xgcsTTgEp2prHrsxNJjFiR5jN2iIb5MGkhPhzP3JUVZj7
3d4rTKI+TXM8xXS9I8NaFzpPUZBUi0b4kOTlYB91NA6G6LpzgVOamiov20TBJATPZKCAYpAbxjNy
yzS1gps9Kw97wdevBo7Od3UER2LEhmLDvAuffr7OPQdOzYWkdhwAWwbTTKFhK9U0BKHtovRE2DzW
qE3/5SQ/rUFJp4iHgR9gLPnwWsOTbp0r5qFlabyD7+WEzO2XxfupKg8bcgrIgszQJuIHODZklX5w
ZD1//vEwNGkSrYL9ciopW94GwpQumJM0TUs8/Mr1boy7K4zuRbRn27+bu4vbOgKsRAJrD6P9KFm5
wWx++Jffea9sZVBRMaLjzm4UBmHxsmmwieB9Qv5QOhvC2ZNZU7kZg4ShtSBQbVdFMc8etFe22i7O
qBT7RiZGSSUq8ryqGdScvWbVaHGjRzO1yLyEdrWh/LYL91ZUixEXg+1CLuhfvHSfR2FWlOPqTCur
370CVpFHF6Feh3w5Yz0sxUhE+0/d+OlQ4jTQmzJt8jAkxYNjo15Ddn0pwPUkW80g7J6kOTZ2ime4
UUxLkknnX+X26A6yWmCQT54djQRDtO39gvka28vk1v/pim2O/V8AJWZbn0ZRHBOYjqu6ff/HCW5x
5Q3jTWlbJdhW1Gjm207KnkH3BVJ4NGD1/T8oPf0jJ73yUZAOtilkAX8yzx9PyNzYsnX4qAGGrlWH
jTgIIxG8SC7+OaOTEx8N2PY4hDQ+ipYPC3kA0T/s63Mog+CFEuxYejEBC4cX6/JG2PexMLHG771c
PKpiXykOq38Nc5HJyUAOeXQac/ratDbdm4eZl08gUYB4QgvpgmF/TKsw05mUrx1ePwuavSmigmRN
lcX85MlwLks2vI1LzwNNE9n4BRHOuFRwclF6BvdtH68yFMKGCPNhc0I2AGgExBosSfumBmeNnyaq
N86W26Mo3ixfOxX5F9q17gq8YAjmJy2wH8iivhCicjGD1A5wqEafg2DzNS6IAKmHJDWWDsBA7tPb
d42n67iZcPfKt3VSoW8OezU3OdgAY6uyj46DaGm7yhIsKqLsqLpgj0kVF0wTWahmaY3L5e4kDp4M
9ggkRxXDk4ERJTooQpvEgdBQecTrHJRcqhEAuW3MV5DbNzKFN3LU7neWqmbgsj/F7bDpHrfE2S51
zPaRBLfJI/hTQ1/wKWWo3hmGmbxGeM4nSuQtTYNnlcic22ECzGsq2DzmO9qxQ52K/7dCwpi8BRkC
vpOHOgywyWOiB0xkCLL7CKy2oDCq/0iuJdo3NC8hzYob48tTZE6O7ly3313FTdm2+okhe6C9Uv55
KxZNHTGABFVJfaeDqvZJ1hnkjqM+1Q/hQFjb16t8AY0mxpfoo3bF2cYuyCAn2FG9ffEFRn+78ibF
xSIpiCMpadnm3J13FStUZTrweRVK0O7WilK+pK+AS/cEmwAS9ejeMYfClPFQa9FiNOQVp0tsKT1y
OlHyv90qbGRSFg7rnU8BUJNGb50VUJrlhRSkn3oyDmZzbDv9HURlgouF3mPHnWHb5UMOa7CXhhMV
wH++OIOMQGiwWYv1b43eXtaK5uQi9GiOrKBQfU0lVD6/nEpjnLRpxotAWfm4ODQGFr6lHeDLvK4w
8YgZpRapjfFmBoRkcg1BbPnOoRkY+YIdFvOTxBfDl5Q8iqnX1ws/q6v4seNmP+B9czPWaP621PvN
uJqcIYQ1LQ93H88N44gfZ3rr20hgg3pkNAih+CI5R27FPM62L6OviO2iswroGegCiX+1aoZaKnee
V4rVMkKqeGRq4Tn41CBcrGIrWAcOnz+u16hDPNxhuS1hePeraOtTyoB1Q1yu0exKVUnZT2crTHAd
5dh+fj2IAHrgc6c91F1hBxQUsWVJ6hH+JWBGiTyFSLq/JXD95Y9ifuAyt+VhVH5HENX2wgt+6vjM
k5s02KOYjaGD68hsllz1xcQ1eMGl7n4xtiJNqJzVVxIIgzYPZRJQqWoVBu5x9INB4O9OaSqovFZo
cBQtYB1uNszKVxOVJf71XoTdzSnK1bP2i39Wrd3e7oijj+i6xqypfsSYuPG4xO1iPSB5X0TC3Q/I
pANqXHoxN0QefNRjhf3gQNCuMnxwzmy3EMvp/qDXchyMMP1C9lYDUZe3UsF6CcpJxCzCguYZRodF
+XJYbcMIQYYBlGIKIhe8sbVdjzXJ0n3h3wTL/QUbcAygxwBYYG1YLkWrG7pPLEaE1pGxQqHBuYyZ
y8+uQUt4QjH8CUcK4j21/Rkg6FZHsoxSAUmChLzPGd68A7GaQZpeeCj8xSM+YeRxxsZr3PX5hi9m
0TnTRc1vm4rpNwItQiKKGQ42g99oQWphPTnIN6eQaVJa/lu0JwbruV5UDeDN5k7DlKTwCZDGNRib
e6TkRhhWF5dXO7cTiphg6wag3O1JbEO/Yle2NBli8fuHm9yxdqU44vvVhaMt/jUoXxQZ16aj9P4a
WrBjPDmeTqw59aesKr2QZtXI9QxoBAu+/aSyfk4x8mZPVwIuDIN/0MyJvXIZxYHbTGjl6kZ3L31x
E4E4Jkh+F2cexjGYu/NOqUQIOYfEaZkR7FAVTxYc4JI4pJcG0Ifgclk5PwoLlBhCF7QH7+8r7aPk
a7TXc5zu5nG9cqIXrUID/m6a7R8uBj2SUWZpQNau6k+vGJVWnmAnZ3202ADLVOypWStRrv0lcjua
cgxY/Hc+23sqvO4GenKW++ZayklP+gJNEPKKCxjTUxiWbX4OvFdk90G+KxOunIS+ASZv4/zQ0EG4
9fNaCESAoTVW0v1h2G9Aitbj749HfZ1J88KDtkl7FVfrOq9CGlaipyrNpIII1IPcsM4/MpfwxxkZ
K9zSOekKxjd+vNNyAS6OSICPrCyeVh5PITzzODgn81OcyZc8FlCIK35DQ9nBCCuOYXw74ZMrOPMK
6XTInOmhQIwUr0WDO0VlVJGhNKyWPsWWX/np/WDQ2NbGeoJJ15Or4Mr9qnTlogg0K2piM0wNJrcS
HGXgt4Vuvecpi4cOhXU+vJpgTI+0XnOAGRMijr2yHHLPF0h+K3ORy9mVWb+pESfv6dJMiLEzcT1+
H3vjqNUvTuao2L+RAOrN7ZbrfmJ+NbTOR5ZNe3P9cms2rJK9RTSY5Kcch+tKLcWm1oEOZk3CBqtV
lF1tEzLRLkk+xmsh79vC9RKV5PZXGgNW3GGvf5ymEjTuyo2xi+af8EJds1zv5x3gsSaws514j8nT
Djn1sbcvUf8r0tiCZyCBILlzfMWx4b07T5ybxnRH/qharHSa/gVLbSMwbMWhjo8XBEoHRoQ5lqn+
a4HwP2QNGqYlxD7qUex3sH/mPKKZUHVVOsa10uQ7HvFVlXWVokfZRCBzEMgtDuxCHaMXJjRCwisA
uMn5n2dF96zK311BMi9XuZIjG8o0eV6f6mqt/azyuLFG193oCj1vWOuzDb1oZ6KDAHB4QTupBfGK
o89DuTT0jvjwDFouhf+XzQqcPwC647FuoJLRlpjNi3bOk9vckg+IN69pyymWwFBecz/SFSu6gBWe
8C2uiwosb7aWw94Iwe8Q4X8NRaVPUl6yge7wA7SJ9S0bqTfsxjwzGVVJ7tcsHJykk/JshuZZPnHo
aeaAnU5+P96dQZ5Joclpgyq5zMuNZesjr9wo1xG9sWP1Y1JG+B3KPkmRiPOtmu1aJIaP5ivkNSsZ
YoGAHPV2ZbnqWOp8lyeaclvv4pyoz79MmH3UhcxKB96897FIG+kdqcUIkpw/zrP4j5zYuiUXsNLS
b3K5UIj4jS9RU6Za1ShPefi30BhlBP2g+uMBl6phcIQ2B+/qYppthe8SWaAIJGg5z5qAOXBchthH
XkXUCv6IE7SSnViHTFkQKceCQkBGeOTXoWLHh1xKLGVTB+WJvsWfBf2VUFcY2XM0ZMW2BV5lI5dR
X7WU9gZbB/rJShjEprBUolhM/H3wDAUcRsXuNzN+Np5UxvJAopePDwr3I+sMwQH9/o9L2hQFQ024
iItqwMdrp/PUnsuiHEUFsv0VPsdk0xR6hgeMlg57KzDPmkTIWgrbmTu5LbuTMjAy0qKtE08QaMaM
ZUfpLX37doVG0MZ/RnV9pO4B4u/WgpMjd0m7ZBrPP1YNdCn1fAAGm3KmrasypxWjnx/1Wuzaudv7
+1TwaDc3tew5SYR86LQxUt1QYhAhV7LzzNOPQ0FornAXg1ZxDOclZD6Ys5JzkkjjxXR7eqRTRvEP
4dQbKZk9jwIlRCY8QrtcR9crF1RzIQPuHlbuoQSdh7qV1iQs/W4Burrdn668IYHo5NNMjyg+rB5O
Sve+yT/BXwy7mxSMX9qeZXirA22UF7LuUwbjOkoay5ejxI1K03jzMn+BnH532/PLDbKW8+YJq6ly
YlXBdWHQNizts7uaX4AJQCYJHb1BrapxCC3SZaQrEfmneQmu745kuACt1O2NbHpeAAgfXcHJC+HN
6OgVy+KFtBBORMUoURCIppJV5xpAFm9JRjPx6mjuQThtFijgMUzELCxJlSPhvS/ZK6rIi3WYGZcU
sIgBWzHHlQngkw3QihUOzIMdlMW0byL9jtPU7NV1/qUt6cvz4dkxnsMMuwMhdUfI6/ZJ76xYZsHN
xLgP7uYGWm0TBVq66nprLprf0Y5r3C3Iar06Qf3pHdfgI6ihP7bnQp2a/PJiYtlFggCUoq6y7R5h
wBB9KiwsGcG0z7dWVoLU7UMH34YwyMIygLUIbDBeVKWg1Lq2iku7TA9MyI+uozQFOeqBqrQfi3LX
2vlTiLD8JuTbdSNWXAYSGYhIFtzP1Bal+jKFSvnrVCXpiSwD57EZNe1l+WDNiINsPS2oU3M40ds5
lNn3huL51l00Z4S83LohTo3HkgKDzkZvDubrQkoCgMn38WA3PrOB4nwMqo+2bfM8SYViTl5I88Pd
J2ZmLs16/A2ETMtc70QyJa+Ez59EBqEdQ8G669KC+mhVdMvxnUju6KxkgtlsgIquKwO76kjge5o9
eaKFgWO9DNprfj7nr+XaZR0t+mVJlBeL1eWgcpGf/7938c1MSfjpRCAwecwe7gUc26WQS8zW6RuD
cMeK0RPUmhYQPRleo/VdAe38sozVu4miW9FBT+MTGJLkeGF4CDoizzxGhutY/VG8vTjVwr6pa6Jn
8bXnGWTJO3WnkkGOBZR6OH1FkKivYsYMwhGu37gI8JLJ3/yBtY8J/NDD02Bf6glLY1XOGB8pAvMH
ukY+ObUFg8snMKHGMLx8n0fTMRHZg+Cusgw6Sq2qFMthDaKuVhzPSClDJDv7VeTqthrRJnKB6tkW
9FBbPJrDSMvyoEo6F2k2/h2fyW/GgGeM2T61/3ugEawLYB48OVB3kQzS2Th7h8+TI49CtyzkPgpW
+xMRf3dqzMfibUXHFnqwzfYA7dnirM6xIFEnyMPa6pfdMvWs2DwY+XazrRhnU2rWpTuVpAWvLv5+
9GpRBhgqCyZdHr3eu8KqkMeQG7YK+VezP765ELXr29RhiZdnsk31UtrC40kE08LW0b2G57Psa3Lk
rKfK8mTr9x6orM2mvJdqyxyREqEK97Sq29uOjqH6bTPf4qxn3eZALrJlehzlPzh8aAqd2OeRrsBj
smuWbVGSbxPQ+XOsQczs5QDc66MybBCVLlZewYcXbX6zc3CVN+arkHM9ZOXq31bRW49is3zLsq7i
boBlILWH5UFpPvSAY3x3T/lZxf+4o7cIjwzUMzBn0AX5Zq9VyWhPLmNVXIpfqu5eEF3F+dGkisMM
LxuoG/Adhkk7L/D8NJkpSXvAyQSTk6R7DClgWlPWSr8Z+2ICxo8fOPSvL3giRqm7UEYF65GsjpRV
uPK5SEO1Y3aemxYlHRnP0laaHZEo9rbjoRlmfq2xk0t8O6sIfYdVuL179C+MeL2HvJ7f7XinEQQY
UHg+5JRY/hWzE4ql1Y9cf7maJCSH12RdpQf76mBDJ+mvDfbEbUIvCszpj/YLg4+Uys1WaJngzzJ5
3gVdY616Zek3WpIayfJoZdFrJEN8+N59JYvxq2/7iKGBDF9A5uns4XXdi8Aa1cvm6+QPQ5LqgDtR
mNXuuzgqtrg9wnXWlmlqKmt6cT0ZlaqYk9N/iciIJQFInVLobSF/sbHoUV2zgnSrYI0Q2r/JATcO
miZsqiuv++ZfWFy7zMV5eBnMxALrsNU5XHMkQ9SGE+XFcdYrGcmkpsJZ0719jZp1dMY1A9+4T81m
324V3CLDUdhJYslc/a9Icc29rWqgDNe9Sis6TxJjZzNScSmYHOM4s/NZ/8pYrQ+vOPGRSaUpSiy8
N6mTcsE2JHn+78FRNWSu3OSPXyPGPYcIoIjTk2Q+/pq/Z1DTLG4Osop2QunbFhs2/qfgztXGNOH+
L7HKXk0+WVg8vdQtfkTZN7zNySkOMEzxugCpyIRofbUDRIC1LrZ42GhBICxC/bMhKRw7Pgf/ga3v
D7ESNnbMcirfK0eRZeJDxltQKS5N75IrrBfNtLZSq4fUrbtAuMvJE94bVfiA9MAy/wTz0Hb/DhE+
vEjP/4hvvOOEO9OZQzMHGr+8cB4ZQ++vNhDg1fCczVboTgqT2LcV8bzDK3sig+ZBYWGK469F/cCK
wJqdmOUY+cH60XyWJ+v8VMYPd0Rmz+MY6dTw4Qhy+Gn5IN2d02mG8pULMfgILiF/ZukDR4LJDHdf
EfvxKRGDgUcrQaTKoqWbAegSoL0BXKJ/z0ZoDspeq6OEcbA1+WRXdGT5RJayHieXzEMGh76yBN/H
lioIocVvsv7CxhEcYjJqyAoayahpYuvHh8apG7H01908f888O0oGHq1mz2kpf65pw9H8Zm6dNAmO
jjpVnDFOrU//IEdnr02BL/uhWDsohi5BFKTf4DX7aVVsW0NPe1+WZG13/bWD4f/SMUhjat6teHGT
AdKbfWUOI2RtBKhPRfqKxky7WE2mpfG5nLX04FcmKyUlMI6s02SKnl+/K4/BZVDhcrzTj1RqiyGM
mPwqr+91dxqOuKPuv3Uu3AJJO0RziLQT40mpZjntTLHe1bc3bqXoinbLYwTs5GNzl32vSNocOT59
AtXGfym7iloyIQ5tXl6w47bKTB8M0McxArTb4HefPc9u9PViXL2owYQmwNnWdD2IgL8CVaxLRkKd
r9v5uI0TRhPEO+WUTA4Ek3lffl6/mHCZGXSHxa7k0uIN/tj0Pq1WA8IVVI5qv9bwXJVm1cY+l1ED
rYOSx4ofBQAtMlIdLnk7YfxEql40aGSv5lA6Ew91E5CiRHA/h8oCBk4YJzT4iyricNNn1KCuqO7/
71Swwr49bU2YF/TzyIt5sq69vOGNCS6chWSUXwnZeeL1dP2b2UUl4jqgkjEXqrbn16aSYoCrYTwo
rE9mC40Qb7PCdhRm8N+VKOcINzALkIDLpEDv9yRw2rF+a9YSZ22zKOND8G5yjNMLteb5JtW3/3IZ
0X/41ISv9dn3aAUfxE6Cf2Sz2zjfhNAj3Xt9JbiqUbeG+5EQhp4TKlavFTO7lVL/ObQhiciX3fBm
PQb5AXDuLD9KncAKOgxS6uknMdurzGwAqlp3nhQ4WXq2r1+b0Nnl62kQn2HWWK4dqsNs4Ot5/+3v
8hViALP0nSdQsoJ9dJDeF7TrDGmLoiEoA5Dj5SaPCmrLp0BG7SQLVyWsJqwgiTFzgjkiwudEglBQ
NHKiB+UcXDXRaCUOIicEEzcFPtkVAzvlWRO21S6MC5A8611VxwdHMctKqetoijBNPXZDrvpeVCza
r7lAbNYYgsBIy6NA+/Bcy6e9xC+zeLpNOqeaffxfUB0bgLylFpWUykGB+Sx8Fjo2yoNLJlfoJe3O
LzTv0Lhj16j1udN+QQijFWuGl1abWrbEm7F2par3C5Su+k8VGXOJ2u5c6qksxqXVNOL4px4ZcjaP
NCOwKwV16HE+Vm1n/9DiBuMgywPP+Iw1hqohLguMMRxT2GWE7OzXGgvUXVtEoJ52oHWXLcwKsIvN
VV22MUys03wtJ/NpkJur2lU2rl9B/sRei9neSvTbUEOSTCepuYTEb749piu4a+Mpo3wh5eU9L0zn
4JUhsTAGAr0DY2zLy7nsxlE4fLb6ehmEgjYbqJ+KYdEVEtEKaiY7rn6M0C2ObR+Ig+YMT3bvN8dG
7EtEbb1XzhTyDELSC2TmF0urBotmM6m+5LObQKw3GGto9oRW9Fbo/Xy+tH00Xa2qZlB7sKSFcFVV
u5EIhAmvrRFa+E1XdK2BXFA66G19fGjab0SPl3hl5cag252mhAtmGp0fWBXDVo+JPHus0Kh82Ykx
2v5eTvHUXZaol3vCHeGsdNUtqDZf4P0hrv650wmA2F0XwLX7zCZ2Zfu8fsf6h34Q+4uoqXMw4Ki3
KcMPDjUbkLRd25WBIgPsh3zPZeSF3lGIUQnkVi9l6VRmJQrKjh6Py/f+7rjsAlK9nVbK3HTf4OPi
n1eBE9Cs/Cpf0E+PnPoPng02hLE0P/LJVv2nwHHCSRKC6zquYG+mI07IJ4XuHSRMnf85UJrOWgsl
Q1uYZLuSBLVKStcNbFCraqST7AD257itUY0OsW/34HpTI7DKEXYlHijAQRVSGSgLs5lSQdwgTHmG
/raNBM3TNUT+T/OYjvfEsq8iMXVXqP0tt8MYPZy/XI6KuT3nGYZZH+G96hQQBqa3hzitTY5KRC51
XaW47oDImc/ULcvJexH45lrB35IYopkcWBBVlLjB/gsgdVguWK6rq/iCeTUyp1ncb1sd07m1zd3G
tTlGVhXF44wOjAI0RSyErpsq2q9bPTWOdAZp6kUMC2JahBWhyveQ34QUCAMnmL2T8NfvJSxdD3Ux
6g2Qkl11kSy3G5IPpRggcvOd4JMAsmpbLqIWjpoZcovelmNHbjMN2V3aMv+vBrAZeemSQweavdis
woIl88TMYT+/1fdQhEW6SeZmtxGy4BhvrDWXAqYx0JCe9CFq2H4R+q3/ZEHceNnxi+VkQ2n3i0tQ
pg8HcIskUy6KZrIAUif60YlsUkeVUXS8ivlSkzxwkfW4RvKzajtJs710CwYC0mM4S42JYC7RsW+e
IU/9JWDHpBGxqiAA5q7ggc/DMNU8gn+52+s05NNpZBATlGYasGMjvg0y79orJaEYCWEA0C1feX7G
HA75uBANhcV3Xm9XAUz4oPwfU31DR7C/rtZQdnFxz52G3oPH6cIPyFUrRdsbYbkeZcIO0Qoj7JyK
thphA+KpFpiu/AJQul8rXCRBR6ES0XtuOKnp38hBovRqua1cqNsdvoL80o99XFFkTmb4F2vkDfg2
BlcDGyAXlxcn2o0ZCCLIRR8Q/c5Y+4yMeC7ejD2vGil5QYwjrX/wfI82NVkS7cb8GATKWIbpuDkt
QhT632goTPF9SaOo4ef17Ufm9NSt7DzT2Vdp3h4RP2d4Tg4bCeBEk75vS7cE6CIS+EhgK9ppdwqz
JtqMoxu4H5p3n/Yhwm6oc+fw9i5fQ6/qYfWGD8a/eoB12JvTIchb49gpQgOCFEYPvz2fTFPSwkMK
rdtAXnjotFh5eklItNqPHZqRfx4zvlIG5SEhcU7kooOssf9257sFXvGDt5t8j0fjckDv7nm9AsHM
OkNZd2MWiOfA0wTI2HCLOoQGP7LbEpJne+TduZJwI8tROZ/12UIpncZQB8LaiyuqMo/4QiDBAv3k
bqvDYfuMk7d2keff9nEuSpp82wvwZRPT1FCXS0rW322Loy+bWzSFci/b2AXPacdeKl89LxYaZdMN
j38S9vKDThEy3qaa0xT1k6qEMuJuDHODJZOi0upGcKM2pvF/hL9hHdpwta//cW+EcPuKSL34lIJ7
pua3sdyspMvqaHn9/XsvAf/N5jonmRicciekyYKGtnMQBG/TR49Y1PR8vXqytAG8zbbCmgYNBMe0
oOHmnxlBf+H30cziVdAVwopd44yBQeQf/q0oN2ALAHB8UXclraT9/qZom10VN9moE9ASNM40ENpv
b8UpdXfAR9LHAbaXiZKCwJjjXoeSvU4Q6e72taoH6XS3pXQflx05rvEclS6+ZAx3ZJzPUd7dpnId
jmqHOsqgS15mgywtEJ1aMCh8ZZTCKpALMSY4VsB2BLuO/MuyN4GvKttnAmfwjXvk4I7X2n4Y9wtN
qEsrZ8d3pTm71f2n6CcMZr6AU8tzX3uKYIpg/JAV+FT74dbjozCQ78xr6vIpjozRRu6LdfWWBwpO
5Yb6mLVB/zhCNdZleur3yO0BISqNQqk6uKyUHsSLCYhBKvSZK/U1xSUO2ZQzFstpqrlm6cNYvyZP
LHrAVlQAtVgdyj1NCGV0NISy9iFiTz7mJgccMesMjjfaqKekO3dBCI70pdqQjXY6Nqh1pIKTYTQa
W1tnV6WGHqX37pOImalgIXkC4A0mMfcJvr0Q7zUFO1WCykweR3Kc0EbvvCFgJkWstYLMa75Hx22L
7YrY1TnaNoZyi5UHPm1HbXazsnI7FI6/bJvYTkx8FTfQ4J2NQfaE2tffYrOn70xliGwE5QxkDrHo
kRuP852jKPo3YZMuicIpkJYBR6bd7MGKQ3Vveh4lr1lygNs97uj2Gh6+ZUGBVNcqziNKnWsysFJL
0/fMDN4nqcDoLWNFhqmUcKP/47jo1OxubUy0e5AgyRnFqzIe0soxRK2yLBzcghe60mqZjOKgWPtd
Iez5KxslwXUjzbqt6csVINspWKjxZD2em8yVGdDiHMtLxEd+GpwnPcmeia4ThULtaG8ET9PSIHIo
CXX/injEuY6PXPEdMykYeIG2nK+y6mr2OC7AfDDWz46TMDZ8I3ijYRg6CqBdoy02Z/vISWV4Netc
Bdr9AgPOhKiGj/FAvTqrgff6KdPYVMH/w8X7H83HuBauxG2Q/9m7ApGp2r1+uM/7j6QH7b14RIkX
k0DKGksSUWIpqbvsmCX67fgCjJvVw+LfTxjSlQarg6sJSd1k/PNvN+MVxQnbiXEQFmVGyGHPeKU0
j0ug4/RyOhmnS4JYzo07wDIXzDHH9DW4qjHxY/UrsWe9+yxPuJ4xGjWt2g3PI37D/ChJvh6lRAGK
FRF09t15zKJFD3lW40hJ4+5FIJYIdZAZTE2/JTzdGsVdT7GIIau91toMTfpPnC27U5GhTfL4Hx3E
/cqV3GEu0ZyYSqlHYVHlQYJcbIo1nDjTVeSwLHghVDOYjuxSN825xAKt3RQU7EvJ9TqiJ5Td5Hen
FNOLGVt+NEzy68vaPhsr+q+fh8lCAyWgneOykYmt8e0c62YpAyI6UZpyo9jMH2Jka5SUa+VSK0lP
PR5QK3n5jxaaJUsbM6Uh9SDCricruRrlHidDODJyGtR/U0CjFCMOyKozveYIHqWOTS3U14tHVZtY
TYFkJ/6XO8aq4KNgBdhDzNBmGIe1tMgwOGYgiLW5w+qOGSKu0HYFd7Wfzh2eCluL5Kgl7qXM6QiG
UCKtM6sIoBA/3lLiCCrHnKyqEu0raMq2H2telVjLcHY9RFhnwoPfNT48FXaZ6CH2wmFSU7vG4B7z
XvHnWb0GUT8O2yn+CkEdfUQD/OUzg6a+wu+ue0KeYsPrWSJMUkePgNDqRe5TNUu1fIF++pzDoGIk
zueeuJglMlRZFxdog8aLrFow9Rv3E8clixzBMnATrxj9Wf9cTk4I9UpSqVq2unITDh8/3nZHMK9D
eoNXYIR40v/EfjXywCBMvrPsT7Hp/y1M/qkk8NYoaPOHwB6w51KIMeEUgmMSUDeLAD9SveYBW8XQ
5G8O+OgJ4oEtwo9KX9xN6kC5eDuGYzamTPHgLLV5uBUiKn/eN1E/y7RraiZ3rKzxce/G5uxHkdg1
dAxJpQllkQil0Wa3Ek+rYdQt2Y0gCzYeiYP/QMryueOXumkDyW85BXUz+UNSZIE2BDnH6ktwmYIZ
zEkzJuYvSxKnJqSssjggZkuvUdPgPIRhyRBhtjPx4uWoo284lYroua0WCam8e5GUtEXBlsc7tkCA
NQOu8UNcM1X3iHh+UK0vujOknlJd8T3AUgcEFEpWqs0X2wJxrV1LJgicohjVTFR0JHhqDhy0uw5/
vIyc0cKkMboWKqUwxUqVaEFh185biW3Zhxj5UhEzErJtRnYlCD7GS18lkBw0FVi8hi9msHWUcq0b
WTaV3/ONQrYoNoeKTqxvQTENjm/xrpQD+BdL9XDNz9g6LNsu0lB1w4Y4eplwyvBHF1bRRkNuOoOn
/hBBYUN3TRYTW8nvBzuszBnp7jOCgkMMY2yoevzddx/BEaYx6sfcp8QxrBVxclf59AMyNCSnswpS
2ApFMAjxW4NA1TQNGjQ4QaaZRLhNQ1ZUJdWWgjlNS8uPUKkROmcCqOCLfGGnc3OmKRJZgni8MVKR
O76GZELttz8BaS+SE+mKWqWcY2YCc+8MJXClGvU0IcAxWyV6eBEhqEy/YVh5EXKMGk/knqAR64TN
o/UfkC3USXonUU3chuv5U2z939vFH7eRAq3vOFlZLhMZbtTtkVEkWIpxVuMbLRU3zpKOUnbp1UQZ
GQipDuhLIrbkgya2DevaUAkEQRp/seEFzO57odaafqUtDICFAC90pap/wWI0+s3wYdo1PFDXr1dr
0RPFIGSVYuQQb0uS+x62WLcuWJ+OKV4lwg6Qmv+XthiZsrregjR4OMi/U1N7FhhO0PEOIQIZRND/
twLG88nstctAJkTtwashAmbMggzLFQfi9pxv0TMjg3iKFxqGxEzhuV1d4hS64/KWOlbJ9FQy0nFz
QQRSWY8YNmw0K/rTBmeaVGqSt3WsGNVhtt9Ert4pZC9xFfdmT/6BZRhbxM2Dz3TiWkk2+p5Jhbvd
lvrE3afk2F8qoXNgouqY+2n8ioPwY0cgw4oJBxe709ptzPwZWQ5NdSJYXgJ6N7PLgCTfAqqr+XmR
GhdjPCBbQ7ynoTzm9b8u16pOmTjLUt0gXBPeWx4H2b2LeImNBHlYDUVZ7w8+vJYc65ddq87DONSN
KBX+9j0srrU7ETsLISMAD2RTmqDaiLVRUnXKbCoy/0d6mtC3mCE5837paL+KUxbs7wYitVdfrfN5
WA2aixycuKkmZZWTo/vdD+aUiWTgHn27izQoQWimtzRMyIB7DVAc2U8I6Gz0SP/GeiI3VrawYeDf
TdgK8iRqB7fmLPcn8oE+Mhdv1r7sPKKzbJf4feAoJ9aG7LY492b+2Yrm7eSE1iIImp+rr5tiBl8B
y+dAqBDcYvg/8w/478KQD1oMHFg4CbmN08S0SBszhgwPwVJhA8BvnNUrjTOZTacf/YnjGla7NrXv
6ckLAKbyDCJhgZ6ddN+FTOVsy/4fdv3ZYUflt8ocz21H5rsv5AXoE6K52r+x5iJ0AKFkaTKlqr8M
TH/4vNzxlFciBm4wmHEhTZHbw+uBj1d+lYZigqguATd16jxQ6BqvJj85s0s8Nr8k0f698l0xsRP9
TnxHqwLRc7cgD7yOYWupe7+vkJcnFpS9UxKZ4Q2JvPWmq0EtOmgn5G+0IJd6dRb5AzlKqDOnU2Pk
LUwX4eOZMkpTZqHlNz7NgagrEbZEuyT6yBpCWcCr6r7ECwStA9mjvNFqDfGVU/chm6q9u3ku4CMr
NCWZmMABDE/ggviodHudBobx69zMzs9GnRd3aohAKWfCFqOKw5IFCAynnBQAgLPTZ7xAtWCPPLaT
+PycwFV93GWq5D/MEt0S6i6dPAu4wfof30ho0TvEIaSOGvEjV4PZ+Ljn0ApvzN4tSXHRcpo3KMMd
8NhKEMiM1PEWAXqI1Vfrci1RDpgQat+A0EW2WHC6rgdeuCQ7HbY1pNYUOT5BdvRfmBf4hVbJgWIv
Fq0+wKWRgbXfddQkfDGqhHuv/33YgcrQ3ISWn0dedaIbhKH6pjajQ5Ki463aRq1uur8M9u83fO/R
6AYS7+kMa2sWDalvCFFRlGFwBp7QHoS3qdRZLg1s5RKQ889i9j++X1AHmIYAsHm9HMN3YqHNdo13
iSarkKG23QnaIJjSDaDLaX2CFWgb/b3Wcv12MKJFGkmk48oEYh9Enywi6/WMCA7SkCHbfEDd+Olt
+8KqrzMOKAi2R2xWu4+/eS3C5mJrXYMcLJ+WxssOsysa/UeTX00asw6Qd57q679muycwMh9/ngaa
snVrLWbo9C9xvAzH+EQCJiWjVMNFqefF8GOjeE8h4m4qIA9bg3l3MmrZYD3z+dPwbf4/C4OMGFov
gMfM3sg5CXXTua7JPUG5OlgAH1aS9xPJsAK4x30dVxJi1ot/pbikiAj8/CnW05sw5haYCHDQjN/e
eckWSkZmTOSCgP6BsxIw8eXFrMtVfHnyA5ES7SLwiw3Pl0egbueyO235XaIRYoFqZ10La6Aw9m6/
goIs9OHn5UwaK1/PK++h0rpX8p3qPBqwMdZ9L2aSIHYvyLS6RiG6zREekJkbGOmbqKkgyN8TI8ML
XKWQxkY0OV+GAzWeWaXfPYebhIwzx7vw733MPzh8XfuheDIMP4iQbJA/HyiZLGI2jKKLOi35XyPX
m3/btQTp/pyY5v89v6tkS7oKr24h8aUNp1qsqp2+vpHqhojn7ysappNNRkURsZ2ZNcFjHTdGT+mL
QcFr8TAQ36vOQsM7JRQmkbQcqX5oTVIrxdBbZ6dIyv0ndc2SGSVo9FQFN8g3uAyQTevd5g+U434V
xEXscvNmCOzC2Yqygq+jxAPxb13rLVLNhnv05lBtr4uOY3ZV6G+9YkrOCPp7mrPO0/zONP+uGdw/
pD0laHyGv7+OpSVQ67rScVJ2vNmniT5jV40nPWiMDglRg87jEpm5xxcR3sQiKjIbH+3o2cvHP9V7
MtP3UV0K40oHgvayz7xCv+RK6yayXGfkDqa9dBlSt2AGlpGH4r1BE3+P8OVRqiJX10ngdtCC/YFG
opQ1GGpJgmSJwcwQrb6LMYltlH8Y2/lDQvSllBr0L/Mbceb0zBeDY7Ggqi5Ikw5ej1NtmLHUll+I
v0TgPsljc+rQpwQnZP1LqBfL6DLN5Lj86L0fUtL37GRwfFjuBxuX41lOxagQ9mHDtBFDSgxUP+ts
QoT3bE9S3/U6KR8ETanqZEE5nQlopiQ7I36H2ixLrpxBorK5qC3irIunEpB2YX+bv94m9JvIQnWg
3kg/5Gn/lf8Eb+t6nwbNtEaFjiwy5G/Ao918grKNQQmbdk/I3AGAwQ92jfhSje8g3txq8dew0N3c
Z5oAdVkFegYjN4YJ6AXHxNJnM1+FyxvAC84rT6TFid1ODTAx+6rlkr65f8JLSpW6aPAQKveA1pie
nTyfnjku7cYUhX+2tzbisptxR4SJyCbGRSBMjaob51FC60ZcDeu3XFqMfo0X1DrgqRVANCKjdpD7
ZiZTLl2FKuFhTgkQoEH3daIH2m0eeW/hmKHc0GmdmkOUJ/LM23UuSszte+vAzaWNjjIsPlqFatpy
nf6qqIIOVBlt+pHlUfc3JYrEJiEebLes1ch+QlKZc+Wlz/O8SvlQgiHVqPLLvmd8sGQns8xt0A54
yNBKYVkJMQezN2w3nWuznnuIFckWjM5u9vbfJ9+FoJ7UEneYWxAdq1Mhpra/b/ou1Af47loZ6Ocg
kDnDwfvhnp30ihCA9cQzvMYFTFOnx/qVtYja83pWsdbSrXdNLdA+9hjw06v0lnvy0nVkxsAt0SA0
FhSDaEUHckxVvTevAkr9gjYdtPJ8bESeyQB6JmPml6K39XW4AtSViVGgNM+oQkyfdRUwXQDRCPU6
fGN54+trjJzCdy8VrhrPh+vPA+ywPS836G1rlpXRH3SRIUrCmRgafETHeNYh0Uig3OFqG9LbF9Q7
AlupUzI74HfY5zuKDXGhn7wP9YefHe3ZkljgGfifRRD46r5ngfco3XBYFxG72d1GD2gcge1/WLJr
G6Dfw8BpCF0QNmgQFhE/h90DcTYjk3XohqqIYriEPoc+pNIhFUEKFWxnyqcglk+uiRsbmAtPzQNk
YkZgHHpf9pVn/5gwgRHpoTpwhWD4mYll4EaYW0AMJs2WswKVDtRqy/fjEpP5It+N4ulXHJk7hRhJ
K8dFWj2NB2YM7BCvaFcQKCvTOol/4KYLmioBpyVLGGz2AAyeMnr5erS4oxIcrfJUKiksmeO1ftSk
qbq5jLK2QR+yozUh1ogAKLOLoUircrXs/OdlsmwNe7SOXGIo47Qr0E400c8WI9EgrT7u9LbaD+K8
C6Eg3iJL/1uRtK9BMElU/j9A0KMNHVcihmutX5zgzVBB6lrXcFMxcKSEg4uonSMZNyhbxiE3TCi7
vBGW8FenWReGTFDFgektP0e/zqcgxe2QPd1HG9OwLGuFoScXD7+ZwzL2Cf0h+tjRuph5fnePwN5n
4T3lj0rIpX7+ct+2u95uoWtzomLw8x05miGz1WNzoSpHN3wxx4RsQR1U33fYKVz8BN0gauBqcKvd
Oi3/jUovnCTNdxuI1un/fTP/lGhQ4m9NawD4A9ebrEZ6+NeFuiewv6mWRTTY83/S8wdIqoy/egup
pvM2Jk0A2pdP1qpFQm2/9eW3olHpl5d8uTVUzF3LqylCcIm0pPivkPk8RMPpxx3FBF0H/6UU0fxa
qk3XeIYZ9PbSvH1f8ccSXlgb8dfVOFa3ioczoRkPiI3jFTaRKS8j0DZ3lh5l7YnlrJ9fzVFV7ZMZ
0cKjynBV9AjyEN9hBTwaicUJxULk3tjmeRwcyNesE5gpY0pVXgars4e9eMl3adoOLBQbxTtFKx64
TWeCGdk/j4ZEGdu0eyM7cxLZNrQ34imgApONd1oFFJ3nhHOlgcZeme86dOszsVaon25vmQHwdxkC
i1DpkjPnY+tODIzjQ2MrECgtX/HsRLqpk1USVgJ6FqVbXh6Bio29GMNMXyOhOyQnIy3sdcBCcFsd
dFAo/CQp4lnMw8bG4reQX9XZTIqevrfNfTrSjRvjKBZUpFXZ9814rr7veyFm/mbb3gGnHHXs3cyf
R9vUrONQli41hdQurISKgOkciLCNav4f4sAyMCR+EpZP8UmRNdf7PSkoJi/+TLSKtwGpps6Clvj2
U36zRdQZmiabLL8gIZoenJKeuYPo7UR/1OggQS8O+W3IKh+SMGjTCE2iR4+vlAulUhIqGt22cJ7i
RM9BHwAZd9/zQ8ItsUQ0PREdww0KGs6i56DkSajX+8MX7sW5p/QYzYd93iMCr7pt3TCz5lsDap4b
6uVB6HO4L0R5xktSvk9euzCKaMrwTDFpFbc/wueCjXwV9RAhyaF8xC5MrQHyUJBxlw6ZLRtaP7Gx
CPMC5bdP91cSbajMDfnaWNw+g5KObtsWyKg7oRbfvrHa7OyMaIfmUzXjVU9JtkzxlZRDa2xg25Pk
lTNpEnhCa8pMRiiUZ/ro3dnZH1aVfFyK8M5F1/SlDJYDUPhWVXb+AwYyGvDVD9w588TNJGiTFpAe
4TM9WkWh8yF+AY+C9RL+1jEgOdsQII+Lj5BXY7oQAVqkkj1yoataX76bmYIt9Eb53aeiH5dXBy3z
zM7+EuWukxLWIrPewKaIVhjfHWR1w55JU2ecRl8jQp46NRSWLPl4wKouhle2c2+pdhLOB75Ix5Na
S2IJ8YxnxECW0Gi67maslzDyVQOIOFJ3Ko1Be4QtYR0ibNtuVcLYS43fPCOs4IkacWrunM8IvY5t
8ONiJBVj0maB2k0BfWWomf7td8pYejp8+OiZBePP138h6FWEbUX+8quWynAN/psBdhqQS6+kgcWg
BPMZ6U05WYno6vMGHxpb4h287Js/JgZKfyhqyS+DEP0vYn1i4PfEnE04tTvTdxtliUd7n5wWnclv
5r1I9C4vOV96HKFmVtphTfI27T8Onz6C30KjRWS+bauP3K/qmoeJIOX9/41dgpb/7I/xUN0qTscU
b9mQepm4OeM0uO8Ng+/95gleflA+6K4AdIaZltPpNnhcMtze8yK9whJz/ZtY1fwA28qycJoAW0gq
2GVWvz+CxaTxR8hHFDRwmiBE+IN/5aD4k48V5XENRFa1EJSd7NXPJeeT4+0iYGx5jLWW3A0Gclop
TlgLz19x4JxhkAwztFjrTtVsYKduLRb1swD5ZZVJpDheKqzq4/8iNEEOZG5BsiB1yoxMWB9uCrVW
mVsq3nx+sSlGLCJFAIXlo81G9ocW3UojqiZndPPQVLgX6AWReuKgJsYqQTXq8TeT7iOGNNZy0pB+
23NauYFuzmklsV9BsffvoInLx0QCTqXCeBRRy8xqZSLMfhO8MeJJ7wF4kAbOzXBf9p4yyny6EbtX
KitBmeTatr/XvSbWm1IzybNsnBHa7LhnnzSksS6UChxI+gNHq0rvR9veC6qcO2NipBJra9KYwhzV
jQUoU5kZZzWGxJhCJdwELZTWnLc05t4zkSfGRJqlT98NOtf9hlWIKFOuoI3/ZBbvpcxVwTYxrVC0
DY8nwhBKfNgIfhMMKGVUBKmkqwVesK7IXeVtxXQQDiasAwwpzyXOzmpIVNxXFatB55a+qWYZS31C
uQgi8XxBHuWQBrIx10eI0ayP0oRQI/rvZRwbM43QZE/xNVrF3n3uah5eaE9okcE4x8Y/cmDhQ3rQ
kQi7Q63JFG6+2Y/r+9QppQT0g63QyeUtdk6rLOqRRpbkiObe8YrtZYkud6VAV6UnC/QMwZbwT8vY
KD+OwMfrWb/cy5T9gR109XRlOHvxnT9MRrG9sWBmfhJ5gMC3gOvBvVTK2cWwV03ydEJR6irsFV+2
kvxEJgXBJCpwuheJogK3B81OCI/P0Ivi9bwAie0xwd3EQN8Oh64yznXp8Pq+lVav2uO57Do4tSdm
7MaJso67ha/R8E39uNf/xtfO8Vn/evqTs5bLmeZ8t2iRGf0X0V3SUffL8DXNFkG4CM0TsU+oobJK
bCWJIo+iORiCBc/wTlGxUdWzTl9bZ0+xdeEY7GNgoA4pOJD0dN8mXG/tFUKufyVtXmvdckZUuVR0
bZQpO7XiSbmTMrEEjZtNBHrE96i5y462u0TplRYATsN3Z3sYbA2b8w8M7bnKnvEJq2Avj0mMTWYR
jqR4ewjrRpBaNwhru9ESaFSI9TcwxDV/1YvbRatWSTJ9f+4KS/Xqc1SxKY851sGpdBukb1a2temn
TSyMv7wpTKoDkyN1v2eDFlb/jjfi48H6xmk6v/p/Ps6XteeweGmjMdcXearqlgI2sBAyyu3NU0yy
CU+lJVarwp/ohmbEw5MSiUfwIj+QyC+0+C1sIpSGXPTS8/JvwFYoAh5KGuSuv8a3MSBNdBqoGuqr
pN1EE5J1ON1bNb6JMC/UkCv1QGOos8xZwgi2uyRAPjOIyOa76ApgNTYw7GDqLVvclYwY4BC4GTb9
Yep+sgVusO/bhi1DIYO6fPNuDbNrfdc8qGbJpV33Ahpe3daR9e3EV+I0TF8gRT0oWJa4tZVbuQQb
zkCMShalR9/dXO8HPopA37YhkY8ASBKn4MMIjuFXLw+bjDuR98dRLgImY4gtxnyO2h14lE6fU0Mi
mSYsoIwtoqU6oIkRa0I+2DVRY01oSXKM5a96PGjAlR1L3ZnjzIgPpYaxrAbAjHDechWTIzAh92v0
VoebasZjzL+ic/QWPoZhkQ8+W8lSw9wht8yTvBKLjgpBABr2yNXf6JUtScwKMUoAfTLhLLOpnm0R
BVQk7ZM690xL60KUZGXTD+cgvCpF/IZNck8KRjEFpi0NW6fAi62oaLT2rftujEnwUcHxiIZut7vf
InvI+W4g0wMLpD6etPHZjW0ziOF83Ce4qFziLvqoykA4+YRuO1xh/7WZxscP77llFHpBhXd8UcVO
CahZgmCzMfReKgRz9L8duKMv6MuI2qR6TfjZnit0E+NB7Fnj27EO3MyPMxahOg7SVtADvp/k2BX5
3kxlYnZ5oYEI0s1pDR89SimpPscnUhs2fWFQ5mKjcd/mCV1DNbQjLEXTvdQIMsOz1RXrFX42mOzt
kCUKRCnPFsibUzMymgRzZokymMmEH7fK1PAPmH+BiNxzSYZJSWtnEahEcA2cGYxjHoKCOaWdu6Ub
DwgAH0Zt34dPVmYGqCc4VcgPk6/bzPNL/2DRLNN0L/GLHD9pRv3yibZ2qKMvYC5KN6yTShCpSY+C
oWMKS35wwTrWeZC2O99R8QR0PfA66Fyt0Tz3pcBji+BonXs5eEiJ8dIboYqcyc0bBZoEfEwy6/lC
bY/oVQJPhYlNjSEIWbHYdeqK+U+WvwbwuvRkjNJ/DggnZU6wsVe23c9I7AglN4BXEt1Iiz9Z8Twg
Qdaux7Ib/CHZAmjuI4obRtaNxp2PDvf3lsP/qw03YXrEE8tGQuL6NcTRCqxy70204RpLZX++22Fj
I0wj5fPj3CFWxLAG4BuFALxhzeVbukbrZQsZPy837QuM9X7Eq/LLWoxQAHGamkmNPzCrFWGsvzEu
/VaVurSeZN9FqnV+m8DKNHCDvsbH6tFqcYasnQaTE1ggMhbKVvC7gkEXmt45gOLAJgS1jsjCLEiS
n60v6tuNt+D9FbpOMDrrJSI1hhguM83ddfvg99npi2CHLJMhWCXEG/NUuv8gs55lWu9BlXMcV4KC
nTi8qIk8ibJjWdwnnqhvH3W/HCi/SkxVvcQ6vQxQy0QirwgVSwOwGaRSCDtuAOyYIzcyExYc6DNm
8iqmGSQg5g+tzhYaFvjvma0ZUd+vjWHprGtCUWVLLdfb225WPGvl+BzHmapW8m0kF3JYcw3xyQCN
oTuaCx3zeF79SAs3vwHdhhxPeaiw0CUm0Vr5/fzo0HEZvhaDahoqYw8uXNNO3UnlNubtc7voo8C0
ZcealPo09DVvoKb9xN+c9mj2KrEGLVzzrrwMYcCglMzWZ+owyPk6/+7PAHxXTUlQswVFqRqV9Xpn
XGGDTmiPwterR7it8Rkk8B+UC5qZSKlsIc0s9d06Y/ofLaYLQFPonDUGl9E2rZcWXnsr9idsr2YN
mnXHY+YwO5XwcDoeNzkfZKd58sI20rFVnpa38xJHwyMEA9bl45g58cA9pJniH/VuCoIP6w3jX0Oy
lLmndksFoesr25m7iFBLCr+OFdTV6+8y54BwvlQCA1E+Vf7RDs3eVJUZjIgTFtuO8xCmqLcQAtlO
tkSX+8qziEzYVf85Y0eAvrtyUNSUVA1dwO7/VfRN1MMzGCS+M8I9bsj8IlFD5duqDaC0+RNgBXM5
yykonix7Bjw9QNh/HJeMo3VJEG0ei2jEBF+asW3tgvwGDnwsb7m0O4h5TLI5gUwB5MgDAGJ6FgOE
a4rmWScdtwDUyThBjrmmsH0RYt06Rf2eHoPzLCBVr5FS2eT+2QCUl7kckou736VYK/xoY43h4RiC
Wvs4n+fn7bPVA0fN1isN7SssGNzZ8y0WVO0qlgOYuIINOLuynI0nD5LkGQSEjR5jSjTMzLrR9J6d
oPaZkXebd3DaaWXn3Nzq/ykmbw145KJ9nHb0R0E0wDplRFO10IoM386RhKwQr+HFtpHom3JCCM1S
bKT5pJDaVlO05qS8cMTuemjmrE3QiJsjGfrXGCD3N9JuVVZHWcAcA90RuPZeALelFUUwO8zYdBpv
VEcZNVeftcjtHOQxZ9/ugn4THP2Q2eHQ1smgME5TsXtjZq6pyxhVMnHmPKBMmxG3+IDPgLHDjmid
f382YMf/UW0tRZNlAH4MTBs92X9OLJMNXqordgi+PibSBg8esKDBbT+YNE7wVLANIzQIvo0LuA5R
vG0IKs2L75VB3Q1Nq0q5c3Eu3vsLIn9HX+n0HfH0Ax1c2woVZQSSX09W836iq9cmCitUVPprRYnV
GBiEoRCpliZWohJkMM3ZWWIPDk3Q/sR80jcwnDo8BLAqJ+4TZrr38eFKCbtdFPbpWY4IPdobsw8R
N60xENtbHjKsuj4WmAuaUM+/eEf8e/x16aBAnh9u8gaYs4r+D5FonM1BJHVEaPCkLIWICcwTy+/M
DHMTFh9ptpOtB/Cyx7d0Rd/257qmtm1p5uLLdVWM/b/hOY7cLdAxgUwHlW2zlKcSSVagCjHaPzgG
PihK4hQ3f+gGGSqyPRFsavUsXPKo3jpyD2FSfev0+IkIp0O6zUW6m9Gpc35w74+gatYNeHDEH2wf
U7b6g6fBNZgErbC1IM3ZI+DQZNVa9TQiEs1H9qf9MasxFoA99Oteq5tvnBC+GoyVuWemojEP/a8x
NVPb9XQ+kX6u2DWYh0CIbjaraaEIyC67RPGQ9ow4TRtIwXQwOaBDMqAl5Ug9fEo8zd3M3skmLUep
+BUKtAxyTnlAsM35ziHn+Id9FQZ08hNFQPHMfafEBalA1wGFtHw3DX+aJOeiVqrX9w+hkP08VXIA
5ovSWE3dwbH9cR4LLiMWtntQJRXCrBJFuKZ7J9btWQ71cIm3HfaBYzjlVAvIN3wPqADFjVeHP//h
l/gRbW9LyXz6JSdZklybVW8xYvvsoLp9UQX7sppF6OilxWrZxrqOg+5dF6QdWBvS/eXSeBoOX7US
lu2LuaUoTZFNGnVjScCtYWjC4mmHrbi3mQZ52mNa/WXgJY9u9GwDzUkhGMb78958Czkv8IxvW5YH
EqecJsgiOfiaMVUXNaVX+ciLdeXimBxVpcTvVKhHCqUmtKxTN3h2qK46rrXJivYoHQsasragwwnM
MHea9nhdigZSwQDgWRfw35Dem4F315hc0ErIlTIux4bFBQyAYcmk9WiVWQq5AOFMWEXqjWBPAVU6
ljAXMi0IHMmDI6n7HBZIpF5q/YMw3EB3NrlEphNYRE74z474/OYvNuVp07xQFDZoM4zTB/ZyhSHT
vWADsAoJzjSiu40pd0q5E2u1V636HwXAzO+ZlyVD/n7YNYLQacdhIEz3atjd2wq/ELZ5v7cMpGQV
W+nyvNvHVaWEj/n8cz/b6PRoc7cO6I0XtSACkmD5WSo4QLrUKLc7up0nh7/1wpXAo0Kn1uErixZl
aoNKxIP1YOQVbz/Tq3tXOqueCZn8bPt4NLMLHRQdK2Yt3ccICEaL43Z5ImWSi+kxdDLXbjc4u6RH
p9z/OOJ3OySt7XX78wyVvR8jzt2Du7Vw/iOU57fgNBkM6Xb32N/HSUfRxV6nCJZBAsOdgdBo0zyO
ppVpJrW5Y4h8aRN+Cx4x7rcyzvOpx03snD8yc8s32voKkSheoN1xz7SN9zxRuD1rBCReH3qGpjZS
Pj4rdPeAUVl0hSGDed0FjY1t+akMZM/K1beml6FQz2wTnrSlCiHbEFiXZQ+09Ip78WiNrniccraG
UdFRlLtvaY53+3h46f5aVbbmSJJTrzxdKJ3WU8rn60NRVvs6HGrWSjXrBd2OvT9coppg088FX4eR
ry9KNU2yaJ5gRIsR9VDMoaHj4carnF65aoBO/UR1Ct4khA5Cv8AKCbpwjkOPq+PU9fXiAUS9Tl9p
hrsflo87sfiBjIvHUz9G8BjTSkNyWHAB11wLZuifN+gHjFHAM8ak3JoLFCYrlG2e3aZxDdFwU4DH
mMfiY8XtcFzyUmQUpH58Bj/r+nW7vxeG0c5S/FXsJPQE8sAbC0qm1zPdL91lkK9ddNQGr6OLUtnq
kIKYGFBDWrSuQPOxdNlawSJzpDmOetabq6TnLPG1gEnMYijSnh4n5y2F23F+pXdJOR9sc5FzoG61
b21WVpVauHVjNIpaQPdRqkzur4x1rw8PPRqPb5Xz7rALsEIfEo1uovxs++Dyvt8CN7Y+IvLtrbIC
VamqVb6HS1+PXBVVpk4QjIJIl/7tVSnoIeKCArYpwakMur5DjGPhCg7r5N0Vq0RetjsdeDwQ+1bu
u674L4rrZEFy2xVAvQEvGfCeU0zcudb+9HQcDSLRZb4b07MmmLSuNX66Z/1YRwf1zfoJcyqZt/i1
NDuKdO/nU8uDejOTzI9C5S1OKP56A5UzTVmAwud0tQX4SJmbKZuZPGOZ05GU5dvvipWZGm1L1XVV
j3R6CYnT5Sxb6XLoWEunXn3vIhEnifmwIN88SCgql/+78hjnF8DAvT8Ms9HL7LSl27sU20VVzISG
YIK1v7XQXhkx1JD6qZYYV+LD7gNHqRdcGRSUXT1oacURbt7e2nvzxQEPnM/ePLFTZktWcsZ6wXIh
0aaGOnTg8LDf2CFRUv2RvOWePX/BhxQNOepeljufwl8Q69+aXlFhyeSOPtN9AgXdDa96jrhR4TQc
j7r+6IdzBSZjhGBr+gn3KIUMsLIa+fb/H6XISqF0bjXEqFWiirbgzES5IYnMlUDw62qvV6We+2Gq
umTyxpSgoxNrNbVsVG4jdFWH1Wafy2ZXJ0aGXG0ZeHmQkSb32ySu4pCIGN+dTMSjfoL0ZHrTsc2c
3tGYA3AZLbv9jQxUlvInCiPAQvw2Wujdv6tlJJKjIcBXj8VCtEoWmah4ochZtPtERGR0DSFbuLZX
l6wjaNRSpPsjQDEz9BWdH2VC/r9+qcuDVIr/9dAImT4i4c55vfGL3FPEoEfmS1Gzcvyr0+C83+fY
s5hLEkx/raDS1lAoSGHM6/mwNrHvNNlRQUTSFGk8s9wo+rbLse6dyV71UyVqog0WaTasm2w/O/Vc
dj5U+1685xFlGTVTQQKHljOv2q+KkBywoCSXqEcctA1a6NqpS9BE3Jf0sJTu23FwvBsjvngB6zqP
huPcwkA+kwliiNCD1u2pCPUKq2qH7T1VTXZma2MFPT8UohM/hANzScqXuqVBHI8G8bp5tv7CHgXj
FFOanHz+ql917tIK76gO3P5uWrqSj2x6aa1+D4QylYejUjP1IRbRtsmyNZ80kBpqribrFQOLrOcL
m/mQUqRhlhs8752wfRPDuXIgYJ8CRJnQIPY5mpB1Qp7Tj1zX6XMObxQr4GwoOZ4qKTW1VMp5Tsx4
RvPrxQ77Tu6jU+zLFqPmzsRncb2xUPlKs0bgfdH3npJmncCUMytDUpQiFWUFz+3K4cf+lFQhngfQ
klZkYaBEQwjEUkW7Gc5O2DOFX4T6bqSb+rcqtyISXH/4w+z2rx01N0zemQX2QYFOZRvv3du/EEoS
jymVID1XPRrLUg2SeL5IWqoUjSE3bv91Cy4uOyQUMl61Caj/reFjWImFL+ctPV14lkd1g+Dl7N8W
fU25iureS8xF6YCaVJn2y4XtM8VCDei4wnmOBhk3OKP0WkyFIbmKeAcqakRvuSLEyDMGFcfDuU6r
tQuOLQBWwXwftj267Mp/PwnVXRzf8at+TccWfy9nZlOt1z+OgWEWztEu7aDZ/Ti00lQz7Ef3X9U2
nnFvjiYQhsZJRYOU8MNNN6rp6b3n20ezn4Cx9EKVqkE1uD7vPxh5EiCk/uXzgsisUCeEA7iHNgte
0iQi/8tso7kG98M76xTSECb2T9G8tRusBpchUh6gVMZ18oDaKzFSo5bVVfzF8LvgVNnu/qdOSJv2
hAHiHnnj3aKhWGIc3xgc8kf4RAdnvhriwIEkUJHpS9/iJ9LqSnTowibocU2MmhXj31Tq6lfY7CzD
G9L6F6JyPey38IjnHPRcI9wjcgT2p5TIzrJr8TUvCDtb6YmnvBgEq4R0vz+y0qcNpTNeSvRjr/Ek
WtGa9ZIPbjJ+hCEUzlZuGYNmS/15M5bRIrD4zKNSZJBDzqkkm1p3pXhtMzemmKIkmQEZh7ptgKN5
pGfb93KrFqlm8WjGCRzog+dIH/CUOpdP3sLcVeG6gWLH4Wfl+gFdB4eCTfvTN24wdW7HgRPxEqQu
fuleib2faX8wTRY2U6etxVOXutAkzc1eMtLshF2h0T8B9lZoE+aNUNJW9mwCddHMrgt8hoV6TN1d
n1lkskP7ng5R33kwzE4cdxJ7AkFQU0i7GnM4siPr3O7rIlVvuSlhbrtg3WF8CYgGxuPQ4eeF3kuA
Ov2VJ3ZJzbrnUh8CXz9rCllNV4dzPbT/y4XcqHS/kK8qfBxip2mrPEjJI6eZ+aoE2FJ26pasoFaL
Oe5Ppw+bY7SKl25UB7H7aIBW2IhqhsYjbq80cIkTkdt8ry9G6lDa3Qcsw3drdl1RKNN287LEDchB
6P5VIJ1SiHEixrJE3oM3YO+zFzs7nAMXq98v3Xe6ousu793eSgDGZxT9bWTQZKJwsgVm1raq4o7A
uoQX+ZrRnuKOHmJbR+3kbHpvsdUcUDdOAWyuWmzE1ZebBYqSS4xsQRa6JTjpQoUTv2qd7AkZkUfv
02byCLez0NstHvwhoGUL5X27cjXAwKMhEmJKGFixkJztm/ObGrySp3iJMD89WtI6GTqX4fOM1y0c
SGDuUMKe66P+ceLcW+CsvMFmWMCq4gk23UA4P8Qsj4NgonP0h40BWDxfFUESF55CmXwnuNHXXeg0
v6VdsyQIYJDxRDl8+zl+y1JOIzfz0IWMnrOIDC8bv8Imy6LDdv15saEHaJz7t/HrcUohHuU1U7gG
fDiUp6M1D9L88lYor9wSGOtdGr3RsiGe2yE2J0zdLP49eq/eMehHTUk8UQiXqfuwTvGS7hGzeQA7
Ppm2VUwS6S4mGuKp8BSrkWXqEhE35VV6LxsamSh4j0eTvk5e9c5mueJYV+Ptv9pVRWYUD2teln55
b1itf1LPXK7mHkC52ncPdqoPumsl2K2keSNFo1vTFKDdud8mCPZlkFwtrqd6dlktKrYDCjd0jUTb
nWaRotWp5j2u2dDObyO/7U3nk983TEWo6w4aZdEQpCG1fYm/i3AJog0s/EWG212qfoYX5lj1phBP
AnVUpi/lTG7qLwDkmV4vCVXAzE2T8m5qRZb/NG6SqXG+wbJ/KmYb0GJBKDek1hc0SfnAkStMcmx1
M9Y9+xBh3BrzR1TPdnbHKPYpoOvtPM1yIdMsjFDvGARUIQYo0XRC3OqWc1SiIjjcigdNAYy28DQF
fO15ODhTwkLOHnpEzqljzcwa1X14h6LI1yQktR37ED18jjNeXT8rp+kSmJ0iNlZSwzI8YilucUAD
TnZ5lYSN8WWbLt5zjrGawOzk5YSSnORl8peShunbZNajotJl1XA7AZ4F+6T19iaLXI6gDUpjD6XF
aZaMh/R4EV/NifrpGQ4abHQQAhDsDLr+5036rlz9GsACpHZ3dHlTM602qRgIJQGNFDAchDWSbW7F
zeNLdk97gBgiOLY9tZZU9R5Z9Tex+0fV9Sq8HWh+L8LxDHS52tFv1Yf3rWoJYRDdXq1Dio4/+MMY
+yg79C894hbrLg6+AOqn5pXaIw00g2yKjehNq1Z6nwmxBTf7UCfHtbE1ZZ4AHIyRWOzkWu9JFQxI
SRsCKLL//0FWO7uld46cOqANMRzi+p1ekmwyC3/IaYIAywqUvWGYjUd5uXk5ruVSxK8fsCB0Rzvz
h1a8wp21y1tI1l5is6QV3hG5XmAo7MzD09FoPDucq+4F2uVlU/9vPeAjrAFwSrXGg0TWnPkmN9qB
bnCQm9LBv6NXJ5owhtzXB97ThfzU/GXfTFO676Qmb50svoTQk7G1TeshNCZmSHpRYvpAFFr77r6i
qfu1A9ChF+zRYfJCaaHxTeGxXIMJvALTWT0NKPSIw7qjzkkYAynLzIQBzTRvumzBqYVaR9/R10kW
ZRM/rCD7H+/V3MqZnj8qmgkBfx91F1lXfgogYwxOGcgC7oFg1jBlSScMYk7iMef1H41HiwWq4tub
hx9jyiTBASjEKHm6idSjrsr/BVj/8hls6kYkM4Q0veNqtep1UouY8eFAqSTSslxEl26b/wl/wwcw
bTkkUaAa092ZIdF3jsDhE/LOTQwYnxOShTBcA2TAsiGIbzAcWnG6cmjMNIdIWTQ/1c+k9FO86AKh
2g7NArOvcsy2WQq6au7U7v2uACytIksRza6+jhQfEntx528SOJvdpnwSv34ynxzkrEfXdJzuJDLb
N5I2zxmk9a/3R2au/3+Yw+w08gH7DNoCyWFM4qH7JhviSIfrB1P2boxWKMDnVwG+1swc1UlOy1bJ
dudFsfy48ifr0pEtPaEzaN8r7VxZCscNjqYnmsqzHAsX0J9QqcbSQilxb4NB4EubH8w7gfPJuXlN
eqfU454mxpVzB8eVbNiOC7sE8uN9DJMn/3FMDjRH4TZMHy/xxE2C1I702BiK3AS1EBZt0zcyNngj
duJxxlFlYUiyYweoQS3CFgSlp7nwjmrKQ+KIj8rksmFLD9aKvRlM36SqQshlOsMkf17Yw9al1s01
yzAPSR4ujVAAAiJ2xUhyo8shCwzScutsTrzTnetjWRsHLaRWRM78YHq8Y8qZbkepXRGqvFAUBZts
yRvCIRW9ke30Rh5Pd0Q0Mu89CK4lY/VUnGH4Mb12P2FJ2z+xrK1tYKJCGfxLu4+1LlR3pYwOrnp1
hqPuxrjnOE8YQrJsny1alsh3OXh+6jpilN63lJa9wjeCFeBgX6MNypncRlzVdtnVm1y/civi8nQP
EnALmHCFBOl9X7cI6PMs4bS1iipG7en/eAomgYBhNKOSwaNTb0zo9aPt2Cnpa6fgBQ3wJ9K6e1Jz
mFkvOFacPqJRmma3rn22nQoGmuii1SWgJzRmRHwNehESPlXNhe+MdcBHQBoRkYF47YcmV+qH5eu1
4VwygKov8V3KG2fgxiwIXWKl33GRcrv3SdrUoqAUjxLaOC27S6HJHZsAbp5nJ3KR6dqzvzIItW9h
VaZnwnftub8yt0WIzCEFGNTo6cyKYmYCSHvc+qkemgJr1sFlpBJ7a93Z/c2k5P5rCP/t4oechsv9
f3eWh93qaOowZ9pA57DN7Zh4GiQRwAs7eH9xOtYL/uLmJa1Mq2k8qsGi+16XZCibxggdHjiZMTRN
Zey2z2h2jzZvlqDqTg9i4P3O9fKY9v7L775bbIPGzuCANshbUj0N0YYiQ8LnFiUMS0hBKNRZUPoq
xCTKjrKw2ePmQlreAgP0AdDsWci/p5989IRKM3m3dqy0Bl1eXR61OBBEDFIXwrLEeL935AHy54hI
Gpjc3sFGzd6GxwbzHXkhI3flF+EYj/flUFNaeyPS7mzII6RCcGeu3jpXAOi5B7n/p5ENNRG1XvOc
ywKZS5cH0L2E114/VD8zBfrBWQrh6MEGXZz6k0BjaP3KjoAT0MTZebrTImVpqIBKGE2cmajakyEZ
8b06P73mnP619ZF+fNZUUu1iKgz/b2KmbJqttZyIfQ49a7h9BFmMu5XP+6sHmOUT6rpP45TqD1Is
rrJKrSdUi5nResHcT22F0PMUGbwGh706j26C9d85liUGF/ZEOvkzjp9u+3IWMeVPOKjv6RVscSgo
xELUWeho3SE5SD3eWXlyy/vHFiQ7nf7Y6lYJIf1eFWSa9/ibRCFqg+Ssi9qlHB6T8RIfrbQlpGWT
tOkXCxhXRZoGF/wdrZ1jzOrz4l3GQZqvB5kam6lFIsDgHGpwc8JJr4M1e8z5odCMjxdZp5p9mxkR
AUs7EZgo8anXnz1fQ06XrKaeSi7EkPJMUGLse8v9xN7goUbeNSLth8d6E0pZtYZ6zmWio7MDS4IV
93Kgh/nJ9DFtJeVaJ36euQBKCK+ij/8Py3TEhNQTvQn9Ne52q4b7vBfGQfHE8dT3Ani7JdeNtQRn
nJ43JkqCrO+RagW1bF4Blin62ddk+hc5j/FIxXpR2Myq78OT/flMPlqhIPlCotxI6fKeAd2Boup/
keTXCPjkeWbsjjCd8ZUfV0hu+fwclygyQqOOhQO/BR1LtSxieHWUkNy1Eu53b4NH14Daw2h3kDWu
Jm+0fBrlRYEjSQMD27eqhbQWFXVgi6SraoknY7rEk+sDuNXwy5DzkCxwkdGOLmV0x69NBoenrbuj
6mFMM3ZiTqnYel2texwpJKAUJ3v6Mp+Iv2gyUhrhby7oIHwdxhtZ2i8V6QSgkZDlnFX54qHR5tAD
ZOn2OmvrP0ThE/IgBR2Tk6B3wxREHvexgCrYnMut9dJQOJ/KJKyFV17Ew5GWRPiwta4KTvzFVvCn
izhc86R/UOTaL5C3qI6CULKFA9UA23miwqEUsTfyS4X/CVcUZjWnO5rrSE2plWKLPwwIEjFfSwW4
af4w927tHlwl3V9DnXSsFsea5KsDWb90RGswgqpdRYrjptUeksEOdZXDeJkWnR8Wmei0nl60uSbN
ygkWFeYplwc5JLY/CEq3Vi9gO0DnLw5wbHOAOb8YL2g/qIMMfFDmJMGo+KZRQ9rjjPDUHaVoJs6R
FQCGtiMLWBT4pt7I37DwSeC2qYjaDhgYHDSAT0axEECIhk/T2c+o/nJgFTtdKyFTyXpohOxDKpq8
1zRPYKdDFur0Z/VZb/8RpJ80CZltbArELB+swoTcXdx7emPlZZn+ayWtdhac9FUgGQkzb3OmmATH
cex6XViMjNxhhj6fAGBI1OVRwa6FitOzvp8dm1z1QcxjDhS7FzjDzG0km6auIA9Q0eqxzZPtFCVv
6T98FoVDZWVIPa7jfd6M7hNwboCUkDcLnusyaGMIxIvQVeFZisVcNLxETLO9SeQGpSObmRTx5RNP
SYL0iNzewfcHvAk5yuR4W2JNMgesjnIlQ7NZwU/G8JYhWc1h5jX7cbkDfuQysvicmCaT9NCegWMy
UFjTqTLD18pp0aykuVfQEwJOzeTTDhVTl6HbbOKsGRcqsHnW4Ym1ORoqmo8OrsOunfSpQWlXptG9
jVtgCQv3azUctD2cBlfylBkuLZP+g8u/+zcVIl4XnkkQ0LTHKnM9OGBac4LuNgxjEx10RIvxat8N
7s/VYXWwu+cg94NXD8KpHtLJxQSGYoyS17BOrZvlbg/j024kIUkhHPgkOMqc+FDP4u6oNjFHGpz0
9QT2CmPkra1w1FU6UepxumqRjrGiqz9HTn+h4j7a+p7EtEnLr/joj0Jqq+oQXpoYzDasGMQKo/7j
4c5iBtYE2wzhH0VhEPxcaSRjtEhSjrFA+R5eUn4NQjvvPD/doolPXM3Byxyg7NUGiaJlYoNfMecY
Anm1ASL9NuZHIPnyQMCuNSG2mRSkTb2YP204KC59WFILC4aZengHcypQidVbsbvzn22U3RYswZ4A
aFVU90NShj90DsANN+aMYciXL/UqVQrl44Wl9TYv8eDJj1sx2DUtf0WLIKrtgqS4/SD2eaL8My0O
uXfALdTM56t9W2evx5LIsCv3viLIN+KUe6QIjlEPd8zDwK1Ia9Qfe64wBrbXaS4aGd3L267WYTjt
5D+0vohQ62O9+nBpdNSNm22Q1knYfjEDDoJHnp9a6C5QDfm8B2uj+LEmqOzwZCSOas5kcgeASFXs
vE5+/tZ9o11n087bPHKDvwxMQf2ZGhkPWkVKg7U+fBi8OQ8BlkH6fmtHmzAv0KGA3FMBZ33N/rR4
NNpZjsLdRjhZXjWTnydUnF9JxGJ3U+mP/XdkafS0yoK+qWmKTUqnfAS3np/43+wLtMGmT1xfr4MF
KYh5rFv58nGY0kPup4qirw3FwFhPWSdFGdvZkZs8UuyvGAZdAWBlslr892H7tClqCCcRnsoVuHsQ
U8OKT1U+BAHvZ/rnhEaQz4GNwraoJ84ZUqRiA+hphCHyAmoqc0iXUVsnQ3G5Rs/2TQf5EYsQSI7E
w5vBgvkpuC3al27ZMtkKvWeYx/SoZx25g3n7bChFTiGU50njSU/sqOuPLIJxmC0Faq/uhdX2Tbzr
K7x3G+ZsHStzlk/u9xjnMlLasxyA3e27f/rcRKWJc8PEYtWrflKV09F52gE3Oi7gXJGymxucoBTu
EBmkrZzUfiRlQPQwJHviTC38PtySO2ka7pvGWQ+8ta8mY2rq46YBG6qx1WvaDhtVEGyMqD8Xz3lA
/Kbyr74JslvMm86O/7xTqoz5bnerGquEi3Ja8KpWmJZt55cg+12JNctBASuF25+xs/Vl/ozVisz7
BL6cWPGsQBkz87oVAvTcG+SB5BIC/mmRf0HkEO3OT0/jA9xpyCnQ62yec3WBv27s4tdGxyVCgpyE
SMcFmXkHhCVT9NimmzClPEUrpaU5GqBF1x28RmNzTFH4TlfhAfCWdccBQsg8ztTM8hE6YsbV1zNE
5sj6fEHhsu9DE5UJ7O7+Mba4wfwZUiSOR/X3HTdfdMhgO9NP2yOUkCBGiy2Kep3UoKImLW2mUhK7
dxE+vDc9uhM6RTjKOIB5dPBAx9XA2MnZpyfHxI0poKD3wmnND+Z9iuTaAfzbi3+ljN/bU1pZXk/Y
0nfYnrLQYnQrABcQDWRzwTxbMk2xvDsBFmCyBo2qMj457syp5NB1iBdakR+digr9kTqPzFq3+dCv
YPSXIySmK5KBNrvLDTviJsTMf7e537w3tOgfwwTwxGVzxfkrFNIc+s1WEXwjZNDmIt1bnCPzFfun
35VMqJQ2Tj4kcR9Vb09Rip1KFWcV7dhq2mlTF+nN7PHQW/qFgiqquvvgS0acMsGPX+RfwOxIZWlX
nu5M3U9/ThbFUglPHwW132kDHuJvj+0P/iwGIgPNK6W1+bwKQw3F+VUcRS1q49tV9QChuPJFiZpr
cMet0Hw5GftpnZYqPLkFHohw8MRl+8D0//Poa3gBrz9TuQYT9FNiqzAqC3vGFLrP0GVrURTtBiQ/
oa0SGkNBVDNG2KWvUYhc2kdFUUH6NenuQ2O/KPJorQkep4yYJ6fXrJLhsDohNcxkPPIB62bOJprP
spfAnfvwy/mf/pXWcwiueUfh8PWCeDZeLJSVeNElT5sUxbqbf7VKlYW+gG8MVkziSC1gJZj8eX9B
ozbhZiiTc8SFK1SGiuVAHbor9tp52JDrtGdCOLAoBXaOBW6Tp3GTH63E+0Y0LoiV+ntwDh7mkh7V
JfWfKsxM5cII+el9pCgM3ADenw41HDBmLeMFaCW5BjX8VxUupamJpk7RAfRvSI/Rvr3cpj0JM+ar
0yt7MepC5T98JGYNwGS73S21u9THidw4ETjUngEwkasyIavU76iFocj6vwc1K16/IFuZ/amAuH95
Vmx1N1GBzaqZIaHpT9J0dbFK84DXPXrZs42b8U4fi/7I7DtBNlvhSvsa6Iz3RFSK50cUtJrAOaCb
q4xLG8ShkFpfrZc+DXD7ooDpTmT82bdlh83WyaVpTtvmKAIGGqVAducunPWzqYwcRY4ejoonYZN/
vsih81kyS3UYM7QmJEVXl7/TxmWEC7aM8fIMRxUBobZgUwHZPCyBcOXPuOPABySwroh88Vn5vp51
JbECrXJgCCzUxTBzsIQzMPmp/VPeLCnPvNqDUYfpfKu6YEJMVIGFpedXQdkChjkDL9sw2ei2BxRN
odbGUQxNKC/Yf5FbwPaEIDxvDFLKqK1ts/iKK51CWqHrkiq1krIQ5nPoJz9GAS49b/5tdQTYhbtR
B63iLvjJs6VIWitddCXpNJR8vPqKU/Mhuc/L0mMYNtZ/8d7mK6bx7GL4pguzQHs3dYykhFChM+lh
pCP+wiAoh6qTIHxczeRrW4rXtdFYGd8cOeNC5IRqIlK77x1MYDxTWzN8qS2Mmhwk0Yd70vaDD17d
QRyCQP5btNt0auhj+oXLhux9P4EcGxPHczjP0EhlghXsYj8L673zlCcLaQjUoZ18NUL4gFK65Ivj
f/Cg25KV62RrpifeuSpoM/cGPA+XawgN19yVBXLmeWEL82pg2lNg25flsJ0uzvBCaphsyNGV2FbS
AysBDzQPyv3DeHDMs1BTaw850BEJKMk1Kh1HTJj5ZM8pjTfTFolIpYK35AArcH2VyDQ/32c8ffil
H0rvBF6kIdFeOFRj2diowQlF0LeosgqLrbRZQCUhohQpbeNZsh18xDjF6TftCEgKexK0uGrXW0/Z
hlco5L9vwfoXNHGGx0meneqUrhfoZFrlRCmPrRlTuaUuWtKZW4PbicsARctedwmJvBnZ4ZhgoaM0
SJ+/SeI5ebqgPFMfn/9XMypqcA/Xkx7f1W4D5RbpglCFjqUHh+uNr/xJxlxVmVPE9XU0bwcDw5ov
HOMGwP1JaqeKrLaL1fc7U9Dtw257iShNITpSBcn1m5NZF2ALY8O3INcXin3P4b4TO4S6ZrgtDRx1
ET0al6pvpfC8kYn/inaiwfO2q8x2Fo1nJ4EqjM68MVXOK/7hevlZOn0BwGnSQHd0JJZe4Vbk7rDr
gztNDP+uM8kX0GKMdMez7DxbB19d4+9+czozUIXWHV9JHq59zv+DFQ/9tIGP0bCJvEfpXSkmHkly
g+MVPUKaqZ8nCKYT80VoEASjnhpDAt2vunwJ6IFdHyLX5EUhuA2fIm5Lg/gnLnrxjuTs/mBG/e2B
UjzNz7/VSxAeHX+ndQb+BU1uWorIJyTyGrhi2pBdDEPsh3jS74RhM7EqfNOVn3tjoW+YKPyn9lL6
ow3RAXPJ4iU1T/nNJTQ/2bQb3ZbU+d7VKsacLL3YKBlXHEJqUsTn7GRrKdL/1FvFL5ucXfIPuwZ7
oLWZZtuWoSPvLeWllgwV0JE65/hRH7HDw3IaRyD+CzuRF6ZzH66Ue72p4AI7ubasuv4iH/9vRjwY
xABPFxj4zHNzWfDl5GsNZFYVByFe6n1NhE4ClgRUMtJVz3zR20Xr7eANwj8SmKtumGCgUdS4NMJG
UTvQUWvV1XmGTzqXdP/6HC0Wy9WbJKdgr0OCEHoyHqOjeD/yHSdh4/xOTi05Ao93Qop9e0+/V/kN
x7piBrHMPfmH4IVOQzXH50LumXjo2eRilRAssOVLmssTWrVDyqc6DvZYji9gLhEdoEOOOH9RuktS
CUNIAU4D9LIuUBwAJ/zJOkxZofQjOCE0ufwD145zs45eWy9RB1VC7YCwLi4eg/tq0W2Fuh4pYBNj
egF6ad8ABaOgOyqnBwtxtwgG/+jXPOxymGbp11EsEoMoKmlymOkpkiAOW2sSr+7pvhuRhWa7dTSV
gYfFGUEIFd5fyYhNSzhxAE1Oewb6oJTQbI1U91QgESnQ4pLRaoO5W47c6aIenGrn1Tc7rioxjVwE
iB9dKvWJ8HwXj4g7OQZ3mtaqACvmlU+sCy7sFAx6cb8EEuqvxb0SsvuCwtnngv8xKXwkXHb7ckb2
PoWxKua19r0jf/XFwjb46BXTdCI+on9jM1bvcvhr3+SS37A33JwY78QXNzA241wNb8PShSznf3A/
fd8ocaX2dU+fn+mFkShxmNewAGWIG8nhIFKSUP/Ijtr/DMypZKhYipQnqqFwk+DK3UfcV5pviFpO
ygBYazPHrhjgtwh+rYZ00+mMDYimRl5N+3c/ANYsKmTaJg1U3g/0Mp5Dte5p0ILGdXve27ndUnAf
gljRAhOHTheuBxrUumiG02re2/Tdb59w43g+YU2skkYjKVyTB01sF8OOGjI9zu6uzgks/OBsQ47E
2uKcoh0F+/AcdbcscZo4186Uhu/v5KJ3CSl9J4amVg9dqwBGT/kW0kVzac8u/dmFh/uZKNyHCzhI
Xd1KVPphLk9rBEo+6X5h7DvYhrdkWAN7jhxlJcpEAjaF+8RE+IJU7BrChFCt5J7p/otZVCjCXyOp
BApB7Uxz+8HixyijXOx+FgJDsB5xT5uFltaFb6iStCyexl5bIa/xqVfgQ0mn5gZuuigitD0GIt4h
NLx8PaK29xgRjY6nuqtRvx7cIDCP4BMSHazvbT49OxA9syT7fBzoKw87sJMlfuhUMNLhwjBaM1cS
k43CP2Sg8m2Kk4LRuz5b4Fft7keqFwPwRwEF8Lb5kMIMn9YXyMDAwR4jb2Z7Jy3Yxo9QxKcb9kmr
RaYQp5yLVdTmIEdeI+RRmDmEbj3QsdoNJWELZ9Qn06qGLqOP2xuj48RkMmdJTK3JnIzYly5dg2kT
YVPd7oSK6AZiQimX/NRFvJVz1m7qfPxp/lNBzHHZXxQ7BUVrQ44n7Z6dUds6jgOyreyHsr4uzv9J
v/KWX/YDobeLs4fKjPov7DBhmrnZnfqZYnLrgwwuV+k516zJ/P3O3T9F+OqXrpnJ90ruUCSfIMqz
XtLdY8/kBRkHyOymFbq31d8PVTFLYjD/CbvZHPWRggQKtPwnf+1hsS+vldHW1hJglpokieqh5eP/
SK+ftnbsyAwKVe/mykVsVS3RXxX6GTmwbUZpevLSCKvDOBfgBTDn3u9LnmCEVNWfd+fLmeM8ByQA
Ht3i8X25DdMY8SD8WKYHTexveJPD08KNRNIyc3aXByDe5cZVqZi7fjf1WmSGQa3ez/SPZrxcDGpI
3JvMmlZZJrdZqytfz/eRbwvR3sDeDpLfuVD7UygzqVj+TGjFJzon8M69Wdxi+GHOBXM+nfHJEMVK
bEeqF8zzeWkPHLN65Yrc6gab1eskwsdXfNkNNlBy078NbwyFUeaY9l0m4MWW6DWUdvnJWZdH8k2R
PvrepWdQYE2zNHNpLV0TbF7E0OcXfqcEW+ZDTLJpJ3quzyiV95ciFNOnY0LnFUbxExmo8pHaY4HU
NtWhmwRIzgm33PLhxbsByat21/4L7tHNT277QL/KxiJp5NBkYOFuwklivXG0WXFA/dyqF7iA9YuP
yNpMHCNx1yO76EKkuE9AKtQoqkUqx+NWkyyJ4nds1a77AdR9IP6czPcLKj9NPy9v8ACxBXLu08zE
/5wOLA6XBaoVkgRUMwjTAIjRZexbwPPZVkWlKIhW3hL+W0D05sehUiI9ipYaDUiZMdLVR48lClzf
P91U2BpvZ6IqWv/rTUFgX3aV+wYwb4lZdv5XeCDNQFN6zsk1e3kz6pRErJGXQnazWQKrkAbASfTz
VVLKJKycvCvk/hCXakDr8NEs/jyACaDpWbq5Q1sjNSMPBm4GvDfhV/xaxHk9AixF3XF0+EOlGkHR
RDnaQqNNEk3A170RDHlwRapqFo1OdzIjT/qm/Zxo4u4WBi6GiAgeHYfaI+CIvjS3IOIjmgP4/KsL
jp4zs21+SSBh7DEzhAUDKiySYjollq+bS4oAGs4NQkfc6LgCLFBpAMr963+H7uwYfcDlFCXIjkqN
w2zsNz695gKFJAwYb3uTllsaf5lnd9/A+LIO+0pgaZiulvd29ziwPPKHptG17C55Nmx0DPjqIuCb
k5d4xTuRPS/ZoPLAEmq5HfLNiWym+1s+WsWxxhBBIhtPZ1aJ/k/AL4dIMgPycPFnutOaFQe+AehK
UavNsePGDozhaobrph4+WZuQzVNHqtreFZqVXEJmXDMZLGBqOc843d6OPS/9duOYBgni+76h3Snn
lmypgbaGJF3NEQ0DfHWFeSD0VfH1pfIhTUXUPqEXQK4SxLWlvAFMO9oFuHgOfTliepwlKem/eAbr
FQAMry7aqjewUUgT306fWY+IRcmpeBzvWnKKVFHYdAFTbwAU6/dQWfn7D+o9YuplkidsH6FvFOxA
d8N4Sq/FTR3ZcN5giao06BVV++STSWi4wwc8xv3tD3EMozEUwaK1Zd3j9UeQy32v15T0NdO43kZq
/nBQVuhJGUns+g7cduxs0+WhSWhdsrKIUPUXkdb8Svx35U0oF8NAbZQgNwYu1wdcV2DNJYjGwzW9
SRI5y+orOQEx8zr0qkk9f8aGRXkx6UKWGC6a0VVXVZVBByxCcvbr4GNOiKct3tux7GG45pt6bUyp
/fBrFpPAxy3ur+HT8s/wseql547eRAmNeS6iG+ZURSuqt7wvQc4JirrcNTqjEbqORxFu8oeakqs5
eBGnPnL3LCEyfxMIYv+p3JD33R89O8haonZbpU2PBxVXm6wTVFGhcBMG43qpoxaDR1TbKV6JHW5x
nvCAMIi8ncl9JCeD6IwcJ4WyDKpm9wk9v/KgmTc7W2jhxlFJtKBCxPW/pIKxepqa65Bdqm9tbrAN
J5hwzjvvWxvifOalOV2c1minrGMZV3CzNg8cnJv2PyEqcO91PTbHP7vAWcArW8Ykz6ntYWLOJwpF
btK7w/gUK1fOgCLo+mf2t2x0bGOOfEhNDXDTgxIqrzPB4dA9WQ3Q6JC5sGPcj7PTAN8Uf/sbK2qH
ixPbCCoF5l2eTXDXjbwXFZurWDxyKdVIFA69qRpeRafcxlH7/pZGufcM9ytQfHEJlViTaJr39rdZ
yFJG+TLwS4dF77/D79/vw4/EwwTb+gjMMTO5qEwtuQGIubkShYUXVLKVhwoeSH/gBOkmfs280LVD
JN2vP/LH4hfY40RDrl0dfXTOEv5uya7Pw2WX+wgc6OWYlHshIslEaGpd8mVNGgq6VEW9kzmxzp4Z
J0DCy6/p/W4NcdsqywJ/ZYVoaQN1rYNapg14LIh4AJRAv6xSsf2hRvJK7wm8eB3IuwmV4yG4Sl9j
tAITb94Vmp2IUk9jTsb1cdgIDC8mrhni09faXEYpaWhvzfKCPWcxzC3X8ziKpafO9Y6ZdPHfL2Lu
0wqXILVe96PR5uK9vVfHSBI4KcYHnVoqflutNlkyLeMlPIbzQCeC7uBfInj8vKF4TvF5y6rCTpE+
rHWfgBaoEBbnlGUVHXPeyHpGY13OPjfKnnit1WG73nU4zBx/lyuCb1oPBK9pzh4Y/gwvu02LLpaO
RL27nrgqGEg6wcvtdidhnQAAxXf8gDWQFMSsb1qVFmt+UefExyJzB7Z138p7v1diWu5DP/tNZEux
f3BxqZy96NykjDDafim3ht1NhMMgSU6ORHd9Ox1Kqkvcf7wURv/cdt8o5NV6kIuSSQ17SKoHb7bo
8r6LfbNF/1npnYxWNxQXCMZr7h/99WSsMU7RysgUPM183Dujtzb8qN4ZAfSE4uuP3+drwEBcjOiu
a72pNrdVAT56igjeqsMJ00c8CIvlQdBb8EwdLmlxgZvL3dqyFkoQTWukeLl7QwWpczwhKRvxUdWi
RGbqC2AHZesEfXmpXc1ois80hrY1Im0UdF7iwvZUmsCQfePTMl5vxSqMK+pE6aA4AlPIMm3Q/wuz
taU+YoFeFh9lns+Al4KP+vzgNiTjY563xMrSfSIOHw+QtKA0TI2zv7uTjFc6btI0ovoECXr2kATr
h2Q6lSSjFIlnMuV4pWj2cRJ2X+0bJs8gtAAg0LmidoAM5Vaij5+KWkMD98Q8IsDYRoDugrsR2oGy
EsJttFVWWH0d0DjgaJpl3TT5RyxlXh8SanjLUuqdNrx0OlUopG4VCCXAC5W3gxFfoBsqIFFunHbr
Yyf/gM3NB4aPApxX80c9MIE3ZdxnwuhQq689h9fuJuIStygHlcSza12Ex/yETQ2p4IYJKuG2iY2l
DG2wLIUNJSNBUhQQO+TEND37g7CrNz2wCUUaaXMBLAwAPl/soyWyDc8WTTzNX+PWupXy3Qp8Wh8X
3o4m4I34hG0cuMYNIH0KjEybGIJu7EwvEX0MyacXzE6qwd2puONEunSu6Y65J6yeKE8aVcP4RZxo
fB87WwjVS6kI0qG3yJTF0D9XpiOtlKzSyz5Wd222th6rx9w2ANbF4QnNY5n74r8Dz8uLu9K5sh7x
Kdv3fP7K/uZxNiNgDQvUHTXQyS80bjhFoZGiqSPPqGclJxu8nlx7jXUCF1hx3Uoj7Q9T6vE6nPq0
v67iRD4qkn8Kcq4fWlAXJoWIlFN1sBwWKIu1O9SbU2dbdIjEsvjvE5yTgF3dbwV0FBetaXyvYn/d
q4yfx84BFARlhMjV9p/LoHN3tEamq8BI2zlPXSMIAnSOqupUqkKxZKWxjpKz0AK4LpII0R99x8+1
6v9+B6hL/7a31yD64YJB9lYtBAmOHMm2U/SUD4nt+uBAE5jCk+ualLcrpcXwe3snY4LXnmkgyaAF
SprM1sCmhtnhzIFiGbjGjU8iNXMJddRRQ8e1posU9vJbOor5v3pxNF+b4zAy2rVuUX4M4fIgUFcY
4y/IrvTG/ZIsRNhvezffX/zMCMkpVX8KYetJRKIynk5cajjHSnJrW0h1NdtyUhJFZsFmqhrcwTfs
+6bJMi6nt9phG8c+LD04Ib//32bkOLNdsbPKU10FqkyX8Nr/ULYH+SzkcDwb2xFDyL0eQ3IaW8PZ
1+1KAUiloRFYtvB0Yf2rxU+M0rwpVFR2l0ugqLSb/MGRzByidBRhKLufSDAsbyl+E/WE5jeArqmA
TFqodcly6PBEp4TmC3wiFzC0iYNbbNb3p2wUElKR/KMFga0+bCxsx49iWvHbBw75pyzZg5AW9+se
hNn63BzFXMW6aXlvotHjPAe0PVV+9ftpQeHtX7HJVrvHMrBwK1MXiinJAmnRUzl8uyy5CFgxVzAI
EQPj5LLiSCSz3r3LZR9YfhacjBX04FevPxOb79HG7Us9/F7bhpDnfMz15uWkMTUgEwYkVjh2YpsO
awUxv3WEdVy0DoYht/wJqKIx8Q563v0G0ECOsbHrJAhq87gcZ7dg3ZUjl7pD91uAy8xSkFC433ue
JnnRUVOXfxs19+PgitstgaVs2uP8Ho7EQU57CiQfdHgI8cpzlao7/5F1fvRwI38tw7LcLO4T4HU/
j9Q+fsYyYErDZ4VSE2zS9Ix0XfYwoPrtPwqvAWl56jFWAprX5XtrjYY6Aqrwb4U+qLeo74Z4HTmH
6tfAon7IOtMM0/nDbDAb5aSBY0jcdn4JGvUfMERWYcpuwWMCeZF3ltoFx0PcUBlFaPe9MhWqxpCR
iiWkj7BFFOcvz8CXHhapnvTrXmFwRTGkNSzjt7csByKVgmBMcnYQdDW4Vs8RPo8Gv7tzR0+HIh8y
DsvNGCC4SZyobK+N0M+qJNfcQZpA+8MBGJ6AG8MVUiULFT7kgLyLuJpI92kwoShc3lmbFJxEZhST
3j4MhDNM0schl8dLZxetuWOevO/eFsKBV85YUd7vnJXQdOG2HNObut7HDZ/CznGQ8RyppnXbli6p
vUyEnxNM9x/s9AjFsbWqfkVJCv+S6T4YJm/o8mUau7QlHvouNo8f7rbErckKgnqlqgdMMRxh6qQJ
XoOcqCEzJt0isLwmMoAWxC4LjZE+Fdz+NqctyYU/rKvlrTUF6oaDK+L2ebxiZlMgUxYUfTYOv9eW
yKY5fTs04ZiYn1yRXLVeJJRyO2Bq/oN/mFDL6Do4AxTgrHnTsN4yemVYZHDNqPq+VOeq6VXQsa5R
FURI0X/TDmjuZwJW9zQNypHdLYQbBUhaeXj/bI7+rEhVAT/9nrxHuVMbjwXBvX9ZHyQkLftoSeKF
knjL0Hhb9cBSu5rm5Z5rH6uQp4jIb2HYkrhpAj/4qygfGm/zs42Br5QCAc25eT98iZrA43qSyujl
8wZKqOdl6VSZpkmdc53pe3ync+QhcYTq+PbOs6afb+2vkjfZk8Vt522B6NGw3WJxkWELgbE59T7B
PPNbGtrT/pbaM+jUC3f0hnxYDWBhbgq8+TadDmgN2nn5RH1CGR9wdLhtPk8GVQ0cAOFWxG2WQMUy
wEn8RV3i3iMSFFoFhD6m77CqYSng+ZFjnksc7hCVlsbfsgo/hburUxaqodMRDVApjywhblhKY/6Z
alnfcCxBwx328kElOmJleGS+FEdoD7xhlDsdItV9QcUeQaIq2265nDsVU6JG4y4bi+84L1rj4WMZ
/yc68QaGUN6/4vZnFV0tORHYrvbFeP0iZ67uOrRc8xkGZtVLhMjZPxqZ2EB3bcCNY2xUy37YMHPx
aCv1pH54PZu9fxriI38sSeQndVf/kiWVISEpyrOYf1D57k2AXtmU614Jl7aEauWCPLkUE1Iif39Y
+bU7ws/uCEmUg8pd11SUswcD1j7/e6bwAJBzIevmTO0hq505tbv6Vs5emj4zkS/nV9MRGrC9Fs2m
D5weP2li6yuW/AdqS+ymwrRIqF10BV6lGoxCCQmetvCsHdLI9gv1Iom21m/MEit/f8upkBNiLOUk
7bn8Uf8G59OjR3ifgkgZ2xrgxJ8D9sxE4zFKxdVBuVVasE/Q3/Yik0NNtPjIp5dN4ubWUOwbiQS0
FzlcHjAePDxAHUhx0XBFSwltB/11AbodutIdpwLvcNMPk1q96Xh7oqvR0GaQPpMlfTDAfI27UIPt
4ByQXiK8E4TQ6GMpvi+PtjTB8mxQGgoEK5v+U+zm95C4GV6//MKBSbBR9OpLyaXPQRZC5ut+48p/
/n041JDGYTEBImy9rxNcLt/7h+Q2Vr1BQ5XZgkn8EhE2Dq3i6Osqctkp5lon7JsJV0FxE37+aThr
YODwqnNwHlHuFYYl3pdbeZzCnZGFSS9QR8DztGDC6NEdI7Qrg10Recr4zP9WfJfxVp+aqCg3N1iJ
1PJV628W3M7EU7kLHlbCQwcatHS3Cd6wme2viz5L96JQP/TRz5s0Mu1SGjWYYnOjtWxi/r6NdKDK
j828b/6/N9mfmqW9ypctuCCpxtZrPcnXRlkK5iQijfE05/pXmbCHPwys6nnc46UwgV18ZBZy4YDH
aex5O81kbKj2mEm5+MiZXPh5PS7PpHq9TLcuIVM9FxIcO3WNshElsPW/dZP4ehsLsuwASLTca65g
lYfWgOCvPCRiMKeKoYYn1fICV4CuRoeuHF3tBVK+Vi+pPr4rPcDMBJfb3yUNkzWtVQ744avcBGK1
dQtwajxKvw9uvoSm1pNTWBz554vm1c/qUCYM1KGb4y44FoD+ztYjC07NYsjvdjsEd3GMEaoMexFu
Xk7ukxibKjnydGBZij853zunvcjf2sQUQ7F2qncoOqjys25n1ZX9HtTZ2YCAPqoiYCT3OfqFL8nR
tRbBUbwf77PKvw5j1wADNKUWSetFWR7Uv6ExTNNTSqSOM4hXIZighfzOfZEC7XWutaVRbmH+s62q
WG/rPbm8DeFgVBH0NxrH/NjZxY/B+2EJkZa8BttZbOijwy0SSINF+c6cXdrSKDvl9DPFwb3Hbod2
28aSVNYBmC0HkgGK4cB/rnZ1wftV2vgXtvz3WkIJj3FbTWD6LihR0F8GHlm5YjVtc3rSeSrxar3Z
rYx1hO1TS3VFvoUMBjycPSSfA4N/SplsgJ3ZRO60D2aO5EvidFiDhvBSjYqDhbPEz7ryFGB4hAeJ
jqK2QWCdMgeZkA+9bhpf/rVvqectLuKlfjj9uW/k+kKJoLplWWkt4VyHWDlJtqdQZFAoSS9W/tvO
yYEAfOiHMSuSI2ydXAfZm8+qyN2cGa6PTwbYPETcqNWc+T7Qm/tPibN+aMEk18COoo8vXqQU726M
oqLodqQjFTiCSquNujZvyU3hVy0RElyiSHUI553mlbm10wKaPzjahiU4DuYRnywCsXV+gwVW861o
7uHH7qPu/POKRzHOWaq5IXpMEZAUDhi0pSk0f7zMSfAHBjALdyDHOVPfYBxw6u0I9Ji3OtV41VsJ
+I1AAtKo8hJmbA45l8EJVQxwhT7mD/RX19MtYI6HGWG0HUC61UZuWlXuKS7gWXo+YTtI9oHG1EEt
EJR8ELpNBEWIpKeqQ4svwb5Sqzj3dgBxFSCf4hBTsGTlPxgTeeho7om1k+foW44mINYN72S2bGHJ
AE2zNnC1vdv1AvtDn5xewvWn2iyKpnFFHMYgeb2Kd8ACra4dGA9vt8TFXa/qShRl4xBjjG32LRDB
HJIx/0dWRUtZ4S84yBopSnX++KrRBcYYoESjU71HRTFWUDsoRjmw1uPpBI9fBZjvu3/SivSze6lA
dj0bnO9GUffx6ElI+d5fR6yCDxMGirG8E+WdS2NnjtJfMAW1et08tnBa/DaTXoLQYGnjCpkMKUvu
AAiSbEJte8yfyeLGWxXM7PxqFGgmfEnGlqIXpH8Ww+oAIvxhl+Y5YElugU6AmUduQqUZgDpuNYqW
3mSxMuugeELsK4kchbjyab2W8ADy66g+HGZvxVnTbaaySvQeI+CqTAq0GFVukhGltoAvmjlTYn6b
WOKRWH1QeBaCNjO+OkK4/FaOHJ3StB98AkeTv/GZN0q36YvAc2saprfqWUutnW/pUfSM6/Wvpw9J
VMf/miiO402Slu9yR+K5HrCH7bzZfczg7n6Xipgz44zYim7L1J9/CLbV2aJ9zrnQ4W5oGPK3S2Md
bZYmjPpTin07/QvJMsvTO1rEHg+meznCOgXa+HjdX5BlbdnaOkuCBGeau5bmQsrU+JZhOJAo8+DZ
ki4jdxOzGjXDEiRmQglsyzb/JT7Zg8Su0FLdkvFk8aLSeUeCrXjPBb+yCNN2Qo2LPi+WZtQzOHa9
OoDTtZi4L07GOLrWXnE93nfStGWokJOXSe6zRLVbbgTCe8u2u86y0NJFZLEBSjfygGEAhXnfLXMT
QRHHTv7GAQkvEcg3OR/DbxQyYjyZt6Dqq7gWpGzv7hafs6aX9zmZhJSxll9YUK4QjAZxrs9+l4Wx
jCqfH1UtBshmpBLyDnfY9WZ8TPxPsYOSL1Cvu/3vTQUOqqVmAjPOI9/8RUxKbNKoyWhLyCv+KRp5
I8Zil3i8CtgwrVbLFvELvWVdA2WTMAUFb5UJEV3WcWrYPEYcfxD+0UtU6QrUY6Olh//eXVMMFzQE
ffdL1Jxh3qM+oECo3yc7Fm9MzUSkcaObo44a5j6CJBkEzEhV3JVa+lc94eac7+cfOcMHnH5dTEcb
aAMnz9pzRtF2AimoYwbGD2hNO3mbyZrZVoWPpTdrBW+gzVY/8Axe88Ybc4MJvHlFHju1QG3l9gsR
w5ptUqmD4+aBP4S1JXdMzCNSeFW2LFAHPZVhdQSOa4j81pHNp5o/9R3knwqpQB7jIa1sw27IlaHk
c2pdj83p/KfA83axoM/Qt56B5nDmdLTSzH1pyj6OVRTStL79hOHv1d1l/3QKUu3wRN6jDdFHUJVI
B/+NUclq2iN3vWi61MoJfFdrWXl2aBzXVCNFrkqaLcpbPjRkFb5mPee6QajGR9XbJGCW7y1pCbDu
ArTSyShnndK22EJAldw0dzaVqKbU9i+nIc9tNnmtpN0f3zYyl3cnNSkhn/nWZzncQ2MacY8LET3S
ehFtmtiHcTtnAPSgE8Hw9Oec4R2MFzhoJTZuGmnameBms1pOB0jVJ++NY3tSBTufSsks55LvyzC0
cG9DWRGyKzskuG5enI7RzRNh1nHxva/Vwg8IAfBkJmFu9oxwoNRfkuQmvSFej1A76Z8p6o3EUDBd
1TbttHVqjz2cDl9D4fOb90O3Q4ohB0SeUdr3IfRFRwY9Rg831TwxzpAAwSinse++dAq7Vl2rYHK2
bFUmanCt6/kgn1+jLoU4Rwb7jdULWX13QF1UrGSirYgWc7LXu9l9nX/RM7KgwyRYcysn+THnm9iu
pSENISXDNRRDYlas5ibXNDZre7wqmRAwU6XGbSDvZp9ttWS4/0NCGxi8yxovKpbd1rw/eTTcwJIm
YUrcOTlhObUfFAOd9sudUjJz9Kg3Nnoig9DGEoXX+N8QrTp72fqkk7mvG9ol32HgrkJeJHDNh+4o
sjIrUP7qM/1bNRCqVz0umQbnoNWThyXsceHxLrDzM21ClxvtNIcQcQdmpKuvYEf+ti34FQBJvHyk
hbu7olR3MeJ7h/o4j89UKmjInad98N2HaCaDeAVAXCr/AVDAmwVY/tebF0ZG7qhcpu/brRgHypa7
nnwrs2N2VbCNVDQmRNGWZuN95H2P6Esvx6CLnlPrJuk4AJFLwkq0v0gcWx78uOMapNFVOLT9IcQ0
WaJBnqsFTNl3hi+PM/wOXhp9m9ZqRXSBYhkB4zFiqQJFh4S6A569D0PQzH3BPimPAVxmdNA8VFHJ
3o58qj98dP2F8vm6ml2fNZiOt+3HvnM65Q7bKxa2cDi+oPT7ZYMTBAs1edJ1H3Q3sW8Dd6Vrq3rt
/Vr/8kVHn1ZO883lBq+4tUzWlzIdP1jKDwWycrzaOR14J/8SgZVFgrOR9knr5iAOV7gHqVy0eg8C
ksiZcncz25XjLWg5r4nWi5VT60Hv56BXpPiwmHgn/HDY8wxxKdyvpoPQn24AYcgjbUA7ZNwC+q+M
dPlZzMaewjKamHE7kw3f4FY59nYkv+567nlnsAE87965NCwHSKyjpRnjeoKiCeBZsC3crolLTjgU
nlDY7awW7uZi8swhB8nSYPXpjIpNKRqtbTmGFy3R/RdKcy6E4mSAk41gCimU3QvH7deQ7cfnhyTi
2XUnvCA5a1BqmTc0dJa1GvaTWHXGverJADyVt8NtBJ/LMDQeqm5JCxQ2cVyvmZwdCuJfvg1XhHhe
9e+c1unB+HHp19zDmqMKL4/J5qu9Qa4lELOD/0Ud35w7+SPmBBYIOzmqDw3dCPRM5yIs5kr1ii/h
fUYPsawhj+ZZ55V1/3osR/HdCB2F56MVqLlZ980RRSZil8VrS+/zOjx0SC+nYU1SFcss05tBGSSN
2V3jz6SSWcsA9kZbzvbgeWBKhXzfMRY2RzTopcPdFsas2XZNT44ASYwxrnjR4dsf79zM+Xs3KyTv
NklEsffwjnBPGG7KT1EB3fM1I01MDP0HIWHc/jsL/hfeop/X+vmJ01+iNPZ6kadeaJH+rwCgT6Ds
NgzFl9dUb0Fdv1arolq7yJigi858CW/Tio4NbXKo1RMaoXL9af9SLALNLIQkTJqmFzWdfGDZWYyc
9Wsw+g9H8EO+cJFYynEbUnBpVJvTl6tRVsH77TTAx8jyp4AF/3NCYeBB03vzt3BIhKGSxJepCB6r
K7LtDRsxMUZsppoPKTx8ZT9gAd1M02Xw7L8d1rtDQolIeWnqTgOPr9HRlKZwB4H3La4DDs72tpyu
8K9mGAwzpN8S0SC3VVQTmA+JYjab7/MrVPrYMSCSDTkGK88Z5xnsQgZrO4WzkbKVeVE949gpMHEi
sYaQL8xJmj911j6R3W3VWBfwX3Vj83a6jlzZhtpd0kgEvn8kk1cnaGFboRX5RGWN/EUNfzuDHkUs
uYh/tp6milyVhcPpsDTTB0zIht50HXcKOZUx9odsc8OQv/1IHQE2jLjU6agUpBNK1P3T4upAinvk
PfKZSqijAqrUKbgP5zzQKB0gl82tU0/hWOfbX2Vwx5GgQM9aXvpDf08ahDHndXI/h5BL+ToO+GkG
yGQ5LBurKUcdPubd8CRCJ1u/NNZAUKdZc5OXcvqL+UpOXOW9kEURIFZDNK9U2Xk3uEWtZ5F/qyDH
qxfbELz1Azimd9nF8KYJab3JIE+r7SSwxaDDXDgsQrb7OeRT8Em0K136B0e372GHYNs58o4JH2Xp
//NYE7d5v0VQchGXDw8ZkyMXCMyG/wVc6YWc/uZO1RXYCiaN9mf5126TTL0xn7XXh6eUmm3lmhmw
qP0NPESoDVwqxofxZdjeEFAokMdY8GKWiHF8DqlEg2d884gmvU++RsPAsEyg9Ty06wHT++8DGURe
ELTrmjlz7nBSpNNmWcXg1VL1VpKqPpfKk7nB4RyEwgIZm0BOkozgkpt1L9kPHWJs4tY0S3nhyNVJ
TU2pY+Uz53wsL67FuA+26A5fScQX+NgKMvkktmCSEU4BfJaYIhdOKpvpN1CTU1pXZq38N6Zk5oNY
OUfYID8aKsP5pnG9bWlHVyUvJbCR+xFQT9Vcoul32rEZ7sLhm9g+JXQMYCSgccT39HnLMLBgPB90
Uw/Dxtl0DdqBxvFSq4wXZU4JkMzQivpTZDNItMNKrF+XWl7tqWTvU9Q3x7OAdfG7kZV3oFUiFLxg
fBPfjAmPIdmxv+z0VtjmPA2uRh/eNMcZ1dP3Pg02Eyyd4bEjN5Fo/9muFjxKxAJpd9FcZP78F2Xi
qnKFoNs4ly2AXlXqjzhRhT73Ch6ujkC+1g2FzT8BJklTpCwx22JmVEIgQdGkhTic4oorm/Gquv70
dUfVImoHvBD7dB1V3AYG0Swoq+SQsFaAXth5EIoGPV5AuaMlgRmcGvSw76Fb2QeCjuvPDuvNEHTs
Drzc6XmOHhzN7MRdepL5akvjHeqhSrAVlmFy9R1+g9G8e8Og40h5V+2Cg0U31QoR5gmS9taDXQeX
WUoSwkaHzm1Q4LUpdgS99Tm8Vi3AqbxxeO94zKPszT3eWfgeIbASfpzpjFCAAkelWC+99xW7KNe1
TE2CftdxocmPgsxXdnsvzWZdDTYcKsQnjdGy75o8W3nV/1fylZaii7LQJliM6xB0h5rjI8UgF+7w
J3HFprmVDVWfiKckHQwOFCIqjcBmwe8SDunxOsVLureM0HlwebbWaH3/EoIFgIMBhDyHU3mIOA+f
p2yO0cPpHu50LRMzjnesCWZsY8IN3D8ABzx0ge24yqBwNDFnD3TnvoQX2JfjRWS1xtKEGNTUJbls
ynGhBgX7TVkMDILZykns7dvamRbq1Ifn4G6Rb9IM0wibqTS8KdSpaOoF40kUs8KpdTCBR+DRe1kI
H+GmGcVcIUW2ED3XmfjIlu/xHvK8VY1Sm9P76RsaYk62C5kxChRbk+oCZ6CmgyuGJchS5I2hl77G
/cS521bUtL/wfvRkz6iS/m9GdMuWtyNw+lkndN6rJLliM92f3+x4cyevfBP2kjO7wlO990TV+QM5
/NTujeBkUwG3+VGga97kKnW9WNPncWewMt1afbo0uERN5jUTIIWbirtBwq32RwL9oX6JkB2REItq
eZLvecwHkvfi60uvi23uIs6+/L3MetlqR7rtqnEhXpqnFSUggVqWSMDgd7gehpMfvH9Zug6gvVxK
bhLuzxh/FV9b6TSjSh+6i2UbEU4xijxSNmhWwdX7yLEpcMelroA19iDUD93SIh4jwpYXUbipthLO
Fex5jpEBp7zvYeiUnWUscJ8M113j0b7sCFDY7Vly56U3Qxjguq3CXfXXqRq4eZKLkJCSoGHY26Wc
2fTZP8iuRRC8Aha/yQ/v16f2PWOGOGYzzq7z3MfVPSvq90TPwsfoPfJNef/6jFYmw6BUxQpIHTMM
P76GOuDzdF+01SZQeKCQ5BFFz/JQgs9QVypeBknqizdiYtomdpapPMYAvufLiEhe1j50GUavYguj
4IAd54L7gt3ZLT3VAZMMJBnDBFF2dRLojkte/A2gdd+nvn6zrHtp1yxJEXo9ZTRCQzk2fWawScc0
qn8Rog1RzJp1MrnndV7XHeTdK6qZkOZ1bD1RXGDgrLbFvvxF2WbMa4y3sZP5E2OUuDHAOr8Gq2Th
JgkUrrV5gMHdNwY2RyGJoob6g4NPVZyxuvIo0F3x5Mv/uH4a5Bcz/HkSdz0fEXWrkaUKV1nMlIaB
wKi/2SBaqdJWYvuBBVBZDm+saSuig4GQUE5qoYcQIareQMi3K5ks8MDHA0lGpbRsGanKRiGvesYQ
JX5Sk8VQ/EKXzAnQ2aAU2qmRphDfRzPifkyI4tXHrMChUGLcY8zZKjW/HlurIsylqpra73y7+wqP
maWqB/LeaMFX1a88dTQ/sNU6971n+S8NW95EJbYEr64fkbhYFI1sHihilAFnbVECjtky5T0twtFh
iPTS/gQ1VcI9GfWMy6IZGENE/ZbKFBjqu8Mr1JN0ClbPkjufDicSSFND4f4zzos2SXMty3jdZmFe
HkPAU+2Co5F8dgkGzVBy+umpiCyCkKH2KwqO/RJhGjWaLXoLHVm+Dz9qZRGct8ytFjmlhWLjNjXz
SdK5hDRvYxg2OAyMzWy3u5KEr5dA8RuFx7UgvcdBI2LWs38qsTRi/jAQDAhtqWJ1UZSpUslKDz6r
7wi4fZt4mNrLXpJdPiEpWA6vDv9VXk2Z9n9i2B6FZo2ZJmfW0tJ87Ai4rKb3AuFz+6sObbeHBLEG
NTwRT9EcYbcF0hDtdbtYcBoVJfce4N2b173qIaPMRJAGFttaa2x2XFJQm1VHik8iPVjq9/LK3Ew0
eWjmyWb4XT6hUDILdoc8n7440lOY3PFGzpFRiCOFh5VJO2opPnDodTRM8tHwGcUey08jMEHoQ+Qo
ReBYpYgxOlsbO30bIQDcQYwWBHNRZznxGUEe3lcgqTbjnlexbeji1E5FH6K8uVPSYRgLGojlR8yL
VRGESaqZIh+pwNSBw2gXGmcMmoyT1mqz7KcDwJLAuHaIPOHnLS7XmwvH6f3yS+3dsfPVM/Tqb+Hl
2eu+Rmt9PrcHlhQrRI8x3P60ClhCFBQ5MQQCnqMoQFy/2hQ7DTs5t8M771gKJX05bWZF0vXLm1sA
yMfr3fa0nfUrkwC2uGqlPnYGU/Uqo+ImZSvTljeknYLKvocN/gIbsvRUoC0/w7NZbNyUWZ8wTEZV
rHkTyWAdd9j3sNU+/S5/j/hRobmuzZ2BsgBuYvvDJDYc3qiDlplrMN98UP/DyTfcr5yI4RW2n1+d
kNwPNZWJbsA8GK+H8x4KQs0oeKchKRp9E0K9PeUz/2TMKN2aFDLcWgCI2CTNSmzXzEP5u+bSGeQk
CEs5rkbrvyv889kK0MZsvdjTAhUXGslhbD1112gA8sNK9yJ1KVAl5s3ADgv43XOoNOqy3jYaWfmE
QJlgHgfdzsEWhjem/JTZKbGgWivCzXCBpqwEmSs3GL8EsY1TA91t0QRsaOUWrhuTqBYzr9vMsfsM
iU25N0NiCGRSdeZd7SLOlvbwvMOxcHNKWh6iJXxz9zmqybRAqmXTBWkr12MMBcRDChFGs0dpslUm
tAMB5FivawZR1uwBxOd4y7jKHIwQBI8iENiU6peBI+96dvMOktHNfmOCYAIpnr5w8b8G0z5bm1Ts
CrVO2+lamBn1ZgpqImVGhjhKoBPqr/Vrrv2bUpXelA7IvGoC6M0BPze13dS3aFLQJ9OCAwHtPPKe
KS+zH9gnJrHXDqJhwCmst6fWj9BA/bV0icNY+X0/E3jqqClU+c9TVXEynYZrP4DExmdMRYQKid1i
nbtTX8snD8dvmgvnwRoS4LiM0hJmIxl3KeMIw1uk5fYFNfGmBCgpl74P+3gKo42TC80EHiEdfQFu
PciOL0MitSzMMWb5dpmNcqiZ4YsXRaNWtqw1KwiQXUmEFlmGtgq1sUBNVVzFhAz2jQ5/YcKJhK8D
02jHnrn4TdqNc6Nd/UlHfuTRL+t10cyAS4pydNroaaPteNoSIeoGhjrbA5pTgzSYT/2B8hSW46ni
ccjBEgU2E9sV2JPxwFlcAipXsPGzzCK9SJmLRAJilg829MV7GmOlc+Kh7ROuShp+apRVy7HIkHb5
9KI2Nj7nhFw7jhl17o85/huZMkFCwcLy9KjjF+Yt+7cPzKb0N+O5Bgc1ZmXCTtZZBhp59nUNv2+i
3PdCuPExMvh9CM5ZjYDfsH0bVBpjC40RXPkGehFeaQApM/N2sX/zlzk9470F1+hLqOqGK9+C7cye
dmLYYog+LG81DKZh5v5g8ItKbDVHMVHUwMmrm1KQwrsAUqSImmG/rpFixTofklhGjpkbn6V/RJqm
Ae40A9/P2H8xqPIB0FnjdqMbRL4OOSFNAvx0Fkh64EprL1E1O3cZWz4TSfhJmeAxZ7xDUxpZMpL7
TAODDDMQIrCaLTDBi8ZWQ7zxuM8EIf+UZN2RxUp7ZnnXSYceWmllZHzz2tkIzDH0v2plDTllnZ5a
67iqXvazhrqkT81xSdVH48zSvEdWXHg8nLJ8MtkAAuKi2fuKo2i2fB79OSNMMAzQvFKW4G5SWeaZ
dYb2c9BbPIsU0chxHWwocFVHeh7bpbVNT+pBJeDtVXszX4nwfeKSroRSSsSx3GBTZ8O8XonMno+f
RzceDKM99AWQj9FriUugsEoXtpBw5WEjg6x1ZKThWNCq5wfMf7gCjpC97Fb5CSj8tUN2mUXl7ATe
1U/gqF3XibBkRDsxitjRE/nRwfvh4CZCghIjbNM1u6PQcEXom+TzkGhDFdJXON1bYJVroREkieov
GJD9i2XtMmlJnN1V1gB3v8f5v268rLyReuM5FcfGQlhwhg5v3HceXHsZUs+rk3CLtQveERLqFq6N
pxmVcB0WgSq0zQe5dbwSYS6vofDP7l6C7qeHNng6LTkd5rSIjWLnQ5gC1bJWFSHPruGObHd13/gC
PtsVhkU2KXbTWy16m1vTuxBGgJfwKjc2sPwUPuBqVOuW9oS0GlwTeKHCcm1jtzfbXCs9svAlCvZF
hkl1Y6pvdYUdCiJh/0j5zC3q9B24sAtTUFOLPbw0pys2xB/bwDczspVj9m6c3YBgZRFyTUqrKnjb
F4hKgnQzFZpqXAeVx6M5RJ5YxQss/VTDM7yC9ZA/21F8eh4afil5kwHfSj+dvDikJkpLeG8kGQhi
Z3TriJdYQL1Q6HFQH56uIxLmvfqR6y8FWmsqR7tf1+OQhfA3YW+/iGsgpIp86IoZBICSlZ+XZ/j6
f1qS3EY/P+tsUnfVglFSnovrw7nq4aZrV19EXQ9v9d2JZvawVm+jP7u+cQ0OBY0FpzfKlcsw70jt
r25CUtDORqMkOT7Z+F7WgSz/Xm2Zs10C/HhZMxM7Rz9eeNXC4gj45pFM7w4w1ack1RTvsltKTTef
iVKzi8X6setdNwpIeMvwNq2zAzNd22yrPuzEXOBmcHBwOBqlgpwLiuFdqR5XeJLfC1OJJOsSan1k
GbT8yJ9/fwsoC7BvR6v8dDe40+ln+F9Cp6Q/+LAycFIUh5DrDnQMID1hFPLlcK3zus37y+Hbb1jh
hxCdqAJGWYWoOW9sgehtMYvPLeiFoSgJFkaSTcX/UwbdVFhettOb7H094Q3PaRG15f0p6RctPpDQ
yFFQYxKEivoiYcnRT1nJCU6AZj3jGf0YF/H90BHZ5Wyp10eB+HZ1Z9jWExJ02f22r9wm7Dn5VgO4
WQvRs7RQ5Z66nyYi6eB7aUi56fBm+Kgo2YuGX65WR0FcEm6QmFMR+WC0GZNG1CPFXfOaySqPZP1j
tK53NcMDl9Vh2v9jpMAu542yJzqrVKUdCJdca81OS8Hds1dFc4q9IN6M6j330Sf3QdomJhPjPmgY
QUrHn/6SptMT1CXhdQSSYVm7JF8WurFPsgm08nvDZ23s7uPsPMlyIMUejdNcmM4YNSzdUJXjVHZI
BZnSicKdW1GTm+XcXx3bufL7rICxS1DOx/FDQKdG59fcQKeSssmef4Bax2TX5KJ7MuD/xiv+zo3r
51CY/gXzvwfzBS8YFFdWEASE/PAr2PWprN/HDLJXTIylqvQU1/hu/DmzWOv11LblZeAyuk3AUuk3
bvUr0vna84DnwDqXqccwrZs19gxTffwCQUXEJIYm3un7jWZ17SUCsgYKDMs3Jfsms1TR15yPdUJo
zIuu5IcGzxAXj6zL2syUfbeM36yeWrrI3WJW3Td5l6BKWclhd0YHitMWL4HMpo6mf2p2H24oiQFo
W/L99a+cabgiMyTC6MSnm3wyCbXdHaiPGseWoI4avGXux9OyFJxtWc8ksLIMl4MWNescLS/O/WMD
SLAksoADVS/dzD2ELQlDVASEtamOI5/Z1n2LR5POZMIP+KThyrw97cHcVWp+Vg2x9qIA7CJ/bccc
zIlP0F2gUNrcE5N3eXxqNJdWmBPDoIf+hfB0rnur5K0UjAecN6Tztxqsbs1IrUQHr7yiyIV7bOYA
Co0KbbF5BIfkkdfZ1lQIDV/9lBt23Zek8bJJtBSETG+tJaaZS4jEycRre/Hlk164CvUOKfTm9UAo
P0UtwaoV+et3+eeasbqSZvGQja+mlk19RKDKjCzC3lRMz/p89M8qAcs9YpLO1ZZCMmlFp6uRyfgj
b28eDIR9Yxur/qghOpi5LraBPlenUgfdVWN7FBGljohWG1ceieG+LOIeqgqVPpHzGfUiNuDo/coJ
4bwpeXTFFhgJKK5K+YowW/EyH7Lr39+2IqmwAZaXgL/Gpk7QCcm2RQuUv8Qzlyk4yk/Q6tWDJwdh
FfLEZmFJVlwzk3FzYygdBpHIHX5YE/oHj//vrVoIu5ZSkjkNaI2DANme4r0c+ZhrJ3ewZBE/2JTt
X5bsKk8zvjXrbV9snW46wt8KMV4RlvBPwhZJQKvckdvD3Ldavkq2x7a07cQNDFXjhrI4Q+FZGFXv
ogWopjGR5rSwEKGOgVpSdgJUaQ1qRvR/8SVSpPAhEMPpG6wTOAYEQSxBkvoedNubew6JGCdjVAis
91frf/1AME3iU7D3j3gQY4arkCV04KeLLHSHDQ35yxmZkPqEgvEf6n431E9pdtq7Lj6f7ovLD5+K
bcZ2jE7RgRoUZbU7FKDm2T3aQLA2/y1ioAnJAVf9ouEcs8RoYEOZ37fyrYz+wfLO4YKfeJvrx/VY
ehXVvcSI7K12FYPGaT4DzWutyP9n3Dn58UtSf/+J3Jv40pK3aWV5V7ro/ZmW5AUrRSCzg2esv1Gs
K2eOW0bVRmxaGIIw0ylvF6pT9DWYfp8s0EzKWqKVZG1spcNAtqz9CJtXhlUq5qelVBecIJ+48CqU
ntu8tFbpvZld1dbBURLb1iKcwoVy5PTYMf9KaMU0fVD7wuyq1zquS5pRAvBEs7rF/Ni08uAP8bI3
caZdJuyOvkme4N+h5+GbHysOhYUo7HdGthTnTBJfe0Wr2X5tlIWle/7gtZgHtZ512kOIiTbDGRFY
8WUp+gC/4p4ZRC90GQAs5bqWEtZOzGxxlXApMdfkH11k0CEWVZEA3jvlHcqk6Fb6QFHy6WjEDRo5
i419XaRnBIEFrZEcPY1UKK7wf6o8GUyEz7IoJcdkOg88MW3759B+n0SD6yg4Q8owMR782cQdnWDp
8WvRwft/nsHcWcu8vF2UFd4fiBgo5/iv0JdGT1VG6G4aGBz8WRboXfAWGa0vaVROZnDxak3RFHJt
n53i824YWVUfO8wZ+z6Ot5cUhKzbtkjBdsfi93Knn1XHljKLL+LVZGphyYakDqsgEfhZU7qRGUjw
gEU9eQcCe+yAHkrCRBQeYYojrllYOJPgpGV+Fk95RgQPTfLEESivlMgeWNarJSXneVuLnbuTWj0v
Riit1LmpBewx2TRJ4RsJuRLC8df4UkevPzbqiTN7kQIFerlNff5ydH93+SS19aQdMoUPht5GW1mM
R4tNbW73WJSBeLRNtA7QBCXYsGWMqp5rYnpKxLk4nmOWKBblJI1FLe2nWSan70F+G2wtAzYPWne1
MSaL1e27oa7wiEOyP1G72hT9z+kZl54Kvl7hx7NXKyn/6dImXsK56Q7n+6sw5hTRx+DPP7NXvCEg
UDU5RaqtHDKDYYjvoBpo4hj8Y7RCXtep1I6RRUlEO6FbLCF2DLde8FLZ5llSYRxLImpjkpVOavub
LJx08xudEpeCU85knLvkI2pUZWVLFB3qoYu2IuScwrWDF3omU+ZzbpZrSRF9KpXLvDmxKxm1W7Ra
66vZJGN1col0ytu6HgfsXbTCFtQB4UEzRlalus7NZWjkUpxbWYtTDI1YOWzoHvcXPwtLmcv0Tjvp
1eFoofzoVLA/nc3HtUmdfxRIM/0Y0nmcvfiqYSZbw0O8OM+FQCfqn3rU+45dF0IHjCCCACfkO7Ke
s5RILBOZsbPVE4c7wIm4+u+kME7nT44xNCo13c34o+7/QvXS55FT3XOq0F3U5bJcmd0lI+znVKX7
Pqa4y+0gDdWm2qM65qiMQ8M9mQI6UjrykP1DDzggjeP7bsVzgFCs4jXYw7PtYAYcWDCJO4hYLPe7
zeUNJvulJZUatlDHLwf62o30vaICkfoqLq0ZQ4/YOnmPng788fSkprn3e2X/Inw375MT0GK5FoPN
mH2W43T5imgxu7SJ8QzHDM6Z9LKar4G9SpRBSEmUiK1s0LHpnw56++eGvfg36k3j5FVwenB1JJpN
oyNw8RG4/JWzm5saZDicdkBhYCScvO0m6y7CvmdLLxprAxJcogMtZ/SN15m87sQ/mLVLU0+QK07L
ZsQ2ek5zkeBa2SBqdrJeCx8TfgGHdql4wr/EsQD+93o4I5W1ivpGWNVw721NqofosoxlAHy3ZH53
pIiTdWTD9xURTpZ32rwI2bER8+wNjDgg/3Gbs9hM5nOCp8d5TQmGAsWZfS14QzZv3K8sm9ikJS/F
hxIn3R5l/gHK/Pdq1S0XmCY1UzK/pZy0dIg+JsaSTiJ4jPWuw8UOJcwcZd8aSvuWyG372br8cE/C
5TsplgIGqeg1a8+KIs0FNnRyJ3Jm6TZcllfz7+TpbjTrbtlEuuAilaORr4GoAxrhfuTlqM2d3VJ3
i6mnE0QC7l8OiZ5KxD26vYVDu3+vpeN+wUeQPHzBfzagfuKK3hM3sMNDRxZJXX9Pfmwx72foGNwq
86ncBIhIf/7t6tQNfFwJ1XF8RkEk9D4orCYH2hSC0t6aR0DaCYsodpbYObESsQTJObpB4lNZuxyM
s+/HuoO5vZdavJSsHmBsPwgJ8Qh3TJFaeEDd54vHSKAZ2fZid/NTwyoJxuThcknyJEjrWGmewCWl
uDmXsxjrSs2HQYBJEXRa4xwa+bc2SR7iyGs8XMSXTWA3vFE44ZCfIZ28xddc3Nm2frA7ooFNODNt
M/pTGqGiDhvkE6yx0XAUXx3ZCI0zmac4m7XUOt+ccAPW58oWSbIHE/Y+bPSvoXvZU+oqOICtOA6u
/GRa6wWMos+Fl0Br5qb71z36CDiJfu7Ynf79YEVssTg3hGz770li07gQkubCIuqnp5T0wN3+XCQS
zK49phnA5cZOwhkOam2Gw/2m6/PWPCh/vbgrJeGp64hDOzYqQEv0xokIHHbBr0z8UZUdNEYeSrbj
JSNeAfPahwIVyl+ynAmFxFvzjAL0aDb4wlNYRYCJEO+mTHX0puzvhHoyBb6iohwSr0wO+G+Nq7Wv
HuZttLteSRuWG/HEk+hBixgVnfBFWKzueUHm8FTb9580eXgM2eD5Pa4w/NBjRs/YJWpU000d3l0c
2ngkqXj+Ar6pZnMQbu7Oz65phREgWv/1Z5rWr8TnmsBzK1obDClrC2vLOk0Pmrn2EFzI/gN0rdpu
rbzgTlWlMnKMEtCLULjwF9ijo/tNUBxM2XYUXeP++9OmCHb8d5Qp0dD7Y18EceT9Xg+H98xOZ4zv
qJYhr0TmMF+GwusI+j6Xazxsyrxta9ZMKzwymxjiSOSn9o4Lzl4Iv2Yhtfn66g7j7EDZ7nLaZcZv
HOO3IxV9p7GPLpvmZy4Nv1JCY8180c+MpKot+h/SF/kNZnrswUmUvtmVwJcEs6TRHSevAXzPsawZ
1V1bmt/RdCUhCR1cF62yV1jdh1M3ngdp6FcTrSh1l/H0oTPv9Z5uO/a5ZojClvgXJlSXuVg4ooiF
gj79juAj9nDafR0Jn7byDP0acNpIMC9dyFPbjyMcC01pbMw+kLzQFkZpYQgCAmvWcdCrctkWJBkr
P8goXkZgmaQhgmMTO9TQ6FAHl0mt3ZUFW+6ICtVS8+4B2pBKgX/IvUCtq8T8DdNeDg1dCs+tAkCC
rB2dsvVr495HONhITOU3RT1Y9KGwcApHJb9oAdqkXhp+0LR2SR29cUKijIIr/Sr7ymejdGZG+eNE
kWjdUiTo9oE4C2DNtT5Bp7Mf/B1rHkrj6weZLCVCBQmiCAhFpE7gwYNrH0+ziKBRVBbYAPu6YDvK
8rxlty98p8DGqu8UPp/NlPMv1YMXJ8TJoIF94g1yGhRT8T8/B0YgCCLBwDEuM2iFwM61zq61Ap8N
xh9T//1fArByVDbpIsRlfJNitJT8GEKLTrpCSoaC17JLo/TPgpcHWSVfLEPFnrvvwFM+/Nw3hELo
ZgL7A5hO6m1XVxIa01aExbz6rSzvJwctQB+t7Ho3PA10VepkFc4ZxJ/n2Bn/cfAYHVXifOgJVcMd
5qPggdPqowzMHmShdGrBc0fmySef0DbKDMDntfPXaudFeEsXKWB5n5RgqVUTdLRSmGxMiSSJU5GJ
V792QE4wvje5Dk6KHzYVBAMinF2WUsI/ex48OkXrc9LEM6FDKEFGKiQEsb5XJ3ZsdDm/W3ipjC89
NGLiQFvPclFgnXTcmHFniSoClGVckfbutjrE5BbpijrKrTjJkxfpcbczMYQLmLsp8cw+KUXByww+
viio9V6k60ZzmG6KbrpeFyWjtIfuRx7gdF75oalAN2MTNM8yXjQ3DHl8Qi+099+HKvd2AR0b1T5J
lxof774/9dAxj/Jnv+xv4S7aMj9/bPTfqs2KCm+0CwslEcEbwHBvhUbvSV2t8djtSTdHes4LEmMn
mVje1AMR2nfBt9lAIDdWgzEkOg6iZ6n4Ny257dUfK0Vl4ILaGosgtgvjCNnIzwZqu5mX7ip2bj/M
B9Ijpei+5Kaiv4HC99zZYCQLft+3etIBVgJD7KtNsh+in6gbhcv1K437BcCBYbiVVdZg/GtJ6uCN
DLpNVW/z1u2MyBo3w6DbLnCuhtVcVXPkQViaq2gQiUm/WsNsKd11q/TcIrk+S60dqex8JDLL8LDm
kjYV1DNm30xzuYv9izGf9jJAtKtirj9kgoU2lQsXyewAv2XVL49iNQypD6w8MLnUfTTpIu/3KGwf
ZFl5iW6HUS97Uj9mskI/iOPQUVJHWwtCI/orxWWQNnIos9ayMREYrnHpI+ZNr6F5Ao44BnnVXQ8c
5x667SjY0Ka1lG1ZRB1VHpAQM5qzR9EDYbj/g1QgHhT49s8gCYhS7pVatIk1FGVdPeTD/ZkWPbVc
FE7sNC2CWGYBDlZ5FlQJLnSl0CDtOd0hWROl/6fmW2AmqddbnKHgoeNPXHBHHaV0K2bMNh5KwQO2
G/vFyq3CJ5yRC4NpQ2GZrAs7DZHDaXiSaJadICHmtUX6IXxlJ4/I8xZUs5iFmPSf0Y1J5yIMSSx6
kMqsMbCXqpqPBi5a04P5ewXVlD7zn1xbpTIeo+AfVoU6hCfQdoS4c3di6XUBKZI20SjcDWhFIfZb
Qm/dv9AgnkowVj+7s5aL2DB8u1O7Yq9+INR2hNO/Zi2V9FNmJP/NJRKAwhxOO3BPuoINDIYRm0GE
v/rmtQitzMR03/Q9dWoxZ8hynwNGpH3pxDccfsC8FlU7uCSk8MLf2c5DyCErfeymn9yZrZBHDU6r
S52DZvSNOpDQVWh1iS11HSUfJy5zDlJetl+9WlXTizynoDqVUDcYoomk4BL+A+cFp42Hw6ND8Fts
GiZ9Nrdpf7DRecVk+7Ia82t2rwaAZI3TP4edkaqENTZ8d64YM7U6mjU3bzIlKbSaULG1ruY07OJZ
r1+PSKZ2NiA98w5F6uqapcWEzlAFoxbuIhYI3AsM58uu0IywmKaYl2yzq75easwW2VlaO9FQk+Z8
i4lyNwE/14UvRxwPU5XPmUEkvFFeNJQgI//iCvH+w6ZDvT9H6UO46TEXL7TKq/+NPtEddABF8Xjm
BpS1EH1VK3pB8eBomOav5+OLqf9Taa+Zy2AFctP/FWQkx8hEZeDrrzrnZVNUuuQqXOaN4oZ6v35+
nR/LJEHHRXFgqc/hbnYReT8rsNmMItX56AKyO/C9/wIg6kLoIMf9RY9GJoaIC0l+jU6832PtlJB8
N3WmKLdQMrJmOMiCpJOu5nSa9fpmSBIRVAt1WWBULBxYn9yic2lLI/hQJyWGjSLdBeFGIj/xAc1d
O7s1ikK2qhWo+GxyHF8AcSOf6uDeCx9b1S5cMshJaCJCs72J4q9/V+4QHLPlB20Z3BvGEJlN3mAS
qQn4VFDOAMUAabrjiZMmrRThrDJUrRPq9Tp2lzEQ3yxRDtjLzo+A5zOsrVZtLGOjTVaYi8pITNda
HL5c8Z1C6PqUkM2/2B477HGwjACxwR0JlFLn+Vi0TVLS2esyk/A6ESGBX/291y+BuyMwScShHl1R
3cWKNqRzrq2CS29QNcMVI5BWVosSR75kv/2SFA+8iJoHJ78XlMRu7rrQrwyYAthfWiEDg7QRFP1W
I9+urBmJIQ+nxA5BATI5QJaqJm8v0vVyu9gTtNUfYVwidfL6jF4g7p81+Pe9MkraPCSb1BYT/9M5
6FUMuXnCoj2cqNvxscO7IVxUjC5i0w6n9WeOAAq6yhEnUFNjYI06uLy4c5jAhhu8Ugv0Efu5yHn7
t7uIKFI/I9MjZOodrH2Dtnw+eIl0pvvoXiChwwZBpBz6rljNJPNDzvE5Er+fCnpsmpV9q0Jd7xfb
A0pR8jJncgXL7NZ4U3ClxVk1GKxEmfumaWmWSv0n4ThaZAQCwq2vXnKmaxHknsBfJOeBo1oioNzj
ee5vBV/JGlHQTsFRpcTdgb9krxmBFI9Ov86nyvtDr4zZRkpNvcRPPuU+AXZpOxRIHv3FWyOzW/Iq
c7UjFhshAf7UP/lVcxQGOS73kg8AFrclz3UEWnwZOWch1st+rxwcljvoeqgJodTVl7B5AFXcMm67
9DMbV8dIA4ms9F5wVuCtXODRE9og72utH6JMa/JOC7S9qLMMVySn7uemp+OkTyacukS1c2zZiKRD
HTQHxA5xh1cMcwy/cR9rCVyOKxytu3Js+x/IgKrRxBgR/QI29Ot7+yev4WfS8WtmOxEt6xDGXBHN
FYehS2AZ/4ByQQbkIRZK48tOc2XJvYCsht8PyFv4fUVcYjqmgm3xc+XwNtQSn05xvup8Pi7QAmfq
d90LQzNOWazK+tUC2ILwHZLVv0JXNRIo9nIhsW3yNCvkE6WwkqC1nCHde7NzYYtF3W4S0C+56Iez
X0CkJA5TAh9Uo4IvUUPPzOc3mB81SfNyZ/vPoFjJXaOStM26Ozz26I9FACDCNtzCe7SMlw3UNP4Z
OZkgxuTP4pPnHQ63ToXbACNFAfef5HqH1AwVki28Vg/7A1O1TLXIhyfscCnywpXy+mccbxT5QRCV
9URgHDlob1X7UUsu7zZ/WNBJIE9UrE7Xjv4o5EF8FI1mDp3bRxZGL5UwJ8iDBhyauIg7N489IyjM
rR0xnl/a9icV0fPNfDAAczmOK3nSa8ae8E6l+ig4ODX4eYedPt6L08m7cGmw+40NEvHHAtyn64hO
OAcmVYPV8X+o2gZAL07jc8XO1SX4KQobhtbjD8HNH2HSaCqvCsfvZaD8TfwG6H8UkYsyaBPMqoya
i+NL+RndNprr2j+tIRjGjYrYrKZHAMtGx2tpDbdmsMbHhsAcsezpv9w2ShOJVXrW9ZSCOhbrHaK2
8dVfCDSSIZcoXjdEjZXG9T+AgHXq5YfLtnEUXUKmD0ksU0UiyHXq7GRf+8Js7evPq7XEz5V29k1u
6efAk/QvbyFoiREFd+brKJ2N12ZHwBGQayp39Nn3tDhml+W+vAOocXIKtljcfVF7cX9kvB7PcLpa
ABKcFfrs5Kpjv6UjKEIvGsajbp2x1Gxy6UEOUto6N5dvwg8CPzaGpIJ5JPLxz1Rt8HR6tPrqaLXx
7CLeVOvnh9leX9dInKjGz3NQfpwbUi93TupHRbcmoGS7Ck4sFgvWrtSZgbo5kMJP62Ku/G1meoCy
gXVCJGXwfJXkbRqzzhbicAl8C3n4lhix++i/yiNnz3CEURXL5E2GTaZsPhNJUBpTLvvhXkUS1E3a
X3D6r/tAoz7jGlXLuuHYTa+2xHJph1CDQIhNDX9uZxLuBkd9ligPAoh7WLeaf6z5P8Dzkvf+amPG
WOsUHlZBSqf4bFfb59SlDOGth0m+mw3gprmZiZM/kLmq6dl+pP4Y+FRTtSi5X2EqAuGl7/N/Niot
eeZmCXN4Y/qpxBg4gl912i7aHwyHKCp+WMql8a3+QcciYoHs1DLqhq2D3G3NjKEGPCWjAR2HboW/
i3kWarWWCfKySeYMdbI3r0ijTxyDglNA2PaFDDnaEjXv3B7gimguHxidszYd4Wz1xRU2hacZTWzn
oSQ1KnoWF/iJVLw09njHOuXyGhCXR1sW0Cpa0up301AhtP67JS9i0sYMnULf5/OoD5FksZIZGOZ9
zNq1aqT8pn1C/mRU3AzZgTxckli3NW60jabAuHJN+Wi92OEjLQLvX6go8oaLYgwoyDBHGZ9Z1kjQ
GZO3HlnKddUFo1PImdGQKfMKgxRs9v+bDQKjhKC+UrHm5ejtJwyfa3XPS398QZtX6NAsljJP0vt9
moPr4cXkjvvOpYWi+pjZ9H36hGiZz3RScdVGw0FOvY0t+UsGd96ComiyJmIvZXf791qyZ8OqjC3z
WsgKoIFdjrxOk7SFYsdGsixDP4GhKmyxdcSnA2JK8fsBusbmoEADtWDgKtzZJtNXgGI7gyEhrvic
kKjW4HjwZ8JT70987cl9H5dF/NUa/1N0CpQmmy0BAr4/0dGs4fDg0jA0gd7R5vtp2ExTD55f3tT2
KGrnLG5VaFKNVzeqKUfc7Y4bTC7a4+y0QNks3zf//bquE+/AUsk3NlZgW6jKn8qQTUcKLW/0LbT2
QCKTShjahW+iQkEmajjiSdjaVSdBmS0S85r8bsoSQgwmdV1mW4mRBiIkLLEn/ihmznNXOf7Vpj4g
xpbOBHlwHhIZo9SABfzs2UvfUs1fDHnIlx3FyxSaFcQkhg6THZaOYjcRxYAjx2Zq0jF/MwdRHEF0
2IFNHP0LQzUBvVxpWhcEYPAfWtVn5WL7NTfuFU2pUU/PA1ivHLYg0BjWQ7cPFugbb150t2vskBA+
REhRWuj/tbIJwVxW/V/EGCbQQny1E8b1FUmujNwtGArOk9N/Et/laQQdlaxa49cSLrg3ZQUcxIII
azi7b1KN3uToaVmqaPF1r3Cx+Ufs/oYKfdBJz2woeWJTaMS3njBkka5QdKgQnD+YAr9JYpnSUB0G
JOXDoGdb+OnPQrJcLyGMK0QVp1QIswXHIJFBNin+Y0NgjMTjHGdhOedwd1I06qaegw8iYIJcskoh
E7HRCXegCrXcZ8P68mqP/t44NVQSmHo2VhHuyrNbgka2FZnvyAGalec1Z3gHneR9CA8tOCMLX37d
bcB/IWTR3pUEU/DHTkjRxlv7MUC20wF5rqklxAsRkQCvsN/ndNYNy3OcAIh28xElYrVjx4OcZQkB
iESalc9jyi7CunPybGFgWMpXBfKKbqncKugFMosR+fdvtbmz2ohTi+08nR4mOo3wjP6AF9cYQs3R
k2yUJnSkNc3rvmbqiUHKRusic40XyKaBaFQGwdVpTEUg8Cjduf5TJvRWvQZnQTAbNAzLKvU3kbvC
+Emnkm9KkxG3dC1xDDxAAXv3lTKiVKibePTGs6h0V4v+KXmjI3QZm/+1HAxsCspPanNc8IzoWpV2
Evmvw2YlG7HSU1vuKjxJOx7abIZmFeVe/GHUovCG6D8nZpP5jqqaQ47lHvEV+Oqnw82kA2jIQujN
6G1iFYRdSHNwTqevX7tDq78uPsgCkYbLf6VN4/ncWNXyHKgc4GKDkgKbckbsw72KZNHMPMugkI0s
W2WkWS5GdKdfktDDzTdeo0OtHYCsL++BJ4XuzzyVHOWY94p+3o4LBR7wuUw/CghDCWwR7KdkCJu6
+SFAs7ZXRktN1WosWhVuVSu23juRf84zUdUfC3uSIauPQ4jqfzXEINrTqW2H19+0onRIK8i5bM76
YrJu3tYI8oPbvP9pJO+FSARIdVbuddTjXulnBkwwkiGkcxCMrCOmvyGM/W9IdHNQEZBhnG5Ta37B
f+VgUM5lYuYT3vS1qGyd21YRSASKNQnrHOH+UJeiTPcukOp/saIvCKbpWTsn341leb9xC97tKpoD
FmbVu321RAgoPkbiphYsNLpa6GUtRksm3/JOIUXlrSQce/LPSJHVgzh2JtluN2NEVqDL7usdhFRD
CH6i2y/ArcdJ5vOqd9lQ5WHEF3xgG0wxvfqzi41gqQ7sNoqUQpo7rtHGlAIzgaCmmhAma90++0kp
0khfXmRg+9RupBRpqhjqUTSSIIIaK65yTfvHD+Um0Wuh2O8axm9IiDahSftVxjcfX8Z8pIaIQdeH
LVePeujzFhphKs3G9kydnrwe+GM0Vcemg9SRY0vB/IYGtEap8BqRIQASYNaFenHejooud8HO8XVW
lxEhupY9fuho6chF/w7hveI+IWNLq6KuAdjFxWum64vcgKk0sqH41mnLXGNXsKibUR2AeRK67iaY
mUYoHT0+wSfMQS31sV6MFi1tNq+2sBRKnWvnQLqC0dVWeioY7rR/JEmkooX+X3Pmrs61Zbr8TOHl
91VMr47G8RRBoR/RHZB+LzommHfBY8hKAoTEQQk9uUhhE6ZOV5FXc3/WqM3RepymK4yTvPu0RNCQ
XeCembAlwcFFt8CjIlZzD/Sb69qjVYHH6YNxGdtrGz+e93113fqV8FOOTIF6Rb3OA02v1h9Fy3Ny
Sc/BcEwf90qkVGGEIxFXqFNt/7HScvVm2UxWcfSp1CRqofWkv4eCkjNkTXuER5w6j5N+AuhP5TEy
/bGzA1EuO9lbABkjvKNNqs/4KGWmZ371+3hhKAhC+vZJKOOBl5hoelv9dcllaMpe2Ffyvx57CAAv
VKd/q1wwR5J0sHYEQrzdsG5u00QpilbmRFLBPfqhFyOWRs+eD84UAQ5LLVxDxJRzFAxvM7Pi/oAl
Sqci0KJHxmNUGAmMxtSXNXA4HHbw1EEMTO/EfP/a5cN0DC+reQKrCmm4kxlWjqMr2KD+Y7lYLsTl
E4RspLuYkftwBpt/cCOoy/vKJwFodgxqqLXgir0QVylpK1gqAEKWjgYy0eFR4A1hY5uQ3/r7mGW9
eR2LgP/C/4N5dJGSMojFCeJfkjJLpHgpo/wuEiHpgAdDcTMuFld78cwcP8VL5wi1FFFub6n0OHS1
gdHmxWDkBaWNK/0fphHjw2ikcsi55Hlf9cObQplMURCPhf+KNlP8sBLrMbEnUtsf+p+aA1p6rjhT
O5XeZkRjwUDiJWedMGhF1JerWdRnb/gFEwqe5mSeFORGy2Pd7HvL+lqSNISku4JkvwJilOQ4SLco
rRdJSQsYlVMqHWj2J1oLBNN0uY1WC99PKyZ2iltRyckmHxqlFCuOpvtQQQm8gDHr1DFwEGVXkksQ
RvmGgblZvcj+05bOXl/iZvbY0ehQVREFZfXw/DH3xPJhLUwA+NdL1846Odt2qpWxg5MHibNSveDT
kK+tU0iPtVGDi3XtY07zDLUFrzA1lircROLsH6L/DMkJIH/7zXQbRyY+vkYBus+ZjWFrAoP+zTdu
qmfrMDlQOF1EoLoLeJPBwZa/0hYq4V0yBWF3yKiIB9AyBahC91cuK6daRNoLNdb/MOzfpeMR9Jpe
V9SINFQ+3NXZ3RN1ISU1/HGcqFqMXia/KL4kUld96exVI+ma13YKUAlWItrKuwQMPEA1/z2gEgIb
NmwSJaz+lE7QgBOZBlkjGwvU1xcirv/9RffiNT3BWFH+vwgSLdnHIkmQ6SFx/evLDDsBLwOKQJJO
UClneAxcBZrMShJBqNidInhFi3u6ZNZC45LBCZaxNQLWHq8Ild/vcPgUxIOMGo98cvcyq3H1hUne
p6NvU5wz0j/gNHbjpNXsK8yUjclAqYu4MfqafTv737aA1vvws+OICcHm70IJL3MifviPTp0AnQy7
Xtgv2Mh9Bh3wahyE2ym52HOBWFz7cQNyDJjnMHP7+kIEDaz6+e+VR22M2AlJjfhCBxFHzWqaFPFs
Pvga7wGbgNgDotgjK2+CaymfYmgNZT4YsYqmLUQ2sczjNM6CDzgLP2bneYS6OfU0O+bo1q8EKHxZ
DBpUlE3TBT0zStYMU8TQuMjuv0N0eZPWzy4HjjN9UTemMz6VSyvd35fsFl07PCliTQzcHnX9zJvq
WpBOtdXGZQi6UUD7z7jDDQe0Qopwyocc24bSMAZ/cuFue9f/qDApJPYI2US1J02IU+dYofOjKZVf
T2FylzWgYHzW352k6Pi8u0uoqKHXldQrxFg6BJkZIyVBc10zcXDuh1oS8W64EVKRJeOlk9jJN3bv
nc1tRO6M0N5O0xV27SX4ZUKBJc7tzUC7jdl72PAoqXMFWh8sKttzoYb6B3lkrAX/B4iLnY4IHgZt
MEuLe8+ASz4VGPO1TPQ/oDt7jm+I5oi4IvPhrzWEOxr8l0NDCeD5S1iaXlFza1fha3ZLniTzcFtm
5QuZqlzJ2Q2vbS+oL1XJrAa5Xf5dTg2nrEMU8I9vZg2lw5UOAkjVm5oS6y6VRz0mjz3QAAWWFeIr
j48kQT9FrYe9qUoaSfDhNEh13Q1NBfQ6tL/yPEv83nBQ/k/ho8lIWcjQQoMcbp9ioCdIMQ6rtzkc
7BUudxSUsUm9mPRevm5X3PRugbggqFvuzgd+0fUGyAzJMPLnmTDVNqTzcQLBrPYB4sSZ94+F5bPX
H1MqZgoghnoRYZncuOO39GRh5ER1vGVPyCOeei0iX/v0DtSnAiLsZcc9GrZ6ZHbg4X6rfA0gqPFW
nwFZjeLjYR7lD6+9SfPTAXQvLt5Wzi5oKHyq1j+MKyzcoln/aLI7IBb8oPo+VwYD7dmByPoFTNqR
ES6MKsaW9OBdCf1kwTT4ezGhJtk3cWN8y67zDgjUhgKEHXUlO9DJp4RdwuOi72nq9B5BAEKBfL+c
2ru4ZhNMN5fdroVx7vFBQ2R6Pb5dWIl9+KHPhIF8oKqfa8C4FYo2Bp+ERizllhWSaqEm6AR1txpD
/+nXxpRqSX7M6GdPfqoIETBuJi9yMF/MGEYncB/5vl19v75utSuXE1FmVD5wk9LZ8P5OXtmXtcUr
9CvKHFPr81quJ5ZNCfeQMKD2ksZ2tASN6XWS5zYBSvvPtJ0Jf7QBEaMJ9RgLpjIUW130yBdNvvbl
+MEFc1Y7Bxy6JHmzwIg2JfE12t3cyu978q6L718RLkAcX2clhig0fqTyAKf9x6o5sCtO98TMc+2P
PZI/schUhhNgHro4AIv9AX2QMiNZiEnMlw/aRTxg0UHtcW+0iAt1wrrNvfgvB/qSErT14cacRHlC
i76h2R5vxZGOqsQ7Ao8DGbTYblBDfBYPJnjuFs+A5cDa+/0JIXuuNGeK/BqBP/Iw8fF/OIleOqmS
nTPvlNbzeOFOyRxhPcyF/OiG6UQBOHtMv55XCPTtWvv7vk03h4P5UIy7O6LxmzsYfh6PdxWIbRyb
6gfRw8wjW7nxRPQDaNijzKLC35jCPENjnJheZ3y4K67lJqNuKz34OHl+ZCyDUNd5KQccae8UvMcM
2Tq3JFQUQDnZEyIXIGlFaQR9+JxZITZxu/iuB3EfBgi5Alkf31O63+9mji5EVy1P3/3fhUBNgsAM
rQEaCXxe/09iNBqGSvN6lOT48z24/5JNN+q3O0waI1VGAaqNlffX3zfLpug4o8nP3dKWxsPJzytR
ECCnjeKQdHLZunypcQCJsyrZgVo/N6uJZUgmRWOLoOundjD42kqiOacxhJWbSPjb+GY9kSTZPbE1
pN6m20V2AY8Q77mf7qEuhSdmoTmvvdhCXxXZlVXgxjNB4vPS8pyPBPJutEKgHYOmBX1SqNHOtBfU
GFYsdC0bcYnOoGIc47WYv585TsDzGYPkvGZV6XQHatIKpyy0DGPok22kAPuj5eFuUj6+VgpqiwkQ
+cvXQ1Ili8IXYuhqsTvWPaC0YsYsq7rPsEZdo0EBs/5qnLJIBspNzbfFAu6va6awPgMSabf2TBw1
IvVYBs/UnAGOK4X19lDqjw7oJyButXGhnid+4qTAo0iXn1Ng9luXnV2od0eLB6QyX2VepfnBHKD4
XQ9Qa2ShKbmz6YjGOBP64HzBFrGCd6w7mtuNQLdKrj02I9IdxDPTQEgAbgLqJhyp4O43e2BDlTWL
uWPhPqvYpmDx8hUBqKN6K1EWiYgw2PV16R9HV37vNimTHq1cxSouerDFm5AdKCDRts3Nm/u0PVJM
ydJj0H5C94NTX1sNjC/hbnt9f0vfgXBqxKuIq+IT8dvN6NNTkhZ5Gc9W+winrzaf9MntCtNKymKX
FYJilIYGbxRvm7QnmO2+CkekQfvwpWYM1+2/Ze3QKFKxSMf+q50jtUHZAFHFchhSDMzFGCa9H3na
On/Z+4/uaZjxAoP4Ya7ZnAlbiYBeThUELMa/QXacSlW/hZTJcQFH4AKNDQZpJKA6iakHFNbzdWXN
cCCoLEFSsXyic9d1kCkF72zK1W61gLRav/+Hg8QSppjs+t1EIaXQX+55MiZPoNhrKBru3WtBm65n
ouZmf29Rwq8Ihj3S8GFSWESpmizASluiyf6HwOwAShBYsce07oAXfS6mtU+eXdt6P7kLb2/84HZy
04Z2nOxF8SZ5XQ2CebxMkMyWDBHnhAfTQPo0kHzRFRIE08nYV8IsM0xbdcmC1R2yKUzGr42GMgEx
B7A+p1gIb2EK5+M318D2o12V8nrS1ty3riB5zmtbBVyaiePsZ83QumtfBKjMt3yVfBZETB2hdcAD
p6DgvbCJQCEut8PIOWSK3YT2TDV4X8RpxT8u71OJe7YytNF7UV1I6t5o6gTIdOU/7Xktz+ncjyuK
WhtXB3EDJylpMvEUtk0VkTN+QQ9jC4ENjxDioJLvw7lBCEIXgWzugbK7Upxgpe/s5fyKHkAZWHcn
ne+fIZ9yWQ28Rsj693EKHqGtUdcS6Yw6TZth+no6lrWrgE9NlW/O08g7pskU0hVn4SNGm17k4yZu
BGXqY/Ihxdad3s97+fhUaxAa4u8snXvNhJNmIaYxrM8Pbx8KLdPxrYgDpP8dL1V7WZNWILHIbxxN
bSI3zVHHYj06bErb0ntO3OFAfS74TMU0Bkqc0Xz402FlXofRNeY74XGR386/eDPtCDaW5g4jEOKh
Pluxrz9tuF/6tc4Dd3aIvys+nQPlvfb5qhysnwGevYHiZkbfGvYBPU1z7VG0woVZuZeE1fqdF8a/
WSnu67qUOHLj9Xf7Czs6X/+bZLIBaosaxT5yOAIERzO7EwjFXGL9kC2fyyu3CZaVz6yl2b4idteV
Co8d0QE445q07i1hCOBPrKaqNLQ48AosUp/tErFHF8uRV402ig6dOm7MrxRp5jNPVeYKDPs24hvC
rOdDX8oV4CvEjxqKQr4gDVwdKzA5G8wQvg6paxmT/pJiK5AFdVeqxDlnqkKK7wtLo2Tk+By8qur/
yOuEC9hkdUPIjzDI5zJb7d8eZDQVo699dpxOcfFllQ6h5XVmQgrXWlMUTZfrL/m9iQe5YhhyJSMA
IB74cPD/G6KRBdEJia9JV7tUa150WycKoeX+8fk0SWR1NFf1wwlQZCIljAgIy9qrHSXo+TgZLqQ3
ONJfsGOrQyj+oiEtECsVNalCZ3G9DToAEX43m0q2lK6LEWfdUnr/efQ5fayfZ4ZsPEfeN7yVnrLa
HKtZ2rt+VxX9UEwXPNvgFa5ZmEv7kc+vlvupUvGjY2zOOIdJnjB0ltuIVffSCIR97iON0VM+KxJG
DocHpQHXfW+SQzJquRuwBsy0nJUasZ5f26IuSEXrx5fU4fK1OAebqlXs5OrtqdvnRJq60a85g4SK
HihMLZbwj5RktSuqOHk7diy81ZNVq1wdl5w7tJ+ic/jZOud0X66MNahxNNJ1/xkuW8H2UY/jVvmQ
HcDGM+8CyC0NpPy2NSxAsfybN8f8JWGxfkCGK/yb5MHII3UEGq665zV5wzxb0fKOT0jBgfPwx84g
C1ADWbwgofzLVTgfxIaeqZqBRpaTANKohEhH/WLun8TubbRNOrbr4NQ9RHDrymnGV09KcMeoMpDi
wEU+QIXrASkxcQcYghb8SNHDB9f+9op97wLAjY4vfcv63W9kVyk5d1lwiljiQAXVyVF16beT9TTx
nVy+doAxG3xI6DA10SXjJ2/DjH15QTI1eZdaljcnE5nUjBn8nU96dXAjSD51e9eaT0snt7MHblCM
GscZ8wi2tP4vd5J/riwLKAbYwHHww/O2SGt1zokAaXhRTKKTDp6DUDijS50MmmhqY8YXN3XckWx7
9HycivvYGwAYn0ueRbBMM79QWLP3uF+MZ9+fpSb4X1jgy8d4w8+PJ4/PlIy6plbNP33gxOCeNZ0I
/AuIySNu4iYa+QkszZhOFAaG9Hbn7pUadSWiVt9cgkIsGedjRRVq4Mcl+CYW5z5t8XiqCkDhVz7q
I/zsOjwHsl+txC7S5lpSnWgL1mvRe4WUFFInvBdjBsNLEEcL3AWX0XR0FLa3/g6h+k9jCgKUrqfz
gc1O+yj2Ip5RwQP1C20lAYLUB7W1Py67jnA94aXPKKCFBIgO+/K+AmU4pqzhWlbxZp9IS2iI2pp3
2wWQb0r6DjNyWsg+e1p9XzK+2Z6vkEqLRsQ1ozCMLM+LPuWbC7PAGEXKjYi+SRXRNQjQkhmjM7bU
1hnw/n12qQiYjmglxQ+Bbf3EW0mSsP2ftRrICvu/VTlACP6Q2c9tQ3MgYUE4/ZnOQMYlGBGvjt6W
KPHjmR+h+lJGXn0Y4Fxg2nwJ3QLoRhSpU+b7zHdPWJnRB3XR1KuqzfSp0KSTCsIkDqF+jJd4yL0v
ZZLXfMrl3/Qec8V3XmklqknuadEBCsTnNnmFlpq1/7W6uW3Zn4ovGEvcuSDdWj6+rEbiFeBJXzXm
r/7OpHYBECHgBnfMsEknBJAZlDHadS6dr0COREnjzRE+fWFI8UPqz7iVRYCwUlPassx17LQBtMCO
Id97PsxcW1hmSuWpucp/5L5D5vuYXQQxAV5bu9tifPRIH+xG4KQhqCE8Inyu4MJAO2Oj1gNWXBQ+
CXBP87NS/tfNc1vFKpMa4fwETrgfUkBUWQaZ+IJlhil88wY3/9Ch38W+2uRmxL5EQhDlCP6NORji
5ZZ9E0Xryas9cka0UVf/aGsvGrmV+Jx0ET4rIjYCIMHt6glOntEFcUpLl53WWIqYBP3eCo/WQcxt
IegrE91HMzqJwADyz5ohTiglif5+Mr83X6yEZNwVPIgMCEhVr7ltQ1qr9fbI2HFBgojpftZLpbws
PirQJ4a7YcoET8WuRp4TnNayi6UVJQHTA+ZU0UPvmmoG6WSxYVmPcnZ+WWaVB44ghOq5QQifKJtf
HZATO5qEom8jwjDsT4aHeaHs2fpmwpMMLtBrQELyioR/jCQgtccBJvbLCv4tC0INYPLFDgsgnMtW
rNSC/aEHbVSkkA5H18f2lr04d75IpMGwMOgfILMIf4vdz6SUSal74dzGcRbHO5W+j3+q1Qq7zApL
wRw+XArxyo4y9YhJciJxdWrwTHAU95PZF0FjQSwE45hdI0vX5S3CE+fTMBS9yzXBfLkliycT7fyY
cxV1FIoN/F2dN7slzKEK5/VsKJQOKZLgxFugpaaUmA+8uMKH/h8kbGJn9DSYUTWnQiTezGveG1k9
ItO9DdllMD7hYi+cHHxunf6BiczdFIc2/CYzCL4sKnQ+2ZpOCr6bub71Gm9lLSdHMM5JMCFJoHVT
6p77tLQTP+ha28t6PK0aLRuxWDQUbXmJg+nVykSDHH1szaSGmiIQButNnxFu8H8rZf/LY/8XP8B4
mjbQ1/yJoReIJ7dDNTT6aU9T9VjlWYbqrgg41hsgZNqxvzL+a6ItZQ+gjhW5WzKdQAWmBQ2XAqWq
bxS88lACA/Z3MiKv35iLqc1+elTylmAqh33nWFRJCRqZrrsSAHC/AVy2QeGQLeKR1+EN112m85Sl
4e6Ob51Gb5G+qlUXAS3yiGR84q/iuVwP72sppKpzTPByBmwpWmDOpWx4A1PM/iJLmvK6IFJNjJ6k
yOfB9NnVOun8v3lMsG64D+cCLaxRaFoPQ6+IsUXgS1lraGPj4mTqTodU9U8SYV2KU2jW1+CPdPKt
kZdx7vAU5xiG0F8bVaxFjTIhfWfjY+0zUJEYklbSjJ0xQTq4ds22IwlIO3+5fjrSPaFknz3OTY2Z
bj6RLkc8uJkpoz58bkn3jo/Xy0ewJToF+6PVBwIOzqJDHwpf7M+4yg883PkbiF+EHTTfdjEJrzz1
E8KXLPfouQ+U7REwuYwXGEyqBT9sTQsoVBS9EoJ2RSbRGL/ipMWvIwsRgw/dZKC443ElwRK7tAzR
SALS/uooSxpWBa4YnkMvMWxAHzKJD8Jbu/jo24S0vDzBuFeWxWdtLKY7hBdIDk/9iSmfMsqnnIrh
BV72kmWuHntD8WHquNp4RrRXntfIsGFPDjfQZbL9nZ1g1woDJFE/ktVDNrplAPGrDVorg3Cke3wi
tQokhqA2ZFxCrn+tLDErwbVg2dcfA0gXuYFVFDOwUk64thnvOPZp5PILQnEE3dejE7rsN/8kBCO1
jBTVAbZPymMElnDHo11h7RQnhaJu5KBKRChTZ0+oW5kdIUFdHLqkZszE5G4tMnnmyPX87WbBIcoX
74UbM8vQbnA8hKBT1YWffpqTu0BPMSUcSn+nauf5pQSs2e0syzmLFvX4EZUN8lZAhzSQAuKvfYy3
a6cQz2247G1ML7F8rC9rlUct2t/iuDKGATX/m1D9j3F2s3hmPNTohNaUTWubRXJIbSLBStHszV3t
a9mUvjB4CO0BI5yjPq6giCZvrI1Ui1Ye4TMUh1AyJQ237K3Sd9Hz/Qje2mg0JqNH9HerHtd8JQlh
fp5zonHgfD3H0K31lV7c4iPhVm/qCYINu6/FFeP/Q1rrFR916+Ngi9eHxeO5yGjGcJdsl+86PHV5
mYKfbbT71IbUaCZlTmojqxoYF1fFUSMQXLNtMnLuReSk4FVret56adqEoj6Ju8Hg+OVaHq3PbWT+
2dSQVYMHNI0L0KLnhRn0sfhgS/yz/loWAucpJ+nH31XIlIQXQptO2sU8+m9Urj9+sAbgbVshYS0u
NNvB9wus08vtp5+KfWsTABXyvREqt4v7D85N8DQYzy7ReSUXPZb5HzxPVB93z8gTi0qDzmzYOTvv
DoWi5wlXEzYw3hmI9A5ShjOpM2SsqCMqMiBcQVTou5FH+ILBhHRCtP+3suD6eM18C4Ie9yWzKby3
cOhk97PVvp7/95CfdGPzvfpc4MFZUB0j8FjxHtoK5MJnOIj0L06yTvItLrVbHP3KtSU2/oZk1gYH
v7RJde7/fL6MxHWw0yGYV0c0I8F6gT80yut2/WuuIYHMX7QX2Q/Ly10BWLCt1jOpwNqlWU6hHawF
72j9CtIMJdfZnk6DK3p0embO2ceF2wdvrdibLpsHc/f61mreoKLC/tqCmCkW8j08oXohTmWFTPj5
vzPh36Bl2wk6bIhp3cFqMSStirmWpdqAi/QqDYRjt+e31gKyNfbTsdqcY0BeirmpFbAXvD0zVbR2
ZlMBo/U3s6uwEhEV8GoeDEW8CvqQTZJA61TAOdo97AcGRf9OiBv/c3aNOB+y3S0PNkIlzdjYpZL/
LorcTG0UpkJFL8+44hCxzFrWgK/Lx9ANWhEy70Ev4zG5fISktTZKyGO0db47ujacQnA99B7/4iIM
OzMffFBNehvNmSOV8rg23TIczCR0M8LbdCkpPdXPLOe3165VHMrDG0+dhq4DmqIG3vNaZuikOC1H
BBdrL8JxajSpym3f1Tgzza8IEQsRVzAZLvyICmpcD6TP8Xmrxsrm42xsYDRwWgyhTFYSLZ4+Z6kH
nPXyNumgiYBD5flpDIN8wchebk0R1mh1b7UGskCXJtHUYPAVEjK2PUOT9DFUNO2Ea4Dde+MHKH99
/gsxoFbDGhJcrh9KJvvPvrHIPC9ZkKftnGGJbM0Ec1u+v5j+apQTwV8C4yZfLn/hhy1nWZkUkdmS
1AyIA1BIS0WPrADvXbn7OUS7e4q3qdHnz3zS9PKRCvhtIrVbrcxrUDNZ9K8Tzxm9Tk9ZJ7i39mgC
9oOgaIgwkHrkIooAM+Fck0tZjgkt8w2sEilUlB/CHWgRhO1YMZ+HGMFDMhGp6pmx+Y8AyZac5/ZQ
IsHHRqVEG4kseSEA2N9VZa4R+e7ntWrgHaqGcschdPjfifDhW/IUw9wLEqABOoiUPoEVSGeajyyy
F+mv4uIi1jgua4F5elxKb5MwYfJvVCPCEHPN2WEjtg8NWHjqRhSCgLxw29Pl2j3oZHpvC57/Xy7O
XBdYsm42LkwUyCeJwCAqc4KITsE6wSDU5hRS3IRXJl75SWrxXkk8OJqhm13BHoc+ttCTSROQKXtZ
GEb2bwfInik3uypvv1dSUzt/RQkSSDkFKbw65ySmA4Lyq+p+ysIfedKdwdOI7Aj8QfLkXSv2QnNB
9gEsMM6GuyhR9YBnVmV+HYun827Q4zjpsyBElVmnMIOoHqYVpl6f47Man63ozIN0fF2TyrzLalci
UgtGSbRCOCJybdBapewMgaPjdxNZQ69Sty6YBzh+8xdLfZE5n4aUl+2+I/zXered8t2DVtvR6g8R
lMlPDNsaY3sjyGn4CDnNSSswZDTcW2X3MUKPYOZAu+G6fi8UDVUQCFh5WWbaXam+C7GlwXhYVsdh
kf4HsgRUf28obi0HsIXt1G9nRrCxpt6eHrQ7hUkHRIwvZfwDaIibrx1xJMSzhfZ4nLLDapG5X3TD
FOJMcUA/wSogJroD+N5m9YJt6+uWwZxMSt2B5nhiO7l0Wu5DTo08K9cKxsVIhFK+g/1F9UBOES/o
oUU40AS2dCwuxvUcnDr6+Pr2Suo/5BdOgQBkUgAcEHDyQwvrMfKOevemFMxpcAiX7x7Lq3X5FTy7
vV8xAFPuWNDc/WeWb0JXsocwWbastw8o+2x/9/XLHTrpwUjwDAx0aKQPKMYBP/6DbiVDdgu9LxKz
kmhcHsqYXaMtkl37GQZu87THtsUHy8Kj1QnuTzkLWrFI1FZL8wFwDiLxrnGWNxYdwRbYE2Z/3epp
3BXk+uLFa07fBGupewT7hSmGcsXM9kVQBwH+RbtAX1LR9xA7HaTQz8/1ujQA6vy4a9CqcpNM3Et8
s8ilo1TNo4ZbtFBoruuYPRH9Yh4rXQ34Ftp40uw2wApwCllZOw+7tiSOIVToy9sCc4wEo5HcDLY1
AXb2RjBvuOoRsryiZ6huVD+TvenlnczgRDKQw+rgdmM9H6ZF9DC9rSt82DxltadpKBiWUloec/Ua
dpfdWpyER5as2vLos7lKdU0ydkDvckbyAt+Dsv7t3sV7Q2jhCWRbalp/6Gm0zsfd4HRHzauIlMoM
amQwYQaTtUnMqeJqxngbxFaG/0UvL5kMm3v0KdrrosA6ZA6aCV3eGqzcNWhuv89imeLPCpMsxjhX
9Y0Ntj8j4ONuw4EfSOl+fG7SZFAcJeGkk+MJyEwSG2yC8okWSZyszKCfeoFxfYdxaR/LVUKFrcMG
RhGtPZhfvtf8tMD+J6V2OkRYRfrIyZMW7cyLzxiAG2qqdQPOEg/o4jvfvxm5Rdyb0st7uDAJfnJJ
zmVCwD94z9VcBPsO8TrGIQ/syMkEyHU4m1ZzDqLVpAdNQAxQZBDnl3bu3Pzqy84uBSeXDpiUCYyv
sIqPnrgLez3bMVDoqm/9+ugH0id8bFtMPGVrme30bZxEf8HciBmm1+o2gcH0PdBr61aiviTApsM0
Om8lW1jORNPAcg9do8Mb5pNrLadM6M4kIXVdGQ9pMnz6zpJ6VKvNzLUEiWOSrML876M2iwzeOBVD
KlhGQmMp13xyJlMjK2bv0nosNAttihl29TkO+n8n/mioMYMl76fTqwdxPi64s6EDRPhEa13iyWFV
zw5wugBmZESoILdkaIE5Ye86rUO3QSm7PI+Oh7ntpWGBGAgkvb8TF393GZq1Fqhg3UWCV0brLJYS
YOCIBNgxasg9Wp8+cYFIyhbA1kVnyilgy7M7LK20BH2wRJ71SEFNgOVoWbNf5KrDeKCwqs047wb6
kATvBu/eFezyI9obduvQBhLz2WhyPIl5ANqJ6BkffhfAgEO5WqfVzNA6ICjs+1mv1uWD+e9rHF5i
WOEYA9jqyO1WT9Gi88p/aqSohX78qKW3D0qAUQX4WK627HyvPh62YSHuAD18ZxRowRFYFoXiYVAY
884YIaPSXGSlmy6GC5LUhMuyA5Zha0FX+qxZA7iJ5yDuo6hKuWRSievTBRm77wX87J4U3QtkX262
ud6nES8ZHjofLOxp1JMuABlFh0bw0ChY+DcLzhgIDn2mUbcccRLvfUeoh9mAmSXYNRW5wgUurrfF
Q4frwZLDe3W6OLlZ0cA53PWkicTJnedUU/LFqWJo1ZjTJA0WGwRcuY6JHoeds3+3aOV1xHB6yY1k
yNGyZekluCwx1Q439Etn8S1is/POsa48zv1IWGW9qVzSRd3EFbMmzaxDWXGmMuNNSQFUWVKrqj/V
4Ag29QC/5k5lYD2s568aLItNEb8O43o/WQtXstDoYDoeeh3eNGJTZpDWzEsS9vLnI/aPFmZp9EiB
yn+pYmwkqqZ9hBcDcuZNRK/zZc2Sc3Yz1+Qiwda9rKIE5wFDJXQt04GkO3l+wM55HxESAJbj5xZz
sBhQlmidXfhg9scC0RE0NE5qzBoMWLfkvzbk6ta0d/7A5igbAibhhW/nialzKQz4pkr4SIpQsDui
9VOqyCQs8awHOOYOPIYmgegs9GTwNqsMU+1sgzDpzEEyIK30PObdx0vlQvm5tHErmPasLeNuFItf
nYWkZxex4BZVnPJ6r50MnhVVIKF/3TjAv+GF20si3p7hjgfx8d0Yd28ls36jl/LPiP2NQ6DBA78a
vX654+z5OTd1X6UmYt0WH6aM/sqfMIRhgfqPG9O7kiJHA4J70H3fJzfDpNm9Uzhi2U0uxGyH1S7Y
rsD9DWAYZUPEXdq3iwS8G1q3ZPtBWbfOME+HsI5Rpv82qXpM7FX+lvNWlQALNj5DV0SflLTDHCgi
GjNaXBLM7JRNf5oVx6Lit3MyQqHKgsOfynpH/EFJoizZOQexkuWUyoUMjZ8TmwNbEvZUCPFHFBTK
uoznpl9cfe3sufDcesgux8mno42ereVMRacPFFjEnkvz7mKaCfNoHZW4zaP5DgdteEFAP+i62bP6
7LGkrrIasHK6lqQ2ssth2x0jprIFTmvEsyqoYxWABZ8Tgl0Mi8ffA0smxLNsmPaliGF9ror0sayg
eJiY90VwtGLqQ+P7PkVwv4yjDVHPEnP9vvFTAEJyQzC7gCKEJ5W0R0D6QiUf1cwL1JdFbqp2fLj3
+s06L0s6SEOC5Mh5Q2Sne9jcfSUK5mpyrwdyMeIc3bOcQSz/fF+GahssdhxltfNHGBQJLOkWC9sZ
l3s85igkBuPlI1mHQYv30OfJCBtvnboq8Y+9Ij1A0RP2LvoOhfqzvo2z+q8yt5nCyAdQ+9r/WCXi
hqO0T4mLy7sUuadeAQVxyjQkeqLMhun5LT9PRw3avfgsuOggOVpK5eOjTGFabbe4Teidd6RSZf3b
r1VmfTbQ4XjuuCYS+X8yTS4EZHNoHPxjxNxIYdnwr/rF7qfonVliSiZAC9uuhBwqLo21HXXzhxnY
5KkEdsQTXt2giwCofCKiA4GQvj+xCmBYLkkNBTRhLiLIl2KegGEHk9rruq8/j8Cg5SQNM/4M0HN+
e342p4PPOiJPoAY84xYmhISVgnLnF84O6S6PMlyuTIpD1H2R1/NSIv9eSDUJ5W36hC6fA0X7El5b
2pSHWYW3Ags1FZH5hI8Zun1Xa2A7llUv6uPnLB784YY3FXBLro5JdWSv1ojb0kXNN+ZLlLce75Qr
7yq9d8QusujQZk5QwKog6v3eG1QHEE9ZYGq9DIeSxEvoVCXYnekW/zQQgR7L2EdCdRa1LH9MqThB
/B3mdsRtPCOq/9urvjpBKZtJNgJ6tLtMQfIg+07CwCsDkf7DST8TOMJxtXH63PO6aT1bXq5I4YN+
l4gVnKSWfTD4CwvrT1o1b9WEPoHNYpfJDJ8PwR1LTaHHKPZomN/JtQBwXKCAZi7NdidCAe9p5zk3
pYsKxOKCD+Ff6lbooshrouT47CKCxueSeLBbWtHxURgXpaYdbeWdkrKNEiqZe7ukGMysVQuW6RG1
nwiIygqyLgzj6qY69N+b/lanmpO0bQq5XINcSDcjYO+GgJo2w3RDN1ZpLtjsJ3tIrsEFyLsDpAI3
//gYnPHtkDV1iIyKm7u91koQTegawZes33/8hfQ7/uzQLkGQvDgG3WiuBFiAXLf7doBj0XjKD3Z5
RKJA21WoBzuRvzdSu8rK1AD95UP3m7QMRtObUXfIqBC8XeTFA4PQwOZnZfi49Rp0AWtsDH+nAkan
vzWCoJSSfHJXGVdikf0pFsnCtoATOieRaBEqhB6w9CvodKnE87BNy0OjI1zMbLJSlWnpmMxqY1bz
i1g4MLHTg3w5OSHZdpDNEPSdNldHSNm9V7ye01H/7r9dIs3gmJq6aoIwLK7IUdKl8ZEqQRcHhA6p
Lhrzb+hbDcEwZGytjRC+SPkpurOlbY9jPosK65MBN3ZwoDUNE3kz7QA/bZfguJ5LRXbXFRgFR+3Q
0xHXIeJWIWgilUeEczigNakenAXBlNlTOssnbpeBIu0nw8znoyUDM5zMHRjHyvu/IzxM3uzCvT4u
MD04tKqn6G5qCh6zKyy+YLF9T5KpZ9HFZEzv8jeYDyn/F0CyenAtaHEMym4TFrEVxb5mQfuUFZgQ
DXZVb7FAkkHWwnU2wEtuq1/7O1cawnBK9f+B19CWNwoz/Xnyr03pxZGPDMiOlVDUb4JCDD7e1+g1
JGpMO96/bcKcqgLyu/SS6LXJncW8BLmUHTYBLXTe+jA4mav9EnoEHdRvogLf8n15P/u+QTl/0iOZ
wwUgWSclp2LH8V2dpZD3ERdtVWKTxlbSgDhjrzqqwTc1RS14pf0Sa+w1H9ZjKOYod01gsVPHvldl
CXAs6L+7/l+aUVwkRiu9BHWvuUEpixzaL5pNwfC4InqrFZJx7xdjFj/+IZx0qudOwoUOLoIAM7Nq
5xQfucCSfYEkyTa1LoatuJq92oMVzXQr9V5GW18Inl82rNSW9nabpvNQ8K5HvSllfTtsSfgAHDW5
1dlUHpQswojxwMqCCA4gOw2W6i+KMIkunNHyYsU8gU9PBKatddFpkoz5DD+zCR04KjnGjLdinVuQ
Muxoxg3+C/lSfWlUAHoZLFJ1qneACGnty25hFHsvjqdXoEv6USe/Togc5kQtAErk62PgftyzkTG5
/0Rlf5QD7JLINqOMRu7Fj63RX4Bg4YNUr63ubO06yrR2fSl4MQoW7UB4SsJIU+vOAGUQrIfrGDrX
nbw3heLVZvMYT8SyK9fEWrEolNDb/MeGO01YdqRf7P3G97SYLr/rFD/bIh0rIAfu4jsH1h+/lu/G
YF85FxdzyS4/T+BQH52F9BihioL9ubRrtDLreAJrEr/CjSoGjhrVUCJSQThKmcR3PXGsG7O94t+/
OqWf9JSp6oMlH2rjibzOOzqoIshqRgNV13RD/h1Y1caxMOgbqeqlZU1UdrEFETG78PNfZRFuWDmV
4qMeoUCHfNhXULg/O+COuHwJHiIrBCnZZTht+iSbfY2iu0KYLuV2VusQjifUmQVdVgC8tpN/Cij9
DVXQJD7CGFDWcYHkwM0IJ+Mo710CfLGHXWC6EaCJVwnJDymx2yVaBEXA+EWW2nyTEVx7HEccW7GK
nRU5uUyk4ALMLLae+TYfQKG7NKU+49AJpxaOryw3TjeDLCzXSvcnODwOXtTkF44weH95D5eBio07
g4Cy2fP7dspZnNbs9WqliLkE7XDq08AO22YASQHYzu37qwzueWTxgMaukMdrH1MS0XlIcWs6vVPt
zG7+24/7THEif7bqWnaRmW2ZNm9p/a0QohgIs699c5SJu0oPEjS6w/eoGrq1Jh/+HZ6bepQtrPaA
StXY2+Xp0XGEgO0rRIcAK2vY/eAqfxkDGHr1wcEHedDTMeX8oTLavJOsh50YT9I2QFXvHB2MWSlv
K04oYgp1i35p0bBudHY0e3UhtdBzD1xeNPALWfkUe2f1QbqwwR9haz/m7R8t9as8mr6yc8yMQlc0
RCxcvA5NVBk4g+UlITFpdpEeDPn6gM8vAgwBKNGtGGUBW+2ub+85h5jZorVgTCSZJFCoGLSUIDjz
OkkjDembEDfPcTWQUtNfk1t3VPNjHR8xKeOKymmWKkRl89j7UAGOKqt/t7RGuUAcTETyO67FSyHv
wM1G8VYH0Kax9K+eyk5i7TKcLwHdf04Vp3BbAcFE/OuXTAVJzAD3FoPXjanc6gGh/8NJScAd6fQV
zvUOx4po/A22VPn4p9YureZ2uQP68XQwM3DTAPBdtkINnnbg0v7qrwV/rF+fUjC49SfxshDNsJNs
7N24ZZZWzNPFiWE3ESFLM5uiX5+zh9f+bxiEsoPXKRHbpC3MeMFGtRKdQQDICcANdinwODz4klr9
MaIk7TIrj2tkE4LIbmyMP0JZKitiD2/M63Kwm04dDYGbm7BUODh+aknGG1QdAUIL5XrtnoNhe6Cn
GjfaFZvwNvm8Lp7onX29/3hNR86s3UnQC99ezzGIM4NSj3LVu1jd/rrnSmSEnzSbLlWR1/3PPSxQ
RP7JxFyN2vJU1QX1UkzbTuze4Xvq4etsNtdcDm8/eoKjuQvmDudMW8KOyBskOIsf2JHjQBdAQ1bP
5zWPvqbpPbcq+J/kTa78h2H/vvjqCdTRZXi4NFbwMnqKB2/EP3UNWYe7I9QHjyoWZDSeXAndqMzG
M0HyeT/UYCu4wu4YoMzmDR6y2F/QPaLjMaai7k/KsRpgYNlSHM8mL4Sk1NWdg+SUJDHcWPenIuNK
UrCYxwzFQVHL+yOui/gskPehocRkEyipS/SzL4tESOFxmhG1rZpPHy3p6C6SV51F4PMoxtWhFzES
WOMaR5m3g4grgM4expowD89+E4i9c0KlQ1/evm/baL0ijWxtNkYwc//izhn7I0+jUr1igUo0Y8hr
7/RB6tx/Vk27FzuGtQLVSi5pREcnUSiUF5cuVNEh/yoZGAO33pQOqRp90+hRrupJLWCuQOcRlJld
TsIZxYOaugX23s9t7KAlPvi/Y+p8YIPavj+5dHJ+HgnxAmZuR6f5ezeioRXhlRPUNzj/KDjLwfPR
4xZVtTQvomiW+yMfLls/Cn9LidktXvIyuBxwc4W0VnebSjWtLhjo9U5SlM5Qqo57yKhaI+zQQfWt
opwtRuU6bzFdAo0+Rj2lvOTwbMOIPu4tB+3iJVgcBcbRuw5eXdOnUCGmIfS55wiX5Rgh8cVrvkTB
4psUfa9ht2eGavndOS4MF41EWLk8qZJNejibVzRzligYHWeS8I9IAAwRY8SZWbFsYe7YwZKT0txz
xwLmMz8pun55278sLtlXYXhBjwihW72aoJtrQM3LuMpdHHoW2nzOi9iFftxqrYJUbF516ufPhSA6
ZGKEvJyBXG1GieS0W6ql6nvpo4Z7OAtfJ4/VD0HZgb24f8YPRv2EYePQg28TVSceWDDbdF5BJzgt
SgBuepaoDKV4MnndjdjGTvG18eh0JsLSXWli4aHwsILc4l2QFqQyZR+Ucd9BeZT1e4shfwPOm4E6
1KtBTOGMxW9FmfqdsCUzUbpddG5nKrhesKD7wy8/fND3xb7he1sp1ZjGyJsnBopwdCWl8gnUjIqi
CBTpGaKeuSXuo/PToLNAL2cgQdXGwdJExh9qH8eZnOS5E6PNdRCBKtc+aoA5eRtilD5eXQJI7SDA
OAsSK1KuD6LP/vSMEj+phMJ/+BERj9cpdhQbnp0s7p/1XMigJ4GdlE2Q8PG5yQnoPpT/NlRG8gpm
oFNeYGatbUVV/cvcvtOiSId3+T9kVPPANxrg3EDwcjJyScnTs1frWKkDfISPeeDeCGBxCYgxG1tq
janGzIalXlE/VsoHFefp/dDU6AsHW+/Vo2clGz09SGceBzcrsaUyvOeHydrDO6NW3dS/RaksNeRz
MUrNqOx/I9CsThEk9HARrKXRgGcZCQCqcudmLxwuDayJcDgfJOqTH89a+0iasikNrazLHTAbMAFN
SfRVqVHA6qZeWfQzcBx5AT/iJytKZg1h6Z9cjOEVvFhg3FvpCDi+9cQNcEQmBp79RgcoAu7iRiqI
y8TvNM2ql9qdRoeLjTS99Cy8boLJ6ytc82FFMqQzJwxpHv9h8FtAiv2CARjWHNrTlsDZSwCUaO4O
Vw+AUyH/DIpWj0/c37Oqdhjjjgxuj//L7UIgVfUxozTkplsMPnuwviKsVLos+OC3tJGY7HHSjUtB
iZDusrfW6QxZ72E6SG7XGg8mGT25RgQdJBaT+HlPIjGilPzGw1akc50IbMcwhuzdG4VokgatTF7A
z1PSK0B56dh9JxhUP9sJ/3aqbEMXJu2v6KOzFVHmTs78RP+JU7N58xrdVpeTYuGsz26GrEjs/WK1
lNm3Qw/SQbnA7ZUHUXYA9qic6GL1OJG+fvmSDrI+fAXlL7nf+E0Mb1JZsrkyDS5XV7zQ1847+mCO
cCya6QoLIJb71o/CyTD4MrVNm7Mh5EdB1P1YjKNCyci+aR/7h84wBGtIbBWdizPPjCYKPaOU4xJ7
rYklURL2zY+LdJLwyo7QB/M2rxSALUBE4/eV2dZxOSrDoMoAvvO7olaDMfdNFwI3xtk7OcylHCLt
w73a3KPWNaDIa0OymDo+CWy1c1ZM+E216fAeuIuaqol0f903hFCRY/5BNg1/frPaN79s+TtoJGYz
2TMFnufKWAmTzsYLCbUSxBurjnOZxhJTpSZcTymhmM9ARqmik4yToohqBM+Y2fHGsqEBi6inkTf1
q+FHKlK6uTfsm9UHfVoQKPrPcOruSZdY5VWBoaLg6C5oLGKfb6d4U04HlzbSbFZKgm7upZvBtUXm
bOXee6ySBw+BfefNSXMbvS9QYRopCaPB+Evqzh/oCm6LADudAGXVh/k/pc7UZHAh+4y7QheLJpRm
mKaS5GxGtB38aRTMkJAn7vKvzcwlnrVY/FZkY7HOEpyE0TMeTtYDvSGAh/WwDzV1vLSAZHcmo2wa
NDzpTjOQSFYqxl4S30Sz9cMhXnZGEiRnXkw0sxMovssrrgWx9WziQZz2thn9N7Ic1xjTAzmoJFcK
RIgvtQWRW+Kva7WbUSvkG6Id678yIx9w4jIsW716DKHojHHsn9rpcE+/Gi97lPuS/I7oSJowWvr4
TacKCBl3aPH6BpspC8l+7UoDek1c6DWgXRdD5EA1F4OOE69VEf/zZNLvxPqyHH4wJyy/v3ba9onu
V5ly1xeUQ4SqAgSU9FQ+3zrB53+QDTp5GL0nXte14/NpO+0U9xczP12Sk8ryaNZj0E3OIHxypYYp
IFGyalVyYylfqKyLqqjxukS1dUFDjJT4JspFrhkx8c7TN666GAZKu14+eSlfUS4Za/2v5aLt81OE
aLJCpTebgz2BASB0O2TRWRxzlkBUix7+QdnVco/eGyfGzAvvKJhZMOuhaRrOOXo6KvOoMF9M3N3V
L++Vetu8AoEDIfM8p0tzkMESm8PPFiPPSR/2linG8OeBgEmLrrQu7K2z8zKclUGXIEPIm0RGyvVI
D71kKuVyZll5GSxY36lEkYFJPaTArpTUyd8MI84Mk/wGXB70puREyamSq2gut2a5eEHPdfHVpoG2
+IsUBzqPJKdtaZgoWM12tKQbcutyJutlC42euKy1m6txe9hsH3wpUq51ux+oqH1KwN8UEtbkz6E0
aOKhHf0Z0AcnuJEX2xq53aPIGk3WeDioLnjE2KiEx2v+eTUXbE5Ol156AGCG5WuPIKeUoBxHSFDE
rN/vXJL0EiYABTGNujqNuLFbUB2r7a/nb1mmeofEF93XVY+kwu5xSAXRIncwFKBXkTgUqdDlyqs2
DmQBULAC/FxgHTNueoXl5dq11BrO7UcNZYH6uVxWi2JfHaIT5hWlaTn/NP6tiEpuffGkmqX+PPvt
h9U5mnNM3T72JOHLonlNE3iittvzf+wkFjgbDljpClZhCS9DJDFHKOhsHk9Xqe8tMDC1fbqgLQdP
PdprEdUqzNwLG6oIni9S8nBUYcEfhIDrTkGfLrVmIW4DVHIyBjZTcCQmGQFMyTch7gOE0LRYYCgX
6PO0Q8laETzilvc3Antx0AxQRP2nhgPp6yW8vEvE68L4bN2+gCPej6K85rNP80rVZdJLzmzsoo+D
ogy7kbdXDd/jbUyua4x2zWLOxFCut5pQFPwJGnst6Uorft0Ht+Ud3KWtFOyx86E1Z/f5xMtsYeSM
YHIxfwuTjCv13CA5xl0LRPdM8tP76QNCtujZkWwyok/u8RGsjkoinxWAcOCrl65b/0e9OKIdhKHT
thIEEI/g1d5bSi9xaOHecCJdih2s9sSA11EVsnrkWPYknZHJWGYMBpa6QHOkLyP8FEQQtm2rgZeQ
unkPlmYwwoa2ujIbMnNtqVXRIR+M4bnNiX/6F50P5ts/Kx4GzgUeZJSlVJW+ANaZIryfYkWhcewj
wcuQBtSmuVrRov4tXd+sluUMDl9IjfNU4koTqtXjaMMshW+4SMsPEImz9PKgoVgsvpzGCHNSbTQI
ZpLM7lmyT3tpD2D2w45VZd5VLnA5CZYZOy1cMknFU1Z1vlsg41Ql5hNzE5hOpk6xtKD6CSWtLq4w
oaOrUygMy9DYJOkEXhADooMW82irrOkG/en+p3aLsoVmOKQuHR5N5YWRCaemYvu/Tckac4ULze5T
ETGYXDFOyB+IamXiOLusau6102ys7GV6cfVEBgpz9uJ+HL2/to0opGgkOUWOLEpAEEmcqPmBkdOK
xhilmZORv+7j8cDYXORafiXiP7h8VPflxbzhzwLB0PCTNDjSGDJYLyxmatfzJTEyMTp7dnmbSwN1
FaVRNwb1pbXkSTbS+1bNKFjK9KXE9/B33r3vfE5P48HXTB7B2YQiEc8IkRd3ZsXcU4f4GgDgZJEp
x9DHj2Oab0e9cSDPapDpZ6bpiZZDitzuOeLU/rhnJEmsGQ86ptomrgBESUu0nOo0ECiHzeO16CxI
wY/7Twt3Biu+gQ2Z9/GbHjX9VL84TEYpX6ciMLu5FvJZSOuGxoAQtPvfwXTnxIPzm8DkVfmoICw8
KSOnlGk2gBnz5meTeR8OtC1RAFa/dvZAUmxjeCmcgSL2icqPvdEKb2UDRAof2QzM3CtE3jyxkfgk
/OqvOORLQRFlXDVXOHqzF03Wp3ILJd2zqRjpaQigJ6coiHfh5+R9hqXUeMtFRWhdAsz8oMvUp7of
S2NUWLYbDcFW8CzYplT+2eM8OMKAHaqjIJKwfSaJRzLqYbZP3KhR9HXNiY5hCnJqHSUoad7iG3vE
3inIuc3lS0aimQj9vgOgIYq7TSJ4AG/0UapWENj6V7ieyBSOlfdBG/BEo/K/YxKfIvg9zKfL+URo
9njLcf0hv/8P/gbPC8+4MYcJ/Bnw68T5Zp+5VLVx7lqofK4F1MUavWt6RaZ7iNqSmQB+OJolsbtl
elk9QqJE7l6LuF694mYYgp7ouaKRMrTfB/jtbMM3B7x4S8oxe3WB5uojDP/jPkZIvmgmnsF6l+mh
4MC7kFjv4qsrYTeUX2KqHVQihTHPWskmJI1VHMAtQTbbFcxZtb2gg9o+Tk+v9BKsHzNVmTbFRIyE
RRG3J71hG2/Vh0vY4QIkOpZ2KP+ey/tWbksUFDi6T7nF7GcdcI/IayCuC+XvFjptvtB1BH73avly
Zgbh5hW9AKFfaIc0YWbUyrGAabgeSGuNz7rygciaL/pXCKr5TGh3Y3Gkwilca44S/yx2eBmodAPa
93FOzZXW/UbUI7cxiFKZBGKrrbeYwcaYIJMr4ljGICwJ+k3QYwM+gRgqEJg+aulrvaq+512cRhQ4
V8js1m/9UiueQJMMF3bxDP8/Auwc+4xOkOtHIFJ91+HTztRRiGvYO0KM0M9nN3yPX0rXM24lJ3WT
Yqwlg8S+R6xyG0kqXg+GnV2Mfip7IwSw8z03oOTHtxVs4Vi338wPBFgj+nSxj6biDSBH4RiDFdOd
ehcXWEyX9PDFVLxZqq9DnVyhG5IMWmHbepPpHuafAhSX2NKw519W0ZMJA7hlOvC1HK8XXvPzGERx
H+yOg7IfJdah06LD3n2Xkoky5lM0jdHNrJ4RBA4X2DFZ9e+xlJuQJl/rJZNMu1kupjHXNcZ6o8th
euLknXy4nvC6HsWlPzDyibepI5k4m/eiduDbTjrd1eAH8aN9o9bUv9xRyzUIghFC4kGCimw9n6ne
8yK2QZr5bnLNBTkaCQq/3ZDHooMIt7jGz7ZX+Kq2LjgNrmF3UM6sc/a1RFGMdP5Ly0cgY7oMyINK
OxU/LMSu2u42KzSEiPT7n79Zo3+nUeQPm2402+GlamQ0OLiGCMFuGwd325esdpHzpFZIg0oIyK6Q
6Tmozq9nGtZc7RrPFzshp1w2KaI8rX8dlXMeucG7RRWLdmAZwbwep18Q1A5l4P3GrzkfR7fcsnqr
uBmjFAsK1QL8mMJ4fooi0FVWhU1QMKE3iL9dgED1/oEixEWqsLBYxwofNkMMi++AHkWKo9+Bltx0
erUWcfzWbT9aGFolZNadSLrl9Of8mK0ARfOJjb7uFfwqarhkEmjtFltrpJh/tasRD5nxmfS/BrDg
EpdGeqJf93cVUYTXg8gw0aoBhz+/TC97FMim3laz0ndgKzlQbcq4r6GV7LoIrfBHULum5VkmSHpV
ZBBK1BNKrHehBrvjAMc2Q+BtbKDN01DTOAor3HVEATDc8SZV/YBzDFXLUke0gOeS747JL9Nsy6Tl
nlHf2ZveCgKYS93Aq2Q7gms/8shnLAFeodmrjAgjTl568VSzjl3lOuf5vjUPn2THKE8dP1Jdw5ip
XfbciT3zZFtep440bTmxO3df9hvh1hBZObOonJPq4VXRTqJXaWr5xaax7omE1D80XV8CJSa7YTE/
cR1TL5hV+nJ9V4gL2mwHgoaGCkMxo1Sq2qYTLb+aG1k1P4t4MPGhbAg9Y3ffxdSNqYzMDVfilUz8
DdArT/kSr1lEF9R1LNl73y/oaPS5YGutpWu9fmyV6ycP8NNFXpP23/ZapdX97cMDFsuBjNjqmf4I
237TYS7+ibIja2gK1QIbBfXOQAl05PRLIo/v4yAaC9MbBAZ/DEVBKp+qGZ9u8gTFChCqyZFRDrUe
vflsYk9rEahaGPfXT3AnKo8H9xe1ggRK19TNTNVREe+tQtyKTBm0SVjoc9vuSqSytcMX2gaAtn5r
V7d3sxDtkpwVuzmbHI766PQWDC7p2u8ws7j1TYlzmuuhYQvLOJC6//wB9INtrid1c0RDeFfqdITK
THwsUczNWeVT1oiQ/nt93C+DXSpsCZSZLOUHCq2UfGZDmNHL5dJrka7/Zd9o0Uyf5RvPoYzpmtf/
n8LR8ooM/714qakWCfvsacn6lXGIvqr9qC1WWlpUi8WyOefoe9sUdM7q+s42xPnYlV1EYp9W8j1Q
XclN5TXAZCauWybpkAPbwgLs2SC0FBCt3ZjO2exLAqP4VVCCvoH4Vhtj/NflQGjGxdC0W8m5hC1M
K6Yx54YoYK6zralQKnm/w0CMnCiSr7lF/kS8BmbSehln1WzLNqgFWAhDVcJHE8HrdLnsB36Q8DQt
WNb+THRXgi0dpJL41Fg95pEqN/JBGlBM9sYTfdo8CzYGHeGU/B3EFWrE+18Ui2UChv0HgeGQnOkX
loqIpgqZepazHmuIeDp1QWoogYZ3DByp1Eg050ezLoOKK2w6IYJUB3Tc0ZpahTiK6bLNRfttaInQ
f7n7mbx/i2kfIsbgAPMbKoUu7oL559bw4q5Pl/h18jyCBsxJ9d1VdSCoF9nRJz8NBZse9+TzVvPj
59WJ4vvX+3al1Ki2jxinXUSNyqatQl4h1SYkx8/GTdcWddFZCVx8biS6s/YHJ7tMv2Q42FKTADan
wmzhYUUWh9xLNMxQnS9Uz3MS3WvCC+wJTsUrlDuRw0xIPKrWmbD3PdDLtgG1APigJ/xKCZSa7KwH
ufAvtxoEfuVzSgbqIplgCyrDT5Sz5dTbyyEfuGWaLXcpTmEWSKCipeQT85XHoBxOE6pcXOZ7eKjz
aGTvSPPv2hyzBU5a9BmIbi6nXPvxptdfxZDjUbLLpwfz8mjdB975QYN3HNwBt3bEGumSclJ1ihvC
m+iaeMDCKNgUo9cyNFLweQEplxVu3M273/vGTX9WaGWP44H+lJFNdOOxSqMnZvpD0uZjVe5tpr7C
JxVE0GhupFVdFs009LjDVaKVUxx/gV1YJHjQpF9fyrI/hKU/+XC9LcddhqhRl7rBQ3yaZi0aXJOw
NEXZfkYpLFRuA9QhRTz/HxQLcS3FfjOer1cmGhpa7jjUd9lYJ7fJvgMpj8zxVzRdl6C5z6Mk/Qkm
bVJWp/Edpvy/pLsCMCjgt4XBdv7ZEXXB/6PPIMJR5Dh7iekeSEYzhz4Woag/wcVm67iRW812DUhY
P3vZ/H4Crou6+OX/VoZw3R21Kq/LozlHs0dRHVjeDUEzf85LRpCN3ZQ6Z1jsMcN7QRlj+Bytjdvg
l8Rf0HiSUoVDt2N5e+HHMj01gLM99Sb4baYi1QNslQ6z+mKJQLugS89pakpjVLVgV3zCHfdvcHm8
tnxbHSTr6oA7qRyzlbHPGxENKDLDNol2Akm+BtYSQIoqWSiX4qthADPt78D5Rr+TCKTR9kEiCzrg
8d3tOFtPDWNOFLRbM2E0ctW9jFfyPOcNmOUn9x15Tz0LJY0NgONYe9Ci+tGHHKx9TfeGm5yLoSMb
MYbVoDRyplMvzF/lh0ioofdU1a6mSzITNyadIUy5hwlLPxP5e+ngSLHN0XySLCC8DGEYC838waCW
X6H3jj1oJjZfRNDRXPN/rETk4o9/IwW7MKKO/cJhGR71B1pXiI1U7yq4W9ivONIwznFPuYgsR7Nc
E7fMuFPitT9xHpmhTaSvRxZtFPMySiKDAVATf9x+U7tsNRQW6DrdmkzkZqu+vOYC2ygN+pgHBtU/
nNfi/KbTV2flQRc8xYjMWQkAlwS8jhfwwjwooiNvZ3ozhZpwbwNBILiHcR4Wm5G2WW7bw8UOkdpZ
P2tmjLb4c2W8h8o0fL8ETUKb9aeBDOghxEFvlDp3MZVPiYXKJ9A9duM8UIVkh6ITdIfGeksqONbQ
utD0bzdcmqYP0ZS6esnzqWsidOwtnqDfcl8b9dzNaEeMxbu2glXcm5BJ/2FioYfP3eh7fq+reEMN
m3EIx6giZoFHhn1dp9AJACtpTw0Rt6JqqFtsqyh2CofIRc7wTy8BEW8FiR2f98Kl76EhxpSAKoeq
9ITipuYFRlYFew/YD4tf3Zn9GxO8AX/Fua05e+GcJuJQxsPqRn5YmAK3N3HJcxwk4P6nWZ8iOYnJ
6LQQAHNpuGRrUbiLTLK9iQPU6C7TBXGmU1p7lrAZHtlGxw4zD7BtLwHEmzLlaEdzCW0D0+pSoGlg
IrQ5joX4dlJUYMgvK3JQttNfn/2KiGMb8u0LqEP6gOTe9snOIMIYLGQMsJrQhvZvd9hCs18zrzDF
doMHysrv1bC5dvQ7ekXsE1GJJ5PJPVzZdufuiP81jAOYtanvqjmKnnoTWhS2rVGHPXJV6AS5Oyq5
vDbaP8R1JG4X1Jx+PCTtc2xoMiqlV77Qra+EdsIuMfhJNuSKtM4V+n+p4gEjOZyM4oi55oESCAid
WDQ7Na+5P0Z/SPZwGAJ7dVoNDezFCc2Yv6Su2hZySycrMFDEaR6dCyr5NeP2YaNnSf0uWI0UrYIT
ZoRieuZtsjtnIz008AYpBwcuXjfMKVYTeUu4199r6lXIrAG1/C4XhICHQ91E8CatrJwb4PdzyVFz
5laEFjMrglqGSIZouYgBh2uuG9m8xFEzxhG0oYzr270B//TeYIbt5WsdKzogEwniKGuZoVXEMQh3
4SDxwKuSbe9BceRn0FnZZhKzs0GwTQ69dJI+DLCQlnJR1cCAk9Ipc/ADnmPYvImWUPFlqSIleksu
fFENP2PhjP8ExlxAy/mpoHj3yEOmQOG54UPXq4NsVgwdEBky1aJVfG9EaNMwLnmnLT09R/6GJ3tQ
fq0r5LW6pmTO68uKo7jtDbTQpXOo+LiHXbwy5jjm3WDKVtfv1b8aY1MvthPriHgPXTBTqq3AXlRQ
xS+4y7snJWpThWtJjUILMcRGWjCeV46krwyJWx16Yh7MPb3O810BRLu7pimyvqiOHpbNxVP9l5C9
rO+uFwrU5dbmJDkMNDYO0pBF8yYhWgvv/zJqod7DJufZ48nLyDjO9Ns8WC1xd3tsPEAzNe21HTPR
6nJ/Jc5KzzMI38/C9qmDgz63w1E+ialF6boHckPND4VSoRWZJaKlc6HUFZsBRdFO1XjLa/7HrS1g
FiPqcbO13bS/YSiweGcmOa8WGc5Q4c1MXs6dJFLukdEcn9S/oIsF/iqZz5A3XSzcIfsPnJ0/1O57
gBTf+n2SFWaUHmipFsuDIHYwIlPGmSNYYveNiSHg1dgjmZZ5neTi+Lh55fPFYuUKkJ46GWqhmGU9
nh0j+hv5O5wgP4+mpmMVGe0B6xnBZCJymt0Sg6s/PA3pO3b7CwZn0bPIWaVv8uLRZUmGYqiIr7pT
bOpFos1fyB1O8RL7Sfup0dRHI3hym0bkWbcUMdqwmtSVcfN3FlGfBWS+QMK34NzP0OBxPgB5tk75
WEdbo4I/vle8D73SKKAtX6FEc21OVG0IytnWmxk7cmsztbQ9F4Kg7BWqeEKjmBZwg3brf78OzA5d
S3SKmP1ZZWUPTQ7cJ4wDqtX/oq3kuV7kV+uJwiPt0bVR5CwRSe8k1mTf6OIl6uTq6iwzkZTeB+T3
6PQmmscPZpAFny/b7bAMwSX69jVh0VcuH1ISGOWsWTCb3T1slKEKcp/s3znJ1JwQUr/uK+Qnu2ba
fW0hsOLdgwsrgcyxX4vf6ldW5151t1wVGDu1hid1VsIGjyonE9oX4TvRdFVKvONF+BjaWc/oyNaA
DOBKjS64QiUKrh/l0IGMIrOW0/O7Sh9GDFua/b5VDo7zWB3w/YjHrYFQ22NfWaOdoLPshU1qpxo0
ySl6DnJAX33sGSe1UjJ4mzS8Vd0lSVPLb1qKoPbD/fpdd3xUz6Wo3JG/Iu2eBt1iLDs3N+7TGvXA
dptk7ntFQRK2AsooO+5lv28xeoLdrfpFzHvnZgVjHH2Fekr1RgYMb5Zh47ZpP97gU1i5caSVuVUo
qWHrvimNMQJu7/GrdKoyt/vP79mDtBG8MT+XIzjeKwInP26NV7mS9ky0v86ctMT7bAIDGlBJQU/J
OBWMpVAqgtmGEuoQRRGAdbjYfx/blpmYwd/AjFNAFq8orf5fH7z4Jnv7aRMoU8Y3VzdgMxoehh4k
tHMJZGCyxyCsYAeRlozoiU3kMDrWS2zxU4KVMmeLNDec5GZ6GbOxr9VWCpZf12+m82e8shdMNAO6
uWD36wAUUEIJQdhFoFr9xdxG0UKIdiDD6815OafpIT4+F9LNsf4wewRQoEK/rILM8iL81I+5l/5a
EaEiBJsQi3aUC1Xv45K6yWOhzhwb/9xJgNJW2Pf4Xyds9a3cR95DYdYx7BihzXR5Ea2Ve1MRoQ1N
enNiEEgzHnebsMC4PH5kdGmwmwJO6IAO24jqhZ437j3nNUqqkpLtXJpUD0c4XS63dkZu7v6Is8xa
HrJV6jd4pzwNtE3+2RAjHfe9ZSMzsKIMF/zvGWj7V2zXH+/vvqsqUswl53jDAq0FS02HoFNj7FqG
hwLj3U34pg+ystVrgLAn93WP6T5CxFzs781awvn+7Y4+f82rlPuHEaf53ZOSmGzP45KEphs4wg2+
nrLDVLEascX9Uv/Ibi2DdWJ0/2XtNgKpW2HMYvYCLYzKryUvvn1W29pbkDcJYu2ObPATO2o0Pt7J
zfBrGiMcADgd7eZS01BcW9LeY6DWYkaT7Kejyk0AT1WXJokx5xnYRmyPAdbWamdalrtMv5/lzVIJ
0EgT24KGfyqy5J+HiKAb5xiiREpVscVXP0/kDTJpF93zpTmrHnkXgVqdPZG437/Rm04nc1ltGP1s
9SEKZj/wS6+EJdRfscycG6Nw5v5QqDBG99Sd3k7EZn2mc+GKgWgE8MjkIs1u3Azc8GxwxlchUR3X
6aS12+H5hPfin+EuhGxgrrMDbpABYpuEFjFfS5B7+aMwafCXED7Esa0U+1CR2cLNmuiorjFCSaPP
Hx/nJK1twNWClL31RpXOolb68JeDFe1iXChJkkSlHsgixsohqBm1QJEusESEm6SNE0vAcMsJ5Pck
fpV+L7f1oVuYOLUmOigMi9XsStWUh2gszdBZHc9551EsiDMlw0mqgarr8h0RGXsU91rc0HuapQpP
oVSMti2hNSjh77VFSOQYBnckKJnpRWBZp+BiGZZGaX1yeqIMmo8p7MUmjSND0Lv3Mo91BWpojq4Q
Ick3KGhiRvz/VuT/CIeF/WBHP6n3jh2P3+GHyV12HKNko2gqJFf5zZz6t4eu0iDKKRJvQufjf8w/
KgK7WErpKeG0mNaeEDMkPcotHed1+8SmjxZd0Y84iBIt8UgR5F9cqGZFYrl85pRq2FYTiQ3T50m7
CVKP8qNC/XIBpqeKhu7p+xGGtkM3i/Nlyk9dOm6LfQO46U7uGRU/WDmmPg7KXmluTfGlua7hSXQB
Wm9wEcAyTbMyFt8QX0Cl4bvYAgqM8n17LupmYV58PyAKLmrswcmtS5Jd2xPoldhZ4t/PcsD04sfq
lS7cbvHlwRwzt1SnDD8xEgMCCrUTu8mQnlOnzaeGUi/5JGsxAr5xe61vKSIPdVoVU8fP55YOrPIu
Qqm1LqQLxsVtsoj/10wxN+VB4pZipcY4TGVZoA2xCekxk86dzdjEFV6quW2pQMjq0LJnnewpkOFM
B7L5xOt2obgMV3Aqy0qXGF2r2X4yWiagZelW52nRbn9Zvqp18nuBJjLntlmUxA6KzqZz5POHpU9v
sx8NWFXUQFSIv98HY6xGTtSbyIgDPTACI1bUX0ynp8VZuDlHCe3mK9lQJBY06sr3tTO0AOVnUGVl
8OWeeUbnHy3BHTeRqsvqmNaudiK1JkkfOPbmetbNlTDchofJ8AIQDEzUBfrf5ati3hBMQsojxM7M
PJ2ISKozs7nrZxP4m4fZU1c5v01qw2H3cIPpvFSFJhZKoScIxQFjUdDLoAgR2Ct1+pu8C/laVzSH
eiwpcwOjPc8W7STFiWeroEgPVGiWgS7Q8WBSp0ulJ4K+Vb//0rh0Y87ew/lPofOnqkIuT4+JFp06
dUAfR0Cv75M3bbgllFu22pBp819cMWZXeogtTLwbimIb9yJMTBGJd5lwfC6wCn1f/9Xw2I4XGiK2
Q5zR15zIHT5YJ324Oyrq4dwEgu5VHMcWWM9iy0eMClQRgMvHc0nc9kcS5VkZhiNm2OFlJumJt9bi
BeQVPecz1LzXqkVO6ZXIbcwLmErGoQaWNNaR0jtfVYtKmebWi+WHwNnjV21tlS6M+1TcikxJbbFt
p0IGTC/R47SnMkKHjY5enNQDNyrtmqsYnHM2vS5JTio7HatbjJWPd5kRUUfzNL7MTj98I0I778Fl
SOdl1SoikaazDJGwaLEtgPwypkKBYuSaMQfjH7iAWtR35yXkiEZKbOu/C2ut6y4yruvEB1MVWjg7
qOoC2DxMLmJOCbGLVwIyxByNmqIRcr+F3qREg/OSaFC6UZbnGnzHwg7jf776NIWJB8p8sio+ZURt
jFOgg4AUUaHCq+QR3tnmwpLiYZo3vzyuypA/clBEvcRkEhnxLlmYwrjjSO5wwGqN5RoOyDtuZdko
ZUmpfI3/UL8Sp/jm84I6byYg6K1hvQoB63gLHS/3wKfRCCeTCHJ8AG5cC9ox5O26mbS1JQtntsn7
qumCk2OQItf4uyI11O1X1RkRMK4bI9Rbgsr9RGZqBG39zE2l4S4eIRplqQSwThZE2ImL6wwwcC1C
ZlJGE1RMcUF5w3p9YG7vM3wq0XzCGyWn1Z/dreah8cmCO9JtB+KTm4Szn0q3ln2Mwc9P3qQZ4/EJ
rTGbW2mF6ixef9QDbtxxxk8MNCWgPUB84KBA8x2hdCVcO6ovi/FmsGigZ5oiDHG+rhZ/yhHivw1J
a0l1l/EfTSSM06u0CX3idSYYCup2eEIo685Yfw840KpO+wzCXrhENowJGzELHKMzX7anlo3kLgYy
AAiXBvUuEHAoEGQCHRTx+BwOWY55CwsCHNjyApAtGt0BkQ4NmK8FOGy8vtRcdC6UITgiDo3pYR5L
j/2uyVAxFet3zyg5NO4GRDapEA8iW3Qh/k+gMWRIYqZoxvyd0+oLXT5N7syjByV4LuWiDfKy/Zt6
//yozVOEj/anRRsevLrkSyKsuOuWswkBCTPADD7o1myxOvyOpgHu/Rt+4pDZbgD7/GyB9On342xN
11/VwANobXV6PGkCVfZulWnwJ1/92LBXarWaYqzilDk4m49+TXRxIpB3gkJiLhVZhUXLYpU4bo4k
5GbepShfNAAC8pV1Ml76PUnqzq66+q1Kpq4zLMFw4oT64BfumfUMLTiunzFr50fk/0TCNHfeDSRa
cOc3x7EQskTEPL4fwr8LhxrdLdr1qcsKua/QA4gaQGvQSlCD4q4kKEOPouaT6+QNPHn6EPnjf75f
YRVVLAbEeFcqBvHfDqEH2O5xLXlM6JZHmZrTEs+BUQDxv7xJJVjDyRGaDuZy3dgYVhuESvdOzJTt
/dpj2NBDxRHPKayeiR+61NvTikilSyonwtQRI8dfGT9uDAr4qFRFkwGa5rCP5PICyFAAPnNskPbY
LKqMLlaSQDkpIGiBW/D+Lsug1/MrUACQHbado2lPFYSx//JCcI5R6FP3PDS4SOzoaKQQvVI/hqnW
n6frdeDz+oAh+Txu17DCGOTD0JJkUoxGZMZ2OvX+/sWO4cfw0qnmDNE1BdiQQTWAmcAdLpeGdS7d
bu3qZcuFBWsUZWZutpdQGOfg2GoyCEJOKYXRVVneMo/NWPh1tFBlXLD1pNc1V8xd6ZHb6COk3QY4
XnLka7ELJFm5ghN59JOTX6s+yFFVdN4BAwacK4+SH5v5kalYBC32ntZAbgsdZRVvgTgdpoeLyPe4
SUI9x8PXxVwOToqjmvRIIKry8sb1G+8yxhzgiv10DUTNZUNRlOtj+CHM/V6XuhMudfVWoHFRYM/1
j1NCYg7hCEWQ6RkUDUrHvY0DmLv+7zj97Q+QSmPpvVFnbe9oDQP5W87RkFcpG6W/+MZmhs25YRjK
Da6ux6xLz03BBYw5qKk+Mc8jxjlmQsTmxZ+OvkITxb5xYfKioCrPR2g3q+mXQJMh+2/0PEhHoZ20
BP+W6lWvd4ub5oFFTKgIUryNDuIquObEBfjDTeXIJEcoKy/K0gdTkBXa4WfBwl+DQ9z5vBDhdtZb
zDUXm/FYm7Ee8J5sRD24QkNVefX4PjUeB7UzIG7cqzmUWNdzN0XlYtfv8NWHxBKAXlaCHSKeg0Wv
CFTigcosJ7knSS7JsRXMSRwmfLyQEkXutCXZfWUqZNkIo0+SphbROhgu15vcSPZzCFooPItKAOnM
1ycLmn5ZGxbuhNkQS6RFj3eyTpXB7BVAfXIY+0KceaBRqO4iVlO65TY2J0bdHmgT7DogikilHYm5
0VtOA+GipeATWDxBnocCtJueXsQBqSLf8vJ73Q1E+Y7/1mA/RUU6SN9s6F0WnZm+ibZ1c0UY8R5i
1mzBrpn6DMkE0LyHEihyei8IZXEhuNVF5wCkyg5sajkr71LlRkBNvPmgqbZjYgzMeMdocg5OX3sZ
HRXcytQnIZb82k2F3FjjDPCJLrbJeZTCztORmpOBUUa8eLLiAnmST0hHb3rvNNZYW+LAbS1u8yAk
HenKeQ4Yn9A8fNwJks63jkmJUwHQpG07nSreyy4gSJeMFC6FyQCw5JFIefU1ycUCz1lQLHgEYYIm
A5GQKRRbmzn5bEeUwMSaNb+jFKl/U+6I3Yk2XMWb6Y6yHR/XwpSDPg1qNK0iZt0nr7nqpSU1Pouu
1MIubtpgHr70zBtfOqK+O0DdTcMlq7dOeH5N++PoujQUTXH56Ru32PnpqiTN7kMw61j3AEj3nMG7
XppBT2yvHQYIFKV6urMhpjRZP0GbnVFhIlGQzCsIQm+yIS3msW8FeKDwqLxIdilXZSXMxz5K0RL3
V8lI3aKlvW045/Tkh9Fh/BSHSME3T+5hK0/1/NNfxtR8+GvLnXlKcgBI9nX7rCqLm0h8VOtXcLas
yzJTDPZOyeMQvEQdwzDUI58xPfrBIzqdXoyTpLEYASd/mxLwATThX21IWT1LjLlo6wwoAwYZNCSh
MxnKJZ+HnQN/Kvzd1WGQckYNdc+gzZ61Obd0JJgXbMK1ebGLgPDCkldPaCdBIBjWt/5RKX77XgIf
8BIub4w1YB2vnMOgioA4q1MRGBc5wtHkPZm4awsQqZ9ru9nGtrYD9byItfT4nUmpMkVvD5PMtGKj
8qpmOtEAUKUa8br5aWnX+6FOEAdkvNqQoNyN42OKJIUlLjgAbS6VAPXuwTPJu/YyiaeREWPJ54Vf
gKfCUUteTvp3YxIIODqKBJKX5FAO9CiYXWBTkEtGaRkWnZkL/jIdG3gnAC9bZ+dnqZXVddHDLea/
ROelLydXJffVERJn7q69cjrmzXdcJuPwEkuduL2Mvim/1ywKragi6QaJxu1mwf7gw4uNeUczNg3E
v3mHlqU8A0lXtcdYMpmTsXkVIZs6q9QNq8XtRKxWJquImr75Iovx0KvAsf1G4IZZPX7o0n6dRe+V
f0kkpgddyYrM0wtEVBn59TES+d0tg+z5KgDlP/yW1Hwufz6hCy32cekQqRJWVMYQfF2A7kONgVtt
qYANz7jVoC4EMlST9SgIk2/UBr3jyxHiieMuAfmXHVgKGQBCSTuVINDte0vQzqjUZdCZ1CUsByIS
DjBITOJpAD7dSfonruBkhOV3MxUuxBaVyGPQ/jT+4imVNl0bdeu07swrcGqHGvUtobltaMzOyIuJ
GrDjrTDAhXmWfC7wkBDMmTk7LAWTDAHlT+JPc5GVYNymlTuP2BZFM2c5mV5Wf96dctNQQohQmG+0
39S37hHG+2jgD+ryS7FguKlJ+WFcIh7X8dcf3EwTG+jv5tn/A8pSEsbj33go/XSzaVXo0+89q57e
SQpknGUJUcXCkBp9lSgnnuxGVnAFzwM217+7EKepcPThFkI2lCpSoObWUAQpwr6+DBx3SqJK4F5B
sL3RfoDuAUmDI/h8zVGYSYCAxLG1eSYtTXOk9c0y1eWiEiI46zDn4X5Mpgnk/YlQ58yjiyWOfyP/
GtL1VOZwX/51n7wMcI2gwPMGrDu6LKXJfld9MmiMBsZUj9lY7N6YR/zJ3oTUm9BXGpJpvbm1to+n
Wb6fMb+jABdOr+4787SQDrNqL8TBayYuNj739HYHpWeNwrBQVq724XB71a1+MSvHqkEWoHJspzuQ
3J5ABr/T87HPiLHmLVSRxq4YGq2XlVPSxJjSgUAq9O8YVc2oTrc+imL3Wxx8Fzr3VitSupgh7bor
qTYfi9GQUQjkYxDbQqkFutxSSL0CiJoseErV2dsRWPQjF+IIYAwwHpFOH0hDYxL0LJSemYOhbrPu
7dncalmycYVn3X8++7CEb9NbS1fBcZWRRRWVFtLXdzyiq+zSjl8gnIB+9w1jUj0Wy2AuB2CLBCd0
uo0PZlqZC+nLSfqqVf/uLyxVnPzQ0LnPrP68ABo00RstLDJqgh7oR5+fDTrJiS9O07ljgz4ulWnt
UdbcTwrAjKufstBVNFk3BH6zknj9PDq0MuKBmSkCOcnjbaOkRk/7Mrj5ibx2uEwcmDCFpiH8Owxy
k8ScBrTIgxj74A8jbwBacAgR5Yxx5t53RJKqHZ+KKTtkV3Y/QiVm5NNk8BqaGfN/nXHje4HdGc7s
PgdrvoTV8k2XqjbQS3oUNf58So8f4OdYk+GnavKvJxytMQtoHRQlOZ2AHkhlQCfx6dZJ0HUclsR+
/pnnEe9N1Qcy03EHzbqE8zaiK7O+KUrRDjv2a2R/ArBVob8/+Sn4R6Vmn/MfMi4marnK0NE32qdQ
xumt1ZdiUW8ucAhccXiJuxbfioKiQ8loaVn3eKW8M+JLVhPuCHtm1P/tE2gNz1K0+F9dzBHnMvnr
j4LE1MXtmeKyBklLGwJ2arwoBEkmHNd57Zf4RzUqJYD54DzAbG/tqopc2/eD+qkOUzxmSAihXvgr
k5h/TOFZ+jH/wH6ofl76X6q/jhwW61fljsvmEqii8GmuOABJdeLEOF9tL3TJZsIWfoeHASc36OCf
7Y4H+WkrQFovC9Y9o2vCnnYJ79KJd5J9DolwLITb7Nq5+oGlOCVu/YxZd1FgPY7Akao3Fcn/beLl
f0UzybMavA01202Y9W7+0SAXGYBCd5Owes3QvFOOJ+Njv9sms3BjJj8bYWp7MDefgSTyFLuBczjv
DGtghEdwbm6cYYYUNWcxroFFHiGYv47UkQkDdTSJptA6G8TJJHbQigAttQ5N96WDb+oNQcvQpnxD
J6gLXJ++mJUK/h4lb6d9ZWwYFLWkIU6E5rh+0m2ZWgIPzE8DTy4zpFhSo97DbGuOXKMOXijXSGea
33n5gaQbLJzAkRuBui9BYpHnuDu/IQu2PqS8BCrOZ3pR7Rc3VnuUkhHFxOl0PR3R5QbDqPoFxkQg
4+kekG7X78wYYUv26PhZ6NnNC/7dFgCI8cB5qQyZHBEWQodoa4C/M8BJGDoIK4BE+xWN+u04klje
TxFqFKM2JDKKsQX6XikDeZnLYxHcRUW6UlB5j1p8JKZNvq+ZX+ReItOvTs2CQXLYM863AFTzqikU
DIXi/euxJ7D8HYCuAx5CWQLM8zn/dPzqS3KFuwzaJgsrqQ6OJdyPZpFMroQU3axGNmtbHxR4u82N
kAtJQ04r1iL9kmqEgBv/pTS4ZIoYDZWiRbMsoZTwlhXBcK7BAFQ1+B44kWTJK/+uPsDbHaEQSlq+
wC9/MZG9HE1nFsYMOvlohM1BP9JYHXBDhJ4CzZrhtQS9mnSOuf/eq3qXnMSxdCVLoudSRk2Vlfu3
SlK3yxgap5VkyEjY5SpHhHhqjIqEvKcstEBP+dEYIWNhxjBasQZH6CFMQbuWAa0M3QG6dKGbWLL5
ePF1O5TThQ3bOwjbHeYghgD1RtCPcfvwVuqOd8ERM8JSWR9potw+EVf9xkKWGHE/5uP4gcuZxNe/
cZoWU5STiePOx3cmkSs4xBgFCtPQmt+Z5M6jc8SCSJU5c9+/y76R/Woyt5k6+Cbq9FO8+cIQ26nk
ckVTq0iZsuFBDrcK3b8H1PJvVguKoCxOr/hhoaQ2EWg7lFMLYlD9OWHPNrGoBRsdeiOIcE0LrcKa
c4FE5Vb93ZKiDfOcFQwqTmoL9Zt63wgLAedCCfbgAOxxra2YuyewPnyHII5DSfBbWi+NecnyMsBG
VoZNNxikIR6XVsDx8WP6k5Jps8ogLXFH2lhkcjAh0mnJxVcgSRBkp/Cf5FxkeiSj7AjUQESTnuHU
N4cxM/1LmuVbjSz3RtQ+FDttOlvqoRzWjvKtEpz1pD37yrnoxP5WvKznAMrnuGfyOIXhw9wlzVX/
L9IbW32if+y1dfQU6nvfBwy+NZ7azS1djEjcRJq/sfYz2/ohV2TzbXpkltFfpp06eBRXKogZf+DU
duzTrfxB68XsYKnt2w9eh0wCdbqU1vls520E3u036TPRgrObuuPSFJdu+3OmgFXGArpqY8Rik7l5
e5r/R+5/ROXTSHOyzCV2FfItiDuzuhYhgs3zpPnbxJVg2MYAlvgn9gGBzibXAGEPAbB0eJmv5jFW
1XPKHSw52sdpr4UYXVO0eBaslo+aWLF3R60ym0bJ+61CYmVFdRFY3L98pieTg1jUA9WUlDNiGsKW
yXVRbGdISkwPJM3sRE8L2VeUU3eAasPKJKYEsLjdU0jxXcdoAxvP+i+Id9Zvv4cvAh24+Dlg0Dz8
V5Pe38ce/WGBIL9waC5EQKLaTM9/zHOex5YxoqzCZMK4ofTDWR650vGwyCLAWPZoR3hAL3HGW08O
HG9ljFhqpK0AJmaJIiIpbtuYHFb2qyg0bU6AikEQADlrUvyvg0AGBRG9kjcV7MMem7mwpagSsbGY
WfLLWDgc2xMkDF+6nUQOFDObT2CVJ4eAUHkH5H263f0iqLMlsv+OQY9HjBBTde5mtMr31QNqYbD6
Focvsi+BzbVtqT1XE/pYBk2fyPhcFkfnG7a2pyE0cnlG0rbN28Zv5fydaxPrO81ZLp1cPoVjiYic
pvo1YhSxNFflJRm+xDj8kYOxoaHZS3U+nYUpIncq5gx0D5jMgMSoCC7HkzMsUpnxeyswcvMXCQtn
l4J5F94PliH1c6rpK94Dn+idxP0asz5v+0s9VFc2uffIJztDgyqLxrUw1W1gvuJ/C0eRAcT2cOLO
xZmHLlQfSXIQSzqOOAw16RHKagcG2HFoIfoTE9t9TjgEFwMA3Q+4B5Em8+G8dCmg2Ykugfs9kYRn
luWMG6Wihz5mJyWnJ7Hb6D+TIFQEjmZ5hZrVtrL873f3vDZRZeXdSBQjIq9Z9SA35NMzNfHkVXif
qllE/H+LwCnm1+/+S7/KaqswRth6qyEi6+t7MqH52WCz0U5LPZ4eebMI78L2fpxlagrFKYjlWROD
LPLxHfyM452NtK2f0Q6nmLd0IxAH7veUr/qLokDFBIr3psG0PlGR2vG/9iXDWBwu96cUa/HIDSUd
RYrHYvGb7qvpsk+w2XT70HgPIly9EadfnBM7V3g8DzG6Ee7zAuYH6wOwjUPw/o6oOhx+UBhkGYoe
aaMMsQn7IT5tPUTEkjjGVKcoPBzF2OKcnsjiETj1XtWuJXcqv2SybpBV6rD0hH99+q4uV+jEEr01
pNxSqkTuTyi4Qq2DXXxrYQw7MhEUMWLtHBsm5/HuA8XXlt97sfME23dkZ9GP2tCRl5CLWJrgPFry
d6gyiuKv9qnyqJaMDk/WwdODtK08cUQNCZd/kTNFL6MwjkZPmdi5f/woCKTSfdzMp86D1AHnODTv
aheH0ZZK7A8cOkD7QOCyfKHL/YArLnrDTEKHFCK0mkuUlxMIXOqOuJjgBF0e8CJM5LT74rg9JEJG
wMQonJ98t5Y5POr9b4XsUOFmRnJbcW4s2FR3lYjp2oS55sS2XFkMJ8Jn2T2/Orj8ck7B9l6S3U6c
IN4/EIQ8E+jRT3Ytkm6OxDH+lrn3QDxmmFh1OOq5n+bIgad5Wa0BeYEcaQ5e0IyX0joJFoR/GOpi
C3PKi9i5ccknf/skDd8MVvaNWVBstbN6rvFKMq11E4Vm+lpKIAYyIUsKSH0pgRwt8Lu2Savzhg+D
2WrWlcOqL70CpRcLFhdziNp7RTzAge3Ty5k3ZPPxedPyaS+Csuw/DXKZZ7KrIy6mEHdrb8LV4m+Q
q5o8ZTgO5Q1RBptcvcNrFK7U7xuBsJXD4CQ84txYRNDIIRXAVoXRHC/YsfT2O+dlGf4wEAtkbeGt
Fzc0AviMnq5Ey3kWg7ozS5k7yqgG+WXrxIdNGzZ7OaG5a0R4vo2Ox0Ggir7pCrF6RjGF3vZWG4fs
yY2/2biVIAoa0XUO4mNJKynzYPMLoJqUh8tEYh6b084rlDsFZqt125EIF1gt1mqf03IUBm4OADoc
TSxGs2Ykujdja6ilrMNwguauPfrNKvGqBy6a52cWFf2YC+rY01sOC+4jy83EP8QDgVFY1EVxcmbJ
4xQLEqTKhZKWJuSPX9C6HZ69hFkiHrnLEoKIhXYSGIA1IRVBhrGcKYYmd/FM3eOF7Sc8Eic3IA6+
k2ixnaTsRmi2SeM7fS/Uj4XSqDDrRW1ed5xqUObZOxz7906pn1qI6AaK3LDZTJDF7HNR03gUt6lI
9/wecLPYLNtaAag5ALRKEZe24/BIvVFis+4lNyXnFjsUTHodEdaQEV5Io+j8R3H/5GUoogbXqPB1
p31PBeo8xIxlvROFU1ghYSGMmIF5TM4Tc8N7clNKUu5XGxKIqII4q2xqBICoNTqKw4xuIdwpSM49
V5tFnPMPTcHqqpH7TCPF2aObVs6hMTJLjh6QhipQtoV9QMPko7vrC+6EMJaQVrOzFXDy8f+CHllV
zhcjjKTlX4N4CEI6e5OF1Nn8bj5pTuXRrUu/SD0tN4Tn8NNEStKBGN7G7qF/XZSP9lbSKoq4DaCK
jl2d+Kq5ic1KXv/t0dCp/Qgo5mOkoDh6tLQCGXm2gc6jFKtglmADAUFCm6hfb44+WUcCvdaBbMJq
DJfUBK10AU1MShBXF5xV3HCeT3t+kuJNiWYx4v6fIUTUGbpiFoMTRPGpLHyqvEqanJRU5nmo1Et0
QX1lhqxkA9ztIxsIv4rE0DLhdPn32cE0KCTWQP875zbCvPm6xvbcA6zgJos839pTR1BxpzBsDuFh
cq5A8ivbizKMUuFBHL2uZvasw6MaS+pkzLcwzh2NGkpq0DBhv4/zkueCd0tXdadwYiCsBbA9u6kL
PWTn12i2cNxFQaTRlT8GJpIC62r2TmX0uFWrtHT7YxhzKDJVdSqcbOwznmJX/f6DlmLWwkIhvxfx
DeJw7TnnvfOJJEKi6xfv02yYsJsSNZxiJ3YC11zfnhVTi7CAac7UFrvZ2fbqjEfZdnitC4BnMoCJ
3TpXfIVVEcWnfX3WxgSmsKeNGD4EsgeX3BMXtu7xD45Q06ekG4t0MxiYNqHr8YnV3z0hX74HVAdz
ZVz+CFPysxqrrhNFgfKwmKyCY9hB3PKYuAAtMB25jnntIpZJuOSj+tnsOVyEnbybhUlAO7H+L+8V
3dfIJwaTWzEJFSHfFjR4M2Yvzn42hhrcoIsxcpd/Arbg7JuqqeK9djEC5cHa2v32torRayI3LpYu
iJUtcDSFq84KasMXoK99/H+pzfvG398G/QG+Kh9q2PUJXANE7OicnTC+K/lhpz+/FDkY4xGLlXEj
Glz+srJeORzJo0tWVQy6arqNhOtyz37FpCkevMcTLnjmKKMyHnkk2Y10Bxy9WLxa8suor97qt0hL
h/7WlGDFTJfdquzhDoFwnn5KMBcv07VWdrP5hPkpIL4V89Mh7YXCE8xkFEVBWIwsPoXrF5KJyOr+
fp0hOqZj7Gl8rO16if7fe6oCcLfoKra5I3Bth23o9B5RAfUfqjhvIahO4loizoFQF6dPCf8SWdvX
4J00tW0LjRZqPsnIgmF/w+5OkZ5ad2toefEz5VqUEyfFusmTk2zbt7aptNXjXIHi4Q1Zy0p+UdTi
70LoDlbGl95y+eAfgaMfXQNCX4oJ8h+t1zItLZQUZebUdFy2sD83/VL8y5CkdtEsgp3D1ysYah3R
6nrnsg3mDV2XlaruRmO1CmzPMSqZsfpXnsRE3VLVBKQrn7V1OaG7oUAdEEnXQXGiixwym2rkKpBG
N2rFdPuFwYrz0C6y5FyX8Ln8uiTfHMO8cKZA3siNZsq3LRaC9sl84H8M4x2hbzk1Kz/Wb7QJbvoq
xk5m9z5HZZN7Z/EhKbZHGL9PRSWv7G3xw+0uaKfD5HNtMFPE2+Ci2qv0ExxQMwQ9uvSI62wOky8L
W7i1xsb9SjjaIhBAsmAQD1Sg/dBkQaGjFfnqLBJZW3uZo9e2Vdvdk1Zn7iKz1dH3ITPhKUnVCqA2
8ymFSga0rBgHI4XK4mXoOGFoWds72KtvnWW5YK9gihHDcDyN3Ye73Hy+34TeNF461Or2NJGJ7+Mf
MNAU1p+ggkWN7/2byub2uGVwct6W5JCuaFD0iHiWh88qM5uDCJPt/sVvfiMCoBOup9fuLR64w03C
U/AeJ3vN88tPFdRxHU/AI4a9H6axaG58zeODuVLs3QLIouodEjM0+UuBDnnnRgbDkOhze2Kodtzg
zLYUA+hDc/7ez719ZE60HyRqi7NyVqvcuLAlG553wP45GIYFFXhlsZCfaIOwuZRLztq24nv554RS
gpXI+Oa1WYNu9mvuShwb32jb3qCOlc3NhAAeoMrcuHxg/7QuOm/tzHX6g+BTBVvfheP0RIS4vmBA
rzhHc0BggQy3NWMFA8svFVfANQckyRNjxOCghR1K+iRhFQ+L3YcMyk8ntECBqNpMaNR7ST8NuFTN
PvI3bwmc9zhKC7Vh5340pTPEBCf2Bv/u9DNCfXakwqZK/cvmTGus5XtE8q8NraTwtn3w8kKDBAYn
+euWvUfcy8fiF7Zm05ZuJqM/lBW71apEv7TDUsL9CIFtJh7NVUMXWsxq2Fp3Lf2srTzAlAa4Wj9l
LqSS/hdfG9wX1bjHT5ieBplmM69SdaMhPBUDd436iSJo3HD1hbFawnFoi/m8LQ0wkd3e6apRUAS8
+Wko9SehR9K4YK2HZKsEcYyJvtz5Lklvbj7xrTpSC2u+B812LY9Ln0Ga6P9xwszDcsQHW+bdcchb
71nT5W4brjxeyagTin0LYIwAOH4UHjaA1yDP0JU6lXXXN/64Nr4E+WDhAmPp7J1kSVTRDVT199qm
5tP/b+HlqDDywc1bCLG47mCAcuCkWLKM8/qb6BtFegQennLF/kVCpuWKyLY2PZkQsdykoWN2MTpF
aogUz0vxrOWXQj8oz3JyHm+O7YuBmv2iUi8r19A5feYKNhUcxXOq9w++Zq8esrilJ59VmWPSsL1N
Qi6X2NZi6hRHXw4xHdwa6gLsh9T2P/juoJ80WixncLm8D9NVIfhRmdSY4n29SIggg5IsTkPuprxB
6+KI+kin4m5Po+VdxWJ2DzSyUwWaACEgsGu3QcHwnqfGUp997Ahm1oP3QVmfLA/veZY1Tz8AAj5x
355O7wQc00XgL/Y5HAQasr22M8Yb60/IpuPC7dfYYEV8sdlrrdocXG2VZsdykrhG/anc8inMDWY2
PXk9YUAn45DvIuCu4g56fVA4Dxopak8N8yLqvgVlAKe3zLhsA3pSw1hT7RGYGWw/hqUtDUMZGS15
YRuYMjBX87WHNi3PPm1UGNjh1QsY+8MRpN0h4NU+gABEEObmRgs/rAnBVWrMD+c7Feig3yIfnmML
7TF0NhqKF1b3khr1VbzQNp75NDPgb+Fh4RTaDUJAtZU19Xoeh8KyaZHeetpwLtN6aAt4rtebgESk
o0d48xykpVrKfmuMbUHgoV4M/MMnEdCbYgr9Gv7qmAjyusckICN1B4xpmYOHPfX3vzcEqdYT2j2G
POXmS8+YVlKUrKx7PnkPl9RlAvWSoXntCcyPfknUvD+yTsgT0TZlvEda+Fs3cf2Lv7BWapArfA+g
1cGMJIBnoll90hmJNBSYQomL18/yEPyxky4ALICpE1cQOT23jrMlelNooJchDShC5mG566TzCZQ8
sXpqD1AESmfz/5HC0E+WiO63AGiaw+VukQm62lLZDf2YthsC6bxi6RcUbVEIfHgcEWM58gw3cfJ2
N5FnL9fQOK7MS3r6yj2E1ejcxKwusnBvEDvBrcjVpvuC6hSHLmy/unXQrRlnGb4Dic0AqShfjZDG
xXfdv6kuDcpLcO8s66LmiQ6AC/UD2d/gY8VYD+Nf/XbqVXMvZtvpdiYK7PnEJKOMC4XQstZ+FFod
v+2ttyXLrzfZ9M+FQvxR4gRPNVUtJ0XfH54E2ZTWy/Wpr43MqU884a0SwjUqKGIvJlXbdLwQ+Vwq
zBWk8+l+ZxAswu/FHrmr9Ewb6nktFKguD7Fy2ne0RhV63QPH2G4SviNQgoTQY43SyBQmIvxbMEo0
rpgaup6QbDB3it+PE4HY1rsA6LPDDxl3g+8DINRT/k/lwEtnkeg+KxrAEE25KLpeixl6jOROfsdI
e2kPGD0TKcvJoHUHuA3gLiTxYPFIbpxTC8B5dqDsEQtut48eDjeUxJESxv1jt7vwb6LKrIcY1VDh
HFtvaMWf5TsTwMnFZui26YTABlQLaz2fjLjEB9edi5M7NKV5/bVWvkTdSRTYTVdK8xeyeza44ZSQ
ZMx6kepCtpBl642IDzBbZB0s/EmCCJucahuTaPl2o9GIumlDaYakrrBq9j1XG3rzP0TSYaHWJ53s
t3Q1reaUmnRIRBZ5bVOMwTXpijHxQ4qCRJtUfyK12dSb6A66V9awtvyeoJNvwbEXCGg2ecxDAaKk
/PPH9JGrYIsWQIuUqFATAWdVcjmhsDRU8OXVE+r98qtSKmmO9970fCYvEimDeRL2SGn/zoWIdA/1
o/Ol7pn0N6ywWDHqf6K8EOT7RI0GVMK3SnD7nAfCHS5MfqGSIppNDcQMX3KYzm7snQP4HoLZ+vqP
pRyGrVwdgYZByshB81vbjtHIoZMOaYqRN50R6fdKo5kxnTiVORRxo+PhGLv603p9IjKzgVN7gYfh
caWwUN1R5rVQ6EsFrzfbsJ9qOkgt42x9Un8IwMm5ljO3wjWju0JQ5Epu5gRienK+RIRFgxu+lA0Z
XOWMjw9zQ5SUvwvc2QA+wnkLAs10j3DyINPedkz3xXZUo/eQJWDj/dntxIb8HZrPStwdNkE+6WYj
lHCToBCq/jArVPCqPYDWv9bdo8JwAUW1r0WJAxmPfo4CfGToTY90kXxWFTZuggFrzVvs/Z11MOq3
vybJ0auooXDAJpSFuvfExZbLTQCOUSZj4gf9+yIUMYv9mPKe/BAqVIncOPJqa5KKg1jsrZx03IV3
NCh3FJNrtI8XE9OfcRKKhsEDuNDZ1yqnBc+6v8VLzYyoUP57D70oytkz0hJoOmTzHOLYwTkGMGK2
gqjllzVzBRTMJDA+xZpqx4KSZ+zRmKmXfpqCGy4sCWzFK7RZyTihR5gRUM1kHBkwyeJAZJErGw/u
cr40m5Mf+XGvVELIl6/5L9b/jIDO6AlyXnEAk0rGkonQHdA8vgsFBTJkQY5SX3QaMbogLDFdqenz
/S+43X9lopthJfW9VyEdgz/2zhO7sI+oi/DdTLErJ+uNA/jLGedqchCXkZ9k0Eff4Op746lfy77D
vH6zavWnPvznSxorZueJ863yclWdpskcTNCqlC9LtVTz4oqGMo6nZHPxeDWm/3oY8DAMIYlgc+Mg
vmVuTwwXvf6LrT8sTbIsrHaZqdIAmCIfj/8oC2vzna1Iy7EhLFMbek3xD2xGtOruKS5UKc4tBFXZ
tJXgqs1c3dl8C/UH8k26HWD0w6yxeDp/8+bJnUQvdOUKKs2sL2Hqs/L6J31uFQRF1cK3PhqpXsSp
7dTcifOgCO1R+MdHEZoOnlzpu7aSN2+nVZCgmSfNdgl3chRsmfI49dhi7fdg+7cnBYPH8TKz1Qd7
fyCqSG5aCrmihpTeM5w7Zq23gM3EZ0L6mPdGBc+3u7ziBqDZTsbHgSKv8bpg4sOSQVjswxhOSxcd
BobsiiTjAPE3+Qwu2QJ9bKNbAPHkMrdOpNShr/NA4bbNUfAKoxCreHmTDdi/RBt1PgS3hzJNcDNT
H093+HIygqSrygGq1AaQcy+6kY6RkWmO4fwSgjLvhj1PhwcmYaLtyfE1KcNxG9ycP5Kqs0GFCzOa
W1aBcdCaaCKcPQwxZc8xa1+9jSJ6tFEXBhiR7wlfAXmgviKq3cDhJQ7CmxTNY9LqSxPbB7NctU6f
Q1fah2AJf+0AJ2nD3rVmyC9Db2jEq5gn8If0VMQsL+HM1ZKpe5aj3HxzA7gi1tF8S9RKFm3zK05n
vNmv0XL+LVtx7iVhWv3Ll1K/r+rm30z0T3bwj9HZ3BweV0KGceqTyWZgb3BvSyPJPC3i3YLtBNhh
m6CV0DkusNWVLzzXONI7u9HJGYXiIZ2Pn/+l4sPg2gYft2GmeDWmh7k/ig178h1DAJ5UIJExRPDO
BJZN8/FVx0DR6rThnsr5tadDzYcdqVw9Cesfv/+b0r3R50p0/DO9ZthmfWzj80syDvLlLQBkj4qm
3CtIzIb3Zs/w75n6xqt6QD9NEgvrS46oppmaRw2mJQ2G/vctR8Xc83IgKe9OupkqIdn3Zr95x4Mh
JwnaiUxSERs1b8I2GnULCoX9yqFxJ4AmFt969/dOoJEeu5IMoae+fef4ndJ7LmU6yczNv/gYL57W
bFHxqqTKHHtCxPK5UKevcbwJLGePa7eII8noLB+LqsnguSkLkfVBmhRHOQ+ZyBJvR5J/OQHGveBt
WiIS2viNWvdlT1ii4gJLWRmFao7TPxS6UjDkwQSCRREb7B3nPs6mg44YeknmllA/scUvDwcCossp
/8BuWzXufYTM45JnXJk+X19YDvZ1P4l8mT0OVdxcTbKMN+0ysR1XRBsLhKIflm2ue2iuUOFDsIeX
RynvzobXmsXyLAA3qp0MlWa7RCnc2tsLZk6mQvluJZguOxkcEUuE0PTEPD6a3d24lrQ79w+q1aIu
xYy6zNEXLbbWLe01cQX7FvqfGQJdbt7Xp+HJqwBzx8mv5Qb0l06dgZRNaF8c89aDbqTOg8+/80E0
H+Iss0GNAnxcCxsowpFShpAI84WAk3fdlurvSXyfLMoYHR46LMHof0uSp/uOt8MIH3NCB4V/quc1
tzaFRBCb43KvYWg/XlTjVNGARGMzopNqFkIbNttiLt36PjK0lvVpARdSzJaChSppEvsHa3ECb/4U
AMJ4aFAONs+BdvOaHWkF7S1ZXu/9E/aiTt7tz2mIf7me4Ddh/hm2Va5+jYZL7Ns+G7jVT1ro8ya/
Zj7mj8di6RCOTcDX8ATnchEza/lkG3jGoqFN1JBN+1ANiTn8l6bUd6hPBVJ087bccWyy3NDM30EC
6iseP+d3hMDGe72AO1/iWemXPAV5ss6IjPQZcOnTMFYWfVfXKFm9o8DT4PpTmZf0/Nri/MTQyUx/
9eSz4tJFu/8Af6iaoCudhvMFtREi5Syp5DIKqGCyj/sGOuWkTUrcibU9N3fyTfgMIybSxFx4UPdf
VC2c1iI/SKjxW6O0yvBQBYOAjQ13iHjHJLrWKIm/zVurA0622gB/2rHzvLbfBik4ZmbiNdhBsb1O
uKKt4zvi48WgR0ATqsPv+qoG3RWq8moOtjWNDn8bN6q/ngjxkgiFdW34/CV/kL4P1sq/pb31uBcp
3sTFa/OxFsyR6JLed7iR7TjhLEDjpQkH/F8pI0xWlAVBM//429Qw3FeYcMcpsMnDQhsH6Mdpd2gJ
Mvi6Un0TiQjRDe5Y8fnSoxOnLlXOJ5Z3fFFLVcn6tTq1ieCxH+hq13PJhIdqKHdY684+r0yCJQmZ
Xh6HksK47TzeU3K4aKq6rhIra/OR7FVdp5VVuW0EepTgtbpJOSo0aCx1+kGLsaA6K9reDHSXlLqM
tBwKL2qehBrZGVXVjIdlJu0GHiJ3C6RnRtfo7X037uPXhtoCXgg/r++h0WSk0EmuJvJ9r79DotEp
9zUj3adjbZ+3NnNf5AeCR/eCizgqlY5AErQfua48mRsn2LfYWTcVVS+SvGNCKJ6XpCT4/xSdTJiR
z8gqJpSrWEvmQcqWHaydhTTC5VuoKcfARy2wEv6AC8E6RfAkHhzzFm1TdyWJBXMcZwjcTLdMYbnM
h4l3Z9VEUplWIQdeGyn9+3EzGcNJhI2DzpCWyRdXEiJdxNjDHMvoEvsKH6kLhI804Xd/V8LL4ROy
9O6lUZxZTD7Gkdsu4INk+u8QdWTnHn/TxYOSyTGhVNu869r93cOBV6deTqEOSNe2Sp0JOyUFZr8U
/mm3btVP/jLx5/tASKCGNHU8l3YY6HT5IoAR8XXbxo8Eh3kdMeKdBmm4qBL0c8U3xQuwdnoXa/tn
HgIQk6pfKHMCYOPrHtPqABzmK/l9Adp+QbliezWe6K01p5Mf8FIhKTq75JQCuNGoG12XpMhhMY3w
zJJYWWqWZQbWSSEAnwNl3sghIlDXP205cMfVDlQXP9zSlfqPT98dxaBF8hj8U182ZNXYgqvSDLop
MxBUCTJV8HHVRQnm95aiScGZGKtKWLzQ/1rHuo6p62yjXGkBZ1JgKKXVXGfQR/5pbHk/TLvnECMS
FV/I8UYk/1ATBbpwYxWziKl0snBkLxmnJht/aYZJZYQmjGQaP3taFtim4Gu0l4lYcjQ9jA65du97
bpWPfzI10ffoptaaEX4ai+ZOeUQwMNVv35G++ZEr3ZzRc3oXKLfViBjHPhR75vslS4vqTVlU2D52
uK2mySJpjqNpRocWVWfovdJ0Rd6/c7i2MogNiO4kjR1wL+k2PYWCw8V4v/6DhdvUlZvJlm9tgYQa
rC2IxNxSFxTdd8BZh80hSAp2SNBrGYwGGwVOHgAsqhTizyvIBucyiU4TI0dTb/tqrtF2BFquJVxd
LjHb0om0HHg4wANEnKTVoqJZXwRPJhPzIlLYNsqLd2o3gOvZ+zC+yZFzLZCMR4k5iQssdHmBUyCV
+4gi3YdKAbzoNeayrL6XUCUXVgvD5dfn5bLlzkH4Kg9Q/B/kPf8GtlEhtyE75WhnxzcPqCvobJG+
a7rNjoBqOnekGDR8iPt211rWCzTQ3Wu5OUKR/bXufKkXzof+8jF3lQiQjHHu3jiPH8Cm7DQnk+gs
uZ9vCDxGitGOnfkE6NOKrIDdxYQ2Ape9TxCyiRzsZy4by0PEpa29SKeIxpe4v9Y7ApwcEsAX7yId
6l/sGF24bsyVbWihxpMdu4Fq5SN9m+2zxE/NDKkODCFiATWPC9/ueUrfaXzJC1/aDRvOtJyqcruZ
mJqkXJAziuH4gWtc69B0YnIH1XjtLGf3yyJzlW1t7Gyus7jOVPNgHsItk+yMW7EUgIVfjfrapaSh
y/IsBT8cLw0yAJ2JzS2QjOpFHLO/OgZ9I008KpKyqVqfEOnkjjfZsINfUc0pzsfPVvbLyuYmiCsJ
dMNiiBecB8Bht+ibYvv6sZDyBFUuI/ULmFMuXrzAe1seSbIk1qa5n4aPGMZj5W74c2AoAyfpoHnh
kKwtnxPe7IDnO3YsqUN757SQuQcawdhXjAqlEOmMCl0QOhoFgNN76vRKn2nmwal9A+Jy83hZSmRC
AN1+/hNtLHv6HLFdgU3DeEBNAO4BeungPdfUlb6uVnM3cVWdd9UJjaZlW7Z2RXmSDxJlSurzRKOe
dakTYS1LYGK1ZuQQXRymdoXosx0G7YTqTyAs2AP4FvfOAg4RxZ1et0l5iFZI9ik+Pxio7gSevJzZ
OLWoK6f6uNGvbkAFt/UGoc16jcw6wUqRZm23i1/SiEogEatu7NQbgkNGBeDQh1K4nhr+BMXAGrrF
fuWB7XAWnJRB9WUPmNTeDd6wfU4BLrQAce6dvDSMZCfSzFZ6Y2CCGqXqFDUgIbooFoftdYE9XjrC
hir8fj1++VOW3hXErbOB4Kx2aeOMfnUOZu9kb6Xfg9YmyrN9KYpN6gNA6xcxtT87Tcc9robMqRuo
PJXJz9WS5oGa7NwQd1G+Sz7JVx5ICfkYOXSsJQGlH2WVZbeQI+3KCVnE5I7YXhNXwhWD4EiRWMFG
JxBGH+YbS/mUCFNPZaBQYTpKaTb06JRJiWPGHaPcTR6r847Ws70WTgfxBDgZohXyQulVHaLeLoQk
RvrDDaG4LPzY0kBfgH5q8Pv4GvHYDEWmok7ENZzD8H8beKqiYPDRjoOghfMrEJ9cZrtB+nDqvWE9
/muffIqvuP4goJyJ1nD0ENtAGd2U74mA4DCRM7Krow3eIOQC+WWOYKUd/B935rljlwbVBEIY13Yt
MqmJ4kh92JmlRTT0TuIv2vz2pce2Ny8rS/BTJQ70bNmw139nIs+tg311gUoyXtKjsOmXkvty+Nl7
IxzI2WQQ1VRBW0BIv9m54DY+abHIQQxAG8MlUFR9k5iPArjMF4Vhr9meqEASmJtL+yvl7VOS4L8y
KBNS7hchdfp6uzcCaMpvSqeDDWaOjUauoMOt+0I0zfrOzNq0ogNpw1fQft11q1v6+F1XPGubxNYW
Jvynt6iMbbqRWYxz7k+pBUrgymH+J4b2NINKt5yuOYFUTfMQEwaTumLhAKziplOHHhTXhPLvJee7
3zvEj+6uhWaXPfwz/3Th6LnAsIey1y7npELdhhHPsdoJ1CZjZvMv5PJmIgsokFJBMl8qfWH7iUX9
onPlOQuw/l7pwTmpROFxtTMXW/2Py+vl0skTYXptcjbGX/3oLLNltzlUBmY4X8rUw3V/yhRqkGb4
/7NciEZuynXjWY9QBIgMwce/3mF5oBuXXG1n7X7Q73PgV957vJ90iQj1FD3/gsU8g8ievF+cRf+7
avnsmXIxo616zNa5q/5pe+uLE2qMXUZ+cbfYv8uzKhwUqfd2wnpflLuRM1fKo7rxG/erASoEJRA1
ruPZ8VCTMDaRj4GXRaOfy8ESVp5ooxJlPOv5Y0c29vjGACEK7DxJd12ZliZZ6L5diICYrgYRw+7l
BgQxzwDP6DUU1K1nNPV7HGItxcWTYoLmfimc0YM9fT4ZnLcScZKuwhWDDh8eIdke0dSZkwi0ZJ0E
l3EGooMhOdJU9qBnM4llowXe3U+y33LgJ34D6WNM1jXF4fwywU6TyzfamhPbHHDAAAIfSQxeyISZ
osM6br2IHdMUtqebeQIfq7+F4OPzrOlXpAOnBncqMxH89EyNo4EdfC5c61mUEzqW70z7OxSESvGS
INesSLAJGDDQ3lgCI/0hJf3PbC7ex8gkmmxsvR4kHu+fmzzIjWRc+tpFp3ec66SmwgmbQv2j8xpb
2V9+PmZ9g119AizlwaMnriUr4ooTAk0e5KrB/RNIP0PjppxU/MjDH39CpDt7UdItc3kHUSImt8O6
ld94ekArWzCnMDLtNhBk43c8ga91zEqaGUAROJ8FFM6g3q2U68FhSO6C3B4yE6Xkk0dC2k3HgWC6
PMGFbvNiVZ9MCmXb9Qf91tlpWNdMVwUX+Agq1KV75OtyzW99L/Vab4rXT+NcQ3Eac2/ThKYSWM4p
7o89ihj4KVy7yeYyhiw3H67d/+89RAf/5Z2C7Aepe1FXyjGd1+CtnquCFSZ8T8FzZLOem/6Ju9Dk
TrTfDL7b/owDIXjZXlJ1L4tATMKabRWKKW/vH75tT6V/8M3+fy6hkoyzVzpGlbRuo9Eoy4wZrMlk
KZ7zYlyVgVJgWec94VBln+PuaogeRR9EUYXbDMI8LmI8Pnp7xnXvVcE8ry6ZdDSSdo9MEQvDqKu9
XcHBP70U9OxMC+H+xOMFwLQQB7BKRiMoOgu3jULXYnvzPQtH7l1K1+kWle2lRkGtTHWTecHeVJsk
OvvmbDw5nOFsHzo3kZ+Y2FBcrcKvYq+kdD6ij8LCAX3AeSd24bmjyOUv7q8k9zmdqm8XovDccZpU
mZG3EaiLrZHBA0TBgeUgTUIDpWyobC8WjgPC/MZjurslVVOg9mtxghDf99H4eJVynnasbhjZQlH0
PoLU0PI8/Sf7SOz5GTyV+vJrGWv2LmsVSvN0QFFvgESw1Kjg3RcQhkfw22hgN+WXH2zfkCjn2bGu
P/dd50tPrRH13M/gk3rhQWytKPp0Cd6Af+uYVmeUbLZZpFMVno5Mi0BCWFrEuxtf1zMArU8s+r4B
dbElFCv+RP96uRKjgKw4MxtkrrMyPtFq/SrTKxL2tjIIjVwLXKk54MKiaAktCfXKV2yaZW+cwg97
/ixfzHrbg5hraTxhjPs1MqoJrTV838O2VrHKZTtkH1C6gLpP+aA1BI/9JuK4xSwlZEWSY80WAZWF
PutLxsVs+yYrNc1uj5eApJuGE+LznoQG9bUg7TkRl0iu1ClSQXg14qxohBiRDc5XcaKtND8H1Dtl
4lUrQLMGJnOODU9mF2Duvvk5RqDsBwfHkFqbl+YeqP3PSe/WCYdZhR5wF+wmQAUpGxdcIlkDNNbQ
YWdEHZZY/qIFigTqYguvaej620Lj1D7VzZeoOQD8BurysdX0GIsmatYVSWgo5G41RkX3dA4rJk9Y
CKl8A9ofkYWl/XoC3ZZmOoO7ynucE6VGkXa7jrVdc+WjhX8NZpuameoripPRpY9GTeGf6krdXKP1
egCO4t+SvNF1irKJyjdIYJybD5c6wywN49mP0zr2TX1oTthuGbANt1hsaPEy8WfyQO05pycNikF/
glUYDzYt14Y2MS/2tiKyK6uaH047lsOylHSC/g1595vJN0pOAcyq7fUdP2pjcD838HUvualemOf2
/AUZHR6dABQfxMTbjvyyqtFGdp+4N+1/BJ3whl0OFhQonWqBHsVOgCQdpGAgprWWAR9QnXlqEgHW
CsaIdTe7IA7SnWKbQlbj0plVNYPM6UHA+UOxY8IVbkq2YvsVejvUrhMM3KsumBJoB8o/+bzTwiWb
iHPHL2bamqdV5ETOocz0A5Sne4cmicvYu0BMh8YRm8WPSePEcdEoaoySYs4J9PsXGabkB/VhxbuH
jijrn47zIlyRA9l7NuVN6iUgimxYCDDzIt+V1jS9ztiZYZ6k+94ynJa2dyjdPEbmSLq5iO8yiFAD
QWXvcp23Ysi0v6bKFyXXmqvpH5qMTWX7Jygy426Y9TazyXGA+mdp3NHzdyolWtVrqQdrFKtD1WLY
vOvS9hmiyOXYlGeW6naKo8EeL1oBwT8RjjYZKkgxaE98xNax4xm7dVdDFnyAt8rvVCnvpRF7TMQ7
NmwPRB69qHyo7eLT8TS+S4xjQLolFKcw1Sp6NdmCALEbKS6rRfGnD2le4hmlDjMjKnbYkG/hwXs/
MSqAzZ5+M9ZYTsuzHIjydydrP2IcoINwseeEz0hRngPMK6J0EoiCG1SLWusx/tNeYaths+MAnI4a
v1rQdDCriiDvpCGh78E/W76nq3TdBMWT1ZCXdsLHk/HlUI8KDKQ+GX57DPl1VJGEJscYVFa40vBn
sBxLr9QId1WC6+JOrCCTXzPs38ysbPr+HbPhqe55edJexpwU2e0MxXXHF3A6mEtYzOr1sCIRiegG
iYzEDEk9MnX4ihDQI7tkHzVQ+SApjEvtNVQI04PjTBnnGpSDjlTaA8Sae9KWx8dX6m2iRqWrQH9L
5raZvuzXkDp6vXpwGMrXefhS4qfHdLm9KMqpWuOdzYlV0honm6cAL9DuuqkB/m+YlA29xleXrNrm
xdNtLCgkByDQff0hNZ3K06IdSgBHOpipNvx4Q32g13ysK4rp058VGxwPe0rEqLYpQLavV8CmuU+L
yMExyziG2FnFpNiMHeS/37O/r2pFBo3CCqhlLFmO8Xm947DMY5EtfqBPhZMT/iO4jzUCUIT4R3AI
pe5vZEG2tCZxs3QTJk0kidyv8/Wj4d7hZnqwnh0tqQ0pOrtHypBhj591BnXNPg01yvwd4S75GlwQ
z+gGMjZiRlLk+UWi1jzr5s6qjC4LY5IYjxNhJulZgH9nbrVOw7LpDdyQHXzoZdYNGUdnqq3du0A5
rd0iejESFmxEeA0q1RrIdcpBX+OfB2R7QkpdTOOnzP5V0P9iBJEIjRbNjCN7gkuH1u3i+Fyjztrn
Br87gnscQTtVsavEuSKhCfupjF/YZctcyeb5P00FaP+s9lycoCDgmM2ji8OHlU7a0vl+zMPe6TXD
JX0odaA1bicQSkH3zOy6onkQett+HbQkPmkAkf12fgVdr2r++IxRPNk7tbDBaJ3brSVfu/XcHlWm
nW9P/jOwBKdzhJ4kMqbIw9eY0Cf6kXJ9g4s2XRjKRwDG397wPapFd3rI1aS015ep78yDJgJxyx3a
NnhULmfnMb8iwscAYi/TU6mp6uIxR0y7U47iRfWmE0KkMhGYAG48+dr3Qg0ji9AZPQY2hTkz3yN6
1Opz9LNFBk8Gv4d089SPa0Q7tvM3ItgGN8ijAKJMKGJeEnOcyRmWHXor+zQdv5BfeStZ53Q9Vqsm
kTTMZwvUvk+Sm2B6A2fKBx0OPDB+THW+pel5bVrgrEVphmyxiWvJfAAjkdYNhM2ws9ZGrcw/gPyE
pvxAwHD2hV9zjB9Pko/AiqG5wMZffCfBJ89LTlo8O+3XE1SlIteAK5LjGC+kfKcTcbUyjQTOKclS
6oLPTcjyrdeTMF95/6Joeh4nji0NuviGsZG0mEXA6A7vuN7nMljQs7srPiR21LRmlnRXxX1chpEI
vOKgEt8HYgSFR4sAxt3ZjxAzRqApQ6cQTHnzf6hDwR+U6lFoHPubpNMK4TID4I+McZHoi/8m3nRH
KP8xngGntd7eu462m40Xe46gSq9GAsW4ZSeATljT4TLp/B5NCDP19BneJlTSmDU3APB2artiOPmu
Q132G3M07XYpdPBg/BhtHCs8CnKWEgdCEtuBs1x4eAj1+Oo3KzxjaeOfxoVlJ1ZxpvU+NQGieNFd
m464ArRZyKWkHjTqVGI7MJ7vPf8X5NSAb25ySlDQLW90XzA2TD8gP09ewQ6/E6ETKODEC4JybN4M
jkw9FdRfPpxWiig5qiHt/UxwB6jVz03VZT0G+MMLuL6ggymwZJVnxmxEBydv6TW4IiiXE8ofIDTB
17sSdfy0LBbVRqn0n1szl48h4RF4ZJ5OvJhaX95DzRFD9grg+z5Zr28GexQmkVJVAqaYgFBQdUdH
M7JxIzgnwlkNuzGHRfD0MqUwDTzdxGxiUe6S5de3UNU9D5y0RhB/vJ25Ur6REsdlHDeoxCf5O4rV
aASMYjpY/Q9bNfs9fBrw19b6dAmbi1ptGHJg+TY+oaEz6uT++Je3xfX2kTqqGG/9AOnjQqC0jqfN
3AV4DogjZsp6245F5r17C2GmthTKapThlnA44cbZTspoCAtLEjiwO6mHb7AxGU+47hltM4yImsnB
iH97BeXcvs4B9dNdz4ILKt6CU/fKYbtBrygtDIAlAd5BwU1gYCe47KA5s+iVj31jHHQm9YwV7ksl
nYfktzq4E1MSnTWRFoTuLrpTtyznP+b0vii6OdBRtkMb59uLAYSWRekwGaTI9TSgzRk3Kgz4op4x
53Q9jL7pst049GzWdXUzlIo7bzpZK5JGq2GzowJvQtEtp3jED4FbgzhjU8whZW25P5Um9dUOiIvD
cce6ViBzAE3WjSL3MMcBOp/D6AZmvYS9UffL9siXlOpflIJfOnrFu5Y+s755cxRTaLqgsZe2jwEw
ZEH01fjixmXdSo70wGgEfxBVfTrsL1Npw0z9luBv3Pyd/sgYU2bjlHgHxZ5TaPcUG5CNnXtFadLF
yVVY6gKDX2P3Km0Y+bPgEOBUn9Yi1c7jKu6LzFS+SQC+3Ox4jC+JhgxDNJkDnoL2vR0Gf+3gWaBk
DjDDuzx+60TOIrKT+B+6my82sA/ZKuA8LAsD0sTi/6j3R0rejoeR9AjVYmaUFErJWJCGB71IUvr/
In1TRUGALqan63QeQwrJrnpfN2doJm8nlW5/TF6/oDtEk+Zk7qayuX2kn96V6lDadyvOVSl1hTIx
9WP3cBzYf+4NN9Qyi6pLpl4bD8L7eJJlXgoMdU/0gG08f4V5BeIrtjdOZ5q8BRjh7ZqRYXxdJK3d
HHdzFOLOfQ7ezd0ZEuWsOUBSwfKJomKgP6ipKXJi1WsDO6ACRy1AO7A3qYrWKAwnz1Z1qyzEkOwY
f0g5BxVO2l8ToJI4VRfWj4k2908LQcaX33kJCgwmBoEDSZsHbTSimLyB+fdnslREjUfrIeustS7r
94nNn2EuF1vShgs6ee/LytHdcQhAkIVsMbt5cdbMyvzty6KsjUJPzkcqmJJB2OAPREPd99lOLJdC
c+Vc6aJ01o++KNk+0wyg1r6mqP88H7x8nO1kBIxs+PZwvt2wWCmu3bVZzEEd+B9Tot7ZwaX9ZcFS
HBKmE6U7fhtlWeGbOVR/kA6gphy8/ThjHG0qZjFtqP1vSvBIurNjnujxNJ0a+wEikHYXMjHvN6zI
sleZ9BeNdn9vtA4BUOUfaN8l/t9tox0WDAtbvHB/OKX+hpnnykGw4PP43D1llfsNXe0nbrr6MRTe
m0vhvM3pkcWEpgpqGCv44NBexjKkgIltg1bD8EyG8hn6gA0FCajOvwF5pvaL+rLARPR1C7Hml20V
dz0/s45H1qNc3jDWC8jbU+QGQXp3UTBJoeUhpRxelN9HioZ6rUi54G6Gbk5PeCSGzB7Rm6VPZnVm
ug836JKeqaDC3XKc6OS3QVWl66VrZ5JsN8b4nQQdDiWfjbHt+PFwHK7FuOrElNVikh9o1+m3sCvB
uukquuE0QPopbvIFSRmUsF079ebe9ArpcSsa8KhgEZk4o8nzxoSa/WKa8UQV4A3nSWZq3L6c9VtG
gWw3gaG0pmvObKnjKO9nH0BxMs4Mo3YBgYZDbg3bxuFbTxEp/gLs0mKQg2aGZaLJIWQ9SL4EtCiL
g6jIgXPXoybxK6H5e5G01aqG7G4r8Ni55zgN8tvrSkEuA0HbITG924CWjQbASpRxbV+fOPnpozKf
r25ad6XbPP988FNrdOnWGeYkydNYcu/mAbDUNMYJLSV/k3P6CtnEmdk8XHPJY3Setx9zy6eQvDG3
m+QO/G4M6otoYmDjSXzS5kwFxIL3XoIkJVDswT/YdR/PKTTTxddlS8vs7ZrM2yR9w0vGVWfyda9g
V0NNxVerl94xhtpIAwDT5onpMh4EcQR7Vg4/0nB52ZKqVs4w+Y2Md983GwRFEajncbYEXnab/bVV
AVTZwUS9qiw8Paec0qxc8HofHx47xtK8Fs6yIa7YZ/8jLDxiTvYrxcib3IzwIgUWx3BpNiPOf+UR
cw+cOqVcxMCc+TguIWQWPm4xTYHwIq/oNGnQ49eCjYyjn31xFJgPSApQF85x1IvJwHzn65k9NU6H
UsLeP4ursK7svtoUGmdopu5gB9UTrkvk2cYz53slkjRzi2OrUg5hdTiXHnwTUczs3I62qFqUfMau
Mrzw2SHgbMsQEQEeKGaZNjzJnn+tS+AKIHG8krWdsFxNB05TGu9rwLm0WkxxnadoO0BpG/bovlbU
0TrcczPbWnKI/fEClTkpyhKOoqpXRqiGx9LRjhviIyAuc5RWuWQNoJimrmjfUissO5Rl0gaHXX1P
E2gk9gTVA5Mf7X9bisxxZ3mVGKsXw12TJdvugCP4UAFhxnduhudWYi4/AWa07uzvSxzJL3bxa6ep
XRuFvXKFvQ2+RUq5FDWrMlEd2YNRw2f3crB8ARb/F7/xc25VtV5gq62McjE/Gw40fzzdwGbwQ3Ru
1+hWsfbRLNlJnsKnaSWwS5neinNq+RCFpCQ+akGCiyGe7DUZpI/Xf6hfLjvhRcO2egk7GWNkFf2N
gzTU55jEpG3WalO6Ng4m60KgflMA2gueicN4hJ30wj7gEACs9FQY7arDjX2a8PlM7S06pYGLVEeO
EVJxH91FD948kE127b5V1Q3e1dUHRiyTSsYklzjhZN6Ea4C5dh/vP9Go2AFTmPrYn7T7CMv++wVf
qX5ajPSciYB6qB9qtnGXzRrBYWcdUQUmYGcWwQIJbYCjEWFsNteptRMw2wDgi7jp0jf2OZsJfqoj
j4leAw/um/Jw9OEekmCuBxkMfKGX5XlMP2jkrIdrfLvCFAXH3qPq8Dgvq/HZ04iZk3dLgVYhoDRN
cwWTlP8EwBxrw3wmPd93sClilVSMAq15bk2gKfw1PcgbxOsiw6wh103AMnbOehv6L4TQ/jjbSNis
uy3N4xR9iOGNvyNdD1cHo1U/Uo0R+uUBI16J4lZp9EUWovsA49XMIy9f3JHaGc2DxCrMmUBTYcyx
+IQvZQ6sJFFRRaPdJDDCFmg0ZLUbjrKYJqgxC3cAadHx2JnWm6Ui7ulJOw34x53E+VBXMfVIahqk
TmWv52ClzB3MGFchw6oS8Tv8m7Us/dHGSS/roYV/UqZWvEsUoBdJCR9lg2Od2WeB/xIjZQK5E+4l
wjEtsPz9Db2s7o+QQARFyd6RjMefqRxiBREPoH8Azy/Y3avHLAtlil87Mi8ph+fPShT/0e9rj5C3
9gTb3TuinhYHToL/MHEeY0DdELxqgaAzviqnhSnlJ8udxkoFrCIV05bHlk7DL3iYDNHvqXEjASxG
7OHm3eV85VFGDGZmCoJpai6vqZaky8kFQeAfrP4up5UTpNzT4197MafXxK7gN7p9wkWOvAHSDbWM
Jt7l3N11LDZCBH0CpQPxaGJq/OnaH7E0grCafzlhiZ3ElisqZ4ZGw+Tchiq9lc49Gf9gCbcPG1sq
c84Q0jmAPWgeKrleslhh7V9JnfwaqbMPC6gCnh2+slvgM2GPrGsxsIIjYUiJrcOiiNvRDd7rUz6g
q/xAOK2FOFPrUohNhVPDdjyFs9Pp5eJP7P+KDhwpvrqV4r6Xd1xYq3ZDz3kbzNNqWGNa7zxrLYH2
wlumPsMdXL+RWTTFk14Fvi6viaJzoW81y2WGFUyUUiyAEaiFBx5xpF+p1TniSuf4FGdRJWEoBEwf
mLahz7pMWH4wkxI6llTygcNz+g258gxvsXYVDHOZzGoBdaTYcGpx/N/WZYy9qRhAkxc0wgcHTUHs
goCGyRSv7b1tqTKP3rxKZOJ2Jevd+1a+n6NHiulOhzlnRKhKOfvGkYYMC2LuR8fN5U0qKfcbSmZ0
wV6UwVy/7EAWFKqRvEdPXvIWNPdyyNIAFVc1VFJZKHoSNJUJLm3ZwlBSqWHiKcw0bYFpKeB4AXLi
VaErf1LU4fQl512OEou8TZTK943oMMQhQIUk4gmTNE5XsRoOcgMEc460d8otEMMaFuwoVXqCYX/7
Q8RNXXlKlBOEbyCSIqZXwzVbV5pbUBhdtvuxxkCl7L3pk4W7DVuE5oTQ+OxBLTryZ1DkM3VdzitO
NXYxh/MkhDU9xgdAjAiWEcGN0zDZ4z/Y6vWxQDRfYrvtp239wJUm2rJe38g6WHG4ub9+MbnDmTJ+
Eitnuxacv/bTNr2MvHQmUKrQYIZK4O1Wbxux8o8SZ0CJntTeEQQiiIVy0wmzFiMQIpLZYiEkn4b3
KttlWMAH9By+W5MYI0AQmYFFKl+sCn1kstlIrD35rghf9pbj6h+qhXGXR9f8UdgDEj8T7+8g+r1P
yoOlUm+WGfvn6w0PZFlhGFeY5qtm8xhLymAG/V/0erTlyRubAfPD8fneRKdIbP6oT3hqakUSzUIq
N+h/I+2RaUnI+eDw2jzFoyb8Nh4O2l03g5HkYcAIS2dEu1X/wIXEOvQdQn9AMTXKJNSKo39S7FC3
PIqcljxejTsfB3L9MNQyalfkKNszVvq78sApJvnRYSXOgf0oDACDRPDi3mtYGB6ISwxvrw4EWZVq
BXYy7LiglG5zifIOW2/BMA6PhYBFwV7UCRhMA9Lduj0ZxiXQN0uELldzaP5ukUOf2BuuwxGCg5mR
U0knk/b7+no80YDFmD2+KJzS5GWTmavQLOGz4QiGalQWmGQXxLCK9hmmoc6JrZuYBL5OB540R46R
xY3FrQla4I/EP59wktKn147yhdyu8JV4+/hoblT2EISMwMa9+e8h5n/V+vnveIqj5PCmEsF+jg7S
egsJdsZ5ZcjolgtlPA4W6JhMCLZhGq/EUHmShG6DlReU3Ko5KrbuYkeqgtM29UKGu1G7t7qU4ltc
lCC4WdK1NBfZsTe7trlkqiI91ZXEWlOKh+mElHGUeojMO1DNoHAZ8Q7AMGiHExjMUKbvAH11RWix
Y9zpEXDqHHVQsitRR0Dut3L+71qs4fZ8UCl3sMXMoQFo2d+xk5u+8GQRVu9HRIQopaS0WrCkEOBr
PzEXZi8vU0L0qnTi25J6btMOm5znuZOxtnODZb9OfRVjRoSHkuxyYJfEvRRkyETapyogVELb9QNu
Q6IDCf0Cr6Z3KYWjh39T/yEpzzL81wFPgLyeowUetaNpXsX1XdkEufO5HDnr4Kr8uZkkUYCmc7pp
tBhLR5/zPTXtLiPPFJaq+DHgPBd3zZAAxcus4lD60kZimIE0oQSz2riFJMl5IRJgqScYEkjycZM0
FJOAbb6d9AASp3sL1hY72HDQoAzWosfhN32gx7CIhY+t6mOEr8Yt80Z6aGdTqFavFkNY01clY8i9
dt2qjXbKi1IvZgn1t9Me10e9Wy0vnciIQvbUQs5Xl2P3iAYaGsRo8wGSU0+23osWgqjAGT7npTYo
3oLAp3LnD1xW3x/hh+zDlEgZ2efmarcCaOJ9XI6Sa0E+Namk+W6FHqtZQ5ww7dt6WypR9ywkfadS
HFiE+0lJyr0uQbY9ESSEQ8JjSODa3oyeRxzOhmIKRtVZx+fSuIeRDcWoVN8IhYHXK6V/4lsdrnak
T6ptwpOmHbOVgxWDLUt+DCe2fYBAAOsjrLR5o3oI32t6B+2oZbmJq5ZnTwJq/rbz85BTfushVTzH
Wcxp8PKnqL7hguMYeEGa8xF164mR/R+I9Q3Z/IPPzkgbKqmNHpdhlCSnclaKvV2QQyd0NE83+Kr7
4H7zmM2R63MP8/tZU+yYSNLFJmq3qSp8lt0yTXfntHRCfD4JfD9KQlMTB6RjldzRN7oaVLveyHj/
t+4vnKr5lI7AQ6/l3sbv+fsWC5Tcwkescj8INNMWQqnikfjLG/g7akwSxM9+r+mubBBHS7a4i1b6
Ng5dbl/2kMs5DfUIfqLuf0k0DmDWteBC2w6n0ZUAC9jrO+B+TJdzJQTDWD6/Wywlnu2IPVvMNbpD
2mzd3uTK7qclk5zLsmqa6RcHA3S376TfH3NGlBKsWJcDFtfzn+7bzofGjybCt4cEker9OkfHputO
Vx8VmSNWaKH9cLduBRStjmG2rLgDy+Ck8LLfK2XDre0N3nr2ZbDSby/t7lmx9t4ETjzCFd1fEgrM
HLW9cWW7RpCZEGNyal9Yj6d2vrbUy7lPrN2zF5c0dkeo5+xOQmXV/Z5+23jzvdRfVDxrB6iQD6PL
LnFbdfQSTXGoj2OJhirrylUkm2/ik5U2MrP7BQJYEXA5kpZwP9H08jQqFOqxgaUU83xXPGBLMo1U
xI5D+8ad+vahVwluwQ36jZ+plgiBOBhVh4QWcQOBNiS4zYNswOQneiTKa/WQx0RsvtlF3u9KHMK0
FcKIG5MHIJ5IhHFHIV+QfiylnomLWrJEkX61Co3ZV2/oVpVJCoZ9B03ufH8/Ox1OqQcsj3cVJBQ5
UA7BV/ScpyYpLFwU9XJaGvHQYVdGleLXaykpXHWlLxefYhqeM84Ra6xP/kUjVT1Lxa6RbPi0VwVL
lmJWPwzSpFA32w/xS64VchdZ4JbHo+wo6Y15S7q6AngRn4xk0xCyI0v4xaWqrZZtLHitWHF5Hflz
OsrKLoHWqfg5sqNJNZbrXnCCJWdQj5F7cOJeX0EGo1xrsC0GPutl9yfAsg67hYXZqss5JkEd61wa
ydrPpSs/zr2dSvfOyRdJJYcF22bbsnhTvv3Yk1fHBSVjJtc8tV3ffE3CP6Tn+upxDf8l2jCx78Ss
jhqpz5yFkNy2fXpxztHJz6HOskGcLI9Atc7t3EXe3+1n0Faq2+eGRz74C01sDR4IxIAiyPYgR940
BKPxoX1DmwGZVfad3tbffmhy/kURcwv8sKXiQbM9Ryyvfk1SYJpxzz/FCu7r3x3I8mapaU5WmGJx
WzQBSUucICryBMY5W6q4kjqFbvUQ1jGGGqeAjZyO0PH4IxxvfnCnrPq+b4yp5RDcnk4ek9WeM4Gv
Npc95bfvm/z5newTy9iQTVDNfOcsjx9DbLR/q78PqjMJY7SOO7bbs8Ro3ENVre+sQ4JivVfm5HWR
7AOXRjjXIM9/kmucmu/rV3nt/aoT9JjkIK7MjUhUlFB+E3+AKqCbkGT8EdWPpbsWbs+eBbQM9Zxy
UtzZoA0CzlC+cvBieDtjZy64/q8g7+k192/rFQnmD+UG9DSrJecUeL0Wu7sq3BcN8alyVK/8LglS
A0OhcQpjz9n0bDpsLRP38L7rNVh9NBO3TOMeEDkm6+BiEqUZb0YArS7ITRCp2WBLavbVEhpbdPeg
VnA5e3Gc02Qh/1Z48V6rjANJdwA6Xd72PMDetW38LZD4RH+M1m1BWFQG5i0HYd/c+8N/6mIisWVt
7OWIJ1wVI56NlItmgyHuu3vmGIooikSNS9MuiJng1AQeXt77Z7qFiD7hTQhxb2wxfFsZWCL+BH9V
LUfSL1NgT3FuzkoGxDt7dvL0dt+CzHMPf99u3eVSQO9jBkCoXchfElUlhOut8cpZuwFquIzqdYrB
sb3fpd7s9OLjbslU0doc7H8vx60ZzTnEWKkomZQzfEdWMJtKxawpw5AsofJKgkbx/v9c1r6R3Zs2
IjK+za4Sc7Wb0Oo9ECtpTevGh324/q/mR8XaNfIkSE3yCOhVdiMNmm4hzR5gVPKfpFDjgrWzbG4h
5zB5HJ4NWYXFOq9H6bZBsxqkEAl0CDkFMo0NNgu+OkrdNCT05Bw3ih6GKLJD5b83TmrfjtilCHow
XYytCuPQ/E9qZrpmUy+s45Z7Mi7DIbGXpmorNm/7YzAZ+4c+xWN38EFeGDdwGZz7wbMiFZXDCCdY
NWl1KGG1Sns9wo3Ir+AxLD6h90pilETVcW7HSmBR6MBLIz2Aqe/5VG8CiI2Imq+j6euP7f9vroq/
I4K1P4RHwMZbvjaJyRCC4aMKVGjkjdIXyhPxWg0z6WLMjAeHRHRUDwTWC1PzGhnN/WA2A57pR2An
tSLlBKJfyFvkiexdg7YKAWR4mmcMXSCvq5uAoDPnO2MyaxNCkG9cqzQPtmD7u2geoGlHf61chkdB
AF6QxTtP6j3ELe0vLfecuRoQr3v10oPL+hGZ25XDVMoVDYRDiZD/QazFj930RwOPQZRIK+k/rzsl
uY8Gmn09ERetreA6SWpkEtJiW1XjrCiZ1nniUxCNwey9SntyLOyv+r6hWpDncd8SNcSfBCb4iGw0
7hjD7tYIAEHb+jr94g6vFb3i5DOtisjbSkKWiv6N+esB5R00ithJwTCz0Yjvp//fl4neL23tFRZS
2ZpEEQkHUxOsL5sqDLthbq7Y149lHuuT1JP2DM8hqbLTyMwWhpIdRqLJV71Z5E5yKxX+JcewCm9+
EMxvQHJTxrxFRQP0I1lGqVMkYSN/L/nelhpXdiwj0KngJ+3M6cOtLWmbH3xh7BgEl5XV5NbmkfSf
7L9JWukKrBNXG7jhNp+7asUD+MqscXg4dwNxyc2OEmlw6sngkbuQOc+rQys1NrlHbId45FWoBTtI
NyGWnlmdBTP3Hc+thY9GY0TQShEfyzCQSoF7GdZOvYd7Cl/9+pgGaC3NSckxjCS7adt9XZWvhua/
O/f7SIlZwvPERaK2vpEvFemXLr+gYl8ZFX1pvDP0caiXH1gR8xEhYvR380pgoXtn/qkrg9Lz3hwS
99sOZOJACdOpy7APHF0Mo0D4jZbkj9EcOCqV3pilN8VO/ZTwYyovTZpfrMNt+xTlSQvFTrpWOMsn
EygghtLYYYI4IBSNswC3cpSpLJB2fw6DHDGeUo03EMhJKiti/S4tpvcTteLXAC9pPmMxq37sM1yO
qRLg+eFya9BKvFS5mg4Qjyf+GC5zzTJ5O3c++wVWawVCOYN0cKdNjH+Bzk8zhKcOOsznM+37uPCV
clufYzxMcw/PUHgAh2cowoISrQKWPv8CqTfJjttPjwqbPu2QIrKXntWXwc0PdCx8tc1y079nkz7i
5Sclb2YnAK1XA5dysnmW6djlh/5fL03LTlizllrQ/DeeIGi/+7kuPfKgIppHMHFe3CQ009SBGxIl
6FB5p2dF3kN+E0pLZ3iv2tG5tOuBFiBBwydUEayfnrKC1J//E/xWyKG8661Ldo9NdZMUH9+xyA42
jRYn98DxHQdIedzyNiQHVwHCXj8NABv235Y02Xo82AW/n7ml6GgsclKtoG0E9fasWhYGJ4OCu66F
1jIrjWIahKP08Ih7mQHlFEDAN8vCF5TXuzpG5mawQ8rHpk2kapcknzXHRyf80kLngsgyqEfTNQ7O
ANyLmSXzChK5xtnyDlg5RKXGavDEBqAtH/q55Oy56Ck2l/b6Ys5Agb/8xIp8X/xpRZbrqNy1Ws49
vsg5ucHUYytPI6KvG5NjoFJJh4FQ1faAg09yWsbb/pN4ZbUR+mfkBPTMt8xzOC7vVyFtivzCoMcO
Ub/7q5EPkVeX0PAvJ0SZNo8GrGVE7TcXscB9QzUT75PAf8huBiSiZRDibY2LhvKhE7665cxBZQEv
gqrStM9Of1BhPEhSi5hvSOJLU4iF5xmGHC9iqm690XFKjDo7n8vDq3Klgr6yIjyFlHTDczT+ZCHz
6ZYKD19YLWqRVjRl9FXOgKUNiUI8rEuqPjtltWOq0yIBe3Pu3Rc3vlKhrAZMZ9Bu7c3V8FAHzA9l
ktc4Iu+i3mUuKTZxu1tt3fbx0DzJ6gIYQDcPpI1ihkGOyKKW2pIkDstPS2OAIs4xxcH5pC8N8s90
XHpkd5TSweFKp15IILu6KOcQgAlFcg/7izpVr3tyhVBsiRwmY6nWsckdZ6VSXotuEtWK4s4ckvpw
hd99cftcCjP/wZKypzEG0cj96ormeGeA0lo87TTfj7Y3Icq5jx+SrgIoRxrRKtOu/4VMZ6DDB7T8
6qSEoqZFAcmQgTcwG9C2dJmH3hc9xnRkdYbR+WboKWJPPzSyy5IekFRyl0BY9bVp0sTBBPmshpfo
TmyBKQNgOIaVf8GnrqCVxQlSabom78qQpYFN0HTUK771VvGiLiy/QPeMXkQj+tF6K+8W0AnoxyJW
wQZZpJPs56SMSJJh6ftfLsDGojD+immoTBNuctNZPmqgUJeuUy2j168ENRQ03qMn5UetkqTwqnnV
oQ/8KeIu8RtEki0LtpX9Tsd9QRak0qvhzurFObXMXG2clrexpkDuodNss5O/wra0CcnYyTOCjQqH
xH0+btQgD1DfforjjTJUGz/ybqinFc66G37+/UVaDkUc767db0S4niDQ26HhehOSiZk68+WR3Fhl
Y4JyOghdYpfk4w77hexetcbW8NnYEU5NyP/BX3xAZu301YpzLGMz0cFVSy8XnZu786owSoGrC2qO
PQHFEG2jyGxuhEck67bWUi5Uh//ew2rrzHNwfghBQd8sbzaI8+hQIaL+lcOdOIAvQq8EjAghuJra
Dx6SmbjywC9eZYJH2F63a3ERPkYl+tiwTsU70Rc2mFLzAAXTdmKki0e6VqFaxwJE1niSK2B2UJKf
/6MPamCaMjgxcgWB1pNze+7XRPKRl85R/oea8eHj67YB8fSxBV6uchuJb/WvcntBnNahjLXwPjA8
3TRTVBSZ/eVkyI+k92qEe3OzIWRQ5V7CQ7tH/3ni66v9GRNI6VDf9rX+PzsrRwG8GOZrhW7BsinZ
kGGs2T9GzhPl9sl4Il4p0fAsVZPvOgQrjwWiRnTsBzj7Pw9lTazRqwAhb6J4/9mJ8aYkNY0eMOjw
cMqeVfeBo1eLpYvO65KJHKVAImD0AuFDlndL8FD9YAr32Uots2rlx1ksAPTIBLRLgT97K37h1Nx3
aM+4w+hdJxR92q0APNYBprpO5z6cV9uYlVRplsJv+K8PV7XZMRqDpSDjCIH7AM21wyf8SytptvzQ
JOoeuyCZYwS9J195GW8wt9JIolw87S/sryLbJ6FMpXMZLKJ8HZkvJW4lLA4ChY26shKFPQ4UZmgG
qAL12yKHcdOIOK7Dv6Bvb2jbQPkZGYglEL8zJo0iwBDL2rVJlPGQz0Lps2VmqJdyTye+z4brr/va
uBeHSAgyWAjrUsdThM2puMkgkxW9Q0WaCt86pvNMoapm7cryG5CQiJP3B7gYAMciBE3xayiTrrdp
AnxxRrzT0+DohJbbwCOBQu9qX8H4DPtEX2WCa60gfnSkGLxqfn6RaVJnDAn6eZIobXnKBkJBaUn3
Rwdms6nZCyKaIRGsiywCwqQ+Zntg6XimatWFYuhd18YiHraFLSkwYgtxA0D80J+Vornizko+uhhT
9f13NI/98nqpyuSeEAh8nDVeO9dB1N9kNpF1711N3cQQaRwi+SWPSAOU3R4L+pkGDiXgfbgJmnah
gNv2hfG8OHgZUdhk/evL+o8BIwXWbxYbEA7HMdgRaNk3kdHNF7N6B4B1GlQXx0WV9S5y8Q4TWzPX
NEFZXOnmQ+BIwGzHx77xKarz/mSqU1LCCqwYlhzyPQjsBgDphfyaQ6HEmgRNITHMhq0e+5MbxtqS
SNfuDv/wHk1fhbTMG+UmemQRxeKAq3DoeqG53Ibo593EpYZ/7q/ca1DqZM2k0R7XjbOu/MweYBbJ
0vK1JBfAqN4M/q1UcD7/tf+QR4vchI0n1EpJQ6pRLq32TqAAyeeyDxrD14Ls2XmkM5L4WrHecQlA
ThDhiXFw1OCXsbgEiwQiQpSbuRHfSyOC4wbTZY+AEic705XbUrzuj6i8GXXnoMrinRwsoyfwLLuj
hKw+4pLlzsGSqYF2kZeabWsSA0hbn0jyV4AhftwXWAHNYeljSTmXVO9oQ7a6HHQBuRF0UnYMw0tl
AASHoSVZxflxMXf6+4CcS1K/YrAA5SKMfxI8oZ0CnFPN2IT9OEoH265L622VbvdDNfiQ3eV5ABbt
+SYK4CuYIm4zqA2RDWXDAcOPa/1Ok1cXbfeofGBV5qEKAAcnyomm8Witujtl5xVQ0MQApDeWoVma
LGBrztxu0VbDB/yJzI8XRD2UES1FnS3EA2cxvhoYPC7M66k8h2s2yrRzvUH/ijSjWNWZdksufWz1
/A92nUx7Vw8UkCVZrca8GUNvtVcYINbpTAI10j7nny92yZgNnIkcEgl8n+Q7pBA1X7zEgGSfD29D
R77oTy/U46jNEqbj5UIuQlljvy0+8MSD0tKCXe/YERdPKcbyy5hmLhqAsWg6cQB/8+EwZ53TREyd
DJUYoSkNAl8b/pGL5APn92Z6AIbw8Xsr35v3o5lw3GXIKLiF9rQsy2nCSTHNd8PQVgQkL4YvW4T5
2gv4xl8CZ1sZm5WSm4C6k7ubnUCuvTkIRTR1czCHozJr6rd+3pzPvcS5tXq8SxImOkZ4IT/9HxEB
t2tNtVLVzFpfknS1ojmcE6gZ+oHytWe6mtZOI+sL5DzXxKMmWqd3LStiQ9hiZIvKheu9fptN704K
w02vOLz0Cpg18fcThJE5rFKXJfdHP/rqPWykbmQtYaL5mYBQmc0vH8nMRHF3JzXW7b16kRvDhN5O
X7XPw0DQeHK/YHYuor+FvxbnCMB3QtKJPl65amHo8LH3cgdS2jBnsBmMTSarkbU/rXVaO/7zzJRe
/1Ie+mb1LmT1936AyQNg6oDLvRAMUNktbcerLn0tTUiXdhwfQ0t8qxhUZW5b7Ip9YzIRCXD2xBkJ
vt74Nls4ipSWBdKNQeIzVsg3KL2ioMJa7CoFMHRNnJLtyZg54HyX67m4j/7EmK1CQwp/ZZAoVb6L
P8FWd6/iAoyB8GxCDZsQ/xzOqaszDFpiio6h+8brE48UWA9XEXB9N7D6wDMAjcGWZE6xLKCjxz0N
N6y1SuVjxYCu6MWR53dIaMD/dOdGh8rYrDfNj3vi1YFJkrnnsWs7AS5UbQGLXryfptN68doo7fg0
Uh2QUqUXkWGpS8Pps3gPasV9b6mPuErQ6kXcijYt6GVoPUZAErSmZdD5mqLddFEtRDPOrzt+cUhp
jaEOt9nO3Ib6DNIfZpGdoYMbL8apDPy7/4LhSnKjZXasiWwmWd7DuNVNsLkLRjAYX8Qlp5cskT2s
raif9mPjPfJ5jtFTpyBQAYe5Cb1iYLBtBubxygKmTinfuK4pT5k00a0XXJX+ctheIw6/nDsbX4LK
OldfFuMNy8OsurDGPHqPnreHuzRZEjS4ouIYSch5O/PKI03QvsEt1d33L6/r1hFMHK76vHhvnEn6
x2ze0C13kctqWMwVpdpmuMzvIFJIuB7f81ZXP+JdRXEMrHuc+uRZjN8m9PkmhfLQ9OEd/3sORLOj
bLagpUGRCpx8su3ruJf8qkm4bXIBYZ4vZPEv6vUabz/aNWF7kwpNk30b1X/6Ch/8u2oK0LmLPp4G
YhTKlTEVc+72KGqlF9xitwGeYyJap5aWe036pE9Pa36DZ3wgRGSdK5eh2fShFsWJZJjmfWLw9iBH
B4mMkPRQwvAQfWGLnIqwPj79cpQqzEnT5C4lmT5DXxWPBuU9BvsB02NqYvH5j6z2EV+6dJtEXumR
dXO+Slshiuu6cwphubNFPKI21k9ht/V+vc2wqea5IV8gidA8XCfwnKwcCPRbiWFYO9fWQwxpVCbr
xKCT1K4NMzFYJdo50IhJjWgV9ClVupu6GkcY10YzOBDs8TOi1QQwYbtFsFadkK9W3U7naya4/FPk
yaKMv7obrLIjZnclmkb6yOGH3NTu+422ktM16x4W8Nk1UzgSJSk8hTQyTv+MY4xSlHf+IC1Kf+xB
XD+AtKIR8qklKssKJWhVJ0o9BBcjidPiXugfscRfBt/8k5jfQI3fp/QNWu4rFxV1MbY6xdyNDCRS
lhX2bubtbVJi2k2fzQ4Esk0Bm3T369pYtJBwkoQ1JJVy/otLaEYPnzkH9X97Nk88HuXfTgwzoWqe
4SdOhlSDeTvl+P8WLHJkQkZM905QQe2KGneR6iK67vryV0c3GuZJaYdKFUVHWLomoSsPPIA9HdHV
WUmZGYtEGy1Ru/pbcXOusfDPqsAFPnhSRRpp+ltjrNTcUp/9evHd8nJtuDkrnjMFs97/zKgkPsXr
Ch07yFXDRnjQHs608sOm/9EDlfCmzt1uVKc3O1RlSq7SGHJaei9iQQsYcEaRT+dXsaM+3/hFcOOU
m405PiQtE32pbcFBdkOeLMV2Rqmm/sGw2Javi8fhEWGjDcs9biIqfrXa4gofjrYUfmTKr2s0mgWE
8AGpheTag7bE9H6XmKj2XiRxlOe4lAmZqvfXJPohUMwk8aFj3jzdqHkbxD5JmYZ76zL5SqAZCzwr
QIj9vMVL/34iFfd9oLoIkh6A8KbpQKdQpzwbYVwxgmm4wWW7QaNRqwc2JYNHkkWztv0A4ZdrVDUy
H3h1ev5M+Ah7QyV7pJFLViz0yqYCGx81H3DwdWnbW5SJ3F/5yP+oBiilyQIYA8iDnPINrw6c9GCn
vCfDUXdfJs/B+yoje7W6Kg8irRAw1SpH1FD8k3aPPNtfoT3LPc+Zyfjl5a655KS78cioBFhSwn8n
DKllma21fO03jpMJBXRzTdaiSRA3ZQI5brGQQ1sEzsYMGSc6p8fnZ7hOV9sfVLMIThZb8MmkEYHA
xDoaXcJC5uC7dG0lXyWhPto2g/kOXenpXBQTkQ3Aem5a+zcwz7xoC6oGfN5g7rR/AGpWgepoPpa+
KBwNrE7LAM99xVjyxq7oBvAtxf1uZOZJTlXUBMqWtZlZBZ8Neze8B6afmPlnqPc4sBqAjCbaOzwu
1/EOUEJikV4wUbz6maIZTVLW7t8uKCwPntbq3T4RPN7ShkUXWxkirSRayYU2NmdWQx5p+VIVpeOq
DdcqxndeDvHJM47guaqbuVn7RNmfdQtrdifjYh+SZkHKrLUtZ0CTZ1OBIuGmdr2JlVKOadlZqt/d
2RnNH5VDK5euBkRSFQkgy0l8YIAq5tAGOhjJaK3LCX4w+JPfLdhn+BDtxX33C48CZgpNYO+S8ep2
yONNJkeXJNXJemjHmu6M54z/aGkXBwX9AIbxHPHxN2SgCUGFPNJdzVA3rkUJWuP3ptRz6Hvffqx8
L4qKYNey91RKLMSyfBoP7ivnGEkMjqyBYwk5IvPxgfVVgHXCUxbhkYLfR0MIeIfLlxmiYtq2248x
bO0Lq0pE5tyLLzMt+WujwnCM28TURwBUaLAzLm644NWArsmEYlbPQB/j6RwsvIrJwTCJZEk3DzAq
iT3fliKKWvAUuCY32g9blXD+zts5l+9pfUAitrQqvBquRwUnjDNZkYJhnssKCKiEFqk30fgjuFb6
H0tLydIBAW3nGFHzvbHwvMURhxQTB8a7n68fhquovN6yhAkghM1pSHqz5yK5zzLVvx3dL0oIP2Mt
WL61ZlNVYiReq3kt8Gkg3DD+N/DTrLST6MXTcaVDMpEwZ6SO7DL1Qdwuh9QuwC4CqnarABiw/ej7
Et+fYHyQt2BNCfuRpCOWnTlXvGL8Mj+HAiPYVUz+b99OQaCoBcuU31b8lNXm8Kt6x0cm6nUw+Kf9
TcABVXRMx1joMINo8TlLKqK0DUQXoaDJCReK45qgknOmm+LC6rVA7D2O6XA1DQrw//pttKM4aMI1
jxzdH93Y64lQOSJNz6Wv8C83g+0SOp3kiMtSzHce6mFJzgRGkdkCFu3JRY1EU2m7S7vbfbdNCfje
oaMLk5fiknfJVo3rEvHAxP6sPbWSKrY3yZX3NsByhRgeeJmP0y7BC5LoXP3Ak0P2biI1WIKIfCEB
mv7zvGvbaXROit7Cz1SZf3DzKwg8UIOGDJJLFHMOyoLPn3I1pYdm+oEJAsaCqvgl33KaA4v2TJ+U
esoRy2olgyNUgsUJ47zuWRFyvOvZGqbO6Wy6H0oeY01+PUW/B8SvhAFVCMxJOwyKrp2HhcE2FZid
GUvMs+VrBvBHUZpN8p/twE9Uwzaz2Nloij7HdA4IUSzjy9DqoHjUVIi3OM9N+XrlbuJXpuOQE9Vs
ts8Yb1g59IItvNf6wWPo9RXBnnqK8yGEe/V3cFwbrYZMu7vzuzwmply1sniA+cRJB/RA1aFTGeCb
q+igj46vuZpXPBVghsGHY0i/eaRkE5lpqhKPO6/SIX+eHk6SDJI1yQ95g0VY8qULoRwx/fLwps4h
j7lsxfTRhfYylxy2KPran+ceWJffONFIMuGKfDMRZ0pRmxngSdWfcxC/uKIyASGs/hIFyO2P019j
AxhtuwkdhglRjMB5C/UPzo1kPD0efF7h99mXgJ+iSepMkfEYs/cMnuUAjeVQJYJJX9lhj6+r1WeV
bLakzt9k1tnpF9MV9/03EjOhTeYAtUK05PIr8q5e6HwTdfmQ0GkXDiw7FkFINgRS1mdwC/yksY5w
bQd8W5WoVCUaqB2QsUJQrdDRQtagv984GwunzIPRac3vgWxRID8hfJqJFFu9XKMXSbFVMHFRgNjN
g3XQiE+uRcG9GGdm2CwUSBsqG3tpk/dXb+TChOKUrNgpRyj1WUi1oamSpR81oZZFMzyT05wAgmxU
Drh5/w8sUqKO7FB/rRkMhnYbCuLNRl0LkCakOaYvdEJJt2kaWvRptxXA+2nT6TJBGdrtMdIF2yU5
c8JxCoqds0B9x3Q0x0cxKCbru4gdfWeMA7xWsVXPTfrYV93SlneraW9Nt6vKddcF6NruYmc7lBJh
Y4I4Jl0VUXaMVqhotC+QvPcy/+AQeOdM5bzfOKjaeH2+0nADQLCocWahoimBKRUu1y5jM73gzlLY
jlhLbCktFcxbTPHHRkJN5VT1uCHA6t04ACml7QN3Hv3zDVvA7ot4kKfaaOda0xlMt3q6yMNt6ACz
aPlXajXR2nPWm99YDDgbwjTa56zGzJVbW57GFwfSnfL52peTwMgEpk/AlFhXCIhKT0g5XOYqoTUF
QmN9GaNFW/hU2cogHmj3cNAZLf6NnOZ0H00tj3dK+w68fPswv0Fr37/VKHuPvjNw4+S+cjmCqMrR
0uJOsfa4l60/q2FYbnpy3y5jI+Yp4WHlAbfJCOq7CBTh3nTkO9XuKgaU4DND5O0+mh/7dkuP5MoW
uBPSho8sp/l0tRPbo9b6lGOFVbz4SBt/FI8y7KZ9u+7rAx5UB+gn+5i/rCaVUcQAvvJAgZIQzet/
FLElExRnlvuaHaBG49KLtRMmM+OX011btqoaRfXVK1iIO+zvu3De4cYDxxfpafOUvSCgLTblA+oS
bWjHwts0X8YLn775GSMQvn3abIAAJOhcnbmEwqCrqvjs9rDm4imWC87J9sFfTQ/4QxZGXYj8KMfL
bc6NT3IugI/PniuYkcZmBm8OsBAVAVZ1A5WRloxIQG5jW4stbtNMBS0YfAEDjSJn9Y7+0O2aGJnX
6QVwBwBtkemB9b8tNoCez4WUzOSsslRZ0UYLnrXLTcIKFjdYjXZBogZO+HGd0S6bdtW/KmhhCkGQ
YpPeSUpDQRT4mEAkHRgEaKEVMnamABvN24Q0Ayi7jD+xEf4MSq3Eu5e9CeQ8aloksfbhJcWdpCKP
zS/dGZAS8Jcmo8hk3unt10+/v61mv3FD1j9Qmphe32dO9rhMOZaIuGZ8RJebLroNp2yRPZBdDW00
SQxtm0xXH04IDea6uoBMdmyo+7ktQw/s+2wjJxSL95ZeX0uetybCvf1OuWJwM7vMvkEpSm8UnYb7
4CWFZ39pxgqI1/GWAFWQisuoZxelqxibpTKb1fkLlqwpoYtOpWtuzic5vtH9i2z3vxoI8zTUjPgO
dYrmFjM0Dzc5hBjpGC14YpUHUoB5jMRdlWRY4uYcYSrCUw8zJrdHeI7kDgLTTImkIcu3pn+dIaRT
EDZ2z/qQsPpYZLjRsDxv1xhyy2WiBE45GKyeCCvi36F8QuymVlLw3KR9PMFLnJTu1Ee694Zn3z4D
c4GC8FG6qFlA98HK+CZKlnD6KI49R8eRHxwUzf8sYd4+hjNWrwoja3TObN6psB2ZLe0OE6iLMp60
PqYfOB/gjZaKWjXFNroVj66g4PHHv+F42bYTasP/UOSnLoQUGsa3UFWu1RON8ZWP4OYjPUY4P1Na
fBDOUHjY9sho8a+iG5jmW3LSY2rIrxrEgdguDGSPs1xwex2Sn0OzWi+JD0HXmcB8XqN791PNFiZZ
o2JFpRh2cDl4J0p6auMg9bBYYc3Od//m5bQcOYjKvReQGePSiZ8chRG2+AsJxhlvPNMFHipIqX4R
V7H4cruLAAQDAdjxuBvjquK1QNhb//a3XsKUbwrPEqAe8KUY8U5rhM2I6Ahxg1vZ5sEYHY9l1N5V
5rcyIHHYxT9w30lPWpxj57ZeN+4EuWx38nJbCEPDvRNAtDST6clIkECMCXWXUdfM/PdWehnjO8sN
HBs+zPnnuiwMcqMXg2dwRMWb0MoJ/G62XG0/k8j3ypBeLJOZ3xpLmloFMO6ufUK1Mxu115jWNf/s
S5L3X51y6SLDLCoSd5Drm+CNma0K3cCOWuaY3R6k3rUMfFKkRLIE39xm6jAkU+/c7wcIDdIzgkX1
URU/Ecaggd2e9zgc/3ujL1mTZHnNy4x/m6HCtJOJLMyS/hA5VlFvdyfmcy01YnVVkY+eDy8RRMR1
juiTEmWJumxT0CDYrNI8oqJAuBZmkhScsahHVm2NPsaTl6rD8If3cyqC0Hnr0LGOy7VkqPWGnAzw
L3KcaxRzzrx08xGipeG3IitBJ2OJN0OFyrFQSBr11Jy7G8qQfdUsOpZu9pirggFApbI0qDoBED7f
R48Am9JnJ1e72VMSwAOLUwZFKPTXsDX2dIMNLF/WK7P1vv0EO1SLDxjyhjd7E++W7sCtFR0x4UZh
uKu9iTi59UPQMsk/riVeMcT2oLExoiik5CkDx2snz2WSh+I5zuS6z1GFqKMcstnd4qzQ2q4ABhxy
W5RNN8hyn6MjURS/yf2zrQ3wNXLF2XgBkxPMQeiiSeblXvsT1Zy/S6CwI6i0m9rY7ZPPMuweGToH
kwRZjXKTNyl5cOFOMNcJoOFST+GPhddg8fU0JeXd6tXcrgtKfKEUoFxe/bPa07YtyQaIb2Gxb3gx
c7+paqYPzf+EkIIK2NRBbdG8HmRaQ0A4XTAxz1wOzkUMeHJNjsgeqZvUo+L68WoB7kIt6BR2bGrf
FvbkrEX1Ms7V9lNiMfBGNslJZg9IsZwK6HAYtxMN3bxUVrusBgxLb8X81ARvSE1FhlKQsp2oWYuD
EHTMrx8JhTp3zJyVNYnGVq1ZFRSd8LW136+7CMuBLQdE/5ut+rmnzZZUde+9ackaYFkNCuUEsQyZ
CX7lpYqGTTu0LWHgkSMzRiWDlYhfrYCI23mzZN94X9EZYxyqDZZnmnhqKqMFdDlZNHpAgluja8wm
wOEo3E1BZiOEXIGvi9sE1JaCUixyYmH1+HfKozCzh7uhCMQCYDN9wscYFc14L0iWLU417ld+Ylmy
VAtj4pS4VSgNqHUqfQaD5fqlj6FTTnozTuVXseFmNTj9ysOD/AnMG66jksC3mwU0ZljUF0aIINc8
iQ6/PB9AkCXVxz6W+xtyba+TK3qtdZ2vBcbs6gyGO4AYuAVCs9yzLJZ+1tu5DtuibKnxEWrcpOCR
Y2AaULDgsc4bQB3zLyyXsK1/lJ/t1SHm/dKhfR4JDG6KfPNJoJ7XS3AWESKes9nnA2Z3W5HK8FBQ
QTKGIcw/NqbzUytwsHn1ns6lba6uEJfn6Wime2RfoA+/mFUFwArWOLRizerPGSfRzlC1U3ELURR0
/SPGDScZ7t+1rU/fhq1A3P777uTQDzzll8EiCVMWS7oG5a/tBD1sxKcfhZ+9p4EtRVNkU9YpSiHS
435yUYbzVI7RmhDlTo/km6JNm9/qPjMg3blM3XLjc/TQPEklMk0cC4aApJMNbl46E9mJRK+Lt/hR
8BRcexo3XRfWU49xu7K5J9KDbKMbLd+LRh0JM8XCZUnLzbuQNb9bek3zFU1XhSfhygtMWjTGqJ+F
4JIYDsfCqETcN2LvfK3uuGiIGPXkecMbIyU3BNgfCo8Y6PytAaiBWIGp5Dr1x0piR0AdeexnZgM+
FSitBYztcVWPfOrPrQ+BWo+eV935g0TD6wONTERm1ythKsFhy2ZQubjBRKTYZZUhanZRUWbEA+aU
Ddq53xwwLeMB6PLMoopNyik2S1Ia6T6Bazd1sZPZ7L1KiZ3ONjkXLDVR9cthR/xeosbMcjRgHuyS
m8Z5DrG+wzVwAEuQuk2wpBWUQ4t1MhehEq7kiOUlkQBULMVsGP1vI5PXWWxVutiXNf84J7Nl+JF0
vJSj7SyWsOQ9LcQgmvGwZ4XGnVUWo+EueDtEbfhAUfzuSA+rhOylI01tPugsmJchZIJqD3uPkugq
UMO/x8qZnWNM7h4LRZ9+x7qEyEU1TrNiHoxVEkECA1kXnTQ0X6m5hGoqBDeS0z3xWgFJkHYvNHU1
33oS6/dAE+CmHtsPT92fFGC6I+1ei2UHJec8ByykvChPCJapnDj7azxcc0UDjlRnz2FgxOxJF0e5
MSJqq/lTAbPLMsYQfgNbUL37ZMdsWT8hFP+soZUf67yPq5dN0gdnS06/wfg2KDPt5FjqSxcxJY9s
eLLpBGZP18EGChmqNGoz6934kJ8OhVK33AbgWvo4OajoiO6Wz10ihmC+bVeIHS21qcLXT2xe4+BH
A4u2vjBkxhYvTQgfzbidMurTgqmvudXsw5NXFsBEwFFLsWjRTCL9k7nCQjlCkkIjs9b4VsOE4FWV
aOfmmfNK/z374cD0Yk4CuyOAR1B1vPmiYtCphickYz+rxC84/tbmvpZuI7JWOBNLSTTQi+XFwTPf
tkJ9JD3mMUCKCxmggBNOAHWoHTZ5hTqW19kMMWZVEDf3kn1ovl+t53hwPHUv/qhDLLkRsN72ZmDg
j2MupSLPxGk5VFQQHWV5jq1FTYf8EVd5tRYXouUBYMIMxNN4f4dVsCeto70Ygm5TcM+0foFs8xsZ
UjIwZ1zUIdKMXhk0+zd3oquVtxRjYS6S9QB4gft/QnZh89nsj8nzZo3QNJrm4+7WyHz5ieTdiCv3
QMwsIZWCV4SOLE+ld3lBSv0kpKTBeaJaAgXQSzZbxwBRDzbnM1+B7DJ+PEl8T0QiJtZUTqRtqJTU
l+4Ns3LAloXzFoX5hMs0o7oCIssgn15bJhKLLGo23bFVEB5lrWe8eSAT+ueenpNVQjWq2VOomcda
lcW91x1U/xqBzseKtfXLdMgu9DL2G8E7CILYDpG5nqyj17SAPegnOB3gQlHewnl5Sn75MbYAeDbK
PnzS4Y7P4ZTn0JJ7Zov+4okYdd6ji7Vj6FnC6v/sTubAc1iCoU+Ft48PHvloGg9X/tXUH+7AsUMi
7/OOr3ugILetySJzzkaYZEML1b0q2lxJSlf/qNyB5pGsTVb+DG1c1lR/3LKAjaNjpahcmSy3d2Q2
qOd3CY2+InVSDdAdkzo+sjcWUJ2l10keY8Bc+lfi2P5fMHkkEPOfWxcD2tUfgFC6tgLZXsHOVWs1
XQd9XOqws/V9wFc7RUSVT6owcctLYVgKUB5kp8ETNvGr6SkqWehQRWunlbbGzTlBbI4wpOnF62c/
gFWMGZ2ewRkxBIxOxjo6uE8uN6ypVYxfpamFJ/yVW1oyfisqIDdjdkB5CDamKfvazdR1McZqrECE
GAmeJTl7fW0MXA5G9ymIGw2mWJFYdh9ZlUI1HGkmVbbvbirUgl8ahxtGpOCOcaAH3UXB20CArW8+
SpH9I/a5HgieaKtgJgxurubXdVGhXZdoSc0aLCSsP9bqFHZz03IU0nsCz5vvHY3pk6f4RtHveZXS
5Hlctj9EGRjw7PX9r4CCG6/hiMCKjmSwiIwjSgNH/3rZubb7kPU+yWH2ujVaUqTDUh7Xl8PQvOQT
mE+JAzDadmZpPMCcemk5SrRa8p7IrgqLBigyxhsRo/U0z1MqJW2AnC7XsH08S7+WLhL1LboXLs7R
lFWJFyT5DcOu13BMuO89SVh/1+N4gKiv0UI5ttTuL9vz1/j71MWXxDtGFgm+fiCCgbox/Gs9m8F2
HLzOULptkenFZcO4dJNOc5gAf7woY42ujIJkPbsg3rni5WfEAx5wq2ePmm3ywIvQIsX7/kERC6Uq
vBpX+wVnuAJCxfzmvw+gLM7Sh4xixb9tu61m3iLf0A0zPcycR/YG5AkkAilKRn90VZNrqkgHmxMU
bBzTSYRaWu4g7G6bls4ysXZQHzfTuDDInxOh2NyEan3NdFfW8BrXjDPrvAPe95br1NFBmDu4EunZ
J9n+ivpxgVR4QQf4O0neh8bxInzCsh6r1dLWSJvTp0D5i2K847oBIfHOWDmHDCvBu+6XileqfQxG
keHR4zkEkZ0B3KD0sg45UiCMLwHpwjRP933vQ+GHO/hDT7dAVcsn1SS93NKUH/zU+Mzp1KRInc04
Tocgusy0CNQw8/hcxOYWQrgidH5h515jmS7sToL5Yw9i3iQ6x7IKT5iyQBM9p4LB8Y4kG/10BmZc
uWsMwzttkLNyD0sY3p7jeNhgeRQnxjHcqoM8Sl7G6MMdPPoY+KY9+JL0WpTLtXh7yyZnINsn4Toy
uxKq1/eOlmFIQFtI3ohyarq8vetCIZfytOTKNA4LEaoy28N1uqPqNOYE7Tf1gCD4p01CwBLkIajP
Ryn1vAdmcAuJYcmNTH+ZxVtSmRq+ELWjTjnVs1dNWhe1cjKBoSWdvU+Js87vHOBfSx7B07Y0uIAx
qfTw0idh8W8J6deJkqGvacHWho9PHeOTfn2Y3S8rQJfnhrSYmTor1eJc2DNDaJUiFJIKwW9GCLMj
XFSaIN+1ViXEFzs+HZMNSRW4Bx3fz9QqxelZjq7mJvDjIkxDZvReDhUT9ESMeaSb3wY4NajF95r9
Um4BH80RkjfQSHantVSe/j2DPbV0Wt1JWBRWPnA/R8k2ig4xzRjgOJ0OURrkTEfFqz8uyI+QiVjq
+Gampb3qkh/nHyDfXHVSj/sYM7sXsbiup2w5tH+NudInaeAlFstizPN759AHwRlc4A4uV6A46hWM
hk6M6Gxl8yysf9IOOZdAWLZVXI0cu631mSjZwCTki1LLQIYkfvIgZsaKk0+PdYYdkE6MUo2j/UGM
cXgpuBT127MbK/CB0H97wAiO+GRnmHk7BFP3MrwnH3Et6wbHySKC78K1tYxh2PDD7VdbGibIClKY
8LczUp+nASj6sprQGl/ZINd05xTe3LIlXp7pXBWvVHYyIMvJypkzkmQkp62RkAErB2rWJICht5W0
QeLuoQkx0//FXrcXmlY5g3hhGzLSlGo96lDmXcs5pFAQsem0qGe37ZUxWAaTprdPXlTFKHbTH7q4
TdndBea5DZkyUx4OjwafZ2ChJrtdWx5LuZYMhnsvoobyDMZob94UY5YE1g4QT/sjZl5FT6zdGm4J
Fct0qxJvPUlaZ7/OQpfr1kNHXoQfOsxX5Dv022CT/5oUl8/GsDdYJadtSZO6Z0N6T55gyaQZguWZ
2FUbgDInJq/5SP/+h5XJ6uR4kzQjOHDRMGl7MZ/xBdwmSeHwMkpXnwACWducSMHFHjYAyVQEyoUj
HZXs2MY+6ysmf0bhNUk5n6rcyIibT8AwUpXBnHYDOkuiMrOoFgg94g0zSn0ZDw6cRE3Iyu9rDCG1
KKvpzfbG4CunJJZLrpwHlpbIX2ZQwzh+RvrebcB9/uGUYfOt/+V1J0Pi2d7yyc6rbvIgeE7ax2pd
B6SOdCqBYIbJ3Qtj1+7+MU669do9YwqOVNNr6/RUvZZdRALWpWtbk8i3oktIc+lG2oH/l2KdLLMZ
kE765KUvAF5q87gnelejTppEYJYkp0MbIbyRfzpdLY1z41OL5+ioQsCiJwhGTX8mmGssW6BaXrGj
bYU81RATvS9HGCMXm7gXeUfDTPnEguxYsvxrNzsHFgGj0DmyHa8/JFj0b11PCIZGI3AsebCQnGWR
DdEosY1vh3Y8tAMR43gWQFWJxlGshUcPGMg0/kW6morM4JRhS6VNHaG7vVYJzM/Vx2MjdsauEeQs
IAgxW4xR4S8wvssuTEhJTqOQY+pRqe7giFkUNRvfp7/5WLx0qsNQtAU6QnzrLQlYSpDnfviq3Wi9
ffGHEdh1eZgGXtBbRyEa4PmffOMHYfV6sEPYXzv2tap6xhUy76Xaiet+lWyJ6HLnpiq9s26gs69Y
Zdi4iQm76E+X+zhTf++lVstJ+zN4w0buFRWzR9rRn7NwqSZcrPyOpZiNGQ5lePVvG5CKQl7AIY9Z
RMCmrZBGxpUcw5GDQW7x9QAAaUpj8iZHYnl0rzvUOvk9SaufqWC4okzDcjxftPLeBzXK4c8ygW2H
YVP6UIiGumbB4y6GmOXiQ/xptSAVC3JNZHAZOiKHjPzPLNZBjK4974klYXIr4QC3oOLS+Qb9cyl+
0/hhXsHkMSsKX+/01jxY0DWZX0tzojqeYcCIo+dYwvdMfh2Yz7Uc9Qdcn+0RRj3Z/lsf6j4t7dpZ
smntcgBsOfF4a61uCprY5ER+lTH9EAsLgwAWe7L7mG8NFqNyfHwvKmLBcQVjlLv7B22pJ+Gy87V6
jqOln5G18g5bM0ZCxzHMRmvWnaXMHste+0+ZVefTMs51sLT26X3JwXeEz2olDBtrWOWKejpnpGhV
FMGuyNT4S3vIFXtxSnvHmjBZ+lYLEAZdaU5Gy/miiVrz7ull5W9sLvqXv/JTl0MZUJNu9MmVCAKQ
YIXndrVklfqprQ1au081VM+FLGTJyvoLaqpIKCsjO4HhqdrMst6WRXC3UqYdywOri3MaVzV0wg5q
sYII/yuQYvT0QZGX60uajvJAJJSzZqiyosNm6gaD/7FsWnxHS0TasquToLgnOnP6qplmJTaFepYA
PQQizV3U88senRBtiAhfD8EJKEAT1qm/hUlc234YnXOisLhUalVxp8LhbEl4jW4n0Vr94KXN+jli
zcddlK38/QtLWMXeZzF/TT+GQxzNs6cJgfegSvDi4Kue1+SX8MaDXsuxl6sfEHBnxevR0UIpw1mc
zsjbdo/z1MnSU6i90HmyNNWSQY0itPh77zjFmgZ+ikoT8UbK4Bn+O4cBRNFsvEhTmKQm5N8s+1T7
hznGr9oI7/4LLQPUAFpIqR/MPdSgIe8i0DlDSpemvBf0bdn02NYiU499JRJIQ6KvSC1s0/yJGUh1
6F7RnnipW8Q1hmvLdAHYoR8nhh5j5mw+JzBRTCnMjhdempd0bPehaK0FAnHt75dh8mi62GeyMjlL
pigbhDho1VIemS1r5xyrYx3Twq9PcAdof4qrfKNd4Bs+16w+Q/j6aYwuxswwvvvOhwzqR981gTtM
fuMmIi3L/KPTSVWTWfITgaxkNzeDU6+4gsVEmCe9nbt+DvZqsDqkvh1dTEBTtU6iLDQ5AWaknWCf
Ib/WFjk5hqX62q/KiUcQjPcHG0cT9N9PXl51CL7olMH73zhWinKT0WijZ4360pBTOGLy7cDYbY4U
28tdbve7fEa0sBUUVsG6pKLq2Iz0kODiW+VRDKNwunpIQMdBCWR7R1BzEBnCn84uUw/LWD2GdHh0
1WxsBfw7F2mbG1dQXMByvBx33t5avqF18EvWKPc6Hsz63Df3yXI1HD5yUqppkYV8ilXa0rCUsZHH
uOhZJ7rrXnsegU9dmRngwFMhVNrsKddEVjYl15BGYfg7L7mA9kGweSDVCd6pNoVQEeq1KMCuBzvl
G6hqMOXOPiiAIa4MqmrM/0MYSlC1L+/LU2sH3Yx3FCIJSBVLxHHQvBu8N72wIiNI37V0ByIJLmQk
BXxguhV/NU4Rl4VONai1GLeT7F9EObg6YQy3pdnpftZ4ndqNPL437K/yCRYEcftJuN7yonAISQPM
flUK56R8BGKkjwMh/kg4iRb0i4UppMFHrcM51dmY+5JY+ZWfo2cl1EP4cCjdxG/aBd4lcJthvGUA
gSvcEjtbkvK/p4F25vTbko/Ac5I+19IrP+S7lECm9b+7eG0d19oAP0OngGQFuWY5xPl3+Br25850
pfhWT/Mys6YU3Ebm+QGkPTRigSd29xNgd5c0lEprhH9xx8iDeS9wk2oaKqIb3iVf14MmWxynO7PC
aDbNmqUs3dpXHVqG2FV8HBI9fFKGBllASvng7O/PDsgt9Ml638wZxCrVMUR1gcGN66wrY4EJXO+K
GI2GfbMQEpcYZhDSAwyUgIwq0bRbvw1v9JW/rn+2wiL/ZSKvS1YuMIh8/rjk6JWRreLulQecFHQ+
Bl1bPLDb/1FJh4mainHnkNj80OGFAXm53NfS6bnaZZtKT0YS6E5KzWou9DodgsZhcgM70oABLJMN
/HbfWky4jUlMha3boLwpdIdTuNJs0vCX/ynkoEgKlsEDv4O7KVGxhhUydJBE9BGkXQromImAlG1N
ilrfFaUmxQhkWPU5NcvtjVgkyBCA1WRY4ylYPT3uKKO1vWUKuzinxI2ZhzimoM2I02z4fn6a/pUb
rANQrNHY6GWszg31SxblaVYrcCC/REqfqNtymiWfBl9x3X5qvAxNi6iUaEHu1ooqJ/qRtZV795X/
dPz6hdbsBww4ThdrNpqkcUStqBUS/le+wmLGLz87CEOjFwjuRFAhfQTjaGJ+G9oGdl6Mc+pZVQW0
UuvhOoDwvNlL6ylTSzZBzL2e2HjfZD6Ysmzv/NLuow66JCC41xRAiBhH88BPJgjF8U7iD1nGWMY4
OgDNPmJ58a9B23fGt4Yjc3s9KqYer6rL6YinYgz6AW4WUbV0Dxla2NuNIq3K4DYITJmWTKFyEnfz
b8ueocMgpDnVIn/knqcZ1dCfE2eEzrk2YS22869SKDmS1BbBqQE99qV6TUMujnlh473rg9g1tDe1
0mVEq8zaEHIKXSe5xdqw5u3tLwkEUwH8T6WVlTvnhxSS32sS9rmKEKSYQFv2sTDrwBMC7AqK4LOn
+e/aLppVid7kJgj5l9UK2xiGosH09iqIdSaRX9Hmb+dWFsQATQpUWLopVp0AbFw82+TQu9PHM8oW
mGeSuy7JBPeya5wN6lQtwax97Pwfz7epuBC6rDSs00qQgFXs16lA5YimK2kaPZ4rv86T/2cLGY6W
jWRRBw4+cb6shSHfcTG0MMiDnVinRm/y9yw4OzGVs/jX04gpkAK9W6uuUKQLk2Kg11HkER6sV7KH
CgfmPS335Ze8qvxSEz0UJ7ddxESj2cmrmgJgInSjBTs2XegDRuz6Ptu/V22759tu6nb5ffzytdIY
9vsERXxoNPuW06D7ummlIpvEeB4IUtq2PCnb1ZCYnzOFYM9T1mPVdOPecRbncookXgCl3g3lxGwV
YoCpeYoiyhNpJMJgA3FHUa7t+UbClyiPSMU41VIjaH3QAtehk8FntDLUvVfXLIpbS6KZHTchkLiu
IQgwGH0TRGIm06HI5Rifap5awAur8a+iafMwtZHLY2NCTgmALbPR8bhEVVWz6XU62KDBsV8dXHI5
bJj7NYwJLMgmiQFzZmqvOhopJaq8r8So3MF2UK074tB0Wk6G29NJJHwLoHnt95Sm2JcsxUUGKItn
HsRGH9YujaW+FbPbqwipQSO5WADK9uhR2ZVpCTuugURX3ph7yU+1rvOHqXClP9TAwIg9rEjpDh7Y
Enx+iPsHYugyzmc0iLuZ3oFjEP9tsEb7yFvNkSLnyUUrGMkyoPlVYh90+/lk/2UtdQtaTrYTJvNc
4TsCz6OI0JXVNKOJ4U77cDSrTYV4hM9cBVXBtTFCt/mA3TKermUPbpdxaEMA2nUOrDxlbA1TZdwp
rjevbFgBZxTyLS7iy5oWR4rr84KNJiRFMhIw5eC8gmHWEEm27cp39ZEHpbD8FUFp83wv2VC3uczx
C+gefuPwj7VmAIuVG+QMF0tYKx44/ZKLHtAl1PNmiSeODbOTuVpJbtH0/1farZwTNz9Q2phIaVYC
UM0PARG/E6/cHuxSRSfPpDGXOboh9GcUWYsiJ78eGWew4VGiihzXok6EmnP5TTskTNgokmHs0mSB
qhUe3S85T4mdAdTKVNXwqAopPbu9TiBHIKKtGk3ktzG3wjZO+WxN7ZUxnDdUIf4ARBHENArwkJJ+
UTyRwJ7LUTQ5fQb1Xt9J2mHW8sJOmLPCGbgRIk2bV6MfCBeVThjAV55eEFTnA7ZOFEQmu+2zO/N1
Pr7ke6C6hmlwkdxw12VSZ5M/Ur5CNvSxYXTZ0+8Ql/mdjxeuPNUjdsfz3B34yMP4+eI0uOcpDNne
EODKCbWybp3blXyF0KNmCXESVYVpczHZRRtRKbjretxA1IxGqlbOcpA4qwsC2PJ/FRW++CuBAWyb
fVzS2dRIok58QWA1tLLM1Hb9FKd9wkFd3riBVsiZ3m8Qn5l3kWuGkOhDDsuwJOyazb44TsdrLRrX
9Gf/rp0Skv43U05NRnAHSZbWAYPRw2p8r/bpGaJ5WouZzXCwyEKYPp/o9z+9+vodyuOkbYFtGIAD
2gOuE3uLsePlFyqa5ar3CA2tlNQ5AVqrZ9Rz4GbkkKxHZSiX/Emfue+NA5iD81PA5QwIbHXFQFa9
mjDanY+p9BKysb0quVqP0Rix/Qh0OeEopFjDBsnR/1AvRlQrXx9r3ocWWn8dePpPgK0IeItqIz6D
MHTYQY8aMler+91F9j096k6F0K1KsOnTQlG8LEPjeyAZK/zlpi9w4qih1uZ54mOZsMdk85GxWkOe
JzS+WZf6zvH65z20x2clLKhY9Cg7aE0egXOcN7RwIU/YFIqbSFZlbARCOJCNkRVkFNyEsn4mDlAU
bzu3AoqtRsqubdK/DsZG5s/FIHBYrN813JE/1lXrmbeKqm6ICgHZaBAmL1UoGNxq/1RGL9IggDq+
GQM4OAeuNvPYytPMXm0Nk/r+VbYa0WiL3IWnnhq16k9fjbT90KJBPzn7Df6O6/33ie2wny8+UDSR
ja5wp2EjlS/s0jvoPbJ9Y5zO2i+ZCwxmS6txglIUFqCzR4/HOHDzhX4rb4nUav/lwpSfkKE/wRv4
f+FC5iPPCLIlpBzi90evrSqQcxAZsuWMwdIgSs5ikbpWkzX1kQCWsGxmM5CUPF0LesESg55nnNwA
70kTxoH+8TOd9Rwx4wfLLK52zPV8mi164n0CDCFxvBkiGgYoatnIhnFwGdAyz7Uf/RzM58PFz+dV
M5ZcMhgmJCC+KhhotAOiZbM3SDIKVXUhlfhcBMGR/k3G5QquzXcn/bIOv8fzcOJfZqPDbcfrizY2
U74lgmGPcjpWc6Dk3sF5tQcdrduqIdot3LFDo/skMHphC0jT8UIBIFdoxIFSHWwl7rhaFGXtzl3H
q39pVW2Ez21mg9FEGESev/j4nAK4gR5zlqpKp1j71DTO9h00/yJoFGGyPI2tqTTW9ltSw5llxSLs
h/lFqMmreqYYBYUhTtyrCZalnLLguYlUsfm/k84mGJZDJJ8pBmd2NfociT6NNqFZgABElGaZtIqb
AWTYlUAGQHoO1P8h42gsmIJMETDweJlo0Ma59sqq6pRHlppzO6mU36oaERdL15Brn0MTJlfQZpKF
fl+g35+Zl/tWzMXzL6wCzUPplqRUVNlfjTJzSuuC6GXb+qvcrbgrZacSRW4eqnjwEaHLMeiAgd6X
lwltcNtv/n+6C6SKLGlPsj2opTzRXP/0Z9RvbKrwJszOfbkhKVRAm5NDmt/mkmk1Mv7mU1dWvFVl
Prh3sn65BY0o3xhrHanqli66R4SrVW24AS/O/Fz3Tl8t08WPXwAwen9waCcam55DtPK8eCTU0SU/
nlgE9fYG/sdCVRVMDtAEcGUxxocrxRitakJIHTh9lP8t89CQ0SXaE7wa948MZgiJ1fSoRq/5pRBc
2np9caZTImRyFVFcHwwZZXswaydLhWkegSUmIEBbwLbSVx9CPE5L3guuhL3Ijj+KM6b1nWuTzoon
cf4H24IiLNAuda4v7t5x8RRrSm5M5za9TA44a6JWZVLK9hebtKxj4ZKHOLhDZiZ3CZfrW5JiPnGm
c8VUsYmhvN20fUVo1bpi5v5nB84OzldWk9LfdQJCql9GZUiw+21qPgc/SVpTnmhNhEWiDzz7bp0p
21hcF+oLzQaic8ycVAiPv4QTVX+WBv3maM1Yg5YZYVzjDkGqNAHjvku/Xo1w7mSS8rLfrGMhRfkH
l78v32P371K7qVaxnM5qUDFvVCXuQD5JhncjbJRWPMz8B6dFPwHBZGZMqtR2Qtyo8lmq+81to56t
Bt6EbJK4wzyKpiZ2uBtWohwQMLEJHvRLtE65Kj50ddjiMg1HofIeT0blSBvwQlBhhx32Fk5/YK/4
YjVsHN+BMDsBl18t3vDM+7PTQVmhx9g5FSz1hKno9kPEYvcYK63dmLYWwU/1GEjzKrCHXPxiD80N
RVD2RwkKimQx43x6chgwGoiMKo5Mt/myCvJxAefmZpP3oLkIn+KA+ZNp7DbXbi1qDob3ssFHiBLW
FxcaIDhYGIEtK74x1rwa+9BNoZldv2Xtdr2gpFXw3xlwqV1LWHbRD9o4fZAB/hBpQpe24xASOPXu
PmjHchmOEozWiILMVaPzL6SXw7DQf1PaMbT9e0Lo3NBnESNb8MZtt+OW9msTD1LErAFfXpBEWiYv
AQdpfU0gJ8xGJmegDO6zi5sxe3MQmFgCYjglj3XSRj0NO1T9mnyHrdbK/tShJk9x/c0LORrWb8De
8xbpfmLEtvE+Lw98u0E3LInjEYo7FsaaQ+A/rlUnBAOc7QBULEVB8u/M6tk6p/OAxI4ucdXsAsD+
b2z7PiP2A/A3ywWMPtJ9IgDnl0A/1uBSXHX5dIp6VxfFkksEABNzBwklYSg33SbRC1OhAWi71XS9
TeTUwI7pg5CUbQYNRUTgGNOY+Xi6Ok/lFvV/yLJMw1zEYJr02Uo+ha7kH3q65JU4wRREvCOHE/XT
cyDoUTXuj+jWpVtDa15dUlrJrIU+VYsUi0ttFVTTCro9ganReqNKuNxvPPs5tzueZMkL4lx13K5C
eluieFGa/jvlI1eGIN5Psbk/DJ0YlFY7CE6o9HuDuYYTlCRQYl2Bue+kMb1EXJv5w4ZEMmkaq2FG
Zr3Wcm7ve2/iyoc9Ws5uvL/trWHld84dJ8rtei9i7eg3q6d6Lv9dd6TFGhEUzPzHFfXCTkkQWqV9
999aGWoxC1GTq28z4U9WEwYptE5V4EWTCLmjaIWMahdFSLCd+4opcF+XYU9YbCJoOY36oHDlmxXP
431mq091l+J61dAJMzPjDXihvHs8cHcjp0NHJDeA8EmPG1DhH6kBxbllPk7rYvAxJZTVZzMyWYND
e/UyvRNp5d9uF8+YXAXi+wg9UeoxegP6J5NdZAbVF8/0+I9wYAz2Qx0ls4Pe/pnHX6EoFnAQELLL
12BGxjV6Vaza0w+YcxsMIOHdDvNAmn0FIB2vxHeu1a8/+9zLOfPoAI8j1P7JHnYCbUOzOt8FUfC2
fC3qGrtaZbrhqeWKOwXt11bf7TfR9eZMJkpJbW0vrit6JIH4olCV7yil4uCwk+mKxbf3/djugtez
IMdhObCUPHHXC3tM6WmI6D+wWN17C91pj/znIw+S5YmNgnhG+GOmEVw8/acMWQO0YtF7WhoXET0W
Y7dT/+/we/a9XqbnL1nfqlCnP2pdeEPVz7VJs+Ywvc3q30+6Gris+B8YIssshLBCv1dufX8UpPj0
vVImPurOz/Gh3GzApkVrYDuDATpK9Mkv2nYlHBzpEX/BqtnZzxiBtGWR8XoQH0ahitYcUD5ecv+x
YZA8as9826CRO5rPyy+cp5+n6XASF9supZI0PUJ3yicLsqEVKx69aSq+Z6maqankMnE/HdXyi5V7
/Je9vmPHA2UdSFVMwH7oLiAIKYV0WaGbj154MTGOdFTKBz3UmSJcIwoG11J/b402Zturoy6qjMTN
TxBi2pV4snirgRhVhl+Rp6pNlrD/ziNK9x0y0rPd1a1X7jqV4IVm6zCl1+Gl0Cu0SFY0WRMTzuGb
tQnIVhbj74MPrjsYY3O1c5+zatGhR1UZQtpiadt1P+JXCNTzIAyr5idoEmWWgtVS8c6YNYEtEq5V
W8TLS2guf3v2he+q7T+34XrkZ73blHOj35vXt7evbkwBg+nFTOIiCuh7utQdTQL9coZl5a2vLwYT
hfwksIl51g7JK//iE29hwP3HNqmKYUfioNTIL5tpGqRPrFrREfIjwG5jKfhF/vbTpbQGdi8ekByx
26eXymYzlf92jeDX8jqUc0CWMOpAynnbp6MN5DqNvh2Cb1YjaY8K7CyK6kATHDhjva/ZRhK+3jKY
lvhPgNMAZj1mjVnweIqZZVMNfSSuGp1BIG8TKy7p1bpVoTiVqq/GeTrDWaAV6cP5J97NxMLY4X0I
DRBkRbEuDFWhSbzsKzh5036KJPXu8IigQ4uuJwGysm+Mhe/gWHUExQ7YsshJ3V0jq7bKbqjOX/g7
S6WSlUN3loqS+fdCeLF3NJqHVt9VV35B2bSSs9pwUNFlMAdTLysEm9GJJ8cPRS7dr9fh39g3iqG4
GTh2dR8hU6XXOjWnX3sauW62++OFZsfjNQtiEwdVIFRpuL7IzMdhCbeWidcfskmqSq1x8x1BR/+u
OxNGjGNE+e1+COlT9KbYo0D6S49uQTMLdrWDznYvuUGsF0xGm+WCEuXS6mCvEl7zc8LcplbvDXKw
XmcwP5LSCS0Z+X35ftwnEkwScH49A86RTY4PBikrJDWHTFt2lbylnDVtMDvu5MVQAKZn4B/MSeiK
PO1p0U9V0LtDvjxSBHM80N0GsFo8v8t5rzGGFqBh/da7lbIaKUqhmj1WizMwKywYOfz8BpYegZF5
4bHntlD5NM8hcIECO5bmYKz7IWi/HLeZSlFDnCk+CYvEbF8PGIfsh7lVeqv0pXD9Z+m2bihd0piI
8vJdxR1ZvrjuDDM35lbDxMckHDHxFp3bLVdXbRotJeHMpHXD0K9dFpGIwtGfvVoauk0jVCtXxzjX
AF7CsbfvOnMHe1UGZ6sIT7TkT7pPsYqtlpvLZOJcx2yLvnfjxShOtt/1KXh2KVumV8opzGMmbMKq
XM34rlnmukfTW8aHhc9RRvY1L6LfZh9NTq82/vhW4PC6jdqA2wcqQo7da/1nlr9+JHWCIw80Ba0b
UY+Sb+oZqHTL+oIk1gT78ntwTg3xiAqSrY3GuNqMUnMmQkmhYyAx6SyzYZuorGZmTkOwpt9y+z70
oV9HJBOw4B8iht/kIiRoczM8f7oSFG1HrH9/u6Ya+uX6O3J09QWXyNdt3CXV6vKdtSw/Fe2yXinb
VzITa9AsFKuPMe4wzIohWYnuEMH7MggmrClEAdcSiUU34IXtFlQYvosT5Uk0JxGfC/e6JucnGPdx
9iZCoGFDWV9V3thEP/od/wMJ/O6T1rNkRb9Z8hwBv2DDK3hVxq0H0/B7IBv821x7h5Kuv2BkYumv
WBzlyJnG4YFXiILbRiTVkCB9DOVB/tsqy8Fv1Guwo39Af6xEVt9Yxsjfn4igVRzk15gCfCsPKpEa
rQ5G3E4EwthOa1p4WQjp/lgteZJPO7TGlwfBmqwXvxfis/wmmWCIvVpKQDmNHBQrbFhRkkISq5Lv
xAV9+n12A6WAyDSPpXOeVmHJ5O49lzNCdxjAMxM/paUKl83JtYOkT5FSgB1Si1c961fbBmVnP22Q
S08JRjvxCGC8AOGRvLO8sxBchDqFpJ250EfBlnxky+QYRh03ul5qr+IUDUqrmEDpjJtSqwNdLHJA
dD6Y+D72IujblbhT0mX13wK9zivsvMyhgTqEuX81jdms+whXWVoT+iXJR3TgWVSNv9xhG/9yi7QZ
5Aj8ZNXuFIcufphMSB5F51U01REvE42hDja20a2bs04D4d5dldGM2Pz+ugwmHMD6oXttymQeKtp/
bPTNmf8mvj328KUNnXo5cy8I6WEU9Y592eGMtVB4wbPwCDPyQYBbTmiLzAv+jgcys1isWXR72D0N
qXESjI6zv6dGFD26/gSAeA5nSbFltjTvElmVyXkwLMUVkSpVWUB8WK965ggTnGALqo8FBxborfDU
UBp3GRkNxOXZR2yaiFnH2DUu/u0rf6ZTybsT/qBWqPvkmEz7XDXxFIZD+s+L8p84nTb8mBbrTiaS
0bqNAM8pQ81VRK0CFNRwECHkm40+3p+njBzevQMAW/isbHynslSsteo2Sua/M+gLEJFqxprcu65K
exFCzdcfcSy8DAoa/s1hfIHqQdzT4G9qQddqdRsXtW84HJBu1ZLoELjsb6aiwfCyWDaTd2498BU7
8FUePpG+CI1uYSrNs2xq807DsaBeN+wGslyXEepCeTzwrXIluf70g7JVqQdPLa7lhJWYaAjgmVop
khuNRxrTm905WMUQg62dNbjEHSrr+wiEGrwXK4+VMUN5ku10ZPGcJTPC3LXBtChby9tUmISSsulZ
xWcNj+YQnc+TaH041CEnnj0Uv2prVjecrPEiLq9CDIvvR+9QIQWsj+yg5a220pSjWoNRHw+x8ypK
S5Qmv+ExRpGEfmeNN44ab7rm4jfvAg0Dpb6mU5C111oivfWOUl3vMGLuRXoIir2velfYQrmXGxN6
GcSqxDpiJZw4ljT1bqIqo8LRQfS+OTNpSSokquVzU8HjJo95Gjjcw1tA8qOcw6W9a5TdvnlxZ4rP
nIIvdFsAV6g66fDz7d3ndPny/+PfuKWuLjzDWibbCOQ6AHDHbI9VreyhC2SHVlpLhMUAWAPEBjkB
uz3CbcQQjTY6i9kTI9UL5USCZH4VCYa2k0qyQ0USnj3xFzmtfBqoBUfyOhQAk6juVGjzEGbl5C7A
dfQnTuYQWYTceHBdvZj+rxkGOpnV/4yXgdaNKP3eMGrN1hQofw2E8SbA1pQpkDzE94CyYcnzYx4q
8h0Lqmse4J8fYmDViQ6x647ikXPpWWjk7OfKAeHJH2aeaRCCCoFYoUkBq6/l9XOXlPPNHukJREG0
1fL8UvvbQCOoKB1EEd2Wg3w44DmMay9Oo5K05Km3nrbBumndSZbD86bkItang3A2bk53c++mKKGr
zEHTfEQ7pxm3UJ1LOcgNKQnpOGjbB0y4XMDUFoVEsOHx+LS3hrreZsXeIjBCEggrG7eBaopSSwvu
iPQs/VPyiG8V35JzfxGGpddDKVvTyd+8J3YUyJFJS2szBJGnsO6+B9H/DqjvDgZMT0KbmbMZQzpb
0V9HuZxd2mmUEO2Lr4BK50ROybY9Ya5EXo9l5r0RH2WhURWjB4rudtyjJQuCjriA0iuyegebguag
Aw+wxlzQZ5cI46+U0RBrwrXaVczggv3XcW7cMxEwTzdCnktfaf6E0Qw2MV60/LhcaWn+ZxWmPK+L
4jL/0ul/rdMNhb3b149h457cuqHXURHU2ZrvLKduhA4eo/4klyoCEb6KaqHFgrTwWOtBnC6zO69a
M9ANV8g0oRb39F12FXFDmMkwOCgbvqgKAU67bKc2Lx98Bg9ULdLJYpWCyGVNQOvb6lNjlKWbUSV+
yZu8sqdBiyepVvAhZKpCTN1f8XT5UIZ4mD05+Vpoh+es3u4Wo381CPIteGogQrWltIPU/1+Apmp0
4ELZjcJ7qwsrtbTXLOUiLkJA1a4viJq91J7Qzb1jyCmLb3lVvjD+og0qI9f+6pUU+KxoFfMhCNr3
NBtGyWoNUNpaK9MehJh8WnYY7KlxFjSjGmsnQUe6aYhQrfc5feE/17Uy4skzRESLg+fBilUdKxAG
d/RmJekJaT9HSWroxt1CanwWSJk2qLXfJ+tcQOkvdkKyCFnaQasdXIxgF92yleUcBfWa6UJEPEWJ
xhjjVGu92pqIGRcsYUq46U8oS0g3+DmOaHNqJFF4hAW7w4o9uqWYuNQ9GlKVSJ1osRgDmoefL0j8
6tJ8xzs1VxbBoIxLoKe0e/M61VpOeCAhKACNFSysyxjAzJtNM/j/Y7mF6P367Pmra8jxVVw/t9Z7
KG5vMoA4rPwqDQiq1J4PeGuS1XxaY7uf3muUZruz8BqsrnMr38wkS5ApjRf3wyYy/Pm0/e2NSMw6
vFdzkK8t/LbpDa1ItzFjPzGBrWhRoGZ0dc3tFfMiMs79SSuaHbcSLsm7bIXE9jWFszU8LY4SGmPf
v95NG7bHxgfWZ7fQ46+CFkU0odHVTU9FO7KDBXvPvmVbNTEMTOpKtloSiy56Yy9UaVcNC4stcsxk
JdNiuvRyFRrvjwr+KHoKGh3d8NoHruWxEsdjG83whCv3M2ukCFi+fHGEkfkMD0H0YKmeb6qb8KcA
kJO0xHLqAbNhwWDdekj8Qp2fZFymLtQC0Ses+dbWUZomK8n87ehi9kQXCYaoIG5Y9ckKh7daN52o
46nQIvLz3PFuLq6Nos02oPmbyasrvS6fy8o7UoDFWncrToT9ex9BCzECzjQJcDxZUFFzu8QfXKMs
jp3s/Z6/r22haCXWoC6SjAdeuCUiaOPuhFMgFpGnNNXsn7KpyhE/xHvd5tm8eUA5NvEvGbPWiw01
ooFS9kYeUks54QY7BHpWmwU7Kak/BtCziXQqmDwddefw51ZHTZmSaDJ3ynpxduNVUpkyP9eof+6+
kcTr08tcOk5RObHXOMI32BsLuOz9C4dvK8a6KH9gruh9VGt/KKb7gZf3OKmK/GSdUnQgpnQ+jUdg
36zNXulDcavsfSIYU0PCE6XAhYs1hEzR1uUSzVbhUJepssa/3AIRpsWK5hTN//OQTm4wv0DEi3P5
K4sXTF0wPgPt+PW1PF90O8j77YEE8sx9BggyOgHZmX6yRy9jBrf//a0nyT8UFnV2YedQDWy/eThd
4WBM7UjT4T/XsReVGyPj6UZUnyLDpCmLVWQKKA045Zsx9VmNx4KitRbbnKCC/ZjUIrEdhazwBCEY
8n0P7DC+/NGCG56aGR4MDzTshRaVplwini4PDLeSqXLbKzExYKg7KVXTB4Ho3BTYfKKP9PiBiAgb
U8xY4azmGxzGeEJwgtn/s2juFYu5QUjLI7S4LLgOPgr5fsJlHhMZGR7wmcSzSbmsJOEx/s8eex7U
m/IR1G5ygyRY6neKqudXgZ5HbjNE/x8UH7NUBUewOST39xsSoHWIU1/FlDqe1GJcQ2C0S/+xsrFY
m9sNOk6QUYwZz3xHydVWD1CaEMBYg1v95W08SAj9bLBZ4l9tf2fo2YAJWxhn47ibSpYJczGmmCB6
5o68iHrBXQJFyPTjCB/YmQ1hP6aquYzUMB+j/9bFfOPiZUHZD4MDMM7xDH4GrsPWdnUli/ryunag
ePnM8/tVFelfDTWOS8AHjHdzYCTSs911H58BqNSyFstkU4CZqJWhvW3TdWoL7UoQZQUeH0tPXN9x
RIiKNAuJqn9ueF08/zu/JYnLnay+rsJLcG2+ABrjCrjwXF+xSD5KzRahmwDRgSGBMct5nynyPYiV
J8vbwCW2MkVNVmpt/1uhhrYH5sRDbHHlDjon5lHyAXpoGLO1rdS0TcBspXBNUM6ELRrLCAJMc/0t
GPCSsKE1U8bIfFicpVsEdydSstl6P7rVjDgglIGhWYXewITfwJ2OexqPR/1dBfxYq/CpdS4o8sxC
/cGEzslQ1yHTP4cGJoyuZCFJ9OCZ6ACGAXsLM0caNUe0U3c6sMq+7BZinTF9KBONchAdoKolaVY4
3/Uq9V2tI5Jb0X1LJvaQWnO4KWnUm81zM1pKT1HuBfrllWAxvn4chRGyeRvxMiI2e90swtKzl7Z4
INBflCHYzkZu9eZ3fiaUqCXBbqBUspno8gKsrnUgXURC7LfdkqmwyWIDQRFhilRpHaFUern8UtC0
Le9RTsq9kebmtcrUEEzXrL5w0qWwXEZcyRMyO48OFa3MJfocXPq8jQJq7eet9ECYJ4VcHlV6rftE
nv63qwZGCVjW0Zrge2Lo/DQofLhocg5kOd8lm6yDVRBT8CQbMnwT+pRVIYNJcthY25sMOqs1TlWW
nm2uoyl2Ak8AoFknI0WvuJeSVo+qg1t0PfwmLlksI10xjTpKb2jvtMUtcV0MhQTdVuy62Q3TocjP
Reze/dhUs3vS0nS3UuqAePPGRDdnlmb4Z2WJppKMYcoRek18WyDP+oE3p3K4xf07l/b20YUj02EA
MIxm+odjM4cub2DoTy8CQCQndodMGRuO3IayjCihMI3QJeUbb7LcTHmGW/uEW5Io+RbUh5YQrMsa
oXc8zAbxYWpuyMXgpPvD8pThKUpr9lYB/tZsiWKAs2PU1KPrAA8JJ+2luyqE2enoaUzpJ+hbOQQn
TFPXulfMLy9XyFzOrHuXtLSk/Ll8qaFqwGUcjgaUGOLE8+BWGD6w0loKU9NZCwbgUvUjSIe91b9W
ibhs8fSZCJ2U+xRHJY7ImNJrZgx1V7AMuwIGgiGJChGRYSzUPlQchVhPeptkNlz2vZxVL5OCF/ZN
S2dGTZbl/LBN5zWcG8tR+xQTdnufT7VHrLRLczSQlybO2Rby3HK8/2+E4u2d21b8ELxLSglrlNGt
XIJacD+LRq6U45T4aKQ64uUgIX5px7YBJXvie5xc5J47/R4V8vBA9zdktTegFOrRpIwGiWPDuIXh
5ypnWho2NbreQkBuW1DaZ3UmoGHtYk9QgH9NEN3Vi3OFhb44XHadUsTwOt3wHPMU6c5NJ+RoSIw+
O5hk9y7atUas6xU1ACHZhQlXNlBqFA4dZBCDvSx6+dMfc4QgZblFdu3PVGFBYf+RRzdMItiiMQ24
cqtQ11R/k1PYW1q/yTBp6qes/L+yos2tWdz8fj3roVQyUqyJkY9LZtLdt5ZDflsMEcf0hDX+ZeKX
1JXfEEKUh+p28fButuumjF5c1YN2vnt7OF0n97ZLa6nD4EIUsDzF1RHHtAlf+luIXW/VrhMdrXpz
y4exM8v0hZKAVZvmln3xH4KBaZiI3WRCkPxnSOaoVZkBB29w66S41Y5NwEySgegJY9LJjjaR/0NO
m9WiqaJ2K7NoRYxAFDtk6K/VfiiG6619foXrZmzi7JGvjAQrSWeEsrDQtX7pIm1kz+dlctP9I+80
zX+mADAzW8LkizvQzJCiOD97aZQqiNDu+aYsEZ86hxNZ73fCojICSaeUuIaFiJ1g0aGsNCi1ht1E
YlNby+ZeKiIB+urMxgTJFTgQcclbH8XbRP7rggOfi3GvJZnDwXPaeoB7q5seIHHw2ntMuE3pCzo+
21/jaEES6bN/+hGQqxesMz39idB+aNvFJWmP/admcUXbjGbb8nXldIftvi9YUltpYRsFVCpsvgb0
xdTSI0GXWmU1Awo9L+pjfBE8TXVcn2qDmoEZCWWlgC9U9aqbqiefORTGvV6SNOHTj+JihsTz/rxs
OWUpKernakLuHGjeOWvQHxtbrNJ2eLvWdh8t49o9T5CkEXNG4OJF+jDnsLQa1+185GNWQOKoVKSd
FqRqQkA7Zd9X9WnDCmhNFgm2LCI9CHzE+hLo5cDvCfhbtFvpjkbeVwsTjq6E78bDNBDf+uSIqO+l
5oUk26qWwN10ruPlH/a8TGkT0KKzeGVcu9mzOC+LA+Q20SsdCBLobSaYrKA1DA4weNLMzaAWxhQK
Q1Kb6YKoXFEw76OyETIX/FmnMwQ92Xy9apICByQf+zmFK+fqPQzxxlDxMhskY2L++3tWOvHdfGKa
f4kruLgjCXV5AH46fqL+3Yx6iUOrRd0Y0j/YhBoQUdXTZoAZKDdXaMrgzcg5XZZfbAWcyCvSUnO8
PYvEGPf8MUb1wiznOtpNIxlOrPJna5FtEEwiy6A8QEC2qBAyBgXe3JGXmHaeHC4y+MzvaphvuRn9
yHtrCeSHJgw6E1wsnjZRokIXFqbxZo3uIPfcRVAlsI1ufmgTFBLXrROjqGJXhYp1YsEJLMUJ2RVk
Oq58KJYOicgI9V1XV3haNoimaSRSsXxwyLkEIYOdqrCB8PyKCnD8aMqqfARYD+FiTxb6hxL2Intj
AWeTN3/7eQxc7grw46VjiQO7EC/n1A/qzlyeCSaEx4O6oOeG8HJz1xE9kCwblC1OofGtf8gEx90h
lsKbSqFYWaO5OHSqwXLEp/LMgqwpsVJo/UVBfpu9JAO3qXoSaOB/SdIBu6GrdxojNtkI/hZtCjJs
JKfQsfoXBcHyA5MnZ3ZhUbxBI5dJJu58+y8Iw9q/YvILwo0a8ES6jcueOjKtw353IgEMccF6W6VG
IIVHKdQLoRKYQuvadJUP21nI3vN9ku8rpao6sKrIRzVzw3+YlWsmRt0xHjKp9iI04wa12YNB/OeK
bEK66KHJPC6VUCM6aQjlyoFYgo3oX+0of1q4YuNWaBM1E9hto9E7GbGMA0cCzfRIEVZm8G5bPnv8
zLXJ5hc0I/PtFh0Zxor3n3eNCjLR3EgzXCHvfd5JUT5O7URHlSb7o2IaMv+fkHQXmiHbAvJZCcDP
CfpCaLlECfNSBec9/SIZH+PeuDN/LfNL0ENmv5p6FUGRs5YYrbN//3MdUTxCmtxw7YJaDXaacXP8
s+7Gpicq31da0Zyw6elYriOl0OBGOsxiO2GcWEndyDqICi8ktkIHDzx+xQqyosHywe6zmUc3ZXH2
HWYc9vw8rlrXbOBfg27296ybQntKSIYoKMlRZmb2/f9HdYXuw42CoFfZAm1kvUubBy8f55ZY3xhr
q0c6BfgZCigLKU0W+mn4bzoubzKPtYe5m9I7csD1wONEP5EUnawwXCJzOQuWdzAte01ZnTHwlKkD
2RnQOSYz9miyaAB2oxyObOa24c7GgfXr1vN0lm79mhp4QNoBKRuAqK4qhgKBFCW+IqX6JQwUpuot
U8a0s4FePR7iUBxwOby9MHHDip9vgta0v2EazLxQxYTtAazBZROOOxbHbOnJ+sT4cjS5bmHphDM1
ydrbqoS9ICJ8hw8IvK0klNbJxy2R5RrmGEqpF6OQjYcVb4hsG+gMqqn1J2yny9Lz6NYkMnzVIxM9
PSRKOHu5gZ6+mIkVVyO7PXQ52m7hJ9UFpJ8rZ48sl8zgkF+bqoKvXOJoUMkAJIFX6qdpErKdyRrw
CRy+OCVNtk77lrpWbSNuI82fVZ3/uE3RO4rYK0ZikfWllIqO3VqeY3MJeahPjqRWx388lCun8vRl
HyQu7Vj6oQitWr/AqGPTLgLJCguenOIpWKtD8+L56mnHYqAwUNDYlzKRlwJ2siPYr6hB0UwOki9U
V0ZU30rN2dbv5imqzVmeoSR6wCz64Q3KQD6y4Ltxxn3rQUi4u5E8pvbDEnc4PLhPl20LjWmSWyqO
5VptxKZmHxOcNfYcDTX0LZG7QFBAhZE8VQoKMk7CdMPsHC7O8ajzpzHyMMluvEuWQYXH3KuNql2W
FH48ppSOeaymc+VNDA+z6UpbNtrHEbwEKr+gDgjlmSwXUjyjIzPJ6jyq8yseMsvYGatHFx6m57pM
KprxKEo02wdM5G37LDS6NBUvwH595irDWtJlaSBHG6By7BwBR5j9PHtdUN8qxxAKlVL55lYYJIXY
ObxIY9Y+jrng+CY6wWas0rxcSmpNvWcBTn88nR7P0Uv6mrR7c84C9lds2JPaTYQVfvNVsq+CTWnd
rbhFLir6UXtgwwcr7/mYlunREupdK+99U0zDpgiP07o99cjk78LfRI+DPSNe/XB2naapv629QZ20
7zfA8B585/s6sntxAWheT5Uvs2YT7iKG22FOfs7/89BaFac2lPqmDuM9LMzGJcEsWE9fM5AHmTJv
DXJ5EPwaf9wE5xcJ84WavcvhNOireP3ewXwsh1DspkjoyQDdAnHJaw+TKJ1+cQULt8bKMwGGtu4N
TE0ApKQNdiCuZdkc8Iip4VNKynHKYqu/sSDfJIlz1sd5hJ1f+NHa7VCYhw/7GMdPkzM1LWtSCpWx
TH91JELR/I+7pzexKKWOAu0UcbDDCxdmcBdi8FJM98ZjYXJ4JkXGdzR3ZNyYWw1eKaoZ5CnNP9wk
/0iF6nS27HC/+qBhpLWt63yGMnSeWuK7X2kXqkzW90S8fGNdPXuAahYdx8zyMX3cJFxNDON7YDE9
ZAcuW+c2Jgh+jH4yjhrlGogIYlIFqh2zbZz42+r91kn2Zyh4wDp0NL1emYnWCio9423NqfGZDmsP
gEav5HqxGmrB0W1ZYAx0W9vwzEhjAjWJpL8ehK5jFSgDslUnFhWwkxFoQUW8KPi3mnI4JatBH8qX
vxk0Jm99IPtAlK9vYZ59JYrEPz8mf1gQx56leVBLZHB5PyrUusA8GaP3FZAO3sATZGyUAJE/CQCB
V+LNUmJS9jj3FbKOoUaA5BjjvyLrDDBJFBM83/rUfIjblujdk2EPXuwAQDety2qAFqcT52aeJLs2
fhqwlO7rGHBq61TBh+MA6EHxshQSQi37VcRDbYbb+0Bk44hOMx3k0I5KffYX4W4/+gsUzLHB3hvu
MVvmlLKWo4vNyb9nu50W3pHeSo3MOgR9HNrP2EYHdAGE8tVV/AggMMXdwP7o3pVHyWCMAE3nSUpq
sDCLKmhx81PfFhLgZFjDrkXmm8WV8uRqH/dwpT3UPO10VdNetVt9FrDoEX9w4bnh7pBshTkwKWcH
frbjG2jeFrxeV6vGzroUdIwQYEPxmzqSyWil69PonwsLlBiXNJ/N2JSeACsz078OqLmvxGKpgF2G
995x4ZIC1JewfWmWk0U1Gk+eFFgux+hDRRQO6e045gZhQLHknx1OOSgI7BHcPEzB8NsqBqWCALT9
69bddhAVpaj1bN953awN2i/XVr6fL6YMN8WDaZgLRAYQXbg6yUzeFahKmkza5PZyfTl2kwS2F/0h
Uam4NexT4tkr33K/qE9+OsF3HfyHzXSt4zISm3U5V2nY6NwQ5pkYCKJzZHIO1HoO1T1MXFC/cGJY
1p1Y1rGEnayfiLxrDE482zx+eBj4xbUdJpz7NidqV7jBuNNd/5lpFEbM6t3sm07zbw4m/g/2arHB
j5ZrSNkOZxGdZfCH296y5mVMMWPtQHhxOuE78MagcPVqhGyV8twip2vJnzqN8YkO0ozaErYxC4EW
z5KGAyjoqZCyT+3650mHcVW1k8oE0+b2zCZ9aGPyZ0lbzV+FBcDY1u52R7olK1aBZ/1ECxOeLYoa
wGytWYym68o341LpArcwwcbRvmXFaiUq81LeQAcPC/EPz6Ugmkqj/LysrTVIUResqerqoESONv14
KZFRVZ5buaAIf7oOA3tNpSspnoYvbdr8iRBEccvqOdnBry019qhLf4iUxjUKN26Jn3w+yZ0JTCpy
Cp9T5KRTGkyAzCt16g6DnyWmCK5iKIBlJC4b0Gdm7FMQEETbxMb0g6Wl8wHoieEoMfpg7GEq+MFg
/6fjUzn40NX2zGDDvq9SNSUlt/5Jtmp6m+qfrgWV/WAVDWt7ePCWZQ9UC31vp744HL0+djeiZaek
2A+DKP8aqT1wLuVqVH3nMVrDaW+40niV4BjAiil4FpuU8ZYRd/0MuJkwP0KKEzqdcY5BbpnA8yfb
LEDFPlJwHh61fYpmD4pr1hmhZtb807qfuvTpeU4cnSkT307DHfLWu0SQvJMCBrDzqHBjQA/AfaOn
ZTHjG98cfZQQB6g5S3pu6YZ74LhjFgnOAKSApUuc9/M9mO3Y+a9qES0YBtC2FvnAIjDMaeNjt+ei
1dNmgMrKXIrKn+hJivz6mU8uQ4xdX2k6W/u8WRAUhk7CSRMcYe7SyJTFYE0zFi7RwgO0ZbTePUiN
Vnj7Esa4SDlkTugVhIbRP0JcaCuWYlGVdfRUQnqoaKkLXgvQprCkzule6XUZ0XVtcPweRmbW0v9X
epjB4+GA6NvaAqgUmmdqeyX73j54PJtxaTyeAchKltP15AI3St/w4rDKfcC/T5ZEXQxEqcmY3/gy
vnJH9p/bD+eLuEJroYUlBOQjobScasuHAbdG+E0rkuGxu9GKn7Ci2TMsJMFgse6p6oc0bWXMzank
TwRs7O32rXWs5Vhv4JGVsFCTUBhnMMvTyQdGt8IA5rIP3EdpmRCeXnlAKxCT6AMeHwatypKthlOM
LVcs3h5SwWV87MPvzZ9nnOVoHRIPGWBaao6qgojg7dK6xc2e7pld6Rz3VuMNZz5y4hMrfIO4e/1q
lim9HvKygaqTcTxPH4RmKOWK8o7q4haaRSAov9g9lTQFkUQdfve6wkRADcThE5+zhyHtRtB/hbPH
YuBhGCwx862aWkZ4AEpQfha3Cinom7ASq4kkpuzL7LWynUUTNGbMYYE8nQlVXV99t4EtIx+x/Wor
j/ldqAWKU4aWs+pV6UAW/8tBJqts73cFlBEpCsq5rK3lbUF6hKw2YB2x1zd2OdbRZDz2T9n5KzLy
tt6KX/rXRTqjAuX+lHNMjJqXi54uq78jv0j+FrdanpACMz5ewWBQsPQw30EEqdoGrFq/Mqi2gOtd
PtrmY9+BcUW0eh+zGwuR2wRBEqTbjrNFE2G5x+Xjnj69WsIbRZkypLgNaOBHmxUMJBP5eJ+6jugF
Fgu37JEnnBuaG0M6fWMkxDPTvqMkBVOrwJ8ynRir84vEKc66WRKEhXBrIjO2+1qA8vOBiWtu3h4J
Cn86ezeqGx3tIkOraOhC03+L17OUrOaaBwlbimIAmTRL0jNtNZLffeYmidDD0Icl4GkS2KsnDASE
3r8l+s0zh7X9pkETy4h4HENp1Cq+SeuhXB0Wc3sHbTTFJJvl1kJzYzWzetLIY6oToW0Wzpt4Abcz
+9KEP/ZR/uMYz7KZUDlTqfC7enJtzcvRKRwgGfKjwN/Z/s1rHRYkG96KH7XoUOkisOJOf0G/GWNt
V07393BXI7n9+Q1nB7O6I8dyYNH1ql+K3gyNPhWMXZ7hYRFXAojZSRFkQDM/fEZjzxmHo8xbJE9f
Gi9HpK/PK3F0fhhMlCsy23jqaaOxWH0CzyEEN/MiGCorfdL5YEJkrkR2E4mzbxDYVBU4xvNkSVfX
rTsMb68KJKg+JZW7A+qmiNxgtKtFnIarOfGUAR6ogyxz4+l2RN5Auj3H3Q8FPlMr76Qsj7NRLXlO
nBKEacsqnyJyYRjNYrc6pI3TSqAX50Yvvp1m1EuuiAo16QbL2OaO8GSCgxNiYALtR75DeW7irG+C
+pO+lzcBSf57oinJxic/6mLDxL0MdB3UDRPLmtqNdLUZr+2ciZMS9oyScaggk7sucBA0yFaUgIJ+
0uJiF1oGF8fwrkZ02MPmEDjyj7ZmCMXkVMnQBRGEhCLLad+qbEcGuc7Hle/Y+Yn3+bdOEvFjhu3J
US9BrrolbqWM1r+Dxtgzkr7yrydHg9ENAbNZpXkOCOZAWq6q7fabrwayQYL5vFhTu90NTX8FpLZP
bToINeYumSYbfUmR8Wi5Z5uis8Wnkb1jWtvX3vrtv97yBUD+TfyJ14CmqEm4CUC5jCqfnCNj+Q9I
opg1kJ+D3qh4L1iwVPhCByHrPZ/wQyJ5MJ33rQNve5+6iEUGVN6R6bo69bXBsj+LrkFW1c6ExLHN
KwywazH5GfG+nm6cg/d4cTX8thFY0r6TZ/WZR1rmoUz2jZ+331BGEY5At3PudpuTh45D5ljmTHmY
6zjwNA053hqUFOruj7d+bWpWChbYe5CxQR9mt261jdLHpvtd+hqm7yN3/Vqx9qqz8U/WS9ywRux/
TgY2AsENI+F/ODvLIv3ni8xwMG+NMiCT28l2WahwTZh00tFd6PQWNd75PRPqvQa2bqqSuCVg92zh
cgQ2s+KdySJcxs0P9OQD9dChYqzcFccgrdcHSeZfscbegujxfo4PmffSG/25Krumik9r0s+PbMiI
1fQZvfZZfomGavJPFNhokQLGZZjtLllIftOMEpkfGoCVtbu4yjXvs+6GKv9MpR4hGoXjNfzXtKne
u3M28RirnJE1tA7z2yNPhI8vRCfMw4YOHgkU4/ij8yvDK4SrVn5HZ4IExbDXjube8/HhNcxNnOjy
OrPNGIBHTr5V1Z8hTa5QWTAsR3HUuAn5j6JM6SA4JGqWojEtuqmeEOPxPu/HE1uGHD1/K7pyrhzE
o2BUz9f7kKWBK2PPQpPAZgTfiFgtsn+aq/QbyXxnlp5NH11jS1mIt3/HyLkhb9U6Tv1tty8BRKbj
V7IxhfWT3Z9aPwT4c6eMYNTvbtvKH0Al4BVUSkkwe/H2eECiVlSVKVX0svtEmrGXtYzRTHyxIjHI
0USm2GqFYqXOlb06rJoEkyp1kzT+aMzHvE72nDJmfgQaO/ZVvluZShFDL6kleJgaaHKVU8NTJs3q
B8v3abhEj+bW7XwPZ/Sp/wdbnieOYagJQVCD5+khja/QZJYN7GhjOT1FyNckKZHiP/El6mPDGimT
UX1vQCr2QSFW88vHVICcsaXEzuEKVFDsW9tb+fMR8dehe+OScv1IqVI5cnIpMj8E2X0AxGnsSptI
WeHTZy+4E9OVZeuSdJROdVCPV/Li1WrIFusJRhxaoHIpq0iEmKkLsGj8AYS8/9iTZh7FX80QbU8E
y2/V1TlgqsuRpbWSvryV/g7nTVTEjej4NwmgelrNVXjDjivHZDR9XHqaEY4bGU3Vag5d+II6FNp6
oM1LXSnyYrwAVuyY4R9kLjwd3oLZbjZyJ+DIxGgMBoRJgbMerUXjoINH/aO6UYxyj38hBCu3R0Rs
0uN7qxgony4Vx3ITsBF47A7Jocj8vZUR+kLG69Nc3JW/G/m4tDY4ghQ81mp5Pra9/GTfmS85fw8c
4Bp0I+QjMK/94RXBK9Ojw6t7VR8Ir58xuxlgurlYyJo6ZPSPdoPth+lcMD8PstcZfxqe6DwTvZzN
gbkUSddsyPS2kWL3qMFjncYbYY4TPsEbqCDwmGMy8VOnZoF0n02waOPgnStiRJlfWDnaFEBbtys+
E8GH0Pwl+BFbPIlDkQQzFB15h8TuyQaPUydA7B54TvTm+PSEP522jsiOp3aywfoj3ts2KjvVSs1m
CyMhKG0FdzU0rWc1NmiiAjKfGlrRFhyO2dwifFH/VodpuDs1J8eF/Jj/2A7XQUUdq3seSscwHpDm
6mYL4Z7dWL3b6m3wMNeTlmPV0EZydBlR/Bz2zae9saQYHLmz55JsiXDRR6QMcG+4PcLSWDwgUZBK
9nXUgTdn2xg6Nj7dPIf/+Cc3Hq0t3zAX9GyFNfkGaNNcUhmb0HFwm/E4OQ8OcNqmV0PvbqSfi7ag
yyqjnNG10OmPhOegOPWqI2GhXRqEMDgQDWeU3K5u1VdNQqNab35JZOjWrbbCo3HuHdhKLGxH7eZx
2B7cCz1chteXsdD1Y1nWB7ow0K0bn8FTA4hxSAU6k0Q2ZmPeKBV6zDZ/nERwxGf+4zhoHtmKFvkz
eR8mZyT9CVilUQK6iMBA3oI2IE+J6IFf7ZtvIynRCZ8HUTFPEKep3L8hKnIOglD/Z4aTZ85/fPMP
U36XICRK8wUvxdvTL5fGsSrvZckTpZiZLTYzJX3J+Wf+m1WSiBxxOoYdDM8fwNVHcz8i2/MST713
ka5t4x5d7rU8pElwEzsayfPknpkdYzNnWx8pbjxGQtn3wXJJxslF42aH2PfQtv5QQIVXK4nlBhU4
gVCkBEOL+7UZSpXCPRCuiXuEaj5YD68rTYcyR/YF15Pza2Acz6hoQ35Lqk6FmoZQzbnMHpmGWtKY
S2gm2yYguAv6nNIyviD/8iwHh73TDHu21fuJXtaalJKgoK4pztYUNJzBTzu4t0IherPOyid7sqjk
FKn0JtNPQou30nNqWbNbNwrtaXvD2clofCaRdLquT1HRv62kxQSmAh9IiHieylLTWuyBoXylrdmB
Wr0VtPT8PkxdG6wgw7hr1BzeUNK9mJuq+gHdBKMdgWaXwy1BR1Z6rjRo+KYy0Zde44n3+X/LF2s9
svIztpL4pzUMR6rQOYTNj290gqoL2R5FjCdH5fevkxbhKzGG0lYnzfFhryeJyrcbWiXZjJR9kIYU
fCf9zHA+C7WqPL5hVr5mTS4nt40TSFSh39LjypkcNU1z51gITyJs7VhIo+lnQX0cMpi1Txn/vbLG
11rAlUQlfzqp6zeNTg9npiHr1bytA5reLdDytpx7prAbEYJgElXWXbsF/6AjnRVmzQvCu9r8cZ69
SvTqOPR11tQY9zUxobXS+KPYnDMm1hMMhBl7toeb/hSDKk8Gnz5WCtQfw5dOMoMDT/+2ZMQ+BheF
keWLJ2tCe2HMC154lF+FzV2MVlWA+UidLBaQgUxSpU2fQrDn3THX/W4XKr+Tv+QSEEEnMyy8Uy0a
jDR2gUWW1KlyG9dErk6AWE9bdVQ1O/4S2eHZ5xxmRsJ5c9bhFyr6BwUqFdVgc/tajUUudOj9TaLq
NO+SI+M/7ZumVZc3OSpbYTIqmTpyloEtYML9Mtv6da1htN7z6ZND+Rkb6ZzNNC1FrWPslgJBWNO7
TEmBKq2jf+XqQjRzRTK1dq1EqsoN3PdAcbQO03SHDXDikMGrdEiJfrC/6piIJR4L4yFgufai7o4c
o0fIoNEXE8hPsHwmo//TUo8yzDWQ9VIm9xJ1yWlv4Da3lsAljmiqvaAJTos+mySUwMdhChzIcntZ
xvWjby9sGw5msa/z1voAcMtvF9sq6OXQ6WCg+0J0/RWdHW3+lXdvLB7S8g59yoDFUQwjeB7iqXfM
WeWL3c0TX7WPi+jzfmht/eVucrQx+2u/LmKZMCayKu9Q0XBMh7UgqZhUK/98ASL9/z/TomZ3MtRg
uH1+glQWMyvSkXbiV3BT+bg41ZNlQyz1b2BaELeu31QRThQeGBb7c5Hq18g8Wqnpn5MREEfrVl5M
AvNwVyba3CaJQ8uuMci0XsCnXzsGZDIs8VfU+aYz1FoOYdagfEN6Y0lXQaS6Xu8QAJU8YkfOFfnL
CYbumV74K19vvN87omez7xdlyTdR+c0yM/FTYea3zHlohsaIXluxhfpISTggfN87Zln3adkHwTN8
2RDQvROpm0VNHZPT2k6VZIZsPklrpuUudC1XsZLD8yaos9JPNJtNEOZepBUhJ4oJXeomgRI91cnE
OvziYpKiz9dK+3GOYmBlO4xl97Tyelg0lOvlZ2g/Mi2Uds3SjD8bPw79rgXNaDWUZazQmPY/IUdW
CuebOVt5ljm5SKP13hQ4NDulqlfGb4TeKgiL8+nKZ+0e/K6mNgBxwB/yLMyu3PS+YSdiUQgz4zLq
r0cO4p+OJpqzr/rkkRuyrI76/bAxOCQqQV2zamXpzDXLwWWCta59pa+oCQS7U170RjBLqfs1l8HV
l5epIC4YRK9wafi4EUfH6J8WcVW9GjQ23lrP88+RR5WMB0ZgBpsAf9Z79AxSY2kFj/qUaqVyi66a
bsgY7hnua9cKFfntfRGx80gx/DKXaovCX0bQ0LSHd4D5VP3ZPc3UFfvr/rN7p81MzALusIT/nikW
XBFRuZB/LZ8cJsV5YTxArTQ8cE8FQk7uKZ3ET+bBY+lBb1m7b7RA7UlXiBSbtHq8sskfFu5SR6Oy
cbMd6PveD+cdhGHiiAc/Mu/x+xvEmq+CPfYROAX5ejiy3DNpgmZelN3Godt1zG+z9gpbMr5CJe28
HSDH3Txg0L6S3HOq2ZR46Qce46pijW/ltwGcl94YnuQ1pMTQvORuqkmZ1bNsc759t64vZWDt+0Ib
U5nkkkfeMCn1QH+ezto5xLAdLf4E/rWfkEttbXRhHCUad4fYD3JAPYdxrv3+MQe33L1HPUOeq1Pc
IpKv/bTUVfRvVIiUaRf6ylx+riVl9EsRwbXjDqxcYvHpoOckGzAvwdtoV+4uG2L+GQRzvDeHVuFZ
1SqkWV0K6h+YbmvSG8LHWBrP0uMIhGFKO8CZ2rBovN3+HcShkjDeIvglkkMvp3E5kMnS7U97MGo8
R24kc1xGfMGLWvbchlGZHcGVbNrBc42qY+DuvpSypZch8kru35UhDV8plkuEPSzsYCTeExllSW51
HpYdUS8dZBIjd157tvQ73H/L+BJkvoqgwi38fduFyyCm9X+2G6V0qQ4k4/GaWiT7vun3RspgovRZ
FethhHWbZ6/5I7DZsA44w0KTOFepv2PKeY2ylmq2aCSt7tCQrfXbpgCKPaAYxOcPDCMSGJe/VIAE
UxOHzBUwwGrvzdpOkUF8OsnD9Tg2lAqB+DmbU/ydRtcZDVqwwewCqrHIsnJ6yq0VjWgvIEFDGT19
h5k+UYhGw19BnIGvhafezPVIAwvR4A8ZC/rQaW0MBOCf6M7Bwm8iPw2/e/Ec561DcKexd5X45Kcu
TyN2uZiGjvJgYrNHBnUc9ojfJiw8NwXXdhqOR9d5xAq691dbBbbfO9AHC/MaArZeSB9GSfJQxsfU
Gy64pTqFA73sTwvLZaJXs+vhGRRfFF7dUGNcKuZPI3i49AN9w68Jn5wCvoeRSElA5ieZnwUix+47
9ctfUemG4EG8+biv8XCvtokub0rhF6EeWUb6yFRG1eLAWKHS/0wk/Esdjghvk7Ule8jMumHA8SEA
qcahfZGDPbTZ1mrdnbbqwTfZfolGABSsfNx7Gl6odPVxYH+XJnyTyIlqW5mPfUA7L62KEpJmeIaq
CoujSA6Kxy58ozyBX+v2GmjBjpwRLM8cAuusTgBWsHxPj317U26MrhAphcXT7MBxzDFJ56aWcPYr
hoxFD8qSrSgRPpY/wKB7zaeeScTYBk2qNPEPRRO2IggHTis0AcTiPiQk4YjuUKCq9FY3+7lk2C72
8AFh5ztRnXGNrRvpXnXvvYvKhliRaoBjih7s62oOglz4dHUaX/y29S2odwwrgbnGu+L1ZzNOuj+g
DJHgbEcnRbfpp311Rl967JCuUW81CabrGhIjLWBYcGxTimq/bA54UmT2ELErc8cVDNWaaJvP+qgo
Doe4WQTEWdiIY9H4j1rj5+sh+kBSzDm+S1d/CTlDqjUkJEGRTCn003IvrVzKnmc9gUw13lyc3Z6A
7/CRYTzRqsEqyRHmoRg4E4vja29N+VrenZRsEDj1+d5B2yh7GEaP2qYZYRbM2xqYisXwj7bbhkRZ
q0fhXDu2ROPjMXbaQZVkfyGkD5xKEdbIzcxQXyhDkXHhGUDjcifM6rlSVTF0pZ7KF3j8+x6/l8lI
1LKLp4FNkHMdTEh1QjNLfs0feHJDckRQpFhAJWIfMTGiW9IUnqmuqqbYpeIaEP8WHCyh2vcXi9e1
jzr4zme2d44RhvwevU1/bD+jE2a7JNyPvda32rAWMCcEeNu5vRHgUd6FzGc9JiKDZ3aMZ5drzg36
yDuTydny8smEA855pD2TGovKXXEjuA/G+Mgc0D/sjDda0AVlmj+W5LrT6/C1JVtjpHKvcuZYMugf
hUYuIV+jPoDZ5MVSzQlDoOsCeoWX8dbgnBP/lDs3t7PQD8b1AXfV265ayF0DwZpOzoxWk+RJfKq5
NtLGM/zv7w5ztgNefV/IgSnoA4YhcrGDAOMi7kjPq2DG09uSpG8kLrOTq6Hdqc4FKb4aBLqBwGKP
vYrNLRPyCC7Jylp5yOVE/of/pw+vY/mYuU5C/P+X+PZnM9ubm3JDvAulcuniEqdw0e1ZMsj8ecFz
1jQeTksN8OPaX2V0TviIEO0IPlOeqLRehlenwF4MWzwHJln213g3i4e2bNcxN7FB67xl3fyowX8N
rtNLoyMuPySECmHbXpUwUWaKcdk6tMWJ4bSZ03vn4JK2sEoedmHjWm3ejbRZD6DCjgw7eWjMUhcu
f666d/xAuLU08bmlUDztR9VZJZWRHjdwYoF2JKcfCUwMlEl7KrpjdMNH+PwFZRr4jCMY+KbWA46o
JJYyLCcGYhQAe3C1zydwjJr6y6GnXfBfTLB3wS/FCm/wI6uCPI3s7zW+36dA0Ngi8+CWvhz1C5Pv
Qhs5BC6KZLiBT5Z1KGDGBXwJ4lHT0qSWHUwOS7ietJwKmcm+2XnRJUaXc8qcP9BDbPMy86ZOvgaa
ZAyrxLXsZ/4PjLEudEzQBCNIFOLjYdh5VNo1r2RUiFkSPaE+yYsq2LO21B5rKVvIvCvW52AD1Do3
L9OL+WqfEZdVeQou3LkPwW7BzCcajv5Hybt57kM1ijL47qtvNXD2pmaYJ45RFuF8ZVkccafU0X4N
UX0i84PrpXi28PT37DauaKm1IWDmgegviuI5yh0nmvfrXa1EtAutPJpDNk70UFcj9gIIsEYFiAOe
p8re6JD8bPxlguFoVYjHd2Op6T5EvbUgKNrmjA8wPEun4ZSL+6zR7t5n4TP/ZWEYFKMsPDZcHhO8
4edchDj2plVXXwarmUMe5Sl4Oerzp1K3Y3O6xNvf38viDbtAdFjhU+K9dJqvDz2CVg3Zw3HBd6ed
dtIHPlNytWZ9+OZSBNu2Bnqzk/9pX8d6G1LBu7vt5UZw6ZNYtRVx8uCWZ2Z0S5iTHUg1MqPbJok/
r8bI9ssP3+SCmO83PMxjt4+Y1kGw7F814Z/WQc+ScSR3yfqNPx4ARo0vr99/AC8363nHY76afX2Z
GjrXyMnSzrXUpCuIgcaB1M2C0X4ZTgrDa/Rvq4q3QOJCqlmmDz/ey3XMG/LlgjKm6hjg3yHr4IZR
+ezPLZ/G+eeR//n3i8Y/2gPRa1Vp+KHQZc56eLmuPk4Hvljfx28OnWLswpHodvPud1f8etjwMltK
5hs4ftVsQR5P0MAFDlBcAmKtzr5DrqDdrfuJ2LnA5rB15SNVsuNWLq7qE6Ta+ts84Ez2mpgW4rHj
AVYbTA76QGqzIl3GfzJGDsMu1Vn1Ks3AlRWgqTkTfoArtDGIeT3TtJk1k8Sv67FJo0s5JT3EbBs+
QZPNadmcn/fNsbaSFIZ882ffpEu5qjJjTTp1LMMHRU9aF7ArnKsGJb9gayY2VoxPTcvZsmYQKpGt
Dd8pICzXuU1hWJdIgIlx9c1Jw4Kd2znTdYSG7k2JfWuy5MWiKYBckzXKVbgeBcAviSq7sOnM2zLU
tLtAC/RYpngClXn5NW7Xoru2udCnsfUB5/LlO0hOS7SaX6966ZJRKkHd3w/YrPWfTJOYRoLPljSG
FfBVV8TfJl3oGmn0bQYFvEfYWgd9FYwm620ZsmLrTfzWNCTpIgJv6IhfrQbUodLgfb+ws/+Cu0Hv
mhWQ+vee6Ku9AWcLrx3ed/6S9Ba5Ej2FeKP6Pv/+tYYIQ6r5+lL0eWahJJuU1BAexeOSU5cVLkpA
RKS8fLPp1lM28UY05+PzQqsEHd1p2owqixHFTAnkKlYvcrdsCc0Wn3lZ7wj9OfFnuAawDDZ/vwJn
FAIsL54kIZwWVASZoyGRdofmvrG6T/KwxhRwX0jWOxWbqcUIVRV//5Y3eoiLuSLgXmwmUI+xvdyS
4sKVIu8TLcCx9MoydjR3YmBTgFDjjB9+oylOu97LBcupXAqvXKm7ckXatFiFWkRC3Eb+/kmf7Ihr
5gE1yq/sCOREPU2xRNTxDFQ2PNANsLoRGPssvwB5KcBtx1VjQrclscJ1WxeOw/GCsge0BV63wF83
GjdAAn+y7u2glOG2nWpXkCRwrgpD4VjEsA7AtXJj1kPpwyPjpEP9VUxYA8NdK79u1+PKizjs7DWj
w6dAmmXxBOZzViet5Mx3A/+0OrlyrGcg+x8Ep4y/o0agIRTMr7qmtHizhaUTo3dta959GWlDhJmZ
gANrdBSesjeqXX85/7RW7csuRzRx8g/oUzfbG+f4Wa93LTPY/zrVbUTR9C1ptVGGSM7hZELq/lYl
QS8fttSLHezrTvGlPsqoTMM8Wpxjj7QwKQoaviYk7qaIkEaYCOYsbdSeGzBBolQXBVjSw9GAP4HX
JGzmKyJiaCmvQUhWcsg7q7iRV46Y8086pQHaYqGXecRSactOZKxA+Y1LY2PlHPkQyy7wlGlKIwIV
NzHxR4O43QETiE+cXXJTuDiptTTkApdjWxCM+1pT8UaQD8Bpg1OnyjEVApf6Pcnfr1yQ3cA1bHb1
nc+Dv0wlKdxamsFG+r92KdZWUK/r4/8ZXjVjFpX9PAGfxPVfAZ0zjxltV8pFZnH6IY8AyCclxb9W
AzK6VWHupnAMOkDyZ/3g4fh7OipYXTaWR7FIMAtzuk5FqApItADUg/s8FnFV2EbzCL0DkoU+hVGR
IDtXX4SD3MfHFIBBMG707qrZvDuilR9qBZqgb1yBGbVcslLHmfRc2+gIvr0GRm+e8EMGlIouzCgX
yvhVNa+1QFVo9PaGv/uJeDgi+PGm52QOKWWdhJNHhVzlayBTRMlGW0HGDSAAOmgNPtfpwWLW54P1
5l3YwqjK4njGXewugCo+6AC49LfsvTFm4+2XkSFpher7OwhoDCP+iMx6ON0WrbNujvtoHfbs+H7V
RmTXk4VcZ72OZ+5Y7QtXNs7KGKvlB6z/ZfcsRKAPqkLtbOx47YRdwJ1CCg4yf/tfMFlcsUPb4FrQ
FB6o/kS93lXVgwxBlGYbkQxybk2Lci2vmi6z4dp/d0jf4YHNx0ExuJyJRu7pcX580lRIccXHDaZF
dzuj5iTn9x2MvtYcfJ9SAVan8Zxe7hhUCVZxqO55y4gozm3lGEowo1gHrIflVvHjB3YCfce79/BU
nJEDM6AVnO+YqrSdtKX/CR/oM1xawCjirNDeS4A71odld3OC8W4vcW4hiwGE5qMpQRmyUJCMTIZR
+qns/LCPMvB/sC4OYKcL8pRm1LjI8h941TJ8r1K0REX0/gvT/qHSZQuGg6CJKFEz5WUV6JAHX4q4
BKlk+Yui/HPM/BfWSBzIV0Pi7Bw5oQBERLB/KK/fjS+nZOwHsTH/poKG1R+wI4eNz8JRvhqgV3hv
F9Uxa1ZLcP7SQQq3thq1egxvdS1mxJfetY6jBBIasILNsbvlnMOVcioJZXpzkbUB8x9xXtt4wHYJ
kzyKxw3ZvgLgyWpnbxe5ycTBUX8rh3wYqqFGetChXi7IM2fgITNZ9pnD1tBo3vCzIJECSWJcPPRk
BwcE950JEmEqUcrACEg7lWW6z2d/0nGXsKBXvFp+kGKWAX0NTI2n6xKEy7nLB0LV2wD/ufv7k5jR
EDwwSqhlo2zHZ13lw4zEAtKNujPDy/JJqPZH8jTiIgX+nIi/4LdUa+/dAQZW9sAErUsaOAMM8qph
KKUEvXoSxZUrVfA6B6k2M6f32SBMERKZiNEDtVBK1BpzkfxRF2rRT3XWKqQSqRyqlKguHiFIWP82
RPoWnNcbivVwIRzQV6wgykAyZ+dmfaC+h+F8YmeKWru3HLp14MoqNF7AB9KXyydKhvFcdwBd/EIj
MMdb77yrYZb47Ph8+UrN2/rCCKiJWMisf0uOxUDh7HI5Sle+DZbIoflUUiTuKhPAi99q//8yTaPq
olKjtWvfvPg6HuRiIzPIc+m3/EL7jg25/rh8NoT77jScP1yLkyZvG4kjDgbx/3fpdE2xNEn44gkr
Xop212j8E9tH9WZWUPg/IxcJPslXvikFG5rn5CBfYI4iMr97v1J4jXYIoXPAsCPrP7pmEltdXBFa
dU9UL6NypIXCOyPRrxkh9FWKFtxWDOz+q6fXhEp3zC0bpug8IWYZHZv19eJX2fftXEYIB5GiCIgX
V9SY8mi6GbE7Ld7xcZviuBG330S6hP3kRhA6342cdRQRtFFgXj4EXKuGNgYnXfC74syVUrEXfEY+
Wj6gIesqsRnPuD8vy+7bG97hZ4Xu25Hde9Gilv/x6hQG6McAxGJpxvUV1A6svwLXNJ40uihBU4O/
HmTrKbXoeQIWJp92qkYNG2mu9T32MbIXrcodx/gK/advaljnB1UNVilsW/hniEAq2+iN4pGqV/jS
822Fu/KgR3NtXQy2C6RerKGwwwTkyab8xtfDxcp2F6loz2XlhDKsCv9/R+E9A2XUuc8ZgK/LgtwS
GuzbnBwER55VhRqEZxzmmZn2qtDFkJVh22l/WpXaHDyu1z0SJw3WJsRC1DLmXd33DO2d58uc7Qzc
Fi064FBytIxiJW9HpNxhBbNaCAipHIhMCVq7kuxEqV2jrDxAaekTPk2viyn4vbplIHNgMmSja6xG
vhzhscu8X55S5exRe7Pf9QShCmCFmk7nXY2J65Bf+q+NeYkDmWJq7TXiRSRoPSK5lbVSIXkf4Sm3
4WR9fzFzuboE84KId5mshdro44Hd6JaSOt76N5kYE3DpV/UkMgLad+xtoiyqnRKtLXNfFzmcVu1s
WVgkFusljkHJ1PaAphBXPuqI6vaj3gqkg0byQ24lsMslY09jnTFxCmhx1xR9OmhlT0Jaqs6ffu3x
wNG3Ja1BLks73Rshuq57/aMKv34ZHjeslKWx6xoE/LlRxGpq27d4pKeoWS9WgxHjG0IXAUXX4iMR
XfaUvorJArMU8zLZwSyaLNqPLSUssv9S3OyzwuG74u57bhOMb9JGEUxXoH/o4wx5xlQAXp2GTsIf
/XUCsu7WMXsWCKlEFYumr19s2ohk2qpP+cV3U2CmTMs/oqcOvOV/gQewuSJDa3jXxR9sD/8umnir
RtSGpfxjJF4q6eIYhtYkBW/ZYyhPAssM7A4o0ACNjCm+a0HpcsB8oJyxktxRKhLNqrmcHs/k3yhH
PSbsqXUyE4zMeYBQwSzd3iJfCWxHeGskQChAz25/vsnPYW6npuu4RcqWP10mCgn6i9VdYRgNKQJZ
GNOpnlzzunRt9T0AwVgYJSQuflWznPZ0lS34CqdcreSy3QS9k1EDdqWoyhMV77ET9zAj3II/Lf+d
tHVE7Eyuicf3Q2Is0Kps6f0nPo3qJP12U+MeSxDuc+BQlixj7PS2UZFC5u7bFGIyXpYhCUQ2BiAU
rpPEizPtyoL9KX2qLR1gJwTKkz0VRxeXzU8NwvW29fSW4anogmIlvNLZOu7NaujbSRsLlOmdhVQr
EUMNADzFrz1Lui3QeTsvLuduJjYbbIBz/S3gojSIaTaF2N+AkPMhcAwr+i20XE2jUnHrSPkWKD3L
XZR2+6/mo1Bikp2D6wfYFuGnbQ9PutesWP2117cPOMMu43FbqzagFdcerW3cMJFiAcCu9NAVc893
SzV0+XhQra9xinJo1tfXzzZjK/ZVvC6phoGz2B7X817LKe3JPYotAd/epAjLNNYcNp9zxsmmXEqh
lv5S4Plw9YRe3AdlI0jss3QVpECwzYmGIJp6sH9uFHnC5vw1fK1/IfV+GlgK7INkMtfXdFQFoVpb
+TdOxOcRNdIw+QYpI2rfif32KF7XVusV718b+8GM1OQn0EYSKGdAa9fI6CWDHFn3vmCnF5ngD3pR
C4LK+dyf+J+MnaoiFHw+YG0UsxczW142oSq8UMy6reV3MAW7J5lBXJA9ogtPdOxwUxsM3t+dar1Y
WXUlm+PBk9ThEBzzS9jfvBR5VE4BKEa6i3jeIBbBATiMksmGK9vEg4HyJwzxR2/Dn8lcC8qqLLZX
WQ67vtTnaZ1n4w7qOEgrP/GCdlcNfAsq4DTBRh8zizcJUXtZbFBEchO83KqESDtrhlZL21deWuIy
zL/XWXArG/vFRbqVo1LGM4DjqcCwH2So5Aw9iqD9ei7RKs8nQzOIIVo0xdTXnaVbmihm+HfafYge
blQErSZ3E+8v7JJ/xjmlHcHypeNkMWEZc+X+NqHFgMfdT0tdtCBHtbSOTkLCuVXRWp9eZAM3z1Ft
G88lT2EJpZZjCU2wMCA803FQGBhSu+thtKk82c1givEFMx9OxuhOPDDQJPCGqhCJb3duNradxBOG
dE4TkXq2rB9qVV5v7v9yc57YK7BKrVVAkDuyL171q6CbyT9OrKNd0otI5A4AOOc4OBIjW25tAipB
48GTt7o1szpifxDEW2oHeAwWBzO+KXbF1qVtUC1POMaDphDgsrOzZXYjMv1UNIkSh/NAeXglIRV5
Oixq0slLXCAIqxbZqwNLUex0GsCDYDz/S+D4/lM7zjdEBKO7235WvJiB77K/H439DI4USemV9Wdm
mOg+QdtbrCMgOTfoL4XS1hLNdnUeayu4X0kE7tRE909n1F4hF2ndf+LFaQHOCOQ/w/7vqpgqgv4n
jc8jlpv7Ik32Cice6Ry4xLyZj4nS4wAxRVfpz1h4zZ7Bagu57JD27f4xggzKzLDRkDaTHhc120Nr
TfkrHHdqcJtUb1jhf1bPl31y+RducMr+DB6XMmDn9wuU4ShFm7Hr6945QuqIF5Vmd8XKQm7x/G+z
PhUcKJ5VYdYuAyGOKH7wsDY/O+bqwlTS/A+wjg56w+Rqtci2cEK1+8e5Q3qb4P/kf2wDI2hWeC3N
AiqBPKZGJINh7pRRiCH/jhNWjVFmX/4WC5TMeE+BlCxZWEHpOoUROdLR0ONtxSbyLNtYG4qmE8Qg
NzWUhwnAPT6b+WnhJrkDUo5FqcG2DcRUCh/FXWPVs5ZtcLdJCc8xhBJwsgBb81UgKGnsYYrlx8Ke
6pu9Jg4j1WvQb+yEeeYq1khmPr34uAO9lS9dfaI4Oj8IUjfFWQ7KPhaJTHAyg7lUxkKFS4ZaFa2s
tqbPD8jeJQJ+51szRWWukmsUY95jVRhYgnpTjTC+0R4JyxZkAvKLt2mte5M88jDL5HDmaC/zRJbu
RqRkiUKR3OFS6xL1kyM3ImDJxd7lk8U/SwfgeEBj/YR3AsAwKU7P7UP0PScBHUdRVllSqUHZfR4E
bidwmBiG088LOipFOXnJYKQZ9h9Nxd5LWs9W32yOTJcHkvZhlrXJ7DYYG4rBcN/eL+tpM/7VpXz4
qtowdM/TRCoeJjsKusbB07D82zlpkme65kxvzs7lCaIGRhO6ibStCcUGagvfzNX72KrpGdDxple5
h72jS1AkJn9foKS/3Cnx8atmwFsyWL3WVVnIh45NInt4+LRqa/m+fbuGieRoDg3ullJn7h3GC3Z3
2vNr36cXaxc1/y+IOyiZn/pKaKzTpqq3VHf5flhIiZ4GY6c2JWhQy2kSBGr8qUM1pXRFA5XJt9q8
FyCxbPQH0lQLhupZsU4zLY2o8AmMKVQXmXuxTXlxQ1a9ifnFIOE+g4CMNJn33XoQNeceGXefPDMr
eDuJTsRKcm+1m84HIUNjCI++gJ+UBZJLVKXR9XkltHVTls1CEHq8Zd/+aqhtWVVlk0vo0HH8TMOy
/BG6I/Y/a5a+/tnYTpgMr9G6dch3YP9BnN1SNlTjVc3TSGx9zODMq4CtVyKJ2SIxwI7+GfBC/sds
iIRIivg2ST+RUQqu0LHhekO2R9+Ozs8snxS7INyjtnBfv+tXDfE+0vnzf6IUyjyHzud7q18oLaVC
0XOZx6hMqYItrSRV0FbGIwea1AkZAvHbcBJqfHzCk0At17ZMFcCzsyUQKjbo5WvvW4FiaKEQsFS7
Z/VEIUS/6nr443D98hV8mVVHXxZieLnE46Ybm2CTOvEdQio7gTue7N/PGfUID8MZdUlpdIL4iGx1
0+hn3nPGE9OZ5Gs12XJoUtu6TW+ugeiUuQHd0CZcNefu1S3YLB++WpGmk7nCkBsJVhGkfzlbj3b/
h3CsaFmTFx91AZgG0KfN6tjYamrF+dd0OogcjFjHpj/jLOEvB16Vsdj9n+BPq1FVLklevmPj7o8M
5uk8j7V8/7NiBc3wSqalYnlLpFjg/LfkB9CtvMeS09PzQAqJAoxYni4eIqW0jiJDdLsHjn8n5bjJ
JgXian+TxEkjc5KKMRz0Me0A/VV7GbLZp8/TH/g1ATOamTgXNRKRnxmOQOxGKbRRwn/IlCk24ugt
tgaTLwP4DmKXpm3X/oIPYX32JdWtpWNEzx2P73Cy5EEUHFjZkm6u/29b3L/zM3nkAuM2Rkzhr2iA
UHaUqOGWJcarqF6nsYa65kMPPcZ8Ez9Vt5UjlkpUd+h30r1m6rRQHCVvNviPU9ssIm2vwfcOwIdK
zcKu/OG9n4ce4ldnod/tnAcmz3duMXewhQJI59yjWUba8sewTfW3U06v/bOteLxzIHPZtzmSSU8r
hohAHFkX4NrWHne3EFUNiZo7/HlNvBVDDiUGExGFBhfPPF5htNV5fVk6/IS2X0wfID5I40GREKWc
WrfL14xQUSyuf8NikT0TNzBYh96J/A+1r03bCxKHITThDJkLSDb68+iTrEBAvY/KgnGiGlHWUiVH
NQ1PQtJ24GWc4P+h6on1RcWIg1verrFFXNzjPY1Jpkj0IyzO+XjWz1978Ccd3iIIcedRorRlQQaC
Yaw8XfZlCTgdwnjHpknPHxx39H28KQzWuDA85dDCdt0HLEi+HbjxA4NOI3dLmfWpWzokxFcMcNYK
aDUqYThrObVVHyXNpOINpLsQxR1hrKB/oSVi6vehWbKdGCeYgidGsA9ytGN4udpegQJvtpXvkZcN
8k2uhX9ujb3A9lJZF6uhfVEJDmQxyHZgSlmacfD2FJxoZ72y0Dho3tCOypCHo3lTGJ98GpGfXvca
gwtLV4h/VY9VNjVEIeBpHtcxvPjsQ9c6FsKUQEdhJbSTnNyejUJXknriM9jJIeV7JbPZZNC3577A
Nj/9Z5jatfx/XnYgxtLJxvsYFllSxbfSyaI7RhBCMljr5+yNZSiUGl7S88Et7JS7vaioh8sBPNFg
J8USE0nBPQ8a9Ue7Qi5DYUWYU58YN1mwi4lNsVf1tH7V4WxnzlidBF+uli30E4HpjDhgJsUnWBEa
Zmc3lu75f3m2eD53qIVFkqsG4AHif38XY59Nf/Ozj64PINZT1IRDelR8L0hK2hsM6mXiQCbxuIj+
LhhoAUag2fkFNLbcd2Ct4YZYHgAlZ6SKXkJ4kMP5P6wUasugVYTfOtwagaslMBhRjEDcLLDE9LQn
r4ZwehTbv9TGAviWVP3bf/Z1i/c5YeQQzT9Oa5nANT0NuwVdH5fkSk7XHFG4P1vizjCeXf6+HHVn
rVjxoEKY/dCm+9TGEcP5oPpf0D3a4QdQ2WFAV55gVIdzyJST92OF9OK37s6u6ZfwCIMJwOUCcVYQ
M5aONt+hjQPIIoP5VxMh1wkziI7QpyRug3pxc6YcKOqfKH45kmn1Z5GREgBQTxrEdTHgTLy7CxXq
vIacLMxPkMkR+wALO2LkTNKsJBugNNrXeSutYFVcc1AHK8fnzYMx3jnYshszw5//EbYmyNOd/QES
ydlP6pFIIZXGlPsPXTjsEDvqIPRw1TaUx5tLnuZ1wvI2xxcAWZYb1eEiU4jf4BqLl9HIdWiYL4qQ
UTL5TJUmD4A223aVJAPEYgwux+6J0DWyKmNxfFyfRgMfqQOmocGo1JxvTlUuPIjztnEZ67pwk2Wd
wtGDXdDhl7GN0lJTIR0fF9++NbO9I0aIXrU6LPkv1bMJRA4Nj6QIrQRKeph2S2LwqntKJWMQeCij
+wgpJl5zp+ceaJFF8XmWwzNnWVBTDgIOuE9LT2XMjVThgybp6/ZC380rhVGx9FKmoW72XCdbxGKh
TWF0dFI1PfFFSgcbRTdBCScf6+l0eaa2seS7UB5suBGUArwlRAjuj7uSeQySaHnSa1L2KDfOP/mS
aR2SR4q9jdOOtvofbyi3kRzI4GBKbKyJK9swN4OIm3BrB3wcsm1iMQq968Fn3DmSR5BTyHg2Pw8Z
gMwfEsx89Ipf1YEtzX7qjuaseA/LIR9Mmyc6UW2uYp7oAEUUYbOTRbBSUyjbMcX1lr+pRaZli9mq
R6GToCZdUh0TJh0UA1rdiP3L0fOmNiG8ScN032trdqRsiLDyqO64dBR6PH5p2LDaxbHdYXrSSuzC
3MJXaDqvHaGdAoDqC2vYAti79R67I1Sn2KdoYkiHH14MPl4plF9tltM5ATE+bV9CjtWx6I5u6uQT
/YVHZlwqAJe1U5OMjyk4Tpyr7j7VVUHWr2bjkkIs2d+rGZhqEObymuZxzLEGbmH0PCY3rpjdFqdY
uUUHu067r3j+XhhFZoypweli6+zM3yQzf84aUaoM+VxybC8Q7J7m6Ez0l7EuoW5nXBxYm8tmZFEB
bPLVmqIB+WCvC/c5eI5xIgo8WYj4wONKBMgsB/PSufDwyWgLuTyoj91JDs+GxW/CA1ptabHcoLqU
8BsfJYFt6Kkfj0m8aVlnxjwgZRGaH1ogLhod9kDOVm3s8QHx08dcseqb0j5aTAsu6I70oFV2Op5X
EAliTNTUatbVoBvMKArcnyJURH8URvPdMpOSOSj4ugrLi1gnK038TFAjVIUZuEZIY/nZSUzLsG1v
THA6Jp0ZRCXugIfUzBmtlCMsQV55Ez9rSji2FlJ8jDi6a78+8vqePbylmarP7yAy8Gc+EntOCrJL
bThpDXXPej2TbmzbOQ6KtX9nrqg9Uyq7PryLMrvwif5zUzglqiLD2IRoaCXAAmzs3Y7nciFjzLTk
dGHs4aTDyXBYSgqCBvQ9FucZxm1Y2pdZVOEjukP+DYph7wNe7LO4Jd8F680hvMwm44pDvz8YMfu9
VO6T9LqMq/DHcxiTJKsiaJByFoWjSflLyi0yWQ3hZwsbBRqPNSRb33oJYoTg9Gd2EMptl4uvy1cM
JaqaXljtiZYaRnAk4VSX+uAX1ZbZd3p/v9GulNZrx5JqxwQZWKiPzgWn6gK0Z/vjxuO6c/RQJgeW
Lc1vMWgbHK9FGQyJrj6Egdz+gwij5p0V8jxH7YHeYwubz9FzXXiRaQrFtT/xjNWngmXUggpoeT36
h7ZoWSBkFphFV54gk5Xg0j+vZPXVerkj3jZFzM2ITBXPu1kVdr8ngevAC4uxPBBCP75kWFFbCq60
AHDz7EdQonaMmJrglsmYWmk6Plp0mxnba+/fV5HpBqD7nhMa+u2NMbBIFTl/NMGIMF3wBGAn2Ego
qO4B73WUTmSFTgzykjArjqC4qYspl7wBsHf5KLr/2Yf/pHSFr38Z3GacxijEYg5HJijoR9JmCpcD
ha3//BQsfaikd4YGcZPptcHihGFhgQOHVtEDOvuwjN+MUJqc+WJSe0hR3kzsWvkrBnUgFkvZH28t
YZbIvMg7124ub2vk3QpdtOjZAn9A0gB2aYEx2nLmjSWIMedUVSUi7Hf4nJLJWO+PmVRaWcXJotMY
X1JRTID81/NzhTY8MNgfX46+X5Evw4lc8FokHPwR9EJsyOnC7DdcuFHPCndClKoUqsc2zdvIpqBb
Eh1qES+47wMZRA41qLdZsjpPxq3BtWwj1QC69aMQkVomFzHj+PxKiUashOLCW1sYP29BVvuHmfYk
2e9AxBIJqggBUt9InWvdWjuJs1SR/ajLz9bFWiUWgn5jFzSHlrB/t6kRY4vs6fBltCFxBt9mVRyf
s/rCd3Av/bXQZ/vjS/Tyl3kr19yN4qF8AIBuagN0uFBHSNviE6d6N9CIq3bUOEJbIUY8fSWvDeZn
IQp/+sHBvy/T3hA4De7F52w5fSa0/ZceeHBjDslyEVnd+9DlJ8o7964n1BNXenJlydczXf6+V3Wy
wpKLew8wVDU6QkKCDbBYuNArlJCiCSNXYIkV4GcQ7oH1j5Q5qxuU5ym4e00bt/ZLbF3D9RVpT6W7
tQhC1sUXaX1c7q+4C1eXxgsG3zJ7lMfkv/+jHTuwsU39pdNrbyDQetjXPr+kOpF1AsnSsSLpzE1a
xgMiHZevJdzcvHtsfGUqxlryypJKlsIsxqn5qoRJ8/pg9N/IfoiKvhEpZmCOwUU8z/MCqD59CWRA
vB7pFYty4S/uIh0pFyqPLitk6Z4OHl4q61DOXnPGik+34My7QGWaWUcTrC966f0nqgV8uUtV2Ycy
gBJKPF75+JZRs2xhTwBz8cze+O5ktitaC6dcrrVwneG7eLRIJoZbskxqNty03BMkGnJA5b7Bsbl8
L655ttSEYwVQVFp0vw/b86TciF4Gi5uEC+ybupQ4X+SkvydiskggtEj1n3ZQEZwuOyxLCFkLZCoI
myAznj1t6uRMFRn28ZQIsOx3KE7E/iRGEj0jUQDXGSGgtHzzhh1m1ShGTKmw5Mw2g/gvxxCw2NaV
6kPY3GvYwhEsJY72PBGFK28HG2+QxZIrkAH9g6pVMfxxska1OHyBrzuV8Om5LP05e/OVqBL0iVvz
tdUNw7sxqicGKxriQVZC+Git9inlQSRM5yn5ScYPdIl1fngNTAnXEHVCC3XiAjrhLTw/yOyiXno6
B5eLyd43L52whLhlKTH25cWTJ7e1nTRzme3GNmOTrZCXEY7HxhMx5g85gDBPHBT0C/BPkHcYp2WJ
YlqVDIp6UYTFTaKq5jf153yG/eQS5nZIQbbV9fCuggrtPozz9g5y0w6aVGdgJR0zs//iecHuvrfX
DUttwbohfxh3gCu4xXQkRQuF+UCCZ2GX3xZoiuUu604HU7i3uvCZmJXqKQu/U6clsBWAljG4+dSh
1x6+OpKSyuNH18ZPVcs5IIeMJp/pkwxEmxJknfaYqKjk/fBYujpsngWxvrXcLKwyv78CdkFiPUoG
5NeHFsamw7AU26Jq4PDTB4FyQzUS257mrljOKpnsHoLy+ckNgYSaZ00ohb9OpMLGBiXqEEwFNUqL
jI4HPZieJxSVmSR2+umlXbbp+KMmsRqmWa/MKKK4N0SvPMhA80jBvbO0cqzpn2DLt2mgSEqiioy1
9QhyeAF9s6gH3o6Cf9lESJg+11N5n8zbzSOE9meQMI5uGrtnVCpWltrNrQqZCGeV5X6yP7i4gBHq
/iTIjrXWMHyI29O3PoSQu9JCeXgH2GDQdMDUsYbKu6OL5nvR2s2AcmpBG40eUyds03spPC2KfwKo
yFUeJSYw2swdjPwv3DEJkPA5THY7eQEm61UxhBJN4Xp3MFtka1NkMfe1D7CnCCPu+sspGH6B9OX+
/Q8nRpm25g56OwbjqFVuTWSKfQfnSHDaW0yOx6rb1EoG0Lk0i99FXjrUFZh8VPzJB0HfjcZE1l9Q
u0r/2wMyAPfdbFtwL4h8Zl/0zETvhdm5f6hGf68TWNXVN0PehA77z3lzowa7vi9woAW5hbm78tEJ
MRGslb4PO+qY9IFo9sKnIBpfFG+9/ZeCFyzXXTtp+NER3neM6QRfqpVdHm4wvEBWvCyEvCPf7JBQ
d6E5sd69YIHrcET9N2XCOq30vnjAyEah4lEoP3mq7hqXSrx4E/+o6Hr38fzC2zCO3Drv/OQF7R20
JaYMiieSZ0sFLbXAaYVgRessAfuDR7ZMsbp+1Y1FVqvp+9W+A5lcwtEfgWHtRB/K4teD8TV1GzIA
Ad+fVnCh7QArXSsIcZTJzzGanMQ/1BIwUZ5u32PsAgAc3Z8P2EvQEUTgF0X8hmOhIulsaov44+cK
SSHGljs+XjepMO+jqWgm5RvRBb1tHBEMdPXXthkjhQ+TM2nyPvaghLsd8pnKxwGGEfO11b3leKks
vgHGRTg+hme9If8iSTXDOibTV8zIajktkh6K9+493x3T7FNsZrormnbOZ90MUyeaDl/KxC+6o1DO
GTZtC41dXCPEBZm7z3BKHwXRym/SF6scTORIpNmBGA7uVPDex6v5aThHTDWU7iyoCsVtT4HwoGKv
TZi0Ig64ZrMDmE5CbyKJbbPjydNjVkrQJn2N6zTnlP+qPohZQaYCb7eUZJ+XwJwsb+a99ITgQRfF
v6YbCUsCOJsrfbfKqVvMt2SzveD6zv5Brzn2OybPNjaLiNF/wY2YE+3hrjZRbEVrknN8Nai2Q2ku
wCBzangwVtwuPhPPSt7zeZ10KXIV/42M8U7aYOs8AIV78ZhbEtsHdg/SNEUU0sWkspfU/tmUupst
tMjboosGX70P6jHq4iG5Nq38L7kDRGfQtS5e1gdu4jzg1jPx8xR5GX97ZE31OPs29d3xBlarrxLG
tgT9woXtOiHuv5LQ6WVeYonwKMHm+PRCP2fw2MFmVx2yj2xeKOcxir65Fzd7uKiPlWms15orfetl
NvDYbzNLrQCVCsSIDYdpfd0uMDOUr/wbxgMKM+a04aI4eJq45EhJSI1C3zw23DaZBfwnNT9MHLAw
Lx5wqq0s1gU5pk9s/fLfSLcm2UdUYogvQMnUNrLbUSO6EQVXY5SfT47lzDk0/jElTAyjwfh1bQyO
Rb/wkmWRIW6SpIuqaizJuT+RYTEuypqoIl2Lts2eHSuoRelY7ofrUzMWLExVl8t1jCbJctqaQ2MM
EK1CeA7uU5p+aqfj0XenDSyoG7Pbllvhe0kohNKNCWOgMnu1nj6wBvMjAuoxE93XDUqM13Le+0WX
5ixp+qiMEAObaefGnGBWPI57V0c9wkf7CZlj/R0YCe7YakGmzMGrFsmjfQQBvvHsd1dZKKOnx/ad
wmubTWjfoglLAojYzcLzk8MFNXqIYVYIJdTT+axUK8z8+cFrbkfTftIUSYQjEn8Mp8abdfwtQXFC
VO0sxIUJGPkVRehVH67WKeG3DlbR8NLtIDx2G/TIucL4YeBsyEeC2osnYvWiNyRLhPuIXp+g5zen
Qu5Xyh7nP6ewn8WK5eZEDvUb1rxCQXHKH/R4Hwbg2BspjhlJ0+PZ7gFYY/RUO25o5cLLi7CYkYV1
ayMP0+Mw1mBRzYr4SSZV25vYFPII9doXD0lp/Aq0hBqgau2LrYxTw3h/WWexkHFTHB5GydMX8vQ3
XH00ykyRi23ISjKkHDx16WshP1HAQNEDx/T3oFMV4+VGvZebXx92XtMFutIX7wV15Hlh5tVSAn9V
XBp/Hm1MIXP8TJ+Anp1g4vIXSI89U/0B+ZU3jLOUJhzvQlF9C2yVd7IPMjdeRVDjRODBfMMsddlH
sdt0HJSk8txe99yoK2ms9fHryOvGOdyLMI6Jz+eYEnYw9R32zQ+Lnskd38h3UsHBMabbAim+2fgl
g/KljJQAEisxSw+pCljvCUHmCchk+G3K6NoClMIdQF6Cl3NYn86tgHUNp/m5XGf78ZOzWfc0R6u7
xaG6gZWYOCGJIEK1Z0Dp+Lo9BJIJLdIIKQzmvee8aUVCrhKXDoVPfeIJM2YEo3CSMH1awCNkBLIh
tFkS/PM1BDhannIsmgZUCoWJDkjknUYaJehye+tqrfDXjD+Zp2Oz8BRQaQP7YpLHyP08YkiBoEfJ
36NwOowJU6ZOHE30jO8ZBQuBZBDXSgGbiU9+x+sTME5p7fcfnPblxGKA0LV8Mu909ReDCRV8NLZA
ERl5gjfJbJH3ru+ouw43Mg+JQ7IejeDwycGzqIvfDixKQZrVFI0qQJkmID5QLB8TE3Un2Bb+4ig7
whZLUKn7iLC5mEcUGYJFZg+UkZYjSouXYIl+uW03sj5+Z4/7D2jSW3Y2peGeojSHsl+9/f+OpBD4
h0upA2kh++ZdvqGimjAxK4P3vG315P01Hog2nNQuOERCIGqbqxlVbb8GI/HUM4bQBr8W5ZooAIl0
ghg4fOqTyqDfIqotDkeCkbjM0p/6yeaPPc4KqUIdtw9FxAy9E7D5p84B88gRE4ur9kzCBTaSMReU
jgC5y7uLU3OnOL6kFjCWWKBcijOtyoG04NLEOiNrYpuU5XbzzE0lnSi+MmkfpZpf/8NjMgi6+kRX
3fJ/aWiqKr8KFSEb0vEdL+zAjjit7La2jFAOS1rcQqZaAafCK23JoifxsiUSFkwD3fNCNU610ORe
QXr6hgofOYFckcv3ym3wEg9qhidDTDFooaWQ4/rgVoCjM59zzIS+5XIDBtmA1txwaAVBqOoiWY7u
HmwP5pWd39IAIf3W49GMZCQfDD3SK8kSngtBeJOjeySxqCOZyElvTkMgKqHf7EVUfiMItB+3hOx1
1TGyhTiSZn4nNXTH3voX5IOh65MLsdyP9L88HZ4QBQOvKoUopoizNaWswEkGM4NmQ54a1WgL2Li2
eb8JmJHiBSo5RejhKDOjDe8u1Io5a8I/LofK24huv1mdM2xdP6UXhKeL032D6uMDth334SZhuz9Z
zzxA3zu4LcjxL/TC2vziURC0FCxLedzzyD7FLrsUEXRrsulP9egpYeERKv9jjv9Mea/1c2u1rK0Q
q8UYG6KKb3ySwjz761hP5KD6putj4hG8Eu6FdUh+82aFQxze/IEZW7YJTrgctHOJJ+uXsYiPpKyk
JxtBJfLoQC40ylnveCrMRCYIntWglLYNLGsba7kvLrnWMLkmMuTBq0QA6DwGDTIcF9ofohRFPWBL
6v3iVOGi9xGuc20so52yobMxhklaNPo/vTzVdP+cNTvbxxPFXGzYNOKD/59pdzkZWywLW34a7Nyf
V+GChmmtmcmKSPqkKG41F09eQIU2ZbMh0Gp+Bffqfd+efcCiTaesvetlwifIslnSpPbgPpUJdwf+
+eflreMiRySZUapANBLQ8vyiNZjVG3dZpcgrVSDdk4CC6jXmYNLN5pIiZXDQ4bIZowmsRd4+ny3V
mZiND3/fVnnCxQqgBmqJFoMcd0Cxn3GA8Gk1vrI0u9NaM6da/3BcS1AZbj2mypLHbYv5hXv0bSYh
bRCn3vZbeF/SZRCDoHK6U6gGj+A8dQ5XH6IPaed0WRWmYf/dV2yigYsbviYXhCWJK938iLaP07/b
OTgQp5v99xQLDy+WMplysCjr0FuRz5LOR5Qpy7rwH4EDn3aOdEUT3axtnuX9hHlEFS7cAnpOduvM
zYDKF8onMNx9hEhzKQVPvVgJZUDBhJlZ71MDS5gFoXpkhgUl99pNlkpSa4ASg+ul7KcNstU8OTgc
tTSOqzcYWzt7ConSmXHKfkUtyNa5e+7adK6YNjeCmV0QJzMzpNSp5IGEdL4weEl7e6kwJMPXnseQ
z4Mc4Ahey02iQ13V4P7+jU+zGEj62Hqdsw3n64nLjprOqb9iaaDAGO/WzKHBpEMvdoacZFsdN0gm
wpk/eBnYAaeKVclWMoLXUh0BELCoYG0PdbZ7xpFUGvzdBS7ieTmZ0e+vo14Tqnay/9xhFMAQ3kYB
M0srjVTTKqBfHFB4FjFJ0pYZsQ3WLRhGcRLja0q1mq+jwgc/mRYT8OKtMCKwEF8lmgG9wpnfFNjt
55QxcyUpGqhXXhuzLvZUuMeYTOwiEfmVTKSTb2DblytfEQiWYfE74ASzdvD/RP73Nba5VAI37OrT
E3fakChrf62JgAKqF1jfgZMkGe0VSq28GbbZODkANY4csMI/w+/mmlcNEqp7BHv+OQAV+LT6mXbb
ZnSwBuBNG9qxCytizLt4J3focPdM8FRLEpfM29CKcPi11lvAbINNg+RphKSMf0t9+efC0ozhRc1P
oZjgBbKFQy2FyLozJhai6AbDDt3+YDkN8TTVZ0iBqp5ihaSu5J6YQsLS4w+uC1tTQZTY1mLoVGR0
AJdyWB2lIrdvEl23ijKVxsMCbZ1RmhUezh/RDVcoZFdor7guK/apzFjsqRebOk+olbeHmGT+eIAF
qaENNk94DlaRFeZm9gWw9/KByeaBJioycMFjeFT1v7Geep8xVCud2qPsVxBCHWrGK+1mgrb3PQGI
78xOVy9Rn6ooetGpDk9Y8ob64LtiXypstv3gTNnMvhrOrJOLDH8GuTvZIniEk/XbOXLLMbSoxTb8
MZb76nAPHVp1fCYYEpvOsbzI2Tf8fz6szIPi2iSdVobr29HJrJQRcM+0gsjU5T1+Ps92PoYMlIBt
uPgcb8Nt2zeubfnNG7QsnNzobMll8Z/0NHbPd6ezK9PkuFEkAKjAF8Yl9foWzDsk8eO93K/7iQmP
UhMrX2eNwmIcNSlP9ES1e+mfAr1dn8BDeUDBV9+IpPgdv9QlyjixPZZdwt55ZW9WwyzHDtfbDrUA
p6pyrC3HumJN8Hs9b1CYWVJNj5ntSy1ocXhHwa2jh5CsY2laZtnjquhye5ZujMI929ldgxmiCY7+
yGSn759G9DJeua5vqnbwASE5/2V8Gjhzvv21/WgkCbnqoQmdLGKghRdsB9hsd1h/H54LV7qqkv0o
pSrxPgbmWB4cP4qtnwOah+Xnd0c8B2SGGDcjFidqnAimIxcZjDHU3bpMnU/XJxD+oeuycGe0UxqP
Pibeq6hAcwIhG+ihwddWldycHg1W790RHnndLmdlywTIxKs/BwpfOGeec+oySRPKll32JZvlE6ET
dwYEM264m8+QWgwWSGgaNAaZIuKDb/uFmi6T/FcRrVOmUKfi0tZtA+adm9Ge8sXCogw/PHK+gaGx
DQJAZvYmqOQZQ2R9UnOGwG2SjHAGLNFzTC0er40sBH04Dk7AncsCyAXlwDHnFAGZ+hurwetXXUFh
vItwpUJhpRyHEjJ5ffBZygCfFb4/cAO/5OHGYG41AWJNJYgIJ0OUbwSpE/gFERlYmNctPEvjgJbb
NhELiIXwchp7rvXPP1YBw2rMqUCtns1bHQm63bD2zN5bmgmF2NVfX2YG8kbk3gupCZB78PX/3Cci
rY/vrREzBIpZ7WfQyElnz4ajKvn7rhWx9lns0t2GFfLOiva71Vj3mLRAA2ztQI0U8pBrCJg3nA58
yjVBY3L4cUVGVw/ejTsq0wTJAhY0Q4c+OoSXxp0+lnWPdJQ7jgkUO03R7hH3wQjty8KC30iyfVJq
rFzfHJdLnvM95kb+fEorNwBCpMu3QDS2cnQRToywhjxPUZjMP3Tm4Nl35l5fP4We9FBlcW0qU853
2TjguFRi3mEUrGqCegsO47GpU/uN6bVkI1ngVBvrMTQ57FDVJREXodiRW88ASUamvtX11nkOysnY
nWbvT7o0gSRhzoXiOrPcn+yqBiM1/czGSv7TbTafriV3BVKX4ny24BL3CT2y7D4IsUF4k2GLSBXV
EWYwEwZGWI7rneDU3Pn/jWjOX0kcZSFz60pI/otiFaJK1tBdW3y4hUuVVYwa0tHz2wFcEZeHJXcC
8EuC0z6oNN+mM7wGLfWrVt12FpB46NM7bMCh5UytYXSQ063SXOJKBqaUWomSY9D7lr1y5fvDItI3
OVuSHUtRtJ87LzHK2Zbh5vsA9niuirO7PNczfTAaQ81Qe0Y9RWUBuJA1wZoB3Fth+/+/Ts1M7zH0
Pux6k9/QzcZKaDsXbMnEcgyrY2G6urs87FEVVQWlDABla+Xea0Fpdtw8BDHafZX7rZFJsMINmNHD
dQTaM6bA37xzONaXTfhMWlsJhh9dqvI+JKotq2FR+JLJAp8h2p9Hrtc1VPYQskvshq8a0hqkkTMW
Yk11vcIAGn4CY2zRxZUx8L0QG8A0zBptgDaKNq3fs0BE2jLkxkI8rPLqtXR6fcHfBH7x+oI7bx9q
ewbPEH7wjDFnSRfcCCnJ5Sdtqqcv817+tHzHlcW0Ak0ssRWbLww0bUA6xU38iCJaTBtvuW10miJI
yobCA+xekzModbLrLtP6O2tb6PfT2F0i6kt/qTh7Dmx4AD1UNnMA0maUWLoFIC6pIvzePHKOhjOc
qe6gDuHciYw8saRi4wG41N0fYka8KnX8r4Jrw9nhjiATvnrNoB6qeiByKauTgz/1jsUWgr68mp5j
0EX4bUfcmzmMLI86RpAcpJ064leXCSFdqEc7FSnhccj5w9QbxSDnoTsCiborKhXhREYM70DrFHDP
EMCD3jreAeItAnMitQbj4C0EJ0F/FmigcgXLWFkN5Ax8sYbMHqTiOSoqG1cWmuQiQZTui4jlTkEz
ZLdC+mpzXCxZUOSjwZWd/PKIXN6MJMgSVAKE4K5bRAbBq2CO9ihJRiWEv46rGnFYtZiZQ4zxWL//
OUmvUVS/qqWBmyb7aoRhN0tLrmV5kA810MDL2gKxBqCOK4Yp1yiW8PbfHDt9xivnURRv8fk5dOB6
mYmM4mhYsdWrTdeck0ZQt2lVfiXdP2VLHPZ19UbQ31gCGNmbW6GVDySsr/mg8aztSzKy4HaD3wpo
dgqbXNx/kGe8bpy8cDJbDyI5SIO0HlLXjV6o0hkAtie2aH7AEbjp1KrrTWxad2NHdqdqm6HjcwGe
rJGUOqGQ/503W7YmJYlKUVvUZfb9euclPu9PWBsvm23UVQL5wxO2EsogHVLnHOv28TCjHS0xqB6I
+VxpjhwFFOt3d6FdfSfezxKYObciNzyfu07ZnoGEzCDN9IsNuHtW5hg8Bd2NG8L7GJp57bnKvsRP
UoYNr6NZqYubqk+xp+Ad5wasAta1u6uSYkcdwq0aiDnIpZjGlGUgqZT1QYRwIGikWXAnwUtnZyrF
qQ3sq0vXuyfLGNE4JmUrRuk/3l0NiSx5TDGOlBnQb0EaTBXSFmOnkZy/fSGPxMhv0Gow9TX5MLhp
TCs2h79JTUIIZreipRr0D5kGp97C4+j1LiB3FnBt4curnSzizNmGtrgVvtj4be8b2S5rA68aFROS
f3rqzw/ywpIpKorxhFOj8qJDu16Y2iTMBv0MqIUlw4Osc01ec5eNfP9eQLZzKHbShyCn8/lsnd5D
63kPXBi46RP0S7g/Bl5qJ5fa9G9PXl6V35bbSZiOFL56GEzfqs3st9KFRUMRW8gkx0zAHwpHHghh
etTVSxO6gmEChNIgLUYQ1gH7L0KdXA3WoeIph38UKvkW/qhuYzmxbEeRSsXaWJxmnd+ACBqAQFoj
GTCJrWVXYyxEmUDmSLekyLIFcsnwYqEqV6f/G4fjjI059NJqEEkEOCOpbupvyzCfA+cMeI+dbNKH
S5NR6EqEVeCoBeDUseRdoIP5eMcskfuS9yl1/qDztquYhCfTdb4XvuAVKwTXoThYWdVBQe8weerR
3uBqO4+Zma+RtvR56wMpT50sSzBwc/SlXnTht+HzMHFAyOeTwjHN6n9B17s3y3WIC0mfTQGBF2A+
xAbkty3xUf/BeIiT6oLkyzPecNw2F3dRZhaZPJxS5wwiVYe34kBPy02f0BrYMpmtXpi+3dcYxs7o
W5zC43mbpIEEtSO/lx/2HOdOU5DjARQdXQ0c10hUWsPasdDAE+qabFGvH2xlkfrxP7hb223NyNNH
9tttLS1RuP/pL6E+IOtchqnd2vnPIOI094zMkW6a8sryQfgl/kCYdmAgqH1lQy1HRkIM2BcDAER1
z8rv/z/nh5iVexalDKdSqscuO8eC/B86BoR30fADq+pU2qC7017nPuGL9fVbwYePWgjSFgc9U2ex
yBAajQOuch2mpmU+wEsIPcIKKlkI0VnxYCbpqjbClEbuRKtSgsvX9t4zVEpC5I2iQ52FHoqz+gpz
Appsq+bAtW0Q6cbXns6o2J51gK01dSoUe4/t04ufUVcH0cLCfbgVYIBIrf+tfGBB/edM5zZY1TNg
ua3bJaBn0sH4hJRAmZNwTxyz6G1RWjOmOqfjupVGsUomPw8De66ERDuWGspxQU4R212BpL4mKIt6
YXAmPTpaYaGQWP2U1Xkksa0/iqut9bNboI8h8gcR59kgcGalYU79f8hDX9vsXwh+9rotzjFD60HR
9dKoDmq7KGF7g5yU0VVgyF5c6S3Q9RzNfaGXaz8afsHoe9zIcIIO409zANY+thGTWX9LmXteyISK
iMoCAsL3wRQ3ZHGWwxLByC8eO/YxmMbRN0KydixDDhXT+2OcFKdQ3YEB47bdgzCNCgxiv9TUzb4j
ztaGwqJqz15fbeq+oV+7H+/VZrktEEadNl+OXYS6OZWKy2UTb5xtoBy0z0FK6zBoxvzo2nqeo43f
MG4Dz3pYsHP8LbTH2EGLtEMaM/EhXMfJOGvf2N2h+27bS04Mf3fiKxTBvjAkBbkTlbPYSB5udDUZ
D1VveazBd+F/LEtFjMRzcesst5wgKxcb//fXT3lgNIPXN00A4I/y4mWRSIkEcXo4a+Ux8917OzVY
cT0tlJb2xcCsf9q5oBHpeiYHAB7Q+A4cgoTx5Umt+vbPQCv6OjpHlcsTd//l4mDgSttzJMDWckxU
4Msn3kOZ1zbtOH68oSQ0SsD1iMg6Z6IXio3gMAWSiMnfIpRfhzduw9UJgM9YdbrDMwmon9XsZVSR
9Ks5s8Ube/kYfytA0MtknAXQe/MoeF3gZBKoaUdRPT90WpQxbI0zLOkCGhCuv48ohr8ou58AjkoS
3b6gdfYKCY77eWixWfkCD/UfzCzoupu5SUrvj7+8LZNXfFGBES0DDHJ4ktDAL5ESQ6UjCVyBQ3er
d5R8D35ZCgo8UagIiW5b+p3NO6Y/EHrkzLDx+zPUu/aWlPxLJLzvAAXhM/NDGzVP0yGSf+zgvAiY
ANqfEgp7uyCb9Egj4zXQ47xMp9JUbU4UMKKWo2yZZRZHG3Q04FTlHvj0xT6TBCGCK9aPMRMtp9v1
v2FqiU4ubWdD9WXhF1iOV2H2f+t9YqJoto2cMf1zOF7O3J9xNYmtyLFNgZgA/BA3I3wjP1PWTiTb
9As9ayurDpWnQBvYy7JkhIjBByjqHsglCCOpXVNSF8ihGNfBcMxuzufmhlNXr9k1m2k/FpWfHNK9
JEKLMa36F3Nm+AUWwHrSm1TlhUUihrcplUJMoaGqyOydzhtyng14qoJBgiA7Srn065CRbqFHFd3x
uudxIvPVJU9q+ZVPrznrDC9echYQ/EeHoVsP8CJUeTIlXKu3QPRCim9M+rpTB4DsBzappb2x2eSl
Hsqd8Sk9YTnOhd8O7jRpOmQavWFdGPz4dea6GS3zXGMMA0uZFpHxfrAkeHHEIBM6rWeBK35bIcbP
7S4TUMACnzX35akB/xDDNjMVldmvzT/VMi+R/Q+SCDP80OM1aag4Apvngu/CJuGFIKNYwMA04EIP
RdMLWvWmZAeeI5DqK3znamCyL+CDw/18oyTsW9TdidgYpG9FrVRRDbOpTU1wZH09tsLyaTMk5uFa
o1RI/DnsQUbPvzIqWB+kKkZgFgpZtyPvqrzGg1iyx5qTStG3D/l8I+bfYQJL1QcQ/WLG1A5lgB51
KD/pg0HxRiFFbE5vXSsfqwKaN45q/Ja5qFh1nBHAVcm8pkUpNb06+adoiqvpESQtul11ggayH4Ep
XrVC2ADUtG3qwPfm/vysstljDnk04F1Q3uIsNEnzo1zMJn1qvVg3whHaGdTyG6991chIQElciniq
o3Mo9vdoWWkj1fIdBm+WmsGEFkRdQN71FQ1PoIF4UNUNdbOnIs3fq+u7hqAwsnis5oTU977nzrB0
0Rx5bMRT7j+Xz5cXs03lZTS8N2CSDkM/9NjpJrJEWFWwj5OqFAm0UFmQFODcdO5MAX8anamsIljV
j6KCPa8OpWrJyR6BZNeupzt6qD1YVy4WbfkJZYHl2egw3KQH+ZEyToARP9kog+nfIy1ynkhS5oPI
cyOGg9jEKJ+iS5LSBUOsrJoOq18qdq/jSrsSrxwlqwtqzicH6nergIpxAypOklbdkr3cg0+Jm4vb
J2M/BAEwd4OtZi7kCx3aXiSTxEVkiEeKp+L8nrpvQH7cMCoA8JcmoDOkKiLdR7R/6tSJF6V/h8d5
k6xIC8m/0FoVfPOaFdElNHmfJ8HaFe9WkyYOhGS2iB/MFXQkbURhDDpO4RDIJkZ9ia0gf29qCzZ/
oCQEwr9V3EugAVWzsRAlZ2cK1OJibqREzS3/JJ1DH67CCR0xQbsO8mGUeiqo/NstfG8ZK7wz4zk7
ROe5SwxAFqUsnxij7mQf9gsMXICldzzMusU+qCvt2ere8fSWDscn4nutmhfU0t6TScF4N93CMPeo
h+3ppcRJuGUvoQrNWw96LXQ6kk2UDAwxU2Vot9OuCJgrNA1o8APzdq2vKmAchjgDx+T3jKppqx58
BO4Vi775KPBqp/44eCLdYcW9T7Km7Q/o7LcYGFEBKNs3BiDDY3BKB3D61Mw3yfxd35qN7HizZG3v
g8EGciGNzqfkbXmVC+9Z8/st9joPoFQ50Nz/IoQ5n2196cQOpbP+f1JZVo5Z6K1e4LfaWEF2Nk30
TOG/REModxL5Ga9rnntSxRsFHfJSEpesZUPjrNN+tTsDhFAOaYhHwOzSPqOUFVwesT4u1jGjUsWj
F83IwhhCouNAuk5f77ev6t8Hga630G0MiKN4yiU//b6hWLPA1JbDgCT881bblLo+HXiwucdC1zpq
T3ZgYyWcM5rPClDwxqcMHAWZW7uDkfJZ8I0TWoQ/JyIM0qz2W09Ywoyv/F+s4baan7Et2QWyWoRy
BL3aFH0V8DuDQBuv78N2zeJfJLhVnVE/fOz+GwnUtuUl+lUDFm3B/eVYBVkz36tdNPeUDZorWce/
Ur+nhOcVHNqTNlJwik40Rz1LDZvEafse89jE/TqJXAbGpnEJnSyynF8PRVwgQfb/HBhsUn6PALB8
pnErmFRYb7zZNuBIegw79Wm2G7jUPRWHdXbUPn5PDLg00a5YYy3ZJ+lJh8cbnA4RUgHH/NvetGl7
XoP2q9ByLhA7QhDPH0jf5mGJBJbtFi84R9EMYs04HRsa+T/2g41nmtl6U2/vkjYvEsHKYuCRlge3
+bTNWlpsq+6VJ2YUZTBD5+Jw5IsBOIIUpwjoDFR4d+3YRqJ7/9lmIqfxaS6ZXNaI+IW3T5QpsGe7
edBtvcX5DrjiD1vYNZ6EzA0KBBQm0UOqCKUVLkMzuD0l2b9fR+E/oM9eHTi4L1lTmcnB+ZMOEI5g
wFXlfKTi1bqybl0AgDOovbrU0mKoik23odzKoTjCmDIpogPPgFd3VkpfKhoTghHN+BjCHs3m1+I6
Uq5M/o+ry3ngqIAWDPOttq+JNEgbhHHe2XLnhL6MNpsQImeW4HRen1PdLC5DrXFkRxdFkwZqwswS
CqAG+QcMZVjLzxZkwFi7TM71BjoiHgiWKuNojnVDiMe09zm33GrEYYLohb4omP1n7Ek/ghyvejMg
uHJetk7xMJYHOakulvEQGxT5id+Rcnchpy85W9pGcLMbqfbZ3KDga++oXnh7UTJAMC+/AaCcQFTA
qfSA64loCUC2IwXe58ztw2r7vBhuWjyV8qACVaC6IPAPVW6RwUioVws8gpFMTTEde4DBXuqGjfF6
lsZ3uqHvYwiaK8T7Y0p9C2/+EjVsvbsr7QRQdCFdpY6nxnZqQmplWCRRafBTnyaaehE3ZRRMB6cz
W6Zn86WCv+Vzd4GGaBnYA3uChT3Ejm8e9kl8WH3ZcQ8iMA9DhuN3Upjeu9fz6VSB3NPAs9KR3f8v
pO6TtTZcn2eLkafALPItNpIjBgsWPXWVfx0dzsnSOde09D/EPQ31OQ6I5KcDoch2J4qpHMmWdqov
wcBIH6jFiTfLXioIl5gkykSpcf9zSWorvKnSJWUUF4BPVJ3dj/FHdHUSsKHc1b8v6qjevOE2ItrA
vD3HgAZaZcwCohMC0vhS+x+0oZpqmPvbcsvxWZHofg3I/IaBINrFoYs3wAzF4/ov00DMMbL/JNBV
PZQp1Ky6E1WweChKjnbFHTTQR4ofEU9G3rQl9WkSr6APvuDNqTjIHd7mjMad4c5vztDhtes5Oq2P
KzuG3F/24R/kjtMt18jikw6MRzmUSJE3qDjy/0pFmb+85CinLIchNbuYZxTKHE9nSxxieYsz1Ozi
e3WgXSgNCnfwYYO1+dlVaMdQqWaaRJ5Ef31rkVIQiLyWiCnuSiUqD4a78l/qROdB6O2tM3NjiEeq
R/TwEVjxEffcnowCNqa/gDfmGm8kvP/uHtQEmwzrTSVK8EOFshaHtmlPY04mp77kh8aa8R1dbJBc
Pjci9F1nZ1E/TdEh+jCsaI+OSg5/hhUHWLryTwWRfljChzG8/dubT9XI/eogJBhKh7IXh7irj2ZN
pGl716UfwURsOdUMhH4ageZOBeoqWN+yCXS7RcqcO4yhjYUTTGSOh8hZzRI5iZDrGV8Zy2QLAuV+
5FFVxQIxvxbkbJDL4G+giVGX/XSLO3jUl3MDHpVnt4BNQeO+r++LG2Ht8At/7N2C0hFmWXeRom+o
wvFXD/ggY9Ya5XdJYkmESb5hurJFBE2rmRWy+rYy2LgtCYIlOAZbBYPruyvhfQ6tMiQkIaiSONlB
BCAaRLU3Vtui1FlcgR1Yq9Z5i8eYyartecB8ueYm1Pu24ZG0R9rZnL8JLPHSsPBHpt4XBJAXLQtF
URDZVcHIJKsmef0gbLE3x0GNS6VoWTGQHjHef98fbZCKBiki7tZTFCiCdZe9LoqM25tYBWNArecV
H0d4Sgt/fDVebaXlrSjiLuIUZN6be/l+OIGjRpKVcNAGwGoBhsda64TxyL7WLPtt/XKXr2FU5Yx8
qVzhv6REmk5KEtVUY7isINPUFRmW+42TCgG47UH9gf1ikBFldv6qsIfnY387YNjTnKij+S8PVEB6
ldDCs1Y0Xs5/lD9LZSnUU+NWFI/kj6L4hppGd7+te+czKMMGwZOkiSfq4h0Tlpe68JhdAHBZ6jtx
i7qOzMSaLX7idM4o6WCXR4B2n76NkPAHFa4Sd/bfzNMDvITBJq0jWU1S1Qxz+IGdWbP12TP/EGWf
BoGNHie7SkAttsPhXeudktd7OOIbVx8HrJ41yYL+pA+O+X9pBFd8SPO9dgbici4brlHYeHAXdLEa
Puf03wfMb2AkI3BrcYA21/T9cGFcOFSVmw+joNWGX5nw4/rO9zKdazMa5IdvL9itm7c3+qAvO7bS
8suecPljTlVBAIKuBoaH1AjAVUC6c1WJkRpt6cIv66iJHIAN7HpHbgfzjVjHYhtsgkjcJS4nvkIB
QvXC/ykGdFXOAHDWOzxHb78l+J33yXGHLh49btNhFOrZiRaW8QhfX9L5kLaDu3M9WCDbf4Ij1A5Y
YLsSheMcBEbnz7/uKJmZ09/BpuKQIzSXx/4R6szP5f4+dRfuMsMIH7W9t+eeXllDMq3eDFsEeK7N
RmRZOMsCxCu8LHv907kXWdA9UR+P3yFrgIalCSExXEsmU4fAMIBGloXHhaGt48DFeyblicxgRsXx
P/qmBs5xsfeGqZr6i15+O7wMF86Bg7Oa15ygGzGIr52lorVQt75xmu4hVf19OpEAVQl8cU76jZk4
VBdov+mT0EvuhI1D2Urk83pzqfp+tFTzNCdBk7xrsKyw5AEYHwAAGOzTL6zVU6FA6yrsjAvxcdpc
jmlrHm9nTtFliJgAEZmeJ6x00Q2d78S7LRKpuuY5hFuVnF7P6szdNNpgCK4OAlrEYJ22XKcFAM/Z
qzp60zCJ26sa4XSMpjR1l235dqfPUburntcfE7NWVZ10ygPzEoR2CWoROBhnHonOqB5W3yMY6wYo
ke5tIL0VEp0U+zCj667ySrv8vjDW+CTFsOUEdiHE/YK9WKG5T1knGGKBs7Q6y6r1+7Frqasi+Ohx
bxPqoXSpFjSOIblh5VMNYSMnQ/kBqmLyv+oBSo1fkGXBgr0PPQwL6qoBHUUqEIk7kbuohwT0qWct
yYSSMz/FrKVq3OHebe+6ngaDsqlgP5kuKyIO9894xP8ozfL4Ta+eXiwfUAEtFue+2vwc+cUkmv20
OQ5yn7wCG4OqAIx+WiAeV47kwBC6a1y+fGDAX0h/9vhQIII888mFMKAwkpKvOr86Sz4d6JlYGdhQ
dYfW9d7q1XzywqHZyz95cZ5FMuLfBHmDFtIvDx+H+MlQgfGL9Zi7ItuXb18Q/lBURP8yxVxbysIe
6aYJFsZYMRQ9pDdfwqH0f+Vrqp1P/5u1ug2bALAhVHP0Oao7CZgAB1ZXxRQNCGxSh4zTSZ1ocVKG
e8lcc3mMdopp1/biEwoY1cjGzFcYalMjAVL5u3Uz2xWVeNTd7ZVt5xSAO3rZSf6z+zgxXIDXuIGf
YMltfcAIb2jQ3awt+UG2l4M83FhTcIUF/+fYnsu1XNxWAzL14BHDCvEhubAxsvTgRSebHTNROxsj
+tW9KwTXagGHvt74jyee6SakohXyMvIrRbWBplgsaEpknl0RO/hIMh7EI6OJyeTh0CInVn4QjI3U
S/04USJXz43g/JnnmOGPlnma5b5nWBpw61hUJoPfepeW11GgvuCoelTGUYWa6zBwKQ+/enBIJvVy
8Um7h5r+UhSYhz5STxCAdTimLMPyRyXkMgbW3caZxe9NUedPQ0HjwTlZILJDYSCOo5v1SwcGvPRR
Q2DRGccOpj7+RhJd9mfQNH67n+JLx4dQAXZjlmF7e9lRi/SEoR6FF5IFhWVpinkQfRCPwPppjslK
vzN+40Cg/51kcKoBR+UMbrbESiL6yDMsyPWR9qnByhwWg/TpZ7wWoKsTlQh2aqREnNJeZ3dsvnHE
OKedt2/cBHEY+Q2SRlGUEjvIv5mCMLl+gdABx0B6JrlKaWz6eK7Knp05xJYCRWAyPUd071/dRWev
svoflvJRay+pODAbri7cRpcTrM47YJpNT5NxA2lle5hEiV882eH3jUrld1jeTv6PDBmzXEJZLysT
9CO9nd5vSvEaI6vIqBD5sIOslRhSXIlQTiacbn64ruuAqz6FnaBW5gM9A3cWYr6vuV/6ENB8ySfj
Q9UrRBcSf+S2kZPKhgraGotdYFTOYwAqpEVQ1J+e0nUHzwPdn4kruujoTkne3aq3Iag2dab2LFMJ
FPV7hMNZGKCEUdy3oPSOQiE+zZLJrbjxRx/ZOJWBTPkCaf0qWDMpOXE9O/aqKSDBfNStVj01EhkD
4/XSrao0Hargv8e2BtHp42qZaNu1la8PZR32psM5rzHCxcrSgQpqcICYi6zIZjs79xBk5fnEMVdS
YP+NDUTmGUyC41TxjhRLj08BVkOcpKiT4PWGLlajeWkpEpWzXgwd/LYvH9TcEzT1MFj2Kvk+Z4iT
EJWUHVwAiNizZVJXKnpgi6gCAowAonOIIew6HQo5E1PWzajahGRkgXe3CAjSed6XoZnlqSwB7fri
mh6V7ZgewznLpLkW2VmfCRgCs3/n7UilleJY2dESHFiCkARR+h6SAIqpq+IxA0wYLUcQxX/cwdbM
cy7T6m9e7iFUKtkZt4KaAxY3ctb6ZJy4n2U943R8gThWyYW84JAq2N/XuodXmVaIvc8yj6PYJ0TG
5/xQh7ZeXoP1tyjL8zyU8KRL1MnOsjuuhTCTggE6Ixv6GcDR9cPgf+wZGEnB487trvuIBm78IA6D
qsVnDs6QNCXHw5cYj1GpFxThRR7wW6l9h9NoB0zGTl5+3EM2NA4cG5TqVTfmY43sXvEJ1uyDZu6U
OFY7wmSXI1sbbcIv7c+JkS97oPmRFXw2Ijz2bjWbV8w0wOUFWOptUYvuahGGhPH7x+KrKRTdf9Yx
1YRfVvQHe+Vpf95icRCxhen5ZXDH18oZYa6mc+Tmg14M0Se8epZug1N4DUELKpLnzAxC7cESpAcj
5W+7UBp9SkCC2JMhXY/QEGMbCiOp/rtOzEL8iBCHxKD9qMimqQATHLHx7b6AMgkIfWvg3wUgE28H
MqrNAEqH322b5M6+ejty9NyRgdgwn0MfbKT/JTGjh54IokpEVu1b8zUZcy29dtBCcIgxoia3T3gK
c2hkCb1aEy2mOreUsX97esylc7SAduHBfpW7mvTwMQH7ZmaYDhqc7Vf4va9i6g8wXWDVBTS23GiB
mnNywe7lzzyyCFlOzMzi8zxGXcBMgU6zS41MfLdQgcVFwOpjXLKLHXLIMoyR0+s72AoM5RKr/EGD
Di5H3agsaLNUpouO54K3mkNqPu96VoVbRrQdGhyCjThYKPDtSJgxDBodRyglFHU56elqtXVVhq8K
DYeSKf57uiTfSRopsQFUtE/wOTG4tGygTokIvNVkCRV35feYCpx7xOIY3W/uhp1C8vdk/oT0h1EX
P0xuogbQO5wRfo/IcOUJtvanXWEA3N37m2/NV9n/EOTN5QsWqLm5h9blTsyoj7W7K/Pf+oLvB93Z
+w3ffcKPYLp4AJ5IXzx3tqYzrxYcdbYiCWG7gtBO8uXh7ThdVNDuv7L9iwJbWgSOkBpnqUgPDtvx
gDVTd4FVAId3drl8JjO3ZfdFzy2oqXVaBKc6Wu0ygBJTuPE4IlBRTqxGzTBPPPpnOUluwmIXqNxd
oocyYLbvpv//yQyNMIukQBjDE9Bsss/RCP1/lw1lI3HT5P8TrQ1L+XIWbqxmnPTfqJo5/du7FpeK
7MMyW3FmwX1BsF/ZG+AYfdDdYy2thWZnIiee1UO+8yeIwZHctnQaZFHV+JNWti5OnXr0LFZrcYf3
tUDOtEDPe4EA6kgrHPOvchbDP9r/8fxKSQ872GrBAtB+ybysKJRMZdsxQcYGx6J9EXm/0wqBaoqK
aMitfLxtlHfWprnFSvyxFTlLib9i90yILc9TzRnUPbtoWZ4J2ROGC0qCqlqjdkcmmw2DpMgdHT8m
kRK5YIep4hiClU2v1FXgAm/LtHptGEgO8VwXTBHeivtnzh0JxXifTo+Tsovu1MKECGbzdjXota/9
B6M6p69V9C6MURkUCO1tZFic3w3jCRXNfNi6DRR3DmdWc3yOkMrTqwkvEe6ttlsFHROdU4Kx+lBt
8otyRq/VahgvWsn4FtFeAIEoTfctG/MxLjq8LgyzhkQyIYk3NiNoeMLM7KKQpP+JtOysjwPUDI0p
iDlPshZIghyrV/7ksf7cCnvGGoIyvot6NhB50YFmVlPC2v7hcSl+imZ6K2Uyl4GIdTY6cXswlFug
fKJYqBjMpTiqzHvD3cDp98RAF2evrAdDt7flUfjqz7QjM+axd5wWoAdtFKGKgr53WKYJ+SRmn7Gi
5Cw8LbZ3Zqo/GAPD3WHyTD3+RHXq3FltN4uWD+IVHAUwvcMEAf4RyzWJdWoI7/jS8ytN5DYW+x42
xYzRmpkdsOw9/nTXMu5oozjWgUtKf0MPayvjL3fanoqyqLyPU0/xDa+Hh3OZzyBD1q01VvKBqZR8
nvr5vOrJ+9TwTFuCwVutUuNrCwP0XM5qv0OldvQH0seHjbrEOlFabaznlaQiFXKVAiJQpxKwsHTY
LWQfw60WBepHEzd7xnz9SrBCiyDmBFICnRl+YGTQnYCA+Si/WFreft2QB8+L8PFGcTbJJdnVXGje
hMUJbwkvlYU7rOOVRPQEVwS1Af062/AYBf14Zw/D9zFtgpQouIbPsUx7qbUibY3dAkJPibP+7AED
G1/aaZMVsHjngBylaHbjoxX689QusQHaPi2jrwvVst6KbsjVtBiZv+GDFjzOC2Lsae9cll1WKJ4W
9C5+X/lXGt8VEx5WgQdX3ACS7eK/Mtz38aXIDEQsbsUyaVA01k2QiiZ+D8WQ3KR2wmyri8SWLFm6
pAjdvvxQnmbj2K4QU6khaC3diA3ilLh/s6xtPIWbxBc64Lg9VFQrI8ZjnivW6jAyo4P5RVGzoVNd
jhbTx5jKnNwlackuYQFRteFDbp5AFb570a5GuUOpQRd7ThjBLbFZjgdzCYKcidGrok06gnzt+D6+
EZHFo/LYdrXH594fFVV87zNjOSbpGCVtI4xxgi9Q57jYt25uS6HVcC5woEYoFCNblVSMTz6vD3p8
N/Yx74kud6Zfo0FaSllLRD61N9qlHyYA0aZ0ajM+Qa0Ye8W1m1KWkRcHW6tfQp3o02qG0WebsYiU
rrQ05Kiid1/hOOZh6oS1DR3V1J9PigjL5rGY5LJh+oBBAFLhrKmH5TvBfAN8MwC+sU0xWrd6HetM
iyJpxKEyFN/0Hn5XKDsbT6f/25yPsoSPWkbJQ8w9Tg/OJCrKonFBIR/r49WXLrXjKTE0ZsCJpjVd
fugEtHWhnBapz7LiRLn4ZR7OaoKdJ3PNeTZ0bdhFrBHnD2ddxSPJNl9s5UNQO3wPcmoy/yzwfRE7
WUX83Xko2Jb0n6h1XYnZj2dFr+BwIE4FPtAUjvkaG3eCicAutVeSU+QJfRioYU6HIlod3KANEBv6
n9HlvP7/xzmPt2iO0qruANjiy+XBj+pwDf+LQOSBZnTVNHOkT+RXajeBYGSNQalHNoDUcPHCvk81
mQ06M3k77bwb5pc+OA1LG2yisvYXEJSHMA4Aa/7al19AQVlJTyM8gUyGNj3GEEQvXMh5Mt02sr9x
aHDPmEp8P/NNGMbj4V4bGIPFHxoxK6hMWI1ruPhVJgA0rpnV4SHzQbzlETtK+l+U/ZiqwH8mCgJZ
ExcE+TBwQ39wTXWSh37b4hCKMkMm1H6nTGRzUkwuDt66M/HBsVwu9CYyOe+1GeGJWH/l38RgfH2a
IurgiQ3JwkskBDkODNgf/HL/OaPOgWDu/TWh3KXyQwerkp4VQO/LitPQjc0Wei1IkpRSXFvfYmtj
ovhxahHPbIhIUEG1QDgR0L4K495R+LDiRWCdI6F7gVG846l7LmCfND7M93FGGM6w+Jm6+vL3WKzE
cP7aR6uXv6lbyP3IURgStgatWpoifl2jb6aOSqUL8sswkhbOlxFwkhGITiRGNlio9I89xadUgs2D
EOAHUiT18SwffPNsrxzUNA0oYOTVqIpy3yDGv8FRCHYd6w+P0YO/fFeS0IgXO56vcQk1kGe+USTH
REd+Th99LvFqtL+iFkAKrVjSlSJj89YXG2WaG6YqUX9gHuKH1+PyT/cnYh/HWuKhY/OAindJ9VTs
X3rZzIYXWaKYD/46CHBuxxLS3kKRA+sUZUsArBGI0aAZ883pNRumjk0GWpQ2qQ5+rS1NyHLyeq9A
BOB1nxA8Ahv9aKQTpDMXvJMN6VR/VlZRnyZdafa6QqYE2Y04aLQRymR4Q0SVfg1xxjqQj/XE435W
FJEWGN/79fUl+0YIqjPfuHxTfoBujwf3azhID4vs9/8uUXqR/pkBDUpXzczkPVzEKdiVEPNFNQzt
k7FhVq0H6ZVs+LDmukOdwKi9clk9KOz9kLxjT/jdChbc/fJ2Ih3v5EmbdGZ2qPJECf+jtOpRLrwr
jExOkoQ1kyxdcjAfzhuT/upTs3tO8WMydcEJRg9f1Tt9Vpfb4dkdq7gjeKorvhoNu0sRl1Rrzmsj
x8AFwcw4b0/rSSuXkRfyAMQKtuPcuhQsYcUgzAYcJ25dTRmN+n6AUCLBogIAITa+N3EQNHBeBzql
UX3MoIYrfrC5h6abHMEfnEcH96dZ4ESdvcTf6bQXBL3cBdkWMem1eEjT6Fl9vRcljQd94ztZFoRG
nm/ErUkxKxY9ia6Q9cVakPFAQnCO/HnCD2pKo7znuU0kBw7v1/RlKkeqcyOQqQjXhUpLvbSmYMV0
eBH/ps0J4ANNXam5HBzykThW7rOjtIpHU5TmDToMbCT+41eW2F+INSurgUEZ25P7Q4UlD7McLxIr
Curhk0Wyli3/KG1fESb+/MbXRCNZbg97vJvUvKJg7OrL94aV8vCp+mI5C12TZjISPVNuareimYM3
F3cjHKiQYAjsK6pmLnDu8vLAXFSjLE5Zeu8DxEnqzzlrS1TinY7yOzJu2dIdMQwtyQgCByA/HH1k
2rhzxpijmAElHB8yOQNykxRanGLmvYWfgizBiVyU3crZTtAJn1QsWKB9gGOdL95C4b9cDB/Ch1HZ
7j7OtmJXBdnzrYqgAJo4yMCirkzIcbZkgGIurGpKAygwp5aWpnesx1JmR4c2/H69EhFFv+43hiNM
v1JRFhMFGF3g3/85ypVFAQRTKztCmqTIqz84lC86YCOrbDOR3i5zITegu97wjMWfbvSvwdJGpC8i
43EpgjuQVTCj/oexxa4WFBQJ2okU/PSnF9kRuEaHkRrq+a5eT1I7zQaFQ3jfOX5KIDJp16S40AX4
T3L0hTynIQsDrQbK+2njy9b3PWvvS3whvs3kZU2mR3Zv9nuXuzuEaPRIUf0wlcLYztHnuJaRZK1c
NaZx7jbk6RfVUIOwFwNkxQMcZCzyrheTjB9dRpbBsGrkO2nxeTzubi0drm6MiAZveAOe0HDkmCD8
J8kwB7Fr8gXMjtmX88gRGX1RAOwMEZ9qZfKwZuXhny0dAnb8VjZ9NuuTgPdUvE7JNLh1AUrWQh37
kFcJEEL1sgkaQvoUlNI7lVPDg5hxja8RCORla7OlKS3njG5Fo4jDdr6gTSTlWal4CJeN6u4ysrEo
CX1h1RXwwOEkIoP3sRqwPqwYtbf/XYI8IF0vQFRNa36FD7IkZcTGSuVZ2BKlUqT8DHSF4aZaNMkt
iuVcyyLKJHfnoTIuGEVFDV1//ASfR+92cr4uYETb/on/amzvd572i+ixNr7d7yS1mPBkTsUeuS1d
sGolx8pR4AELqRJFpVtWgn1VGo59m5y+7+lQjYcuVfWZY+/zNoialZyX4PRGRim3M9YnOak/3ucc
LhR7IGsqGtgEE/9LekK/Ofo5EDx+sGCbw0YPkW4r/193kd81YYqxILmF8gCY3CBL22LHuCWGsbgy
O4ZP6dZV4lfgGhlYlrV3sHDMWaDacLML5wRW9lAq6xJJSvFnOOLxg3ppGQ/BUPDEQVAkzCUumkRa
awIgaB0i8iPucOlon2WUf7br/EOuqtTDL/LPtXZ8u65dB/IW5iImYUdmGmTKuVBhOWv6E6Fq8Eg/
cc7JoL5ep2PP+QhRf9s2bpuuSRcFhsLMsg8l6JWYs93RVMfhXy06mY48NKnPNzC2g9iPd1b2CWxt
C5lMJHhDj0v78xmj3yjOmz+he6DoUJujuSIrGBi4roRaKXmo9CQLhjFM4Oz9VuAA+OM+kfZ4mZc+
AVcklu5W5pMp2nRydRsJzDary2w2eFX0SkK9EUgRuFurG4OgTWWHKKA3E7MXidW5DfDblhl2HP/+
QLdSQX7B1a1QGESti3cUe956ba2X6JBlsz8ECb6D+0HDesvTj4p5E3b/1DyorZJBORdqY3xadBHY
ZpHG/Lm6UFYVPxK1hqqz2EYIjYWtt7cY6fQj1iuHyByXOuYyk1jcp6ykSTKBCJIfR06KJHthKLNH
T8ytOFU7TQQBNlik0A1H8BkVmFd0aPt3Pn0RUO8PstOoXCJMNS1snYc5ADwbg7uJLgpYjfY+Ioyy
ZCH7+IWH2t6uc/haz2Ru9dY6UGNweWSEsGD5zfdBEG4qON+/JBZet3fbMvWQ2mhlxuVxJROo2o1H
pzqx2X6TzUdsjFtS9/81EkRozjx5qwKBn1XUiJGOAAB7D5gwgFu0NfB0OHhmL9V1vV+gZKuJrdFg
/ncx1gvbCf3zKG6UIbjzyzppIsG2VYSpNvLK6TKazCTYcXXc8v1vOKK8I1PdiV5jopWo9R2FNixP
/DXGfpsE/KIWDqJgs8EHtPzOOhXU+hH8FK5VvkjXit/NPHp2UIk+VKTJGstu+koMD7nynbzTNINp
LAjEEdna4JT4vZiPHTTPbTP80iavie3FdTUMowSGIMuzfkNy18fCD5BDvHGjCdPW6+hTSGYNiU35
98z/Sl1P/mlAT2LIXs33uSKm2b6/VGazGj9y60KfLjONj53b3kEoqT5cta0JQo82v8CphibSS2zQ
I7cmHDZIeZbuMtC1/DrS5htbFaRYWkKDfgLSa3rBa6k6c9MZ3qOU6FkeNCJ79BnAN9MDDvaginDx
EoMpzriwYMxQbrqIunpi6WdDLOvY8VIu1YXh3HB1Lk8MxaDrw9hKigZnbKcE44QBx6clZ2/pzNgC
ypyEAYHQYMFbVR2mN6o0644GFd88Uv0d49kinhTFPHpZ4xZko5HbgMLxGyOxOq4OpsowzFXb/KeB
IcITskJ5owPSnhU/5/aXBtWyBouNW6uzjd4/joFKBxkobuGcH/qfSkdPDXO2XVZWOdu1wQiDyI2H
nabrt8eWLvrJL1HHksO+owICeCAQ4aeEZR70XHsJeWmYVSz5BpXTHgg02iVdNIKkcqLBDSGZ6eui
A7EEB6Flad3KoNyZjYc6FARcQgqQ5FXDps2e6PH8AT//XIKkVHVuNu+FjEJcSZNA91JiFAeULZPW
bm4Hi7a3R40gkhtdWC/CHSPXrMekilyBl5I6LPPML5pbkBYzht6DxY05QdfjOogeQIzWJFE3J9AK
LMpuRSAvm4jGj1IxoJY5lmOWyTvuY1znZrFQh2fZJ0oUTDfXu6BA+9K2VTe/y6LfnoeqqJ28BK8c
ITk/AKTtyIREfkdLT88b1a4FHXaXuqqG9aNbDovTK/8DE4gcjIzLoK9gg26AlBEza9pzLHVeV0zo
NFHbfBMaqIYKG1HVcDoukeeQx4o4ebJSEhDKQMLeZCDqQOdwlAUmWMFiNBkbNcJ8nTIE/czquyvo
3jAbxZ2/H66MYT8CjOHmW5EBJU3lPItWxlLSTIqrwYvSOeYJyTvcDWryEbKTL72qprFZGQim+JSu
YV0JIL6s3I2XqCt8izGBsDQx6i2stx16cgp9qeDNeCZPoDXEbUxGkxTH/00/N6nN8ym/5oA8Az53
kDNWTj0SfyLopY3OB8yZD2y4JilfxnZQsretmOSfVVz+2EO1kOnUrWh2YHJvTFX1Gn2+HnYPyDeS
mUAk/ULquWqrEELtke5VGhCNSNZxkSW74umtCihSa5haw9WEvDPeSH7lgqV1SZaFxTD2WHDqAzwV
NBwqX4rq/mVFfJWGP4pA6HHSRnhMGMw8JeDviTNZFwX2qAe+Y6Mce76m4i91KGVNOxRFWmxL44sQ
cxnUWzZ6pyBrffwLsHUQ61UC7//QzAHakFCl1PSpDAxgtEpJgT5VJm50CS0xJPO29Ira1L0IQUby
L9OLNQ2409c0Y9AiNh/3taJVpyFWxq70o18JDLDmo+AjU+X1+g5HTvTjSn8qYbvVFW0QEyV50Qwd
T29dT3YOXy8JZpVy1FwvTSKMHTSNdqGmjwVGHaEVQNDbCcqh4w4eIq/na2JCHI7vDmbihMwP5Rzv
zJkQEIPHGKqXo8SWW7ZBjidZt/V5BQRaq/0W19dh6btm4gAwLjRY6tW5xWxXjgtW4qazO1u3e4Yw
GuvQCLaPXuPPo8vShzAlMq/1qn0ATGf6l0IL7HTLtH0pZZKFjNLpt0TiXHaISzkKax4W8KoN+lpa
6GrrL0v97UjnSYiDH2Mb/mT9Qa0GgDJc2X9eEnNQHKsIqIage7ZBV1V8piT620kx9oZzRltP7Ux5
PGXWAYcAlhgjYIfmfI7iX1b2w8EfZ+7a3QXSL6Jve+QBiht6QQj+56T3oWhy3jM52vcnmHu6YabC
TNCJFu3dpbR+qZmhSr/LZLhDI6fvn5kz3YnusRcSCCJgmde3Ta6ISUQtVulvXQJu/pyuutZ4FTz0
UHlDbGccydWZyMT5aTktug3DmVcjtd9DeyZghBBcAoupYIh22Tl8XbsdsT+gaXsmCS1V818VQSqF
TDBactsn2ph+M8RYJGtgopkauve5iV0OoQZdqwOFDh/lIMjm6mmb7zzbVJ5OKc7DQ/C0jR9B2W+v
c+HC4Fy70bA+NL8Z9kJ9i4WK1dk5QUREiXRRV78H0aiBj8M6jc/YGSkVAWktQNmpO+QeI0sFY18Z
gaKRI64XWKQQ5RL/NNw9PtCG9gjKCW55FwdkOOCEroCdNdsE2Z4fpSE3/44+VuqK/Lca+6mTkUQ5
xNISqYqwWgJhxf4MSRNY8Z3SWan0xL518G6LMcvr2a57ojdCGCEN6v6Flh0r+gxiTMS7kB/FiJrT
rU1xvS4oiHc8SZtjlpPvM92J2z+FGsWqHsLeMxNV/rosII4aA880SxmvHNflztt8OjkAHntgR3bY
OWGlFW0BmSOknK9jpF4Z/h3YlYxwlmKC+IOaC8b7ywHEnQu/9vHoGtAjBJEh5a924LKKBKeGoauL
CC6Ey06ObikkrJquyeWSyYY1zO0hJh/RmOcE3/JB6r3/GVbr2zByT/5SccijnTkodaWLi/w/jokS
/D/T1HZ8ahlN4OIfh/GWkuV8DFOk7DJ7RBy0qT7BozBQDl6V3WyLSqMI8JM4p6ynnqB1weCgmALr
h2JLKPu8liFQ2L2Liym3sPt4mvZ/p8k8z4LEstu3DOGEIL8pRDCToIChIPAMjUxcsg4I2A5hSyVD
HoCjMWb9iNr5QDBLr2CJFNvzZ5Y3ftpd3ySuaeFDJO+uczQKgNJ8cwKcArvgQIxIgfosapXcAZxW
zWkFtJ4r3Xwwyy0M+kAy2eoMQ/q5dGWpE5EXP+LdAsSUw3p7jmhxwMvsdKTwIEukwNejaIJ9fHUN
3aJ/XIea+u7IgkS11YtTQAUv7+7tRmml2YosVIXWZEohYuyt657PYj0bcV5O1i97wV+GLwLc4ulU
5uleaoAvhFqI8145AH7XZG+i4YtJqRW+PR6/2V9EhXPKXeCXLVnJoaAq1IHte4BwUnc8NyHBnCMY
il9NpSDT8etRpACvmLDLn1bPq8I3d7njBc4PoAjSgoxjwSmCCg164dPxyMsd08obOjYSqXQ33s0p
frpGtfmNhnE1ocQIKNza4dqcIwMNhfI7diFABMtjfb/lkauwyC1sr85ozq49QFO5OKJzqzPA0tos
NpFh+KVBH5FT36zeT39UOUWDPnz+nCDZEcbHOu5H8DrNxwR1JsjzK3vAwwl0kSw5uNO3yhnVX5Xr
qkEkXHEhHLaZa0pVbkBbKpIqMV/k9VQOk078WfTuXLP8/Q5jag8Zojtqo6EVLzk4j1GfIJ9lVAz9
MBqi5/M206wHE478mJpLooovWbVZ25LSGekuudsgcyGKatX1nQ0hheJW5O9EwwD6dhoI6Kkx0wFn
C6/9OlrncxPPUCkCmeTb+Sn08q6JvM07vibqV/hlQ1DblhPTfajDdLU2wsDkhCfKcf4hmUIf2Acl
zZ/Ass+PT23knVkLBkovXaLiosB5OR18ikOCw8oODbmbQ3NQky+xqib7+rcWljQAZqd1L3fxh3h6
1kdqoebLX1gJMEhCl+LSH8AztKZEJ+RfqI6IeE38AYKDTw6Hs3Xm0so6bEurc5Yi+jnsOinvbglw
8X5u/EVP2T6P6QHAaSNWeWmMno1hggy/2240/VGebi/WM6sCE8g6iaWU4Xy7qcnd+qlwcr8Q8qc0
nNR6uXzQh4/+EWdnZxa4V1WyZUeVAiTCVUQ8qIUspRAv6xERx4JNY0iJjy73Pf3nNsOQVEkuNWYN
Tgh1XYcMWMVXkX66RPhXJz+0A3TL0As9Hw2HySfLhsodQesHp2GeqBYuNhkGYjGzGMuc3EM0ssNb
VkNUaPqp16ImSqcliv5eebmdjAHZYbq5nghQqQpChiGO8wRPwbDzGGc6S20I5xwqk0YhMmx43w8d
WvlyNxYTiw1e8plO5MaqlKWRVtKWne2EEVfSQG5EJz7PhLKoqeuCVBcKuXUCymLWuaZLmgzK2gqa
//Cpq/7dQ+f2ilmzoiJeb6VsSSoLmrGz8JIoNuRe6YFuh8U9qFZOM4Ly/qAtZ3o1R0SW867WG9TN
B2sxapYrs6ylVHPjqK/jySG3P1Vck/aI81L8S/uPKGXCpdEPIfISkzmUCSxMzyhbJ7NSWan9vJLw
djBaE7hnKsNIm8pssY+sr4SNTCIKMhOBSS1q1K4KU4mh+3hgq/4BsstvglEP2JCAGXGzUw74RL3F
Lg4xeiC3Q0KuBht68gQ4gF9vuMBDDVwrZqLQNgfpeJivhn4cCuK1txqzbr6glBIliOqvr/YfLz42
14sfk5Egjl2TS2MLpXlF7x8jmlTSYlDnSBwLaq/n8GjVNFz5CeEFXc2d0Sl0CWhIC6X95dtpkr7t
pNqbpqPSeqFyFHiewyR2YQn4WNHOJNNY5pfOoN8HyhQEmiqK3M+1ABlDhlj5dTPg4OD3BdnGgrvs
LLMjj5fT0OusXJfeC+uk2fR/4B6KaG/5T6JGQjUMQXlTP5TFRUyS9yDg/8UgMIWacElTVsL8n3td
fs4zI9TZGxUFIHS/hLkyME9vVaE2gNs2LGQ2OM55/NwE0ZOtKvS3R9ZGB8oNjcrPmqa2dLQwh+kz
suKZJj4i8R//c3kxHThugL3Nsk3HCR2Jvc4WTQM8DTzLJ9LV2/Su/9lYkbg2mBPVNHxC70bPgMDH
UkmhOyI/i7+IM6EBbvSsW0NtLuwuLEIyWIsmH/CREeS8RZDCaqSzoFa+QMRobNcSVEgmj5puiBbb
SADDweVLIwxFzJLCdE68hEu/8l43JsGDLDswGdZbdju2iPgd6SdcqrOJnItAvZhG7c8iSHm/hhIM
ejj35O+Sf0ZcezmEQuW1azkSUcE3XXCRrnPigQD85eRT1MF0xgrhREnMWgODST3QVBOj+u8ianHx
fQDh68K6OU3xZS4+qJjRhM7clhcwTm0WyPzF6xD4AJzXrqc6lIuwNaqDn6R6fm2kYA95PCBBMqJo
tnHA9eO4k6Xi0rTbkkE0cpMTh57FJehmEQNuNDSxuhB0VFAzkahPmoJoWXdHbdo3t1EuT3T9adOw
26yDsBddz0bJjzm4YDW6m9nA2k4m59DMJ9nLoY56fvp4TYnzzgP5QQYAMAdvs3/mI67kzS7Ayy11
y23yYKGvW4JIbr79PSviR826Qcv/Anhh1cIjXNxywpVggAkDtt8qQAOTf7OEmyZZY+YZ/MlTmk6t
Rz9VtC/5rRKZ3WjJEbsw00V7KZxMsfF2PUqfXj5ebD+oZjYK3tMAupagBstSHp8RWEqsG8V6UiT5
cG4E5lRdBKIGM/mQpfC3LA1IwyNB0xEi/XARefnAKyldr3kjwDv4P3HDz9cfGIl0OZKhV8xQsgAZ
RGRag5gR+0dF+buOKpyoNkSaKmUf9uvSiNPWqN9s3N6Mk8pyG1+gs+2rnCcZ4XVEX6YU5Aiv3ksO
PIKJmdEmryKlZMMZdrJpQD2udIB7tpRjXCgX0f7RsoL9KEnB9eNhlJKu5OIXURrczX9a79UZGTO9
JVnpmgp615u28AdmgM84vXlqrnPrL9zlB3gJ/SGxHiDmZwNM+rin4IJlanNRu1FKouH+wKjN/ZPq
NqLD4yuQXHMPPTkJMSn2ElqkC4L6+1P92V1tXpMoutaYNMcf5vDLxKfJ8+V1CJOuo0o2RgMMeDub
AyqUbcLZHqGMYdB5PAatm0T35FTzprQaR+Qjb3gR0eHMSMbRtv2TG40sY/ActEb4j0vPX5Z+nGG1
t1a8sg9G8X3iuHxc8O1huTbzILvqk3Gb2di6/CDG7/z7afAqAKOOCQs5z9gRifjY9E761sLApU+c
o4tHDAuZ61okT48oGE7S4JsNBZPa+DGvJSmgnB2GP66TmO1vnaLld2DlgFV58Op8z5DLluo9i7oQ
swIPbnU3Pq60BWmv19dVO3wCVh36dXIkB6vI+fC7SncT83RXSme7bSYdQc+Beg1v/ONcHzG1duW0
8AIVvZ9XyjkqzPCnbVPo/aYCpR8wTUfvTBfPi7qGjpxYYDJMe2EYUs9qqxq1ZhUDyZBdWI0LNkoT
JDHomkp+M96WZYOMN1E7soKucHyjz3tVojbRfTAeiQqjZRFRMoGp7zE1PASL+Np+bVqGKMoaPhNA
+9f4CpdweUwsaJijnkk8WUV52RG9QunuXGnC0TePadaiTBcfPjMFVjUBHeqI9yHBEP/EciSd6D4a
18aMWHztlHUi+NCSPtIHHN4avcTfS4UqA1L0s+JwwSNylIlljeFkQRSmdBddHeRHRfB63mWacekG
zsFTYj7TyJlD4k2fGV+bzhbQa53TKlsbM1SvrnLvYlU29QNda9GkPOU/wtueK3xDtEL6y9010X2F
29OcSg6v1NGe6xTmTpad5PkEoAUFG9g89yIDaxAXchD3KZ+rYDU0SyBdcjVjVXMIG86JCGx0HzN/
bn0gyKnKVSL7AzkjVTMpGydisQX3b4fOgqd3Xx/Afa9aTLHoV3SISQuV33pyf8jUTJoWQZ6hxWQ8
uBUDRFtzmlbWfTsT/kOQp1wB8LREKcysCIgcBO6bFw0qCe9GeGyks0Bb6g713d+eNs1/3sX926xg
lhy22jg5q1Y0ZoZT8noV08gj0KoC9ZH+p9KgYRhU8SQch1qz+wYwoO5M21r7K1QIyp0jzXsfqWo5
xBk3eRq5QaES48clhvaJMOVpub2pkzn79glzkW3pBP8pDJNk4p7/dw6Rrwil5wnRkrxjep6QLLVW
whWo/N5HRC4d5YX7fliRTTKQ8im78gadbuqnWzaI1LXCC7RAPF/tKecATJNkykDaeA/UwFM6Ccvp
csSjFx8ouJQhX2NLgc80qkVbeWHq3FsOKYhp/9p6Fmg6PAgfis81/oaOLBisdFyx0FSrxo7RwjNU
HyoPlS3Opsojb4XGHH2hRJfZwrFkeqSm093OCTACPhvu0XfJGEvCn/hTMW5m1zv+RljHXbNAwHOU
9Y4YzhYRnm6ZX8IDKQg1Xb4Tx6XZT+tFrKMiEDnvbobZQx8rMcCsT7EdPiZ0to/OuvuLB6fbsRku
uKqNavQdPnoPRCIC1jkn6zZklLQoh9sZ7c3XGgBcxIlxh4f9jLjQ4VRsi/E3tCZrfdsvXDTm22XZ
GQLYndrPafT3eDs2iEJxgTNpv00f64TRgnClZnTkfyaQBD0xiev+5zWbtoZzA4tmD6l2j0AQ91f3
cF/r7MzfZaUzfaAnZgbirOH3PuVBzKs46jHIvX7hTrhgYYvSyh+lp6EU5kK97PLClgsUaTrT3p0R
5225jpoCR6QxuhhcblSAPTWnUO14Z+yPR6T73r4pUOorS290fDUyxhFJPOcW8QliMCd1G09fO2Yn
htIfHL3DgCwo7jC3+tiEe1cnni/EpOvI+xOWSay5KaFglsGB1MoO4Kx6Q6MNjBCeK94NgLVuTTT/
u86LpLF3czF0oyaHBCSbHcvp40zRdka2sm4t1cUpDXCD8TcSUd2z1JooFNa8y/pcOqCEb+axvM+Y
rsi9keY2WdCBAdcE2SN2Cn5i6Qxqu6n7rH/6ONxV9jwPKKWXmOEW1xJPx+tJ2UMJH7x4rwm9BqjZ
cQ11jrkXD05jqeneyL7IrXPUSSv9ywSvBgr3QsegftJDz6b6B2Qd2cm6zMjIoesVQPWFxEuLYw70
rn9l/nhlpDrgz/wnbIgYRG75o91DjM87siYaGbaY2W+bZqHsxnEAnEpKLJgd6C9g2yQdbvB1Wy/q
GzsE367bHJDOhH+R8ZqpSpTGFJTWbw/SuzO32xwYDutKL1s0KWszhF1krngW+zNbPYVDkflaVk/E
H9yjgvzcTlOiacd0Y6AMu6/3wmQFlugOXz/DETjK4kXLjhaTlJXgDdblgziI2CyxSPmIdM0X9M7P
miMmHAVTFPR/Qr+V/C1H1R68vNH2Wejgiw9dGsG0w44RCgHwDQEttEBu5G8P1meWUJEL4LD6fQnk
A6J8wBGSoXhCLr8G8T+ODXPVJEAo4gZUyKMbtvTk83zjJnaR4pMIohZ/fwt9qQRV9f1JRm/VtIjk
Kl8ONOOH95LCWa4wSs+cpbZKf0m2z/xtH3dow6X1p2QHJG3waiQC/v31hor4tPz9HHIPbDq2yjp2
Ane/ZJGYGbT6mKfiC4LxuhwFizPLMxV3RRpkgY4FrtfaGySdovmM0CQQGwIv30pn6s9enleUyG/I
E5i3swcBdCq0aLnm8oWvbob5GOaHk7aNdGXV7ZGk21K6CI/G2F6wGwFTEFuyTIKrO5rOf1pQ4Wrx
HP+k/1xxdqLT1gd1WizoOdfJFoHb6Hq3fQ0ra/quomActjYkzh5S2w1ZbNmMBPpBJgtJ2h8Uy9Ud
/VYH/5U2O54MSpX5hSkhd3pZA40x128asTR32SvWo83nr463Do+RFSqoVV9+/tu46rLuRzgCrDdx
DkmTr/SZuZfqUHEq2tvgg3W5K2/1J4NlDFzA9YvbnA7kLQmag3OXNWhiMZ1LCHgtyt6I7hAy1T+J
xhcjfmlCkLXdCdtW+WayVSKV+Ux4gZEfSB5Oxp34x8tA/Cmq0quRaVovrXZo4aRpzm1OKazLh4ou
gNTvxCWfV0JTlF10pWsuNWPzFhwfgzd7Ff84lPK1VgOtWIBYGCNuHi76X4vsBhlaxnvXDqZzvN3w
lq+257CnYPvpWm1Di/XSMs+FIvHyx2c9gNEIx8Envm2n3phJ6A/w+V88UrssgnQkWldzYIBasJvD
awgDrwkTrUWy4JkVi1CWYrDSx8LoXSv1eDYiOxvLpTgwFxe0iayII1ftneYJhLciOaVix7YLWgT9
z0+gSuRSVVs0tjfxi+DPmKd1ZMq43EYcQhAHnwIodItrL5UZkpTolBtrA9jGDZM424I/8zzu0ZFf
ufxZdd6GACkewxzHiNFsu+PRqHclmQxsx4uUm1B0EkDqIqG86CtVOoVElm8A42Girn4IIeu71AKE
xIJYZZWbv1I4hyADCVFkzS/r5L7OZOzl2LXIoq4DnUKvgk5ZlK9ZGiBxSUt22fbuU6PVmIhvHKvF
oZYP7GkZaeWF5XfSJgJkGpvdT2A7r+MhA7xwmex/zBXrLI06OdBSVZSm8YGcPaQsXadf/wO+PYp3
Mhlm1/FluXcHvu6R1E4J0/z/WqyiIcPmYPNB0QWXNY4isSbCwSxjvVAYubEFJuSJXhHYqC7m/CC0
eG13Nv7TVhChwjj5yLfoaeEO3U/OjPvRnrMuyF2uM0WZvto4WVrnZLg9drDUN5a41RHV0/mQNCg1
9WijR7s72GFS/IkT/wPrxXLHu90zcRbTaercqjAX2krcq61VQamZF5+UHGi6AkKQlyBBD6Qm0Rmu
VDlOMz2Zo9FHpU0va/m2WoA0REK7e3o5fAFOR5CVGwrjeUJSAFOLs/IWOMJj5kzWK28QqSbnJSqk
7RboPQtqqHaMkXtiVRhP7DALTSn4z7jJKGQGQS8KfyTnAyYhQuYc3acT9qgpI4Fz0ZfRRK/eCf8f
N1+wrzc9gIlWOYwsN2lTeDfD6zERbrMxoNZxpo+o1FYJfIwNtWpD+CoP/xrV+z7EYfBZQIPvVHK7
f4pKr2azl13T/WFMuBsDNIBKowSBsaQ/4ZH6jBWcjQHHCIjCP+TyrBlpjNPb56JGoQ8sIPJMz0qN
emZ232im5qLU+O9fEJdrTGsWV53vz+uLtrILoscY5xtPiryzitLG3fcuULjcFGwYEy53mzlN/JX4
xHDO0yhU3lwoAbcubeGMHnUP8Q71LFfbW3sU4HSaF2Tkn/kv9DbkCyTC7ChJDx9lCahXDaohkWCI
dCmnygH62/Fnwwg1tIxeqhQa8KuHMKm2ycOJKZi09VSp1Ucf9gYxXj4jWjYkZfEocYh0MOb+5Ij6
bLKmy2Ls5lsSf7Zr45bDeeo4k5jVhUsBP7jE55+dNQ6SG8lfELwAb3LMBg7gP01PKugrlj/v2Gqj
qvijrovI0VgbdvsdDBHpNImRsf/7j0iYoOb84sGILvw4z56gum3NIgP2XM4H7e6FJheEr9rv8Cuk
udAE4pKAUyyZEYW9J5s19ovNNEgGqp9g4vgXKeNtmfy/2zYIJLpWMajLAerB8ZxVcGAH/YJa4w1n
zccnusS1dJx9aw/vqNxb7w5xemgsPRE76cbBVeHxwuPu0zh3CfC/5D+a8zfD7i2HYt7HgkVaJYOL
CxMolVFWkxh3tKRH3JPqlfsHOLN29Dk+RAwmuGYEpD/wjFOTjKkoYoQu9nPC6hDp2DxH/N4FZ5IK
NnLVnrezRKygaPbPobRT4WJ+XlNDDwAThnkAF7C7smBng5KGNOI6u1XkJaLbjrNvVoBT83JNCNAU
+kZHm110KB+gAIJNVFXPVaZluq+so8E9r5370PhAWraboVP37EUfnpa/ge8KD00AXG3DyUOWz6T0
7HgX719ONxIxd6cDWfDStHepHMn/G3UW2p6XM4onNkxnQCvS03QsRsQWXRYfUuWkXkT2aHT/+Y4J
S8WueNmWJV0SYOx+SrJmFarF3uwZ8tw/dgPRr12vgYvUBVH5Xjpf9/2OY8gjIJtHDu1ppJ0UxD1S
3zjtLP0lzBnBEXL5adSeJwVkYjT5FSVIrCAwu3kbkx3EDhwZTzAYytdbV68TMH90XUuLlpGgtjxs
NQoyNqYZERO0wq4HKfv75QB/lfNuQyZyBBFvFFqQjUTsYm6kOjj8PIFr8R7LXaJBS5235KV/+mJV
JfeUasbBCvPfq2I9IaCjCvWIP06pt/AYXl4jUOI0hut+u6IvDmZ4SyODRmprQ3Y185LZxz6dMqW/
mSQnmTre049+NNYnDrSsRWqHmzXPaHJ//NXQDjWJPvIacP5ERvjjvd7FJN90I7ubmreLKOHPmkYG
WXbpP11fp1amHXNnd9/vd2Mt0yuRSxavDuvPdFr6EfsHkkTrWRXicujDEk1E+73KjnYU/F9wIllq
lyl0NfGX4T7U+FXUYdwVtkLt76He2HP1EUCDreOQL2Pxo9rKTckPqCNdGkJLKGMNm5FE2S9t5QRk
OylT0g999+MBDSj2vil4VzcmAuw1N43BLJ9gLo4cTfeN14QgbFHQl9ahi9aPRCivwFisomcUHMV/
wVxdnsIdJ2maRF9Vws3WSbKd4Nb9a3KLF5cTGl+k5rKkjKneakh36WfVMrZtj6bLdUa/Q3t/G55H
2XWqrui1pj3ac3xpW3nUaTkNMN8Y+/l/Noa1APe/RcA3GZ2cWlrg8XpBDwsp5DCR7bzAi1ylOnm2
cVqE/9EQwGAQjBun3MWv1nDacYDMyaJ9QRwwVcte7g7EcsEzREBZJoNJuGKUNttgR5zbusnOVxhC
LZzliE8eZSYpCWidC8W14H9W8NINDaMSZBeZ98LmqEG7rZz0bPaBiZzqqC+uiIlclbQYTZc7RrVS
B9+pyC0VCZnwo/DSk3BnOfNo0fKqdotlkDmq37CImfZtVeihkZRwj5R3burPA0rPHFlvKwAaXe6L
mkfnFy2KRvRuxsaD1ldlaZXN9sxHQqv3IHhC6AKlwoVY27bEy40y+XyVgtqJlotL2NRN/myq/4aR
73Q1unIzezTkzhuSPxEbNUq0lVvK8CIWuI/F6iPvmikbnx3LZclt+j7UxENVXZAjykGPlLdJ910U
b0jAslnkkA2SceHs0MWjV+ksEF1PFNEwpmXmxoiWtG2lCw8CMjISAUmS8Z4f2m+XRYZfa+Nss5Rq
E7hinU+06JzpZWmXLeL9XDY+rE9os0d0ppc5GzEtjpZo4ulmzqPb9mmrXGyl9RYH01OixyfexGMB
RNkHmiijYi77KtoDdT5l9KQAjNUybZSk+Y0UnwcazBEeb3H559WNIgb7w6Mz50M2QYLeChgn+slH
HBDGrxEZ2S85uUhnsw+q6Nh72v/Nhkkari89irWGf33YiRkl978iaawQMirNkq4SgymgXyv2a7bP
C7gW/uiUD3Nn4gdkeBaUtdo9SaOZWoOieRctXz3Bn0um1x5PLKYc3El4vqrFxsxwyEnKKp7DPT4S
n3thsQCxaMTg9xrCvWhgvRHFPTyMlYsiOa98o2GFpFfhCJtAN4VMCU8XHNpIvpkuwHO11GJPRMKZ
XHs1vCLfoj+3BQoByCtBj++6xKZMA+OR1DrIDx+ZiELF/bdCwYsUM5t8axR6aub2TdDX7EvZ1H7D
eFar8egDlgP0k8H9/C07aA0by8IMgi0BIQ0QaaWWWQLtr7PswHpRkJrBsf68s1SiJp8ID8q6ar4u
KCWzSx863sZiml59FVsp1/F1CeWNi+XEcxWSPXWwguY2S6OIlzne8KM4+vG30ZHHSjEaZEKoSteq
JWg4JxxfBJ2vtGXekhwIKeMYTFZ+3ky/pOs3K3n+g8pu2P+br/rCyUh++H/ll10KnGY7dUdf5KW3
yuFTXs2vZR7jbVC9wYmteJ2WO5ezbO9NuWhRQUaQuoxWgObNvqzVSSlJJJlRVOzfLda8SQw01Tzx
tRfRozEwTIiAj1I2HfS6i+VIUk2DABcSTjTWEgspGyvJUOjZVk/g7sPAHDWZsIYA/BRk8ypFAzYr
BH+egRyF1oS0oi9NiRT3asXEc6G9FzttdJ4K3KrLJ1GwIfh6zySL1jzlkJ/FU1QZzt9iZyqsqizq
A9PYkcJp696BrrOEk4NBnAgdenK/m8NE6JDahDdyb/SFMdrpRaEVXpLUr8NKH4QrA/oYmw4X5Snk
ZGFWBJc8aWEpUqDIUhWom7rEAZqdC2N4KGLJz9xNQ07LK8WCUDjUISC/XGkuFbV0ZTh8u4pmw+Pf
t3pLrYd0IgeBmRH/sbk/j+ja76ZlAEYSjldTtqPzVYNYIuvwP4wnfMri9fdd8LFgOQT3EmBhlza1
UuDjwqwBzjJ28EdCPlnWBhj5Vo6Y7r+EchGR7JnzU9IziDsBreOqZdXTRljnVf3osDd34nkXc+p7
iNgjr9LzJxZh1GuQU1IdnS9Y9vMMwvF3Ijjv2xDZqIcdGkXAW75Lej531Wl7BH55WbX0VvTG+Fng
lEzYZUsHpbIkVJ1FsSN4RCAJ1J0GliGPWEGiBy2W0WdJD6+gAWz2DhGIJIEYVlT/lxAL9CicQ4eX
rhjm8/w7H1gPFmvQpBRQFN3h7GDe8xOjrcarh1SCyb292T1gYHlCy/4H2IPn/CeVJKxoPBBYBFRO
0PsO832bsp2FFqLZNR+vQsGjL3oXkNuNeMzKUs/aZIspoueJhiQELy5sYB7aVEg0+4WDBZifY3I4
mhKvd9EsyyhaIBOjtrUIkOqQrTifPZTUEhuUINOw5+OQrDmcyRACsAIrDW94RyMK7H4HiFc76nUt
vXSpJZE+K75xymvXUvVnpIkEAcUZMzG9SjI+UFKyVc4fq5QP2kHR9Pwk8i5DT8sTq8prCCakBTGB
y9HZCL11Ecf0wL/pFMgdArl/JlWt4ox6mAF83sDCYNVOgD+wsuyvtIzcduQTrZWo1D5aKLXjbabx
ivQbOlLxdQq9JzPXF4yOlgO96trc4lPQGPaNIKECBXtGPW0KyTEcgLv1/ZdLwJhbi2Je4zWvWRwa
K4mu2aOScv2E8iTnK0XBKL5jxYsX3sUN8pj30MFobQtgs/nZfIlO5K4hXmys+yUkU92+ojx+pCpI
MxX3jP9jPw22zxCgItTjOVf2IwiaVirH2LdH3aWLt3Iw+TRIj8tiC4iLczyEn/hlYjvpOfXlW4nu
jeEnCQfyNufFeditFWE587DAu/hJLPDxq6bwIo6NNj2AC5NR504EoP3AJi9phaUKDkF+tFDA2T9W
DbpM1dt3iirL7b07AIBL8pTJ8lVFn8VZiZGgooppwF0zR5Avz1z7yt8pLFeYiEbT7ZMxirdZa3EX
IPUE/jrom6Exr1SJq//981hfJrY2YNGbOYzcL3epfCqokYt5lWPpkFl1MDb1qkPktZcwblAIdf9m
aKFzTN85HeEAqiCtIikArTOpyWTMvhgQDCq6qZF04ebSGIa/KKTzCwDDZYzhrTrD69BX14utdNjY
9qOynTp8FnMtdo/iSeHgv9uZNxDwYeQNEVCgC85WCLHdb/QEVUJF+1iMfptNStCZpdgOQExjRNu+
RhAKNttG0SrQY+WbJu5MPd6qDo9E3yvf3cSqKy+I75NFR/6+WTU1VCRSW/S4x6lDiM/BZ4qZa9if
ud3DB98cQNXYviHrxXxl1h1w8UNIbTSReb7ffBviOIyMRCyFD+2ImVzWd1QqkCo4iqbp4lfuw4wd
yjdJxPjfMkk1V0CtsSbGaywKX8Rf324ucAjPgVWN1TFc6ZZGP4zp+IKLq3mMZCZs3OJoa3H1cM5L
J4n9tfqqOn4HVYsZDULzp82jVTt4Kzs82LeHmJ9JjEm5fMqmasXQy1msJIB8C0NAQ5IsrLQ4/Byx
MaF0IoosRb5kIol/cF8DvckozlIeiesw99JASOose//f4c0xkPJAvppT5YF72RcH7obhaZ9zJUtu
NEvMuFVU8CpRJHwJ0It0sHq6+6GoT5HL5ipf42GbkHtrzOxWkXVY/oVaNWShnA0uZYzLoP9uRNet
BIIpsnbnBalZ8jz175apJgQz2iYap1mHjgNm9vwErqL+IikPV5Q1K3YV8i+GaoAOh1WDFoL4PTBV
yHRinDA95WBM8OrhUTvKqsubXHI3Xbj7HzwQm8+lhU3LTuO6rjQXW5ggS/Np3g+85xgnoRUesUcZ
Upj0l7BEfJnKcXm1YLD+tNiqs48gUirklughYLwIQT4I77w1CebKx6KAZw18ubuA1h6JSBpjtsaq
kWTLl6bMhlpL3X+hyc6AlLHKzJjHRVOBlFJP4eD6AeoSiDQbHb4PjUHl8ThvDUzKpJNE+t6WPQp5
u5Mj3Yd3ridD1lmYUTDuwsf7kadx/YoQyYZVuIpqYRn+vz0+SDGXJuDAlHxIfZ9htzHk5ZInTn3R
tGXPfl7tNJyvuy4VT37PYkeCV5pSS4j7Y8Qo4ZFtmyxpW5VsH97kBiht2xtbbSPZ496GuvLDAvHu
kUEIPkHuQdbNqT8Ptc/0QPXdRTHhnKOPLB1s8KBrwxBlnEgiDKhIDEVpi707pkr9DZhdQ5EJCMYn
0+AUsn2mzSAJfi9XBtFtFzm1Pmac74sCEiKL3+A73kaXdYTq1JgNhDXQf8CByBYUIHKzAYXZYMNF
KnqTxD2PbtNfAmYmBT/AEW1LGUoX+WlGOSWFgZk0ZJWzHpzhoqvsFl+QZERaC85phuOyt0uQAnfC
rorPh9Qx0dbBoNyZMZU2Y6S27y16IvHzs1N2ZDhRltTgwCvogSTS2cNH9yHjNMmoWi3HcpsvJL2j
b2YmBfPfP51rbW3EZzUS1ppdn9/BbOGQCzxKERT6A7qhGLg9jSC316BNQY/aZqD7+rFB2mZkDoTG
44t4VzJLw04hjCZc+FoK7l6PXTBVQkN9LC/te0jn9vJpFQDefDC1TkMEVSt8/3q8RT1G4xwyMg1l
GnYoq3KQZedvDphFZM5Y6txATmt10MOsWT5dc8qToXmd5znB8pCWFpHahlQNsBH9E6eB55mAFa81
O+sNdLEqcKvSwsd1/s5xvlIQ7zvGd2SL+3e50cM9KFH7MVEg/VAP8GmlHPRWyRs4bSk4pWcUHfk5
zMzOvVLkLqYY2xIIiPAwC6V6ca85Ki4/FDE68SC6AKy3jOM9TfWDM2LT/BE4ykVHMQvGJeAm5ND6
RjsCWiFUx7Nb4iVt94Bck+SeHSNfrEXjWo4glRg85ph68zoOHtl0gOsJTe5gn8zau/T2k2deoJeK
TWqxTCEo0A18brRujkQkP9QX/akQ/d2uyY3a6kNMmn6PByuYLHLMaRTYCfQMOocRH1u4r5uIDPEo
eX9nuHEz5RrFJ+ujLpIRuN4+Ew4xORbSqbdP8km8UkZAR0irLHWVpXOqf4ad7F1/MY/vrIekMhjp
tBRGZ0bGWVaomB7tq0CuvRtwYsHhv+9P5mk7C2eGBSwajzd/Yk49dvPnm+dUjQQwrpa0Udq2Uot2
mS2JoUtD+4ySH6Fb0sjC8D4HiPvQtulBrp3JCw0T8rPcR0FmKmd/xRtlIigCcg82Ktd3fWuNKEXk
zqAw2T4/I/3wmNMg3xuCg2vuwWPlpJcdUY83NowUrgmM30wnwqsLisHRwEm/OyA/ZLXiLo7aUqE1
s+y19e/cZyaWru68BAOXlvbAlMvr0jhq/XRY+FoKVafBdIdU0t5Pw9mmUzNfm2NaCPpSmcgivbTY
XAtuAnwVtzD3LHOU9dYbgypoETZla1WaR41lZsRvyOSjZUETKXWCjFrnHeQBfmCRjfoxt7LQ17Jf
irh3uchj1MSKoP8Xw9ipdUVsqQMA46bFbn400PzEM1mxt4OGDX5tygPs9a3K4X1IA/1btf+UcUEV
nGLdybrQhinzgnPGZKaerwrR6I9pVNT0ZWM8Y/LkhKviSCflnhi3xKsCa2EP1xaYGj8/gl4FIg0I
Y2PzlAGsU/+UtIBtO1OBGp2qB0Mv5f4uH9GgktiRiC+UJ/fpxp6bpJcTwS2QTgbPUKbmzi5BzT5d
5bpY/25WSBpuRKV2+tidlGh13nCU4kZH0LghiMqFep11Xrli1P7DVsR6zN2ty2u7U8fAR1GN/f/G
6q8i75Wch9c49KpXqQcO7ePNwapt07EjWG1lzc8r051lNuFLzKus+0WrhVLfmzTAqABayKYVS1xi
oD8htq/b8cudiESg5P7+pMYj/UkY6uoDEqrAHVRpJNYgpMvIrnr5DcbsjCYqfNfWRPWt9iyNELUo
dDxqDbqqIo2KcJuQgttKLtRt/dvmP18L7xYzlImdeWLMuYqE7TkaIhG+MdD0sFKSwmh+CchJnVp2
bpLjqVCM3q/jQHs8jd4v04ZUdJbGWdyaWF6EWjWEdnJdl+BMS5rOZNFU0I83DUV46LqYmzxMzmSM
cnho56bXzk0W18oRmYQulUze6dW9OJkw6azIo78B3km903rGTYz1SzvLAmiLRbbBc4TzC8x7hv+D
ikH3NExQYsM6hcJ/rcNAz/cYfSOA+mtsDz8gRmxiJFEesdJKld6QJ7Kgj3CApzLqwyR2gLoYO1AG
Rrn9AN+iGAlmsNNod9TItoc5+fegoLbpnqS6twnuLcoZBpRC7QYSK3Gf1/BIbKnD4dFWRUHSfSsj
tGd2JwyCurUwEjQCjowZysKv5lJoqGrR39iUVLKjgPF3CLUlJXiXUcJ+tvMzpeFJCvsOnD4efB9S
HGrAfGJkngmF1AaU1MuYSGU/ka8nAN5ZyEAd1Dyv8aQ+E/DXP4tmfpz4xi+dZDLECT9t61GJDx0y
rQKJ0f5IJzJ44MB8tyhP+K+XNkIXsi9rAdytPp3Bd3BKynde8E7a8yq6kRjgCwIOYkIcFptQ/st3
6nOCTZT7v3UjLItYpQdaqAX9aO6OgSa2nkDscxtnsX0lV55MHkN2IJTxb4IZSBH1olinUBMrwnLz
MLP6UVzI6D0iAL3/L83zHjWTCYpfijN2MvGjw60fMcSoBvCA6xYMDKoPkzQ1aSnMncBgOu2mFeKF
PaYVpOzHxxhz6960ra7Qghlazve41xJkGioXiM533mXAP08vsRDRXwiBWTbXjtLZQicPKWMRa5if
36jOIVtH/sQWQLdyNCCapClM4oydAdXjTK72t97Wz9jwpfSIXFUljhPibhZ7YWaxLnuhO3ghrc6r
im0Z3Yt8eaZtOO5OSKmhc6MdL1h03xgGdB9T6+bmZQIotuYqQLZImnrRwS6GZ3X/0yAUCDMnD4GU
p/dfNCBrbg5FYwKX5xMqGNx4693E/NnGCAMnGPVjC1US6S8MIgTGzEyzH23/oNabdlzgGyGZUab4
5xpNas8Els7hRZt0NirBZeHh22HPDc2Gd3BUwhsyfIc4f+NSjRgryOZNYChBSzae2m12MYP0PCaO
Cgnx7rZrhMol/hWpKvlA9itCYOz1KJY8P/9DKMPUHgSbnLjDT0pKBpHN4MOnh0ue1fsc7Sf5KyVR
K/L17YyCjn+EOE224CZ5pZ2Dv6SVOukiy6a7lC8n+Yt2uCnPcvOhfJ36WdjFg2B3IBBIoCMRBi/Y
8FzHOY13WiqPl3TjOX69RyaI3dM4nOq1V53Pnd+2SjWE6n0DmgP+HaejdOSlpN8EqjxreM5DofHf
z1/I61KLn4BN52FMBFN4XOpKGNEcHO+gSVqi5Y9eM6VAaQOv168MmCUc8nZd97vTEH9zemVfqemi
J2zrIUqhbllUaGgvra+qrtJQGME0xKSfEUyJBW17mihFZxCqbG7GhIZmZMw4mMtmwKpeIZhv1wZa
ydkLngAvkdjUBiSy7oT/hMb0FFRl2VmVsrmC6/PUFxPVF9CJ10Sh+PePoTBAiNxC20UtUrmCGcA/
/z2i7ydTZXcBRZsiSU5dLO54A/Kp5R4XKnF9LqXazB//vNzMzx/aN9rVAHp+nMR2SlZk4Jn3jJg5
LX8/CdjirDxyqz3u7Fo/O7So0Nat4zXZIH6CYRGvw/w4eC6O/oN8Y36yP5Yst1LOqrbn8Sea68Uh
mdbySsJlSi/1ypwc0Szb53c0Dx7qTk+JgEdMeZ5uv7hGG+DB/9yIKMXlc9OPfHBITDy0EELk5pC6
BHEqDUKEEGXH4LSAvf4kp7gr0pg792OVkpXKEf9bKIihMEAAisRKIyF3GrfRvujF0WRUPB5Z+Wdb
++7/BmYbBnca6vAjkccIqHKTYaSOEtievl9Rf1BqPipQp0Up08XX/yVlqIijkQtVTr3T9Yd4is+p
LgtFs9gGuy7esEF2r0HmO0TkYzVmZLmBv74teeOlsMrQAGRKN/tYRUjDylQYiSOCoZIbFtXl446I
V0X6R4KPbP3y/T6xavG1wYS1U98fX318fodkHmApzrKZvKROFoqXGIxrCRPyx5PuH5OWuBOEuIme
J9zfAZcSC/NA0ckejVEVVMujY5KRjBnEOmygENzTShpTYgMjCEYYJahwjwknCw3L7sWWQqQCsz0a
hGmOCrzM0hP2bDjT+ALifaWmps0bZCY3ZD8CbmDwJun+tlnEcuGlZ4BhyLRThTS0G765BuShPZAO
8z/d4BO7gSgUheRq02AOyJVeTcOzp+hhqzCneouGCC55ySnvkHvL+8IaNgsQmG85tXRXU39N9TiP
ya5Z0XKXEN5ToCZspd/CpCyO99Sa8sIjNSmg2xNbftxHYEh9JqrBDrk+mtDP4VQf1YffmlqHJmmW
LgTpQbLS+UaSBqB272tEbFUgulfWu5mNwh7HeINkilEMzHq6w3rni95R1IZFtWKxcQuTUEC6Xw9g
StqVMM2QcjboSelvgJ6EzmB37HCZa/EgBp//0CaX88NBcM4A7e+suV2j7TV7Jp+AWJAx5bnwukgN
9NlgR63Nbdh+yrpv5eM65JgtLp+JTtEK1aOtYna9nDYe4QRZsd/D/jsMbWijpc3LfeBHxYkm78bz
nZIVrx8Wf1rZ12PD3iCad/HWDLX8a1dEnffZsE5rcrEw2uZbjEp1aMJXnndDUc9eUEEGoGWxlq6/
CebsmukfCr11GCyDOyFzEsdOkNlOExpbqmA9CgRU8DGIo0nnkWJXYj+jP6oTwMZmjPef79d33CC8
E9hQjoBUnPeKr22hJCJ7rXNm6XHoEfLvkNC0YuapM6g4IRb06soZQcXr0D2sxt6rjYcsKxSNI9G9
1Lia4B3GAzMQqVGtELVY8uXinJXVlSNbO0wwHhfdMZGw12WDheOEht1lFdtpNmSlosb1Z4202JD7
FOueiU4dNb/iei8vtetjFkdcLBMMSwGUMsRA1+xLQQJUyH2Wef1SdVavnkoYC49J6xGtDGqZdGhM
rL6ktGCYj1IBQ6ysL6Tsm6J/Nz1iSWsJtCWfp7feAw7TUFOxrM8egn51f4G94MCaK3efCgjax3be
8/j0fQX6bEO7K6p591pzprpkek/FC3hwTkyNQsr74QnRzwYXBQKGLvvLq0nmd0EMhIoLzcD4iKSS
vC5hAiknJPPOw/l2OMdZFxguEV1421mBzCpyYUCWu8yyTGJ1AF9G/3tRD664uxytUxbz554MkA3c
DEREIueEoS4Bd77Bpym1XUNPeQ3qcn9FSeg2UuRrHMEqazoCF3TeX62bjVWZxIHI0CWsLwjM/pc7
kqCQh/as7Y2vIjZlR7mDKPb2tmIBTuoSyQ+gC29dGsHU1MSJ3LvNWiI3zz2pgYKxAWYDa9G6bRKy
tshSQH/TkKLbu5YH5N0csdUJYfV9bvUlwouzzjU8zZ0EO6ka5aFsjnER48DRRFPi5X2eAx3P+rmy
/qdmz/HPI4b8gCtDghqkGz0DV8KDXE4WvFYZA1q+gGjwlZ9SFw+SMuSkwrtnpqfSq/VVjjeRprd6
21hwtfDAvgOoPxj74M8owBUjhl6EIjhC73ruHdUEaa+pHTcf+Jqge+m+boc+Ym8U8uINBQLYM+xS
9bJzx3HmGQj5qt3/TvIugn7XqJX9Q+En3NcYoldfMNduKkyuW9GP6l3ePLaVtLPgjRFGnKVM4OBH
272rNZwwiBPKNBIGYHcgNOAEaoaDEjAzBX+RytHz1Gr5Sc85grYTBEly2b5Mv6uccYeCYZcPXcKJ
yZYQ3alYO1bBAkgw+m52/B27Irto17XyHSSF9Dm/mcFIwRAAT6H40L7g+cPyAk0ylenDapU0zJIP
IFeNIodW36EscddoOtjO+zar1epiOlwq63vP2W34N7B8JnVYo23l+a6q6X2OvC2LjOQdy/2vRcUT
478Q2Bl/s5e3ZXX4Ng4lI7eRQaT4ox5mdRH3UPnrLIUb6E+l383mMJWeWh7hPBEIeDOBqhnDGrUq
YP4I39YqjUsU+XQrSUAuC+j0HEp4qjQ7P0k3qGVWFWlvXp2VrVKa6mu9E5ooReEtNEbiB337Dr7z
Ptm9J3wR2IJ+r1Ah7lYbzVoX44kcD0K4Hqvg7rAXXqAFsOu+Y7IrAYu3rQBo13M+Jk8ntk4wzbot
4/QvAUNg2eCxhRYigIw82NrBDz5QI1hjxPogLQWX1jfUqOhXCYM5QP1LPy55pJM8vMvfHYF47u7N
DgaVfjVjUQOjFvbziWBjxF2ll7gx7fqecv4hXOPCxIomNzk5Me/2w15cp/Ex65+lL8T6ORL1j6rK
dxo8aGjOdUHB+13ppZoBRXzEQzOtQoKip7UVw/+jXfTwpNblJVGC/zXvG6mrCVXmEZqSloggHZ+S
VyvpSRmS8s8/H8UBvJNBydZ/T/6qIKmzkkh47wqlzbMgKz6Bmpb7cA2pDpZySihzwB7e3zvuE9ZZ
v9K3O06y3+Ijy1UZO20nxNzAP8i8ffZQHtedLm0BAhKWjAixo8cIyGLr/CMSyPD7kLllQwPDxhN9
IbxJOs9Q9PCNYEY4Ke6l3emzbjBshHYNgY6m69LMH1aX26hV83GZaIRgWQYYMRIFerwZ0na+B1w5
Wz6Olas71SrP4TUQg+54AjEQ9TF/CMH8t+a/OkrTtZ1DTwGnuDKJMJw4Y4OoOa/lfH50pF5v2200
caxbZ7HY6Pw6hBlnzGywkjAjlm7E0ZfoEFQDu52Wl/wOKwkGi/DEqvuf73dYTxa2jyPupiFdSlfl
Bl3lsUshj/1MY8xkPSyx2w40I4EYukcc6JQCcRQ/NZdHp5PK8CsdIctPpDemM4nQIoxe+Wvp1sW/
be9Fl95w+YAadGY+KSWTbJb3ajRj3sDOc0e7bC+aqcfEcshnRKfcb2zYKSPUZayge8zPZcQQox+5
tWyu5EMtEQunUGszfaqZ6cXHCuo0XYr/483UX7/+9H0C1UnscPbgWHxnXVpN9IwII7XgTw+5uJA0
v6v338GkT/ccyMevvHXNmoJH1mNULznfMk1FtMSSAkDTTbKInhzdUHeUtI0j7WNtJ1e7LycQLSv0
X7dXuGd3wufsc2BsKMIbZeZTtUKxsA/iW6hRc6t7RAfNCbUj7fEbQCiUbmSQgYBsSJ/yV5gw5JMD
9Xa13DGmz9HUCVRWLN1m0/Vcu/r6sU2FekKdXLaz/Hz0TN0cgXMIiblNfETbKpiQBmt2bE1hJsuG
CQ4FHPR/I864j2Z7AoOJSYL/B3BUyyFf8DT9iokVwMD6Qxv9l2rbz7vOUDJAQD0hOOuXh0H6kWGV
t383OlIgRTXK389CEbp5XpeUadeTfyN+UEWoFugNNjMGIn8h9YOpzJnbKcWpWrmTsJplGfXm88HF
Q4/WMzY0AEwQpHj+C3G7BTav/Rpabx0r4Twb3Bsj92zfKuJxNeZN2km+JNDXQJwHBs8dF6CoNJv1
5mzhDNygtxKmfSZVpEz6hpRIApi4ZpoZNxBHA1S9tYTrMj/kM+wlkMPYnUTJ9jHJ5lzx+54Sd3h5
xu4k9ZnH1dDOm+VIna0nsgQ8SjDGcF8uLuWTqwABWf6ITTiUk8Yq2aAAT5Ay96lAe2Jq8+FprTIA
uAX+nTtVeqmxnXto2g4I1J/7owCc6RtLOf5WGsAhIZEhNS11FFYUopwQ2Af+jKrp2RjWgU7pG6LL
kESNucm3wQkf9FejrxIoxeVNtEy+iIpVL4l9aStavuFBiHIhOY4BsaUuePX+1noLw5CTKH8PRH71
q52ZcZNVh/FgRgO7xiaQea7vqUbbfeTzFyb0vb1j6+9KCbqQnD9xbS05deFhl1WxFiurO62niEpM
9bq7n614WBZXkMGWz3qC/ptT3YNgYF519L/XVJxsG9X1od0RT9MQHyCGqvu3UFxYbGcKgAjYnhv2
MHdpIPGM4M6fGi/TSXgzf+t2GXR+LIHgulChkD6nS+g2p9q0NJzAqcnGd1fsew8JRkuqUiHJSTfk
rnI5t2xVyz9iKdcYezpvowtbQqD5qjjT3FgSB0ZHOdL02S63T3vttQHoGaqB0LAuGCxxb1l8PN8o
emHqE16xRAHvsD4MVh2Uq7rxQWKHheSVab+PHhRld+X0rWJSTmT9ksqeG73vbMqnyGYh47PD5lbu
s1qs93Jz7PIrU9W7mIsan2lz1imxx94MBPx6FUAd3EC6IlNTMJ5rQEvc9x7U/LWCLuJUYy4YLXdH
h44ziHZUJp50IejeLIEw6YxJej/+IPjH9Q1RlA5/juQyelQ15XwXodNwkXiTFh+PqEEYT0LSMeNh
3Iv+p8wPHuYx/jZW+nWdRGVZBPbLyyXp5puTa3NSgzEDI+g1Ki+vgPXKBggIJc/RajImZyDwe+SK
o7LDOpNPkKwZ0KYhy0XgpBSdRP/mYoLx3fZjWGO6rf59bgQ0kfLSf9i5vI7WTe8dvtj1fAXG1Zqu
nYujcrGoNfBKBiqeIPDTJKTEpgr95YMzJkZ49brGrKsTl6y+1v/1xK9ipaaWD9OFX8//C6oq5j4m
wnkpVXyX6FkqkaB4P/cE/ss8OS6Gpju1+5GF3is8bGjLcYcZ5Smei+FmPLCcxVvFJ/WKtAhYlix8
zBogOgQo1olqBCJKvX7xQd9vNEoAhg7tm2LUf5lIpQvs/7R0Ul9DdrF4sjYWsT6Tofsl4nAxPGak
WAGc6bDp39b2N4Am4XgU0s/poBlzlmXYkHppIDeN4xocUJD5pYZMQxTA3HkuRVCDhMF5wn+1VoLq
NMKdhfD8w7DR62oq7AHT1gmpCWEH6CxYCEq0q5eCvTS3HOyKwV0QbzWAysLw0LObST8DkxDfD5T+
bGBEyijyBF4PJntrHs+NxCdkGO7baXZyhusPfMvN07RPVK+kFyc05leyZkY/aFgrLhafY5qD1gAf
KwjSx27Erf4Lv8pQg+dRyssxksMgPHojfMZgX3WavLXFH50cr5WIZvuiJVaT86GCQhkgrBceev4I
iKFH/Efuj3Ecb5AfzpQlTVjRLzMqGHYf3klXRgWq/zQAXQzohCkAJpMq7TFM5XhsxoRORuMbHnpn
ys+4QjnddxWiCffza598R6ontbBrMWOxa1yoA5ZB5CQIEsU16YtkaQcie8LcnFXZ52uUaOao3BiW
evnlMBYspJoC78A/L2KMltkH9yZPLTW0sUZRucE4ADNd4G9upo9p1c+n3UwA+I0apQZRSulFa3jr
2L32YgHCbroYV7SEuIzwwtDVZmZNKzwnFQ9gelva5RYhTUf6W2EnLCUVVM657MonW4MUJe30jG6f
AjEzg/B0rJqZhtwOiCMY7S21c0Ob8cikX1MZAxRvtYvvIWwPs1RGd7BmXFefTGf5zMdzrq3hA2Oi
bEUootJoBGEFCSpS2C2lni6jxaib/qOynmVODB4+3Sln1Gd/4kVstPkqNZMpBZ9RcSYpkuwcSLDl
zGXaZ+2QtYmmj/QXgGGcgiJ1y8h13YzcGQ5nLCx6mYO2EwHdqp9jNxQO39Xz40Pa4Tx50h8TRqCh
YNjgAS5sl8ZdpivTMCOoqNIo3FYjGN/Y2diZLPbhi82+fiEoZqqx7UyW5QoyhuqhmPkvlbGH/ASN
uOfb7xnymkY1by2W89nccRdRFmqAB7SgiGpyTW3WtM8K0C4lp2pgGYQDM8zww72CK5nURgP/PjcG
Zos73jDWdNOJyLsyOnwpcsl+Y6JyI+8r9iOwdz0n5iUw0Q8hA18U6/5qH6g8KB+4iHHL650h3RNS
42m87yuerUdv1jsL9RHS+pAbHB7aEjgY/FrMCfwOkwq1i1g+YpwKDSb6dJMteELqU52SpP6FsEoN
ZRLVbRuoumrNSKOTchit47AAyOakKJycAofM5En1RNTcUTcQ6BHtWROXD/EwFPa4Jr+RiZaNj3BS
Qn0czMrN96BMqJVYHUu2U4UhJzd3UY6UhQOfkSY9TMC/ne63E8xn3fVIzXpfzVq0nAHtlnnBVnQA
SePHQXVlCuvOLEj4Fvz2d5tveA6Bq1J5T08iBgnlSRdTV4PJuS3aPKROR0JLNG5Dkr9vT8nASh4P
bWAaqLCO06ierqxPnd5jYGJbYmUT/m9zjLmfpzz9AnrR7Z8GFmP466iLUNk4gWtNvifuGCWTdxJs
SrJ+G3T3uiFTkYqdVtWf7DTN8cP8a6wKgIJQ/7JTthxn15RcJngHuRd0b7pqSh5SPgKOKaZF2LS4
KLzMiBB5tOTL2apqpfYLd1cRFlKtrwOdaM4N+Jy8jmUTysBJ+LVZSGyINf+3h69quzIpzwrPjkCP
0RLh52YKOyN2bH4Wqsh0Vz5fmVPB8DDJXGIXNaiYcDmEXCVwdXbSaV60fRnpdYfTuFDcpDSuaVr2
Re0MC+gCLfe0D/PEHlKGkFb6g4pz8x8QhKwjHiWlodtQBnsgPek++0+4B7ToGI1Mu7hSmKo2WovJ
Y1UVnOU3wluJ44yGB+XM17PyG6fMm531jSFpLx0kRnOmYc2vX+RLLBIbjiLCNobpc3c+AKZH+tHC
Ta4TTmnYVYfAZ9oUANyTEGiyWZaHF5KPL5ZkxWpGnQFNOPllu4Hs29J2eTsrO/4Y3cbC6OCCoNvp
MbCpaQMprJmmaF7ZzD5I+FoYM76/GdA04bS2h/wcsmMDEn16r/J/f2vVkixuFDkJQsL6sIY12v2d
QOfH4hVDMUzdOmxqlmW/I9Z54YpFo3rQRHQKzqmw9bVhzmro6KkwhHvsAp7zN9u1WC2QXfLGwVw8
ksDj0NntnRyt/z1Gf0IvftKFgKDwGz9/p/sOBMq69YIm2EF0e7m5Ws1Oc6+gPDVrsvl5OeYUNwmp
K4eMcQu4QdzU1zHqpAi5HF6cHBnGni6ZgEr8nD+3W2HZtlnbseSXD03wms1Z35SR9UiHMjGxvRev
URY40CQepLG9iPjLxFI3ba95PEz2SAOsXYNBvqPHS8D/Dp+NoVbfrWRpHiyT66Sbqquu+2wJRfeL
x2dfUk8ly753DAIFy0Cv8sUx07Cq4qBUxSlj3P+vnL7L895YBYjD0FHQenioxDMdKlA7uvqW8oCb
ULZ94dDbSzltWjm1NbcHtbkstLM/wuPWgwiQ1s9yXDZkGfGZ33SbL8rDLPAtfDfCyRzVPjd+gTiU
4NBIySvWmlOqbmYjRIZmj9VEzALnUyQ0KITz3TXs/6wGQcGJGwRY6AbSKyi60rolFcL2jbYclCL8
fvjoyhgTjS5rYowkVXo+A/t1b2LaFAJ9rpluSw/c8vEqu5vs9WBq6ATbPy37cGwGfaDiAQpHKUwd
A1K9ELMYE9xf89WVi/qOfhIiVQZ1+9EWj8lZ0qmxKhVuleRMkCQD1xFa91mCygbm3xyIK+7CkUM1
31AaTiCWnBWvGTOZgAqlWhQ1KqcmA+kWpXewzY7o37fqcNvyIF/PP8nGYywdmfeanQ1Wjx+r1QOP
8CxWxGPoS0ULVQdo2D7+iNmxZVLAPzXmxtaUpEyaJHSEFpXaVzsTQsvapFG8JTLl/XeB2nPXItFe
2lv4SJz60BQuPcDQITK9e7//pGn5G5vrnYvfVCsTjnVUzyGnIIDCatidmZPppXXffxflQlOOpEKT
IV5wdzXCBI0FFWj835KBNRwQeF4FinsebvknFHi5WVIgWl9flOyLWqwVnv5ut8QpWyQBo8bwM623
pbmJSw0Aam/Dbh+jVxRJbLcoebLPRM3LYJ8Je0HWSlSKwMDKlNNZjc2qzhmlqx8zOtAp1G5fm8xo
kr7xjJf9DY0AJMnbCTpElQyoRMiqvXGgN0HmKLN+8Awn7FeUeHKgIWxHwv9HKy3sr0bhURobbVfV
Va6girIz8vz6TrNwx6s6hJkIJaKnw+GB7F7hJ1McFmAkHWPMXxwYzDwW6ejcIMoTunYGDklOwv9J
1n/xeMjWNcEFGLwvKjUp94rdAuleIquIfK3aiK3uvFtEL8g1zOdVLUgEl2YDeaqmJj/sS1+YnWHe
owEvnhDKSNMY62QkwYVKnqIcoZjrjLpeJgW9tsngtUXEvjkmCqVJrTXtsPIw9fZGdPvWwgkY8Db+
9+Np39T9oQGbxx3CNtibe5Il4MuEnAtDrNJcDe44D6wdHoPfDBeSD/NzOt1dm9ez7ynGX5PeU7RV
RPR4fMundQUQccoIdZDq3evyDFTGR026Jjo+uUVRm+MhxHPbpk7jmvItjGsbyrzacJE26XcwSk5I
wA6ZdVgCX1G0gJvnvcVJQpGPsr6qozQ40cV85oy4Rm8ukaqVaZbDlI+GEV2pQdpYNrsi473NxBh1
fnNqJv2ECwSZ2it4MAFlEQCYdVUzidLUC9+VRgUr/MWkkTYklzoG+yL5n88Wiz8tcnGIWi6GCfPC
whEc8ClSgQNCxTwLka7OI633kd9P3wYby3jsO6GCvVoj5pj1gJvKj15sbQ8U3shOO7wSzrc0TBrT
xA7WutmtOwe0aI/C1mZU8AzyI1s4VLPhMbMRJZg2eHExQ0a536TrN5rVh9bQ7sFdeAag3jC4InX8
elAjWatWJb0atki7tPpcY7fWUB76lN8z8Lhh781LlvKBWejtGLaezK2BI/3lDnEGsT5D5VLL03Wl
QxN5MVK0UuCJD1yqLng2RPk9PRum2WxmaCj54bE/YxVDQmqOsgLQmS77wp/IgvKEceEUW4t/BH9y
KhgDp0Dx2lqDhycgtdgnuqmsgcBtads9puXtNNPCWCRDNdSHcBEfx9dSqeM7DUV2nhltUJ/60yng
fHf3QWpABeYs8AjcE6H5uIvomMgFAc5tx5PYbQsW5UC2Ydr9Tg+yN55PsxbGVQJPSXCEH2Flrgtc
ypVfOAtmkCAEBU7PirDt3HG1sJiksZG8DyoIamhcAdfmT7GPNIs9Olf6/6VsXgKZG4+cABf7KMOC
3C2/qpbeRjpX6k+dT9S5MyIEcK7pAXpwWp3RKZ8pXeMGOLb3lwArshMllCyMHHU/bk/w3IbCBBCc
cL+fS7zKO8dgl/Hpw6Q/lytCpv3ZQEYIRwzSTTQm5Ss8EK6wjMG++ocXMrE36lFESTxEbMJ64d7b
UYnCAgYaqgVgfqLe80k/32M+sJj3jJhjzTP11Y6UmYpENBRwQzU7//urWdiFRg/D59ygEkPcKpaq
KgqSPeIindQkF8udN6LM086rSrRnybZUUADJ2WonbBX9B6xw9kG7sN5PUhB1wz8OFoOXCGPSJL7n
zXReMnk8+EGx3fpycYLtZRygNyujkupza1BCRkozyjwCTzIAbYNxRsfHEKlahrLbPrgpQOQK3PK3
ODStCDk+7729f99+OD3UDYmBRPUXnxDGa0woxCEJcKpy77PsG+24WWV3z8r/u0FusquAgDKB8X4v
mF/m3zkGmVQqtYO6W91WhUXHIHPLwATtEEoJlYyAw/WJEAOcj/yjIFBK0iUeUTjMEOd8uEzGWU9t
kn2744RTz2YET7mROce/xymiQlormggqUhQ+vqFRjtfJdbiyZcXBQanF3OBxVSMpM4EUn9Z3vnnp
yslPC2kzp3V3sNcwvIwCjHR96ZtZ+ZeHJCGL+uOd6lFReiRmjam/TJiP2SgmAEwEF0e2f7pJ0Wtu
KtwtgjFctQirVYfRb+xQeXRCPqr58OZPdMd0Zt1c/5w2DC0uKtJlmcZcN4BTxB6E4p1JZD/tQIR1
kXHKBoQlBuOtdX/cX5/jXlFm/FMwxHNHB+CaKq6c3IlgG5SUAB4or8xG/2CGyAfrjr68GoBWP9NN
ERVBRE0aFENrfEp4twen5BAKO7GvGuXBin8Q3fada1+3EYCAzvvCF7VpzfPqnoCPl2Ca+1IDp5xJ
zc4M+K/wFQwldljA4q3RRgM9Wo2t85hhf/8Suf20f76siK0zmh8+4hWgCaJyTcgU2VPFMpExEgjl
XodK8ZvD20EYMW3Gfv8tkY/urzofuyXdzExnIBIv3n57AR1UylkMqnRyIHoa8O4/FaSxZ9/Mrl9A
BmC3RhfIOYFXVdJ/KfV9QKYrEqSPBgb2vmJSzv84I8JUluSr7WPU+5T1ChkQMGiQxN8z2xh+pcJ4
qVUNZ4iq4y7U7vVInuYougtkeJGscx29sKq1rM+45buvYRIDti8/BjxoXtwIdS9shcx4hvwnv5KL
wz9HC8FXgnxrqm1zU84ZrjJJn02DEWTrox7r2cdDh2w3SG4oAJuIf33fq14Rj7NdfOlUVqF5hhy4
H4PbT5oeT6IpdIbn0uLjsVxCRX4vcH399NwVBvgE/Rz9ILAqNWKDSPSfIKLstU63myJz4Z71DK5t
Vr19pDvFejGSOKWaFkKQN+WOiYF0C8Aet04QiL6B6jksGj2O0x+WOPMVUEAO0tAwqbwUNkXW05lR
QDro0cU1h8rm94YoEQS7pnWFwR2IoM0Uba1NpBAnRw8iPxvYbjOe4MM3Y6vyodk+1LZdN55reLzJ
+WYEEnh3e7l1ahl1rjF9HriF8C2MPwVJMseVwmYhssn4f+HctfhHynCpX/27J5xE04chM7dylfqW
QnJv/PeamAQjwi20zRrEHrpjqR7csJ9vdsdUYe8INgYjAprs7DgBH4PvCwyPfVegCitxyukmnaw+
/ykciyI2gmptuevw5n6wfrJBtINboCWT5e2VHikbipXhaVuSAmvSqs1JuOvR7WXiBNsbb0VCJoRi
hmDc5jj40eoe6cKbE7pZU1Azo2mTLI5mFAOePWoWpI5sJPEwh35kSplURr7l34OMRvMfvZMraMBY
PgyC2wYT+ZfLPly7nX8H7YIvtayGJWo3imZd0fXn3WiHE2Ykmf2Clj5+zfRi0qdT7yPnvVsyL+Um
j5QcRLzitWlGH7wD3JqdAFwtbNVdc1emomj6qesVfLM97y9jFVl2DuHNQnpUtPxAzsG/kQ+zLGkm
dQjAoOx7zEtxJcTRNG6U2l3VO7SJfEsJdRfMcPQ4Y1KqUSh9rwGXh2D/gt26o4HKZQq9QY9WXShd
U7s/7IRA57M9J83gOs9hEoaQhkBEmeqnWavMlbbhhq81R+gfVbc8TtdKes4Jjh0oU/T91CMz/qB/
HziK/lx8UDHruhcKRPP3AMJ0XYp5W03k+Wq25t6jgcikU7Qe877Cr+72YLpOphtW2fyMgN+DPQDo
F81hAj08cdOcowxkzPMt4MXd00GEEOdqUgCZCBHmggspe7O/mOvJDvpSZmqXGLdch098xOQvQcnD
UcXuVGws9sHU+D5dhQujSH8LPU5pA2m/6ood4QeHkAeylFPs/RYI8km4zQJmn9KnLCfbKAoq0WGl
dSnOqFLkcPR//kjbsjdO/3A4qMSTxJbxM4uaW7SvZhFHYkeuLmLg+zyjztI2tU0ZKz7SwuMd61aW
Hp5t4n4LxA4LuWwQvznze0To9bV9+Q4XAZzUoQV3seD00WI1kBijvdUaekByfamzTllpHCUUi/id
ZSUEQHvyHjumMT/Ysf2X1tYbE9GtE+9t1p9npgXxWimWvzYCumoto3qWAMsk8K4QQimE9KfrANhO
B3WZlVG/JGWExD9rUApKOCWjrzNFnea48qsdNUejeJV6+MfeOfxLb6pXsBsnJxymmx45kjOn5VfF
8HyRCrF21DOKooX6EikY5Ndb8sjjPFd8mBtVgqHsT0FJXg4WNcKutEFplzysEOjfwSMs6+9yI+/k
mWygkIO9lV/ngGToeFgmcSJ0a/ssnqZiOFRNym1paFTs0i6vJ29QVm1ndBaLMg2n1YWu9fLOQ9tv
FXo1vU3h1sHn4G6Ht4ubFGy2hYYb6GCoZr7cCC2EKI7kS41e38VoI8gpBeRy5ClYqzjQ2vxEM+Ue
h1D5BRHYppDcMFgjsYuJ6x2rtBw2+4nSvJvZr1wG4ged5901v8G7iY8FpCNurAmx9UnrlPlwxP2m
YsjGd7ldymB9YuL3B9uKyzRlA8iKk0XBVAbYGrMsRUEew7IU0tNgVYdQUYjyNurRpVuL29ifOog9
fr2QPFupbn70hGI+KP+PyKnQTq0zvy7bTtXH0P50BoQkDuIkBY5wKRLaUhOtWBfzbETljFiTssfQ
dv9+jSzdwOjk3ebF9pvVTY9W47Fk5+nWRg5ONWPQjDYXot2OtgnycEUjks5ZGLfrOXSYgMLwKXFf
0OqMAQPwl5nRm2hNwyC6mYOvz8gGZpZSJkThbFVX4e4k9lHQDIkhQI5+kAPZduFmiQwAL+XIfPFc
7CJ29D51ViWg9Tq7e9p0aTYc0n/QVP60b8EFQg5jjC3JcgcY6xSMySdsMektncBAs9z1NneGXefe
WnEmRO9ZJnjf5917sFOjbCy3lcEJ8LT6jB0twtp/z6pVM+Uzg6BebfMvUja4q2f+inK03kCZM2QU
QUW1jQxR/1CVMgCDR7aHW+ioAmbFJDh8TiCvOvplmjf9idE4MFhO6XpneVmDUHBZ+W5lP0Ct0Xwo
4PKZTm9SsOfLobeupe/dj9whyeVNplAzP1PCJQx0cu+8rat0YjPhmuY+QPrkIDgwPeBeNN15WO+M
Y3JBqf4rMaKwUuz3rahP3BjJtEeZIo9dzuLQ5EIzEpp9baTZxBsIYVz/dZSTP5XzohWWIzsa1l3u
3d1h+ptqckk42rFNzaNXEiAjOCmCe9FR105rZF0KtiC9V3KOLwmb42xuiRVtRfkm2wsXGLixp4QB
2/HsqG11UnzBQQTCP8uLCV1XRRI7EFqIf05n8Lhk/A3OBrx5cuUeqNn8xsqeGWn4xGHhPoJo/moJ
MSiPtSdMuIFHDn2PgLOmRPVLlH467xIkbU4SPfhd4Now87CXqBnOC58k1TYpFonBIM2FIUldSVLp
s2pm/5ZLkSAiNaV3husgfqJuINi0SBzbumV6quO4T8Li3RWWh2g5d5iwZ72IHdnNnmp4tt1scMWP
6uCu3IHEPL3t5qdZXZuoery+FGk0FvXaiwxLsBPcA8cYKCJrS6XgjWsWEYCd2HYgIaabz7weKse9
eSi8P6V1vMgw7iVPZMZlmdGsSoJlv3VjSYsIbW38CuR7FDw3YP0qScu8GmKlIp0Rbc3RM7HlUrQ+
NT2ZVeryZSAMbbdxjBROrENixZZqcCK8DOLA6vNVmpq/05/IaACIPhDBPFmV0odIzZ5n07bEQe83
gSHJ00yXMe5JBXYS8hty/O+vTTdiZ6m9+/3t233GxfmeeZje0LZPSYXS1fro1pw0AF3Fc19XcaVt
yl6qR4UUN48mPTJWewWV24Kbv2g+RlunWck1JlA7aKjSQCaK+mwnNXe4X2Dhxq+RqLBX2q0Ej3Z4
bhwWfYBIyGFtSvez0B87KTXdDPsM6SC+/HYZ5K28TJlb3Afzb47TNamrwovjV9za/Bywx8yqqxpM
J7/6v8IEO1Yz48kVd1umrc+ANkuve8JINVNKYPhnAg//mkOSy0GdeoRpdH8hQGjHeh11ekcgAgux
4YY3yqlWgGAlxyHs4oOTI9VoGdGUQ3faJ0t8ADFEqtBxBmqmMpNaaHPjI9FR37xQje0GcwLe833l
vGISv5UxowPYzBOfvcublndhruaW68Nf8OkipifpnOAmvlANPut5e1f4v9trPu0S1nHs+9JAabz9
I9tMd+8074hgRcTFmq5r9KVBxkfnqsWCQfqc+zOz3UUVs8WmBDOv3/WF2PfpKurklgWIjv/GfnoL
YTgMHRjkXA7wBUlydcwjcU/XvSkn/27pZynJIrFlk23PzfDCKsJC5NQ2kt0FYDCRppM0//zFjt5m
g5L7dmE2MYObjfAXLxXi/y0BBB6pbXqzNMtfbMJPb9bcQvxANCQhqwX4ZUo5WdSWDfV1GBi9WF5o
UtlcY2NTpC/Qb0Jt3GXYM3hR7B0ubFeEyvWXvgYRWi/LEBYSMruHyKZmRfeZskgYmGXOeU3Y4Cz/
qVyrB2Lo5M+jVdggdNQMLOSJWyloc+l32m4jVK/eoD2v2CgMm7YL6rXsJRDWcWx3+AIvErm74gqj
E4nzlbr0tggKjVVEyrzpipcgkljeExhQjn5VxWyg1MNWwOY7GWhYfWVk+T7FtGfdioNCPVPbF6AM
YEznOzHLleXWrrsUqgHhQGzuNlYWSIFweCIHFDDCVMJKSb4hm97sJxnHy+td1ll1lXvbfZkGaF+D
IjeEkqxfajaruZHoplX1UEKvb7nwNPTXi4MFLrlzqOIJuexuOaSBzAjxOiJ6O+mk1IziVApiyVcu
VLVvFyGOe8uaJRxeZHbAXO4hQCtw9oq14iszVx+4o7/vVIOXl7KpuRQkkDNVTXpKIgKJIJ7qUf3H
rnjhxYh5XPa7cpJjs36vwplEE91DcNbc8HpATzV9ujCPMTu1minFNB6ubIatnrpwToPTK/k4dtr+
bYDw5gLYwO+GXuQS9Ay3prJgVHajNgdi9OsLiR//JVpCRr/PD6yRPdKIjD4xf3w1DSVqz7qW77Jb
W/nhbDnYFrb5DRfZE0O4s1jy9wy/IbjVbcYgnc7LcQ8tFd48mofm548UV8xKzUjEdlqzCqXhIeCQ
iszAVvbp9vsSaAUcE0LjClnYC04/XG3cIYw+SDbQHyZmNoHOc7goOJ+H8wGi1thGVRFDTN5srdXe
8LPl1ZXucKaNHfRDqLY+QYatQBg9DoPWRQRAkc2PFqERdK0ecFlVKr5yMo5M43Hx/BI3/al1Fzu7
zZ1Jotckar8reEm+f6N1kPucuDwPzE01jvgGj5y/7WxBtsNl8gXMYO/k4wa4tUlWHaZMZrjujhpy
aRynEJtqSv1jBae1FL1VW/VvugBtmyk/Ee1x8UDQ3oMCQ+a/5KTNfhiHkLmiftBP+UOz4nxF9g8q
i8tXl1789yQntIzuploJW4qozU9Yh0qhj4qeMtEYy09/XynpFgrMp77msKInCQpDH7vlNJZvscKJ
TGjke/Njc4/fddTOYbUiN6qlLXh9P+FqKBLieGQXrXYp60j7w+DcQ2tFysr5rXWv2HAVbRKBlnMS
m4uhvg+cINNq9XH/wna5a3+Abw8AZTI5FOoNn7lJmlocJQSKIG8NmdjAhWM+E9Ex8n+Tgbs6FYeQ
wpaM22zYAmu948QrvQibNvpedqpBTMSVL81dPln6ZWlv7PfFyW6cGhbF6Ky1HK84siN5saRhwqbd
lu8jvsaf6rHguCP+nyNGYVf0OdrUaqjPetRLK8q+HBsi6PeD0M1PpoIiArXCTBFu+trDWRzcw09s
xNoSDA5xYZ1DXTMV6tS1/lhfp8gw2262RQQAvHveC0mskn+e2UcAAKGm2Lp7gy9Wrb6qaf3IX2vB
Dqe+8gncEKpRS7reaMp+XZdxnYb7YHkgZBs9ywHRf8CpRLnJphN0Uh4V+eBvm6VnthoNfMqEyNBs
2Tn/cSD2ukQ3AnavGHs+7OXWHwi15Z3E3b4XlTEuSQL2WFaVV7g81hd/+JuCtxPIzvL4AzDzQgSN
V1RvTWuSRN4aaCofWshadsLOUlaHY98PPVU5AgS6DrpawpcDUB2S2J2jTMbJ460dkPhUH4i1Gl86
LdG1EWp7n9QmUey4DPnyULkOQcFgsKA9g2GqxowCHUFRoOudy5gvWciODa+WdS7JSDKfrJBmI3Ql
5GHhWp+axQen+sU8xeKyW6PlFCWHww+aVuj7GTWyk98fmedqCxNbp2wabbcwEyeqhdqvF00JwcaT
ol1Jxe5GaTSHL9Kned2gdYEOJ3T986EZclbg+i4dGI+aVT6f16swmPdUNtNCYpcxHpZrRwDVdwvF
HXOEHH29tQ53m178B1VFAdK12tjzM/trIttAO883QMedrBKeLU7KyePcvLRvTBu8w8x34q+BK+RG
W6XZweC5QBcyWuBwIJArW2lwV/Wj/0dX98LVf9YC6zrV4NMrz9YjrVpomcxChejFNExHc0VqO0jl
N11Wi0noX9g657mAcVov1yN1IRDdA+S1lX9h8+yL831zrIlRFgCOKWCoZYGd9MK7TDchFOutrEDY
t0j++ZHsxgxb/Pgc9sQGH2/0gO+VgsIL/zBQfkP65Scr6HYzeluy6uGZd+G23PS9dRi8tgGCp+cz
w4w6JgTlH4B09p2xEiUB4SwOEJZjoKrP+vcdbDUHejX9C4WCyxiUuNa/o816ee3A/mFSUX+MaqlH
hvB0Bj3uSKl9Aelwr4/N18JJLsNg91BPG2umDhrm4RiPPCt1uHNb8wKkVCdTH+72QFxWNGuMKwmA
XkLG1wecaI3IZlDCnAjXv5juzXOwhN0kKZ7dVAo02oIJfs7NGENQ0luIvkWzuil4GRtSs5Wdgjek
+lw7weLiwXVZbhMDsHr7XLIrKhrKf4i8It39FsvUkJ6yQegLmTsisLzYKuvoV97lDkvJz71fyxCE
IUCRk8cBhLy+dkAOC0HOpcMu72KsWkhuCt83b6Gt0l/WIbLwtECafDZgknemfo/byZa+u8FExJQD
rbLAmeTo1psIHGguRG5vHcBIu4k5BXqPYNFEuKkcz+jsSXZLJST2rN9ZD40BwROFRLnb5/foD2bJ
eiG9JZGU6QW0kRKjRY7HoyjCwbwSoIWqXGhLPQVVVIyY8UVn3e97QeqyTYW0O1BOMMsBvaf+9mMK
pbKYxOhF2wD/M/AsYEKVKvfzavuTbJpdtf/9fZX17Wl2HLEOAVxLbj333srC7MPe8+aWqRThnfzZ
Vm0sZJl1IOzfUHCS6IXqorzp/t6ESltpvpp9b4KCE6V8EYr7HRxrGhcEpNKuBMOgdTa0+vlHHtlC
MEJCONIPZYvfsXgB8e+kC9VGawCH8X1yz2zBJ3ObE+5tV+RcQPDODf0kdiHMPZxgCCiMi3Gr7IqS
78t0Oi1pP8gSKXrUMBlBBW5Qgl3FVwIHNqkF+1q0Uu9/Qmoe0onsZFYJS3dl1kJ41vwO4IRHyUj+
v4F02+03+KCdvC0/Cm3w4r/u4OUkxmgIM8bETdF2Ui/4TnhinfNXLcW8ksVw7ePH8IzI8Wu3buz1
b87Lpxfl3pGX3sZRI59M/ONxBZsY1qCkVuZ808Mkd+cDNxUWorzTMY7VG+pcdPWd7SrzamEQOLjG
bRoUGBb+WOpVOUTv9Dv9PeFR5NoUHse+vgbpEs4a9EkaCk+2FnrFDDYZ5vJiumNg1qcvyJlQuIMp
7rDXC4OkJILaJaq62J9yn54EEtGCpcu+WNl/AgPsjKlylxLnwS8vswPlihImtaahRl5OOiwQdv+u
T3JCz1gvmzV8JluFhtoTCsjGNniGgLpGF5jQmOG9u7VYjwD8e+RpLG2G799NA8+ZzO2GW8+rmgDr
Sg/1i9Kz/J6zcNWdIDBiFc/vIf4j7KsQOav7D99Ms8+KYs+lGoxSG/KiPTndiGWh1LaujZuuJlZs
iItAPEHA6sVn5d7sTYcNGhmKliqOomWJuAvCZ58vW0NxDCHWlUQfdf5uhMCInaRIEvugDXLL0ZME
57j4OvLinstU9CyPy/S/B/r3MvG9eE0oMlYWdpF25PiUBQ/wGjAMZAmhskx762V9PmP2MWrUt6m+
z6L8LU/viroqVZ8kkbUzPE7v/q39NEqn3/rU42b80tKFoSWjiuNJqfgMOvG948hlEIvEkuP1PzxL
FnhvfZXY8o4z5yTxtG8spPnKwoIUOxfVKR5oRfWrNz0rJkk0VpPa2v2ocqkADAWRTfWiRVDiAdfo
Ucxj/+PkJCLEQlCooKywDILo2705fXV1M8F0s9GXHBJr+ZaPJOu3yGsxgydh3EYQpN443F4qHaBp
EznpcG2MM/JB3Qo+8cAAzhMiBb0iBjQCN2FLnvWC4HFQKcEZSeQI5mwDSlJNrFlwEUP6vHcUcwSm
kVpyg02QLTEseVQNMYC+PTG++qYtlkqk8ibsR3JLjOp6LHnKXMdUYvI5jrGBOW4azhg20hP30Wdw
23WARbbT6ANeCz3tN8vC9BFYQxfA1eFv42vYE0TXrevJrdfnqwWpSnXSY7e/4sTYeC9znwRDysxW
F5f6jvFuK876KAy1xi2Qr7j3z0oJJaBgtzNNqMxbScLnPLCeaORs+ZZ2U4cNZuwgNJQKmfeNOGGL
IrLeI7YVrqYhGtzvru7qzzO3v26AH/NY9TUDSEN7g3VTLLLgTkLIhHkscub0wwPy0qYRhVB7NO5v
1Uw9WOdvCsk9jMAxeKrHa/LmUvlJGE3SAmf7HwjagVGJW0tqcfT/48NhIsHlvaWHTNbjArOGwKE5
mBQy0c0pstT0yiH26tC7sVzjYxGl4z3Bhkm8QUUbNbrx31UivXsZZQfJe2rVeqv1bEUojFOIKJtG
Z8Rj6tfbmiL1OMWGT2gDCzwYl3xS0MJCsG0X03xcM1RvsMA3D70keIvZCKgip5a8o8R8ieh2pOsP
MFKErgIf1+duVoD8hqYhRw6Chz0V7r08jASkmc6F2+adVrSYWuiEtt03Am1oTRB4BjFQaESO5c2D
B3Wz8Cbj/5f6Wg0NHEbThwzfA8M25SdfSrwRYwn7P57WYzKm72k+YVKBSkkS7u0djyqftgjkC5pV
PmFvdu7DbCZ95AqKQ+6xYLWyC0yeYvP5RoZVTYHOzzST0kbLtLEYSlqgOeeI5eI4U+uHwMLtT91L
rSOcF9RzekdZdeLMVaFUGI6a5P/Mi90+hTGqE/q6fuiLdkQgFPDkfdSTNu/wLIfSa8JPSn59Eb0d
45yV5FyxadwuVJtX03LqPssnMVDGu3ZAHrv0EgkiAAhu9rDcLbvytbPOmYxKG9ThPfei4WHdzj+e
zg3dwG3ydF5xKLDXUsaoxtnDET7W/EqlFCEGsxfUDCmOnP/fgwYVXawM6gStuLghjiUNh6bke9cu
nJq0cPrxoRJDF0zhvEt+cjW/irQSQ53Akw/nobUQbtkLR6rq+0dpY0myd258u8MSTpI+43FImDuO
3g98w6p8PX0GU5TYVrcT6wSNa525Az277yDjo09hMAUij+/vK/LdMD5GRm0duWIv7gOb5YJI68kV
25OymQxdKOwul8IBH53bnPvlVHoiA56ScxKZa7BJIGwnnoHFk7IHj0smhQsBvwKkxuKYPNnVWrJk
K259LmSkJpc6MVoduHmSFwMndTt5QdMNG1lf8xUwfL5UMW+N6WAnejBUYsJHbpb3EKJjkvQ8BEpa
6CCCIvWJyaRIS5on5vJHEJQ78zC4A4Z+duhN9q7UtwZYnieRX3gsjLfrJwrEnac0NuZz0EGV9X2K
IO2drMpMuaiS7NxlSByglFNpHiK70b6Z0m5kmMMCvgLm+24x0SDnYizi8Ag/4W9ralrJmEiV8ETK
a5huE0baCBzpeRNyt0UZg6jh++o08sfLokc/Wtc++ists16W56l2SRirjy8nNSMuVjnLuk2VrZ0+
6y1rGFRtuLLvTTiZ1TR1PtbTntd2wEGgJ7kdxwnh5F5PqTe5xsDIeCe6ngBBtWSDvjsuofWiaN+F
3/j9PO2P7KA4UFNSnm5IfLD7SKWlzcAyJkxsbJfzyWy5cJ8vflq+ojOsGCztQujIoq+Q/ec64YO3
dKBB80yIY3rGM3ulE0yCCx4sybPO3ntmCSOsA/ml0wzwtxbB9aol5o3/DwsXmA4nOUAxJWtTnnv8
2R8hko6Avy/79yBaW/3x06JkZ/WCJnqWtT8qkbRrN50xY+9I6nioYFaWVlrdLBZWrWBGh8nxBCY9
2M+SZWililjQX/rkV/YaijYcdlX55m4hfspZ9OxqTArUN65xW9/kD4L+wOoOCGc8ipoTDtKOxUyp
lAjuNfqcPgsTxhwYPTLBnxOJi4nv5iG3ug1358PUMd3zaahm4ssqx4Ii+NNsd4sre2Pc0iFBONnx
JmDWxW/d8HyPPUxkjk+5VSP95KBxGSzdR4otCGLEckGjZydVJEYMTEpWyycPwIvAtljzTQc0OSAM
xsPqpG6x+jvm4Y0b927We6kkxny7xXK7v/6mLB7+yE50dkfNv8IoMc4oXalgo4xkAKgS1qxjydeE
RNiIl0L9s7Z7sUpOoiAb+0uXlU60HikiTxIbmrxwzYRONf4IJlJqgk/IHgvrohy8bKx1rwQhIvzG
EJvl8yYfy75LNtAcqGiWG/zExHCz4eMqIhY9GgsevriQx7635OgSZAjM0WBLKHl/1oDOe4RJQJSo
ehhLHD6pVo38rfK19H/ghc6FoCq0vTbxKfeBsmdZNHCUXuHpPphOBD9a+N8CTu+rYEREDh47zLg+
mfjQQ0HRhUHvZSRewvsoLvMcJdDcnJfOG/9mjEmmFNoyWw1udggE2RZUfs52kPdcvwVg9G6xZTEY
ePxCakqycLwzPNo8mIanhQE6oVWKmK1y3UT4QZWkOBIcxp2fmqs5pIzIDXrLg4Wiy5Nok9CAoGqC
ClVnqrseA8/A9kjle5xcmKMf1bqqI0L2M0KVBv+zi23YcmWRA2Syo+UUfnbcv1qg+AllN1ED8fxO
Og8ghpTQ/TrPsT5HiyzrH9ByZPsRNsicmOyRQqLmZ6cvU4Mwj6+Io+gXtZINP1tDbe+GmokZSHfQ
SbJG5nkCJXAJMVrEwhai1H5HXMrH99K2U2mytS/ULE8vY5JDFdwNHVr69YiUCCP2Cv397ykFpL3q
S01cB2TnLTDVhuEfwkMW1UeuEZiyrf3BWAFRjIUwlLTlWeo+AdDKmt4NpEtk+j1rS1//MMT9LBLp
IBXyjRuReKXMvBfC8WlgRsakihO6yU1AWCaDWe8WDxK7YkfM2o8p8BSAJ5nHs3vgASEkPJO8Ix5n
fZ4MPtpOKF9/m9MvZx9vTDjR8i27FM47gij1Tt9v8QeMGLxBG3cPCe1Pj53rLHIPewcVAbWP8WDk
dHiAqCsTBEp7/RTRTBCLFBpgYHUHfW6iDoZVEL5Hm74FbgKkK4zQWMAfaALC8BMNHcLp+OMFSdk+
AsAnZpjupjPF1376MRbgodDijm/fARzE8MgiSAHjtltDdaYBD4yRrQI1BQV3LKV9fWTllf4lYeRf
zEp7N4xYjAuBWvz7WQwDLV7T8/14072fi8biz3qSjj7pi/txyCkRVpBb82KJZichK9G6vAKNyWvk
OPA0mlQZwNjYMDkSotenWHHIrhbUj0cFmjXVH1bkvpCgAjcrf9XsPNy821srmi1FggeHUs5inlxj
UrqG5UIyXVDBDBRmE0F0tUUCnSxaSwrvQ+XJ/j65Qv0lLgPqPCkKGTWEJPexcAn1R51PJcnKysAL
TC0Y8Xla2daKrWoBWXCPwjee6tXwAEvuF5xV3IK4yjnCsQaiXuuH+revnopmnuvAEY4CnAAceCd/
Z9nlYAHNj3bmH2dY7abj313qKRXKD508PSwn2+fUIFHhPNtj0GkWOPAbZJcBunY7db3Rt+GxVJxt
9Lzr/J/wNgxB+JPLZI5wzaIde99HzJlkyKqYBlFPIPBLuNpshetkHdbLQAs7D3ruqtEvkB0CdDSg
1rfMfy5hFSwwFdyfPtkWYx+16WcZ/hwCM/3a0nKO9CGqBcncnONrAf81ixSByU3u/cGaFuUJLD2l
BQpeXCGvcurw+spFDnpi32te55KsjivzlyNNI6SCR9T0r37cw1vN32cRSpezFE3Fe6DYDxD9GUEy
HtGcRfAyW4iM5mEftHBOS+3A59Uw4Xl8hJ3lKKIw3Pe+ClzZXK83km7f39aNvPESSpRxJg4/+/73
XP2U2uNWNHr9KUTtaUxALtSc/QZvy3Oxfx501x4kB3KDHDqnesZMp1UfOdExTBKVG3pJjlddqugl
UQNNHevh6Fb+WZQyM5dD6NWXzJkCBTQ/crm6VPgLq2m69i0PuKX4QhOppdfl7bt4dKJh6b7N5cOO
Su1ota/lIACmCMZQisgDsZUAatUvz/3FAjXJ8UUWG7FTS/apgNdOVd6czDqIJeGHA/wMEG1lCJMl
HktaO45zXXrQoe38rqar2AvDFyiPQVBDmu3B9hm+bxxRQ9P9yEkyYBWJFY5Qy9Fd9QlvUcDXujbL
rIcwDLv00iBzsTeA5Phn+BEwU2mBgqnOYSitgznhL+5HadpBSjjHhmb1rVM7BpZg4uQ2Sqz0TGqf
bLD32vYsvXRVTZ+KW/UBKJLsRVqiTWWsNPGezbvWEndTBcrRa7Ot4tJfv9EfwGwJ3imFQwBFbuo3
37KESJ328pj/0yPHE1bvDGqVjhpRrI9sTVdT2TZHyX38RK9dCgGTj1+xQwN/DIYM6mRLystpWPgN
zvQZh3PSPefng3a0FZUf3uh6YXKerKfsb6TKmmt4xpt95JA/mD6PZBWkGZoHW2aObOcj4+4tPcsQ
ltqcLTSf61RDdfik8jXDSNL3Qiz58mpmQTPep3wymIg62jxEmzZa9nABeSFvBTQn4xUIPbzc7IY8
MaRH+n2MxOf3++28ZYKa66HpoRGatZe8gcW72tpOANztHzHevw3CQ89X62F7JpO5QhPB51sdYZXz
tnWFvbOoPZiafEXJBjqF/EPe1Jg469nPzwKSZDA5oOmk8OnyQuZIDULhd9qVoBRUNnkvkNHkY8Ww
+w4Kl/psO69Ec7zdnR8py1Y2/zENXSfXaW1SESnIK271OGuVzP7ctD+ylX7LoszidaRqIzrg2G4A
YktgZWiAfZVLSjWIp0s4f6LTsx5bunn3dZRcRXXK5yQEyeBgX9cz8iahbxg4gFSsCAMYQKK12LDH
xDKCquzD48VfaZ6Ne72r3BuJeqwRF+0Ab+E0nYqQN6ocPSEdLdTl5dv1GuqmuyBuKW4iBOyJ4rue
ahH11w9y6gogIwBnnqESPzIHvKty7I9sUgEi8wneLTOA5FIHsIJm1X10FNeOlPBxM4JtqLlkrBpP
F06Y7Hrwei28xgYpHZB9s8wWt/WrS3beczSClLkX4rog58Yjor86R3vOGQdb8Bt8jSVBTPXnIIIA
TlETjvs9H+iG9fSlRrY3lfhKY3PpPh/KCQAoLSnyUFlVDAEgckpZrNzY3ExcUJvyjfpCxznad2GT
busvTcc1+XAnYxDEzAOvMzbZch7/tqScAD9Y46MhIsvFwVaBHemavf2g0WJL1ddcg4xB5AtT5Lzj
Xj8j4vVxFuTwc2wHYd4yM2oNjdmSYM4PB6fbIbtJ8qkvL2ydKE26LTrfd56xNUuWFOB/znABEctK
Ab+NcozBRIVf00ATdeI4A69PnPfkkrkKDQATV5ZNZUO1RRMLS1ribDndJnthdidC8ozJ496ep098
YgaDRWyydHDdO+Cmf6Rk0wUa0U4xo1qMtDkZAThmEOOatr1FbiDSS3j2EJyrtBV3e7gBYTR67CwJ
q6Ne/oesG/wlxhe8jxsFwOXexJdYhjpObHS4O7ovZ4TPtanb7+T04598nClnK+Fgyj3OvYmIZ3fs
nUuPbLCSeH/Y6qkpGWdJpWr5CF21Wen7EcwCMEnsjm14NTyIs5OnKv2S6Gw2ST3Q4mBEI+iYz5uK
xWn4E5b+dBr/3FKol7KNT4RqzZRvd6/9mVVvk3LCAKeXQwL1MVVnG4ThSDIPL/EHcV3pl3OGqhh7
7ZFUGa9m51/fLc1uJxqVsNZzK751bQPlmiguMoIxX6ewuzJ7x+zkssrMpXqymgw5hPvSIVnqzzkW
3vuWakP1DTR9ugsRIHnlFJg3NRWs96mvVrvjIEbHqd2BaIAI9xOeQ6Pmpb/fVRsfjRn6y+O2YqDD
OFxQiDjQg+GT1nZ+bbPbTyiE1z0vFxlZMHaf31skLNHhSc20djoFbQLDRI1/qb/tXGrQNp2o5BOW
tsIhnSkAXNPUXCzavgT3/BpZsUoaWX9oLUBIaX0Zfw0hvhCgSv9jG8Dx4VOZDFf1BakD+OnsmtOQ
r8JPaoolKCPh3/UWkxQGEcMrffFLrxb9RfoSKoyTmLM+HJCulUYFmO5QoSDux+I87MPyuec4/vvV
DpmggkCG2H6ZajuIfTHxAUhK0DIbLDm5+WifzMErRHIgffoCvuP32mOD0mb01i3Rdsljzc4fiWRl
eAed0w6PtA9b+IYL9kFiDmWi+r/pfrWksEJ8zwzI/66RAtmImRIkyKVd6gcetfbendfhIjZOLcJ8
9khCI8c4wZOnVoDpzs5OT2TgXaHOWlY8FgVxL4Lc4GVzyR3mZjcV5VYmEXfX2IMs4DB1VHA2hG8d
Hd9NrqajE0fPU9jJVw7rfEstik5ClUMX1Hnz/csC6zNrsKm/2DVN9TkQnQ0QGdnxgBja4HWG7XNh
MfD5GhSGEO+tP/2NypkxHBoUNvMJRJ1jhOSguBVDB4hDFkAmkSCT5iDTebM6CZ3GSqOfku33AMa8
YfiUVRSkkHLpvBePO7GbNz37CM4kCsqPkk5uA36B/qN1qVSKq+7aliaJSDy9X4ny7Pn5mPhNLhDw
kuf7QjVkY6dIkK5r8TxDWiW2M4m8fvMn4QK58cventN8gD3qkE0TKUe5YLGeVvBfJzTNjykKzinj
swX4MmTMiliZP8r6I3oIUpi5UkpFcKzsZtl3Yl3EgrXhZe1wYciGxV2HFdoiHbbH5boTPjYnAOLL
6i/aESEsbZ9PHtZqfov5+FieCjl1wKjRl4cw6gC0Eif0XAYlUPmjM3hBh82OPdVlksKEqS/+iKW5
gkmWKEYMiTpWxs8k1nuf54F5t1CZS49uN/QDb00P7yye9GUKHHHBOvKNiDrVwcfEQG7YlnLU0S5b
FPjs17CvrbTMQaJG2rqk5fNYmZ+gA5MbrVcAtW9DiSO7QCxzG6N2weRumvmIAkjQBLoGdH7YTmQj
DShpxSM8eCdYx+krHI5WA/CvAwMU0Sw5Dx9Y8+e1ujUlXEPUg6UHsFtqcsxTxqc8/bOz8NWzymr2
hhEDgsatuLgEq5aotrUAXT6VhJYIXMA2YhpqXhufbi99Pk86PZ3MYcNRDNm8aifBMQ8fq12JSmlV
wANn8fiugNEhplbTwkHwjR2Qd1I38sh3U4fLzGtHQXcnTEQQ4FMZNgQ3tyRLZw+zCX9SQYgUtQk6
wS/Adk73ERQ+W9fSjxK4qwWK2FErkh4HmZ8F6w0O/Q+BQjOE0zY+fTTUZFHxkxxEXVm5Zi54eKoh
YJdKbIweRh33Wt2LeZkV+2n0QNOZt7S7p+1+5JqUNjw5dCT6QZBMuqDBdV1palLNklM29SUccr6i
7Gj8SZFWCA8TlD58oes7BIO+rIZJbxCnm2rBXR6KMY58/ySgWmWX3LL76YbUdQzINS4j8+REeIsj
EffzeY3nZWVXQlQs+4vJXEkkExfiZhRVRRAryyOZw9uktmdQOeEodJosA8MK0C6a+K66FvCDBrdk
U+l9Cd29IrvNYBw6hvIYCkLKJx1hdzyjVeoWhAbhGcfP/G4Y6ANsSg7yPvY4QLm2u+7X+VNFG9MZ
8JmeZEd6WW42LocwtoaDCiYyeDFRWjitwxPWMpdSXgmGaMJbVYzdifIiXXwEwVcYdrDbABNSD/H7
HJA9S59ZuNM1mMetLO2d36G0ldN0qswVipLiF8qErkPM9psaxJ2zgN6Fp4l7jdZBo4JpYIun6q5G
HT7qhvMAgjWfg4PqupRnPJGGHZ40WXiZBpxa4rqBHwdBTvoFNpvARjeu9CPdG+WEpTrpMtAd5hik
sys20Nk66xoDK6aEWwzOvvSv5oA0s8+WRXwu5gN2LMfR0CexUW395TL5HGnWrcg9EtAAYsPnJuCO
/QaOsTd2lg9WgSEz2Hnq+t5wssi6AcrXHRotnC6W/qFXQkDja/Zy8kbAojjiNW3qq8SM3iSMEFaA
qAtj+CyNXDlRwLK82tiSkarHS3HUWMN4vCK85TO+RV4ZyQkkKVXwyxx13cOlqT3aXu7KQdMdIaOf
vCLQRQ070dzjycXrmWYGcxO0xm8SD2rbU/rU/GRXM4ZbR4G0q/1iaFZsjU+If+KOa+T3gC9OWmSd
kPsBoeIp7Ke6V4dD2FGXwMyI6zu6egg6gRiC+ptz/56v9wtqMDQZMmJeBfTALjU/fOtO6iORpi6S
mrd1+rWOyZR2QjkTRMqtf4HJQpaWA2hN21WGiDKa6QLauN1Ti0pWBaz+gcV3jdKg98f5I0sEyrqk
KlfnmvLAUF8tPZZwwK6zORniNxPEvuhFtzNpcQhSj4hdjnEt5v9VzzF+ncbOME1UO03IuuDNVLYG
F7WL8NL424+3Su6lG7m+cwqGFdXqVQojg8xGefspANZkDNTathmIeR625ohaHb2XbMuhv27P22Y+
niApWUcNvCEC78zha2zUH5F0qOYYMW9Zgc2RBnuF/fir8kIDqsU3RJe7BBFQ4jCnwO1A5TkYZ0Jv
u9h4Ta1VCbBxvMk0KeXUo810jsftEgynQFyys6NyL7lZHb7Odv/UEvClo1KvaP/dYi11QtiVLJ58
8YvIAO3XMwvcvzJp4cSVOc3FCsz0pzhOL4Ovx9vzI5mxDugFtxrLYIjBEOa08y2ydTVMvMwXAcCn
kR8WMweFwUqUEzQwTHa+uMhhDhFjYGLdpqiSH6Kx3z05cNV+/pH3x3OGglNqQ2g7dxB30CSfYGKr
uBZLufSi5A5M9E9PTXMTWTQGXpq4eEldfOfrLeUb8Tc25787840jm5ZzdFoQ6F7THin9760gNOvX
7eCk0W13uIex+6v26i3NfNSwk/00MBRym7XlDyK/xhMcFvqqATi3l3bTMzj15r1r3t22grvpNJeg
S+PFzHqx3HnVNtorGXQG08CECw88w3usO4bLdlDnDr08/hxTEgCLE3kEP4dqZvOYY3xwJGEsV0ls
+8PW5fqwfL0CW5MQOToqbgmW5DOLZ+wopxVu8wdhcTovvfJkLuSja36MKJu4NPg7vL1+uEaZzSPw
82k9dp/MTnXsb7/SVDvpMAO8LtQUinDupKezU7VvUvDDRIs+ifiMKkBW+0Q7mfcF+HYZmusugT23
vnAciEf/BwcH/k30AJRPFtIfV1jEAoD1lNIE6Kpvc5yxjHnPaiUetwynZVi6KzmL9I36jLT/Bj+4
U8NE1aT0yv3Ch6pKRiP/hI58Wjpg8K6jKv9F2/anyLDhJu4nHUkz6zZjE5TSmVu/BCaTASPghpE7
ndGezcUnDZ90oT+R+CvMNvaqT3FGWSI3J5XIph7xUo0VtXae6ZkxNlgWoHdIBQDsPn6yWhQH1XWL
REyunBgxWjJgoeKcVrPVwMeF4Wy6kL3qK+6aCmSwMR+8VQdjmTfKiMYM6rboQMIYJQcL5eqj0Ncd
x+wBE4wij17xGgDE1WioXDTk5eg8JnDolAjVBs3O/ymxFdUUPf1wIj6ESzbBHcCWdEl0qReXEd3t
OGCU5BYvhNe5zif4zGgpDP20ThAt+rnNMzdTHH0HaKUtlll0RWnYu5fmym/odlsu0BGCFq173sbS
w3YglRYpOMT9PdMZ1h2ix9giCfVQu5ezmD1ikMSGng97bU/Er+lbuuLtJ130L4wR4vohgWEChCwM
x+T8rW0R4A2jXVxVcuRaD7klQBT1JwfeXI4RbQYAOTFl9NWXe4W3t9nUPrvIZqYXnngJPOHCQocO
UNjJ40asPZ95JlAqCfdz6GcwYrjV+J5EetZCotuwcFV6emNzCjp74NajjdjTYsglsfAk1PApsSV0
WF9KnTU3zlU84TrqMbmwfmrXNSr/kwTFFLWynyNKBWZzucRt2vv9L+4pmNdZ7LJibEbd5lxHJmMB
hF+JiP4eCN7t92uH7t+9HmvxZpWN/Y0niJOSFOyzfdMZFUsLunI7j68wnoQugxC/CP5JvqIWYYwH
74cmqTqkSFixTKXTp7hYotf6melzzGfGt//fjzQYKrUGjcivD8DQNQMVZk5jDAjzzRwR4Tam6ijm
KryZTErB+5DQvNLVoXD2rum7Jssq7l09RNLAOd1xvYo9iJ2Y0Nz7XMIRpcZ4cvKju/57Eio5hcqF
Q8xhdNGG9cDqXEugxX47p+kfORkscmM3kU6zreDzjdCkw3kBACu/zjl85gyMvxtrRZKZPk0v/njC
y83n+2ZfwKkgUk7lXnu7L6ERuvpqkXjDY3Ya58gYZxf1n8ldTPNjrs48rltd6j8CjsriDaLoYnYH
VRYr50qsGjv1++J7el+XXyFAVHgI66BGSKMdIfBAMYWsn6KfO9vF6TgTeIhuRo/HNwS3WzEvXOIT
CiDQbyL61CmbQVO9ObZuLAt6TwMYR83/0duQr6+ur+dseVkIZvX5Gl6iYVXMW/ScwMLllJvckRcw
XX9ue4DO8IDtBUTtQkjVJqKFgn1QC7Nn0iddfwQuXRorg8EV52j0KzxeQQl5U7iQToiYYKV37kLU
zrxGfW9T9ADLu76apkVu7QarhPAWj6cgAJUdDcmkSnJLBqaQBAcP9G36P9zqNsHcXTY74TOg6s/3
QJwsmlPIaRGuCDaLO2LAIutdEuawejeSN3L+5wPio/ib0P3Y8hFBNwM3iwcPwhWA8W93OuiLShU9
fISLuWvGvV3zq56v61gRlffOqRC8W/zOLnyqVQhNK7aU84pksL4K1xduyDH4sdf+vDso0OHpLRnJ
CrDSr74wSAyvhy+xehsv0Mr9aOKtxFYlxM+W0Of31vSchpegvjb54q2vCx7R0pPHT4WtCfLcKVH2
hPRHB9qB0QAKl7/P6dXa+UoLx6YvuP3uQzM16g7/JBu7eDn06y6aAVJ0ASxtjbuZD51HSHHuHl11
f4plJWYixJpSlpXmDGnzNz48JQP8pVn9CBhCjL+Q+/RbMKIdFnZwiZ9KQtH1NxW6SKUqGRX/aeaE
lpBT9Iq8mtr4DGKdFDsqDFeKBahWM1HVP3vPwKdZKU2eC4K4Fflx9sxnQmvi7QKOKLIBLvT9jrCB
o1zPw6eBFjatwVAEKDJYNYUIq+MEvCw+4vjvyTusfFOk4cGHKH6wlBWHvCWwRbwbvQ0fRBzUs19U
RJEkm9yC1SXJc6Cr9g+PUt6GmmslzBMUMlnXAWunUO9Y1dIL1AFZwn/LNdtcS0c3ZOr3oHx6gg7R
2u5bPC4HdavTO1luAr8NLjQ5F9lm6pWAc4bYgIlFnbF+VrV5tNreU+M+IL/+O0NnpjKKhpas+I9g
YDhezP3UM/nG1cMrWisd177ObP8IoSMXdvBBEbpGCCnm6m1+h3MaVoaQ+K0y5PDj7c5kAKWWIRwM
VGkkPKzhn1uBUTQtiMss9ibLiguLg9lzmOogCBvTqa9hVEDR25Y1E0VJpUcRJgBmH23YIOwqz/lU
6I76VZ2rL6W5d0Nrbf5wSoFNljOuDjiiR8g7uBHYacOYdEwZy5QwPfbtkvAfay62+oJWCVIqbC5K
IWSGmZrDbWIwc5qp+X3ld6p568ppEACOqZow+a88LDUkuNEWGQsnwfDpW9aJNvrE5JNMH7AlYW6G
lNfGUS1cxYgguW09m8i2fLVhUJyHZl79vhBwgD2SW8Q3TuzALJgQ1w8BFKZ0Q5PTVpOVuo+cDsGI
IWt33rnPGQbgGaftwT8uwLTwAknK4z6wq+E6N+ylmR6b+6uw88RBgIlU1X6uwyDgB4/n1IZGgqHm
j1fmm3YKde5YHG/z9aIUobSAi7oUQJ9gb4UVyNZmagAtI6uCge6kt+vesynb9T27adcB/xV6o8OE
s7jZYskporFOI5fARdhcE9rF+F7v6wjVG7hm9nqxu97rOnxnZyr3ByUQCT2MmXNnunPNAuRysg/X
SGOJAHuBZaxUxxD+ErVULFDy0eEBgBbrap1dFqKEaVUyiigOq6DRNU+0Z6pfShNq9O9jMtNYLqed
T8FhYwLwcBTEpAh7jNzkYE1QAMbFO2VE6S/QXgZP6fQdtUAY2AmhZNEvao/xta+tQrQWpQDVxeQh
BAQVuGdE8Q62WsGxmTEkJoE2VuqBWLEVCOczRZM5A6hdAvjzgvohAf/KcDjRRaav1J9ixhgDSNkC
thCQIaMnYEXecAYGfJZ78vmDwOd3JhjB/l3xqhnFeyIgeVxMCVti/ZVrvgFawZWVqhrqHUrBgM4+
Bpxcw2xTbbDlLhCTYxi6l/bpz/3e6C/LEqjGmb3gk6iBWIyP0DKrq2gPSHUBzIeyfRkCayR2cQH5
JwawZLJbFEEiKf3or7+n2z+p9+uhB0IK8YC7i3RE6p9OK5F0gVDDAAwsTYuzL4vZhNU10wntmKwL
3MId5531L3qhkXtjkPwiHZ9sEYnKhtg0NbrBux+wS7i7x3O5rjjJHa3wZSwKlBJHErHt0+iSMa/O
MjxboQJPYClYkaJA44JzFrkxOhcEfNBWVqNokwSNGH5dizJpME6O/j2+Z4OGpV384MJO2CSo44pF
i13NdBIL3U1M/9tSfyWEVU9n39kqgwKI67SVutu82tkxnw7tMnXzm1+R+Z7cEUQj+lHZ3iakXhyU
YydhCPcO9qn2DmasYFXGxshf+MKWRg058Nr4ugSVEIUqAFWt3N5jDNzYTD67uJU2feQtxlqtKAUE
jJvWXiueSdmSBQjG3tugqITR3mXk1B1CabhYFrF60VeMAhEGQFvZfPltIWmIjFWsFE6JV3vEVc8s
QVVOHNHAO0ueH2S2ut9aqP09y/EaJe4RG8a45DcYC1OUEjjESunIpDmzu5l9czOW9DjuOeVcqTC9
M1G6DBI+n9yT6u6epqAQ/ECrtOWH5Kh810YvlNcDa47FFGGzxAcOijJ4VOYo5qacCpiIRXd8TsN3
5G8Vn9Iid/qKNC17/V5ymSkpOKOFf7GsmPiLUG0LZzcAXl3EUvwY5V2Al+uLZsOBtl86UG9D7iHI
moWZbhwl2F6hGjFJJIErvOQ9GZqRZxmwYjiaxa1CL5bts4MylkyYoytHXrcJDEK0IH2NKr+t02Eg
W1ClbyNLoNe6t3BIjL6H+ydfLQRbSBCKM4zC2z0RyIQcQJ5b0EED42qfozhJiFVzJ1e08FFnE8MG
G6MPk2jYwfMuJjB/jf7sVIzjnpR21yU5j+W79KeNgS6sCdJ0fUq1+lRiwHpCzRcIbnxfIJUR4GAk
MiykvXJGF7cjblYGP3MfQAnQ9J71f+AuhEmpJ1fKp0Cthc9U+dk4az2B823NgcsINpci02XXKSdu
1L2YXOhjBtiDgldaGq8nGz9314L65wxPINvwQt3SAifMbCtuLLrGI7oq08P9w4KqrraoyAvyj+pv
3CC/ciJYJoypT8Cg9Tsj1m5NrfaMsxuRB8t4Xh58XhoucbjNj/M7ZARusWvvGCa+ZfZ/SA5A++mw
C602zogbXEtO4LqoIavkgt1VeEQP0IE/lM5s8P3X3gI8bNozCwSkQLlEWXiUo7JCsTRy5sZlxq7B
eYEsY2yyrT8BmQKKE1YtdPdMornP8PCzXAsY9V9vOO8YFfYqJxKOBUnzp+Zly0XFwiI8Z7MLTqY9
dKf5wNMShMfcUZbpSdGHkgxdzg6gCMiVrjc0t9Hb6g0p7dWb8PknAFRHcYCzniM3PifTigWBBi+C
304ZE1jOGQPMh4SkyvvgHb98jYL/6NIUdyTM8yF9eh7SUCvovciYAXVyq6LhJIqXY60yzZ1OxbCm
Y2WDCOiOtaXqH4wyqCI1pafZri++Y4ebqUm5ElHo3NvPGe5JmRxh1H+DtfG3EJa3yklGAlZ76ASQ
G06vPjEJaR+iZFalIktXVZxmp8QqaBiNpTkH/P+Z0Iq9j4qass/JpsUrO0k+OZkhgd6CsTTQ3CRx
JOif2OpfQ962T5zaVzj36izmi0reUjoh+TWqABdtdzc+vZPcYOPUb5xeCgepAjvMi3DopH8iwNz0
SYNynEhSUnpYz0dYDrTEsM3GFgfBubiT4PzGy2qvpxESj2bf3bxvvjLQSluYXxyT4Ow7Sfd99hm2
4g2h4/M+HC/3Aj5ArBQNp+1HM3+8KKXfyX4p6hz4P1YICH8JsbsSN7sux/J/qUKXGjHxK58YtfBP
EWole6McrEtRhasyOliAPoi0jmAIXDNhLsgXG8ZuiT2Oj7CmI4v9nEb1QHTzhfUfNI92TeNnCA6e
V2LNUgTNWll26j9Z3pirrd+kdAcGSlESsBusw5U/EBnibttcEmQMRSZmorXeGN9j0wJvTYWK0RZz
WtK27G9NmBJd49Bwr8EZqtlTEF0i8nJGnBJ7N65aYLYCos5ehehajbxhyykFWCJs+PoRo5VJLNW3
TfY2uhF2BuxsZO+rfL2QgMGqx/CXesTL+zLYRaySfwoh+aRweD6KxI4IPi5YlZF+k2Je5ug7nUKW
NP3mvO7trmW5XRIfedMv530WVkEktzt1qvZLzv5/E2RKyGp4Wd3sNoa8Daaaa5EjSDwx6yLCHKy1
SUKs3wAZX+L+E7XlwX3l/ClC2lSNVwyJvaw8wA+cBJgEtCI5RVuzq03OUAWKf+MwM0PnFjg2POtH
5FTVg61lnSyxay3VlZjjkOZCLEROWPnvozPk5GdFiIV/9hemGMRjmRL2GgQw8oAyNdpmDQRH/WHk
YlzP9sbAHnEcYVa411svJgyTR9s/Lw3OW72W13Zpvxj852vD2my+UQrUWNPIw+OTDHl8UpZzfNAy
FN6velC3WakMlfqyZoni8goqobCDdJNvPgk6QoHMybKIOlaLFGFq8OCU5miKle51a3Borup/lF56
FY7cBG34tvkAGcf8WuCoKAECNk89GG+FM9g2eth9BJelFR0CF/Jc7p6pEBTuOASR9MQFIeNJSa38
kfT7hemALNEyPTtWb0MSjeHcZkmgJ/puXBxFQoAKe7CLsRzUa1lQRWKD/Zn/7ZlIbcoOSu+ey4/6
jzKy0pgorEkUIGs+Z8e3UVLZtMuM22EvgO12M1X26a49dZRMWpt6NkPMCFaKzuX/H0899m4Xqmqk
vB/g5HtEpTVU31C5rH1p73q2UL7vHLlGGaiQ1QtQffhxQAVuafsHiPH54V6ZmdXvo70EFrMqM0OZ
xRR5uydOkyJYwSpQMNRYU8lKoMbdPth0obbETIwv4vXTmwX8vj+d4paVEWbT4NRaX4Glk9t6rGtN
+tpfOLpLOgoCbS7hWRIjU3Bii307rf7VO8F5CN8IwjdHi8GXICULtTS5ugU48DWMbyG6yW7OTcoL
Mpd7b8wvUjdrnmh3FjzkfrTzi4CUzycx3K7buIGAtuZjW5Gyf1t4Kfr82HbqD8VXJKjrXJi8tf+k
8hzkTZ4UgDuPucboCRep0t6wmM9qeSJz544QCbF36hCg96pndSqqgsiiW+s4Y62EVdQgmzInBej0
gforoclJBqMKfp9qzzKHvVxq/vmx/4Ir+jJtvgUEkmjKnbELFc6s50fNVjxraW6VyrPSC4Xfg4Pp
2iaYEL1sf3G62dN5fgzyN6AUp1+4FHyXH01519Is+CvrLV/RyqSheTvtl1qU/FzR8YUiMl6aSS4j
n+opBp/zLyT9Ay41YeB8c2T+XqZ6/SoVFQzLc/YDSr6+M/wNEvWeqCprTnq+0XhBFrnnaUah0paY
mFHn693uEMP+Q+smkPlPcAThi9UhFt52+LLRxDCtaZgbyrA2urYZZVtqOoRzFdbwiEr8++k/0LRG
BC93XnvRANM3NAbQTtXZI8zGxvzcwC+dZtd8w9aO8Jv7fts8LImvUxFLcqduCxAO8sgD8ogGA2KO
NpmfJLgOCGYHdPPBVCzrJNMo7kdC6CfIv5eqnwLQig6UHRrm8D5hUqudNNkYwfOIGLNZrz3TtiXS
6vvtaPz2Esz1jLe0/K9Y8aFgdn1xKQ+hQbkEexAtpCMDHFkxDues+01Rlg4bfMSqUMmjFTaMhLGk
Jtmmo+1aqz8YM13OYyCKUiziwF6Isl3BUtKp4fw1dgMIT7pRCUXzhBmxoP6tZ5sXjb6FIFTr1xzd
fgmBHkfuRtym+KDzp/yhN0kHOiwcMxc8VKS+tO0UFvsKmGqGVCwfm/gu6pxbxoUrxZMXEPbrjMq/
Bok8tq2LQFik+z2yBHPlW6x1PAxBgsSN5MdL5O9c5yrTO9QC6819AFMHIPxRz1/NPSc4Nzrw2Ycn
rEfSl1ikJcxGTS9oiMf8Q+KFlOl3DxHIOSMBgk4Lg9p/47HOa+oO6SoeqdhZ3e2Rb/jBvySjMrDF
HzJj10r4DwAMJzgFHCq+C0gRQfjyAUyvldbN9gNPhlRLMwBc3NFsA2MR19Sj4kKfxG2SINpDE1rl
2BBzvO1qW/GlVq8TA2hHls4MTyFe+/wLobTwr1wgquZWWRmyojR9LduyZwDit0z+iAfmUlmD20W7
WLQetJLOhmOymrPuj5Qw3fb1EJ8KOlLtchtnagUpZ7xvLlxkRctQ4U+mei0uig6UvqEPLGhClJkv
/qgGwX5m6XzyUczy8p2xxipX7jiuea+In8z529LPnoXKeSZG7qSfAGzOJ77igHcgfx4RXXArwCnz
zSgSPuntQFY32cdEzEpodboFhb64/sYvYLCYqqWq0l6O5hEQtsdCjIT4u2afYLj0UxwpWF1Riajr
yp3JUDhVvYraAW43pIRlIaLnFAuZHE7oRHXjvcW2pHJMrdZFTBZiJCAgmpqyj6YSNqpLJJOozyTi
RJP6KkV40tCn4xKiboaR6HyR7yzc6eq9c59wLXEo/U8KkXQCvg6elbGyBw9hfQxwRqODviilUHxn
cUatGSInvWT1A5DHK6TIHbulIaJ77p+9+94QtFx9PQzsWbv7kAqMB1h191vzx7UamsBnaDQzDvRM
DlVsbKLoT2ymmYHSMD7K7w8GSao94y/VKFxOh7JnOGMUKtj9aUjtfTs59/yJz8UEKCe5wqT1rXVv
AQOm7mdtMWYZhzVIcvqErK+2a6dIk2t6WsVwV4SQ4qBJGdwD9KLQeGKXyEsy62mxZ+quLGCjcapz
d29Z2tc4rqhSySAHu/OWYmTleAyFK15UFZo8DNTtlm6LyLfv8Nq6ayoQcgHdAHGP5aaQ/DDXCSie
EpubNo1hM0y2D9vIYQ7xCtQ4k78veE8U60V6kgj214pCZuM45PpLqMOFifU5zs8OT1U8jGB4GFyM
9ZnA2fguWyQn05K6gb6f9D4oBwS+XyuWRYo4dJbuH++K5xQ4zbtNvubEwo95i4KqPUD9GhwOuWO6
zpfMnG2TJsPvesaHKcL0HyICTjX6ZNR9LVwspi+dkMv8hpJqzGJaau2nkHvBadVxjZXOM2ldB/j8
D7+iZD0BOpSjRztiBDcr5opjdvBnimGhIm+IWbZVB0U6BrTNDRSl+DkuVHd/8/v62a5OSuBXhlhG
ukdLO0kQgRLUq3nFVUH/BtxFNIp/tPdMuGMq+dImpLfEzYF1LVlnvQ3yrO8oX8nVK1vvUlFv2x7X
dnhzfQkOkvK6z2ohen2VyHk9f7lK0PTU9LAJGhpClRGMcms6n3Wg7UI/rZs1yDt1X2oso2FIIizN
kFKS+ycAu1HouFupMb5/KTSU84vTXL7+Jlmn9mIhcd+aNsV6rMO4hewsy4RhKsj3Ua73kuiKYPaO
Tn1Ycv4h7uyJli7k3PkiOP0kBR/H9mhbZKjgT9zFZULWhgECXauUz3p5+8Rq97iVMMM6KykXQ5eo
4b7pGhpzQKVt51hSzustL/DpCOkTb2HOvFN9DZQDUyA/U/mdwuDxOP40Crb/h3/qCYFvqMEvDkXQ
ENx/pcKwRkuseDF/OYPnGGvsmR3Q7FWW5EFQD8Ua8QxpXV4Qq8KVqudp6DYroOI4FEmxYQ2lu5Jb
XajTu1H5gbvahBmBtDX60SR+Mqhs3o8ZKDGObfWOMi3MYPlrtWce1AhuZxOiaB60A+gLtE+Dd54X
U/6jRrBM772LVt4i6i4KMEibAyI2CP7P4E812Mx7f33ckQ9HZETPgZhqv++f7wYESPOrI1dHA5aZ
y9ELY5kntIOX2aKC6ONpiPxetbGbl5ArLekmgCpyyGjDDbCmhKuwBTlz7T/qWGoSeBk1Wz6xDC8W
HemdynGHqXkihUt/8oe9ZynNM06eMENdvXWzW8Dn4wTNuxFWF1Do/Kd6AKtm2tRaPkOPNP+uzJ2x
A7tT7TFGcuLCTsJOkMQNOERM2GONtxvp7xgJpyfTyNUwTVZ1I3YpsFuJkS0Uw9FDJZ+CPdTtspII
KJRyVTH3iPvV3G+xKMEjtamDTcIJr3jDArcZTQNSaNALJqL+e5UpKfoFyEigOZlLGqKyw8U1+VAE
C7t49rnbW24qifBVtgR2CCTyHHJqSnk7Vj9+kLdzRimxIDQG9ybYHFFnusOElTdAoLEUMXfpDo+D
0ywtgnxCC358qGH5vH0PrxhAJ4DgeWQ66udpYC4RnQk7Ma4KMQXUu76EE7YIOrrB+4r9WmOazil6
//HtHC54dMiI8/luKIUB4DaCmhGtmCXNEkQrkNOqkyed3Yjw7+mVl7kPMjJTTGkfNqk/0TuQgqb1
ERTzlf8ANMvAIAk5VsZFL/lTKZ9JzktTAW+T3NEmONfefB4ArhyermlLydtdqRBqCt1PjzR2eh6Y
/iW6SiEeH9w1V6ek4gzNAEX3txlexTmFQ3gGlOWLUPSmqtVr9Dz8Avs0UTTTF9DXiqBMl6xT7MtP
FZwAI4jkEZDmKMh3aJzSPZxymPQwaFaVoTV96bgqwwEK+/epCqKVWGfHtfNZrg//0AlU+17OlmP8
9/yty00UmFBe/55r9kxbsy8uCe+TF8bDE56vSe0mS/4oojZqKO91bpf/NNSiV9Emp838/7xLWtUf
rAy23RiwrdMqQitmC1iES5bAYL/GWPwYfnZycMPgMTBSncixZAtiV6AjPbFsBb246SxW/2L7WqcK
miKdH2zboq7fLUVVEkduYLBqTMNP1aJCsuUlkeWQcgKXIKVcXDbPKD7gqOGnEneGT77YXlmTH/3t
bnVvoZxL58XBs10DoH6En7tzgKQCKF9ejfq2tBEJaylpessJOWHGA6TEuDu0eqlV6lWi2Sf4ms9P
H1Fo1Wu6Tf5vO35LQH8m54j5OjIvg08PQAqcW2laiAPssB2FFVF1pZI+cQNc66ZhjaRmr9yQCvNm
9alnXWFkqyVWhvOhmdUsSG96PdjeZaU58M6PbTstIV4ZRRQSfYwUPPEWyCOVcRE2xg4eahzDTp2c
Rt152V81Ftb2IdmxYME07/bgNs0kI6pTupNBuPp2pag4kJALJSixhvKSW1cAFFtrbjzJUHY70aAU
tixRqsPkEW8cNX7O9WhN9/ec/5F0+ns4YXx/nNzklVJbv/OlhhC623bAOJNETFJOhHyrtSvkTmab
fDXHqKju8vxNUP+ByGDVIKBZ0zDBFRwtoGKc30var4qYANShzC71d83nw5ziXfc58Xlwg6fjYtgc
yPZIJg8k4I+b4cW7mhXzkfNi/TaEiaG8o6h9eyDLUSI5cc8ixzudIs4r9NW34WFWr5loacw/Qw/s
9ffvKEVLENhZ86EVPoCODAypqk8MGHmFYYt1YrXSB+HtuLgTSAyRSUiYWaZCVN4SctkOfw0EP5qA
aL9VLUjFr10TbE1Nc+Q5vKqwKL6IzYXpwRSVNo7GKdd/Ok9hRKYttvN2nJvDeI5Q6v5xjv11M6v1
Mr259b8W+wmFOEFJQntsZVRBxfxqn0L8yUyYCwhxBxUmDtRusjDUspIG9w35tHqeEXCU55LXY3jV
eDylVwIVlFmSTl5ImtiBYXr6ftRnuEoskmDhudqls1U7Nl+DmFWhzwxS2PjpHmdjjXrs6sKp9iCq
KP8nUavmdtMBUtZXUCDG0S9LczgwRqizF1fE2zAb1H6iSSqOSC/HdBSx9LcA3JC9vpDAp7+BbP1A
xNtYKaZO7v6YxFHFaWGH+FY9BleCUTCVHCcnyqDBUE3VYMSuU2JR55aW5NJoWRFpIrpvTebTzPEi
tbex/7neSFeJiZaZvOvcSt17E9eH0tuu7N5ag4/rdhEV3vlGJ3q8tyMTurDSiDj/LRSVHv29U4aC
+SQes7U+sZlbRY/AoXOp7UXCnVPbpm556KLlrDFk68v8K8bedWR94RHt6ull18MMgyMXNWRkNItf
ACslIQETTQxb+dWodRAUZxA4yktaJsFH78SKJSyVCjzBbT2ZWScg5QprgeEUdW150rdgAaMXfglI
16mW5/u9T72+2V4bP7vvppLteE7B3QM15MOCUQzuWBQGw9UPFOjMkg8ZNK4TWa52LCh0wnyK3OCt
cQF6l9oCe4kymhzq/lurXB8APJseBuRJZtPPZYIqxcV8K55tFR2T17+Su6hJwQPR2ees946bpvjW
FWlHGKicvs3QnjEJElpyAwiwjgd91GiQL+P6WHjoJX6Y2zC6bLuiah5NSreGhP1t7i5B64tjJ0EU
3rEnHcynRfI3vHA2m+CsrXc6fkpowIAHQVALtFppPLcmqQpW6k5Gp6cVCMNywmz+wWzNcRu23Smu
CYhVgv4GyRiZaYd0bnJz2cuzzAkwE60bQs0Birso4BuFTUocVir7ALMgft2vU41PADolgb4+lxat
6eteI+E96I9CWucLuDMEDptI4XiMUPW9i7kOnW4SKsQvnlUsc9++/LIvnZUJ216evjL1WXACDd/f
oZZ+H6IT3UtqjqLrRGD517ouKSO7wWfNgrilu3FqcR+/9G7YDGC9mzEdQb2TUxygyIO/XdH6BW/1
OK7k5wKIC0s5rRq5AjTXZl3vfhQ7VduC3/SmsV6ofbybUgYFeBjbOKe5Dj4hdGj96om1yznUhlzJ
9u7/nD9bAApsTscCgT7RmBCayt4qsFJxvA3Gsk70xPt2aFDuZK/yX/J+NNZLhkD2taqTglnyiohq
o3E4ax9NNIL7mvhl7dTR15+qL0kQ33GeDQ4GiblwjHe0RqLh/uW98szd8qceAsuscjT04vavdnk+
OC4zKIDVAol1V42bboCR2QppLs5Y/Lb/3O/B1z7mhgik10YxkVETtu+RC5lmpH3tx9i8C7vrq+P2
a+1I2rIBAaid80jDuLx/BdggluJQRVPnaRgq0bBK93o4mkqb9tQtMwNTTO089GdkDCOKBfWy0q4Z
35pB43bOU03AZVIx0uEor+MOwF++i47tJkM/2DveStuzbAxtaxhzy4RHjtfkyRz6gEzTxqcSX+fc
7PO+PKb+5h/iU1oxmdKd7L31vcD4P622mXoG4uw7Ia17iF90679w45S+iXcEAs3SomF8WlX92LdS
Ccd5rCbffJHOLjcceLHCX8Yx2XaJ7w5RQEOOz29yJoat/ZQSnMIOnl10qe+JK/gdQ7O0Zat2DMmF
N/P50DIESyVKV+Tjx0HtJ6jrme2Tj0+GTfnweDIvqAgXe7HtTxK+Gtia8nTkIKi4BLbUx7nI7yF5
zwQbpgedlWKJtsPPSenarJ51d1b6kZwX6SJ+vukV7aORfcUrjXwmLZiowGb1wytZPSQpnPTKm/Sw
opUba3FMzsd78hkS/Taq4X6OJ/U8zr5SSncMKC/rv295Au1SBUQFWrre7rJj+c6t/Dbmm68Ebpg/
ET5+yzbxkwia/Hjwws03X3mAwFdkucvZuOPCr1Jw6N2B4gvNyiKMl5ZhqfWm+yf8ZmvHcrnduCQY
EOfz0RAr5REmd8Tr0USFcM2bJsOi0xZQ6ayN450F93i2rXh3YbtXIZEZsJcrz8ou4w+cs5RBZr2h
QBJGZcy1gnqWJKo5DgZcuEdC0PTQYQlsOsPtedi8IHRlZryLRAD2GxvgOUXdpagAJGZ3akVu4Phf
kHALgL1Kbz1ku79BBJfh14QzTwM89UYdJ9ZHbv+lXZyrUnsJdxyUhvviuWmZTirbY/xG7tzwej8A
MsBeolwPgUUBUc1EQ8urssDzktWQqdI4AewuNa54oJsrCW0UsxJNV0+sAwKWQG4//45VNZ/wYeEA
4rKzQZtzWNu3mcJoogSrlwZJf58V6XK4zv+OFH+w5JaYIhJCak5j+UL4O/dD4wOeqbTW2s6NSiIF
w+Ai/kqc+Uw2niZWagqzvCO6Qr0+8D/AqHJFXU3uKBv3yfj8v3Mcm7ajscRJWkIW3IjnxdNxkuQM
N7wXo5gBeWcXfV1D91ns5AeALBgjK8YJrtCGJZ0FpZp9m7Cfk+DQ0AihpvSGbTaBU5JZbXwudZ9r
HIQMgJGXEDFWC2mP+CoPkuAUyrCBL1Sc4SK77OCvTZNQgvTLGpFrBJ36UWYeybUEEv4Pjh5UjvGV
nqjU5S941FKaAy03ecj4b1E9CKe8tS6Ac511yXR8njyyGfkgXvcBMgCFX9V16WPWvKpe1aBrdyFG
3jmXdwLdLp2s5kpBuBUVTjELweDtf52d+zEJj4sIWj3pUTIZZqv3U9eHEbpqObz7ule8JL8m2b0A
5TtBrjW0ZQrFvwk/hjcDz+yAi8+akXVakPmKZH6B0Oy+mZUkuYy7B3qAXv+5vkYwgK1V8Q2jPRd4
xFK6IlVuk4VTXAeP9VPQUDe0+M6XoTFZ4cPOSIUMOTlD+2Xy+GF/oOJQ08Ndb19GkN5pKmN4QXfu
3DwDqOPy0fioh09lrQHypdHzbw6reQb2Pftu0pvbk0tinVUjdqo39/NK3350G4WCiHi+jcQw9+Ia
n9vfynlthFGLrFj+8jXP1l//rIrUG2BSWmFLnuwbw79JNebrxOH8JfYHaSj5ZYKf2+SlfCRK0vwE
v2meSbcv2+oD3pwevjn2CoxEv5eoqNWHehFTS4PjbqyV9/aGevPhBay2LEHOnJmDxplXDahLRPPL
wcXXo4Deys1MAIBemZKbl+Q5YBW2s+kATvqFzbVeeXCS8SGAqPjYgGT+6wdNWE8Cu5vo5fKAyRfR
62msXphd6RRAvalwXcgLF8OtTNLVDzPUNb66hwFt7f+Ymjqpf589kX5mkvpWa6vKx1vTKj6q2mHB
lZ2l7mutCGv1HgJYRh14Dm0cxbAGTZvfRWoAhKzEtP3PNchYJDUIrfT3iIjXfftC1zorgUpT/4N5
05Z5DwwcB0Q+7E6RUdrTKnEUYA3DnQur3O4/Rbni5EHXaaq+z6bMSUu0jtq7emhKb7aHZcHsZ8+t
9DaqzgCgbyGyiZhn4J+xXlbXSTJ0G7S9oa5YQBzS9wqoxJ1ANaLtY3FExwBeF6zN0wxNbp3l4Au+
YQFg2ysfv/SVIizvslr8RTUffkWpxA5MEPLOa61FqcOCNc+BcMxoXm396PoPcgWYlEN9P9RtQWNa
ecBc1PwDmtvHIqbzKlu3VYpKnXJ9Mm+CQ6toXcCSiU2UrDw3UD/dPFXQYEA8wqIBFdgW2vz/UaoX
dvoO0Pyhi/5YH6eOUzM0tbB61504vtPAwkxv1nkOFJ7T8qqck9H1TT9Id0WoTLwQHUFZo8VoD4Fp
o8UFYsY8D7Wo0AL/zCM06yqgGSp8ucbatEKE1dSSA0UZaoEzeP7RegZEm2Bv16L4jrUoDPWOZKWz
SujkjxHU71/4R/et4Jh2bTKKqhDfjytMPskV9irp+wLJunboLa+pyAa3loK86z5bvdqMrh/Z0KFH
cQj6DkOT98pWXEQQZAw1rsrbQir2MEc2W3gZdpBIeIxReyRDqlthYzbdJYE10oKZBYGUN2wfjcoq
fzf02EoZ5IHgtoORbmRltFi2o5mJoR6QmIEYQ09ghdzWeRumc/6Ro7pjLp3AJXiHb54EB8/yG7yH
l1HN0xbOzN7sc29gPEXfR8QZnSdTP8lWey90sA8f80McWu7cdS0z7ByloycjpwcXnS5dArDzuVZh
61qet4Ka6J2t6xJMdF//fU10QxVfgvO0r/JCbJzVxhrWHIffiAqJjJyszKDYCgfGnezz//oz+eLr
etXAuAee4Bf+/d4aCILqkLgMsWVdDfu3YIcSwAoswg8xRh0fS69D9C7g72ihSquk5bjS4dF8uEQf
qvyJg0hpSr92fy+Yl5SiObLcUFRd41Hti2YkKDOck0HLScBPUIiu9TY08E8cW8/4MJtT9+oSdaVC
SrF9uJ95bchwrUUAJ47ZrmtR2kAHZP1X/uAtzkPSdxCj4AQoaj1ijPR9LH7gDLbSbWWm/KDg3mAA
UGe6nqcZJMcjGBCtGGD47NZ+eFkATiVb+dQ/+GdiPotjP76oK2Iu0nmRat1bYtm2jF+iCZq1Wnbb
FJ++vhxTaO1ecEOcrtH3UAgZK9CcyM3nlFUjn39jUYv7tScwMPZjL51VCB32vM+zyqKJy5jyAoiA
hGocyY3DS6DuiXCorA+u/ENvfLDzXSSOnEuyw5RmtBrHufm5zReOhRdI/6IOI5y68UQIF9sI9YdZ
RJzyZWutYjj8NsYDrAqY/Ak3YjmZMByLMqbidsjbQaxfMeBbpi1m0Uw3DOGHrIyUKLESuHNz7KX2
7oK2sTGgovSvODFp81SLychuO3orduKGZDuVysA+F+l5BfKJ1Xup6BRT43LoY+6vP/cPRLrLX3LX
63V8qDLCeCuMsMyKj2l8h6oHLlSZ/uynX2uwHjCsSnWfiet6FGImbvmixaxVOiV0WSz7nAET/U7v
HurUBPIC024ITYKft8zXX+7rJ6Q5RsztiDYH3V+IrbMHoDNHQD3YQN/Ur4FlePLApHSaJvj6/HvX
Gpod2/0UEb17usBPogphwjwtHs9bt7Q8djjIgLd5qLFCZFnlGvVeP9aieXpdJox3vCdlOPkhB0lV
uDFIC/2ePZpwu0SjNBaUT5uE/Hw2ppLZVYn72+RaggbtWAujwMeUmNlITH0PdVI5+DrO2ALyCELu
o30bS98NJ+I74/VufI6gMXwD5BrMm71ckd5f1JKue7nc0s4mrNeYTVq3CUQK4IyQ6ET3/0QjhzJX
GY7ofIGQN2UwgHWXozGrkkTCygyiYXoc8ywxoTbbDTrlwYKcDVatxUpcyBFUMYyQTH6o9OyEOYbd
6/2c2JegZqlBVzJ992dbbKX3xnlYI718GrJgPKkqnJO+ZYxrRr8jtlWtX7Ku/Vy7+3NqXb1Qem5g
XLMIVscJ1RFmqaMp71N+It93wLRuBqTXZM1iv0EQJv2DUsUgrfhtxm0N3M2ug0fwjqdiBGNiCri5
zPs6A1u4bIU4LU9iCPPegtGiJAThd3jJ+/oD81x/1BN/FO2pehxQLjqb3mbMpjFIioPWC9v3VHpp
d2+qYNPDnyoc9vwVr3P6SzWwajdvDWFxV90DKWkTDbHP3wqbBo1Nb9iWyrV1fhoo3VoMPaIe+Qsk
P7Q7nm8CBxglrC++d9WrFngjVU+N4RUAtXsXbPlTYzjTBdJSxfA4rnXO+E8xFFoIf/DgdbE0RQKi
PKOPXaLAZ4CmPylh7UWC4Wuo/P08jcoNBNY976y3fD9OZ6via/w0RuyRy3DK1QnWmclI5trH5ZO1
elJ5WKsa9YVbyRdpKp5SQtxF7I6fuTJVQyMVC32kXXzhNf0bjO7cxtRzy5Ee1sVZwY454RnZGWaM
KkDODdYrWMybJWqivsG6XnDQsbr0m/l31MwVic2thPMScN5l+F81IwHZZEJH2AnEs7XbqHRgQQ07
FMhnBd+BX51qDFTpmR+l7OMEP6EsukL/G4X9r2eETUqDuHlfUWE/wAoNmYT+WvU5HQkjknWJI6XV
ibGicrajfNMyokEnSbfbiz/CElvAGsR/x+aCI+3jymzCM1W2zANFGaJFzl9xHRfAhO+0REl2CNFa
v7iCUoMKDT3CWj5utYZVLilSo69SwgYSSPogUVJRQtLREnymlScEROEOw7yIqlgvy+b9wt73vbwI
Vs0r+WQNpyIHMiOo9NY8ZFAce80ih+9DKcNzvABKU48/zd5pQljL6JFiL8cHO7khpgeD8fA/w5Ls
9aSas6ob1Ox45Ep4/s5JZGUokwososIMBTog72RrjzCt7PCNUXhm4ouT0wN6wML0hRHnNMoDBJhC
cFPaaTelwkRhdLuszvwYP2mUzZMMSpsPu1sChCa5kdYGElm74REHqb5ldPxi9mFAL+K4UTIc3d8n
8J5clI4knTjXwepeZdSc7UsWw4FK/bqFNpG07SgIDoajG19MyJ68S8+afwAtweNug4SjbvfM8Gx2
u39esSQJh1pQKF9bCQql6swe10kbgm/v3YcpZG844Zd3RjvdzXK8AaCFD9/qof9GyzCDFBm3ZqJm
Atbj5u6tHSkoz159XDMUgJA2JrkdBuIATRZIBGMikhJ9COXc37Bjl3TaCLzRzyaZDbEZOOAMBnCj
PbcteOURDiXqb1tdBgKFXldrbfrLY1KX54wNk90/KFOrN+C0goqUAflfptoEiZdfBAuwAJbAgy1v
PKGaOPnF5BTINNFeF/ze3snLI+bb1X9QvX0ntjjhRAd36RoqNbbLAz0ww95XMcJL3DjT9Ux4PVOI
zbYGxAfEM4CnrdPcsda0s4rsURrd3by+kmG8vorYoYHXPbZcWG6/iVhCxgF6y2eoIbLIjGHjTzHJ
ZtmZJUMG2ThgfOker1nnVnmuVOrrmJH00kLUcL6MA17mC5n2QAAWsQOTSI/yGNDjpwNMGhbngl2w
MqPcnWzKAKpvcXqMabdnAKilUOMyrM5bOauiArvy3qv+lg3nGSKBBg3pGFD0RKJC84n8/nkncI9w
XtUkW2Yn/txwrw1Xs9TG4fZ6IQywBmLrN9wDXh6MVv1JTOTKkXXa91sHbA+CdWvTd6eV36QMJpm7
vPHYHxrewdORcTmAtI723/Htppjbqe9lPxXcdY1NByT584nPV7Niow2AGhKZIv5vdkgsa0iy4ik9
n1n0TbNP1DyRZhHIXzcfAN+Mm1yv6Ooql5wV1Xa+46pNLH1EcP4BwWn7HXRB7VPUhE24H1QNwNcQ
zQGgZ3CaUBkbYck5jlrvBnCoMEf07QMu8dddS2/Irm7okizoOO4TZ0UCLfMCo3yF6x7julZlDiHT
egoYE1ZI7T4NFNE7Cg6TlI+PFoFGFXAmEcZWBaGLSaQ4mTRpGQyf0HGJAVRvXAOq6E2Tm4grtbaj
hNUUr/XO+bREtjz7I7pqeAi/J7s3ReUce2vUNqNx0r9c6gxCyncuPA2veOJGGDdpPb0EyCRuhqab
gmwuHrRDeoCF173nzKOtc44pIkEvS+hojCaX3O5LXF6QeMfbHcVLBPrUotLMOfGfdKp12UPdcDs7
pbuBngUyDuHmr1Oun32CDKe3TRi504CQdOHdzu5W8QBYQZBJoRoflaLuMSpOl8RuKG64SBNtbN+1
awZdxqcO1Jn10UOtsfoCln0Z20F1HUOXyLRweaDpEui1lZo8es4QlSd7xIyqToGozfwpTO5QAK/t
j/qxOkyMGgCt0IDm6foaMSfE7/eZ95EiXFurYw6/O+gFvINx86KPSFuIuMpjPkzIHNw5E+P3jvfr
TMhgO09j207zErS+bpoj2QGAm8IxGfCOp+vOANn60SQ5WJDZwej0Yxe0ZSkEsSEZE3bMWEYK/ufw
+BlnhMvdeHPOl7jnaBoIzQsKQIl/4yJJnpWAHcsekoBquAEZknyfspUnnWHYl6mamSzV9Y9vMBUU
/L95sa1Rkn+V4khDKu3bCxr87VtzZz8F6KN++yOhrfIPk8XIZge7djySx3u1ojU4bmyDvJnIXppm
VBMuEU4oOOEwn62lzbI+XDkdKI0TX6UQYZz9LcErJIbwgmPHZIftfzvGiCa9f4hQg8nCIk2Brg7U
izPeEZVH3HBwhsPlmo0Mx3qYsL10SFtTNCIq15V5mHXq5zwhZmDcpdw5RSjVsAAbkNapcg38vJbj
Qk6LY4/tfkPwwPO19iqz8UPX3AJUXkrzIl2CQPPFTtRyNgRMLDx5GKsTPZpVsIo1Em+jHOe7VuUZ
TK6ZaHIkhDug7AR0bbmDtbzhkgjZX0KQbTxENWVwX3jO33AF7VPRNwbRokDIUBO6bN4866lqRu20
ifFLqOSg/vmplUnoTpOzWIl0N6qlOKTaQ8ygkBWvdxz7pXpifQI98T1dkLl+MmUS+Z7f5Bk4kTED
dPbgotb7Gs+HYZ/dJogzP7I73RWd/DYzdSNxRdrpzYUVmxjWxenjSA/frg4yjJjJA7dqtFX1Zr7n
k/xsPI3M9AO01rEYB+t3YWvFF8w0CvTZ+EJLkYxGacX/yCGm3Evfg4MVgWzqbBx2gOt1Jipx6Gki
kpvBf/ZNA0pHML2QfZTlMVE1epqpbTb4SR4gxfoyGKGWMj+l9F4eM6bOTJMSXI6AKMHFZ470HbWp
0wtBxP0X2GRjwu426N9S3ewWhc7RQAOlKXMWwze6oix97LkazJkZ20YtZR8g7/ionQvbGSjslSc1
9XoZt8PxsMTPukyJRz4DvGFeAeiNU6KewPsJd5XXz3NH/bAUwryqd3vL06fUPO/RLlwq39Tn6aOO
yqcIId1W3shiOfZEt4YqsGTCZt577EOklMAFgoPGJaUaZXvaW3E488RN6153w1g1VsKrKgIy8PGR
4DDz34XkxWUW7DLh5kMtCHOBFEcUvBSA+WQbE0SIVud5pIx3Qx55imf/k15i8Kq+RFZFGQIPEq42
A4VhWneFxPi+P9ZHxxglh87ho/GU+MYQOgOhYSI3sRLAwqmJB78y3LlDjK3vHdiMuqY1JtnNbDpm
UtMbLjf3UFoUUYZx7V779nA+26S1AxEEzIlXdCYHl/ZgfhVmXTfxAtJh6mE43l+gFwGXd/q5D7wb
0tcqIDRqK/1qzFuQPFR2BzyjBRjNv5BFmM/9+JQmPxASOr8SgC7SJrzugb3w20orcI/FD4f2qTvL
ksYdDUeC/SalQOPXQuX/RBza1dCXueEF0DkmASYuAz8yKnCAri22B0wHptgK36tYc6Oh08lA2lU5
qAWUdd+z2rHW7sCc/CsNy2djVc7I980vwE6BrMo+gKvMguAfbnj3nHKcVys1yBV4bY7Ua7DWrfr8
eYL9QCD2beAgsSPHWAK/BBXacKEUa91N3yBYZ66k/Gyo3gHypg/P0i1rq8niCinKUa4H1H51vBlZ
LDlTo7nSI7UKTbVY6TkBN5Dig0/6RAMV2aYXOo7dACkm3gztMOHEEhOwkAD3JnEgKC6QUpYNCxNS
o2TDpwHQCvphWZPbM07XKpaRVCLxWQn5GKF3st7n3nMrMYotHnGlHBtzKC17PrNXg9SCJhO7GaHJ
/ci/TzDlP1NyisVAIpLCRj/Ug8sSCY41w0ec5kaA0dvsNfwbznpjzRz3MTTD7bSTv+fbugGkqVmk
0PLmyELUFoiPZaU0pQvj6XQ/OP++Vz9Kra8/ubjr2hSB7P/g+1e4l+nV3+QYxPmwlMXHlaOexiZs
wpapiD1SpaMC+05ftlepTgRzUiL6ZH3fLnrhwgxdd9daFOiCqS6qcCmKX/Gdc1JBY8L8ixD5nLn3
aI1fggElzW/1858OAI8grsQT2Nlf0IGaej5eidtLSvL+nRMo12AwBR8vNVDum7JF0fvNO+Pg0V8+
G8qz07wNFX7E5xXz/W/xOhtPvGmJ/OD8xEBGNQ9vcsZU8uWwf2afg1XpNlaaLG/RAxwGrkDGUjYn
mtZ1x/md7ZJBwPVnDAC1scSzztemm8FYerAGhL1e5ho+3oJHVvaZqG3KHJUcn6upqahEblnfxT2V
C9aq10ygXGIRj8YoRmXccfk4nHinPpVKWEm1igZJBP+vk9uGyCHMfNzGVpMczh1SLVZ8rlrgrg9H
K+/53YPbKnzBBgp9B4uNaT3rkPkO7kxE9tb9CjUgDQ53jvurJOxyIGBFnNsLkhXBQZ8qXvk1iJT4
xq/7zO/8hUo7hkbz4a0ehqIIULl2+mocawKR1THwbSmY2jnZ/OgSxgLNsqqoKA5bUhzszZ3iuUlU
JzVIHUq8MHgkegepOAHFuZzacsZzM78H5tQpBaUmkL7QPhltRZU8ar2RNpRvgqHxIMUXzo5BdOwT
jyZ6YW+yVJjDU38emv/wLyKFDoT1A/f3y+qQXVzcJCb/F8u0kSKw2YV49rKL7zsjaIKeomfSOdlG
A7zi/TPMLR7vwLx3e6/nGGq/3fBXEAMiU05hix4kPDhBDm7iA3icKM0BSPM6NmAh/pcRTZQBc1I9
HRHllA1oDihQmQF60pOxNgEcT4tkwwhTVxmuMxXkD7zs0hJE+cB92Dg6tfv+HMiR5xVjI2lgFtKI
Vsl5v/ddOumGLLTDBzPa/ZB1NFQ5k4c+9qiNzGQ2mKXN+Hq1srrLP2zY/sU1sem+uDB20wmFvmt4
m47cRKGc8nGOGUmie0auAFN5EtQPJn1g3H+npsv3Olrxdy3yywVN59Cn4TeeDs0vEivN/JdDNU72
AGFQIH/zjZyqLENH7gqej0hFC0Ur+UhR/7gp2zwjp2+rCMK8Y1kkFjATsCJDJbAndQ4NRHbRqVCX
P5MYk3lndwaDh2kMGJlmQWERyIGeVaIJZJIybgNOEva/JaqjJtRMkwpDHWU1cHol44OQcngYxl1T
DSeQ+A4VuAu7pAT9j2Bl7buJ7eViXrL2bTqTB9UQPk+7bR1Yl+PYFwVS8zEmA17qU+nD7WXLf/s+
ql8uplIkNxYa1TxvU9q2Sncvpig7lRf02JNLgcSkXoMSKg6bqUyXyzajCTpXoXJiLTZ2T3Pmlx+j
iR6bcBTOvxj/g4aHMW9E59vlY/HTF98s+Fi3bGaiVvf4MTuRd+AqBwrZOlndRGv5jcFhXyOBRRRB
wlvDtf4flGJRy1AWEwZ4ayLMc9NBhcjKOy3iSVTJ4XoqL2NGm4YfyKJRO5PGwrTTQ0DgR4PcPXe7
zYJpWUH9lDBRhNR/levG2+rF+RIUIHmUOTuHDISK5Bm7om4ICvWe1Q4K8irqJtRf13OLHV/gpVX9
t417nDZ+FkezldDJUyn4KCf7+Ugo877hAtHbzXmE1Rsv2mKDkmH+YR2Yuxg9bL78NIaYcoh628vw
lt32djrwCPBBjlWxmVnnt9UZ93V5HyXavbVC2QpvNEe1Gt+s2kabXZiyPXTUBHtaal5EoHbKhbDi
Dz/JGxtQyssCD9Lk2q9cPq+paduyPXwmk7SEjc/Ydkz+8bknjIVQuwlOXCppZfyDT/+80425/JXI
7Jk3OXVL9oaGGTXc2AfYFQf2vAQWFxyPpuHleyc9HHSjMOlKrmyWb3a4Yj1Tl1NV4t+DMgI08iZi
3lq8YfrauYCIzMvd8Hz3TdxzGqCjR7q/VFK/UjeIj6pyQc2Wv2lpVc0THmLQCIDqBDXytnfwaYa9
ToY497LewC7YF938AkXa/2bvGx+FuBRIDgsKYZZLMfuMdZGu0pLIn0nZBpjkfdQPFaAxl3f/z+wb
OJ4kwFGsTpWaDtGRCdX7eNeMhrGW5PDpEhOjCm0D9QhUjK2rRSo97BkmgjfJfuXvxSzgwgKLzxa2
NyOWow+L0RxF7Mvlc5KfuUYViYE7rIJ+zVXfeO4DiK43OCaGPLLWbrUDPbTpdbtotHTJb4SPE7sW
5fl5XcMM/ysZr7W/LJW3UN5jWKWKVx3YQoCDbZxTYDGJHXrcKHVUFwSejQlMjgMXdY10ANL9NJ6B
KR83RXmiqxB9r8uEF039vNJNU3KcS0JCtsx/Hdc6J3NS6fLxQWU1FjQvruwg9R1zk4zwSkoICBf4
n/8L86MBhvcapaXbzWDrIv8UfM2e4jtP/oST74meJukrb6OG/t1hf72iZpcpBCqcNN8NOPPjWFkm
JbgXhAXeDSLve8RtIH84TY7D6zXH0pEjMEArEs9bxdYCL5BpWurEaYmPGFpLu14niLgU/+vBZ++2
uIvdRgAcLQpgP8TeCw2VgKHqCmoPxnYkbEtDCvgND+5bb19HRt9S8fu0p+Yg2/EPzYea5Xum6ODI
yWZYy2f8jffJ73lBCGutMbYaAfIp86o3Xui6NlBOKHjtY7EH8OUT/Za/Xo540SM3SwUd2lHV/GVd
kU3BwJ+LCyKaM9x3EUgrG+PMnvsSt+HCO5wjCS67PHHJAciGQsUWRApl2KtmeCpK45E1POYGLbI/
QuuTz8iEVPB/zUQekxs4u02GRMxlsAGyXMb1LDF5OGi6KQAXGKh5TB0+H711Ks0CLBaUhIQHH6Ux
q5vANXYzL3A7A2iDAeIUsIPmDSxZc14uOfXBW8Ko8a0L1DQOfGQoqv+3ZBIjYFh2DfbOL+jT6R7f
UCamy9fnr/gaJ6KFmAXte8AjzMclyrUx3F3yov6GicOWDuFynnhLGwyZQcqk8sp3W0Dbe/wH8d6a
QNV4iWxjEVoyTTpNyPXe0rGBWee1+lyWV3ilx6Cr4S1qu5Vt1X51SMofaCyUroLa6GxzHbuAoBGL
BmqwPMczRU9zCjsZulie7Ky+AJ8cloToMASbdVujdWp+xVldYfBcLCRoKyJnC2noGFnpTMerz6Up
az+ihfemEnvG+rSWW+RttSEBsJQe7fTgb+HaFcxxmirabUxgoqRKVnJLjbCTsZNcqmLten+UkLSL
5Ji8++NDXlIjWbSDqQlZQY9VVLzCn+ex9tcdx25aVtTh6VK4eEr8GY916Ry9oHkiGLhJ5qnph0q7
QPfCNr0Jl1z60uRKtFmDJ97w+xs8lrXP4jf7ziUOJP9v7whI1LmvKIc35IConFZ12HcEdm1NPjsM
8tO7+eoYfqtyTGwiEcIWyCc+Ysrt1r9KQbl8HCfHeR/aoT+fz7MYZOkkTefKwqA+ulBo/P6sUTV5
psYsWp3XIdSdPKS87VFfI+EoBUOsIz+0DjBmCpHs72VCDCoejbXmUTQAxjLO/T8pFq/yjUd15HJr
bGeunION7zlJl7BE9Xxffb0wm/g5h65YMSx+5i2LYCqQZX5jEaMU24X0Vvt2VFphwShW4W0HIVTN
oaqFGKYEjdcb7lKhg5AuetiuEepidqjSTSgZYiXs9LTp0ElY2uZEL2OdDN9taamJ5M905ViIerWe
049aYU+bGk6Ly9jtgb3RTLpIHl2J8tzRLTEQdqNQNgwztj7CRIMdJVqOayvoBMpOJOF/Fs/McmHF
+LI6qSO7neEeXEihC//cIdW3P0x7mCgOrhjLo7PO5p4BCF9pkVjtH1XQZ/3AAuOAjc21XLBIx9Px
KBhmpNo6H55Olkf+YUi1/O7lqeEfIpCdq2n+AKEb+zW4LNl0yHJV1RCgCVCXembgom9T37tGpnbI
JIGls1Y00BLFO5fP8rIB1R2yRJJ1QAf6b60eURF7x7NQYunqOeFmGecM5xJr9RCHLAY2hQg/fv9G
fBlNOg5mg3Bgge0iWSgLEiAOH/z/1SMd9VObcXUEXHE0aien6+WwY/TiiISDUxkcVVqISwX3qhH1
nmgcv4Vf5NWG036dnmRfTe+tETBe/o8F3Zlz/2tqU7z4ca9SAxltVDTQfHNtPrVK+hMf+uDu72lh
j0aDJYvzcja91UmJLv49U/pns6qf2YBPOs1Fa/7psNXk32F4U5pZ4zFmzmyjlK9eWvjEzALNKncU
d5kr/jxQ7cgISdeRI8hgKrigo6VfqMEn2bqGjlwbuAAXau8IIrqA243gqFHfKHCUdsrXF0jpURuz
Ae3jd6BzgbwU12FO1HOPFbx1+FatQfueP97b0oKFf5nvYzPFtE1b5Gnvoy4Hb6kKhbUpjLMmtPR4
KKXdjHmL6FPMrHhUfeR9d1p1drutVCA6/PfZEOubQ4swEYxA1uw0thfp1MtTmXKUSiFQNCk/y/xb
C4+XRhSiKIJX2vk0OPWCdLM4wpiVtqU65GODDGoDHHasNvmIOJJyq0J+qHARY9CpwEe+UB5grhGM
HU+fjpzb4fSdJdmn3PvbXTFZPhNN90PZHQqnHgwfwUvOWCTMA+3GFyab4C4TEmUURk5rXS6CWl3f
jGWFy/byM9Y9twsgZgKMgYkIKAINp4Y2mYLTLiqpDQEiiLmjvl0jS7mMW9S58PGZsnFwkPnr6G7+
B9e8prst0GcajMMBrWEPlrd4PHnVuTnpDF0bbzqWYsDz65e9MA/6xXIbRnnjX0JC8FsJvr2A2jGX
bLVKUb8bjNstfA5tnzHr7XXxVKnGbsel/U2siV1EwHFefSV1h/wXuJInunXnA/OqDDBZdjVIOqv5
xpAtegJaLBBePoZ+Ki2zS86lIqF5WuJzMGlrhfkv5C6JPem9iJ5Orj7/C13LPcApBcFnW1maXYLJ
9dCow5NjvTCgUaYe/upL6r4sIEviK6DmsOkpuzAMLoPNfz2giNODN91M27jqg5O4SGrZYUgGbibt
bPkanOjHt0ziEUGMPWhC9cS7FD+szXSZwZTcu7Z6OvLNauXCuFqawEWRrTs2wq2hGQgh85NB6qpl
ge2NTPrahTUbNxXVX/YohVSa92sYYYJtCLAzw8SMlui8ZjJrgv6Zg9jsHZva40HNV6ZQM9VlBKnn
U3GHN2PQc01wlEBqpwu3zOrHgAjVp0OSQhIMMtHvY6AVMTKQZhGwAFlUWG6KNrsh8VokAoL3ijZZ
bsPFjzGVN9EdS1TC9y0uTS9R98Y746YZAUTjG/22LGpAQ/ByRZJa5/8rTHAD4+8qCbjFjHg3t91D
g5dsBecgXhqSCvgsqz5YT8/4HPqcd6BcYNXRVeyLD6P3FGYWKb85lIdD8MriUU5219X8ewbqhYFY
dTsCHgykWWq39s1TNQd996dnNhXdHPLk+IPuQ0Nng8SoLBomOFJg9ucp0Hml7mV7EN/9QtVudUFb
su2RfiDhnvcfOqKxuqAL7aFo5DKNn3p8oAgnr0nIalaWoBaOylpaUR60bO4lorv9z+02BqOGhIox
r4U8Pu9P5PBk0CmytvqrU0x/IYNQlc74dYH2NDjbK7MG98olNfdl7x+1HIt1SONH3IwVHai4IvD4
cRazXulePn5NZk7opqCzEazkYWUWZrAHk/vyk4kT+6UEqiUhbhiqc1rMT7AMGWswEYtdDHP7d1+c
UVp5QVLh/BhFxpRwiy/wC5R1jeQKaUzm5AUW2MifZhtObW+8VcO8iMrY7AoqaugrGXInG+cMED9Y
uGP/WWdsdO1CVJuMynBbbE+e8Xl51kvLm0udr6g9ZWYpGaJ6nS683qZpJXD4xwgXybLtn93Qcyep
270zTZLb6uazDx3fokGJH8wkp7xVki3eEaMEG+v9cfOtZWXSzk4eJ8S8HojV91Rk2Tph8D44IqzV
Twr1+TMcQeoHMWGzlyV6Ls7Tz5lMNS8GkUK87w6lVRS/WebRDSbs4oL7OXl41BfFJhezqc4iDORC
fHyjgGNdqvpI2ik0ppgVIZ8/0HZXXxujQhk2vGZKhMRLQTKCuGWzduE5Oced3+opRPkQoFbSxDpC
I7solhsvLhzVUVawfqOC0Y/ctEVg1HPh9Wwj6vPX+yh/DnnOxrN0pWHGubXjpyEflrZi1MXhZ68z
6Rl23pD3dWgTXPYqBkakOwhsNJYgLqMudok2ayT+fd+bmJx03ThtMGYZrqWEFqQzXBhZm/Zt+IbE
FNBu9iGGkcMQ3ppZqWkq2SrYAuwc0n9dI3iHBuxXsuCzwaJGo4z/3QEmHPI6GFaF1A40ojUUVjVo
3oUcatBBy49xRab6I4iqfbcGT3a3aKC4Rz2LVf0Jh5FjBVkMZZftkWXD94WLljIuEEhFEsN0G/kV
fVUu6wmkIraACpeSxa5/MbAEYJ/kaKMeeotb0jtKJWvgmfp8sIe5N4bEu7Z0AnoxT3CjTCGrVLtO
g4weOF8H/KKnn/kJt9fdcUGrt9Su/W53+wgfs6KTFmemAVLq00P6kAvNBVeJd824fBBNSaQLimC8
nk/HMNL17MdIi4hG2aAWrwWuW37P/oxglOJ9l2Av9rWnYorHh6HIp+VbQdbTg+TgHn3Gex8zpkq/
JvQh5gHqPiLybR4EGS/EftxDq9u8ru0A+CqV8e10Y27koPN/r/lxTH5UAo9l+7Jl/0/c8s1aTj3i
4aOOAu9SDUNT9I4G+QdMkN7UMKWryrZg1OWq6jDGDBootg7KiwrR1FhP7WL5XDLr6FOpirx+2bFT
8m2DjrTohm8g/akE2s9DdrItpHggD+vksde7kreXWIb86GWrFikYiS81mNQOZQpvPz8zUC/8sWMd
3gFFg4TA2XEhvhdaHnjaH7YvHqjUrTkt+w6w4OzPuXuoZew6c31O5+wLMRixrlvhq+1lDKVUWKzX
lKfu1Wv02bWWuUqeBQ3Bc5I7LJEJQ7yNLv6NOW8GrGruqjFOCazzSZPgn6F9KUqiVdKqbcPBDW16
blRctc/NgOcEd2IZWVM7HeG9m9YR3GaJv6fbcZxz38zdbZDsm5fQn7OSWA8x/EJ/fkGDk5kPeznj
2LC14ULSmEBfSxEoSg9lDv0+5h8GqcRx1i9xoKvjv1DcnZMwU5Nk+aZTxFFFZ/ZpjdcfTwoy1MmT
tV6SDmyArcgh/AhKhBAUfhH8SGYeu4FOxU2w576VcNZnROivRTnwGc9aqKmDhjkCDs+62IQ/lzUL
W/jox3NmohQjdH1Aq9iAn0GCy12Gz1aIuGsimxS0SVncMJkvE1iAp3Mka/zPJyi4u0IrChKrn7Lu
mNy+y2ldewjZArDa3miYKnMXWM557YK+u4ZbW+N/PBIsOxJTtGcPmFZBrjCf/dcsQefyiwRXIWIn
v2Q8sR45PRKHBqvTzT2mAkSnYTrAIEZnmo2pevLnB1469GaZKkvbZdGgFlRuAAa3FbJN3Co97qsj
xw1/uiGD0U3WaSnou3yGUhnNL58mjsW4LRe/i4ClM02FCSnncaAD0naD0PKDvBRkRsw4MyGBBj+c
Zve0DsF0Vvhzi2PWXwBh8LgiFyNurcwJs4jA1Y4FCX1EcB5AjVs5Cpc1vCQq7R71fn5BosJZp4tc
DQXNtjfWcHR7V/HwCu6CQ7pft+tfOLHTK++2PskcxlNcqDDuS44W4OCyh9Mb8FwDpnFm0EDGd3Vz
xvR7vCv3Io56QuaZEeDXQwk4L66HtUpW6HOfbiw9iNH4vw9SGKxXmEYu7tyWotiVkVTp3A1h0T5k
Pf0MRI055isOtCr8vJAHNXshALM9D1wDsXkU3bN+2m26csc9ya9Bl7UE7ZdbNJZsc90TTSqSMW7f
0xR52E79eThIz/VfkJkIea4axoJIaZT0HyMrjRkPMZ9Zw99oNFppZJ0ZBc2WU4BfocJ+bgynHCzz
53TQxSh8oA+vx4z6BfGinB3v2gtCvFXT6FnJyhWYYbw/y0I9Jd1C+nf79+lY6CtGFIslZhso9Cj9
OIynwPtLy3gp9fTxH/yGXQTS9ULi3gnINLKMt7KqJyr8QEJM5Dl+juNRZVYNJIZDzUKkAJlzz6zQ
aMTtahe0GLn5Tm2H23kgC/MZZZOk7C1qSR6tuVbuWDNfKh/e2w00SegRDGW8q6OibwMKhNPJqch0
GZIuV/fqt5u52BcRHYEFoy8qhR02YpC+b5lfJTW9sismghsQIxUYRu31r+cwtr3AMI14U51d/SNR
6la++HPrG4obZl9vNxQcsCF4KV5YvMPCqVFt/UqBDtIa/uH3kEvYe7Px30zh4bPOCKLXaldB5Td3
h5651IEHGlpz9o+ji5pfUljgWv77CFai+0m9W2ISMdlBB2FnqnhqUMiELJfkCJATBSYv3h7oHKc2
2H/0h3pllVU4FWaUybV2d/GFap7dULSJT8iL2JmW08Od0G+h/qmRnX5Tnm/n3dYyprfz+bPg2h51
dLFQw+uOeVvP2AhRKzb0Bi7BigE9KUTTyjkOr7pU1nvY7E6XnKdgxIU5ywO7y6nneOXtTi44jKLT
pHT1I4wU1z3QKWn/ubRA0ezfFxMVLKjVsXdaTK2gEUXdiG8JUKg/avhQX6/5dpDQ61n6Dux41+CX
HaTUC7cVz3qhUdTjVY83FSytQflVknPnSboTXRC2KwMai0legY/igke5TtJn0tNrcng7/CpKO4X3
tLD6Nfoyj50bapu92Y2vreX/MapO/yiXYUle2Z8fI+vy6vQa7YSTqO0v4fmZZmhjh2sep8qCxiys
orn++A5QyloMeurjJpazzY8er/voCPwQFcUTdJvubtGTE+LlgAIDXhAUKproMB6KXqa2j8466Tpp
Wcjl4VVurEIUAIJpQhF/1OFBkqMo5zwDNxgQOvzhUqb0nxngcu42m82eLCs1l4pk5s383LAehTcj
fsiDh9BSFedCl+H8wQdChbG8pK7nCF1tM9NKgw7WdWS8hlZWtqB3WqlPiTq7axYe1biL45649bbl
bNSfxwVPDyNjvjH9OHSyx5y9luqhSEU71fqdpyaJYgj2RD3+enSf8JPiFm9Zvk94d2LsCL91CpAP
fvh30DlBHkwC5UbQvJJW+fpeIRv9b78BN4liBwbzygDhLx2YE1PvcD/ZiHl5TawpcehiSqZD68Og
wQ5HSOq9JqH96TuXKLpSx4W23ThC6UYnZLLa8jTFnUMxjI0dJInF6X+/XsmQZeiOInB+3SobWaH3
TAS88myyizq6csC2RV8DkVkSlhV/YcbLrLKUizgYCUuzJrmQPyE2aKuxaa/KsceN/7HM+EgFs4Y8
EJOgXwnNqMSrn53dN8ORTwwXQQcjI+ZSfWaHBFkR5ms0hEINjUxSc6UcnVWl8hirjDufe19RFQUb
G70FGi7bl00WYyX6muTQ0o9xrSpQ3+/BAgggp9V2sNT+PH+Hu3gkhIqQB4ojdRH1amCXtTV1lrk8
P/2/OxbGWqJQ/5P5Dw2Zas7lzAWe+k5ryfMJP4UjHMFcu+WIGtIAUa0Pl+EX9f95N1S5kl+Fyf1X
w7tOEzoa9mmWveBsRvaOwBTISvYz1bRgL7IRgqAS2DAPFKL+1VM2edOBmUIYgM4JeuqKpcu2jKAM
inFSDTPxdczJNBpYFxxQqjpKG22xK3Qy4oR4FCaQWoSo/3lBGsm3ejC7psu1mlgH32wPuiTYVjRP
ThOdz7gHHU2G3or2W/Y/nNhT6Vk2B49tZHH/euhdrnxutu4DfFS8OVVQySkOyCsvJs+JUy8g9d6t
FGHcsfzDvbCz6R977nwbcmPU3zxPYk+8jRSIVXXSUmVDV3gaofrB9H3tSspbN208bYNUyg4/1u2H
AGiGNJSLV8eVdY/KYPVRwcEMx7SfSqglAm3N4YRUqOidMGRV29+vXjfhE4f0XPtU0r7m4kVGfyLm
9GhWL7e69VLoZBBBTlD2snuX3/LkoOCfabogd6OwIa/JawrF8PrHL6UD2OVDBF62JnLLrSRxtESw
FNusRs6+BbdtKrfDieVznPqy7iySpKsKWD+5yBQ3XAWGmn+cO3hPGVNcuyYSA+STZfrLtJJeMnmv
15lZbpXI3dgBZWX4ceQ3jOPE4Z2Y+86KwZPj/+u7c5skNuE938pB0ftXfZ4SyqxhfMjHieJpYyG7
Iji1Mm8u+tW4qfnkodOyqqR0QZfllTMWLlpNj3prUoybYtc8GdEf6YBySAGlU6aFUkQ5dyk3oIKC
HBgEEc7p6WYHO1/1AxcCYH7fYpDbGLfNfm/VlrOt8lpauTtDVqxxi/CmhjLrl97cYaB/bTPfL21F
z2DTmepZuBTvsMdj3b8T+KC2cTCpLjFAEe2dpCILhiTzQRpXmo4B2TgZHwGe23qIeLWmDyzye+4V
0tzOZXJVCaNiGm8qx8IqlmO9wJys6aFn9vhmT2LdJKMijhrQ2sd0R8/Yr+6q/FZgBb7eXYszPtSN
EyD8SGjVy4GE87C9gY86TukgMjDkp/2EhciJqVkjpkj/N7TVgbGXOGwTrb88Xcb+ewbFKwBkkCGm
tX4vPYX3t3qj4abthCbUXjrHtHKRAwM9fsGglrKgm8/flwB/tDiAU01cCy1l49LGQ0kIh6+uGYsE
KffqDVggzbwfJ+gyc9mb8B7RdDAiylmM6Sn2IVrGqFmJuwPiumSpg3GLvUD9coYZVmc7/05i4gfI
l+K3gNAdyHujkPHz2EHA8oXvlHJwpFLFvoMekwZFGnmsN/9nYn6br4kCI/7kdCOR1CX/Kfhx5+My
tVdQV2M2C5ZAgn5AkeFeCd9fwo7X1VSgS7NgMh6Q8wdG04Wlbg5ZFF82z58B8YVjsjJF1TE2bF9f
YMZ3qivhFUMX5cya0KOmlxnTK90no5lwYt5jSYZPcKJQ0p8Pp7F7eBN1xCgFMx1QOulm1bwT85DX
xAi2zIlgc4S+jpCchhDY8og/NQ4ZLbnPTeAo/7LCkvOH73RBWvQ+CXI7VdVFGIsvPZX4TkoYLi/s
/bKJk6RHwHa+JGuPzymjwYo5+lHF9W3ntTMAye8y7cJsL1DbE32xTxva6pyRhJ2eP3tE3mBMGjfu
qljp9uWTPnVsmIr5WKzSu/qrAfn7hFxoLogu2NIaCmnwi1FXcS2UV50qoDON3X478ygtEuRZaVFq
l+ithO/CTNwOVb1Qx/YUxw2IrGywyPiBMclK+mB2SG3sH7qX/n20HLJHLbIHrD7JgZXsXY/h2bIK
g9EwHqBfUiBzkRLGlc4mhl9MY1zLEGjc7XNQs/Oa+XeYQWLAtpDESPLyrBFvnWoo/toPEbWqN8FH
nBb2FAYMsYu4eWNA+dPlUyqKNAd+wgCKIdR0wlc4B1EULQvrATuEiwUKw1bx85woRQRkpTvVcVEC
xt2SI1xrHWKkaJAIrd+kbPFB+KktM/Syu0AaAxA/OTnLSegD29DSnXJBTv0jFdme26BBUvwEXIV+
3zpRSWtfjASDLM/y21+yLAE/3t9J3RsmQqYh0kqGG9cpk3jCaaj7fikG4HxAiO28C3cnCXTRHD7c
2uIlcyrow9meMGrTD+A4rzIaCclEb6J9AxA7e3LzuZYbgSpUJLX/WTF1ifmhCJ0vIwC91KYf8HEm
PJbXX8kKDFhvA/5S0HglGCsGIxJi6CrhD43YiVJnY6XI/x+g3hPbaqH9FHULc3x97dr8qNhW+b2p
xXsel3zVWKnabW40SCg+3JQmBM1nfg0kyb08DDQ8tE0HeZ6cAM2P2TTXpkynWhu7iKnzfeqHg8DZ
WQ9arXnjI0n/SbuG2MNlGDT16V6H/PN2AoRa1eBFdMAo5CLFoptQVFEWEpCsSnsdWZKnob5Zs1FD
LSKoTybFWxUNEhsbkGE3CKXlfUu3QAi+7xTGOToJvYchL8waDVz+HygiR52sM/J2WtJHoQ2NDfx9
3IMpQw/oE8ciEMVMRykzvJO+IYJDzBx7SWUWNgsTcctx+Bn5H2M6p2/PV4yBNl7GtTdoWQlxu6ID
bpeRCIYCtpOEr1JCIGA0+T+cydprzgnl002jgBo75eh4VpuGcrz5X7N+u/7gFd0ISkTPngqDO4O7
XAW+tO4kvxey0HYbk+7ofFdm89VjxiFd94SRMlPYbOnGQjxhhG5Q+rBNG2kiS3Y3poVVowFSo8Q/
qwHuv+t0NcSWYSCGn51Uka2wSVsmKF/0+lFxq1p7oWRQ/951MuKshEB6OOusl8aFzCQlR/B/9XE2
/tjYN+PYJG2GapU1UXV+lzzb+oGv+jaNwSRDha0RAR8vIedmu6JXgalR3fvkbTiw8uKsz7fyHzS3
hO9QQlQA789p1HH/jYz3t3OP6YRm95teE30xsbl9n5EObFnUcC1HX5SZ4HwAWISQCdI+C0UpQJNI
ctNpr9mQkZ8wCxqbodane0UFQTComklH5aWN8KqaO5Ec1k5brnfbw9OOS58hU2OYl62ENCV06M6B
5r7Zmt2LpowsfTceaNuuSxL6Wpf3eCy0F3u5gu2aBJpRt0Q0GQqcq0icbuyb+ij7ZqSYN5akSuE9
e5b3Rjh+VPBlJjVGkDj6q2qvLdvTu/7mUOfn9q8WkcaHCQ1GwteVt9X/Qxs96JvT5KbOI4PfRWjS
ZJAY8U8CVPsayGp3hcGTpIRBaVt69GSXJzfbncUHbzHfJcRfg5Jmg1FGIZtpqmDLB1Y4pV4ROI8P
uZPaonRgW9UnDiYQKtfEy3YZUQ4DhiLyyJdwiCv/IGks/i23Puub3De200IQXoj0ZUQOHDckazJ6
dDKZrzYD5j9vRX+vC/mWlET1BXTq9k3/d80DZ15XmsvAGUrY4B7luGlfSQnkvnlwTcoYEyHckH1M
WJjtg0i9apJNoB5jmI+gttUPqDrVzQ6z7QNlTjtT8u1ZCDzaCEzPedMEeYuaAfNzxI3OhVmLm6IH
Jv9DbSVNKzsSw7YpCSb1VTE3yZvh2hLodZItOmB5ULmHwk1FQLYdm+I2G1xxnjtmGagMl9FOQK3U
d08RRB9zk2wtVF4Z63AfxaPnNWkAcWRCAiZPgaksW0ydKRDd6s8aopHiZbJnf7FbYi3emenyvxVh
Fp36mJhLuT3NE7/xvldetomQSd+AImeKOyUrBuP4rKgk2Zv4mRl09+8rDHA5vmfLtCciCBRfqIZi
/MaFr6XjNh4BdR9UK+9r9onHhZ73fNnzmKvobBUNapBt9NjMIxAKvndtSsvVtt2qPbYcppJQacPi
WAADPa32FWLEN0KSi1ohuWCSIA3AvvXzQHCkKC78Um9vzIx1SpinHUfzfrnslblwnXJ7kjao9MAH
k82qRybXPtCT625qOuLLlq8HdZN+yL670WMKblst2TzAn6lpzAJ/bbdPkbvvO4xeMQa9eTIPcAFD
bNlUQY/wZkYMc6eR/40K6NWDOmwO8H6BwP4TG70h5oQLEkh1FJKYDQBPHMovCJHM+ttM0/ydM6SO
GX4xfEyi+qAi9l25j3702tIn3y/y/5A/0tHDEMkSYDUMN5JdaM1sb+VuQzM1mt3i82UmVVPeYZ7p
35tzIoWrnn/kwTOUbhml2gg7+wHJx0iOPOYXFygzGQ6ULHtXLRaN8nt24A3XAdhiQStwAUlOppVL
LNwiQSS6GdzWWas8p4afopq3zK+bAfp8U635p3Rpvzm/0zlKK48/PHXQH2esWghzWMWoUeVitGKR
MYQy/Ek8Y61F6vaxEYWClhT+7Tw36uRNkn+/DbrtT4RPz9dj06HOmG2L2NZhOkzuE/tackekfn0E
VmHEhQ+9zPoxInMy6Zy5to7JiTo70Vyy1bycEPwoq8UV+mOUe2bEBQVLpBy5jiM8odJdL/aVVFAC
OOixlR1g+p9jzWIu+4yh+BXI+onWABi1AbjYqkkocVUHG7mqZpwDLg3zWoyn3B+fCt/Ih4GINCEF
EEz8/XqKu+m1x5OaTxqnhkWLlrsfqaxTJtiVHU7yj/e4K5MgSjncXyN9SWXaqaiYKTGgyceaymn4
mN004eUROMwm4db24QRsL+IKxKaXNSIBGDVC6oLvrLiMyq/QFe4MLQCcqmI8EIii1WD0Q7rzHJHq
GRLxLr5t5SstMtd6LLt+AnT1UEZWC4Bd7sBYjmaR8FvtL886Vc7XtPhCug0ixqhMNPSevVLDrfbs
3Hvfu79wq19KoIT7kmPS/CqFbRGxukpAnn3TxtwO15XJtU65AvyrrAx8/1xA3mEdX4CMNR+uvckN
rsB6MTO+1H67f9SgqUCkV9UYEulFR9wgx3CyUHDRmgBCB+AQZMDPNF42Z+b30xTRHR93tHfyM6WI
Oht63zIgTvD4XY7TIPhFJmwW22dP1USD5TAkSAIPwikDMMCdFVesVI5PiP/VtKh6WPiAvRBO7dhL
qI3UkrcTupYXSSuuC25pzoRSY6tc+Ymo54iH1wPtmH1lH1sAf5C8YbO6drrD91x/kO/m3Za9mmpK
7tx3IFHpJ8CgHTMjRMrfzJFxISMDoOKYkUTxL+6yt07Sd4WAkERm5O2z0WiZ3N2OaXvkknsc07D5
Qiv5cMfbjJ8BA/eMH5edwfj04Ucb/NVHP1qBnWoCsC7GYLf72bW6myE8HBtOxK9Y45bxX0bbRBXw
KVRqo/YiiGRaUftXdC3G/LbXpUwZcbh0H4qKgPGzqB3HmnjIb3y6gKFjyhbMPC16Yxn6/jrtMkmh
l8O443AG36DXo+oLHz+NUhg3G3xlpNq4bqRTf55/tCgMz2rb9v5p/msv6uBkI0HyrthAG9yyo8rV
KdjDjohE9t8gsrF1RyPwUJSt8HSl5QjZVbjHuh5njd9qAPQp5o5jXRxK2uY3ccD7+vHpDRCfGHvU
52bViX6xPt4hfGeM0PMEvtIybP3ECfYBCcLORrJGXkU0LGickhiGebTN746Q7eaXG8JefKwPVF/j
vaj2utT18KKNrX56XIWJn2iIT+RwKc2UqmZxyKCVqIwBImUTylphvZZFJORD8DMugt7JgkwDvB1C
Hn+dfsxhoWK22bIrlLXKQVyljSWMkFviLiay1nbeAXIK2xtAEDGggFNFGiaf0s4pgZsxmncQqR/q
oE5Wzogx4acRzIgoXgoMBuSUbpk6cpRwQeAEEWKZmYhAkT+iYxM6rANJleTcx0a6o35wUsn7BzRX
qkPbLnQQ41/nEUcx2D4Er/ULHeZr+x8TU3OPqQIVP8iNFaTcf+Ya4X7CDmiKJUjahEVj28QbDck1
T3HZkk0hYvf84C3ecCVaV+ZhEhw7G66MwkxD1VQF5LGXwyXKpJiqMOa8Uol5uz2WzvQCh86dnNuD
flDML4e2Sws/h3mIVBxg5J9w4YJH5o79NE1cfKH5ApopSwkaZyK4W9VncNNYWmaGZdjWc98n9h0+
/oM03KZHFEGXmUoa6jtsn7y6M6P6YHkNzdtdc3Qfxd84dbCln9CpJsKxEAcj584KTtfxg21m9pL/
6Jd8jtu+A0YA4NW/nIFhRudYhWAws1CjVQcvBZLnqb9g9b9k6j/wgjbRCwjZ47DhiXHUNj9MJFGy
/VGU1k3V4nNFjQYhahDFk9DYDF9rnrd7caGElbRtTJrwhGD0wf3qAuJNHs+EUA+Ft2gWp1L71OWF
9QnNykS1ffeIgWHevMB5uEEEGblnGRJrvgc3G5akt0T9xWqVXvCBn4n1MgNqHBl+ByKUM3PkV1nJ
5aUCdQPqU80WgeNXz/fc08yo5KOff5qlAXl6wfVpuIgkdn0fYPLdqjtqOn1Oldh0ToNav8MZX7F/
svWB1baR1ZiERKdBxshBeYyBej6NITfwzx0Nq+Wv6iqdIs+7Plo8ICf11E4mvs+RZkY4EOE5zFry
PCRfLwoc7mz/fRSchi0Fqc7ymn1jds+a9eMc4ZRgBckjSkU4wuVOwdXDHHOuqc6KOOGPPYZtARBo
obYshjOFdX5ND2QZlBk3RByiljaoWZL1Zlr9OrBKUsmu1GMC0iIjrAQzqX/VViJRorc/lYR4W01o
13P8Coex8eADI/lyY1d4WDwFUshbC6ymGCtzMcC6R3kpeknq/R3no4jc1HQCtioyZyb/bvlPy/Y6
cZvAZ29uq1IarMK1Mt1XZglvpwlXdP5uVHS1t6KlqUbXK5Qt55+kDj2oD531dLlfzW9c4E12nmFu
BGeCKUo6bmqdBJpoTgcr4dqsJHocO281vuoR0rsj367QJwdd09zxCs6NXQ7eQhqDIUQw3rjfwE7+
FRSoxBQfn6E/dOv5lBd7BkIE5yYbvqnRGrBSLZIUm+6xR5PcGC2Ao1soPV9HfZh+0vEzEbA5+i7X
gST51DEYhTamXe50XzMM/tm6RyW2CQFts/XOBftmZhuqfOjabRJKQSe0ZOpL92I3idh6fz33qGRM
DymqGDQ+wjZTd/jdQkIxZkGRd4N2zGs8mWg09B5WVsS+bLh4qt+y0VEAC0LqQlYO3XFNMytwVHz8
EIL6Y20guantGlaecLN/BS2VW2KRjgEkl5IBwSmW4lVqMgi4YGbR8uzNrTN8av0jPx9KGvZ1iZtG
yRXTYyDnBPpOfIskIrIr4rILvdHCxCPjn1U0YE/sx22SQtmrgQE2zEjSSNy6IRP1imu+hJVd/LWE
mHJslwu9LgFNEd7oyL5GvV16NCJJCzVbCapeFShju9nyXqewo+wEUoKaK5r6ovlISnW+/ArIz1De
YC3lidTKbg5hXLT2Z6Jm62JY143E7ohtUfsSIyO5HK93o8NgSUvaoU0Y+6uMpDAAR3FxE0UOT+3G
s4vhfai34sWXENuJlWHWdLwjvG4bgga/KI2N99pb0FsrjFJwGfYsDU63l4lmoWGBOVHDnDK72z0I
Z7QlytwJFVDF5BcUZRCa0D4TBLBqruVgFxwW/1ZBSwNSgle5CA7lgrXJgXqmdHUBrYWj6MrT1rMt
huL+vk6uqOh3s3jPdWCx7wPVwWDlcRrH4hRz8RljBhcK0GDXR/SqQyJOf+ZBEE/bSIZq6T/xfNPe
m5orR8cdvJZKvGN8MGD+E6xfS1WSPjLlaoHbtstT/Ff9fUwQhfRo+61MbKE6Ye2holjSUlVS/FsT
pQfUtD/NQegtwYvbwaHwuJUkHbROwH1r+IUmgu+5yplc2PTmhQdI6rSkD/afzFTdgIatHgFgsuC8
i+ywsxyFsxoVOtAtkM/Z9C7SQFSa22nGzuDTAcRRQXb2Y43+41QsdvCYu03fJJ+QeqIOkIpFTpxV
pNHaXjy84kAdlXTjNH0xfwYk85lGjGLm9pjcfZdApH2kQuu90fdAxI2FxxA3MFoxqOziIgT4JeV1
EjxC4Q61eoKuVLA5aXv9EYW11XqP1osKuWvLrLmmnqn0nSYds9hqN5tZaQ/epy+AhbmHcR+yTdxc
B2qOP9fPimpXPr+rkgj/JQGwmCjfLkkqipz1UWHiw8R4mIIdYzZUNch1mBWsxtZq76z4cRwhIZAC
Epv5WnrZwpd0tCFT0p1BA5aw8vJbK1n0qQ3Hmw+ZypcZSdDhLfPV/xhyyeFOk+fWJ7chf8nIn7Dm
etXZ901l+Hq+ArAnQj7qHNAshhkLDSM6Cks6aXCGuVEBlQhe/DHfJvzFT5tbZ4+LCVFTm+Q+vH9C
iQBdEH5Jevx6YVUhzV3mMbf0B4EKqvZvggLDweK9SRgm9xN+MBs9DDFJDpRh2SmD+H4f9oYEpiAd
LwZquM0U28zz94oTY43wV9zEeg1gNGXP96SNn3wwdSMnftRsz9jnV1J7FZygQUwK6yx1VpDefdNw
PDECbQ8K1rguKsIP6zalYfkUS1aIQnd7zVmG6j88oNfaKeIV0UJHdtZTW0nRY9s9quucGikUFype
057PP0VwSSdNtKueRPmyWTaJF98CFfafPgzmrpBCjdN+jVsLo2NO9809xgqowrvAKCsJA4vr/RHA
TD+W/jAzJCOI7Tz7SH+vpcE+ia953SXk7PWXOjzGCkQr21rlvib/GYrekz4MEXE+lcDM88u8TZhz
BgPtfz61guFYF1eW0Ef6q6RL7s63JhnCkqzynt7kXvMOl0G9QuIE9gB0vHGNdrXYEW/GlRIWgZPf
pVOSOKxRfOd27azkkkRfmCF0HnkiQw8RdLvr7uYzv7AJemq8mJCH9ZCeCIcndE8psVNi9W9gadB3
GUtxNva3WEf8I7tiSh7vfmondF70OGpVKrrAmZpHaPkf06ueuHxxKtkclbTR6QChqRP0LuP7PGQH
a4T5D1lvuvFHaZ+Kghcy3Su0j5rMEqnCmcQ/7sguU9L/Fx4azhasg9zjIOvEp1V1MhMDSiCm2k0G
ru1xrqD2WZu+nU/DqZdp8DBhgEfBPlhrPOyQ8ZHrv95T3QN/8DwyNtvzdw1v9tpyiq8un9xBfXKx
vFkkAj4pzj/e0dl1+b9gBwlBn/M7vTWMz7XKdwVHb8RGYpCUYiVHAtX4CmkmIJ12qsJrVPPSAEdU
zIALDb4wy2/wvDdY4FUVgSFuDd2yeb6Q9anpHHWNTlhMeq6rOrVPVPAW/KSmWdmXQNhrJc0odTrI
DcvbdZHA16u5p9Xh+crmw8KuavBMcXHdEulFIttsRgs6+ev8h+Rg5h5v8B/dkY4ciLuMTPMieQl1
mVXK9Zq7zu3QrjEmxK+J/f36xoAPapf92ezR/HZ9KWSQcsCiIinSGayeYXGOllXkWAdRUI+2QTWf
tkGUCCOMQRD79MghOtKDGltewWVMBz7p96wUKeZSCj0sxamqlpZZgYX4LcLtnyzeSOeNJmVhBtG/
UvsPJc9wixwjT4wPhLQZ+EO0oUm8XfDZ+8p6XH3SaEPSsfEJWTJQ3n98Y8AirrGg1RVKZG25aZmT
fjYLA6BVzAMCO46rggvqYvrNw8DueJD4csVQItFLHoydgSczT6QK/kVCFlEQLK6E/EH3GvnX+vI+
kYkBtTebmP6b0VTvdaCFpBM20fbiAgOs1mo/dIh+J/LEcQkp+KUsLaTMt7IGlTFD7aATjjJ7frCv
A8GFCnCN3+MipTkYYUeJen1U/CZJL3W5HsM/0JxUvd1UhL9MP6VlXBedk5utFrYlD4GvW7+fQYjz
VbdGYErUS132kbDPdmwd4Du2CrrOTH/ylOqJUGV6i3ratYlpCcbHWA6V4W383gE5bZgy2hX9qU1r
U+hdORWVIIitaSScZ1zM1jf2zpHIzoU+DFCmpiEHtFRfD72z/rQX+oQfWIQBkHfjFbwHkyU+gNHL
LqKkW+9Hxwe+KvImreqzaDYdOZR2sGdCJKhRuY1eVhkNwtPpA0LPrr7u/8TCEb0IEYJnFZX/wB7Y
Lmvpe45ERErXamwYRzhluY/k8flhJv4l4QMAALjJ4ie9aniWGy8RHsjvXx+e0s0TAzyp9wc/SXBF
gGTDezvWgSCyFpZny1UGpclDXnBihViJxrQPTvGfNSzGENlyjCTBSsWdnNR5Zzf3N4oofw7mvlr6
c+z2ZBaqvi0b63/Kp71HEBS0iHWXU8RFwFxnf/ni9n71FUUX3yRGKnnqPD4RGjLm38JJYjq/n5ON
wp80pQxFRmIe77FYdkOx/7d1ww1/G0pO5q32r+RYMVzfhu7ZTB/Ab/DVQM7qof2PkNhmRr+4tE+R
ec8ZqNvQhYkfFYoguQoD3Uk2BE8AoFgzN0GC7mftFXqQADvNGRtpMA3vfQno//gb0vWcljZNmY7x
jUWDISIcN7MHNp+MNPoLnh5w1j0WoVNG3mYIVgX2jPkCPXmrnaiG5ag8qLJtyE10BGq/FlxNeyDz
k9GHqN7h0WfEhei+Fwmy0VtuypqHnZxZgczZyfuTccmN/u1wPZmgbM7V0EGmEEE6oC2ZuOXZbSQ3
u/GkIDbx3ehGs+mBycdzAGiZSPbRbJEs/4zhQULWVp1qkTR5eoWkbVW6kDBjpuFJVfrr78LDg77K
vwWnhcp9gOhOI4U8IWuwt+WUJiZSG0QuNYrT+s1kePi7Ee0sAunRv35GlxR946gOLxrL+H6K2CSj
82Ie8KFHz/ANKpBh+Gt10qqUWgWy7h2gsOp2DKGN1dUyWor/vhg75s/69TMFbftk/KeKTs50FQLz
+c3A1/asr0MF/ptMndPtSgZQaqXdCmgJhSdbVNEqEpriyVIx04ISnVj48/E1iN8F/2/9z/w7QDpC
jfU+UyrdnvobkHg9vLEaVaTB9xJu9VI77citvZpcKwrbZVSrt95/dnHR5PIhr3KEneYuXkLWGEhT
wG1tLnRyPVcZjSv0Ys0z3fnHt1YK09iMiMKCU6DYlb9B6jFNM3oaWx2M307/3kZKg5S/mM0tTioj
A+V6s9gzL0HRHLASe+i+UxSA65HSIAdL/kr0khjHTiKrMqiqe2FSre/J7KZik1ymzF6c2+1EFpPo
elwTfXYDlWoO9hAhNoOVD6fyFNx99iNxeTIfVxSTaoNQuBiODFZ5h5NFlIGN3SMClhAMX4o11UK8
peZc7e+DMqMKF+G0CmyD9sHUDIHEsEgh8wd67x8XvXqSk+m/7WaCrONuHIItoALoGeQq/FFg4mAf
wivGvq80M6yXnaSX4RsMHV1hSp/bDqqwQViGL5VX5HjCcpMm8cLX/n0fLGUGsLLWOE0kioM7YF8G
/g5RWuZTY02pNDeV5af1KfCEl7mjPGQBID/GA1R+K50zOtykAeidHwKTeLQPT83PCMNpebHFAg6l
4e8gCbeMIFLtDHt++f9KCTellZpQBOJA3bPFptpZMRHPo5PXrQIfh+/OCY1yK8vAtD8u17UHmjNP
qFWHi28U045KkrF0lxG2K6ssDjDgvvCsP/oIGpR8HEylAcC6CljDGsYZypOiS0rNW2v0yw9nXP6i
qSPWsyFJEGDBi0DzBCvpHRblzQ28wuHRkgBMuB2VI3GD2hcGQCd66vluwWxI4F5E15Fmwj6wDkMT
mJ3kD1hMrJSlivNC7qEDaTudbCytlJssqg1Of3fjG9UMEoj5LDZn5D7OZEnEfWYcNLf+lsADfTpz
V4sLQXyq3gB3v+wBgctpCyqD4e4onluD3UUAYhJqw6jEoBdptECNdMF1YLsjo1Re/LK9Aj52Am8u
0YhcdWkWEcxuIfT8bxXCOjxvYWFtlIe66sS7xJccyrLuzWjLwxLVVggUlKp0DTKZncCbN0Eu0tL6
8a5T/GLzFhxP4mt6kiceppeOhURx05p+zx9x36Ja8Uy2Ju7WZD2EFxqkTLGcTicVTmb+PY8wFGvI
BK4cgglDPlN3r2ywcFf8dkZlFIw3BXvW6obqC0kiYXSz3YKk1JHqmqV0oe4ISjnmx4ZjPvDZOD6G
N1X8hKhuwEkQfdHkXP2byOaE4KD6IGJvUD2Z77+vJRDla4skGrXiXXzMtgmG21fZlF2v8jcLnRfY
aHkarnljFbLPJqcW5p5AEzjCQxsxQpvxETzmQK9e4rZEiZC51uMol8Uy9ETD4H0eO+mN6v9mvh6i
dmmKhZuuZkobQZswlsah18PJZU1NNgxUyFGUIMs5ScYLnF5Ps47srD5qiSNwmoIp2fnJvteg7mh1
TQJcnSgCVXq1ijBcEHAvWMoBLtx0giEorFHtxEmGRm9s/O8fyiw4j+cW/wKWnsIHYTe3/TG/hPIU
pUYz0cG9bhXU4Th2yl5UntIeYFh2Xx9lbMbPCA5nwjejWIUj4H0Iw3038PdQnmG6QZaJXnSNJgQb
PnPXIUCatN5zzJ+8bIgCDnD6jes5X3Dyc2b2OimYUIPI6J+VJnopwt8+Ds30lJtcHDZsh7H2Mlml
udezCgc/QlXl0FMdqnazrHvlK5QXq5B/kjTy4T+CxY4AgXfeOBWJ6JyNamaNIABEfgzT+4hiDinz
FR3HVA/1jbL00713tN2hgMQD1Q96w3g7TPP+Mc1AmRaVTKgK6cZ97K665idHrT7Zg52iHQJOzlIs
M7zk0gdAzsbhlOW4Dka2io5W+AgODGzP8kkVzRDEgQEm7lbnSigYjKOr2owGosy53l8UF+uZJCjx
9YZwTsjLOQpvCaywzJxeBr2nNHsxHUHA5O+rITPi/mzu3p2OxCfQ8hJn9+Pz7CGLx5kDDoo30hu9
c3QebQs4MnOm5TD0ZnD+CauQsH5Rnu3b5JYRgoyNgKxww2UCR15UN0XBBtEdSKZZy8tmgGfefsEK
dfsfBuL0Z7WChtFZX6sDnXl/kSkUx4jHpkAfoI0XJquntXcOlD0is8OmimYf2nN9SHTKW6hiKow0
kw+fXlmBpzAo/A3IwcwnYHvDi8nBnG20v18jVKVKDksWOKsqg39qZKKeqptsouu7awwPVzoJO6oG
QBfkdipfNImVlK1YQMGKfiLHnMTwkFUwCaQHgcN5DklpfF13D9afNaBF8NwfV1UIq3uTvvV13Dgv
koIluEnSwiUKpzXwnBe0nSn+Q8lE5esgD6ruJ5OFnYU672Cw4B896F58pHVNZPdD43KLfTkULE7f
yzzH3bU3An3EIQCf/9Bf4ZYRJnCv2huGBHRnd8dV0Mrv3pXYXNc2bDGvlAtK6q0jeVsb7PXiU1VK
CmLte0j9wpFmxJz22PBioumMeqyPAb5l+k3aLju5zIICTcibbQV57Dym+atH/0B6lWe0Ton2vDKK
e8U82h9T8AVR1e2MM0h3hL4B0B+VJSrpQ84YWNVSEscCeq1yAtUIs4XfaRnXqC9Tz1J4eTQiBzlX
gKiJl9OPCeEOF+N8Sku8EX6drTFyRgG6+DjoVYlaURwre+DYIz8ONzEj3pPYB3d2MyZWu1H1aIXW
+0HxK57gWaPUTAQ0KWuMW0hzixBL43O2ivlTVBfH96ISGp2i9FWGUValnNnKDSX7Nkb4yvFef0y6
1c9XFra2CSeaX0mSI7nIxXdVNpmSc1Y4QpWRAH3CgC5cQQKvvGTG617AHzFaEkTNSh9UVLM8Aw46
YKYuMZx6isEqVTWoNQFs8l1njlCdj16cfLR4ASbzP1xSZdj7zxtuf6i8AEZhlZt2Y5IoJUjjMDaT
6jdpCuOWZMk9JaCDsq8wnpZSFkqA46dPMG4TrkI31iIVAigYC1wrh8ri5GKfA8g50tHi0gssD60P
zl1Je7AlQ4uOqnvFSBGNaIplKcpmOgV8Ru/94uAfSIbCrqj+L1F59BDBfvq+ZsEXSMcyF5YCJa4g
q/AK3DGgohaLcKcGJB+jtXh8hWPXmgDoYyyN/0fgrQUkdIvvZSAbOH8XB9iLeFScUOEPwviDk13+
OKGhVHpxM9TKx0rx8gPGoV94wD4t1W2UmEiFstZ1ps372GxHJMxL2q2fU90H7nvdTTY/aQw42nFg
D7TkMWHq3jKeOFybSICNfq/xgVwDXlDM4x51dyp2TuW5dGBYSehCMvWtz52Pff3TDmwGfmRX1Wc1
oioUwj8kq+I1MxxJzKJyRELBubNZ8M7mURnYyIxkUUlyBXHcZG0bQkC6VyxoLymc/FJF7OiaPML8
D1XSisLwcd/ATlUmX2ybP7qcD2Mv5X0bgeWIn6HvCGEFKSpsGvS/v/OgtmtQvP9D5n+gX9iYTBni
mgQB7Q79Z+TwpJWe70SJDq8IwoyCIs23L3FivBENVtA9b+I4/j4eTu+6DzoOrg5rBkHTDytOTytx
GVFufXKb5inh2tHOp0mRCJeBEwdzT0oW0jYrSc5ezsY/5vDPwtchkZ0e132hne7d9sxVhLWd4LQa
q8URlblWX9oalDpujRieGbpbprWgER3o23NXS60h+dKYXqrIsWaxCOtJBmBL4zj70yUTrx3BqYOj
hhnZEyDgwxO+HTLmoap3EYruZoYymESf6IXjJfjnSaqpX7WqpZVSXfawLzDQ2tzh0rG5m4lIEtH/
iCywnGZppO13fk19GTvTYwBtDGdkE8WEf/sRtWdBrYiCVXJjLkWZAY8orTeGcSG+gsRaEKQY5zlT
XueSQAev+4Duh5ZrAyaAiwxsGsiCPxNGYYfD7AFwtCso1h0p29fZ04JzVqYCa9jftd2obHfMuF1j
WBPC1TS7x9/SnttSmqbtInbAz4D9CX6ZxdVJi3h9+hxZ2OlN4gZY6NRZ7xz7m0MboyJj0Em6lMLG
4jH7OEc97UTv7pbeIrZtu6wK5dh67X+fs/9oRAEZbmy1Vd85b2ZNr77PU8DXqmH9LbiP1B9DW0xj
oG6Mw37k73Iqb1BR4UyJGWAgsiLluPu9CAsnRvzuW8QNw3L0lejeRfPwvnCh3YmntnFBr1Y8cAZk
R4oTu31yMlu7Mlk/ZLvvMPGY+GjmP1x6DJp9y8egFqLyZkVd1kEhiV00ezpgNZ9fNR0j9ZXpUaYE
JUy6YPUE+3GlPUgDGFEVXxUIZDdjYZ5Fn0zH1OsvV5b93R3BQ4YKvx76NQ38Rd0ngga/24mKT4o+
g3f4FyTObKrIxkeqhRcDdo6qgeqsq82+KerWs33MEnJ9XKncbPz0m1hM5110/C0De5c/GhR0VhLS
uu5j1uPy+5ipERCyYcANDeuxhePCI/iyjklehfb7oMJdxRho0AtvQMfSVm8rc4Dihtn3gXrl4PR4
MIQF1KHdTqP68ZBf+PQBTnWfbuWC2QAKBN8iPs0pCgGkEYx/7pe3dkPIFTNEfZy082IUx3dmAh54
lMODWn0AUeBQ+ggTLjFT6ns4nkUvoKBv7wsrP7AKWsmL6bda8qRkZKOKlzeJ28l18/o/jWZ49V0u
A5PvnK+ns0E+X8F/p/iQu/VCZylV/VzcXqIN1kXxq0vV1ip4d8sAT59xIGzLr4f/mTMRR/ZG1Ws3
92j7jvxAT87OWPueKsym/q3Q/sba0fH+qPkSkjTVUe2CttlJV+p4F7j0zAtrcY2XWq0+nn+2CM1a
kbH6erUMOx/4bwBK8j1XHJ6Vp04Uof61XTX8DIP+F/C39m2bPUyqd9QGqb61a2ZcE+1lrf8E1Ntj
D68KWvH+bzyAm/8+Rs5j3F3fqekNLEe9bQWIvNSa6gjHQIn6xFrmWhF9edUCAv6btrfkPxpiiwNo
Gpz0Ig2Jbjn9rPV6aYIGB6O9uPJO94p9jXgAZWhQr12HWgMHMKLXOS9KaHdzGUk1AApfinr/1yUs
hSTCNxv/jNpV7l7fY0EnGG1Gb0Jsf5OyR4PfORR2OEFbyVIJKrVeZ9kR1Pws0siywjKa1KhLt/IE
QryJLWtmewlCJWGElLxiRU2V69yTggBUmrFlpGnPwNHd94FUsfJMenQLQer8TFA46/8zgmnjE+sX
HhNLIP1ccMfoFQQnh7xHDP3Mfb+6E1YPeTAvoyT+xtlOaxz4jod8eLYn1uHTCqq5xziDymF5/O/r
A01TooZ9iINza9MQZtaMSKdFnPKyFmcG3yG+ktqLpnnHZeAs+fSeIdFekUFhVH+Ci0YYWNTmVJen
G7QTGnHypOkaupSh2salTpL8D19xO0GsFLkDJpvtO46FpEID1swL7weNPfNr7TY0JnSHREvb5xdJ
FThpz221XUm/kVYUEcUJLf1dt41vV6Ze4rqRLC7vSRNSE4wVT+BKeJRzdNxdH9FA2kQHgNPfNkFZ
QIkOvBCQ6Rie9vpE4orZzv/jwguJE5T3mBvN3WRFEvxmWGYAlbYNOd7lg2k50ZVjlLMPTSXdgtNX
lE9zxef3s4/y2lfkeYBI1D7SRRTw01JXy6gv8htpTQku3R1sJ0JqR6byjUlr7A0ToFfV0iif+cB8
Q71bNmfBvVUpnoxtXd7SE/dCimvgtAnJMH4wAyW5GiEpI4MdowCe49v5eWX4FfFgAOgAqLNyA+Ei
BPe7QKZjHMTY5glcW58vN5GW66R2UMy9OCTRiU+VPgcjGKGICbeJSrv98zgfps4eW2i13+uwPD+4
x6J/MWnQx/1d4p87SCNDDq4FftgEKWOfhdkZpq9LG6lGE9EQF4OmkeILDzRe3BgLn1gfBKmVPrOb
AFA99fqK3/ZGSn1zDw1H1mUh/0lfNckhiQ4beHxKBkFzfZvLX+r7O/jecbCHoxUwpSXsa8oof+Ao
fcYMC/R5mMNpKzPWkKM/sk8H6RVtYRoHM22HKA+TtiT5baFjKfWTD6djpXvps1BY3KtJZggASXET
+YhF7gDiutwXlwahvze94k4hAqfU7H9szzt7pQJR2x0rc3dbm3Bbjz5/clZr+NygF54OGzkEmaQ7
Uokdl6dlrzGyPkjku1teiOjEYKZfbFSv1n50KHTvv9AXqS7i+mf6sSFoHkuwvqqVAhyF1w4n5deK
cI/iDYwZVCtjitv+mwOX5N0R58NLg3SKF5YHLPcdB/nm41yPCSSL6NRg7B8atnzxxpeuQ1xrlFeW
CpPFcwG20HTCpm7D9eNTNyGGqaNb4S4daZ8H5e5cUQP0XCaG7kBS3t9dYp8mtVUfjj3f5LQeP7Wz
A6G3/H4XdoEchgJOWubx+s2/19IP3x/EhY3GGx6dz1pwZWyaktX2kriAn/ffmsqB5zsP9hNCMsJQ
a+mMXtgmOEMlGWQowG7mLf6uH6ykvhg5tFRJOiv6KmWmS8k8oGUDJcR3lAbVN5OCFSDbwPzYc78Z
iDmozbNTS6IAGOyGFGltywWKU8to1hnSDIhTSiKo2THP4C7tyK/wNnpjrbNIO4MxHeXnGdk5311c
8ziqd7kNmEioykinl3gHoxGlSkBA0oIceOPInxDghDiR+Z90OSvRHixfzxz6TTTSXOyu3DKgtnBI
FpVlftfg9Byj8JtsmbN/m7Sit0zQKsPUu8TWSuvFZ8qoQ+T59FOO1S7TGHskVg/KGzFxlN47MNyl
xgdKZlWBVNZxlC5oeOd9mKiclYCgKROxF0HxzKhNOSGKR+TXBDu3bZTyPjiEJjNyEzPdj4EXQRU2
twD36ymHVlQzXSFRmEClfieluBqQNI0hz8x6Indt3ggaa8qFV0PpWWPNrE+tESf4gyZAySUA1HnK
Bq5ejbOIU32OK2HoI2J7K1NEM04MsDySfpq20bcRerXxNN+II/HwnayFadjRjo6OaKxerTz3ZS0X
wC/n5dXe3Z0jvmQnsZ5pVjov3JW0T4Osef3k8Ul9ZwQd0Vn68ySZmx4/e2lexvNxYvipUShue+Ii
Hvtppug8ZozTLdmXbjUre14U78bk23vS7OtIygVcx2TDYst8QQHzNvtxAQEZZmCztLvC1/GSJxLT
JmghcwOIZVwsokvCOGvbzhFcrjiqG6g/AODBS7Z7pPuG9uKSBbS+DEa5QlvcFcTae6CH0GQOMFnP
V33/C+mxEDrPmRwlUQ2SGfX4HqUcf9rc/QLUjIfsc+iRmphpprCXV8qxUyye+7WpWGyZuv8RnJPo
oDfg/GScVFd1nMmn0hjSuI6MzJGy0Kcj84L6EPzwEMldzFuU5qNaeocwdboZM1G/NnZEb7ZVvRBQ
ZiXCU5ghp0vvtH+qgvUeut7T2MTSHQqDWP1augMZbBswHKTS45ha63uMEJsTUZf6X7vk4BmCv2//
ib0/lFT8Y35S6wSOyi+JlDNvMzUSOrdH/JnL3GFasjLFaju9YLCyHlB6a3jFI2+UcUQkYBHiZppl
GwKJZnfpvT9cbSCgUXH5dQAbDCM2dehoQ5FQlTL2VJt0gNuPc2hC32LpxoijWfZbCA5k7k1ZoxtD
xtlncCgMZ+IdBJREPlZ6h0C73kdiXXjfqs6h1F0Sj9fJXFbrV8lRKMfx80HJ/8AzmrL2Zy/9hw7y
QPdaYJb6mHjA+lku/mr3Z10qTS30lohurVlH9OjWpSGspp7GG1lUEmDAu9ikwI0O/1pj8x5kmy1D
h4qxOHHRstnXgL2WiEXs8sXVp/SHKiADP6At/MoyJZX1C/bqOb2N6BS7lnLuX0ndbKCqlerlGsX7
A5mA4RIqSHeHsE3eGHxAo8M9y2JclBEsaJRjnXXYHvPRBUdXsiPVO0k5TcLsFhJ+1lhbF0kNTo+s
KiZTvX0IV4TiBcU09mGUok1yQ6Yj52uA39zM9fZRnC/8hNJEX6eMzXXTsplDb1HNRGU8cQ8P/VCc
ncWDrNgtTpgsX3J/hohlBR/dPk/8w3kI8GvhDqZFZNFhh4oAz6TnHKVegZCTpfo4DNsR1adxuetG
Y+v4q/MUXALLVWXJaGczSrFh25JyGYo2SY/Y1Itn76M++iSAyOT4L2biSxVjiWPycHooUS8ZskcB
ZnpXx+AQOo/BXSI9uubOd2fgwnAKlKXrsQL/EJsA3pG+gF7iT3zv0pfD7/p/dm28hRAg74KH0Ox7
0eam9UeNra20DoZaYnIJ3tQLhWgP3EI/6Xa0i+AihfZgI0SUGG4l9x3sys2aoovpiOHbop1JiNcD
yi2FSTWEKU95iLgpaLSGTx1xdObX3zrlG90S7cec2rosnJ7PnS/gnGJ+OiBnEz6Q3Ncd654NZahk
pK9nn3cbmPY6oGt51uhm5eaIGF73bwW+buCMJ9oQDXn9+PIRu7nhCY0C0HHV7OxiriV6ZXoBHQSg
16ktwH2r05vRKwloARCTz4+JHs4PEST1LSGaWCRKTfLQoSGhTph6eq5zq8Hr3j/g8PT8NmuqfuAU
XVcRTXPpkvxnAsCMoCOX/DjxiepAgi29fwvpFoS3SHJ4E2yMNW73EoeThtF21zfb+P3OdmATsBVk
85kNq2AGIZT0ca/o9ZKTAtk7pxRMw5HttM20pcskWalkB5mTbiRPA5YDdKiJkI+0jN3/4kV3d/jV
cErhlV9xAUExbEMsbmlUcYoMacsAgINCSVE1vva3LzaQlzKPbHnLeiCuuLTWMfCOLX20tTC8tKTJ
O8U+QvNAHfJSwYZQXUsMkdw5+1+kdJdbgl/JBjZcNmwOD8auSkwT5urU8CIr74yQyQ+r3dz9R3Ci
d1zzSysrZYC+tlRW37XNiT7TQTALuLQCHfAijDyw0L+WOKC4Z12Caumuz34bUxYE+m8jaFeaYgAu
07RoI6GI/Jiso5ethhBgPIlWDDcqTrEcAiI4PkCnb/65xBuMVhQvxdifz6jGk1xleRIj3iNCTW2C
nkqHybanObGKMp951cOtIKekb3b1B0UphKGgNnPytgyZhPhPPP/Wn5V+EHnGimiDm+uWrpNakYS/
NDNkRNK3NAjZLZdqgof4x2ZPg8NZUl52tRKe+D7ThXD7UkxwFohpVzBv51pcqaiv1d0eyy0kSB3K
CT0Y+ZZYHC4/nN9OeZy4zYz96zs4Iznc2PhYFCfMUTFMyiW8Zq2f2iWGLKC6CwXV7bnZzzzD/ux5
mt81KV6rPsLx9ytM1135yeUJ+/iQkR5WhNkyOQGVfvkrsRrTfV3r+NK77B0YGr+L9a9h3GhmHo4K
OHzxIOVuFwzvc3Q5RUhMq5R8g/Y00eE9m0htoPb14kqc9XgvOuCowuE1K7wq+KwULCnF8I6mUEVj
QyUqeS8NiUr7y4ttn7CxIsyugS0s1Dqdy9xBQSvC6goqu/vNJCzjzx8TiHgyAAkcbcju6g7euswR
vaPjh+SeHKePaTzJY5mT3V6kPjdxRhJTgNsyfi9Q9E97IkUfq/ocRSBDqwdq8MzJ17WdPDJS5/mv
272bAscYxTRL591s0g3tD9XLhYLv5hfd9IPogSUAMIHX7lmatetYg5lH2q/1I4GWEkSBxsEak75B
fHf3aOhWOhAE8I4KHO+c2rxC4rnrxo8OqpF9iPCV7sc8w9DNm1y2GJjZZuDiGYX+OA+Yao/kh6Ei
locxR322Ungfj3ZynWFF9GOWezGyVnhXfzs9qlo2PW09M2sC4LeZeWt4WDWFdevHTS0XMdR8pfV9
88Psc3+ValY9rgM1js39HGmloBpiKbBPTBj0b+b1s/psCTB0H3y8KKzocxU3o9cAJhXm4kvyoCt4
6NyAX/T3YX4b4zJYCdyZfAh+RTqYeOEE0TWkGW8sVTQOaTFiC/bSifdwAm55PAlBOczp9vq3JI8j
mAzIohAIC1IB8Jf8XK6++m2wKLH7NI+AE/3GRxgXI8OqGZCnpZaD98HaB2wSHUgo1Di1JKLROmEX
4Xv97VHkcNZiDJ8GtDN7lrTiv4egv7Dvqi8rbTXKIJ1PqB936CcyImypOSMa501CvtR+M2vPj9XC
QKCZFPD6u9m08W41GoisiRNdURo3AmbjHYvqwLu5k6Ln9OChX68+d9bkei6i6rev5NKSIopiaG1Z
OKTcV+PPe+7vnIy4KA+DyX6KH5lYIrVtTM0JpowmchyDE2FFWlhHknaMtffiCXN9tN8F7fIYiUgH
218r6eEMPxNx0V1+XVf+gx0VxIEDiqvfHvJCczUcM+nbLwaSUYjoGYe4CLf0qkAZWK7GkSOqhBbd
pDFoqdpHY8cEw1p2HPO0VnERHUYuQBYwFaVgCwEbZ9+KVXM9bkDNYeYSMZ/df4wO+1fXT08G+LDC
5t8RII8tQRsRDCRYmCN3ic2lJ5/GtBuZmj9ruAHTQfraLlAwHfX9GbJfFKZVeUzTxzXYg3B5QSsN
0RD8sK4WgGOb2BkGvDMXPUy9IYYtxYx/1HsllBZvvS9kKSVkOOqfE0Kcfv2Q2oYNpNTETr/pmwDf
uy4trCk8wXE3hg7b7tG+D0jxhpRqmTFlpsEQS/FIgwo9lZxi7X9XweAq3ra21/BYqyCkXamuKEDb
k3GNtBXTBpT+fmi1B0HvhMKg4MftARqMMr9H9d8an1EE9Wr9b1sqJgPD3bre+Ext1ZtqWvvtUMDe
crBspgaCZxWStgVFrRizJiO8rDd5oE00lMeu6QJyy6JDcoQ19fEBe1HRiugD0joh/7Z+sUJLjRN8
5lIbhJYQ036ALeNILuhZN5PfH039dIVweACBSEq+xB01cYrOPAB4S31ztmf6TokzgUYdDfCFqpuJ
eRozYyoGRtkN7S5+ucev/PvNeG4R++Qbqy+qOBfqxcamDR5EhKqSaKkCV8MSJQX1JikmcwZC+4jD
LQ8jahvzPLzInsGVHgz+VYDIyN/+RQrCsZfx5yQAmpD0fo+0ie+w9DcG4G+juzVfJOy4q4BwXhhp
kh5Goay1czltj4k9QnEB72jrZJrZEK+G0kXdbJq/Mc/ZP+Z/UnUDXgtY7S1AMggoqQ6cNblZwQ7A
KVAOFJrtlH2mggr0RJl/TzghgQKF7GCQXVl3+BO6TU4KBfADmcqRnVpe0VXBJeZjuFh0f9xTGvf7
Meq+nak0i9Rmh+kevcNmh/OeY8w11OlCB0r2AL/xBWiWPGNkyTw7AjPrNDku0iAl87Y4Zr/TiiNG
p0f/hDzs5AxBCp2wImKi1LLhFhsHM2UObrFAFMmTGfcefv6VUTK61bGJCEdtKPUciAFkE1j7FcDF
qoAz7TE5BoKojjgMSFVzvkZWYFmUWa02IAdgAUkrZjrL9onltL5PXEhxnmuFLX+4dYvbmKs9+24p
X+upYmzdxHRscd+Yl+r815EQDod+6F519MJuLADndFPS4kAcaeUDKvYoCjtJhcqHRRXdabQKSEox
qr+yshlyKRUu2oBZivfGH9ZhoDqBBvroJj5E57vIeWhgWB/+7mvdk2mNrDnPoAoDQe1x4hexJVsj
nabGNSUypjxjyOhEjG8G7Q+OAmVsBo6rbAGyvNiq+TXt9rQjBPiJAlN8CeukYxkqelvRl6lbqs4o
myzGv5NEK9U94HG+WpvoicbSz5o8IF+KMd89gBFTWf1cIPQJPXoAFZQSwaPM44nrcMT2N2vveIzF
JhdJC707dQkT9plwlpthR/hRQdeFXiGMcmhAY3/KZQHmsDUTu7vernwR1VVYDUifGkecWvli5IGs
NZWRhANVsxauiHdOJIBCWBxq5uJRwwWt7/529jcX37QMDUmGgY0yJr1FfTTAoaLHe12XRpiPAcf9
8Wca2ddVR8uMyY9+owtE7yJ+OMmnwUrTlxuvXNEIRpIW93brCfy4VrqVYDKp0izbPAUa7vz1LGzI
YMie5+26PDUowXuEuwBwapiw636USD1kgIpFE0znLFBwmElZE7mblHEfJ9Rz+W8qy+3SUW5TD/YN
9Uh+m7LMhHVa1xGzvNKLdQg9V3JDhE/pPMD431KRtnSaHDvBj2onYQ92Rr9w/A3BnDmZex09K89B
grCOMKeUcz5p5B6NEW6cbBgwohLip5BytFagoK3EZamTxgWrQCPqFbSS40Ls25AGLMF6bafXRScL
ympyliQnnJ3ZJZiRGHq0AnSn9W+MVEwjbd3vpu3RU5bhO8LrY4ROj2enFO/P51cnKfj91YSCXx8S
HsF6ejllkIuk6MLnuyA55gci+SdigCFhcL74l2N13oMv7aG/zh0PTmKkojqCxfA8t0zYAPEoVFBp
LiS9ciYq6kKEiIvptczs/dRkgit/p8oBwpHMPLqCi92ei+0qVe7UDqokLUgmDy+cnsvWbaroIYgN
udD5CbBmKcE1vojHYYatRKTmkuSIN+kZ5zSRrBHyNFxTUW9+Axw6x/TL+22yl9SOUcUDxB52Qxob
2cLW1GBl60LKHZinm7ppCLhR2Ua8OnxkHL3ApIB2KVSQEsfub0ei3WR3tnOylLsduepVQJleJMeN
Y2jfHfVfUYAtjERW5zHoshpmjJspzkzWBW8l0Rp6BxiiZVwdG3WLaSaVjQGz40zwCCfbYc/dWO0w
KXEx+i12QCU29HLue5WRg5a2D30U9aqbcv8GCBRUBgcsHsHHvOeHy4K+exAXg6etCANlwpN/DlyN
kFceSa0JMNMlPlOZ0oU9w6cC6Avr3aHD8IoHl/i10pjHYq7XqZ4ey/Uu4a/7wIXx7kLzlHQSJiVY
3Qp86qOGxvHWuKhwzeGiggcDnRYryCQgxakeFNGA0Sen9xcyNh7hoOvvPqjTM2hfhTx3n4ml7b0h
edOoFcPvZ9q5JhTsbWIRZ3lLq3vaa6TXdVRwU6JELmGLBNPFrCdBQ2eLKLZvhWE57jfPocHvfo5z
qDmdx8+261EcH1HVmAaKuylMDfqxSeCSUvT8WdegjPb5LT9tfA1ymX4MjL3glT7X6P95u7Fj7Lqf
tTmPgvKwrDkNuUXF1oFr9ki274EssXkKSgKsjhloTz+NKyIEiGHjTiQzGpknsgkuBffgTEqITjzO
ftbL4sU7rXk0QGn2xOWwtbBV31CBXBPBfNB7kgxW860IjrItfxOfIE0aQyH5jsze0iTSR3xlCd0B
CWOnxm6okIkndq9zvDFaYvWcmEGhN/dvgEO94BtG3dzvEuF5cHrYngwBSUeQNYAUIyMy6Gx8TPLG
4L7Ackzg4uymDY6p746axTY5VwDYcgwsZxtP71oTHe/wSSrpRUnTJwQxhUE6SD9IyoFmiW01MWy3
xYY/sdlpV4G4uWITvZ1HR5CQUV5MVD6Y3wIDS8++JwDGipfyDMADYTOyNOnM9AenQbRQlDfs0ZpW
T0Zvi6NaFvkswJZgdCBJ2WO0rnQP9sOj0rIZGNYu0JLT4ZBrxOcYXvXL6wkpOtieNIwfJmHIqXId
sRxQU0biUczSpOpn1eBztKw7KwgLbLWDz97QiX/8n6Lrs6MYrUvKWpSXpicZbtUfXoudSRutOMtW
tsQ3lnkFBtyZik2G4cpSYeIoPLJSV20EsmvJiLMYArb/7VOheS4nJJhXHTUZLykmC5tcijgd55l4
uketCVzncp3LVLJlMCpwvbgBhUqAu0KD7CJJfE+HVB9fWCQ/C80tBoQ9TdphXTqYy0hWTBdd6Olm
HZqODdwSkH+7aBiohcVVlbFEZ7kKZeZNmrZqVH+NMZKH0vX+CvyFn8ZsBNvu9RVIE5IiRRUYDTwk
w8SuzUcMw3QHpMja2c0JR+Sy+Mi+PV7gnNeXybv7wBwe++/cxItFVd5aQQ+eltjpzXd2bHRFzX9+
Zlm+IIutNAqBEsaGZw9c4L2nRFw3IgK1lE2wl6pXMtl5n42MtyXohl4Pj6mJngYda4jnFEk+F7p1
LNaT/Hir3g1rpP70UlbttimaTuzravyMXFU1G/EiWqhMk+ozg0lCUn2E1lGTkP1YdIUPncCmy9e0
Klzzrjq3856UOJ4nwU+3vU+ddj1/9DsNVUvCqacJWWELh/vQ5HQLovDfsJeItQ3ABfkIGGVqBlJY
CukeZZINWKJEST0PUqyixrzqfXilNKEUUtfelu52enCchOiOaCOMXOQkhJvFvmQ0uVJQDikJianp
Dp8WZkdY7j8SoF1rjFY+3UNY2cvy/Zw9b5ej3FQBS6necaphUjO/5K3pKW6ZJeGh8LPf6VIg3/uo
EXDqHwRWA+6SHkRdQWqCqS6Ggd9zLuDY2MhsApDk6L6PA1DCzicSkRA8g0lIOaaIin0b5lPAAh7g
/LiUlDDh0nDGlmCrbzgAH+w9a4uulCEKmuHPyeOPzSLieS0d0s21GBdVWWxC2Dxbb/mFwG/cr0mJ
wZJBWy0YtVXZV61/eOXtkFpiiiGSHa+04hDwcUzyIWJFFhEaHIpmJQjgMwwfdzbmRUyQicQ3DrQ8
0N31l5GuCLLktxrx/aR1qsF+5cULr5VuuQbbiy8eR7UrV4yPXuqgT6H17z+CPGWh5gbfVTInnCu6
zi97Hy5/YEHXiU2Q+3cAgB6Il1Ttm/dD8JHpVCI4W5YaVs1xUWdIHQsG+jDXOoJBBozsSt6e4CvP
5Sf6xH0mHit8bKfkE1K6DxDbpikLqq0l5DmnEGa3ZuZ4yiHsJPrqwEODKgKJOCiqm7g6lAbVhzEw
R5Tr5BtjEj85Zenxtiy7sNRiJVy2E4mdWAT0pK0UWDaS/M2GKse26wtI018rRrCseXAzLigu+lO+
pvwzWuIlxPFOHsniEXcLuzWoUGQqKr/FevNCSscH5Zpv+/IJ19JMlB/SMYbijmQU7lNc/9ajb5Yk
Wr+3sNER8/tT7kW1HjgcbWa8fshbLykYglizG03uvAN+j/OLghqVHKkHuGvX2GFj9r3d8Mg8rCHW
7HJgZUaisaPmQRoIWUPKt7r8cqhegWLAn4RFvF3m6Zb5fxTyQHGekQ/LZuEsF6TYG2MnEhq5sjFl
ILb+rtXC5eSg4XhnIgvTY4WK0X8iwseQIPY/YXsr2MdjHGgPXolq8voFcyosx4CQFrktL13iFN5S
/ghj7M9FIdfM48Pr0/UfWyXOPAAX/ALQMxRfV/w6DaFg9o8pUdbx3NLW5dYauc8pta2ZdeDUnnk/
qvMj8VLEX22+he+tx/SZAoWqahKTlJ4/mgw/lpAH9NQtuv5YUbhyKvBilQVTWbt8tfWhQcBHipHO
TVGxWNBmYSDEylEAASWJxZ2+2+8MWQIfw2ZBheyJvWza1c3lG4Ha2OwqaWkxA0QkgWgJcryAfrRn
6PSCkVjT/dHttUJc4ldjodSlW84vjE/C/4zLaKkyHfL7W0vu4yO1/E/eAyXhJGczW6xveMaGtpeJ
Hb/uU/qkBzGeSdsd4RPnIYBAC38L0qqW5LmeEU6LBqqw4/O3eKxMCXCDf3qRt4StLsZ4aJQl2zIv
boeriiYDNyvBu21hB3arF9om6MSWrhjgjpQjXNVLeWrFtdZFoBmd4kDH03qo1w5TtnNFzeWtPQl/
jTR63NQ9HsjA8+8DchRcXZvrlfrjqofxvy/RO+BckjJVYVCJrHnqCTG/EPcjkSNQYHpzhgGRTty6
Z7qXtAMKZq6iqqpBePYCaKDXeyH/mvDzL6xWKuUBv27fpVhqsFFxz3DQ/i//1EaZ29TCYVn6S7J0
/YGcLWtda0LKEtcSycOB8efaXarJk77V+Hu/4iVEOzVwQTUWHbAcPXonRspEV3z3h33Hcx14vkfG
EUXgD3c+TXQidKckYtxt5kRS3E81oQSvfY3vo196OS66owihb3faG+TeJL7a0KrDt/B6S9NX5v6e
J1FbEqOp3n87//G2H7EOQTCAYBb70DCKNYX4o5MvaE1DwcuBnTO9idmWeNFbLyc31RN6Yq5Nd74k
vooYAeEqlYQPHR3xr2xIBFaLnayKfodBAS8//TA2Cg8nUFHioB5csvI5QtCKtHkwJMh3dH6TBgnZ
inhwufzVsN1uVIHlCasjad4ncLjcNU3Vxw68oiOaZbT20uaknVo9qhBnYya6SKJzsvRJDLhmyFfF
djMVj3TaphhLv4NchSX3p5VOgJwqfYiCAtirkKp7emaOnnlyqBuMg+m5AZHRylYoa8BYkh+ft2vQ
WvvVl2OQsWvZCduVA/RAG/HQzVBpQPOiB9cZCogAX2CvTjSDxHDPfygC2u+Y/eTmw4mgX5NeQyqa
3o1t7C4/Yx5LlIRif+C7S9PAcWWL/OZyGkzcZr/cFRCGl+dCUYDWQXz1lQbrjaSQzTs5BPH2ERCM
09ZkZyBenBb7Dg6b1+Pq9l0/icpuB4dUBh/LCO0xdr88A1+5D3om3YdXPoW99xhhm0ZNfEQ2tEZz
M89Ciyt+3WWLS6ZaugYn3CjYauYoQ3nNujj88FsxhAqKg9G+P6q1YZf0sm3Khx6VuECkPicqSzjD
NWRHq2ML7qiihqzNRj0qMKRStm3uZPjLw5ljXsoA9Tnj6Qjy2Xotyuip9yrIm/W6JgxWGQ0eyYBM
lXLbl6dCwOV5ogHM6AWxyfNaCabD/e9XloUnLB5G6iEI3XUZwiYK3SOII2ls6vQ1cSCBHJXF1MoL
gAyQnIJBAIPJVHYYQs5UMJO+krRY/NdUNn2Qv5sVlQEQNEBrSQ5mNIG4fgMBJEtUqfAhYC4DjtGm
sNmH67nA9OvFfLk/ax7OgG+eQ20zK1Zcd+cntQOVSh9W/72DCvKmgJGm24efDAqtxCnTWlfo/b64
D9+OT1mazfX6uwrBCsGY0WrCwMUaU9AJzDyg+v0/UYV4viOIdyS0h2PQgYIxNyb+JsYsLs9VsTmm
VSziovy/dfs+NwDXaEqG3kMK0vgTJ5PvDk6qjXM9f/BkozpnUFHVwWoa5Eh3OR7Op3yCaygQvB7a
giz1UKW3pHI80m3Sm+qLviDEbgIWaWzoAd14NSa9Rl2sLY3RzEq07RBqm+Q7sM4oidkoch6HoZaz
7NKWv3aaPQlElO3mGG22pH0njS+OHdufCk1RzcmkQHW+sV50wqocucOryUwKlpIHGpE//2bPjlY8
XqzRrX9spVBjM8j8AaY9lM63738uVebkiEosq5laDyIqRqfg5K2LPeTpbR0WF4rrL5sbCT8tVTBL
UUKO+l0d6WOVuMyU6J9fetEJIsNCKgJgSZgoyWx+jvyQHfCrcd66KrnTFC+2nwS+gDXgeKDTTQ6k
AwepnTav3tkaH73SLV20jRsNVWa2eSIKs7aH3roGQRs30WB4AAW1UGCRBVHpuf9VBsOQYbsaOBs2
/8LA/sB+RLM+PSFUaHZXl41qjPhvMzJoflAn3UoFtgzZkBy+JSgKjG2J8GMG990M9NCVCwto3S9e
wutFDnWwsEnzY79ljr8g1CiR9jZXLMpwcWwOcjtEBUGn7g9mqxbJZjNjrPVhP7s8mNs5l4MoDUXc
03ezn82ihmPflsjfudhQK9W0kiqIWzatWTNHWWE5iNkTEemCITsLmgWskG+ZSh7rfc2842r1S55L
FlVl7xta7drVR5s809ZJ0W5e8vNgVCVckpvtFuqKape6VkWM6in/kZFK+oy4VXYDjB9fybd4+28h
X6Y3zGGpDJzki13rdEbh4PkHV2sf8gH+xRI1qF54yTGiypMd3P055Srayu8762edXvRRJkCNM7GW
n2a98B/fgxPO/h0JIa51zhZbwtQHnIu0tFa2Vxun4kgENTZxnbKV+xlAHoj8yzz30FEOf2hBbzua
bvEM1cnHTncQucpfxYzZ9IRti0tujnYzg6d0ryTRHVqYkTrfwVVCh8iAWehb6QODGy0BQajxpO6T
q63mL263n0pFe9hUxyiDZnZUw83BB0q2EvIUIOVZ9odLaAgUqs+TtmQtROomQHYeRvC0NrOrBF4a
g9X+h9YjxnvChjbxDtyHOH/es3B9r2FLtAC7uKuO3NQkoVX3RcJzxAvTGW4q2qj7LHteQjhR69gd
9YWE5yTFvNZRF6oRiqtuSW2zA097UzVFHTJ/xewIRVJvaKgbs78S19zey95ZWMvVfEAs6yX+LWi9
eXnVF9MtzLw1pNeKAK/BkldZs1HFK1X/sA177TYiPgjmdA2Qj8lx5pzsELnF57jVuX1CQjFzhvZ6
8C0RGV2ROs8ndk7tc4K0tNRyB5m+vVS0n997mNQp1mt8bqcoZQGrrOH9ZotXi1hamAbN2Toa2wJD
GOJyPp4K54oXs0HxoA1t4JqDkOc4ViMw1eMBx2+pH1j96oKxjK7quRfUvazkfVbLZZ3zNhFkJI47
7sNm3u7ZxIw9ECT50MZTdLOGU0saliNfzGQ5zoR6SwP/eXnCodA0ai3a0OmYB4b2eaRje0JQWI9x
cf/hYYDO0/GOLJRAGsQgZREFtMpxU24deQkkiUDaAMeUj323vde65/Xv+jHz6DOOcOO7OT4LzWvD
voKDsG1vTepsRp/rtP0Ke9XkHJr4sHgL9iFMqKTEDJwceAVW3cQJZolC6WwdvAfNVUn0HNku4UHd
MPdGMw/aWhArJ2efmI/zFMPCc3km8CgTk7xgue7q4EThfML04gUakK0zTQWENCAl55n478YVe4Do
1lsToDXoDN5yZ4A8ag/hzOzXf3WVPCuJUmzAnlM5VV74fNInk34Z41O5zls7+rD0fG5Yxgi1Idpf
fQsuoPnMdUw4+asIfQCTQhmTWMOF0gmJH1aWJl5XKxZYApSkfCJhmQrQVnBVz0TBurNqV+X6g96I
eaC/R0Ta+T0F2uT8xjimneCQ12jS28tnEGYzM8Ypmv9XaFpgz89y710Rp7AkNf9I+0rJ1NwG7So9
PnArXNSeQcouW3IIX5HnMV/bC3rLHY7Nd/b5E0N3pbfCohG6R44I3sEvOXgSeHDibb3L7Dr6gDF3
sUma7+NvQUR1Ntr2jC52n13qu4iX6Lk5BwKPdp7F/dwWnME+DmqdTggjKYKEZxg5OC1AM0HENcS5
0CFE/cpfrMykfPtP87VGCS0w2khlMmVOWA8PMq1FbfNUCnxgRAABgrLakg521eq6GnRrtxXvhco9
t5l2sVJXLIQllRQFyiD2YJ3VhKbWId+2cjcCttYj9AY0d8yLsFWkPAoefffvlEjoFzT+PJPRIi8f
Po/AonDcwuLE2+y/g/BfgKGwCNraJDgHu6/RgIPpW1eK2BkGSPZnw+PPw2xTXO/CyohQ9CvDYHi8
UdPF6CD4/ibFWi4uHrs7a3m/ZZxdevNbCJVC7DeJoVby2nWat9kdTA2WkdMUbCWZDhAv1/dYJ1BT
9maEP4QxCfDsLfeRPzBzae8i13z6v2L/TLTLrxYWHcBBeHxFuda+khOGPu0l+pPGJxXd+5mVbt4i
ElJ5bsYFHerem9fKyG/d5KJ/PWOnL1yykZGOmxlL8nc4Y/1dFhrKJucUUszpbqYf4kFWUVGA2P3E
rxiH9MA3wq+TGzCtFEXW566feGIXhOFr362cZxbCWlcy6/F6meicgz0JceuLB6FxboyjTYgpUGTY
VE11m1Qhd8l7wrShQDdNCmSBOOmIUhLIoNTFyeBYNHEJg+FHTj+RntUp9lk106wY+8CvS3t7rxEd
gGZX0O+WaWCkPio68iBCj1RnEj0U6mQojW1ZT9HRRZ1RlPbF62seGxldSwLsu0nw3iW+icSpvRP7
xwaWnGE0giVIEVFLGz4/z8bFy4fDSZ4RvrBdzP31y1q+wcNHbrTROFUJeNQ/vD+z8d2LGOV6yRkM
raGyxPdCBRJMqzydULvJz+8z7kuHO7xPEIavnYQxFrSwgXA9iDRs1TePUg2Pkk+gTHrDshI9IcVB
HLcP2wjahXCp/FZIz106ODWJkY+QlliiyDFxnnj9AI+AF5peP5Nc/YN9bxw/kRTmTPdwYeyp7f5E
YJrkLeBkmLdr30QnfaDYbx2wpH4BWlNczNanphXN5s+FtQfmvfrYOTh6uPqHVXWyjr/oncPlO5qF
lJ5tscg/WlXbQBSTiOJGm015b+/Z4Pl6yDd+Te2KssbRFUFjFuwxYC8/ug7kX+GnNhJNGNls3WaT
Z2hfrn/R03Vt2FNw53DJg4xGMjpwU99i4nZNNrPS+gKboxuwLTqbWDoSQVhYni1k6zTz0kvm0dIJ
C+uXFdkx2MRRy4N8jFIDTGiXhGiEIl1BptwrT5M17bQNykpbtaFHkIgI09mbNvaft6neapdL3vAY
Ltf1t5Qu/V06vW1nsmMwykviyDRIoSwW5ivxDTjuAqk6mCVYetwAPcNPYO4T78Ei4TC2kOaaf4Ry
lxmb+MEhnA3RicmyFHErzqEqqwjW2ZucjpJWo3xhhSeF9cOKQWbSBeul2Qi2lsXtMe+xao9tV9v6
K7ZncC5hckvvd/AhEzTamnofoKTvno+wpQc1CDL7pD0bIlGp6Pxu3b1pw7VURTgI+ekyaHB3BWwZ
RlfB2XGTV/HZMUTG7xY1bRLV8v/1mhe0xpF+3G3snWjjwPdvjNp6xd8rZWbxuLckgIsrI+9B+Ry8
fCg4z49wvcTgTY9A9ZuhQVHBXw4CLzeixE4aWMRcOcD22H1e/NZA5Zw1HqAkg2cr+HFqi7NE7wvu
m5iLgYbu8hsx5kNCzAqu7BPtpgDtBuigzhWguCQ64KiqJqBE/z6dijOYOYB+CjA7urzKDN3SKP6W
wJMLlsaQnCGUemRsY27PFUNdljFasfhe67ZCnSYZYp6Ge9IeGm8/aeC967MomaePKvkJMZYz7CKt
YHHOGYVfuKRhtbrjFkKeq5UZdS7VmR8wDvvVrcJowFA6DodaZw7FmU3oVQSIX/CDXP8MsszrpNHy
Re1NQiUR1NZjoJtFS5UsGLQjPtl9dQBm27dL+7NW2cQ2lm+2DyPkzbUsL4PdI5+61Au/pZoHkK64
IZ6JXQQLk2kl631arSrIt9T8y1eOKcaKV9/T2WqGWxmtQn13GZ2nTgMI8EezRvNlv7y69zcP79u+
lCBZH/4D18VLMIm0tQozR2fLbQefxUGisfavqrununYYPljYAF1DZugbwZs5s2m20rEgg7X3JW/7
aers2PuLjCSqe+GanIFWb+P5VJ07+0Y6nMJDiTz1NEAOWFH6kvxv3ARnIZ7wpE35FXoH7wQ6FNKw
PuAb0qvfx09JAzyCVNdhf0RUdtWVhNQyjFCUgdpCqyIipIkOzw8DGwa2RjCov/QLsszbmSNI7Bm/
/UKF7yFEov5nRI3+IWFJagtnqRMueKFBN08mvmr183z9GEh6vv028kicC1Mxe8AueFLsNeYuqz0r
RnAd00/rspouWh0kwpSOyq30KlAVMSCSzJFVNT7YRCeUlW1LJDSfPRTf7HaQqYzYK/cyFI4Q2M5H
2BzdZb6pW67UgGD9sRZfRDsZ5q4ma5KnTTJrWIK4XkVulaiUn4sTp13qdAkukAXfTHA5KSh8vpaU
dtrJTZiHTsnhQV4bBCzD30MCHg+JP70mHs9D1pW5hTOmbGL9E+1tzb5S6556hI8BZGdRbaO9pVGt
YXOILyPhOnF2j96pcmv1CLsYXyFF4Cz8yI0HJEXRi66bv/4VoB+p1REFLgVflGw30xYbLlGvssaS
2MIHCA2H/7JummloXsV/xTRhST7Kx4y+csCHT3GJ/BeX3mnDf8cFfT/2uUP+abMAAZBlpLgvT0EX
afk4gAmFDxeFlyqfuE7tAdNWxTtljwHOOS+ylriH/0eEeE9DFEBgGj3SzACqKHbqGxQwVQAbBmBu
xWbRBRfes0TKxXAiAHeNTLH4+ClirgZPEcWAs/af6VQ4xAqV9i/u5mKa4J6xKuNgL6u5+cVb4fMO
TRn8DphdVGxfR0zC3VYaDvC2dcfqZjZfJJw00+M/WGGzxvvaMkMc6gAWpoCimWhYEHOvR5DUMzlx
6oyQraaQvQnbILMhI0SVwouSqeW4RbK5eLOWHnlC8/I+9ZwQtQnj7a/OG8zUsDSAGOYYtZC7wBKb
M+ZUwzbSw2Pg4jXk2Jp/jz3CaliLlFzTW5RPmkpE8aO79usVIzXQhaawSfxEVCuVfxYnW6oO6Eel
CPcEZntr3O7oNs51foEWkTSKSAxbWOAOfro6tlyNXQeS3gX+aa47JFqFeqQ96zUWDl9Hg7aJoFQm
5Yp7TYH2erQ58S6wU0cNto++c8b1dDnp0mp1XwU2TRw5GNXklCWdNUGee/bjj3kd2TaV1UNwak+A
SvPgUTxWnxOkuoNXBmuIOrvQV05wRk03zLcMK4atD/XZ7LThH3fbTqUe6Uoz7hpUqb26bLY9XbXo
yaQ0herq/THqoHrsIz9ZHCmcNSJY3oeFf4inp5aEg817fRLtOD94QEn7FdHM2w58XUar9O5x6GtS
CEImSa1rnP4VJdQRL0JlX8WfcKqUvzjjubVu1tDyibKgs0hWTq0KPIO5efA3/uZ4CswQ1+l0FuJI
MWft2c5wSz3iJWyXNjtigOyIaDqUWYGFUwwaN5KRnDbo8F98IkfSROQU0QTgGl07DX9DxMjHFavU
5eI1KY32+imaBpi8CwSIJ1I0lJ/6BSbjvwClfBls3gHyeeq9kHa+TjUXaTkoob4pVmCluJqXRtb9
S2C2mAzuM91hDkX5uGFmwWotfyZPsCAtl0y9ZfHabw2e4JCCDgQWlaO353DHU3ftkEXPRHy3efbb
F6nyLFR17tgh1hgygt4hMWFEIvhQWFTR0EZV+N6z5BT+9t97uf8sp0Ttnt+AAzc5fbjdMUlMvf2I
nraIk9Uui3dxQYUfg6c59HkqyREKgRIdVDqoaZN7oFNljGYfCM9Ro6IIfWS4SwOzeN1hpP4UG+md
iGJHNmbb+G14mdkw17kWLuLaecljnEx98ng5v4vehJEiaaHZaRYqTdRd6FCHhHETjAle745Px8Uk
0cokodg94Ts3Gy+cy7xHTxkp2BRtOZWVa1AnAH6Z25RO7aZT5YU+gQGZ3HqKl/sgOyIvhCywusMh
TuGHQ/NToLwmKbxCwTMrLm4ktEvtBUxJHom145Kero9Mok8VFYrjd+4cW4vLWj/ejcYq9Tv9uQxz
/aEciFjSM3W8B7YYpdxR+EthI/J1lLtjr3bk5Koy3q61OKJOKFSpcgmKNknnL6IgBUyh8VPCtf2u
7aRfoPyWQ1FzSE6T73lDuhvnYOBV9AByFx86JOueIrwmIEYN15OdJIqEnl7vG2jh/pO/g+3Nk4zu
6AgkRKBIxJRBgMPgrGbg6liNqIRSSOBSXRU7ErvIq+RvDIf3QmpFtfVpWNYTP8Z4W7WTGFIEKU8g
OTflkv30mNOzj/NSgORxCOadad/aUHwr7bkZOyXG5RG8DhIbCy5RBD0sAC43Pyx/WjiqRg7XUOOL
YN8cyupExwm8IscDp0ybcmADDRjoDj/EfAr6c6nXKG5uM9KXvIgI0lR/X+PDQDKBp63rmENCpt7M
s2TG4t0CZpiNf/pBcnEMcgRzWgMUzVHITS7zJMt4sAXIXPKOyjFU8lq4vtMwr4Q18iIfoTFPpBbQ
u9O2jx6piJ2scuKyzHRFT0BAQk+WSGVlYGMPWZeagMv8jK0FuqSDUgYEe+QAwxugrxuSTXl3W9S/
TCO8PGh7hokXX7yj63KCzfA/0k+R6zzPGOv8yKwMDo61Fy5zC3PRvW4iExh0jNiceTRgAvZ6hPMW
1yopOPte8y6FzVfRE2bFjXRpDgh2XBjGBqso3d6Mp4DhGAeJKsOueS8CwYfHA1eCXm7Mnh82bOQ+
3vpGgMjdAQeunokiE9Fg0zXVeLyZA5vQHFGII7u5rp78Xl9ZWFz1iPJomomfHnE8pZGZkJLBOSey
dazmxhKztkB/apUq3SoRjEpf3g+SDR6f++gV1Pu+ULW5BrdVgIhv/UifqWVf7tgMBOoEg8YPY559
VIdN9vuLoLzzV/h5gkoIAOQxTCmXrL8AKjqzkMJduz7oveQcy4L5Pk8ceTlEDxs2Nd8ZRdyaMxFW
85KFIDtvc27E3jtSrfEv4civErJ/18mmsnVhQvd1qPht8qohQionPxIMRyfQ7WLbBUh1KaZyjDyU
R4RsbpRBfX1uOghj15sW42MvpJjK/5Yz/kFeAdPtgJIvtv0fk/7eeaZ9Uxr20j0CH2uW53bVOTMl
vGaUEk3bmDyHvBcsODFiX9bsRZ+6L+zVj0xUmwxmW6Ch1sX4EcZDztIEBsCX0T/oJIMLuMp/tJHC
y1XLn4Ec8x1InuDZkECn4VRuXbopzeGxTUzq/8oqjhz/3xMFEVT8GXuTAzthe/kwMYTEhX5boJMi
8yvSj7GRLKJfi/htodAUsBChltHJImz8KNOX4dAdGppUhXO9lwuqRolxu0S6Vu5XOdmtn6izEEOj
8b0FzHTZl+AJCanj3/y9hMcA5I42Kc4Panc8llU0YSGbpna3rJwoev9tplX64e0rP7AVAcShje1p
6oupxIHxBMw5gr3a0nyl/BatW8EcJAbtym4nOGuGhopyPv0i4G1UxPL7nhgGYu+2F4cjW707lw6l
J/pAUmaJPCTUXj3DRAGntlhi2R7HkQXis9DC/xWAAi7H75qhRWAyWoumZa9o2Foyj8HU3xr1d16v
GfUmBNYASJnZ64WjjfJ7bowwj/PRea6htYQVA8S3vLsw2ck3nZS1EpqI8uYT1dGQ3sGFT32QyuAN
wWYGLHwLgV1/O+Hpu5jGQ+1E+dabX8y72zIDpWJ99mrI13MuIouJn3L7o2Tlwc7+bVxgqQhQtaqx
sUm5aN5+g8NKA/vtqS1P83UVWDvb9UKpcP+zyjHu0xwDFnrCGX9l40iGW/44BElSOC1XlIPUsLM8
f5esFhcPdODWWxYfE0pVCoPvjVXD9/gclP5+ow+G7FsZVfwde3ibMeb0hg6u71RUvCTzgOFUuaWd
x2Osm134YnUhWtd2ZvfqG59G1xtRj4m5P+Wt9l2kE0ue/TtF/FeZofqNoi6+BmZHwDyLScjz5wmT
NnSo3TQNvIGFeEWGf0fVxNS/kHhmW3bWvOUTKial1eX9TY9w0ZWk+aJ4XLaYP2Zv55b16Whp2eOA
Mb41hzC0/Iy7SAXPdwPnQcaHE5mIeyCoLovF7ys20QhB8m4WH2V/t7TJXHgYbTwGvKDRn2u6iGh5
EY2Qa5rIwZVh+8Ou3MVZQG3Ad6bqUHS5qP8rrKbvyOL6xqsNxBXQs29fTmtjVjj73rcmViPKhlnl
s+Z3AovNfSqByuc5QRDmzM0LcXa2iqBBLXldYr4+TR2QWD6/oUu3dvi4Rdp/6UZ2qVrthvPljloF
p+qYMOToCBjU5Q8Esf1JFoRQOMsKikJBOa/9S9i2DOZCb66sooGnub8ePdA1OmClzMCVPS6XwFxG
fzLEt/TZHbAMdS2hO8xOi3jH9POnnDNCzdaYQPhP8Fk2d64Wx8qg0+0gjOkuL51yfrGmq3mmjRIb
BP/LtQYYpEXy7vIO9Oh6Q3ESgM7Mvl4lw38hrPDGeoONphMVvIc4CrKjzNMxVIYxlDa4LiWttpAS
XbXJ2nEAEKh5plf0Thi/VJT2k5scQq5DeOD5ZixEb7fzmAWL9zxG8YSpaaM4Gy8AOAKSzJLOQMLc
KK83aGueICtZKMbPwmlDbsh2AxT+gc3TcEs/hqPZvWfjkpJo6Kkd+IhSwE0Td1bs/2ui+Jj1nWvY
dAJrxFUX0zFw2x/wzSah01b5i3BjpnCHpEVKLU0uLqxNL1rhDGaKc6zXvO2xzSg2+WwU4fpTkRG2
qHuGBLryB+vW182qGDBohbHmx5i0mT8RPxxO5F6+LgSn8kWXatLk4idNCh5bAbL1Add3ifzYXaD9
7/xxSVbWmsC/wpNVG7sg1ZgG83rWYM1spEr+V+v4QIScJqTdrdAv/faS2pB3VmvpbCAip35P7EFW
+wutacTLQRYMF8DTNmw7GqdHwq6culhGxNT0UuRm12fFI9XrU2eR+vbAzzZZQe02w3xIwOqcBQDM
1/Y2s2AEG+j9ZsZi7aTsBKIfGPAumjp/JJ/Iip6wodd8P6/FdaAqz486gBpXFnmAdDVWRR7VxnKB
zvcg/qK/y26pfdiutXh4JwbSq2kEUbmWDE1S2kla+QFqZSXAkfbiIxfqY9kAkhhb0rIMo/HwbJWu
XOpiZDAtunJ0ve0BWfEHOc1JhWBzUFPaa9AsFJaCw+zJmP/CpZnuuS9NehAToTXCHMkPolhX123O
J+GdHQTy8vt3KoWLFLyqVSyTmmZffOHk1FfaNeloqCZt5sSQbqOWFqqPnujl2tbqrjPZz9EG+Ul4
P/yiveL5qq602CFChAUSeesdzViaEKH+GjDP/G5yhsgwshQq1a6P+yc/s76yaFwEtlqh4+RN04pq
aK/p1NbP+ujzEuV3lD9BbQx0lBJGARwBp8ja5E+PlqPld5Q/V0//11kCnRiIi2QZ2JqOhuuYlOEx
oWl1WnTdzVeV0B2epS2uWFPq4Twj5NQv2rCJQvBUrogjUWmk3ZO9wznP/ls+5muJQwRB+khUJy1+
KdYdCKXKrmqhQqfCVFSyDMllHs/WLZ8RLHpcf29zDRkVmizCoBOEnQvZe5EWkC/4Vvx4xnbq0E1T
T/7YIF8LqZ5csiBSKaYC9JjV+CDW5XvsMzmi7Yx/Kg/XUinQP4uipw8smNoPgL62r2b+076M72kL
SeEET0SDevysvohYymVV6e7+z7mcbN1vpsDjy0MyKDekG5gh1RV5Xm/Z1b7SuWe+uHRhKvwQbgiV
WuHoJWwE8TPvQ0NbS8DMUFTWtLRR4Gch3ZB/GwXq+lCN7Y+5cpk7B4DDDDFlcFsfzePA+C/Cdj5f
LvLHwvI9Yn8zGqgG4rKx0ycigzS5wSTlkyhujOb9Hk8im1rO0Hn6i0oGwVfWyphLFA7ss311fk7i
kT6uFSXC4swUOnYoCR+zVI7p7MyWW79MONhdcT2z1qJ2ne4r4pEXo8QX80srT4HPDQFMv20n5kKC
FuoLSlGGPSfA7/CNMSWqmgKKLAK5+ZvGwqjBN6a/t+1sBUr1IboO+jRBX4/QPGSzTEe1L+i9ZeLt
9J1pm2EUtIr/AvjjaOWJbrO9hfz8a+DEFzdV28oWNK7HZmHTEwIM2gRIvmhXmgkMuZAcBSAUjUPH
urRjMSIc61eRTHxuzPeSdDusiYxgAS72exQ2dIw+fKaXNL3jqhcmbNRy5Dgd3NLdV0CYZY5NJmf6
0fGcMkiJaemz8Xif78uxYAwxisUn1/IiVmOaZbiBWJOq7nuG2fJT2AmTE5PvaGSv5unGr2eYesIy
93w7CEKV1dAcTAlZS4D78aSuX0PXcsSiXeW8VDu9pHIzVIzQ4F/YNyCUrIqlOakr/rSBO7IZJamC
rl6sSgCTceh+XBltuUvg4tqSj6Q1txyim8loO6g3+5cD4MVi1u4+0U3oN1nzE+OzWRB2wMqAVbrt
+0DfMRVRlNtY2gEGFyRJitPBAgWANxJRx1u66OTCHEh9KMV9E8E/huNe6v1jNN+xigJKFk5sui9a
X5DBC5lDP263JnMsZ1rY/L9JiMAwjLgYTDNAfHePXADtpeUIVG5EeYfBhK3DDYWbcD8lcwr6jFyU
axskj9ZY0EjLHvqtHwIRa5yyKGgx1gKuUMCjxXKZq7Y81EYY/cD5lfs2c/qv8TXci0wGAnW6KaLs
7OcqcpUyc3YYWDHS304zeU83zNkrFw6hflDVrFhuIgBPFX8IffUDPdcsGULO1Wz9nr8+iaStkCbA
J/RaEimGMl0adUbwJ6SXIuLyys3lcykoy2tczSrvXCYmgtW/t7tQJo6Ov/VXeRTqyiDdEajDiE99
RiI0xcV/59s2oy8Rrw85kmg2MpSdUp3P3aPWTldJfAX827W67RjjIvFkIy2erZoVLlUGyZeQrh4h
UKXVaQ4TRbm2KCQ0XWml6CvwtuViHhFHy+qwuvF9P8zlFhd9w1rG0huUFkM5WNaHVHwH7IeKgLYJ
Tx+sHTIADIxTApK+LTeq2JIQtw4o2BaSIgQDPP0E+r3f2jT5nO1/Uw/ImOf6UVLV+B9ab3br+V6a
fTKqWQ/eh6sLPlhSvI6ERJoDyHOWZSFeznJroGZYIcDhVoiSJStC1BMqgOBFvi5A0rNAjro19cr2
6YPD3VtTNMGiHqc7ZX0dH+lsEt+VUmkQKwcLr+pKOIDoYXbFYXAwb6mJU/kPKrSLEgQDO6aVFfIp
Hnxu20A6OubduiTmluqzApeKQF1BTlmmERgXYMt9wA4PNeStl5sxN2KqWQxZXxKzXEbR+u6jPwlW
N0MLvcE2if1OMYsz/WKuWwra6Pf3LRJU4sP3ThU44Fs1gv0fPn2S3IRwvje6gWrGIkoKpQrN7HOq
SdeIaLqrsyFLQFdZbMkJBwIeNno4HvQSncZaLmNWYCIfvQ/amEaWpzZTP/GISgW/fjS5DxyaDbNB
2T77MwcSCd3zqJHw/pcve4dXRxvHq1tj9Cu825QFE0yYSzV+43XfUVkeJF12S3pSUH13B0qm5W8o
M8d9jd9WbMXvXcMEhJqmtRtTN//MB+9p3mprD2jZkeGnCdjnvj8OjUprTFSdh9enOTt6xa5CILKA
SUIQ2D3MLjEdEutx6VsBZcUgq520lfA3sfcZ9VezY9qMrYuoFnKAMwxlXGreggWpQSUkx0biR2dI
kfNNlAewgHfiMJWv5zXg28HuXR3TlwvZMjgQjhqQLXqrxkrG9HmioiWFkSN86dh/y9Iujufy6CDs
oGHsLs0nKsQr0Ux7EqyhvRl71mP7aHUJco74UNNYewx1JBCpIijnFoUrRFj3gkNuByyLKxMEhL6v
gUs/XZCiy6vp1iPfz8bwpBIuZFa5XOGeosdMGEgJyRk8RJBCONpIRekncUZwdnDWZRY/wM3s9Dec
t83eEHODdoFxBr/aS0v+8gilpT4fv+Bdh9+mIRRfxgkohBCuDF5cUxybtB0VFC48gC6/k1fp9Uwi
XSzTTaZI0uJoa2lJpyrUwbfq2lsXSSZRLk2pJDkf5nngEFNSHOnYO6Yg5jTwNpnuzU3KxI7kZvUr
6aLrvQip3InqGC7RhEBgmTqLuj2BcmBCOTp90U/talzGdhgHT1XjBhYGxiGpCOyMtEaJcDJDjSrb
zl6ja0s6Q1YVvFChROFvsSj5Wnxwl7jD6OcAyWH4QyZ0Jil8VAs5jlOqJGbTpDH3NC+5wYdckflT
kt6ycgAUuX+lIDiy0NiDZuIX+lJhTCVZFQb6Ty/xEJs0PWpiijfsnVtGVT9YNRPFtEIR9xf9dyJf
nIFNblPjAX9JWWRnEktcBibtDQ0dyVr44tdCj4XJR3tMNW1Le4pQBYHfayguyFQCUAnDE6mSSFZG
N6M4wWnVMQGLzK9cafehGWQO9N4YxFjxHSJZSYVd7kpnyD4gl3ulSA/AAbsF8sJrG1gaBOc4UEja
mlCuZh6vkwlYiVqNUeCvPJf2JZehi0Ldv1lsuT4dTKdQAeKanAInDGFxzgtdiK0Ykl9PGMS9WvJz
yJUc4dkYDv2F14VXiULzo7DWXEeru67GQG/SW9LwCcJtG5glvP9iotYHF0nuI2qe2mNnfd5XSnP8
7e123dvGf9lPcTBflyPcTcXBDsK7FuUgztPIcURM+kQ7I0FF8r+9UGU8+P+OOY/lyggh7l1QFYQw
A677SJjMOZ/UV6KiWU8Dtqz0cmeU9oWSag+yt1YYyazWl658ckRo6j9IRaUh/ppjhHVRKZvK4x3g
uOBOvcTNWpU8rgBVGMx/AzWpj2eSzMjN6ut8vdx8gIQERJ9gKIEResb2ogHhTyliaWMcOrz98K61
mAnr5WHlGW7WuNuv+MtZdocS1YcX/zsVeZ5SvgaRIXf9jk+4g348brPZJ66gDYAYCZ7LZFuZbCpj
mEzQzC+Cm1vxTgTHWsTEPWp/gEvffIlHhUZtV3i7YlqiIWjSyODj+RWeBAxk+9J24M3rzEspyO3f
A1LCCvVOmmT5Gdn6GCwOPSCHb0kgN9vDYLzfXOnErqqmB9mRttgKlY8G/JarHb5gtoNzvR/ZE7Z3
NxE36RaiFB0FTVA33J05Ohy1wdiFffAd5NlYamNdU367t0HBVouxARCi3qsP3rucyaBvE+mnyPDf
dN0qJwjVQWqu126eoHfNC/zvVXzSIaCEc18k9EmYAi1p4mXD/6kOORQ0EVm5hxCl+vPXTa7zanA9
d/uPFovjCfq210pDrV14raBRrc7RGDVb3vAIpqtGAut8SplpmwpaFKTc5laZ12o/a8S4X+LdGHXf
4FFO7MOMItTWOvry7nwcnMRaNF6EGyI2z/Ki8N5mYP9QTu6zzrmpTTUVmp9OJfPWtg5VcdBnd1uI
ZTe7u2ReZM+opTZpaRlgGqLO9Y+AOPpj3aimea1FxrBCsfGOYjzmuiZRyp1+yHIDXDfJ8pvNB0gP
xQK2uVvb+XAHfNdunvt/GHlgcgXs9ZUXsgnReGHVc2n6wUZLOqGl9hUF5baWrUEbpXUPNRM1Ppr/
sXcZPJSxjCDVkIIa9Ik1YI5OomDGR50t23bXHAEC1zOnlFr0J+4GqEIZRFJ+oLsa/Ajqp9c9xhyd
uxtE2CGj4UQZ6CP3aI5FyZSrHzItunZ3SNHU5RNqVGHNq0goY5bya1lOsisFI4LENR/SSgwG5pZq
crbzHijJ+fcgk2V4feXwAgArX3DKqCE3VaTSLFDvC2O5hgLJNlKZf2PkVk2H+sNHW6NgLcRBKb3x
Pt41UV/YyspQMOSUTmz61iLogrjECFkeRO7ejB3/LKMcmROrZlM5usWvGO2wBoyqVtt2kcuYQzkp
w1rMcK7w3k6Y4gfzdaKsSIO/l+kJQwk1zgmTuJdOd3WQ/v/6Zndra4W58sT2IPCTjIM/Y2rcoNZr
zx2nprrg2Z35zQnS6b8SVdkvNHggYpQf49Q854n4Ob38GI6u6Kd5s2ZGKwOUy4Cr9FPnxAQJIq6X
6Zk9NgQXmFWmVwmeTQB7SjuOBFe0pw+ezyCjrpv1v/5fHc6l6jqypjP1NTPw67q9GTP0zHkEHoGG
A4SGw++0L6qIBo6wO9JP5Nr+hZCuP49wdPWxklc2eI6OqJ3hrR0zhhtgLSQprZAWmv9DEUKjyAUa
eTWlTHz1uS39ZdobKbR4e9bZw0mjXhLhb/kc40KtjIJX9PeLPksDA2s5R6pt9p7vjKAD8aoo4QdX
6E2yjIAiVe3vezFNiH/htEtsgpAlD2yWDfFlGM71WGmQAd1ZcucCwsXcz3TgMyxJ5IYkx0SZuE3G
QuNZf7vW963h0NL+2Hou2oqhZ3ID1zFvRVJyeRdzbXFLTklN9GWDblVNfa9IYR5LCZ5/OSYyWQIq
IV7Z+7Dl9ZIUyRSSZ0Y92YKZA7x1pT6QkFZJ26r4m0JAzN7IKEd7ZPKHMAtbvsLDTw30gHU+06HP
La9o81GgNdLS1Fr64sSuZadRBu9DY02NVgIx99b6cE15z3+WUUR76AfzUNnSN4IXldxMyvKHrvJO
bRKt6rqVgbX1gy4ep0hkcCVYDtQ5Z7JEqEz/em9fFeSjsSMnpzllTwKaIvCX4ItWDilF4NJMOBZx
WaUqft5S7pYaBZBm/4W8GIVbm4R5zQIzbpuy4hjkNL6W3UAeu3n2vgRSN2P++8ufQpbVfLpJk9oC
uMRk9U1yp8OEfHqSRjwmdPe7KrndjHe+mswJg6h3EjhUHFbsRtN8QJ8z8sZBCRmW7tZNMXGSJckK
vFsig9CygYffSnwaNXAQsH6jzB6Me22gD4mURh4NfKhDMxdM8fT3tszpzzE36YEcgfulzuSrDcez
X8OOqlmrT+gm4tkFFaaIBp8QYJ0uPb3AYQ9ZOzFOezzkDVLh/mG5icIkpwbO5Da2mZI/FnEh7Or6
m9kCWY6zo5VopqvtykQOBhYSiDnMIl29+BsP2E5Jqum6N+ozrS6raPFs+oUXuTJNPdpxpAekhGTW
cYD4AHP3jwM/+tFhDySCDVV4b3DqiiCjAuenCic9fVh8+x9Xe6q8u+V1W1kbEvm6UYBNyJc9po2s
PY47fiDTV6JheDrr9vRisL4ZxpeyGWsODxZhk/7fhPv7k8Qk9uT5fdbus4/pDTSMeusi+riSsq+C
FbY6AehOzTwRAF0SYlQFnNtVhIHhSHYRBuBw8S+1KJWQPLS8V0Xc131GnKvLuOoEySMTK+rHN0p+
MA34GwjSWIgegjK/t35sYlQ3FcRk5a1XGsPjIruYqsraoPyEYc1xxnLF2r/HwHfYIyQcpvDhEtLK
urS5700KiCD+ftamI8z6wsHggFQ0kqrqir+TzQnXGpzcvJQ22gt8qYTYdDJpiUbV9WB2iOtZjExY
yWQaDjoYx072nJmkj2AbWM2E/kiGfH0gfAK9uw3Q/4pDe5UXBShdsm9dBUZ1Sur+7yDlBli4rliq
gixSLhI5HRNaRKlgwy9PkmXcc2zimqosVwvIz3rvI5cLjy6Gh5lDCyJ6nRimtmO2iAG7tQap1K4h
EHYHvb3Z6MQYudu0a2HkBB4RD2EZhsNu1olb5luqLwFXvLxZ/gZbczhb4oT9ii8m5ptIFAUelA6w
FZt5DYsONJ4tr0lmnYBeK+g5FaOj0/N2LZwqraiuwUmfhP2tgKrSKC5a2hQf64Wl3FXZ0nrUs/Eh
iMM1j5aF8lp5V+3RFJ9VlXA6SV9agqPTjkxw4LzWHi70V+90Q2lgLCtoGu3pAsNqJo6Uc98UUZnW
WSWQ36Ix52uw7kRpgMpCRJO0EqGhvnAGrzn6T2eYRas16muiDVrcaiMkP4iwEpdI0QlY2Y6fWU5/
Jqlpsu++8JSqXlTqMnqWoD0QjmWrZBUcDRaqNakhHcAs52tMsAUhm44v9tTlMD9+to+iX3Weja2j
8Mf7V6jPnTX1fMeHIoDRl+4nc6YjtcNxH+e9ujHlhFbGTs/Zyf0HTWRObstcNUaGgQz40LtNUxm+
KTGAPtCm+nuUESyE5iv3olCl9SxfkfLF20ocWN/hldP3+Pzzo74FRZFQYBy12Ij1FB6YPkcLExqd
hW8+SwSH56eIAFOSMU1AAZjWxolpjCpyEjRWAgmuQIBH6EwwCY29uoCoGDWRPSr6BmkKRu2GUB9R
cb3cdCEoJzKSFi7eYd4WmBObwSJeblk/ACM5pCyEhLMuLRo9SGkAXZbDOA7gEIdZL/8oj9YZKXCY
M1XksYkjNvKjZEE/Xai81N0fA7+od6+EpSjzIuAfZCs/PDLb4X+S/gBrHF3MPeMk+O2g+JTWjUU1
BtapLo+33vEt1HOnq/nVqCImfOf+KxYdkdQNaWYmgSAw1C7TFTi0ANSXQHQSLMInKC/umMIazx1g
0109eOYXf6WU6uux3uJk6vQBaLapAvhvM2NNAuzbsLR8Bfy/wcyZR/5Fr3GJbQ6UnXT3IMsunEtY
TPfLgFjDwdSMuJGEzwen/yp0PUQ9hhDZlaawpSjJKfOeGod06TE8dUk8g4lFZ8B+OE2ebB7ajlHK
jtbjqQDRoM2scW4b1fgwqrq6bS2PeI4M7tDN/mLcEPPP9Nwiys1ihrjUcOSzcrpaVi4+QxFKalzz
OKv4oJGXeyGKbGvRqra7aH9llo+N2TcZOnJsfaQ77HLcy589GPes7gVsaC56pewxwGi2w35buZ2M
v8DmCxNsXApJw6m3GHjE17r9e9ditYsLjfAQkEidq9/FknaUnwRurcweLURfX4TM5t3zkkWmg4is
vzDcaiTn4XxFHGlofIB9FNbBI4HMksCC/f4R+ZooyokAizyzn1pDRyN+EQ0SfBTWFmJYAtH+O0Dr
XaPEIESgyuDZPQNU2ake5qbFisGH/DSqa6sxJaTfdWqbBwULvIIYubFw5xNusb1QjF8RL3jt262F
6B7Mi4h632ts/536WvI2SRp1r2d943Gcgj9PIeASTw25okgwiuEs6O+DfM9V6eHh9/rHTMRK775i
fMpl6cPG+8ALivWxV53AWUVjRWK0ERIHU5/371WrY7rSKCg+kOAnrDkMkmXs7NzV7cE444NmLXi9
WijyTBRSlS3QeDJeYdyqH9M1AzLnZ6ionM343+MY2gu9D/3MpZwZu1e/DRuyIUEBLJAomX4n8Qle
iXJW6IC/lCsJijEBWOrfPZDSyz7m4AS2ILv7l8/MeZQqZtVdeBkW03/oW3CVRDAhk+n+tJBgDAZg
bBP+9cwPm5FCZk1vupkSYxjTX1SOT6lFB7MYhWLhUOqXxHMpSFNtopwRtT2mHwdcwDn+GzxuOq9z
sxaKSNm6Wfak/OCkwA2jT9Kp7tJFoBTmZ2VMTIecgL5skstfNssGxMZSCzt5nJr5UK/1UjpgnRa/
hxHQqXcPjy/qB2ip8jYWmI51FSPQzOaaeeRtLzAcRm74aKWv0JNjBRpZUUQbA6A40jV7VDH9IogE
d7P0Z2a13GEhEcxLcA/1tnJremj8jsI8uwjnn1SFzQXgECkeBzFhypmK3Sn27Bo6ncaSTYNIORhO
dXKHp2wlAsyesuULrrnGgLD5y/uC8yNJxNHPbeDfQwadZjjxLUMSkJTDhujwSZXnxUr/p6W2PL8h
QvFexZpAymciDdFdNRkHSoIKqQtxvnEDZEPEpsK66uAz+lLX05vFcei1k8zPgX+J933fS5+qX3DQ
MiNLracl3i3RbZ7ORfcmjmRaZTYvSSI/18MiwvgpLBStHhT0wTqHu6TN1PDg87DFOkepjcZnNQ35
WHKEvOyOD1xUdTh15Qgnz+n6TPmt0eXZkWx1641tCNpbhHJ3N8UtrE8woQft0htA2n9SG5Q7L/68
+RqaMDeZ7uaHyTnYwtUxs/roX6c+VOzhVsYvYRvJn1eIvvvlWEyvovrtHAlMuefooClAOckAENAG
XckqNnvFV35LtqZep2KCWvUJS0FH8WiTUGabzFA9kx5B8CRE/Wpxe9si2y5Qsm2uShnoCcP2ccKn
+p/8mMEuvFVRy9bR4Hrkw/BgHx/Jyf9Qr3fGRp+IlrRTivy/rmyshScIkAcRsRS/YpE+dxUMnSwM
fgD9BsSlfbsgDri2xyqncmY9XyVskGLr3GGAxXHfyAynYs+oiAyz7Ex2D2pSvVr9tUm/6qMEulbf
epbq8OHRugT5Id9EnC4pTs065vtymfknaRJpB1bze+hD4OPcRHJKlOOTugRVq4AuZs2S0Eap2k+a
bez/ZsdaVhIVjXbhVQAySB6Wrzuz1tDTBWsZEAu/s+J22nRl4t6WQnXml9FhavnhLh9ua3fWVPdz
qLAIAOxlcR/PAd3ZjJ5pnSQbvGQk2zB5JaC88L0fLVa9V5wTyLOOa/QOFUl4QgcyigIcCDticMQz
uQdoY1o4UIHoRqas6Fagf06VbWDVLMW541isnT79zfbqJVVwWxybt8stuDK4at3Mkekqjhit9osM
PUYDPZyAoktpoTSxN51lhWymb1gaH1asoyTGvSu+XzHGNOiqWPln6FwPh4KYFDatPDpL/U6PUa4c
YAy1UDwBo2KB91LrotzicOL2kfhCRTXT8R+lWn/rRIkkY5KZA+4ByW2TMOjU+A5R4yPibrzEH/Yf
6XWLpDig/hkMtwLJqzv7RM269KA+C0ZXfdJlLIb4DUncKML5G/DscthSpsULyVdpkczkD6pDARVk
uphTOVfIUvx0YQCxujYS1OA7LM309o68zJL+FfbBh/fJ1ZzYA233s5/pUOmDocMkzMNT8uQZvhcd
EyI5fsvMjv2tqT0p1F3bwJyhSPJUhRb6FhDNIW1PpEtsqEuNqvgbFYsM5QioZwID0SEawf9PoIlY
z0WbEdwNpPbBed4BnLs5/6EqEj9K8mqW9AYQMQTN9CRsQcdL4+z9KSBl0mQD8d5DDsb3AgPRgS79
v3o8cZ0RlfEpShZYrQ7qUDBJ4OgZW/pktq74J63USzIbqsx1+xOwBHp6ws2amLuTRjRAVcem6Iwd
kyHsJ3l0YwihT9ATC6f4Gu7cI0kQ3LI7lERZNznVcQsMQE2N3LoTf5rjJP9bYa2utVfGf9kOdKLQ
ndbJyiUm4oEr2HeLTn7r2wXEer0feJQetpdWMsqwqwb/SuQe/wn308j9/Gj5eL84DNSPPGn8DK0f
9IZM7/wOjmeyJsVXLP/Nd8osmn4zLSyZLZDT0nLwYuMEPTL+ikl9HqZ5L3uHsxSM+HmrJE6KM5GC
tpsQN7Vy4sA6WIN3AFpqAg+wlNPa22dfHsi/UKeYFHdiwSnOO8NOfM8jsDe9eB3J7SNvIs8CQpv7
ov+OStEFlCOzK8q8L/nAGNnJDy2uu0ETt4K3Shfzr8MCXt7ALKw3H+A7yMeP7jXwFnnyIWu7dATV
erb6oNvf1JIho37Ue7cCaOQkPHPnqconrqDpA6jh8tRI8O2ilaBn3Pq8YVGG09wfXDsq+5YYpG1r
7yBRGTNX7rJ8tWZVmI9v4A0tZIWS5dtfLF9cueR5flK7dnHGpVL8l7bQDFPHL2AAyWxD48elQzTF
OXzX7VYu2FPjFX21vAkgnRMWE7e7Q1Vj5k7aVwtOSaKCaosiD3VC8nfboRfNIXmXK+WnIMZ6znLj
C7HCK9DJFdeuK6PIcF+GzrAuMq7dJEjsUGklgwcuMbK8XivV+OwtskC59euhaln8xZiYP6mWjeRZ
yo7FenG74Hm+aq0mWv3Mp1jHF9lkPdjxHTywfK1iIJSrsLqOMZ9TCfh4wD/3+YwBAWuWzJp4+G5B
691M+65BHp0UToELl9dzMm5YCB1+KCbmwDbZbj3B3qeEQ76qSpYQgU2K2ARocIQjNSAeIJ9yWZlk
2rutqY2g604eNJgs/Zox3e9G5wh0Xs83W0Sz87GudSJO+S9KJ90ObIF0enzGM2IFdsJ2k9feuABh
PG5ONqBc0foOOVKJI+/+ghBaqH1vJR/cGfuAVRh6Bt/eqIOVrqKR4+lWym+KKVz1/bDVwESkUfNT
MTgbLvlBU3nEFxxyDnUc+WGDwpmgNxI9Xd7kMVcU59XcoaEG8z3VJYUCq0yYyV/lOG+bVJjIz3SE
ACLMCPCJyUWreOIO8Y7R0gKRo+JGA7aiw1rArSYYYvYlZaL+jvfjAxON9IIu0HHVJsu1gYKQoKyZ
uanBgMrOB0+oJQwNjK074I5gkf8fbts2K9pMp7gvnw9Bp5pBXDuAcbhEZBH3nR5bnXes2R2W8mHh
HR/jdtIkD9PDIxEx7WFPaKzvWAughUD6b9gXK9XfAwUjOXufAqfkxPprX7TdiSRnUHiY6cR/BpBW
+0a991PH1mvv1FeWavGg4Nsld8xiVchqteUPkSaffdvidijY+UQ2EPL4FuV8hSJN+WhQlkX+rjTy
io4f+CDxCcd78YEZSV2u1YvuA7asB79X8ijPlGn2594NBJFLadMCQ8d1G5Lu1P8F3JSTqqFlXeFX
jKvkooyqW8ky0BME3PC3sxbhzkEzYi61ICzFAQIx0xs0flWKFfOtdnt9NnQLe0lVBgj1WH2pwU15
r8K59Ik0Haa79rVJg/+YWx/sNovo/H2xOoqUFKc1xz7hsZdXhQitXSze/Z2iBWEHJwqo9T7fTC9h
QPfaGqAdCs17765+qbYxw337Uh9V0o1EVbL/ki8/hvdU8KrswJslteBt6gj2xN7hJmVSjyDD66jq
cstpf9Riz2IIUrzoohyFUxt3KxNrjakijhoIzy/+mn4HSvcyo4eZ23MLGyMDD7l9l3hwzr0mqucy
mwDircKO8aPV15Py9FwF9oDpslniIhfF/Bc52csjaSX3E5VxgSRWeUZUWOC77kIODm9v7UOR2+Y/
/TyfsXrgwLlPipIfT0gYcwouIrY3EcS1hDQ1HOnF2DuEepOtc10iXXZdiaUYorNCmHagNf3qdoCr
01XR+msyRrBLOdOofxssnMy3IUuA4w7iiebekQG3MLsRoY7D6vdp58HxjwXjdFv3tCIVfHNJSrRG
p3swPDrOVpeNnELQCEClCj/5ksZrz82/UmBwhkZ6EIKH5ffiepL/8eiQ8YI/08eO7Vcjs/5EB+su
yQi8xlTwGlRtAcsxkQzYzK4yfOk1gTDiW5VxzoW+1rHmhJCfYbNYT0iB1wfckwWkyEXPIx5KShwQ
dQHW/D7mMoiLUVTTzbJqZlYFFnpqmcPBo3FhkgNVo03GIMX1AqoHY1zXbe+BcqAho1lmu61IV10G
CZUUEqE4TKIe/MFhb5DNshGzGJb+nhrCeeO6yMyNO9wU+FsbJ6p86UKwrs9apf/1yfSidC3BA3Ev
FKTZCX9dX6j0r5hhHhgf6QOCRUfCQSDGOPA9R1wbqx1rgM73kcsWSJRnpMNIrHoYABu2MHYoY5I8
zL0CLdfM4uCkQxJxkMAMFtxyc5i3zzYEi7GJHooCNC/fNMk9T7Rwy5Z8myykpZv6laHY9mJLfLE9
obSr7kTCas9DHmY5nmexuOUrCxiJ7azhn8PQhEyI6E+D0Q/tUhvZ9l6FGqw0rpfNO83raamQSST7
yQQJdOjrCsqQEe9lBUrIQtKx+vOvWdG8OX0vLZyHSKDkSri9RqKI4k4WhWtQ6aRVCqkJiwtq7FbW
IpzlEpDCXHpOY3iy5fqHABlhSdp9mz+WAL+QPKrZPoKzrJ7n8u5i+qBgwzWDJdLHPwM50OnPnwKd
gy0mOmneoaI3HLbNc7g77bWo6fg/GKvn3tAbwqKZ6FdGpXXHy78SQlw18ZpvYUs6OKahsj8sm4fl
PnAIXUIiIp3sS4mFBtom5bo98hyVqZuQCrRtf+T4x9HYxDs6AVmBIATNmVj1sNrWgEWJNGOk5aBg
KlsamqSCaBQWlVAktFjZkG5vJNemn0zUL/16foz1+IkocS/lT9Yp/ZuKmOTXmiGWhOsnu061PVol
85ewLm0gP2rWDq4oHQtenhAW50p2eQaORZ+1F12gzcNyBSG187yEd8HEOUPD+Ck7tXDBITAd4+DA
YDlYmkm77nLgqUxxfdNszHzXllGdVf5RzlKCPAPeebLlV2sqjYE1wWZOGsn5mHvp0WRx9NBZASRT
jtdSezV7RVnh+nJ619vpiFnVEB4/pQFPgtmSCwZuZCqFRlBDuHKrXcE4ZX0TRCdSVke4J6oXNkxy
/WqgHzdQAC5LGasoHVP9A/NwwTChzDaL2GutLibutc1hlTKdLnfPv8GfhFGISpbb8ztuJCGiPkqj
1cdktpS7qiMYMhisxPdXSeJOSdSS78nDWRbUmstxn10JZSE7+z0wigXJ+l4hq46D7OBsUgsBBNcc
wnLlEGaOoV8IR7z5runL5Ccv1N1BvzPrp/fGbizKGW1HW+Ct54SSh2EzsoPWiLJjAuYCCKQ6+Bfo
b8a3HcowKZsQuv+C/bqaeWwad+Wwo+KLIFR8FCth2wfuW52zIEDhWX5MGGU9EOimJkLKDPkDzmA6
aPRrA2d+mrM5jvL4HebAgA5kJtEThaJMdSHBicT70TvfT/ndaN1Nzx50AQoC4eYevpzwbSo91G8W
Z0UBMkXvCWH3nYwsLSjqOD7L7BOoqhj4NmUuiTpKlEuCIgeplnM2QvXlb6xg9RvRP6Oi7E/xPhvl
xGz142Ro3i+ZaaCWYtbHz9g+DX2amgD1ozushAQQl5dMHm6FFJ2UfL57iLmlH4x0L5C+A5dn9gmI
O1HKrpIewm3NCGyvE5OaPaOH1NrUAHfo5X8vuL1u+eFu8XAiRRxv8E+usT3wXU7tTMWwaT1fTK5e
VnewjKliAhxJ0eElp+4lIDnSLLjxnE4efrp4LdqfJfUnq3lHjeO3eW4AcXmndb0YGfB0zgVWQJOG
Rg0bEOaskEXyl8uNakl175em/U6RONxr3aeSyAv2UoF+NNDuz+ZTifWFD7QwVOioAkcKaAQFx34C
7AZD7CgmM76pEs304wHNMcFrc+tEgoWxU1RU1oGkLYsepWuHExAaQjmOuYV7HHqVaAgkI7qCYttY
RvNWduPUEiiFL/KxuUTjpL9CmfZK+Dk2zJ6f+6dYxpfXGC23gx828geDocYpQ78QGQq8i0dn5te+
E0MoAfBsyCbO5GZmfbgCbzaBzKAXDhmPhCLdka+/liaXkkLch2QB6cvVlz6CRk458eDvDEk5oJNH
zcj+p55MRrRlCB+pA3kRGrxw9xtRNe5kD73rt+Zd1dGSxVrg6zZX7OJH3K5QtCGeze3qE9VFHSAW
1gSytNib/BKUhAKFkmGcdeSNguNw5tNQkOxe2R5Oze2k36mQwEojRn8GdtLfIeGZlBU28qWX7/M/
BkHyoPtekGi/kB4qM0CatDLl77MWmdzdDBM/Za92b5qK/KhNa5MfWla5ufhGxqXGKsgbnw+Zpm35
igd8GhDZYA85D8/SR/ncdYTKOe0mjAMkclOgCsYzEUsqHQp9AxWD1YRN0NTFQcGMcH+KV+sw6lE3
xkOQMxNQ8phWgPV5tkuzOWJE9Q9EOgqG6pqug96yPxD1Qq/TUdiLPSo+qOzBHDN/4UNp3ERsHgai
MFl21Knq6g4X/MG5vO8lxFY+3o2OkatOEPQtNiYDcuqiZtZmKJmUKq+v0eh4M9HNR0TBmiDk5kRk
s5DWaH+KJB07ppIuPANKROGGhdIEU+f5BbTa9OhoVHAa/l54889HjV9ip4HOPCXCarFfDXRZOksi
B1ZhRnueB5xo7Bvaf/y81vb4vjzjvQVybGPCPW+x/mJZekyKPmYcAGLn9XMn6CdV0JPXUToqAfun
46MCXX/85k9hZBQCeBNKbc5ELZ2hpyyZ8QIooqADIx5Jo24YWQ+90sqUfx8D6OQOG+zYNOXCeQL7
Ga3A5/sxDE14+HGb2gWgWOWGT6zVeleW7GhAuuTOlz8/l2uZG52QSsHtX6oNjA4iU7Pu89hcd4OY
QzUuDmuG1YrgvM+uYxmpwUcNCNa5LbkeSFIXKc8qk1EbvIhs07uGrlH6IhnlU4QKINwBk6zRRoGN
nYuZ0DeRxBJZkrqOWbSXbbFO67Z3SrpqOjLkoTIHWrKWUsefZ+ZZKcqu7kI3BK9uxoBRUkXSJevS
irTZ6ssqlXW9+RkGOUjtRyQDWw079PeajNXyRuYV8YqJ9izUzuO7S9AanpMq3GawtPW1nsxnSy3T
SSvNQdGgi0STudGFiYSiezQGEb0Hfdnez229IAJaVpAwKkqmsDlxhQiXFhmBrW40LYZTDMiXG82e
CuoKg1DdegpVONuqvUlEopYwU8XoN7C35IaBPPwhVuHPrA5rNk4cMy1I0F8lIR2GXJiybuEgsU45
C4XAqnJqQQGgqgbfrwY05drwfmIJ1TiIr2U4zvFshCRO5OEFIo69MBeShHds0CPevCk9lkXkfXJ4
g/Nrngmkna2Zb+9aLijnuUUfFv9d4SJGc2NmptohQxxh40MHJHl0FWmQC3uYFc0/p8NS1Nm02uNK
7tnrXcjjL8ov/nIKsuGj5qnli/7ONBLLboMxFpwRx4sEMEx3qC6wpVn2aXN9gc/wA12d/Z9pJFSL
tg9LvTTJXSCPoLafjEwAUvKdk791kDCbaVOp7+jLbN8doY6Xzh9cYOnlpPslkFmNfqml9zdm9ofW
SxtK1Ov7KChmPnVXIh12SCXPXfKK2vERxMkSijTPi4BaJYKhisMecDC0SooTNkdPRmEa94+DLBO9
wQNMDBmOmiW7GNhK7Ve7lM9+zdEGZyrWUADqdWYnALd9iw26wBpmRfUqvn4TliFBVxcQIzNBe+gm
cOXOnGSlHy/kdJ3se6Z0WMlS5V2rBbwQPHXLiwZ3V0Bow2Cx1AbFfjIsquH+36gXE+7kJfWqBMx5
XVGQp+vI42kbHT+eYH5dhUbYbJS8xTm0W91/55YZXo1dbV2xnzprLhG1KSw+FSFcc7Sd046FBcTt
5rJy4Ow85ezJ8fmQoXWRnOwbcRGl6WLQf++YLBOP7eEEWIAVds+OKNh+eI82bS9Hc1oZ0I2M+8va
dZVU8QETBdZABgYGG3XbpmAPeq7LEYLgFqbHjx8QSDq+HSHrV/DWsULlOH1mXq9KDxJiQX/7oZLp
yGW9R9mSphl2bozUGMAeqEKgIlbzdUBcLB0LjMBh4Qlwt0RvxpMPt9FqVUTQJViDV1argyOlDubH
2DBkE+HrhZgygv8JWZjWcUGsIlCQalCm9IsV/0NBzYpSuzGbirLWI0tjiVW9IsRVgsIjUO3DX5i+
7bqI0bmhEqtM9CSFKb0CZuvc7dzUI0hXzSAc06oPW9K2mctxOi6391JYljoDsyilmSJnk6EHFA1l
1Mrd/WHfvQKB610ObHA9pdNr6Vduy42PuZF9vmuZ9Qwsu+A9F31iarYU1a19Grhbsilt53rEK4ZE
WL8ykf2hmbKzdv5An9DWEcMpadue/EpyTVT3Eu8B2uApZLJr5tekJajsqrwt071P7gZs3qP37Pv3
7sHi0LHMAShG/GBPPITbAtvOzrMd8KmXpbiVM3i3+vEg+o3Lo1al0UKas94lbWyrJdTXQvt7BuY5
1RNadG0CV9wm6xfN/R7qbnLshtDPo7OEzPxLJySIsjLpdjzlA1LpMecZKBKxSCi9IY2KMTk86PBn
UFb/kK2IwI1u0dDy297hmE2HZKMzlYIB+39LqFuSRv69IR11HTabkEA9sOBY+0pr0POi0L4ekkhH
2o8QUCwUAQQw+whg282ZH9rfwhOQf+F8eNEtwuEdWA8CQbSeU2zJ8m34nAl0YJn+tTvCb995qupe
WYo6b7zsqJT5IJ+etDmyUeSdNRdecBlXe2nKA0Fn0Ve5DiEfIAcgJs5LAAhXpKhNPgNZEtw2G3fb
K5eLYNrcV9Wziihr4nDC45psWCLZoRVyzOLHTnRwjVOrksuYMKxvJioMxspj4qNfP3WOZ0RiufZb
Sl2v+5suiZDLi+57Wm+hy7eimbljvAXWcFpR7EaCbUAqFCqxj4Rp1B6EAF+iZVOv3cz57yg/+g/N
lCZBNKbbbpn2ASuuBNvYFA4/s7vaZjoTFhyoq+wWnvtARKYalhLCVXRWATIbIgoqfkmBFnZB1I5R
0ZADZO6E2TzPYm1bxOq82aWKs1fSBw+ylaFnflMW0vGRTT2vj0aouIIAK/t2ugMNxtCXJJhmX1YU
SODrTLyjy41A7ZDylUk86U5nft+pbeGySSmKtTePKc1wswTyJAURk04/aJf8sdiW7sQmIO6XpFSj
FvodOzpHO12zUlPsFFRim+W7EhdTEx8xXhXYeLvSkfyq8sbJeCNOkm53QRb5WXaG0pbS0TJ/NMjr
+199x4flDYNgeszpIR0d/Uwv+BFsgb4TSVTFiUQRHovkx3g/U2rBvvYeOYqPdVteu6I+dYAiMV0o
5HsUKpfVx2vDPXXJwh2z1dOdhIbN8uMS3lHiLArwKE8akGJR+fDMTUrjmXybACFHcmTV0kioJViB
2q2w0hwVG4mqGfx5xnFDyjIeceCc2KWPRHULf6fHo9syVe4pCUW5Wc53L4jEwj1+aoEKVDI7vGQs
+oNhju0/9R2EK7uZnsa//GQcE8eJggsDC5uf8tYwVzf+7hrrsi6nI7zJSxNIGcID422zr0SUxzoi
Ad8yHSKsHqigd4lZHybxHfS6jsLoRnbBYP4/1YXsupD2RIydOPJqtMJBMW0KAzvX4/1Q9ZiubHPi
zSEiB99JPtzcnFxT+p9fbTsqFHlqXKRl/WrVGeSF2BmHpRuu8azit2X0gcJHX2vkCf8lv4XfmlIc
PsVzb+Du4fOuxra0IdaVHhRNeW/4/he+c36TmkOK1QTndKsEHTapKX2iKatn/zlNg2eqh7rTufjb
ji7KW8yjQ0jXnnD+UN3pZwA7OTLgxIZ+QGDtXE6/NiflFsh1hEcZTi3bbQGjNYQHa/cwvlvalNLE
8GFKljRdjap4439prQTrBHuK6zCQBg/vOKQ6VuLhlkaqn6oKx5tevB/GbeW7gkR/kdFSLeTM8P7t
5GUIDXDjxwQhhMSphvj+FbZpdkNTjMedkuXVQe70rBnQpC2Z5knT5TVixZwmRESbaAX+rxXVGLCa
c0h18StS6CNJodrXOXGuugIS2Z6bh2Nb8lq6lcKTHVPsO99WYpTsozDh03qVDaYa0miv87UPHFkv
sJN6JUZGJxK2NwAUaNxmBlX24VDMxqdNVa0rKsSank2qSj2RyFSyJeWFj9hW9zMOhSmglNuw5UTR
NR/tAjD1dmH/D/ygoEmA6m/NaOcK2QApHSl2ImL2GVpNF6k60XlvfYrQBJQKKsX7yG597x4Igf2N
8SAMvZkT4xF0PRgSfU38wHR2Tuf1Lr6t/SFZViIx4xZmVCUn24ZcQzYKHZB8PCnKysItjW2tFIuI
JQUboe95j1QElpyBQzatO1B+Gk6lqI01d+fACU+JbnoR0jmQ/Vo/+MAUCM+Cx8vC1z0gC3dcHZjF
v575j6/DouZ4TxR11vkVIXhcFzoBdhmcRE21i8F5gPWTX3uT2hpX6Siv14TSY4NKbynaHQDlnNfK
an8sWXhl+0SOIj0JuvfPfyLyvDnT9y+0ndzHcWNBw1eqgqjXZHzxIxpAKRKqFC44EC8E1f8+1XtI
Tj/nKoMO+uzqyze6WXNfrufYk40lfCHYKJWEncp209/tqsWcCOKf68K2cF2TizLlqLbHIzV299BL
nNep6E/dJIz4bof91YyXrBNHv+Kni6I1QBuOy0OMCQDoATQWwcU9HIghUYurxvd1ourEIFabSAEh
M4fHmu8c3PSOS0Zugba4lgFtzIS+O6msT6N1gM2xNGMeY6+Bk/LhaoeCRdjHYiKc+1h0StYETiop
Gfp23MyP7+3RNmitBnw2/H0QVGgBV42TKC4HfbhJP6GmDgSvk5uylCU7wkdvGUdWJl5qPHJ0i4FA
leIK5z1Ax6cEotHMhu2OyfgZfg7Q0V2LectW8nq97vdLA5r9XPiStsEyd1tXignSUQeUhD3el/vZ
oseBbVlyu1Ts1koYnI4j0M9kISgF6NynT0qvM8Ijda5FyukCUnLJzB35oyZAqxX++Fx07mVqnIHo
xEdEEYWDp5dsLmPunN9AOPGveMbbaWPtQtH+hIIH6XRjPqWC7n7o6YN8wARHDOLFCcB0FL6MuRTH
w5XFWPxYpxg2eUJt002wxYM1rE/N450H2fcFpfgd4aX21gAfQ5mSe3PkSZfpM0SVC0T+S0VptrAK
NVor8AkZTWRTWENZBpXAV+CFMjAqLxRDs5z2PvFRG3Q+tdOBpC5XsjRYuhD/SBk+/wJaGXqDYdua
JTeQxeqRtu4HAokqD6vHZTZS1+XZozZQFHFKr9lYcuTvaRA0ecUWCLAOQHRVe6AZgU+KH61LWl05
8TjLqeRdLfBNQ14jRteQ3B680bOCpkdUZ9ZYKv9AH8UPVRq5W3KJ6boftNEjOs/YM8DUzCwVyenj
ewCltKCFLJaQsJY6Dg80ejFPS8GJduRnX9GxJBz8RYIZbjk/fzN+48Y3HXXtbCmt6FEZ1vyrBmmZ
p2kzHwy4jlaFQ9PmZpEFkTty8JHgAO65LbRtGoeBgNBlbnrCFYiUNeld/eBgVNJTAbZ3l/2KCbyU
o78SIO9t0E0GmARxeFjZjDf5iIQtIUIifCXRswe0381TeFWrdJo2zSXTDQ1K9ABrvosELIKRgn72
KYi89Rzw5VZazWkElCu7pHuznKU+H76MSxQLdH9br7SUxkS1WVwnVcWcOsLM27uCQxZX/f9eiqSB
VzGwxLkZCe9+qor/Fdv0ayZhsrwS1KI4CSPY3VAuQhBTLgaVDs+AceORKlOuWdJc2ZtmzQEXCPOj
sRfZ7i3AV/FfYMpG0k8UwfB7NmBErCeaCVtXmyD3e1cjhAYDhjKwE6sdGV/Or4DAL8t4hrR0il1x
pq6fNegIlSl1oUVMVRwAlUp+HtDyktBMipnegV6dYZZ1Rc2uiRjQSo8eWULeGGvHiwsebp6b5XW0
h5+BlFm4K/zUMwufkUOAtLT1z24cyCojGYndmgN459rC0WlXzlRFXGThFa0+JoEemH6g6gMOhI0r
+N1DwAdqAecIVlnEtRHtb7cxHJzbQ2mqRw1l7WMRCoXHR3JwXo+qo3GcnFop+JZDQHd+m/zxWMa1
Cgny+H/ynNJGmglF/QVTVMhLATw6qs+E4KpPsZxWNqRyrRlJXgp+y2sFo0tJ9VsUXXzYLZEQWOR3
Crvc84duWu50AGZqZM7IkHgmQyoouzJEXpXiNdsabix1zK48OG0Mj768IMSxGnZiVS6UX9ARbXBv
mnoCv1SepBN9YGlRKWVC6Cfxizz/s/FPY4c9sLdeOYIa67LCnMzx5dXsbHy8TQGVAQNkDacY+iHj
cMJTNoyslV7aE5YQkqg3m5I7JODJZQYYkcL8td7/4BLHG0bxAfd3l8ET+3IbNpzZq9SkvMtOBOsL
CzZHLahx8YoglITGYA1Ld/7z26exWR1loXlmXpNiPcZYxcU4U3XZR634hkEThqQUCwsjsU9wsaVc
zRoK06rlScMxiGT5bzudjZZd9lvyjJ7I6On70CBO5ALiI7Foeo39hCH/O5TvyIUOatKDEQtFBB5l
eNV6jHdkA0J5H94ehvdJAixvUt2v0Am49ITiaX0GBdYy2wws/mI6gcHLnIWDIfrE4/KrS0KdJhTq
up9Ln+BcNbxjl5EYbL9kuZmlwEE0qMaqQJnGSKm1eseVb9e4cZRMmW3Wy2GTZ5GYhpB/88Bi7VZF
I9MxdceFMqLQhlmbhm/NYCQ8QGR/xGnJIIq8TXmds1TdUnI1eNVD6+eGizVxmXD3PKsUgJURpsn9
leRO2yMZRfFFOd9CYSaTLVYtodX+V8wMT28DidXeciVp34Auid4fVVL/8j7uOXrRpZslDxsMy/62
jDccHsaXIUpYvBJI4TF15vDmN+QXyeIJcDlpGTIeai2liJD3SkcJMwfSgU+t3D2mWst2GXitEMsO
b+WSKfksvw4cmRWAgBcS2FO3KWfeWIIlSgRZsk/X1r7iIgmB0bSDU35ECckVSEqXrZFsXA+kGXyj
tf6/EBXVNqBjSK9/rdUiTzfXjUk1ho6DkPj45G4sG3NWiAzlVsBJndmEj9EzuMbrOtEM4BiK7fFP
GMUcd7pZipxDBSk1GlDSI6k3h7SuCDShJuEonYPLwP7K9ss/H8rjIXz3IUj3Ki8M2BYkF50zlKzO
t+RPNhyg1UeJTpSv9xT6mNxGxkQ3+0xEO2WS8Uz+zO9yPinI03i3GEiuND7BRzJGWRs8bWdQ9tO8
ew5rx5L6NEgwnzwfc6HqiVLGhGGiTderx8Vt8zz1C/f9UTKQ1IJUGrEPfpk5NISUyic+eT4l5w70
AcBnjs5hDHChrb4rKTgI5oNDF/jRZ1m+aevyzoroSB1kglK06uewD4/F6SacByw6BQZc0wIabM4g
SEUuyQxO1azJwVdXs0Hib9oqkkJhENac/YVldXeWCXLPX+P6l9+iptBGi/OMO2PLLHZhSn6mQkQA
qhN1ZwOZB/ycArBpbkQTl5sp0DfniryCHY/Yet6bYFtDbVE1jfUm5oTqg6EYtMePAhGvSe43VPmV
2rlIt0HdVvCuakInMSBSUluT7/96/nY0VeOK8KIy4Xxxl8590ToS7REMnmi4qjEU61RNWzr/rWrz
VP5fDgxSCAawJOWVPPFDe56TJhUI8g9a8ngFtmJyH/kvoqhLux0o25BqRFnRIklV3QDhMYtk2kjU
Pld67BwgA1qwICkm4c5rBrtR2v83vuUdqSjCJJXLl6B9ITGGBHI86oNMbYJ8UAqd++VshLbdNi6C
su+X9jLByAU8mOFLvmwvRt+nLi4zp5DVYDLMEitnYumo8vMCnMFglRm0TjrSlBnxwWyK3H89Clrk
7VSCv+Hf3unNNJQpuiEBkkE9f2HVjGdPkzRphEHa0M6x1YdB/vYdB9OhxzPLe7aXpVsA4BI+27bV
rC0rVkNm6asFcjFbojcnSrwPS7ZOHj3rSjWlQf3ULy2TNEFeit6wvsHVxQPmLJStHKdQBx6mCwcE
y7SEhKRZ4DzzXM6jfhe76j5dxGtxljt0dGjG7f8DR++m8CDaAuLf5IE3RS2MKDKn/dKdOPWjAAft
8OuzPElrEnIu/pGE4uYCfyFU2Bo3ehy/QMX9+KpYJu+ga+tYCVbRPMeUs9P9iwuTAYznpVTA8kvG
jRjol1X+HSzL7UzVjGOMu174hyL6gj1FmRQS7kvSgzlf3Fb9gg/YEy7XsLKYk4JdaF37bWyeL2GU
o/kjPuTcfaLb5JPqfsyfZmxHpMgrgUY+iCtzWmhSEGoL8wbCPEyftmNxGrDIG1X4y5shOG2c8R6I
UD1jtUOOaw3tH5vEQCZKDPl87ZB/yZVhwKwNDh9IptrQA0d1tpfvnrE6UXwhcJyJyFa6dByiEGwX
4S44hNGpG8k59WfOJpfGp8A1dq4pKBFIl6DgcTgEjVGz/PnwhPCDZdAyoVKe3igWROXcVc86Fg2H
aHrnqSBWjGisPZWHvkUgY5KOPirEgeamVFRTJbnOB0oO5e2gDv8o+RVT2H+/MGesg4/j7AoLvIWO
li+upPpBAZm/hvWMO0BPYlXEIW7EP4RDExo55PZdbxxdW350ixRJsDssKqKMEVqbr6Hjueb3JZgt
q/P2tA3Smyh8aLKVGixzHCVtuJxiDiYServsI47sMluopxS1Y2k16D+cFTl7ceL0aJrrZfVKGcJJ
kUrjWkVNJY9SzvNBkLzns7/4SzlpiR25KbyGdQbvtO/k2iddrxB9ZX+RFduG/YiBbMDRsf3glwfV
nJf0tsASjB8WD7aknKICpv4ydmA76s4nGNjwc4tfhSiVgMFttsCNltI2fyZzf1T0rsMLZAbrjhhF
aDreiwzRKlo4O5YU/8cOQdAFKYMtSskZ5Z/5gm2iQb+LRSEw1QL0KwjRAdmv52NxHLBtwy+kxT2h
0IsMG5IXJk4aqnnaKCO0VHP+4p1dkHrlfMeyWes09eKgC9j5Dj7Mxy8987ZbzZ3Or+4WSXIWsLaT
tHrziG9Jb5eNPS+FxpBKCr5uAZQn4G2s14D48Wep6/zQC/hmBlV88WJX4Weqp3iECx5J0HGPb2yc
Z0vLJehIX3Gp6O686i/PUqxD4/LI7xtlQPNlAzceQvw0V6TucsTrh6RxtUWAaGjNlihmN6n+okUi
+UIAeaBh8FJNAl3dJmOn72F05Rm/aDH0vNerHw3JEtJ79a6DnmUGtuDIxV7BEyOTj0XHMdtNuttR
l1Hfamcc0Onr9YE6N/UKBa8764YgrkhpoctQl2DjGdCl4HLYrGE/idYl9L1+4GN2vapN3hD5oIVQ
54VEjAQOeQsSy5tO3oL7kXeTilJcT2cjds2fDl3i8uNJ/2Sj9lBqsnzAlhcNHTVVEM2QPwOxIjam
/feX+ZD9oKC/6DzZQiS94CRL5lksBoh6VpPW3ZzvUOycL3/2/6bYCcLkp+PiSgigwEVW+aEf0OG7
JxC2fKphpj0g9fvvb6QSxtRzRXvYrY2YABPKSdlz22CGK9vFrcnNmWBuXcJSYVu2ULap4C5jupV9
UV4OZ5No3POeyPJjjUP/51/jagBbpVyA20e5wkOeGkBDSOtiMXiT7LuEmu1uN2XqtaZeBLJbDm8k
ToN8W5QKBMdVv1hjeWiuKvQDR2YcEwK1rSW93ZtIbxMjrTp77B4Mfsk4YJ5a3BaqnKSER1zyF2EM
fQFrGWtPOoyKcuXF7sWFm5E4jcnNGCvozSB5vhjmcZuR7vEdy0h5R2M97Z7OqgDt9Ck8mKhS395m
j+V+kgn9iM44TsIF9QxIBX6E5RnDmYY9BnvJh3UO3ud73PInsXdISnp/m/JyGENphR+c1/0Tm3LK
ocmX9lDmejSM7JL4pA4I9bxy/IIDWWMzQEjiNdXRbYjCEttwn0tCW1u5apQBIVzd3SiglDjWd4fd
JOgw1A9rWQoGuYq2vYLOUSEI49mrydTnhAXKBNJ+y3h0Wo4go1TPcBJmBHZO0sMUAdgl4CxctLAG
ddbaZnu0EganAtpgiGhoOsvgc4nnutWmOhPhAwzv3iT9i5ujzShdn/g4pii1c02y5G/m7/T1j04g
nT8XPgfrdF1a+r6G37h2v0t9NMFOzHzgCBqH9v+XkddMeZ49lV0EBwBRM6ho0nj8wdg0j1gr48tp
H6PHY64ejwfbseHJA823KzY+r/FwS5sHNk4O/d3auCyEnqpstpMQ9KR+aCM7fodEhqiMMgPpeC1J
UC72NXpB1CM1V/weuAgRUeP5+UG4VSEE32X1le5UxsU2rCmDGNH2FNWIXPQn/k1Pz5iQDMkRatCS
+t5VwPAIapxlPrAPZE1gcGRtaGdirxpgcuHmXLx8QqzHXoUuzpwzWXkAK66QkzsgEUT7UYkOnFL6
hR8GaCiDVOActORobYkMRO46dAtSAjRMrB2GlZSRr37x+zfaSvQdl5Ugv4MXmfe6CiJjwpQcY5QB
HHYgmXv+GEwBsPRMXEB+Uvg52GdtGuIOM6NopNkDCxahnDbY7x9VwA/PRp8A8FLaQMXhcMHoGFhQ
1pzO6XpxD2x8eO4JOl4bQcdpBhs4HpMM9xKFPUDPgL2NU3fPzwHDwK+V5NnFviQbzWJsOb/eyLJs
ONvq6q4+VZXTX3MwgZlkeeBbGr9tUp7W8m2BIkSl2gcnMSzd3FaW7Z1faJa7bP1Eg2LHcNRvY4OH
xVCyJF+3C6Oxvr4llqvXi9dCgSuFGLi/pBgljQuO6hVf/C0UgYLXR5y8JRKne48BAT+ZwXg8XHhj
OT/eIvQsdUFzuLqQ3rMlsCMUL85kNOe2ng9yRJQwlgbSCVVgp09y20AjGbYZ+AFrMv6PHQt6q7Ce
ma1WqelhmA4W1kp7ba2ifnZt6gY86J2iP4z6gC4N/0LouuPpXGXDlZRs8MZa8PQkmcWw/ZwB5e/h
ptes86etfp2pfCeIEJyasSNvEUzA5ZqOxxwyr/apWmA8ppQYYZUxNDk4+XiHSWzxbHYyEzuKodmK
eazjnrF9XwRR734m5TZ1JJo1hUxA0JVf8hqQTm5fAUDoAvxjEmhF3qzT4eeVVLEWRCVHGhgVga7Z
BopyGaLKb6/KXUSjT/Qt0gKoKXXH3lBl5cTse7Hkz4DbOlzHgQHnOpOPzGKtQxYkmPrWHNo+VWNA
v1RixGUXEN+sONFtmPolIcBt2Fcz4C610+57hPLdCC6BXK1q0aqSsj93VWqDc8ajqY89m9RcX4Gz
wTZpHRRhLkO9wdNis8s4kTSDHHjLnLdb+gRJcpTPjoKZmIst4C0cYdwtpbQquL2xmFRpUDbV0tFg
02MMgPGuOyduOIYDLHNUt3IV3OpJx+Xhln3+aqnvpC6xnVXeDKRAoAZuWv+RsfVEYOq4V/NeSQRW
7BDgkFCdjJYrbdWd2lwgfbKXTVLOqWhWXh47ABupclA+xHlSoG6RhNfzX1MlbIYNyS9l9XoxqDIz
3YrY26EXvGlKxn0nf/nPTLkJ7zqJItU4Bb7TGABRRZfpOQG97xNENgTa75SczHPcJHWIQ4gS44GG
wC6fl31L2iC8PuB+35ZtrQMROkx2+4jsoq8wJsBWOQYzqrrHGqQNikxbZV9wtfbb0SUUgxObNMQ6
I2f4l9nvv4+Z3AmXCjj11N7NzhHfmNybRiCUs8JJXo2CQBvq5EEl3U/XtF43WN380rXyX+xpl8+t
ViqASNrmjuTRttCQwoNNtkrFSsMDvbK7oXxuHwY4Y+KcjPRE8JM7Mbqhp5M/zyUQ0ELnSrOdZNt3
bl7PmfafxRL0N7cGKzimVYXUlkSsV2JbtSq/ZL1DyRHxBYJ3Gsl7LUKSooTDTFE/JSu5w/eR9O+v
xAmxci+/azC+vN8/n+DGoAF7kTu7i49L/c8EohXQiyn3DykvWO3ec4VL+bPojC04UcN1HhMutD+G
5cL5AGOy/mXUDKqUEv1dGI2Rc/UL2GfcI6Owv5AoBddZfPlGKkxq9b0ggmv9RR6drUnvU2jOJgCZ
KXpEl+JeB/RT71vWu5fwuBUDvvRQ27hDFU9Y3vfaFciu6IZP/pphex0ij/jazq5tOWxnuynv19vJ
njRR8+8vChwvDRXztXGBk5Yuk0E/KDtssRWpkq3DoEogw8wvkfTdHTd0u8F2KF2VkS+K9U9pYsaU
UY9EsVfJ2tdKAQHUe0TjgByoq6R3I5uB7p7Pddb/kjgCj7cSNmvQJLaHoUdNyMQxZTar2Vz9UVvJ
Dpf9/qpuJ/pLN65jQF87n86BwkD7OxNwTbY0QvliOahmc7Fb6Jf2C++FOBly4HsJFXpj228e6ebq
O8MzRdiH7k4PMFQ7gNaabUR6XfQ9MQOuwYOFLPA3WQj6g/HwuzmV3ByGoLDr113NKBUAC+eXGRUs
hPLpUdV+DvD8oAepPonqwS88Y3JQpMn7im9Epkyq7iKfHDMhucY09IaEkfIXIyjyF1mklpd5fmed
2EzpL3aIGqlzPKFI6ZyQ5jkctt4J4iKcxOIb4wUCjQ3kZLxTL4et4GmkjaTxD+q7iaOg04uueRuy
8l3ADQBkoV9+ZGI0Jl8bLKX1EEc8D7KTVugPG4aM/dYwEPvVcwNLdgLV3zudJePNWmWJYJVy/7Ck
BRLaYQCvfJq/8uOfFRkuKDBltjXsPUNooBda94SVRx0pZkZoXg5oOMlRZsOZsCw7ls+vid1nsMJK
StqEI8oOZSta1LTep+ScZKRaJ9b0Z/J9WC89qmFXj/SncX+h6jN5Upj8VirzACRRQg98zlcG6cSp
PsUBf47S1wlIPiqFpfXY4Vz2bwtAlt+8vbdZPXNO4sGltLrx5Mkxwfn1qspA3snOEQDEUzSbV8R9
VL11wP3bt8QiJEz+en8Uo1OumVNhHpQaBDmkcDDVQfxzo5aBR9S8r1s2En8MVvwbHBQ/zKqF9DAW
n+lp7qNhtzf5USAXOGOLfak5SgHd2odNAfEXRNN7tMmRYkj7DkQMw6SZPQ7GbehgqE7CqcTUuoR7
g+9GK0YbRAghmYigOZE3xJ/GjLZvw5Dou28ok9PcOeCQad1dy29DwlEo18Ij7Xsb9LgGH00gKvLq
PsvY8yMBD3ZMczz7DTV1LyAB/H8htHkQggwMepgxHkxC9u94lFGkhM5WD7bBjM4fCnHobIyTrlFi
O3hog4RyUgPfLwi8AtVpC5m1zP3tWZXgld5YnjZNLAWvgBgFY/wLApQ9Ur4tyXUZWeqyPslX8Lp2
199J9WAjKNdnKci/O5H0fMOvRsZl8YGxByX252ybs1pvaM4Brug3pWxlF9WakcrsufveJ02bQwVH
TSqJuwPI1bmXH3beGaHNzTWju73XaGSNzscwCSzQWShfH8enPQIOwCocyXjNwpZ/TwuAtNyvh+lS
JvZRMISA/W76KrUcZ7pQ1VBFAzzMSaOafXPSHdjpNja4yYfVFsFXELZoZiPki/75qbxg96s7dhiH
hcOeVuA4ULyvWiwe0Ho+CPtFZbfQCHunj4aZEVr0Lxr9h61ibn7M31gV5Oz/CApCOoW7TZYF/pPm
FvObPpA4O3hMbTp+OMrWK5aROSU3CBMieqUVJMXSBFG2nbMWDyt7GAYA6A34Je4yeYQ3t10yXdiP
zv71difqfHBo70wzrHUNZoyy896KZ3rAzUuChVpu6rPEnmHvSBIuEY0efKQdhfB0NmuRpEEumHQa
YAPC7ZLCfhHITjhLrOnQ06/Jijrpyra75BZmvHwtLlooA/2Ng1+nCkhwT0SK/7FF4fWJ/eoSjg8v
3WnF3VUGnsW9NLyLRbSkvX4SqskKp5cRlFjkFkKKe7UUAN4mPYWsjT7+1qFtsXs55OrmdCHaNTfH
G+Kiz4KLM5BcMubq0+DViKnPBJ8AjyTBfDv1a7jk9/BfD/3+6wkjLjCtOi1QSK3RdyBjfQk8vhI9
HAehLMatl5rC8nvwjzKQq9AVxICQrfFdjktwUsjh4du/5anqYAqGGHZ+HXLUTeeFQz7DdR3ptwp7
ygyOwls0gyNZITqrKPy2/mAdb20N0hZJbePyx5nbTMvmU2TB4n5ZdXSSrLWp/BHh6MNj0vJfWeqH
SzhYdM22Khb0UcuH8JjMJJnbrKYatGdAsF5vNTXNgkeDbc/HSZNMe+LTdrMHg9NDU0PBdSr/HgfP
RgxnTedazX51I6w7LvM9J1mSp6PDOWXHWKRTgju5vpxUUmFf82zB05BIdh0uNKw8QvEmqpbnnzaD
gZTezE1+Zcem7t81LDkIik2kQLRj0SQXAZqcNbMGEaNlpgJfLdiOVq8qBXHMvx8MyZzZjKuEfwiL
GW2+xWa0mudCZWE9fzOmNQKrrPfAsz8rXnlWGZ/DrAhp8TbqOuYeKHgIG8MCnMb0gR7Jr8JfUPCo
4jleHRBB+5/D1Rru68G/13jFJalYAoGHebus+cFnBONpiW9hpBCr+E3N8SuVIWJmmcwqqwZVWuiX
sR57ZfTx0A7uUEfW+a2oaPIKdTUNcsR45uC52buVpjqma0GgFNEZ12biftwLz9I1t+gf0vpvuBrr
GXPQptahNychkF/88jqO2rUF6fBgIM4ENQ/eCPWmAsl1drj8+gntFtMPemiA0jR/O8Cxuu5jn2Z3
tl0jR3Ysbxgi364U2/ys2OjY0lGyHbzMotCio7W4aiJH+lKJNjGP7EfNTNdHqehgh5VuGHawfTfg
UzQhP5KetvvPXWHW26wRGqKx6TdEgrQxqs5ivdw8fG1W74Tktan8ipaWXLEq0+TIgfmElkFWRKHH
IRi0iBFm/X7LeEsQqlQXUmfKRmcYG1NrNmV4c7VcMHxBn5kKlJAjqN7Hs/Anp3G9HTw+RPqoOWd8
5B+qoNvTr3aSHa64HZXjjLriAvjaEx3tdhHAoP+LStt4O4mknwlaav4eGz5cJUImwhyl6la2AfTN
OXCYYFojwt4Xly+j9gH04YIKMnTjosBqS6H7Oseb8QT+9GwStiDzRJ9kdajvvLxXD8xDz6M4WfSm
KLW7VcYAJeSYk8oE2br5rDctfJiYisOmbdtR2/WmDtfw00WglbKnketGcPks2OhwVyOfWpMmD9Zs
RMx7Y9EAayls0l6fplBWW1ESl6MxMaIgYV25ejgjmvwAbJt+zLlaoJcS5z27SGieTQchaxIAdmXh
5lupEi8Se6LtDP7DooXEJwoh2E0nJ7LPlRObqI4CMN60oKvfB0kDUf2vpl6npTFpS0JPLjsTc9uL
lCmIBfV7bHeMscQ43wNOArE9GyciXqnr2XPZ+5qp+13gh2SqcsVvDYq4woxyDxaPA+ELyAUFeVRo
ae0G0E9IvGrYd/HPWICA5mrmm0zK7bPWzcrlaFSiD73nll/dFHtMwU/a7VM3jy4lVlIrGswuahyH
nDXJ9tDLa5Z3XDSJcAx3MBW0fR3ePf5nBheGuFWzfz9H8FXZKhZwGWA+E95zgiLziljVaUI/cpHb
QaD1rrPvQ2+nG51t9P6qjYqZJ23X8oDYeude1rXut3EtA5mD4+OhM4R5Bdz/y4babTymyT1/m0Ec
JjXDH5yZ/3jWJC6NWM1OWnavOATn2TuL4+vSGtC0JsIfbhKSO/K56JsULYXfFowAsCjabfXUIqai
rZsqFAUxI9JEKWmhqY2pNl+98DwGr90FL6uJCHHHMUpzEGAtudT3tab5gkW9V1wecPknMclFhpwG
O4zBIChiNjmaksGwBYGBlwtQeopyFZLXTzbaMjgbFCG/YHV7x9CVCEKxnMcLDbcML9TE1A7Y36MP
i6Y2S+f+Cnyo4oziL1njmNSpbIMyBMV4oxuHvIVgjF4XMma6WuUmopBkVUcMF/Ochjo4wh/G2CRE
PDw7+rtc9V4gpAUvphrw098rUxkMicu9CUlvkrhixUuMmG8f0oE9OsBPc4j/Su2jReuTfY+6PByI
UCVC3nFbeO0bndAdsQqM0tSJoZy97h8ekBSN9Xpgq47lYWlSeTxN7IKd1qc/mywVTGqy6S9c3lbq
PNC/T/zVhu2GGidYqldIeV7UvN/DJZX55ldEzGJKBlDhZe4iBcLD7jwolnecUkeGdLi0sO5DfDcr
5gibB+aWkztThOs+O4sitxzQYxhC1qg4t/UnK+R84qEbihV8nBQE8dlfTisGCXetYcPKMpft5BOl
FSA89cEzu5rErbX8M1z18UP/Qxms0uupHDyjbmOxaj6JTzQUGPo4yjlSxP7fgkG06HvjcMBEj2Dc
t03rnyQoGg7oeqW07mtjluyVdmj73viC14KUq8dgg1pSMPphuMffpa7nFvHLsWMj+2QT99Y6NlZr
6eoiWLn2vx2154ead5d6oZZPy+8Rc6UF++eK6xLeFmwV+c4dAPRqma9dh5Pz3Ze+iwY+osOpVpxM
SYPOmCv2AfdpF1k+qUjeqENK+A2QHzfsuJW/fKqjXzE4ZTGFIdCPeq5RuLGfAxLR981DtSpYVW7b
HAR2tSzmf/UrHBs2j3g2u5EeIcmwZNC6EVsC11KNtgxtx5q3jj3/a16RLvwC4+HBSh3ndOs6flDF
+FaUameUUCLdolY/QM2o5RcoIqYKsGLLzxNsH77mbnzI6Mb6MlB5U/+UTPFL2l8sL9EV/VsYEJpl
7542Hbg3yFXdbM9hpuuQpKBUORXSHxBC5n5jVqdAlakDdrOMdSDtMVoJvKZtGg1BptOXH+hMFBmO
V9JprK8JLg6vNHnGsDLIKmvdqqytwTpq7acYiVBNZjv1dSVlgxqWQbbK7POGLsadM5N29LD1BuSZ
jslOPFZ/bh7wq3iwgUtOaBMhqpGgbxu5hVuVIMlxRwOH6vlSUoqTESCdeeyKRMKzPiLpaFal0dtB
d+2jsO/iksRyOAqBchjeh3rxTYwgx1OA7OENIEM87dVQuAJkdjrOZvk/DNcp+gEdnsHrVRGWy+XC
FTXwRy2THeMhFnhFUCyuA7+r38WCrC/g6e7hPg2zBp8C27DSDNDKIdoJG/ATSrOZwrfK5baqpblM
NUTp67ztl7AVn2a8gMs7e6sJ9RobVkpGjjao4uQyrI7toG3ARIaqOFgrH1OpoxoK7JPJpBDm2O+D
ul0beDWunxsIZizsNy/ofJ2D4wGJYqim1wHWMV/SmDLjLJW99wtp+KkphBHHeHNbOlnd3IvX6ZMz
+1jWrwsx+KDeAjMJKGTbRyAtluvrfw7rCW6QgDgc1wR6u7+uv/kGLkLqsXaYMfz9098rUeDYzbEz
huDR2M+/x1+KgTpeZ8/nQHEFoAvvHPaSV4igoRN8VO/v7VkxRBmsvkBlY+1zKwmMqJx5IJH8qZl+
HEkiehajn/ndnzO1XclA8Bpq7Eli1sWmAxqhGxzUvAhtQ4QmE2CX+w50IqUqjMSNKhqUDMwNUxKy
QT1YBwJQrlP8Yjt3Y39nuAzupcOFC5fVMjlGHB9hiHTkIhm2X0SkFN2mwmMmfPQROWLXuIVAjmfg
n0bl9436clUbs2+Bwzai19Adc5IAS9XBTzEgZMZD8xCE/6HGAahzUMmaUc8Zl1XCGO9CM/0pjn0a
llN7yIgSTDPXgIdpWfCvhGF16vfGhurrX0SGmrTO/ntAE6Cigoh5d6tE6BJbH5XYmEQlz2ERW9of
V9fEiQyLCL9Zl+yX2MDaIkdxiX4eiV+8XtpGhhKaIjQoDBBWkqddH7TLTcap/X35+YLdWq/HtKdJ
ApVsX4jw1M2XBANpQzAa1Z//CnOq90bd5/zETi8VWIiDEyeiE/qlbauyIxwEuw2gkc1vu0760iAr
hWNqIDzgcl/E88C1TZDGQ+GKw+MSWrDSsV/gUqQ1jKUTIx8XKk0t++y9zFcAb578puydj/Z7QaJB
l94L0Fnh4VDsRTmkXii0zOv2sAOMFTFFR693w5ae8B59Upmplk7gtiZwH9dMUc/KgipUtNVqcIt3
CHqgVikJJC2EqNp0Sd5bYvvpix/hiC4FORIVOycc0C7LtQzi1whH6YPTwCbW1ymZtqksjqDESBo+
PrXx7KB/5GBVL+bMAi1xJHCcgglww91t3ocRo1yoeFtFNVIUcZi9WfAv5XcRZivrlBqitOv1BNrI
gBbYtJb5/ZeuyrfaNjqsQ8Lq5motowTJmBIiQOQiwWgSvX1LHqIpoekDSWtkR75MIH0dV1FSjpsp
Y4KbldgSolyg49QE+wu6e/DDnCgz2AHoCgoyQgG25tkbpYYyy66iyVYfE1lnSKMIWJttPt4XXKAl
6bWLWx7moAcbwofgC8H7WqfXlu4eECoszCqPyCRI0o4vZwnv/E85B51/AOGzS1/cL2eGZc8RaAZS
G+d2uvGtuu3V2BpHECngjbIuszf5cUQdyt05lahawjqDIgrv4og9+klW/bfKnJDlX53ekO4d4vgu
mbE0y/3ObKxnqqiOtw8BjtrqZnOUrYLJhtppQqPezr1HCnEJoJQh1DMR5PA9JeUG+r47NL6j5zfB
6nOQFm7Ot49PE5ffeKTozrcAtH3ly2TxOJl2BN0naIc6sX2QGsTsroOwwpWKCozO1Kvs/YSoJGLP
DlWdOevPKl2RJ0MAjWe7y1w2vVU1yHnwe7iMg9d0tCj6wo/XPAGdY0B7X3kHlq7eZAVW6hgIPX+7
5jVAw0KaehNp2HB4gmF9BrIKlHXch1DOOhBku7YjTYxoExD8OLYQXdEftuToF6MvacSplczSvyEH
jiEEcWuHYElWwVbL2BFXaJ+p3s9h2LdTaNQB85RRslgLOa/L84OOy0pOtfP3Qp31izIMc+AeEX9b
MUoCaTqiBo2kWpk/tdYrkE7iNTfxTlYZGkAQRQa4WNjPwGLg0UC5Bi7i2I8aacs5CPpQE4romNqk
IzvssyFfblBr54a++0MRMObRKe5zzuUSD3v2VI+EH7V1A17C7iseVFs+w1Xc93/uzfsWXUJMkLjg
ArmftR2Z9MCmebO81gFHb0dj3nSu0eV0CiAQELxPsowkqGpx1Br4vTUMP89bR/niC1xHqish3rE+
PDdf+26cyBDT32yrFSYG16wHYz1rCGKQmNyLgmQcCsqrmn8TiHWQ/glKNfqEfwDyJ3GIwOFjvLpV
VYChxggExYLVjsG9yPO+zCwM8iUL70kvQabI5IvDLSujD/ba+72WKAvJRLnG7VsllkbK2dbEwS51
ps/ceUu2Sonf3CEt7lHUOf9LYVF9/dnZKNAi2G1BIpmLg19Qzw/bomq0M8QWRiny2ZBrq11FYv0u
Cct8I7S72B20jKRodL43sKSurtaHavCwCbURy7cshgaofMmF/fqvMVN4eEkFGkFIlaYFqp0H/rq6
c/Dd7M2Rgo9FiJoKlry0R7qnDwm05DVFrpssIQZCUTMObj3Xc3lRiwGbtYeIrzmSJgaYZKTjpw7r
n2JRmYdRyzeFQnaZZpZ8oWXVZIfJ//IBA9zdC8UFFgi5ZwKqNBUAWg2NY/jhoTmByrAx4qIoliGk
cr/wuN3IqnZUVtrxT4+mpztbzSSArBDNSqPndKtE7l7DQgLlX7u8ya7XtQw+3cSs8u5tGZyikgN1
BWEpOMvo1pSmzJlg9ZnURxonF9MLtF+mzDfSOrBc5J29oS+y7O/+VWxZkedbR1lGsU9IhQXjETjx
xVC14AaiqpIzr9ZtOp0WuCX21EIUWLsBUFzTfEBJz8Rof08y7Mxs8NOubvJu4LEybis1sE7HmFLP
D4tH64ZtlYBbqQU3JL9TMtIi58f9gZN3Fdcw3oOoG7U1APaGI/adX2QuxX8k+5FJ+mYKHUdZu6/4
i6poDt6MqanwGZn/M0FEauv2EhrbPDrGJVCbTSHdvOirjEmSPhINiSeNtt5KfHxJ1BhWXkqA6ckJ
2mJjgkv1z+JrNX88hBYw58j+wT0CSfcqOoseSMSC9OcmYtd5bj2JvXfx0e3f4wH/daDbtN8MXnhg
pa8FPEFlV3zex3jx4dDYecIaQqHl0/DXH3rwLSKw//S5vPoNyOfMGzboF4A8s/24fbpeaQQoU8XH
34pN1v45jNBTl/KlhX/LYdKvgrwyKEC6J69YtKiLZKaIxoszXb2DWh55v0KDzhz3DHt6fSFUVkoW
P2CTOVhELr2OapY1ivFxVfGp4ZzM3/xaFPtP+5IBgz4sO9uHW6fJ46dmoTGf0/FeoxWdRzR3Y4Ft
lgt5+XcskukXcEk9MgfSnL6maS3MgMe5bYYbUjR+MRwydoaQw1w2/FyrthOUhneqfBrmMCtSL/OA
0b/XFEcwlGxYbk5/TrmwZYNMyuLgskN5q4oZPI8HDLWPF7efvbj4238RRyV1S/m6BeyfA5WJbTWF
qJUShObpIJuazjKVXYrtDNNiQ6R4PJKE3g0Ik+qrLyki5ngA/Jif39IDYB+pChgBG66ItTxmqsKe
GBmlWftWfbVorKNR5Y6XRViLuAcdZ0C7orHrzr2HQB6sFpyZMfMeIJwkatu1Hcl0z3X3nuUokHcc
vqoGkrvXbtOfD13NaAANZp6A8f1D6N2lBasgjArbl7KnBEDhWtVdmtRUQXt3fHEUkzubCvQbAui2
GFmr8fImANr4IdsM24LlIXFcxCXvz7II9tHKBINn6wbBt+4rToWQ/vG6jCZjNFuWGZafE/Ir5jM6
S7Q0JF1HZpvQRQYuPEOZTo2SeBz4TDidoKm4xfuF3dgoHbwflQXEi7WkN3SkWWARI+MhU53NZVrO
SHQst8fD0qraquDPhcEV3MpoI968MvLn3SBTUkhqRPsUAb5mm96tl3VQoWRrndamExdWVPbUu7m6
YlW6RiNEQol5f8+iMoczDrLA3LiNDG7zTITgb7ZswqiA2c4j4Wiir9gZKpiE2NNCjr6q7AyyD/sD
CbwzlJFRKk/hmcnKkQQt8gasHdWManBE2Y6xkjYV73KHP+40BbS51ZdAGmZea6i90/Xz5OlguQ5c
pQYXeMiMmXO6U8dyq3itmsZQDW3eW7IkVJPiRwcHEeae1J4VFWbSKOeR0F5+/xVjW6lCpDwc16Pk
Suu3UpHqNxVjZ4I+dTBp1f+kaoku5fHJJPN9x7f1QkjWsypKLL0qnnJ1SRYfQkiozk6iMxuniW06
pvTD7qKVeJ4FkM8+432U0aPvEsS0q2/dF/ZR1WFXW52rynhshDWRFzsV064G2bo8DzvnhzaxXwlO
ENArwVkrAql4Ne/9W6DpFQ9DvcKAus5kO3JRR9ocPXvRA0bQ94uSlse8di3a2hTfTPU4GRbMI7Z3
hWU6l/7ng6cEkJtazhxsANoIzLgnlpD+c0C1RsZYdtYMaCi0lccTVUZmznzELx8ejmNUHESpP5Fw
WGJIqguRSyubIzhPLx0BNbe3tAi5qkndwZZOBuSFc2eO9Dc76FgxU8WIVtRjsyP1ObRqkKw80yyY
7s4yoxm4PtH9KfzwnLQK71Z9kThj2u1wfMc8PE/6zne24HfgvIULZDA6CE1ZxM+CRTXJxsSCDdYm
qbQRY2nsGwQWLrgBGahj/YSFQLGoZwt0+o2zju4QpglpsG+NDrB6WbKUxG0jQQc1AajNpeY0yfvc
ItQ/ycyuYF9g1b0nce21GvAb2efPfyPvfu60wsW3EHRokfQdhKq0d1ezBZTqu4va1UHSdOPzLzL9
byHJE9xhx6Yc8B3UOVa5j2AeS9HvuTyFy7A5bZiwRZj9xgV0eqTksOn8I2CpdCWFEKoa1jlFI5Oe
n6PHemSKOuvfp0kTa0bUnDce7ZI0vJb8kC9PEkxci2cTz1qRef+8vTr8IWpEBgOkeFUsjUA2gYgY
lVyQWCGMjJ9JSTSrwacb8y5Uc0s8PjWh02k+e5Sh/3GshRj96H1dqhkPSammVLE24IQZRMNVe6kv
6+usrB9LUEGbC4BZc+Wtevmpw0t7aGn3Evvx3a+7mEn84JBkoO6Dj78USmR1CKzarvFwvRtLlzTN
Xxd1T1PVcOUNgZMyshSmn8vaPEPphlMZM7aRVnq4te9VDI3LkPjdD+p1FDLVEB5r034XmJCWAygT
eVxbCk3sgUeFtPhMHColsTrt4Zlz5mxN3JU3eu0oWtLvrtAVZLzWnZAsNplbunmZ/mFsIN7SG/ap
Odf+rSTTLUfbM571kBp/qODl/143e6O9uehU1+lrqrQ5A68nQgwrV33D0dgUAjliYUxpiRIYJQ/9
nbuJx3OmQken/TVsv2bACsT6PrpUS6v+ImhQOPkouNOFZLmlOytGr0yTMo/Gyw3WX3rKrCnGMkOU
GsDKimITyEnY4bth26ceti0ybtVKmBjQ9bH1T4iq9VD9zRw2DlbL8zdZ/QKrGNonUg4cjr9JLvOJ
q+DYooGYCU3zuAFsHxGJsGPbuRpLVav1a6mPXVNeisLV2vlQNgjqiZ9FCULg8Ud8ULWhLi4Dd+DJ
T7XFNAdyBSRZdjYKKnUqL4SxF8vzTTPAFuo7bj9Ava8SNzkmkWVuAY3rIP87exfeepKPApgrsT/E
6J8WNZNEw1VlV//JlcK/VJ1HArHxPh+MZHXaAM87op0IUcXICfeWrGWR4MA+xLF0gwRkaPH/KNTG
2kNKS2JgDIIJsgGA6n6h4zUNx33SQn6HbVvDi3azr/TLeHrFSoTosg7K14ajIGjzk2LeyfpLbJ27
F1mwYydPB0R1pQsshntBJRthzvgio2soO6cOyC9925So1NnXPgijug5Gy1Ysu2qyVs5XVyEDnLg1
5aXLjeBCk7L/S69zX5C8J4546o7N4E/i00DYTmmB0gyblIKEJaMG8Q9MUMEqXTGgm5szBkASHwBJ
1xar3UXYIw0DimYIpFAqHi7J3Y/mKJtj04YMRArYabBAX5UBQePLwLLRGfHfVAj/Kc6+hV2x6CMi
cTvC0AeKBK6yPLWJsEL6Fuh9A7JkC3AyJDUrA6KS76anCvQG87dot3UyyFyrjzuDda4+ITRoC1Jl
/5/W5zz+ZHDZnQv3rn/chIMDsdw5+x3mIfDasazuqpeUcG3CcN7rDspUbXiKVJMXOyJhoOsu8Pw5
jfT3TFj4Vpq2my/PDCZLFmomen22mcfgc8EcqlB/31WK02lmqQDbqWaMJgeGgeet6PCJi1po1DUT
2+d4Z5+TAot7vgq2cU1VXXvM/6sSdkdLkSl+/YjYcnOC9Qr+NPihHKD4UV9kWTYNsd6epTJjTYC3
HUnOabyLqUHxTEcRB/UXZ4vRkursWeuXd2mA3Q5YOpNNZ2ild6pUCXqYpNgTT/fUuOnzwwLKYN6k
zk2C1m33St+grEudpHKxxG8fW2nj6/O5xHapNN4gejHeiS9ONOMM9crO4GRaRkD1f5fr6zCh+5I5
o6zoa/Bh5AvsrbQyiRld02fBm5TnXJqu1MM8R+FSnzPbsn3/DDV2Nc8AorDi/zNHrc+Q7zB6kYrI
yD8DrnIq0jQI/COfHra1xMbCHqn2KR3usbedrmOdlXSlO3ZsLYW03GmkDSi0NzY+Y25+UEIS1d/f
NOYVH8umc5+r2Oqcy8Znbh9CDKnR7VKsRFPTaesXJvrQl86dznZDnO/DCoHl7JLnDh1M3DGLbD2U
hzdJTlft3HjAN52zCnrdzq1iccMjnk8FcKpKXK8A3kT4Lyx1xCSFx/kTFdg/aWy/Tb2R8bEDAmzy
0VXHvgWoq7HvSCTGEQBJACV66osktepJtRc4Ee8rMe4mlsejArMGLaoOkZ1DIb3KUPNdSc1ycc00
/4TJ38OzbMrJBxcWKVxgWaCn3jW6ot4SfA5BAGHJnnnAVmVBjkyxSQBFNqvoYY9SD310vn3YNsZ2
5fiP2k/OwQMqYnoMPE34OYFaTJtx7cp9a9B6PWMnzmICAA6w/oKrOgqk9VJKq21PvL4LoByTv4QK
Dd2FqwuV+oSDyoaP3y/HSnzJIunQcssyc7c6KFQ6ZN1jIHEYLu9IiYzRMGgGe85JV0nk430qCgfX
ekCPFjPVbijGRbhD7oLKHLOpfxqqUffddNekTYlzDqmmFUNGRsGSnNttZ5BZ740reGEfOj/iwDkr
LV+YoFxyEhBAopSoNCJDByt0LmbtVf1bNKUCuLFQBnTj/lGFD+SJo7fFQUIQo1ECmPQPnLRAj4dB
SgrhM9YI/yzXkCsddvQkH/QGOpVlsjYa7TIWE24DCvRZvhQsQzuPGZ4aYK72NhQEK9AZeN8jTBBe
FaWzIY9WjTAl0DRMWGjmJqmcMbofDqzoD8GYW12U7EDDEs/xZRT0qQKRvslsYoNzWmHINS4WfIwx
it4oXgfiBCuxFaOq5a8BtIBHJJglobWCUAi3MFa+htudgKuCJbsgFUFQEiJcYWy4ahJxxOt65I5B
3cPwZ5y/j4BOjYnto7w8+G4qL5420+ZT1OwYPKH0YGOAIHirZu6esRNx5QXULK2bcAhYZIILj9If
kBohV5XoiYkfkWRhxsOIqnp+tuMJVISSoqjzkY/wOiVHZCE4amy3GSGIpAGGYfKaofGo6Pg+lh0U
4TUEcGDX9/Un4RDXcvc/NjbrGuDtLrqCDf80hp1/KavrmwS5qvVlzQSkct6JxQs8c/Sb20O8FQb+
JHpqW2W+gyH5V4ALygGKPiD/jdnPVghC8Rz++ieYUjBkMdwCaxVur/v7Kp7RcC76FvOoNzWSk1Ya
6zTrtDW+WqQtaRHdXzhjnmscIwu+pPDxBysdwxvr6xAIC8qxu8jA2q++XjLBovGFPrH88btBQpry
aHnN7OGKH3R5gfUnNiYRA6wk5cxRZ8LaKzm1u4YP+QtGsbxJtGiTrR/7LhLzvpkcFbuA74UC8tNI
YOK0nCk8iLD3CpnZczpsvH0sGSzwCh8wsdLMzKt97T9lqSAo36uQ3wvlBJVhKuH5pMQJl0iAhKyR
QcdIHfcXdzJWGsEm2dztcMnuxzgek4SSIlQG5NH4J5oSCj3SCaZ+4AgZImmksote77Pvo+zRK2rH
mXoY73QNgTmOme7EVZuE7tz3XbwTtKfEQdzk8szqmAX1CRJI4m1VYHKevxPDrg1glYdP4Ot4XC8F
BCpB4VW8p/G7fEzpF1CAO7EkxDVKZ5B8t6Uwy6OF/viF7IdoTRCUBzr6pDFqVF7v/tE05tvi6/xy
jMkWRWmwjfJxnjoY4o7dQpP9FLww9zK1iuFoCDWz/68kqHrmSF+vG2QX34rX9V4JKjcFl6jbpJv9
b5hM7/fuP7X/MF42k6vdtXjks9cE8EDMaeE1jONIeuU0DcOEzwwPerFyE7pvLaGkFfie9yqPIOqC
pioWL33ja/GIfX0htXuqX92oZrLrK5OnNxqOmIuOrTfMOkBi7eMwdVRVZU4uNXIZ+9m2s3+zuFPC
g2p3/m/uSIQ2wZQnU3NZhQA5qjr6lguWzlx9dq9Bk9BFQnCrFDXXvTQE0tOpoJetgZ+kiOvvBame
8krVCIIkYKsrRlJ7WVucAdhtSOLyXjNdrZCMO+E4KNvRGFRWnGF2xGGC4S/WEHSsFyv4bycreza0
M4onVISCStd3ktL8ITqyGPORMdti25/P7TPlowtUJtZfTWtyjcjz1fkQ4laLWW1beBpos1uYvd0U
MWGY4VwjMe7OFl+W43KNHK7lHOqT+r/ALjH4MkmrAmWMjRe19sK0QRRwQnj5gDVV24Sh9+WWNbbP
ndlM6yq1+sdpzeR+GmtTxUTYhoO5+GLKvLXq8hhbmcvwpMJ44KGFVMp5gT/1zlcKqKPzeMeQTrQH
JaZvhpjUqHMExbQP1DGcyVYBmG6aQCCulmMLnBzreCrp/n0k7R5ypech8UVTgTJuMCOf/14O7wJK
leHH6Ik60TRM8fAyx2pdLB+3pdTlRPMMnL6LKAf1DGD0Em3fjE3PBOTlDaoQ5DlZkAUVDx+vLWMO
cF9cczHs6E448xiSYWRLDdPcE9htzM3S0zfBz+iKY98PD4JKgPnA+GVTgRNyeu4COKDsOEeLgepG
vk3ngtNol8bm8aSoyFF3sM2TrfR0XxTxSHvQfMfv4XFJnhMH4faMLLOn+F3Wpb+pwg567MhetOJO
tT5DQgPY0t+4OVhRIduwRsWGGMB+vZlTsT/ASAaC3AYCSlg+N4yGhRqL1ycsadCPyDEo4Fq52rnw
RrKiQZJI+TqBk66ZqlV3In6u8hIIEgZtIiIngKIEFUMu9GRyZCDL/ji2nGOhJfgo/u3P1XIwSGLw
Qf+Lr0V3gFRiTYal/VI9WLVSgVxZAyMxIKZAzqvemncIDEBbtUGhN7bd3GhCXe4coqLzbpKL1Su+
KgdiUE7tzmwT5bfcQqINmNYFFBWuWxTmf/NxZYqdPEenqEWK0iAk53aBtPTsvBVLkAok5gvDh3UJ
M3r3V5+TenS44K3ZV3JLTIVq6HMBqs5q5frEJ9SWi+dU3abYO7yAO6VGqjC0OPHHHbECRlN/TELC
88gfAD+ZyGAPgjw5Rihm1zE5ZZ68fbf6Yso+xukznrGSXrxMgv8VUd2LdD4qdj218lsnDvhfSpHL
YRxuVn5bBt3hbOPIe0Qkzrpl/6UDYbznyvm53V/6sJ/yjDKaYD1fnxzufoxGz5e5sW5J7N4oW1Yp
gn40dG0IgYPzDed5LpqaLDAZHbIQ3UNQ44LH6VZ/bpbnThZpIISnawWwrB64pxKFG+bVhe1PPTao
wdJ2fi2izmyX4pUjpB85cc37/dPx4uqMZS4A6Fg77E9q+MPoAp+mn0FtILf8evWp/BAzTM25sR/i
/B5oQ7d/Mt/QDADZfsihxrkE8EczgJRPmQfO1h6RrJG4zFfGsjWqLk39jW8ueeJRITTFtXdt/FAn
rfXEbTtWiy5+QeiPc+oWjvqsKHRy6PnSijIJw3MfLiBCxw2H6GKdKAciz6t8SoFZgo1DPtmEYBoG
dnVnXn24fPsgcH0z75qiPr5trYnNl49JgMDLnmrffvToJtXNyakR+QKBzjAlq9y2YjZRH7WjJXRu
WBkB1BIyxJIlXsQ+4v68HPA9CNTeh9nrNKkMZaD6mEHsyRWHRlNQLuN/LpOdpWQ9KbcKh3L3fgwS
m1rgjth4TzEBKUI8eK4/h2/PGGyajP88pHaF3Tur5o1db6XJVW3w14DkqiI8mqxzqfpfXZCL5bMz
MTwr8tsf8vzQvtjm0NhkOGvBPwLrZpCuMpo54Tvby03H17CQ2PR4W0gdVzAhjdDwL9X2J6WTv6Mj
aHIG46c2AY8TtK7mcH5xR9bfG/T+Gwo3FESR2GeoJp7Py1N8i199zXP5/yZglgK5sFDCdLzos4Or
fmpeRrJt9DHvXbzo65iKDQo3lZtCHtIwdvbMPXR7CdclHV3BOZTrhNMtyJBBEximLM9nca9/ACc5
rV5ZQQnerFENdTly3g5t1dbhO6Nl8Mz/Bt8LybY5gQ+hWYTXWc0LA+OFTQvjGTnmS9RFsNozU7mG
k657I5dFSdypQRvwPD2OKjoaMdGgYAaVsWodqKAV9TMauj2mqhS24nW31rwHyZA/B++kcBOTX6Sn
9qviVUAQJFOv8wOpy6XfnVMEmg7VualfsjMWh/sbbA4tOrUIU7cDXsQCbsWw5xHGBvDbTTTGPtQJ
VnBnvDPoO2cF3ptTlIpfX6w2OTbVscjnlXJRNw7yYr+8qK91GfOaeFC1tk3/hThIQzZgaoQU7PRJ
ZED1HREzipA22ueL4g1yJtZV7X2LZgIq46vkcfan5mfnNN3P0zWof3QNecD0ktExpGLB4Mzc8UmJ
1VbKNOTldUjtYc83iwjFpccejfUsj1Gh0EltHYOl6wxCCR7SAI5BnT+/NJkVFg8SA6bOSmTAqeaJ
H26HvFxf2PV8MsLE49ir7fE+rABlLFhdXXU4JZQ6sW5JhwqDAyNCnOx2bVzAYfL3XIGqiihOF4h+
EZ7jcu1/HeZJU6Gf2nK4n8OSrvu3vKP5zLd1tRGFnXf256VgODUdlcfgFQHR6kOIaG17DFGjavKO
biIz92aheRP+XRqbSNvH06C1PvlwRUv4WGmg8qeMwtsFwp8kNlhmTSoBDOcSotH2oVDpH8YcXwZA
EQ3dG2MRwzw+iA4M2jFDeo57lkNnwzzCuZKZ4Wt8AykSsNonkfs7gmZjvEwhULP7b6ygAUIQJ3hh
GoV1Zs6JZAD6W45iP7T4XPBqSnbfI29nxp1dOnsJ2SSP4bAtbdjW6pX2fFHX1VsSpt9aIYMs7DWn
CzVNiuN8noQdMFdNybgQySF26OUHSFYTm3QjrTtF8TEEO0Q5sxgNwG+DfJGsxar7gwpYPZyWyEjh
3enugcUNMi8JxpttnRztWofOOo5ZTYfHm9RCEc1H3YzWIIMSGpBpPmWkx45Z+qqoButWxDkOr6hc
YmDZvlXoT5xGAVye6XLm2MsaxM+vP7xTYCz+RYwi8LX1dW+VdrGZoL/Inl7PJx8BV/b/XCqd323V
FZQYPX28vUEg4ihXb8jwsohgfbK6jXNQ+m63hia5wnyb09/2yNyDYx6AmYixVw2Hisxn0SEh7Em4
/gnPCw4uPQfRtl3vAmdPObpDx4Dasa/eBoBWm0BBLzb/evNpclZa3bmBX7qte+fSPB6BBYSTzYrh
c8Yt5Lrpg287VcKT1yCLnKd7zSjwPtAtsNmJbbmIEe2nSIFvjV+1+B+h3JLnylj0n4KVpMJ7rE2K
+9eRY9yPFNd0JBc6UNRgyhGZhhxPI1ATMPxwcxX+FdL8ipSreZRIiXxSK11JnqX6//zCzvEqpn2T
T+h/Bd39I1y5yGSUXrooZRk/X/25kmL7KE0/eYmbuHTPpTn4W5dqhv6Kq4ibrqkoQDdjFYp+iLlS
5LwN8opsw/mMiDxF2YINwcKpozwq/krCJ4crrUfQSZzX9NAEn972KxErrTew9XKJ1ajxadkx0nkX
cAUBcTfeZq79c5K4XhwQI2sPNRlS3NiFnK0rjy0/9tKp4lpo7cWGge7UQpTVr28M6h354caWQwM5
mAO/1wBVencw93VnyJFDMeKLRR4IJZc/j+yLISmkwwHys9aHQkrXNVUj8oLHHZkvDrHfxJMEFn3f
jOuHQUKtMpDkmoXa1wpDgAFZZC/m1b0220SNMT/Gx/wLAFwyKpLhqZK++izyqYnYF19NIF0La4zF
nWj7lRmPg5sahnwejdwecVWMFcYtR0+XSFamjpZlmoC3T9I57PBthvaiIOBKzKxxpDViRDbd4ikF
38HvoBXSxq1k3wULgWhMR7gvKPO8tKHXkOf4OMQdcOiIr3Ewxn33EcwZ8pS9YZieXWYOGQjFtjZj
uJErYj8mqfwX7lQCX9UzuvYi1/XQ8v2KspxfJ9v+ayzY+3h5cHq0ljIqeEbtZSw+7XqSxgf5egii
X0JjtPoVcReFjYnYCRFEtvrxu0bxNSXQaMxXT4cf9iJyHFd4vBfq4Xbt9sVxAOGMnKUvEng/bI22
ULQua78CVjHOTo64SjsrHIK/Ub/mKjnBewWYXODLYelWQAjchMGJtCrgXxXw65DQI5PSDHu21H0E
x6LM0aETxf22bsFgk/qY5lp0HeoSEOIS1HuwA8cRslylXUwL/sbCb1RCzWb35LO974rOsM8V+feu
7u+qVte49eCzbFfBJ1boC9wqYW0k62GBORvnIpHA5dGt0frqJ7nGSA3WdSWkdmDlk4D7I89XZAlN
ip5qCD0Z3fkhZOnz4DcsIoKRrUWmsiC8kkfgQoaIF4W4L3Bx3nj9qFWlcrYECn/RinW6hOrv2g6l
sug2XHtbubOsDBebKylsJEwIsSDzER/djwPwoPB2lEDYSBzd9d3JNkFmKPHyCTIxD4hl2eU1Tsgg
T66oFegbGs3enW4ZpVmGG5LE6CoI/a0gcw7g/PQU1tO6xHuErUwxP5qqvkVD5/cAAsXjkqxo/DiK
sroywuw1L7LqRFXlWQEJ4I26H+fY8/sEKYO8p00J5FCpV9hT3/7+POlqMMUCMTwtez5YQyIihwbX
mL799BAvKU/kEyDoU4j7wKiSyYOQ0gNxZ+8EanmlJNW3Ib0LQxrqKoW7VDhEAWwCmV4mUtvbi0Eb
UEczsF3Bug6H27eM2yQQcD0l4Lvvz7AdPbr/7hyEoYQsCCUUmPyrs6R2JznaH5lFZ0QjnBP51V6u
vfabl4EQGJJkAtZztV5bD9H/Qag9FQUY2XluJcTKXBScksbzC3y2uZG/767NG+zlqOo/JG6KsWGC
kppDgjb5dehTlJTvb+zvOwF6D33kn33kueu7V5yHN0u36Tjv2uvxPpwFwTiFEiFJi8gWVMFcuhoU
xiZC3TjxrSi2//13SjF4T7ejRKqqxkKG6HhG3xmquZT8MwxHnoARVRXKRYfOnGwrpz931kn+ntN5
AhFwCsIQg/rUGIPIgtKOfGHnbMy/rE39MjH5altF0IZAxSs0GMEL1P/OoxE6N5Q4VNki/a+5VDSN
HimA3CuMr/u9Nks0Sjbsyo/AERiJ9+zF+FtuqasWXyprpMpa9YUUrVyJBHCwD7VIh3rAvmkyJtJY
apBK/H5G+ToioUUqW5HL/1y+qmx7Gl2hOIOKoTo5OEhN0Ukt/aYxK9P3DgYaqHutZqJw35ipCyKh
o1PWPKZaHrr+kGDYwFk/FENuk02oTbVfxvVOodS1NB5bKzTJIz0EFa/+WywWn0KOquD3YhZ3VdtT
p3J0LitTeLsoSL0phT5eNhZPcniFjdLkHXVZl15SyBOCkX8MtD7z9BiX6HW1dUBs0jlyTEQGSoL2
9Qb2GFsouKEQQofBNYkHymnk69Ntm0tlyYt828AC/QwPUjCc80I+FVnBihWm0gkwE9/ROXXOQlKF
L01e/FmrvWw/f7k+5epEuZ75tLe1neUyzrtQbhKqXgxCvUZWByakO+O6kkJLKzPE4wDJb5RytvGV
ao7YTyuXGdj3HgKCIUfzeCDDn/IPXGHyPe/ns8Mvlg0dhg093YjW8gK50vRdc7BfN8fasywW7wMj
D0/ttx+OvihDx3+96uTnVsOM32Bg4f97+Fh6bnSW5EU6lzrKwKEjzB4AjDP7l7zcDs/j8vJTilYQ
GA13u6VB65OJp9Qunf8X8QmaYmPZjyhqMCPpTOF2ZQdfnpgDtr1bONqXLoXHFhzuWz/1ZDAvwUUI
dR1aBgxEmsx8iTtJMH+q2AaOR7rrFyCPSmIKNSdItl0JBzhWx+lB0hoAJ+lOWt0YwY6XGxjFKL2t
4zOVLJNPLQh2JeF+Wr70ZFvy2z2YH0xUDzOy1I1xhfCrCbA8wrS7kg74FT6TbpzzmSe9c66u2uLn
lsgd4TTELaypvJGb9rHvkQXRB+ba9tl9/GPEmD8X5JI9/L8d1cbs0I72AQxM6VS4CH/mfsdiwEoA
wi2Cvd/H+p5xEp6wU8Nl7j6w93kJ67dR9VVZm5j2htEEp68dYVBY7UU8u/uFqZ0LohaIOGZGNzv3
wSz87Al6ruWtVHaXQa5Gz9XdwyEgGQ+IKzUEHDnwPo6UDu3Vl+0QNfRrvT7ODs5X8lq4cdQJoX2r
qBv/ZIt0gQucrsYIDaRpPMj8ExGblXFSNg7g4dhqNy+DNPH7Dp6Pt3r8zY4my3IAjut5J3FomDHF
Yv7WF1HbPeJ45uHRxrbRAHUmUL//f5Lhj39Edbwy1q+0W5kuNz24TTzQULoDSXgVCDYoqiAlwDc9
BvMPPuP05B//cXDbE1UxNS3FLBfjKFwBbjPqVs0dC20QGhPfRjb+pgBOakU1towHY0ELMRzwKxnB
W/LC0NQQckeBfGPLaeQuNeVhBPpdY+GKX/TtDDB5BqWmLx8Tn9E/T5nyZQYKHsKJVUdrz3HlmBSp
XSivbs3EGeTfNMVyOIrilqbxdRsjX3iZMGfteZi7v5aMtAhruhozDC3gUKWL2YREJcCsFqd90zzC
OMUh3G/G9IeoBc7j9nUOZF9jZqnu1+571oC5/+KU/mBG6JngT8dmxsgrDrt/4mCD9hImonSoZqGY
CmYKFuin0zx1PFmTp70CVudHUj5bRUP721q0pGtg+Ucsati/gxt5Gr5lZG5SXqvgXg9be/3YszV6
Nh2FltVarSMe1Sr8XLEt5dx1JI+ynistEzboiCKZARqZn7W22NRVJQEyEN8JabAdh6WQ1ieJoA/p
QEbeOZYrgQx9+st2isNarNCfyrnVWDWPdB+8DOJVnnKziDEoIfrUYidSBCaei7QI/yTUurynb66B
9CE1aNteLXwepRpRbK1dzsCDMZV+hS/s/QU+MUmmWUj8UXEf813ylFcDx0/51qKXsMTI5e5tUdPT
ZPhCROGBT0maudF5rafrQV6k9BckyJaHqJvPHKWlGkxqgg52S7E6kZMN8xb9iyiazQxzGcYyVP0e
cw+JPd2fQOp0bDtsV4kURhIIaTfKH/jkrmgG4Lo7JJlljnOlGmJMohgmgeWM5stWPQntHJarplqA
F2sJ6x3dTpsxU+0mgeosFSyfS2p6of+Wv2MX+eNZ+VdANXaU1mi1alJpg47SL66m+8LV9N9J4zCZ
ZJ6r6nsO1c0JyzdKGkESOfgqni383Woo6pV4JQKCQsgCGPghE7GIGUYS4EIQkDdU+ONBe96pKj3t
3iA8GAoQ08lOjb9Jt8SCQ8ca9u5XEafhzulfLPhItMR7nAUPR3CvssWjkNmAzcyogbTq3QB/jkeV
qwgiRh/Pv+4TcRy5ltGxq7PMJoYXdySW817Cx6eYXYmwtoLKqjGVGyTPhcNLFd+Gpyez4iM39BkT
ibh7FDWARUbzf25m3tivRHwOOsdMYJL2RMM+cyUPQmLpRV7AHbG6334MwyqTHHqRJOc97SL23LUl
JDZgEDBQngSx9eHgv9SJWAtVfe40sn7vouXo+6MQIy+KTFxzbiRMosjqvvdvWRin4jvvwzSswaiv
5w6bzEBnyBw+bHv9qN3pHNYxpQAphDfwzB6D9R8nuPryn83SN0msmvo6ZMSYiBGjHrI+1CtvH2D8
Pz/gSF8JqJUKk0aL5XtA4iSuvu42SOJpk5zlwll0ESP05XwR+XrLhmUhjBm9BnDxeGNlrvjsjRgv
EpkNFUoyamyXNlDsm5tBZBg0DsljThPQ4Gn8XTSc5KcchyrvfF5vhw0dAumuH/G5mbf3oZiqtL2B
r6PXgsPsoU0fug8qUSqJX/QuViD2PWVTZaId5Yc2FQTw9DktGSM0EAN3kJ+2NXELYBv2/TCf3E19
stDym6WvLdl1k0RK4GVNFqp51K8OPBbt5Olbs8NXX+yxu/7ZF60WTYMOToOWEHaOUCf+cfQI42pU
sKbesncEZv4Ot2hySQTTWg0RG2Fh/wyfKlu/3jF9Y08Pwj/9TxAAPbXL8CNQaPZ5S7Z+hwpb1kAC
beuw+2uNPJzmP8YU6InkyKp97gOoPLmTzhRv+FhKHvBZTcHZZYX7BC5ZuJi/RS2uhMq/I+RVKoN+
E2oOkdNEyvX7JfEacryokU/fLgNG2mA93AA4F8q6nRef5eoq2pF4iYxH2gBNJVJCPSNGozej7yKn
isRB+RB9lo8gD4Go3zFfSO2b8yFsxIDSvxspu/sXOn6bOKTfVHb019Vw+n9Q5RyMHLgw1jmvgYnF
nLOjzSTuknlPYOXtWA9mVxwfQQdMWEEF1//YC4AHiD6PIeGpJJwH9NTjVHzPNHI66Jiq8VEHQHaI
6JK29d+8ChiBj/2QKkfFOPJhyTDq8nG/ThQj9jvPak6emWaezAA4G4zZs/r0dhb/HO9GtSMLsKWC
6lm0eUCUESsePG7H+DRlrd/nwu9zhskXiPRJ5GH3aoSp7LhUy5pGNye8agps7/zoKG7WpHaHJR6f
R8dAePGmtykWb5Rl5OkwmW5yFX4z5hKgZRf1vXZdjEvdMJJk8Q4vnQL+XFH8K15NeORPSECAJP8a
IfrBE+DX4lC3d09h3K4yNVETa8PE0bpuwMANlOZLYK9vh7OkZz8R3HzQIx/fHbsEUYsbbXyKh5t4
uvLAmF5nNfpOPq6in/V2kgqcoC8RIVLFuja2d3/tVsUViL6JzGKegVQeSqIpb17QsWDhtxVJwINn
J/bNf5urW2tsoNm1Tc2PuEvKiHvrWYMBFQvMjRTBLxQG+vJCobIgNs3ACrlXPy533XiPqLvxnWX1
HR+Su1S4eUoDAg/T5eyVnoNJX/GB/Mk8nyAzHf6HI9EXWkXbDaJNy2gl/ajlYtjqtCyxO5XK0buE
9dr8ackNTIyclk+TUMmpzFMxeaWrO5uaBVx8YHcwrlbHPar4W/0McGpf+hUaMCdli6QxlT0+Yrzz
aTA+GMdLym9gWGooIJglyutVVbXLY+Tl0JQX3F5p/H6AnIeukkKEvAckWcsvY11ixiOVfWnKpzI6
REvOizxr3CcoJOciEJIquSB7oQGLNgBB4hkK/0Dq3c9c+I3CZpSIzs/zsGeuztutIeumbvj0EViE
kikkmsjDcvmDd+l4vvpkbRl6myGrnALAMQkq8rQE1KcNEIQjD/6maXxKPsINnhVZkWZ7LujWFKjC
bsf+UH2HIZTECfGZxdUOA4jqAtVgR3KNbrda10PlE9+eK+3novefP+XebhwefvVoe32JFJXsBcFA
8HzQTLeRVFas7wv4GqvPmSP/XI1eFnaJejQRra0n0q8C/BPXfHIKm2xdqgYBJmgVS2dYKCjN5zEV
NA6tCa0C20OmDIxbMl5nDJ/IDmv0z0tTJiCcXhaSUg5W2Z/zt0jBQWMkR5l67u5ElmDXlmygF3qf
/praoOiRN5EBEtDPyT213e6GXGHr+F2jHM/tI7cgY3EfUE+z+ejZmnGZL8GOev93jFFL5WbtQCrw
YvujLwFBg5A/loBP2l2LxoFldA0ihFVpCxtBJQQjoSggfeVJOHYHi5JygZFMT0hQ0Bci3bpdnJ/i
CkDfotr7XCzLjVX8b3s3OXmVHES8GNtOogQMb3YQgjLm7m0XIjWyzLqMnaeQH2XdRMzebJWNlA4w
5N5QgNvqUF8v4YRFpZ9xuGaYtuVA9HPDtbwqYJnw00ip/a6ptFE+hy8RjCGdKVbO3i+HxfKwMwVR
hUZuLTCZ2FYSRQr7Pj062b3DaCW0cQc3qLW+5cLEexmycyne2NCrT6D+FboNgpnnp/NPLTvPKLXE
h9kruP0lxdCN7d0zp5FdXPkpDpKVdZojEVmYlXVuf8foH9xsfe4MbpccZxaGdnbt66YbiMLD39My
OrPZAopnn8jyZOg8Yj+vHNGEwBPOC3faT+QTropY0q98nu2hZ+DHNF2iQ8KGs3j8df49KSOcZVg5
wNZaHrgahAl7tNFF72ewBHwj9UI5qemmmBhIIFcQtIvCGuUzzHWhR6xtC3koW6FyoyStS6kpvV//
6PUNMm9Q+sRynT4FrS8S6oa/0FVSdAvdtLVKZA8fuHGaWptgFTKF1F5fDKGTLy0/rxfFoD32vaqG
cEc70ljLr4XJAipxcGh8c8yyIBBoPAGYegbwIxpU89A0wmbL6PqwWloVWcvHYEUhxMb/e65HKjwu
Cokj9g39rqDnlDGHknC6T4plY6/h9qXDMUjvEP0Dp6C0Vc+5zFxr025bdbAvMXp+k89hfS/tA4Yp
BqxH7p8ZahaVliY/m5USKKacWGia6g8hw2HCBPU+nsXKid4dOuqHfzD2YYmWxc8Q5dgQK9fA1KDw
gURxkeL87e6ddjg0yrjn2bc6GiNpANOicMKD6aeppVrxcvLM1e+Y76YQyxxbE92UzTbyNINY6zAw
ITiD2wGKTQjsRVrK7DvcvNvjODclZoQiguGOSukXbCJroG52nlwKq7gfm9NszA9WuOU2ynUD1ACW
xNbXtNdhy5mskDXtkJ0K8qVCnn1mFdu4pUmTc/RutKXg1Jja7CScD3gZ54/AlGtme8Dw5+24FbL0
41NW63LN9Ogo84VOO+8QlzTjYVl+CJQS6dKQMAz4CcqDzC3YBZdGYJ9KUUDpzOqdVTDo4ioKKkxm
Ubb+gb4sat0NAgyNlCS/e0sB+zUyqp9IGr3Bx5OjLQ/h/liAV7uKaKNkexq//tyz+M5Vn+g4EfnE
VGiGIJ1iXUpDmDt2lG5/DTBGgNnQJXII798OgA/CWjIqoY+KA9g1U6k4zWmzhTJcZzw4B7szeB6k
FTD/dpX5rdmEqN83rtwmYJgWHos+YVL08DpzFXTaB0KBA6d8iMnJ28B/l+GBs7DYTfZrvP94CuzK
lFKbw4Kgxfq4Vh0tc1mH5QAB1ZhtDKXCSeyYmrQzyoimSERnk3lH+QqIcI0nwEzjZDKHPc0/L5HP
71Qz2+Wz4P89GdLoGRkEIVyL7L6O6Jjk5Cob5SRwhacudn3K8Ul6T7y4qAg+L5xnKZyiBUHAnaRM
6R8FiEdnY5ryf+vzd5ByoEZiZa+2QhCvEOLZckhr7kOl5BT/gxbVPllxk4iEOk4BRbHdNy32e24X
tvKNRSYaz14lEq/RzTWikw4PUyOS5fxxMaTUg5kRoxktLxESHAK3XOlm+GQP+x/SRY02SUSdO4wj
lZ79KFiGmWzp7IUH1kt7qa+6/cLdJuVuoWk7xdUXcN+izksKWFgzrSm5d6dnzgw3Fo8rvbzWkX8/
3aashtLAWMHBt97vdT73r6PRrQtS7PVlN1RSUjstfpq1HOeRrWdDe2lMhhSjewJ2rc1H+zrCr37y
G1IfMSoUQeDZ8EcJMIYAd4tWjFyQwqWll9R7cGI1Hrmoe3JjtPXen1OprD9L37TZZC0RPY7z+vUx
zKnJnm1SKI+ybP/6r+QD6WvX6gYzxCpO29RFg1fVDSlUe1NgrpV3o6nMUyBU11+OQhpcsZsCqhnv
S2mPld5yRiS8Uz03L1eNR8LIECCZa8gkMijYnGdcyb0QWaOAzBDcbgTIUiO0PZaDRTRa9SenMWLl
uFqAxWYnJ7UdKLGJANxeFnFR4DnV7SFjdLETi9uC674Mwb204nI+TpEnNxQhaKJ/FF5zPph3XKOj
JbgFZRpXfk3M5FBP5CjODTzcB3jxU2mknvtWHj2YVW3NTwJBbv+H1DFPJzarZ/9mf0lHCjpJQbxz
ox4jLhuiH7DPnntUsItPIEBOLeUVTDWdv9N/+gy56FxXfQIz4MYtshcZrQz3xUmfjARsKZYtR0wq
Y5T9hJr4eGlCo2eRB9aa+Fy1U3sKF7Zy2gEC/wUKO1v34bUvx7JbU/89tIpkpGRYJ9inIMfC+oGQ
28y+kaiTgcdt8tJAXDjxCYFKadGkeBmHNjkHwd0bQLMPbfgUVptO83jM3Gh80mpFptjKOFm+Cmwj
jkxEB7yrDr7PJZoCiJcS5dYoxaHUwAeaBO69+ExgIizuuSwM5T6HLfBNV0mwYKvGu6hxTp4Thzz5
OECOMZXylfrRCkfBsSlSPeVA6AZhPzO0RK5Jm0Ev7R5hpnXsH7+pMMrMdKsS99HOFPx2CcYAHBfL
juub02Fhq3fYiZZMWBHlcHEEBohLx0xCZ8C48ty7oglSY2823L6Mb+3OfoWWcJqubo30MpX6SOyd
tLeTm5++6xYt0rv50bzFKursvvJeG90DRSCjvWtfW0Qx9+avBoueDDWT6x1K/xoSBmqtEGnQ75nS
+FBOJPhVlVgWeFwr+yKUQDUgtY2WSNu9nHJlUWqo21+x2KDXDe7ANM3HwkF2L0qdw2Q6glDMDzqO
WVgawm6W20V86gqZeO6ZS36gu5b1xbgZyT+zlP4GYadRreDlEujl4goTttxH6hcJaPsKbhTe7t6v
u9pDEwR83rvCGcQ8bc/+la6W/gtS0dVzNGEw2kj9V78NWeYrNq8rqhvow7Xb6etcAJ4jwtvXlkjx
PGmFONrmXATETSxe1UsLCGqo/mluA3XDR0qx9cAPSUsdV8VqiKl8goh9YU04Wq609tICr1psVHOG
yZkutRyiWUwmuV/4JbjwfsYqZgNVRaXk5MBlH+/R5xaY2gnfAmBzuNkm0dy633JWKvntKs10u8z3
+ie+qRMGEaFSFnXdrrdPNv6TjTh3R8/Ch/bIPX5IEUGFr8kM8kgrudFrvCO+8V1bfHdzdp4CSgsV
ulxnxzHx68cG8dFKFRjJ19Uk0utI+PxJQ0SulwkTVmzXOuS2b73Dw0byL57FBXCWChAyY6E3Uw5C
muX/Yc4XswR9rtlmvxr3GrT8gCZV6LSjWPXabSRGpH+NYEvYIgPwd8dpXprhVzJHoZp92XWfqUOj
ZpHu4W6LrhaseXBHPId6+kiEP9w6VU+d25Y5I4qWjeQeESjRTvfvY5HSq9Ik7FbgcAEvgxqSzjw9
Kh26sau/ghC7xLqDDa4B2G45g6mLg52zgWHNu4fzNKkujgmCNNpc7CBGaZexADnmTUeZ9yQkQaSn
sixii1+0s/WV9oCAb6lDTrRX4uiUJnoUqr7sM8abzFl5I/YQPsIgPJsUiVfAwrg9ksZNDtdXm/ha
AjgIq627G5rJG2pQtsxQ12unO/bJABy87GQlVOpl6NTPHc9pUzKFHl9AWnCUMha94Ok2pY3RIKQj
47RxqhrMncBznn9Kxiw3jwrfXSyHHvf/VXyXN8fYDhH6Y3ikRBnCkVM1Ca+lJFyTUdTa88pOfvbE
6FZMX08m2uK1sh5FycD9eSTsoNMVsOwUw2rmdudX1Kkip2kidTidtwFpC5s5B7WTbUqFhtwxygUc
jwIbNtZel2F2mLwfdZYhm2AKwbeuAQVEEkOF3wAJ77k4JfY9GJRhwkHiD4NIQyBc3xcFgKkTx6hX
VsCbzFTrsaw1RZOxTGUJtnbLQIug/TOtbRKTlO/u2KP8NZ+r+2IxAhQMvwlv5sCXacQYaedvreLQ
W89g/Rzm7bdwvbTZlHHDONlYa9Znw7hxV+Ac5wrMYyb73BcwPkgh7ST5uSlknhyFOxZuoC5knQmL
j1rK7s9Grcp082qAO3egA2OxZnOYz4CY+50g3ucS06FHJBIc6Tn24eyC8bXZl16IEf0llhy3ufvR
Dy3CsRyvr65GOyI8eL3e0YNtPBW9nrkU+4Vo6hvKqdvCoc+GNdiyTuk1ptrK7ETswzpgIPhm74Nj
n+NUnzqrKlNEV/Zzs7lA43pfncZ81GzNqYvwpiBB//u1eY1rlhiKmK5MXK+xMu6wLVgerNAthPib
FnF6E8dscKzEgIVszpHgzbWG72DuPt83jYTGQo73JXOV51LR0dHqLHvqIMrNTYRYZOyB1JLwmzxw
e1q+4Om1/KhkSgT3G/5rujf7/dWkF8PYUCCCBKDlmrcOHBgg7fWTmssovaaAIsBXlExV+59t1Cse
sbq1ftelMSpxKaK6s9vdBPZblGxuoEiKl6cl6ezxSFjoM3cFdohI0nAgXtdG8Z48zrAICYGbRZtS
rc6yryO00oEZshd0p8VA2CUBDDZ7w3Wbp19My7ldi3QeswfSIxhqWjtCMa2sTuUyIwX7jEtOB9/L
zqjMIQQ9qS/0jmq/wnlLhhdujDnDLWvCtsFjoBctXHC2LtQPJ3IleGngHnNmgIi9ILZ5urZMiy84
BxNUmg10cyp7TsBysCxycwXdOPW7LpDG/NGChcJYUlTzehxg5QCD3AtexmNHSWAUxjmm88szWKA4
Gvw5eCn/BdgOrba4b3zDKsVDdykBj8qo3oJVUTVskOS5Z1o5wHNMlBLrYy3eO6PeSDbRrV/s35HD
V3cxdE133scFNrfAiUiv/k8+GwtzVvP4YAHiP4KdgAguKr5bEXkgo26kJt9w5AXSH5LTp/ObM3gB
nswkqGE4i4CT0mLhJ0j7Y3iKkdAQjpJxQsWZ+5eun4maVn06tmxlLMwB+p4VNSudG6mSLlPn7Uav
yyZ2GcmrLP7TkEaOn1AWtrkw3z5aWL4sGDFvOAou5CKQvPSpHfjYS2ukdYzLSIuuwedaXEV419k2
3jar41BZ3Jy+aRRwm4RJtoaRppvcG7dog6AqeS9gEE+heruORwd7n/yTNtTadrcFhM6SbCw8mVPR
9fOFMYPYLZm9FkfdfsyGwTOfOw3qyjBXZIdUrbsD1XLfwxEYHpjHM/OpJJzH0ru6ylF6JH3VTUbc
KNiiuO4nHwNrAHxa1/Cl4+ZuC5ImlfypSxwznjdHqCJOCMfh4wKAd8UmyfHR/vTJC6rE4wW0fHbI
EplxQmoTLByH/3dds+iV7b8HIzsNOPtO/5vk/X3Y6ZQHyFpless4glrKKJoHNE9E4t3jbn4JTe1S
RYxp5aW4BchPGzZPoHz+soPCPBh5IhceaLbz0KUGzt8JdVIqCSfy4fGRnPycukzTE46W0TqpdH4T
Z7le8IwNsb2Kb9dFAdDNuDc14I64V3bP4SFsWWM5/ivybLEdLgC3tR+xvaZ1SDdL5kBWKiU5mFAF
8DyzGvMsSdsMSZQ27cfoDX9B8c0CA5+H/A+hZE0e8AwYyExMZdmK2CnHiTZgW76IuOHesGLtAPtc
BW0NZIx227TOqlMUMlH2NNxPBAkqZJ+k2h6p8vMQZRdd3jajUkKDeRraISNkNmyfO17a5vv5G/ap
B/d/kQLMnWO7+pvS1BXaSxmzMTABVZ9BW6nkbuspwgeprjP1zFdeEHpWrtiIpakqZytMmVUUslyb
gOjrAO7MuqNZ3U+pjVRkWMMKaeaaJ0KV2VZacFvGUZpODMBZsVMeKxNicvHdVXe0O4pPlSblNZ+E
3fqL7SSnmb7HSpTZJAIKwEESUsWwdf+JpbqZtcEi5OioMm8I5YQpIhkQIhN2SWlGzFA8jr6IXsxt
0O1syR0pci+IGpnoDM+1g6S7S+TPVcebP7e4zYSuWASDonXmFppGRq5j+AM8bQCFrWdSMCcvtctP
YuMPW318QlEE2wtokemmlu57AdD/kals5T02T+8KwSMjLdFueuhCQ5zbOJ+xXATX8k/0cwmpIes3
avjx93DzfYWFs2aepMlrB0XM0Pj2GgkquP0VtLj9J9eyPJkfrJLXYS7XXHq1QHNmBx8K48m9F9Q2
qisqu9MgMCGCPvlKLs9AxFDo1SYBrDMwbhcjtnAaGU2tdNXFzNI8XPoppraa6qiV2mN7fMR+F9LC
1Ykj5Kebq2ipt86uwfPpqGWbSqrVk87Qu62trpbnZ7W2QnqYdf6XTtmXQi3QxNHGF7+/tgy/9Xbb
3oYUZmRsRkJaYSo58ZcNTVpq/Gx6D0ifSzzwsCrk0bEmQBOU/7oB4JZHrmlMAwqvSSlROb/JKU0a
X11HKfiUxfLIXLE7F2fJd95q1jmFq85TT4O0OWnl3UJT98cLwL9oACXC8q+zS0Tmlr5UnPirdKXi
mIlfhMAHO5ztQrUKvIB83tY5qxIhe58Bd1G9+ccPchz8p2ZdsoCtMNfiGZ6HxK+xWeTRrwloknkp
HjKPf6TRphGFfVCF9wsSlK4EgVx7lWTDPp32dRmq2HlzUZgHz54IjdRUEXUGSA0IzECwss5WJlOa
0InAryLyETTlo/On2C5Z+czQmcRuxKwd/v6gnh79Aa7H4fPWxKxpqvnBSiwaqI+h1d7MoMBblyzg
qpRdv9+uvjZZ/u2OYWV0gab5i5hAscm5DrhbtZYkQG7RPEFc9GhJLuPCLpqNVJtf4W9JskQaDE3N
DBGNNohk0FW5e9UyXsbxtd82kVLt7fwBXgECWqea572ZeP91uZ6e3GCt4PQLWlr+CAw65OemP4SE
89TRZMmrPFNqiPFTgO6RDUr7Z71GIbpsELSOO2/OxeA7n4Lo9dcSmL3+9fzq1TV/FF0cfXp70h45
Z2u6Vu4OpY/9DoD0N/PduVYdakTn0mIM9XlhjNSNO/C1CQC28sl3QliGG5CRIhwYtxgLvxXTAAOe
sEu44j714uuSKjKo2xgNoqW5Lowm8WoDutlNypuF7fEyjBbeWaPeVHaZ7ZzpbwFsnNBV4AqEQSEH
NTrSitLtRaSGI3sibr3YL3ij3UtzSVkF8CqYVlhacsefT2AyPQ/CYQK3Lp9SB04Weotlv4R5heF0
8OLkGCPeK6/TpPC3fKno1k5XYuaNDC6T+7PYliPCDOYxyUrJKcaL1vRr49GUiTDVM9FbatAmt8P5
RC4FJSpAYntsSCu8z5eg9Dt9aeDX9kPO082TEJgCuzkqRjadKq/5yClDv1OZK4VD79TjLimAQMjB
9jLCxjpkEm448WH23ukBqYmVOImwxxIsEGvrZVkNoGabjaoDoinr4ZBeOnnyucCmxtmG5aOeM1A9
lu3fhOPWHroHllJFjqsHIxq+bgH8oIXMF3BCLK4rirpED777UvJ5QWG98xKtiya7MyBBXZQhsxVo
KoMsb67w/mkhpiV4V1k54/gPx2oISdDBj2NIEl0LYE6iaKf5q0EzEvvNBP4xoDLpz+eHp+45MxpO
B1dsbSzSkP7xy49xWfi8QGlhsqfMVV64Im8ik5ivqyq/JmpTD+EherYC+Ira2oGkv23NPX05O6lF
UlVcp13ASqtjHgnWwjj+7/sDp5cyGCULQkmkCVgOPpCdMwipIK04EsEmwmXqPGr8sNeXiLyY1HW6
jcb3yPqwNIipOAfwwgnrahM7yLrEaehJjXG4GvBF8mPYVcOvRiQfiU/9L3Lmnbukf7Pkg1D+e5nP
O9jU3a7o9d3FRgT0uKgd/FMq00o+sY+DImFG6M+POS+oTCVBRhP1xY+jLxAXNiC8pXlUqU2umAuf
NHIDGcgKm1lV1FRIcXgszZnyXkRYG5BQr5e1+RYIk/Tww3wmZvCuKOj5kcP8+cZAykKt49q04M3G
EsdRVaInZ6qSXaHbXsOkklSTEFYB0i61N+mCXK7R4LgKfVST01ou45E1kBIs6AKO3Cvu5GplH4eJ
IQa251HxyWa1y7hxzftCqjF1UbOKtazgh2iQDI0adT4Ar9GoLXgr1+DRLJgkid8jKOEOz4JszK1Q
/rAwlpEVF0L536ctPukb9ApCUXMSeIF340+zNPXvK8Var52IPta/CykwBpoD8ffvKUZp/7xrT4ST
H1QiJOz2jzFrUUiX7WTG29rXNBn7lEWHAoIsfE2wA7LA27LSoG+84JwsVhKfQWHNNswSCGcOCJEb
qDb5Zxqlm6evr8iyWiar6x6rPJX0zuJ7HwN7HD8Li8b8ejQT/D+huzEMJ9CYEG21ZzZVd1MGGNRv
SMQZUByNt79hl/gdPsLvUy8uMm+YRP3XziAVGyhE4l/ouVEtAtr4liv7FvulIloEKkcPjdoEo2Ub
VXIDcSzugZVl8MNeP43SmhnJrdW2i+dr3mDYpCYT81Aq5UCGb/dhHZUbYssJSgZe/SW+ALjElo9J
oKcWKwFhKbdLr8j16JXLIqMJl7mIqYSHz4S3Zkx3v4onvOPLMyoAkCVQ36GvoH/tBssdiDvrLZjI
gfCqbT4NkPzHA07sV6WHzICI03F6hUyFdNlMnALbjlVm+H+zjFbrpaROztKoFK1xiVLQGCXgYsB/
Tdopwa725/4N39JxzjSyJjtZu4HfYGtK3qP5Ym59LUKqTPNq5RL+p5hQLfZuAFHv+4nHvMnXoKmf
piNRdjvCfooD9ubPlWbDpZTZgnbgSn/ytSMGt/QoUde7c5QsXzlc2tgvVMbVQPToxGdzT84H3vsx
wH6/oiAHF3ZufZdQkLKd0jJZEgZ3bNkmxio9g4k1Fx1GKAJOQUFTyl8+bjnc29giot2SHnMrBvC0
SFep4IzRFS67qQwU4eWZJTwjSKX3qUdlU2I5stko9nF/XkooBrr3EXvmwUEoqYiRdnpFuQpfl+Vm
4Khm4gFEcxdfKy2rgqn0HfbH1KeugxK/ZrY7Kh7TXVu0rKQA5z2W7C9s1WTO72Cigd1/f9/d3K9P
EwJGLyghfaRZEbJGyy1VHNe/0vAtImHntnUSuKlOZLJO2KxuZVDt2vy9+gnS/obfXrTeLPjC4nRX
sYyo32M2XBnfgfLLr8rOEsI6o6QSKVlHZk4x2soD+xui++upjsNTN0WbclFiQD3DfqkpshdQDW9Q
b0dVxK5aELHavYn3EWeT1Pv0qOYSWutHjtvl7mfztx6uYcrGOpID6CFPYxbJptK+TmGD7eyrXdjG
fTL4tufeFjh/4mZhBO0qcG9veI2Is7hOjO+xZEOrmiCoWv4BWctjEua967wby5LD7csvcvLTSvD/
eY3KyjvESMOxeilTd3UtZcul2S2ZLCoDImqzvB/m7wV5Jpxy2luLi+vQamFNNRPKS6j+FAkFhJiz
rWO084F6lLeBLyblJap1qIKuZcWaO/nrXRx17ZhY9RB94kiDL7pP24VFN21BsTzlp6vT4YTabH0D
/yzQAQ6WKv2OPrCuMScwvIemnku6bqQyS1qTT97zxo28GKRClYWbxP/gnP3PvslKEY27kytY/q6s
qoYWSYrOVE0Nu/qYqw0Wq19y1AfqCX+V6/et1CKOmfToVOc+jNS8/GJqDy0xVKpywQxvd4Rxxv8w
K1SOb5/iU0FWeJ/boTdGbf9+7FQLki9rU6lLjoT87biOk4ZlcTKZQJnsh/mTrVrPEjfG2r+Luux9
hL7merRPFl/maacWUOLR/Mzcj5+smDcBERe/yXL7Nt1xIWu0b0adxbrDibjXN8MVppCLgkqS7F6R
CDXswkUDrJ0e91XPK8sVusd1WaQDXUc6ZeizzZBOOzhQJo125f3uTN43nhV8n9SKcKF5M3YjoLHk
Tm/5hoopWv/jpzwkpp9BP11uoJs5vuBssJdGIJ4oMpgI0RHCac84Ic1vo9fEufcoNzN/2lfyC4BU
56CklRwXNZgv+beTrTuj3BhdwBOK87rnzEdSjcXQzxtI5meT4PvARPGW4qGmSDrO9S7aCJM/4san
GuT/3eyv8xq7zxv7qEcgkjSOvKGVdoryF+qYJJv7ta7F+MoHJx7GBCnvPNlofr7yV2wxKd7dRULP
OYJP2UX993TcIjwcf9hw6xzA6HQGhsMbVmHzryttL55SEnlgQ+fG9dtjsX+XJQXzG8mGvi4J/3h/
hoZly0sqc0xHhpS/gOEhEssR4+sTEJvHO9AkN/kXf1pJ00j1LDigjiBaY7BPPQLvumIyohxPIgrW
/viR122PJ435MUr2+imRd6UVWx7IdfvuKp4YjMforyb8WaVmEt0qgBS3ITv8SgCPSVA/+6vldXsa
kSZAxsQ7cr2Zu0yZO/daxcScV/T6Ud53SHPwGM13dr9lrYqrulQjwOuwuVL3yna1+fROjfitkPpq
Doz23SjDI/zOinqa7k3XMkZQC4Vf86bsrLa4AYFISdZUus8OBWj44Mh+fDUEz6LTbgnxtrB/gvQA
RmEDo1vtsTRjulYF69hphvbIwnnBccyBcVloWolzckk2qb9OBMp+4c5igx5jJPleVhouanyu8fDG
D72OSbmm8dLS3rWVpkIZwBOASm/0ak3B9QJmLqQH7LMDTlTJLrgOff7SCLNCUSV1c9Fo6KVjT/L7
6UHSc9kXK7Du0mgBeSkehZ/ZPAqAyRJGhwEEYlSJWzKy8YjTwsYQMdzaIvAw4FTeXNJvWcz5fI8g
7YnPX/jL85I8fFmEI8TJMQ1Ap6drQgsOjqLdo5io8gmb5lgeVyYmGOFAN1kmXKXXY+uEZsptC1zI
Ejz9zRHlMzVSe2vrxJLHv35M1JMgW2R7rJKLu2T16zp+JYG27InC/zDjOfrA5qCQQoKenH2EdZdW
KYXPSaftke30Aqo9iJ5dABj4C0Xprc1Dp7DS6JiIw5k34VfQTsQ7b6EAwV2fEHYB1sYr6emi7c6u
0JeKAxv+6M5L89qntlzaAIcaNHT0dIIorenlFxC9YsYn7CiS323USCQ5VZLO7jAs0QY6Mlns/97C
+Vwa+8N18WryeWvzK5x6yNCeREz4pYaOK/S8GOhletQbf4ZDaE33Y8KMk7Oi0H4BLQlhdDL24ZUP
lBHoDvQeYrRdOMOLLocXgDnwfdvLQ/u9aTVD7HSNRmP+MW7XSLt1JR/fJavaUChIAQMT0KrWt6GZ
TwOu63kJtv19a9M786tmm3pyAkVaxJXgnIBCynElsK3qc2IzEkHA4oP/tnJdZOTxA78Gbren8r3s
fOb/yGg3zTcQqw3S8FlCKdNrgymc/mW4HsD0uvvbgR/BUygrmqqD6tz7Zy5BGgQtp0oQ935SKKmH
Ic+Z3FINqV1P83f34idi0vJXWfhXgxxnEi0nTWmjUv0KS9f6P5yja0wAilFbOxbPHlRw32mRKkik
f4VvP69OdEoyElF983/fOGkzJ0FO/II/J7fmao4OjyNW3m4ayHSwqT2Q3jgFsOI3sxZafb957w9t
eNdyfClJJ8a52JEu0aa91EMQX/M5Kaq3Ocmc4u8WGuqtusJE6TSbKrN1DG/uPhd1x+zu5BR+gUFY
qeWrhnxBTN9StAie7qJSYJ0i1b/nBcERd/cLIeMKJctQMrLRIHYZ51e594TprO/fn+LUKbjVCOTB
TFqCkB1jRiEcPX8BSffmoX7W1CpvJx+QKI0OobwR5NVwHa9Khbb7muKL4HBTWnWIPKJaWKegN3t0
lUBv9G4Suqwn14Yd1zVrNaRgNE3B1F3pbEG1kZvxRzC9uDnCIp7n5zMmR3sqNLHatiplHVe8qnWU
ECQwu1DznJpDeRcL+murde4Ufd38x1vx7uT0wshBj3TY+hyj7IlmcsjK1eEmjgdafYK8kwHXxYn0
box74d4GPj9bomlZmJbYClNyGey4P/SEgHKtfIfQOfW+Q/wappiui8ePwDQIho9YYmnc+X37q7Ud
OA//pXXqb+uA9y7DcfVX/NGa5gP6yw2GC0f1MLn01k639+mNIE633CBOZn+qWTd19+MnmIRdk8gB
zMjspY2i0WuYlM0LsBz0bKb1o7s10Taei/gcYBW6spLA8+fecHbnCpt+dUDuF7nLo5a1HnWR7u2I
WltCye8QETi2nOVNK+0Cvpwzkp+0DW5IpopKwSTolwiCcc6zIMMsE07IoG8XWntM3FqE2w/tLoTQ
BBbp0lE0aQuY0QtaGwdgZYMTIJPOqklhXoOTd/fjJCq4w6+wIS9x+D28YfrcsistAcxp6tHY3wst
OEYve1kt5E5phIrarPnND1xGhr3XPmmixawg797jXmvYEmATw6vBSE3BGDV7phbjsqIJXPGspx6+
or6Ki2ixr9aMe1N/9K2IE37qVVh984JPT5i1OL+XzvkGsECyT4Hv1Gfoaqnfd9ok0afbUhKen5x+
bSJYWynmoB0f9OnVvu8GXjlqHl1k78dqjuc5ltIEpX1PwwVABKDZM0f2qZT6SG1x9s++l1kKTYLp
HV6yzbT1AUmYJiE/tubR78EbC8ZpWKoQZSnBKXyrEIk9FGabHUtWNK4rpU3C9v7dsMP3wHLoaubt
qgutyEht2cxxDXzsu3RTpiC7xRJNQs3H8xPTRWtEdmPgt8+bGth1yaC43SFf6cePqYPZZLHLzkJ+
vz5yx+Rq2IRwRxtiY/gscqM7KbOp2q+Fm7uQQPco3E1N95I3wmXagOOy3aSRD2wiw42YBL+Mkgsa
TV7LJi4IIvjx8J6xUWI8sxeBAJM+HUZ4AOc6T44Pr0ZHO1ziil4J3jx8zCfsoJJLoSVkJRUcWOCx
gFq33XFnKY1XalMEVPrP1Xceu6JsDXfUmMTcoei7KY+Iz6RnuKZ8SV7vJTb4qra/qSuC6HMP4vqA
C7P+Q7mH0i+YzaU/AYi4jepRh+L7qwaz+Jsd/IMCK5m/BTDARmqQD55WIX6S8xk98KPhZcwvWF4i
4+mTpHBjIBC4ibSehWnBbbIYgJNQKWkHU44qwMp4clg2Xg2yIFC3rhTRhZ7uVVY+9kLFo1VHXw2O
6FPaJ+9qKSq9zSRo5Q+231oFiYtniq3PtSrGbF2bpBmHLMy2LLR4lPuIxVKxTCS/cKMjAPWM4uYW
0TGVGBiABT6/0TF30+2ZEf57P+loWBkba9+AJ9WqywU/RcjL/T+hRzmtTb3nqZGiya9+DiIVxB5p
iofVfe87zOkPZ8b4VQVp39qeIfK4CCB3ASsIIVKrezhL1+mAIzXwM7HyPYLH0f1NpPO8bThwZUxJ
ltNw1su+NncPVfb+ep0QPhtrO3p5E9dPlJisTHTEAmokRjHiZEkZrissqzh7Yzf0wesqB3aFMUwy
OoH9uYyFFiUO1Fv/4/LcBXw2/1oyJi/3sGJbslJpracp2G+3zW+8LzgqdL3AxRNDdVUTYclkSwd6
HjdvmPJjUvPbSPwtWUdE/cOOI1jsFwnOYKleoPJmAQnaZzJ1B9MlKvAAEkD2SKdPxcWcktdm75Gy
TM3pEgeMh40SZcrjH4FNca62bTj1JQoqSkBps5MY/Vh6Z949l8QkEbH03ehFh4uYjAr8KtiTE5Ei
JrTKGSRIcMgXL5wO3xel8sbTFcM5aaJ2+RGI5cg8VZ72Trc61IkmZZtgRmpFfH/HjBregZ3Zycpz
pFoJozhKBc2dYYJxX2eipPpgluXekVVnQ+mHnNuarGiSkesuA1+s62mrSOYLJgTuF9APXKjrntqW
B8LYne7aEtlvyvTuk+pCy44YQhf6bYZgGRPYYGy4FMHFERy1+jGQ76TwMRRaUW8EOzqjesVJQv99
wvto3ut7kbFHYpdCp/Wf0z5NEiLTvoPmeWuYMaRQUx110MRL2ludJzhCLjW/eW40sKJ26MH9F4Jq
u9WRkrYKQxv6Lltam6oRPOVjz3RXq6oSw2s/z7FEc5fsJqlZk7wz5dDK9IkaUwsrkUARez0OwMD2
FWWTXgYsnFEhCreRTS23bXWrXdtMXaWKT/Q0zG9DqYwQYa1excfcWHVcvYm1e0AwoHQ4eDZZNuFU
8HbrH5r5ivQSr1/E69hPXKGOeqL/+Ei/eLzPqA3ocBmgfncstOT8WXZ90/8YBfRFGxblwvPP2AvR
gz7MWwfNlSoo1a/BFs2gdqcUabLETq8SpK4L+BiY/HDhheaGjtjclphfgWecnwoIzAPIm4pcFje5
TAU7nELo8mwljHRypUxjUNCMS2VdGNiQHtFFlsGcR5R+arBhD0SOy6PSLU+nfg99cIePmGRdv5ka
H4nhRvVRa+RMt4D0wqef/tNxx8i+1PcSyjIzxjWw8EewudbjHO+oegKVGTl4boFJNojN0MWYy9Po
dONYqVeA6pmKsbg0gtf9wGo+AcibbBF5I7XcQ77yq7/C5NBUrhQ526QL6nt5eEZu1tDIRdhVbLpX
4DGLC7n0E+/xgedGXMED44DIYxuoLf6c03pDvSaI51x7wgpq5ApQj2/Nek2NnFbWoli705v8qUqJ
fLbZpLQ8oKHfoO139UBMMT8RX1Y4xaTRrmW9nBizpdgaBWcT10i4y/pp3IjC9c/HoihKWVVZcE0C
iN2/e94jy2Qw+z7R4PDa0HsruALvYd5QEOpK0+MgRYQ2GYgaM/59mefRH4ZohiJI0zoZ8IFPLdCM
p2gd51zg/HAnJVwzGmP77lQAssT9kJO2yNpEty29uLKnEW3acuMVCo3YREW50rzZRNK+fahi7Ql2
TQYUggzbaRBMVCS/i9vTrUU5aLKI7mWKdTbV6dzLMPQLwwwKh1vEv8dTAb5PQK52ib8aPxA43fNt
Y3ta0tiwlARylyobk7KS4fN2aGTI9bYJdiMu/zHIGNI16Q0B6+aIsKMiUDae6nJKUaQipuBrwqZ3
AFV90LP/fbVl+1KLp2SeWQ+NgPnBV5CtKJt9kD/hlVOmevL80S9Fk7jXrWY8J8UT7LpnTcmfrp5f
Ja+cgyWasbhAKv2lXHuUBblKsmg5UJjwgluX4m1lEG3Y6eODfs+E2LjDh9ddaUZu2T/ifuo/XpTN
+XX1DlLqQrfpiJw4c0+YjRPUx9Rj0ls5bbTH1xRylvAZbRZnlU9sVtPUQyys9oqu9wZhTegijsJy
eeLVsgT3w49//WoKsyoRPvuVqDjHx1HxmCgr3e1OXm7Hz/9LhJJ9Atkw3K7kt0foElxdmXYUEmwN
j4eqxgi+XatB6vV+2WJ7XDUr0+pacwQdIUXrC+OiDCn0IxF34GKWs4tmc6ZnJ8nVEQDXR2QWWQqJ
U8GvRbDPEzni+a9mlcVO8C9mKUuG+OyM6GyHr3W7B40exn8rFbfJ1HR7m9sdy5c5CulzXdeHfWgd
SKp1Nd81jL78Ocd54sZ3GwsH/v8NtdhxI4XOHogzYqpdKK43XoP545XMmXw3EpGJQeRnUvtRHgsc
ZKsyMlyOW2nbXDmIIMZg2Nbr6D4efba1/yUZet5YKQ7cRBwMbayb2kqW5oNHXZUAgOGzziHpMuzE
dEmPfP9wx/g9R987cnZo220Fvi4kIHt8lW4ncTZqXkfcnKqvmG3v8auIiwRKPDmQogP7mw6Kg7bf
2FsoQHYAp8tLBu38Az/ojGCOGdwFED+j3W7n8WCiwjLWzRhRmj26W/9ma3YFyvFEpfDCFugD9T0V
TVaLg7i8cbAdkPdxiD4X9tRpV2nY+x5oiZW+SwvJyvx6X18IFzyf6m+08bpv2Lpr0B/kEQcIM7fD
sQFx6BU1b1f9mLb/TXF1+b5yPvgP5lnn1EK8zcf0T/uN4nEhipY/Egn8SAMHpdpPV+WxtbxU6VSZ
B3O2gEt/qvWeCBhUF1sp4XNSmTYDxyN9XApXx0iaDNddAQRyOcwMcPhngryOWxlCpRna4mmDOA14
ujwouIfOCKHPBCJrEbdcTHJTM+FPSeB+7Bip6hTk9zwMGTSv6cubIkG2w8rFeZn+FgK+O9ZGiBLY
sGUMRfdNOrahfWFBn6572FpsgcyXHHhppHlIXkICupvy53DlWV8O+rIPY/orTuXrSTb/heo9Z1td
90OnVCbnQ64cdXSZgmJL+jWKjUeE+6kHPfUEd1w0ZwLXYeQOEasarY+Dvbz8AUDrCepiFO5y+zxE
0f5WyAgHRGtlOimL0AgRkvdz0bIqOVl/dhVwLotUOQoPOGwe6mLMaiTFjfaS4fy+xucsaInHyKPs
DzyvyGbnaCBchCRmyJsAlKd38OSjPG+JQNC7GGTTnFRrYmzqDZfZwXJjOJnzJG/t1m1Wf4i+kt3K
sO/LmAcibf3aIG7yqdcLRXl39t5E7mMNzYg9H7qy7yH97XAJx8wOE9kdwLyqvr8SNzo4jDy6twj+
HDKE1Cfuft7X6JL8djtdAW8qH5YBcwhi3aZJtAbpUK6LHLYVZrePYs2UkxPe74AH0YYzHo2n/jLZ
2AOZCkiEUsMHl6cOI8f2W+0FbUBruWDLbQeoK4GyV1iMLgagYkdhuBGU/DxAxEvlr38ySjiav9oh
p9SSy4gOyyYlK5TcfkU1PJvKozY9c9zjGGUggs4wV13UMDDgyAh6zGjX4Nj40at3IPlkHSWGrJma
dJ4S42U75cDkGRSzMAu48DvGQM7/R7FSCaIJ9+Dw3mNeml5eft0RCUTFdEucfabrq6BqMrqFRfBh
rp2e74MWvbk9jEjiLV/KF8PXo5HVPWYRH4u7b9uRATYmW/pRaPZh4BcrEd0SfQhmaKiei9KC2n0c
O3BBJ+gm/chE54w6Dno6wYcKaR1LeyLfRaQSnDpKqS2NPi4QoD9c6xHPGEjeBGGvwJ87nEXE1w6v
w6Hc3Ig0mmktt8wQPjVXWGPy/wtKeYxVlNVy8op+UgYJzRwCEDtp63TxHR+Fxz3Vi43dojCqpp8R
dnY0tU9qZ9W7sF6gZ1oZkdS8WFiG0wpaXgyiR65IH0uvIyAkXzYnj4IZhFvnTBli5dYk+jHVf/+o
5tBHTLkhb83JPO+usLhJSyFF48nbl6soOfKyA0T0PJUKHeEwaaL5O0B0b/XXi8NxfceD+PJ0kIbz
LrvYGh7uNj8bt8mOF7PxYoqCRZgvsbefnFj/aN8s5zHaIliCNxOQK82axq1fKV2/TNWzHFbSt96+
6tc2qjEoN4/mJjr75KRDE3KBQcLcPoLwcOhdKsrgGhINhAlM0GUOVT1rELyDNX6j9d4bWw6Z2Dg1
t4buv2dZ24WRJBQbvNpNtF9wvS8nPoIzbTsBCZkk8NzhRtSPnC8DF2MFZXltSeel//dcksPEmATD
r+c3eYTXf9YjuK0JwlxHwoHGMBdUBCCFhfOWxrpQg3DRIoKkWPrhz/0B14JPzbA6XCcvedBk7QHo
l/XVhAzg3QhhQdGi69uRH1Jx4DbUHEMKaropqGWdu2+Q1KKPvC43t/ZfMj7ERYjgUNTNEo34p9Lz
B+/PbAaZtDTVFAKn64L/oGQrTh8R9ppwlZ4heL4gqHZGn+9CGoN2H6gPykUatNEtvX0z5YVTUWQ+
L5uNfa4ZvF2vvDDtYodHDlLuQkNSP4pm5vEy8D03/6HIhxIloVlZwT90ImiU4zIzribMwmcc6fKM
Tv2GUWTc+0q/Pz5BXhbkedYO5cKxzSZPuRCZn0GXZVIRyuM+b/65sRBpaAQhUcy3IOBTq3WuZkTo
0KFR25NKUfJmkfGr5KgNpjyZOE1vezBOihpW6DzSrKjH9aKuV6pLyuMdKg8+wXGhQg2uQFDnEtaz
td+8xhPKGr6AE0d2hYjlBtquuJd/A5XMCzhWQjAusC5txbqZoVTXUBeMeX8p3m5yCW+awX/6L7Qm
hxZn2DDWKtacu9gDAdM0NcI7Pb73DSR6RrPFM4OR9d5h7mgaYowlT+rphcAnaKSSS4vziKBzW6+B
uWt9v2zM8aVuDK5oOpudJFfFqF9UqqgEHY78QIWMW/OWhT+DIhUCOtWHA1/9fbD4f4wuDe1KJb7b
d68f0kGPwceaV+D3jJ2eOrsH6gBhCuK0C1yUCS9pvFg07LqnwHWZM3b+oofxZ1Z3g/nI71/Ah5mq
ftTa9gySEujpT3tEc0kLHTOp1vhc02Xr30oMB6ZJBly1LsavPyGTSSi4TB6zgXz0eHALF9iklO+p
mGpkdxfp7PvtXdKyjVeajDLG8QdJ4yGJ3dA9/AbCe+vcWtIV1e9Ccl+sPzpnJ+ZLHRd3QqPM/hYI
1CAB3tKg51EejfRWh5bkgUIJ8EoAvqQiblSUiyo93lyfz02s88B7vAF2L0F7xsnc/Ho/KXF+TSpm
QJdLgCzoK/pl70KH9V6migP5J7vMITNtYtHacNHI9AFmMjFt2KwevrF6BrDQRcL8nYnCossnwSYN
QcJMZd7X4eJnYSAMfcxEdr66K1cqV1okJzQjQ0R9AnfPGTeLABV0qmkvUArNfRSbMLKw+v3+eokp
jLBYwMuOuIUkWWCjmd7IkHZfjeqb8WJ576pe+R24MuX11Eg+gkGtMM+ra80R6oaHzWFLRhF/06on
fvQgAAdMbaFpNqQBtsOZefzrIh/XEhyeRE2TNIaptFqpmRaH2/mw3hle2oD0QZEWpfoqK9ONqXhQ
02/ggSt0a4DNP8aoAhjkWIrflbCWVfwnWT1Cw7mzrIH9On7GbcFByLy7kRBfQXzBEUfmBEkvrcAw
aCrWznHYVdGFyhYBtrQ/0rT9N28KRW7Dnx/AR9+e+CMMwQ8A7mwQJaxf4T8YM5tdigyJ1S+qBnXr
9nY3X0rlMVEiMi5WjzYY4qStcJ86pzqcIFvzmE1JoQ86W4uURFSmJyxn1FFPBL19dTjB8o1RKKv4
aYf+tvXVfT8fGMeXGC7wOZef8QXxfF1cnQ6eBKNzFb9UoyVlKmGocWaD045VybBK+6X79zy4jr2y
bCZDB4T1AEadvDr9r4eNpe8DQD+0kpfwJTOvEMYO9CgZDsXZs6p+7EM0ebFU6Il2popumXUnAs4G
2BBu1F6dcGcRM3ZWGl8kTpzWEGkC0H849d9W1rLyB0j5a778MaxiW2+LBKixeSVpWY43yygxSwj7
gA2kYBKcR718aKQEQhiUU/n1NrssFSqZHBs1Q4Yqj1y4VDEvXJDlFNJOu2ww72RVDPui0ha3xM+6
xhmF+lmVf7Kukk5Cp0K0Jb0foJDPPCYl9+9NHgutjIIZ56DD8ppO8kWiumErjK9GnMbmLy6PNSlI
R5QT2Zoz97SBqQmUkRx4iX7vnLUD+lCdbaT9jkKS4B3XTKj9FKYj99HdEAHVO+xojrOnJ9cyTih1
awL8M0MVL6N34SQOHh/zMWJkxwDztwukY63D8yxAzjo1yD1dwJ6TwsMoIwDvYjAaPxRUyPEu8yRC
MVh6mXb/l+BAL9xvSA0d+YNp/6emtzne1lVTx/Xs9X9sMzSKOw6zEA/8WSSiFEikkq2cZHkLKFYw
V4RKzGiddJjX6xi0yYpTDQ4oWw1x6CIDBogwQM9v0jKatKLj4ce1L/RQOWhaCDYZzmdcnLXa6CmE
RlfaQ8If0iQfqzOM+QxZ00B0uuJ2pSR2rNUFymSocoEXeL9bNw+acNVofTaYNX2WsJUj1Qu61SUd
xMoVXdVsgdvb6kxa2nPSiUhQ9kYiwhfmRcFuvV/ax/j82kFYHkeMudZFyanjtZRO9mutPQ36rHUK
BzCta8mPWDqLRjID4U8Vo9Bx6QnbdV5JLBsPJRiobD3plB5I2JDve2Esn4CGRYgHTmaB9UPU39rg
tICWh56Vw+LRuZsNv9cxWCtqn2p3lO9qH/o3GD+ygPAg+e5zG6HqSjwXHptPH6Aer7C6Eo2SU94q
KlI7yP/4lW5Mqs1Krw8i4WiBw4eULQxuOg4+VI2z7Jr0/82ikdvF0nEheUeveDswltRdCLcpL43i
92UhijOCz9G6ME8BjCi/Cz/3HXJxFlkBEf7Epa50K/f5KurTvR4DmJN6a7HGCT2mqK8WwbfdBxO6
wvGdGnqhd5XmO+c4v+vIXudYy2CRxX3jcgT/prE0aM9quE1yFipjitg2nCBNAfx3M3p9Z2WHYOjY
upXtYUrT6rvmOxpkF+wAljZlWXjzTM9orMTjO2O7dgVCn4M4l1gj0gk36Mplq3jSe3/Oes7qPyVP
Q5Sv9SdZG5VsU/GJPYU95IQjY+HPQwhmkbjt+v4o8TB4A0ZDt8LbzjXcZYPTSeU3trXJCSn/AkkA
g9sihjXqBnIIf6z9CX2cbM8hpVMhSYfhD1CRbMj+C5QJPNLIatcZgY7COZa/9YJqYByo6r9tb6qO
KI8e/CwHptV5PiAY5RmFaCPKq9uBhn4n68alm4gy/J+VDwIB0aTcjCkIJ0BOnFDYjKGhQwav98LY
UjlW4fhfVAYswzNJW0HDJy1b052eybP+7lIhTW/Kb3owofyJ2PaMt6Q+akdKFL2sMlOB0YbZ5ap8
pUEPAcEZFk7hjA98mEmewMQtHNPbzUylmvSakV3zX+Q63raCSvgrmI4SPqgMXO2xXbSnRZP1YVbU
K89j57h2iLySE93qHCNxuma9qZSCHPW1/JNt/7fbhUF5KGjOkYADkbAZ6OTSGECjtCgSZgBJBBB/
IFFfYLymvwHA1kus9LAGP1kNb7ttfQMn5iCYFIDYUU+Zrg65ablNdmjcMw3LW3kFJdom3vXHL+An
HMmBbrfDMSwUjHrgNPYwFSntob5/W3jU4agO8MkuyUo7ry6KcyaZZbtp7acyxSkKPq+jlHGr+Dns
vntpI0u3ePkyn/iydVHwsW2tLlwfubPJtqu2TKvDZ/bhZrHHGJeznvMd3mvlEWYRcgVL9VM5vj6m
7Qmr5gxxhMlb6hrdV7SgvxZlG3N6RLxewIQM+bahemDl0Fc0eQ9ICyfFOFnPT5aKW2uIGbiJffFn
hlnvSPFUK7O23IeAB1k9mPbd7f/fCRxzq8t6lrIO0Ovts61alQIWdaPxhB6YMdQsdRHxgR+JH3Q2
UHQh8Ub3aW1z1WMPvGAUIWzeE2ZTI/vx4Pkbtgn4ftkiEczTTsFBqfgdEjLjKCJh1Y2S+rdM85O9
SiBlLscRKOOJLtjkAbHDZGf2e6x/UwKLyAyCRQmrMdamFRsz8k8zuqtiezZRMMYWXPN7LLB3kBCf
cRJw1wo+OIz4CQ20731OEx2WuXuU9yS7seQAYOSYtF9hwcNoqPfUQyVsjrkPCMEZYYlB5k/ctnkx
D2y/Dd818FkVVJyDZOZlbXnKUO/ZlBNMcBdQEMoCcb/YDmWZ3+bOjA0HEsLVgHtrWlZrxKam1aq8
+L2sWZR1oz1t/7+dw1wtWaeKyUUA6rIHI8F4CVJW09gKjWe27ZJt5gap0QvPk2esLXa1FM6JDE2v
fkgYE/zcqPOOh159Vznt60dlrUV/4YOI8VMxvTgjITCNTE3kF/PgYSXQQDU0mJoQXfarTceDK6yC
7C/aWCim+4pMfpy1yxELGfzhYzicox4cVQABm1MIc36jsArGI7gHBOUQ2pbyEn9yCsxegg0PvH//
z0boqeR+lPJpC7VZ+gg6lBvNkLbOvOk2t8NqzSnBaWjPsVg96hAG/8BFHcZv7tUg83oCgBSZiWVX
wzZ83AG8KM50mDY3mbTwxmaAhYt3Sy0AzlV00HvWuipmfGVH7SH27hBgCfl4T2eUaI4xH7Co6oDh
T88KDzz/0m/N5/s39cENvRzmy8vkbw71hnnCAA/Vpdzzbag85JVIVv67Z74I4BzTDYQ52XbEQTZk
fS4rY05u7nSgX9lvlwIQK/bqjt7OkvwRfFU+ypLQJCc50Tm/8iPiXaBAwArb5IsNLyc8GDiNaIar
KSwl198ny2kWd8W3yk5rIkQVPGb4WDUO06CZV2bzwiHFbiPVSb7opQCZD38zkOA7c/S0fTMptcLY
RVTqG+ngcsrZSRb1sZmqZfv/HRxcTf7oc7ezehzqOPQH+YXbyFT59OwEi7shgSXdZlVK3YjlAXOh
00i/EgSfJaOT2iaipw1VWOvr1oBiVFa3MVWoeH90DZcW7CgpleaqG7Cu0VMhxgq5HZ+BejgDokIB
gktFWQpCWISMCIFEbmQnOwTL28vqGoR6qxu8ibeKZ8RpoPg3WV8YaE+fHpuPDYc/K/m6tsaron2V
Giu4pjU8eKCHRNGn+skL3oRKnUNAW3e2cI6o7y5h08rcvewiBgzg3thsoDM7jKuWJL/1eD+WI0WS
XUwDDoe5cHbQQq2DoOBtbt4Cr9146rpKPJKuuUa/2uuMbuizB02LpmTcnbrqARXy/PxccXv+9gEQ
PtsmKMVXcZkfnErh80elqwOu2lr3I5d/iUpmmAKPoKEYf3irMV39B96LONepJudDk2MJp6SEbfXL
c7YY5XjckfSOf88PzSHDuGgXkSSGF1YAlKtkJlpq/RArzlUHEd2nXNUgt3So6vwfL+nuYS9f2JoU
sp1Kz5ZR4mkk3G25x1+HHE0DpgXbmKVEhY03hLoVc0hmpXoi680u+MSk+o6LUWi4RuXEeKqCKULj
cQy/xDn4iLFCaYbu7aLJMvt3gUk3JrQ71aY/UlcjbXVVMh5HoTEohfBuLGESE6PO8IjE8pyEKqmO
7VmC0S813RKhAUJfa8s8hHvy8lbjwaIik+MQJ8l8wFQm5+Ll8TCFr47vW2CIzL7l5bFKkDPrY7Ed
yj3GaqNmHDmxzp+PKLilValrQIJmtACVBCMEXiTWbQ0Tspjpy0VUvkMi+sr7F8sT11/Q2HtzTmo1
WmhKy0C9QinLKUVvdlSQ2hvWDDdL9YXLHw/u46nn+Ie/Fh6CFfNA3F+TP+IIkQGHRsGJ3QGAjBdh
BUZvOq23hLebDC84tRzG2mXE+99CiTWPdHo88BHA3rTC5Kq3ye0fusutqQffDgvUpPoUsdOhruj+
qU2jBN7FueJuYiAexz03ebvBu7E/7ZXO1lQAiICmOL9c59RsIvstJiF4xGfcCDKn4OWqeE7M3Hf4
877ZdCEuWrsipyj8sLOxTqT2vdigY1HFhDhIK8ji2NZpd94o+KxPSpuuRvf2Lfc/LNP+TwwYC+b+
FpiW6y0LHZw56MVbSYbjUNMGGzzB75DE3lb6zWPzrcze9oJjAFKhL/kXyNeoRF3q22I9RA0QeG4A
1x5xsKsKopF/ZgMz3q6d0BkIaExePfBAba4pXNhk6FWxF9MkegcVwI5/1y7uj3X0vh+6FTL2RtYb
WCxzc1D7ODRLDP06scwbUTJNu7EXQj2FqxxRDPixzOegYrRoKSjDylwtW8cMB0Tam07goIopXIzH
yVgNCvql9faYxRf7NQSXoXmEKq3EWN/gSBLnG9w+WwnrWhjHbLcporJPEdDuNeM1tLJeCNC1afdZ
8jaa88wrLTbxhdEwXlSEkb3qinVuVqjslTunEj73O3wlb8S4tR6vm4a2qg7dLzrE6B/Erpz4IWpg
yapeqmtmGiGor3lPVIR4HsG+Ipd/mYhL80cdGlrz6Npp6oYu7TN3+uwE5FBAAVq/RgF8lVicI/5E
ptKQ8YEaIyuO1zGUrwpF0vAxK9e7r2gMvZYgNhm3UaqvnxxvzsmZg/pa4C+xmELwJUN8j4bZb2fS
0znjguikPXq0OM/TzDIW+gajc9x2tydZEJE5kA4vJh5FoqvP32pSV26PiyDEwnF/atAXEPnE8ycN
9moEKUc0zBfTTDpIp6Vq1v6Uozs1SqE1JTWif1NiSkpEgs7avmkZ0iKrIF2EfUCh0L67SvSCkFQm
9xtcmc/UHKtmloW+B2MU2Yw30GwypyUC5DpOYULZlNnSN6Kta5ZN2eZHdNQgiSagmeiJuyIOD+d7
5vj8MAhKjwIP5czovZnTVZfLv6TPPZizv7HjI+xa6y7Q8fVhrvH50lm332cjZ9AeY+F0LnAO1CU3
UGIDRUJ8/Dmnfjg/td04a/4RTLveAqAzCEghSq54SriAh2Qb1SZjOF0wuXp8ENnzd8RUmCstGgra
m7dKSO0N71ByADJOIDDIZAUt/0+p8AZt+fIv9R1gc+mtB+2GwgeGXhOMQm0hd4LW0MR5qKoyK+yy
r+Snfkl0GVynX/gSlaFUE+2bCeqSsJu3Yz3wJqzO9Ct6o1Q/pD9SBEl20SjbrGoFg7Qtza4KBqdJ
LyrhzTlVoz+Wl5mOJgBK0glbBFSH/Hm462VTy0PE0FzNKoZ/fpBe/w0OdvAxzNfvjEtvTMlt8209
GvfH+26DUlkCigr63p+yoA8elHqHHE+dtX3xvV5QijSs9Ivo/Ss8/zwEZDwqRpG0Tiw1u7DtsnPC
6aiNhXBt9jl3vdYkVEXvRe3khat7a9zyZsPAGuUlXNtBW/tGgOcdPTspaQt82NciDDeaIoldcVo7
JJjSumZp6Pp4jzMRE8yGXeTMCeMg5xvgiUbtgJPbaALA/JQk8cDHSjkr+QsQjfugHkk5Z8RYpHTb
OprsPSrTiIBavTpK35sZBCjwcR3801WPKeBJbyLxHmPvVUQn5kSFEKCML2LSi7Ifjm1s5EtrK5Yc
bETd42wSc0f4svW7JSz7kfQpSjfAZ/iy/CsPfH9R4Kosyc1IgNeWLuK/P3RmgaQ8V/Npk5vOkHxW
4+E0+/GU9NmDmBQbgex/KVV94F+WhepQ5Ij7OCbdAu+FT+QD4FPX3ic0EgzDo80LPWwnnbQkYCzf
oWeKbkwWOghUZ2NTNDX1ST/HZnMMflCTilrQ9BarAJMSNunGbWCEVJ5RqEC79kmSLXTG+xej0GMw
nQ+BYy8AqKIOVDQC8bqktfVTWQXriYgocKWK+zHkeaf2ZuDqWEaKtvMGtgYUe9z1jL1JitlXT3hr
3im6eNubrGkFlm+TGqjZ7oS8Z6pUbR04qM4TbLTgd4nuHwTYigPa1haEaPhmNWsScpMMnDBCgoIj
Inj4081Y+Vq1mr9QyBrE0ZmfM5tbPkW+EGOdMry+dmaw/8zAJP8jffzr0RBIzzI8cEn0ArIlaXjJ
Oo7dgIM7ESI4FVEMk/cmS3iRiVgoLe74g0NKl7EYDbJsZDwZNWnSdOtREQFEhI9vWks9NBF7Veaf
wFbPIX8XKN1Cn40UJCE16WjbSmepDXWIPa4+FXAlLF3uhfUwg8FIqB4tucCAaB1ITWzbFEdWVSnB
URhtAKA3mwrzYBChhpeXu2Xm40Qlm62Oqhb0CPWPnHC2xnu8bmmEfIjj8r8icRbahoHF8Tx32E6S
7xwQMLyjwtiwws6G2bX8QoBct9oSwkryD9w3NA/0dw8Ay2hL6jdywsJS94UIrLOxMacA0xi/tAar
JcLZejfKRDptKjzrI2pd4huvzbdYIyj05Sdbk1+OrBeZROwSr2EHcyWTO+V8pDlmHmw4+OI0nUUk
0ze+nu+eK0GgdlyQiiwNhajWlq/o4rDI+h4JWENzprM13/1d6HudO+R5RDjDOIXK4ORK1GiyxLkH
2QrszvMdkaDr27BYCjEhkIrsPxDNanzRQv5sOhKgFrAVcokBsvm1mOYjB0R/wFag+xmNgYxT4kGT
aFYA5dbO3khsmV4939B04ZJ5eof7UuUi/sDQlcL3zJLMoaUQADHSj90gQaXxs2oRcvCBUk9q2eIa
8fNSvW878tKVKHwZhVm7fe9Hoaa37kTYuyOTXpnA+pLRjYHlfQxP2M8dZloG1fU5J//KAGKYfukO
tp4GRdMG5TU2RhhYO2o8sdwBAoz+PA46pstf5X/R7fSjcPOaQI93hI0aliIMeY+zfus2eZetvYJT
k2qTeXVNxNTWS0DtXWi6FcfbDwz/yLJUm39CTy/bORE+yOEG/PXAsEoQ4SitPL8bMKkJ+xQvGjTF
ot6D9KzkNBPR15D89XXYPNey64ecjNSTrZolF+4t1VqjUULJZI4PtfTFQdPTqZAIbJ7D5bWlp3F6
UsK/Hj+uAasDE6FxgbDPChWZ1Bv4pH+M3HvfM+IgtgfPOIGeE+DaP19z7Gl/SdDwvOSEL33J3Pn0
wfv5LvBI5E4Nmc7rcS5TXEyxL3Z6ZgudKO2bIMTEzwBr1B2G6Q6cZcy7/Y3KGhn6orUC+0Iv8SS7
iAtRukQ+SdxwjuYsXNXvQa2uDYIKm3IuZDZea5XjyiGcSxDTXum8izBknJAOeN4H+Ye/jJ3DzPs1
nfmMym77wuy3Vd0BOHaC2FZ2fOP8nOe69+gQXgFAo47cOL0mPk6pu1ytSVPRqpfQ0rqBxEtXRke9
/z1bfjEuDVu6o7c54NhgtNK7T05pVB07iJ14IxXLNEcSeoa6G2k45Q1pqDla8pLOgS7MwhagEtrP
ccu/AmS1/9H36pfXswQW7xAWzL0r5r9EyB37gSRbMCHfIwjN1Rx8cHsLXAfahynlhuwz2Fz4LDlX
676WSg4T4b+EtKcOK3+istwRNNRQsgtMOhbHgIyk4nHEXPOywQOu9IiUq/vHpkDO4r+DkG7wSDna
CXZMwtf2HE8TwNkHwOq/Y/AmmuL9AR0Vk8OzER9WOjj1Hh+gR4OsB3kVBOo/2Usy4GMAFVGasDTk
tx+NmasM2kQ0IqtawKpB3EdwcnA9Qexw3n4l613s1V86qgwtx0zKJKeYTdTg49qqiLrHQ+GeP6jO
gNiCVGRANeR9qHGw6mApuKDMNW8IaQCZoJdocNMWwLI/wHFIahwqwtspYtejH3XuWcdXo2EnTXC0
6LVU95cCvKoYAzNdNHzv4nM9RFwWVXyvIEZrJ0pe9HWj11BFlBZnrQ4ffjATFQ85OSO2+/Me2q3w
bTWLfPyWNkIj5jfcvlRv6yHBNNFKWw+k2aBi+P+7UQExry4bns9XwMsVbReIJbWqPz/kUpfN158i
8B/V/kpV14vI45PAKFMw56+Bbdxyn0dDxXE9QpkW0XtTycE9Gj8sS0LtsPAAblLuK5OM/KBpYe4s
jeJMekz2KmpL1Qj8tzdDmsTwvhZqhNnVolp9po9xipho33dW9jL5bnKBLgmv+KpxmPp5+Le+iyNW
NtFPq5ExhyE0wzR2hBe6zjLg7gPQUVA+xJ+QO9Hp7yeuHJJZiprB5j3vm//Po2zzAEcHI0vzP6GN
ik19mlll9xxmhWLvFFf7zuaiGWVswU995tt0OppdhFtM4XBTw9ux+InvFw6JHfbuxgXcdZIhVPIH
myF+T91qGkLd8Vgrs8iWmNVp+032W6jxJMDStPzm1/0mvghfazbD/yMfU16qHldfG4jSXjLudfkg
mPFC69ZgqF/DJuhvm12hk4XmysYbb/HE/uNqKQyho6esXZCbPjxOIprfXuPHKziK57fjmfYZRBZg
k4h12rUbrwVeJBY2pEAjS+/fck8l3X4veMqqsD9H0y5+2QSMCZSqIFHq7QMKIEOvraI89pmu5SSZ
ctqJN9I+CICxzCkLh9s6v2PlNtLfWBrzfaaEGG9Gc52d7n1iTBJyBSNRAzSWuMQ6rgFodwkNl9ms
tkPNTbg/SUDP65b8i8B6QU2cJbkTecqck6x55wJ0zQSL9soLNVBoSwN6mXgeXG6NPmQXLy5tmbAn
0T5d2zSClt/b/fAMJeXuOQwONOFeY7AgHhu7dGjtmvfgHzFUlmaZ2YzZGvNb2UjFWK8tvN1Y9zFc
HGVjFw/7pPT0JejuMZ3zx/PGkviAYTYrmj0Rjlk0CFvklFHudu2Uym6f+3pPFunQKTtjZm7nlLIw
HKbRvBvCNdYPVbcFrhiqcFPydHvRR7Pb/Jkz4C6HTRCYr/AlJSzh15ZYI1cdlsZGrC44iyAWi14U
mnaA/G85XH3/u0/51x3pla0hVDNZywLBChLQPS06ccG7lHCycsjhw+y1oyANvo3edxyTE9ZSTkjL
2zANdb0eK9ajFMzR5gf4s3hAcp9PBh6/b4Ys7F4BZr5KPiK6vmFIAOKMiE3F3OvNF5yPIMVSLR6d
KP2szMPpQLQRwZM9L2i650Z6wOF+huiBNnMDyLd8H+4abrNDvp8K4CjgCsj8uHfwhfvYSxFA0KfB
neiYpOlM24/wxZXarJ62ggc69acz0y6HbUA3oD82hiF+w/NtDN/bPOL7e9LsF27Xd7rMjUcz0M6g
qhW9EeH52SbTArbe+QIVA06mdG6lCWAMJ968aSUn+k7KNz8efJMk8iL7cp86dIuOnhyAki1qiB9D
qXr4Apyn+14wzhKIFj9rO1wJyA7JG+htaIKJCuWr+aPEiZhC6Opw93icu0n6gc1YCxG9SN+IEW+b
YyOfN41mWsulITBPfEio9QSxuBtHe7Yf30Oj21CGPvgvX9SJMsf7dk7xtSPlNPfaCUO+WSEaVClm
jiYudmS7t2MHfh9uoUEJ0d7WizrS7RDKjyQyE1fxiOIAEMDiTNhqR2tOY14qlm9TNddpZ4Qijt+j
02WcsPXNlTZj7Xl8oiwYfVmdrW1+Ngjwl+Wh4K0WlCY+ZaNhj8y260OAYHcv4SDwFsKgLJqPMkRy
ROVdgLsxsDTtCUT7vje58ygCCe5zWmGBM6E3bnHwOUH564VXf2RbTs7X6M+fuzgF9ZEnHlFVl8Aq
qcCMYDYtGt1xyCixWO8KUzymPj9y4jZmgTa7IG3lTbJm0DPp786DikgnKZnlKnVrzeZZMc37+mpj
+o8ahCKU1GzMuI8OujuWKR6Cgwd1RLrHS+LOptdyE2NpZDYSKby13iBXkSMNgyp9t8eVY5JP5YsV
V6ezteeErBqiQa7mXV1mWBDQtizLtYJ6kHKT/5oNp9Mnk1HUPt0TQWsNeX0FiiWexezuANMG8x6a
AqlZJ41wTa4NszHsI/6xOnqv4kBqlvYwKr8ori3HLZ/v7jnmGFZgmzdQe71PQgEOfh+1zkGFwvUT
/q9IYA2LiWlhjKrFWZH/xk4V+4TZ5WsxotlRGIGZ4cDQLeLulOWu5wuV8D/jD/YpQCl1314CcegP
Sjg/OTUfm0gSx+V3b50m72161OTwG5p0s4/8mS257u0LUfANZ4ZksUmnYZppGbqGHona+BYpEaKT
Bq94Rz52QshaEiK+ovjWI/uv7I1tQme7Xho8tCtCtBTapkscsaSm0mBkdtBGl9nB9gGMYrvAfGrI
QeQyzY+PjTv6D6ORBdOiG1saQlNMwUKmT5xpF39KQj2m7kxgnnaZutGyzAR0Ju30HdmhfphnUX18
qCa7mRuuYxfgwQmpT9WuyGp4nauwbHiy0MQRHT9fEKjxzadh/sLAheBemmZZqVruGGvfSJqcUnsW
N28Zj72DCGApfrycX9ThSV3nanX1TyEi046dYkwi2aL7EFdN2etfKgZQPh+d35G/i/LYO/BBXvpM
r8zn+DEaMOXEaoClU1TBiyvehetcjZT7jfQrZ3IIkPtdPcbjfwCk3T0Au6REW9jdss9PXuqt4Nia
lkgM3m0HUHu63jDvz4b4VhNDfedUY3o1J4tLnn823rR9j9VKpmpnxEB8ULtb1l0eH1p5xak5Bgkv
sfM3muc3oimBUUK+P1lr1/NbfvlZT2W9JQHDHQsKXoAM4M9qQCNwQJi9m30mIXyyu2Wetr4iglj0
9auTl/ht3jBaytaBR5zIbewWZQm0J0g9VSBH5Yh9uq5xsy8StTKPl2Xiu744KeCIdh5XQqyYX0TV
jRkq5GFMDAgW2MLlhgH2C+ohN01AAO63VLxT4wISlB9k0SZdJYcQ7VCQyU54jRFUqdJs4dXB/BU7
z4qBTucl52F+OZPa4WaXSoh7yqJ1zrotB8Rbw1iU5g+dCLHNWU22nCoKRoSUp/Eajan6joTFHe8K
eHx1xaiFM6p3cBs0rP3TobdGQJM0ISgxWqFQX0BbYuDkFMVLkzLug3MrrSm4QrLRa2gp0Y9JYw3l
M09yyZwq90yNhJX6DAK1Ri5ylYIrUcG18mwnnbLKpj8CR8FDmnALm+Cbe/T4ME3sqsqex/IZo8Qv
SowEB8hBiryb6EVEZVc7QxjrxHzGV0pHvDvT2Oasv9EC/5UmsChz3eIa3mmqsrhgDO5umDZ+rHei
AxkYBRSooLZ2qDzJKknxXxxUPdjk5f2szZncq9FeDFazzyt48ZuDCND6ht/gGLfh1oQD+xBRRE+v
aljik1tQQ19XCcwvCCwYuMPyFrR0vurKlxwIC/Qnn9yfR0vzO7zPpYgJsH77g7kw6aHjtLFLSn19
eVWBVf4jQrW8BglhfJZQurxwONd3WAh6bTWPhdC7s5dvfy9V0rpgB/t3umIF+eOgeNhIaJXCGPPo
T8Bb/L+KvGXG1M5kB/+3plCQ4ZYw/GNe+DLz6QhpxsZmiwtkuSmduKrI7uxQOHPe8mpQvFfBsbS3
lqu8fUxHCzoSlfejsFs59lvtqiLWHyjU0ctz18aP1syKkFXWHFUuPk5a/caop3f+arLqw/0SChlL
/nAmIZ7KE2jYYW0qZoeylnBn6+KBDBLdiNgdrJYMrcj/Z6NoxOs+QwxKWPYmM2k5S/6PZzoxk8tV
yk/dsn+gjg8SpZoxr/JtLRWhQBf+oBlzEd5NldkhZsVh04dR3GL1XMqTr1D7taM/kPaSwGS4eo4+
kkakwnbDy1nCzYYRu7a35UPFNm9Cs93czUDfIwTojrtXmjV9B964mEeWq9HSshmZ/lE8RdSm1uGl
DIaq7owbsCTPbLCHAUoqWFm+8HhkCZbbZF6x/S/YiCadtu8MaUOclnGRVl5WfjqAJXRoL/+wZB0r
Nqm3tjoDDP83Y3cAqbuMs+FBZsP5eRk9JHCQU5uiQPfZzAiV5qVgoLjKr4agN9OAGyfLJvVw7JkN
dZHfZy8qsgvJb013jxyv6/xrMZU651FipFJOOZp4Uen0Va9ETupBAsqpv2X9a+p8eYrQm5jzdPPL
ruAj4me2avLRF7ByEOMmTCzUwxnFZX0kuC4sLOXwXLmzb2xWTVBcjh89y0bDhOmT9MTQsFR7Np5V
Dlr0yJPY+QDow3okEqMqYhymaB8bjOt+hdZ7WvL+uWuX+k5KETMTXLTlcjGRqoAf+o6Lmg6jonnK
fyPkcq+h9KNSlXvZ4i7URzAxLkyipsc371OmlHkI8codNSEYWonv0Io9ytL0RINZgSKCZH6K5zgk
qD+5GO3FFDgyOy8AFdUzanO5uieZX6fuysOZ5Oc3/FUdPGElmPmwoS75155okpdSqrhSiKSeQrND
HGHk7+Z5xY7R+PFG3/DUZG9UjPceU4/ybgSA64LeBg5gcqr3bOyndytXaFBFXKQHreT9DxSucpla
PBNdp/M0TbloiwaPMTf/+FRe5Edk3TUVyos5ZQLFgnoL70UThrVgGVAMNi4zcOmx8sI9PzYftRdy
a1wDejxcL6WBdaQhsQj4MjegAHgw2t02tNB+w1Kdz7UJZbXfke7O94K1OweEA23XVEJsqeXTJe5i
HJhyptoWFYNpQBhJ1UHDGxR1wcWeYQ3iKcDPQgM5D7xXys4sER7Gwb3lgHw2za3Ut/hKB2Rq3EGr
T5BmRrhkn6v8Ul09Fs/PjOsauIlnueLk5YFPqBor8Put40emqmgEM5BVSE4zY5Vkzh9Wlrb0IF5L
AXm7iQTicaJzK4ZMGuf229ZkAq2vYshbdmcsowDxGUi8CQA94+PK7TUJFcJefMKv9bGUZzCoByTx
th34b2I5iAbVZqlL2+ya1FEOCvDwcXxYE3pr19nSPbszO+cTLo3STKIfCfUOxnYcBBRstRo/nXi7
v9K4i/g+76XPsEuvC1A6u4GLQgRyUS9iRsO9T46EyjFHXSWfU6bsHA7DFjbNFRHjDW+6IuVwy7Qp
JsAaKxUnS4xTpVe59bFozpeeUXLSJpmIweKv/hVIhsdtBMB6NaW+WaQmA2akFPg6cbGVRrTrUvwj
sWHNRXqd74z0Yz1H+k3qdtv4yePbq1sjW3KYOpXWl91L5XZKCnFZ5nSunNbpw96ymwjeIVFKZBXM
GU2QA6da1IjY99o7f/dC/S5TfRcun3fhhvskuFb6K9zPjeW7rGny/pWC6g9FlICphMEKIQaT2Qu+
9htLbXlopon6nwFEgxxwKVejP0No3jIlF2rS+9DNT2ZQt2d6vnDlqMqa2SzqoVQrqz7N+nvb7+AM
VlvhI1UHbvV0zlOrCLH6BvAB5ZSU8ik/YrUhrEfYFGX7k+rLQANy0cJSWdYxLkaYfnUoS3xIuRHP
r9kWMNP5Tj/fJdIk+MvkOxw+u4ViWWgQj8RZCXcpZCxxJiTloPWmAG0NzhBiaWuhiq0B10Eb+0SG
qWR8PK5TL02OvXqZTu7HGm8b7Einrvd3CYYz443ZqjpA038An/DbKdYONUooJST8YPlzGKGgpLBi
PsAISfSjfxg5if9/ly1W705sDO4VbGb9az5nzqG1qPlP37qhNCVIqwi3AT+vgvbr4U1nHrq1MK8t
jfvLM+wDxh0cfuElfOhuntADMUHlE8cMV3fK0ItDes36CIVMrGLqGNefx7Tl2mHUfM2bnjwxhTIr
9ox368NqJN8gHroyb5FYLyUGUFzHRQt9o9Lh9EIEq/zllI6lpIZd99I9/36VcHxbLwar5XfuXLjS
TOo2/Q9wz3Neig7QaFyf66Za2Oq3cA7kh9T8MDObiZZV0GZzaUdijZopKSVX+jGxQZtd/SZpNBsW
e1b57ndw+PNaHP6VKkIo19mtbJBdu2cNCzm1maJsRbphdJi0R7yf8KVe+R2h2fCzPbYxaOhGNjpN
4xQ0MWtcZiqqDKoJBfkF3zGgFz2KapZK0XUrcGhR9Ky6v27hafOQoZoG9okJccSfalp1a0JZYsc7
r8gjlK4v7QZVPQTFDKYsLt1XcFcaEo2ZNZcL0WBTe7I6KQCh+F3nLiEg3paCQeTSYMs/3DCtZl/n
xdb1W22ujRvM3lLluWz8evFzdisWZYXGNw1UXBKu7JOhUCjrM/IqpKTaeKjop7pkYklPKUlPl3Ia
4TlLgoZaIX377ShYpfkBHgm3HMQVXM6EM0jCwhfqBmzhgRCwUF+gv5JJ/YB+OENuZ+fBidRGUIu1
tHfdDuAc9M3dLmfLCsbpnoxX+klVa5OafvpHUjjJ1jMhrarEoOh+nMMRfIpAnO42LcmkIqQcUFvB
J8R9ztXvESc1AfP8i3zP9TGP0u8OXRVD8zSnJhY/UxDxKGb1twaq3WikMEPaA8HtxVjA33iUF8M5
WzzhGhq4ZpXf+PJlzt40Z9zEwX7BrNJgh238I762qJvt6LM2G1eT8rZ5UAUfP17TuiLSHE5j4CLZ
0bIRhHTEfEmQybyJwnZKo87EaijUQO4vZyYfyRtg17rLZZ0BYlITvTjO9ojNtxBeQLC17RULHjg+
W8abzEufIjw8mr3qZBRjWQ8hRjq4AF9aMrAHubiyGuQay4QAv5pLIe6nxv23Qd3qetlbTBicwZSS
X8uKdB43jrCoSe7DKA6N5jaaaRYqu72qz/4fyqVUer2mDoxMDem82pVTM8BIDjjK8xKQGVARzBFV
hMZxDhnhc2Vgo0w4ZqUS/DcqOIPupvV2VApHQ0edDSuSPy8sxmoaJIPRI5ep7B/0hQuKqnWSs2gm
6rAobJH885NfXXkfgPJ8Duw7LYaTal2W/BuWak/c0KvUtNybaorU71fL7q8GqqAdyn39kuYyntwU
VNwrHg4gUVNw/XItOFqyJGpa/tA/ka6YgjThRUD/izdiMg9mUVT/G2X3lOLRbumhjsPKekSJkBx1
9ZakTX2zJJDV56qs+h07UiEF2/eAZeeTNTf/mvG3uJyBqc2BmD7RrXywFtDnywolFTp32eGgWpXp
7I2gIqAjpgwWB+NavGY46KOYBrsUK4MR+w/tB3u2JqqB2/l3dQL0ZxoeQuPoexp6TChvii2zPXI8
3hOzKQNp9EKFlzaQjpKtRJpP0ruSFYJADoMNBVslgTfI5VvxT5RPZZ9iTCNARhCI86kw519iogPM
7/ROLoAy+9rQJWKiU8iQXdaTBJJmbktyvfCUPp8/xGVALQV4uXJKmTHS0Uyrs1flEeuRpZCKbPJa
bppjNTTf0jAr4j/PR7eJnP2aGijdf6kEwvsdo2MahqNnKg6URjdWf4nPFeYbdhFEIk//JuSTTdCM
lAKGrChdQGygxwurLkExJyBbXHjUHRbCv8bHzj3abiqs4GQS9uAg1XjAysJElMDm09LMNC56NpNo
o8QwlUTGF6yVyvdXkFCoFf3hB3+b0LLgxrUjtMJ+khabf8pWdLmrHvdDw2RJgleMknj02GCFMeN3
5I5vDuv5rhrAaBEAA1q9asqxDF11hcjMFECLlhxR4N0v2Npla83qbhbgGw1oYvDJewzoLg88o3hq
qw1GnfOxVSjEq9mTDkwDzcLIviXgAWzXUdxV6mXwd0nAqZAERu6eNagWe/7+/o+kEf5KIQ7auJQw
B7neCFTUuBXhU5CBkVqWHbVmKEX27ZicAt9pWq2z59d+GlsCUP4oZ2soVp1IrOk4tK7nan7sYVnF
2o3R8/7LJ+3X4hGLxG1+ZdokIik/vj7UTXRQIHt31ltfgkj1MEBgZ6W/gTH9ZLoRu5BTH1KXwWNI
8a6lOLo/PuHMIJqlI5jvIF056WgfuLniiPmBNvGdgciICQ85hdcmcVaL4iOA6Xjo+SMdnYH28ZiZ
8F5of1spVKMes+82wR8pDmVrYHxpHRZPrXBSAyFGjUMeLgNAoflmpkRVrqm2TxzJdeUMsFsx/T7o
C6EYT/f7jxmDjOiA455R1BPRo+AnqeY7sYurCmGemvdGxdPxCSB3h+EP16VW3RTKoe4LlJY2GWa1
3/mECifSZUSwby7VN6A6BzLUssMerTwFiupPnZ9jZHFYUBsZ79tDUe1lkW8IUM08s/1M2OF3gqDT
HGaWBiM81PxEEj75qfEPb7Y0Wnql29Il3zmjwS8+1sCuQ3CdnZ9Lj7a39iHiajWxl/tciJkIi2SI
sKK7TM1PLn+XIRKw37Qx/sK3vbVt5cAehBMJzq4cC53fweBuVfIOVohIhrIBnRHAJFg5AiiDIuic
zObuc1jT3gIZldlnkT3KGGgZgMsgCKQBph3MSDysSiVXyH9hL5z8IUF1FvooTiG65uB+aFjOO9aK
ERX6ypAlCzBuQWbRG/MsCIQP8LG0CtVCQVvfCYt3UTq9ue5jeMcnHCa4Gzou99jC2EP/TBblibJR
s61LB8NFOvS03LDVJ81dhUer2lmvowXOF9WpU3ZWt03CDyZkix0i8qkH67r+mvVacDzju/HE2VH9
tt8b1tKUnsTsGrTl9V1yZlSqA0Li/IXKLKswmByFiz4hmhxXHJfWtS0uBqC3TU4HLThY39MAcdVL
RNWEipcRSJi8EVnwtl2s9jXYheQhn+xhryCrYc7iBw1hTj0bNt/HPOcagLuczO3p0TBZoZBNZ/2c
aJE5hDPy4jcIS8Zu/RRnB7grAB2uCFJsxDee8kUI0bPE5HEGRkUXCuffDDdco+DQN6Yo2U2+XDGA
WGl0u5VJfHlivmYUo0D1amW1W69zoI2M0R2PTV4jq/G0D2xlp6U41npOcScMU4FwT2pRAiWgAw95
YLTOEdHIIw9Kxopfc1aC7/CYACPqkjXU8+TG4CltS/mj7N70cxo1UU0+Rgm8nRIJuAl8o5LFX3qU
n+s0mTNIKF2Maq6EW8Fz6y7aJ6YAE8L8F5ilx6+tHHQY/xEHBqJ9QOcFSSPSzNgHc2juMNOwQU3T
4CMSKH4PyAjn4IDhLHO1C3sWTVU79BE1+qpzq8+n8NueeFvS8NTeWY1VNqFXqe+KrpIUj/MbOkkX
ffJL9Hc/NqOxhGV6O2H7xSZfKocdydXkzPlZFvzgr/Uk6E1JDMVXEcECU+u1FAebLYI4q7ohSlaj
IHvy1Pw9uf74VD6B+4oYS/hf9hMRudytG6/14I/dzpkxRLqjtQ3mtFqCj2oJFPM5KnXLGkf/f7tX
JExicWi9lFz6K/Knfi4XPJ8B+0vYXXaasPscZfBHhC+MMltPvS1xKNRGty2JndjhF833KeZgHic9
dy3gBAgn6u+etN9+nQxTWSt7fCSGwIk7vEotmWeat2wHo5WosrtLIDeg6LpYMBztBmXxZOp+5a8H
wo5HnzklzRIw+ugtr8hIfo8+YStkj0mqbmAI7pYyDo23fraN6+nYG2Rfx7BPrWFW7HnJKqDeFWb5
G4VZCxuC30h2JR4xsiA0t2z3pxjQ8p30i+xeS6Mj8Y6GHEiNkArh+rIv7rtB7jEB9Gcs/JM/EQ0+
TsghtJWBLVPjFk6rUe8+hbIHojiVFoM5vEl67cUiF9p3Pe6ZzuRf+7r2IIh9bssAvMvQjQ0qFIf5
/ObvOP0r7vU4vK4a1mowJj4WR+jgQU+din3ehAZ5TyV+HH7VW0z5TO6BJZByNERXKMvjDKd0okr3
dyCRa7AFDEYEvAvNsuXhNPoCh25X2ZiQsoAu+XO+oeuDZQaHHc74swG5jlznczPNJaSUM6v2897t
fc+69VJVn5Z8R/ljWaIVXa09UzGK0irwDVHCxvOa64TEkq06IygRNWKQQ98/KH8uhkG/bu5mdYq1
e8EO6sgXI43owpNGVkAfO8CRm46Hss0cf//qjrG0WJx1IsQ2BdfFMpODFkVS6wFtUVR4OD1/04xV
HOGvNR+GI3aToGFgwiS9qS5f+zFOL/TXFq3U2MZ/ASzeloyjyA1G+YYbuWTiVTOoNJGVDECaRSWT
BU9gz67WDO+ePCb4Eed4KClh7101aj6CKscI46Wd082StPrY5SPcxaYUX/ogvoChcIYcnY/1HdeP
09sj6jmxv49M+Leq7/SMM5cPQ96btImGX75i2BkevbltALozl5dgUqRmkX0HcCYNrQC4wDkLG0xv
lewSi6HemHRPlSt9FWfB1mKjzADNd2BBPsNFJbPyP6bKOg4g2ooIWbKD5BDVq9QJNa7sk/G1dkJs
+Y2+NUNq2DG2zxv2cSHDhRdgeYKJlyBbFZhDLd+yc4wBDjrBi9S9FLJJfozc1zQGLo2YUUL+eMH0
1UzRZXBQcb6fvvFdA+6pB+s/ENObKPB1ipbQJHua3+aHt2Tm/0z3SXeE5igF26Q8lS2qUeIbh7Ke
20DWetqRO22z/9ae7I1UwK0AbgZAkyLPbS1ofu/KuCx9EJwyxY2tHnWmCEA6uk2ZJ3Y1e0NL7375
8FnbH0LvWtYtX1CF2yndfYG2J0x2ZRdLbp5n/c/APLg9LkRfhU5cUWrLOo9zhJbUjhBUvLlpFoWS
C33W4uvJsoKhxdVnCRlKzeJaqH5XhPhmSPC3XZ5+Ps16ZGtq939jTlfgjX2y80OdZa1sINAXiKkc
Iuuz1uo5Fns8TxiDjPPr6fkLhsgK+/Cs7Gty2MdoaLn+eVJoX2txypKsnW5ah7dz/2POivrTqwyA
lZ6unRq/yZhg02NhUeGqcGfAy/1VFVuMFwLhoeLoQfA/I1dp61aNtjbAsVY4ME0I5XtJpFH7lU4u
iRYNy/vZQj+uY1yPiKQ+UsiTmsL6B0Z41tpz/kQCYes2nNEhydBe2reOGnRHJcMDt926EuD/CR4g
TXRnImjC1eZao80G/WzN/tCLow0DNn2c2+yYJzKhPB+N0nbBlVUsd1a3EdAOvPKtoYsfZn+7tGz0
hBltaT7ODCByBo559ooORyhW0IKWl2CmDkk6aYhaGtOHrtbClThKJDXc9dA2yDMtvLsM5HPTGv8/
bXD7rCkXfnvXSC/0gPUO00puT+i8IuTJ1xWyxbnkWC5n/HXyr90uOYa5pO979HCzzN+sJFcCOcdz
41SycSakrqfzS22jgX3IBHozdHnU/yUBYM4BqAXq7ESaNHAhmy9/osCCOBQAp3gNvbKJwxitSvN8
Wm+w7LmtTS8RzKEDDFM1zatPdnHYnu1kYU6TW/tao/S1WSZabRD6k0teYlL97zAdvtluAdloZLKI
tb9oIC8FBiBDexfWxKeszSSrVo0UADQNWq8lVGSXuzcKCkFgwh1N5Z92iyIau52yi08NY9MG8ZFx
Uy5pZkWor307zo6scxz1sHGK7p/9RA3iwB9GbcbrcySghi572Dt36DJJEhkul20+j33qvmFgJRM9
6cxR3OmO69ZzKOlDQ4bd6Ar9Ti7kwoMmjbv9n6tr6P00igFlJi6CjC34fbe/ePE/aCW2ixbT5g3V
ffj3pZxtdvqxVq0j9Nqv46oRUpdmgzLc1cZXpIVVJM2HqTmjbPhJjSpZXw/6pScvQpdkHHAQmTwN
Lati5TyWBRVwx+ZrNjjTLK7HHD85Qs7aDCu2SH5N4q1pwDYN+8pZ9diuSGNguhC7CoIxc5u7G05+
6zGK+8W/dL4sqfm/o1QJ3B47XAygzsWX4cl9rMa9DUgSCTxWiEVgqNle8R6alFdbeBU6VgAbotDC
g9uI1Rs3LoSnxCMpJqeXB8ioCJbhHTcDNGRitunONDt3EkaVgT97DyXE5eR6dbQ3W/42KF1n9n1l
R7ZoB01zlugjpzuY2x8sq187NOgsAQD68ypCsDxXhhaCrQ7Dc7cM6mEoyVKSsd8Uj1V53fNUKLJ+
5Qv84nFztJuHQpe9z6BLrO/aMVt6aVbZinqXzebuGDa/PJPQhodeQt0HXh9mkk7TuLeFGd/dFfmb
NXv1AN/6Bh0biPrvKUp9XJGvzw+9yQz3sWeMGgbCzkLSUSJgficIDUVDcnxDOL2XnPVohPV9Jccu
VqussQmCA1d3qVAt2VO/s0CMY3m5+Cc1uzsAzu1um4k3Av+17vxChXft2FbtkBaBnXwQYs/de5xc
BTI4pAWvzSXMikQPTFxdmsRJNPQAnWOwIRHXMY0Pe35wtUCfvpeZM0JEBM0r6C5SLPVOVMDYJ9xW
0DhSZwICpFJDM6HMqXrmm2vfnjo0oG0T1bCjbY6Mq3vFSzcyFpLcx27KXjCjXxF1b/VVSRtMajPS
eatdBvGJ6dVlAqlt9HtJJOZnJUPXZntQH4OkgeiVJntjJ9sH+p+LX6fOdY097W/2BQI+7BKBU5al
c2L2EpymoZagmF1yuOwc0PG+59BuqnlPOgFvS/H/0B2nUZyOg9KrwFUY44QIcQb/IMobC+euijIM
sqxAWo2FBcH0B4wxBWsc3Ip/nLzXPLzQ9bpQdYeYt8bcRbmo9t30b9dqOQ77EEmNYjwtcwPa7Rsv
NVBU5KiZgXLHOH0+HHa7XX1AdnSYmyNC+qDq0MBTUhjskjJvD6vLHjsTbXwYLtulKo41tmyXv7NI
JSsTZwMwBzjd9/Iw0k2N0ThyE51EFjxmqe8DmwwarI0saO1c85q0RCcvdH/+dZkwBLtCQASnVK2r
e5aEDRHwDhBE3wXwVyLr6Sly9Dz3mIDpsFD5422Q7dVusrQlFMZn/7E+vHdW72WzR4Mq2b8Xbi/w
iPQnTWv8OjYOuxsW1L61ZjafeGR1Eui/cxCWu6X1PG0SAcTqHc43Q8b3CqB/jVzH4JkKvLiqLZMi
nwfyGmbHCBZpocqbDjgbQUiFVS91wpZmLhpo5gOM+gSN8iju92EMEygmdDKiSLQeSskxtRoHjgWc
0Qlp3BzE/vaHwnxem8qim4v6g7UBaJdwk+Q/wKHzkBxOUCmvp6c+Ne0utVnSsx9aIT/K7aZwZaId
C809I/SeXDpk6pWJGg0Ubo3agIynzr8ZSlakw/AJ0HG3QpqoIWQW3S/Bw/WIji9DC1ykANQoQuFN
OIqRVHpBlWackqboBiOcibRkd6yRg02z+EJ2LP8U9BsR61LuBi+VWKtil0/++C+NXfCxh1b/eOSI
8lxvWTJ1cOPPtHqC9noZteQE3iP0nq0ytI6rP85a7cUH8CrPA/GoK6+4ZlSMnhhFEDfSbpY5xRUf
VsXXM1bRunO8T4tv+Nkf6c/h8GquA+PZPBVZwwc3tNgE9aoufTm0uTNi3wHMLmFOdapofEawnSQF
ogOoXuTIEQschA0aLdt5Ovsd0Mngh7qBLGAQv2XxM1ZdErXMGQ4c3BYkzHqvohTyn0U3PNml0PCJ
8Pomjhm3VmTH9DsfvMTIPo4GWaxWw5/ZeQrQt/2YHh/LaTvJj2eYV+4fclcMDNo3T4xS4Fjrzvzi
AXGqjqVr7M4GWj/ON36GH6oaRm9caKji2ZoOYQVhqLXYAFBXZ6HfL2X9EYsajZvZwR21wKxuXwyL
t903VkDeaDD9pkQ3G+OPCwC0FRw0zgFXv2fYswkQtMsXZrGKS4NP1g+GVNzS4VlUAVjPCR4I9uot
x+0VsYbO8vbl5fSe/uFJMO5fe84CmPnozIrOrlGZB4TjQ3arFmSgMA0KgI3ks4zcWbp/3ITj38RD
0KCYFiLQv1cCKQi4jkX8FUcYeJpqhZPnXALiE8/2mWEHvzAzi32CFfTeBTx+z4Gp8bfd2E4ezcT3
1b34XKFRBLQ/Gd+yWrEIQR8Kgeip76RHPmmG/JaYLWqxzvV76inCHNtUzkcmFsKlMs4FtxtEkiqZ
jwsbaEj4S3MCxrX8/eStxhzphauadYxOjrlb1cgM4XsmMALk57L2Tj8JlPKb3uK4Dbm9nFhydc4L
hUk1SEUWfvxOhJHs+HzyLfbQ1wd8yXicKpPhGUaKgyOBTn8OMb7Fyq4syA4Huow5h9QOrzkl+jAw
z+zi7g1DRjQsWqbOKC94dt80pkhjaCY8E0hwpqM5KrxVrHZOwSTAa1HHsX1TB2qT2oV7xoJJYaDN
MTKqjrGvSWAfO44E2VTdgvku7NSMEqQstfOA+G74U6NV3KApWn6vOjV1zFD7EF1ToI/rGioPkHpl
jjXB2snEztHHuiFlXWqQh61szQtmKR7PNZhkg0IW23P1fW3AugZ1UnzJfWehkj4QzTSf+lB2UwmI
V5vQ/ywa8i8TYkKZx65/EK0WLQn0Ggm2wZF9uqYQh9sPZoaTmnTHbwTwy4UWq+WSEhj5GXwkvVcn
wmPMivYrytSU/09vLQSKhDdSd+nfw39Mwlmp9zRRrvYNBYjTuSXVS0F3XbiECJmcr5nBB2AWPHY0
sz5FSp2vMGbMKS06zQ+I82TX9MC9STiOqEIIDmcXwJMO0sasSx5vKOZ46PHM/TGeKbrY0+Q3wQ9T
fXp/ofo/moT7/C+xYinkuQwG/T/TMVJmZSp7jCA2IHIP5QMPwGB8L8lxUd1FTTGZLnjmrkmfwW1V
Fg0j98SYEPxpJ31ghkMG3KX0xZ2CiFdP86w2RycjQRcUHuy7JBLtYteoTJ+e5ZKFJagOcgshCt7R
GE8M3F1z2CVmsBFEL1Z45Ie7lH9lT8llKeuW6br9WK+9OyEs1ukU8xFXNy92u7TjMpRYEoJGPw03
v4x3q6v1plPXOWxfx8QZjVVEicumgP6/69UUGObnClkCpXsUhZxyy/wtln5+1CxLFAWfEkEIB/MM
4sUnh7v7+6Fz/wS0DzZvZNFFyJAtD+8KUjz6KLC5uIFIU2p7+67sGis1Cuo035Geddy01OK8pfBW
TtNX/xuWr4YILeIMg9pj5sG5MENASdjiCQiyPlsUfdSZVyXFEAXLcIcrQgskbnasBBiJbDDO3WW+
Z6/QiV34xhWtqO9v0ekDCMHcFuakTqNZcpFB9o6DW5J0aSRR/RhE5OEs952dpkDe/gEM7Se78gR/
5HdNetC47AUlnXNHFY5S8TnsCjLkMa51EMSMrwXJaqqbwZt4vCswUonlOgLAo3nmLmJ7DTXPAe1A
HU4dtQrTjUk+KmVX/K2idaXOgvofn7xhgKCPMIqvQ8zxcMMkXXDNHoQXOlmLDxEtDqi9Zp04n2tb
/vHuFyX3Tq1OosP1MdJE2yqNQFwDbiyKGH5Hu7sp29xKzhI0f2oYA+w2HaFKwXVsLq3ZIuiLlDyf
xIt9U3DyGR8q+wCIGZqrBZC7g8ukWJHPo9FieGAmhO6n5lVjFGaUoaAjH0xC10adKKkZOVK3Y9OQ
5xUVZlJOK78g6WU1A3iCfsc04f2VWdv55NWMI7DeFknnvkMKq7XIlYnS/E4RFrSSe2qZJkXICAqe
b7JOQFPE2akYqyaa6IiJo+Oyogbn0ymvgDE6SY87QXOXk6sT1b/w/3oh3reSP461OYR9kILPkh+c
6eu1lU3pMHSHsQVTt8QClGoOUwBRbABQXn0qwyg14f15AczTvdBMM0nxvtOTHq6OvHFPPuEYnhTE
1tSad9i3RnjDw/XLR/4qq7x4ZBVIkbZO5Ixo1ErNGX+9t6NLowEkmYEToPu6Ybw6Buwb7dsTbOKV
Q9L/0sxv+gKou56V49VHrlIdnkAv42/4YzVfFoBbN/YFCIb/52dScx49xClZSagAV/HVSLXrS9SB
K9C/wkUVwuAPJMufdctdyXvDvdDoh+ES0XoVgqAc7FGKBdm6TsGRkcmfzkpf2ln37ZavqOTxrWG+
PF0YenKmE0ukJMwPOOcIvFoEfoK0pydq6e4mZtz/y1CIlo2MlMw3KSRu4JMkW2fIiYdn1WFXFVaH
5BvaOUJttnTGGP7xH6FZ+4vEYJQKgw5VjgTRCgM3CThF1XztVnIjv5Pn+uU4s71WpQZC3Sl/YAhj
9HCrWWCTeup6d+8x28pEKz5I2gIGrn1HQMsgkWSPO5JbTwkdBc/qDM35NGw4zCtUyr2VkMh2hloy
385tt8DsN//n99gtS+nDhzAShbNjvV0JdtU7o/alKYFGNbs5c9sc7isJjuL1aZr3uQAqArcHHhgG
zT6625PE8IQWdnNWvDPr7IDI7sE7s5DYESdrRNtj7uIS//DaPJZw4MgjHM96X23wuiWKrLc4/f59
8nrJJUHLf7UhLfZpWaDo8jKwBzSOMMgrr632nT9CegRvJ+Vs0wUkwVrm96ixb0/I2b4tS3KDajbw
Lfh9sXQv7QW4XynzhcMiT/OkIoPpugNcTFSttW8eMVCVuA6Zk7iok6OK42c7Yi0ASXdBKddvQviI
q+aJ6CVykWBZA480kKQhCFDUnqU6dtX1J/lMIWAuzO+HxUDFOMXbg/2FydgvouDk0jz6swX1C5rL
NMvcZxM/KVU4P6QLxt/RdRhkaDwFMMkDSdGAYtCXdncrWyyeiok3YZofoqYoEYDS9cKmHzlhwg9p
DTnIJa2ANgL0cJgPUNuihpEtW6ns3zyg1CX1H7wfE9kmFgEFSjOZMZFI0kAS7y6XUXBFK0qYDuTr
ETQlfEM+VeL1akXms9vokbnjslOYPTs5VmNPJmYNKMMPhFbGKIXCX4euB+Glrjmsi8kqLdUkXjEB
ti8xR0TGu3CzAna9YDHhYjzlVYw6iwzqKgs8I/cydqT1QSUARLH6KlgU67ub8rQa0tvjwpz7aLnj
ZdOQkL4R0go92caqDz+CdNNRydQxKnJalxGFtMTuDL45bhdeo7Z1I5jKoTuhf63H2FEGV3ce704C
ezkbapq5ztE8d4dnIYz8CKbo9rfui/xEsIpZ031swjWbKeiDxZX+tfEmm7fw68u/I4jJscH1waZ6
vBD9r9fE3KSj/bm6NznnbcHoaihzNTqi7NKjctDhMb04guwF5SuZrPGSmky/RS9SzN43yNHhrnth
sgZqi7dxta8UBXqJyEbX1dlQTQ8wizkecoBSePL+isTa74cPt/rKjbwPWuy+208KhoErG3zeFc3n
vf7jhUPwMERlouF7AsTwE5Hv4oRJYVgaeLhRNVoN5k2z/ZUzwMIAMRwJD35+f0ovShRHCSuHpJ4A
E1v9TaL3/K78NrX64gqFeCh3wFZ63nSoI20zOJwmyFDL4T6dc7fI2KvKXYog9L2ygZw/+ZKtjLJH
dTfmHOSpe37MOkK5tSjcfAYtGl5f+jHkieIch8lu3MOhaTzJrW1w+UjC8eIl32AAYPGRdgcdYEvx
PtOefnvcakew3BhW66jjoD7Eu61h4zgNLdk87OGtAyIptbx8c83eqxcQpsILpggR0a1cKcKjRU9o
5G5yLRNawBklMaKksbjWsh7NoHo3Siex5u13gETWNoKIN2PjAqE0rnuzk48sFZ5ja1iAFkF8NSWH
AuEYUwjrQa9/QwumgSLkYLh57GLbEL64enoX7h9pAgdy5MTkce9joIMrrJDquUI/0Zi+aemHqDkD
eEjJcQ/6gtiMyVxV+ncJQcf0pv/GzRNghc1t5nNnx6Ub/ecCjRAza0V9UlxvTJ6zvk1xVhiFGzjW
gszGTQLZ4i19oAYJe5FsHdK0qcICgelTx9CKs9SV01sfU4YJKGdNtz70D5YpjGSJmIVnohxYdakC
xgiBRj3uxgfFrLO641gEXboyQcf1aSKNF4vDisNoSzQXryNxdeWOiobFBHRh7Dm8cRtiYw2DluNC
jUsSJ2aJ3CNVXS4Ea9oNdt1KixoLvjd6NY/KLl7j+OXvBaUkLoyxbf97EPri3m4dIX9cqd4Ea41e
D0JMz/3gFnLC7YFKqgJvgwtU5ZZXZZQkk2RxUU4+m4mj5QjqY12TdGWO58HjF1fMbXdPk12IwpKR
6Jvic0cf4rbANrbpr052th5vLrOHcCSarF9t05BaFUVJMgIuq9Su5+2j+rcdW2yVu5A7yAn7pBfw
bM+M/kpAFmABWZ0dye6rfGWyMQATK/T/Uf995hTyOlYzUQfgX5nWGqPAshymVYOVR05eiV7sUufT
jw8s4gAbpLcp42ferfBy/i4VuMTEe3hWNgke6H0EdHdHKpQGv7ahqT0zyucuZ3xS6ncrXdOOaNZ0
y+fvZihK/00hyanaHG6RvioUY6/hOnNiOaNgHP6qyodbHFMSEK9aCobeiV8ABiMvOf+TnYr7wFsn
Vrgd593nGPuzDcBF4xckXYIJL322JbetdeFvS4hjke16z4YGVOXf7CfQEBcUpReCDnCbvYqCCGMo
MMUnBqhLMO2KFPXdCXbcBDLnwojVdXelZv5LqIaQFvWECIClPDReulOBQoNSjGJ40LCAZNEzqdeG
5zcV1qVRD84qKn7WhW6IW0pZYiYC8rnfa58a0pkHhsnS4pahNJ6URgEcgcTO4A4Ez8mGqMztIy5n
c9qGT7JBXyMvgNowu6CarmyeozXL02Kz666abcdsrAyVWB/2EpzTOUh0PpK/04KreQCwELSpidQx
iGs9fCs0EPiSpjMilQFShx8dn0CT9E0BEfGBiJ0Qu1xR+piiq3dRIgACSE8l1PDJ3rS5N6pQKS5s
vA6jYEtMvoyKuy1468vcfXqI6wy7RUM5qsB6ELQXVfRuo51d/RVi0+U6nSB6fetUX4eMbbiT6jeV
Hlsjb838eQXcJBdKJeocrZZwG43IsFTFK2l3Lih4bhS+BcgWzRjY2itP62DessxUL5ixMKYreQ3I
bk1JMzbS+86B5oEbCVBPF9qECjRNk1WIsXmCUWU+wCL0oMTaW7XURaaYLVd9lso345ufRBxQ1TG0
0qy2qYRepZjOe9+snY8Xf536rW59jmD910L74jsuI85hP31C1bcQWc95cuHJrBGXFVFbLXUqlIE7
Uu9Hc/Fgav7OJpGic11s2jUZMBwT4Pk4+JySPuJKnBvGTurzRkz8xqByAOkpwncK5nCaLoI+DMF9
r9jI18m8ZJLBQMzOceZ15HdeQqBcXfD/NMEhgx0ERC7w64tQVhjodIpACDDsH8lV9TLsf+uWGgpj
Nul7EP/J9NN592Vxt2gW9TlhIJF2Y0+9lBSnnd6/oxrVwPWTBwYyfgY5XCNlI8rnbbDvKLx8QvrZ
jDV8KAgYeonvOHmCYJBIZFDSwFmbt80XQ9EZ1+DXvkwH1sIl0WO/3994IrfwRIV9/xkkcamCJKUu
o8PFLmrAeAYcnTreOlE0lGbhH7wm5pi5+2VWE7fBOu6GDeXgbErWoxXSr3TKcI2pl+L2NLUuu5yV
wZRtC0A22nKDEDBKS4X1XDkc4cpYYFvOIQNETxK4rTuB9T9bLzS+/s2X+Q3uUnwfxTIg3C95eFW3
MQYUjsaVisNKkdM5ttpccrfKzhHfzEZbSTwTESK74ENZAJXpcY2MQDv7Rk3xYZgPIGL6b3XfmaPk
abxf+D2tmxJChSjl4pydPFBfAbCc7zb7rZhIIjJD4kgrXftLg05qrCUnshCeWJb6UrFz6scpHWYg
Xt6XI/dKeqjSEFmZSIt1RsljLr0SlobhkLTEeir0juJ5VYM1P7mt+iI/5NLcSEDaegFB767gnwq6
tYMqh5fQFUwCmQ8//RKhHK/Br9v17Dq7mCSSPh3/pBTH3gcg/rMxJzTSItD3MWOvFDPfbewrabSJ
wFRMyqA6nKaXIx5Uz5XJVQ3KWgd2yPiyOnxiUwPMaUwak+CnX/mDBLJliXm8uWldkDRBvRPVczJu
I5FrZ25R+25xQVuL+1hFow8Cnm065DB+y3a+VeFPvplnYaWqvLdLCw8d4cS9wIHGXsLBvtF6Ft+R
c5LJtbKG9qSboVMBq4Q6ZzO8cAviERoW0C5hwaqJgc3nK/+iNUylYU+YaQ6j5RuaEwsB5KXKLDKm
P7jDkaSUt6GXZqain/q6mVDCyjtMgef4u9R478JFG4yFmL4S9+ltHv5XsKF9Xw7qHZ9WsvWtpAz1
B3+8skqL3Rq2Gecgghjdumv4lHihIUNgtRom9WQAky9yDAekrrEXv7ByOap+h30oh1IXV7gp80MO
6UW5ceD9qrU9hm9igWDU3vfTAviTE2/jnrQKSAnI5FVumtBQYcDZkKasMf1EP92DdhWSIQqQ4i7u
dKz1Hi+cVi4fZLU4FEkV79YbK2G1drgulKr6FPhXioOtihWnrxIJYAmiYXx26dhl2QYHXjN/qP+O
n1dVsrUaYEfknGArA6odfEOSHZLHc79Flox0JP1Z5n/LcQgQiGfp58VIhbXVdoVGxM0miCdSgjDp
PQ+ZU1YpHWAuRc7vjwGpBU2hH3JwiGi9uLieW7qwK8sh62J7793FPK90werG6xvbsnLcuTYmCDCB
M0uBPbHgveRK9qBdlTjQCLBQmkohLOy61dKcOxR4BmOqXJHoCsYST9nK+2NivZR8wUPHRvgTNOxs
Be6jWJCZDSeb93EEjkToCIzOr5pECYNdK+tQ5RBduZt6l3XsBvJcx/mJsf27hCCJkQfO+M0GyrHq
BdSMSj05H9hqvdk42zkoUqsLpPj0kL0Fj+uFJRndZwlysT6tyvHBch34z6Tapjm0TdfhqrGmswBp
DKiBGJNZmlvLHHk+VOR7s2U979w3AjeSIJnuKIeNGRLRm7BywapNFDQXyhnzR+ExFlMzH0DqimEb
/FS/0/AHi+I+kPDlFWbL5c5xK28miYiw/Jk/ucZaYe5NSNGx15dwUVGf1RD28NcE1KywPQ7qhBV+
RcN8etIw8J2YqfGSUT8aspL/ieeeMA8djrgXZYp6auOskEqA1G/Sv2qGf9qgvbkvcPrMkWZ38AZ6
COulSeMYjI10XeDUTF+w6kS0BCvrKA1EmPoyLwfNdXh7K4rfzI4WhoySehH0ozO8FfqQWmNwj1TD
0VqMJ40UtSc48QFNHPvYFrns1t8U9TmYuacZOb1wUnKrZjN3g6+KHUP+89IRDEFTDuBYeF6TRvGN
Ti1dgaosCb/L9fEYr6kRaZ5ThwB64Hmhwf+ah2BxmC/AwYe8ktLyNEpg3mW5GZ1pOChla8de+XpQ
LY+b99bOWhNxhBvhnO5RzXN/e6aylEh9qm6HUoP/giw7jrO9gfmZ84+8/wqUT7dwdN1lmIHgYTiK
6wTv2D4YMj8cyBkhFstYwZFjcO4Ov2a8C/RRD4Mb0DplznvndUTOuF2a1btuMPJBv+J/4ggtcRvj
glSOVbGsYbcoN+ZF+tlDkxFZcf/ancCIsPbRjit6PSvXyJArLHmTUoasbp+x+t3t4GdKxFRxnrZa
DHZuZwksafRRgzvswJqfNgt7CF8uWtegmN6v4CL5+PfAKmHh40PUM1M3+gIfSO7bXJvfAVFec5Cu
bliYJCRgk67jha5EQyd/rEMFzc5I87tb0K6+TDyfTyOM+xtDMmDu9HuTnOBXLOYOt8AHL2kZJMrE
Q1BkvUxVUPTKGcdTA23cm2z/36SI5Qy5ba9vgPBvz39pfWPFeI9PFQiyMlfCVpcCucESdMgSU1bb
nePakjBRj7uArA54J3tGQL+aWils2WCnLUzWBNz/MlEZRc/TYg5A+7zn/ZWO+K/C+ECBPkjEOJZt
4d3OtcFxCVV2f24SySQ7Iup6sORILHBC6dNdXamSTo6377FCTNRMKyfo+Q2g5KmbtJFilpQm4OSr
FBTtjCRoIJItjmpyAmpy43uHwbe3a4aWcaxflLcQWbuJqhopfqKrOPMKMdKPDGLJWkE794V9Itgu
UzTWY7dAEcGByO5Nq7XjVugH21Sk+06D6z0eb9k5AbJV+fx11xCGSAARJLZw661sPzs2nyPOntbz
6kMkR/P1C/WU2Pz+X3xdYPu6uX+ltCa2VgpxwNrxJp70D5o3Hr42+7S+gEmT8g8QQ28orlAxPATf
m6gWPDLCLktRmfIRd3tTYkWCEbPX7PyGD/DiCwkYL3g0eDoqv2/pF/tuCuWGSsQu4Rp/N1KEhOUv
ujZnSV50r890n0myAdzk78/HdLg0n6oWLBuuVL0eh8+pBCzNxN4IH7F6abHr6izLAgKnEjXaT6yz
IadyVO8s85EfzI9YIxgm3vZymJiw04FFrJk4//rA314JG4mkQSWgwsLTJu0aXqMo3mJTBT+eOB3K
A+HbuDUyurAh8bdlFXlqwA8JqpOZu8JJuiwZuUoHEoVfXMjm7UwD13nLvI/NXMMsobJqnXWPJM0V
mIz19WpO16EkSIIfHwg8qdK0i8PtO/kISN9YibYs2vBpUIyz15fnIle8gMaG6SYk4+eDHTiQ1Aqf
7kwVXsw4k8kfu/yw+MQfNRNrCdUfvsqlvuRvi4GioTRZMdOraZbW/oWWXEz3yGKimxjvl9RHfSJ7
uAjHQabx2q7WZDNu2EI/1idqjQZr8QqzNQmnmxx9O8+2sHi8nA6Wud9IRVIe5f5DaII3PljnJDJj
5Bm+eluWjqiZjZrWQVXedgTYeGiShurPF24WIFouuHGpZAbkx8z6zMwith7QYDOBIaNt/G0D1VOE
PbkhXgSuyhBXERIY08uxngJC2vCxNu5ltfA6zSESjYhJ5RdrhkWj4N8JMfm052U1kP3l3lwn4bXR
926dedbqxJg9czwmkgN6LHQD73INk/NXb2pTdxXHKfaiEq8dVWgAjTAN0fYIm6hIYAyw4xDuYQW6
sUPLFXNNw0xt9+bA9I4bk5gU6rFoHp1DM773w+BCJtvtYfEX0vkg5UE8hIyDAyOUTLhULSCV+G3y
L8VMSu6b/mFM+cf6URMEpRAggWLbGmsN7ADU9dlTdTO29GTDR1Sgx/qc7m/6xCdpYsKHRbVleTUD
wWCPBJu6Mlf+CqD9/5XiJqtWkzU4OVUoSYBh5IvTizivkBwulBBsn0wNIvZN1Y2w+yEWxm4IziC9
d6hIZc2rIGa60HrgEH6+QHphEbpkdg0xwuTB06CeIuQh9WkYZIOUt6fsNoAgQ/0AR1b/rAUZXau5
jTx2q86d1xVfda9eZCBvnMwZlyipymCVq6TyYaQ6TAoev6tKr905k3K/3lszFHwvdrfwfHDgslfV
HXOCFsAD5mykG1fi1E4M5GwOTrjRNaI/EZNiFHUPhvZd1z0IP0ksQQEzFTqfr2ieUATWLihBmXF8
ZJSQiJm2P+4L44Df5sDZcOSqk0vKBIpXUTJu8QWmj5UxgYNgubJbQK9rlipp3YD6ti5jcuDO2muS
diRJPx4xkbMEW7QWmsuhGyXX9rOJ3LNJGx+11QqPt2NQTbrAtydzNDXHm4j14XPK2Nymd+uN+Fs7
h37aTVisVWLqjeqNF+0DLYJvkeMknYueH0amxMKyIiY4UJLLXM5iS862t8/7GdAj7xK8M5xUHUbe
H67CBKKaB+C6bzNYIJz2sKgKAnnFL191mL8FOovfMKTRtHxxRLEfvL4QCc/yGEOrVHg+lm1pfvxk
xTnEhQNUcx8P3g/4WUPqgseopbG7mjZm5a9/Mr1bANouG1FJIeEmSwyLVpzP6CHXUlMz0QUG3M0w
2aoQy1816SOzyUuLzW6LwZX7o3ST4htnDxE52puwezLfzzOJPOiO8FBN6h4RZsXjGCENeMuOSFlr
KemCn+upBjTiDtO/tk3Gh47jazzO6Vswro/aAOzqiSxV1qoyP4Nn9606vjG3PR3f3alaEKVXA8dP
7IXdPmDVSEJjbEu3qmQ8rBn1c3Z0zE3EefZvCUIaQCPBOUO/z/H187rQ2PXiLMuGBtCQ+l+UVNcp
hBrHMh5k/VSH4TUWG7+v49k9Povr3+9D4+paPtCZMboFE0i7/cXbYr0+lO5cWq8iJml4K1UE1MoW
+zB6wtCj0YDY1aIxrOxCNqDdTVOwGII/JO+RoXccNn9KDnNr6UpT5d2GSs0Jedp/e28mUHzcATnA
55apEsI4kgHJynOFnTZ7tc76iYrDoJN26C0Ty5VbM/4qTo1r74dHWkPXaGg0mHchohskTl7YYJue
IudT6aYGvTxmFrtOMDDnfKHJ6jIg8KfyeQ6Q/d2CUeuq/SY01JH3MxRsVQTIPt+pgnyftMywE1d+
y2Y7eFd6yOsp7JJfJmu4XWnLgzP5rH5fjAfZpVXfo0l7kJBBLWri4a5hWZl5xZRGJRVf6Q0fx65T
jgK0ETVSYn6AOIMS0VGvfqKmPX8RysO6KE2l8H+0Iy3YzhWdddz05gBJxDAULK1eEr/wj2b7vg7S
nQ2EI57aGIsNrMWMD+vy/s4YOpg6dvuwKLaAzTTNrm6X3b4qB719nVt/Lfgf4fKRgDab4fSaJ71S
REK6O3t+Unefa16gF27gDqvACVsrrCTTa7I9ukgzcys9Q0WIVFqIHD9a7JA+Ff2GjafLkkb2pxAf
zn6dvC5jPLq6fF0p/9oEZev/twRb/TweP2aFrcxSA1uIM71OlWk6IgpbCzsIRJJvZlS6ZS+2sNEO
E6WwiffFZKOlvhILoSDDDszhB7xcptKAsuONYN8MX9bvtiZjLf6Um+uf/dKrpJDfUUMGKHOktR7u
KnVBUGU+Q7P5dDbxICF4aflajPTOf2Wcg8QfB2CWYv6soztNizExN7R7pSM+YoA5pZBvk6CkVFkl
1WWdDnI1tyUtSnrvqCoGxFe8kR1CiIlheDGsOQEsxO2mWIxBdjDz8hSrqOHKagTPpMJ9JVXjMl0z
aqBhKCguo6ExJAnkNaOt2idbKnCWvUsZn8HAdGAS2OQmzsfrc7+THZNd69Z4eGLsLQsv/eSrpKs5
Rj8FX+Uo/Rn811s6G1d1ya2Itk/8mh2q7v/rAIQpX7x3aS9hDSGYxwM+MOykMuzIoSpcwcE0YNZ8
245Hxs2NQ3JIUX4w3xZ0jOgW5sTUY/Wu8IrAhSHbpVmZUMx7+dAl5r6/yn+SxYE/L3DYRSaJmhA7
0wME1ax0zPu0X8/BbFLgRIR5Ozzoeo5ZKq6+Kn4/jcacYU18Ifc6cmwI/zucbdOA3/aS62WPxcZB
JrNNWx6OvNG8Ll3fVytRRAaPuoQL/be23xNIRT6movYqXu8r/trYV1og+qx9AITt2AGcOz7HdAV0
hvbktqk8XaJywPxybi5naG1q71kH9WLc+wNgi+fNtdEjUWifalBFeb4PkVHGulN7CTe5SktdWfB1
qEIlrbIhciDoYUjay83Ll4ZmoBQx0pR7C37kBTZSF1u2LlJhcZB4/GhzNp0VMr2ZdFXUDWh3eavw
452W18p41xRcX7/sSq+Qcknw94fCDGS2rL+GzlmFXIdRNg5zjWRjY1cwuiQK8B2WmJXbZr/puFtT
DucY9BOJjN5gN1FrBq6/1kyhWY0CyMIsoLjFabvvnvh8QtydGpbEyPrB5BXfFHaR64i1OYFfBm+d
SjSQcq1mSY4pH9wxj4EM7JFdM6vRLEDS/xstFJw/hHmJnd87sknipnhuHiIWRmLn1nrS9JpCF+s7
gFN5I6A7yEnr+53/KPFjVeoHK9zMZ+pHUzEPXkTsuC7rW/Xv/F7/6UtWAKjAjrn9KNOl7TpXtf4M
HdqxaWEeLn6dSenU76lr+iDX/Vnv4VOe1ooQ5V1e6njr8BGZca2kt/vhG8rNWNE+FuO8Avwjm5EY
WGGe5yjQ/Ap0e4DL2RUrMkvyHjk1OhXnWfzZuhIqxfnR2fS1jK1sJVRQJO0KZWjy9JZWiJ0O1Rvj
ToBxClHidICTUEUAwJOEZr3eCRnyxfXxHNlfrUpU63y43kMDxiPDyazXjR7Y0rEuELj8Xv2ozrJr
m0JeGwiRgSAAXoR6JsHaWOj0O3jxb9l/mCxkl+NuuK9qZLGGOhAi+LcQvPr/AgYV9IJhBv/tYMOV
OVjVs++psAuY4lU+1NnNMtKKjVnTQ4kSe5Yo5SO2dURk0qWLTVjPp9ZBOXX4PBh4NnWpQPFU7AyP
QavXWV1FVVGpRWM/j1JByxLHWAQUVIRH2m+geSFNgtvaFGXe2J5Dw9cQwaJDHQu5w9MFX2wOD+dn
IcUdaPX+JcBbuT5tS27VwpTHDJBUP0IWBtTRjqurgjYh40YVoITaHzRDlVAtbVmF+vkjZ5MGiT+a
I3mlsLpXS9L7H52eNXdy3Vw2WXa4PjsgLjuQkKcM62ZNiOlOf+j7MiX7TEu/gxuqhAcnOFvay5xr
2iGFu/OagiKcWVHV24KWmkwWY/m28uPeLgNjmmtAlxxPtIGBLv/hEOVf9xhm/E+jZflm1Bg7Utw2
xjUu3YwhrRIipzGYu0+gqq/222c7fGJGQ1Wl7cM29MGdX3CU6LgKCaDWBYD02dy7YCHJGY+2fo+9
h1bdhbcoDAWFzDXAS/iEiWfLyftTiPPD7EcCEty2xnfobZ+L7PxWDM9rn7kJVoe6fq4GAE53IRn3
XENBo0kUl2F0bcMWPWtb6l84x9Emm0ENrWh1phyITrGQHplrW4fqcDdSnO7OSw7lxsa5adP+MhAE
UYNIlc247KmuVcF9ZYmrnmVcIa6j095mbQ1NTcj1cUx20sdjNWrElO1eTIGKQZyt3WVqcBZhmxYO
7TifoGVAhJp4z9OlBvoGDbNSfviEPA1sdhKQ5/2LhYlXLddF/KEPXAyH4ag+vOGoSpDI+sJwcR/J
LHJJnoAeklao2ZPDmO4JZqTv3lpuv8LNGiHr1egJnuzrRCRc7WQNFojiQ/YbIXiuXtgF9VOZL1mn
My7MWI16OdwemtmIOi/I61lxW/2gOL/NsrBsofCbhyll3JIMNS0bQg63S07Q/hBBxGWIl7iLSeWQ
KMBaK25urv4P4+2MkUDu4kzffpxC522uuGVhUpakfhEsnInsWuSNc2bhpjnqufI44uQe4icuzqVm
ZXFH12HqWJKIQaq7bcSEjOQcub+q9HbChCUbbRK3WM6k9GpF8/LNeTgJfOW3FGsTlqPjQignWB7m
LMc82P4OQYzc2MEdIJe/HMJfc7dNegKT9J9RmSXtdqBfuS0K5JH3lV7ZeIfJArtpU1ICryTEXgGl
oFvol7oxm1hgsmZ97o6bedas56wxaLYal+uw3FJAYxAijSEPn9/75EQ4wtJomtsxH1Vo2ouI4YRu
XYv7g1cXEY/NwQP0Gws/TBK9QKKBgHwJMocsoQa99THV/NYJpe4APIiYDtKxaiX6PeMu5jdVGzFv
HLNB/2VPhR3jmlFsoMYJEuFkQgB/fInPcNjXW/CxuX4wjJmNfgEuxiJEHDWjzGB/xFoe/P/SPqIm
XcyK62/S1qcElS7GhwRcfqIYCyA6concOkNoWjP5ZNeaRS4jsz3ERhPvDjhSfmgw7xrZBiE+RVum
DnXbFpVViOvH8bgjDXrmqjwxDySvhABr8Cl9qW/Cok637+/YRSwbh9NjlUkzyo3mm69b8PrKgIba
PYMu8IaAq0VoTgyctVtCSUoWgJsBZ7Q6yJljBrCAoycy1YYh4GtG6VAf2mv5bvci6fyc8/uBqJ+9
b5NLJDMlIuPbeA8ZrAtq4e/zpA+TrqoYuHpBk3jApaDQqNA/asAc2S7iJ6onF7J5UoloNtwfRLGM
4LMqbDpVDs6egoRtzFlfymJE5U7hZTUbG3zA08Fmy1vzFjcJkH5ZiRYuOJRtx4ETAxdxYzaKwHQ3
eBOLcj2IWLn3SRuCSS+hVicIrBXhewEyq9u5Efkg/xM5Gb1eptiUK9Esg4uqj6l9QIyI8lKeSEXJ
7zuNCiY87IZ8QWQYzNrQPBtsQKIrpL0cvBi5AoTcECTatqPNVINF/KD35JONrirVtRK7CYA+pudA
dv38dP1/I6BVUio3dSwDlvEP/Zvcw1Q8VYezKBO+nXmAm0O2lSKFo0Q3NWupwZZMxPVTw64kuUHx
JrPAd9ZtH66XV1OO93yq7p4HQgzQ5OSRLOjiI4/L7Cw91iFkTkzqOwoU61yAEOz7Fe7YCBC2vhZo
iJSsa2sc2QL1MZNSq2yPbAiqjsUCyogqdrL7a/kKQ6e6Z2e7/L8liQsrd42gifKE2xlvAqTml6Zn
987wlXo3jmj8ilrhVGAsCT2pzB/OYajrlZ6k7TmUtUo+ZvxlI9U/Djnj5yBZcXXZMF+LtwDqcprz
UebRr5fL4u746tgP3baGnTipwqOsx7O1QZ7GSaMYmUpa/pzEjCRuW1mdLsN7oSe6Wd6xlLb+wpIn
Hrww13banccSqybgEvWU8I7R9N4aacpF9ZGdCswAkzNudrXLWGByAYsYwdM8d/LuZwn8ygVrlyXb
go20RZU8pR65LSBjMPz/JorG5oqklShFWrWM0qZxc3LIi05QgSw5YTipGoLImTiQU/hTXXt86v1v
QAPa4pUCaFvxQ/ubnmE6K7uwdh2N2mwXjrqOS5sHtzzsAzWml1of1UHTZfCKGCsCik15JGfU33lz
GErxrYpul3g9qN7+JiWw4BjqFzOOXbabINdAlK9I1UKQM3EokTsJrxjWVFFbsVIsGZYImUR/q04A
T/P9qWZ2laOZj3HOcWRL00KfVzRItGhCFKb8EVj7XXNiiv94/nMcqcK7DCeefv8DSoXkOaBeYG7f
V5kxpYkR/OKz66u898wMdViEQewdOWPr9yrnvGajKa88p4T5CpCXF+JLVU6ojbt2OUyMvfzVPbHo
LnZisvpe3EHP2uBav70+jnrSPbOoj0vZ/m5v2TMDrimKYtg89lyE6TfA3COzo5YrXihQEDtC5RNj
fOY3A0SndxPyt+EKx6HvZipfNCEaUCt8aGw4WtvkPHDJM8YIKKNzUZW9GKB/FkJqkKqTvjRSv8PQ
YQmcGXkZ3eEVctFrnh9ltBVusGEeNA2vEN8FBAASI++XEyMLcY2DxPatKx2jyQpGWOU6SMUAr3r6
eobC441mF9sMY2kaxlxUYiEA7Llpp25Ne8tuDRytP8TOFunQjarIuA2AbEkDHhlJ3DX213lT/8NR
fyMmFrFmw9qTExYgjnnY88pYw++OhHk78XDRpOq8tpPrsKyZFVpLSCaNN/c8rKpXIrVHbDfGuWMd
2OCCUfjvnlojeb+ByzKOgjzNNLgslVfjlmgBMQOpeACpMXPXhCM2tIFnFfxz1pvLG9PjhhBGP8eD
ytpui5hUfHmukv1EMWK+ZKvqSep4/QEPms9FMDIDXSg0OfA8QVbV/JPzrtWST8+6weAO8EXegg6+
Zf5NGrRFayPgH2mMBsvWS9/uEwjE8k9+YLCyR97wiXGmk5KjVwD2gLEGiYKb+s/yEc160y5AL1eJ
iMeFDmQEHCbCuH4vc0y7fc8mvNnxdD2jtFdnVP67dJHIHyOpmEzFkeFnfZo+oCBNeKYFAEQ4bg0C
2jVgGKHZEo0m0QQqOxocPIJDjd3+QNW+cCT2PPH0HFxCP+ePTC8cJisuj8Qc2AIFmXgNVv6BR+3z
m0ZLmwco8M0nzuCcgPHQWip777R7/r5yIWnJRhuaKSWLHDT8IMGmZQ/Aa3wERX57pauphVQfvyhz
/uDOvMJIAm3UZItaocPV3kZ94mkz5itcH2wyrJj87qxOrWXcTTEO9qP9HPsYO2NgRp4SrlvaK5MR
BLCkP0okPh/3fwhDHe5Pvl2ZLscUZ2mj06nynY5QNvmyBOreeqUZrx/W3tzhRp1PJSTObqzdKhOb
P/pvWSHCghnUpljiunlz0Pn2CQ3WmwJAchqeOOOZ5T90K3u7b6RUoo0nJiBACoSxFnFrCrnxaTlX
Rx1Uljr1srg1DkStz27j+1bFRSX7XUGkQHZbSmHARaSOwDV9uBI6L5MSRdU4LHQWE0+U6E28d5I7
KPnwKOkklZYlyk91bGZ4QMr/gu3gmVydOmRz4xQ7k24qj/np0qyBJgrzJjKVgSBN22dleidbRgDj
vE38LlLIcZYq3eUNLW35/hZs1TPwG1VjlijvAX7Si10StXU6yqkji1q/E9aJvshUnDVNK/DIWZq9
iu0t8wFFzyPgc8tR9bd5hicIY3eVPZuXpxe9eJ1UJLUgGsxcnygzsK549dOW+Rm4gbG4mxZxklJ+
FeBIcmCpvzarbr5Px9/O9jTsug9oqiBOTH/aDFbtdtgPkb4qi4aUe2VcCWXlgLXbLVhx9pVNT+t9
tJUgzR1UWFkEahIOZwJiUkoZydG2GR5ef6E9wVxSXN9zOkHnq06YV+x76ZiCQZ+JiTgceT646jKd
Aw3tJuwIh1ygUlpd7EkaxX33gptoKstH00ykpft4cB5Gv2AEzE8xwAgAuqL3ofxLKLhfD4gHtvxY
7Qx+GwlO7uPqsf4wQBjyzx6o9j0ypv9hC6YJIm+M9PX029G5i927RD8mqlSKJ3+YciE9tyjvKhRE
8asNn4VLq8g6LQgeiRGfK99sbUfrHUUrkidZWI7sAiYuCc4+iG7t02jekoSkjy8fs1Ip6acf7X2j
v6OQa9C7hxfTQGb8tHH2qlhc8QQEz/9KkAjhM0HCipNk381LoGApoEfkYaCr5LSbtgeLhq4CjpzJ
48FxbcGZUwxJp1Hl3vCNBM6TpEAZNppBNC7PUa/5y1M1VBj1TcnyNgvzrXYHyPZ6llQTQoejX517
1wOVnXJWpos6QKRI3Qvj0tJ6dIXbiAp5bz75QL5O7pU7uK9r9foDRmfxVa1Vc1aGYNnS+maPAIJM
8PqahyFZmQYWbyd4NtOWQyNLwy/0NWUthRaB6gsVUcwOunv8QIlwHOG6XbutorP3JkdCEkg4PsKm
W/v4fu6mXJ5hJC5tq7L0xQPlA0TVZUpBG0JBfMYCk885KZy/W3cc6glXVO55hF4/Jf/g2jteYOBV
gpNZrgRrxZHFLhtt76xdfkYhzInnpDcpL3Ak2nqo0RZ6H9R7e15xPnTuxsHV309OQMAek58YLwQ+
XRyTTl2HVzjsTvnUVsynUb3oBkcH4XGUkxFaEvSju8/yFdLVlqAYrGszqsnNlCNyA34oJFCE+aBY
mqCeq2IAya6+jaxH1lr/i1DYR46MF6obAx/V3oDBHnPqx2gmPVEtq6shieS78QnvW5HsLEp1MxSb
VIaCj1kBn+68kvhbK2iHybyNoOKYwpovi1AvGb9ggQeNYM3Z8TtrszaJlZ8W/KnMqpWek9aMQoK+
tkbUECughnzYtby3hFNLgSWLne1DTosF93fHuzY3qEgS3USxAKIKNRJQkaHa4EapxUaE99Q4FExm
lq8hAbehbzU5rwNLaVGGxY52dX1rrBZjAOiTEWmqTOrSrGf+TLPyt6j/nXPpDpdnfoL+GXJSo08t
LHIVaa/Xlt5DVmdGK9IdBJr1Nt5wJpblQ6jeTmrfQZa8of0KQxuh87nuH8msoxLoBtfT827KSoMA
3xNpo0QsKbWcC40i2v8kFkAdWhxtIShkrYx1W5HgI6VWRZAzJxOjT7GIjQhX5y0DcOkxIaV04tuF
ZuySjY56GkaDYatdKRu5/6zNYCNLLZug91Pq5bfOyuStlkCk97qVNI8xzlGms+YRhb/5Hrt6tm/G
utDUuD2mANOBNodEwW9FFP6NtKAaH4qdtc5lNJkMHCFIFEBy9qG8DebD2oVt9QNUH/Dvf/8yd4xR
Se2pqqeJAUEgRcHL9Ys/VPbs+Vzzc17FbwV09cFZuAkMp0GlZ5ZhZb4atLw5t5upyK5LR2BAmyYp
Is8gW9sIMm5VzaWd2KWTJUQiMuFjR06/VO3LmbOZYI9+1coWefyWNmGYbSGMWFQ350hCIwtbHmHh
bm9c+oeTNFi0TrCP+6OZ1Gr0mP8IZBAJLxg9atEPdX46yi86bGU7h3hwvcHWKouB5z/dkBdJ9vET
eQjYm/lnSrrwigUmM/UDYCelH/jWrdJacEDa3JLanYgiLoEWeUELjlmLfZdjADMCbWPmy1uy7mEF
+a0cQOZynr36hLFhmQuyonCn+Pz98obWCWFJ4rmAhASYDIFiQXgrZVahFsM7OuoFxwvMZuB3K4aT
9xNKZhaZ0aUqrYaM6bwqmKc6KaxeaYLp5GgSs52qg915eeKGM46iASVl03CPOUxo4F58HWTC4K4f
rhD3XGNPGf7/IU+cR9Mv1kqlrIrnq9xQuwa0/zilAAcoFlWksJT1gZaoQ2/S5OLanuVe8YRmpt95
Vbw/QwHtrxj8N8eyRw+W09MIUNColk4kQ8NOKWGMaAloYyu9FZmhSQfE6rraQlDPZ4hRewdVmGnT
HJmEVSGW2NeJC808AxSXXiwS+pcbW1GgHUYoBnLo8v1tBdCdlqCq0KfQS5aEN1SCxMEZ7VzDbOHE
t5If7Yd26jMSc2RjppibVLleAnFu3biVdD1GH7NUnEYbOe0Vzq1Bn8Jaw7kxs0/MXLx82sgS8Db5
YAfw/msaXvogbPj0q+RcXzPLRIJr3sP/o0pst8JC8/B1cbxwIJgeXXH4lyOXovgJ27YJL4kwmYjz
jOhq9hswPSYnzov27KiMub9N7RVkj5zHXFlO/kxZFZ9ME/VjqohaBbUAYOnczqg4gv6KVvUxI2oR
XlxF9xgWllWnrFlu2A9JIGEoqCIwUfLEqTO2/Uw+8ZyNBy6Jy8bHDoZQv1dlcBmayyGPXdTcUCaa
xpWj8VsCbIer6NnfjVqNO2lAOJwGbB1GZbZuM/ZZKVwRNfaopiRm9VgmG3kf/qwsc9hnmmq/FD1d
VYBiPXF2NP1tLsRdepVhjrYIY7jN8RZdaCJagrCoEA4781wYTGE8/XfWRaWQh8vYXjFkNtq5I/0n
+d056CgxCVUUB7TDzVj8AX2AvWWLypQYRECUijRVcqw73O1+gfq6SbH9XN6yn+fWq12wrLkLJpFj
UeJpLv50olCh1Vbxb2e3GTHHAjqYdGfEQ3ILT8jTY7NNSdiCi3zVDj4XV0SnfpUVyp0B2wqPcEX4
1BkF/ccHh2/023cQwL30hJWq8hABzYgG/CS3F6e12sgecNNZAVlVjsHFADZ3PhfjqIOs+WLlBYWF
4BtKn2RrOoa2Quv9hHcI2lxHAJ5RpvuNm0s+kcUFyWBnlY6VU0l3l4nXd6uUJBMLbWZFBe09FU/e
uJMkqKzbhW3wIFOfq0E0X/UU+5s6k/KVMv80/hevxWInImQbaUEkYsM9x5J+VJslYxet12MjBLjs
cCt38tbh33yAXGGq5x8G5k+S9Gqq7HAkTIqaXyzptB1JaiHjgS/7M/37R4X1fqSvcKCCFlp/iakC
Kh5rSAQIyRK1TnMBeM3RY1QOoReyva5BIfaAKbOM+FC6jU6fEV5ZsW3mksEzPUzR82nIfujpvBoO
K6NhBUy9j9ZBK+XpGK+Ju7S+KXpnIeoQfDlptJMCIZeTj16TQl4cDneKNgP0vGVyC3g3UwOHoSEA
IkKScGLPoGJVwrQiM2aDsXw6aZGT17EEcpEv2yX75fliExS3QejM1IM1/F2Ngi5xvhGv0y4/8TPR
6QSrtALTt7usHkv3VDzo/TETza5NeJtaqz/R9OK4Pt5CMTdPezvH30kz1xPffQ9ZVGo1Si12Tdfd
UdAoUKX3p3fNUpWUDcGT8KJvSga3eEbq1k1cfeYrh/0JUbJ979MKqhc8Us0ps+bAP3bCWSxkmIzX
dVvyOk7KsF51x5Srt3vLjXv3rZx3D4yCJzRzyWRD6OOQzSJSIjgjy2VBNJ6dOyOQHJc8GcD2tklM
/GPLWWKGVllIHybTDgcqefTMCdS8s6tbewVmLgrV32ZnyFxOqdgQITz6MftQgRQRVUrtSXsiBPUO
j0GIYjrOLhB3X2/eMigZd+SGjERxE2UCiFL+zQYwepB401JnIkU+TbbI95Jb45WQvHoQqeMhonPk
J3O893yioJ6//0vbhKC0jD3HEsbioSS9t7FAwrTAX4FiIvwYUxK8VBHAJ9H2E08HuWabC/MtLeFv
kyBu4O55yKQs45LIyrpxiOcxii3d0xTwNZbGvlKMu0CLz4M/+yiK+bp1VWkWlZORMXt0/xZKC39W
XJEU5XIFo5RQ0xIfsvpFfHr+ni7Axqbz5TbpeZAFBq82kNYvwMIxy6Tl5C/TCq2v06MkjFCQD18F
DS6kEp8ScmBH9Rnwx836gw0jBZW6EbHxOXCokKsjedGJzvcoptIgIFzAUIpakaZNzWu09wPvqqlY
rm7PEa/Yrz7azq6tnNjELZDAN01K4oVDSROKovEvDzX0o1PTf2wdy/cn6AD1DWZc0RHz2tM9DH7y
LBbXZoEtWTjPJHf3n9vjDcVOc2MAhHoNV0ROa/qt0UjBWbrvcKYzeNiIxtrF4MLUxqqUVCakNPbM
sNnib50CW6a2dPh54GyYJ/ShKhf8niVDaSdErO6EUg+1MhHQaieSgLplI9SUpu1wPGaB7jCdcKfc
+SMK5a+E72tvjSzunLa8R15zVESoIxXgcP+826VfQHP4Yu8ZWEazHD7xDqY2nDREQ1X0F4/vss8R
ZoRimfK/0/olVPi4gg0bYaDy9rRU1Udtks9oCOABbm7JGJzwKBItnz3awc64HKBfdFilXvh92KXu
B6ArT9ZG0s8rIpc2RrBGzHUCF6MWTXMNoyCVeytwUenyQ3KW9lOodOEBRgaAiAIcitpxFHU4bdhI
1oYoY4j10840FTTvZ5IECEvkRtXdiqwc6xKAIww3bJBABo1MSCU9exGej/lEI5uKWRduleOBnjQi
X5mBY9ioT1RYvngI9pJ8cL5Bxy6SUMti7f0Q55Uzlty79EdArGCcwXXDyrt+cvl2mG77JczaSsom
NF6w7HPUEQhfxdITRu3QvvWTzhTqd2uguFRP2Fs9ILwtXWbRYdhBKnUXq7sF9C4IVhcdyRTd78K3
T6WZUOXQRVmLwIXJ/PpTSwvRU/ddt+E+JcKiFcVLPuqBaaPl0zTkn76aG5uVqmky+SqdXEsIlb3q
jnB/kW0pj4nkonG6LwHLhsfwTlXQXrfGx1tYWP4/Fw2kM08pVR4YTFve7CEtdArBBndD/b9QamUN
2dHMth1Unce2iRuLHJKHBv9nZ7y1Ww2X9Th4hL+iMziuwYzX84w9bh5KwUPzQkV5WenG9W2N//vY
q3Yl7y65XsN+5dDV1qPoRdpqAHDT3aLfEYhLF9tZwa4rxWwLmQEP0gjk/sIvTbFp0dif2qdZ+u2W
foFAO+9rZQBsoryCewLEx8MP4p5ByENXMRHl4WhwIhk5Z/bIxOIE0YVI0FAE/veXhHud5T2I9Xln
fEJpKZWDPi5Qm4t9+dRj18Stpb9lcjrwvf/rM37MQjdNaOD8qyy4K6U31/27T1j1bYgm1BDZ32N+
Y1I9gF67OMp9zbd33/tmlM9bhw80R7UWDClQxqA/0nAuwAAqL67XzeI5/c8GR+bCvRTw6huVTObP
cNAIppAvDCrGwK0a5g3cMqb6NcIFb4gm3RMJ4A/G49ZVEUhIFyshVnI9K9dpCTLfY5xDK3tsChwc
ogXixEUYb4XJ7rkPm0kfLecTsG2wRXRifPppEhjjMbBT77rDd+uiT7lw3OtR9Z3n9cPwmvDYMUQT
hu6iPJYghV/4iyh5JI3ZJARCTVZggR+6YRCOMH2FXYGV6ykSx66spgo4Nl1ZWSGRJfBgyHyvo0uu
bIRpHQ6dtAN5F1Nf3/yabFIEpR/dgYwrdREDC+6bsfDcdEKDmQY/Z6lFM5MR7Sj+SQ0gyTT0bhW3
Tu9Uoyyvp3mQmQteDtV5HlktcNgjJblgAfSGih6VxK/e83jZadKpiDBQ4dpH3AfC/F3eIbiI+zk0
0xj+qEnofeWwl7C3NIP2L5I5qwu/dJOWYqi22DzbMVHqUx/CozD1bTAmAj32uTyal6m5C0vLx48I
YoWaUkuWxi1Lgi9TP4lnlO8mDdR2zk4cK83ohV6CbWh5gAU/ZnztBW5iPNkNJCUvEqhoUu7zCsBN
HuHVv1SeVnQJvwLgpHAjjjl1A14KQVJvpQTpRM+889xsv1d+yMgZs0gFj581+C3hRG9JS6mLM/+u
uFsP8S/jUyuV6E59uFvDHKJuNokgtMrFfgldpjlCHrhZyCLu5kGIfowe1njvlUoGLDKA/FeGbMnv
N/jAWgW94BnvOXXKwe7EiE1NcX6ctcHCF8hilDa4lrouNZCwuovXROPgmwbh+QuTxbNzL0yJohlx
JwqL8lDellsgTJOH0Z5M3auRCBaawk4/lLtcRhHNBAs3czaRPpOl16P34fUunnaZKJqhzsw3gXff
1iKVCkNG31rmOH0Egq6eu4vFS9gGTnusJatxu+2o/SLOph+11TDWcp99LIWVXtTqxpJKWxJliB6Y
3jcluRKNZZkk5zk7b9bMj6000j6zhg5rpuaUURFMh+zA+7yBupG9erwurvoT7IUceewmmlBM3Otd
/8QgJLeVmjPElB2jYOF7DoHEYkrre4D0s8BlatcZldh41FOkmRGNx2r2zBDq37+aGEv6sB3ed24K
rLP+r4RxBC3T/GaAWlrQNhj7pt8WfIPJPV+y97EyTNfcqjqoSbOvMa8kmOGiMP4HLdMfmFKv8ARh
Gom8n8Z6vW9XhJx5O5H0u+6oZFwSvZTwZZbymemYr8YlTuC3iGhJRDwws+1WsZUPhJujAycZHy4s
8eMcPZdCEEMuAby8IX8NHHDKW02dOil2hJqYNvC8WjRp87mXuPzUuc032d9BbBYFbJaMBMG3VGm4
EsPWANwcLeXLKWlO2OfNHs6Jl3M490r5s+Tr+90ARetX7dGtGkwydEzWSo8MNW5wbdIMRvbtw6Ev
Y8zthX01DiIOy9yV2HvUPxz3NzW+oazqnXXXjQa8Xj8oyARkExM1ajPhTo+i5svIDfpt0+nQfLep
qfK+SM+FbNGJggyK2Llf3xCT6OX6xwjorXg88jXyfReA7r3NTKHyrA0zmHxoE7TUvf1jH+ym7Slb
j7sSym21mkheWn/OCviUaMi7z92ZSpPE3Yl/KUTueBsLWCMndwFTo1gB6Ms4uOx7KE67/CfXii1m
xGBgEykY7uMSOPPBUmOX8pCJl8Wn+hUMjJRxPzMFoTuQSOKkturpVX6zRV1BsXPROMclA7XaIzdX
BDdurAILJ/GdNecYj/y+WLpacXMQ01uI3KAhuTgTkTMJN5AC1pGppPv/f9OyvmTMorJaQwFRnb1E
rBU+Udo7jVp6XsU5vTnhwL0C1tzO8aJcMs8KBGdDjA7aZoWoU7W9ntDNsEBqjf5puXEGM6Gko23g
VEiX+YxqvME0B5GfuxMFav1fZngVaBcFpJQoI57iI7z4rfQOf56HGeMFtUw/JzQGcYh7UuciyK6H
5ycfy3rG6BG0HtIJI5A8CAoAAx/WYbq5VvdptWlVWkcirY0KL0WNSzSrgqKn7kWRrQ747uph0S0R
8nIqqL6RhTaD/p6waGrJjSu26P6E7eScDOdEsg7rujUFT/rW9tf5226rO666hl4+5tJIf9qlPb49
F0q091rxll+JYseSNEIUZrMq4HmKX6gH1ZL79byeC0kBRT8dzPzhbMb59iek10G8NXrApqt8IjKx
IrzOL/OjSNf9zEjSCzbUdlob/jgkDNERekQ1ve4dV2De4mv+RdDbOUAEwDeMYeWpVnCmcxHViHr+
+om74fe9xssgY2dn7RAbeBN9jMoX2M5Xs9ePPRuK9J/ztaSH8a+UdgET+e0jmqxUpy5J2KRYiqb4
j0U3DkxQ3MXzTQX911d9kX7/RKS6dCWtu4gMAQ1Pj7ovPE6GM9Y0BF3gsTWtUp1Molmkf3kRV1mg
v5m8K7dNZR1u94AVpTmlnehLTDOm/dry68ARCZN3gYvgrGLOv7v/MMiUjCLKn7/7Xp9akt/6OXCh
7v6shFM1VCDxUKQcsttqMlqJeNmfjbzX4Yv/iGPYsSEZizKEGJcozx+0NEE3K/57FTuLjQUbGBQV
9wfZ0qe9/mqEE9Mu28hHUEBZCW4OQaFExikDJ/OvMtGv5VNa50+4GWAuohuaARvhyoXgxSGS5owx
KmFDACNSztUQcvKaTvXGOgcSV88pIiyeXuFYL4Goi2Es4YRe+nvbaKR+uv14jt2B0MpX1mc/AfvG
PujWZCRhz1JVpwGj3WEBMm9euv8wvwLbZGS3dVLfXvEtFCboz7lHsyqz2R2oUd0x5Hi0rio3uxn0
2GUYK27EQl/XVNQJMrF/cMaNQwWI2pbQYZ+t3Cc/oskk53yUzQPOd6oEjwNhLUI9SpNR2ZC+poN5
LUPvcyDFZhnSjJSI0VYzgJepVoXwDdAlMSpbSPLHVHpyCb6Bk6OLJddtZun1dQP6wEkaAUL5ANjj
QhGCEeeZMYIRWBQNjOzvhNJohszR5gBsqD9IdXr9fGB81Huk0TkrSH+RzGNRxYJyiwLVBZzemkau
9b0WAZPUveGZomT14U9CAXxro1qeM9Ir9vlA1/DiLflQxJXMTIFgSRtDP59qJg6/P385NS++IS7t
GW4UlSq3AaJ21VbxoQdie/YA8+RnSXSJxNzD2J3lxSICNXzpo/sSseZ0yX8lBkaq64f1QlwRCqhz
PCKWrTZLdV2uRluHSMsGhI3Q6YqBcP8vreAsjJ3+kXiuh7pjFZVP28nUOOaPP5oGnUX1/OJdbtas
ifYHJ7Kym5X3OfZKnj/EBa2nTaYub1vBJPDywObIr/Do1Kh0oQONER3vZsp6iP0GSllEkzIxsttH
jhQ8lVPdSyDEfj03s1cGX7S+6Setg9ucxO/LdWKul1GTAVDCSOYEOgjeX1pJXJDWIiowskw9q6/P
CvDlQiUdieACUYsKD+ZdyY4Q/i700o6N9p+ZoPyyp3rE7pi+x5hJqJSF5KPYcShPflNd8ZiQse9t
7JkgXrxqa6xbfVTLdTbb43iOzsHj9xPwlT4/+N0isBlSA4RbyEmwKTXuyvx7LyeErZlOaZrvPPQm
zg31aj7EVi45L1z+fihR/St1fz/vGwECt2Yl9apGElsnWd8Q7vfTJO7+PF+npEYDQm6xG9V36dcM
Wt8SgYXwaRRR9oTMu7flrU3DOPkzsxbDbFFpldSqQsjCIvUkg0yMVrCjle2JE8MbdaX8RLe9mHCV
VBovPOI9sMnI0Q4r4UKyROFgHRCkFJAkF/e0i513MPlejl4eoVwGhE/edWP2ivWiAZewWQwjFkUI
y3piCsqrYcf3z78sS1Lzsf5orfbjf/dXywN6e1b0em9agMMX683NjXUTkG+frJL5w5OVUm9GhR6M
6aH5IYrNqyU1hbsdOOl0IGxEHaSLvdNDi2z4a8uIqRDqkphFy9+h7KNsBjJxqtFmNPkYd0WhqOcH
W+LdCwOzea5+gsXjNxYTOasKSgZRCBbztt9VkPZesOrx9mc4EUy4FtM5XSlnbFmvSaaAX0/Vtiba
BoA1Mapp1fxf3iw1MSzYGjMlPvAYMfrEM+c/kU+HiFyruw7b9JHfP6g9SNnDVkiZeNQD58Fhhz30
uGCeqQvZnxyAjFwpikr8+9A1zYrLGrBl3qeHoJLuNXOoayN6vt+WgPV3+z4/yOmJusQBLNCWsgX+
5XENkSaDrvhj0ZNNbND/qPAJBa3Ex2Tyj7ZXu3E4Bgnxr2z4z4P5jxJ2HRtj90k8YCsFGXM5yiRD
koPIlc8ULFchR3T08HI8qNNOlgyfpRAKNRTgquA3Sgc0jazRZoKApSAl6a8lrHpvNa8u0Asvk1qe
Vx+ZonbEbCG/Yrdb/fZ+ZsIPZfYCosz6JYNTyspUnyhBkz7jWMWvqt1Ex8XA5KAr5QrUKcyVZe0J
TePEL5+D0kdTsae3Y0wqTj3jC0uVsYBLRcNeg6dFdv8QwTq10pD6REZjlJhEy6Tarhlit85jkcfi
7agSq7YNcngJk+7+8EG1UE7LkY5Ao8kEKNARvhKOzM4uEwIeWAoWYRdTn46+J37ryTUGIubq9Vp1
o/xz1dVAcr+xnhPw4Gq7ThyWqk9PX6Sys7stP9aMrw31PvVZxd1UX+8HIu0bDKgLZ4JdMwtI0UDh
toKPU5M3Jp7dfJxibFBWiukt+bGyJ0ZTlrYnxbJycFu8bBI51DE3xym0r23Vd1q9RMhC+9IYaYDT
0nTGZaJO0Qa6J32tH12j3Sv8N8Ke/F5qxEk0j+WyD1F2c6W6c7NqC4NHO6BfCk0rn1c/k8iB3nbp
n9QM/4o9gbsPMJ1VuTY77mrCpT6t21Dt5ywngZgYOPjGOe6mNNqyuchbGVeGIpxrHPkHV4jMNww6
7WhShFofLVhz8izqw11nDpv2hE25n02q4U/nySAIt9sHrY3xZSGluihMpiPYHWs9dGdQ1eKl6bQF
+RPxm6N+o48Nv5kxdCZXJRwyAs41KWmgRq3PiCtiLK85HyM4QdS9xKK0FtxNF9AUgRY1DmnV/07C
ifZYfh4Jw2YB8+M74Jzx0Z/S64TtAEQdYSiOWZiqfx4NhBp5HcB3BAJXw7tlg9TYlQmfLsLC66R6
kRwnlkxNJvqvM116u/yfSTKzU5AfNFFhFqCVwPBz8x49TxzOQAwEqE00h+Zj48ZiAZL/ZAPzDH4J
Cotwi/vpS0N7G7WgV1ihPXml+BbUqf6W5jVuDpHAeSpRHqyvNNDsMGqTmMKuN/8sZMEohmnSTiHe
de2iCpSy7ir+n8YNWPGyVIGNPeovRlxKj7fVGp/tMB3L5DkEpDBhebl+Nx6STHLlnmXdFHdD4VW9
9kJ7JCSlypFGykZyjdWHtVd6PRVS0U2LQdnSkiQtV1/DxukiIzUnz/I2Djr0pLFzTveGACW3qu8/
6PvV+g02hX8lgz77dgPJJdM+/V5/qPKPjaLc+F6aZ/3hfkyeBuRDduyIPgsqXltKg/U18+T0P23z
67kymqfbV5MWUSgK34pRdXFdzOOQkK8lrzutodY96HWcz6X2LMUayAoVxj+0KnIoacNnGvZaaeR0
kz1Vlag2il9Kx/8EFrahXOqttGcNY9julhWj4ydneLodfEWXsx+3PVIdSaLLoY2l43wsWg+Ff83i
HiRF4kQ+otJvr26K2mg3afvoXr/XwncjNysIUuUmo3TyOHFaSyE9oluJBSKkdQichElcxQZAa+o+
yA/Z8ayprkTBVesx2xp+/xqR/F9+nFErCT3EYPP99Ixz8rASQ+aNSicXov14amAoMMWmGCeS16/o
cwg2hI31MUTDhUTBy6ParOBR9MWxsvKMHBzCtrwJ5uR9IRFI99ulUEP5j8j1izzJCIstSu/umKGH
3ym7IKSPvuc3ZS+DJz6weHb+lyrYVqo8pbGoPSf8FYX8B4bXHDUX11naGWaHo4TnXFUAc2j3YE92
Nableu+5SqhzRDo/TFsVWX/vyfbVHv8lqMudC1I+db0TdzxyzjwwEykpFFJfWIo8o4FeeNmy+yal
Kd0l3IP8N5UEYB4kpRVJnOJahBjweXj0xAd1x9HUY4hmRoEpWyTZD56wDlR5sdklVEu86nbmGz1E
893VpRN9GZmwjYlQp+0nIi1xCGxqHIxV5yyK0QH3gnDX3i1smIdgboFOUlqmF2D6o18UZU95FbFy
6ETxYkyt9eNdeFTbmVsbeBCncQNrQ0m7f3xDQJBcmEsVj3RwaKWJ2lH17bBhjUwzsuCWZQUrPnCT
0kMSPB/h0iQhtDkxvyJvDY/ioYcWk80zxoVacUHWHLYxBd7wnLWKbLa8Qi40Bbf1jTKMjCXtu8hN
1ULbrZCBt8oTjgc+TxWrFeFp86HLN+kEjuZSAZkouE9ZymjHGNHUAQ8RzZPjIK2sOebvcmcR+/HV
e9nIwJSLv8iOozKfiUImLNaQz+gYGcZdl6P8DLlTmelBmGwrN5qWsMdyqtn0mCSVGp33VFXUTa7k
XGyQ0jUkwcM5BKJ0PdVNL379pRoE6xGW2mRl+m6DByFlvCKvxBjc+QEvzHz7/ASbdwKX7ACqYrli
zInbHQ48qt30ik7PxCxU0NZ7hlHgqcq+xCJdeVnmCpYAan07NeKS73SzXbYT3H3HnjzKjFRXLBfa
m6LRD0OzZw9Aeg02cza98o+KzxJPEfVfK6qX7R/G+HwhVuyIF+hEAiTspthcY1RaLOySkctCiMo+
5sUjDSu2CdYAmsHSo+E5OOjdolHXwoXW+jSleGy0GYMoYG6Gp/gsdKYOdQI43Ogs/fvGhH8n/ZLd
rZt/QrUByi5E7Rs2uqpc0YUGruqQSWSxW2S39LvzqrbXqHFoUYon38wL9WlwiHITHDynr+EvcRRs
VtvwK7o+pi3kxS+sv+5YYaYNojDeqfYDkStU2aPJtJ9ojv7hWTXX3UIi+xycEtpllK+VIy9AdKjv
YbpLZYAu3ww4SczZNfiOdqwSUDaQa/BLKjvzvazkps0dHyEQOBFfUzecpAxro3nZNaNuXI0AwXPy
4x1ANUMM6sPagh6OQDrO11qY3BdKgkZ1x6WoIL5Tqwc8qzE0ayDejCsoJjyv+Vwi1LcKYHSMcqz5
XAKl2yNbNl8uUrbIUBqmnUwAxZaCrnlaCq2sjSXl502z7RwbiR1y8GyKkp/5fyv9HOrrvTN/Ordk
AFQvI3AgnwOI5PsJjojXY9/X4OFQ/3+bYVamZyVsa2HyjNRq32PbBi0zK3uGnQDy5i4GiCqB9Ks+
jtnhQcMH7Z/I1uOU6hEX3nydX0gCqR3zjX8et7MO5LsK0x+K0XSBciegir5ZqWr4ujljehDiVtSJ
RrXkYh4NlmviXHLyv3ftfbopXxB1M92eSmt9chxlJoyd+hnnr2wUFTbXud/tLLhbcZUqhz0hFc79
PFzgPsqeMsIkXmJe6Zea9nEogI4oo0BFvj+qTWDI4WdfhHGwU1PMUrkuTP0SGe1ojuswPk9ClMEy
YOxYl3ClGGFaQyfFxKwV8UYMqTgGwPbfvMlne0KJCxjD4zOqUGJJRRIbzToab6rgNoIYpWs1SfgB
Jj5lRv8g4t1YVxo9hGRHyXT74MitIp/ouhZBx0Fd1iAxkiMWrytJ3ZSkzHteviEnapNc0RTqcEOQ
sRf+886BpP7fVAkXgMl01wphvbFjYXxG2DrC0SpgwyE/9LippSLjz5//Bz/ZExVnUZYBJfoM3ZNX
C+X0q1wnu3QE2q9Qfy835kNAA/RCnUbBrRlWtaRlJdAA8rpHtzjqbjpAG5C60Dvk5NDA/TlxxpDV
STCXt9a7MNGPIAzib131iu7o94XJBERzNnU4SAvl4HN2QzmWIPvKkTZnS5pjk8lXKpPZtj43iAmA
/CI6z33I9QVrjL4Hb0hmUIfzz8atF5PWQ7SQ7GGfmIxzYImT9DrH30/qwgXlo2AWtqWQR64o+3Wk
gqvUWdvaC+slkL/GdTzkCVcQkgzxDRuwThu4oT1Gh3Oy2vbn7OOb2Lxp6AdjIzmYx+coKn5y4iqt
v1vxV3icBDTiq7gMOAgV/XUFR0sSpDs+MvZ7q5kWpLr5ZQ73XT6Fi8YGZ01Fo8kJqXsfmMa2KLs3
m91hNfLZhKq0brzWfRU/n03vh/aw/4FSL+l7SelkXm+0tm5I1k41H+o1ii5DexjiWBt8aXgiNWFZ
ND+K3x5aw8Ycvt15fC2lZwb4oc/wHjrLroaFvTqTDKe4ukmK0+bXy8t5LAaBHt8kr2UItFpBlZki
IGUJwpxuRySxBx12bo4EwK28RfYkVCzOF54QOace1SxXuwr7IehlNdOLo5VYfe/Z06VMfY7mISV8
6UCwozh8q6cHsAekbT4NHNRdinpjCPSySH9mXO6MOkPU1DLsKe6MW3kHxGtgDREklZDGiHq8Yl31
tlVQY/k6Dp36x1AHPFSvGSlCA0XqF8RZhc3uzNieeSmxd+GTtcluK+PRjMF31DThRIYjrdZWyxTz
aNhTCYukjAd0JC8szqlcM+1dnXW3s8xDw71EjTeEAfUaf4m7g3sKLHI7+EGQnePBXfAad9hnY+2h
wXJAiuUYv+uJ6t6J6xl4Ilmt+TBwe0Yajdxcl5L1jA58oyo5T6xrvsgaU0t3XvclBD3ipR6+z5qp
HLJkrRJ5VVztyYcSsa32bwsN13kgb5J0fVTWqFOL29bdrJOikvv1trUaHiVk2DinUBozYYPoEgtn
AxrnSKgykHF9KF9Vqt7ETHT81ek1sDCm3vmee/b+4dRDzlxOT+/+3sM7V5HZlr82Ex/jUom9tKV2
4SIkAx7pWoH/YHLt8XzVnk+QDtYpgUrNY1vBSX/phm9OcG/OTDnPbO+piKbXjL6glsh1tlJRZWMw
ljK3F8Lc5syi/jfjuFsVNvN8PW1/0ozWiJewZEMjXMlZhmtWoyblD2fLv9MxNEPelDsnc+wjbMkg
sGCJd4picWQFMFBkVDyHkGV8sHXhnHGW0FPOSgDBf1HpmPei+w8wD3FCOPK6pC6SGOGETzjLcx0w
82KbL7RkPPgr1UTTFMicfAqwJ2r2MdJRR5BmOXjnXQxMOg7L94Af+pa1k/fQ6rYPPxJ/7mhys2Fs
oBKrqmlLsbugbAGIHu3ESyokMki5LxjBwGoNhP91uXIoT5s99fduT6bAIcIDcxd+CwhwXm8/TKv4
w02pee9ZAVChVP6Cwo7HiX/ATBOSCXasAAHbf63wqSJyUjxD8VFP7bpgRJeclaCATYTtS2xH6HXe
rA53UYM0rN3GerhZY/t53j6WvItKGb9h2mFDD2vvSoq3QIEuHIMmvYbmTssd/XyzmUMKi8vGMpje
t7jsrcV+pnSba4i4mmcZs472e+VBh/JRq3wwHZBfBOAs97jYa+habIwYuJo0TmQUAUVxGmtbVmTL
dLKW0xZfd1nlwWCFb4FPyKSYC+/udI8cRo9DWJhLmqxPXZA3kb7c0vpwq/76iR9Ml9pySGdrz0P0
iDDu7qtUxjvux+UbRF0pFQd9pHUngQAbkg4CaOw+f2486Y77OkZW4vDc/ZHmmSB7RH9MjZClPqY/
+3cjjBs8q95d1epKYoQ6YpIIWSG8mnuPPdZiddXiXaza7fy2+1B+5Eglmtr08uZmzLejiG+wXHGq
ngwgLeVWeueXmq013zmGrDLnZh7ZBt3RxHHk3UGNJsP6TzOZc4xnwt8hVUgxNlO7l9xYXV72lmby
+plbzgJ+e7ca2S1yKbVkpZgbhcJuoFkdfSfKPOmhT0ww9tdluCuea/5K0HcYY5O7MubrystJy0IQ
2FObEUawFB9SjJ4sJLfGwk+1kUsuVaqz8QpMTMBJ4NRpYdRGWuFx6J03ycGsolBlLrNm6q5f/gsv
q1oRvPgoSwVhJqrc0PrJKqGNFR4GTIu8+szxTx08QT2+OFvGwtUO5nFL4ypcEuMyyLVbiQHZ1cqf
QH4MyHbWnHEvvr02++Li1a2MvdtzSyCdikW5in3ZpQv9D8pd0ibDfRhMPuqElAaGwEEzASAGfZf4
RRv2gGxq3JFRgdUPdMYSWmuBgEgRjpoyVZ1XTS0qQfl4usO2Ug1t/CRmuDSPEgw4Yf4vPF0xOOaU
gZWnH33qikZ2Mu2eza831hSkY7BRoljVnVP0IvcsHXIeEMNNgZRDxLRLRUP9W3VEFB5VMDAGXmAi
1NiFyXDpv9EvV+BVH0byj4lOlwKS8b16p7RijL5Ydpk9l2J/cF8OLZWFV8IXwVLbBsRGnLmZZwTc
q3XskB09k53dcEg+ZAQJYPMSg4fEE0INbYXfW+LEsCv+SrOCr//rCtoFdnEnaqWLvscQR8N44ZFs
LIrnbPw999lqQPxfYxKz6UF1vz7naxV/qBi4jfEjVk+yCDHCtUzW9b5zjr3zgw1nL1bpQwIvzlJ0
jEz+wlrTQglydPrUZ/oyEBe+OcUds6XNXaT2vwr2uA9O0FO2bhnW+5jOlF/7zZHHXevJXD2pvs/u
DENejYSo4bb6tL4yPkqyXRSlzgOl63iBrlTXbgH6llnIvSzWQ4KoJsNsdvSXQDgWVbTuuYiH+3mR
QGDZbYRB2mj23PmHrXbMuajtmhiEJNn+GCwzT9DHKIlHc+QjHnHmxxjwAgVigP0Xr0zPQP2mog0r
Ij8fK4lpRA0G35qUEbMfNCqSruqD7AIZklu+06K6KghYOQJurfBMhbOXSJAfu0NHjIKZT+mDpXQh
c1j7kUr84GCoZ7U3qcnPkieVumC/hvakQxo5UFugnrxeYuweEEdzXcR1xNdaYNyWt240PhS9pB07
bsKMQa/JDYwNfOvQePK6yp4QTzIQhBkcn5IlgksFjcaehkL7wXnMudj9jK/+HtxcIop8rw/a5tv1
z2tAc7ZowXbNNi3eRHB8lb04ZCQO+itDDCORi6crjvgVZ0qm622l/RQ6KRCG7LpV4pQ4RiA9i4hc
nN7PKInvPqyk1fYPIxh5ur6P1GGX9I3Ybgb6OH5sPJEUh9hrMua9veRFjirNCvjzKqEVEWrJVXhZ
c7OiV49zYmTEb/z38LqGnj4tD+D9gZhlz3teRrECpm9Zc+ep2apOaCda0SkKpavi/PBuzW/+uq46
uM0p+y0hOKbgSC6njXglMT0un9LyFa83uTPl8bzWbXTzvDStPb9ew3IYyK1QVbc5zwwadgilVHCr
CbdzJzTsxpeu/pHteCFSc3K8TnK61C5CLv1igJrvTv882nIY7OH0b7SoAdX63LKi71JbWZyC2Bt9
YBr6QCNHiOqbtzqyxQwYZ313+roAhHkvEsuLyXzfEFRJjZPUE8X8hPZ8gVR1uflrsNoFtzHdVTBs
Sgq7gzj5iXbpnBPKDTufl3mX9mjJZ0BtkscyyBixGze9f0s0RkIcv8ygWoaJMKNKUhLh+ynNI71X
/f13L/btcv2MTKP9aB/b92O+eMUYhZUAMjcIH5jf+KyjHxXlCnlX5A9SA0Q/QWrFz5yL/oD5+b9e
rsy8oQtPce2jsh2xvonQhon291U70iYdd89+aQSYNtGN9cXZAxma7CU4bneWS2/RyqXDH/vn1fC0
nyyRLCJ9v/rx8sJNcoG2irFDj9Bu7tPHDU0N6BYJhdvPlTxoQTpBPDeAZptgOhxcaZnKlX0pP8oA
ia0StNJR3qVc9FHGwLSVZatRPA7n2SbznowPoLh9B6KLTQZF1QIGwfoQ9y51NFgTPmn6g93cvVqb
CJG3hxpYpo6CLj/m+ODhBO6cBUcSMNDvcHHMl4smw+NRDHVEWkqftfKEcp4qITQUy8KbGbVl4G7a
pjl2HI32Ihf5+l6HO8qpvgY/8aFhZavtphRE3Q2TWgb30H9u/XmlCMfj10O1aJcIAF7E8YS3rcCC
HOLDc6I/b1iSyxlRE5+NRe5wSlZ9vJqgkU0AkODmo3Yt8u8AbApL91mvUm+K/oyOjClNXHypYsnH
lFGlOm2lz/t/X/a6q78/0lsDOmWdCB72rPOQDExvePrHnnRKP5HBH7xDCR86XLFPIkombFZF1Ckc
xhYkyDGkIj8QSBA3K5yOrOdQd5kTVw+ec4jdDK53hxSwrN1JcHE5DO4xx2BbknKyJMu5/eOMT15D
xPaEx8BsN5IntE4Q8ofWmjsOXGSG0ktemUzSqOUv8Czm/dqViEUS7M+vKRNXgEeXrWsu6qqtfcxn
sVjI2BAnyauAK7qK3sOOKtsvs7S6CazQ88Tg+kfrmXNgxMXhbcxfYu5w51ToWpKlmb9QUHS+TbxA
jVcEkiAcupJ/HfMBiJ8sxtJDmDK9YpWU/HC9DYm5CymGMD3T7Xiokp4WeW5VBNKEPIWbhvAuiFEc
nm09k/2oo1yV0ws371A6+NuauUO3Uwkt20zsPas3xtdKmXZDgd19uIhaSMrZRQAccKacarp+h0+H
eWHg0iZW2hdKRxpBZzBhmdKFW5hw/bTqXB7Gl1pN73e26s9p88/9qVLlroGS9p6eqoVpoNzqam9O
Tca3VBm+sX0HjDsdXQpey2FFBDTdpBWp5aINkur20bNBv2YQe30QHEkUP7A54t6PeaA2QQbt//mG
SPsK1OpmRq//IRLOT/b/RD3cL2rN7EwzKvAzDkYfrNoYhwHRLzf1tOxxDsG/QPYOvcnMKkqtmIUd
mTaj0nYViv0HcZ+NKcR7Y1hZzxfS5ZUep/BRbikSRUNnOm0CvWVGvMX197CcfUro2dcF6wSlgIWt
AXTyCIHDca/8JcDCJiHGu0UDfD2hT3rB8ZSY693CiSMBq7kJ/84+4PBBkwxWW4BtJH0euKTBXs8j
O8DMGsZTL5xPLX6iaJrAqLPM3tx6dWREVP+6MGj+8x1lCfSm0w3erUWTDmz2yY6PjQN5vfdEkPbh
1/5HjqXlyRCyiRcv9gIOaSZzR//yGME7DTOplk/mgpIGDUuE9SiaTp+ljnWDySRQudsNm25e9f/+
iw7ejQGNqGdavAR7xdSJ+nnaNl50LHdewPhFcbfZV8ogg3sybEErIG6WPX07LHEs7U+6H4AtHjuO
1bTZmhZV+2KGTtCKIMfkDRebQIyNwcV9G0SAwHDPSp7BSlOaRXE9zKStT86KxrC8MqeHcyy+Kl6D
X8XkEfjL6t5BsWJBnVc2ATdLz4nxQmFJ+rJTCaIklxpKebDITurrnraaRWg2r7CnsB5GkOOdk7EE
EAeKPwquNFl317cGQ7psuzqNV/SIDij7v9H2Uh0MjLCDrRIwcGrmM60ZITJyRg8NugFz0qRxVBCU
F8Bqy7FV6KlM/X1MxJtiSZId4vIViiY5MfOqoCJFFkCPcRP4vQYjI6Ihy9sQdscI3kLEEe7Zo6uz
fNhVnf0QU8k3zaSV0R5CGldTPbmjd+Pjg836RWNnpP2BApEc3LCr/uQQftwtb+q5muvMrQEBieb7
plIJl0GXyJXveX/nStLLJmFqFEr1JTPxJM0ee7w+4Bds0wvFgI51B3Bv2PPoQGWv5xzEgoT8QOPA
bri2WJI1SyCQOXnszZthal3zG1LxIUZ/HLHK3ineqjenk3+dQD0/XHKy/bqg4Hsn7rz9bds9nW4G
yh52AGozi8K8EVpWYbrFC6QuZu4krZu8+VoBruEf5ES+1cbIBJVlwWcwPdN4d/x4453g2WXc8Du/
Fm551v/tGwGjVdxFuHucYWdKogDnKNLWI64rLYzDYaY3ta0Nm0SaX50xdkuUfJdo7d6VAXi13RQR
gjwSgJ+cjAO1nUUfNijVzbNKRb/0sl/R/SiXJYJiZJO0chThhIWUGIob8gBZQckGpGtInnFPnPdH
yjIPKP04vwykMRcJteF6CBysElVBVRmJD3neUxSyU5S7y3KFyXiJHCa8fBzHLfBhTuU3k9Xl1kwR
bKtKvKth+2QbBEFKZzW62MVk57aFmHdnIdNFOW6AR0eC2wwKWdn4KXpJM9MlzvzAgpWABzet0Qsg
Zi2MFLSQjnExuYNBxBWv0qgSJRf74/iZA5QnKJvxZIQT7BstOVFnHQxlRXRuUKMcLh0DVAsBDesb
ErWnA3VC0Qe+mHGZ/0/PGziaVAUB8nhDHd2CDjrKAQqF0LW5u4xvgCAL4knWOmxxOyj3pG8K4MLC
qToflUJ+zhK1Q1UkZ9Jc2Ihe9f+TFvckf5aF6gu3kwvGgzgYhkPIGXsjMG73DoGxkTgNXoyk4/S0
jWogfPOcXy3ZjVcqOp7FmwBjy7W3NecSdccIl4ySkXNfq+pbH1RBhwoiTHWlVHj0+h6tr2a/A08U
HYkRqNQeT3uvbwd8n5t0KooMKg9RMCtv5HFBPl9HptZreiGPZmWfoiCvc+DSL/+IiuuaV9ZKfRDJ
W+AChja1TB00RXtDXDvYountjpvE+YxBEdTKisHFaxX+L7fbZTBNyrqMe+4VFFvmGXaGxiIwMrPz
27qhx697Pc6QA1/d9bhUMYIX4V8xXhfFXI4tLus/eMqY/bXA43eczLJlpQa/sfjE7ZldqUiLcHFj
KzUvnukeMQFea32cMKpCUWTiiaKtgH/bB7gDkFHd3AfPTp/5m5askAxtHT5pD4Eh/ZfGkYACy2Gc
NxNDN4g+hKOZjpp+iHO8qcK6LIhzt9+jEbSgmRtbZxVFGtMc1ECJpEzZTIRMhBbuePqKrHjEtFd2
jx2N5mkQhYWlGRnCIwRM2BNjCVUyCCqn6E/Jq9qLlbhUsTIzUcBzoFdPlpSWDFIyospwpa/rjXus
jzDiOZOFa9yDSxPDlVM3tv4x7CVV874qshL7+EJXFHiRPhsRetHdyotkApxCB9T+7cSMndheI30V
0Oy2ppO2vQRegNKuTSQG4BR52y2R/w//n/wgRq6X4dVF/8yEp62prFmYDzdmzJkKbBd22rI9z8Ai
JyO4d47pZGfnhIhtoGjkS9E/DorbRAownbK628NP7J4krnH6r1lPC1OypRWEGowRs6dnjR6AepnQ
82DFToMyY6lH2vxlBddVSMx1KXJUO5GormoaDTdkSTBGkBfGrHdhikVPuJ/WJL65SCLZpMX6/OUp
hCzkZ88SPqmI3ZpLWjns/NZjYWdAusD+6VqFfwwGxGOY5K09BJH+/SvlFfCz/V81FTd8awhYd6aB
z4OlVpIGWdQkdMPCeLdoyQDy/XwLIrr3zA7pZ37q3wDwbfV+MWEd7IY6Fre0M1Lzo9NSSP4H2zH1
vKAQquB0Armsm1PtONrnb6Pa1edwUcevCcuAPF+3IQ9CD3PrT+1BjNlwM6KDNrih6hjjtvWk2ALY
Et+RM+YgJwCxIbT5ZvWYWSnC4pKFZ4lW4OhPsNVzCGAKZef4Qxtaj54uS2UINJLjoxw3wKXNwBPH
mua3M5aRS+iVtir1eCL/HZrtwmPfa2+qzVWFd1+6cIgifBz/sXH+O+3uXQ+ZLBswDepNI2+qNMqR
zfZWgE51larTUZ4q79KmcSD6ooP3/XOed7PK9z57WtLOWydxXe0+MHyat3zNvTgn521o3ukSB8HD
ry1e12HeMIYL3yVAF/8QxButB6axuCKK/veEb6a8/NhZuZjJqGTv2rFa0WcNJiCH+07dnH62gYw8
TvNiT1cNfI15lORjMvmyvgoAofO5fpvnlwtxLVch1weCz50qOvFwI8LrnMlwAKzHL63k2S7bZWfe
Rmek+kirNReXtPXghMgxuEHjlIE6C1JEQtTtMX0vht67TyWWkpSYd0XtHWe/TLhRxUpIb+uFWhid
3Du3AO7YQvnEg43XKRyZe1EYaIiY3Z3rZt9F5VYpIzK59wpkUT6vxAHLoa9qOtkW3TM2wSQspKfc
sGbFawIYW0w2P0QfRIEHHHmEnLPnCUmtFtBf1PiV3aZlk34WxHn5dub7aDDuHUtJgVpTz7T5IPt+
Kb4FB39g/egMBgZmTVFZHzEkys1QdAPitdjtOQEE6f/5kBL5A25zjPpv14683USEPWkXsUjczA9/
HuzFdNgpZoSEV1sX5Z18sPrpGohjeA7PVOCkYOUTcrE13DPo7kgROWAPS1qiDpsx/r0H3+C52IO0
XkcqlLFGRgxaodwbVX622TzVJEHsgGN2dN69lMzEBkxq/DEji/N2xrqFkg8x8Kc3oRTn7QHqtdSx
tFiExxUNlbZnCC3D3OhcHp4E+qjDty0AliJ+EK7gR6n/R2U3TY00AEW032i+PzR7jL1VPNwTNn5e
OedmB5HVKS0a4iE7o2KTdLGBHsE/yqHofY/Udu88vvWHtQuNat6TUWAjCjaDydS/fWVgbd38vrok
sZLqPrNLYbhJdayFUbk0oBjm4QILRdOXOPUH/vIxvJbWLT8xXdwLjHgeTnjW3W1mRW7KRD5VUVAc
pP0MIaeXuyVesQiJ11xh7PkkIYm1jZRWpPl98pX2SUdmQgT+hRTX3cV1BwHRTEwUB+vpfiiqwEn/
ZkAWOops4xH+CYTq7My5QUfYQtNkTufCO51OT/TYV7O5o74VgRsfMzV9DEJXGnpj5wXpOwdxP2cc
2Q6vqizzgJzeAd/bSNc8YxxO1YhRxyzM9xnTqhoQpCUspiIEu3rxY1Vf0BMNyb2ss6tmX5cCwOPf
t0+C4h4pZYAGwD6iTAKG1rZSLl8bKLLCp1uEPj5RwCPI7RIZT70FuF+PqJkSF+wDdOiKiS88rwfu
gbDY9LW17zel4Y1EdxU1IYUcm77cPLdUEioRISLoG47PMyvVoikmo62prAqi+NDNkTMuNb/ypz9m
XEOuqR774CwM2vqFIKun3vALtUpbQfJa807uOcmY+YbNScsCfxPC9BgSJBTbdVaEjLqha46ZImRx
J3n4FDI64GO3YnblgByXnzzayGhzKu/VVc/M7deYYeHW5WRiAxAVHE2n9vc6iWGT4J1ie+TXyQja
3NidfTKbNjLxLNr0+uW/1WEhceKxPCz8GaEo4FwDFFFOg69PwyauHTYj5nrz79EHN9UgWOAsI85d
078KK2c0Q75NFpSE/ukNaeNUBdAAFekcdcMwEAQLM9uYFQ7M2uvaKAAwhSWMX1mu9e44l8choFJa
BKLpFqfG9hh1ushSey27G6kkAg9QZo0EegaOHy9PBX3mYyFTcDH2S1WvxZ7tzuliDdpybaGVMIfS
CNTKYqtAtj/ZaO/qKB5ZLAP6pU3xPo1aIhF4kV6Z0WomCxFBHGm/B2gpxyPgHcW7wfBvkHUn4YzX
HhEnjz3V9ETf/utEGO64qaUnvOED06RE3AmJU0VKMPeDXDpm2yZDbpgDwCcJUc4wafhyd8gF4KNo
qhKuIwyx1Uhvgzbt05AKtIz30iHxZ/tCOwRN6vW3TEPqjHBkLCZ25hF52+6t3COuQITW6yh2P0+/
jZdwKXjcEp5ehI59YcHlO+Wu52eVmtdTd8vXHS+TnfAXeVksWDgc/oyAodwz1bnFFTlwWNztmu2N
HOmLalLM99uclRi1GRuzj2gTfoyD6aKUxyU45XA2gTOqMutoMep5sN1rmPJmfT4mf79dTg/ftKrA
e/oL41673Jil81F5BCmxwXp4tYSmq73xxxBfFvZbL062rmky1OOwavMlH4AasIcfGcR1hVUfPOzj
85loC7boUuUsaJrzyOHrRGf59A14GzBbTQHS2LVxwTz1bb9bE29nwwOkuEnqpBVC0NXottIO/pqe
2yyjkMdpwCOxqwAC9k0tt9jtCS3RzArdCzNY3uBVYLnUKOsHNSAqf9JE/fLv26WNOGZFJotsjGrf
ozXGqea9N47mBkCKbkO0LMbx519phfG2S7whZ9ZVLdI/KpHZD5ERUx/bY7IWUzcFJ7LPGVbLty3v
ZFxbYXr3sIzYVCyu4JXWDPClSb8pw/Q2zfSsTep2vntQdoKaI6kT9Hya/7YgDewofeZV6sUCt+Qh
8hZn2i/DGr8598R9YmywASNE4A+yBqVFFlH0mATQgBkmsUhknxVgBFuC7WR2Q0c22lGBGwfBwxw5
CccFOCFQiJpPi3BE5a2o+mygvcF/lAG5CTBDBkmk0Tr26szA+AyRuNrCmhU/u29Rb51STzzPQbVQ
7rwwzif5+RfKR0TlmbiGK11qZZoKEcSC0ScHMtu4Ibnv1sfffhKvaTz/OrBDZVrVPcqguE8h4RVo
oH1fXiMg4f0eFD3WoK3psCF3M0r55BHdv2olNYrkheD1j4t4hm3u+Zgi0T6hld2QrNOrV0MbIc+o
jYDGjB+x90XT9sCr5ZqAKraSlbQVub0iBr4UhDEDQBVQm8xy5KhsJ7Bd3kmqIGmY3fnNDo3ykbFt
Pf5+rqOjyvA4xeMT6nvSSm8WdLj0fEJFqWkyTwxSbal2Y2W/XTjd/+WCKroMJaRee+hOMCR2zCs+
OolQddBZHboMPRmmMy1c/FUNDwB9LFgr946a9A1hIPwMfus+OlEA1v7E/sPojr8FAPeIHnR97xKz
ipG/lo4DQe6KkHm3rZ34uTPLrtV3/5HIL85Y/Z+6kAQo1tvU2ScaNEQxEmbzf1yeyg4vlF5UxyCG
noyYzxvp2w2CijQsRzf7XTXuUclfmoVVs133LKNZMTy2weF9BD9oDu679dpXTx/DKL7N4d3YOhCQ
FlXe9zD8q+SYYbMZ2h8cT+/EHIhdvfPPQ3K4ex23AXO1FfNJVITA6xEtnJguw4k6X/UuamOlfzzt
3/K4IKYdmEcHMWtyQp7JnvuvdoN/tB0XFkd42AU4+ix2z4ulNb4WnHNik+jaSLsK52aVSZKbiPZO
m8vE/MGm1ZApnFa0ajHnwy9sAJ5/7fppqpDTpCIm4cKNpER50YKvcKtUHa3yz4r+w5UqfZ6sqtPZ
6WDTTH+C8ry7ckj2XB1H5DlOpi/4gcaPJwmYRSuauC1UL+0bgxVY/C6+hkBpdMVDuX4TWcu8FgMM
FAImLkoUXltBH5AVQGugUFK5SGLatJw18oQVWjRpp35XvPfa8MZuEaq6yF1AzWpud4IVArK1Imhh
kPEXfNq5tUnUEwRrzb4fSrSrFv9Ktp5QcxmdxfpRHD+fgJRHWavoXsPp4cGFIMDgIs6I5BkwQc/R
wopM8kO4aIBKE9aSzVGruuw84qAWT4/hUGjWmZJyuJLb07ve05LibyU/TeVKasqLwMo/fjcTnQ4C
+/azOjEO7/hLti0+DrYMkaoZKEU5vr5eyj865YwbISWcA9wGud9xyANVx4+4OFme5HjeiCWyRU+X
bBoVzeYKcCFJfBriBGIApnyY97xYlc1Wqgh3uE2iGEAiDvY+WBHzFKE/DbK/rNd0KrdhPrerH3ud
jtgm4D2YShOzi4yF3YC/WWDyGXcFem+dm9tSgT4fT27yl6+DJ1ditom2LgF6I0e4OzToN3+z5qbS
wW4+S4tzD3CMzoneVh4NAiDFmKqX9nqfssuGyEGDJhmDYr7WMYyM2Eica6K1dibg4ec76qsjYVQO
v9JKISlOIr5LSfJ2INXoCFm8aWiLyPI9q8NHxQa0+Xh3KrskAaonQnNfWP30Hq20OlfZe2W0xqk2
4/vrG/Ss0ghkvzd/l0Uw5hg9gSazTOctSm6QiH4ERuJveRCbL+2UCcSInwTia/vJvHl0/3NnmiVq
WwLACAxtDUJkiyADpCiNWUjdxgMbhZvM/eLo/BN7wDeQR9pXKnrNQ8UKUV3EZ2zC29eBTVbint7p
ONFW7kGrhEqV1sTzCIe95SXCvJRkTeOH5AokMYYV7aSD3Hpmz2IMp7/1waUqar0pCLODYJKaNe8M
gQQuqTjbH2OnlQP6s+AEaCkVzsxsqs5LFLS0u8VlRhjqguS4XYZ7RlhnEbwELp1H3YK+ZZO4VE6E
gpShtJbee3FPZnNdtSCvGoAPxhn6sZR7gUR846nBMyzG3uMblTGZLszU9X3smQzn4Chh938+W0jp
uvkHMRij4+6zSTRA6eh8fbM08oegiMjrtfsPUkGAbyRCn2Sl7ZzpId3w59/yJberYKXjJGOUtc8W
TwHDWLy/gMqkSythvhPwXPv6/jvSRkievQAqhcHD/9AFeUuSWTnoCXhzSotrR6EAt8s4cs7sEqsM
JJN8iIQSHV/lRWieGLGJiQ5mr1Jgk20vt2dpD7lHW4is7zVVF5eUGVOiBgpaunBtuEx+phMCUivc
/3RZa1YoEBnAlYNw5i3v7nypPiXKWxbA8OqUe4TZjY6CDDafBjuRuMUviZB+Hk0x4TQNSses4l/s
4fdG05mry8QfTnDwMZllIMHtd6nXk+Mnadtyl04DohbfVoAqb/Nq4E7oEllCOTDtMU7bIIEviPg2
/JKgeuh4dyKTuUbFQZNpU3AEAGJNx2u6E3MjMfoYDuGutPZO17Rj9rMeiNJrKon1sqFgkcH99tlC
u7SqSBF6OuD2h6Kci34HHBASWrjA9lIJiNUaZVmFR7esmn/ko4KpS1tid2SgSgJA2RFGMjNMJmZm
zm5nZLNLNHyV06biBeJLrVViL8b8ZAb0AL+0cpolhFJybtsnUfR1y2TsTdzFU/I7OgtyIgv9JINR
r29zwmAoh/Zg+a6nP2rwlcHpr1anXZ/i/gXP/E3zu5rfZCRQhb6jHcZQw+qd26QOVL6ayfgnuO4G
bLtXRGCepRiHxMhs3XZfEQKvCRNt/bo4fbjyq0OfpHYIKPJNb+hWzJJSxZXuCx0d8Gk5iMr31Qo6
DKG50JTjKT+0RqkP2XrA90qcjnpytBIr44lfFJXTGw582BrBoMZ09+Jf52IBack2oRx7nsGPebhC
kvJ3Noay0ohDgM01z6RrpEJkZNgL9C0dgdTBYmbvKQr1i+rS173qFDFdSBSyPuc/ENTgp6D+INuh
kJY5gYvG9ExnxvBbdj89bg0BLhBrUI6zOa1nzlQJZsJGVc3tOZDhOCHyIgs2OEvxhVI7FP0HVk8c
1asChJYow0H04XLw/6Xzp6e92qVnEtUv4I5Yilrww5P5h9R5b1aiVWFEuQuLkoyeMS2DMsCLyjD2
z6h/N1vvqbL9o7Xh6oyqTtH1FBLB6iNHo4RY6a93syeBqwzP6IfnLmEjeJ3flgS82I7Awfgax2Z5
8PSf3mJBB7+oHat4tN+8gVMPnSnZ0gfQxUw5SvdQ0Aov9Fa3sEYO7uJLJWjliMWx0kD67h76Skej
VyGioXp4bsyeRAN8x1kZOerrk2DQkHUAsZ6uqDrLC+cx7oaBQ/0iX6aK7Bru4SldX2RZBxpXLE8O
nmcl+v9rrPkDJsOF8k0VirqhdcFMiCNQobiKlQKGI+lFYIJVqh4NEdAQhSnYSuAOwDHKuQdCKZRo
V6wF6KElMijuCTvL4cQ2pOyKXjWsb0dT6Uztuml+1GYATuzd6MKWXZK/uq80jRX0IAvPLfVk6ZUv
FbkgjF22mYY3jHqvd9n31D89CJTS22REJaoAZY4ycYr38xNOLE0UbIgKQtDy6DpwNR027Y980v8x
4uu6Zo+APyOyvIKwd16jGoJ3Xq8r03IEH0217ENLTANcLDy9/K9A4JtdM5ng1vwu0UDUNwXfpByC
BHaPUNLDqocPgBJBa548QAo0vARx2svan5BB9NOUkehh7viYRL+1OBsbtEfYGGQsytaOu25t+Fcd
bdNr+9AY47LDk+W1Ej1tml6qpRIt5szFy1lb1A77dn0qKQHNVyYdHe1e9NyqfOYm5HkTMcpLq246
W98kgUUAuo2zSo72vKYrEwI96pNyt6kQj8wLJkzxdoPyoSLM1smIFtTt1CGzJohlqIua+JHd/L0f
FbMxjRjTf7s35aaF/RDVKZhWRJT+hFud4tikdySU+cjuvRoFX+gAf7JQUBfdzMZkFh0HAtIwPgll
jcHXK7dEeb26Q9emPnx/HxNzfnDWXn3OlFv0gF/NsOyS+I+qhdrgSCYiGVePZG7v32IPczb2zcjt
4R3akFGRA1hVMYx1TQ2am8NLfnD2+psIx8KX/LoO3uEZOlvWFgYMxqhX8GEmysFSsHTjtPQ5yl12
u8H9bt+cUr7XwCplLHhi/0LeFQG6dEebnkHHQsU2bh8o4iVzz5VPZH9bToJ8KiQqZBzuhsB9ZLMj
VwuM8h+NX2idid3mVJFB+FQTVc+SiscASquMHrzwbh/YC93RXQunWrLoogk1rMa1EuMbHBcbdIKF
MtNaq82cJicCNwFFozBWaInxJZ+ABPX5jV7Dj4a0GLXF1MQS68H9/rUsNTSMgNbEa7wtLftWqTnq
FArVDiwpwRQcBqKnWqMAGc6mhr1ubVSk4DhR6VrNO0yElO65axDSrP+dXLXRIc6t03DR+Ad203Z/
gsOtfbTymvlw6To3IpaZZAHwzRFziYxtT1xi8866eyYV9hYTYYEgm76QrkJJ8vKxzIBoUOmASyu5
WqEp97Nr8cpQvV50SiMTX47qH9bcm+C6X5zK9CdxqcNB9j29x2e1G96q1ClgRiUMAfWT+N5WIpAn
D+/9OMiQAoIy0YiWvvVvFJbTrYX1iKyfYKGH88ZAhA8X8xw5bGN/KesGBNVC+R/ANyVpPlqxSDt0
s95VUvlP3MmRLNmAyPzN710SY4Q88U716BgUwsdsIvJxCZnb77fOxXt+YAHPVf9U23CkRXPPIxZS
28X0fLvDsQxyFk/sGFh3py39kL0dVUQerMub3zkgPjkmnvwgSeyGC9l2l42TbrtAADpXGbbAlQql
JYKverPTMMnYxMp/GfS2u7ecLOfLKXo2h480cIWVyVYyqMfunUkxDcudD23XnWcK/cxZsnbzbqHx
kn/+ZxdGmUfbAcx8DzbClfW30pYrABeiWQokiYrB6ZW4F4eni2oZjX+Qnx4DS5K7ZbLx11+O9JqA
4R7JOytdM47aoJHua9HYIg8QSTzdUDjoDUowVEDpI6ILlGNE0LFvEcphkxVk30cs5oAHwoL+HPbh
VED6luMrxFE1Dr1frDHJDaMhcXHCJBDrKZzGg8LuOvb6WwsmGVNvyMqag1pDOomlZIyDh+huE/Oe
QTdUW/aCO0Q2tB1HKuY8nPMshZ59tAc3mnDvkd4la0eHTEpAn8pJuM0p2Tl/hwjy7YJZ34JeWkSI
vg5UhEJILsP1HLOE5VDxxJLTYmt1MVPzmUckuDHOFYfIgppl2hWwd4WWWmnkiPnQpjGjXmBCDE6x
XC8GRcavzAeSyO1xZmM/sxvY0q/bZN4IT6y7tM69ffxM3z5weSpYi53Esm5BaRsiOcVVJEBhLEKu
T7UTT5kMTzGiUpNv5v66ZL/qpY3k9IoBqYy1P6FO5bK/a1IJ4fzeWGgM9XzvvHRaoZn8O/hPzUwY
j8wFVRy4TWP8N8hPvfCZuaqq3TbUNxFRgnzrTSD3wUpc7eNlJoDQLt4b9HebqHvuwZgs4sOX+CRB
0jmzHC7RvwWGFwd+Vjb4ATU+3das0dAgjwiqQxcX/fH3d77cVYaN6bHJTZa4LAyWR5Xox4caceD4
4LQR6MRLdWFYXgZKFEW3yv0Shiih3eoFA5DUsUxpMbD7VzPDTinorf/o8e6HqUYTxad/UpmSMOAA
wqpuRddS/CTCresexjYXi+s8PMYZ5WCFejIUSL+Zn+HJJqI9TOkaefv9CdVr7cDmEThjqAagyixA
1IbC3wMm04+AkVXZQ0q3tCgmWm4oVt/v6Fhp35XcuXKnjLNHbcly6PHY8Gsiaa/UASsTpMoBN/ik
45do9g+02d7xwafaJp7UQ0InvGWGCDQyZjBLBXEfrIfC9uFgsKz08b/wf+JgeM0haMyGB9NDIUG7
A537Z+GIu8QkjMgg0IIMp265T25jmgcA2FMBXqBMKpQwj5Eac7+12iAZBLm7w0Vrx/jVRAMtOlKz
kNCKxjSt0jpETaKG2nE0tA2WhY9xd2qr5GlwIvafImqydUvwV2+K0zrDehOcucBK+4iTCYYoUML1
SOifiRGaGyOqdt2B3UCKeSBqK+/cE8YU2Xc+UnPXw/pPq3OZ9ocMIUGoFeX0J+92qg2LBX1pPP54
nSoETcvvXc7NzOEfLOPr7tDGXJ9KfXvaGcgfUpSNJO+dCo8MPkAETeoOWAJgLRSRvxLYkKblwLP3
nCXC8gerTJ0cZCTMX9aNMBA/G2Yr/S1UQFzjOR8dlirhLDe664A3nsijy+/IvLNTohjjI57/ZioA
QIcxfqPMqohJsiacDDfvKYxOPZwgl2SLeqmoNcKdrTVJ2dIyZxmPJdp/LOwyNEON4HmPuaWCOh2g
yxk7u4bgTegHsx6mYE3YASD1+ZcQkx+1EeReneUsVP0TbyxhHrVe4ScTBfUjzdUcNoc2MEASkxzQ
pdOz5sDoxaW1x7TD53WpGUl+VmRye/EYhHI4yolfP6v/xaQw0VyXDZlRdcTOuX7dwUmu9cXh+MYh
z/mfN1dSyZPB7PsTVbAU3HH1FagwaTkLWOHhfYWZdmkGm+xVaFRpr88E/2lIS8+ksQaZ3ggtzm0m
6rg3hwLsgTrXUzxQBLNBmxXKcvvtHFUSPZ5oamrxnhN2PPtwh28gtsb6MAkxdGem5gzLaaZUoF1F
SqLIbQP39B3JBo6r6SecEzXqbHqPgKyOs6IDp1iV1C/4Mie5K4Q3S7nUE5I/nvR2elHGwZ/bFsEu
48RgkuCFw/lTl0gxeWLGeGF8R9t3ud8pBR+OQ78ufL/oAd0Z9DpUvG9cw+sHzeHwQMmoixKA9fZu
pvRxe7U/yKxU9j1GAAwmD5j+li4K8EW14qcttzDm8Sk3isHeH7NGqPC6OGiuV8oYHukMhBuk9knj
bMEHxwe6etzeb8cmVSwVfNroQOCj5PteRjlOJ7GkCJ6ROOvQSkSSWaTJ9FBdRFKKAr6EDKh0kW+m
rGXdHMsfcZxvK6abU+I55MEIYmKowpd/ew2/NDt7iO80VMgDvb6ytzp+Mva4Mz+SiFgbx4YBEz6i
KxrfqOxrode5CUkNXcEo/C2+EqdydLaR1Fe6T1TAuRMo0Zxj3hliOwEtptX1urC/lzzA3hEdtddQ
z83VUPaA1grJJWMWCbkv9ZQ525pBA41ZZpNiox1QZB37+XxpkJgVhMQ5crezxsOKM/b+BIB15xAH
Pd0CUEhRYdlMVg01p1ZMt7sRJZDUK6dlj+ycS5Q8MvC8JIC9SkevewgLMiPFklu1YhtGtughVbL7
m2ZXR3Zz1YqTLgAj063STgx4eJDlDMJKUH2QL76ydHDexzzK5OCTPQU7F9tp2YNT0EuK7dpm6nwK
oP6etjPVvrTB8hG1ZW+qGXDUELsXTdEAegwjY0mQ02zq8HRdkT+d3uXWSRaDa+vWzyVwXbCRBfCv
hqugSXLA7/F5PMlPuzjTiVvxl+c7SGeF6da4gfY66IeYP7d0LnFOEpl5/m97cGKfE16Rug46IxG1
/iJxSICnWzFS80IMAPmT+b2jFBHPGTI2dA1IHFqc7t0tttt1pi0H+gHFUcRrUbI2kGL8sTWSI7kU
AkIjcG0NgwNrj/7/ybI9z0svtGpSe86aYYwgYoic5HFLDGQYLKyQZq/D0bRfoyAHPiiE8tyGHTyW
6ksxGvlohfh5lzBspBCaUNlhZ53SatHtAK8DKstcvptNEc4fKeqW9OPAnQtunsadt6N4f/WoYy2s
61ckW/fxmtFlFva2iga4WE7Dm/xYMmuZxfHsuPiugpBUyxIxYkVS08W+vSOYpH7OsMyJEzj3BKqC
9E7WmbrhS/9hWT1nEfPhmvcsn9mIFsiucsVFoX50pt8zL5p0dfYxIdykM11BJvLIkYURv3v6MNLL
ly81oQUB2rkziK9X6sQYg0bjxdNDSu5DwEwmUf51vgHifW06eUkyIktv7IUG4EMrTdGgtsEbCnMg
Fze/j76iAhwlXhsotny/pP/p4jxkH9uRvmmZwv3QIY6kQIVfkIO5hPBvsGetcIIfhDLeOh0Muzu/
OBiyvHn8HJHbZ8FfZ8O4q8k8FAMjl+Old7aYoWncdb4zRUYWe5GufBISchj1ETtgGhuRjb8+8H7V
cgUJdzy4WPW+cRb4zYjZKV+PnSairXm1pV76fH0a4rZ9SZcBcdThtn3xJGdTdlq3tFNOX1zaL+gA
vvdUbJty2fjDfhqlZxYNKpeNIXhZdw42Wr1eAR6+QsNxzDUfyl6hONOFwLSvhRNoBJL91Q936jFj
57JDGsxNJymfXc3+tAKqYIyK1BplrVTKyhG16/a0pkC29Mp3Agb0Vmzw37XZTbj3AY+QzXCaoXNO
q5sMH0x5+KKETTMkGbj7pWwpJw6vuTMckNSe2MR7K+9n9+eKa5WnnqNpWLCQje9f3kN0gOLjczTP
RIcewaMyMNpuFnHueWl+JMLRJ3XT2z33yMvZX8+sLCAbzdX/BG063CgFAXwCa6vq/CUiIHiN+jyi
5Y/srojynwghDeeD0MnOYR8JJKN0BZu1j8ZVOfyZQ1gFaRRHEHAraKQEtLF9rM8qm5D01h1XTGiJ
mWUYZvBZGXamURbNcAL6MdraOYT2kvdt7fqFowcKl+NKEzj3Q/zg8t88AYiynoGika24SOjzCmTd
hrEilsEjFxvwKP2Y45ZsItOqIXTwtLAQ3nPJUIirz+P93kw7ExpihPeTYSvfcBvgSPIUMrVzTKye
oIuPU2cmDbSSSWyFvcEGtIum42HNHfyg15Fpnnnv8D7QZGF7MrKsqR+7ULSKxDbAL3iIy67ZwY+T
A+Xnu3iIr+wXGxqZvjHU5G7wMUrN7c21DXwlYJD8T2UCjRl0+n3rKXsfU50/pTCKM2vM10SL88mm
mPvEBpbEQ1yRYepO0tKb221nviD6xV7arObDgIMhCaFcXLE3UIQ9cOF9XuxcuPIp4frVRd7Tx2yM
xnhb+jpNIMtWpb0Zve3s4rgSn7PN1nvsHsqD1RcF2eT77ITEv+HWS03mRw4Jk9qa04wChUp8RcyX
jTavtu93aaRSN2N7jKbSaLUtgrQTxDTiwFkbZXKHPLihes2sm09TsU6gpRVMnnIK6o+uvjXX6dmK
g86MC01hj8rSjYrd9x6BkAi7LmtxII6e5eZo9wNmx5JvGiWorP46HvQwBfdsWfXV1f0msW4r24LO
aF5vgb9IuXVCFbVCLzZdH06PBUeeQfngVDuAEERmWq9dTPxeDTzy0OzCtoI5GsVFkJltoFu6OqXf
lCUl0vuv1EmKMg3EwJVUKF8gMbqK5Ef3qsqQJ1JLEIeQUv+bS9xQxOjL/FF3TwiJ73gnJTgVeMdM
QYDQjYlykBSjnU05Yo9alttOhN/enPUYsec/CYxC/nal80HHSLkFnv5+YKIu4PIFBzb8J8vrVBM+
RsJ7QodwBQLYS0k3u+NhKEeJs9wcZvpsNqw3GD2o+R/I/R5Wt4BGAvirX5xMf6EXbH5pTkFL3rqH
2bcHMCje7xlmPsrMo295ZAnmHZ2B6KEpyDIusEqDg+2oqX5LU5bzm6B9tUeMsN6ZVT6NtkjnGxr1
Bp7mCnXcYxLyGJIyNVwYONriBu1X6s78mGDBfJt3IKBEZndYu8KP82heA5kMva9fEqgKUKjDQVfW
bKb6HSas6NwdjSxs074MVZOkv+LLPM37csGKYlP7yIFU91zSXvz/aUd0ieYCHQnKLVYglmAL9GjX
nSNgYRecqQbtJBcKJyUbqAjQJH+toPt1dkO6pgwnPlHwcfIr9i3Bs+4r9QfjArcSmWt21W3XCuDf
kka+UZ2EkOhGvqEa70xuUiu/oxfz5vldZ/pOjuvYEJx/lbdn+360OiSD82jfQyNKyYp4p37KTBab
mAgdsJyKAEs7LjbyLIMtH238TJrJifBLaEH4/1DNeWu9rjxLjwxfOi0d9Us9z9fEhn7S9cbXnPRx
dnCCJxwuV+wzTTfUiIQ3uCRGJZxiIuacYwhT6edBiqvUrtTwLnQjK+101okM62meLaEdCWFU9Osj
SNGvVIjExynhrOCDrP1P7CTw3czQf9qZ7RF6f3lIa1hwKQZMDVuNhjkZQIwnevHs4ySvKUm0OnZI
WfmnBNa3iGap2YlHgDLfPxvO4lKgpNvmpNEPrsfhQHxMkNgR96+7WjB8IqwH9BMKYskqPh7jwli/
7ZtD1uRnlMUq2poH6tL5KVLhCerDgZMGmxThHVLd73BQXEi/k4O2onp7XsrBe8TxwTCf65+m0Dbx
/dbcBp3Y12YpsiRRpU7yhenUoYl2sBipfiPQeauMBmZBPbf/sHmiN6IRq05yEtVxowmH1LkbWO4D
g5//QnAHVeHzv8MdRYVNIdGij4bTHMtlFpWe+CLcWfRi3f2v8q/p1I8Ti9MPvXt3H8jg4msnZeUJ
k/WMAFBH/OVsApDKtomD8x5W0wL0iaf8KWSZEH7cCNJt847D8CDY3xP2jmX3L41a5TLeqsoRCoHs
R4EVngqoyjDI2GhWEdygMMowqGUAAQeZvBakAZbfafT0m/Wss7mUvf5eGwI7oxBkzuEIXpsKTY8Z
w6KLRXlpJboMFQ2JEqN+BNquEZxo9UQYGesyh0gpd320uimXaWStSN8Fzdwi3wJcdUwhfgkECyH3
tvx5Fbps28piD7+ovUwjm0WSVNP/5srUOCqgLON6AsPonild5xJK/W8W9qldYQbRfpbkt4lGhZLd
sgxfMe6FnGn82yEXnnTXiZfnCxAHvLG1g82x23LywPp7xO62LyzxI+TQ+lsSY6cGQtawKs+5KsUX
b4kn9RbFm1Y1pSZqXYFaopPX4lYVW3sM9VDxLujQHMBkaektgNUCnwiUOSXnpfeoSydQVASr4NAz
s5pOUYpmuMhZmUnfrUvcRyqqHD0Aj/Nl7ejEA1A+VfS/R8HOYdj5doF8m+Cotz0o3FEdOJBLxKR1
G6ULC2HQMfleMU2D8Svq9ekkMXBjS4x+PMxe3LKUJK73CgK73HSnyY2iQMzV+8a319cCyEY2UPQd
CewlKuo53lyNXwp1wriEF3pb7xly25ejrKVSDoWFMF+rkimW+abIgc75q2mHC3iyHyKsiHrMBDOU
whoywnUrwlSjYU/HxPkGFY0qh+7CF/vWgSTzeLYBc8yrHYWCiYsX9zTbZvpwruaYyZofNYyS9sQB
AgRZjp1NfFUFQE/dGlSt3u/zzHGJ0ij6jmOeF4DvtZwxfwEyuOnFxXX060EuNDOfPTAXxF4Jeta7
s255G7d75ZD/xpkUlbHa0zdZZptVGCFP++lN56pXGMqkzUFqtWD4K3OvT5U6cJuBAIgjAvjUXfGu
+cqlmgOwrh5Gg7+c1NNGWOnK5NPsCAK6z/HvqApQYL9kWv7dbRyjEEZaAFkD5sIsQveagqcwn+k/
iiotv67ruZ3ppctbKsddf2EolFABaXFZ0bv/W21ejcPOvGzAIh8hxSAo4ioM4kXeku3JtQj5OsgB
mS0G/xvqLfOXjDYJ6+1fKaNK5up+QC1zLansQUOvz8+BNJdAb78f3GZNxf1BhIxWy56imLWbJEtB
4mcDVP4bIFTkBlUauHYh8SYudvsU+07IeUUJH+AZEnQqlCW8C1PRNB3upGAQHjQb+pnP9YnYx957
P4kALxKy8jLfRvDTFFUIxjSYrNzohlz5dQXpL1Z+Jf5KUz0b/cOZcQpPBEJ1VaZAi/zLQek5Ft6E
LXiel9BvcGziFO8/VVA6FdhGkdi6BFz0KJDsGCZXjL5pgyxjCYxGkb8MqrjOfevCbkuu/RFmmb2b
R6QGzLKT0hZkjB9Iw5cEr3Vx5EcizfNMoSWoZS5cjL5ZXPDqis2V5EbuO+I/EFMZ5oW7Sv92eyhS
SRNwW3/DwRRXYUD1N30bCXpPy4tJJe9BhgAZE3hPzJ0FrTPuWaf4KSp22cuJngzBmdyMA/dHDwFz
FpvCh6+p4wICf0k58673Z8afa6z6LnIx1buRIQwOaISkEjypLtNkehtd0POpTerWQdA2Aw+Yy/2D
rtLoLh/6VKikq+mFR/10gxngHRT/rT4grhC8cKXVw2E3nbJqQfzATmnm9j3ErBeknUNhNPliGC0O
DViVGthTPhG1z5ou+R6Hw/Y76Dkva4xP/wCd//jbKZhwUqmdHmE6UePRsenu1J2sgCEZ6fWbwwH2
wdfd/gEaHx+940NWpIgu7841RwtdfIjCAV5aJESgyGIUi4846z7cPY6nH2SeELP9X/reU+UHsPGH
T/ZAND+2zMeusVLPOI6B7KU3OK57j0Yce4hD2XYggzzGk9e14sJpkU7b+vkjY0d9GBZCT3PHCEYn
ScH+z09RonfkHdBJ2WuRLojG7QtltP5qvS/WFmnDKRXrAbA2f372qs3V0mikCA5jrmOIoDiBwYQR
SDFkMoeVsf/45V4xfzaQ5ZX8+zqs5fg0PhFb7TPbjCuweZGFZ/+eK5rs7wvFIChIyTBVi5Ir7CpF
M4whX7roTgKJkI1o5bIRETqNbOhZiyhRWLlnN06nU8WU2UD0Voc5UHMB/WmnAJ96lSFp1g+6Tn5/
a9wEz94GSr4NSqujwuPHMHGXTpJjqewq4tx0Sf2RJZVdXwh+ASej+pcux4Uf7xnfW93wE1Rpto4h
GYkLJaol6Qav0smGIoQB8FL3mAT7X+Qg20NJhattLhxiNq5kd8NVtNOPYG8mrWjqMMBGiutjo+bT
zWUX5KEUz7fwO+Genx+407P6vxJLfM5HoyibpHYt3EWzsY0jWpsC/o0AXxlCjA/zwtWKdS2x7ugW
+7NEk0l9Ui5AkeAPZwhHmjdkK7lx2g0zSPJpp3aNzFD9/S0vtVzCpmiZDmh68fFeAhM6veisqMjT
2UVOn70Fel4haNkvLLIZE77ZFwm1ngMbwUtmv7xPjRNxrcPAr1veL2TZhozSZGmeFDQnEqSSxqha
s+HkAIkOd5tA6AiYVp6ZhKV5Ped+T7N1psLAowZ1v7b4N9cf06wFSkejgMIuBUn1O/E5hBZfbdkS
WVNSw/3qk3OnJPiSlA8UWH/Z7dOETd3fURbjbnSQl3KbA+51n778NOyJ6LXWLD6hIc8yUuWUdFpe
Jdo0eiR3KWuIth4/7wjkup7KSSX2D12pQQHelnxR+iWINgybZ04Tnwt/ypX0mFCRJHzivECGKXPO
6rAB0Rh9a3JaN8+08fgdmqtjGPEsI+VnurkMd9MUf8tnI2/v7fvZssDR7OBCkHLyp/p5tWr/KKoF
Pi7OtbJaOIMVQydN9LCxq6VxoQXJT5M/oHIEql6/XTJhi2Mu5jYYNL8MO/OmG4omnikRQoKD+ncM
i3xE5HyQZkTgi/hVrNoHUbU3iBRspIBZDRhKOadePWGPtyzYnP4+BBOP+9HRQIx+M/nagyN6NwqW
I/anQzdonKvWDhMU82gZwP2RtcZJJ4FmR4JCxWOTVFTxMrVtV+eYl2MsxObGHQpRjObtF+0JXXBc
CmxRkO3nx/suL7G9U7xVf3de/G68c3unfLxL1rnF4AH/tY+OdIqKEcqoAJQ5wrvMjrDCobYt2fPa
5tp3BdpKFb+/7+wjPVUi7U1+31lk8ap6xOQkt40Nicl9UrWBzwjtPmYmmgql++G0dmsPez0hAyVC
kctihDnqE3HmoaySS6MJvVzl6kKiWALNksK8TYTXNAjveUK2yhbTDJZRR05UumlZsa3tCfxW+doG
7cXypzm+z+BjbwvwmXsM7EDBy3OI9mXEuOwbzoSzCzakX4LQ1FcQ7dQ59D3PHyxCCC/BWGC6uHwG
DqS3EDQiCWjOxP28VRnqmQ0gJR43qbl1STB+ka7SlAQPdkZ3pG0uME8pyOeVFo+cLD4vfg5LM7GY
eeRYn8/acfq8jLENP1N4TXPZbBRnJ8T6yf2JLyALheaRhgUYtTz7Jme2XElq7pV9Jr7oZ/QUrgFu
zkv7Ahq6Hfm0MTp0F1RfzELV8/57nD22eE1/3/4LEMKlRU7XsAtShFwdey+vL+CN9ZaaXgORh9au
QdruTQo9bRhy2MKDLop8bsAa6DGKdkQ8RnofvcCGe7LxZmsCbm3xg+SOJDQy4sK4T3X8YcOGBhZi
TinHW4/mSf7Rw2/2oYEHnVzt2g5gGAPiBcUkYcQFajopFlC7g0GonRozPR6ZuT2+SbroQYgHKpLy
PX+L7HYJMsWU8GRHAHCH7bAZPCOg++MkRztLgC19hJPaHOe2iZNmvoM2riQssrtEp75ENhD7Jg9C
HJw8AE+D378MT1675thkJ05iVvMH2fb7tFxMvrq9WsUtebEBbQq+4LZ75xo2Hgzspai1ovLphZyS
o+v1HYo0rJhp/0AE/fJZGU7VHXNfieCzidqIB3trt6W0VLUh9MoobxjP1elv5MXXx4u8P8GU5yfs
fbqo4D970S9Ky+lYSNAfm/CzUaRZroIaMWqJuzAXVg6hTExlUJ+xuTfL71rfdCWtJuufkifvqjZi
cVBnOJY3i1jK6Jm1yqnCPk/wvH3l5T4NX+yZowSapg54n+NMUFSOPL6uYmYwGEnIyvjD/XOhJ3Dr
tRK82mWhSiRAGnrQ47roFhd/D8/j87NBgqHgIZq4rLUJ52RgD5JqDz3/6FTz62vp+/CR3cLUUALg
A/DbxAtmGIQBXzSu8T2xOnzHsEFITcGxMcCLzd4jdRGHK1WpwZqt9Q723Y+xkIeBG/ix/Yx9FT9+
UwbAo4II4skzhAaS4KMNDddO/49dwRJN/54xnkRH+HiVDLXDWSi+Lv4I4JGXCtSDB5B+tjokTbip
qK4lJGuk2tw9aeYnxQm/9fCZ5TnRmBjXHu136YrWVrPHu3uWxiGRjKNZFcLM9/ynSsn6iykOCQ4Q
2Dr2RzF+H4fhMighWdTYtK+xOdcwGqoAi6ukDbB6srAw6Exxnnbm+4nvVwN9AkApK/ZR7v8RfIFY
b8JvXTwlVbUG7fSq0nXcT0gzxZNuIPdOj7AqvN8AVGTpS+55yYf8KmwMdveIJk8kGzOt1Jj4uOc0
i5JL7SGsGPWPslckbS72CAZAryL2BUFEO5Op5p7PiDqkOCUtiEL5/vhFteEMolgt4NCLxpyMAW4B
u3LBMO8oOHmZlF0iyEByy//1oUfD9iTM74TKALfkf5AJVuLNlQ6STIT8k3aAjd/tUOkZNnzbHwtx
4w4NEAKxp9ekP+4nFbsxMM62hLM4cPyOWMP1gMt4+QGd8hSG6+Gbn4k+x3nS5nC6HXw23U9HaOsr
ZhaF5dJwudsGnE13NWo4U2XiqPXMPwtGFyojf3k1xxIwPBp2nGX3MJqgLR31p8PR4ubgInIb+7Fd
yzpKRs9D0JyDrks0K3GNWDttpfFvkYB8cv77RtdifKb91jZXiMzn7in9LLqcrVKVKHE2qr6UP91x
1veVPwLFw6Ts3m2CexwZG/ts9ky+g2HWffkfObpsMg0D+B+CQHiCfvMJ2n4JIwnttzdfa6Yi8YCT
ePmRkBXXyC1tCRouMG/+IGeJcPhfihZDwrSQyySVgNviTJpQal5+7gsoTCG0GpnCI/K50MXgmziq
Wt0brV0WBR40oZ7yztBjp5W5C/8swu3L08k+5D25m7R1lWHU04/NuAMZkeV19hP+WHM8E++M69Nf
bPSnW6hhrEMC46+tFjLc53y1KUd7mIy2tn4NOgs2LZk0dqF/HSmBJks1l8tQoE+dwyMKA2BVU6wO
pACiNCrxLzZTogniX7blnIqhz1AWyseOJFWUtwVBQODTWS8NzT9MgzDL7NFWPqo6g5rb03dPFqLu
qyWmSbJpg1zb8WpWQw9/Dw3fmDCIn4PsfJKouKtn+TQTH0YmCZ7hcpjL6s4EwPKOzap5SbPaTJxx
Y7VrcwvAiPOOX/UaUsZJmdypjnLy/SwUic1L+iEDVlyGshEsbHwoZGFImFkkPPvfZC0CSWsccuvg
MiMTed5pD+/UppWys09yrQXsE8+hcO6K4yG5HQk+GtJB3knPlqcKBT3YFe6cTjIii+b7aE+l2tS4
wSbfBAN79dcF0EwnIBfNskUI0kcfsi18V5RkJcJGJ/9Rq1RcnTyszm9fXM/CeorbcDdoesO7KQHz
yigArtHk38GQkN+2T3ZX9wg4VXvSJoZ0HhpqX3xapLu+O03O/2uSgFN+M1FC8M0FWOsSSOCquc9R
X76TN6HKsHtsPYvtm1NgbLiVG98T5lIWsw/7f+TDXBMmSjIXgN7WmDp/OPJ9ng9x/jcDhJ6SAPlK
oxpebUqg462aZNDF+lCn5JVS5qcjejgG/gkYA88TbMJdZNVvw+p837tt2QzdmdX6l6G3iJPbXydV
M+Lhe9dD4kUNMPUe6I/SI3CdnJ9aXkFz7sYHMNMBUytXK75mFn7F4aark6ZvpC5YJOzz7z/rF9nm
AICEfk+7xwoCnSfYdWsqBJmry5RpIdIWV5fBpYNrqa4U01y+d76jgpSDVupGgxJJMAHSvFAMstCl
a3Hn1GJ/yiXNDankulsHzHwPGpTCpIC+VTxL0+cqC+noXZ84KOZf/lo3LSB9UCv1fF15HYjZdDU+
6rnMhDAtxPEOzX6+Him7/cxF1R3SBZwwWIeBV6PGGa6Uqjo5Yn8lrQGP4CQYS7Qb3oiUSJiQJ4I4
qTbvaZ6EkRWfN4BUeg/f6Ipe+1Bg10vw6jGYtTE7BwcoGtFcaacj1R+wQvuhdUZiudL3Y7xegPPm
pi0z2RuMIZL3o2rktkF8MpI0ugeR2kIsORFac4Ki1r+E8plmVglU/HoorogOvd7hyYA1BgLDwAIJ
4lVgastX+MLj6bc0nypLGPaFhL2XTydf0PHQfbi7Y9r4XFfmAt4sYoaik6DgvUFgf+wV/WYiX/6l
aXRKsTtCXTyU2ZsvDRzxdDKlGR8Q/0nJYtdZmNRM8WYgGL34nYD6pDhMJPH0pKRoUj4/wOVxXI+d
jf8TwHD5zpAXblFLoWMu5CpJr3LJAE/y2SwR07iz7GQAyF/ia7egOY46lH0A886TxmWZurZYx3tl
QkURVMQG8UFdq9oWp2Gw8d/aHn+o+S5YjTgGMdmUHadgvoeC8TD464GFSHwoC4N8enVGC6/jG/Fj
V+/oVRni0gxoCNSgs+ki872NcmquTp+JXiYSu9k10tkR82+JaIj/X1hCQWRBbANJm+9rlrBN7P80
Qwcfq6tOb0nmDIMe4aAurXYGaFfQCjJhws0n3DDhoWLjNI9EgVZbpntIlZzqwCSx0rSNO1Pi9VP2
EDi8bWvvFg9KWZIvUxO1BMgLDSzNU08x+uatqkh7VRyu1Dv2cpxJkjgnR7Jh/h01iEZ+jhf8xl6r
TBRdmCUsB3FFoW/Og3WHVSq0F7LxNPiqu3U28ItaYKOlM2pvsWpohfU3EX+MWOpAi7SiZBpdkHeU
I5gr+acshJ2WWa8Me1iC0DRcuf6zqHkjV23SdwQ00D2hqotJGCozLMb6uk7M6/mDeR3GHb3xYILS
pVBbWKvSb5ouJB0oCW7/yKON/uCh7xmOyWKT90irZuisNlRMYRZopJMtPvQq6IUW1zKEasla0Bhq
Q48AkZyFZVhOcPV+wYsBRb0lHYERhbAnoxKIjz2zWPy6Dwm9dsjB9TYG9eMN7KyPRp91FE/TyVO8
XfBjhACD+POUvMB5qdzOnB+mBBRWrg7pB8ghFDcszRHnxFwOabOX3brPr6LEteG9Mayq+ldFj9MO
JoBOqrgWfj75aiFYxm5hKVpjb73MymUdlO4aCvQOk7Ss80Sr3oJ2jQqn8tPYy3Hi6MlX1c2xfzmW
XAF3A8dABMS5rJNtVDMtkPT/dhgjpcbZt41ZBhXqroC89rOThQxmeJB68uuVBhAondSBU/zQKJxb
Frkfzf+hsPKRRQuS6HNWIPoYg0rTxUvL+1CrCv7316nEV1iGHu+HBqutI3sTZcTCx/7INiVflohl
8JFBgxZx0ZQIshB2/uokttRIMbFOiMpFWWHqlK8AHIGpRtJ77cAQ1ii0a0FCmZ/GAh4cUIgU5ttM
AgEHRghL4GcsdLjuuXss9nv5xOP1fHa044HNd7oNeaIpiYIxzLlZZMSRl1e/vo/S/zLDCR4jPFA8
SWhQTh6FYRDC5JKW75mr+KlX+Q03mT4SlHeIB/6MQHPXZpH9uXYlPKT2l4i9b108FxnnE8hSFXLR
tJ79tCrKSB5zM6si1QXsiL6WTl+soMOBBLB5cYAr1VuMYA8MIjFgzyNzQqTzL5QHYBmr6CeYVivK
Cmu982m2lsc4tC3us4E3jR7OVvALTiVudL06j7mu1eglu+UyJ+LBAUd8QZ6NZYrVSHeXunpf2or3
4/Tnj4JF5SM/DHO4fSoSA5YC/mbdc2m+OmOQgguzg7LCr+otST1CseYcvpQTHjTnlH4FVEarEk9s
UrPVLUG2WBVdD6MKrZw4i7tWUEGitbgeVN2AQyaZ0Gqqgxuwj0mU3JNAWkKl7qnrEaQCKhl7qdpJ
expSJe9YvzMKlcNe8PalfvRDRfaHIbxPhhP89Mf4G5IdtfKTFmG4xYe/S+PmUU0kRmxL00Vucty6
2PC4VzGrK3DDBCti3MCDjJLg4116Q6o7pyxTiLZFcqrg9/1EhRD0lWd+DTDsHX98EWujiJqRP15E
TP84h2bPqBS9JTzfJcEIpMrNdWHgFYkfqEUz06XuYjGECBZ51a0e4xe66k+RQlowtCEdv6mGvmNb
7Rm0g2c87iANaZBCGcFShI9NFY0tY6kuvTe4PuUoXyLwISypPJL76crC1hh356DHf8RWImcNbDlL
UV5zJjP/hl0Tr66FvQ3UqzSfwCG+1jXAP0XUm21euZT8uQA2vOeFDHnBXdLqIqI8LPd33sURYT/d
1/uNZB4nGb5LbW5ApIuz9k1hT+ORhMmEahK5+YGkM0DbhjPFDMM3QNvOCOejdL6S9QEhM5Tvi+/X
OjVps1SvwxJ5RG302bA9WLX3bhyKh8aKfN8wz8TKYYVfEut2MUpXrmorXDhIvtOk74fGrK2A5Dte
oaeKK2fF0zspxk7BiVPbL43XX4xOp/zJEpSrji7uytfeAGDVZLPZ/ryCH7aLRF/trOyJP6ijP5ax
s+m3rsio5Kq+CZvWiJdPvilYapfarFROz8XCL588O6yLgweC2JiEDndg7RrN1W50MB8SOXYqvjL8
a2r+uFufidTF0QDfMpne/VtpephuXHogAMG/kRh3uAkXv+jWXlvRVVs0YpzZys8oxWQzIFWTCUeR
B4VIhxRLFsPK3bYCctcdVfHxdW5bb5bxbd7GnwzZpX6AvyCv7JSNxpXM3Jpp9/zaH7tfnf0n7/jL
LqfE5WlqX9z7f4aSrFiBGkAI3Fdz5EKtQBJQRIxTDd6sZOjprXjWxTzMnrarbq7GJkbnj8AVFzNE
FnNu69En+5V4wV0bxdfbnHScylxH0o/JuKZ64YXWUI9+C0YKNiEiO/S469kdudjd71GwF7DVu461
i3mtflpb9SouT+HLYyY1W+7g1fC5EY9cBYEdRVqkelsO77upIDIH8rx4EOM7/Vtjm+BAwx5rmqfK
qBS0G5+hvITHKlYMVmXU3METWWe1Vcnp4nd2kuMMP31jtL3umyYKeTjp/v+5VLsYHrYKY7Yu4VDt
rDYe7iOMSHwmNpK8jVcfTkjd88JHi0s19s2WdInAkWNt3Egth2S+zXL5DbbY3EZ2BaFYT/iPWy+L
pOdRQvz6F2cyce2N39lodpgAF0dKUxM0O8E4U3Y27Ozqy47AeeLS4/q5nC6U5lscCvbictRieunG
Q2iPWGjyuGmwXsSltYQCspCH1Yx0UlGitvrR+DRtmaW4wQdL32w6mz4YCYk/ZrwXJgSUVoG+Fn29
a3/4bADW3c4odq3m95UEkokE36PZWGhKfS5cnFChYu01VZbvid9tx6nPSTe/wRGHcdZ6beR6LDww
oTfAdLGKDwiKrNlrQ3pcL98B9Y+U/uXgAcRlMPCwaluaDwwdSVKXGWKWpKgCb1g+MYSruLKBbgxD
dt8+1NdAyuo5ybfK3XnWFX0zPSJsLAEBsWF/W9TcLwFuXpVR4Zf6Mfvr846Q3Qcd/tfVf0yqRbO/
IMDFu5oS6QCbrYi44PVNrM1oSofOOMVQL1wQMm1PgQhemWAySKIQWLaqGcHMsqg7L0AX4J/NYFzP
NdwPchZtV6yejd4I0sJM+V8DDSEo/6v/ahNAgxqhJSS7ovBo20VjIIUKqV3EcTXhrbRgZ1tCqbHY
RuN5Twl7X/tHalz83qB0+EPEuJwKIV2N62TK6ACW3x4PJ3EDa1m6vlULwj5KynqE68TQVsmYTbcK
UGUCZzAfaw9l7T+Cm0lO9UUZfSinIABDLWpx7BpCFDNq/WYXXE7XHI+fVDR5o0PonHVw45kIHA/B
a7VGcQjb/2IyFFv2g1ELnvTEWjlcCsZojChhy1lrWGdazr8nUJo3pcuBwd7truaMIZbCko7kyRGO
tT7QWkgC+Dgkg0oiJG7iWkr0qf3NvHvtI0YCxCd7gKjCMoyIw1ne1ZycvgLnAlZSkviWBSP1SelV
223jUtH/tsc+IHvy5Fhg0HHMskG9uoTE2UPJBK/PU/dEND2aYocr6xjsFTDqBw0jSYOnnLhASyT5
EjpRd2UbTqeUWLo/PqGJr/ubkB228u/y/EDprunj+k/rael0tjz9tIGk8jAlWlH/SFH5cuE5wFLH
lT/vX3mWlNzDydEH7iXv+zZ7g0hb4nV4BNer4FC83EZLFAdeUaV9vjZ3glHTGegDjbME+jQpUsPb
IK6Kf4MsO2NUFB6x6q4oW96fgNeL5vbl2WDmVaYy15Fti8p0YoWLeMD1tYik20dV5Z3Dh2wL7JA7
HV5YVuHADJb2zyUO2isSiLKNCBj0wTZfzi779aJ+zhc4LSmOpTvxMLaDNX01XpcetdyxPYbMgiSy
E59IdiIC/3cGbrIPTxTSKPSh9Y9FD94QSiNKw8fcX0QqfDdJ1p82i8LnVkXWoOZ1Bz9CatG5O+NQ
b+zUY3wLeG41k+9HTF3CQiZxhDQ1nMWnEtMNys9u/RUZ2WZgrvtJ3okLK1K/Dz6W9a8PEEiZztuY
lafDI9ea6eOFhsDEQhI2OuVskXgd49ihZp3yV4XWxrUcKuQoEe7AHkr0jwjwNH+7VouP1x9f+rMY
DYKxwSpAvLxpIlmnrNFPT6We6VOXcxRVVw4f+mUwLLg/rOux5iJ6NqyO1MTAVnmm2KjWVnwmBP5d
uDZ2V8QZLMhW3eOn/+cyex+NiVF7Hgo9uUYtKdIZbY+ElFEKLwX94c/RSfBNDuyxaXcqdlfp01xH
ua6HyylJ13yYGLcFZzKPw40jFpVAIlL51xKWjQfA6TMrhBKxCL1qYCmQejKmJSzcxaKTbnusoele
pX7CTrvijiVAqApGkN65o4ZHDtGR2HRuLq4nBFJXS98FH/OxMY79a3vHSPpL3fjMBozQqJSBfedu
bonkRdBfPRUoaCollDw0APNrh/cNBYC56pDoQesdjv5Y1basLR4kwFWrVUrccQFpRmit1j3JUSj0
teVFNTi0nwbX81mrmtFVqYkzGetX4AW4pRUKylrLB6EC1fdGKXUH1Ui9slGuQjJnDxZKL6uHRIuv
v2sQmDJG7OYwm6IOmxm+N1hob0bIMWqWaeFJ1/Ch3YnyrI9frq+iyEQK9eN0EAMKgLnbKDTdwX0P
tEIkPtrE5z1nQYQblLwhkrIydRu//fjSN7WmHaA7YUV985BxxT3F+LzndtiANOKls9tC2tvTo5lH
rP3MSo/c6b988hVkrJNN2IVo92hzpaK7uwtPcdLMpyA13PYUCYmklHgsZzALbcQpv81x+f0YyhEQ
S7AxfDdgTsHf1/dIM3rpQPmhUKF+OU4Xj/t0mqeDmLY9Wx3p6XbKpHFcm+PHpBdi+faGsXY4uUWI
rJq9X4Mqig+KPqRnzOiEPFgQlDJOz1wOQJYV3QMvcM/TUpHKcagwy55EFT7aQX2YqrGGCOS62ia7
JTIfFgdaclEMVibo9MOAGgyhdDZa5/qhi1srj04VdEzGbL15PNXwo7Zyo807pnGcvhBuS55Wbuhv
pHoQ4aXE9auZeUTKQ9m0CiTOtardMQyfWDmcsuYfIbCylC9O5iL3ZMj4oWdEVaSxO64DgGk5y5Cv
CdnTEoL8tPICJ5EfobmOg6TjU1sibhPVGuj5TkaeAQFNJ8D04n9bUt2RIY6h6hiq0370M1ebmcvJ
kwyZQniZW9lhq7aTc5Uywib9MturTGzOXtacCJL+eoV8UcFohSpWDl9TLFEuBy0YQIl9IOfhiI4K
r1PcfeZNAayEVEJSbIUKPU7AHyW2g8n6MWYRf43+oFinP4jmjBqvaK6em58SwDl9wj5tMd9H3Jkk
4wgaaTOZaFrtnm4r89/SKFAXplzbpJzeB9Vpv4Z0f0P5f+/A5Wxjp1HJJfWufT058yaEBGVWEkww
GC0zFA4p+Qu/NgYHmtrgU28lS53mp1dRaoCGiy6lLOGQi64XOqiBFnokPu0WcoJ36X7EpyJI+I1W
8PLUkGQaKqG5zRjc0/ULM4eSju+Xw3hsYDgcpQm4RZUvhst9r5oRjntnB46+BrwukIzZMhwc8xwe
Xu2dpfauuaAq4aQArXm7QsxDxnwBOe/kqVolZb4++pxkxJAVcAyvW27vL/fSOcDbUL0WzV41gyle
J1PKLi9/ToCSVtoXEEZI4BUOfWZ7guzilPof4vL2fzBbTqe8gvDIdZL20BsW6TV4PATxfD0dhEoM
F6bmAH2R8Td4Co3w1gQNpkWzrzdJFYOFY+4Qg60reBz+2C3kLwYN8TMBgCvGfzhrV/551jIU0+op
KWPSFVOXPfQq9y6w+KJ6IFYWBt96G63ITFgPrYS0ji/yDSpe0Ru5aHgJWjyUo6BZVJOJE8ih7lU/
AI6RCVzfFVThFbB2lmy5Wspyuc0TkIHqu3v6Pb3y8f7BMR0FsOl2mkUCLmzj2Czax/0Kty4tuGR2
Fb3Ai+jJgiFYzSzaxsTfEfbb0P5A4M7sYhoegl2TP9mjCbR4fRQd+rwBMIrzCApMiMv3i0Bk3pWj
ImG8tjUtSYxNxyyzVKag+CaKenbTgQnTVEp0qG2knDgFVK5Fj80DMn67mdv6QXNXoy3OUuKDhnhH
rjGn6S1/0s3Z1t2JkM6BBvhc/P1JXcB/S74EZ5M9UReaY5rmCCrrZw8EVgH7NBwYiMExPmr602aj
LoD/HNdLopJoYhaLcQeMN0oKk871zOc0ICx0MlQzuULoUadPy7oE60/4mySFt+bh+jizj8lSp6x5
nB1nAqCKgoevSvLvPjoTcN1KBcxCgcQ01cqM618eEeU1k0GWjVHD8TF+d6OBDEIrnkELRLqlb6ma
tMzMUh9V7c/lyShtGBTMGY/Fxp80vImItzIM9kFrypVVdZJelPRWwnO+Uzg8nwzMrUPaqPnjFxXG
nTGmINWB5KI3yNuszbeNUFmdu6vXWim9XLtFGTAZdUQxt8Ue/Ao6X94a/WnpUciBlBUzCRZLu2Xx
bM8C6wffuxKW/tdFwBm7Qa40xenYiDMd1sm9NXPSQR9SMof38oCgCD0s3oTzcF0/QQo8SQaBriyu
t4GMM5Mz04bg2d2UH1q57fbyT3Pkl4VTS+tC8jywZ4WaykXxT6gjOKo/OXKP83UblJyxLlRE0ZPj
SZlDAkY+CJV1Nw7g7eookzBdw5ivw/UtcULG7pUVzKvr0PSbtfebPqQtpBYYnYxzO8WWL6dsdWvN
3r8NvMjLXlFFDex2zBTgzCWM2yYy+XSAa+vxDCBrW/4hH0fZnvyZsK16LOaIx9Cauvayu1rF74Ra
weCs5YxyXJJ1Jp4stvZSON2IdtjrnSibmA3jQKgcVX8Ho416KyrSWiL+WqM05J3BG2zTF6bq5MQN
snGiNmZcIwxLwqcb32DyDvI4pf18kEHP21D8YYTY1/J0rcZcXeXcjA6x1xkfOQ7XCpIbtMzFsS0L
KPdDQtwy0/w31bGENT9KFSypD+hZpxOg/naMTN5IMjHn10kqovQbOFnr7Bku0jzegF42wjcTeQsU
o5J/5J3M6XrHaWg2uGPzzAShoizHX5qrBEkaxakEB4pmHY6BjqbSIikcbfEkvuxgmqR8zxmYBsX9
Dpr7D2dt/OyQ13CmzkJbR6vNLqnXjOKr8dw37mNxlBbSn7yULYsMdqvANGxj/xbuSMt401FB0Qom
OP8SvZxN2NM+8X/3yi1tZvr6GmmO9aIqvum7D1Tjs/PEktzSTSJMxQsd9yFTZIpAdb++L5D84QFE
qoiczaE6RvytBeJlVZ7FtSotPGhCuURv8FRlgCBeVceTyk8W8KxJ4+cD6TA9OW3bd7Y58RUUuOEh
cslZ+D4qhnNUDuvvaxd3/FCyorpySxdRT7mTZSQq245zTsExHneirda0XYuONYISgITurTaYuOeP
+kVra0an6L4GMlVvFge69uBSxIINuTPwL3oGZLUQTfcRki6oZ4PMPq9AAN3PP6MYd3fxIbA72pZe
uR3rBBY5RwbFbibtOpeXe6EbXpnzSZ7ri2otEg/sHu+H5THSi28TEkL4nA5mIWXSsMhNY1w8jDET
0PH7ADxs66i8M8zg5qnsX95O3Vuf65hr/69g1C3IBjuj89G3PE0K6C8OD6G9iP54agglsqBinw9e
mP2AmtOCuDZg0I858plXhiFW/Gb3DJfasAkS4N+YydxjkF6nU5TrCsd1gvNJ7VQxUEDa/cI9IkK5
7GCcuo3xEpMOfgTtPf5APPTtZ6P7u5xGI0oyvLbDeLwcQipcARwdqXjR6LxchaKKWEgVOCgO72Rd
WLuBx6Af+HATypt1lylpNE/eXHKWRRSg/Jp3WmZzaWnvF7XeWPGPUO2dPhxavc/LgKWufx4eApRc
sE5an7j6Hsq3/ZShibmlNsY/0I/4uHnfwpnulxL/9g/jMJyTKiZMvba+xAnqRk9wi8tv0QL0KvNH
Vv4qNU2GmfsHMBKL/AFj5BFKg540BlcHHcUiI8lwOM+G1wTy174kJRoppYl/CWNT01oXlB90BmXr
Nh8OqJOLFBxvauQRKPTlftQd6Q5arKTaJJacMdzm8POfUg0QxifFE2+Ebe+Mn1fI3TPHwSnT2wA3
eqhRyeGo5n8tQau6WMJYO+/tUYHG+wWaIdMXmIqSnPV4PAzXDD2ssjoQEPhbhhHQaOZKkiqjo5If
0iDRDkNV0hM/IaElvdC+qu8sN2SjBlZ9hFDqkbXiLTdR9Jm85sf/q7FPtPt0nh+ByTxC38pGLmMR
NRkeR1OFrv2JAwkuJ6IoeBWtj71JPlSvBxtinoGapKL8xvlrVrQfX2nXOvikCosP/+jRoyabxLkv
whucNdLiZm4pyW6BUv3RtL9HAe7B3r6QS0cl6Q2vR7/GjDvXd4XHvlfYFMZa8OLAK1lHvPRMMHAP
S17c1PrMYbvLHBbduhZBsvT3qL/49rbbfY2w9PIEbvvMAAL9uln0gA4NrGUZqL9SBcTT8/2lj22Z
NEsPp4XbESS4fh8wCTAFtV/iNdtVy5jqapAnlKYG3gNM+l43UWEqKK86izS4lBbfvljXWIL5248M
Ew5v1uUFrKpSvxa1C29JSrCgJdFjNWrOJKTciXcOJAuhizqdM2zmnC3M1oumSTjPVlMQZcm9yjY/
h21vnXTz25fR5fkOKjzK+fGriFNu9MZtc1AjRsVBR3AvwM7jGuOM1xS6UmYrRpqJwhTfFPNdzSsq
NgSGiyZ7wrC+rwEknz0Nf6C1PDc5kP9Ct41wZ/og4TK4HKTMN66Nz5D7X0jpnEMJKzEJEuBO93b1
aIzoJDGre9RarCbhbDU5Gz5n7u/LqHQ/P8bn8sZ9nlc2OS3pt6wQ64CiO22SfW7Ri5EwpyKr3Ael
MNxGXoxX4IHY/IsqWNOdZOgjcfg7ewHOO23y+eaI4Jc5B6ADZZF6d/yl7kjivje0MFcknMGFGApq
uF740oAjT91pRXpgsxS2VHfQl2et1Jq4ckIL2JSeFElW47KHSQVulnGJmpcpMthav6kkAVg3SMdl
PX4rmdpf3YQAuebRc3n6s0c0+TTzIIIAJYpXiRYzhXTw+G6OLcnBIckfsZlDApl1LJ3VOGr9GHIw
FFQ9EXUjRdjnBu+g7H05+ufzgDMOSWmcodX6VTstxA3QSu+qsyOBq/7Qd3UGbTb2RcqJEZ4vHmVb
EcYm5fSOGB8yOr8K6uttrD4Nw+eoENF0Yl0S0vGAWbO3MgMqeuN8Cn1GgVH3Ig+6lwWba+0IX2Ol
dcHpIankiHXvzma4Nk57fJ4OG6NclMiGCHkXkLqWe6z/riR7XtPVxarwoCA+i1JgUuPIEGeXxP/z
pIWSlp2llWZMBQ7VLHAqmCIvjUTjOhfKWWsZk4Xy8sQAtQ/b0uQYDNOcIeX4wl9HJ94bEO36UIjN
RsMMALOATb24mVlpyBfh0vKoV+s7W2axsOYhWZDEH96Oub/YBPkKFqOkaxCrNIMNS+T52Tvi3Z/v
Nq60DDykGjPH/FN6YLZwdcjfnOyqdidMfJAnEwpZ9/dVTL8rp0XciuTb4ybGBzeR7L2xZ6R0mWaM
yl6qggO4N3QmNKVfHfLlFpKxlHx3RN5Tfj9hUR7Wf087HPBI7DDMw7IxAAD4Xf/HOCsJB8a6QG5t
vNckGeXEePYdNwqAoSfgGfsDqBvasP5zOr/AJyCYpGmMnZK9RQWEPb/QFSWySod7+ZhhjzNTla57
JRgt16MklD+r6hLOO+K9mnKbq4zKi8OQKTorVB3QJQCP3OiKw1+n+sb8j0Rw2XmyUUzCeyjyEnas
EdIrjRmthPMR8RutPON8I0YJ/gydqmIj6gSAIl0eJq0keJ5jdc+/mWGPCxGCGJjzpI2rLkagLD4+
BYc0+Ivh1vJ8ca3sE+rjVFrfWGvi2cu0ZTX/SmkZZZQ0NF3LpSrfA2Ku+0S4BxMcCi4B3KPFjYAY
YcBSWLkRnvd53jAq9Ncinj7wYS9K//V8oZHYY8dFoBd5wt/nFggVFxfKSXGmkj++irs7E4NgrlZ1
I/2yvvUA7ae9p6mFwjf78aJZ2wDICVTZJfVfcQ3v/btkSPZ2EqyLRUuwsbeYq9NjtbLLlmyiY6Wh
8ODxoFVzU0V9F8CvhHYJTzqkjU3VuS2/znI65VWCc9AhVP1qJx7ruEj1d6KBl8QmHNRTWKGdm6Yc
IiunHiS+sHgxu86VbyScP5L0oHCoGz8a0Zz8HWINTdg3M/nN6XsfbP1nud+Lbs981pFmyJGf40HW
1+SeejKFH+DuN89o43dJ9luq01icBdOGOlfBHttlVVcB6xnW/3GjKZ0T5YTs0l+RNjOqOlyIiic1
+4YJYu41uyZAuSmn8QHt3zjBS1CiLRuQllY4o2vxpL/alouEPVqzJI8Lyh59Wx9uCANtTySOx3hD
BrzPY2Xkm8IkEjBZPxbsvM2sg3j2+UTuEnToC2U4gRuzIQBDT0FzFuRclfAfjGLELcyTI67+e7hR
NwQ6oTbZsFiHR6sZNWruhNp7eqV7Eo/J2i7KcfEKm0NzF3+3GvylgT6LXV1kD1AdicdzM6k1RqO4
8WBQ5rJS+jBWEca1oFkLbqQnoaXv3WPk2a/u5eFzXkRgbIw+gydqeaHVEwCaNwIJeenrqNB2P5f2
ceITRHFiOzVVGJm70e5FVH/kOh0daNr4OgxrDihONhXRyMQ2Wp7IvF8nkG7RsOO2lIOP/P7xu5Gr
+7aTeONp0uFn21SgxY0zWA/mOCaz+e3tmsjWNNQcXbDtPLfBww4rd7ba49EyrHN+/3zhFA7HO+Ug
W2unBjYLpTanTk8YYc+s6bzbP82ooQKVajzFRA9UjY6+4PY7qiZljGSz10mfH04jypis883i7KNG
a+9T9KhkrvrtikJmcnucbYpYlL4ZHCUk99vKnwk9/98BLjcsWuifyIczAsYJ6SBK/XogSv0Pj2Ww
q7bqEp9qPCAHU4jk8ccoMGGBP1hZkNUK+wPauNUxs5xOlLlO9jrO93JzED9Wuv2gVOLOxaWDPq6j
gLXQL4GjAWSYvtiP+vusK9XWZxYjm4F1np+5qI282fSzYt19Tcw1zkho9/TT82oOHdZfdZq9SO9h
cC9eM5ZzY9BslrZA3Qvho6FavRNQc5z5un+gjB79BdmNKOPyTyf3/zTKAJQVV4xr8G+gSJlGVvd5
4ac2HFmE2mekr59t8pxH1B4kyJYjMYPNmbouIRgu+5hyKsyhQIuvU8/8aSf2oYlkVYuI/xy/MD1h
AAwzdJQ3JXfcUZittBqQMMEtNIi2ZPhZC4Poy1pu6L8HYapcHSxQyzh8KP6A9Ufg622V+0VHNhQE
l4ufNYJZmZBh0xbjWurBF0nlCaD8pIgIWMrZut97Z/K1pO/x5naQrEuoveTKxjaHmUDZ4UG5mL6n
ibC091hOGaV9vVk6rCAAqQjIaZisbk44xSxZ+tr+J/MbDQcjkLB5XBODpPDpjiR9Ivc2+RF8thME
0M+vkWod9gwKsGhGWcoAM2kIrPmhImeKp5z2jZ4IvdGeueYnWwPctqlbBjjt0+yT1SIb45xe+SOz
sltKwH1hej03Sb8wiDtDSO+GRdOfex47jgTqAXmQlcwmhjFkeiBghrCfK15sn1bGmdfFoedhRrko
9XzFpZ1uGk8bwUD8GufRhvuFgTQt7xhaZ7+1+CnBMFvogunlZtygyeXiYOp7ZwDHn6nAZg3ZTHun
6cQynxhvBMCVGjd0t0euYdxnANJ9mIWItnzQ3rhZI+xuisggRZ4hREGWH2Qa4XmPVyCTzYgbRFas
hEGywLojSlsrkB3WAVhoBCHbXKSbFz0xLMuYS66M8XunM9GBU4wFZDWAikIXE9SaBdFT60R3JgRo
OSR98wE+0AuMLAkdp+cxYXSIAuW4N1Hhd8jhFpnY4o/uWA4T6eZC7t+SE0aFxTQ9eTsypvJnlVlI
7PPKiWm8glQOiDHVnuX3DSuAFhmtg2+yeu6S56f8RuvEF78KGpKg7RFr4bri6HgO2HnyYEzEO0Mx
uuKwpgS1IKXQbc2e4rz2tlNa59Gm1SAdTA8dJVlFSr+N1rTpLeRMVOduNKc/ca07yxTlFYC+fR0Q
4lkZtM/fslrHyDkhdBlGLWyOs4NcnsX+77s7IyqAFx2zfRZAeV4GxVXr/JJ4yTh+WkxnSZaN6n3L
lBqk8yLef5+ae78PwdBSIBPChlpzeAHpNsBnn7aPxLM1kAo+/JRULSB89kY3EExnW08ZRxZji5IU
2vou/olMZ/cpHEDXqqmeZsinzKcS4rGJcTvQ/6qnW8dsbrPILHo7KZmcCuLKfIm3n1DkvNTvgFvj
UKrxaBx3tNQ6m7957aoh+YRXD+8JWHQNq+nM60w9ZA9r3oXXgquoONTK2RQ5WWWnLihg6qQub7hr
SJo789rgUH+n/hF5sDBRDXWONrul9xlLuunTZoZOw8+uAU2q2Tj5mutsrh9fnpmpilGrdjTDvIqU
ugNqwhLHDKJej/IZixveDdH8JUruerbjF8FMiJLz4PozX2Vu3jpWMOfI79xpuLYmcLjDNcvQvHtb
zLUtKqUzp7BW1yVLRLiMO58E50EBw21WzGURYhxGjAJveSBJ2YxDQb89+FyUs9qaFGnO/AtaKuoY
MfKOpXcH9BBj5ike8GwkNgInpTzIRqyKogCvQpWjQBfZLbyxQEj8Jfyb0tLMpJ+5gCMSq+nVkkEB
bEICAGijpkOTrGoifAR18r6zUmwv0b41BSYxIiMIY/Cc/mn64uGf6g+nS8UYoIq1dpwI3Cd0oslF
r1dDxYlx00e8YccZ4LGsQObtbWi1ERac5LOoJ7/ni4QxdTpaBZaPU/hUntOfNvavRl1pBez+Z9KY
l3APDG/ZG1zjCkLLDcy3uYFGzIqkZ3CSQ2/Xl4dLChAKg/ngtR+mXAqSjRM3IfXQ4ZG7iTurJPWd
tENOXIAY64t8jwZTO1osXrR5FcaaTn+fsJXLpNARDaiFsBM/SqQX7drzzyJyVg4nAHPJVsuslETj
fPcq8Bewkg5Tgx5O3efPE9lfu2Y1mT5hHKfIKtNSE+gIbP59kGhgd9wP5sFjk3JldDD2GIA8BxIg
DLiSKjLHHTJPJdveeEGXN3L0EmCWKblXkk52yUfbLtcoepbXLiExRN0doKZsOFdH9xB9xWa6nK5b
jBo5c/QUt6e9zsIB2Zs25g5GOd5PpXPM2g1G56nU8tcFlzPeAy+DLjXcffiwhmSBQDBV2gsC+NI7
/fA+H6LR3yTR/AgXQgbFkKZY4/oUB1s+GO6mNnAqYWrQQuZb4gMzd8SIfgItUlO3f5f3h/kioSRF
lpKTWjFPYuBy4KIy24DKBFYgKP9DkcgPTzFf8UdlLf1vHeeVOQ4Qd/6aLUmKLk+ckcorm71cE+zQ
b7rowfAF0r4ZzQgricEJHlGM/MWIhwBzpe7UGiGFBU8mAaI/8RJmCsgLSgCL/I0gjWmFpn2QyPMO
QaiOfcruJHQFgyrjpbq6CZ0kj1JO3sldddBjloQnDM82f0ikSQwivQ86f056R+HBBV9o7cL3Hjj7
8JEhUsMCtKgZ8CQFc5SYZ2DwyT63hbDPQuXSSrWe/OjWtOWmhBzHb8qfEeRBJNi115zUtVztSsfY
7miH5KKFA1kIEWm2bP+MvGzRFh+guqHdACbovQV8Z+X4nxp9/2Q/vgIo8OIZwUbxQd4AgYa2vBTj
TE8DD4I45bEtxj8f2rl5N6iFYjlfQTJ+i0sqtrWZmbmBU+FRV7iJrtmC4W1nwIdkHSBCSqtbA5mI
jyRNOmbkIRQpYNCJbNzmdg697zLtbCSaZ1mC2AtNjFRqwffGiNTIOZvrss82q1NdTEDBdaIi4cdG
Z0iUqcRfMuLgx2yl3bObLpu5Y7ss3lQgjFM/n6KsYq6xwRTfQprYuyOrbNi5jCCjJaMSGrtOQ+k+
xIAVi6Rtk9edA05RxVYnoVM9FurL6TULsJwrWJYbPNOTS5OapmdDInBdGmEQ+GZ/iBdY482gKeRu
UMePwypu8OIGRl31fzyDHzaMLi1i7Npb1xcFlnvmNNEKQrSf+6QgK3YHIEYQrHVJ0p+jHrV6e61M
tADNCjBF9SiIfiYoBB/wKdYnpn0vgp4cEC7Q0JqDkB3GssSX6ZLWBIpiZun5EaFPySoAJRrNamVE
ERQ3tssFAe7IG1OLUzlERi1S7qfjQneSmltxCC8DxyJwb5WgCOSf1Djv+xRZi1ARlVn+2eSA5nX4
yS4VwILu+3U/Q1iGmojvoRYoT9IT+USUWU1dLq/v1XerL4ddmCZm/UqASUtydkDMOrnKOM93VY0C
mzKdlKiZS80dqCjBNXEaSm3IBZyCQe9Iw/Ge139qoEx2NzjkZw39pGIOCNq+rBSUyARMFX4awahz
T/1YgMcitl+wvVMye5ibQLfToD9Gm+9bBI9q66glF4LYFGXBKzjxCjIs9E6y9MYsY7194Mbffgtb
1csqi9DXp/gsJVM6V7qQ5xfFDDG1agNso5xN3mcgQ1WGbN2yXi8p9fH7PZnsKwrKOxyeS3VOsH2k
VQ0wpawpRidpwQtTIRierugYyiiH8CBJKHf1UPqdpx5Mwnk/g/CorfuvpeiM4uDJfXIsTpmATFZc
TFpEU1IYF0xIhOsQhvcgaOPeR1O2AYI16yO6hYtRdvGzqX3TcFU38dsc+utPVfBlCU3fSFEagl99
xK2A8+jIkNRARiTD7jtWrmVo3nA8fsRag1sJN3Qrbg2Q5CSEAd/ia1g0w3TpYcTDqVcii2gl+ORb
FnBRw9eL+hai+nrITGdO6EXSOfJKZoLBr2KsfON5SPEPYjKadYqF2nMa/AxZMriXZbcmXhbI+y9I
qRH2TB6pKX8X0GrpMJSp6ejFXvRTobEAYaK/3XuOPDmTXacnrIXTktebGAdKbPr1RHN9jZ5iR3x+
yCBR2KMc+lq3sDYp3YHguR7GfHdZLildf3Zp3FBIfdRZu3sYGj9fuq+51/pQm8z6MzNy1U49cBGy
+BNfZ7kkhNv/18r19wxzmMPBv3v13tES4LGbdTkMlTiZ+OGllhsXYZ4bg7RM66N3z3SWPzt88UPh
dHjaTKTXntW3xciIMKlY3lbZzW2D0CUWyuMUl+sh7QkNbSyiQTmCujFVrwi521AktKazwpa4jotE
buvfcHcmPAvwIeCSLSvo9yoVQx2+H7Yw5EMWC6UjobfsENifnmuCQKUpA/T7MIcPKJubewWfgo/I
dUGYE+rSVznrN6cz/GnW0ud8k/4zljIOv3WXLWHydVc+esMt+RIgdb8Y/NXVIFLISu+zdYJni9Yp
JuNqRwiLIjatA+2+wmJyOzJlOePvTkct88b4Z8vk8XYKiTEzKPPPddgZLSWiyV1QM8XvmhmgDK32
/ephvPNWeMQlDbkW+9BtY/iBToQJvgHb0+yIKcMlQl8g0ctXpHzrAYS379A+pbAvh+cAuV9DHeTI
OUJ+vLOqRqs+X6DvStEt7WrabdglynHa0nTEtxxPHg9WPXm+/mY2aL27/6BwtWM99enb6oowwqDd
aCrLL4sh7PsLQTe/pU/QxtpQi/BtGtYuaOT8/1MLRPhaG0eauRo3QNKSm6EJbNeEuOyEK725HO6m
C+5wppGia9cbmsqBWi20AohssZ6fjPdupKRu5aEkyzUSuhx5WSzq2FCvfklJXobsIdmY1e3ZGANz
78CZH/eVJnnSlMM6AKIyp7zcJ0GJNtaCJe5iMrRkAmdfbTv7HyUc4x4N3qtvQGYK8fqUUjvjBXl5
gOeS1ORv/sHCHsPqazrSWV03ZrsKnvollnLGgcN+52apC8qsaPTHCGPGvI1qFTVi8B6ynAFPsuX9
jVpoXJ/TnB+h3BV6WYYPqhPjPgP/JyR0RIhoSfpo16piNvQjzMPuRDc0/cyz6v3gerIztwJhqMAa
HUkz/lwpUlj40UMcdMaRGXZKeH8o1BlUV7j8JPTAxHDdJbAgKycIzNetYahhlVt9w7vcmXALYJfX
OWhBae6d+THP/cpK4uiWwwdM0RyYrbdzl80HgOHx9UnoUgnCnmLH/5x5l501gE690Tp2bg9+7kBP
9cDZ7mx4WQLL+2E9tvDFYr8ahfUladg7/n/0sK+FElrIkPpCUT/uOLaYVozTHYqVfogwn7GP/s6e
7LuZnKY0xcV+lff1P7YaJq+/3AycJZNPRdIKNF+TOGUkz4V8TJZtwwEyCglOZIlKCMJAMYL006nF
vHtfvujLjjtnWYFFybnjeUa0zQXL+OhgEz1DR+svlqB0zXC51C6CiLsZbnmq2HD7B+PTdP6RHlFF
pUDv8aSPSZzZKoaJwk6AFMZnq6AjknzHaRpv1fV5gfocUclNCfq/3UHmhl4FTDMVLtRrZr/ld5wA
Wm+FFVubCmPDCMphhDWXAcSCQycNGA/UEOpfjXQh51hUB3uPF7FIcXzd/HhJ/F/jHeGjaRLYUVui
5d+npIX3HjROTlEVTkDUChGUGWid1W0dbWlu+b7s9hMmrkElrnuXTM9ne4MZKPN59fQvMx9+s/Ft
dmNHGYaVXz3SQU7cOqcp5sr/uKZ8zS3f6BOvvAzjxp7uObbzyWvZr2PLBdbXyTgY7o5Exh5V5pFo
j5EcLnSWzWGAi+Cueb4R/wUnmKACDBbw7uJNJIaEXj8tU3RTx5OhW9Iq5pnIvb3Z5Do2b+4h2RHi
0Q23UjrQ2vHo6BlnlwrNj6wniaw2Fo4C/64P47M1+xHnTFrIKhIaqAM+/rd3Ajsr9tywTxz2aWsh
LI2DH29FZL6dHrL7yj4rfGR/f1Iyfyje25MymjmEm7nQBK9O8I7WfvKyS9re8TdUtkGQxrOGF20E
cdMdX6smUm51RjyILjRg8nuddHzYKaFbEMLM11bxPowfFd9k8KO8zDSmZCE848N6/PK7o6SQvMl5
lSEorNit8ze9PPTvR72+KOKVdG3mEM4h7zYrVv2uGT18DDR5b9dkaUT0gvfdR/sqiJ8HMvKK853e
e/+l1iOJweiK6BIPmVHxyuaDsp0KGwiwCNiOXsmo46fi7mIyzbzN3xoVPS6cRQtOxDdTnSl09mrg
PYhZtgWXYJlN1sOvbmUlpLQhhWDMWwX08KHfJuIXXj4ftnFlc4s54FexEYe5FmnGTEnp3RBEVmEF
apEcXvO+Np4sp+CrMZve03NoAWb2D+GLbdoCMGC3MAdOqcy5fD/T5b10uDURHJCrXy+CvooIiM6F
xumEOot50lvxZAJsY+N4a6uKmkD46F1LLiPP5KPfCd19wGABRdfsg//mmvvo4WvPJ3sOSnqnDf44
7Z2rfo1wW9EC4/phb0d5ZRtA0RkuPTNapTsOHxLU+IlpG5ya3dWy0gLrdgvt1Vb3+sipBOhEygMp
PNUf7YxYKTHYzR6h8Z/kZiZ3mKu8Zp58VVGJ22h/6rh0GX2wUDVYeMTasMcP0uShE1IyVMdB3J95
fDCSk0IQPa9ucU2OCovgKxb7g1+2NOqkesembMH18hNJEuyUI+XLZG7cvubePV5rDVQz+voKCQwf
McF4jMzvIG7rShq+gtoNfdpatxhyPCck6K44Ea+7aQ60b3QMecBcUvFJFTni/aO2glhEt2zbfMfg
2bLMJSZgDWOQ7TeqoDhgJCNTRSSzvFf+SJjAbyshVFsojNdsCN1UzDngVDSyJKDWpoXRSLfH+mWM
XZz/9lKPMm6sO+jM+kynQqw0wMizdClLDf+uwpHtp6+FIOU481LchW0e4BJj5iIDWND35faIbUoJ
865fy3H2W2oIPlGXSfrifWiVLoq9dXrErhM8zhbqodjTTJS4pWJocQECa9uafBdAS190tUQ3AgQY
XSu4/U2/PQkzb8OgQAvWC+WEKpT+pv2xNgemjF/4o9E4KZURdVH3FUEXNCP7w3rU8jHzs1YA6TLF
72akxWwTygPdh7jTLeYZN5TBjVGHh86OypHq9HekL7rCfgujwumke1w3WYmhUe6QgeR8P1vWQ8x9
aXkX2pVsWRb5P8LKRfuoI0SKyt5alZ/EQrhbc5L6av8Za6676xYqk8UnvALdzTeCgZi/LgkPoXk0
UyY2Ft9mg9GbTBbq+djUPpoNBymUsuDfHj9P7DA7L6WJZzraHhJR8MVthNcXKGqCEbxlR+x0x8U+
SQagnFwji5RhI4tXFeQasb+nicbB/y1aKQdPvxUQQ3eOzAzQJKU3IPMbWXn2cZry72wos5K9YgSu
kxqQfdRIRJ+IWkjBzUZSji1cg9BQIua8CFEfCfC+fbGZZSe1xxXDUeEJyKefEkm1Kp1CG3dYam1E
A9a3KEqHGr6vuaNipRhAsD8JbPot/4llOzfPW8L8YedZWJUi1LMbhl7yjnOu4Pm7Y5g30FHBeoSC
rTWugx6ie2YNWLL9RQKLs0qqaD1zx2GMYNjsAXfOAqhFwIUEvBRJB0HaazwCQZ65WAKAjR/dlEop
wdnskprn1/5TjJYszKr8NE7qHCcF71smx/va1OW93iuNWnRnrfkz6cPFuliSRluP1Sq5PFU+10Y5
bDSWRjDwFm0sjKwDfxhYUDHTQ7mZxLRhcLmyOn2YKSGh+fAIIAZQiF1qbyXl9yLGHJlVczc+EVo4
XZ8sISSmMdZdtDkDcD2uGpInWvbwJG0IxoIyQcIdTVoCEuFCFB8i+xu/nyPIrLNhnxbiLX4vJuIW
7UXRXMB1VcjNLJPHxT/nzaJLQaaDxK66Lr5uSa3XeRNw2t9cMCsvFlNew8HlQe23Gi0W7HLN60TD
u1pMsmGwb1l8gz7DzozZLMtQ1HPIiRaj72vCZJHK0ErZH4JwVAqmCEvhIw6lAlrIQVynb/eKinSu
CnSwJzOG66JHYpDBPSkk+MdeZfJjNLjw26aHEhKAizegUaqbpvy3pOZY0Xw/0lrOdylLtzmVqKRf
pRRs7CwsfaXjjKzslsVIuYaqNfbnXAO2kntjqXI38dzkw6a+4wDLlilPCrjcOZFzPeBPNFb8RHcB
24SaI/5ITUN9LSJ73GhwCj4EqqvNuhDDuvo3R0GuclLAeRPJLd3x93vzencER7uWnFuq9qYXlmYK
uHlSvUb1WZ2Qgp3ezlRzhHJd4qG7uxiTd4X5lwK/5x8qQOmHJ2eNSf2VCV9lQu+SHcefN8YR++2K
vCU4wfoP585IL0A48Nha9e1gVYo2NpU27riPh+DGrqSsnMrb8NpTmXBx16yixz6H22t9DqOQyBzz
bYvfV3xYpAA3bo7BqOVp+UQ6XxO07vpDewIBF/jRbkCyuTr2ogwqW1BJLvOP3T0ikot3E+DKPTQa
Y3rA4eBSXPl1pYAABIyrbbHasjbCPeJQUQgR7WrAJDpsZQjbviM6F+ZJyusyNbVgbScZxJedV4DZ
PylRAld0f+CfuuOc11VYvRyZj4uXxBPd3F5AnFUC5qV8p26bs6hySApy/LLHptLUSsuGwuINTpKH
6Y08ry2t3DyllXioVy0g1pDFcVjNSuhB1ITTBxcdcl4b9Mq8r9JyjNfdwjKcpDGmxLbfvvg12ddH
A+kZIxu10anRbN3aWED+UrCH4CM1sxSDoGUtQH5ubGFcUQiUaXcV/rXV+mnprXOfc6QryPq39rhN
UIc8sMynL3LqeblsbEdwusQBa5OT4hSRSE/LSPw4u0PWG1D4rveYcSqpetSNZ+wcR7XvCicTeyv/
ng0TJo6YC9Nk1lYPyvxD3Ep/22+l3JENtCbcGtHLF6PVlKDZYJxBquFfnte6S8x76TntbsRVRvuZ
qZmbdvYmek/qRXYatpIbFT/ZAdooIQapgBcixX+MsHEc6xW4eZTtMcgiIjpAgqD5B2uYKrkGmVty
ziFBggsYkln+2dh0vSCSCtueMOCRJ8P77Gs5NPUFQX/y+QM2RksnlWDHB5pSIbhNsSaI5YbLuyWh
TKsoy35b2CtuoiKQKqoMS74qzQWSVh8bJkRysGFnLleHBGkeaLUD2cp3+NVq1WRvZA7DcUm+V90r
6viOefii0UICFLI2KV2ovZAIfgsF0dhfAY7CbN3YmWrgaH/Fls2kH8kLEGGHToUw231Sizo2rD13
Fzo+iCIAaz9fgVP4Xauvv6+O7rzC3uOQXw+Zn2+YHWuck64Mya8WYwfVffA/5X5mITn2nuuuqXx6
1Y0A9FGfy0j9NxGkqiWjtTJf2ZFYKu6PueMEA/TZWvw3qCRyRZl7yXzMV/eSVE8Yo+1ExevU8x05
TcsXD53Ph4puQoWjSXPsEkVI4IQQrOkIDzZ5v3YzgWR8VtKPGbxVfpsCGDZIOlwH+RIjI2LlnVGq
35XX4OscNDtjQG6NE8OL4aF4ZCNKL3vLIpwQWY8wi5blPTdWr4oUyMoD6GFUYzsOSBPkQywQ6B5x
kdUuwl2Eyynu5alx1m+lKAH7y1lowigNYuOOQ9b1dwYFIex3tfrIVWX2DsvTePmkmQZ4s+Lwwle1
/wuGE17tOSGGFUXHDr7gOFcF4d4Gk0AaRQLouZDFAFWzPYVUMKr8cOdtAhgj3N2xI5qMMU2rKT+A
K9nEGQSLMobP6m/KW9mAAyC2DAK+zkQPjBRSmgfGVSH47H7jET/CgeZgUfh8ztIbRPOuzCMSg9bU
sS7WMm2yHVv/Np+OyAxHFkzpsskaU4M57+LleG0QDNeFyPxq9RFLOvN80hOJDQQQWdRI1EYj/Grv
morBtU1pw7dYAvwbtT9M8wufLGW/vxLOfLxwOEeFrAF4cmoBLAMuldJCO7BAC0AWei6ta2+Dl/GH
ek7Qlp1T67N2o2j8f5wOp2r/qzfROUFsztD2sp0/IchpQ4h0eeqdGt5lL8iLZGuEwyE+oYbp6z8Q
iHfnU0kU+ZPVNKYWiSlIn75KUbUFzynr+3jVHWrGpdNs/ygrZJx0W8VnZLgqlNP2zu6zxoPZwe+i
y3VzKxVEMXO2mVyKPuLkbbLweLqoCX+Md1v7HmLnE8gmTxLvh8XA7Vd4O8kNihl7+AikkcDqwk1G
mEn8nNl36lsvdb+HwS5Q9pjj0VN0fTEkBy8p/oRagwVGoZJ1u6U0rMdYdC6+Sz39GgK0eVz5MN9j
hW6SyWbJdj0oMCdYkuof7SxmYHzi9RF8BG7CEsUKXVec+0KQv5R32ZiXSh1FpRLOL5Jw7VwGE8Nr
ZWKxuo1OVIUhIApm8bVahtopqd0bZG/ZDFwG8fPOPIjNmdqb+xeNxbqgxwvu1CaU0WH4BA3MpqEm
nYXYLHOlq0tVZsRrVm0/aZ/OnK2uvi1sB8s01NCKUAgWbecxSMj/VOikW9Plyq1Pod8fNjHslr09
7Lg7oM1LyObUsYXg/OhcATCw/1ohfz3B99t+peN6iRI+Q89Ovn2gYNGuwvGiX0vJlDP90FnzeV9G
lMOwyqcjVBkQe5YyrxaJxwiT2JKyeXeAKtRzuUxvYt08h2dkD7UiGx8tRA5vJ0pqLfUswAQcSCGp
CnEuL5HKHgoN5KyiM0FKYd+D/q4kZMdmmtQbqjoAWUlU1at4S7Cnoq+FbMWbbwHZac3e6GyCQJbS
WqFWQLykiGJKj9nQotTcRIMcZErFkEo+oeMYVpmV8TDsZJ1lZB9oz9r22g9kDV/5XZesZL5OT599
EUVeAc+GgW/ES941csKoFzEx9mLrKgNdhlxCw+rvkL/xqEU6Sr2vcIwOLjEpMjzwWG95fldCA5nT
18OHqTHl0Lbx/53qXb8X2awgjX0DWoRa8zDWv3KxIWiVQC5qs5Rc5DKI20lJjHKVMoZt3VrdLh6t
J7qgpyHS+hYIhrVx4Ucf43GOhX73itNR/Atco4lKITT1WtZ7yhS1Xk604e8MDjtc89Nm90nUbxD4
DUByDiuSeqlWp9YZJ9k+7iRqoRbGfdKIZP4ajDUDtj9sj5W1Z4eW/DYwWdLsb35HZdlhnPNZi8ge
7lqY1dQvH1XnJYGZ5VyUyVc1sCHaXRR4IaR1MjBLBQbwlc9n0zwXp2zwCRo+opbZX/wYyMX+cMyK
auEnWVkEwy7jdy9wY7ga1Qyb1qeYDcSC+ZfYP6/vtIfG+q3cxLr3JPPzI3Wk+v2ZND5ZG7gWqbTb
S+yqRagFQAe6EzHbGjEPYfE06QZXV5+nd1+rWoHJ9UMR5gHClEyFgPC3P4DYTP655LiXLRcHkvNt
lIIIHBuLZL1h72/1qS+roPc5YSMYDG50TfmF9YfkOljXHnVIyBQjRoXmpn65KcAYfJF90hrXxuyI
nVoLXwk0G14NXVAqe+hC2OcV6uqCWx/qV27YNerzWpKEauDJBmDlvbvjw++fAqlF4D8G1IsSUNUu
/3PfoTnOrzzEoRqpNgfYWIFHlMSows+6N/zhYz9Se1dILs0Tpf3sgIwkrdRpwYUq15OYJ7NysfG9
6pHP/71BtHMFdvg17DxZwUnpT1KxDF6TPSWmBmUiiPuelKYLN4mquI261NmuJKwHvEqXm7HpnViu
VlkfAcYrs8YE3/xyTqGskvS/TZQ4k/nL4QwmIlqDoQOTOwQWSNB4wSw6YZSUlcr0Af+O0u51F5WU
kqBAlv9UG5bhn1mYdP2rq9XuSEcj3+HDj8hrXb3jjRbNTSG2LQQUECy7xcorQ0IgbiJ+PECtsN8J
+k9OtDgPv1FED0hV76DTfEwJK5xgtNE/fCCrhC/48jSWqgTDEkg2gV3mKmwIVPsqe9MLk7ALGZes
RstKwyXSjp2zZN0fjEDBDiDuICaQLiRMwZiZxod+1ay3JcSWjmQWYSKUH1wyJ0e4nmxXPZ4QUZUi
Nbl5JJfzUkJzCLOGIoBqTI8KybvjEl6JNMkgOiuFMTNg4T1BhZvJ1D+0V7F6D5H7O2snj+wOSZgq
IfCQQ5jVPnQPJHD5xa9UkcGBlLeBOwU2CWyn333vzBgrTGDL1re2N+dVpiJBnTsTQtM+JB/3dFES
QjHU81uBFr6zhRiwVEfaK0kJ/dtA89F6CdwYJXmJWiPyEiDzGIsPaKMKvSU0xTVr/fwo4w8QVfFe
TVfAOIrxqsX/t9nr1pjfbqpmHjjWmFLrJGJngiT49a2ihBJNhUzVsbho/3X/vmZAYx8zFdvsQeC/
vdMpMuMmJvRa6m8CUn5zzGxZcUM46wpEnKFPjJ1PGDb4eTWega6eFOBV62qreGupZ8LZu6L5BepF
RaDdRNq2GhWvWPTBeimWDs/wPc3IJMACIA/MTPiGA+rbSA+3kgZRd2irvH0NAMkH4ZOItcg9U+hY
2O+ALI+877ePgr1wgh20Wb+vP+gwLNGLHt0rTfVbkqmeghoVNoBPsq2PXGWmjVjbQwOcwuLNVvR0
e78mQZ956Cxh2UnuVRMq4OUReIxz904zNWC9adEvOLQnL8m9bAQCncn+xclbGw5RA0HsqnUSSRiX
CONrMS/C2LdjNGlzjaKbE/5jGdBEAPcN6sGAX4pXUWWzCIbkKXJ6YZxAxY55KN9DFPxS79VODuJF
m0GlpoHjF83D8oOZRxBtDgtApypxqramldnpX4pN74tLaGIvHy+hkQZRnh8mBl6MDfPPBFqQRhMB
ebJzX5QTQKp9YDtn1/N9913/sxeqUkxR7D7UZoyTlR1JAqyxNtp410rwC4T1D0PH4eSKLXkppP27
zR1XspAydQMQna79ckzN+Zh3+05Nu09VgKjxmt6ynvrJIAcd7azcO4rFILpehgCxrmzqvGy+BGLM
8J8lTXQo+y0yJASXmKwf6zskn9fYD17yVfXRntfSPcbprlCLRZPXVoGtV1yyN6F/Bx/eSCNXJmn8
zj691ypafQ4jHC9k6qxyGgT2AXC6iDt1BWLj0rEsRIfGv6viI5s5h+8Vi0rzlaBXeHcOw+0ShLpC
PykmWHrKtn+S94mufu/lzmCH6WoUdTfWTPdkeH49gYjsGa2TgVMIJ5C1m5dD9XpfoBfnFM0fse+6
H7YS5JnC4JAWVW0pm578mSUsxuS3tapwSWVeCNWNUnz2FjMMgOAhLGGFdYTvU+hwd13dyxrU0Ydb
CxdXbBi12E4Ywe5YFxhMJuB47T+jw9sLnNQMGIcly9FB0+wVsCnbTgRj+A1+0qJGjkMWIXwQiVlQ
JASBPzYgcTy1+IrMD2KFFFneZclxUiPBGO3Ak1duMm19AvfX2ioK4wRTN0JMKoT2MpAvF6FHXBNn
QJ8OnIiO6oSHMJ5LE7YCFQiuoAFvHhs8ChoJVwTXSA/vvflE+mchEgpjvC3Ka3ezYgo09bJ7l7w8
CE6eaUu3YrozMZ2P/C8Jpb6Qq5ia84TTIaNVAVIAVvC9budOJAqqBtklKWODJ6y0MPUwHMKyJ4Ym
elInqVNdwnnOpsaZSyro0pUb2D2YEKxD8gQWOpaO23xDO+RlRITAcFQgD7IljaifEM/0JQhphNQf
hyzvjcW8rsHUOacYaw1p9W/nyAPjN40F6inr9UiDdGoEAGZ+/qkubpW79DWFNk2bT4LM3gQ9uk9S
YiKPaeRdA/+KPZ+rod7OlEOeFh0eOthr38Ui0Q9f7Nx8d718LEOBK3geX96Dv/zI4s4QKTOi83A3
o0VCWST3sNPRI2UGsGAL4CMYSdvj3zTTWXT78x+eVyn54A9RbIbZDgHEkEVR7A+YR/b2Zja8N/Fi
W7QuBV69Kr5WI+wsq9rRlZc4DTOj0EKfJ5zhV9Bbzf0B6ZXUltPvFuA5z8PHiIYK2641jiSGIqmV
NWAhtb63AGFIM/YsjxBFbt+luaEurfQyE07wPNyyzg7ZmXg4DbmydOi1xim6bVf/MGb7eEcrXZGp
eIDS7R6HMuEcbkTm+S9KReRgWY3IeaQZI0YoGm3As5C4lH+yv/1K/X7DZAnZHe17A2SyMODERAoO
pUhzm8KbBs6EOGrBA0UwwzY51PjTXQJBu5m+kkqGbn/AYOwF1ZadodusYHsDtMYRaFUm/SwWI+QH
RDMOC+DDsymMCAgT8yfoqYTedBEPsU9hvo6VDxyofaiKJZQmAcXAqOqja60ehEMRcNfKmrus7nAl
FPn3qq1Ivf3vQ6ryl+D0OL8DSgC2+1SOIj9LVEH9kOJNjjIM1cpO496tt3QPZB9ZRS7nYEv2GAIz
s8LClFbm3Yqb3SklWFWbtB3pQrQkCUeih3sEnBsv5KpntPci60YBdzWOVNHjj4n94mvemBQf2Sjk
l54dez/8Y3tHNIbN+N4cmPZbXN0HDPGYvHBm6qbBdRSjSxAFyssYwpOI9WDOncQPrYcs6fLiRLjZ
dQHVm0HnaiXJnm01piUYU1BYEJmCknKOFRHFfSjY0wFLHxprjg4X3QJD5iCjmudbdSL7sOxMAzcO
/jBlxfGTUuAEIVEIb8gPS/3zKaJ9GQ30baHu76vd7h/+C0d9nkhoZ/cfrFVOAvkOULXgEcNYhkcK
L6Xozjvl4BO4o97F6/aq9DPRCNBEYdQ8GTMOSNtjdqUXeedn7Zb2s7Umt/6dR4v4NIkWhqOW4NeU
/zZuLv7/AahS4vy5PGCtWGNkTpnqTo8mgw7b6d28soaj32HP2SY3zSVrNktfbjV0VeFOQ4tuoy8w
1TWpXZ0YnnOaTdwN+NiXM9vDRSZSEv0tUeCV8Wd9uc3oAaUl6mbXrp9wjE9N4LwvSrLBwkhLLUIu
kqhS1FpItAJPCqKzBCQIS65p3xwCKXRkeVAoZCwtyQl9gQrAMa+Rsmm/ttCUGe+Oi0flFn2olhDh
3tBcb+qh7u7zKUTaAIJNqMWSoSWBwGAAFKdTC+I2A075abuqcKCR93Jq/Y8o/K+/IrDb/GNFsmDx
SQYbm3QkfG1M1yUoU1EOs+sVIhdg1TpH+p+0ZuNZBMFumW8sGl1uLFJoK+m8MXvLI3iq+jDwzjI/
sF7B4EoLdH/4xON426OwojHx/iW3yqPQlBlY7E6fInXUvXEWLtdHEiF7eugnbx7aCoe2C1F8K5rd
7HuLyFN259Qdt3TUn2L/g+AUFxBQoiUb2WANWRqVDRO5y3zas8EtOMXOa4HivuLA/2wY2rN15W21
4og8t3iD0q5b0nPsgs90IMWvayZ6NecVUmnGT3NMrXc9U8wFtbZSAvSbFm9I0sbLZTBayrY74QFi
bTg0jJV/DQ1RZf7TR4EULuLLPWHlPVhR5WXWZyLOm6NgW4J9LwXHMZEblZ8Wf7hsLGVv5VfFdkhQ
p4y81W6B5xnP34aIBj1XT8toI4o9AyelV1lnApV2NNj88JbGt2xgPC7/c5C9Z+W2HmCogAdmtdyY
jJnaozYsx+mSMWgMFw3Y1QJElKUqxWr40gcee7NnuCUfg8w6kb242PBJAFqxzjKn0IqREy6m6odJ
QWX8/Q2/2/xjGD1DSO9+nK3T+sMcy4w10TMkJIWiVJN25nwHKWmopo9yNPyXnlJJf7XqKFtk+SQK
XYdBUEN34uwY4WU2xbMptBnz70EJeVmEElrluySePRjiM03xJT42zGvf0cvqdF+hWlHWPICNYrGp
GMN01us4YrN4+iGq4xeYTCcJekqph366qNtQhinbQ7eRiZpRTsyNa4sEBw4pKU8uwF5WNrlytWfP
Q+5OoINk7fNDGWCZfI5IlxIVpJgJzapvOPHzpOKFEri4XN3Z5qxqG3O4ttx+Bybw1Ly3MbbHjSk5
Juc6xgWHeCWZhCSL1trOvNWcmLcTz75Gk+/nlEoP4Z0ixy1JBk2Inzwqe9fCmw3DW5vQkopKWor8
b2/XTY5JfuctQulCTPlTcIkJolH6zayycYl2j2wHqMha/IT7HC4c++0clipYpfiXTjrGqvJAOoYG
sbrZPKPrGRVzYILKuGDPQ9YfDNjduV4zM5A8jymCK83d9Hbn247hRJ/ewpT4DkDyOfamSfPhPp9q
gNjIDres9RealLE+hOt8us9KBiWbEvLCJG4NgaIo3Nwud8k3g04d4rMoTqMKzzOve9MoSkXJQpi8
kCMzsYb6A9GrGda/34/WxPTDIcRg3rqBs/FzUXP3qLZxglRi45U+X3FBXC/zIEGHTnLopUzQHo9U
xOwt0974Hlw0u6I6OPZgodHyeLA/Apjxcr9VafeIJLoEMeKqEleF9re9zPY5UJk5MTM5rXqwnkI8
OtxDd+tIfljI44ktg9bUEcyQ/mrj7ElfDu+tmTu9MBOBMOJLgEsDzBWdjsiZx1PSspfQiCkoU1lw
tbLH56/8itDy4eAuRutdPx7Fs1tM8Cz/MMsejgb6TUWJpuoTf2KJVelhAYg3qyNwIpxiODip6RIB
ZmWyZAggwUQfty6nyYMsm10rnNRMTkAcwm/FpHx6ot9ttQush3PoMnGJaFdLMkgOiZtG3IIW2GNy
FJdH2hjAkp5PExFGGOH1xN+lP8tYd+Faqng9SCCQwDvsS7LCBNRERHUEaUCv4ceAb3T9GuI9C3o0
fFwl4h04d6rV1uO2e925cupOoORQ+o7Mo9v+lccIAQcn/57z5BxcRwObcsBxaWTkSn1ZM+lNjggg
r8Ca0Eo9V8JCGBAJXi9lL9Zeb9qW3fFBzDNWHVrEEDYSe8EXAho5fuLNCO1/K74If9BmXfpP2WbL
TVJ6GYeCF43hTN0cPj0OJp+58UoxSr4cEFqLG08nDg2oKogdnUkGanXUMlvVQv/ees57JKbu5RaD
sp9B0AiENaMN6lxyfYzTJ3wt3u4iFrSuUIkjGbNy4PkrRK291itNLAlR6xMRCFYt/59pna3je7Jg
D2IEn5pcuarkAfKAQ6ExYJhRzpDQ32iG/t0It/pcaUwc3jjcQo7vvxlo8tre5mTjRfMp9I82cIOl
5j6WVhItzsoPW5wWF3tRfQf/DfE16XMCoxMPtmzP6X8CDBVGsU/aJRorgTTkk4nmu0JS9B5cCIVs
j128vH659eLSuI3FolsVPeqOy5D4pYTkwbZ98HMSxGF5riq3lIdxrtjPnIma4Rdr4cieba2RfbZZ
FvEIsnxNBXbJxPgPkF/yw0IH0Yn1EoqphlUhsAGSAQmBxZO3dapHL6uyFqFqpqseO042/TijTveh
ANfXLSxk46Fefzw5a/2R7MD7fSZWA9+ST1Mi4bjkEBD0+S+4rziOSrVUUq7mtFP+bvYJjByFKm2h
PQAOfB1rO3GUXxXsTIczo2NK2aZq8dtgT39ZtGVLoZ5V8pptWUpcwq+3y6A4HWHbzjO0iFSaqDJe
Sfh62/YSfnaWZSvDw4wnwcLaqZo1WcYqlRbAs/lDuskifgdGtuwmnMJwND1/8AM13N7FiNuCJdh2
saIOY8sDBHE/l5sV8wiqgdcXAmJCM8RXHYjrPtQbmID7ZidHinG1nUQ0xvhmRf5taMCClh/d5Dmw
oXFiAqrA4MM3VCeQ0LANi2PTRZJXKy57BrljDWds5M+lFHci/aqcWJ5rCFsZRaoKriboFU3Y2OsL
XWamMFP/zoVjh8hudaJGeyPzanmNl0hH0jfAP/bYUIRzxinYhPFAgVJvwdwlJ+NSB5Mjq7bmtGPM
PKN22qQwfnlEdLzgrS7+QZcGyohJcsh6iEEKPfGFKgienL6+SoJjabkhh5nWC2flkROSNWOHKBoR
Mwg2VAmhNPKTBUq3qwk8xtUMhFuIp09a6NEOd5kKs5goa6nMlYM6oEDi3cnOI1P8v9VAbAdCQbzE
K7rBtWKHGpR/cRU08rnXxA50kbr0C8jaRAVGUVwt0PPeflbD0p0sh4G1sUL+sHM14n04MdM2+Zw6
MT4FZZ5SHCNcEO1ERmzfM9SGxlhGbSISddVCsQbaXmXQS1AnenlG9nxkjiiZwj0zATD97FXl0zIX
PC7l+F5VHh2SUJ5UnnqozwRU3Zco3n38sONvYGFEwg0T+vRYEhlI3zZ7HtGd9VkZ3sxzzLrgxa3p
k+/dVTCftlgYaOQq9kFtzITgOiV9TH3MSsZ2h+C10TCe9pYAs8/kSOAFFP6WST9/cyYjDpe/bX/L
nifpJUXF1Nk2SKq++iYa5t2wP9lIz0HZHwNvQ4FikKXAdXt8WeId5n7TKPlEr52ZCh7B1/flmynb
JTopqX5NVoFAo7AAC3mxl+thCQa4WUoPhxZaEfccC3HScmN9BKX520KzMQZpI0sy7Cco7VX1EH4f
WSOHFZYhO3sSq89Qfmwypy8l/5X65T3VMVVbeReuUVh8tSNb9nmM8VGJjgpS9ZsE91RtX6n2e+lV
Z3aofaPwNbTNkQQ7h9ucV1TNaeDn+RthMbDHUhRelo99V+JY9BeT+je6g8qcuUrTrCjVbAEp/lpn
qBfWo/dScc48n8uEnpObgJLFfboP4zE46zg0Qanzkjvki5bBunmRBkhJvXAgYdttruIx2tr65Vf5
S67Ur9CqrNAjaTBuH35nZG2GWGYKArybxogBZHVYQDx/VQH+vynpEkF5GWZd9IiBkcPFhtsYnfCV
82Gy0hCqY3HVzMaNSmyJUBW2a6gmaJ04cfkMJ+5KfBelCuCS7NXCdzV0uEwrs6oUjNob9OgPDVAt
WsCFR2xzX+5C7M04ieoAEJEkbrmfRmegOJblKplZmUGjnXQGW1wWxjn31xryq3nrQrHy0NCfkVZe
xVpiVsxuXXShyCzwCLTDV8wOj2H8Qw2LgSBrTqCz/AWQ5Xz2+f7r1NgMH6yrC+iUDrwS0CnXwEm9
G+yVSNqEasTyn9Je5H64KTQhN/Cav+n+oEU73lhm6Z8ZUQtNs5US9eSTQHcfs/eQ+ME7dY6XBzXX
U10daZYOlbCqBfyqexZarcBJ7j/r0WkBxDVcw1Yf+K8UZcRVPyTXC6a4qmncKo3dZMm/BYBK27Qw
wje+aDgl5/k3A1n/VvsFD7MifcItiPZmTCJZnbhkUz5ldnpghETU1qMTsuZCeP/zM5TFrrBuo0Be
VnosPygcIIL/5uScMp0dhIBN6iu6c+tDUL7HUZ2XgK5V2sj/u6RQt6KWvOR5i97PG0CVvi0iezz2
/SshvfeAxehl29NEzZZ4NY42OetLli7aQa5RfZO6Pq/vNSOFBJFZT/thcbtLQ8Pu3MnNLjkCdV5z
SVIRyhlTGcJ9WAt8gjd6q2+DO/NOH+d3mlUJJlI5Npz/C8HQY4z/GrPl+ii2wjonsBuOyDvO/bG+
HPCPL8hyjXsoJJE0Ys7DsJNS+o9omT4fje2zW6gtf6uIIBHOiQ1RVSs1wvmh/XUrxse0hYiBs+Wh
Sxr9sn2zSSXtHnnsVYoQjwsyC+1HwUcSGFVXQySHvAwx6rfr+XeqUTRwR5lrpeoRKOXu+6atClw0
qT0TNWh7NsUuwjf/DfiUcguqWyX7FET5PtqmbilZjTXimlbmQ/ON998MmV0zpV1+n+eBoKMXHY17
5b6bwqRGkHRRFsSvy7REqvTZYpCtJJ+UydwpcKgyyoeBEHaRoGsEUsoNFRyx7NCqRQa8axEWX5c2
6JQlohkrY0n/emEzylyS5XrUIIuDRjh8ede68esCw+rnYChpwbwxrHpfzjA4Vf0x2tHimzuajp54
z9g6tCJi4H2yFOWMjK1RsNCo8Jg4tTE7tf+vnmGqzKCK9dfRQy00wsXIDZmdurHC3cizfj5msWpj
8RA2tIW2SvZqRvG+4UBcn2XKcLAK6mI6e4XkFrF3EnbnRSnLXji89piAdUYPA4OWaLSVwW9318dh
GTk33kTSDLfAQtNhRUje1SsAX+bpeelWM511rnp+PaFrzlcuvoaGDelEhW2M8sM5AB+6pedylTTy
5MuBQt0YRQ7DEDxb1F+4s7j/AtE3eXcZFJrJx3depSZER+Wri0mTZFVoOj0KUy0NrVzDQOwUSc1E
a6txmmxmPkIuvcGJ3loMkmzHcxridU6tDKhSB2QcXUTiNwVwuuE2S2Nd0AGhuy3U/xtsqhB4B9qC
kAqZ7kwF0vTTuG5Cv2aTqSZza2/6A1yJCtEZTuAT/HxVWRxnnQAG0kMDhPJ9oZNK2nkbKgD93qNZ
D0cHcKRgObuyL1W6V4UIWUkiwPQ8DnmDobZ3I5nXawuRiOwLeZwYT9094x6ND+TB8b2doJrgMWS4
oThaWUt5ZMN4ZojwzmAAP91oQYYRYDPHKUUL8XxCHRTxmL0By+mzqTJN0I49szWRn6BjjlXTwAGy
lpnuo2YzuADGZ5m15KoNdvUrcxI5stKwTILnuJxoMlfyL+EieuHvtPGot580G/xwiaFCT8KtIjHc
dGBSwyIgYw48NF4kh/FssSjy/RHmafUxqDFIV4cCr41n8AO3bGB+zZLJjp6dGaWg3UtgyXPrjnqJ
fugk2HnEWZk3foY9bqWwmFuuP9GU+JFUYWjO1c5liUVqc1dH81Hzm6ibGtOxWaIRgJgbugQlHZEZ
h4zOAdOcjw8CTkOoJKl7ERveRy4TA6PXENLAdlKZi4ES9tY1OCjAqJMXWq/Vvazmd+f7nOitT+zm
hk1rXhlrhyQ55n80/VdiSV+Btym7OYUkShOAY57C17uUyuB9thnpFlrlk1Tp6eLqSAnGyakkBwXe
4OmtV/krt+FrrxBF/lP46QkMvvnkDVwSmNl2G18NcGbu6gquvV0+n7GhQ/k/DX7qd9lkFhbKdCrg
fUJQqiMt6zMlz0UVH2ld9+KRz75zhCBS1JVSoDMhp7tmWSf+NvRgEhSyLZZZT6o36xntzy6AbkF3
sGb3E+UBrmyTOG1gNdTQww+HIuoo79fnL9jDhml3dFdPjryT9XcNS0SGAmWTYLQ2JOFPndHlqBTx
xXj15BvONbPK+IBXwPmd8nmZXeRaVOaeFQDyeeFF03bTP8htZyxPhHe6XBchjzSOC38Z2Y9fOmH2
uQ+AIy4iFmXuXILGTIsy7I6vYX5tge9614fAfQT2edB6904kHwUC7sWkiX4tmBZGmIakM42IOz+I
aXf3c7sRo+3oExKjRUHUdVcHU0svS81SydzgHKZMV68KuU/oZyBdouHV9UTz3Zlqi15lCQWeCarg
qrZXyn/UNT4DdlRIY66oiMKPTYozNJyCiZhoRztm5cWXXXeNW7yxWhz/5zI3vNRs+DJk7GMxjnS0
uz+p+Z8GIXuX8OmVPIZWeDUea5lpoaalpF/TnqVgwtL/v67NXsXaytcgv/KNqRry7an6FdGbFx99
CAkowaHA+64pOd4qZ4Vfo0oJW+eL6hUHjOTqUtGpDevB70NNqf3Oqf6LZMD/oQmhd+4b0GlMkcEW
FYxQeBOQ2g/AioGHfzABsSawDcrQbA1wz/1VRtASZZ2Se8HbZBwrhu21G+uvdQBZYUyoQ4q5RsOn
ETnKwuWnIBNUujcsltxYT7fcnC0+bFOEHfev5JYMNFInTAsvZpXEC8vvAR6TVfNpHCL6o3Sw1tmF
iHZLdmmmxFeislj0QPRH7cp25gqrP6IYshqF+aLDUnin4HiVHcVAQL1OyxZAjndNvqSSrsZhLW9m
NR0b6+G5GRtPCSROQaQxOQ3ePI0p+911yDiCLQKGz+Ca7dnpZAfs+f03nhJI+ztVtZqLBRzNWahs
Z36O50Bp68KyN4UsAOVISFKJJnK37JNTz1qI1q4N1zWKnFjTwAFP5mMZGq060Swv5yWzjRja3cqG
cg11og0XiXjPJtMfc8v/Mtn1BWULUp4hvbeyiUbAVxFCY5i+vteRBY/uVEHg5weDNblISdxLlTvo
lXNvPhC5n33321rJFq7OhzixamFWYOkdhzosyYrdVHMLKS1/BadSv4wMHPK3SL3GZ3yWHZLyesvw
d9sVXi6gsi7W6fzGiIi22JiIk41rMPstfGtfx0fHF3Zntj5/VCNX28zuI8b7GDfPmSs6hJDpP8Pu
NvYy2bVVEwlYL29KKv8scT0iEIEKfyj9ZzEBQjxgcwHRPTGEwJ1+wOjUR34bCD2AT3hV9N2avWDf
Vcms4PqBq+lyh9vsgmQHT0nN1s0bRgYdAC/nGQpa8vjiY42PVMxtbrA6kAqoxnZsIvYgii1tP6Tw
i/mlonF51brK8DxFHErkQkItdK4AmMtlvOsZLXzKS/Uipkx1Yl7O/S8YlME8/7EK/Om5lvbNpup/
eQ2voBQXkjOd+P78Nx1LLU65KN9OqFIWrwUvjey0aqAu33Qr0jNEoshzPZlw0lye9iiF4/YBhNty
PoliJxvRmgIiN98dpUfHNMZ+s0xP+WrWLm1XQ1Jdtg/4vE/J+BZU1I8r+A/w2RYKI12CHcW5ama/
dqA7mXXrTfyhoYriX9gQ02X/uIo/R4b8E1Ow+zv6glBiDQJdobXGr0BNYnwvQUay+PTfiU25gqLa
jEjyPzhrJNKyYimJxgbVVLZCuc9hrx9aZCPo/u/o2a+tF9Vtp9BInL/1PvSNfL2HdfyVTMOCYbBa
DJBwtnCZEvlILooAQDXP/knlQYuEgrKoMJ3ti30AdSGJ2l78PqU5yBWh+5Nrr0asezI+x8Otu+Ur
cqzOBDU2HKAwCXje6wT0owLiAWdeN0rIgyMaClsXwFk2TAbL0mU/orBQuw6EK5uXbBxAb2dx2Ec0
3k5KRfUmOWa45W1wcXsUeZNt/NJofcS8wbIh9qiXDyLgg1nDbIFLrBFUpxVE2xwSvSsDmsGN9gVO
N4Y+5wrw+Yr+UqXyU0lQT8T02Q/kzRss/6dOKJEmUgwV4qhFCWRZL6eN1qVJNb6je/2BAzjDU/MJ
tCi6zqd0IHpPM314/C6ZMAi4g1oHj3q8HbWwH9m3zEkAY9PHApADAQGjeai9+bQEMD05w2651pBJ
WVeNaJQKBSB+wgpBUmq9037Nu6EtfnXUM6cwJyO2FlXYybmPZrB8BKapquCm/CkpWTzMnBHoQqzE
3O2XEb7yxBw3T0UECaAKA3AeTp6iatuFnoMwzNNmbL1trFnamj7d0jhJi6m2tUU6JcjbXTeW80jy
NlRCHNZZRXwWyEKL++ib5pE0COrH3RNidaIdJ1lyNI6/wufmYcAmBzcs9QcBGPHAWLXDfyqqK6ew
YO6CBiYZsJTP4z4jI7AUwb5A7VrS3/CkOprortdpAwwZv7WBf/izBCfWrGBD5HYBmxgxmZMYE+md
amyFUTbl82/YGU3XF/pwabRAFv1jTJAF658F8PwKsO7ZYHukyVwEkS9jffB2S8dAZ3g44bSOZbep
m8UXWz2khNq1nm79CCbhc9V7904uwA58UGUKGII6u8cdmzNqp9rcu2aJDuxV6kwrrgXUjUkyd31c
mNjTKJluz0hqrjqC0CAtreWYBa7jOvBb4SuG1m+0N3mJPlgxr4JIDV4rJAvmrXFCNbMxMYyp9yo1
3wstSm8W6P4uaZgjF1nSFub6jhk/KjbKYkLHweWa1ilEUyuog0wt3/ImkDK1iFkbEHctxxlHr8g8
fX+iBizFy8iJLLXYMwQrlezz+5YDcQYUZfSeGaZCtrBH13ouELsk/GCkAj3Z8fK1UTMjBPw7kiob
bgcinrn6GUPMi4uTBxPfVhmGrmaOWb1pGAXaBXXvb6mKXrA0cNqsJoeo8xsVSTtp70YjmeK2P2nR
XBnYPrIhQreIaSwYt18e3s3zVnIIfXwc7hdJOYuXx+kh4IaglSrSKVyPKzmZ5N+XrKZq5V/rHNQ1
5oklhAwY0wVep3dNJGzLIWA+KBiCxdRZFlsnr0OprrdiHy96HPSpzOP50e5jK+8fVv2jI6Knkoub
TuHw25JSVCP6ggOS24ZrR88ys3mLP64V1mWNNBOFYfkoY8KigKq2kgaAlo6bUNkwmUOmFaMECLAH
XawXj2dHSeAGjhbDzZIsA65O6dSPEHxgb5n9cdCBF5A1xRVSCcefHxhADNf8VXeDrKngSmvlZulm
voXOSBKwndhREvQE1gkoeKAb8bX9GoTzXk1Kf8kP139eYo2pd4G+BJ6PfTPF4kaunj2Nuhe1XA1i
6Tv7yR0QqC8z7D6x//DU4JNy77mYiicACTyDHo9ZiJVy0sPv1lWTChazkCIkRAvasIrb5XDUb1fX
6FNPZBEvQaMgjUVVyk7YtykoWwL/zdw7lA1Wbd2ledqUZrfATRdf1YIDg2OzRYeHEh9kHKh2eQFp
i4ZH0oa07FbWCj39FdFC5MmGRe+PpiNCcJZOj/6Vv7nNCzuDaeuzBfC0CraNWQ9q7jP4e4qyXEEO
Ri4Snnphbehwlv918ZPAxGgexVAoBQnp1tQ4CvZ9IdRkVsb5thEXnEGC4WGoic4JhpiFS+lqqVIJ
+s7Fh2hVhBYy2swiboKNBRhkH0wUvwIDyNU9DihMSoCYCvEnNdlFUI0eFywWXmegrK7nu7QGX506
KYFTNPA6lufdB5/MXv4MlesPluxYV3Hrt+E3u5MwLI06fLPOflN6ihcK16GQ5pIMsokCbMXPwNq4
4Sbg8cVpG4LZDwR709e0Vw+8E4VLU2tioyKW2hiHYSPH4MwM1PfgOqRmQELaLeQ/P6pF/vLHn4hY
2jMtDtK3d0eRIlG+J985l6w/Wkrk4eq08nx0k6fdOX2MkOr5pZpCT9L8emLeSlzItiidR55wmUM8
aCLd+7PUYU9cFizWrP1VszU9zbycnXbrK+tuVHm+DtDXa6mXb6+dJuy9vhH0UNBojMXclmEu24+4
ndVjF0oYYYEurrJAPYVEzQpnCWCrxQQwGuNzsg72/LtPPolu+x7bC1tNsCymEsfVOAduvTbHiQUy
xuu4eWEqnLWNL90YDJuEXp6PeaM4jOeMcg71GElisGE6PfHovMrFD4IL/QPQkBYnQlh1r0KlExCu
Geknz9PKJnIUK5Q3JI37/FQjX047EXAAOQzYM8Mi6QGHHvuv2n6POARCreO/tzFy6uHBSMlUehDQ
P5plae0zNjUK48lx/uj76agKnxWhogrX38Y2jaJk6jfgdZEFmITwOPNnQDCZgoG8gLaEZUnz5PUX
KleEmUv3DEAVrk+h/+qDTK0ixYTG3PrO1GGD2oORurVUXY6D230pnzDrwWk750lIu2GG+Esihcwl
Crdhpr5MjjaGf84fP2OqZTL3eu1G09Xw6eulYR8cJ07lZZasd8IPbnYU5Go0bNHTWp3l0aUODsCm
QScimvfc3EcJov0rCYUaX3IZtHiWlEQu2KevYCoqLQrXBg1B08DBa1urkOOly4h5SzOFr9AJ5eQ0
3DiFha6u47jMT6ArYL9iYI3Qc1bzi/iLs6+SRUtm8d97juigbLo4e4wCdvfjxw5GMMalc5MtS+lW
x733ZFDnRyWylzZOW9a6ZVBqSTcHnAdelGkDR+7l+e2ECHfnbB54nyF7E7C9lTDYgbzX16hDQkKN
iDsnx7oppYkQc6dlK8NkqlWM8xUTcSilIl1UCPxsDNIPnd+qxrsr2sPJi3VPSzsQqkjUeuMZxeHU
qb43pfzURUN5okUf7ko9bvvjyBxoT/V7yqH/SZz6PcHoxf+qcG7YaDDGU2DAKq94LeNGQm/ZVjRG
xfezYh9+85zHCCWRWRQO7dpDKEE2xKhtps5NV01QDRTh5OkDeNCQKjaidyae0gStm/ikInkVo+Vi
l7IbaPxiY6qBm1Hl/hslZXORom6bStDO/QtcJSu/x0E3TkduuzAVovraXKApTkjejQe1IyFA8bnU
ZtLXTdjXJwIkCZK4+dEldg0GyEq1uUst4cJzXl/OimFCaClzIT1dNkqN94zwyRxl0eXHSbm82SIJ
bKobcBXtCpb52clkU591a8bC8QeTJMX1jYlPXNFryeiIawMyJfxYU0naBfxH2LzIFCXq+bPhQcvk
OsdRvDJrqiYPRHDlt9YEoldCUQHwBhC5ypTa4hLvPfJB5odr1IdywMSttKY6joxlLMCZD6YLCJTi
N0YO8f9x3Wi8iznVnPpHQgnkIwFxjkDQr1A8lDjODbxSpHyxjwkv2T6Q6jipaT3DNc/qhR23etuW
5ngWLMk5Y8YqSyyyzKJoune/6l1B6OYWoW+NJ7q83AfTqsnFay9CMq7/sdMAM2XtChWFWbdPyl7i
LGnPper4T2OmEbPxR6bEc2/fZo1R/lyAT4BF27e/l00yeLy+bb+qLWT0C2lrRwce/TSuKl6d62UV
OITusOQ+YeTmMWjBRhf73V3KYJ+ljxf4cOJWxj8tIc5O1sqFxlAr2IDbYlLLw6vqfah11RpSlitN
WYWvimGwi4/d2RZAyCySDLPGuSQ5OdU+40PoCnhPaeqQXBJvC/wZNv+plrbsGHtZo3TJUA/5cHmF
nr6Izpce0k39l6wRqBZGQHhMVs9JNJVmiM8sgymElqpLPx3y4WywsloePfQphmA6yL8FGuX/KFZo
TOBTGtBnAdzLxk49pSl5ibGxoxRqPmwP3Qe25mxfR0ujUuaUxwvxKrGneiXtWIWDewk7YjnPDqJN
QP4/JKwOsidnx8/sIUdx0rHU+31K6AM/u4tEqFEtnwFv51dIeDDxbUm1U1naPtxg3OQE4mCGlJVm
iOoeNwl+zts2YDn+FU6ZE5n0fAuiRb9URbRaK1jYB4UXZd4fFE4Wvqpr72XOmUTOPVq/Ky61lK7b
+xf6PuztstUt64trzfx1lkXjd66vaf104pf/HgiL9wTuYrKKyx6Lw+Qzgxr1huVcL9J/libyOmeN
ZObNVzH5MDiVWhLWxgpLxfos/JiAHMrgzA12arPUqrpjEDXpWfedaZ2JuecM2BHpU1QhUR4wHWD1
8KH+Gd5QnjfsxQXNlCO6joRHzL4kWWqP/xAiQ6ieAHXfBkO1HfAwOB6guqALERCKzQvyE2nLEPOm
6AsqwOyfCbNkl4ckBURpxLDWANjEg+19U3FRJB3jeGVQcyQtfybv/Udlwv+02LesV/MjxBDEM541
opjjcQIDHT68mNhIIQ9/V4JzQGfnRAbAc9vK0RTsGoxt72xl6lM73hRsXDi9T9WkflFLtjRzVVAh
Gz4WOb/OfDxfQeyJ6SDoto/sZ52PZol/o5NvpeNOmkiOj1N7lp2Yd133mkpIky62InOmf+NzfsN0
DIPIcNJ5OMwFw7QlRaKrTz93RXijumEDSVT+o6zQlkxPjkh7KoKHjkcmoI01JR2aGH1az5EGUSZ9
877rH1nQb3rsah4roIIkAoZAXmSC2uURRXxBu30ibaX6a+krNk3gGI7sGTG2VhRxb6hV4OCaFRyi
3eFaM4sL3txl1tGzfuAIZScIACoXH7Y22sqh42gEW7hOUFfoDdk0t5+Y3OZOQgOp6KZUE4gG2Tgm
1/F0IHrnxK341nNYDULyqZ6Q5MZ9Ag+6fUq6XBgCD8RZJypD6HCPFYkRx9iNsykhBozNSr0DDJBV
92BRSoPNGer62FvTTztXwos1PrjXfET3mkl59Iz1nAURKd3P/aDWFJetD4mydUlU
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity divider32s is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  dividend :  in std_logic_vector(31 downto 0);
  divisor :  in std_logic_vector(31 downto 0);
  quotient :  out std_logic_vector(31 downto 0));
end divider32s;
architecture beh of divider32s is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~integer_division.divider32s\
port(
  clk: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  rstn: in std_logic;
  divisor : in std_logic_vector(31 downto 0);
  dividend : in std_logic_vector(31 downto 0);
  quotient : out std_logic_vector(31 downto 0));
end component;
begin
GND_s32: GND
port map (
  G => GND_0);
VCC_s32: VCC
port map (
  V => VCC_0);
GSR_60: GSR
port map (
  GSRI => VCC_0);
integer_division_inst: \~integer_division.divider32s\
port map(
  clk => clk,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  rstn => rstn,
  divisor(31 downto 0) => divisor(31 downto 0),
  dividend(31 downto 0) => dividend(31 downto 0),
  quotient(31 downto 0) => quotient(31 downto 0));
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Wed Feb 14 09:32:06 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/Integer_Division/data/integer_division_wrap.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/Integer_Division/data/integer_division.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
q13FZRQxCOhYe/nPgauCgPZlgfIOl4+McJHb+9qBG0uUanqGl5fDcmpBuHyw/cCYDL99x5vXs3ur
uqoqoom4DlVxhuYsGVrYQu8k0oV6LuCDxeNt36UTvWyhMw1nV0GlIbdK/BH0J8nGwktyvl9kMGN8
uZSMgPsvSXkjSU/vE0KdhjqDU+7nGLXDS8P8QQSxqucNIyPM0UqUiZvA5H7FUAY9uMkDUsRX+NDt
fBWvC66uvC1NHLStCCX1HFaDUdfQ8qAHGyvR4BrrU2tiqBdjaJ1pmqGo0xZwtMYjyQ0THkBqrDkc
QO8/xGkFg7tZCKsLKvkJzlsKt+1rxuVNBXQVgA==

`protect encoding=(enctype="base64", line_length=76, bytes=449200)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
2g5OJEyIreHKNHZcFV4WYEM6RevWK89OefIMQipsuX9IiYLeQ1Dbw5fmy8OO3QWBj8POzG3cs88H
FjXX6kqEmetB6ZEX+mPBtU795oYbCLzU6rbkX7aMUBcDQxOLUYA9tMf6aM+OlAT7Tl69FKwgBvyG
TKHvefa1KgqxmJD+caaHDxXZKwqq/i/LsfOGL7h5Bb1bRCIosTLlkSpoae0fCzIoDTGESFZtWxrv
bWbvVB8pvlkRcDRBMwtB0BVGXh5KCsnp+s6XAE7BgvjVZzxKQHQuUGJf8FeBwhL0dh9V2s6sgSwB
gethPFhP3KtIlzNZ9vQ2z+PWJ+HrsqLUJbvnYRmjn6WNHvaMsbmDDKiJkmpl4fIukcsgjks54HbA
aJ4C2hRHZ27DbM/ZyUsHwO9Rl6XopwS+M/TudhWqxErN8CPW/j/vzd5500MGc16CiPs56omnyh8p
/ez2Xvk/Vh3CK+1PKcT7/5pqhhFG3O6HFHsLocLlZYfrtJlQiKDbuGNWDh74E4U5BlYA2myNrEHH
tUiBHKBwZ4OxhUMCtWEEp+0M5zGGD3qUxlufmTlfoqDy6BugQa5Ya5u1xLJqJB2Nobt2A/u+merA
Mtnyd0ZHhFEzTesoo3HcqGfx0FLhyN2osW0XQekA3doFT4Wuv2oLMGQ3I6qQ/85ucZUYt4NMqJOL
F3VKgVhaNJjHSGrY/1o2Wv9302ta1Amt1nc9eyo/1lQKMng6AHw3OCI4MMXFjmAm2Kcjy/INJETz
1/heyjOkwRl0q5i58CSyzOIQwaIF6Whmfw3cO9mlXmEoILCvYVjMc/2fGWdLJ1sbCA4XcA22ktS5
FpvK4e4yHsR2a1JTuRQSBZ66ABEEZienN3TX+JMnRt4dqzru4y6BBsDQFCcTVlZo4geyrxY+eIvo
RXC3jKGdG+kcO1wBAGbiEgF+VkC0xtRuxthL7I45aWp5m/jvnQJeEbv3CV606f1HU0jtM7Pwv9LO
llrzsezNG1P+lHl0h6YJIFWyGY3qNtLth1XP068YNJxtSmWYRnMrqC1Si6W6qjD4QC6rV8Hh8jZl
dp4Zd0j8FeRRjPZVgMGdDQ5zGTRIjizNuiZeAvsbpFaQ8V4EMwYdTZUaXffwLkawOVcVXS+X1FUY
6KnbhnqxTMgBq354C/frc4ICYkRljWO3d9wMlOduoM0dWAGk+JK6F76spemDY8NUNkHDaVKFTFG+
jFp03dC/d3jb6oY7Xecfo2mFNNClhHLkoCo3a6Yf+WHEK43l/CgGpID9l6+RtzlGpZHIsewjj//7
RR48mSAgWdnwDmt1353pGnE1UviDaD8raJkm2i1/tqymNUyW0IdvYVVMeJjJ6cSsfvC8GWMYOMlP
CU97Wj3LhE5pNkTFosTl4jg8hU1+CTBwYz95oxgOX0JeQExnQEXkkcM6//PZVa+ugj1m+xHz4oYP
5mSdJlHSurPeRrVV5kgulH7dP56wwpZW6MB9Q11/hUQ1rOZIkr6wii5seLiaij1H1TQT0Po6J/OO
qXh2GjiSyxz7QwD67NIX4EaVIdPqaPh2wpB4Rx9rRGWVzKkCc9qJJsdIqOpEILgo3lEbCOuyxjKc
+xk1dEZfq/EEUKsyPd15bYcgDNWJMfk59true6bwqtfZEa/KW0vdlOalgQ4Q4vxjaSrvvEuBrmMv
CbXDUwseAqh0B0NDPdvpYFO25OAyTTkMdj/O1Uc75pkY99T+6cypJ+US33f4M8lJ/bhUfPMMIayn
f2KtLb+IwJisuSld57JTR863hWLccoe8tQGM7u2c+CDvkxJvYVNWxyQ1MGLzf62xrAEjeYqEVTtw
ZaaHjvlYK42zcQwczpbuGSOmnCMKrFeZ53Hd9V9hB2wMEvy2Cx8WwSyQfgL6qiVAhq/0glTsQ6Qj
t6HD41loc4Ix19fkZHGVpUdjfpR0bBa+In7z+9wI5rRo4b+30jT+gLR/4jAnuLNqIDVBmxdk+dHp
S5wc8vfupAgexXLnbRXFz6Mq0V7Kh22TULk2EiQI94wd0HWBAFrsRFY7dEzkybUt5cu+vrwxbslr
vZ5Mvuw/6Y+Fucz8cPv/5KG2tS87gkwFsidNixD82GbPRI+t1dkxtMAiUHUZrHxGZtFseFIWoBrn
RFwFvOT2eyNU4lUV8/lUDNeUyqhuR3LeewX2NGK2Gd9/mkQQ2oNFc2G9QpOw7H2wmSjFBOeF2NDS
0FB+JwDQTal7mObkcP1x6LdGUu+UsyFC8byhXviCOOVKZ3FGZISzyxeosLAx/L4VuAQVvpyHk+Lj
e+FykTvCoF3fFyKBFcrdooeOD/DreWz2yAs0awihxp2TFvNgZwc1poY/1RY2hTWjhC/aPHPArXV9
XuVz6hErXchkPFHzeYPug1LwiJDuiuFFxMq8E6MGIwm6SpOso3vYT4XBbV4UZnRw1ITUV9ACvMKi
SmNNlVmUj4mB3mctYGCDrGaMww62I7qxOyOh+wM/5l6Al4ZoAL11lPO7+Kzr4RhiXotEwb574Or9
ONTABUjoQljHxJG581x72MAfEtF3bDTCT6OChbnupp3Ti9Kiz/+Of1umvrZyWDIFBiSgv7owyi7G
gFYvbudxWuJ8fHCz0eLXZh2v+VVQrzSZQG23H+qpgsFlH8iFYEbXU/ujXJmmCzEmI5BjEEUCwZUC
yxTQ8Bu4cT7NxhecgJ22kQYjNERkV+7CU5n0sTLgMBdMWR288t8SUjDcFf7gN1t94Y35KzU+dAnZ
46I3Oiey4eIqMiQFUz+jC6VDY822AkJjxm6Zp3OCYeibq92aKBkS7qFL2Ix+JCvSZjKUChjT59u0
G8tYk66G/oSSfG5s265Yl2BWGAlVQ4qye6S77mHr+Ki7xCkTAP8SWMtL9aw80QuZTasC13WyMtAj
b0hXGNjRzOCHOt4KwFrGqSwsFSZziFxiOnWmzsUVdg+sHn5YyErC06vx54GGMmjBepEK6848dpf2
ZMyNiSnvM9M1lahmG83JPVKw09Bdi5JPiUNQVJSDuWhAMjLeK65ibkmkUq8ltPOHGJ3MEE66Kf/5
cF9Cflkf3Lza5SqgeGk4t/9q6Ac37DkfDSok+V+ENe4unIapzN+1GYbUMeNITkhVsnoeEkr9Z5/A
GSfX1rAb8+oxKbz2PxqMYjwBwAuDeVpZOh9LktxRlyj2s4WZtMwa1r1kLLeknLE7VpJTENgs5MYa
rfP7jf3KYgrAjIiYCAhwblSkwvVd6aAw/VpsTe2AdO+ECh6G2B4RLFrV/dZP87sRBsvp+dCVDu7M
//8qlKYIe2SQJPk/CKrcV99uBxYQGN4SU0o0S+t5wUah89mCUx8gvqLsv4LRI+m9pYM9oTispjdQ
SwB7yRgSja9LwCaKH3a13YoAWoKnGE7RTT5MgoUG+vgIIT4venmW2eX4ZQqlJN2Mlzqws6slw69F
xG/NuX88FJibNp3rXu2XZ/VLXrZz/gseSdFjTHndRjWT6J/6HJN+LBofB2gcVcMxOfAZ6BXKw6VW
2G3DC66miNUq7coy9uMgRZaSx3DK2kDz3Q/HPuyQDGNdmwm3crdD345a5iMB4mlK55NTF19ER8XU
qgCHWcgQT5N/4CJFVnxCQG1ZaVxOyGUqpAbWQtYo3K5W5yYnCJeWCLjaJuj42kkVDCLFZd6VfjVL
05UiOVt3bCKbFdnH33qCpsFp/t9DPF6kng5BJ88b76nHRILJnCNhe5drrwBJVI4hUMMvI0hqH9/G
L8nDKyryMiUp58MrXAA0Q+AZDeMOfX0KlJNo+mZl8djQEJ56TNY7g2ADRMrqc45f2I5rVGmgHqlG
pqsU8sN7ThfCGerO2LT70LOIsim+hZ4fVufMAyAmoNuuy5nRltSUGp+KAOAO0S3iHvYwyEQqQdVY
ErWFHGFV52pggKTQT7dd+AmPHdHFA7lop63l4sAjTg3bn9eOaxXNaz/BBVR4B5F98YSZAw02sToV
TdeKKpqVGA4+gDqIUH3oBRX0iGhR5KcRxW4dfXTv+Q9w77AK7IJO7v8wmMQJHMrcrOgDO6kxMtbC
kcU7qi4mA39S4+vlHO62aEMxoYmDbaLkW4svb+HruphV2w/KeNtiZXqS9eQIGoRgNXC1dmEEY9LL
gXYKHSADbvHsvdd6s9lRn6WdxoBic1rLDD4tkJg5FGKO26mSxAMsRrdsmbiQkGRntUkT+9elDT4R
S1+9qCaA22BLh+pghgfvWiwACcI2ytcwtSyyNbQip1p6BIxiq2eGnusmszGQsfMQeLYEfPj6YSgb
nb0nzIbBBurK/YQGn3vyawRhVewNsAmYTO/ATAJEVUcw5Ey7PkAQ9VkEmNvpye02PELTkXdMniV+
6arDTiw5vzG8diWnaIVwrqewwn6I8Dx2WxV1/k9ofA+LiG+HIIoyXrJXsGDkKu2MUSewyRYKmuf6
xqUt7g6nisPXHAqmjrnUXLerroYH0NovT91wNebd/RFl+35KgZo5STdZ48/C4tq6foDd+W9lEh49
rIsjnOXW64uN/wsJPDSfEZQr4aSgXxshq9K7erO87E9kQrjPlhX+FGrwcuMo85SgCaTXb7e10Rxu
L7t3G/KJ2Bguhyv6z7Jsy1r1B4s6kQHCTAgH8aXu0jRsb7QpMGSidThq1N1hWQVAJmumbLu0cmga
xGB4/T6Vl286kBq4N9I3emBS4/7+cqgIIMkXSsa+RJWb8njx9hWBNxEw9KZPYZ9HcrL9IUdWB6zl
d8ofIAXH++CeU/cQWYJGeBEdZAmH8qHqm7xy/5cTZEJ+tDowYe2eh+kRmP2qj7O9UPqp+sylIX5p
HPWwevSyuQtOBw8zAcDWlzJa1ujuHJ0JbZcAQsz1OvMFNvLEXbRVFhKFde3rvp93FNvaq/o0mTc1
WFD6JnVUVPWpQ/BmX0Xy+KYIvT3OtVLhTlNU2tph4sVgznOEIcDqYKyMcx5BuB5Ys42/c/DidzAD
OLdmDsH8/ATOEEx9y+oz+xe1Ff4tVFd3pT2YRiHs/W5ndbkFRRNOcr926SUJnhsa4aqgOIlJPGja
eqQZSfjNJ/28lZMEAHaBwU9uNU5kkC+S71fcdtM3iQgSs88CYqXEUaXnVdUZxl9KdSnCyB7DZlIR
NpltBO8sTVblbGXfMywhH86cApGMHfNDN158T0u48jldLaNPW7gj5LRBGczVyJuJPZEhovbii4Qr
8o0bHJlmNa1opLVJe6ChkETmmaeyIX8P86V8ZMjXHjOQD0LG5do8sXJ9gn+kyXi7wD1QI96bu+8z
MVetExtCaSLva5+1ZkvBlErnhr657MKB7xeiNhUWfBnlYe5xTxGRaOTsCmwQLx4nq8bfLNumxx8F
EQW2jPPyT6ai/6qBGtoEQENE93ibMGi2iCFwbyWNRY7fMHljMuP2TLEKvJHzXDLRqs8zmsbJdA5N
T9d26qsQSCLDBAbD2zhYpTqSv8us4zOo1BuUoZ0Oj8qpulNBwEyIdTuc9gz/j1cBKJD8DncBSFY0
ZRBMGo/mxIsXWLbE3yAYZOO7Ft5reotLiVRub9EQDCa5PxY/rXYlp8n6c8VVaoJ7Tooz5OTbbqv4
+7pXwAoney4ryam+Pnym/QQcrA/AmaHoI6BDwUQtUEXB5fBlpBvAVHHdKA151qErsCCkbdKleGE8
Ju7lwrM4LGSGpTFzDkTD87qisOxkg90jwKUMp+H+AqqP15ZoU/FiBUm3BiyIzyjZ/AtM2jqZfoXl
uBqpmhNCHRPwcaHBzoCs7fZDbn5I2IDipJO0ZoBtrPk8RVul0F/Z17l8RQtdoHbefHTueSn1Q0YI
Ba3Cj5ceyryzfW2pkeBE8ZZ5pFQJwo3YfTbvCEFufcfeWWKXl5XnCqkx6GG2zaP6Jnelc1zXJFXs
5jcdR2KsqF81mC25WLA8RKJWeTIjdgiQoOJecSa35FSD6zqDPZ4dV2bbFSqGqlMbFDVK7eARcfwr
Snu7x6ORRXAgnG0ir6djBUgdF/MdTSqXPs2RQlwUaD9xKIrI2UV5v31U8K8eQOnuapYAdd/ZoK6p
O2WPAX7U9dOd7NSnooTKTutFEmVmgc7mwqktclCHF9anH8MA977YnJqMMglA02pPvr0lXNsj0Eyd
k6w2qBEvtx8oe8H+OH5QlTiTrDB+TkNj0nn2GWZru3NevBHgwfbE84lTCoMdk38RS9oJFL2r5aQt
1dkEHFaEXmasvhnPFSuOxsTemExUMkSPlfCryNj+Rr79WM07dL1n0IAg4PLJHMEfWR2hP3i3IUMd
F+AHQqMLdWLI6dtjRd0bbD4YST64QiDTR5xvv5Fili6Ybc9mjvtk447O5WdXrcQGrvoui3a3bHtD
SjW+ypEEcYnFvNaIXlxRuDobb7EES0DYN6bUF//bFm5WhQm0CZGjg8i/TLYW+h35Grb1tcJsY9ZH
1T1xVQkHq8P4kXSJpFCLzn8XVQyoMcScgv31rQbJK57ii0vhX3+t5OT+0B2wl8cpCysR3WErPbKx
wZNvav6Q96pEO3tLk3z+WLad9Vw6+VU3ZPsn0u3gIyXO6PKvJVvZCuVeKC8jkcpZePxm7CL3ycAH
ry5C9DYDmVJA6NI6IKYCbEiQCeYvckm1ulv19SjvM4e9D7WmmGdHsMAGPN37QyLNijJ14YHOZfxq
AKB5Nx8VKsPAbDJ4FTGDw5TQozahKk5cYH4E3KVVekEq2XnWCMxh6mCu7uncqAnNg6vqv/z+bU+o
QfAJScN/mddwYNLbBRR5KOc5DIF39gJe0gVjmApNGmHkugcdFVV+qqqlEjZMbg0ZPZxOf6TaYp8K
abpieydJuQZ4m3F4Z3MaHSv1t7c5c8/0EkpEQxDdSpTvjKdkeoDHAmNXGpIkBs65dx+vTGsL3NxK
wXDYB2Ej7v2yNyPqj2YUj780V7PIkf4JTlPDNKMt63Qb8aNMH7g7jctUGJnIvGucfmmWg3cCu+Wz
8gHNQY9SytRGh+FdI7+EHK9OvYr2DCmZlxUlmNF1SEOxcBi4wmNgjjEaa0qu8Lu9PglbEWnC6dvI
pFBeFv+RPxyK1rQeIFY3a/PBcVljM3seJd1t8NXwrexKoipTdCnH+bfLqoB2gxoTfxEcka0x/iVI
QPlZnYQXFYpF/bsqkiD2Se0NcYZjscIbiGi3gtGYc+bX2LsXH/guZIPioWHC0H5BITIH/5Zi/b2K
CmU6AUe48EIy9lXJjbO+OQ89a4cqU7N7tuk3IXrmusZ492tECGHQEkNdUC0oO1eiB3w7cIOLxk9T
SkvGhXWVbXaHBf//2doGDa4jqmA0NNY51VZncJCQWg1ZRhb1j/Cnx3sVHDUyHQw1op5n2ia5hGv+
kAro2ZOVEbO7Zc82qY6kcXQeRuq+duCCT13Q+rht9Sthcg71xv/7geN66rfOV1lzr74gKl0Xo3BP
sQ/G8+YTbohL+tGq6Z4+67MZjv6QtpfvJ1F/0sAjY7xiVN4pK5bloXObcfQGQL8WoTXFqd20D734
s7rXiGlCG9uYKm/5BAre64AE0V5Mrzo1ch7ABRsxFYav64WXwEBb4d2R8EI/NZ75DrB6HO8iw7O/
L3fU22BB9mcQo6CHjESMmgp8yjVDkbii+6XeHeU+ue2tm//tfr7thK0xSJ2m20oyEHbPwP09NtdW
xH1pzo77djOOhq1XKBUrBky7Jqmtwkdnk2ma24SJIrwWY5qSzWoHTG4eNG9a9QuW8lJNWUbqP67j
LZ40Pdz4FOBF23+cnH5laxRDaYvsiQlMNlLHmvgETNOmUtAfC2irPkx9gStKzCISTh5r/Cs8mf2Y
SREWVV6fo9pEe0/wFyzd5RafuDyutz2n9zN/SDqszfnomHOUFo2ExjS3JOXMKkKBuDBqWW7HYU6b
W3YvADvP4zLbqN44TIYyCqalp7F+BCPyk7/wjvFlq1w3rl/blWZXwmRzfgMeqJK3yfW6Z8F+1ii8
7ql47LkYG5CysK3NjaX3+rk+Zofceqm8kvsaqYM3Gmh9zO4Que67sj4z/boPdGiKvepqOl1pV6Ub
pK8nI99+9o/uUyjjjnQgQ1YorNH/ZwBdIS0WclVl0/p3m683z8qgZy+BXnxG6llyCaUEk998a6OE
wnEVqVyQsV5PdS97VIH7GBSQA0R5pGL44lEAsQl6wPXuJKFbLO9UQzVzk0kvQGQyXhbmFz0YIpV5
wIMP6xGh0ZbaY+BHB+zAFMKThfn1/FW7n0yyuTH9kbUDKCjhbMD8pJaSV89b4qh8trxpA9rQOPsF
ZNhPYaYoTihsEjbDknEZwGCHOEIg4foT9AC+cUB8xmn9umbazTdd1KC+emf+taHVAf/mnU25yVmu
vsh2JZmOwjrsmU3AvyFOKpPaelB4vOuP5vWYqeJoAauuUrcGY41JVZwDd39jVK8xyewKIBQXv5zj
bNCG/kuFRdv1fF29HO7U5xMmvwc8pyAaIOXBYdLxQO67fVfBJEbIWYIoVMzQ0xRK0OBIOvMyMM/Y
zLM7NMZcHEcrXPZXxRzMy7/g9tvIHvO0NGUd2h8NdhajJGGXvm4EkqIYkAgHeEGkv+l9ewwrUwdz
QwmLgm4YjQtldoCxDhyNHuDHHE6HetSOy3A1DHrgvRt5+xnSxGbHCeKMp4QI+4wGd3IFswTs9NRT
DW5Yjl5ImDiV2uaQO8MoSfRtQceelFZPdaWS7/jOQRViuTqua4vYECVHJda/wcEQl3p3VN9r9rrq
U3OcFb+0YR3rVsk2iEBHp4Yi/qutqEoc0s4t2UVzqCQC21vRNE+iGEOH+qsGx8iHDFNqP9Tu8Br5
zydOm/R14kC4MZX89fsTXx6tgPj4pUsQDlsuaGc8K+IrZDN7Z9tDe1K/Fn6q+Sre8LyMtS7Va/kv
L5vlufpWNn36eGqvVBIcB9sErgPqu4P4OkvkdFNjAh1rKFG4MnpRZF6TEonTjNaQd2FRf82B1Fs3
YuayEkEJxZvBJKmf3vD+3PFWSK3scvX+UAhd3rziE5Iob89dCRVf0ndBqF5DupSnL6MjAGHC1XEc
/QwQlr8n35ApQCJCkNypevpEMu+p07y32rr0ecUFAfzO2pkvibTbxTgwCBHG4/gWGEoGPaLVG5/u
2LQfqiKvWBF0mQ6CRLDn0BVlvNX0bseVUMJheDYyfV2BafQ3vlHJnV3tO39+JYlZib79vBVhOPhL
3VT7wksvY0nK85NJCWeG8HWWwVtScqIj1nkjJSAjQlLKnk4gRAEXrlrzzkAgwyf0JDYUxYG2OsFb
wpbBP2E9OBG1EN6SqJlRWHKU6amuV58uCJ+xVV/2fxzOTorXn2KyalI1MXyyEj/lZm80S30oXVFF
vRepgKw1bFXAYPB/X+5Ny4K9P2aKPofBlDXqq3Zg5IxosyWYVnNfPjI/deXEhMZLHoQa94O4jjY/
KTnkKVT+3ZGlco3YwDRZdHYPaEH1TKrr7YYuohM/494aF44nS6KKq8OqRIqUGEojnoj7UQbvoA+1
QudRs0/G82+QyMWPaUzNpVwGTv8FcG2BaKhEiUtc+DC5jnupjrhI6ziqSpcUan+Gklm0F2to+dvy
dG1yP9csfPmM1WKiOa6eT1SgMMq35Gevh9hWzp5vkwIS70BblUMKOHuoCINVzFGcoFHyS5W0Z3c3
bdiD8JXMVshMfcm4Ds+c1k8Cl9fDL+rVs7uncdiV868SUpp/0MsI1OGqhPNAf1D8fAuJceHJzB1W
Bw44k+BH9/8N4eH8vw7jZ28vq81XO7ORGkb5ItcNLy1O3HGKqOYit/S5pBKmEvcDS1iixERcJ8RA
Uu+fUFrF5R/Y2Dh4V/vUOQ07u3qr8oO72EOI34o4JTcQwpTB2WfHlrJOFPsArzXm6L7tl1ipbEU9
MDLhKUz4I0aqB6iUVjkS6rVktfclTk0pskkOpSAs36MTTfaYGA1KtOh3aQZUS60qbBuz0pu/OmOG
rejtil4OAAJep0YccRebuTYynoUzvuDFmMXfCnHUzFSWfu8inyk9uuINJCnIdzO+ScS/wj5tyThN
LNFyCJcZ4Fd/ope63DAB2cB5XaBsImceca8QDWlXQx9xqjPWgbDVpKGgpySsqzG/cmeKyMdpRktK
kSr97s31vLJ7hAsoezNbz38XT5Zj3txXqdYBExh7v5wUC5S8bvKImMJsEL3iaC7EpcEwxyshxHm/
4T/bfRFOSMMkTZEKeRsw/OisOg7nB3bDAOfA8DmWSYPcYQUO9KUus72D0yNibXYnFffhgym5oUSG
OKMTWcDtilTUYByAJHSWddeTgALObeNBMq/La0/co8/ZU/z6eRrXJAkL1EIo4xDVAoKAoRktxL7H
gGd2o69ekNRTFPogGv7rryeNsUc5xUkNdAbfGqxryc7OcqnUEl1Y9c1mMH1FQeb9orE8cBGW4tBt
deAf0nvGQ2tx2cpQdbJ3KWfJD7j5/ID0KZJ2EGwIt0HJqgjQcFxyJR/NMUqrgamqMYfcw5s+2wsf
lbgufaIuKFgg/AR+P3RlZY4oQjK6bHqBKrxVrILMF+W8BkB9DM0TuNqO/Du3mf4tV4zqWriooLZ2
h4j+bn7B5UPv7IjFumjCiTbWHPIWE0B2sTylSP6Xx0J3ap/3bpcU5ZzM/UhMz6p5KedG5urPPpYe
5tsqFGT4A7F/ll9wtQWNcgXGxgm8UI2ipudYg7UuZwa6ZcjE1Za+QtGUu0bqSjsay5QzaorHmbUt
CYsmW0ZTWWvm92SF9uEPFSrHE4t9fEirhVPuEp46K3JOQeOaLKLFip740eTS7JAA+gPaaXt+R9cL
sXhPFj3eO1PnC/lm9O9p3cyK5GpCQiKx1HmtAI31FPqGHRdeBZOvgaMl6ZwB6svJRYhfMxBQg7/r
fv5Uw4u5QUd3VlJdok3AdFnlyk5kX+vpJcL2AqZ06K5L/lbikrMy2odWD8N70NZGANt48gX5Jrid
3JFO6ua2i7ZbP0HYPIZPKTvoTEivCl9xuN34Ag/PVa+JUObomKy5eeRmaf9F0fDpNwxWrUWwrQr2
y6ejS2rBFt57UwwHBlmvNUonPlAbkEMZ7G556W4adue8IWOvBQvpSgB1Nyfirodd6hJeaxKoe5Qk
N2WLAi9Ff9TkzAf/K0mWxDpLvT5Rz0nxEI8YthsbOezGaLATaVYNVQIqSnrp7ijJNMbMyamKrHKO
cMjhqnGFFY8CaH2qEsT2ErOVNav6aAEm8XpvYzlLvSsnhC+x0j0NXxAB+1bJsqGU7IQKaw1X/jrW
LO6iL6auTITzNtfQiFTNPG7ZWeWu/MIMJanltn5OKM1AkPSpSs1tVXS50kqBhNBWoC675arymbQj
nTFa1WVmoXifJThSem7wYnUfxEsOT17ZF1u6lI26XP4GbV45aiq0mF08MZ8osSYtk+dQTdsKb9QF
FGv8mOar+Cs0QQ1V/qMplI2XJ8IJx4Yi+BuPCKnmFKRq8IZLi2LdV2sWtipcEQA1SRAvVkRe92Qi
1brNTQSRoS6JMSij3D65aeqyUShw5dxRREse1KIXbtUYF1woB7OzI7Er5ldDLSLImcqb/VcTiCRu
jvmFd/+DR+PzQiUhzsD85or66libB2lUX710kn7kNs6KemrGijkxQJqQWCKcuVF/fTQ5VZA/e6TG
pSpoc43pWu9Fy3re0J6gDJ0PfJgTxGNXwY5wYeTkc9VX2IaBI/MSWjCYgJMbcIQ3mqoFFQknTEXg
kmRw3ix+FaX2zL1sIwVE8lGiWV8e+UpCvRRoBODwhSolYPWghHhEoAP2NQrZm3BThuthKAZMk3uS
J9eO73Pru1hC1qBdMhLXd7RaZbm1T6fJbHdvqiRorcJdFMUM8fbduBaTEhZB/p5zmbQ1By3/5Fav
A+K8CDS6EuNmd6VQCM/SpjxyYEj/SNvhMu8Mo0k3fTwc6L4VuYYheIN9Tch3lQuRORyCBjDJ68OU
/x6edZEw2YmrJILbiJRpy31zAYLA4JgdnmfkdI6lQsps7fdJ2sqf0lQkEwmHvQVllKyH1d8Bokpn
Oe+b5+dxuJ1Tl1jnafOT79z5ZgQVYH0fP6n4Qn0bicdT/opxQcgYWkOHZOvFVKTm5VVcFOVBC2R5
fEHL0tUt8ujHSfhpAv+gGUzhLuWL/FlvqDirG1/muLsnTTswUHFhKmhq92uFxwX1ifr4ZwYXBf8j
/h8OaUx2OK4rNjMSyd3oacCuxtoljf1fR7E/ybwIOtBy70vjd8OOUscXTtS+JfEytZe7wM6g5qdH
YvoMjBjfngnD1n02iXdLrbpBvW2glt9Kjx9HQmE4vRbW8u70bmlxe/U7ta76w8+d6GjG9bL7rKc4
zsm/zJ6r9Kmhpt0MyylXp9lZJI3/Gzel1yRmo4LUOB2RhqGAfTkDBJQUjhkAXXlEWgxjG3fPMBmZ
S6neJ+Rh1XFdQM+kLHnP67YB6WW80nZ9VjT4FGuLyJWBvX9zt9ovhgpQKh3KmsahcejQuHu06eDc
cCotapGaKAJpUVO9vDRFbDwMuYKnPpyo+UH8T4aoOPfRG/PC+6/cWzkJkAye5wTHXBkxMrvsqX7B
P2k8Mzo5gW+IcmRiBfID/w3ra+ReKOJskclU+gR8qWNm4OosQyFBUgpxg1lPZCldNIuaJOWLW3R8
01y2GsMFHd4fdHkh1qTm3e4Vi05mVN8IxRdrGxCerWAFyVr0Wlac3nshDBXp3PpBxh4jH9pMrGOw
Sa+Pw13g68RwnpN3SQwtTaBln25dE/XnfgI5wdcgR9DOrKTMZow21K3ufCCjMLtetwE8hu7Jk7aT
ZL9YaeTCAPWFZzADfrg0sXbTy5xhusAC4kscdeVv7RagckssAn2YTBGVejBnxO5lx7lKdaJa1YwK
i/JqFW7H9ORHpdOsKs2u64K62cvOQqu0ONJ4vEjGIYLfBwfKV8a3OIWMfy7Qla2htS8OsaeFmjrm
PrXydOLsfQ7HbfQQDRhicjOsYY65QPvtj4MHL55yxCQkQFxHFudl4+zJ50kYSb8A/Jow8XcMENRQ
cI7bMxduxUoTtI7JG40qMUvA71F+HNuujNXpPu7DF4GBOgsldi2tMzAEo9++tnDir4ovYG0F+xwr
imz6ttNFGjd5OYTta82jICrtCAmlaNjR+oY64mD9g2lQ5sQJ2ZMuPqKdldSLxR3VfIpa9OJTtlU5
nDNA1tmefA+6sJFVQappeA1sKX9dJDQZYNWk5iq3EUIBRpa1PYkTyHpuudnZWNrOgdpezRtVQXPb
S/fXeLpnFceUp0JviXh9OWEo1CC6mwMbWcZ1tCsR1/EiMUX30NwMMT2nmvV6FENmKP4+vYb/MUom
eOxct7JEkULBbs4j1W4plIHfNf8rWe4kzZ19rnZlqrSDMi8XbO+uPqz72Z4DfnDbeFCsQQrRJ4Hh
yLGgfCKOUbsTFuKpUJd2NyI2G+3SR2vb0PJrAoCIkwUcmp6cNFd+bW+gL7sh1WFOVT1QNbevCvNG
NL5j1jQAiHBnWlYikBWBr/KmYDfHX9El3AuOZRtKFYassSd7MI6w/9WxpMGWWsWc2kyh6pmgVy9h
F6+BxANLXCkcH22kOnMToQnJGztQxx17evyfRVnxF+3gpHCRFOc9QYzIrNcRZzJJUqZRX6ydC/fG
sSWzmjkWSYSmNHRrmjqIcDDKw7qzKz3SZeykCI3PH25pL15xoOYB0sEDLHzFvwucD43T3KhwnUfa
PkQ/Zhdff4S1q6O2B5W1y1sGi1sTd7oCCLSJMqVFde4UxDnrm7BSbRxWssPmS426EU3IQuBsjbHg
WG6n1sKank3+zAoOJYrXqyMAjo/k2VGcCg1KcA5aVMeYmiTUgC/DIIOrPs3T5inglcCxzxDXp0LU
ZNcrnNOYc8HD1+I/DejFvQr6m7MPT84Gw9ke20XWPbx8ynRG7CQKCdzAu3nUnly/GsVoyd1ZUdsh
JZ/+PXaEy1NVDWEinFxWwfXajxbJYfwwlXEdODQyiwl9BwSqlPXjafxvBcoAzJ9flpLYWhwAEuik
IigzD6zLMgH74dSdbrHk8Ggm2CAG399sE6czLDV3hICjUSD2vtxku85Ll4A+ySGIukx/xX2eY0UA
VRV4eBDQwppphsqFTrYTtMCl9NiZ79XDC/XNIxH8VnSJG4SC20jkCTk20Rahr5XOyQ8fz4gbAfw8
sHFVFHPC4OI1xcqJN4vtP7yguAOAPe0yWMQD4OrizhW6eC7V9Fx5P0sK/pf2rWZgnsZc91nA4j6i
3RJa74euaYAPkKSvlPofXzTLUuFMCxko4s1CrbgVW9FU5dZq8evqRxiNlO8/Bo87t83bmdma1nTb
IvMqtpo7nEx3hwK1BWQLHscB6W/bTpXrFEmKSb3gKBdEMe/yxB24iEEnXpByP9298K38s8EMasUs
2aBRW3dOXJlWcH4beJ/ziri7X7BgaOV97smWH10lxv2KjYbGx+yCYDQGkBF50oG4/g5N5h/INAlP
NSPoIz5lYPJu5fy8ABexjpkDZuNauDakDt/V6sEwXTXNG2Qm0HosxwEbDT6s26z1uZWrU6MZmdcY
BUWgS15O0pG5JmFlNlq1fvfiiLo9jK07gD67cFNjVMWzsMsiq1M8ywiI3B4InIbrasT1k4QxNqVy
F0VyI9wtUE+N8T7XNMT/d/wELzhUJMs6F36vNpwvayltiXy28uoa3hZ+f/jmBIEeG3J7AdCPhO/G
YlXe2vutW3Q/cyNRZeuG18p5uyX3znVaKYesRXmll2VtQF1I8AP+TuUeBVCqvITIRaEF6vZ95kVD
jEkGAxqYJ3H5KJAoVae4z8QcauvBmCJrtgwprjuux+BGlUzrCBWmMt9z16A3isnCJslPJp8Zrc2+
sgW7Q3DPhEXosA5FwsjHwuy7wCB+7lP1jpQb/CkueQIo/EnCUmvY7U7SJIUMSS+lLcLN9gn+ShjV
KpulReMbpmOUpGBpOtVfcaHBFod9z94ddUp4uCAWsRkUZ6tJEt32FUevw6eoIc1GhPSBaM7fBxhX
SUJsXvdfU9sZ7AVjhEQZEwGZUoYd/tt85qHiu1nULiRjVOrbTQZL3+aAWmrD3x6rNNMNF+vjebJl
ds+31oO1SOp4CtF69YbXtBgzwrFeg0mf+R+mRqbpPQniWTk4hDLX7yCdm/FQKBHtVB6GOh1fXd9V
urNsoNWWg9VHgx0OChlO3abOhFrIA4Oxf8/0ESF5ew6lgWBWxB/Brvj6Md5DMS9WQVNcMHwoUWki
p+nspqlXECWlyOYVttxmYe+O+5U4hrMMq35u51SVoYqE0S76Dwj75AogUnnkJlPPXt0cMrHuvLeQ
462AHpodmeQvOQuCtCi6fLOgfOB/BHIRTlw62IHvlTURv97j02yoLucdgmSRhx1ktZn45gfYvtx6
pnMaiqTxvKlBEt/+725VNsaoVW3K6j28nxNVDh4Pudz0tKxjxsDhYaPsWamLy8Za9wUZxWp9B+iD
d1zZ2isI4doNA0Y/D0LFr+vHp2v8mbNZ/5d+qo2vY0yNic7Da7am9UMkBBQ1Y8OT6H5VssQrlVu4
A96C4U+Tw/NHtrRAgOIJ5LNq77sAZpTVkSG9GCXrHIjBHRYggwz8aXLt8mR5akDXSHWGnnnSP5Ds
quSZI7eoKkKjFj2KbXpfZMi7mvVKoHSd8lccA4ZYeHw0V4PN0w9N0JsKNtpnnBbaPWVbieHX7h+r
cNaMcuVG521fc10KmZt9X5mPuUQvAwiQI/mlFMKPlYEm71x4Hk93Syqeqir64+gUTNSOeyQoPlg/
sc1RETaeu0V2FUTf4EecXX3UGg8c8a6Yh4DbwKrztSBZpgwrmTIWVVVKeyc6ScnIf7WjSoelqJic
CqITEYKyJyLFVkXTa/dgUfTmnJ9xADCr/Rgc3R4hETzz2819oP4G5p7Hhah6r+ovtXibF/bfMJvT
BFFBaOFbGjk+7H/Zdu0aSxot6LY/3rKYbfRK7GMPuAjFNokoIcY2Btu/iwQdlZSMznPcZyDtS4Sl
PBEf6zqCW17F4QDTFKgBsx38EMcRWDLf3sy7vOzqvBO4KgsQ7k4pJUSMglsqgrKiCdB2fK21uWd4
lcHPqtrn7RNdX4lows5sylKgu+vtEpuXCC/k/L6GW3Q3yxqtZs9WlQ3zA9yWhjKyUFSrSc+BlIvv
dmbIIDZsbMyPHKwEhwZVEE2DxQ7mpk3CIQ0824zEH3D7jcZAOk3BCidFzDVCR8irPqD1HCzjFsfC
UOZW4QFg34JVaVycm5VSoMUqVrYKIHDw4Ox/XvkFbqoqPu2JvaC11pQHRYgx4bcB+YtU99C6GAeA
jxjDCk4l44vNJGAHR5wNmfUfjCBTY17BckZ0MdwjxvFq1WhDvzfef0niZRlwugJyr9TFZlkPYHPp
+J7iXnopmd2CSvGV9d0qju0uURuHctIdF/IxyDevRq3XmBMf6vpAJOqIpRImaFned9AV0yvFeHv9
bNVqkkjBi3JCS0VWHng0BWP2q6Yvzd/t++hiGLAQvt/iLJeLvlTetEnZHby/I00D6HmMPN61faED
RJL44nXfyNMsbEi20kdvRJjve9HTR0x4H4g3ecfSN/GHOvehzoH2dCwka32EdDOnb7PkVMUZi1kA
quRxsquK9KXFapEPbkb59E2wsaRPPFRpMODZXHP5FLFcoy/DOPoBg++JdU3R9gnWJJ/i32UcRySY
LWZzOOsv0liexLLF/aIy6FwraGhFzOPYQ5KXTLr1pbXgdX+CVEmqkJwMcEo3Ct4D1OOLcQGAwaTX
eO1PbLGqPwbWVKgsCHC60qrVqk0waxRj3WyVp+RuePWFgnXRJ8mTOoBZiXrMvQbCwMGteJGQ/Bqa
YeLQhghB3LlNPZXr5ECHsi9+tEwZoGOksnZe6l9HUOGDfaMedFbksMZK3dostXcY/E9UQcBKFk+U
Cp6llbn0hfF4JwEjNyCVjAD40VOOWnDf+H3wU/eWGtDiaN0v9k9eTjwuCk+cuptg4hE3ch8J+3gQ
VGPLqXj3CIqQpYcWa9isrHjCIWX7F7RyQ1eEWboq2jqbUnuEIoz+IbFgFy6O4q6xinBPP+/MWITC
bcC0dHhPYc2tyhO55M2bdNJtBd1LvUPJG9FnLpZ2zqMg8cQFkpl5nBc3OAuk9YrwXSFTREoaGbRv
oYYOryneBeg+bziCuA8ZDaEbUim6L+ML0lHMllqZlTrJ/7Klaj8OMp6KIcLG9ItDxey9xV8luvwX
C+3oWE4Tcom1AmJkPOZRmTJl69IFshAYPoF7z6NwWnZWDYrnHzolTxKtDOhUU0SNb4Y5QQtOHo3R
R96zhs++UlZxSrG/gcqAjYZr6omNgh+mvOJm5WwDs/a3SvTYTTAFesyvjLcRLP1yhX1i5XXTPyge
5VkHOkOCM6pA/xLIOoZ1pN6xxGXcVWrvavzzVakeupvY/eOcHumKRdozm6kWEmbC62GNPDWv129F
a/h8kb0J1hKWtQizgWkI0BG5F865A/GF8JZZ3AthyK6Tqfec+ucqQtE8TiL9Udfj30uG0ftShgOt
H5q29phYG4bdHt6WJVkjaiAUrHVUTKtp3zbvyMRVul5CXyRHSTVa+FGt17Pn9fVHmm8+mqV7bN7T
B74IlOknYZbDTft1P4gE1wo4Y8RC4hldfCQP/nhGcBaFvVwpiWNQEbLX9XPg8lS4YllprbXe5r0d
feLQoPN65DY38JJFNgBY/a299sTg3q+Lpjs2azIbcGDalP05uM20O5rtqQLNvYeKbe8HHLOZkAqh
DqH0GzM1uzr4iWAop6hsVpupssNnSjwLEsTIRgWNXX4GHuFQu14GwLpTQ6vSC1uyusB0fQoF8wmm
XpybCS3ws+24lz+IW+l4gRFdqckJsCJwk7TL3gJHAMZfCqZrIySt9MyktEWvscGSoR/TlQAtD1UR
Gq/MlpjUc7xN+jvExD0istRI14csmV4zeotfZ4ZA2+7O9SR7zNZHqmheYgC7HtDLiQwk7m8f+261
0IfyrDlyMggRtGCh5XTVScpt23Hv45+VGqAJUFrC9Lfun+UCErLEF05Cx9BpNGOsjI0xpVgYD1Sh
dMvWFpIA2zpR3nXN4zuIKWju7Qt6LzW9VcIGanbZq3cHophnwTZLXKwXl4eulIvq8++wJ1gpI1/p
RbH9yiJ98MAsmMuNzQe7qjIQzqlFkqlJyMiQKYoGqIBsycJzCfQmc/+su6qI7zRMLHSc4oQv+AYI
ivfrFzyVu5C7NrXamYNYcxpobnc30rbvIAAUnHk0owSxa6mi0X1jDUN4sdX2HTUhDtqFi4of9YtM
ZylYf2AVkzHyH1RZRWVNqD86/DBnwTN4qB8h3/40MYKyEAPsBZf11+uihijcnkdU5b/50tZrY8yq
swIl/0ABSlUGT97yxNd9hdNoz0EtclEXK+0joTDCJeKNYxFIvefmfSlXKPqOOt4qQvUfC6xpkeDA
yoH4DLhS5J+PztxVa6nSTc8r7AqVRe6MNIL0ljwYnjvNmck6dS1h8GTRcrj7PwxJZVfsbl9AjnFM
Pug6TmLDFZen/xO5UHvi8SIFAihKjkEt1alDLF12LUVkftu2VrdILZ5Hf5KaLFCvVsxj71zDPpO+
NNMeF2hLHOFfjKKnF4Q6Gzbq0ZArWaBYJkHft2QZFOgynlBcFh+Wgt9ceRVBQC6fxxAmlaxRyz/r
QOl91c9lmDT9R6eE08Mh3ettGHWSWDXkOXQgY1mk39iKuPso3EKIzsT+ZTZcr2bbSgc0aj/3Dk5u
qSlkQhLHAYR2C+BhCgZW7FIVcNex9AJmS/b6eEJPmqG5tGMohPAc8+z98QqivxNyqr94rOOvDbbs
dXVWWzHuv0qTwBoiwH3tPRGjzj18LXFpXTIFmzj6uUYI1BMMG7tZcp4Jb/cO4bbj+CFAd3ADGXQd
e339yVW3KXe+QbyKTDDelZHVlOfxYWpMPMpvhpPrXMNRjAJ6lW6ZssYLEwR7t/LjPXip9jX97vuZ
KcxE3QNtxNTBk8sA8nA8oJj8UCelrWK1StnFovET79DAbmvSINPtZPZ/nzqUCpFjHzbUKpYW5sWy
6bOHzF33zblFcGgiNglPVgcQQO3xtrA4GvO183CtaA1FoIGVSYqg99bfQ+26TTmxP0CMnmQFo8vs
RZ4KgUQ/y1orcWb8xGXmu0mUEdrZGTdQweN7JOBeuwZ1l+miHUUcmGO2vio5EnDE/NYQneTTeDNJ
D56ERc/EprkrL0ukUwBuoU71uKgO0ENas98prZhR3ZtrLTUlBjKVKblpLdoueh7dIrmV8Goc883/
8YnxQXmrNLpt+QrVm82uJKYV4d/9ENbwWiVMbnQrQPSF8vfwE4fwT9SfAU79q/S9aPdnf/3aFn6u
htR1OwLyvCYElX2AvUNVA36Pm+/j8o5K4RCCYJwx/TM9do8tznXGEuEh8JGPHm784q05ulkwmEOA
53JRxVgQ15EmrL+alkM0LvQji+1FV1eoH95BcBk0hfojyf2GkWYqLINxFE7Tq6ZqRhNxQxB7CsYi
5/mXFPAj8E5T7pCzbg2rfwdPh4nTTuvC+W1gwACxsenpomdMEfOTaOCo2Uhp12rgnvUkZqUuCphq
0EFv15PKi7ZUPKqFqxtLWpHdWur8vdlfEr+d+WLixroOHV2QSuY2KBU57xeB3bQHihep384LfCwb
meK/9c7iSJd6PNLdbNQzu8wU6lq2Om2QCDB1wARcnF4lxM3qWNFG3/yRela/4XzoU7BsgyeSx16a
VESN/fceFiv9kxzQi/QdbEihDw4fWaHv/2N1lbT16L4Pmm+5GX/5D6AsPlw7t96N85ck4PpalnzW
MAXxgh44jmrIMXzuss83GZNk2/puD+JLprufyNeK+kS0H23DqNKqA2PZ839f+Wz8IxmHwsksyN9e
fI0F0XnA9Nh8lmNt8yFejaeAfF8V7e/ToV9yZ3kK0lwbpaodu9z597Pui/3kMw9DBy0MU+YZl9Zy
1gFJpCYIluyquwXPYinuzsdCUvWEP37xbhnYlAxPsGSZRXhO5nglJMCP95G1LtJSbKIQRQmzk6dt
9MfB3aA6fwvjtflEMuy42OSs5U41rF1FVak9i8DfEbq4pkGRrp5p+jW4FHS0w4J1ZtxtKWlbPerW
W9ZGh5yUZW4aX8dnClUWn/reRFS8/EWGAp3uHcoHX0fF2rdKd0stFFEwjPCgWDf46TJOSRd7Wic8
V0YxH8SUjSmgIs331hJafTxjv3zC/C1LtWb4rjPrJ7mmIXFLZNO1yBF7dBXfHH77+BV8fsOPZfkZ
8maiG7IstkVlGfwhAoDfFnzvZCoXG7UFEIwwoROgV1NvNALkKFeDc+/icpke2PR4FS6WmATY4fEt
u9++GTDNDHic/K4W+DzbcNiUsTha0C0h4dcYEMRXaBsRasn4RARM0oBdXpOt+6vG8RwwgnmDcrbz
S9GYXGFfVA8o+ov1sI4dl9pShwAp1RS3gMvy38EHPLKK+BgFqM1nW/N/PH9FNr5v5YCJRQhIUzcb
2yINHmjswL69s1B8tAKenwIILQSl4FNAa7jOlxUtkpMqpTFmJ2JXDiRrIqSQjeg7LIxX6s+Zcn+w
3KC3Q6WA6qDZJjnU66fn+sIH1pWX5DEBwFApW3LZcKT86BJx7Y7PhxtvaOBH6hiTu2EnWRE4QNLc
pS4Jjkb9CoGnT3FqHHbpuP0BY/6+QRQUTKOHksv40VRWSwCiAxQR99N86Z/52lRHAcGIFlB73VDA
RbM6G3vyEo8gjpek2XCO6SXW6Khn8uiNnInCpavwNxkmXN8ZqfksRCm97xfwThttvjMCqY/hcby4
eMUc55Z9qmqNTqXi6Sbdxoc4eGpAaxayDJMUnx6N6iHmIsDZb65TjVhchrPXv9IqDM5EzZr4698c
qVaXaovsDFFlzsDgEyv1eslpzcezRtRZlZjIyZCpFfBvl1WxPQXM8yH4FKkkIEpvaFmLTA5BZi42
7+oifSEiorUqU5nvJjx8+kGh2YqRfAUhNhb11da7crW79QTjAVkJek8NSQWDrY6qvXlflHOay918
OdRRKjYZDVwMYjPWRlkLZOJJKhdEE0eWOzatxMvtAPlSvQIt6af/RGvTUu2cr7i8vgz16LspMfLh
0NM/wwIDg7zRanTmolukMz63chRM4o9mAznj7fU58trn/WBsMnN/9M/bauyyydr1BeZSe2gjoutZ
VaYxdZaSHW+HmYIETRI9CFcQICPwe1He2V91ezVZ5x9MjZS+jqaDMbl7pL5hAi+3gZ++EUqYLwTN
GKnC1XoggPbA5JyE0YWOoXT5V3Yd/uhnZ+QohkzfYcIUYj1YC0679kgbYkw1fJCwiYgoUsAsCuRw
LgjNF0w+drGt73uCoFiniDXjPM/V5/RLTbfVRVCY3ycKaj0e7SCScPvF9/2oPVZ4OV36Jqo3GCnw
eS5ylHpxHdHzbpeeR++vzrTV9h4YLPqVqBs7RGMrtU7sujh9G6Etbhy9wk86nK2I96GZzexKrQju
hnWaX/5ehXv59/dH89Dzgjccukf1yhEnTTbbjyMXW2R91C7ONaETvfxabbGQCY1Q1kL7LOS8U/3s
OExJxrnJOyuQmsLXXo6IfTzIgHxD6fLF7JrgFZX6uVbF4B1UE5pEPoI+sj8z2Tp3XQXzr6nvxQ8m
0llAAEsztt7PY0DY0KzH87l7G2/GsnPrcSextVMATtTkaraCoxwWoc1Ntom7/o8FhqWt9tthdsgu
Pd2gjEUi5yjoJiE2C2rTBYpN7u9F012z4qW4HdXTASfCMOICsLRL6TIhsi+zkx/qDSVRzKZu44nH
djlLSR41OUP3cQw6h3DU+P/R9olShqIEDnDmibd+iFpYvlZSbT9EMaaF1IJhwIpuzq7q+Brri+mA
xZsH9DqgswRZX8YoCKP/ZxWye1su0g6pESU98QdV/YFOKuqoFWjbtp2elKqoUHv/AXMFPN7tfJc4
QcqlLrhSe5ruvaIyLGIQAPSB3AM97dClr5L+VOUZRy183F7tLuUtNzKL/F5ACftTbrMeeCGcekix
U1Gb2ft50wBi66RV4fulpr0JFnjk6CqH0jDq0PA8st1y4zljh/ak9wHadrS36XinOm3axaz/gcDj
hQV4V2WCXafjz8FRX4aqHfa39/14LmoMwXl7/N5IAqKRJfQq8+MzmvHa1pnRDl2fkfXp1CxJ9x25
svkkttONHKp7CC+vHWKCcm55IFwvKb48oMQCbdHJUcOq5pWWYFTffSqZzDS8K/uFqu5POHN8PpMY
x1kQ5neySBOy9Cgy9f3mYmBa6Wb87fhNphurNWe/+JR9wd5Lgf7Uezs3JZSuNEx9R9vsnZPBmB0M
iPyZeiq10mrk9De2eoFSiMo27vDfXkkMDpZznbhRvn6noR0pwXP25XrVOgyFCe7hN0nK1mfaDiV6
Xd7qExsU6h2k9VOkrf+VP3umUbuHfi8JAslUsfnsqPdc9uvt66i3kYyeHO34unbxkjyTu0vdu2Bi
y4DXreevZq6PETPI0oyrsOmLq2kho68I21mqVg3R60eWcNcVwwPgHD0vLB61kFLbI231jqxhB/pT
sOuBWDVUM1Hpe//490xoyQOtitGl5nlT4o37M5eIknh4zDBfD3z5fK1El+Cv9mJs4l5bXaEbBRcB
/OCu1b4qjt81HUZP8UaEq3OobVHP5SBTKoAz5xjcLmq07c7os7c3KgNEHmRZRhRc+NcuHVXLGdX0
uzerjLs7gFVZjHz3ApC0jQ8ZG7TYYIsLXp6BT3ZE0cLRchzmeGO+Y98m2zIc7p1/YqSCRVJBAP4k
er/wK+8rtlPA7ff2ktd5t9Ht45UTAcYR72fDAWn5wxF6DfYRHeCcjqgHt/pDs6lg+5i/zMTGRwRc
O64mgX+smOtQVvvq83/c6UPLxopZSy15zEpSWXV8/JFEWjY8Ggbb0NGWYLankIMNq32MMgUZTn2B
0j0urRruZM/5PO44FrPagUh1cLKsMX7wSizmuJAOoKe83e+8eYoE4lTcI8J3PwT0xAzuCTUR4WQ8
rSJdyDkYRBwqbuIR/Y+STyttr+0kkouj4V0P5oaR+c+i/0gbCc2NsagnC8/8w6fkWQR/0PIQSiHO
RWR5ZpcmH887TsB9+IKJgIV826601wdq5syfAWp5ZwxxUHoTnV6LjmjINQT0ghP1IKJbWHMY33yM
zsff2sVmwuI0CyP/qjxRlw/dy/drQR4x/sNSN+TEi/kkQewU4sUjNzy4Y9WFAj0Xzhh3MafeZMQm
Mj0CCLA4maP5n6DkRt7TJrLccUmBjywpo3WJRQRBQT8Ncz/H2AEDxrkP2tuUwB+FqxGANjJ2BAMi
N0XOZicvRHZmkpkI7FdCpeOlAKzwo/pBHkMylTopy5e7cE4gXyJhaHJ9scicx3O8TwwT/Yfle4As
h+f6PJ9YhsoEj44Jst6hfmKHCOU9KgSkCkerw/ImJTw1sfygwjsdAxi5g0Vm/zPo7fK0Lbz198UI
wlsjcayVuIctYlp1moiMSqIZTCbO4ZLKjoETcM4DA6q/ymlo+ZyCJ9Ec1jAqqn2/XIQnP0QQvafH
AmCeonNth3JztOYiDcI4Eq/k4D7SBfkTWkk0ZWXGSoOOOcjh3DNchSuZDUKqRaKsXxdSuH3JbqvX
ceGfR8bbmRWpHBnbjYpR4TJwAQYRrL2gsjWV1B0h910vxmdbtEWgIjX6C9jlmm+C61gw/5/kO4ij
R5aioltJev2UnixB7inwcXjhHdrgOw8EJEUfqvsG7CM1v8vEK7v3L3Dp7jp5398w7sRgKe66ORjd
TFxYvtFdJYFsBYAIv1tkQeD0ni124Iqksf/RZKOstxTL/oPeScSyeu2RP9HaxSCVfXlahYMNt22h
ZLk0F2Gnf1FUjxlYgd5gjoExDwJ9zrLhsxwu8VD5gqZOkFWnFZKfL/21T2oukx1oUQihn2pV/tRM
UTl8Yio40A61eqKtt23UssuOYpTKVRZA6S3YqrCVr/KBLgzh8AZRt+QD3MoQ0e/pBF4F81qq2p73
mUcsapJdVJ/XlVTpELCn+4CE/ZlJWrvrGcwtNMgOxf+K5/wpLu7a9JB4my2fcFhvispBUl2b+t6W
VvRqEiHoU402vX5u/xowo5vf4dZ606yoBQYrWT7Qn6gUnTiZfO10pVDQmrdXXeJ2tk9bt5T2A890
T/xT2UeAhg5uBEMRxS02webAdM0nZcCBo6MkXlYxDdSGI0hxxgY576J/bN9tz+ZaJYQdY79HwDAD
ijE4mHFdfaaii+TlsORmo5jpH1CNZPLiS7wSHSIUQeO6pmRGsvzFpd1BRpASngtXSHBaIerAcqVh
ZJZ/jP6sjk4b9xc5L+PnHzW32lUNVHIMPzXrPjkq10wSHGto7diK4CLfk0F6wNJHh9kxHPv1tJBr
jpIEiEkDpgSDitfyTVOrozt430wRqesg0AQIP3Qd5vRlHgfunXsRm3ilRVQsu+SnZSAiMC/N35uI
7T9RR6b8rdupjGsB+FtxGSH5V9OlPBz5k9yEeYfGisk18FXqguGA0ACPTFeLBYHosiL87mgAojvD
zSAry6/Tj2V9lRyAc68HDpNw0A/PrNyDVm16AVNCc44rlz5FGkQ++pigPVbUgoncMb7dHDCGnpZE
LVPdOXF9DswYRm5szz2l6t/jIkfsttui08vK2OLiBZmU17/EWzRsrAGZmda566yG8vW3dRIdXkWv
hyUq5lnm9WF3gI/nL5oXQ1P+xEouQETEFXLJw20s7ONQYm4Clbt2jQuu2BzS/89/Hgf6wf+EloGR
u5Jg4Awgo4ULgzU5eviEBEjat0Ca8pCt7P6Aks9jWXErvvRJSfDqiixFOL3crdWAolXYwE+QUx4B
wuKOzDpsxe3Q6Cz2khtBnvAxk9hMqBwb4q8MOumMJtctA4mOIib0Pc43mmLFwlt5pE9usK8u1XTB
eqCm6PAd4IANiZ1OMdGsiJtedbYUHMPRM+4C/AkeG5yxmF8Mv/or8clF6OK9Iuk/H9glyt35zDxn
NmidODvEejqXnWAkuRN7Raocit6qD7s/+9nknTkGNE9MwUobq0EnUOLvNHJ/Zxy8RKDZ74dlylq1
/+SWQ+SK1Q7DLxk1j2A6C1Bhxf76XQezWDyKIiLw5JwsLyJnS2A0A+TbD9kMWGCUcQ9arE31455L
vO6X+YMTlgCOWZ/sng1yEzWa455hBqhYouVFVsjhPfSVG+2J6AHswREbY9g1OTRc7QNnvwaUQXdm
MH3rz3l/Bj5YzRd5zWWq4nO+1qbpA/d9SGDOIYUpg3gEoDCVWVz6EUbxaGN08Go9x95MxY2JRmlm
/4KR5HFm2PAD1Iy5b6FqPIKIc4m8DV6iA/zcFvJnzbZrI0ECs0NUcWoxima+OvMpElLFTZkFz8oy
meSc9kZ26HMkGDl1bpOzR86imXcRmBhd811k7KnD+ZWaGJdfqwjXmURYA2PQI9pXY9YEFOPcqM3R
qEmo5FSBUpG/mO1cK3YVJ+hz4oxd9RlSrmY890PxELjF04pRI4NLVcWBO091NnoAZXCb46hvva86
ZiJb4vUZ2tyybg4WF8PC+IPA6POQE5wYSS332n3N0TMioPAv+pMzvKgmdVDMFuvU9feZfvkqxkgw
WVRcpmtUYCJWT8TObHPuVExSzz0i5uMI4FtWP8NKf62Q2pu32N1zkYT9cdahUcxzrv7DY3YdkWuv
0eSyXAXEwwHO/DShAH0kC11i2RNVPCXL/5JIyABnAJX5O1TBVWVo1IBLZ/2hZ/6wSsUXR/JB0gMA
MxSbpEpEz3nER/NPdiyDO4Wm1se/isAz6mPUPClvQxnkIAiUF9LQu/C9wG2S5E9cFHUC3ZHXt6Jt
rjbcaWH3GXPfWXhK3DS6/8yywhgUupJb0xM8I/6SOMngPrKup7A9hO7YMtuVPRHkRufn4Kk6q9WP
sVje7M+dky2326J1+qWUxGsPDv2A3XIIMJi1Vj6PYupySBxZawGmgwGktWMM021oD006titGpFwi
PnaQ5RhYdFgGT6RyUkDKseKYy3dCjWIgrweczqEnmAT05llZ7eallnrQ7YqeUORl9kKhbHZzzBx9
8AnVABANQUKAau+a2Ik6Cl0k09toSGN/Mml9EZFl1LylKxx86U+AGz9iLcKIxvuwpGRDKomwH4Rk
6RPsYUlp/JAhr+43Ug5WuavRzVzSCYcjooC3G/pES4h2W6acapKpiog/jloVUw/nGVAxoAOpJuVt
CsLVLnIxgcfhk301TOyX8E4GgH4cCiIxeYiT3pvLtjVj/NfRWnLY4JDD+BsYIq1Ntn042CzAZe24
OCqeQdyHLDL9IhPeUG5jlV4QyVOaQ02wyfIyh//UX/mxYotaK3fHPKqDOM5+0a5kEovjeExhSwUQ
u9XyxYSLjPCI/jxVYJa5jbuDDjxHBh030o7irRY3AFTuno8yrv7OIZkfDYfR/4sjAkmnAZtrYZw+
g2I2OlzcYaSKNRXk4v1ELbdlhYp9IubNF/ht8eBmHJuyN7VOEqevVoQe6vGqgRMbhvy62V9WInNE
McOsCDjy96AlLiGISO3fGrcH5q56shl0gT+J2ZQRC+oCjo3GdoUjxw7INiVsL/AGuZB5P25IklHp
9y69IyQjMpL9bMdU91m/xMYp83p8xSPvPxeZ+zsKSziJEtggTYtS0cNC2IlnXSbxo9guMqh3wcNa
iREIrd/srT1yJYZfx+Lp5AxkQeCQc2Nu4jpoka4ItsSh0L3xi/w4B0jNOO30BQw/mYOV1DhzJMwL
5CDhX6ZDkiIltxt6FD/TvE30kxAmW+aG7aUruawoGnWbaKZ1zRqE8xMeg8tnAfgwxyKBk0UHeCjb
N4QfkcxKhC/ur5YGwrUqxu8gjSI7RHdA3H6l1urzYwztcG4J5YHkReX9fZqECWyPE/n7OE0aYsPu
x5mNMWnjEYCkAE3SJY2f2elNDw3kzoKxXolpxm10rXuJHcKr9BdcPLPrGkmU6KpXN2EWc74U/kRH
hCrLVRCEGL1nOAX6QlMK2+xMd1FeA7v853AvT8qm2TcB2mqQkyjEYCIGPECghOd1vq7SzbYiWDe5
+q3rJDz0Rrke9UtTV16ib0Zs0zfQeYSbHhYOswS1RYQ+fZKD5ozsaqDqq92+C1In9g12flMJGp96
2SVmjajaei89YXHTLsoNEsBn+pHRaS6N9Wb8zfZpQXwSJ8b2F/HE8JnyyPWd48WTmhXXoLCmq6e2
jB91E824o6uFkStoWZJHFSPn6Q/+z8x4Tpfl5oo5OMQXhU5ElUllagWLyRRLsSoWsbW+86PdqHe1
yAcRormd/LtNjXN6FgYDJ0dG5NOx4YO78EV4GnMBMjmwd5/5a67v8asr6lbf/8G5sy208U0KILIw
YiCQNUdLwqZ3aAC5mekymhGJJf7vVBwr6TQW9PEstBApcOD0tRm6mncAmgJNPOlooiL79yeo9Jwj
Mnwm0bjNMDUxCBHVCQ4gTw747g/Ce8gL4AY+MDaQCiHo/QremJOGyVR+KK6MV0ovSlMSORksNe5q
wrNaZFkPI/aGSH42zcce2SMrtS8pD247ebiuZkaEPchHUyCsmtymClEXdy9kZTFTbd8GRXAU8Y58
K3CnioOHr1VVhNz+V+TlKyOWR6jRzD4ZR0PcRak0hcbxBVB3fxFwnQn0gIe/RyuJ316BDKxbwHOk
lF+oybpBsuci2oviiJZwJuaUVuU2uqFrYWAZ28O/gPDlU2/mDcMTLtaXwYR3QC4tko8nRkL10Ltc
TNXnucgDLOl8NVr1smYtY9UzFHQpjkNZxobz6XPym6yiH4PgXqBu5jcTzHD5wJaIItWeFurS/w4O
rIIAaxqIrc4UqPlDoHOMMgeIhmLCPXrSAypu8cv8hFtM3Xlw7n2j1ynlPz+JMzgYCKVmI4liHtOz
hufLP6Wk04if5P3aXbItlt6wW3UuRUQso28s4BPNG8yS3n3urkSJOpDPXJWg9/4eN/LeWSTn9gQz
o7NpDTgqE4fmHahB4/TPZxMDQqTVrHTYzNmdrttffAQMXJRckDOVJYmpL20BYSvpi7dayVMqu8w7
XsxjX4vSSOsKTxKnuvbVNWJFbTuBXRB8StWFAPHttymTYZVfyCJGNWxVX3la7+zN1gDG8yGOM0Ij
L6vlhQEHtuYQZwm/BRXSXfy6mgFjy+Tdh4nlR2hDYpizqD74qrThyc8eOuqbt8zcYn/gRIAJTwvq
2MxxlL0JojkqQbjBQJS0Vn1gNYaD0PgHPX1/WwPpDigqmQAPK1oARtbQ+C3/UCz/1IM2oUKuQWzU
/M8+0baNWwIoWNNrYpw3EIGwtbWFG4gYEgDf8RgGsWuswbsY5XH/j+l74+h7pr4k4MFi9t/5m3Cj
BPs/c5vVH4CgmpUoBv3uU4aXanx2LEGuBr6u+bGWYYYoM9zyVh3wyVJtFUQ3QlMLQtHqh5tIHrJI
ncvd5yiPBNP92Bzt/I86GIVGwnfMi8Spg4XEh1c8WZlVjaLHZnf5ma/XQYfssGnXcv72rggNrSJM
Vyq437txkRRBhXri1kjjzvtAGgSf+uXE6A5b0QkHZIOjS420xVP2wVsnM5pEq4YYKHZJ7lWjcZOC
X1JOH30cRhuildxPiMjAC08BYATlp5vaThb6zTNx/gHrjQ7mIzKRIT5R4UOAvoiHi6l2xe+QXXdr
lWgPhFLzoNln6Bf90JVG65ltQ65lWX+MPuUdDj6Sd19uTR09BCI8dksNexUjHOIHPTKrr/2Ng63O
ERSLXF2V7bB96BAsmhNT2YZjXm8xSgbEEJ6Ribh68TmDJFbAD+K9362nVz1r+j8Hzo/zGKbBM0eL
KZ/c4oqfJldb/yEAE2CDf4yHTsszS+bEHroBEo2n7Yahd231oz61BDKoydYfKo+A5dNNztitRJIw
h7L7Dsse83RLdBizUEYQsncp97LGRCDY/Vi0O/gEvQDpW/056t5omFtizQgAM9QjXXrIpMX4QqXg
BR2B8MchM8x9Po7pRzVaKc5BN5tbv8YUtV0F4GWFCEju6uK6gFMy2SkI+GXFf5xe0ntf+WKDNCfK
zgHZT+PSv7fVcm4zvxyqnlssiO1hayAx/O7pIsx6/UxdTUPmx0aPEAY/w8Mj07FMZ901VbdINcYA
rNDdBcPc0cmFUfscxpmDUclddUqw28S/a/i8pWljbc92THS58XtHKWThC+io3ajuNnOK+tn16Q3O
ZR8HU/FU6SKnGc85aYIDjpNlvbrQIqmmGvRPPLLVmNZZjLIWVUh7GF0mul7ql4UmXotpHcSoNVXT
oK6TvIPaHL0nY2xuctpF7ox13KH0RuVUeRF18SRlc3PgEDhqFQhobZP+PC+Aasr9yMwyU7yFdc8c
PkIXBEdD8mZcgOzyguazzrgh/y67RjQbJeu/gghQFfsc8InF2oGRRrP8eq191MOtUtF7+jNqUGtL
2spgQhvqn9I6903/L2j+qUqoEDAyOgbMydYbbd67fMDNthPoGMgDzNUPNCw6QUVV1BxvpDtGM0tn
6yKYj0/l4jGu87q1HEAVt7jMxZP33vdvAtknkXeDADHGfUEqD15QQysuK3YItOJLI0GjBrlD3bbt
qsqOavdXoYXxNMXJIPRpSMkpJU4GIJcNEqZkbfbI1MKg1EkJ4TlDaygApDzULYRV/YnaOHrxdFiy
obLEPtZLM3GfcEQwEzh8lVXhlitqRgqnzdoF+ilAmqvZ9Z6BvX7GE22Rjbh6q5QfV1Z0Sj/OkLg+
WrwAjeIXQz9Q69h6EdEMN6JFFPs8Q0nH1r6cgMHG6lC0BhaQ73Pu3TyWIz/GjPRSfqaK6EExp4uZ
x9WjlMbWp5J8N/O0wOCVaLhKiTNvEjPOk1mhcIm+hhbA5LVk9iNSWyuUtPpDbOiO7OZjxtSg9xue
its2UMgTUtsURBjcpCxcCAt0pQyGuWA6lG+NjBzryuueBcmSG7pG0ljorZTy8n2TTvog2fd3Ps7G
yGtlnykVr6Rva8vNd21wZWcSrSkbxiLtfus2cy4VjCgeLpK65kfLBz8d3VLau25BC4xTyXRyrC3n
uLQBaIyM3I6SK0fbAxl00WPFXho1VT5FdGPYmoswqr7pn0SxVYrvFh7BUuk3EgNgBNvdLLMcfzWE
O8y+pp1UU1wJTkYc/QeWWZUUFSpw2+Ag4T1XR+T05RaqgZm3sbc3ZglYAmG2lE/xebRZGO5e6NHH
fbZa0c4c2eum7aWxGK4p6rI8DuwD2TDb4e711V+gh2eT6uUJuOuhDafpLQdxBgMnGrIo73Ub3Jbr
gajoZscz3mHe71hGM4GKfa5CxZvI1piKSXQT9r4PZVdAy08BoO7K1uw2XVeqwd/NGmXYWRSGHM31
VODPfn6TES+ODc9h6V0Vh2wxgbU2tuGABADKPFwvc8I6ez3vq9HTwkWjFgh+CaGqvNf1t+ra090j
5yZlHGaGEpDa5qQrFOXfhMjRJgfdNDpDoVzqHZIMR4H+GxhPe7/uHRML5us8NLOlbDRekfGUDucv
HemOrCNkxzZuyIFpzFeWXzOip9thvBN1DATw/nPYEnXpUG8vUMIS85DNVW7fhYV2mY7qkJqlncWj
rJGXjbYJen9TY/LCFVxBSfGFpg3JZNJlAcBiHPhj8wX+z2QOTfpRGiE/RyEVIbCjDZc+XFpIycVP
PfVXFbM0GkXdsbphhWox0sB90dEXnkKXVlhJuikVMR+deo8JV2obo3b0Qf9y4GeE+rrEM1bi8Bs0
i3tL+y2swrKf/wm+jQH7dTZQD95ILzPyLdYze9+SV2zp6fcniE9KBnCsnwrdZPwS045MiVa2qvP1
w/SezjbiwYF7cDLJ7cRLe+1Zd9rDPZXtSu6mRqkCQPInIY5blA316PBz6mJTTIQ5THFGUGaymxU7
yAS8IhZtYax/NMLurxpFVvoGTnh3fbDZginV/rtnHkgSt7QVqQDIfAH8P3l0Eukx+JdLZiXquHq4
fU/ShxVVSsYYzrNzQvf1mGVlq0h6G80eNZmANQ1AXsRPYvSdG9PoLy6H8MuYXozjzFDXGnXQj9Ln
SKj8YKlAkRR98SRkTX44TaWo1RzKOu5owmrM9jUmLh6xvOksLlvL31AcTv/ZXhEWJ0c/yLRgMvIv
KQR0sxEctGQFsQ4QpV9AqM6n+FysSKg1detqfSltV3tv66FPV2hA3anajwgB2bMPNR5fRM4E3JiF
8wlh5RuMVlG6rUkJFNOynPCDnyYioyTa/bFGJC8zFaH32AB9iIMXALRu5gbS8fa92QK/FNyDhct3
DRyLgqUV5s3T0d4mOa6Ywcy0NxHKLtReHImMCGhjCJybjjAlgBkn1peuFDW5qG1Kh14E9cBEqimJ
P7aj4r3hR6YGG3xYRxuBq/+Y8jw+G8zXL+GBC2fegcNhFEu4RY53GgQG7BkSr5rET+HuQBc0xg12
+HJpbfBnOae5luK5txq65krKiSQ1J1DshUwoCXCeDXKJ1028cZg+kMv4Uo825611odJ+3KXhltoW
in+Ca8zf3WSzYKpDGsCQ/rz7aHsvYmldVJQGOi85bNZdVaBrIBqvW37qIu8jDlPyhRIeNCVEPebi
1E1csfXA69r99eiLA9ALRylzI/y+aQ9zrAnki9jXqwrxbdzVgeUMnbRRAQ4XfKjJx1Y3ACEIvl2i
pBZQrOjfrXLygyg1c5fiwtVfO/2VaYUPHLEq8Fkm3xUV0u62t7uPoyolmfZt64XqOsfkvLP34zVb
IAfmEgTP2bcR52HU5hqJ8gLtF1YgaM8nQVDsWdYAz397VkpiyJpNHZZG5JLEibFcaMKJlOPeArRc
nDpyXwxgN3kKypjtltda9E3WSS6Cro+rTHLVpeZNz/H/8/36vhPQMUPX4mAcMf5/8q79VMCKq55/
wvGb8z76og/laABOuJIm1/pC+9nfl8QUst8kxO15Qy+NAjLNawmn3UmzdrLBLIVfVK8NBHbcN7r/
tYbOWgqQHVbdewW+MkxIxSVT8sTlve0WMSfY2o+xifhVPOjjrSFYuEuAbDuvRBAH+frJv7T/FC+E
0XYF/PCRSXcOFgLHnstUp/mkcG6DQqrqu8iIimGI4ZF/M6IY3DrWFZHMg9LNlkIUZBCC7vYFilgZ
6JFzFiC7NYF3OD/Q7JW65oxY4tcK8coRWsTZlKEPK/MofTglqBk055vDaPWW1RwvxGYL1rDxBJEa
JcRQ6f6Ix5NygUU4hYjCHuR/mkgvacMXm+SNVoiTeATZuLQ/yz/TV+d5s6rRVJ4B/05cdOyff0dW
DzVxZ1/KbjReDGxAH7UE/P8ffZdE9Nx0vnu8xE1nb73OLuOYAnLoKXq1/N/en95IcDziqvMr9A9y
/7Eqm2+wW4qu7qhP5hD/jXBjcVLDJCS09a/dZmrL4xxyw4EUj5YKxjwd3ATofCUoguXtXk8ClFNZ
uo5JREsuddBL1PVwWitUMRKzTYmCkREIs0ypeDQNkYrz2XrX2x8HiwEaM2mpLmGG7HZ04TfvmDvs
8YXT9VLGGYRviSc5WLWM7Lxi+ECrDZDhdTNX7CwwHbfQqsqd51psynPZmtKu3oSNPLMa+fp/kMQ/
wnpnhQs+YxCCYpIFP69m91lZJ1inZuTPjZgwozdvTuowqjoh5HZt9Cfhct2MLDlM+ycjnUMfAx6L
ATXhA1DkJH1GYsyPHDqym2G1lqoFDBWjV26tyCYWc7F6pGoz7EZVc/N8LSI9HzjbAWSMoS57nhdM
HKN6rHKY22Ayj6qwgyfLV/p+U/6ju8uG3sOdLz+CNm6U+n+JqQOcsoBXMvrJKbBK577EOR1gS1tM
Q10J4Jcy28gflvV6gQHOp0CxQS2zcIlF5QuKLNCwFzmmE7P4jFEmsuIyUX3wBD1QGRPrS2AFCDns
Bpc5pJ27A3ZY1vVCiHVBXXWV4NMl74VtOIrs+C8qeaWZIjdEJVcPXOMH/gfk5Rh+8yVikqn3NlJW
J4xsOgFNwPorqA7y4GXKYMGVjONYxigr7hIoya3n8MCmcoGZyhxIfLKq9XQEUzmSUvEQUaP4mDSU
Ki3DQftVGaDSAC7FWj1wRQvdZBXTz5IUQJF5/P2N0ADvfVlpxVVjzdkdx0nYuFtAMpgacXqWs7oR
9PXv6H8KAMuwzyIV+nnFmxKToQy/NCrhaJunxlFNFSKIH23TDRmbHrTevT5g5HVbrHV/9zD3eqeA
U3Sdu+/3Ty3CSv2I8wXxpFgTy4lkWdmyyPH5GzlwYY73RZ35TmY+FpZ3Jset8kCbkT4LyGrdVc41
W9mHe4VkgDibgdjVRsTpuP3WKJewdihR2/CY37SA4R0gmtYdZ5Z5hJPFkDrAKGIuLDqFWxOeZZsj
C/S31yb2uGUgxWSb3i7TrfFRKRpt/yphbUC89Nfyi5cvycidymdFiy6hXrGmYC+NBfVz8pOiK7Rp
brZPUMGIchlOpUNCWIDRAlb4MaTQzU5fpvnDWOolJc1VjUECkxhyObEGKI56cj8cI7gT3/6Wb4js
wgg56Y5JjY5rxbOlj914ftaVkIdCMv/ESNLcw4b0AyurpC0B4GuRsc0s7jYon9bKjQ+VYYbRlDk9
cn0JefFZhjLqKDylIrefhCj5TItweSWl7QgN56yQAevFZJ78Ia0LW1aC7PavWvKkqKcoIlvFeVWF
KdlmEWZJ69zmLh9vJ3xD4HhWSe8jO5QpGPlu0Uz7Gesvvd85KhE6twWE5q9hppRqIaeYQa/92dJx
gfrH0EwYuPsxo9fu25HsQbXExQn2Yg2M3aFzRGOQ7N4XZJ6NfeWjzW0peMBRCUgxbXsQ34Jj01+s
lcRBGIU0iygrMbPyNPK9+WfT9rFWII0PzLzZn4bR0KMfR5bUUSJleJ6u6zLIIS49BQobD3X2gzYL
zpOto3VjopsSd73xaAQ5avrMidDQu6m9WRZOdQGdPWYazMYYthoBLPSdppek9Ilp0jMMbhcDqCZl
4DFY6fexcqe0BSvOXBp9HAZSGPYkr9HocEMN1dvrUyI8oj3c8LTPIk2ff4+5qVc9YayjYkz2gOHj
rcJ18DjeINwKR/mHxDi2rk1hv0eR6xEKwsBgc+MKOc6boPnZVoLeUlTE3prxoY5IBroJtbkokTro
WHFW4xPWiGlQlKgUEZ59KadZx+rSMO/F7+Vu3AVxKGuvla7SM+wdRLUBM/hPxCAssJh6xRB+0euQ
gHDHPmyt94BN2mpERrrczCZV6oHVkcSY3e5j/lt8vs4PLYZNCvldx0cxJlnBVng9HFN3INS2V2PS
ZS2UhxrUxZ0G6Li3e4cAajLU7nbCsiqCyb8dWtRVuJfzsCSqxIKRSWsMoz7g5w8wtMfsAixIhIVb
OLs4Ykc/kTk81S5tn7lDs4u5B5gYG4OGM6eXezq8hzbu/tOAUEJdGTSDMCCzHfyOTmDh6BoFNjyn
IZmuNROaaHsD3yMYd4va62abVL2rf8zSxsddc35tln3GVgt77mv/ZEQTfqYGOjoIuX76nAqAqzA/
XwDsRcRxpixwE23auezJvdJxNAvws9Tf4ps58+uIhWyk1mC4aG94n9KmfWvNchCdYNRzJ6u3OLTQ
2G+hFz/ttRkRbl/GbFi76MCnjgSUqwo451MzqNIQghocRyvpqdyZVtmeAxW/yFI23SZCaK+8WFey
ftgxFNG+jOy+WVB/2D9R3qbjyubwy73HkJpe+wsfxUStHaqxbdt9KdTVKTI4bTQM27+ge4BMg3t8
FyeNcD1HiOPl9B5QsjwkYYolzDqoJA3owpwPX/KZyFeCAtGS2HSShr4sxL/JWyUpW8BOJ4bCERWm
T8zyH3tbYMJ6SNNOgjcDJJaltRPehjWshtiUhcMdUXi4a3DaB+3M+NlzYAtgfygyUhD39/9hiIar
qRp5r1depaw0uoRtaRgbrL6LlM9VcxXPYa+CPKDbfhNMkb98pT3+KR01zPAaMG3nn4LFB6uZvk0C
bBuExsv3RvPzmj0c0HgCcb1ABPJhgWsaQtyQtKy2c4CHXCs86+pGiO0AcCysUcme9Lqz8ds1sqBg
Nn+mHxZQE2Km7kHQJuv80gOtSIE0fJzILk+Gfq2ceeyDRDHuYsY8tqLcy4ScpugHVYTjBwhcM3Xo
NJ0sjPUrp/cl59gDs2dVWdqhZegEtr3ORP/h6mYZzKTR1Cc5bIRR8IiW/LcYDQlKKAqOfokcXDKZ
8MHXE2JZnc1BDuYw0JIXJt5l2jMFPcYu7wEdUThXF4ckJKsAWDvDQ5BrtYyKuryzCjdtB1MpeFFw
Cnnz7buspXOBDxPo7rY9hYlHAseN8JMqmXiV1dcgg3yJlIQT6Ghp1XcsyIhF0N1agDQ57b65iG7w
H5tklH5ZnSvnRwNLMHuPtvzG5JIvDml6PPmyhkk6BCIoI07ubVJE4PWsLV4Ac4ka3pzIIMVHZ7Kv
VM6EI17FKhD7k/H/Z78iRtjAKzTu6Wmupd/rCh/Kz2L6MsjAPZSNAZr2MtNNen3L6t99tk9H9rM2
FyptSS0bgsf+kiX+i6f2gsL+eyWk4+yX5T5Ey1gsp1eHLtj+as4u35oDL/24uwSHxlVNBY6ZieOG
t7vn6gg0zTk1bkNG7ikKiBHjWZb0xx8YMHNgumNkj2eJSEE4JMsy2JwDXNS+CI9LC5pzkCb0LuGL
PyfC3MdSH4p52X5MO4z3FeMTCzSdvPyPtsUYFPQN2H/y6kxni5VoPE5R6dz6E3bm8ZTYq6emI81a
D0dIPRtWHPQcJG+DgTUSGkc8lpmM0kDDw9ieSE5WhWyWg2Nn0wE3NImB9COv5nBYI8RJqPrOfKzN
K/CBewXJsV3NH4SdGr6hmROyHnLpivOjnkRri+i+3oSwYYsX3TuNxPv8aiaMm7ZuFXX5vA5fry9c
5O2fJUEBQmx7sNe6976SJg9HlSAsXmqizHcOMFQ0fKiW2XA3LmD4bL3AMvFCg+MbyCXSjeo14qVy
IHSTYoGQLQxybc3RFzeZUyVIDLRS3PU/uKzFizHPlE0vXIWgYwVwx3YG/PlLbWYzaz31V9VD3bk+
R+CycQMGd9AjAkiJPdBTEwKyAMtVYRHWpe7cWQ1a0/D5TpHy7yBXhjZYCjEZKvlc69AWY3VV4KQ/
K2p2RC2FLF67vS7wYG+GhtgJ9f7DFiWZTXJv2NonlYJeUgB10AdqboEFstGvDfPqrmhNB0lFdCCP
C2y4IXv7Z0ASqoB4SPiRQS+16gA+ZDTIdJKtBgs60BE8K0TTImhhC752uGBFQ8IB3iox9GhxQ+LS
5yhRQO5LeJ/n5Ra6DgO6MzinMse0LmXgOoQZ9KlHRSvjd3aylR51x6dx0pmfPYlk7p42mko4vSxN
FDHC7PQ9AuFOf1/4ZCYxFvldDnCDr/GkYX9fe8kQQsowf9CFdk3G8ImCj9XGVsmTIftKFp9JRe1d
eMQVioVM+YgZeIVjfILapBuorhEG11iggg6AIjdyWynOb9IF3g4Aq8mLSGpmGOvflSVGLQIf0HEr
OC4Zl+n92VLiYoisK6bZ/NfQBqy55UQ9yjI/kuDuamHDix/3ogDX9KB6KrdIbUjGTd/l1kYHXgen
wO7EavZRfvzarAEGhiFE1g9e5Q4TMrkgSd2Hs1uKeWC8CaqX/1aruDb9A8tHdV2bSalQtfavJ6qU
a86YM1UhqeLWF+akXafmn4zmQL0cSHKwZxb37m/w2w3RO/XboY+tRTdjf5H013UQhqrfG3OLij0+
1sRes5PVkySY2m3+w074djiyYGfGTddsDBwyp6PdtJXiSmNggZAkHinIOgVfm7+v52r7xyALy6n0
wE7B01Lwj5cqGkIczoM2LQFSopsx9NFbtnojNhEFDPu4gAisyV+OKzd+fe5OsO0Nzw37ShiIEU+3
LS2mxwrIU/oJJjJ7PrTjHTby2w3LQ9ImooSNHKKN3GAxnj4v0xbJ1Bmm+DnvZoHm/IO5iztljRkR
cp4jX+MXqRoMWB8yRhPKrS61wrrBgw06iF16t3JabIWgKwqi+3QSRJqavP5dJSBaC+ShZU223eus
KR75AtB3IiHEQmaQYL2V6/6KBNBKwR3l+0cwjiCjxxjzoorQw/s78SJ3HY5/0Dd/4/3xQCrOALtW
bNZRvtXiptBHQZXvjNUOmeigvr7WMG8bHrvEzeexriD6MD8Gr7WJBPKKELpjbhHU4IQL9OYhmS+m
paCPVODFymyzgDu3vfila934/kaqDrv0+ARlzARFZltdoRRIjJlS80MRjXwe+XjBVa3C18e0Cko5
qq/t1j+BO09cVEednaeXcZrISgf98ZziDnYm9MeDUx9SPFIlTeMxkZd/TGwb/0f2YTF2lH72ljho
Nz2zEbUzv2coWj0Ye8YvnYPSWu3av8vSguAprlS6jen2GhZU7QQ1UxTAY4k9/+qKUKf/CutJwUnt
42JhVG6ilLm+Obn8BasLj+NqU07Ybs6ldsQPXlI88FxAND7Qk4KXcBII22/uFGi+cx9RIReB2aZO
W6vcrxZtauj7GyFeStPFxl+yG7gnglLuObzeXsBZPNtnVvwB3mqwLaJ7hmdQkTqiHQlQ4MKBOW2u
em5OYE5SamfMznuw8lSN97ApYy4dxeyPdHJa+BLAQQE/KUlN4lmMLS3qPvoEnnafLGWqMhH6iI5b
C6wWvxepC/R8wyoJqC3n9yst2SP2Y16/c9BHcAwIj02ViEfAHuzfwBrtL8SaloN9PQyOYtHNACVa
w/WJH2UgV20IxzU6o0DVhVcN8+pyndBjayYhzTy1tl5UxAOpXP9+pPPNRv8cu2pEd0bGluwKeg0P
Y12EYacCsSUOwISa4kMJK3wjnli+H6GUKW7CFQhIp22tVM3UBsDVimbP4vNoBqa6L9lS+kV59Dhd
oSb8qsYYi8ZxQNbjdUU2nW9Z/dYEPku6bqrW0Ta0zHp0PpI5GuooftHvFLfskyAOVSMOoQkuZ5FB
s12dOL9u7X6WhkjSoNHT5vVhr0msBbsscpzl4Z4vVwmkjPI5X/yGVi+UVbeUpoFloggtH6qxclh9
Dbe+gQTXP5dgrZkIpj93hypC0nCVYavIcpYMqluHpwZUxGaBJDXezR5NSO77uLORxPGO3b9iEyy4
ssBgi//6NT3WC0qtVrfSXKvOcM1hf4AGS6hZbTLuuXK7u3ZGufLQewi/59Z/NWOjcIXJxbIvABEj
YnZl7zmcWK1rwfAkt/4oo3LNoN3kQ46YGBxfeCw9PZOc3WvREc/VA3F0UZjFMSpQqPKh4DzyAgr2
SxaPBgIYkCuGZYxU1WnDRh/JGjBCP/XfDyYBA4w2b/1aCPehNgMMahv7duSza/HyrYvogFPQuRoa
wNgVFxaINDTi213/AQXPQRejuJ9glv4vB3ofhKSrkgGKbPLqMpxlm9yWPkPtEeNEeD2xAfqLLXWZ
h7MCfB0TfQEKlolX6/Eu6v1Z/sSgJacleMLwbs7qA9oeKO80ahsrPnERtzORwx68nYB4kqarTREt
RRyRaqHKH6F4ewYI13xVcU/H9MEKFQC1drQinOrSy4+41eHwUx9WYUg0+du+xSt0ZnjYWIFxhYsi
yDKB+FUr1zdh5GSwUYp0FYPnJWHFNL8eMBOwKuH6jlYmXeX02vFOkOsYR8kZjAKHIh3DkmaEVyC7
VXPNr7eZw8kO86t4pir4ZfxFXyAPbSUiAux8EKZtap1XGHbXvEcYHVwj0d7zucdGfQOnRV2WLYEb
n7/ZKl0TbUe7NMx1zuzK21SvzuLAnyeyUEJTAUqAjLRnDoFLNleJBVCPZzn+MJC6q5RdwFjyO38s
zsx4KWP4x+8zhmfFyJvNCtmw1Y0d5k2HFPLyFWHdi6M52pqSsJULVS7EytTr4QhtELRBGQFM+tNz
z9V2Wf2Y9TcaTxzTcmpjbJEpvtCZ1qvCN+wmrWuB3owbsAA6DqbbCiaEzR7AFbyWo/+Y5iET3J0H
AA4qbT32R7+h8bf7bpnsN/pHn5FMcvNYAa76nXeJUQXbPH+5sS4K7lexaaaWtI+6LRbJ17OAZ+TT
KHvJdjqzuyCy+Ky6ZrtypGFDxNcYns0guYxc0FwoJD72ss+X3MZMTCxGMz8PyyUeKKsNFBvODDgV
xufGzFhn6nEIaVEr/kJpKdSrDFEt/W3kb/cBEHK/evVkhL7o4w6p7Iyp1Kri5tw8u48kgMcDkL/6
EhtOJvtk9fNwLnGeL2GZz8gSaG9N+yMoThqZ9NllEtrgvE2Vz3bJW1Uk9Xg+gl4bWPBW6r8A7j0L
YyGCfruxAxzzpb9Q5cI1P8y6b4HkY1JG5CFeCYQhumRzTQ0oq1bxXePStvJoXV93LHE+1tZHrVYQ
C4OeMtRbnGBjV5vKOQMvIQOyzMCXb83k6t+kd1TtqW6X6QVfzJ1CJsvY9vKAFa53D7UppkkKdY7N
/Fleg2wh9l/u+e+W9w4k7+Z1Wtqn2vCMf9C9CF4tuThGft1O7t3OSCmon8zudIRj2NdSHCuzHddK
zP3OMC+dIOtN1bekY75FfTFfCqoIHCZI7SHEmirs5FWijJqbPLoCCXnLk5/CEIU7BF337Y1puYUV
kBwnREioiOtyau9y0sQa61bIVICaKvs9D2F2L5BYDni4Nd2ZN1gj+V8D9D43Rsm04JgXWRxPnw+s
LhNQ9UMcFn545KamlfJ7JcBSqO3Hj7KqHJh85FuQHPBZODdx0xh/JvNbLRGiewHP9tWmW/oJtjvv
tHU4Qx+TKxpV3U43jvnJgna3Pawel1hOy3jjJRT91ceJEofpc6nBq3jREo9VqqkC/MGuSNnMfP5s
nOL6QsetCGAlox9dOcZAj2xpu5gc12+BVDQLAUd5r/HsjjW6mm7wJCaRkqPgxOjiWG8/3bUcmE2H
3IxZvXot7iRUYUrS9BYa8t7d7cXJ3QArXAAa0de00SiNn260UeqbDQN0HYcV6njQ3QI8+9ax44ag
EMbb6KGM/BGPESLxwwZJxg+5q7BoHLOfGRSu2JY/l7Xh5Bbd9U5lqyFcVurx/zb/6m3VnXi4CjJi
vIMutY5tve4y2/dug8Hfx2of4qzc2TCAdp9v7FVXTBjKeN8Qq/ZwcWEJYKoTwtBnUvgeXe7UqJsY
Pes+pRFymQEtXKcrljY58dJBcj6zlAdPRRBMsJQEl7HL4HAKcVVviRdp6/7wFG7qwdrvvxZqRhms
dOdtCYa8SQnmRWAGdZlQZmg6EpVeE7QHS7TuZZKd6YolKAPX11BC0M9jXI041kZ4i9XIfw6hwBdB
kZLrsk9K+S3/S2//d/chVKrMlfT4u1gxQgwS8Mp8dj4yIw25zNhud5oNxREZVH+h3fT9qvAXV5cw
7GMo1mWY7VJKPI/QbaXkPHOCMaYRpuXY9XKfgR/ALVqWDXO/HaQzzX8Xcg8E5gyvzxQ16ohT6FIS
SEKDd9ro3hXSZ4+oq54sm1tmV11y7OHYWb4feOWi+mlI8PRGF2VWWCLy2iH/c4+5X/KvICa5dFCm
fMEXh2NPSyq1bWYY8LaOX4Hv14ZO8qLPF5bMadVcVNvFfmTjQDfVPDF1z+s8kp160SzJ9NVqRELF
AA1dUVMnFPxc7MEL7BnOn8wCrO6ffacOT4KFE9dcd3zwcvTvxhaft6A5MGqPS6ZjRbnNrhOY6mMv
Xk+WllNqx3Gr7J5AucQ76yeTP+eceGdzA8c66VRP/LsxbQRaDc8VlztmYK8ZQJXKyp0nz4uP9EV7
HysLme0WdziMPoytgVqkc3xsoH5TIR117eS1Yys0sL7+afUYrjOTAUdTUzO90HFEpyPy+DkB7Anl
9v4njrHa+DidC2IrjQz1CLbZDiJGGUSe5dJZwXZQD5YTpfQSq/y32qSTzVBVWHnicJcpcBAQHFWR
JW2BTZCNxaNMqLWu0U4XPKjlLRJxpGCUYZSo8d1CYC9eqAC5yzoZ3+ZnKAjcCm5DhoAnMTyY7d5r
B8/WqRzrpGEoLQUjsnLxiS37OPMo7UCdf+DeRLMmkoKklq19BpEGfP1vgoVuU3Hy3A2UeAgAeuBz
V2Vjtn1S+zC3WM+GKffPd+774c8EZP8tqEiVw3hTZlYGyHBh7aMMjSPg0kxDRtQqFbzBjGYItY7K
bFtPjXaUId9OqTCBxZz8MliLkX7LLmWHbyhSy6a/AQITrU2X9T5Rb3qaw8IFI1kqkoi2iN0z3IC/
1SVc4rOhRXePJDCb9vjCEo/3foArS6Q904VC+a/lMyNpqmhCOZMMx/DIarmaLnkd8e/4HDCj8OJZ
VJGFl8hO/Fd2gndqpeuNuYSP68ALFCk0DghlDRam8nTssUTeEoRwVVQ7W+WxhgbtIkn3Ev0TxrFe
lYiydABCppJhI82CP+bj2Z39bY6ON6cdumEZHvV7xyQ3ToX6VE4rTZCRhqaE/4FJ4W/BYG3ZhP2W
BG3ze+8S31QFOrk6Xxarab2bu/SgI2udp8GxjOzJpOxpHi0wmfMxYbmXhKSwEsmorED2+ZkUhNKC
m7cTUWOog2qkKfCVKbbqY1ioG6M9SFqk1PCyLomk0d5okQbx9jPe7ah5C+jpukE1eQ9ZR71GJkGN
xBwXIXKsA96gfL+Uzmg+MZRKAkOqYmtQnSYFYFcY3OL97JcDDL5VeEZTAdG6j6LjEysDvpaKJ2E6
yYmDvSq9XYe1/ZmF1K9KDbLYyaBRbbqFU+narpDSAKeWQ6nQKDRmbIUHeJc0aWHC+HRMYzjiybUo
FkA6Mv4YDQe/HUM1d4C7xxuKaLu8Cs9jsXU6S80GJygpvtjY9Of4LQbLRBosXcOIQV53iceVZ2ZC
Rl/TKc/KI4tBk6UGPSb4lUxftV28EdOHhyLSoYubF7QtFZh0A2krJzVZ895W5oZ86lg1gOJK5ASA
zuNWQoB0AuGPO9z0VOOzjUa+Cnvs9r4zr8t8BqncMC30E6xH8YDgv5CaueofNSHLzc8SFJCK4Flo
rj9oXuPpEv3jPVY+y8poaHws7/dcGTiII1cNuHbip5seSC5hHiHoXcNaD3uAKtVltcP9TKzvxdoc
7j3gLeNsJbZio+ip7lz3XxOkEdoBV4L3RQ4K+JRliOK+IkCxZm+FUkV1gGA2Qiqs7w013P0Jc421
qGcXsYfQrm0mhQ8RHEYxS9vjSMD2QxQJX/eW478zeB4zDGirRthdzTyL3bth4YFywn4Eoo6Eu+DL
c71ig8TmaXUTbp/Ynqk12Aq+VquCjnar0sLggUJPPDkmy23mOrncNY5Vylxo9Toz+l2LMCMHjStp
3zu5OPn/TiZkmO51XoJChSrfKbBJ2OyijReXndRnkyf+z0EUwkA42il9ZkmyMoSdmIKqD7NpyG94
2H9cwjNdOLAmYOCgN1ggzo0KAf+S4nypHRtmtrROUiSvpXKgQKGn6/CmN+sDYl4rRCJU3U02CUZg
aIAOHR4cQAVFA1bT9SB7ifN2qYYvynb7F2Qi41HMuNNj+6/AY3Q/3OYY5sY4NAjgVY2YWpcsdR1z
zx3joVV1ha7V/dW9Gois34qcmsM1U4MkGVf/flXyJw/OaAo2Uv/mIzGozBmV+/Zuvz78oA5QKzWL
ieBZeSBYZApxQieG2h4zFZ67mJLkK9VJDLNh8f2EPIxt3AiSV86yN58YsEwbEiSHlsQMuweDlXwE
vlMBLsyhpqWD+1aLGzWt6jUQyXzlT/kKhR2GZQbjSaZ0qQScfBrcUEJl9HeHDFL7EH40Y3Dk0sn/
l24iFeCXPTxtMAjFdQMcYB1E+VsO802axRdsuoYa0/FGDy1TOplhIhccuxFViWSGYWFr6R7P5Dtm
wv12goq8NGqR1L7wbslJbDnB7qQF5+7nstcrrK5FPAFlxAkr0VSxGHgSM+GyeIjYiHy4txGJ5FXY
kki64rMXvNR5v9jWMUuUdSfhiRxzn9FGZQEgGVJ21ux1+kTPp/3PdgVSPuzm+K7nLXKJoq7Sbx+6
43QeK44wzgcwtCWjBbJ203kKPcdNHlQtxohHkR7kgSmTubdrD05x0H1lLz4IMcne2SWcf5ddtwqz
FeSmibNPBh3wadOyFZ3rWXHaaQk1FRine3k/FbdLPnytYjo0lJEFHfxaX9ZzU+rOq4yMrwhxuvrZ
RfhMWIt9t318OblaKtgZd0p6/XyNNXZceC3LO3osFIbXSWmvaqHyRxKUV6EigGq3XX7bvL2N4vt9
Tsp9iXUwnFDClVDDTVF8sEJqjU95GjJKCuOYAj38H5oZL8+OcFLtkIq5FlncOz/ul3ejMi8QkSc6
W8sfdfJQlu0oHUQFBfyR19QRcvXI5n47So1O/DUxNdA7HtgdLJfPhgCi6XGsAyY4mKmpv5RK2KRq
07OoHhyUUsT5X/UU88uh98lp6pd9RhEoHWKFo4ICe6gfE6HUZmOeQQQw47UbgQVdrxBAfQN88Clk
vJKjhuZN1iY4aBto+YuGno380LCChcgUT/FrNFQUgbWskiAxX9naAtpKi6aj1L1AU/Z340hceHoq
0tkctcEAcMgr/Yj2Oqoo7LkArRWQkeyTRphHG1qAEMiEAlbkDpd44shRVru2W6JTgI9ZP5T5NOHC
xMrvF7ejD+DUxszvwsZmW7Y0+A4C+AY2H/RITy671rXdtdiIv2FvITAkVUmygFh91bgDzyRkJz32
CcU48ZjMkXXNRe4hQoSlRhHmcSkEzONsEaANjOPVCWQG/RrrRoKKXYOOc4Kyas+lYaGeAl4lYRme
6y5VYWxIT2UR6TJi9Ff+3NWcsojPpCEA2sNLH2qn6Z0AJ5GlYUifoPe2lWiywEYnqzqswmKOMYKb
++axCgjJAP2vA6TIkJtdRKE4guamuA6qKi+CPwFRIaqY6HCByb+qVGKIBi3gujZjXCKkJaeEom0+
HdyrHcyQo6O8m7MZ819cCUFQr1eGqiB69EWu+A3rpRUO9i+8c/E24e29mdequn/w9yVS5xr07mu5
mC2PZcYqlUU8YNwPrs9yQKc+fc7gIL2KeD/j3K2jAHy+2rynSaOnB0slt1cDvPFhgJUUQUYx8oTj
7Fg9MliB57tNNfMgXb6OBbddskHfEbvhokpLgvhz8C48MfNrUBZOdCK8toooUQP4hxHplUvhX7EN
hvuVK4bF02J+ue3obQoKFL6DhS4Z6uDzz/OipqipOE8qAD6OWLXD0a1Y1iCeOx1u81fr1/pwDRlI
sXnlhTMBVMsCeAzMYNpnWsr0F2PiaSQ1Jp4BDdSCFu7wuQCEYFVq+la3lzpoTIllmpUUPFbtTYHr
dU/Jk80ScugM5IBUHC8YM1WuPxE+YphqPfPQBt08A+2XdrkNdM46qyduvjmzVXHwofr5KIdJNv/l
avS9E1hw3q5u1lhQgAzQTk6JC40Yf06HZ+XS6+joJDGY8sSywvJCYmXr0opPdpys2BnI+J1PyzLL
WPc47JaFyk+E1kmfvv1e70uNzdqt8qi0apfn9i158+YUdbXrs5fxSJCkhR8596ZhVLpdq1MFyM8v
WHTiyw2hM3IAmXTuhyiZ7gwie+wxxTxinRQD+KpPc4oI4ciMHU/0x0D0Cd3PRYEadoup/ekX+jlu
C5bkn/O6w2twRDC9f8QlYICn+ozaWpO7q6YxW92iehcKzGZvuW883b6hbUvH+vFuIkalokJwjbXC
rHP9Kr517x/Mqb6XRepBC9KzW8yNMOu7IwG0ZQk/SgcfTqELwTUyvJCDWO2WbzxN/o93AuJPl8QR
Q3ABCBUZ9kTQsskO1gzQCwTVe2qh1IqtXCgK2xPsfWisEBB3tQclWMJP+ccFM/wmeqtXXFld4OlX
xxhO/8Ezol4jHhQrZRRGSTo7cEOKJNsiBchjq0ZZRlw252+JEXAZZX6vvgPlgmEVgoFJhvDABnAZ
gOCdZt+bh4iZ4Xamf2Xf/vYXuLjaQAaHDbYsrvkGKpev79VQjVFJJyeuib8tvrKJHc6jhO/DgKOR
L9GuQkYJwyaeQvgNproVSda5J31XwXSojaNcJn2MfJZR7pvxUHFX5N6x60nlGOF/TJuYf5F79RFb
fWjjn8zIE0tnx3n/rSUuI21Wc+1V/KFYu1ocRbjN7Mar/VmrGsNR85aaL6mz28NjbgxA6+7zKJHm
rNxY9l55PRmHvasPF8Iz7R4pdHWcGsIOAAptUbmygXZ06H3JOes0HlG9ZmIfLx2WNjVm1M+CcCzB
M/IhAZ99EZHopmsTeVePB2IIadxRCxEwKgMT5+ARSmDaztKYQZlIaRNo/p5iJeNJvTfUf9xsi7/H
mDMIKAzQr6X/oE9CPmDEsRzXlEXmm6bY5Nsk1YHYqouDx6a77n6yHw+nWXI1qkVPsHY2AG6nfmHj
ZRh9zhU6kR7loY6y1IYvF1r4Q/XALVkTe8Ap6iq6/09k0jVug4uB90o0BNXh6OIESauUKeru20xE
oZfc1gqQx3RjwKU7RGNbgej3mp8uCR678H7TKIgfGiVYsevAFoTTQC5OQRsK7f4Xrt0MuaMmUa3e
753aWYxJ/zpU1UWO+zuphr4Vepp1eSANeUsAgVslIBvWCALSLlhMu1uHSTx07XwYjj+jaQnO1CHR
AGHpIhSq0qkgm3fvUIcAaNUCBvjwJyZuDMMAPCwzQIZWS7gYTlTofF2PaGxisdZzxVFNIThD1S5K
OybEdkx0SM6G61P/y40qVk82gUvBoVW3uSD2/ZdR42jFarT4+RJGiJugSg9u2iKn1u9dY+lneDuf
G+/BWW6I3xgtln0BMEdWWCkw6nqKAfSYi6FysV9yOb9UyTsqE0EN6atXOa4OPhG7RQQI9onOaFst
sgu+MKwbL/LGSyy3x/I2uys6YnhDfswmMZGfng5vEaXXY6Pvr2P95PNTxR0rqt24t2jSQ62zzSD3
C1YjEFK5JIlYN8FEb1WiGErIXO0bhe1AUmRzBkOzaw62LJfwYEU2LPVO/7evVVhW080qrqgFmt0q
wcgdHZ5Ys7BlVqE7klGNpj1EpytyY/Lr8c60As2qBTDyBVpPZSAPaaKFF+UabGbAHVIE2RP/4h0u
p7sIUAqAEpoxpmfqHA/IfdSh4mvfwt6HoSZd6qHIPqOrgRtUIrRj2TN2A2soKhnD+zJvC9nzNW6O
DDnKZs1F0PECFA4hVv/3aWj4mtbZiYTndii7J3SXb8r9abp63nD/4ZGgGUZa0oi2TBpZcLAdBsH6
lAON6fLghfgqETqrw/Hgx/U/VSzwA8UFukw6E1uE646RG6IMSfsdBGYnUodR86bvtgs/CyUOE88L
CMGho8PkScePngRwtB5hJgW5G9K7CsQWk5GLscdH9vIk3P4HtFlxVCsi5LH0HJGUFpyBrRUPzH1i
avRrjRGsZHKrDRmEx0aRFL6QRRjufMhYaxxVO2TKz23E9GeKZycvCoAoXjs6s3tcIlFHLP1OxiHf
WuG1uSVQjs9Dr9u4lj/LdP4YOA0+omGc4Dv1GZFkCufhorpRquMyVWokAdPYo1jm0gVsNP0Pu3HO
+MDk0HSknI9MeSs+XRRQRG2UYU1n6JbhbaUpY/MfyFODTiWTLZ+zXe/TREKBS26OOCt5IKQX5ZZH
12NIpFVqg2OzWZIQ8kRORz2lgaA/uJ0Bo7qgCjD8KHI1eviI8nO0WQLRfowc/dyhTOgZStr2wzx7
ehLq3/lDFWpzkV8G8ELCwJW5xbjRl6JsDN0ObiUuP13m0G17OSFhwdlatBGdiu6q0enKcArGnJgl
DkUGltTohoahwHRoQ/wc46nTfvRFDkECZMqiCKaipHENFylqbufWw+oOG+gFDkRLB+PV3UJPsP0k
WwwPPkPVkAmI5oR9645l7yV56Lx74hLIVvjTnJFyOd2i0PzKv70kW4mxK7JF8HQ5pJMjg1vDAhCW
ZJhR9Caw/kQEKNUwXNH4HUQLJ6Pc+ZfD5lM6fyJWZIambNa4hyCjAht+NaKbgoafH0ass6j3SdI+
2ZNBh6T1VMU0kx9ovxVFlMcM/zmYm4ky5JIAD/W3lzNEcF0ypIZGW2Flcm1bw/HoHtOd6KH5hQJM
+wrt9spAbL4PPcqKoWUxToDfVg2ZZpw6YTLEwgOCTVkM6cfVpyfOHBKFPSqOKo5sfXEgx4u5vt9A
/eDpen0qLHaFYtzGgcVO/4e276q4gWwXl+FCO/tQxQYl5g1kfc2D1/WC81gJXZz0x6T7hVo1USTP
mHsRld5BJfK45Dl9sbVXnTWiDPZyISeDZZlgCWxNNjR9l8TR7/K6nH0hw9v3/k3GPuN2rESEHPvD
Ahmqs/bGWRA2nSUJ87K5ck1dbwfhmoWnUTJY69o9aA0bY5Smw4qf0Q3lMbUPegjW4RhT27NaxSz5
7OyaueFYhyBYt33uEG9sh4e3HOQcx4Vf3c8oM4FempyAY1DHsEadrx7xQkb2yTxsH9kwtCUcIH6A
iGieUtL/guBDxeYzx9hHXPwy2Btx5wTqbRNbiBRYKRZ+j+lIqzr3PaB8GyQgXT4u6b3SszhzGWZy
qFOzVFId6sbv2U1a9RtIYT78WNOnodPR0jwnafzt+64FkUFfRAvB31fwxFQKxGpDqZAMBD/nQ0cQ
EmLU9PwVPdBBFl3X17h03uFGljfWTJnRW6md+9Ws9h2Vr1UmZI+egW8xzrQycsl7GBlhL/nodws+
28q49Har7qSgXfVQOY0aua00WfKq5RR+Z5Rf54apORTWh3uqzQJ4GbmN/Rb+79gq3Lp7FGDZR0oO
Ymhv9hp6hJEmbp6myBiEC/LJ6R14JXCQmiYnN9qEV4gkb4Jb1USiqPeiqVGGbk4AjTphLNWXR1Ht
QWktzczf/0qpdzAZ3/da2dSvrpSyBdfuPciOyi6DQTc+4GUTYDeLrKe4v+efWw1Y3NhWgbBUTMP5
XJI58PW3gYNF/At/bxyvnqOe9HWMTSZgas2UbgobnjJ8SQEF78hg4v2J9ZBHJTGBzfuEw3l7r17C
W1pzT/q2Hb7gO/SxiH7yvCn2EWgSZEBiJ/KSM3WYrlSrYBfxwpfv2JuLFI8YDMmTdIFKaRHiVOv0
pqDy6U0/I5wGthHgu4M2p/6RPv5TQST3VMmO7E6tG+XRaKosTfGR3dQNq6s1JFRrtlHryZeDBUpX
E2Qd8FXWankCcNhVd8DhBjHdDPWtSOsQfWB5b9mdfkQrmQINe0tCUL4LYScevZq3ls0lBnRMOIuY
1O0IKN1CE6j1EklGJEvQTFei3FBAWmZDHVmjEVw0gbYzcbkRtYzUFlSftFrEoFASaIBnsJ9GhHXY
gs1uDQERW6vl4YuB/ObWvfr9IYpT0SJNTVis7bvlhBR0+P1+Oez6I9iRN0yi+qUrvTuVHMXFE3p5
EwynBjshR5dEOwad7OkKUUDr+fiPl8XJFfbB9BZyGTLSxFdcgh+qG943nLJhxrczqpQbipylfO9y
Hk3Ua6KEm0BJt0srckLWJG7uOajsyhrCRynbjMkB5U9gT7Pq9KQox9oCW5kOlGwudy5wn+kvncLn
1DRTj1z5LBgMFCt4oMxy5aoxwXfbC2mXmRQJf/k7Utf0Zmvty9Ov5evuQ41fD6r0gL6/r2ppk0TJ
BSCehCtZtkDKMN+ZyZMbLJ1BccFYlwIilJZTTj5F5AY/4Ze+AHX3LiBHlij3AFNlgqKvf/uAIzqI
oq/qf5xRDFNTPVv49p4GWY3CXakVq/uhj0RUlIaPKcJxYRWdK6OA99/jEeBspuEFgEcxUQG9NG9F
dl065YNYN7ibbpEoEtqfTlY4FpvaDM8rmpsvU5HGnKyFhZqF+qWi//g5U/IjlBYZNQE8bCVYGBpt
k/6yfczGHJBMhbkZxw/w/+u//wh1cQPQJuD8Br/1s9L5MK7IgB+EnPh7PwdOZMmhydoPR1o0N6fg
M/NTldQIW1QJEltfdMFPhfbhT1A+nBcIDn3iHcvauRn5HuCHum7oGlx7oEkdjnDdCX+aXzIsLeOV
ENXiiSV9Y+rLkdD047KTdJWOQTR4UOW+0prHi3uotsJ+pNcCMoOTMi/xSFWNTud7BNsXvfFYQ0kT
m/V0s8CYdPrGJFdXaXmQRVFsNThZDBRwuCZZtkbYxi1+hHbtUFinmapr9aORNWmMQFY5WdhdRy8j
Amzo7TKJCwiZXWAl4sjT6/Aegfbw5CiYfv5DSw5DTwwVaj+5U3oz/ydxnjsi1wr7TfdaJryjFCL2
oMFLUv3jQ8YPTifwGHtNVwrXowX2aJLXLmf4WX7OxGTDIE1plczGX7IVpLQFNSW/4l+tRV4XfLVp
jajLxeUqKzKvUVFr25I+7AVwYb6XvgoD1wzIXWjEjH3Gubtn4E0XP2Cn8s/caa/7mApetnLNEEK0
E+CGtURIbA6ZwDrxa75/aGYxBAC9C4kWuEjmIENkgS4Hny+5ANV6PIUA5Reicm1rbCfOhPmKE67M
oeWFkuKNMHDvgJko6RCk38rvr2eKpb3r7h1WCQ7VFp06XIkTLneKypnP91q0Y6ak6QBOsDK/H0if
IthQCHzdhgJ3syG7dWbqiIjr3kZLHnaA82hOJwr2KehhTLobwUmGFKNVdOzPlmSLVSkb3ilK922A
u6jex5iGiGGUAuq4TYXbHscTyYytmk/Bij42u1qSbez/UUDjqL9xd4xcdFoIkjjtItDWdxPo+hk3
3njkAcOzPXui6eroxQ6zT+u4h45UHun3Wz8v8qe6UBr2PrsmA18mKwUJ69HLxQpwlgWPTd5vWNqY
OFQsT8O1+aoliigE64lzdxVaJHynK7yjk6Uwhwpo9hklFy1VKz45Kc26xFMXCZmVHKjxJdl4LYXV
Anyk8vtSBOGYOdgJy3lZpe0MzImzDFA4WQCIyhgrDC9q4ORkWjvkv0Tx/ZyoSYo+oh6NHTP/sRik
05HtpN04JjfZ2xmQOzK2KP20WSYuRuXa2zfExFSRvd4uTc13wAB8RqUBhdCse38ScDzERFkH+LHz
7zp9y4qE39dgxqlZVIv5zTsapkCqISjD2CadUbp+cG3crjHokLP+YiK5Q6mTVQHc+2BOI+7y9pvF
MzOZ7ZGsFu9zkK4mlZUFt6WTzNusDUDvzBzStHUtv3X/422966t/nZovfIrWR2IvcmEDNDVehfZC
M6Mv+wLMwY3mJsts7YAqlfeJGupP1EXB6VtHn8CWlN++Sd66cMKZfugALCZHT5Icz6z3pxMaJHUG
/8wZEU3XRGXwODY45hDqcZUijaXcP/91oFe/6seTdNrCckHPqshk/lOaJQTH+h68JFiGuD+00EqF
1McS0iajJUfpjV3zSyrdgXClb4EOb3P7iYBBIj5gxZa6usgKTKKvFpUmr91JSLHLE/RNKbyfZktd
h2VrW3FJ5UAYDbM1dyo9l2LmxI5SQYlrm32Vyox/5nNR0DNcWB9Qwl5JQGcK51p+QO7dK9MnVTpb
c7U1KzXCY91qQzlX/RNuRScqJByFV8UgzoZFL4/kvSgERfdbNfKyAUbmhvHUA3GRP63lxBX6RjeT
6Y98c6DBuzkKuD+2slnRGQULhqMFYwqeKf0B72tUD6hRglXLrvH0tVXhkAlub6tKae4Jn2ll0DMa
e7zidzbJ/t+z4PV/iAgY1V5jabTSaA01+U3+Y1lwfxFdq/KDBHOa238ytdK4JubbZiQGp05CsX09
tpj2iPPKScSlaaqb78udbom+fQOqiti6g7JyYi/80qcyzEszbro7ZlMvILa0gqzLkVdg/hKOwBLh
Mc2iMILGQORKGVYoDS2yYKzxXDzVYeFf4drY9hy8cVFjspETI7pg7AhTkEop0rEGn+7pXF0kOsw0
lYwEhoW8Z9L08/X8cZvI/cujP0BuU6Xgd6dEHpboNQnpl2czoM6g7YCM3wLjeb8MneR7VDv6Y25n
ormwcx1IuR/0LBoY5UE6xzPJWtjpwpZnSU2kvdN2dNfzOXrZHQbUANeZXSP3+RiNgt9J7nq41wWr
1qnKkVLhN+rj4n7axZOuSksO7dWDisXGE/GT2SR9VSGtUbB3oAH22EC3CJY0tj/vWd/UvaH5Zhxu
kb3xNW4aRgV3Cv7Bch9p4RDUvKZADJn1DNz7/3bd39D0Qbk3zZ01Lkm4Ndi7Ds5L69ofs/kovGW+
6O80AGD1lia4CU5UQR/aApNJ8AT/mjP4DweXOm2+6ufoR5Drh1xaLAPMHAA3BRxGPSdqjV9Azhcz
i5MFW9ieoDUu2L5W8+neG5o+l5a1CYxmiA4u9kYaM8Nm2fvKx0KmYzISuw8PUONNE992Iz1afUU3
yW5+tb9QFxqy4Nty7aq6dzW0JQpbqY2H0GAq5+/Yqwt/gbp4EVidR8TncXQHjlFx7Ce77zdXsldT
yKvK/wlMMREklQIECMSB+jUd/OKCvBavlr7qc3za8Ll/y6efS2TDBvrG5vIRu2H1sG0PMJHzdY/D
Vn9KaftqPbmn/+HFRqdh8FxsaHR74t4n3YmIeN0p0A8AD6eXLSVnfoFbjpp7zzN6sGqKuuvKMWIY
+iPrMmRQxjZnB70r7f5SL6wUPLfboPhBJUZpgk4gqOajCdVYTC5HKlaIK88Pke629qouv2eC4iVw
kfN1y+luTC4NPglhIwgv/MczQmvKAZri7zvMm1AJjlulMphO0NwQxv5vjW1bC1dLAiDhEmSyRahx
sewT7oPUG0HvdiqOuoGiYKwe/MikxfeZF+1iBRjS9UmtijQFdSTV35tnzGasv5cdPKCRrDPMnZ3A
JcGDJopyjHB401/vJEeSLB/K8F7PLpfnHOUVaefSnarHpVGmxsDgOlFRmD2OX4Slz0SHvx12AabI
byT/izRrf9fcb1/RBmLZwOjRbI+66YQEfM472SboOUvdgdgn61v2nv1ow4KT9bfvDNJIleN6ZjNC
luuOjdICmHzfSJWc4giaZGC03Cijp4RL1CALztDh6J+6qcP9SoclGbZOfm3XjkAWhOsznV0Q5QMu
4B6GhOH6+I2rx+sgDm8XFwOsNszcTK+3TmrydzpXoxXzg+U0v6KaL1uboRnaKTTAgbu9fsZ97dqM
89Km3WFdCvhXWubbx61Qqj82EgrwlQbuF05Kq6QaXxgv8x/WonlikpgtAtfX9FviloVml+01ge58
9717TM0Mf8g8wwHW4gS/JKrXsmRlb+H6Ez2TM6uX54jMKQDr9l7EnIbfKqIDOQAGJZDlCYXv9nBl
UL1QwatzZSE3xsB6BD64QRFYFJ6UjiGwt/ikcSy4J6Yi8Psurce3B8B4jsntGSg6syVt4824yLU2
iNgO1kbrB5nJK2ulr16g3kO+c8iO4/Nnq82dU4qF3uS+LvYKnQRLYfseimFsRqh+DfKIwaLF21/o
uDfNrdn2WscTA27CnffkhzGLMyXfrVp6q6wYj3jM5XDuHMHkpOKJw728+kXm6D8d4Hy00ofEAqT0
Qy1QnCfenkOu7g4MYOCmF7LBQ5ZSdE/RoVGQ4v00q0N74K2YgrVOnJgSSildI1mZed8wvMa55nHI
YO0kfVg0nNBwCaoK4IK0yRvtvbx4LC66WoY1MDS4/dqYm/LKu9d93QAB7Z+By5p5QKX3SYWDRxeS
+Jcbg2/Ut65cxz7qRv3jHvgQh+t4L4DFY9cwkDenYdSQkGq0Pia4NplsQhVlt5NjThfhaIPylqzF
4pyIpCqy6FpEh+Yke6IRqxVy8GTNARCaYRMRM9vMfLSM67CHWnRLSePUkOmJUaL7di7ZD95rFqd3
xMWNSH2i3MxE/hehjJQkZWecM9hvEOfiRvLdoiNmFCWRsciYIlogs2lKTEwPiMdK0ThSpA9KgvzF
jtPLBItlVdmhIuhewVTpoApZZMYlMuF7K1NF+bdOWWWj8XbUDI16DRfjoHqd9LxEXPbx4HoTA4px
E7Juhgz7+L1RBOXFaGQdb8q/XWY2CoX3144iMOOXS1GjvdwbC4JM1U2+KmeG3W2Jpa3abWsT0CKy
wIwjWEmjIhaIJM5xjnb2gp6EXk+V0vJeA1UBnRyyv9LhkuO662B2jpjTNFMoUwRv8vMLTDj4vm0U
9a/cK9WQ5c2wFCNqrIET68fU7rbgDPKw3xb/fYVr209ByKdUC3xgali7yd2RI22srwWIgC/IWiE7
jgHhntBoKNsGWPP2UyzEtZ7+Y7LezO7bxTVe1kSd5IFNylXNysfANLMYBnL0AFNu7gGRk5MYYITe
DL7fQFmtynHgLKf1WYtY58XwUDGG7M8yn1uXxsO8jMt7WiPEoTLL8SLA2c2iRlaDMxMXQLJKqZJx
lQp/HldGULET0DWkhk617kp0wG6350/l0hv0nuBG5ghJtXJO7UBeO4fDfkYlXqu3s37PfEnWlRPb
tXrQdSIR5shjnOlnYcbOf+iZo+FLqWaIIxsVqSlHtJ3g1LeDu00JlFsvdCernqaf1WwIJUvovqvL
mcqsKFI9DQO0NogALhDgKbOGhM0mPPH9vD2G/DB8bwNzYtTsmDa2TfQohpx0lEkE8GY00lLrAhTS
3UMKqimVP4A+kbsgB9o/eUcHOUF5EitkYgPxhTcPbBbb1yTDpf2VQV2XYBbnzPHkCUkTt2ZLhYqN
9YCdDmVJ295yVfzDT0MdCQrQ8B4EvypdGBUkp+84MYiRScF8Noy62fp5U7ifD7pPYBcr5DPeysnQ
SBgDYUlUVE4NiN/aM1F+qf17Ve+SUPOVdZ1gR9ilEb+V7OEZhRmhr9XKGyQZ2GuN3FvfO7nE4KgA
bahOoxZSXDrvCSl2Yh7qGxiiBleShU6xb9YPU2JYqrRO8S7O52BnksMNmufQ8cO71XlfnO8IS6B1
JFsH6f62leE550rcRmp56DJQMkcPisookR9dVC329nIqrd+lzOOV5wb0+MEEChFp4SxCUX7xqolU
0O/obBDJ0uXRRKDmgVe4TKAz4/pQjMTwYJQpUFJzecDBU3rhMjbB/LRvQD3BsXaxh/yfLxnXr+nl
hVnG/VpVY0Yu1EU56vBxCNTRFsXJ238FC+Tl7Mh77SBL4g4KnPiBUBWEchyxcgOewt3t436qJUFu
fN7sLBxgXa9Nwuo0zFMtCWwBWhBU0qU4X6mv9b5lLat5iDSrOaL4Up65ijsiDGXq1HVVv/k9khK/
cGf0M2qvQ5ZiksB84mn+1XxPcrDoVuVvkyVWPlHkMUw7C6f1DX6JihKwdDGA+X4bLQ9kzzfif/X6
D84vXS3C1ADtOc/MRUGb4Laf9qx0vw8xS0A4GKPFX+YlVhLcQLdagtcy/S3OYx4xBCODpr5rcZt4
2EdqBLcivMK2T6qO3iRreGQkuB57ClR6cBbHCO/2aKxsFxyL7EERgHHRkr5jJGe+FyIChqM1Siqs
hY34utCWWRyVzwEx7FQNg4AhIuaH+nWmrlBxNnBrKS3o0473xAfmKg0qtTWSaSBasWx+bj4Zp5MK
894wu1qKxIFI3ccYYoK10yja8Usj8Kf568jiM6mU8FidA/yWQfcBP7tstIKvDgVjqGjODn3WqCfj
P2AmRaZa66hFcmg2By+jvwM4/tdJ22lxGhciAx3t+538v3m1mkwXZi7vgNB9/fkb9bIX+SKAvHIq
35bkQQ2dUrB3Dwe1gn30j52defWF0ZCLoug2UIpVZ68MwLOcT8uPQEicUTXYFqxxg6CmsK3LRPP1
wiPr++WNpSwHeM2Nlc2Z33IjDUyW9Z1k1q1Zn7RaPATPOEDqC+7/8tQFzN3ePx3ImqFeiN+OQI17
C5g+hHAId5uFznGXU6rh7aRP6JUsRcuhxZuooGdL3hmY94wDaGb5KxgjPSqSV3FKTJpeZ7+okM2n
kN2CQcHEUfupZfeyE3ATymrkebu/WR4X9+q1ak2I9HiFMybDpLGHe6t8dj1BbmP2wjdkWiLnvb33
FCiTaSWRPa8GynE6zuW2LmeiktwSyo5Jv9LXjB60O0oC2GMKWVpQeWpwJ/ZnalvT5c6mQZtyVkRr
wtmYNBlbpS0d00txnQqpQZEtRfrERsOUhrUecRVJjhh8K2KX2QzZ3Jd9frgORIPDWZ3pvDv7kE4N
by1j3fjtEpb013BH4yBsJ/3Z3PVt6ghsXEvfRc3XXayTismwtm1WDwb7vnGg9vf3C5KHTfAaaSI8
Fj+lmXl/X7zzbHlSJYIAzK/XvPUjFww5SYdaASS9nHQpYwznq/YzWQlZGDuX67SGDXpwuxR7cVTb
/KAa0WHR9jUHHBm0RKIRdZ7NEKGHKrbzy5vOjLIOpsj7DxxruXmnnHpDSuhWKxFxO2cGL1B8zXmh
Msv4594WMBZppjTNF1giXbI7EpacIOgyG9QbJJ59E/nckzaZUmoWaweiYkgA6ZHyngT+ueClPQnp
SJ41FB/9+lOW2/ruZi4DoIFNhZlP4Nzpyc9zvaybRkFK4sMSZfVHko+5o0aUKAHWBjE1p+4CphOk
EHLQA6yZjh+ZEKF1P/Ud2wi3ojOY1Arf3hXPk6XJpJBrXaOV7XJBFvM4/BWfu50j/JvNtrkH3wgw
DgxmHaR6OA9U6TrentsCGT0MnM8S3ZPnhwm/3DwIktyiAZfVNF3WULqSA2s4+p5U6dKp3HlDMwlZ
lTpkfmLO+YMak/F/jggR5HO9GULFEvkaKIuoUwlDBmL7+Y88WTacNRmd7iWT7+t5W2qQhBp7IyWT
UyUt4uCjNrot192k5vitQmxHwKqLTGWag7hqtpvgyeqbGqIEr3WLQgBstpzGGWvKpKKbD7ZaGxGP
MnEaubYFxVfEb/ijZWiiNCipXedWtMJc9zA9TUqOPLL0aNi/PYX2e2IjK9BEw+qSkBD66kClOhw0
V35LcmLZp3mpYHTxu4g85AnpkJMWuqhAptvVUWw1rkpd+Zx7l/VYsr7urhCG7M1k0u5C23fpp7xU
Fg0yjWjPBuAwxKNb2O2nuoqEEEz+QnGNDTEQvwfleeh7CnHexSW9pQ5RK+dTC7TcAOrLepUUXZXM
8jizCbUjQpRU8sv4p7KdUwkqzQ719vj82xOs8dqSQ5LIw7b5YA1Z0dp1bQHQRcefHrL61smVFzGa
yU4LPTcvmPoOj6qrHECp212+73gFeVGmahHTNwy1J6Ur88kl2a0/80A6qQx1+omLxgg5iuD5LkN2
1YlzVXc8qVoV9rfOTrjY/S13IJcUhlF+2UEJq49QIZ1gwJI9VV3Mu/L4QMX0wIgHEI5FIksFOr2A
DUTqqMm2S/RFZFpeAWD6/yqEgB7EvTBjQCzNTI4tCwhcUxzAKr/V+KoCQTk2W7YAXj4UwZvIvT6n
93sMgX+DanNymCFgL0DB1yq8Ecez39oROLoIAGLMIOT1LWC8PIuhd8goG2dwmtOt/QwUA020o1Bt
DNA0mKDLetis4lOffIBs/fkYJOzUcF//lFhtOVtUyM2LP+jJRXIQmATRV0k6U+3K0FlBuoIHlLvg
C9RuZK/XEPOFzRTuNYymbVXDubsg15NU/9Ga8i7cC3HPy+NsxZthnzcHDnJxP/JlZ1ozi9KTB/iR
fUAr403xJR6e4UTVvI0nwKQGeEbxN1yUNpbGB24PdN0N5DVNn2Dn/YIFAQ/5PPExWlU3zUSrnZqk
1miWgGgzlD5Ej2F1wEpLZLDe3h4V7KbE4WFBnAF+0PRk/tmyEsCFoo/LG2P78flUKcEcw5+Q4A6I
feWB64+QechB24D0U1A9yldjvAAvJYeB6P/tumYh4zg/tJi54bqikHRpIhZyJDAx1kTzbEfq41Kf
vrrDAlctxfMekFzq5FcIiJIzVmXSz/kf3QTkSvItZnjYUvcy/OeMU75QDJBMh+2+IXRULewNbVUP
JfOdE+7qNz1gTgQuUlp/8Z0NNf5cYo9+R8W5Bx4bAsvwEdVSWBZvRefE+OSUOYSAi7JSgTxUaYiE
83c+bbp2t5feqL0RvCVft34eWV2bffio7zGq94T9cXGItPqkkmIhCD+iyoWWMK9xvNImuLi9M/WS
zRdsybzm8kTstzgWJDt55ZKJddwmb2zbPune2e1JeV074+oQ3N1VL7+84IoXIK2ZnpUKpP/Pi0YP
k9nQ6Z0veQ+Sgz0xWRBJTTsR9sxggV2HYBpjRTiFmWdDZ+Qc/WmF4pY0RZSZLjwNmlufhRK0Km+7
2FMVmy+N0qT5XvqNCXlDwoAkRpxZx24JMpSexBD7wR38Q244DZKnlZFIsRv+qwZXyKiE3ax76KFi
OzOs9Xw7N0RIG4LdfUdP3G1BvbSyzOtyUTjl6DiX0INIJcQE08g4oA8eq4WEwZKHufmu9Mbq8Eak
d8E26ArJKWyHRQvm4JBeLkRCOPEDVQFfR9//y7oLx1pYsWQBUbVFFjM+uMevrC0oQ8nWAycSq0Rj
V5F7VOJRHT8uBnM2opEvbVi5lcSYayJM+lpxE9Cbd1zDKZbnBmX8GJuuIXV0STLhVQXVHi0dIfZn
BkCkJFEIeGUt3VCxC5roPe4gLdsm71FIPGkd4B1uHIo/kX0VobpCLEjQaBXYqxo11gSuYiY+aVkH
t2CJaanJBOfXfxGGs+q4gIkabw6VWmNGV3lx4JZQxkxsk7+k5cfZq23dNxbdnnT/EhAMC5SySsKG
0psTWvk2jWgxP8fXxKnK8J0AZ/rtjWpW222lLzHtB2DXUTjy3oXKp8VZypZ2jw/62Os0/j0Xe1X/
onpA0ZgX1NqDO3jO9R/+EJobUn2aZE1eP61ZVIib1KrMO5DEv6xmLD+HXe1BlzZAqZuyDG+pNJMK
1f3AnBEa/SVSnvukpGfpv8V2gIFPq3w3Ym1abnxMjIeai9S2Id5uJJX3AKmAPHNW6UFPDe/EzGpD
/P+JUcXzkQapkIGTSeCIkOvwjRzuHgyFkbCat6EXQUQfQR+X5QbSu96uHGhY2gy6KZQYZ5ZRWbJa
4XViraNHy1MBR7gULDCbhO8QyCk+Fo9s8xB2gHDvu1hGR9jYc+BpWJQuvkoByPzPz1sHOssuDeR9
2Waw7vW0YI90eYyUNXSNupPr5mpqTO8yth8CxZXVnqXrTObiAT4WORkTCEz3MbAIStiQ4v3XFCKA
UDVzPscpX3LVCIAwtHYGR5Y9BjPa5LSWlkUy5V9Lpnw1sKnxIF5wlWWRYaOgqyv3ca1u6Ez5YihG
5lh5qPMIOETxWZlc0fAoAVWx+bA9uAgY6OomVtd3irdJ4ZWhFJI9XQ8jezWIzSSinsbqp/7QhQj3
Wn09c0HvoYvekzhQfRnqphowhuP2I8GNe3mg6/YHDqz0ZWGxcmQrfU7o+x/bIQL431MMNcZfVOua
NuRl5Bi1N4LCQz7wP0a4fK8y0QCv7SJl4+DbVTBaZgSvIFWHDNGLIraonJNvvqNSuweDiJAGXYSs
C55rm7p7g82ZA2SDfC4MyQjqP8rAPj+YGLtvWVVZt5vJ7uhBMZF1IZpAUxnO5FqVK+Uyzs0PvYW9
8zIUs1/1LaOZ9QxibAH1mw4LD/3i5lq+kiqhJNvhxbjSl3EssDlJf8VO5jJVV5sowjbWXFgQYT72
12H7X+UgsJUX7r8XQ283cHCfWsMusS4cso2tw8rRbhndedkimSiwJFI/w11whES41fUi00xBYhB3
G4G0kJ4dblR7ShLoqXUJcJmQDxcMdZx2TvTfOVcO2j+DTdBdOpHfjcNMds80zT8UWBIuJgWFTh5i
+mBbSgWdF6KQOBYzJ9Vo9lVmzd1UurYNnDsGuOyDxI2rSQv8DhKXl/DIH3MTZyiwH0wd/k75vVbF
Hykps8i9Qy13PDzWnb0dFIoIdTbOR3KQKzno85O31gQ7d0hkZ2IpH8GoRvrAUvdiEVKA59dFgSv5
v5lDWRXnE6/NaDW67qLJBfLVMQxVVCC3YHj5zK+z/AEj78TJ13yIU/Uo1DbsZJ77kkP0G7JlCnyG
zgUWa+VAW+SPGVaH0AN1jyD4uXpMZ8MlxiNIawawICvtkbAfY2MKPJy29fra5oWsyglcrv9B3MQL
z2gEdBflQnS6IQIEoEG2NPN3CfZGLGOnoZOvTPSGOPgLRjtzzadDB+7UXZ+D6pMfg9sLzuSodhrB
gGKpy3y7DfAz6AHRDVASSLpROTuz6UvFXWzosffKMviNK5WIrhSqlDGOa4hBwtiNe5Z4h9G2MVn+
NLWEP6/Pzw3lVC2k86lXBzugRE9Yd+Krc5Lfi0q/WzOA+o9ge8TBzHRuDraD42g6B2oce8gIssP8
fGDBg7uCSAU5VfNDoIAseufWpxbL7q/F6IKJQ/8MS4cXRM7OR9bmDRykmqYjy0BXN7I5Qxc1p+St
iWoS26yJob3+iVyqb8SL0SdIo6kQHL9cR1m6CucGoM0ELSkXKDgxf6m9NLYLrGC+OLNfkdskH//N
c1iNK94nppu+YJu58LdG2R6JQouxkIq+vrjLNMX/Av65K3O74tnsOczGYfSguiH/j+nuoGUESw8T
OuRVvPI1IrbqLqzv612zhsGHARj0OvTKX5pk3XE3F/01BXZ9OXkgtFZYuoagj6XmFuBjS2MlskLp
I+ACBwTBBf83FJ/HBMDNbWgsGoKQngR3TGq37Gvp0KPlwP/PWu79JUw92JAQeEgcjUJ2tsh3+LYP
rkFayrUuBnviQ8XY/Af1oztN0C+cbEV6Abqsy1dcXmLmQH2GuMBZui0gEVOu+m1Pj3RzeiAmKH6k
X7lt3zBlDdxWHQ8syfgymCrR9Fv2cpAjlJ1U1c03vm0IZA51Ysjs/BQbKpwZGbqX4l2JDHqtYtIy
IZs4e4mbiZ3EBY2IfPP1Vha7n+DShsgptg4KbqbZHXUZAtM510MXkaRWzUunz1gUbLN19x83pYrN
tOkofNPPDei3PIKm6Vuo0ydlhMBwM/iGZ48UgUUrvyJ4E/6c/JCtIz7+SJ/PPwj9NMeY96o232gB
gzxhPHGha50Rx5FXfhv7UXCT2znGO7d740bojxi77FJg6eojCdmz/+yB8owwOaPeHQt6pVoePRoE
CVOEq4DQ7mZcgxhQhJR+DUtX1cfn+fgySPLdIgMAEGAptj7IKQqU73P4Qkwqe42UX7pjNpSSPjaV
1DHgmLTqZyai2FmsQnwREWIKeRzCl1727FiyAL+91VXDqfB1Ba5pPuZ4UTGsJiB0FRzhnvPs17AF
AWhFVOPulqSVsMr7uQSvifL10hHkw297ApKia28PtTls0GvxW+AD+7WYYiRas0gsk38Ymob61TFW
RsUkwLgRHjpb/oAMrXSeKiyqGTfYGTnn1BNotjiPfm5j9O/gb71Be03/pCCapjfXwam9l/LwOsGi
sYe8DNlGRFCV7Y63cSPXm5lmHuvt678+h62R/o0adViIjkBglJ7PURm4a7UTv2zcgqmEnH1sssNb
Y8oMvK6+kyN2DSavvHDCYpOjgSLbW1ZYn/hr1cGdtZNM6d9BHIs0krGQyrou2ehKoFzMXsBMG+uk
otplyM3tAsy4tCE/aO+pwzL87NNEZAML+NZnsZ//1WF4NV2DUtQ3WBUb0aT2JrMevnOpGenlCpAK
16TszfAOFL5Mbw0io9F23nVKim3qDiVdsYg7tozRJOEEqM0UPeI4Q4C5YfUrzsTPAYX4xl72wFk2
1Y7g4m2LvyFL66kfYdsq8b5JNPKUoboSeG5UK09mfY5UUG4rFe0wmTiMmNk85zjIWef147C/z6WK
pbsI5AraH5C5Yq95304Yq13xaqEY/z16LqNZzE5BRJ98akfigekS5M9b2IpveF4u92+I+iNUW1sV
xjVJKnieWWCnYe8MzIRISPFNRK3QylE2glgvURfAeJ70TfF0t+UszUjSXDqYoVu0+mIKnXaoFWpB
rvYY1WODzkazk3glJwOenkDJDw8IF/XYiQ5JsgzP5AZ9aKmxmDGZ1p74EXDBgeoHUWRii+fZRaGC
avTaTurdPdCB+JSDzrTxkQK4AZokUjZmqjEjUIuLxBouDp1U0JXh0MITgq7IdvKuOrkHFqn3EbPJ
uxK9icQlu5SvdpIcwaGLmxB6hIfExWZE5b6D1ShndwW/pNoy6uWqJRl8eriPI1dDAnIgmlMvpRJT
+Akf1RbkUqNWjTWhadhUTDHfSxEls+PtrfmWF+pWel0uZ+WpmIL61G6oRfcWYqw4eypBstITWlec
oqzZoLzQfAID/wwbSxetGpyx4fTJxo38hB5EmD8EOUAOG5ZW2tB6vjx2rgBeqDKzBDnqhgFpaMTP
Enzu56/CM5m9j8buSXOh/vRr7Uzn6WEvtWrlTGgk2xLN0Njf6vhTWzZIj46eHgFPgrbwmqtb9DEJ
bTfx7+GCuMxfYjFstCg+eL0jHlX2SkyiacgnV/a1w/fG5Y9Fo7fPF43RvLJXaP72+x41OKhFCIbx
UucQtlsek5zKW4cw0I+g6ZT4CFW6jiJHB61Y2Iuu/W1ef+ac0s/9dSvvoFtczeqCLOJ83ox0Mvbj
SmBZdYx3Juy7K/26WDUamq78twpU3rRew96pFGDhNiVQdVITuSrGuwuR9EBDIvDB2qMbaYlT61dj
LUlyMltCSd8V7DKUwJok83/Z+3nvn6sE3S35H8O3/ohv9cYjJB1EFYngPyD7Tb8rtL1KqXRDNC2j
Bhtbck1V++El8EFK2FwsYV+XyJKPqxkU4OOil2oN/2czo7i/UiiAU8vfbdTxibMqC9/cNgEuz5xf
nK8PWWjOnOtYymCiiDiUNV1I2afcgI3hs1UQLtMA6q8LycR4MHdpi6icSn6NkpedTTky/kKMmXMu
5Nc5lVdzj2Jyosfgv4C72DbIcecRdWfGNXzMhhqfZ6FxZgI9w7GzHy6rXNI78w1ADzlVs9i5i5C4
+V15fMCaqVK5xaz38B4KKOf1je63l0yZFy8wv254lL+FHTTzxz3gzpjhnww1x+cLpEudEpZ9IgWi
SZ8ZXNPMF1EKKxNMjTg8algNwSt8JTfpnDxKbplhFKN5XEJQ6/ETr8agMn0ODVmaam/+B8ynCbo9
GfwkVLK8W8gsJdWTUtm8JkLlUEO0mqL7PLaTpsUHWTK9VFYhzWi4hZYh8MpCSeAnuAmQDQpEDJGv
HV1ysXwEXJg/1kfMH3H0JEItrjBBuxJBAzH18Yavgt9G21Kta4L2Fi9fw0BCqGvbllEE7mLE1Ms0
/XL2pmmGeVzUIgLRjKYf+39GpO4GFcllXt2P3tI5hL6uJZsyU6hY7eHbhJymstW4Pv64UbJbTmYJ
v5z1T8pog/F6SlYbfeRRBC2CBWGnYEuiQZVhdNucYYsSfu9czOTYi8tMRFl2MEdbC+u65boSpLAQ
yT3Ssds4iumLdBgJO7ZP8N+vu8eHDFWySrqoR4emNVB9Fb9VTJYF6QHkp77fHb6TiztZ/hCkwHwE
mk+nzMTLSGx3oq+h9WCt53GGWyziMVIzTZkjK4fi6Lni3V0sa8O8J9zWRIyjCGAe6SznLNAvvz+l
LivgWgyDABS5LAXZeLVTJ3+DGHKy7iqtMOSt96u2qBsTWsHhMQkklCsXzppVA90bNhRvltGXy9Gt
M9Y0kxz5+ZEIb2f7x//LmsLSOQk6fQ0Y38QMu44r02EoHRjRrFvfDC24owLxXgw6iO2sFn6hWz44
JrHfcCucIX8FdehkGsXE7mnWM3nXCOEHZDYGsURlStkegMSjSCuFrCmVJBptNnig5cFfLwS5ZjX+
WEROnu2FF4BdEe1gukJmFgSbYLu5fkbS0gb/m9b12nJZZZ2jiKsmM8Et0r0ivLqAtzM/MpxtDI6/
t5R4FdUyHjVgVffuzmJ4Eil9x243KejKryxgDici70vFQx/JgDUtyVSQfX/0y2c44RQOd2lz4Y96
N8HFwablA0bLpVzWfzPXVi+QNlHBtLyy1HUH4UEXRghgPOxJrvzkmX0noWqrlF94ISIxj45khZd4
68jNwEZWclkMoB/hQNUJAdcCFENOxONqB/WkY3dJ6VWWZWAnkqsMyg2b58k9z3iBJ6DMtYq36rn3
Y3zBUnnsuOPeysvdHh6xx9NNfNcJcDvC3Ba6p9UCI4gxmvSjjQfrnOJBxrLuRqInD/AF7VjmoQP+
cyGCVolFtM/C2D8AaW12YNSopcAYHs+Ww1ufiaTJ+d1/aKox8AiA8EdPqmtT7dKBFuBwsU7ljhA3
e+gH+ZVyt4nGrkJwvKVyWmZEayzJawByAT8LalkmreLxAd9KvZRzXZmMji48tyngiaprZ5wbHp2y
YuFtiwF1E/QvdBJAFrja+JuGLNIzzscb1RKqaSuw4m1oQOnWLkLSTonuisz4r9x0ZVNDGuIoCegd
EMyT5eFXx9mYEyMOgb4k4dnFcTRagWA2Wxm5Ds/yynrh6eUHaI/8YGlfMbf07bdN+2lDpAGuw5op
fAwCANHyyJ/CSeO8vC04T80G2gZjARupeA54Xoli5mn/fXicBH9kXwtZT4dGEnceO1hsrs8xp+Gf
2sk/WRhIqsoswrZoS4Pcv7o4ZycKSrzUPlN4SLVwWHsP2wXpi0o0ILPAY+Zn1058HOBo61ZJsF5y
5rJkytoLfUF5ubBCOj8fmtHNa4qPpf9qLh1f0vsVkP5oCVflhHESuWUrQIafjuaHOvbDXvf6076O
eTFqnRDbQxs8ioYLBKflH/b3cvg8O/i8/q/4bALKnL0ok8lE3nYUzAfNPXDE+XN9tYc+vsb4Y4lf
2vdcB6liiVIH/OauuDImM/5kthHKiuqdlWMJolJZX0K7fH0Osxh7O2SkcBLsTt9vhENWEPvFS73b
+K3U/hO+2L/eHPVtZYKDwcFsqF73Xk4lJPxTKpxQoFtWVsKeLsTD+XPmj+vBSBNvKRaqCpUXBZEo
VzDvX4k7+xICj0WYRCyPz0cn98cjk+ypEGvEsMEW2VPSF90cCbFT2iNJ1P5MeozkYjQbMshuhC2O
S14ScBgYXOcwroC5gwLugdRx/J+M2JigCfJuV8Sw+U9RnV9QeTOeUCxdr1IaHvSTMD8j4vrc/KzX
lo3wzUzmuZRZchB/1TEe2JVN7WopmWafJlYla6za61+rShYB/tseHcW8lY28MlMfdRi9+7VyU/ZS
oJNH9RR1F9U8lrtohIYZNuUhrTz7hepWhJ/uQQgU3l1ffigbEfBrofiFPI4D+QBHGuie30xiZkIE
AoryID+DWygb2L3rJ+XC8HBiFkXzPUuyiXc1qkBaQwuaz1FP20H3baF8hnfaq9c9FDTlBC36JdaR
9xWR67ENdj9NE+tG+dYzIPxo1hiRbb7AMVIpkwxxu7riZaiU5CiJl8GVyXdXmS0vMmVqlvN5zbyM
+wdWWjjmbtDnX005fr4ts/TWzan1O0lExJboGvMpzeJEtpPmmQQdemO2yn+/0Lr2NEYCmeqbGHGg
pRTRXCDDml/aoAziSFuJf+HCDjvNhWNF9t/TVXCKST8JBTQCravr94v1yI5fJGpi44/kdNtsYPoi
+iEHhMWvrzIwTp+j3kMG7RXpfncmpkqzTsISzwvvy8NUFETpu7XoMKPh3g7ovriLywLOLyqrYpQo
0QEtgU/etrA7lgT8Pgx2Xa4hm1KiwCaeCHewJ+CpvU0aGNkR1NoDpvoCkIkhtwjsu6q9PS3vxrSw
u+SPASfc2HqtpPqHonDbmxFwSPAqnz3ledHdUfeBDQimwYU9mdDGVVVpW2O0oTZ78McGtgdq/KTX
VYVVRN5ma+aAZmpxVA6tQeJCW14Lk2GYPCsmgaIbdqbyLEz6SaUBQT8mWHyKPpRVDYxnRJP5kNda
wfjFHlcLkRbr+wkDqFU2AkdvKdvZX/u1FjXAkHe+hP34EWP8cydnNh4tRoCiTzsWKzMo5eTfx7BA
JTObH/7qrmbu3fPj5btmwjFsFucZS99bl3Mo7N+8/2cNzI8XK9VL4tpNn8mz1wt+zj1jOzLxupmp
/FKpoOubfv1vpT03XB02CTm9evlu2xkcl8BtJ0ErrcaLwZoO2upn7/89482n3I23KfwDzpzCHuLl
NaQnDrtEbCiGW5gQW+fgCc2EjdgPg2mHjQ/qyo+iIrCvGbT9nR6C5sjQ8ODPcOfKfem3MN7BaB0N
HP5qNLJgOzzC6rXMskGEobmYNWFqBKaUcsjEbTeRHZEnAG6siFWI1Oiv0JyYIMzlnnz0134hi/2q
/RAhMLzY/fqbrpx28639pwiu4Gy6EshSNuK8mUPEHWAC82zrYuKUTLzespgWds4L7UFxgKHgvnmg
oqXIopxfMziNleZN6uAdzbaCBXDKCabwdmDtAxZF6jhvbIu91J4yKuKDJJbqxb+q5ao+y0lk4JOI
yWVqmyVUHI4ATl24MGngb+m6yCX4q8O6sVT1gTq+vCKL9qc0XMkgxcjRuzW1etNaqfwKYjnPyEkz
6eKMBTSt/zyjlXmdCsYsn+5E3uwFkWzh8uAn4dfu6lHqg34EV/e2ocYdQxRZnLW2AuF7QI9sYYet
OxzJPgNKxQ/BqiiX4iS6hLe0pZ+g+nVxkHyeo+sENP83iCcnuM87QrOnhlobT8u6znysVGX1STxx
GAiHc/sI3HUEoiv3vcawrTKPh2M2VNyzxWTR3qIs+CnlYZiVoJFNQZlH0IsaCbRbCGhf2e3IRNTN
Igbz0CHOpj3GssJWOB+zm9JXiZhf3S24DkM5yhd4pq+49rRF9RJGhKjzgR74jQ8FGbYWwNRnMiU2
oktvzvt+JaqCJUQ7vCBY0fc25LJ9UwSBnO93UFOg8+gFYT+GaR7+n3Luck/VRihm37t2EEyxbqM/
nYVqVfO78G9tdXPsizcTPWAvpxuu6kXbQa1QCKfHnPGa6/Ic8Y+R/zyuA3Ypm6LlkT4Fxs0vcXj8
FOHmXqMO3PwwVrs/wQ9uNdDTudYI4jy3xitBsot5dRChfDt7+icrBsE3FmV4hQu8lDqL3X6TsVf9
0M+eQbtge/UJImiwqpem49Ab21T59BXpGE8Ty1lS2O5WCOksOgmXcm0gietCiqTLOw3Z4MyFMjQJ
kfLSIHs51NyQZ9BNUpCB1xq5+P38nTw5Ghe0uZdRS1gNkrDJhN7GIwvieRc6HtXnezO2cWI5136x
adv7A//Z/WbmEUC0F6pSw7i2O74fSt7AW0ctAr/hudhOB1CxsOdxDJi+o75IfsZfz/UOqCDHTOZM
Z7qr13njXGeZsAWCCATzZDbiJ8nbSQeMUVW87kISFOLrujXWcfQ8/dWXbCLUJ2vwoBTx/4FGExPC
8Zsvc5riB38NyvSHJNZOGzeBtLxL9epFJpBjNCdLfTi6NsRYJU6Pv22yAhmf9xEBw6ILkpjQ/3vJ
K1FwpM5kmqR4iIipa+HTmq7ec8rOihmFm8UNzNgpqzEeZIDz4RqBT0cfYIqeDGNB9myhfYRpmm34
9WvrQon9C6D18+WVNuVmMgZSBTqCfWWc3aAXb9Ub6oGNlUaw0Uojbth/m83u/dRbP+a0nlx+MiBE
QHA/sJLR5me9YDCCtBCHz+kqINliMovJa2H/L9bEHAVP0W2WeuSG9zx5v34V04RRPt63AeUqCfrq
UUojokOyjM22HOPSgkbJbdZZp9+WSPKTDJWYQ9S2bGYHhYTY8SwmRF1/HXoQnzydckO3ZxcobBhC
NY4WpRCN/b8dd040CMS0WKyEsuAw0IgvebLsll3EQXc8mRN8gRi9AhDa4SnwPpBtXW8YtaaVzNnS
BdNhCO+fOnBwKdZMSUwlwF3TEb3go1nd7YFR2GoFKdra7RqLB2cill7tuLjE/tGaB07YqIKWPUNr
y//jISvOwDMm1pwgh7Hkvf4ZiWnrYxLo/vBH3OOSsuZBAVrQVNnq5OC51VT0h5yWTvRagIdaAdbb
rYBPoX0PDOHGlvPm42gus2vJDi9zzKJ/sgHrTYa4LbugGBzi2NGExLNYFDgu2KiLAVRocX4q8Fzm
XxHkoN9t27UJsZx+2ROSMPyRiSFyecP2wl2HqZptCLh1WMeaaPZ4BleqpmvKWzAsKA3uW1f2oH2Y
G/RT7sXPKJq7YRsvVYofFceIEj4aIpVH94fxwR6eGU3PAMd96+kDeCYXlvOTef9Sylpgaydn4Y6N
JKPF6CQULK+araaGQ487ObfvsG+W/t7MftBRxXXWo7sWiplI/bu/FwoszHM/5x7Y1dYxK3XIOHCJ
5b9wirsyq9+NYgsCQPK4VODra0nqCSTVwdkCuOFDv90BD1nFpaawHc4ufi8FFWiPTefOjbwejl4L
497jnymdRUT4yweEWe2zqb+eft/CbY+K6Ua1+yY05wz92NXWVR0UhBVojuz/BqPrvvt/+nwa9u5Q
YuU24SbmTLGkumKICtgwd55pbc7HizXPfBLDRf4YGdkoXwRoO1fEJHW4ecMcGv+7MX6yDLMrEc+Q
jqQoPZbWptVAdosdIqqVZ3ZW+IqDuVvok9cRxUesbQMoB58bMu21jKW7VIxyxkaCXlHSuTOSh2Ue
Q67Pvet4Z0uPb6vhwirBZgfDH3Icyv4NypQ8wiljPyXsL/CoG6teOAYByt07x7fXa8ThyLOE28JB
RiSWzuFxDD0xWBdceRXiiggbJgBXKyZlWzTxHN71BG7hl1DunJGJXeoKIRNzV7NNVRq9m3dhfS++
wWlZMH9F8Eda0RC21gOCZlt2eSEZw7NUHrFThCNuHjxzPPDyzhVgnMvI/X0+SfcMEnM7pQl5VD6c
phGOjp6fi8ENXTyIeO/2bU1pJy+OVEftiHe4/N1TBg8IFKS9XyjJg76BoVqTwG7mrq1DUhUxJ9Pf
AsTX9gV2Rkl5n4Qy6TpCWPgDOu7ZsVHxvQ3nj5SWvZEaPH6saS8QNN/khVtVpHTNgoLtayTAK6D2
pe8AVNJFLw4u6Q7nMfgJ1AYciFa8ktumr9p84DpOzGNiF39JqcUszTuk4LlMLKwXMtNWKE8YDshp
XyI8tXdZXy1fm++wPEn3Coy+oHXwSHvfhvo2gB9j7bMuKXBOeKNtglMKknhU17OePiFtEAHIBgyh
kADqadf6enwqewyJNS8wlzLKzmICH7vLfXZZ4yug6Mx46SdhBweZt5xrEKP/qwCOzgLFOdoEP8hm
sJMixFZPGiGDxY7RKJGFu1gQJS9mmBVo4PHPDQMraLzGyrV8elInPUq/rahZWLvmbvYI+33RDrbd
tPEXBCjmsZfJn2GT2DzfaM96gdaBP7G68CBunFOeRg3LEDM4q8KFZ+dGVddaKKRXfYUogILCLf/6
T723FjeuDREib0BbBZHGvZpLO1K9VR3zLTnIMe6mocfZcA/mk3/97/RRfNH+0uI5MO/HKMxPtibK
OsTzOtb9bpuvUcbIGvncJq5IXh/42ZSiMk5HCMLHJuY+klta8QcGvtJXqI9YfXXk9xgtc3+lGg+/
A7pVgaDDWAc7l2O/Sc0UHkw0nylvZxiO3aOkZBtZlipSqtwLZhSdjL6g3xZnDLXdWIQJeDLlbadw
w6cALqQ0Lv5TZp/Uj/EhybHNPhRfZXZtJoW8qG1XQPU+dMmFrmmv65XQXW04n95CKCRfUCsycRf6
ee0iSqiLFZJFPCABW8Br3G1o4MYH2KZGwCL9VbXMWlI5TABVv+lhu9SF0wXlMsAIXAgfQy333D36
hq1Ywnf8sxs4HsL+chKcV6cV4r/6LFLnR6p22DIVS10vVI8rnehWG00TB8SYpxmra+HANLTyWZKK
UFYC2PLDmWPREYozIG7dwcRw+vZGX5GK0RFO8drbSrvBlbvG5LhpVrX63UMOfz5vZacCIAlT2ogY
iwNl+nHDrQMg3gvMbuxp8zhQVgA00y+DGZAll+Ic0QmmRsNcomPIo1OzlqVz0wF8qh0xTI46aZj0
N97jMHeI7UVpVChEEWrgBf7bUqDHshkDoG3RUhKt3kFKq2Yzkk5mwMuPnOB8AGLIKYqY1WI8F4Zj
3eTyDBEUyaxQqql0lheiElscwxAfzuFvkIDamTgGZzPDWS5TtCijrrzs19dXRtXBZwz3Cj7MnSQF
uaPK4DASB9FZ4EUkUwQfe306mRx9ovfddo+NEImLscu2YXPiH5ITn8i3XJ5zqdfRP3NbmIc7wCUW
aK19QKF/8ZdLnxnt1RI5P6yMTP58rEmKgOJKCjFI3dzqiceOXAf+3nMZ5ZUFUHaR5LriXYjNVYT6
qqwpOaxKyE/+vfuCbvsIhlFrCvKtn91WkCBuoCerPy5qex5kB33HgeuJMaqhyhOC18xtzGMgQlnH
6et+4UVA/OyYRNh4YUjkXWGucyv4MAb6dtt+wBaoWHpIffOQl4SnGzxkXtg1oqD/otiyRPKJ/NbT
9mhjCH6rXtD4E73qVx/Ckuob/O9e2PLBgGPzC8zAlu5uw5lsg0D5WL4QF6qnyc4maHEiEdj0DSbm
S8EXOr22xXj3bvEAmq7imEnCRnEQXtLyF8BJChTNEdkSUlpAnsDeYmrxQJnCM884jrd52X4MSsjB
azvNhZ4cpuczRYdB5aaQ8HYJfuv8ncZWdDtyQDmjJnbrdAXPXu+k6pwBtNGbHsoP3b06aoQvfR3c
QQCG6ICW5SkNjA95lrfjoXIUFwH69/KFOmiELn+24zBYTz6jV8ASPj7+wUQsxDuYQnsuf/4ZOall
z4M9bfd7Artza6L8tRlW78eaLgDwph54zynrpu/G360VMwsINVxr2lHGTIQHLlTVz9/JXKaHQ8xz
+l6Nq6dd0TdrQSwNuBzjyZPeNKheIL8XRR3zFoJ9AlGfeO8XIYFwhq8JHW2Y1zHTn9dv7FvKTAbX
3xMir18FS57r8hUJQyAsTFuj66mmp1MYIvwL0TdEV2V5Q1NNC/3Oo+Fe/gJXjUuWi7QwZ2Pyw7uA
RJTdxylRyye/wI2Ca8MCSe7H1E5hLJaS+oFCt68llXVnvuJAjMADPxgdTFcukS7Mbb/XoXbNMHvT
mF9A3WZ8dpmpD7Wo7FuLN+NehNC43scfS6w5YZf82Hifoj1+9kr7RsY38aLE7ABlswjDo8uQBium
FQSTGdWx8M0NAK/q+nXrIRVBEwu/LYZ1xGEyvY6c+rllW57wzC8U2S1fiPthdpbarY/WUqiUQ9Qk
FMw7Ku3dX5nyFi1TnIXZzUCloe5AJBVYetLq33cNc2KZsppV9jBOsLPaBNTGfuN6uV1d0vJUxPX5
DhTdY+iatRFG5O94MJzQ8HY06z1qhHIaJmdVPznO3cGJVWxBznSU5CcGJViZMa3cA7CK7cFXXHHh
8tyJcEdUAIWJIcf/6ERAKPmhf4JTmOJd/VXcHM8W9KdD6S8mMObGrGtp6tkbgSTV6CvLJE7+Of4s
bdTlofupVMQvCk04zaRw6f7WO8fGv0ScO+6ChyyLhO1SxALUWCgpGsN5K4U2eC2YpMNxtygaS5jG
hSLQxsg6EZFwfrJuoCvTKgkHFagj3mId2Oih6StIJJ07/P1cdLrIBHwkqQmFe2hm0ZoBX18HVJYc
UxVcWPpzhIMb/qIqztAXDksng/efcfpAR3JvcCaWX658kDD141H8NU+smIHHC0tye3rdI/FrchFA
qJX4lf1YzjqqaQHq+wmwEco/WYfpzfxIfaCBjU94YNW+IypHC17Dk+dQaaJnjmTH5Uz8Y2tCNioM
AQJae5yvKxWeFGTQYTRX+3Fl+jJ/PMrq4KRVwG+Oa+4CjCbtG3VlGMfLJ4iMqlQkZFbByX0YzaqL
AJTBOyRBEXe73hI7Sz+93uPNuNvwQUrXjV+LqZJx4uSed4Eafr5/hbFcrq6ZEQUv8JpNa4wc/O8A
bLUW0CRnR8c5LuATM3VlGoPQMe3s9itLmlEC6zN0ZG9hvVjC7+agNvEIYYZyHMBQuJwT3vHQTLQA
IpXbd3eMdMq9SeeUaIaqPn5cv7jcMqmwfbCfGEEPV2izML665LLV/NftkkeNOrOXG/C/fUkEqjvY
0yY06vsl9LMgd2oP+rLeFBB0SPKzdPPe2JnBVrulTEBzl1McTywK2Zxd16notaCTycBbVewnPo8g
s9SIE1yooP0AQ8UMnmE1eXswIPIudHJC0eevO8wZiIQU3zQ00souptQeb7b/VbimdzzDRHMfTW9J
AaT84wj7tVI7/WespZZ5hAV0LHiM7wKv2KhsVY9+2oLhspdKbtF+5C7JIYJSRWagmiNMigd5+fow
yGunVPlOXY/1U2W+Ds/AvgEYp6x7toDSvflZcsgL8ie793ptkatF/zu/oHYXdlcd4fBVKJSQzKpw
YFpb6A3yJ8zofRJOQj4qhfOxgKA+ofjoEscyKD0lNJPUqlVSe5MRhb3xr36ZASgH1XrWiD4gD25Q
dhN3g9tvGyDybHhTGYy+ScjahjMtXhvT5QE/a7mhepf/AGMBpNlpiJ8c3ekvYxa8CE0fvpY0G8jw
o/EBZZkaj2ARqsdk2nQb8zTmpecB8S0ay5/CgZAv0i5hJiohve1v9Z9jecJStag4289UbY47mk+x
Ix7l2lAcaqpS12T/8LDfl8i8lBS3PMzplBVnAF2d2ArUKn0waBlBvaHbJiKrDRO8h+hppuB8PQXp
zkT+rUa3tLSX69AVsEN/qi1OK+eaFDB1uyIttXHC1GxMjhSAEm4DFlnrMoUe3WzeVMOT1YtSZbIu
B1r0gIKF8TgtXS7xY87Hd9/SSo3I2S8TKcegG1hKP26i8Vl1fOgcuRNCMVYvYsI8uIkgZ49uAlLK
TibN8cH6Ze8Z2gippKqXiXu9NV7CwhwgxsvZV5Kx65UezrxtzT0cmq1oSdvHf7BgjVfByLiN1rop
TIHHKuGt9biLL4agCDBWrtzy2tv1hpD7ZNojfkQ7phjRxpmSSY4Ntqg0OpkCnCZh8e0rIPMu/Y2h
YAzAN0dtK4dIZnp7gpxuXFBxll0K1X0j9OWvz1g+c2TtntABwXQCGaxlKDBjb2AmkZqA9+ISM54+
TIGh+izPWyYdnPCvliFg4FfYY0a7ng1NvAbry/bp/U0bD4iKpTtCNad8QLyV+zvobdyAJJbCRjHd
EPSoR+4fVyC3pye7VwVBP8FQRcyK3hro4JstgtMpTrjycS94liGFsG55x3BQYuMkBrrMlDv2MqIH
a6ACdZGT14HvNLrc5+ob0T0xUzuct5aZwWMmWAtJ5DsWKsZMIy0jUCo3oSY5rbmT8gxjhVk+XtB6
YgJOaIYBnefWVRCAcyNPh70D3ujBXVHyCOlR63X4r9bBjrfQMPMrWkSAPlVQUOorCJxmG8lAJ7Av
OipRaIpqym06RXkFQ2txdIbxnPdBpWh9iqtamnQDcEfiS/fV1ynbZjk/es1Dg2Xod7PNALKdfsOU
q5hoXWE2uptEI9jpKtVgSy0vz9tAABTR/io6UnZovqcha1SYTR/I/HvQTIv/m6nKKBMhoh+zrsfd
vnzb2EqZ9Caey2kFHRtyrBl5oe8eMuosTQQtVeF71p8Xzegwfe8KCZa7u+JYOUwBMuhwab/jFyyN
ovVSdkmBwmx07O7ywariKeq6KdVE4sPMgIIEqWQnooM+YHXfCwUVS4k15BcV5ogKTpUWXUC2CoEw
h+Stusf40GExeDc3cxblrhZQYID6k5XX9kyjEG11TyM/XPbAujgapKWbxDeCX4ffEhcIkihqtwn+
4B5uhRlF3ABLyRjoCUuaarFM8U/8x/cfC9bwPC91p9js+zR1bojODQ5LloWeVg/7AQ089FNLOSDE
cmKZ+72Dk9WZguiAcrfZj+hcsPh7e/rbN8irQSFJgvJmGX4lSA0zk64WWYKRaEN075Q2dszLN1ne
/IMIh92borKsxKRueL1ri5kKgq2KIgiYsB+iQCSGTsPH8sfLQhw066w9ZM2yzEnr6t0hrbCk0/TH
O5/Dd+2//pu/HWHs8/XRB9ckk/UKekf4d+c2szqA+GIMv8DNq4+vWOmMZTdxiNF5TR3N6ZCbv1Uy
QMgGCnbBV5rM+I8gnvB5UX/EoNYmss2hSmK8z0heNl3lgUSGnyuVjyDByATQ1SIQ2p0/dip1GXAw
7smmHUqJAv6zS9rVbS2uxUWwleRsvKVj3aZV/KTkOg+4SpykVvPEZxGkyjVW+YNBNX1VSG/Wih1e
CDOz8E6JJYoTOf8PJDBtudBuZ9gXtoxJJU38gFwRsu3DCa4Xtoo8BOnYIISlNXaoWxGr1xRipFYb
8HCTYHxzAAKFCz++6piRm/4nW2mOimAUEC/lDEyn22sAAXqGCLvF3fYNBA//aH5HH4TAL8hPu59k
V9hDYEkdhqTiWB5r5sv5Az5lY82P1IrzhFGg+ForIuoUIex29UB8sJIaSQarTABl+/cPuemZsw9Q
MxefcGrGqJtkitqSFkAQCVMrNB4xpCxWeDfjlSzYG9wbd60DPALRPTQojipksWhPUyUMR3rmz4wE
4QyaLFKtA0ZA1bwkkwAxbit1bkH8SklRIsCdv/TgFXYahwYnRso8ygF/cJ7ebzN0Bn6myNx5oeCV
MtmzOl6Zp5twIdxR7wJobwGArqoC/y5i2W14+kjCZxUulb1ZAVqWRf0caNyJ8VFG5EMHpijYfar4
I/IaEyKPnyMGHoBRyATnoG6Th0sNaNk1vagNpMinp4OyxA7CN60pPXo4Sw0ZG9XWJKsLzCj5FebU
s44gjbB/UFJeBF+zsjI75rFugQM/3ChE0IIyr/hc9hyntUCx6X1hDYCxJeFwp+8aXEc0lCgYc3hU
VQPK1OsK/HWgfNkDadjbxEz4x70GD2tDEtshgOtBeo/l4e2iZuFHzVRt9zMT73Lg7egwhJGLhs0p
diC+lNYqD0C8JY3j6/fa8M2rRdGluQCtXKOD1vgHgEE47KgNKwU41/8WMmx3UKSssS8U+aqDkJW3
oLzvhLE7gSDbVHzlnzTLlzWrk3aodT/kTac3jX8b/NUnryAMOxiiv22zYhE+Muk+mNokCYWx8TPv
mhv7s3lkY0J35rtZIV5kTlGgsHjNtWJZ5MDjBYhrHNa2Z1ScigifGT7awdJuvQ6lA4xQoHLGrauI
mLH40rmB9GmTzzhJ9tOTumZQxilqSTuK4cUUxl0WWKr5yri34NhFvCrJoCJXo27w5X0dwE2/rhY4
Q0Fh0ttJOcvzNtrTm/gm+jMBa1K8/qCk+bvHUDbD6NyKx9mr1iOYOKZhcuMJrktuOnPTtmcgKLkk
0aiQSYoxQAOOrY6Ch0IPWce1ieeXIjGHxm432rff6jIrJKpOmm1D16BTYyXxALTNIaV1KFmiEWYz
wd6Nx/8JN8+cPNN7DELKPOcMkauFf7+2Gr+72/YdaJKbhP/9zEMlsljWI6oqkradL+kDDTd7b0nk
o9bZxk9tkW/2BOyGocX3xb/8KAvF+CjdNpJtf2f6X6hfuI0BeoHP61X1UasNGJmbDPLkfD6km5zr
qy94e7zkx1xR4RuXzK8DvB6YhSz48SgueGlghvD44N/TzoYlWl4dHQ5xRW/0/7KCAiT0jb7FNej3
u51LpM6DwIlGsVX/VQU0rldnLUW8XxzaFVe5p2Qxex0g8FqAhE/EfNW9GYa1uHgAhmfBsoX3CcRu
WNHrTkvMrzNsmhTsUustl0wdbyPfxhieB2DN7L6b4JTFFn59b/SwLAbq9yO1BJb9SJyqq4bhG8MM
3DX//gO/rQ903dSGS2ZnvrU5Il9i45MNkQRp6M8sr1VI7LtDA9aF68yYP/6w98vsfbirqOEEMzcA
1Yc4YZZ9V7Du7qpSETq5BMEhtPycTDrAABBBkONVDB/IKowSWjAJVIP09HXA3JASTdYfl7lf0sW/
2ZFyIQESg4uCV6y3khsxsPhiWPePWdUhfW00Mg66YQyw+T6zVwI+NYiZBHWNSI5sofpuoZtmFw2b
RLYkcrFmc4cYd5rGiuvx+2Br1txDMzjBS1W8LEaqkw2yCXaLdgQvCfUkQmmX/auqwM3DEJeFtwwx
D2BKeV9uvYjB/LiNA8GPTL3U3QkgfRm/jxfaId/grmRFYO6MHBYVThEsPD/gQCHpS4XjfAmtH8Qx
zPe2FpWR1Hcy3SJ5dJ/7hJ5rnIFsiVNGm6ozZ5ZAVsX3kRQweFAAcziqS1dSrBV9vpOVdztTjSJM
T1efmxkhHcGEHFs326hcwj1WNDGG3aaftFvJs6aXbei+MLQmK2SYi02J3O1N+e5XZudLw6uXgMCt
wYdKuU8NYiX/W/WMMd86vwp+0E1dZDCLvdBdOqAaoVo2MbHImAsRXyn+f9MzCI8lGxoLSyu4kAHG
NjLS4G0Q+Uu9+qykH1diN8hmV/12JpF0rScscQShvIUiI93EU0KsA8a2qF0Ltgre67XV2fYG6xLO
d7Xae5qsxSSXRPikAb8Fa3Kmppcsd6orZAJ3TaYtADZYdmIl147IaxptmAJs/Sa399z+VM50JErR
fxi7ZNb3Vo1sXaDBVITJjAvC89CrN9qsB59u0MBf/KUbElH+VQAXRc4kUGgmwj+W1flNIN9+SXTl
Fl2khhtjwF7KL++BJV/RKd0kbh/4ZebayRc6Khhc3t84eoBIoYwiY0E41YrHEPK4QpSyfoOdkR77
E/dCQQLmZ2TSWz9YeZ2F2lkpqI98DE5PvMQS0Awb1Ut8Qg/H3iIYwpIKZ7qy5AMVh7K5ulNJkNUI
qS/hunHvk3enoQIvCNlYM9WmgF5LgwCVQ4I72FZpoc6Bk0/5l/KjLciNMl7/MxfolbcPG1ldJLZ+
5oymkzy7BjQsOotPmGunGhKeTFHAQE7tPoh2PgjYOugcz12cHrd5l6S9uWq0+CbfYx/6tiyjPwYu
U5NFzC+8NNfr9gTiKFU6pSHxSzHnYt61zGYV5uCRaKr54FSZlhU/2mySCuQHppugHce1Ng1D4IXD
2vxXRXwXoKEX90Hm5su9sRV/3btDUep1ZX11ZK/Sq3fmjETnCUiQbMgv95ot+ujRe/7CRpDqSjBc
06ioval5JW/X9h6t/wyCt1Qpae6dEy6z4+9OFdSFa7OeS0w0OsTiOV573tPiv0IXbkrfQtkp+YEI
A4sNivDfBRiGBxuxYB3sWgiLD/TAd4VQIQ/aflNch5v4nCypxoRJd18GnB1OnzLcqgLn5S0l97qW
A/4rqbwG1h79w5LQj4xY880pbvyxGD4wQAabqGtXpZyZ3YFlLKqC9MbTj2YbF+Log3EwZpTiL7rC
e1E+tm7asny6/u0TWp/9Y/NZ/HeMH0Ut/U2k9ND58HDJnAWtye+chRpzuN+8NG6e7hQ978sCYuee
clLFSlFO7L5QhQ2nZprr3DJqo6JAV1enftZf6vUniagje778T4paOIRCr/hXImVx88phOixV2DQq
kkcQC6SBojHCjBudEV+dZ463fS216nPWkV/KfJ8mAsN3dO9Z294IngmXdpiC+xDugJWe3Qxs0DqG
+mSA1OkXQjuOMYv7id6YfU51qprOKmM2Awtu8MG3/szgNhVQRVS7mR+6ZTJSSNLhGlqypdUyrJik
/XH+i29kR5koHBnrrj0ssCwhyMqE6pZPSmeOkrP934krpynyish1fgDtnTQ4HoD3Fm/TuSFi10hg
KtG5j5h6FiPHPYpdaak9HldWozfcfUfSwJUwrGKRr0PrVnnRst6DAIUjO7tk5Q79DqN+l93axD4X
rCP6IcJzUfZsR7dLZnhmCF6J94JWFd5xwzxy2B/zYU6TpluBnk6H0f+u2q0ZE7tH57F2w3cc0pJP
LfUDM3EQt/cyZnI4zAAJZ9M2Me3mb3406YlIkGHQDqWEj0LQMlayBBH1pwBerFWHKpbDO05iip9S
55SeTDeefeIXTKxKYBhlxkWbol4bJbM3Rir9xrRAwBDIUVnP+4LtD2ohw3yrffU9uyYzDVcLCsEX
SYrfJS7RIG9Rr5iouM2nUmtQ7mUeud65EPO7DcGBjTWNl1n2AhbVcaLUJVD7+wL/y5rP6eF69gef
WvAX0Rta86glKiItTidT1U2z5jS0x1ckcgjKJpDNvkdYWgBE6rPmf9CdklXaSFyOINfUxa23Dc5l
ReHyLo/4Pt/95vt3IXhi6z3VUjJVMjkmh5SoLbvQYvooP5pCq8Of8rJEBtMuITxZ6Jsf1GB7qtay
/cT+wSY5WA9kN+XdbccZ7V/CxMT5E54/xdAYCgD06mI6YJpSCXU6vqLrW6M4tEnK5z0a2wPyqXYM
S3raonfREcpxWMEFEr7dUteNVUnCRdI4ZWb5ClB3aDQqpMtnfrcVoRIaTeXGNPB3Ym2ArG6qAgCE
Pim+Px1jfLkgl+n3zqzBEwmFLq3YYpJ6mWxr09swtVyLb2PZL4rXcM3A6QR6DOCNifL53KknbgMj
0LS7LXeKOAH5WknuoEDMQDSfnyFd7JdckXOF/Tx26G+0WTIivDhRGzmDxU1EHG3IrpkHHTJDLSm1
9oOxeo2LW6jLTNHlFGTZGcUtpJQyjOHTu+1raa7OzmIWazdbpun7mBQ8lb24P4ponrTE7mcJFK06
Rr4kyhjEdO+f7cCW1UYWe1pSJrzv6sDg/6iZvCF3WK3I61pCZH+68xD4XqIFwhikmVrlS3A7iOAk
afIARZUC21u1s2tEonpCZ6nsXtjfa5uI1VOElYZDFpLUc8dPC9FRVTiXOOauAIiQjD2KOYiJoUpD
Tc9FEih6fBUjVPYjowU3WdzRlz4djj9Zq8JMDljLNQGWMmguF85tF7gFFfTVPEQ//Fa+vDTm+pzz
mn93V9J1nwWzO7ztJP+2XSCTg9qipKk/9nRQkrkz4Bk6ggVS8n0DMPI6doA/aSTjJGLj47y6pnIm
QnwEZC0APGfACsTeq6H6B/FWRatPLNYJOVgmbnlQFPjwiaXs8bk1/8elG1tKbeoyrKaW3gk2DZmx
d0hYLmNyp2xFJ87UdBQiVLYtxwTQYj4P/+oNr7rZFs/nB9vOuK4uuCOg5WmJ9zxk4wQBAphbzt8F
Tnh8ItaBKD1RULcSR4QNG9ZtEvl7r/lDr16X2cdqieDjWRgvUF6B8xOtkl8RsJH3DdGLOZuiZPQq
KsqcYCVhOslJ03HXyNmOelysV1FO0n+eF12+wgDhFf4WaeQFznbUeGKsVkVsMfF/yCzO35E3fH58
efTtNG1hCDsfjmHtJGvOwfCzsQoS8YTxq8/ze/wRfnAtZbfldo+ABe93TNg1xIgEeJ39cxBpoqKL
OcOukidSU18+P1dr0lwq4i65v6N5ehhlSkDXArPUNYkx+WnVBmQasCEKcA7LIKw5KzIPtQD/IUbJ
IWC1mEyK8AnltZJGTjlYfhF4tKq/dlq95xkHouIjAI4tv+s2cbkhTwXsEvpjlcR7MJKWJ/G+BN+H
KQoTJHszCnlPyuZxd+wuZ9UtiGKuYsgccvTpZlqkOIbjB2BL5v8DDWdMaUQDcXYcGFQ9rNZg9qfE
7RaiLvP2NiQeR348vrr7J0+FeuRS5dxURB/0yu2QUhU7+sylgmCREuFp4s3jFfqcuGFj814cyVG4
NtF2F18l/KhMRaZLg8s92sw8B/zwS3JaA4xpWmeUirD09gdQPCZ+dWtLFYRSK8Mhx7hcSOdlY7aM
D2oSQNArGu99GsCt/mm12znQU1xLerxKq0bYbqk9cEBtFtN/+8mUAWGeCe8DJxOrAlPfjHO+ftfA
L4UHokHePUvi9V2hq6L7jlEujID+Yd+ZUnKzjfH6EKFJb3/pPJYCMRAwNMfKGbf7V8XT86Ud1Pbe
sbch3kev1slt2nUVlEx93efQ/dmZMa/gLtbiu9eZ2Ee9+IOXWVLvqV6vSYdHfnVW4bVJQFG0cUEu
BYgRaA/ZLrBlI1E9ylNs5q4P+bS4EmAnsheM72jtLaKEt0qIedGUOnhIysteqJenqj3No91oAObR
INt5XcB+SeeX4WJV/F/8ja5vRQ861t1NrYbE5pUlArY2zVE7KNryKrfysNFvXDMUelt+qDjfR/R3
hxnxkmyz6SYBtX9r5F16vznnsGM7viHyyFMHlO3YCyds0qOhmWddhZM2i6q8sjjpl3/nl1gzqpD8
jLZORVM+36xD0keCR/ZEPrDo4ReT5NbvaNkVXSwgwKMCi/j+MZFsw9jd1LTUg7P5ndtCV5/a2XFb
tT6Ofv4lw5XgJRIBnAyDbSn0OzbMptdk1Ot0H+soV9UIkWtevbgx1BvTfhI6pZXNsIKZqf9/ubJ4
c1oYUc0TzXOAco/fdXv4/CbtUaW31LDa2oOri8uhH3vgsRCwobZfwor3RxwrFlZ8EPbCP1Rr91j6
/wn71XmsiQBaeWCwieYRSvJShvEHMPxycP9GUP2GAbH2o576bLdIZ6UfsPD8SN1z1m81CmpnCR+B
1yy6SQPaHjxzrZJQZ4IbKpu41IpdzFKBpYFjJ+F4rAYypai6vqpLT37ElkOGSyWbDgw3w5U0CoxD
bcxCklav0QZrTBTrJ2QWCQhrjkUNO5VGJm/kAlZS6c6lQMrsxiPKNcet2zL/riWVOnFb9zVaw3Qc
0p6D/u6dhyulMHJgaPuUpLiZgKCAh0AbePTwexsYjHOtKcmgRQAd3aofaP5fnuKQkSuuUpwBpx6M
eoVHc4BztqilRxU4eKwRVG1AEkpsiD5KF1Ini/QFFSPkt1qU5phUajb5YdEA5BH/cDzVlJ3u/Djm
uhQH5Mw3bmIg93jqI0YDAuvpnXW7iopw4b8R0crZ57vz5p6cORk8SzHdjrd9GFi3b4CrXyHq/Lpl
qKG3iQXCOQ59yiuSDHGtXSrbHoYmyh4Xlp+Yauh8Tp9maTTLMlDl6QRjmdoRhgv4GOqDRFiJEiKo
gyZUloTzi3oMrimDAKxOmW1HQJ+uEsUhq/ZtmgoSEumSqPeCtD04yI8L/pkaA08h+4wtgRRQlOV9
wWIYgH4RodX+bBm2efInQJKOps3L+rOtmJVcVekwhJj5lgkhZ0ToiPPTH8Ydq11BGvabXucZeR6i
BCMRUqo+a60xJwmyqftgmbrjDYis1CB9lZ49ulTOQTdxqgWT+8ykFCSBEZPAUmp3I3UoCdfB4X5z
Fmbhcph6HePg4BxyzdjGgpxTEx84SiHxOHccyOySWZOg61TwTeNdyWd1hugH2jLNp8SIUZy+lb7Z
raE6v+i7jkdMbO4uXuYpV2COq6ZNbFjjDhky72Hy7Bqn5WSWLnxyD36WV9uX9agLiZVlfGdYzk5n
IG8Tf0linNMCnzA6gasbtDr1EyOzELT0aNaxUO7e2V69yjfdgvOgfgUZn87G7SrtfySJ9pZ9qvjU
9eMIFVaK3g2RBQINYqLJAZPBt91J0S+0772muBPNVDUOjZO0m1crPxKhp0zYTJm4CPBJ/Ns5GIRH
oa2SavuANSGEpnNxCx97w85ui8XR7VthQ798o8Be6V70t2UPiU04aVi90nC+e3hAvzo5dNyM73vm
GWSvmgLQzI1OU4dA287TOnPF4Geg9sx5rMo1LjYkDI41OmBf7eitnfm+QJWCVoFLYsQDqgt17hqf
n8jnDPcG161lnWxe2IbTFvRL4dZkxzusG/aHKJrOlGoqoLCbF4sk7gelO71/R4U/KEv9BLDX7FUn
NBCHFDwlRmm9B5N0msaQc5ffvT9h7gviRC0UUZZIDpNLvjOAqXlMiNCGyDqIK45/PmJolIZk1NEz
8R1853ztQgvURAZHVF/jpyJRxdN1jlq18Dc/ytEVOdX2xqcckEjbeDt3dPbkXOIFop24PyGEufK5
meHJuuKw73aqWFic/9b+b/U7RQvi+0Tay69zyHg76GOQoydqGbrxO6MKLBtq7pVJ4QJdjPFdWEeJ
W02eyalSYB9FkLwkexo+8KWZbMiiAZoQgnghADLHaJLznuiQ2wF7Sbjt/v2kAL55CpZWsJr6+j00
39xlIUK5RqctZlUsyqa4absJ+/MEUSkpQS9Il9dSa20XQ4julBdBMt4czurb7yOXglFK5+afI1xY
QmJ7mvkrJi2rNdaMT9k3Fbbyb2SyhX1ukSgCicf+0WZ0om/6AtXVZ4GcxYDpzxzgGwz3W+3jwN9J
AXJC17q7eS2xj0oe8u1IsEp4aqEn2xU8vL4cM2gO92QA5/IhcA/3m2ByEcOzissPlhpqbzo9ny/J
NdXYYPnop5zwTUSsulvNum3YzMXG5qAEkJeGh8gk0k9sHqBQYTQN7TfIo8gUjH/2Id1RMPy4yFZL
kcOdP4nRw5ewuymg+/da83dXvSBxEPxLr0Y+n5lfyxHNLD53oCfNUjJKu+Ht5OlavulUVGcnH/Yc
1tBnRvE5fInP2paE1HZlFxi3MxmvvhPPIBTP0CEB0GE9lrLiNj0MTif9oFCMcft2JLzovpKaLZHH
jI4N9HckhYcb7tBDfno4oiaoDScsZy2TfZ8+fpzNnr2vb6iPKwmZyBUkc5dUEFeYEeWm8v6BOVO4
v9lwwiv8cL5RvfUq5YEkmcCFyC3mt19rTG8J703QolLKdSC8VgWYN3nrhIDnWan73g3zDleOiQNB
lysohv05CjLKNtlisOcKM8rWb8zizBSufFZQJWjrw4eVb664Q0tJvCjmyyYbAHaXZtW8uYULJs2E
XJZYXYwIOgKxygBCMK7NVBnm7uWNls4lE4Rnel/zi+WHbR22BcAdttexJtCYg/+34UxpKkZYPBA+
i85owXjtv+dHH3sGs4W2bM5ansIAynRDzOatAVxIjQH96TCGIcwyA1YIx69+RrG8LhgixgxXAx9A
Gvf5lNPCmtnVGuC1PoaRpQj70yr7pID1056Q37HqHjA1VbNDOn7QttBkRpFkbct94+ycw1Tz4xT4
7oENMwsYPKyFkKr4ptJ6bVnhJrNgICG7BcyuCaDaRfz3Ef+AUP+37Znn6qV2SH21vgDlS3eGiEcP
oPcAlwcgedqnvE0e5qxFkPhlJmPYToKdt9gXGGWQZefExFXYzxTg84rsBjYZnsZd5lHHG4Ps1WCx
p3SI41UW3tFPZxTyCzoLerqwexgKuAsdVqJSsYGK3B9DqzPNrvEGIcGP+ncu6svowovW5HuyoQZb
X6CLC/e9AaQgPhjgR8fPuWJuX2k17koBEMpk9TzVbZvrz3nKMfqW567797WWrAzL/icXJLWDqxFH
0hwqJuNeAK2qSfBE/O0BI5GovZtjI/vDukOCqyYMbsjnpAdvZ0XIvcpGCYcU7OX38/qqCfLon5OH
TY9V7CPEERDjSya0jFF503i/6KZvwolW+yx2Qx1dy6tTQsc0XvSwpWPOLOE6rG1292rFIRO4B0NS
RSd5uLXQQbYQxag1E6nkQwmsFLydqfNye54ltYGgdoaRMKm7ABnAr37n48AOMCHUaA3NyA70S4up
gyBFiUeZV10sEgJCHxGJk+sQKiL/7brHIRxdiCLzu31zbdPMlyOk0Ua3bYkjooLODDANXXs7mhjS
SE46YGn1v1S0+BisOcvS2aUh9J8w4/UrIfM+Wvo0EqAhX1cqSj3h1cAEzzVCnUZ5oRpZIpBDYXMm
2FHbWB9roLG0sF1ULMGRy8PInPHOzy7wX0M6C6822s3f/cPSzoA7F2oiMNZN46GkjkXoDvy1kysm
pCLCgtah1iquFhsD/JY/33WpD3RkTucqQBbUdQBiBxTXllbPYCuCljipKcEN44Pc1P4IoFsBUcls
cMJHTA5FzBMM8xmSF2XWQDplrS8Ce9L6+AyHGuhWc9Iie3TIvGS/Eg9W8uR0M1BOekSvgVkrMYGi
m+yTsqkgOBJ21rlRA9fWBSEg/ofIU1l7upWHKEpfet3TMgLAm+MpMX6X/9TnDZPvYF6eNOfoBI4/
0b95mc15UWE4/q9tp8wSOPBdGKZ+McCP3D2PsdueQWAXjlYP7OQQtuGac6slfIGObAhdxQVLjbho
nTBOWcK7jcVnwnEr/35el7EGnG8Mxy7CKBzhEOPyJkyqEK+Im4N6H8rAzZPAO9Ok8eTpDRPJzLJz
pHb7/6eyK+LUAxXAaLqXky8Yq7nlhMTHbxDWv058D2iM73+p/j7dbvVdH7XDSd89VhOdCnqegBkQ
RPH1lrnBgK9oVO14lS1Dq3cHtA0o0oxszxvEqZbxsPAvBcb9xwHQT2D0Qaj7L4Wc373Ut/Ple4jH
BT4REZi/fGxyT0E3mwvGt4SU2iheqQCxvK0aLdOcaP+DCsC7Wja/dmOPflV1mIMpxKGiKrrCuj8a
tIavF3y5h/tqsnShdtR0Nu4hLi9O5MzC8rRYciaOuwDZJWhcV/8D7/A4R8cDQavFgAkyK1zZAZRU
HQYpzgQ4hxY7kWk3RLK+zUbcGc5Feavf8098rudIFAKQC55XRoJQ4Si1BgpLtrGzkwaG6XwNzRCn
/PKplSXsnHNmjOAlVVDEgEXViH5B9QpmwH9wKc8XfvF/cNJk4AtNgpFsXiZsuYiUwhQCwBzhztjh
Ne622Nykl71ikP//tfEGqFnb8RLhSD1r2UkjAz700TEK5hrRyjenyYJhYXfCJt1uuKk8YzxN9oGB
/Ggo0xzhzsRXSMGq1X2hmUJxSJFgXpDo3xiPzJ+LQlftIkGAMtUW4TsN91oOaC0VjcT81tOgiXoi
6eG+W3nVxSlvy5vMoJidobheDNgZqIJTU8OhgJBqkqknPq2KxbMoWXdOkFLZr6W2W2LQ3spRI2Iy
3i/ObO63O3wKFoxRxEaTn3xtm0dhOWoQ7gW74N4yD7X6j46Tfh2rHqZDuCcQPs3rub8He0hcFtZU
8Ja7uCY6t4I0k1HNfSJUk15HQhJ69cme7wJ+Jba2YsilsjR0QfTR/iIYlCEYAdtOIXxTmnxUm4Od
2cfuPYTVC/58L/rGZxE3LSs5984HaQExhD4aF9thDuwynZ0wBAuQ1/3RT34KTvr6GCCAGeCIg6TC
0Bvhq2wrVjilGrSIzxW9/dhdIs+Ez1JGGRC1Cn66xO58k3D39biZuA4ycD3/ef26Sgx991MscVGa
TMuO/pM3R4Dd0OC7oZmKd96eheAN6vYHOIBqKf6J9wanVHSQuGMGE1X0HSAWJ8FRAj8tIGK5BqBa
9dLRM8cZ47TbGuyTbXfzFsj0zbREWux4ZfzaOb+ebRx+kKj4Gdyy01Vzw3GLBNRAvEVn/jE+UQJz
M/LbIYtwYxUNAzlazpUW+b4elE4UqtKmSAazeDsGrHGVzqQKZIzJkKm5jXJl/cZ2BpOtaygv6alE
HysQoy/rSCLgjHWgZzGrHzretjOYiDFyBw98rr31r8jjWtJ1ICiH9PBrz2cZGLA1zWMsZw6cf19d
umvWywUmfxC6PpTvWhgRunP2M76ZOfV2aiwpStd/wsfVP82TftXqn5k4VhrYG+y2KrRmPjxIB2od
5q+R7R12aJdzGkbWgVF3WQ/IqkX1vg25RoXNXJ58SUiv6wSpaEL0qQxjJktw6R9lelt8jFaxfUog
TooRz+CadrE4v5RYzoSm/hH9dH//dx3YcxBgTDMxzkoE0Uq7axkAtzdw04NKfIR2fjf8AM//RACg
pcXgUKRzCyvgFG9a5DdyLmNCdQLq4QYCDUturT/Qzgego+I56ZmdoZn2Y7PGNuxmHD3vMhaelhI0
15TwnyyMs9O6uvtE6zAgI1YPzBFMQkrT154y1ozJ6911blASCsFOwMHCZFQoBBQXhlf2osuWT/YE
0oVfHkcfckZW5dU1cu7/30wvtK1uO/C3Wg1CFCuxPJvqLpviUjhoIVUVExMdDndkFxG1gcl/BU7x
weJO5zzRA2xAz1TG2fAZ9tec7r9n7IZKAXnWcUnnvOdAwwCwuUsyy/h8pMLgsoWNTMGwjiB6LHff
eimbCTuwTOsbXumakF58gK8MU9+z92FwjSPbLZJ7Vx4s9aSne1+x4cLu+Ya09/UXXOStg2JQe4ZX
2BLhv26bIxTzneZEEjHaMXnxIYccq9SO9nbORX5jYfajjc//eo5jypT29Gdoju1XQP+vDDQirK+r
A79u8cy6S6vhw4V9HoWZntL2mwuaV5/zIOEzwFJ+3l6Stn/96dqZA5D5E2nv37roOsVU1l5HNV4p
p2xzQgrKZ3W3Rs7LssxKneic5QoN7w5ngiBqUfkTMg9lT6h8EGPh/yxkOKSF8+oqRthyWIHu9XGd
pk/g5EqIfMBlQuhy6rlc54WR2qdEc1UDs5qPOdz4j9vfyKdOq9nZJe89PSfxHxDabEBNKLLvEZ7s
j1dbyeiL2Kha8SMDuSrPQVfdYhqYlvI99aLiMq5w6nxFdrAVEgA1x1DM8WNuK+lxbhHmcDwKA9UY
BPf4gU6hoiePhEmosZ6BgxMLH7uFSAPHZJBZrxcpc6PwazbJJ+jh/+d10RwwqzHWRnh3IvUXhWuW
qD/2VMaWqk1UT6bVg6CTcR7mwbCNq+TNMU7fLc+JUois5EWPhbPi6XE19EAV3c5tCAfTNLmhHJBG
6WVl26bNggE6i5Hb7EK20GL0/hhWPrDTsS/Rkp+IxEHXTpE6FrJgarvajKi8flHx3GkU1GT30VK/
ZhsMdhOCtDAgDrqGBMDHgZSJ0kMyzgp8Eio8YjM4diY1Ljn8NkQ7hswu1xB41Igqgdtc44vkC/W2
XlkA9QfGP8fo5i72R4lMD0blWx3BztHPCKEh9cSAjS8JnymdCHIo7ojTa+RvumWNH7CVN7OAcBOD
ygBl7WpXLegfqwL1+VMHL9GeYrX5LuUg3csXYIJheB0Cg/Oyzy4CHFrNHR67DjaJF+jPwnJSorlm
KXgm7xIPFXV4AWoGEjyquORpXHdHJMmI4Ctj64yMa/RocBI02nwSYXdfXrC9g+wfDeXj4nWzDcUP
lboTgpn250Ih+t0cnUTFakq536CbVDHVz51nBOkKzXG70wGVpnkhiPPcOBLp+PwhXMOJkoaOFqQQ
FWbfwcQoA7FZEh0llwSWQX/1zSlGSo0Y9QvCuRmX0pc3mPbWFV1JT7iNCdPb46tXjTXDTsgMWcG+
+WFOoJb7uOiOj9PhfzBveCtwrBUXno8EigvxIMK8XzzaXHsoNfG4RKFL3sFbx0qW/DYAiDo3vtZk
PEETZX2JihEb9NzogjsuR19scvOY584ZVZD1jBgRmMVDS5Nx6H6Q8tU8hv/ECZL+uv+cnLt0Glnz
5RCodaKqbwnaD+YestypsP6f8/0SDF4SMoIbDhbVaalBbbmrYBC2YN1m8TTMIoM9LDJ9PzkRA4iH
nNOo8sC3+Habk0tPRMoMVc9FzGjR/AQD7bImmxHOHvyGEzoV6TMUd/0Ca2bb0W2vLUCIj375FMe9
KkbETxS757CkIJzzC5nxk8dbkLkB/awX0pNRFvTjL7aN9t/iiQuFskqzgXTc+Hn1uZMgRjjLUvLu
g1WFMC8Ac0u3XLRHsGbzQdtv9X0CUXGb0nv0N1DwCqTy89HfVg1ylNxwxduoLERcfJ9Ubz+1Ezoc
CtdwqQBqYIdQcvwTWF3aLYdON+ucFHvPheOzYm8FXuyKEs1S2RApSUsbhkyesgFocrG7qvF5kHO2
RSHmEbyUOCOp6mIfnaEstRSdQ9fs6wPE5T61yXkpxBkSRVpkFAxf08M8oWVP9dMvwDXahJNhRo6v
jvBjXFPnb8fYLBFG+2Y9Kof6vdQSZtiex2ls8bH3hdfBY+u8UYPBQCPZ3wUxxladER5SytjdLCsZ
e5z6bV0PWxMyTcnf9fjIA9FhHJ3bdFRdHSofOc15waAcXpuhyDQ3exPW/kH6k7wYiyaK7/2vYIK5
RUyyRypN2FLeS8NYvBfj6LCPbliNTeU/Z09uuV/NjewaoFb+/RvI0HGGl3IIcT3CMp7z/oNpwc9/
zuhot+/WU11RynsL8PfhdKciF4YUMdmgDscXFPiDkzKUV535pcA1HRJwSOnt6psVhuYd/uL1616h
7IgiRgYTbuTlIs/breeqWKzKOMLFjPenU9GNZ+gYdnShfBMbb7gMyGnHW3OQb1aY+nVTJfNWh7El
iRgRhZT+hRTxvjKy4YExMXHNmb+8NtM2QBolqrrWKc1INrj/zUsFiy4sHZocUyWFnoQDQf3370YD
NgmD1LmuJkBeQ41Ry1bhwK5gb+v/9x/YWsbs7/Fjfv75Rkwb+ytWQEVEdXXg/GLC8OiMdAqbfFJb
sXcS3Xc3BW1lu98JdUhy2Mwfy0+uOjAdJ8FXBr6ju+O6nIkd5a7qz1rxarAwCHdkCj6QayZ2CUyM
erkdiOYiuHXvetm2p01eG/xrg9xXPTk7/5hdZDRcnt2KKyKNrNKIc92qKSm14O+xGBbZsHiUG2W1
SNk04O9XssWFozB9RlEVbMPUtHo8Fs8SNKbWwHcuvShWiY4lRDOUg/J055awHG9VSvzzdGBeH5WT
FQr0kWo5C0LsqdAFlKyxEhgr8IZvHm6OPayhCnZY1BMgkUlGqoqbOBM2BBQtp4bEPbjCQTjoET9u
iehEHYD5pOv0nLRh8pI/qetVSGQ4i5UqDTUri5IDLsXyi1GMFlaf7BmbPYRy8apcgQi5DbniHXTd
YihIbjKOHY1FPE3JXq79OAOEO8jMOpG0cYF9LrbjCHCGqFhsKvffG6xzfeD31cx54bfVEjXl1Ov3
wYw2bB42UP5OtTcBgXkUlNELBOtnMwM9CnNQK7bUPAbj62VWjzuFQ40aPeIbCdGgGTScxBOvkQSh
EGj36oXGjZatah6rT5l06Q4xD2fLTA8CPNkxEWWIiRfKBuzaUBAAz0kx21TEbqXhryzAoJXC3tB3
96KAHxludV056CoL78f8a4ljb34Kh7lUfcQfESt9NG+xRoL+ndTd/Pb9aXd/sZduVFq5gd8mpiF2
ddMxgcZ58kyWLR+gdkrfXuhh8lCgS07JX5hoMi2Mz8aeTA7maj9JfDWppl52T2K+GEDVXME+F9kM
3MFow+TVLDhL6TbDtqbLzNDG3sTP2NJjNiq30GKlW0ak2Y1KC3SVpiHfRL7xflTFCoemSYaBAKME
Y1DkfGoGvMsbcCXX+8h2Qerf5WkajuRVJavrOG+ABIs6TdURlumAn1KmAzQvOuSfueavJd8SS6PV
Hto1b0Ra3oCjQNxeAPs61lN7R2plgtxfICXvvwLXcCQT/neF+KgiICdvNxg66XL1B5oHl+xmCbti
wmgwpH+qWB3aTMoxgBI9xf+GZEuHVKnIE4Pl9R13/iCeqiraoyCPEktTAHBGPDuHi/rN3SxOL76t
EqnVcl1f746KdGlSJZAm2U7pmhgarCVRKlyDP4CFtss7C2/zlzXyTuu8YJfmSggqr/PifaFPLgF7
h9gSaGyqlwqAMKQH7LZK/4h0vf2wrR+T8O6J6I2qEMiufRs+2wtw/zNSx3xsKTHpTYTiuDCNq3La
7MEQMB0Q3SmvzjVl7xXpHOrG4ikZtBdMbU2g6vNFwGofFofKVk/PV5w6BINtq5gL/RcG4CTaRN+U
XLBXZYq0yUya22M2g46EwNiYaoGV845vvPPpSPZL9FJh1srmIKT9vrO47ctqU4r0JCnB4vJbWb54
4x51ypUeLy2MF1NH8JRzD4xSuaX0ivLva1xa3VQXBzzKhaLUFkRyVP3Jtvu9JSNh/F9odFNo1ABb
y8HlNrB+xgI+svCAUIA47FIE7S+QlawEvYxOPkz7ZStFogD+wfjCIHbgMtRQaL3K/Y0YqwOwrSJf
0r+KWyZqBbJhN598v/E5C4pcVapYdzv1+MUMMr3A3/zYHm7nNJThSY7Jv0+tk4RA3l5ghLh/YXsL
ujXksOGMlT3y/ZV4yMuUSJoEqLIsrPNpRi7yrOxg1YSFs4x40yYpdv9Mriu6y8R4QutttKtiqKoX
EmlNeBn41zfg/oRznw9691tj5hVCotxydO9YmlvkSBAUJ70o2Y/LcEX5QFSYiLrdaZ3qLucHDpHT
nWMm9RonL4p8wSD1m9LTXHo2EITESH5OqCjOKdC1bxbndr0uHIfg8w/rHk/ZdH6Ph8shDfdoRMAn
Zyq9QXKLT4d+lyx729QUrJZeALFFiFpcK+Vr9NsVGiKvseRtXtlyaT4TszgLsBwGD7p2JGGPBqDK
VjcmWEF9oHjmjWY4Vn254QQp9t2+mhmqmjNf5v7A8G0S6BZ2YjbJDbZJ8TiM6PS0SRtlywwCVPIe
gQ7lKGby4e0595tksnVgTUGJjjgN/PmHt8dj4As4nzw7gZHpvyN1W+L96HYp2/80jXzZpk1xWnlS
jXbrwvRw+FpF4yBl4Npaht0h3jEsEoZJERz/TOIqp10FcWjRLiMuPQVKbM6P3WR4OMgonizDaked
l5jZA9sD6Vq+jVACE+Nukt1nBpmpylgsQqne6FFbafEC7rC2b9ZCkG2/uyBKCJeB3gO1eqwYKhro
L9s5GqkbUFc3U/hZ2XwlJ9SqqfvWSlLzFZNJI76cwwuqgwalfvFI0hPG9dB8iXaUm4ErZVC3jwXy
HfpWH8VtsoVFJMGO1HjEf94FfCkZeuYZ2w5iQBmjBkbOLvP3vjlhVn+pK30KD8dcnWacMBpoUohW
dxblMZV+fRdMMaMnMbnk9sel2dt3xyx5YQebsvmpzqJJDizUVzAOs+QZgoIERHO8oRN+dCeV9mCD
nepqDYDj/haI4M4kRUUvQlJPPZPy+MbCUkoOBEuGzmEPof94gjxW1UD9chbK84VnqtA8PZmhEc1u
rIAMzjiOHIDv9ElLHo/ycA4uEg+4rigUKSaPe50br8cKqdKMbwB0/GkeJAfgi+JawBOo1+ROpNHJ
4+1pTkjQvPfmivccc4tkAOUUYbXrW01nH+L/otKpyEhDzRchLvfPGZQwUX7GLbn1lSNCG/ehTEH9
kUsole0vXeyjgYdXv3D+7HhxOnHeeDfLAZ2md5XFQiewBGRzlNSJnyAfrz7crhuAAaSJEpVzkDVK
eybH9U5OgdWXAQ+nJDcGxnHma3aR7aLRubTPlHe8cBSF0kLQcTTRidsBeptLjLoa8T6lvBFFQ4p9
rlE4dvyKZ+o+mHJ9Etg47GUgdE6FBQU6DlU4lRyDp4hu5Au/znH3FoiP9ciQAPmCP/aOKxoJp9v1
pSG4QrZKaQiKGtp0PAbb0hiPZcfw2cPplIMVhcAUbQK3fQ7iME4buP4QoDt1ZP7Tr02oBxoj5OKs
rxHS434uTXZA3Gfj0hjl0dqY8Vff1pAJ7V8mxKuBpCb5cYNTGT669KVkOavGcI+q0BIKEHjJqAKP
gX1cEUgAZiztwiR5QQ6eu7CLWH2178NbUUi2IocVL/+6CO/7q3VztoY7Bxs0cETsJVNYTk/rsnUR
ErYBuUb3NsA4LAFzWPATVekv0uPRjvXCm1C1IHJZGxuQFj57VuYgyD9N/9BXp2M/LJAh41RelWIB
THjeInF3tx2rxiMbHx43ew60At3kPeZMBaoDgjpHmHPIZay8V5dY8o+5Y0rJV8aVBWuRYjZgHaBm
e1URq7S37aC1X6piB4AR/y5wP7iEfAd4WBw+dDc+pCKGknfNu0g/M2/lmHK8Shs6qsdH/qNzYct9
ebf8U4CI053dKW1DC6GfRXI8K9+StG07Q30QeBnsdcil2dBzlFvu6g/IBjn69ucS2MiAZ7bduKvx
l2KyzT6/rHbnOoot1oxjLvXuwZtn44ydTInO9QfrL8FC9rc/b1KJtuJXYzHOVH2VHO3VYorkdKNj
4Nlh6+AUZMEqpwADMRFnuYJjpYv+Nb1OgxPG+EcQs1aR2d850avMozsnvw4omsky0bm0wcnbkPmN
1IyR1GVfB8AXAsK195ncGkZF6/ROi3ZETh9w2WJncTF8kz1/6uO6hrjMgvJ2kx1FWCHlaXsJKWzK
x6UuoNp+yk9EXtwQyIKugshP1QkQElezWYZAw/hGgru/JZnhOsQf+4e+rYcy/qGsHX6wRRSq0uyY
q/le7pjgszYwAp38lWfHP7irAm5dXJPp8qJ+2vHWqPGDCRja010wbkBv34DsxG2NBZ26W8L1UcKK
ZtEt8FlYbhT8SxPO+kxugERc9MF1kDJk72X9y2L626dnBRs+tC/Ysby9vi2L4Q0xTtRMW+EnYKMd
P6JqPIaJreZFIctxGVZK32u1vVzaEwo0BQVNHyMm52G0j/FZFZBR+UFOBaMjB88LxOcyeBfcVBBp
Q2nUUnDVfEuuUdjVBKvwmSamK0Prqm+3vX+eWG3HaqxmNph14ojTAwEJj/gRzJEo7aseWZLJiZWz
jzb5sWlUoHyyxpu1SvE2YkwSqUDsWXYsxtavgIgLg+RHFeCo6ZZK2S0N3B30UegW+Oz8uJtWZill
httGVdcxbRfV5uBJMaD+xUr25oUoDFg68GloqiUjWkyx5z6k+f/Q5DVWF65cToREBZ0LbzWJgcuH
AQVsNE7SxgTVTgiuvA5t7j6CnUTq0bHFLVtrKSCBKfgdviYTpso+jp1Jq0nqp8+BGZCliNTeKSo0
pl0pWu8LhtTW7qSpUt4/4Wyq8QHKXT3ziowJOGRTyennzB3csAUzlryC5RLH+w6o1O0r1KVWOWOj
qpaxb9rXypJO6qShfAmGIkmddniQfKdod092YfbCr4T1kefCenHkUmi/tew5jznl3ZZU/rfD8gc6
OqHFy+9q7L19WV4OumfD3gHtLscTOuWA+qLghwlz0z82kC8IHxHPJ8VY7dnsqc0SlsuIMqlxf5Mv
RKoOVHR3iYZA0SEN2c2iMVQpWLd0tzFtd7KG11qtZOu2wUi5d2P0JU/MggorVmUmuAx5+eYO/J4E
xFIQc20ARZvXjcdeVd/pS1CJn64j/Zb81PPzcMkPDwoFkOk609YnqTN+Sdl5hAwRChn9evwCDcws
HsNX28bMaXCoZzLL2PFlii8CGZiDg9JP+natQ/PyBWjVmtycPiYSSce7mxf7r3XgQvmr1/Ev4KnL
pt55rWLlTiuc0GLtfguOvTCgKMzra3an36IEY6b5kWVfM8bi+X+Ty2qyVBWSFhxgZoCw8nw9E/H5
JlwxkRNg6x0HqJXzu9BF4qIljj7FRurgcQebST6YNZ3rbMGcuARsYN7EHeZZhFyJvCwVaEjLIAWT
Q6MEMqVD0Jo5bLiwouNY1ABQGN4MF9STgNUdyDTM3UHeuD01l330d7hltfyszy5u0ShqfypDKe8/
/5AoePbrzSAA9A3w3OH5FIsV9ucYR3P/soF2zJZ8udRPvwvP3BBikodP0fdiT/R+fSYjvmPjwLmf
+B3dXruMzvh/KINTF9bkljI7h4RgaeZ9MzfQFI1uXYAtdDkoB8E8fNVagv6CRPwAiBblC9ij83XQ
bwgH+yuRKpAyV9T779MA8xZ1gFC+ABwzxiq4KNH3Q8vU6p/50QxZafH0r/J1vd9PxMjdkUhT/ZVc
tBVe/9zBrVuksWY9ubyZb5IvMOs1Ao8vLTPr/FlRkjXVmrpIaATp7BONCTZgSp3AjXONAB5Ya1UY
2rq6QJioTQUFFhEXB8aT9jUjDmHNeiOuRT71pGnrMpSmm5XLD0RfVl+J8zMY8xkfKXQa91emSb0I
rxVpwXq3DFW3uJmskiB9AoaFKJh07jPQOlqEmxSYWGuc6yUd1kC8KfPjePo+LKdE8QnHZ4KlK2pA
K/xqWs2zfegU+LxoJMwdjSmhn1HZLdkLlChSGSFdjC9x0tbvqwvrUHEsiDyrFMiSrNGqdflEnEe2
t4O6w7sHf6gIqfVPqZwsEo1zSYIjPXoWb+Q95YEvoYqXHSFpf9ZSlVeGRtEE9+BWwNueZ0tewldT
Goh+avQOWtQCaX3DHl0hhRyJ3lnBrTRPIXuLxTvWyvxQPElyBiBM4Fo0b4UY34tzFzMB+4u8MdSR
pUYj/fYwWv0GUhZx58FyVzI3P0zciGsgArH4M67l499fdSh6KB6DqGrX12b7/OKjlIhwYqCuQla9
fNGDp5DveOH8H94Gx49J0u5suSJfiAOxj2aC6M1HuPh0WVAywpcJqfBsH326rwfZv0eK/ZNTuHVv
KC9+l4rVL7QXrdkw1GHT3xGOFKsSN9vvI+bgMg7DNNcuCsFe1+00rb7FL0RhUO2TJcvmhip+VtR0
qapZrmXbD4oABV59lV/LD+1VNixcpoHpW/7Ql/DiqXBaJkGPl5IHmJQ/9dcCMJ4v9DeiyB5QPG6D
xTXemtl3XfXgfZCbkOxzK4LDYYdLpPyG5yw7JnvcOCtQirprnm8jHGhSWKzuxPbO96nauEYRZs/R
GmwYCDYbfYQ6mgQ2qm2o6rlfoXach+uYYTK1okcypd2b57baB8J9qEJ8elo3g26kDbksG+BbjSPk
umjvDPyk04UZm3Z3ShVVk5Rwc59gdBwIOtkK/PAgN1ykNvI27BFIwJ0F4+wEc3gbVmhuMb7D+42Z
Ok8WHNQKNpC0rfuDwfBMk0bA1cT0WT1pvzzgUKu9bh7mtyckOBpEVkcgsATlfJUvwWA+k1HoteJT
bHyTT4wb0e2M645PqEEXWlEUDue57lc4GdD4FanOrg3jeXBjcFc+K2Ge8ogHQGyzTTXb2NeS+3uA
RtNpOOYSXqfDBaRCSy7gQ0Kej0Efx+mnpEZJn73N5FawOw3rGOn01REmsztDY91vftn61rU4jDPx
CsAlQuEQJkgKsTLff7TrttQPHYpv1Eu+SssL9XI8GgvqusBIX44iCP5xSGKfQ5SZIPNbX2rcQLv4
dQZnYZcSVvKEzEr2f8+ye2dCLTjI9NKQO5T7tDcLxGTDWZjgskNM/LRSAU9l/KRWih8VaZkPynNy
Y99dHS/dDy1PJ/JmvvLxW4i/3Wb2SiLb0HPvKNsTx1hCatBXxtSF7FPiO4xNGvm6D5jwauzIb4SX
ig3CkuWYi6f+P3IeowAnIxWT3RYmHr8Gf1UdSaw7gk0XiSQ7RWcDyULqMhVPbiH6WRmkzKlB6mxU
jJczwdnN2IcJDmN+V4naKcAUDvNoe202TDN0gIksyXmiEcKAJYSDtwKO89ALxLxBHMRabrqzYy5E
62Xz5qQbrWjN8jx8HjzqmdZIIL5y/AS1JXrq6gD+8ftxJ7jpHnnfEhjA0OE4DHcW94i8psurGmM8
r7N7TlqnhIhkgMc42/EB/e9B0f6M6LAxpoiiCfvsjUGjPxWieaWl8Gd0UFun1guNxt9lf5Gp/6Vx
lMgYTzSBhBkrL2Q9XM6CZrC+v4ji46oJs/MCysKQkFDDEZdTlt7wxq6EcM7d+uXUqDxaI78Bn4fw
Vr9uJKGvymZjXgnaZJSw2sb+5d6wTudeArTKnF43f0Ibw+jkQ7MYfZpwp3dIu/KcsDUb0++uY+2U
Hu6UvwnYSaWoB9nb1Vz5zEfKO02W3K/GNWFTajsZj5TrXHgv4T1FO7g6jmkdeAp8kkoSXveOIm6P
11iXHYjOIcH3kUyUvh/1zpHdrjpvDssGVIsUnNh5zJoDzoMXx6MtFLCEaSsqghMP1VjvWx8WVTgy
VDhTRhTw5wxl3OPSPcMw1H0CG5uZpwEt2WA1WNsmUArCbTF5IKuPpPCa1xqsF6bbJSPie/+UmgRp
7FKYBzEl/YRwDjAq9c0u4/5lBHGa5cOfZ0vkKX9No2J3RggLlpyPZVNivhF41T+21r3Px97E6TVv
7XUdPLD4UdEh+kbXeJ9qqOTRXRyMJ8+eqzqtY/BXr+Ial2osQR2bE7VlG7b+rN4PKbho5uzFXU/G
Yp9Mj21uyemNIN+V4wDbkVL4bSEPLVh86zdTRByUpjzxFwf4m0HrEInSjk45mFV2NKv+CiHv60Nn
WAJPulAilKWpxgUFAkG+kSZ9MPskr2S+etkIlktzytVGfne3gzYMgGXdwBcVpCBvrET7luxNspXV
J8b70SFacs/TBrGs4GP2KegmbglAv/yERkkJQvuVJqvggwonodhZpWheAIWqGquDQwgO6kbalw3q
/sbveNG6iqnkLwZHzUKdjWtZvb5sxjZbffJA99xUhpGfj1M804PHFBH/7ESQdhr3qYHHaAIyOlri
YSJM8md/qYz++3NHjVJlOnSBq2d2CW92MVg1Yi/+0qKtIhYn2bT09af2F2qIIhgO8RSHpKVtkM66
t0+m3ycq0slXVvL3G+AbvqCY+iabOjemydjiWqpwfpULkwDt4LefwyZXYTmM+nXcwDIJR9AR4PIV
xZZDcT/WvLCi6o0LhPIFEkVFzbP8KHgOR8ojysSHIb19lyWs2qcY00j1bO4B69GYKsBSKrBYh3gj
UNTMmxN5E+OHi0hanldEEdGMfwv+DmrbvPKsLT/Ae1Pb11jZV8pjDEfDMTR4wbpK/t2fsKceimq8
hQk18nl5bhof29LR5PVrvOxztzIHgqXG2DI8z3nA/LVHmDXthRPuL7z9OdVbbixJWb8fodXbQxTR
VVVt5lG5ckRPUIuKqYXntD3HDwTYStiqCKduwheAanwLf5EmjYdsA/cCXQVuwRq65Tkh75zYT/pt
qeFWzwdDPmEXmzl2KQa9rVx9NHH0RD4CqP4f5wmdFX9mr9LQbCHIth10MxGOEftz1j7Pmiqv5f8G
bRZeGeAxZUOTHfxbxyN1rm+2fgaz3c/AzpjtYJWx3bSu9WZ/4haY0ViT/u/EF1/15EBxA+U1qz4N
ClX6zhwny3GGo4jm30JtTy45OG2gd+uS8OE1xLTMZWJOJwasxr+J9DMqyUKEewOTwVbA2wHNkqKX
mh6ULT+mQ+ep42lFSlK/i/QKyw9+1BfneKPAGXNKBJgtldaqvqfEki64GELt/lGDkAHlQuxLywGG
7mm7cQpvHqplYkJ6cuxrV2RKxXiC8fBm7U1bqsvg7Z6Ot/SNcdy0z1DRYs7UWxPglzkciPmLyall
fIQRgJaUn81ytK8T6Z4sOs5cWzP3Sb5rsGZT5GIJpvg5KFaGv7l/DLV5c4ZIOsl2OhD+pWmkskOQ
+6T6qxQTI3T7uaZGHFplp+w6sJVwMn8kwkLuBXG3LEbucN0wiKTprWbzqVYwAt9cvpK7vlqF4QOw
dPc9ED23wy5IRYCLnT3h96o266xdrPcm0l0MJF8pQGnii3lxiG6kBJzBoxTrTtYvvEGlKlNm9QJQ
3W67S61Gu+SM9NZJ13npZ5D/TkzDld2lfKCFsoK7jP/gF/vRj2rnX7Br8M3+gNKEKOtMVJqLqHYE
+lVHuCiaY7/em2Y2V7VkEIf670yRRUBFG/DDVfvPnEInkOWEfVSGPqI+eO21ZhMsIU2Inr0y0+p5
qz0knA6jhrGnH3hNV3zUo1QRCAXxG3QSlNoyAbIazwBAJXgmhvJ0lPEpDKls7lhTVXOKUFaHWFki
dmeAXsRl4nV5QDutcg9EU8GzgjcCAH7BWDVUxD8jkgcWuDGyaSnX6k7KYkh3gIpC/hrnY86Ty5Nz
GvRQhUGf65nJT0Inywgq75FuoeoqNv9JgOyKVD4y7gmzysw6qaTvKa/+OtJgT9zfgAhJ6cItYxV0
ErVyEjPYtDgfLYyjps1aGHgx/yQwHh89UUEeFEM5zPNVvXxZo4gakXeYJmj4jm5+XPJYGMn+j+eB
q8tyZMMxg+rsXBmnFHxlHsHmGccB+nxlgTTCPF0OwaYds1nYSm/ELjwNUZSA/yZQyVYjzwMSsHvc
TZyDPTRngGBaHELApkdZtlrQCAp2CfWc3gJnFsQOt1whYQtH4k0iNt/7QP+oxLQlQ2t1HXfbMYkF
Ia8W1Pz/lOhNZCsa8uOI9EtCQB2Mc6cPd4GbceQj7VaE3cEL53SKMT1Bdz32yfcBJDsPk4m39whI
1SPbGn1jkuUCuTo8DjzToOS7ZYn1nzpgN5Cbze5TlqEYsObP0YCM+F0pI7qQkj/ToyMDVPwNfXsF
z8BzpgSxrB1swAhu6IZpThbcAAM2hapuzMzArArQMs7qd6VmoXs3WrjEE1uUAUPkV1OWUSugtY45
yVFys2MhadMnhtejKaDl04bUuKwR9Q+Ys+hgdLZoOllAklo0LS50iDaBkEhriOOP0li4AHATY+KU
eaLIpgXWgAXN2FGkd5bKYTwAmgxhbngOt2GN8pLwjeNbL29bj7f8cWdQvMTVu8NpEWxqZmfR9YeH
53X6P1IDvZzAorSQMDp2QxOhMNWFSqGKfZlyCdoxQf1IsBQ7VDZhUnQHIZJr1C+ta+n+N9eCcsUI
0HT/CbPP38KlgnYRGdWIsEmKFSJnx21WuoWuH7jj4UJ7BZQNsCJgj8opDD+F4vt43e6BuP5DxtlR
0D+slItqcuOKKoVrf/in5b3qsHommYGAfsSL6c+Wu85BBQkC9lHbCTrn4ws/+CDGapOiBByR+JEd
eWJ8nzaAkdo5CzelQE2WZy4zvLr507btX8E1XetVOVcxCbjv/LMdltazFM+qucaq92q2MczJMIXQ
P7FAa21lAC7HufYvcaxxLjQkASgl+0br3jY2t4U5oqtwviPtZGD6Qk6WHTdUi8BsMZiXUfgB7/e+
I0Zl2dIZSwsFoh95TI+umAPMwJuWbhgnlTWo+0QJE9LRP3iBoJj7Ef/3HjGINQRwVIn7DYVKpB6u
W35yhB5Qr59zYZhzRyZS/lk6EKWVInhLo3F5FY1vkJ9MAu5kv71gbAsA3I7e+qeV+x0rxwxdCjLj
1pK2jPhzmfV0rSJ48ADjAO/kPGO0vo3Qkn9WaxS8zutmUv1Oc2Uubyu+L0KcRUM0jvqtR+1YC44W
PZF7M0eq+b5kjBNN+ZqUbYMd1g1qpgbm2fG2YXK+AVtNKkwjM9RByBU4O9C76NgaQnXlk2HaInyq
KCNYLW9wDM90V5WLCGXn2i2r4c8FEACy+ALbPf0et7IYScbzRAiJGbr7ofsngJSRdBTzHRQiqUJt
sdhgtcalQ8ceKbcHlhebPWInG6RsB2J8qkKx7lnypTBN/0wui9FnoQm3fSN/zjbSWmo3kt0Wi1FH
7vXSbgwpIxQKXFYZyA6uZkyllk0wmeAvOJHWVkjF3DNpVc1briaXhIPOFJFT7Z4XwRjgHSQY2ujf
EJSpLr68Pfgmcc6KWtgzb37rUPw7/tUU4K9/Y3Gm/GauM1Jyqp77eZnqsahD4DsJxRffuPzmc24v
kqrgXvYhuOTS3/5hrO+YQC9+046d9219BPxR10j3suaT3OEhrp5A4CAEmkIQOGlCAo8nL/zIyzsK
VPdFS7PNqMQbE4nIdAoo/C4KKHRkobnBIYreCfmJUXUxeIq8MwtrWO2UDqXf0hEVHuFvp2b4gfsa
o0K0IlUWOKe0suFgJvKponR/+YC71kPqVjiOaTCBzx0XLl9t2DNRhuQgVLNYuQWEumHj2n11Sot9
RG3YV5CSmAHGwm9hYc4YLNMmTre9Kdnlgh3y1aUb5GlGE9resG/PhhO2H09+Mebvfs8uevRpLRxq
xg9ah5+z72vxoMD8thbuwn17yrTgAEhvZeeVSObWCGoRtS2f6HZdfzNZMOz/mXw4WzYNl2kuNbdA
rB6XLfgxuLwv9OzcOqBAWr2Uh+M3j5UzUM8ToMng5RGQR5DLc4jpAqKbddN3DNKoB++u7zd/ONra
K9J2o3NlPgaBY/VVh3VA0oieyGFrrPlh3JJWlL9cb6qgYysnml12g7aXg9f5bVftiVKBd7FXJLyc
lRJ9f47uUxXzzHRg+ypb58rtT3q5gYcAkLVzCjJ1DzHKvcytWybI1eSmTza7t/nZQA4lcNZRmpVb
Bvrj6tGm4dxl62sjxwLgSjSK0Zlt9l5kxyrVydralGePTcs06QVpl/MnbsQ3B7dQj8I1S3ibxhFF
rexNqpIa/CrCLyXME9ungDjWVU3vE21s6Po2Wi5wVaaTMJGwatl+4FSrxae+IeSpcMOnI2Nt63ys
LEIyoVCo8kZPzTAZN4KIZdQvBliqc5YtjMbeaxnRAtiQg3KPCZqZhmdd2qPGLB67IMkSWFEFfxK6
u1Z60CGmsjnlZlLkWvktJaGDheY+9Wvs/0linPYseW1MzDaf/TqTReq7Vi995nKHrExgpzMyfiKZ
YB5apMnRUgGrjpg7ABeJENx0s/y5nJbN7lhNsVd5lWEpDtUlpyohaTgPcRhwYw9oNfmcAR/89kA4
JCTjernO7wu+buwboVWl3XYcRU2fE6+77um1JLdCnKMOKts4OusM40BAa4fD6hIMK1FGvPxLa6eo
IbxKFAn6Fek23dDajRdbLzDVBYzHwgeYP7QT3D4VsGWGpEjPPctN5xyfZ37aCPPtKW4hZTG8k4NM
U00JC0rlBDG5l7bfTG+teknuTit18qBG21oWdfr0lsryP3hHss2YZDL6A6Igv2fd6llbGbcdSByQ
D6RF1R8KWf/BZhSjGl5Qxnh4RCuQMTin4IGsoGeO9/ZOmPvFY08QDOupvOlwfQPqegeUO98d2Kje
6u3nH04yRP543/sUbaZquAuJnX7QeTmII4yELbScuePAzgr/iqbCwdizU+fCf2zc9Pep1+W7ziYf
bWCrEIu4wov0k8r+sq9kriHepplvKakGjXyChJn6DAAr5RUUljBODPvr4RmtGuQUYgsBeymAR3yj
aOYUsRoNlhVBSpSdywcx9NSX5gGFbs6U2xI87V6jMqNKzb7nCLpmMO+ye4dd18FDnccBF3L9G3B7
c7NAUhrOS1mQ+CCI6fuvCX0Zrv3lqmdNqXEXqyeB3m9yzTfd1m1zggmqFSobTAx2ZQ4ccpb/KvGD
gbuKGZAtii9pQ7GL3iMuvVRmtTfgYGCpHR2DzVJpXiHZNS3lTxzg9UZNKYWCeyg2FnhekQb8LyoD
65+plcQfJKDl2X9jRyVHOb888YKUv6Lg49clQUeXRy5jdhM8edvLZdFElk76cr0euZkR4QDf6yuG
EIcL+WgPD4EEyVArhpXY94mjNe7RQNXpbWfm/dKuxVJkqDFOB8CfuVRZ9KMibpz5I3dr+aY4EYai
B4z1JdXs2QdoIY7Pwf10muhVfgeoURVL4iMfTOPVb/slkxzgcdAEAEzwpvITS5u5FVIq5QtwS/Jy
h/zvH8vcm6NFUwVBKvsG2sYHXqnytWvc2bfJ6mvs8wCOPJyd2xCXrMmRhWtiIqPAb4Xuxio+4nKy
8OHoOK5Vky2e6kaeMHcdOqarRFcw83fFW0SJNab0U/WnUnHslWIcR7KH/HNptzsRlad5pOspssk2
7q1bqwTr54Yd+genbT7HBoNhAmvC52K5jBRb5F4oCAYOMhIu7czpxFL4oCuzBZDtXSxs1DceR4DQ
0rh3HxkfLzklXiqLcfNlMKBLWGvBtrXT1PMK6FUueiiL2JyDr30m2nlVCcUuTQ5v3NE4RaBbL3o4
AxDSO7TOXerNhETMzd6n0sM5QHGY9liTUic6aE8h1JjyeET+OUyG75Dlz/31B2l7VbBdIkcMejmO
TnujuuaYsE8rEjQCvtccMUbZF3hTTJlFKOpK+0LJi298EYDLHsXpJmwWmfEZWLWtHlz37fUylVut
jdxiO+1HZVQmyZfNcFroU5XKMS2tvxIoMVLPnMomcluwWTA41lp+ocLjVq+6XtyvnLM84iUlCf0l
5RIP7ps4/jCag6AEqGwZeTRDafzxQpwM1pXYONKQVppKqJy+b+tXq+cBw311lFSsS1BH3KpjCWo3
vAWM+AqslIo25nGLhRU6mi2+fik/hs0Vr+9zyDK2lRrzqm4W1bnfaQmfaZ6HU08CSj+cvFSTSakm
oA/025N5/L+8DkPOzYtj1YpNTZwDAEij9hf9R0dKGhlhBCo2CHn7S210HFxLD4vKVTN7VHSAvqYT
ljy8db8W7aBdM+8WibWDq8FbHB3cn5xGgNbhsKJNeVbIvkF8tqCnXGFSPCA1M9W3q5zsRQ5i3bEq
KDpcphoND0UWwUKY8iGveZ0/4EzDaYdM5s7fMRi2GkPkgT/1fyQwK7GH+9/q2DIB1SNLSrf8jTg5
IQEHb3IIKz9JjjZsFidmWO91TChgPGKNdJ4+i2NVbHWFU9ViRzyj9cgDwP+VIiXeCUxYEBY3m6sv
oUQbIRCXHmzauF4GqZoUr5qqv2YXS71znbsCaRId+d3djcNW5/gpkmn9oIbS3xWIJC+avQ123N66
F5AzBLoH3hfsrCu6eXjyOdplmx4gMczOLUQbvfNPH+DUB9jq6lmu0ttgOOgdH4qyZlscworkCyoZ
WZP412RwNzelV+evbn/n9Tfylz4gFUwSEAgETHPBc5iOPYl9PkaMQuBcxmq+gnebXelXIMs43eqp
QgWfQp95TsMebtgfDSnro3Zo3wCQFajvHoxi2cyEMVuX2cxdsXGQ7JZOqsuhFadn+vsv45Cfe223
UB4PIDZkj2gurpURZrk3RocZCKXf/P44A8oEAfYik90IcMc7Ugp6mTBBEqW2WFI64I54i08i3YBY
UG5Z5FLCrlVg5r1SsE7a07GUl9DN+mVpw+PPZFvz71VaVdbWgtBLETMzR3N6pbsWzAL3Kjx8u9Ad
jS3jl9DXIMIWf+DOOzEnrJ1KfWz8iuYenkq6+gJSoQ876zf8FiZ6wyQRwIa+hGlKSuufJBZBISmg
pzN1RduP6q9524qa/g1NxFfugGlLmmWb0JvBR8yIGImL550zWnSUhQTGcPwrur5euXTdJGXBR7Xz
a346WQFuhHSkXcUXGUhL5LuqPIfAGcDQcYZw42iq7mwfZpy36cvyAMwheXqT4vicg91RIkey0jVn
QAcjeVPzR6+G99J6eoa9SwDGZfLc5VXCWFczTDvmqTk6BNBBkr7/UH/Xq2VDiegKCnB2syGnPiNJ
weyceFxzBeDr3ryHj96zH1wgaPHUTOxittn3Cex8UQ5VLZW8FQhEPhHH3k8y+DsGcs0cgvo2DpCS
9SkVeKMGYpuzSR5CKwh/y2XtDEhVxxiUKriDXIZWbJnksjzhIDL5FPAacchRZEgQzWE0rljrrEAZ
f+qgtxWdHREAMF1RVgxRQCSZxQw3zc461hn/dWt65L6UhknJU10rK4FCPNXl6dPejDve82O6Wvgz
nGh4horQbMLWifnBDDc4ZSEVsbwgu7fQFiYE0FDRKS2bO5B1vRme7Kyqk07Lzx18TnlEE0xuZEQx
s39WtFXM35BW+Pfi3wtjYbtjTapx02E2W2DkQT6eRE0FvrcceyJT8eVhisLuMB1jXnt+LEWKpWLy
6WOUU/m5THZtXkt32+ZQ2EliesxaVWhiA7KNzxKrnm4KpC0hGsEVhoRB8BF7Dbw4YBQHAncBV8ME
Wy/fYvNBxDgYqHVxstEFXBPNtn4fCb5kkXIqeqJ6F1q/7ZkkZ1v9zMNDWJ7yNpHKDERKgIGucggR
e27Aw4Y2fzgdvjc5SlGRLJAQG9+pzifrhuRjBmQ4Pu/eVcu7IezCvMlqtcDsNM5Te4+K5QXmiSEV
RlGU9N+cK6nFy7i2E9gEVB1+4Rjn5iKDx7vOSY+WRIYUiSKSp7LWWCgP7P6CB0oFeJ89CHQMzDN6
lhhyAJ78sQ4LDVFVFGGRUasmno+icw5pn8lx8/BENJFwdK2EDr+qOcKl0zSuhbuOSTOaOf3EJ+6o
9DivHFj1UCvEFuATz3QRCn6P3UrcH+h9AbEaBi8lEdgnKXvb6ZHj8Wb3sQGEQg75bW/xZKg6xRqN
W2mgCco5xuWTbP9xpLamnlpDVBF8e3yjrX61nyJr+eA5fnCQwzgMa8OGzGud9LM/BIPL+81CIgqk
wOHuoMD7zsVgFEFXmHZb9UX2OqDW1a0F+L0zJaWd2nq42H2KNaibhe7v5tkMsGA+HYQ6HbxG7b9p
l8uYvQzQNW5ItrgNyaObLtRLretKAJz2IscbxHxkfNXMb2xNeJoC3IOevg8ijMBrySujWhgYWWYr
keMe3p97FfJo5kO3m814eec5o2hlMc7n363U+pnZ8t41mMnFRDfs1M/GZrK2crSgXaUngp2WEAA6
BTMDbLNezIDEZfRvbDJO1sRnUTyOThI3ns9fD3NHBL6oCfGS8wb5+dZY13qlxpVs1LQDs40TM4qs
gT5DIqEdzKUVwGAhRrpu1iaLbWVJVs+n2L/LwZcDYVbyFXcmqmxIXsxYuRKc6NhPNlDRNUUOhBzj
BBk+yUqYdQya04xXP2h7cPdP4t7C1c/FimsJ6cUU36XV6E/OiVcFMtClLp5KTW6dYl0kxTY8sPm1
qmw82VQllD2kytAHaOdZYOZS5S8LL/dOb0LsmWo2jWRucyqNdQAx6Sae9MC42g/3sx6LiF409C3g
PYWL6t7DtAlpv3gzVlxIQT2/Ul+jjHB+00EcWOt31z+X8/w3E7uaK0EIUp/uJ4txn+rn4trHTo2v
2sqiHlARapJt9LTCDL/UE7Ul9B3h6cK7y1xWcC5Pmxy1O4tBgmlmElguqgCOlxAGeIR6TDg2/krL
/hwGerBC52MkvUM5SP2diFl+lN5j6xPmVLCuw4dqDi6tLW+IWPs1XfNjKW4u/Kc5o5PjZ59FLNvR
keLT3oy3jsJtMc9oXe/dR5Bg/vu5Uepr65vPa3+BiOmQfgRKTjs7m3xwTG5kmj8Qy36X52rYz2Vu
LG8L9Jegt3HWXM7UWZuH0Za1nPiTLb8Ty05RnP9HSbFeknQVP6RDK5cMPGBRxdq4UJt6xD14uoLP
ePbusZJpzCMCf+tWKpa/91Aju7WrUU2Mmf6XXgSw59ZfuaFS21x1ibfeRYvRv7obvuXfHMwB+uSJ
Wb4WAdwJy8D0fdKg+CjdG1Lus+Kit4B1hDCeMo8yGiAOL0Mduolfq7yycZlic8QT4smB/nUI0KaM
ifgBKaCTBsKmX28HL1umoC1fAiHRpXiaVwThkq2RTLCXIxpbqXJyTw+lnW5z24/QZwS7yj7X8y9W
Sgy7Nqv43PRcCUyCCWJFd8CSTnkCxtLPQK+JnEh0QT+Wp2RKgNaK5qhNnH5gqNJzV6WHK3rhQHa2
Z6I544SuxbprTzNmdrD4PBAdy2e2FEPfZ/dKqVhJTili2JrZhfCHKQ3wiw4bbfAQwEY4oIbB9HPb
hTMn/fpzgkXTIYJeyLIT59El8lge6Ps8M58MlFgbe59TEEtPd1xm68LMyePk5ZZsxj22Oa5IO/CI
/MDKwUZYxjq7YFmCLyU38JVdgiY6qbh8q87LCLPp3ndvIt7S9fpzz5NsPNn5toZwLWyqF91p6Zq9
sQJu8HqAo4PGTnj6Ek9A+Smj3Xw9RDUFWGPAP5ZhJoN5YmOwzwPMW8ktsvy5Apl011hrXffK1c5Q
lQnXHWzfHfVE5rOksaGzp5JuYIS6P57IG8AKlxTnIX+7/pTrFeni10/ZksJ+Co/QyRfL6RIKMQ+j
y2eu0u7RaVhkchvYZ9TfO2HbGMQKzMjKtZqur6COKmja0wLpVlp3Fu+xKn24SDshtlEFDeSqKJwC
tO+ykrEsNcCNbUYYv50HMmgf3ASEMH9HGQOBZquLOHEROQjRdNYdAfGKSG5ItWdlA3TAkwPlVTUz
XGiISwHhMkHNKARqDJPA4lEf7nI568jGpxKKMON/1TqegrZH782LfVr7KpQW9hOwNKwu0iCZD8eZ
G5Zj9U2yhe9tS1rjcshNqfOOdHEmPY4D+DxYL0Ir1fYzsq8C0jgK2VryrxKZKmFnajw6+crh5S/S
Vm6YIDYYNhs7836kFSLUVF2FBKQdAE52AwKhxYTkyi048CfwogSUbQ0uJyQVfNJVeIBk8NdHgZsW
cHDpJKX3HaMubeHivkO6jG9lQIsPhe4uemNNAyuuCIy82zx/zjb7jHsK9l3gzNKeRb3X/pWmXjsO
2uKhg/Otz63Q0pBfNZcnBXRedDczg0WYCCUzjd+c1uGvHdOKtLgPfU5za/DpY2pmkllopnE6od/D
zJuAurm2GSvX/E9yESAwPFOeF/y3A9UI/Hz4hqodIaINeyyKEQoPSKC+eHertaA+VKAl1C5foWqQ
UPg9Gta9nVdpFmM5pnlc3eY/C8rw7KilKFlkHKlVav8JoM5RmqL0jbWiJwy2og2zmKTGiB4EzS1O
s8eJwsEXMmOskSRUksqi1fniduiqBcSw/OSDncXeT0fqqpMqQIGDnjteeTeOgtIYkWg0VGUuK2b1
PW3eu/VkBbKa8pbUEPmjaaWlUwexND81KHSEKypW+qil4+Tm1IAk8olg6l/mcumkASJ7KjdTTc2x
Iy3P0FsFkH2XKtx+UAdGrmj404COkrvjmDwZ0jKF7QzVGKhZfszkpnAkaAYILTRpeIRokIbYB1B5
ChA0F8NNf7cU/RcWZbzZeUr8KNy4fuTkBUGWNJkwjqWZZGmFUSUoHFzMZSii3TEQM9XbiyrqnKWi
ai7myfmta2YOperUrXudXjL5l3bovuJz3ucHLDNQuQzbP2nsPmEcxyonEhv+Ju8Gnl590hyMdywX
98V+GqRy2j9W4dDmfq01HqOr0OlgEx5nLOTzBmbJstl9bJADx6Ox/+b7RKHyJ0BXelgDn2MSaauR
kTLCX77JC77dEA5guAb3pC/h873B5S/NvxuzGuErFxqOxsAShcQR75OBsUSzJxK1gpQahkxzbXmh
01PjwqTAWPD7960/2NQs316j+pC8dOpRGeOyyGDQn7i2SqbyLVHYMkqrMa1/jZSmUk6daltpCgNE
L2GAK/zaPxWugSLIWJPgMLcsF1aqgYK7ExE0Gvm3uqfMMSqUS3cH2cs9K+FXiLY5ZG+WOH7DpshA
o4V3JZllrm9JHHe/ZCUA6A454rmXklyPN/orq33szXYbuKBDxe2lpXI8emJYyvWcBepcCjaY/3xo
NqxprqcrdaO3Gh9j65P5LBRYVH88kKxnf6rtwJN+ROjaeZa+hRHeZWb2RbyltYYviMu3Uf220F/y
4vOBgrOixlO4Wq9V4X0y7zCUeosSrvGsKKQALzSI3ptrV6rR00hwmMVtEkwRW6Xu4+v4z3F21Tfq
k3LJh5AQo2nWvIQKa7EGi90MLS8nVptczPd2pXdzhtt6D2bwvXIcPQNAPxkgrZUiG5KT/2CsXQbD
LJbvr9zooB/1sdQPhQXEwQaaDofkNB75iJYe7Mj9+f9C+ZnlT4msR1KJe7xw0wBnWcfnfTpfGKNO
BeWkNFd19rJvbNaLN7yJTjJWBiZpO27U5ESKJL6/YAvte0B+G64AoI3yMses0B64VKaxxhyRN/1g
ANNGqyHfoVhYGeBLuI0aYotn7+3nwSthPubZRXCBHiXASMzz1P3D5GiiS0EarZUXCSCMsLc/Wh83
X1O+HqHrbqDKpB0df1z920RAyEhYsWDufEKmsgBH6RvbBjjR7uj95NPm4weeh9mQjfRSz/lvWyQ4
dmy94ALBpKxM8QLIurdgstBr9wXOdq/NSx6PHiJ6FbURNXhcR4BoJJjYJqjQ3KiTt9QljsXK8wGS
QEDA5BwzFFkY5dJiCnqjV6egognrjqrmj2b43BBwG6XVcSXPhw8SiodnsavsLQmcxruxUcKKiSf+
yHJBbS4hCU84mj9MZvJghii7xt6wzJAhR2fVqYrL4Mx7F4mwTUl2qi/dgw5DtqFbqgg9lWv/M9ym
mUoyITFBqorBqWFBIlMOI3yMoeg2u5D6KparT7GNQZ1TVav5dLuUQDR6sytD4NVh3H2gFYdFOFc+
hIvLUnZyzWi/BruHMfw3q6EuSLa/ZnsA/vTKv2JWI2N2TUmS0af8OKHcmr1mXPLJvEeaTB3o6Qbd
l11LzTlek14cCkfbvpS4NthhsRbToiwZ7ADZ+uOmA4eqOHV2PcKjhSdK8WJbXALSYrkK3ST0VXri
fiwgH5nlQumbEgxdZCwx76ZXS7d03+QntSxajEhYt1s2EwQoLkv40/DtFb0pwbW7dJgq0pZBQ2hA
mMqOfWUDMa+W3+3JUdgwpEu/P1RErH2cHymeU2jhI3bYkq/17kE5TsiB0Irc6m+w6MYIxo+85NPV
vggbXilLCOijXAT0JD7jNsrULxCQFDOMBpH4oVPE+Nx8+eOwVmwclNizpszytDNmqoMSeK8zKmLy
JfEgtGL8zKEEKgh/nA2ZgnhaYYDDlBDaGf5NSeRTz9PTrioMrN2llpNkW5vz3ljZ3+SMQd2Zx9u+
HDh7FD3MwTshPmTpiH6MCXkM4X0dXErW02WNTPCBibR9c0VmpI9K74LN9o1KPENJv7tDWCnBZGzw
FBHzjrjcYMItwLt1FcchVjRCIGvDJWNaDmZN0f8sbP90x80QHybB8omWxM7pyYoA7HoUm5lSvmxw
Bp9JYPCz0SNJ+CQUb84nv3h+VxIMsSZocSBb15jdTS1CTYZYC2B0r3XSxTij+kWLRf6X12zlOIod
CMpKHvMZwS/juoCM18kGuKKeL/aanwamDjetx3rKn9KwM+bsOp/6x5QHxr5vmgu1iuXkw4uJNvLy
Aynqade5Hze/byd3EIw8DHrVNx3IzNq56s+ngWUIt1z2AWTSRoP6LQ6+El/f3xRZbXJzZ+ZMnHte
f0tGWjuiJkIwOuaaV6lvxPhEweXknYvtq6VR3RJhviSrPnFOV9cZUYOqk2vPonT1b4hWBoY4vTaD
IYefq9yZiKmsqHmTNxU3gvh7eiplIhA1om2FG1k6q00t2qgNoK7vixalHydPE3Nh8MiP3CWClCQy
NHhc5jIddCYfIEcAHrkNxUdrfjgXQXKTXOifzlI94AljO8zTCoEHfBTCa4J1Qn9mEuB5Ym8NDLjP
24XVyZjO42F+UGz6kHyO+nYHpDqUORpmm+nRiEYWtAV50yAcm2d+ytiKDY+rxXXHSHI0e+UnySIh
HgyoW81IyWDr+F3Ug0u7x93jYvBhTmxHQmMuIfNcTBrEIP4EDrXKAm5xYqSUWxFdPuteKwyGRmah
rf4JBmI9uVSIh56ZBORYB6sWKpxplMh1uSD10L0GJXQbVu9WgCh++HZ/+ve/XeAWFpiEcPyKyJ7f
WUuQ8udbLr+nBQS6BGkGenKNWjQSIgKMEtXKZYGzDnOfCGAfRpUHxHZYdDrQnnxDrkNJZHuUcGiX
hJJ+/oOnDWB0RB9pc+zScheNfqB7E8BJcNCJh6A9j0i/YZdUYAk//VW0OG+WrWLYCoeWqF81hAMO
iBCptQl850zqjgTxAVWlO3RwSdiiHoa5XE7pu1for3ibYfJLYn1MEpL38SwwAjHwsK9tZ8+4Q5OE
RPNvkhci34/hGQ7fBPxXiGEdEn4XGWIjprLoXmBPrH0TYPrzMtAM/HDXfKg51+IsnfNYU2JAvNM8
9boMMNP/p6/mdpbNlcL7rh6br/8LvHJC6w4UrT7e9H5jUYJ10JcU/EWcVpTIFX/ZkwKHELtTkzV0
Mp8G5MTHTS+DHEtGJttiY9ELdl6O952zlGLzs9Edv/+atB/0wEKl1oKQhZc0Cf1paAvUKE0l0ts2
UCRsieduIo6RcZr486D6HikBu3E4SvkJEYY0qxP6HXKOAS4x4B95qCMvYhTUIiUF26F6e8sB3p+m
ZZe4jGzsMFZUUBe5V8bgTu0DwIH7ERCjbGPEt5y2dqgcA7MOZQb/KjwCBqs2EpL7czBWflT3+YKx
zMC+1Kwc5aGEw38wPxHiWZ3C1M1N59cYv8y5TftDbH2BIN3baDDXUc6wzhCTkukVZZqw9ez7wQ9p
Cn43kZ4iolm9ygwiA/rfEZHyZ+2lglr2q3vb46cPro8+jBRBh9tJ6hM8fSusypHNxVf6dHytEDLc
s8IgvPDhLmdgbU5uyI9IetEMUcTQXO1+fZz9XnOcKgFcQiU/ILaxkksa6a4MZEdRCPwULSq58hJu
nFuvt1j8zOcKjCZYZC4chsJ607AwE43Uvt/72HFx6smOOm9faN7vl1WiBmUk9ZwigfFn8MeWwHA1
SSc4sjNQOKBxJfYWIQlalLFsfwMnkFnQjrBjJxCDz6POAKJRk4pvwgsnPgScJ0iEXAp+b77NVf/7
+4LtpN0izCLUSC25g3FT/TtWJRXkzzJBxw5F72dJJCBcgXlFgXaqgXtRQKXoFZdMNX/zxEzxeQaH
MW0ZKlh3JUBZcOA+hzV5OKPP5yvKpFoURT4F2LL4L+SGDMLq144z+SQ47sLtRdWCi7N8npXzO4dD
VC7SERwi2Wzn3JwRU7zjlqB7/QXaKtVTUlAlkdzqbiuscSJLHzjag+fsfblFTVq8UHi+fcj8lHpB
1qzCrVuchDyYmP6IQeoF43CwMM5EzBqa5pMxxHsFl4AzztoIY7LczbLWYZSS3XxpAOQhciAWxqei
p26JlWzJvpl2CocDNum44dhj7po+46yaUrAvkokByDB8EidU+uzbOJbyem2JGsTdH31pI1EYbiJU
hA9OXenakr0XV1rKQsPP2uWn4DXFfweIiWnz1OHcrbt9r1z6HmYe+Vux54zti7qoFC4uS6NXMmeN
0F9mct9g07PmnXlEpAKLQpo3+3YLDygd+FnRwfRnNqaSQQO36uQmZ4ABMpcHMuV1bd6/9RaONd80
jr8XK9QM0pH0C19Mig854xGIsY+5ad1iIW8f0QI4e8RqSO4s2md2BycmHP0eLB3PtJHk0klLgk86
kDPyKg0vNgh9GeUb0+LokQMlBHitAtXOAy/XidUPIcVBIZkd62oyvuRIdLg60AZNMb2n2BxNMmtr
U/+ymTv6vKwkzANr7we4EcM1tSajL1iFk/p7Apa2jh2UxuAVD2Fc6EmavvqEw06D2VhhAhTsE2SS
qyy9mKzn4HWBi68GzWnkGaqNpISyBEBv3ZaejCnWSyaorqsTm+Pqk5ZUTU4S7hYprW/ciPjCxtJ/
oyvDE1YGQyRWBFZd5kzy/wBcpgkb+4YGvZqS8Fentp2QX40uoS6WYeBDlKAwNm6qUlA4vTnFtRYT
Z19e+HPrVJ/ZaR+bvEoMnmgS0/3lEMn1W4IhkJy7Bbc5cEw8peHlLTHwxfb6lQTexKyz7j35kM9C
aJjepuGQXGAPg2mLi0IR9yp6/NkDbnpsRXZiX/lptKSlU4m6opWxbU5Z1CjenmUrwgF+HsBcB9jI
KoSwX43hj9wKPY5A1ObGRFzpYG2TEKUWi6Y4c350Fdbsuew1mvZdwyo941FMSyeYP1rczvWdK26G
eRFpwlXXwSZhLqWrayHYNNtMzU0AeLKIdRALWBau3NBV6XLJQjLYwDBPW+nBdSvtSLQSe/XIpuwQ
7PaYl0ABhmuFFlJY+G4iZsVu07n57uBOzgmL9CASd+n4968+g48OxMovgTjOLMWTetin2m1NwZ9u
9WW+rFqW3ec2G8ExWozz0R/zH27J4BNzdNmttUFFaV/LwfUfe4fnCubVLxPoPFOr/vhjFvnrB0jM
sBCIWUp4zojHK0IZqP4DK/scGn9Msac/KvEvQwmcIqQs7tpN4IRKasrT/i5MxnxiLDsdw+R9U103
rkMJc04f6cR+RM4/mcl8ZrjWoI0CRX+M2WbijuoJMd673hUMhf7SN33HeiRrpLxo+4rr6VIRdGl3
fdD0NgXaxMK2qQGZA03i18BeUf5DQ8PwA8lZ26AS6x2U++2roraDmbCdQbOXt1r8wk+E7nadsac+
uN53w8mjphl8EiivOylGXzcqTBnyeUZQc84egGyWtaQnhUGIZCyel1btLp0Sq3dSJOr6UmUDtU8e
QZjSQ0uslTL/3z/sO6vePCM/X+PJLx19i2/AwioLBxKHhWgBP989q0SuqBxgvavnxwMVg866C8Gq
Qk/ti08sT4pF/9gMaWd4bTAhH2WSs7zm5vMyJR9grjp8zmGb7QAr2rRE4VBirBxv8PMD3jQ39beU
DM2yA3PPKPn86NgwDct/0vfpR6mJE9De5vr1O52WSmYg77JKdW6nG0juDLlS/6LHpNuhTFmvLTfe
yT0nGPwQGb45Yq5McP3cNbNwZmTVfjU10FORtwXiD7SNmqOT88QO5aM1M0aroZyGTlZ9NSwGDdll
yI4rmbueRXucLmpowNmaMWlYLPaGjMLIboXSi/bRwbMAL+L3FXFBCwmRnGj7fpaFurUJ5rGzsNHk
li+mRmF4IBIpBEKD/tyc7HbuLSpDcEP1gyAD/fW9ZgDTOQWeWNd+wtFKpWlw1ElTB7pujDnj5Sc3
olypyQAazZsGCPragoetYifLuc1fyJFY6caSWZHP1piTbhAumf7gAn9uOxdtt59aQ67k8Dzp3qhI
bL3SdiiqGjwkhAoIz7IpKT9PNXwXulE/06Q1JFUc3XhYiiavRWo+AugUtKd3Yph5i3GcE42STFE6
ik7ekiPXDMfyzbC2TO3Ofbg+00av1JfPYsk69xRV3kttnczZDZK1bfgDcsTG6RcLexMOYXsIowvB
FzP8ZByDPjn+hTRZQ9Q8Pln3Gin0o+5NZ5mJenDQieuc+IUWDCNqJtlOb+P76aLfxOXUfu/oDzl4
lpq43+oEqOWTFRzfZO0Jq3rISC7Py3gpU+iMLHoSyj7/YR6nE80vI+jq/XK/PBk1KlMwNtoqmUwG
vunSlAy2/ciffoqADC04Iecq0xFs6WcGY4S2/4mGz/SZ5QwVVDOBRnxqMPmJjHUG0ejr9DINXNes
0WwszRJX7CC526v7QlWhkPOvBALADC4Plm+Mj6kjCM3S9oujSsmYfkG3avLY+HeCPTDIMD+KIjO5
NasO4KLQMVoScHhOyM+b9r55izm/oWFH1ykrNQSnHBZCsA4hMycfb5XPaxxdYbE1Z509Pn1HbXog
C/pbQgU0HNOGFB0GarVsv6qspimwc0EAX/+NcxIE5CRrmeMGW3x0/obaryT4HPfUCo4yT/ytdIzL
lGUUe3Zb3Dttp/8DC8eLUu9l6Xo28vcEMPZ4b/54I7rUWrvmH2q9GJefeaAHJ5wvfwwbvwCXTwf7
6anyPQLHGC1fhFQWAsvihA4YkqXrPHPL8QmkPD7FclukMeyH47942iDRvehLrDlFjc60i+ymb79Z
uDy6QDIxlxKsAmuzVfSImwnIqYpYQCbTe8PYZ0FrOu2zXN/tcVxXyPYzFiwJtuJsCpkvju0uyOpJ
dN++B2S3Yx8oWbFO33zhODVkBQQfaBDnpQrphqNVkhFggL0imFxQV8boXI4dr2bEHmgJDoj28zL7
/7VQlpg8xHSI8s/g6jCKuuo8plIAh2krKWV2lyjZDcTgR4dgcuuzTHlXYgl0P2Dka4y4Y6cJA2y0
ALz3imev1sl584YG2AnxxP0oLZ3cQRi5HDG8hGc26PH+t71rvUARumyK5GcF7SV6inNEV80YOAbN
6xKwN2iV3h8um2Yoe5/FJYmDHY84Fu35bdSJrXMdfZD8cgzVXTLFcuZk+0Ellmo+I4/rjql3PKnQ
qeZ2OF2Z8jlNPiz0X5ud5mY1lpmc9EAKZpL517gJK4wlJVuwqffo/Uis4mzkhbUgOHdi8Ohb+DOe
YEaoV6ObgZR1Jb7TaLlpf8FrzJX+/PXov5hSG4G9kF8fsLegQ7Cl6VsFKnY01i+cIpJl4vDtBdF1
/qQCkKwkVSvpsWZ2FfLkRKdHzRg/Lnbwew357dQRowK9ARxPVvZL7b6F6XMFZuxNcOJneOXk7wLn
ARrrNSQihdmVC+xJpvlYYmVpSbo0st/4QXQEbE4rPD5VrVln/gONrtETHw2d9nmbdZqcJAO8zoDx
aT9Y60zz+R8FIiR9/8T/q5dTtUI0m1IWAaoHTRzB6KqZd8fO21hM9/6kpuGc8MFg6qS+i/aHJCFc
l9gHtnFa/J9v0dCUbGFS8fuOIuLQjZRWj8nE4txyMQ0aCSV+6I/jgKctjEs3OgBVdB7N2KXNYvrB
5mtsI037LKVjoJEJk+0I5HKvavOTKjTiYkl4OP/cUPdgq7i/Cmj8W0lzEm105v25tY2jDXQ1xTYz
jkTjhPSyCdhfIVXsedCf1NeLzt9YIA2IDix2bJZCFTIpAy3rUZsoIvod7GCjOvd4f/2ZENYiA04E
cN8lq+/HtHIVzHRMbLzc7QxvCpetB1l9V0TdIKCKvnrhZcsVombESZsN59O0MbynDRuRNWhae1co
caWaEPwLyn+joocEw5zAXIDq5fAHxnKdDFwUrN0FJadzYIEnT9yISAGQs0ddjfBFDmFK9k+TLTce
pQNvyuuqQm4bXRUlKMgcJnQjvmRbwqZEtaVHjfJGf0S9SuSHJCQzHyW85WfW1vFdAj+8Rs1BSh5s
DGsrIzc6gFu5xJJ8q0MeZDVUKaNUAaVKRsmvDjQFDoQ3xExE+OUSXHXeEspgONmBd1sTsz36dV1r
0/7WslC7PfXL3ojU+akq2u/tB6/mDz0sUwb4ofOzm5933FMUV6Emb/A1lMQhthZsAbnZanNM3vDb
GqzQf+GeD1TKa9Fk6fKmObwGw4mob0BcitKdyYP+bgjmEjDfDSVZP4v2qQDl+hdZDgqSOuBbqrYD
+8KdnC9FmVa58/fsdHRt5XEbESCkWKDs++hrPBsuSpMWgUMsjQKG+4ovsFLXPLf36TpCIZJXFesV
KVTMpcBaPdAUW+F/Oe4dstymifbm9aZ2rUJxXqa6AaJYTJgJzlhKtwl8qU1zK6z+GVuqgHp/kGUa
bzIW5niJWQUiLdqflCZw4PdPR3pUB4EOfG04P6nW7LjCImkHeAz20JKYcjY67zHtaHmd/7A83EnN
qlmgj1zPDvbzu2oO6djHGPdn8C/NWY2d0LqaTBIcDKdQRpe7JG0yVfSDM0wbITJ0tNRAkaWdXAXG
ffqqAKhI0qyngaBQSOZZgkO8cM7I3yxArAx7Bq6tjry94L98ZaQWb1eBnv/Jp263qRYPE3QmNinO
fAJIU131/Xh+gLskti7RfuJ6xwSt/86P5QQ9g620usCzn6rICnkRJFwJQlKAOjiowGXkCRpMac8s
TqWYJShLCLxv8uh0s5loqPxZnOf4lPw7sfPmoEpfqRcrATcgR5ti6cHeGkUfs0sn3fCajXiofKUC
nDwa7k1mgiv2Nq00nEzUAOeEmdoWLeQcBbsNMWz50wVEydHlxpG7KeLR6JQ5e4qKpnjHRnblEeCi
oDIPKqoU7jZGTWoIIMCss/iTnGPUKc25e7fKruHYX0ndsCKbOzBz34r2Nf6UR7Rgdap5JljzOCCa
BVA6QGLv12o9jCVAQjI71/ZniEK3n3wLvXWG5hCA+ZlHaV0TFK7N0qTXu76BWbOrbLFrS1L7ig87
PVXpGeM3s0F2nORXd0sZ9a1kXYlIW/tIwCDoGZl9E6naBQhkJ8xwN62NU8C3iOx5NDp7w6dLbsQ3
vAvV+3AZN5xZb5urAu6i/KBV0w+zfju8ZVSR/cYV8GAmHEUgbWPHwR2eFAerOgPNoVhJZZeqUexM
f3+p+M0xtPUq8PViYnVN+IQXAvjhB1TMXKjgs1MDmxYeYdXaIzxqz95b43F7oKEZ0Ocs9of3qBrg
qutIse0/kFyBOpcA1kabjIDz16OlF8xDdXKN9YJgwHlmR8Xk1kcjSJf5+2yE+qS0NNpSYpr3yFJa
+yQijqE/8P2MASREEVClkPd1Q4brPpsEjNMBuIedFK7+JhwJ/2XicpVHXeouiunyF9em2u5cepXD
X0frSQKwsu2TaMibz42QBvGmWtrGjXYhemdpRfiEu7jkHYM7mP+BJrjQdBCDu61E/GYEaPv50qXi
no6Vh57zTRafDZiNLvlaFtJTBkmX1ZnWgEDxKqwuCIR3JJFA7fO+hwekBMSWemUYHp+oZvQJ3li5
4KBqSRgpLZ90k+AN3h4ci3+ENsGoxG94CBze1pRGj06KnOfdhHNeb77AE4i4MLptlt1xeSSZhR5h
Qw/ND9NkRIOUTWbuYKl9to9FJnhihmluZP0YsKkRzzmrJamPz9OxuJyNTUmeI+tZ7AcWpB5MQqLV
QFcGxOXw67UCe9hdE6mLMhxVdtbdEPDSTYu6XX07OLVWjxv6c6vCWz3ci+ImwBEobfx/qoWI5LbI
GmNu6Y9rLqraljULJIB7rJQQ5fDYrzx6MUfleRvH/7O4JVjTyiROcdMCpwssk2SoiZtLkarxF+ML
z+orPbZpHIRTpkDW8sQiVRbURh6I9qkczWz+llQuRBuA3wFiD2g3VxgIqPDpPBDA06aNNVk9MzyV
G6XVbw+0ePG3z+1ZLcCwiWhWjF94uS1VpkPpKVjgvXN8IoqMXqzIhEWaW4s7lOYQ1cBrRX9bxlNj
WjgvyWmggpUo1hHzrrfzE9TPp/23MqeXt+IRJTr/YnvAgm+jU2lZn0gJpu56KILqUs/xxZSdH3Wv
CaGVXSouy4cCRC8xOhKS3fYMBeOAPQxMPorHZBN7CxNIQ6sy9+x6YPnIc3w/+oLTbN2RIluPUtwA
UQHzwlJTskXF0rl19vwMEnXTCL4yjAg9QE/3p19Q8SzHYRprMQv65j3eXd9f0+TnaQJSkmODzyOB
OR+enfpMK7//5CzTp683CfLTufEDzm1nKtca+pAJIdRnWdjE80x5sPo3GD/525SQ89BU573uY2m3
mLF6EJBJSlrN4ILIsZBp/oJ9cvjvpyo8D872LCKW5EjLDOpFYeycYQAifYw/trdOUJn6sT/nXzkz
tKzXoBgCza0Ptyliqzix33lEWjik5HZzCuRWvtgHkrCm/PA7FFnZzurW+dKiUXRoawurZjYd3JTs
exmWofc6CDZY7chYwha2aIwFT5Th/TEbMee8vCPnZrDM0C2dn5/60z0w216dNZvWQoPHc5f60PLu
VACJFhYXIzsCRen2KJrwFqSU+VCe3X6+UjRXDznegVxwa2tKeRTKJ8GiOQqtZLP2p8KmkGA3Oz0Z
4XB3RD32Gf2K8FLoiQCPnARd+z1zEoSbruJN7VB5WEC8SRWtdPEY7Y6CvlHNRmSqr86YkHVoNuQQ
PtQYnNtLHeMbTOIk5aghWdWBxW7o0r0SVlsivGEUPx7yWdbampwLGqUNQg9uiYrHXCb7+Ix9EZWL
jrEZSdqOnJ/Z7E2UpNhg8Xzajc4s0YPt0dmX7jFAuMf7lpVIOoB9x3NN1Y/1e9jddF2AFYMCcJ/j
2GKf3gYOt0A0U+KiZKuNiFPKE8TgmOiSqB4GRQyq7KX8Ep5kN0aeuPa6qGaAgnW10UX3W3nytX+7
MxnzJrt4Ew6q+aik0QZGh/8X84XX3PuBy1SRPsdIWMxElVNeYsKhV5A0hti3FMM8pUS34lq/3tVH
zT8vdwXYbot7e5r67xQFlf2FbnNVtzGQqlP+9Y6lqB0/0C/k6GPgpk4eIvhPzkCGkpvGEFGrAaHx
Ld7uoxn58y7hPQOdaXWC/Wfc4IzzT6pG9EE0FpXuSpIkQ+Hqc05xUPstarOV1OAhpcrDRlEuONXK
khrHL2xDOtv0PkmGRf090Hyf+0aUJSR9LSSU02lTCCoqnGzqm7NH2izUjarmUQ3v61RvFnEnlk+S
I40LaBTtYrsHuagYF9N6p3ILNJ/j5kOm1bT9HWD8V7PHwJpJOapjwiB9Miyo3Sk/QmCwCIJ6dBvV
F+j/N9XhuFnkd5bdB+w1LAsXTtvaVixrIjfSgtlr3pL9BAxT6bBYbYiBYZ5hy3iHoBcSUYtLq1j1
KkzLjwqNMMTN0giou80+BM9MKoEp2aDH1iiFl5+qhxhkXvtL+nq8dbQBfe8fCs/tsq+AIiw3cDMm
YBp6IZ5u80H8oS7EwC9imcEsAO8o/dhGh7C1iL+Q3HEHIkAD4UcHGHzx+Z+Xg/FWRs3VKUGNvQM1
lCZJCVlKk1D6/6D4hgvbIIAfEcVQAwYQ5jkAxb1n866vW7mzUtYk+71C+z277in9VSnv31HzkONi
VlIeYJ4dbD8givxWWh/5qjZfRl4ZkEIAM31Naicm3lspD4AuxZ3LfSOo7jDcsEYBglR5Q4YnxZ8L
Kr0FxOafrjDgdmvWTZnmk2Jd1Vk8hLvzvyYkuKTGP5oei9umGLlqDYbfXSmAgyYwZP5UMcJJpDG0
+QwF7wWAig3hrZbejoc1XaAZ4VYA8xmdumMYis85lSdt2NN929512JE8X3d2ZczmRn5pA+9LGeVW
uDQ/Ua3coTfsvixqOpqsJ7etAQAjVovvXM3/n7e2xIeinpAq+G9BySqfL24kaiFqeWsBaiSiJ+s5
Zt8k/lGweeu37LpSA+NR8rAEXw7l6EfBfwgLHki6nPUsCM8hKw4/FNMu9zvrcHoRj67lmwCr4ulY
slR42NaPZBCQfnAQvNkdd7hI2zDLCZDkG+CYpT4yDTm4pq+pVtvzIHEdbymYd5zLUcQkq8arjau+
/bsmIrHvLkmB5ptg8hzfRJn5E5mB7re8O3XYVkEUaC1vOWmMp/Kt5+63qX6MtJrDiGcyWdSU9Z1B
/bN+iNe7xWgXvebUDOkw15EvGXxPycZif2SvOTPeNJPjKG+1lNBnwCRyAMlCjS0zMNIk/1SbNBkq
/8GfBftBxje7dcjjaDX5Kf0rSpkv9wbe0PybYYt+B3yiN73/cg9eAWTl/vAfGtjQ0inhhO+JNB+F
TMW0VvMrgJk4mTLBOI/R0R/L2FGrTAqOos2L40oWF6oNeLd+DnFdTIx29SszlVp9hK6NY/0CNW1+
i/0B567UM2y+60xmZ1T4pgVtfBZWmk/zRyjn8oKSmgVaLevDf6B+FqBVjQujLop2+Bg0SGskobkB
WVt66yK8nK/qdt3vUc/LRPAGex4rjjIFQiQiBHmOofTP7xR4AvDM3MyLUXw+3GBGVhnLgrciBHxS
y5y3ONSITmOW1E6CLOHtc0V2MospeJ6sT+FqvTRdgxAtzP7CTkSi4IBZM02BZ3k5WPtZq1IjE+2Z
afdTu2NgIda1VTV4PXZ4RK5QCq0b2IbsFrtrfm3PQdsfvYJNaAhytU5s2PWqzQShbPxJcVFxRJzJ
Ljnu4NrJr7FQ9TslE76v9Lrf/oZiHwJTI6pj0ozvOw5Z3L8yOI/dP8FzqkHzN8+ErUwcQ+9iXFYv
0ILf66YftMmkWhky4+wSu89BoMaZJykhyVh9uju2hvgX75/wIffhViiYFpkiieJ+O1LyN4wpbe5P
KJzzi2jFQhqXF1Hb2kPmPqXtJR3fRCe6rPMEIVnydmyK9rCh8J3XmckWncX+JXGCRgq3wMf+M0AP
LdD2j4tHdJqAOWLDbLtFLfkW8Uxc5KNXm4JqRQEuaMXiycTPCOWYPkwhqGXauOceq8lNQgFg39o1
JdLp7x5nzJFw9a5coI2wlZj8P4A/tjbFxUaqkALTL/JwNY23l9eo7HR32vA19eKHlqWLAhzaLJLz
3szyJTS5XawTVuKcoRMVcFaRuJ+jETSx43f39/Upzp+kalvtzid6bblprCAVPE5b6k/E6s5Qtnbu
6QzvqfRP9EgqPoGLLzP5iQAW5Bw00DFJEegwoskZfls2kAffz0DKnH4yIV/PL0fJ4D60uA0FYEFK
/Y+GvANklWs8dRsRQOpJAvA+gHEkteKy42YWqozQEhAtVmgCbuRkzBRaHF2O+KKNURDQQ44nDOR+
ZkxDOCQHX6ZVs7dQLk8uQ/8BXzK17HuqPkmrgfzvvMdskK2EaJoLSmKfllVg3tDl40dYudD9/j61
RGOdEwa5kYDYRp9A1PihWvzQY/+KSTwodm23IITwrk6V9rIIZ5DdaEWsZFY5NwlsIeu+DqPzpd1j
Qr4n2Yas8ZPDqpcx3BuVCgnGmpbe4a3EYeGgScFQScu1nHvj3o5fWFKIk/KmmA1/tZnZjn7uMSna
tGrsJfYDTWjkWJuqRtM6Wy/iByyGBtJYc+2Vg371mkfRP8FSlXTMeWxOxeOY3ANme6lZH6sP4B9h
PoyJFK5T71YA4SrMZRL+HByZ1FqrngnAe7TQKisRZ1+Zinz1WP2PI8uUVnClB+D5CgJ9Bn5qMYfN
ATG+z5N2/504xolVlwS0yj3j6s3j+kYssv2BOz8lbvymXoi8K0B8RlraJeM8lLLlnUnNZ/8tJsPS
5VrrRAOEYgbqnPpK5rwVQoNYoJvTKF9okYwr7wPtsZvqIGxfJA0f1bWN+sVSpwUzgMsweM4bkcrn
uVibh9WUXpSsjpHagZWF0Iyoi87WYa0xOULSmRCE7fJssVDpcfMTOXV4fPbBrC2kHkWF45UyKJ4c
ebrpmmhC+rkFzV+SYsTqXfdgawrxJzAk+XI9JAuwJVd2LED/WuXGTRdcuw84N612vSbf6efMDqf+
fsbwJE/deb8N8p/hd7IR1PWTI57ALkktCVhGmzj5xF0K5NUFVXRt4OXxLhYmxVYfddPX5U9N4ZKt
8nElKH32FDKLvOxTim6RxHlUXMsQ4e7l2fBy0A4sDXngvaYD/+qGxZi2+Qe77tz440++go+3hvYt
b4U2HDJfjxsfNOk5u2iN1t10RJdixzSCQxP/RffdUyBkmGzuvzws4Yvme2rx9gboIQtxWGK7z4zX
jnZuah8jAYFaxab2ENGGq7FzP4cC8p8GJHSwLyoYAy4E1eNMwoWQd3YPZ8KddIth5BS84LxKoA4f
bxx+3ruvLUzfJrc8VBeAHD3l1jaKjFLCwuyZvFib2dE6TCx9MxC/H9sCOuRaWhVx8z4wgSxKPMkI
IlwuIDOO7HMOST6GlTLul/cSJG/k7rprOCr0hhiRnuIJ0UdtSYIb6c9ZBtDuTRBg8yHMxbSrF+fe
ImEunVy2qZ+NE8s1dUO8hyZlBW6k1Ape7gzZHaKRbXe1NzIFXzZXC908lW9li+8Q0+Y0vzP1w2CN
LzM3v/PtnKVhddO7iYnFi+SoExAi92by/wCEO8MQeIN1s5EpgNdh4ZjPRgroOrBNRsP954DIl8Mf
LBJz8SQG7uxclQDhskZ3jjsjFbPS13mmJNfQQEX6SYzLM8xCtOI6l1ElAMqriNeTjOg1hNcRqDyC
hn+umYwtmGv9wZ6oGrt3UpGExBxbamtKlmlPv5WKsn6S0JqjoQFjLZT4W1D1H4PLpNsAU89G4IIt
TMDxkAlPBzct18NynIqwtJAo6DkRmwEBp9F9atyN1Q8YRpuvHYolyRsz0zfIaEAhu9Iw6T81zHAa
ir8DvRKyw+XD/aFPXNxKLml72jVT8ZTrBv+oCqERPIykoYWf74ZP3GtvQKV8ppvnUQP0InDHi5d5
UYAGfK12bCSACbR/wZEgNPP5IXNoylojXk0kQEjnkRIQTeZXoZmZjbQxD3hwiqMISMICni4iF3to
9SoDncXVgKLKybz/HmXiC2xxuGFaXHT3IbidmBy3c02NtH/OU82k2Sebhv6iYs+V9x641kqt8NJ/
Zja5CrAxzb5fEVCyTAG2lyfebZsSB4IYP6+NwG5R45kUiJR9c5VmNHNXXxGllxVE09YJFsmWDEei
k7aTOCKz1hEkJDlQobSFQKD+ouM4Fp6ooaG+Y3/NnTOGy4NyoWZct+DROSpSRzCxiQjypAvvXYGZ
+XkX3/YkJYJc5a0oLlpDwJ1lUIRhMFTv8pP0yHt+FVEocIxcp8qBBinJm16V9lktwZer1n1gaeVB
HNg+zKQUGUpzxXy5gMzPSdzSBXQ9pwTGPvrZxtv1BkGpoOt2xNvcjW4ZtivOnyQGEddaOmomYuH8
eyR9HE9iZ8ia0ii1I2ybepGunUOyJn8gRBg4ivtf/aLPT9UUGaGuxC6YXB8idmpZQES4ClGB+Czu
VSqrTckaUoFhzakYOd4+awH+rihEaoB74hRn1KusIXUySgNneLZfXUPCTnJOYDC7TBSGMchJ2EjR
sWt/9iT/D0jI7dEvKhT/uLCQrGKByghUhnDlrhL8Zal562X2klkO+MLl8sxkRvjm8OfERFqioPpK
c2IeFSAJqLan6+3Z++bGp2OWOEziImJnKUc4U0z7WuEbJScFNnf1SUmaCM7iNntHVVsMiUr62Uto
BDgRYBmTQxj5AQHdq8/up8BexEJ6uTu5umPh/p91Xx7BdrdKjnYIrAgQ5WEqkCa1L/V0vmNDGIk7
qmcx3b99cBjUWPI2gsR/jhVyN6wbk7qIhKbZMo7A8dzL20wUc97ao/yrz8AIfUb8k9j8s/nxTnAY
QK5d5EhgZaNTIlcBRJDNdWntMJiqUKdKvLJELdxXCQCDvxIo0pnR9r0jF6McMPVTM8wsS5DQat6o
zjzZgdbubCjR2fwrYkwo9HVXSXD6Dz184bzXuorK/KxuvEoJPFEd7PAI2SyJVvfyqT2yhPPvcWzU
WPJzVrEnkwfHCy3xf8DwNRaYX1G4PjAzV2v0XVyT45H8vDcE+8FbhsD2NBko9muIUN9CqUA7NSKj
fuskW4SAXCKkadvG6p8X8eaQ3s95ZXLQQ+iE05jvxDIvwS1CHRf050L2aEzlAbdsHfmS1kflc9NN
D56yfgc3Nf9oH+Dav4zeyFLPKdwlV4OFUB1KFmTCV/TXR+4dK60MTGrzyfCIf//M5QrybCKH+gqj
Wz+Wk8+j4KyBLaKILFMiEZHSjJnYHhLnDsGQLAXkqq86kMt1h+UHFbBdgbYhjEBlt78bwzsNTghR
bEDJ0bdW9kR0H/2pazgbG9U4N2w978iC+hb5Dt9vI3ZYihEBpVPCdE2I2NtXHw+3vu9LXM80xXQd
1ajxcke+5rOvQM9DfDFXTT9BrnR3RtaF5VDxf/KwUx7PDqRMIIvmeJHuWw6tV9n4BL5zKdlAvnSJ
ON2kCODq1VtfUVusUFHbERirtRY81vHk1tfuRPgmiTMss/CfwO2cxqWt+uQEAEAlKvww9IskItD/
weGCfxDZo5Qk4lDWOO9W+Pl4pUrbwg8QjFJ+T//NgKvQCWkCWS4VF/vuv238LTXXMw6Gi42q3YYE
I/0oV/uHbFDbBSJG2Ak3ohRJqKWa8Lm5WAa/MfJafgAXpSrqoRH+g0FY4hC8opJ2AtjCozt3RHtq
i1TXkl4SoA2e8UzQuZLwAwtru2DplUT/sndBcNKt+NWqFJ8OTm4ECNeYKAXkMA4sQvPN1jNKdS5J
lAFLW2kWgCESwDLzrCFaMrJHuDnii0fH2ofes+jd0EXJFuMPU2/14aWLslxuzFBWNxyYdABWMcAP
S/OFTknWuqJ2hNy9p+5ccOjQVbys3guj/7MAoiVBgaw5hjLk8FpKyeKNIL1svPtMqbb4QFPj5Aij
AsiG+4c9CFGmJfZY9//uKGB+RBm+bTj1hkRNtN0KdJIxQhjGLcrBkocd0ovumB1kcrJ6t00L0o7l
i/HiLTQC/6qS7nvLPRx2SFAJkDhXdhEtMjwo2VVALYo9XWpf8+v7Jnb22+6aUkii8ll4rt/HOXDT
rg6+5EnzMRyCF0eiMv3idR/2FZEkNusS3hn/XdXkUWvnn9rnDMB89/C4ZyCfjXFGL9+rXdnq3BhV
t4fhTmeJUzTeAtn9pREw9I1vt/JZ03nQRo1QVzdC+Qimdv9j5sEmhW6ZaaAtFE2stbLuuV5kRhun
+Sz43U/MWBTLE/gcQCS4PafCCabCoOB6BFs3RnEQGgQA1wkq0RCkfM0NP0lwI6ls0ouxhRX+hoEx
oMwY2xD4Bmi7UNtc9qkvkweuBYXM8B9fp5rmpK1ZWfjDebOADbhsQrECAd3+tSI2x3a5KVEW/vR2
Wlotc72SG45//1A6T8OwXKIsSTgW92JmSbSLRdAbYkDJ1szvwWF85MZzlEe6qIQOTwiTMOr7c84I
IHvuPmbYm7jg8NCxhmDqq9PFAW/jycMntcveLhcJoChp5kaAorRf4CrWRtJqYJVjFgvtgSJGSAUs
akeOcurH2YR0XwWpde3L6IgWssFweaVvZD9R165HAE2wKbJw+BGa7Rax51Bwdjdy0YgyMaYGuwmk
uOt8iX8ScjOnEmw8Jd16ZZRVQRQh/H+7OIqswzjxpn2r8DPxZhoIUaBa6FFsirIR4dcNMZVM1eD/
Q7rxXjAs4bYNU39o6Q8eWCTsa2Sl2ev9ivrKxceubZw2opHvhuDVM6u4QufihTHo5VLJvKmuFHxh
b+4cFbS4ZaV3z+q8hsdN0TRI2DtUlWUWp890xQAPV8/gsWRuZx/JGQT1Negd1Lbzwr59cHP8HBrr
bxsN/IG5xmPM6JqKY4KP7rc39j65P3dTVD1udaISoOqd48GqXdyekdmVlnp4yvQnPLx3OL+1VNUe
hfOX5ICobgMo4YRSv6iqZCfwKj/nXb5XIC6l/GwpuIa9oqZsbvvIS4JyQhXsXjxMhVe2XHHmgoFg
Hp65uGZupk1oJZQztf/0TFSmmpBURULhpNjnRrR82qlvpoQoBe7J4LUDyO7wxIh2P/t0I3eB97z7
AeK9RWTPktLfNT/wWDV2maOAsNKyT+wkU+Bl8jl7dXR9UGGx/6KXuXjygM96LPTzc83TTj1VAaCh
8f0ofAHYsLhTJ4aonPnwkY1+goZBD+gNPSk1oWIka/WFMX8gjkJ1vq3GUaJZ2mdcXDgZe/BRPs1k
7/qNXSdSXLyJxVSu9mRhBZET/RDCtDCS+03P6ZmL/LI8W8cUeNO7DZWinKGrYOqU2Ke0AaNlnyuW
QGd9uab+J9hWS+D0pXvOxjJOMadXXwVOLBLtwOvNza/rvUqBT+wyej+iawSPB1ZVut1ebjvSksoL
VSqWlePfPSR+Sma/8t5n15hJDnpU1BLHPeBMq3O5lhRdEkMAW7MARN69ryOHWjVoWNsgzIqxQQQk
ITyQX6pNUaa3arH4ooj+GsAg5gbMutVJD8Pl29OSnAVS2C7i9RPKEJiipRG/dw6HESzf+FC1f6N1
/bkKvoQT/rU4+5Dx0e0ntQezoZmO2n8HsVptSSTUmI68FqB1et65szZbENi1TCmj+DADQ+HGKe1I
kaG02xcNWA5hH+KrcvKuefmmddJUMD9D5qXMouQ8L2HloRsCgnwQKf4KA8czTFklpf8k3sSH6A9z
Y0VtvBdl6PwOKsB7LQsG9HzYNOU/CwoyBlaS2hw6x3/ZGksHSE/QDYa4CyZooD46nB0DyRRsVWmc
+JMXkObewP+416vugYzeLlglG/5o4vtmn4jJm1l7lX8m5hDavxDv0j8votHgw0l9QqZHVn/08+Oh
8Q0EToFAVDYFYbamK9s1Gya6vpWhaIgkHAm/wiMMhX+4ixTs0XPxpjSsl7xaQRm6w9eh2IsGgJVE
iQxRgi4uLnkX3OJmyoooXfipe6oizg6nKjR6FnW2lyvNnZOO4xKAoOLhUhjFfgJ1Q5+llhGe+cKo
TcKbwG271ytHqYeRj40q2aJD6ye7vQCxv0mexe2CaReGLXqftDBcUmKAZW/M3r/blv5Xi2z4Fy64
M3kBRoOUK7PQp82BZCuJrWYV2KV3U6TWhvV0zF/PH5SqmBiq5YEIFdl/QVgKtgezbv1ktJKVHvG7
ZAkLvEXO3OTP75Km5aMqHo6/nczxBwklUklPcmmiJwM9QZs3UXDhPIlVZdDEhQ7d6f3CxPItVRUQ
2tjpO8fKWOj6uzFEwyoMl2EYv2IMB6Jfxp6+s4U0zlr5+dtjogdnUhPUU2a6Q81MgX0ix/kAoLFC
HPqEi41RI6gkrbTrdRGGo3hMDfnTiEHOvEs31mzot9hx4bxRf3QNYAE5Y7LxFjJ1yI6mD3vpKxgl
b8hRekYja4ZsuksE/+Ss+RsJZqYo6hGBxh3yt/yxmAEEPeUoGnsMXI3vxPg3WW6tXeC75ao1XYe6
rulqG8ULLX6dkEX5Ndx9fVBw3KkkWCfnY7larAfHpPGUehH6fBdIfim7A7e+VBQgYcfoQm4sCxt/
AUGwq1m+kpG2BUYkEOZtn9Rq+qPA67soeOsMT/zdqzNDt5r5ycmYDqMyuIFGA+L98sIR7nVbthq5
y0Vmcl7kgdoi6FfCYV3WFuIxYTaGB25OQCdewpu5M80zKrX4rcmkbZjzfBXiodH8s3sp5h/vU7At
qcz2PeGOjDsk0FtQYeLOa9Kc5HCuEqSagn7fCyB7Bb2tMKmk8wD9QJFcE3TomloAxhtjVDfxrIgd
rpc0XajaLtVDC2oYUBsORUMBRY9bFp1tdiWqt+DrTGeKGnXsqc/ZU4/XyJXsz8NOSre+1qJ5ySuX
1ZVyrFC/475J9+vIt6x2JHEh986nfIGpwjCcny3cxNHiKGBCDhhgMhYHxtfjIzi4NcUMh4WsTcVz
PxfvfOAPrnWkZ/WIq5OZoRV8rhPKsxPTpTJ1k7t3TQUkt1EdjxsWV7zvJBeBX4sshVxigmuoVmOL
f1FvR+MKYYBEBk1DQwRbwJdkUiN5aApHYo4vifLS8VyJPvY3B4McBa66XfYCgC8hlt3ZbAgxxRfG
dolhs/TMTXYnp4J/rysNAcJFGLLiaL2z7mc4jwB6tZVTQtCKZFQsTdlw+vH2Rl5SgTa8OC1vnLUl
gGse0bgXHvnl6EU0QyjxNYM5MXhAFlNfzUEztbJOYygkA8VVjD+z48loP5DmJKSqHdslJVte0x71
LtvXl9yWrFa+Vct5yTNWbKEJgNEjy6Fx8JrDprSPHIdluNJBD03aXmbBK6zuwpGynuVUu5yYQP+f
z1IbNFwgq2XyP8Qw/jFfMXsk7Wq6VdjhoSB4+Ig3gFRTc/i6XfWB7UYOWoYrzGWMmaXjc8WXmLWC
qCmaIvdMSrKDrKW9ZUWfd7H87MX9ZCVVPLLtNliv4EwRV+dRFbB5FWojhectEK2fW3eOWgCXUGZb
EKotpZhK2+0I54yQnAueRoD8SRTigdxd7K3fQ9c2unGhh29MVd9WwKPS2K887J7IllD3aKLLxDZ9
piclh++Lg9q4T3O0Ng/rnFs8kPFdVbwuvNuffsIdwIaS9EzfbbFYcaUkRzzdzU1IO/qKRjE2CaEI
a4+8KL0FDg3fJRTc8eirgjwHaj9KvC470z9StFfzfqnpuheYsa4IQzhbC49B7CxkTHP8C9avNfKt
EYRiCfYJUYH8qMH8hAYQlCpDY6OYbziJElJ8yRI/K7gVslDdyNEQvW4GIZaU5T8xx/p8wE5fptcP
6CN4ni7yMU1bjMVHGRzKN2myjG8XUioVDL9U6jv4b+261EzuluITwRBlJ1Vf5BN7pbNpiq1KA0Se
zk4j8qatB0R/oN4fnEn4Dh3jmkq50yozugY5c3ys1Lm71SfkCaTb8x82BwofU5LVJ+CGJrzXOXxM
br/IRfZiTuVnCelgI2zCHLdNM/UD6yAB/KZRq9v5q7wYaFkb0vGUm7WTvfKj4+KQ+o6sSzYEBN7r
VSaKS2jt9tZO7JEYn4THsrqrk5cI/UYsy30va/5kZOBxQZa4NabEBcBkl8uz/V5vxElXDT4AqBfn
xgcc0tHdjq+pNPaE10O1c0Hfis6mYY3bSlr1iYCNCw+xqWtxtnWOGQhAYfuCOhWYLVwDHx2hVkGQ
YPQ5fgKLnGo7V40UIsx70kedNkZKoSEZ16zbZr5LLLWTx45Rt09dQLFetonZg7RiJTmaqRgyjMpt
JCTzixWaei2PHHTy2jZ+O/9atbrfgCPhRMlalxS2DxVPlWu4D1ppDxRXHN0X29RYDlj3Y4RLPZV/
a4DsCPTVy9o7Bk8LaeCpO+WtmMuxozSNQNCxa+h+zG//gqrVuw09oOyFt+0nC2vZnaUy+S99PqBf
Mqihzlg3V4YuRIhJM/AdHfd0Mu1lP/sUNnj8IeYc4h69QZ6H4WXNrSsHT8SgJAquR/jS+h/YITzD
izfpmGhJEvpJQPYfxnQ0haFWjVBO9Hfn3Hs57i30MhY2K0biv9RwBNhoCRhAOjtoAlqRexFWp/79
fbbMi6F053iV6C2ihj3fws3zF4dpT12Hcu5/aBZq4pU9nYdNe6n6tTW/6K7kBZ/b3u3Fz6TmBwjI
i53440HBIabuxXGdSprl8R5Be6aKwWgE+FbDrkp6xdHFePdX552rAxeCgRJhOAi0fxTfBTvDKZdc
NSmnn7DXCfaXxo3Qzy9SRuYbAQQu2dqJZBq1VYXGZLvXqj7pULVIE/7Lw6zDSSoejYzhI3HHaQrs
C3o55s/uFvTGtDzdWlAM/ZYvBTqmJfGhB4WhB6Ybgnr27PeI72LjZ83KCRNdwKXBbZz3Lrqxur1z
4KnXxVC/2ar9eumnXZkIs62hh8bOC9NMJ2nah3u48paz4A6mabYn7cwwuzA/WfFaMaDUb9WH51mz
buBU/cls0Hb0qAA3qN+2SsQLwKDnKbJfoiqlH6HczPOV78rF3RDSSIUZna6+kDm+RgnVVnhia9Kg
ehmdlPUoEjyTlsCxBibWL3nqG7heIB+FYE3vADgyDFObDtY1ihFtUMsVYMFuRANYrtjzO0pI01KZ
zyOv5F/7BSQzKP4/T0Cm29S4q1qUJJpyYUPXmUYB0r4Cfp5gpdJuIpPIhNPJjs/W3wl2YwAGcDu3
aT0WSDax6nlp726UQLOtKkeov8sQAhYQfxb/2fNf9D4L+5HMcVrxr7kg6kphsBiR7nVHU8+sDp2P
qfbRuFiBChDoqyHx9jxDH1fSa+XoZvuInNPclT6tGWQ8GQt6S2bC1I2CdGlC6EILWKxQzvGcp9vF
lcUbDofOZQbU9IBtyDlPOeCcS+DE+F+S+CMg61AOAYpLCkrUkqnqPIzOj8PIUxyPYW49Df9oHgEM
jauzgD60CuSHfzLTNWa5FjJuJXvieK35/FV9mma2aOgQmvctVE32Z+1qzqlsUskWI+SrVXmi4ISx
oiB9v+QZjhp1nJn3fj//cs56lrvgEpsGgdlh2EeCI/AuRNuMHd865FWNOE63maI1Y5WfI/mRQC3F
xpq5rn43E9xQyqzbURGV5DS9G+i1OANc7DCE/uL5RGnuY0tbPDNKUwSsUOdszlFMtpkjzhbxPxKw
jc8Q4IiNoP+jNoFyNF9Sfd77p7kKU33s42j4KPdmtNYFfCi7RUL5o/Cdfn+AmsBgMP+IKAMtcxUu
/tRokwlXdfbvjGjXKhiClltgEMzxclfS2eCnkkLsluigWdm/yGI42z1TUMSygrseTX//sMKFLcTV
cchNiHiiv7LW953lWNKo6Z+dMk1pgaQu3StneyQCPSAaVf4VhNk+TtnFp0C7qG7CUY/yKPBE/IcW
ViZmuF3EJO6TkcScy4WAQABiVX4ZILThtgwK7WEp4Ke+tOHYKsTihzBWThYlMmzDODTAtWxdapsU
bKsZeT7NSm27oZ1wSGB9waasMJCGr/wTqaIsOM0vYoa4qF74MPFJPtlA48sh2Us/CzYx2gMbGrae
mPgP3BBlaa8+EHHu7YQbO5wqIP+CtnBeyLnMJ5e+el82S4vicDj0UlsCtVwKMcnBizULuw9fNjVk
CwzWmWbovt0FjQPzS7vqLFdD/T+hdxd6JLX7UeDq93MT1JMb5zVHbDvr8jFO74PM5jtJs1Et/kxm
IDD3bKtSr/crA/KCPLyt5kQNm290OekpSLLOeJd21gEdAasSjROnDCmIuWDdmzhpK6h6q3h6EUQp
qfuXNr8sfp9BEHBVc/7phdf8iVNVhMAP3u2q4KtfR2wwzRDv2f9PWSe6a1CVnh7G3JcASJn4TS7B
H1ArKPnSN4TSpPI/LRDihA1NyGeyNHUgY6IhMA6AIjiYlWZ5QWlw7dQbc1WStrT9yK478oV42f22
6ag+VlYv4xhS2l+85rau18N10EPZYDcOEU+9UIR4eM0KE01tymaLvNtAXY5aHI6ekQVtziIP0NMs
UwgQYyFTb9bzkaLkLNChyMsDjZ0IcYQ97kMTbSoaUvWggHgVc2+nLJPLbFo7T8qLxoHqbxhK1nld
FMUZzTinYik2kbYW10oV4d+3hOkbmXKse9zNuIbd7FeiI9CMJcd+ke+qHCFYBAJrFj0PljKJz+bp
Ta0j/jB220CMuSTLreo6BQtjAaZPTIybKFzh1y/zEQ0KYahcOA4NzyMzhZ2NJw+QUJ6OROD1pKuU
P5Gh6ce96q9/fS++omOWK5XrG9YfgWEODU93vzJCMaTewatn80rR/Oi5LznWTf+AxQDKCcLGbpGx
zoLNQETB7yT4s+KcXRqOOr9AJ23CM6gF+MCE3/J8b0poFowtLiBC4nwmldrij5wNyT7uBCJqKI5B
PDiTGrlWaCXEo7ZFEhEnZzhfFf1RaRxxmgDSI5mJppXYjMbXt1RRyXYpE02tvrN62wzjD/6h9afW
ncdR/AN2NGSDuXytR5DjdOZOG3wY4F3c1bRi3Sxbl6OZRlH9aVxkwnLUNBBkh/CnKzMr+l+oYXRv
X3pdH0mYJgRQLgxWjR4asFztefDtOnIyK6/QW2dAiccKGsvd4CTKU10Rhgmk53ZOH3Pg73mqV5bz
E/Bqxztt0PBImCdUFEDgwjdYKmEy3ahDLmfqrVXBKSoRTC9B+4lW0F5vaN0hKRGDfE3aO3eBg0ES
ko43DTXaTUjT8dJKVsDC3YRovO691zEKTKV7EXhaV7Vj7aD/ad6CkJ5DiuTRpbJryonSfkEARwSX
7pYj+UFuEjqIKHdKLvyFki4YRaiArrQgxInPy8NQHLD71xTWU+0bIhP8yq0t50Ps/bEqT7ZIWX7k
8snlz/Mq4+PWYDOghbjTj6mRhMt6mSInSMANGpnRvG/LkCnOih1s0hNniyyQNnmheUDAsrkDAcBp
hqh1l2gqG6XFBJ+IXO6e7Fo0Mf4+WMoXJcLbzQXMP8u8ZKkepHlgoJKbm2MWeS/FUA+XRWsXYZNo
VBr8yOvR/SC0tT0RZX5KtmxlNn226SPgUKw9nJZWkhWDStBj8tb7WWmY9IE44dbMzMkJSLgAEmtQ
xFfsaYFc9jfCNNqFSvDO13uldqMJeN2VDKl+luhh36lm6QLzRp0pN8AMz1s8kTbTh0qPcjRYk3mg
BQyTTm//xzETH2yoRK8STfZOydMacNg4gw80EqwOq7rGQbI1ABUum28C/TjswCAaWBJCyJ3EGNGq
SBhGQRsn+s6ecTtWM42ZWPaWqylgI+dUL48QibxoPAq3hiVRQcfPCP87S1WYFrnPIbYLImF5oO1j
RhvFdfAgpsTBPsc4vLP+xrTVPgYfkF60KK2JjYwAxNNqC6PfesSGSv8bYnp7gW0ZK92ZuoXojlHu
r36cFl5e3qZSsmdOR5VBu2aP6Szji0TRVPqbf+9lWqQbXpm/fHo3iiqZexAW2pNmKznv6IH3F/Cb
4D4C4MgmNgM8zAI3R7gNvsO3DyVXrsnq9zhC3ZburBx6IeEOqK6aMsqg7zAmJ8WtLd9Dy5Pza5y3
sINqU1dwacV4D64np0K3+drQ1esQsUJMAMlhwRlL4Hf/oI2Mc13LoQQvMEF1dwg3ApSzxm3U2dq0
cR4jimQVBxK9yx2O8eapiQF4y7R5jnzcUWGPHyHvDKQADN7btdmDST0yyZfTebPRD143RR++T8Ne
XmQPg4SRA5BzJD7cY8irWeu3+TuunyvbW88PZOL+0axjT9wtN+hgB6J7pYewMdtUDMzNoyC7AQr8
lCkhv1amcy0vzlYOux4dMAzgvsKCW5i+Vu6VGJx/PwKvMKny4jEkSiUMFhATBqyjhcs8gfOCURkI
/FHvfgvLmhaMJovHoV1tCdSryyZC9mc/yAz0b8RLzbiJrzOOFzVLP5U8L6YV8u+JUsv282FrwMkt
MFpa6iYWK3KXmBbEqim4k89DAg4x0s5kWyKrGAO5aGh5sriFPkN+ubQzPIQpRj0FhF7yylwfWEn5
xlNQvuH7SDgAjuQfdwS+++JZjM7S9b2F8zxz74arXNchv86lIdskkWSnTmo2aejcaCk932b+oUsB
7lbIXPl0pmfSSdpu89V/nuBfMgdIfZu+rOaYXjyhg83zsZVJRbDKizfDVEaX2jZ97qhYL0Tbr+i8
uMdayMVlJoqmswk078HKEKq7/DqXi3h6g7z/tImwuiFmeq/RjjPrIHHiM9UzRykMMPreQTGJp3AZ
/Admn27Yt3OyBqo1ZGkhvSlBvzl7HIvI8gUKBf/7HZNNHPYGs9Hl+Avw0sUEQsqD/LlDmtav8USD
syu3zcQxoBpi/3fTCXSVvtsVO9gX+grtc47uQrTUqEsm0VRebL24wyr8VtUh58HXonzm6OxfZAGs
N6Ym8KQBDyJ/GOChcnL4EQ8xRRMndfaBDezbutsBxxGH0mPlE+mG/ksyR0Cu5BK1K18RnjjLdxL/
QMufhc9XObbzr8mt+xPMtJc539ad70k5k7uArCpwwHECOXUIBQQEb3rusovNkhiRA18yEcK+M+uG
Nr7M7jJG59Qa0blqo1yP5i3lM7yS6MS2G8L5+j9PemZgoFWzmd6iH7wCOX5NO0TD5fpeS10FID3c
fbsoycjNzpBS49XmO3Vtq6pQb8eIGy7B9zxl7nIGjjLkw/LqKvftJfs97PmleCFqhrMnxcO/mnwP
o2hXwev19vsiSAtV1MnezT2rqUi4MCKx9EtBMbRJCVRG9Rb4Od0GIfURDjzegfopz/1nZIv2lwic
4tVvjwXjbTLm7G/c824UJS2MciiK2TePOD+1CrejGKR8St7i0gU0wnplEeb4KwQvbEGhityvDn3c
/lp7QZPrxvoKHtV3SUFRJqbb9IIeXVFS+1Appk+FKuwShqiFF+ZnJcBJcPHNzm2H0rt99H143tbJ
2e5UihCXbrsxKzdC9gtABK85SWcWF6D+mXNNvpVkG1FUxX5t+GRFBPoyy1pqzdjiCv8HC8PUdRba
zfuwgDKP5MOUxf/1LrEge0HKg027Pxj/iD0mzdz4LVDgsYHU2SMlmwbvltFV6oPaSEN20NHav7ki
o+ewKtdSRPhPrFW5QCYQD0gsdT3R1axlit2XeuoXIeExlrNrswFfS61fgWjc3D6jbo+FwyL36Kso
QQIhbMLHjGl6HOC6e5MOfAOZ+qGGocBvPbQknKTNlNsmyDjtJXKH7B9tt0cp9GXhsRviPkq5M/k5
u5SMj/f17SDvwjcndzFaacSDBSYv2mnS8i/bu9C2INbjbuhvcOpoLv9EhEIeeJIbOJy48cIKVy+I
4ZMUhNuqrFR1zvapdv8xR79ke5xTVTCIS7qXH42RwOBPH5NfBui3Lxnbgg0y05r8NOZbkb8t2cks
6cIMAX8p6DJjk/xsXxP89r/uaWUgXNw1NHjwUNFamVkJLlql/QFE6Vsbo01Zg2d8zeFztC3qVwnh
Q8QJTZDQX5+duo4TqkTc6u0nTUJ7gqHhMMslxnUnMz5s4mVqXVPiriBn4mCJkGzKCyyeRbfaJQsN
65VQCq5KhsthuiUMXWF20EII44zqqfYxztBvHs6AhjR4gA+QYFgnUZn08/MP2SUwLtStXkFqcZUq
65HMYp7S0A5SK12jCgmddtyuN+wDZPUPvXWXnfbtRjSMTLgEnOQZkPqwi/jYJTRlSNLt4Xvu4q/+
RyOrwyy1EZruWwS8dT/BjBLdZaac9lvUCN74zTUxCcYPOmi7ANgTiZzIqzjhu5PysEPkBNiDRVF0
nn6aR8lM74/EyrtdsxngIk/+RL1budC8pT5U+9EeWfZ3mPGoDYCAIVLeMqL9NgJk7RyPeyG3/XRB
M6BnILi41aKrbGy/bccQs8dbbdqHdjeK2/1XhaDM+TFfYwt+Kx0xy7N+f6DWChrG3TezR633dgDv
qYnLKTUovHo4JzUOjizfpj9EIdXXTa0qHwbhdxRn2Lhr9z0FZONVNZ7tpLEkM6W4sPEpqIu9B66H
ZSb0+2SoOcqi91GS4GQ+EpCGpW6axLRRX+R4tTb/JCaKuUcKusaoapi3OjthgjtIvmY6IKQeVfE4
4/UW/WSmkBJSCg4/fk9VhOhvW6UYOmKPr/tg9u8DFipoqmQNljKDXM2ZIw4Obj9QnKhKWYRDSxzI
LQUK5ZTNDaJtbJJOIWtnrdR+g+wCnX12i36S1LVIqDrXu5+/ZwfoB+ga1guBjJf7m2PBZD0VIjqi
K4Gj05xOYcjtmz10l7HqVifPYBzGOeXzERkBlTgWPrD/PmqvUjBQ6Nc72Rw1d4eOPC89whezqHvI
wiuFmpV91zAQ3KKiFlMo9MbX+bWRF1RJrQY6elU1YQUBywCB/wNDEosR+hXMIYtjGgFec/jnkw7r
lL6Gz3t5f5bVYYWA0q9YrDLpAHUxlZ0Cwgz0ct+Yp4DL5cxIgHbf6Nd620HepLiSs9s8oHf0+V4g
PYrcldCTHAQSLd6dg7RvRWNHtTghfFKN34jm6AxcvyONWhcT9B5icoPQT1VrN5yd/m08c9mhpZZw
x2iJ3aIaVMekakHfG8+hBKMxGS1jWIJzQMxgsdl5CSlThqjpCQHzlkg4w4FYUe+mbQxKmV75hsNG
7SL4yjQchiClqDEZyrh0Ew1HixnMmBh1gtmqtTtlWNGEQc1CKQHqmhLqkWdXJZArYUdMslU+xIsg
TBdy9mJyLZamSXY/sd3r6SyhJSIfOuz6j0jPZ25ysI/syhg55CoRA4w6T1evJc+qU6GxPUXNOHv6
iDqEQis1eDmOMObtSHeWTnGnOxcLzvB48TIhhE+D1N6XM/y9pPtTgXSSB7tJsxgJP/HDYDuSTgCS
ATXeK367hQq0NtJVi4wUuhY+oZy/Qco5/Z1W6T8p+ICovsRGO/gwdK3vylAECQDeZQhP3E3RiUuh
qBhLYEWvWmmv+yfM4ihyvAO4nFQuMc6Sek4bFC+BavBDQg6nhZzWklvhLSeGRVmY9ESXb0dMFw0t
Nc9Tau/qzCNlIp7rBj2kyq3FeGMN0heH53ce1yUoqaYF/gNxSfj8QgSQqA0duePaINQmNtO5ZLZV
gjfHpk49LBmqH5hDRJ2HhJAC/MOyZM4dnvl5UDJsvEf/mpwLXc58tL/cruHcC2uZQ2HTWbcf5ClR
7LmKpFfG4XbPHIY+AyUJiYoCkQ5FmU4ebCXq/JDJ9N+iaFKdXBxwB1iR5P21wM/LdyE6kQ6paaAM
/RXoMLxoj57AhR2wJO6cZzvPvN0AueXUnUS26NlihRWo1d6LhlwtGMb5vtnMXns6YKC7wfxi3G+m
PW4dJEtJ5M8elVdyovzRBBR7yW8Oyu0aN5ig4XKG8v3lFDkUD9llIVH0TwgSCKv5eO+b9vaiizHm
IbEkI47v5KpvkvFW+rULTpHsUYhEaKI8/pXNzOHl4UkXJsvMCNLAHr09E4j7kmeD4HEKLsXgUijr
ZYExmRLKVt/urynaUR85vCxZvleYFyyz8ITlwhOKkbu4G2Ng9QtQY/9BGUmXt/l2sf/hfCTsxEgo
8LhLvkX6/wB/qa6a88yf+JupiVnU8EZ7vdTSPVCHlJqwlT1UL+UNOGk0D0rikkg7z1I/WfI25R0a
ntaIel2meQXGwq1AZFPn1yWDuZDmg1OgafQ52vDp2iAJ4yQVccUy4EdcJm6evSqaiJ7qHnjK6qM4
+cjJwMjuD3KRTpPy3lpVtyXlroJkXyQMS/yDZfbpqaR5PnaLupH6ZbhhdG9peUvzXps03626qZFX
ZdlvxGjaADdzTaAB4cizKqpflSa81dBHKeFFwIcZGurS4KCC22IDZu7CDhfBTOl2p5DuHTrGEItn
mO0dmYH/9OFVEG9sakzVWL/QJymcgbAcRg6Hf5x/yaDFl1d2HHBXvI32t5kKvV1TcJNIANuB0bIE
Pa9bRwQsHVUx+f6UDdTAyI7GwdIB8N+dyqoMYv8Cp/Bs2K7MSAEtvxvJlbHaAJyKhklDz6hb4Zkq
IaX1u9c6CtN4e9GhHrb11bXNANOFCwAOoB+p5RLQH+ISi8oOCRkSBdjflqHBEK33CZDW4pxSJNQM
7dnvEZCHVdnLc9KoQVRk1qYFaRaX4S12sz8jswyicMkdNyzBy6IfiV2LSqqwxJP7Bybl0fE8OZja
lw/wc5zfcGmmcNMrHZIyoVc/BmA3MW8JS3JAG8UASmNEaxd4sqPmsL4KjnwLBqI/Dk2+yyBmQ2LY
F9z47fauJkn3P1sqEe8P2fqDTlpc1/zdoIqxc7ynPdPfPxKvoJ74D7UJTFwhMqMFaskz6iohC9Qg
itN61R8OWZzXU86VIlnRoG1BXlOCPPX3qjsfx917DYHAnhAHG7GM69eUy3qmHfWaCZg4pJp6V0RM
T8226G/EoEgXqmX6K7cavSnzaNzYPvn0mlKSCovG49ACXAKb1qaOESFNpHKFUTXlV03LWNduKUD1
RXQ8185/kgyVUNRGY8fmal4WQkn1Q8t6G8zl9viDCkgXayW+eQ0cMz0EDhgXF1m9FD/QLu8QwWjE
Rg0eABJ77GQdYgHRGLZMkPaI3OlTe54K8BkqgMXiOv38mqfyr5wvH5MsVr07ERhMKuHN9xkBOIr1
Uf1UW4qxc7G4Roffr2jrawjtyy8cR2HVDCgXHxTmJ/VcAbv+0Cr4lGn3ysTgRQc6LSHnWx4+HOzY
7McRp4D7lqOav08vkHG1p4IV2CdPUqUZVhcQ5wSjdxThx0jItydowAS7Vi5S1b5SfJPS2n47pGbW
bkW9MsFrhpaVA99zArSNNDRPiAOExN0WG8CBLN7+JkW9IV79GL6z8JBJEyTNqhzHv/sqRwfRz5yM
U+B2eXwZpvLzdAR/F4A9KPDW3i6c1/jIl9zowYlwK1NP64JRgSy8PoKoYVyV6qXvVdEN9swOo24G
0T4YtpGwR1RrgThrBajLgWlrNlSh6elJRorjvPLB7QSXrIPZ7Ap5oiH98JprWHrvXMlpyPqyVdws
DvbLffSDbtSOItA5QBJ59l2DjyhL49NlUrctgeI9iurfCo9qJBdrje1Bb4Q+42zxGn2l2N3i1UVm
dxIbRHsDtvZ2Y6HWlPFVHZonQFBHHMql+nQFOPROcuXLRgjHyAYgdSChsC9fYTt1Cl+to1Grb1++
EHhN4lKS3cldMmY76AerLgo0JCajmRCONQ3r1n/gxofIjSr2iBxxCKrFYxB1Cp6cXNBU+ekdy820
JpkhLmeQJ/xSXZy/rlzFRjGibhx2Bef+CfFGn8igHRn4ikSexcifPnU3h9APwh/0tJmF6Du8Z5TV
W2IeRO9xOhXq6Ztg6nbBFB3xYwMad+YytJTZKTxABcSHe+ykCJdYXSHw04Rm4//YOtzLrWXmPt2n
kf3YjUlqvsKCYC/yDkund4kyMDPsMG+SppqZHF3Gzr3M1UrEXAELyP/0a1TT1D7FOcoPJJf9BEQO
pAE0G+POGj7ALTS4jny885C0GjKCkWpOaOGn58+dpKyR9vZQepX7XrS4KPwFK/ItY50yVahn2nwJ
yPXqkgc/SHqbIO+bn+YFxI1Q5s1XKfu0VvSPqnL7nQa7vIdTaBCWz4HriAbP9wm/9KK95ouAnpAc
HpcDQiyijWSc842NjcVwBMDnShIok4v8thelTz6CuoUCnm0rm5U7ODpkLYUWC+N9ey7fHr35HPKu
ljbu3lnyizb8jycucpMHX7astzGckP1/3JkFJpYZe3iSkR6t9r8dgBFrHLpFoY7hTH8OwNrMcGde
G8kEPpLyPG8X0f7Wp6mB6YKimP0iLbtH1e9lEajKZ8b1notMqxyUIx7Rg8aw3T36nN/b+GBkupbZ
BoLNlG7Q2D+0Sxu+d1cM6ua4WiAEgLN7cpXDLcjU5nxOGLPvrHE/rFNRPCYuxu/3rjgCraR0l+ao
T5kPwmXmDPWkWtix4TcspoYImH46WKNCagFqDOz7SWnpJ4FyRtlEXFTOxR3fIxAO1O6f7KPvM0iL
1difr+8f4XxCUBJEPgv6PmT0LgU+8df3sTFK9DmBOEEQu31KzwNISHPym7msz0T/SdnWoDRmcctq
Rv4FJ1IAHjr9K0A0vXz6MTkiisQYylsrG72B+UwDMtW1K4fkhIGYuHHsdNwnfj4GxLTsc7upSMYG
0+XqhnugnazJZ5wzcC6ktbxHd09VXAxFaPjh4wJtvfZ/9MHEfoeSmQg88DIF8ik7qReVaAZJQ3hh
H3fjPEWzOaOG2AmGXHF2PSF0KUwLMMN+L2cf//Oushfuw2lqWDXd0ccP13ht967g9MTILdB7fuhp
RCOpBqrt6g8F9XLBFRXC7cGiXix9wTp9Q1BKqEQR6HCicJX1UjgOEY2UlhQ/mlPAwk4lAtmRRVMI
Wk/ccDpjCmp1jQNv+ypOwUiu7CRGgmWFCWUqBafiZlXF3PmXAy/JJ/e76tH0J7vYD8MpffpD85wY
fXNKgT8BgGiiRZH/DR/z4OL+y71HWKcN5qz8U/XjxaJi+3/+GWe9vsXQObgJXZM8vvt3G3te3T/L
J3kNr6YBP0TyTyOrLDUZbyKRlT7DgwH36nzN5HoWV+2jgJVj5g4+daxwRgqRaH6la1lZyS+PBndj
HT0ZO+j19hifjwMeUp7PMzwiUxvW5Pj1D+vW5wjb3F9lhG8IMRRxkdXK0kZheDIuFFImThkIm/Kq
yadDvT+OyX0wZPBpeq0CIIViuKRHSdSEGcIS6zEeU5RIKdlybwgG4EG7NiwCguLCfOB96v2BGZE0
NKxjf07+Gljk5R1z9KDDbC7POFN2YdMDdn60wBCN8aLsEA585q5XE+b3SfEUguWIlptepTtiR2Vp
VLoApW63OBhkkxqWqhm20mArSrgz1WIR+8hVNd4KFAbI8Z6rMusk35jsYzjk1gba02obgzyBCxOc
noR2y1UjuEbRkOQVIdHlMHpAOmEFVwurDIXgL0rm0YqIkRZnL5Fry8DuWdm1IANYFOOn4YAm7yUZ
zLM5WlZsYr+pwze5mFn8bbm1VQb8eWzyMkyvwdEQpssk7kICq0R176qkf93l0mYStok/BROB9t5i
tkUUY+EtC+MZQduaPe3IFh5CyGhzjktJFsGIN7azPMtg5vrWtWy+wbUj7k1jYBkgeAzhov1uSSRD
wYz/9jU0fzNTDWF1cUNd8t0x9egFTTQbUEniLSaVSp7CKnzKJ19G8wJPOHC07aZQhDDtfI41GZoN
7SU2wF5seqXJxGAcJMldY0nnPxker5ZOFHRNF18JECs4lgf7PEriaVpJfHDPvUO8l6joVyZa/y6R
f2UFVCPQuyURsDwaUCJtikzbymtzvjIGXiNASr+WtkR9iTOWN0hzaWO29LljxhHLHgw540pAZFK/
PR6Mz7Q/mT/ltxoYbsXcI9BeVQn3Q+yuyoOg63rUUjhoTRvDgT5o7ET6OvzQXT41Xz1uLBu2WGpD
AN0OEeLR5DPvvodSOQA0CYu6RLDs/DHXQEi9ves7OJeVeifIYEj1sQIQCMfngXnEMV6Xn6jDesxH
Wp61cMwg2TfC3pymJFE2NqccS1yWHbJRhd3TIVjIXHnuCmxXOUhXaLbbXgAruOVIoQ/cBvcGS9B0
BmJQsJE4JJUR0b9YvVFFTwk/bVLr9UVSi2f1/iAmEGzEo7BwtMZLaG4xFAY788dheN8ZVOnXqC+q
GnUbEKagE6bkNkOhBQtw4k1ZCFVCB3M/64X4FbyDckHqBUn+mhWbdJZoyIekTOZ3ORONcpAoOouC
zSpgsUjTFVHcGctdczj/lIb4/qP3SF4iOf41J1NXJcqdgJ0Var8Z0MC7TCQQmUnWo3tTsOHb/M8C
fL/mMtRmRBbe7Atldu4/iEmmezDeDCQ3hbPHR+qRJGJnmEXyRQuK3hbxWWD/HDNxzoTPlE3z82bE
Pjmwy++Tplw5LGmnOAw4PzeWAC4iuZapaf46r51vbV6yQCMn6affj311sLZsg0oUFJx6i1BvCy2l
endfJa1mKLpvfeYsatKMf8K7XEpltbUaK/kJFd9NUSXw1HbFq0aYf/p06DmSEseA2LV03r/NWWnO
J9SobT2/lejyII6udxryYA/osZMy/XZvfjVsRxBHTZ03KoVFKz65sVd+J7gTvxFjFZwvjemY7chT
QrFlFcnk1tcC6bO8KH3L0Gi/iZuUAHFDrSd4VTwNPrURN611TrctvoYKV5N4HG7wKIF7NWaksfgQ
Kr5T1tx1wntLtZQTkKz22I3VAUittiJ70/bzbsy7zovVmmEzPWLSmNoq/8Wp5Q7hlE9c0M3EuBtk
QqIk7m2snOWuN9MrcW9jZNIoAjh+MjMSDVgf/PyU4y4nOsbGmwHj0Q4nvPcJHA6PKMwtv+130NrN
RYZG19qbIUEoQk1D0LYTYDRlomAUaVuXZSAIlyY1cFc6ZP3VCRm8MHjamoGmhmboHDgHO10G8qUG
uy5R5sA/3uKXBQW3gcKXZ3WZmi1eiqt24WTfxxxEtiDCnGfFG78wNDeJIT8ymRSy5/q4uiJ1+/Hj
9i1CwqDLjBG85W7mHgvyXdIZeTQ4Ey3xqPQip54gqyrn12NcPQsa4qV+cqlW3zYin5Hg7OTI2zef
qUVwMX4uVKwvGNzHieU8nXOQq3VaUKbzv+WOST152CbeEwyUYHgsrcW0ZX5hp+4eKfD8niUbpo0Q
7H6/gFjgGfDerUliHCYGuClPKNQOaj6SNH9JIhz6vlM1hgcC7DPNICwvM0MTuBDrjWe9uiefVgoz
0G38wdzlWCiX3kLQUZPe4KtsnsSK58ueaksmh/Vqp2DyWOtEoqv9ibJ3CoFr6+Th7miKOD3VzBlp
4PGfboi88aHMIXfvYEM6vI7gYBdpwJqTNAqgUWBLGR40WGbbH+bwaIumQ+8gtRec46UyNhCGXMzD
qzXVEjBkxrTTxuOpzYh21qyFjlLYUd7g85bPiyOZqr3QkmeJaQPHmBCmUzQfPXu3hPsP7nG1K2G/
ey/2vtIU65sK4j4Jy6c3aaQqyD+EnrfrmmSUymhpf9nKEyKHkiDr3itNyz+XgMa38I/60LvvzCTy
vRPr1PNWHNoULvssmXFE1FpZZTvq8au9eLLKd1JLgYtpLPqb3zhxyU9VI/jw9OFK7PeYWrRm7mVQ
C2whrrabxWN5ymmWzLEhW+QRT9uUeeKGJKcQUInQCIQGDY3IPHrooEe73ki0AtuMph5QoBQkblKA
ACaxYU74gzdKmqiQxmbZajx1Cgp1BNqHXMQI29/fa92eeUI11VNzu3HLGkfnUeGJ5c668FaFiD3F
znrPRrGmdL8I57WGp+0Fk3ZKdWv9HDpWo4um2Rtgbs34Atq5y6VpQShqwzUNna8f5RbkiMUBGUnm
iHf9YOPKQ7nP9izOw/Ccn/0h/MmlW+n1sZC7FClI5FsAhjiXCaHvku1mKVvMRtE1QKVVDdK6CiTf
Kqjq/kiqOXgNf6EzFJIqn79W2JmqPWRskiEoXiQufdTEmroJJ9KyOgvYz0I3A9+6Ov/xPoW/C6hQ
BPOFmNNigDAAQ6qBbcyCcI+2PGVELUnCLToBkaYohkljMR3NaxzmwDXCXyTdj5Jf3VPEiIxDWFC9
CQKqMGqi5cAXoAhJHjp2PKwLIBT977p3P5L3rS28I25eBfKX6hZzgqQ9m9m/OgW0boFrRBCEJFaP
UzDwK1NjOBALQbxVAzx53N7r8IVNIdP44RHAV2RTl8au1O46Bfbj1i/0JkxSwdwRY/D/LJeX3SZ+
m5OWm+n51CHVVzosT2yPrru86hNU/DrziqTknma+PZZKMAtFeNr+EbQTOebwV0uYOKvzAa+0ZA3o
PGQ9nR/DLcUiHn+pmS9H0a0lGLe7d2+ctkPKIPNZaEDw1kBFKAl8egpz41bYQ21ufOoWsYb/hNOt
fkB7ZqTJMc9hEJu5rEiu6IHEDrHFI8XWCEhr5pTxQWDsPQScSE+CFSO4KPjSr2AiKiM5aPre2oqO
Hvg1ap1RqdEdUA9ZWSzqaPMNd7/CVQnXQ5u7V+hS/Kyey9QGfKdIaLZCEPOZwwWDZbLaZhRHG32H
HBHDzUuSkyWctFgC/BxXwqOD3NLP6m0+ahbhZuNSIDGrtVErWApd83umjUmhsEjpJE4zCHH3YOfV
oZn7pf4lhCPO3Mz6KMkzuqWTbKk1qfOPt72ZOtDE4VCJMb0Kf036TitFu7uSLHScbsBwb2s/ouwU
gMI0itgS25kXQUwJibqAaUmZ98YygVK8jHrq43yav+mbGoJ4h1R2jvaOHenvH8u4QguuOiBGXCpP
9ycvSgknG1nRdhCsE5IkHixYCXVT0RA1DFSSBmWDX/2Wd0GG9wjHjc0B+ig8yOPhxY0waN3yhQ7q
Il0i7TeO0OIA3RZVyEXxattDayaOrNtEd86Gk2ZE76UzMR4uxOYOxtcU/TjYagapv/y0gFmgWcq9
MEjncWpPynfvOhEQGuPiq2Bkdy0X/TcVqhjNb9PsQtuoPbCMFKF/cIy4vNnv6YKfnDoHua5p9GLr
I2jSGq12clsRPki5qF+1AAzf9JjA2Pq5OkxxxBgY5Gddyhc8V7hOAv89QBfCF5ALXRS0ex3YtKyx
8j+kSL0/zKggBOYzfb0S9fhIvZK1f1gkGNfKtNUoUYxKNpFQxNgI9rSQ79ABLx2IbCehrK4z2ZOL
VED1UdLqC8loR2dZLbDJ3FmSn73cQUnwSoe3KRW1DOt7WaXleThpnJRh9tWjttN3KzmUmKtYzVpI
Z8AFaMdOg1Wn6ErunMMbbDlvzQsxMa5O9fW3UGg/RNxCAFiMwuWL9hOND/epm8sOXBOrKDQzHH+I
847f1fbPUCWjHPCaKsq7+kP/FGZad0fV9WJro4nOQtTZHq77yNppbkKHFykLfvJsPvWXXfgpWQZy
G5suEWsSCEoVZIwBKlSn3Qu60xM3OXjKusnPiwiGVY9d2TirfgnYQY85knJna0CmzvualIY+BGbi
FU+2WfbDvL+bHr8X+AggTsVJF0+Xd1+dNjXHSGwSEY2iQ7C7IL30aFI7x3YtH0dGrRMDu6hXn5GW
kRQuks2nEvRFpvvVI6CnWDSThj7OE1Qyda+YKvbQdo52cFYPekv64msdOcjeVYq6ObP6HO8pGPg+
Sht1RaEPSspoJkdCR6iAv3FXzOU8FnhSQ33q3IE4sR4cyuZDpZ+QKZz3gz/NKfUb4u/EHROkBoXY
aDaUkj1Utzk2MKozgcaxrzcBhkNQzZ0in7J22fhF27lFjua3f4i1LzTdlOTXBLugcvEP++2uJK2T
Yc2my9nJk/uXxa+p9ROixnI9KOlIVBYwuvFSbeO6RjcJExHJtsufW42SVHysHOloPAV6kEri9IIX
FXQuiO+JDEXs/Srg/EIUv8gzV5qZ2+OMY9ayngYGhRZ0W3cKAb6JzlcCCv/4QqiD/ELUv0NsM1kU
khxY1od2wrqH8dwUWZJGdLlKJGbA7c1GH93yOBaDhP2/Xti7qyyjQCuvrW2KPQu9eQyEJkzAM4MS
HAVkcFYfiTUNPHpreI7kAvxyRLAXfp8oXnjPsApDuyBui17oZMQ6LAGkvySN3pvX1yzO7MQF5nt1
Ggb4LY4SUVaerTkiaXXa7vOUfBfKEXDgV9kCJbEUwE2U2+QdNZxMly3VKH4l6tvlBeULFW8v6Z27
wJhN+Uv+GPv843546uWYXIGXsODByAzMOeBTyS7GTg0Q68EV3Lmtu78zRyMZuU28GhMPiC6ESyas
JmJaJCulXjdVZ3yU0thjHeB4TA6G+euhFa0CP/jEWuy0kvYFgMbeu/glKXpaihfAcfsOoAIw7gEc
lCzELBBVX7QQtXZFYaGE7iKu5qtEccuyqpgMdwIvMgPWb/h2MJX1po/OU5DzNAIHFs0Qj8HZ/Scv
sMpFYw2oN7osOUE5dti5SZUiUH6R+SDpumY8kmdSCgOE6naxoRjcaVlicZE8xwl+fkau2idKBH+X
AxNaw8oOIzN1wCmjIghlQs/Gx0p79r9YVhAgJPmO7wppEd18cNTu43hzChjdwPLfTWY4WH8Uz2xW
acT0jIeY1LHa1H/B+hWr6genWIKNZ/GP1XF/wtVNTEHIcv29611iervEtPCbuGiDuCtv0C9EcaZg
EXCqRHJ5rep2Mhw7Z7Jobb0LmA9gOfJTqxoLl/jeaQIzzWUiWV7sfi61FHZZsNgS6s0BLB5bJw0h
q74DUWDaKO3OQCbHoCYY5qdQvcehqJ/e9DPipXyVW3jDiQGIrXK7J1Ma1oU0h+p0nCWPcfxI3Gd8
aIW3c5Fhi8CzFF5yUStLhCe7Arn6YxknwAWXwWwYzweWElVy1aPkkeRgl75uAM4mGCjQFkGtfAUP
9tGhz1t8ywfDLU/F8Wgyqb5fCh9c3fUgf1cL6r2P/i65ftE/RdNOyl6ZIzI40NKAQvffEOaTwsVA
qN8ZU46C9KQFQrXscig2oEMFAZbve+UdCfyj92WWOgS6y85giwNih20Hc4nrEzh+jhYAlRyVihfS
y90KlEbZ//I2VHNDfFn/ttRUGDFHXiDsmhUQKdOw7paxGjV/4hogZ5s2o3ntP41JLqp0W0AVBEhe
z2EcYrB8cbLENINaxdNbh8WcyKzJ8rVbrzNwFfoEeK5IReW/PITifhUofO0kZTF0ITRg6nMB3nnI
oEaxaSeqIameJw0d7hMdo6jinGv6SqfLHAq99Q6LqxpOeN6PyIOlRc1Jfj3GF5Tk8eP6plTp/bGh
eaYArCj/sYz8E5zK8+m2UHOriFbLjqjbz7IGQ7W+R+bkZaOhVKW3ryxFLjjJvO96i/KrvEECAGYv
5AXSRi3HgWBi4bAkmLZboBdawxLXN62rr02Bhp3WMzgjSc3KPV5ByQB8PFIkkIkU52SyMAVSJKvc
0U8eeMYZ39ds+FMxfFopnoPAxmgIbN0fKE259Y5PJnNqAl9nSrAD/6/FBcHc/vsXK2FLyNjngOff
BAjs6wc7ef/OozKdPSfYuwq5bxBTslEQQv7lomfkFRlx6NR1BiN+kkuqtJOEhYiSXzrkxlxBk7ud
lgYlMJomhM1+ZCDJxnhpcWw8jXEMvqxo2Oh7eHFqq8oms07JDpL0gGaPzCNVs4tafUX9LZ/IOmuI
4DS33li3CvT1FZhc68U8nbEjKtKgoko7chT7cuRsEx4dHpGhdvjTmdYLfMzx+9OiEnzm0lSwIa7C
ON3beOIvPUvgkQaT5EN8dVnkOr6dfG32Sxubnws79gOQs6uulOC8zHKysZyZqysVY+Cp4MEgAcG0
L8hLAMzsmSfgX6IvXE64MEZt+5n6qIQ/iopIqMXcsCKpBaz+BAKdbFKCXgfT92JTfFqDPSpTfYCw
Mcdgbc8W+sFQbBzshrNs3R28gTaid+SNuUSaow1VaasW3g/uzsTBQtq0+vWzrmsZR18eJcfQ0C9U
OwcIcykFLQZ9OFYEFz60CbmI8ovEmUFFEifbUXRB/hFcKwYPHWn5LuPJXEkFrWwVS3do4QElw5fD
eiExG2k3z3yTw3D5t9YWV+zsNQMoa0Z6ZMZIpFeVb7QLe/zAuOhXzZKsT/aL6VJyM9V8QM6xve3b
JoOv9Xj5v/qplsFEODEgM6amVjKmlMTrm591eam/YXcdeJsIdp0o9CNDMqom1uUtFzgkB54sxWTX
9wCs8NId/LOk7Lqj6TeoQCQeP9mS9SBMFhoXS015Fq2nyYhPbandhyOlr/FJAIxvdaKoNQY1wTSL
L009dUFKG/OPCjUVaFGpu67W6zfGMECHC02Seu6XsVit8M9UhOj/mV7JOT8PsKYV890LnOxxNLzK
Dx/+rU+DGHams42sYSiDfBiLMeu9FE0Lzx8+mgYjMS7QOYKN+X6ij/FpUNql4hNA2YTR96JsivY3
vTTAYEHgWGf4xeMoov0/4ImKeIAocFlAEiNMeta/KluyEJPWjIvGAPkNBGrICpkJEA24CjjbWQOB
HbyeyqOuk8fTUqlOWbC3n3V8cvVGw/G+ywRkRsJnB5lqvD9AyIQ1YvP2ikWQt0CF3fdEWtnqifT/
N3CIzIjSARSiyDFtFOo8J9eiYl2oOc39XDb1BUyyPi2sIeiEAxbfq0Lqx560iIB5GbCcxJIkzoy3
czz4bOPwr3kcigi67W0I9AX/KkJ4OtI8VNu1Nc1f6cie2X/0XtC3k7Z1orXpGoYhOKnh2rOcO4a5
M/iG2Vbgsz3tPrHWg/ipx8NVcGENzPv3QuUIBDKp6ZLnBUDFcCARx6s4SYmBLPuuZgXfZSZ7sSen
dDpDt1xkyCZPIxqfhaP8XmUwhi8arRuaTAdIt/K+6lKv68bW5ytyiqq/eGRUdAR0CvasUfgumvnp
q19YKlEN1LuKpa8SO09vizovzG8ZgiDBF0wWcA9X37szoqDWmOc5Bc634p1KHdogDeO3b3m4wb9Q
80+bOJRgvlBaQqlwV7aRGEAs2FmDb+wx9GlDK44G4VArE69vaEUOWQJUU1VU1gh6FOwHkZJJ7M4y
DON9ogc9fS16SFdyLnhQKJqGwORnhZZvoDDnU42UkLV+ELg9UOa6lyzPcJxu6QytvK02oVy3/zDI
ZVHUjn1Ved1yn8mXelf5z7Bi6D1byB5TCkrGgWp39rFMahSdpS4d3/l4QXf9a85EcY5P7NMHhlrp
GbdrhUxQhGn7N5xmu+FHcNxWmP2eZuxn4te2BIHl6fMWc2LjD/wzAH2OoWodBz39zSpm8SOD+jEu
OYULRxsmUp0BsQbdUozV/x4pIsGRpqp4Hnd3hTyFRtC9AUs5Wh1lzwYLKU5AFKWO89eh6QBzxgFl
eF/4qUweirjBFqXoOAaHb1KRPDQ1BzM6Vof2Vj/Oc3SSGqqR3c43iIoJ6/wRrcP0dcnAYHm+0got
8m3BTRwVCvwgGf4spmD325zqUXfNCFdeWew69uQyLEq7kIVpl5nl9uFcuZmoiJZdJTtOneGuDxzW
pQDuBpHzg4USkZP59zJHMy3NZfLT5Uh5d6ZFOFhAJJdCtvimwQbjiIctqRLuZRfuM2m6BgQbyn00
RGKAriUf6GcBbb8fSB7qjsn9bYnbIT6XWLsQVPHZarAl/4bFYtRawj6JL9KY+3iASyb3s2t7RSHG
wWAxtwuocCq5mqDtgcYso19E/PZzoo+o9Vt2uP8V5y/1v8seKZzQd97oN9mXczA+IeTJZa+kKf68
kcZR95+gsRjbAgaSW56jpFulIn9xQ32POesPkPo27jYHWqwoobuYwMuHuHcMtDgb0WLOokxknqR8
nfJMk/Xxeq3YBGzukNJ3ldtg0hAZUsnEsVy720vjjENAltfMeoRJPeLtsxr0M2Uj35FrwFVj2jX5
2zZFaS4kncz7amsrVv/xX9F1+Y78Ug1h+1XjhqllLM2REGzLtcDS2DeT2djyBMbRELit2q/oTO/8
YICYt20R+rHhd332bd0fERnszBOIwHoiBBvM5CGfABWSaRWi9NIuiKCVwTovFUQP2iwW2yj0hrYx
CBzaqocxgnvBUOw3+fDsoglc0Ebz+CDuYCRnw32KCFwplioxFIYooH+RnC1xJbfcqxJghPlPUId0
+dSd7p6PnOCiGwPwpYJhW/vi89pgrs+38ebuHEPrbLt9VGgF9pf8mSg83K2HrtKnlEBkrS1qkwj0
E1l/1+6Kk1MTRyHZMfrLSMHZ05bKatSlY3dkqf/5gO3r8IqShF6pWcNXYVpXTIp2mi3GbtujpOWC
8iO7hMmjN7f2Yq9K5YMp+iPxhpSkBYl55pvTZWPOurG2VNGvArDDYjkIDJO7CcLec41g/LaRG2IN
yN0RUy/D+0XrmxAke8NS5/1/q6WCJdfvM5/W6hKV6lFUoHN7IWLGM0hqXBufjRCaMmwTIeCXgc9C
b/rX7Nd1ySLHFE+wYHWLq3Z43tLDDWZhZRwElDrlwbDLGJx5quOhtx3Y9A6Gb5xAWWiQfY1jUCQh
2rG0lsGV2oSwArXAb28PFOM70vtoc57apBpfgIa6ZM2vn+2KIg2WFUdv5ftI4scAqPjl9rm/98Sq
SkbV31HdMAXD/emoXCHPmhK8WfmFaukMk2Boa+Qqq8u6Q2U5f3vWKjIxpL2CpY8o8J/cJvPclqri
FejsCAM2S3qZYkFnK16hMKaGNdEtA802O8n2u3cadm4TAJ616nfbpsGt7+/JzCTBzMqC/lTjtQOt
yY0jdEa1GPPQsz5YK60OCwMVfxve+kmtbbUP2JBqZAkF5w+dFkY7KOuTZxOMLi6/7naJXSUeZ+p5
LVoKVTi1gIs2XOPJaz4IQ3iLXsTKp7Cu+ojyI1fREHh0ay0L81KCnI4b6HF6uyzPdjg/8ljexybz
5vSFGq5yObBQ5n20q0hSpErrdFVk9rLklF14zGYOQhmdZVU/hWbLclNBJFQT+Gzs4j6J9CpRW6ss
x0UoDyYs0nxxhi+u6AldpEgYahkEoNzN/nxHRMU+wmaFK8hNjJ+ERWZ1z2EnPj8ThV5p8v0pu4Wp
apXRAkAqCdmBOeRdpknGOvuSKxzLS2hXG03PWi7YhsQ+gPWWN82PkvsHNuEoVhQLGLPgpJxMRJA1
vF+EiKGakoOngWlA6Cqjk4CgYpRrmFyF9qGg9BSYgqM1uMKu5fqNxOPo7YbUCNW5VxDJpHackEuE
W+zbRxNqPdEFjInKOMgfk+x9REWnOvS6k30A1lm5gapqQmVtUUle/s7qXMZ/BeYXXcjTkben8Ia6
eQOGmxviG5jDVEY8uTYtFa/+FuJilCWLVMk8HZWf3UZQww4YUQNMlXpdMtoOlXyzQcJ8rjFn6IAL
g5YQ2X9tMulV7BjK8L8kyvH2+NsLoOcAAsdcNY6ohjpJzkBX9QwE6fx1VCLIvBvWjAYc1erUYqhx
JdQWQHNj6QjVuphWuFSi866uRg47nYpAHv7sWkXb8prq/92dwIFENvrGzhrSqIE3C6FJMYXkbfah
hoTwuzYHdQ+ioHPTTFlF2ls7YwCeXHnsbPIhHicKNgxjB8FglxmCqAxxqCXdrAQOPRfDJjWdeiHY
KSqJpx4oA69G8Dd0LX3oxbv1WI0kjtXAp+3xatNwA+aOBV1caWF9UZR0s61eWoqq/sy4k7jbB4QG
RU9nccUKA7Y1c5PrJQ6NarkZwo5BYUDGxXmBe9Tx29c6vMcdCCrj6oromvxdqWJJgQGlWcTnwojx
mFDi8Amd3Gvj2iPr9meQGNL5QlZo9bkoFyzKe5Egv49Umil4cacLgjJ4iDg8WmWMN3/fjdXaxq2D
fuBH8aTe1SCYQrtFwwDmzhkNiCgNB6CBmTUd0rG/nIRL8fvg2EupGyUHhs4B+zH+giMH4FjZjSqO
E4jvn5/AUwrZfJ6k/Ypi3xHL+py6C3K3wc8kLklROoQXgjmxs0B0nBYa+8G4YDNrpD68KXiTTDPA
g77cpTtnA6p3JNiAWkLJe2d1iG+jwPvZmGlNzA9/cADrB0Nx8B0G60Ff/tVlZ5PABYT/mxApOAcf
SaEA4YBnshPTRrHok9aXzZ6Lz/I76iU7rrXanQyQOJc7WoJQegcQ86gWTh4MUp5T8/ity5qWSiEx
CRPNdXKoC5hlFna2E1kjd/j9NkdVYI4Y7fQSeRl7fRStjHrCAwbFOgtxCLA/DqqRYxqZCtN/ughW
HXF6sn3b3R9l0qroggb681YLDgohv3KPwxDTYDQnFWX9sibVm0Yzo3UtwzVgQ47AHQg3KmgFWxYM
6H2KkMhFEo2/TScKZpiVO75MohbIQOh1X4UIYkDIgl9O2gvL6AdBltAtepcuoF2JZMv6lzB4LVYx
9dzXcn0/KsVWvsrrrDtgFOaHY3bqvU7YgJEoWsi8m+AEIHNc3TggNSVc8k6L4X9Kft5w8iIoUXxu
//hSKcp7L5K4FHnox8kVWfcNzUP9OduzNHQBAQlM5Q1neq1gLCKDmZjCFw+6QBNpZG/w7fKsnzf0
f28O1TdEoU8Oj5ECK8Qvy21gz53M80hC5hKHf1zoo9K3oLu9PehN8WkO6WFwhqfb+HLc+Un8nN47
oDd5zfEAIkH16aU5mgPgc5nRro91IFkq4phTXaruAriicFoFPI8sUjfMcGcqVwUkT3xQzPwxrApV
CRnNozLxG/ROcTYWv3JcCGvFoJCtoJ4mmvBsFSlJdas9kvBhA4kL/NmRk6B0Ebunf4RCjfhaShG/
A0InmWrpMnw1sFB2w7ITmgfzNvzNUA6GIfk0X6iB3COCwG/EowYqWz7SrGA0Nn5JsR1y94axm4W8
Ms3e0ULgROiWMgJ3/0Z8Dangiro9qqH+bCdjNHFxNfHtXbhdMotUKfQOIFYF65y/YrqTUy2oGAbt
DT6iERB48NfevpLXjzm9gXKeBXD/ggCxDLh8Zkkyc4NDMwWepQUE17R4NhALJHuavHu9LgYmaetr
GH7JX4DVJPAR4bKtfmdiIkMPjuLCj+0XjXM52YnoOY5NtfD0YxAJknpopDQ1YuYuSser2TPPE5cC
sV89zepuNbehyszjLyyd6Mth51T0k06otNCv9xUCl0KguLssAM+sFsqHE0Q22FpJlY6cOrZvTuM+
h0/a9D3R8qAcbINfCdw3t83fDXCuhTqn+qHBzhitmsSdHLilDQwPUV6ur5lkgcm91pqmN0CuGsJQ
LyhjmT0ljRm1V5QhRXBDWgxqSbB4WhyAEF0R/L6vW8GEuyOtG7XdbAelSKQcv4vkN0IcZxIozSqv
VQTWg+QJYBj2m26ouYN48L8ruVu8tyncnXiQkZHTBioTosYA9Uzo3yyOPDoq4/A9MEnMMzZygQ5O
8gnsxaKCAnFBSqBwO0rb32r50SqEWhu1u/ODx9XCr5sWv9VIdeg+mbdF0gJHga/WFRwVn5mT0oYO
VhRMIhCztETln1AGp+J22S61QPtQ70eX1BWNHgMo927Kw2XT4gYiLxnLxaOR3PStyW+nGnQZHmB5
57QlzyUxG1H01mYyzx5+Dg6uvOzxnxuRL6kllsdv6L+b5Vjy8QT3QDz6YYbkTjohxxYRVKDqWGgY
tgoULHnUXPP9UNieFM65ouJe1r7LNBOXZQsQWZI4HV51vlatbJ5L5aikFg/d107rau+x9kPxJqSq
edy7l63i7vJ18ZEiV+XMy1eimXzGJYvM2Hb2fFG7TjbpW2MNyCkD3mCexIGBhps/U6jeoFGEVqjr
o0Xm+eSj7YTfpB5KhiskL75mDbh+Vd0t8MnTnkr97UBBrVmEj232jfJh3i0mNr7t9aYX46Tf/h0s
G0T/mDRk4jG3vBJp3HUP/lkt+gvgB5+zhcRZunr0o5IqyD65JdmRz0T9JGHbpm6DlY72EHXVmIVR
FPIwiBI9RDV58DVjNTWmAjgnxt54vTQVW4ui03h253JWlaT0UGHGVM/BygdGkN0pwudTyHcysrDy
yLe8hfHizf0VidzibwrA5puqKjTszCymmIP9HDlbca8sY3V5+LPFKUnsfA7AJbvSNKIjxLkk/FCT
Qfk6w1Y5673SNalGYrv2p1li4Qrl5Xlr1I46CO22hhZseDQQpUkmomKDGnZGBu3xlCvI3VGmDkxb
+nGa1+4tfErMQTzcZjeubtluHWW/Z5yqNhhs1MOS92Rdv6MFc276xbGrnZcNVaAy81aYLctHmiZu
IinSycH3aLu5NC34l0xgiAVn88Q2zVbSrce989U8IuimRC/+Z3xzdV+doWndtOEkpJSl2iQrz8wt
8/vJyNrSSCnOuTQpDZBXJ2fnXmI7cMoqdcO+yMyN8mhTA6Afgp9/OOtVszZHCGH31fwIgGQiAN2Y
tCH5HrBKx+qGFpsT/Safpr2sd3EfoedGc82LKwsibuCHgS0Bw1+Pgg1kk9qq+qxreZo+fDVEVwaD
RpxZej4Y0gJiL8gQjN6J49NxlNEDtO4TkhW5QZdBMNAUPS13MFw2t0j1/EPZNQN1KcKdTAqVMwxK
sctCJIqMyj3KSXicGTQFBPvVGTL/mjwDNhxLwM0KqaMraR606aKDV+OYOJbKoHbyGSt/1U6oMPu0
wLe3aSYJrL8vZON8IbB+uv7LtMTYBtArWCkRZ5xgn+NqLgfXMtzteq/iuBeuVg+McfjFNFDvXH/p
eueNcuggL0oJfelXq9KdPyrrmnHajLhaYaVbLnqSMiFrn1Zb8/LhGuiO8xR9xfJ+D7y5KTG/Hnej
DeU2DKmY1HntUjDrHDEyu9BH2K5S96u6+ui6k6zvyhsNQKFSi8XAGquiT2nLBslG8MTSbZxPX2b2
q2LeH/tMGQiM8m0blIcKHjFEu7e/bQn4HH/jb93y9zRVt/I943wR338vLRXtHILuHBbETHnEI2sl
lXKLrDeEooKDcUXy9rc23YQs9umNCrmd1CgmAUEYWoiNI4a6N2Wr24c+qNrcvlDCuwpI+aWkMGfH
DMak1eVs/myBuGqfxh0kRUg0WS7atwBmYUAYUFrOfoeOdGFnFW4OuME06IJrv3doMyz4wft/negS
6oIdC60nh3oDFZVx7Z8gpYuUozG+k3iam1HC1lIYc79iNXikCUnFAcuKQIcjh/VytYPkTe2qbdnO
o6RqA5VMCZJ5YC+S0rBTCVymJO+TQMgRGzjnZwb0JWKx7FVWcJhCKAgyjjnGgMBZ7RKlm8LWw77s
oouECR2/xdMTU1WFqiFQ097eGUzM38OWrDNrzhwM2aFDKkbtyceJFSRmQtAzZANfZWMm0PVWs39X
Fr3EmiE0p2KIyD7SL52Ry3l5EUSqtOAfikWvlKC5iR0//moQvqFkhAPlkCms1ZpaAfulau++Tfu4
Q3JyHVlaPjATlk2IeGpvwwZ7o3JZpGIuy9nktPE9Qm79+8cbEKYlicZNCvKzgFR//dPmaQuCrKiG
AquIlY1BM/WPl5IoVPzI4Y5Auq3XMD48R9gNEaUEiBSGj6zxVYl/EkbN38A8+Y5pZV1zrL5Hp5cU
KYzfoWE7hOYz0ebVVz29n1EeIFAkJ397Ai8TPLl0umTvEGNi+tMtsgBYwNR7LcB0awvcMJqHkqyY
Oc9svznZAlDygpk7tgtxZLbOAQq+J4nePguJv25KQk0KD9X6WOb+U0vxjKODMXuwr81cxOFqJSdk
L3rGnIlBcZQpndEozmv0ZPY1SkA9JcxSIq/8frXx1pwwk9QGKNxsXR4FdBjsV5UhSxvaxfg3iRqm
uq7Ve/GOwkTqgXUn52NBM4kU5l/Q+luGi+/6TU4YBY2Y2RvWzCgKYBsURuifDm7PPqxfI5XCJHSV
DKa5mI465bGqmgL8T2aWHE/8kOiXLLAIrZ5HqUePb9AxTcKqN01jJHxPf81xBOwsoPu5YnE2/HFH
HMJWk1HFaToA6yn9fE714kSLNf4UELJNzklq5fvU6xVlgihrvBYICjYobyo6OWDBO/zY+35NgXt7
SGh680v+9rFMvIwM0lBouto4mgZH83C3gM/kRQl5kdtlynDosaiVt2SjNoaBl+qW6YDYI6F4gjCV
nLVKBy2Xzm837Mi5AS4CnRbhja30M62vRo3Nefn8ekqfHVms3wIG40XQAKq9nDa3bvXYQ3qLT7x+
af8aqNoYRgoqwnPHZuwG1M1cQK0q+ilGonnmvK2UbClHuO947Td8rUicG5snCNYTQGVHOVl81/Xl
H/fGm98iYgDXQRWMy5u6j73PuFvLiX+xD4ZPY4+gudHL2TBjKO0SutPjCAxGdo8XM8LTxl5Y3BRn
Yw9I/NlL4FChHgB0zBgddTaVfT4skOlxAekD9XYG3ljakqoyEbGxp19+bEh3tcWmNm4IFvk/OkC0
zPb6dXZheqPQgUXdSO2UldkLFzmr7F/VbyWdWPE0umvLRca3Y0Y072LON/yCJq2xGPsanRXODFHR
f8OBzR0Ycdr81nsHAmXvgSTkLl/rPCtG99Z0/DvqTVkZfZI314rL6MZYyoxu3DXfIWClqiU/zdd8
yagGCXh1sqaLeCTcNIzqTI3ZA00VCTwgjyByvtniqXX6XLqAQhSwJ0UW+ztFCUgzP9xkvpK3/Whh
afDf72HvwYozvFfWmRPrGDo3knekVaI6K06ENarS13RGTaXSqIJdmufrCrlBU8biwyPlZ0ygLm1S
AJgeJLUPEEgSHJtow2DmCNVXkX7Yc0dCe+1VeKxbdtfLt2S+1ULDaylwMCWsCycWHPtyPKzPr6rY
Oz/WcnC28/Xoga2ODicNLpp5Z/AarPI5uokGiQMI5ZE3zAc0qf3BG/kuQfCNw6fH21OSHbfbO/CX
4jl+6SbUQkzB3NnG+b2zPyX3eFuE4qr0hegoGcR956bPuFgzptZzl+7LCG1CsGeTDAYyc9iUr5Wa
66CS4kMcwGIENrhqsFlNLBX6/RjiK5UwYmkBjwAamJYVrjD4DJS4k2Tw6fVPAAHLeMRyQq5c15Ym
HIFtdRMuwDLH3PVC7wYgQo6FlcO6KLIJ3BZN9r7BfOtHpHmDSJf1HUXpcaJUnSK/hbSxm2kvyiog
S5kM8lz+uDtOsnhZu733BYKWrbsDU0co3KVOhVB04KHX1422vQdAH9AFJE1kCizbf2TJUYsIWt7U
4JZxsFIwA/q88IxAXPx5E+3bQ3Eu5B1DvYT+ajjNLVPW+n4AKPI5whqbo3nmwyBL97CvPnjjovz4
1YyhsHhXNWNPd0hXsrXnLWNnLRs4scrd/ub+pbcE3MUtSNMszRoQsP6HgKbJgtQcYcMwX0t4BvRx
4m0wsvHcC716fQY5lqwoUzyDPPEatDwradOQkZRbKVk890N/dtC+JPLfE8tk8xrdEzwy0+WC4C94
6D5GHf5o1sbvMpvfwCBhG2X0bHZnVElqs+BpqPZE0QmkdY2hYFogUUxkzb2IHo/vo9nA8l+UaorQ
tX/AbYSUiqbcOtrkZ3R4KX4tVVfzkZFdMdPZCmL1kXQAvAm67bc1ZYAuMprziAiFI37HFBRYnBFe
wtAAoLwhfiW/6PTaBl8I8zJ34dU5d1jrFgvBaqdzSU5HQDK1PwIVlrbO4lqCo3FhdHFlXt9k4qdu
Ch9RYV3vIOK/zcFStvN6YU8PaWYt3HWYd6jcPio8EzFORM/3QY/Ton5hnM5dKkDS8VGbCGYygPbE
18KhQA8fLovPlj7pPe4IM6ABImJ6tGhAYl8ZMzEIsx1v0Thk57XBcq6hdfPVuZnY0S7wAgSyPrAg
TxWXlRCLuYyAfvGIJ+xmXDMKKltrBZzOOkZFHaxXTITEB9ZI2CINQ7Rxv5F5y8kNVgeaLw1ACEOf
+C9zZxhYy8HUl1ah5ZevCkn/NE+44LxlIjL2BISKcW0nV/Ury4/62M8ndonau2Q5XATO5e6+pkZZ
Mo9+bo3c6D74FUNinFR8XMFVT9I+uHSWDt4vgjTD30QF88BgNLEhvyNSbS9isOyDWMoq10xKWhJV
9hHKyRi5mcFwvasLF+AwhMTaPs0RGtFEk73scHl6D3dNQWjVYlCUhtE4iYdWvDHeX9X1++I7oGqM
r4J2Fu7ONwQraKrwrHcT8f0lR3lWb0Ppht5+pSIGeTnh2Bknb87fCZ9lWofFW7pJ8NREVaLXbKVA
OW7yeqxvPPaPJPbzTEoqev6UXpsNS1aIjBN96MIdyD6kAq5OCca2J5XaIKzFi5139bHXZhTF4XnI
jWmvGYxAIFtIr+i4aaXdPg7iL5GJj7ysXrQZMv3FKR65uayskdCQTK38dL2YbFBSi4q0MPbZefiB
pVElyqM6o8TWQVxahMR4tMfH10XSQ8idMB2LuSf3leYrEZhO+sDcSFrJPnzkvsdMVH3F55ELqv2/
ybdq6ivfri5ZHiL43qjOrWYfImleuQu6o6s/yhzFPuXd4JUNBmoJuv/HyFiTT0l5QYtawRwNpkFF
y2OUVBtBqgtjVh3q7r82ZDzf4MWzSzhdnBSPherqfRFGXG7Z9lVrKar8HIdp8uJLvCqAEO2a8Xl9
zU3z1Khk4XpGsu49tsq1c5WPZRu4dXT/gZ5fEu27N+iAGPFBehtJCxAa6yIDTQFjhl2KWzhpuB3d
2Bd8yVCXtcEIXpPPBnVZwESU7ACb2jrl271DWk6twvzqN0hy4sT2PCruFfZFGEy7s0TGSGDqsPx3
esoWvc97AlG1UbTtbcuRwQjWDqn0PAxcbJJBX9NMT+qSjeqUewaYPEeRrI8QYivE45UZBx4hm4nS
Q7TEi413V1mrYPpF4JffF3kTyJ+AiOezH5Vfhv0VH+p/SH4Lp6koqvClRRpkqea3TY2icCKN9ovo
DuuoTxotbVM2qHbEGCeJFQtDhzvIJMkehmZd5urlouBzsCVlH6mQpWxtmCtk6NaduuQhq/7ZZHJd
P3AnjiIpbQzzvQEbxGa7+ty9V9tRgz69tDJ8LPRe0guWXKf49ZSvkvNpnBkTgd05EomJVB1jj+P6
6RJQCF6bQFXnICNy6pUMYBGO+71e9M50ApHfjydtGWJkG7fqpYFny7v2Xj4t8IMC0b9VBnELDj5H
qrqPbguAKOYd4DdQjCQAkzGxDg60IyL86X1EPIHAQnHg1swVE2IGHCYNwQgATvA/BdDcPK1BIhcz
PrkqHlTKXATHuVne6sRyCy5LkAAvgAwhPLfpV7eg+GhcmcQIKdKpReN9vozSFX0lGS8uA9Zcwa8H
Ernd7IzUk/+nDF7cffTmwLIzM5QrW+HsYovsk8pgMFpa6cuJg1LjHUoCUNZoWXlc3lfVJi4CWXUz
LONnJS/6krcFCQAE8uvsqFzoX03XswS/Rzsgex/AMTYAaEalf3qlU443yw9hZMUJCewE3EzIbegz
smMNwZ1A6JRc4PQZJ3S8cRP2uOlIj8+PBkRmUTkxpRF1B8lU6yI+o7FHa2ACVYR9/13IEr4o3PRm
N/dCng6kHydy6mzSrS/7FhXDvP/cKneyMQBhQSgHdSQvYxzd90UZ0KzvwCPEbXOUf0CBjPqRtRCd
gtN6nw2SBpHu4CZcH+GQLxVIwh78dSuq2z89GITXLHI9D8fF4C8zOHvD3lAhItQBPa7TMkDunohQ
nOt7KRT3l6xsAxZUhMcxo/CLJ0zEctuale8ZiXAYdFhTmWT6MHAKPROMa3rkU4Bk994KwueGE0wp
ZvfFDJq8YhujDHXIqnYKaILxXxefsqb1VBn/w+edIR/Lav6mXtGcHEkrchtBqAvFE7CihNM9dfAj
22SSxsavlwzM6jWrgZQMf+NIFm9mmnH5FBfMIV2CXx/R5ig/9VHBLkCazyXQUhONQ5AkmnSkzZIe
djBgUBDsKxpz6NujK+gqrZcjtXgAKgOxRsJN5IHUxoQb28c6KC4i+gbZwaij1B/0bsO642r5UHtb
22xuO6AeTVLA7lAJqpHnHL2GQtv0dOJdVHA+t39pTRv85PINWFwqe7hszYjI7bxQhZZDs1po11pT
eE2Z6AGl8NEAE/zEz6By6+s4QQm4t/zTm3Q6C3IOU/gpVbXmBjMdoxk2asrlc1OB8XqoR5XxaftA
UaMCH4W5JLpnbiC743apwgqCYuedieCHXiBOu8R4gsEuv+jywpo3pjIjKLc4C7oAf3+KEa4PtVkj
/XbbzLsHxMqtwj6RaDwZ9M09tl8faL79/X5rbNjWo1yJDkDtehFUkYNaHGqhBBLR+ZotOOuk7kxM
ljjMr0Wrp3jk0aZPoM3S8OHAXrpiJezCq1svlDuDF1cbCWVtrxCC9DPOj+ConodBhVKu9k31OlXY
kzd2+LhsmqIIV7WI+UAlNs/sDOhRsZZ6Gb3M3ZsiyOmbzvbpbspoKvPyFgCX4x7WLQa9obsy3jYq
wbT2ElMLHToff3foRkTUnnMhjbJcHQ19jZypgdRDkp+4wvInWgT9gSks1GRBPXGrCuAdxW9oOrZ3
8rBB31f3zSCFMTsLKNVMsMdWFd7WABE/uIQMwa8WWD98iy4GvotT07zIheLY7IXTUXUxlxuTdepO
TPHX4LATghbqhUJ72HyRDCqI4JAeS+GG+c16PSsu5kMKbTPUp9p2RkUum7HCLwIWCAxoD+o4jq+o
yyUdn88Hgr6X3QrPzXA8Ie6XQK5zTq8mxHRHy3TW3BjFpqSRdPY6vyGa5iGhRQ9EYkWTuY83pp1N
oi7JPMNUp2OTdyC/Nq+wqe24o7A4+7BO3DN2oob4y1GYL34s17n9lqx1N4PTF9rS6kXeQfG/GmdM
qvSrJZF7+loDtkVQM95ap9zb85hbjV4KYwU4tpnUPQBZhVexQGCKw05UD4foUnl36yAY/dP41LI/
N5dIb63f7cIZhCZOLnrSi2lFJ+Aqzea6JX2pMK5DRXKXulv69SJ5gUltOTT0u+2J1j/QKcpmECv2
b2S3Pb+n8eCNxXf4JfjK4o6Q21tdHT62goySHGdTiBzzZ6fKCFsASGrqc1Vx9UWwUy2cDXukCflQ
yr3nGC+zSYaCUDdMizrwCsn9aLuHUNnYQlqAohVcBVtqc41WNbnnHcJGCA88vA2c7sYCoZGnVFdl
u8BJ6Mnooqd0UzKiZ6S/7LKH3oJSO/iZi6QwbitO+5VsNJaJV33E9OhRm2x/Z6iPhmuar5dHAlSd
8fJOYEoDjIwAmT8TbVxjohHB4408cGycyRnRqn/hjTgC7WyW2NhpmdrQYUHAD/FiksLDFgHDHM/w
pUsrfJZcJ0T3hLKKYLFfjhytMOC3lVjzqfP6UYpU6e5MrZZig1xrsRv+wuLOsoadIZdA+8Kz6F7V
gwVZjWwaCZYKYVfXPhPjYGWdfRU7VrYRxSoqdF4v7gkYbV4A4G4vwYW6G0huLeb/9wP77YkTmp3u
yXUZKj923Z+cGQBqvttaRTrMMqXiUHcTHHlqEZVPZotBs+oh7LeV6NSUfC7hkFzTr3DvrTjvruT0
QXZtnh4t8c+lrT9FBzLJ2t+nsSYoTHctVPftWzlqvJlxdp5EUr8qfGLkIx11Yk7hwqKY2KGq5GYD
0EUP+lG6FV6Ywx43OU+68OM8baUwcCgjlNFEOsvOkF4uw9bik26Y3fThaNchTQ0faESD+VqSq0s7
x3rNX7oL+XqeOH2+qGiTXlNr+nxO3P3uXqfMcgSn5mdeFB8/kvMDeKVUDz6rr36D1yfLL0BgrWEn
MGkrYU2Q3cU7etrRn8SpyfIwCKBwX1LiJ/6AFAIRJ2CYyx68ytx2UBwGdzN+6cT5teaHWSBommMB
SI27YOCGrlIdIzr++AhhIjNIkbgrKqIhVL+Ot79YoW2voAl8NBRRp9Pk4Sn3baUFnN/t6aG7DmUx
PjHl0/TVx1Ti0kDmxgwWpXDQiN/cIpY7231INcG8LTaMGtlDnXl2HRiPEMZo2nvYx/hJqmFawcjz
ChBwLiiaXkdW0vfTqfJBDAvuwYaXPhn6uzXBznc9yxx1EFsttz/QybngembhV1hfHiVKcSYBnkaX
LbQpQr+ExPKyh5xby609nuOgBGkl6rri0Jx+PplUETI+o4MqV0WDG5aKjqxoBBpR2Wm6xU+r/cOg
aMobC+NZs9tHt4xeXK5aGyFtjZ2IalnjoOlQNMuZHybXa/B60kZ3h4mxCNYAbZF03j7p8rYLGJKI
BawE6EhS3hJD29jIuLtvQ+mvIk4D4RKyfK4btQsYeqJY7//MdV0YTlgYaRkU/2MDG5dafWtOWGFJ
BXoi15kW4BuewQ4lzUAqFUGku+LFgMXSa4Srvdwt91+6cG+OQsVkq/CSGAUOFyu4YopucQEd4Mdz
rb4LrQhDi6hER5tEDamMX3HDAEpA0XTEcaP5LFfdTpfTVeSmB+Sw+C+mXFZpneZwGFA2tdwLj6gh
wAU618hbLCuffrNcIpOCj0O7qMbj6I6dH+RrtpYe1CJQdM1SP6uUXeMymfvVxjeFBYsLMJ5P0R5v
3+z0l1+i4u/6gKKlvSkvf5eZ0HmB/X4POZxbUFR0XYm02x86jI3NccwQNNHrtUlUwujBi8ltMJK4
OfEzvYGvlvJxHh3M5WZUpQxmmkPM2jD/mfS5red4IZ1qsunVe2HKB/cXP1Nr9kHBdWFreE3mz4od
idgSffDmBjqu23coAVT43ufTG7qz5SwWD0NcDI0ZB/xAGODX9APZyfkTPa6SKyuNzBS9fYh1Q4jx
4UqoMtdoQyMFUn8Ay39BDS2Yj3O0c4bPN415tYOTGRnWIPyKATeT1g1XRe8yxb5yVSLrQKZlnPOi
jLfmnGD9lp9YNraPbZA17aMODGVXe45NtpSjnFFwJqPgGIg4bGOznj39TNvZXcasOcnVYbo46mM3
0QndNqSHMa1Y+Y908XurjlXsVa/lD7YtwgHCqMhUDhaTYLN4a0Wxxoj51dN08Qrxqmv3PyGafkek
BkhTtYQppmNRvJaR/CFPteztqc5NatRmAd4LpcXpPTnanNh14ytn7YdUFUhY0w9EyGsdIZSI19Ne
cQiWUBVumbFfdVupyq1EJsJbyNW6dy08iTF6vZq0lUhU4zhb2NK/EKyqKCTY+Nd0Le9yPWplqiK8
eItZzhXngCLZhoKdrGH0mRuxmd4yOB/ul1RUvbhNC+QLdlbf7QVzgCtk5ujpF/T6FpzNi35A1git
gstFD7LGNpqp3ueVSk4TmQH0Qng3Ag6K17UCk9j6iV77rFjHIktyJ6T3CSTMshpzqlvSIevybFBm
ih2FJ1RGlqsLI0EHoytzHgzVuYIcckFVv50yBEDKzcjV3I9cJ92xqkMfX718CDJGc2Gko+AooJ1M
ppclMlDBAVe9QCy75MeXAYiH4AoO242NVoQXQ6BJk5lWqnkcGm/7MBHi11veSYFRGlfWCSd40+0m
BF53IVHXHcS5EGJvW5TK+GdTA+Q6hL7mwsoQVbsshCJLiiqWXRgjms6dRm7uuX8wbXCeYdkpNQqd
WiiPLY9nICbOTSlrgtP2QJFf3W++59sarnNvkFhm0hrs06RXSYu4sj0qJEWNowgRyn/piRMu05yV
P0xW4KE379L2L/kG2m2Zx6bBDzmFBmKA1jx7on0QUSV0+kmpB8g9h8JXni50izdN78E+LzBtBThF
6zZOtom39M3ZrWGv5gysxzg8QVijeo7364hHE8MSvJMLArfwmdOACbSNLcLf4RKNXigVWPWB9ZoF
PPqyxb+s2WvhhDBCzwhgP4cPNx6JW82SmEruDjsrSDH0cbaLu5t3c2gAjYYM2g8wUzzIXcbwIMs8
gxRD65iy6xlcVavcaeCuR67o7njeXdPA23LjzdjqdU2SjCfi8CSpWy3xqY1ge/TjtqhN3hIDqDHT
uvHGS0009SLNPGrAA66selbmoTgh7s/K4FKnlW4xVByzoj5cqg+0KlogN6JmQr2gEDkh8ty9/+JJ
uoXdGtMB/3Ug12coUA3jOVhVWHKRx9ubIjXcHtpNIsgX2mBD81MzwwFt+c0i+bN2OenLMTeoytWW
W3HlOb5RXeo+1IimBkzhnfTdrBLXri5aiHT3BJguT3H6D12ucGT3lmf22x3q9hxSVgrdSi+2jsJY
OF+Akt4raNM3DxkRAOatfeEKAe2y+0wQp7MOTVRunVI1KRHNY+KT5GTaoGgl8WlBaqkpU1zxdE6t
rGzMamdgqkDK5QWFuH8B1838rGXelwM9KoMoxpNaDC4zdQ15vA8Vbn/1rHAv75Wwjz058CRkhBpT
AAigXbiPEN4ZNocDNnAWdpFYVLrHk3wmngiK+XZ2RjFFbFcr8CcCsogrftCVD2Ivc4sIJk7aYXEz
Yw+5TxSNtyGHQzMRrxD108ZqPQRiripbG80ygwIuCOHeDvHxOfnVxMegp2p9XCOZJk5YSj8/xK8o
o1ycu/xaVR2LN/KK0JB02HFUWPvUMS8R9Segtt5SCqVLBwd9TdngQ1OMS7D1nRx6+n9SeVmVA9tY
rksfr5h8W6DwFYuXW1K0O8N/et2bIvo+LphWmlt7ZaCVmQhsqv2VI8C/q53t/tAyPU3uXG+E/jis
QyfokVVsykoRZ24JvkzwQ3m9ap4KZNWGe/O66g8WmY4VCgGA8sNNE1IiHsI1noUWPwagF1D/SZP9
RUJ/iM9FemUNdcYnGHzeKgCmaGJbmG4CcwpGYYn2SLIYmLa480vzn9owvLueJwHs33GmvPxIvhs7
40ILbhMUjjnBQDBWvH8xJUWXIf8zJp/V2z+gzSK0U++bQGgtVtdJGxxlj2sGfw9GRCI+FpV71HQO
ZKdtpOkEgIZUtZae6aZtRJNngW6FNAZoZAHEIiDv5fQwOF2joSWhwJ0qGyx11o7+DRYrIxZcfRXw
N8FbkGWZ9Gnom8Oz9p/MDEtQvjAj3q0Pv1szBenXqc3MgLJWGh3mp9i5FAAGQN2+aQ4RMH4yIpiS
bJEy/hV92XZNovT1lLWpajKiuMALSARQjIaUkWAwPpzGbvqM9TYurq0uASwf32VPBhqyOGyXsPlN
VKNFl3Ix9nJDBevodf7Z0a5kOGg82/ZBe/5UdhejPXQIxUTwURYgA847p52HNyyVntz7l6p8WsDI
MceZm/D5ZI24ARTyUMAO75xgJFsfeXHjO7TMVLTtLQUd0FYOzgbIkZP6I3FqPkSmx7RlK9H+fJ7o
wKnY0CBMRM2xdudoAagRgxOvbWppwkVLZp+RignwPtSAv8rcK+ZBVyn84d1EziMOVo2AGsAMgqap
OHXHWEiQ0hBBxksmQDbOe6mW1sBHA/XK5Edmf+Trk0symodceeO4pzYzP/hv2qJWO/bnQpha8EXJ
EVMSVUWP1Cjaorv+F5mwDGvr69FrmhJX2TvzH/HXuvIliQ6rjAJmo0Zb4Yrt/lesHViVwTHzmZCj
aazv0bKqySpFxANcSlO6xk+xMvdfMZ3CU3hij490HfNzsdjZHE/J0eeBxNTzKDbvBEB2LQ8WrINj
yOQrf+y474dqSrSPohlmjdSeKa7sVk+p+I4XSlPoJGlA1bP9Ff4uRd7WuKaKyoxD/XaiIlojrRCE
JT7nP4C1c1UpTCVWX6JZb4gGk3aMkXHoH5lZQ8QwtQs5IfCugTTJ6XPn/9LgH/U68h+K4hggxrMu
u/AZ5x224nayjc++hxP5uuFqAcs9Sl2s0Zk+hU/sCI7h3w5gh5tHMUzEpWWynco7KetcGKTiEmuY
xEsPtDY/hcXB5VvyHpg2Zc/UiRwb0LsKWPiLQ87fV/D6AoR+dffLECz0mVYRifXJMv3V5bLM/nxZ
bt4MYMcndoQ2z/VcEdtgK8O4krfqoNF82aQyeVZtC7DZDNqkxoc4hxuWDvl3Zjcc1kRTcv+ofZ4L
jkv6imM5J1ZwihY2wUmPVAnZIdqIDQ2uZpPcdZJ5Fh5OapcCSc1rQarW9ymVm0bf/CzpuV+LEGx0
I9C9LXsiTpFqtSnU682EgkJEl/Il0BVrIUHYsIAMO013rZo3aOFCm9ktfevuJ7szqTckmoksJk+V
ycjFfj8Jx3cy6Q6y/POaeCmt9fwKxux+r3k8jp1hLRAVnD8FFhJYLgyeg/CfJwpJoVWVxH+Cimrl
725m10kEHDjvDz0gyirhbjKm7bF/T41GJEv5bpAlOn+zlfJoCg2JhHibsKHGgBSmvZr7MIIbTgjz
XFg6mJS1z26VT+z627W/lrCA6h0Kni4QnWnSEatbcDSkanwSUqH+fuIpiqa8fBr9A1T8TTplEFwX
bqatSdfUwS7VUrZsiVs/21mkiyBA77tHLCMuo03esxXHRuY2SgUCT00scB7QRlTBLln2f17LFvZW
Bv9djrHoA1gqynsY3tJnC322egw9Gvk3w9fKW5t6cYzrxdEZ4Gxh70gr7yZro9eKvYaTxO0ZJDhB
mnnRRKk3wv/EH8cA+A5ky43oaWRdrDW5TJ/Gi80Xenq3UoqMb0FtFgZCKvNCb+7tMSm2qChr8qBQ
GXvl7jvcSQc7/dj/6HKqROsHeYeqNqeWHJ9hYsrKsHL45K9t9rZ+EUxoNvAtarYdypG5rN0KitPN
RPr1BU7ZOahX+CcyIxl9wamIbP9u3hQIg8z1QzY3wIu9XVUJyDsgQcDoqYcwyvZjSunxX9SYK56t
Adk5vYSp2AWucHj6Rol+Y/uNrhNat10qvzHf++YeWiECG38OXQYgcAQOWIR1/IuBFO2OM5d8wK+3
JHvUtCZWKCIErBt69dAf2uoeksPGUGLu4tp2uYtwcZR0mKn+G7jAC0b/ZJzKCphcCksDa7+uU+f2
VllXDsDZXIHkI3Ao78h2u2EZdHkh11AB3TOZ6JWY4a9ZBpXgICI/zM3xK9nIffUQAdaYLTM3RBTW
83h1TP4hZhllrniJx8XAjWzWpRd3bq6mEre7/3kBC3tZONRb/R7WWKJ9UevrTlAoXTNiI3Z3iB8V
g18611ipNAiCO0HKSDDYndD+4Eca5ORdH3mhiu7T/EeGd56YPNwLgIIhGR+uSl0vlpKi97OiIO+n
drxcukEBFUy3ipgpzzF951F01VJ1t8XMw2+j7gDIQq0GQAne2P5XHVi1ruykCcdU1PDLcQrI5NZD
XGRKMgyhJEX4KW/ZbL9emGW+qulR5Wxsdd9nK+gCiXfG9MgLEnJAw06GDl9O2sahPTqv4LtBshw1
YA9Aw7ujJbMuIwKtv2TrOOmcX8MYt2oJKhCBqJdRdKoXGVvn0RoIcf2BbZor7h25y/MRxdwqAREn
XvxvU04gQJkoqFc8iWtQUqXOK3ZQqsgKwXJ+QtXQ+UiNQEOOvQFUTPynkO+ECiqik7CJew+mRDFN
QtC9qWwVF1qdsMxFIIbwo7VxO2/O7quvhVxFBJ87j6PhqSW+SB91uly3VjevxuOSKfoTBT4uMgU5
BoVjnPP2jRmDgRVvGtR5lIuTj8U4q6f+HCU5iOy42AxvlwlPRRRo13tnSR7/3B+MeVP8Ehh0ybkr
nxW/wk507xoJ4sXnWa4D7v1rLSEH1VGeI1unoBcPv5eZtaDNQGRxe8fF6RracDFKYtJGTFnhvDH7
tGfd8al3m8uplztIFe1Gp+gzhxY1Z8MwwuI3hqt+yXOxx4oMUpJhgfbeqaLNj8GS5J6n3iMl2Mtb
ft76741yPeC8erLDKIB5mfqiDOk+JImT+2U/CGjYqrNpd02lHtmLR8rBgJl825flvwLuVePtONQT
Z7uuOAUegB/Ba5G+lEoAr+cEGy5K4JxnzeSISCMYWHRg2RKO/mPHhoEHPQrm9Znt3EvMTIxvEt5E
G4BV+2Xktb5hCsHDs0Uh+NACkzwj/iOIvY4RoqrtP0czhLpldm8aIrjVG7DuYT1yFXCpyN7dQFhK
FKOcCJkWpIUc6UDKWnSaP2r2mTBPZTBaLOdYL3IdmxIL9EW5N0krvSd96ySHuHzICtFvzPM9pDxw
xqCsQSpQ/5FBf21OcF9Ie9xURslQryXiApjC2JHdcrhkDeb/ck8oX9f/oCTq+hhzIHVQ3AOuOvTU
nv/4vvdj+RiXRVseCzmrkmOU4VBAa9ILmw12P3th4hCU6DYfgMKkjFKJsTkAUGJLmyqV9Tq+PZv6
ze+UpCdUWwZGiXbfyjI1ZheQN3n6P7/DrZs3DC/0DXGCAWVK+057Df5br/8qczhxpdX1dn+OXNNf
/Q+w9RsCSdjBuRvgyXaptmnHv/LWf0v0j9xWMSiDWwm6CcSTWKFKLXjW9O3NHFapn4Jd2AA4gzx0
L8zKZ/4Y7XBK5Y9bWP3OQv6c/jTkg1Q3nlLvuSsfSbm6pS5okOx/VOFV1T+X78lN2eAZ72WgHFTn
5mV/AZdlDalXJpkUlEKoBlzihagTOnOTV8F1yILxju+6gcdPdQ2MgKezPxmUL107Nwew+1V5MS34
d2hSOXy84R+Hf9bVSRmbVXVBFfD7Ue97eflnuHRL4IspCZYYZGqrk1EEgOJWkJT3UUtad7P+iPcG
BAlHj4+lHTX9/o6gHtVC5TlKWH1Nm5Mcl0Ui886Ipcb2wwwKga/6XcKvvtg6rJqsgYiy+fyTK/Hn
SskFeFFJuUyBnYS40RxNPow2ppPuSxMzqOYRUmblkeBefH9taNDZn/j7JQ1/Chuqy5u6S4WrGNI/
7KJ6LfEPFX9XgFXxmbQvFGQHR9B8S1RIxvMbdpMef7cSi95yH/zlkbY+VFrDuZNjNY1sKUaIyIZL
0xcME8AW+wTT9TCfarmuvnz5USon+3xg2xPk2T3G14ZjjwW795Ffa/CAi9wtMTg7dfkpo1yTPtD7
J6rCakGeRNwt70TsqD9WIaBOoj5qSOWo4Eojn1qk0QhfLQxq8InvkiLjipXiqtQyVw8ozAess4/X
Zafkl904BffnZZLXzILbzbxj5otoostIgL1MEGiYGh+YBkIPXjMKxxNaQ9RpgNeeGjkObvfzu8ob
8bsuILYAmrFXcnMHxjoMSjeExn8ODZNNZpBU2NY0v3LSeRJ4A5jfGMi5XSHD2/2eq1wy5p3yhbS4
tLMrBfk/08XchavyLoWkcinWn1KzmwtYbctR3XZKn6vdpXo9nXhStoMPkD9GISS24d72VebIyGPI
A5O3W123CZRp4eeqW7AI25SavO7o9nujtGTvUJnQstmpdV5n6W7iWLVAcBBx9kymH80hrrrNGzRQ
CslTw8JVuasSiKFmMUNzd6x9OzaQYfU3aqFD6tRwG7akhaHesgTJZmWGpMuszkESjKMJbBZOOts2
oH+xM4WYtku3xG2cnDgd7ZD8LHwas/So2nkDXFX8c1PKOn4ATOIx1eltjH3Pm0hvaQXMwF045AhR
uaxfCxfax5XzFsi9ztSICc/0mXdVNSw8NWJF/3TzEKEtHNLqSL8TWUOoCcMKJn4E3sj8btY1VmF+
3ERroF2OQsJxQ7SQn8QCdZ++fEiI40hbJsMGsD1COgd7Pjv9hG8MMKuwRRtqcPNtawpqdBWhF7OY
rWcQ3T4MOOhIa/3hKayHxGr8vvzL4wpxYbXkuAF6xUiz1eieMg75BUkr8PCDj0rBFfTO83QFjtPX
V3xmfmVfqHXdQWKlIKbvVSwrlZqDpf+Mcpe2DFL3fFdXu3MgjfD27rCZbITzpllQUjiyly5njqg7
8RrV9SBFQNM06wBQZvvbCZy0jm6ExE5RZvMdxpQjcz9233jsDVzR1iBfhqjoYlikC1vx7Lth+BYo
So7r7VMZ8EiwtkTGk8mSIhvyW6P9eI4CxVwTrhOJN9h3sWo7M5MEkG/7v52TtcowJ58W9fieN6Rv
hJ5LGQ9AgtKuDal54cLgVCA7pSLeHMY87abMLlM8r6G2zPBE1yCXxTzsMzrr3I95C2hfQ8OQ8Jjb
5e11BktMi1AO8+IEl/slLbdin/Rxs1I2Yf7+B2r9RTglaaJWoi42+Q/PPMTTsWocaqtop43saIfY
8EBwnLtrlRS2nRUYxlK9AfX/pb96qmNFpA+ttJ6HWKlgfAi/lklUjuoutGogscfN6MOS7v8MDf0i
lj6D6+JEf9xKqZjCTEgEsBEns6nURF3w4lg08mUKMg8um4N2S6G3vEpapv5dobTrWHbmDYcjIyWe
2YpZNh6sHrtIHgLnRqibVZFR0UePlXcG5CmqoLva4+u7wMwqdVza9AkkRWJV4cAOX7Ixset/XzoZ
rOG1YMV0hsboC1zgGJDzQCjR42wZLnzOdrbwZFjqMUgfh4UqA57OTVG+JuDVGRGQG0juORKP8lh8
fX89Ylqs0V46Bb26M33FuMlXq817n+FFgFtob1uh/uCA8zZvQYZeQQLmNNf5ou4KaPXTOy6sLjQR
G4kA7wMaSWNTqB7TCaNgbFSe1Zy1l8Bifkc0kNVFSLd9igAhqnMupIaLYFZ2znnc0270oiWvGZbo
9C1EelcQQkTjOs1FyIAN2WzlNzIyNFYIuIq4Jj7++J5tCwG/Pig5hbY9lXnS/6Gs0IVYjF7EtQIA
xbXephmhuMeAW8QcSZbKbj5uMIa7fGa1r4Sa0dVWAN0sQrZoEdruv89wimNQkszbkbPZgOvobsLs
HkwvehHffFAPsS8FfCp+J7Wae/Rrs75yY3c3lIv83n+108Sru22pKddXD6X5e0WM6uVi/6CzCviG
7zY9D4sQ5F/RLl5Wj8FVNGz8T5lMrylnMHPq0pThEy3gi233hnwLdz5Bb6kOJexz5ceKxFuRTlCR
8KorfG/860uaTe0893riTLuwFB/P3hvv8PMHezpYGJzOyQ02FjsDJZ5suQQDDqIbNGgvFi1maQKs
uyKSG4CWy6CBCgwhk6Rl9BVMhEyFvkbLNQLUJR3ipKNpiQHev+HvqADZ2x/PZLuUluFNDYc8vkme
wiT5YRZTsZzVTOOpH+LpdXQ2Qi3TAsseimQnnS1mbILJY8/sm+hM2K09xWsNhPq8Zn/xkGNvyBl2
pqP5gRPENbKKn3vgHrA/yX2hYvMeshIX/adNZ/+5GSGXvE3UDQivDkon5GWRAS8Gd8zAzZkBuo+S
GG4E+IAZRoQn6tB11KEvK2R8pVFJ3fmJ6p9cDZhkdeRtzEgYAGE+7UnvLX28Ndn6ddCgvAzTrOTa
vqzlt7z6ysLpFR+2jjgVCqH6Rb0jsvh4UM8VnJ/QR8HeZFSicB9dHNb2fVsAnzMrVtGJ55HJs7ll
C9MjEdlFoekL+mEz8OFymla9k9HXRqAJQKDdoMOqs8Pk/dSfcdR52GhIwssUNBtGpNUibdptVeWT
OgyAP9IMQEL1AJexFB95RM2Fr8B/n4mXz/PlKe/1elk3yrak9M7/v/Mfhwm8KDMTqd6HzyhmkPaI
bOQUWIRI/gRZjCvjvbmEc++N5hHzidNFMRm3Cw+XUXl5CSuI9g+Gn6/d8BudPLilk8mgzucnMO9V
H00vP2AaNXgUndMFU04JkXW4BhjgUgxPnmKYrGgJ+nqvlSU+N8PMnY4I5QRnrEn/d18DPLwIcS0s
jQbEq6Dq8B8Ul2m9z/m3o1sPoDScOMePcwbcgmKVqOZB3N4FdseKp8xULRJgdwlM8s0iHRQomfpk
Cts1FkhPATuzvGOmSMragp8niuUA0WzGGHTUzSPBZedBJAFvF8Csg+sw14xqvBLBawwn2vMaGKE5
T+kvhoLlaqeZ6Svpox6zXXxRZVhZYlIGzpP0FeYX0ThIhNvCTDcak4DkmK/SdOXx+fMnFD8SIT9m
olu2r29kacKR5H4zDU4z8WH7vshgpqpsSMGknksbwv1PiZeUO9YYHoXzaSpZefgBLDeHxWk3+JoV
7vlYP5zZuB41ZMNvII4jAyyUEUD7jLO9804tU9xt7xKX83TQPtj8bVTQbXuxScnV445KhBigCMI3
qXPTuIhsjKdZ+mFga3lRKy3MXd3XreZReizlHoviTDb71PWUZRQ2KZEeVfgRU+8hPQ0Eh319anJs
yARfyO3EtaMgNDOpwFYtTd87mU1OZwlWjcU2VY8yKpRIsXsSg2E3DjZSavGWk/M7U8jDV8jm2NwH
xYm8jqxoa81fe1wz6l3TjdWnXMB1auwpw1spGXM2NjiKFqSDCmnOzjdPBd/fVoN4N2zMTXvjuWu0
m9ui2t2yHpew8BYhtAmgI+0iCOrTPCe3lAriT0s/U7kmq6Kgoqbjh6GCsyWxsZQvKZXNJxCAVoLG
tASFh1pMShvMZuJrU9CjWzBPR2Csq/H8PjiQDmWTAmoEj/pz4ypEf7ytwiMsODM3VmK2Nbq/FfzX
VWN6UipJCb4r1JWZLdMUOStA7kjo/QhAtrNYORQKMkwdLO5hzkB+xcf7t9L2kD1tX9XceAOGI+80
F85EWc8XeeeE+liTsYblrPEauMuD9yEpn83CkRHiWBL4OcBlmmKMpEYi+U7A6YEDMuowFz5/Grwy
7cG4HWPGJXJcugtdsM2bCAH5VvztL5ytJjPgru05VGVmmWotYSevKtqEdWHSoUEGrG2qA36LMt/t
4HeTMZMBHfQFL1IhoQLNxyepLvGX3fDounP8c9OnWpWngVbcua+kS88VhBBxEVQMUHs9iBYIvoZA
fFsdCakxsSN7QtJCMkfhxy7jJa1IAvJLvu1PlN3EN5Eh3VSQ5mgAr7g0qEY8+wjR87vWDLYxzdh7
gE895Hd/7HiTkl3+nALx+ho5pQ/vQ/au3CmgWxuCbKZPGrmH5UoEf51K50ghFxyOMAbl5e7/Vfxu
JfkKxozCpJSHd8UowAtaKqDZ0ZR52hOc+jUK8LPzK5tkD49UozUvpyuXBUallOYz5nVK+n5jUQ48
8FdzR46agW8O7K4UEc86jms3ha45beEIHJdwpOSlmYdjnsTVFuWzyMnCmEzwpIa6102hpSL07NCC
F/O4ciXTRZftJCmtOCr2eK6lTtGyYGmke0QrpRYu95BdmBu5dtMqWCHzBvkSF/zzzez+pq1grG6p
50XJM1OMvLgjMr4Ah5sp3zoXERX/7sqA55l7t4A72j1LNwjMV4yoBVfM6KosQvF1rgh8PX7vH0dJ
Q+kd0pdxHTtLRRPqjL3VHJs7/H+2FSwxJDXaydX0Kh7pXqt6eSgs11qtyMHyqIyIWK4Uxz46hMfG
2MJhlx2ciGb4yqMU2qUXZWG9CUFfZfZd6ee/EjGc9AS5pIYGQPDM9cIdPtgrL7p/ZstpaG+A9yVg
Px3pqWBN3SxWTpnHsAo4fgdZjlBUbPgaiCNvfSNbeFBD6ddKXp1Ote+lHhawcyTnrndRM0wrfbyR
ylm+zvreUhvzzjFVMUnOwWA0G7k3mq2lZeoVVv6dhMMDLPf7ZadvzlM7+evydCD0E45YHEan+Ac+
G02S8poij/PjEUpLzIf3Y1aWCm5nc0ukHDwV8O+XJR2itu+MgvjixAAfF+EMwZ73IFakDPSbxcJ8
FiY2+WdQeOasKEn+e4toDzUB3PJUsX/7zqFRkWJk2jqP8ORHN5muaFXM6Jui/6x6xWruBmCROgT9
3AKXYbuPMds9RPNzRxiBedh/75ZkHF7KM940RD8voZV+HP1zUVqfKTIdkMFyAsMp1haYh1FGHW+P
etGpNGh+UO4OBk4O+6jeL6qjQrxrG7ySI9hZV/11NqWFZqaIl5TaEX2ueLHMFjnALTWiti3hHKkt
WI9sRBYfKIkLRwUX5vyTZzs0vD/Hx+JXbOR0WQ981uwZ3pkq+nEwzK7HPlccEdl/nkwtvY4UG9ga
HFynLfKPQu8pps2eWaviMWapfkn2aW8on+e/zxh3WorxnkgkdllmOfE/VuYJG1o2pzloNc5ySdOi
VsvKFvPy7ZDU0tiN2rADVXRhETs+NLQ5+HTVS+1TFs96c7SRVI5vtuGwdmPMlYl7Lv/u2ggU1IeB
MRO26FrsRq0pXeifiJOFu+29YMRufTLxzGix2BS6yC2gzMy8ekWhys9r6mL2rfqS4+wmbchIKpiJ
63z38KtRq9xSAutp0fumDsPNxV4wxvR7Nn0oNsP7glylLHXZl+TeAVDm23czpj0FlosVTuLU/q6Z
mmOSIDk7zSLbTBXtmyl4jROaprMv+at5PINiolrS1Vld4lzT8KjxHtCnFo+HsUBfBDmu6pwEUDLI
Ld9RKPfv32XiZY6Em+kMORJ55wk5YPJ+xsN2W8VXU3w3L0KbOXhZdS9FQX6lSr0401NRG+eMgRI1
Hd82aErXMOLlc6OMdQ72bKqbmLPIFaGsThrz1X1j/DvXc+CwKuFHXuOagVSxu/OKFWdJbc1hGG4g
C8RkRxgPs0tDERuoaM/2odo1zbs4yEtiT9xIWWLXI2qL1qhk5F1Hn/MsJ/Pl20HSr+YlBmVcmtn9
tsL4FHID1iK26DzMzBI2z5Vs15HFGvihFjNnVZO33Q7/1YtU7nVp7JzT6dC+hRVxGXaHx3v+a3AJ
4d4rQHena+qsaky9itYA6klHji//qeEgK3pZv4FCeJpG++ZKGj9rAYlW+odl3EBU5Hv4bSDCOpcQ
bWqa3aWD0+Jywah3H7sNcngTnEMSf7sIR2HfS6lKUHPx+kFAE5OiREOArjBMOlZe3SRty2rVECdy
M/Nl/j0WLCWc2hCSpg/AO/3kxoBmLADJOC7DbXHfVRclCMi2wXfCTy7DLYDKjveR51udS39/V1Kf
SqZQnoegsdUBeMI9yKPO7/jg6YjwmLwZ/GWLaHWYpogAJl0gkwBld7TWIMhUMMgFwXdrQNRQG8ew
iRVtSSPtDr1CV6ZJbWiYkDSuzPr3ua5rFHEkoyya69hL8TFaOibS3/5aeNfui925RHxZRH6Phxga
nqqX2YF3e1Im3j0jGt+zAdNEwhgIl6SoLtbGb4o9EQaIOJvRaO1HfbTwBh2yiDDFOcvKgouBWeAG
LnNwU639Ay+yVo5xfCzM72PUj0W4rBzVfmfw/TDrL8iR5hvwUBPjxgNV25yXFwS34mhAwWXS3tRN
Lb5vv0nmG7JEb3oVCZblZO76Kk91Mag7ICbLxMlASRUCLHZ2oJ2Dg8WkLfCIfHLlHfmd7yHqM3kV
IYZq18dj8Cviu/cWS3yth6j1fAfhxwehqM60yPxLVnPXeI7/FwsxWMU4E6G5UaH9O7wXWd3WsTGC
1w1kSIc7g/AadjUkYQD131yO/Xen0o7I0lf2yjS4Z/z/i+ML3xovT7u+i9Jom1pU17LdUDe9diiO
6012A1a8kbYOJpftN/RN0/NoyDj7yV/zvezolFLJX1BPnoiZrTpzT18eYsG/MPf7Lb+uxqYMTjQU
+3UNS2GKeVUNmQwFNSN+cI40fZAz8FPOhClxJ858bw992QbHwkemPQ4Vgw8SizNL4vMGScRRYWkJ
ItaJ0lkqA7oXQd1ctU5lWMi3MkkT4Wd81P53QdKs8WjdrD7SKxfz24XBeM0YoLH8knjVGrWPZLae
FCbEbTeGbVL6mMHdyPCcdtCqg+gt5vVeRpKXi+myI/KgO0BKM5dUh4iVIahJTHpV+iSGCcVrawQB
OBusXqW+YgwMZjkAMSIWnSoETBCkk+pU6pDXfTY1oJOtN7N8nSg5STF68LO6mKFh/RdAbuZnnlbq
TYID4A9OfAaa6PV4AjkmTVMAtw7d9RZo6mOeaQano4kT7nuv19gmM4XDaHh08JcMOy5BuFb8vr70
rnfEYjBGhW/SmuC4gQf0UcAWwrRNdK7MHQDPFJ99gcdtj80ANDRaV0BB5zl+ERgHj6q/MzORZXR3
gWloN1LMxktE7KkeuUdfZ87DSY/io98Z9u7yp5o6ROFT1to4A0j1wtEZIR1+ybf/Jo0CFCSU1IS5
ms6skLrSjU74m8b3/i6+Pf/55URs6fzegWPPWcOlF1gSVP1WvpDicbBpXwBS7iX/LRMVZNOSnUlS
vmQMLVCAkDubGjtRx5MHstAqDDFDdFxn/Rj4RxJZV2cQX+ZPJjHDOOX4dweY80PbUI7zLeKZ1CHK
2OcjI+loJlkF86sjhBnnsueBnulCQEh1nrX8RUkeYF+ngT7ZKH+vwmhDRvxNYNEmtklSyexXXdQl
p9/hZuLZTHENmW4bVellB27eljtCA0T2tTB4k7l2Z0oCpVXnh7GBmwpuxKVQtUgusEbxY0hUSOi7
QgaIfrqmCSXUhCrWlCfXsASa3JG9huX0fTA0UXxGEw8a7hHeeqdPCCJSjICtCV3zgrnHLMzkY8IW
nuiSYmF7i4sGlCKLD/+xPX8Kci5G7Dp6SG2qiCi9FQPGa4V3fiN8eecuhXWzwhZSRp6a/tuUNPFy
Jpoa+vm1uUF/k8DtngzF94MIRguPY6kDOTOjNPZp/cs21Nb2/ZcuhmdnDf37/hnoWf1AKb1PQxO3
WoWapIQI/M2+lCWLO34TWGPIS7Fkis1CLZNNZPOH5HZNuTv61PD7D3rsUeqJBHeuFAt2QOtMCe1b
RARBtTH50uiqy525kSSFb8uA7pkFE7wWzoRSL5/IGLz8IbobC0ek5ziY5L6Q2kwkHKlhGKiTBJk7
0x/jSzQRobILCsLz+CodeYH7KV1EQUw9oCf0SfUCPIANMzwrb1H/fQT3o104PczurPjqBlPdwz74
p4oNpBdClw1NP3aGyczF7XVIp1dgxf9yb5jW1DV2J/JyFZry4kuxeWq1dX1oOjkoTgpsMeNMdBzm
83ZqcSZRbsQiy90mur87gydRz35BLSCsIZuu5J1XwhJjsUZ2Nx6zLE52PGz1W+IuOcV/Tt5XUcJ3
vLZkapknzU9CO9KPjX9yQ4XjjQmsZ4Qul1MkHu6zurlI3vN/WWzayT//lZ6mSUvjQVvYIbBVpjCD
2NDVgHpoYFjnEmeN0F2qoOe6W+jdoxAo2FekMAJMKf2+Y9hG/JXArkN5vgqfb+squzXR4X+3ZGNS
k9DzTAxw5iQUK5A0/IrXOKXNQrPBc5g+YbzZNlX+MKUfwODGK6EpAqhxL3HsvTzyPKzhqE1WLtUZ
Lyx4H/Pu+SN72OVH1+91gSUnq6rTrGveX0FGYxd24GO8hhpt4nrQH6QVKoCjDwemuTY0vG2bUWhw
xuhcNw6ZnVy0evwo+lTlQvnpGCbXucFXIPA3DFcsGyFDWTZDr//E2o4kSzy1HcfSsI2bTHzGW7zn
fauN5tYtuWk/ZZXwf2V4NqSdbEfFpGc+4VDwvBSXLgyyrGGmY7CLeCFXAQYB56NvkSeWXF5+zkLD
wSD76PArVySrMSuvncSQyCGq5gPIW1qQ31ae8zvN/QXN4JrbQJW6ktDpKCePepkWRgyQDhr/fr3C
qufqCtvk1aQrOFFbctJlw/J3PQu/48bPA42E263j7uPU4fkfvw9vkf1+iUDF/dy/+fTeCbEKvlNV
qzJduHvpE5aaWdTCLwh6oZPogqG3s7H8ak5+limjdRc27dFmFz4PNENjalM0qwW7We0VL+4zrV15
Q6Vp/DK1BC+Z64bWH5A51ZcH5q8I7E71zunWMw4wanUZUwrN1HSBfoLnqBZBjegEtIBK2xVgNhaW
dpbtAOzb8hEopidDkACA4S2U7KQ8YkH30lBC8XNGzSS1lzoSQ6BIHeMJqkv+xLouh4BufcWtmolZ
4Q50t41f+HRBEplKQ98mZ2ZTxVK69SHg4J/gzrRrPSH55ZDEpsgqW5DnuPw3kNPS+HA/HDJmrqJk
TfUghUAgsfUAY3Km2LbsSGjrmtorLdro2lSckbJpW7eyv18R1SzUsPcL80++Uawp4S/4tt1wmOO4
DdF3btOi0P7bkyLdhEf3kVlBTrLeiFOa9K1m/rd9rktd+6yC90n/yV8CZDnIHA3RfKDRGwqM4QOp
SjskpEDiihTmDK0Kz4vJSj96GJhfkqk/J0jgOVkX+4ITmsrmw7aE5aEZhIutiNfT0edA3E80U9pS
2lpS0keOIIfv3x45npSIKka7aCPVoqPV3a2FLJ2psfT0sMW+0g5nkGqkgR0sfnILe+4oaO3lu1vk
f+JmBipQ8kqTH8/YpjGb5VRSEIIHanX6s/823dl9XcUegikfA3TkFkBmtSKZGgpYjBuzXmfn5WDL
AQPj2e9GNOa0PQDagLjaRQEhDKVQWEpn8HZ9rtBxaEydWOj6lBtWWo6U/rjPc5elhBtThy6wcV85
4nQCS/EE+suj3lP4EGPFQHAafgl9T4JoWM5A06F9XKGABBfnGKt5o1MNXXXL4fbCjn7Sw2Vbh3iU
RR4leqRNIudQxxGN9OthdZE+ZUKptEWeq+laKlPMW4NHgznl5i40RJrGru7z33wGhSeaRddB9v1+
ZxkKQTMtM3TfQZkzItItK5bQNM8ErprXz6ccwEtumr//MmMaOBh8YrgPb6Kdw1SLmghXEfUx+XKL
xPBnI11CZpkayhg6hC3QDICq+LFibi0+kQl5gB2545cbGV8/Itt57yAVrS9VFqhJJQd2hyPXujgG
iYe971IuJbhuPCwCFij5nAlAkTwx8RfTH0sqUjUvv8B8zY5Q9QzSO4LU07Fq4wfUJEBunHAfy57z
WWfq/BKgLhZr2EzOoUodDmcWAlN86GHpjxqk930I5XIP7mKezQngL+LwZPxXMF7OnGw1TLPLHfZd
YR54y/LmylTL+qMletl3Q8/o3oU5jBhFYnYiQzo0NZ387YFcXXkHA4SJZT5c8eetM7BpK9Trknhb
o5VGdvVCiqI18/5szgpGNCZNh14y8f9gGw5n+GL5H6teiS7U2EXPnae7/CndyuQK4WkL3eQAhi5B
5QcE4LgKhkMiLhDDga+MspujyGSS3JxqmlY4eLOnN6Qk1E6CBvpd81NidaE1Kjo3hbd/k6PIzKb3
2U7MmizyhWQvdlf6469uj1qqUun+CJEVp/7WPecgfTFuTD+GVir/GThvbdSRnz8+ACkoaPeEDwY4
UAqzUdryuEkQ6lDmF0JXSOGhuFlrZ1gZ8yMhHWRt5zMJhFx4/BybDZybvpVH8yeQ9peWbHPq2EEM
9y7A31gwuSITWK28JNLUdoK544C4IM5F/0jTjTfZI3DwBNDhF9LEDxNXzqP4MbDQsbY6Xy70DTjI
uwC56KcVGSMv/ZZ3h578fILYmTBtWCpHu0mBLi5RzPbQbOKn+zk1ks0iR1CjBG/f4I/O3sRE0zFi
DzmK3iBwjMmRYH48zxu+2juiSrM5BAA5Gwg+uRWFBpQ3jMKIyjtC+BgtsiAkMlmNQD8AD5btp7Jz
28z6pAevhCSKzCVtSna7hZanexIVR0UL2hHDe1A3GFVZBEAZggKIVwIR6sWAaLGg9RaAYRY8r0MY
86QvemuL4PLk+OxLGEbyHllI3LyRK/+H+LW311HxePjjNCTjHhUdPUnSy18dslisoRXowaqinzaB
2ka4A0akTMf22uXq0/JmEcFD3bns2BCSwZqGNERTDm49gQR/jfR0zy5n4sc4Yo4RwXPB8+zwmSPs
R51DU+QQW4IfD3xo54lLp3P5HatsJA61/jErA6CXWFvGl9CUAKFS2NaVcHmbYxo9Q3sprs/0+WyI
7nTZZNQNMGTgGufuS4tU8X5SSbnq4Ryor1GGM8yR1jzE0h3vR7v6Y20wfQxRFP4TyQET5Zh7wdYS
NRCGA4vWArG6xgOe8I+d3pN4yKsscw43SmHXqUF2Tz3zT8Nqfn/mfS3FW56zQ7bTGTTTvvE2cxNz
WBojmw6RlluJm47IzYkm8Iitw3dkOm44ibzYovnVEPjwmXwWRakw1Kc/DrjCgi/AuNXlgVgsWVSQ
DyWYS3ayF191QxP6izs4oyxDMDPIvqCH1JE0pnzpPmJNGB5tZbGoJLJQ0MIBXlFTwag9MeOugzgP
4/poo9+JaTqgbbkVizu1oOQBVG2kdfysD2RhPagYGXFSy/CfytbMnnlYFTerIpodA4GNFBgWMkgm
BOyu9fhvjAW+/Fh/WvL2GY9AVQal5gIb1mAbFLq2uRojCaJMb5P5MOrAvQ0/jM4ALzBxiLJ3w9je
2Gtl4jhRvkD2ZKTXhJK8xxugCHClYyjHykLskC2h3yFUJdJ2z/oYNhHlobp5mubFxK/gD1c57ZXV
jaVocAIdLKbstzGcdfnnw7pLpipj9JjmqWdFEJaT/dSvM8h4UkizBDCSkIjSJmS7Afy4IRJ6sT0i
GyfA+vP1l2i9gmXgp2LkSFp9JcpWYsuxBISO2PS5EG5lATZKlGiNYsPeEKNW7uhUtaTc4KSdFdGC
y7ZQfvaPrEsxGTZ1S3iRtpjiXawIgFc+qNlH2iYzB/fBWk1B4RRv7xl1zEqkd3dl110nrChvKLfJ
SK9zQ15ns7NA5uExveVO93gTRL2SbMGDxJF4jAAPdbrAuxDR7U4dTV0puU1UkUZ2/BAbfoOLfe8B
7IlHfiB9DmRBF5bMamhHjo4Ze4iqCN+7vfdFivtlVgYmtcNE/vR4f3DqQWgyU05miSY7limP3JVt
+Qy/UhSPt4jPkDoLA7JgMDZn8rvCatX2pJSlXW67FIfOLC3GPUXDXWKj5lJCoE8JzfqALODprelU
mOmMz5EETPh3OWz9cHL0moiYzqPX/VyZF8Rb7GwI1puYsJLTcQ+5fr55/TRcP83hM2sK38iOuUP+
NNwze+I3mVSAYYs+YDEf4HReV41V7YBPqnTDnjhTr8cQpY21fhlcZ18JsMnYEXPYKyNZ8nYL/4rX
p3koanR/SnlrDrCxuKYrxkVhCEgWA/bNFWbPUMlGc2gpCKg3VTfP9ttYh3g1obCSgq4Yqsa/8sXb
j0a2UdKQqhjM1T0SXd2fd588/83T0tUuF03YLY/qgxwK+LVVuMbBb+lhGqEt7gvXEUvTvE33WiRa
YrfnT+mcvZl3BbZ/wi1O7HsznW2D+qyeQNgJ6ZI3ORawZpPvIqiFvmXGD2/6z4HaYLcumOeD/nHv
Eukol/7p7ATdJyyVWptE0O9N5VzQx/my08zvW/Vq8EiDy1QyDE47HetgdqCEXIgXgl6obi3I8FVL
cqJtusZ8iEuklL0W9jdKRTY6VD2u5P5W0QpW8/Kqm0VINxJJm3WTwRVkGNINXufRCD4PgMYG3+sv
6wPUMYsgnQxTik4OoIzXvju8/L5nwKHCBtajVu9HYw5qjuxTMKq8EWzho2HugHGPeVhzC13dgvtU
AVP1WeklM8Ec8LZlnG68bnZLj229MA/dxlVm9bLnN3h8saTp0hbI2Tb/xvKdwwUhLwgGbQIQrTBN
BnZ2Zy1XxJkDdZV+W73L962yPUY0BpnVAN5XpjozLFaiqqHGRsNRNxZ4UMsTp3gDVfH4b3mI5TbA
98bsXB0vSM7nZDdq1DLf7bJy7NtQ00/Hs1JgGITPoyLdK/DH31jeTc0tN4Mne6o4AAIIClzAWidm
dHPSQAghsLqgPQqTxgYcZsd0216EdRN2H9iUqrK95KhEYdWF/FZb9axNuO6XqEnPHbici9biYn5n
0CV9cNhRxZVYTGn5RA90VLryJb31T0Su+b/mGpYTE05seiDk03+0hJIGlaYBnzB87E8ahLOCDfHJ
bEyfNKH/7t5lGW6hOkdu66ZdPIOOQcrnuir5eZ/jSnxMLhkE1QopSonlKfqOHvPADa/td72p+GCJ
Z/FillAcDjlWonlNUtmtuSsI4L5R198wW8X6wACrrtVFbgJHuxXzd1E4NQDaEcgePYeuhwZCfniv
/ERdORdwy9F+pMv8yYvTtAzk0f7DJuBVt8dbjrjVhNYiy8paB4fhazLexQBuDn7q5urqMHSDTmco
OFUUtGURYma6/wJwWk4eSXP+0Ye/KWVZmhoajupPu+GjChnMEMZDzNXYRs2te8ieea82pS9YTbcz
gLISWSDg7ABvBVXlwiwHQMDTBTBJ9kXJ+18bo/JJJexmzI1GnNZcHrux/TV8hJ1FTDa3eDoXfHmp
KxOQ8KRBTQUe4DXKPPDIWB+CeOQiZ+KaHSD7p9oLirGnxP/qUfVNkHp5eTMZm8I6JqMFjwNytDiu
mvRpW/AyVKlI8DZURn/JBzzl0CypXTQY+2WJfxR07H3ja0x/ypFaM2CqlE7gJ++bLr1GQ6nZZ20f
OwDbGkBW840w74ymdTWU21trXvN0w8o68qv6voH+3NiB4ekltTT2pvJCvONOKS7Mj80BcIGiRPJN
lPiYRIjZ0OnnYHMARKgrP5yc6AHsJqT9okDM20Iaho6bw+5ubNqnBTZJcZeB/KGC4tXTUW32QggW
MQlugV+bc2f3KqO2AxE6sOUFRuxOrjS8B8aitymd+H3BLF1JrPKpKIrqznQT1KnGp7hNFfZBAv/e
E2AOUil1IyQTCi8XzhBjv8Y5SIiyqMsc92uc05QOh584izqc0F1vlzf0+bd+gimVVUE+jTUSATlQ
xUzUQcYXxVeh/iHxUCWqc/nL+94OwrCPOy7DIqODcLJyNn/wPke8bonLP4XXia2CFTWl6myN72gv
KsvDU1faDT6axa0uCeIztXbCCEZ5p25LaUp9iCruKixYCn7wzu7WX++3dkX9Illybjpzzv6KU8tD
ahdO0mnsloYsHQkmlLPmHFXuQ3ZujxOHrGT5456+57+9g7Qv9hz3WzDc1QMTWYGo4AEZ4i3uqABO
3aw37VetXlbilvuIbVBbAqXdqH8GnhAt8bmctWJqF37ND7l6PLJ9bZhzSZskkXrbXMJ+xdezwNCe
EO5LZFa/jbbsY4JcTj/aHU64SukhGOlSDxzsLd7qMlavYR26DLMptXxD7Pkx5o3JIDbZtykFHKvs
1W6ndRCN5Hdlf8cWdXVW/bPNrRBqXZZ9xyFKBt9B4oI1VIuOOI4emuXEfACih81XeLaZE1Tquhv0
Dz1AYsounPoy+NLYFsrKo04qP/fYyLfmyebVoo2P4CsT3f3WOSFPHqV8Z35KQ99sA+PogmWAdAFe
ew1t8xbthyJOIN2/7Bdx68DG2qr2nWOLAvE6s9gYUBI3Lm/AvBHpHSbe2ZT3uLpR47FYJQzy/EMO
azevH0YVSgrysHt+WvY32ekbQyzLzK6gkHnlB++CK9PrHrmRM+C50kLOFXYsWNmgObak8XMaYllm
50/MZ3P2ncOaoUiXPxeL9xYLypucBfgyCwtMuObXHT5W1CEXepEyY+B97AjeHpxVBSL09LKTllJG
oV4t65ox/YVp52buCz49x2C2f0MuGzj32KB2FueIbWL3CfqR1LIpIvf63+vaCfMm1DOmqhvLmpYN
0OdIY+HYflmsHXs0MYMf7DnVMnVJw8v8xyqFt0dK6EpF71FLq7RAreO++rBK0iZz+s3zOq+M0Ey4
qTU+Rt1/4BGkbXuvPWnmS4v4dTgl3df0cuj5/Kk6vGGmBQsrr5KIlqclsg04to3Vv9I5EBtvj9Ac
HvDeS7/jJpBpfDe6+CJUTz2nzSXiaZfwxrxC+wPKFS1GTBzrYfeDfhu1uw9l+bn0dzENfT9MxHLJ
OEDPe6BZmhhbmFD/m5D2jUXFTplQnesPjsc9DlxvXpxllVWX43JcVZot8WcEsyR2p5eObTf2+9z7
NDZtF6eg8D39x/6Mw6BDfQG8ktc21c3kuDWuh1achsKTejFthDT+J2JP7tJDT+tvDcNcyvhTDrtG
oPepZB3pydhenJV9DSP4py7uVzaID7SRF/0BO0qm60IxflDN/ha2Qdb2Ok3QTq8rW8hfl6t4y7m3
Gn6508YmGmGqrww7/VxxEaqUMDb+EQFtDBMjSIRM8nwdhOHIwWBL1WyWnTfcAnpVx32EWoQ4l1r5
pCNGKkrEm7CwCLk509L1rWTotHYZVj27FdIMc3Rf6v3VOPv2R7rs3ukpvc3ZK6aY+rGc1Q0mXPZ8
nk6Ttz4qq2MEFLzVgt9RJhm/+gicm3q68Rkq+UI+OKoAK24eEZrjWGTwEQ9QRudGTuvPb8aCl1do
N1ruFJ4D5UAFKc09utUHLN33b4wsVUfqG0XstoFZllevZxKWiY1UO8xow8djo3YG+nmwj6IEYQD7
YdJsVqjIqzhEy/TxKbBAOcdiz/W1QaxIY1nkujbHZJCmE3tzQ576kro4eBfzK/8+WvX1sgU60UHG
wbtC0/lT2ga2JJJ1SNAzOncdrTbUoRbSN74vcYO/JUpLg/eN5de9SRGtiNzfZ+vXYtiYtFUcKKlE
Sv8GAwJZmMS+NPRPZgDBBsnDr7t50f5/umkouIv/a9H8K8MtyaBoOlMSNDmE2FfXPtsHM3gxBgl0
Efyz+aI0wprbI/qBceOPCZUTxfX3LuwEhke6vYE3uYnF5cxNd0WJ6N5QrzDNhYN/HDOPwKB4+7lD
4TmPjIvBo9+DhSVOaE/8tLcvSENubfE9i4UUhw0G5ymZl0TtE4wqH9U6gIWendmhzhRxIQCcDs52
1McTwaeIOC/ZNCdMS/UNM7WuT/7EXNAnFgOqSuRc0QWiSRb3MyjAMy8Ss7+urVqt8gHAHUNroHv8
8tXlxIY4PTfcpj7GgR0gYHKT1GfhyPSpb9D40TIFYO1IQdMuxRJ4HBKE61zt8LNlDmJPdpdbLo1E
CdDcEYnTzisg9ZdjqEJ+R+Jl0L364MlWyuIIGaaM+6+q1TO3U5Faw+Fr9V4VEcCuynmEe+2/L8gP
0toGbVBoWbxk3/UTu25F/bpttCASFpHVJLHZuRML+prM+2j7bkItJGaKNYe170+DbDuKLLv9BUuc
xPU3pCAqFcaLyZlpkv4MGuiutBMiCZM7uctDHyAyBdaxPJs0C46EK73apfBv5vqePteo4R75eB+x
nMOwD+McgXucN6pGeKxjAtGvpruMLi3yR278FjNPQNaIwDgO6rpN6AZPBrY32VmRX9kNKGfCzFcA
B3jc700q4wI9VomZeeJtAbFS/HI8twTG9eKbnuhRMLm2zFyCBUXZ9COVYRK9LF42M8xcTEDuqqyw
RyNLuT2tIKcFyPc71Hd+m34oq22MbkjrjQT6OvgP+ak9Zc1/YeZ0+l1c9fdc56QyubYORfhj/UZW
UIvkr/WU2ODJQIigInAbbGgV+ZpKGeztSlMRq1ptnZQMW9HIBMLGewIdQOfTZdRpTm4bZyZoCyoh
RUgt5EiU6c1SxcFr9Nogk+tkRsuydASO0K54fGdzSL9kbLNncQeQWwKloMZIes3x9hM1R6TAr5a8
d5Xc7LQ17ycgCNXHOIIgnQfQA+M3ahwIbvBYewFDOj4n/1OC4XBQEOzSIgEVZ63s5Ebn0C5euitP
0uAh+pPYZbfRiKbzFycUVKw0xkPHdDchchcrNIWplHJneZiYMME6zemnjAlbVcLGk4lmjep82HT7
CjoocTswxDkB2ReRF5zeUFflEZwZAhDZhXy2uL/cSg1OzbAAN13Dg7Sf1BobTA4pFx+qaPk9RBGY
x9F8TALT4y0Ng/9REKXIkmtiTkV3R/nCP3d8Y4AHuxH9fz9eE7TEHemqeCvUilsHKU/0BcDLLJYv
bdFLxJuYSl0s5wLBIRVEr9triCCLyOF8o++2RgZwz6Z4Kpgr6f+1ZnkQKpLzb3UAv2HV0CLoaYvI
Cc8L/EV90StVFrjbXdC7c7ZbpSl9BAcw9PyDtRkZMb5VdmRAmNry1x/ZUK7Mz0+9FU56ljQ+EfMq
KZ5Ab5ZmVtI9o+oaNNIJmeChkwVgQ8A33Ao+Nv7Pq/5/kRPi5jXPw3wBibx4bOFnPcRZSVXIF2PW
ZkCzVGZFFl6TmGUjPlNBNbS+seGgsRKwBf6dzflFCI/mgQ2ZyYp9dZC06bahHd9n12fpydOQnHda
dHynsY1mA6W/zjFGEK4KENXyHnI9fK/oJB8As8kIRNB9FPMK5ViQuVKAzybR+ZHlD//eUWhosAxs
l5rh/cKxqgsYzcy4aYOX5rTFw2d46/S+4qr8Tzs4KjNWXCboWYIg73xq5Qb0EFgZt3Oq9WbfDUZy
8oiV2m4Kgo51jY/rKTPPAuDH43XqmiP6BIj9595p6ZHi2ez/pF7DrOco3Q0OrD9oGJ+Gxa7mg0FB
ZFZIIbAfN8YzslojhtPZM1aAxBzwwLUcnF373Br0x/aTcqztgAi6OjTmHvaQZQwXhObbgQO6s88I
j7xW5wE8X3xbIJhpHaZrTDB1qQjLRKZXME0aNwNMB6XPD7hfMjPrly6a3NaZ6SJwp2fJwAJX0vyb
88lAABB810W1oljv0WmbAgd5qOg+4QiV0qJejdhk3pYFFnDnhnSs3dgvCOPIAG3SXLEeEVCF8ADT
WybmgLJ80N2+P9nva7RJvRb+ENASKQORWQ8dpiNMmN31xsMVmGBR38jF9dTEurq4BUas7bxsB0v/
DKnm46hWv2zN1w52e8qrmi50qHmVWCd5/yLsOi2UOcEtP0wIwawRS6jvFCGGBwXh0Mzd5cvFhEm9
k+/ExQPKs5kvb4455hnQnftT5uE/eRE0cJ4bD99wrn9ROTjJOBAecmx5T7MO1Y5XHwWtUeMt9qV2
hCa7oDMxLEv5PHCnhNS9ugp1IZzTV/xcd/FU4NwpRZ3kQZuRfkABZTAruz8OxZ9f+hp3hJvrsVXX
pcCmGIQI2X6eKHGtYHJbW6IhRFfWplsGWpYjqujP0aU5ZonumpWOQBOjEQWSqpS9foyjbvvTkuEG
SAfmmOEZ/P5lgU/B29q3KfyRRyE3TzrkBfmUrOLmx6cI0JBx7AFhb8xZsFQapvIeI9+2MJmsY6L+
/HqHxjqYCjfxSP0B8xGdQ9/or52DUH5VoGvkOF7tKrEdfp5AvgEyXrt9HwDzMcdf0LRSfNaPwIEu
RZ85dtdaefQsNxkh/CZCGoRRkFkmMi0UgVkm/OURlDmWoAjhVkFDcEpzYCmykFQX+yg7vrSnQpPt
bFVd2XpfcDJwJTHeLcwRWVfuPezL4MvepnRz72yK4zhLUCmnurnjVAo7fw+mNfykc5Fa/Q+ikQoP
Wl6rDMTe2QdBub+m01qe1NUvXUdQqMYSpFrh+Uls0vsSfY6hMk1J/MODTb3f8m2SCt4R/FTKkrO1
wtkrpOLhaClHZJnTjihy88MLWwWIFhjshxIf7SySnYXhx+sJrfJYh+YgPny3D1cQInWkz9uBqQnx
bUZZmRQ9/lIwoLBmZE7dXblnatwnwYfk1acjvLDvhz7h09lxVnnRRaqxUN2BFCPGpdI20rnT/Eq4
Y71H+yvHEbDnSy9KnId/mrNLKyI+dOCXnKYJeMcYp0M8yvMFQr/EwiO3ZDLBXoEyeQQEWFbeda7Y
vdqwfoC7fZXj/6ZcR5gposhN0P8PjBefNE5mcah+JQL3dsAt5oSXyEtWeu7m6774LGgoQ1Baim4p
YdM5k2Eb33h5rZckT3REpnYNyh3j6hFBFR18EXO5hb5BG/Z+bpDXdl1MqkkwpPUXDbE7S+GjuEPh
O9Ni8DTh0UNZnCM0X/D6NZcqx8nGFgWcS7/5ydmLDBaV1EjQXpoKMa5010qkv+Y+HnQeOu9xjfi4
11Av8dOTmHa7AE5mBGRBKnEXubCSbqSZLrQKB7ZViXRrJJeBlpursHDYkuxZ2coKrjKM4Ccowlql
eeQ3QEhVt+QLeM3d0RLx9u4ZLS90nGoaCE4uprN3VSlJKMXxZS2KTCcN+EGbH1FZEhZFiYHb2ZBn
4xIqJHSrzTFJl2YNksLQU1cOMR5F0NfqFMC+8093wV7NC1sz5Oi8xdU085HW4DZCu2cJipIE/5Vg
BoUtTWS6mPBEe+/Mh9xldhVvLX7TJDOfwbshcgsyp1FogpsTpLPv/ssB+tDvlf5KxM6TNtwrTgI2
IABxL0fXS+iUD81u3N0OpGlr9XqOMg7YG0oyXsq39v4OKkysp4zH+tSjtAcOE9IAiXN7rqxo46Lz
RwZEDiXU6u2QrvPegIPhsEmg96EnACWHCtv0QQRC4+gQhZLZNFPG0+aA30uU1ZJsvyt0d9XE0Ajx
u0HxZcVqgTz1egFogy918B1CFTywjCvrWsMwJcSVlXHYSBmUctKWStCnBsMTvickzmD+G83MSNLj
4Crz01AQTKS3QSvaQ0G1jujfPtmwcxuXmD+LtbaExwznnQXuTlpWBcm/xS1n/AuphUk3VwaC5lwS
LJJ5cix5sK/ihvoMk1QOhyeb2QfPOHxNqP5T+MPiLH0RO0Kij3Yhj3zPVkPRVpltRswxABQgbNVm
oPMpFhPxa7EDqu3b86xfa8Fdcqjd5a1oQM0xcAUxM2UmQ6CWAOfgxoRVG4MtjRhAfbxZswJcTIKQ
hlkkHfMdOcaMmBXv8prSGY7WTOxYCLUT+bUsEZLZwuAV9nnl/qJtBnCA4OGLDFkyRxTJMxP8ZeHK
Z6FXUz+MmfKB50hcfUiBuspc6gr8GgzvEOL+vGAOM+zsk+LXsyuptzGaVIAjMeb+TiZ1/8LuBJ4+
k7qSS5bOSBggY3u4NJQ+mojXHR1rIwwnjsQur3EbOd8SzoRTD8rT0rG5/tYyohOHaDZvyVfCaKmJ
KT3WhyoGVUG3oA8drW2l4OCwT/XiHyc+q7xZqx1RfAVHxNXNgoebG/J8ykssZH8yuThObaDMh6VX
McFdLa7dcgeanNSMilAb4bbvezIoWvtvpZE0z6p16ptto80MEBn3ElTrUK7oNE1XZSozgmS2aNWS
wnj7nNzkB+s21UBZiBZa21UsVdPjsRYzutqZc+7eZYK9j/GbKm33r3YVboR5PxnK/ZpWfOu7LeCI
wnB2bnzgpYRLd3aQ1MPfMrBjypbW0kw9x3ItJ8Ag7spshDQRUdu42a059TtjzetsEeHSROihtkYL
Mz3e9VZJ1rKbOSENrWIV0ZrutbwX0rGgXfCvKpxQzd2CZUfxStxlEU5/6acfmjGQXbiZ9wl4aqqQ
hkMTzbiWtfE7gIv4bjCbT1dyMlvZ6tEwQq/OT3aBalFEFV3T0UGRexGxyb4HFu9CoZqykJomJDcA
0g9ZPHbJ2UHcX2WD3hGVh6u+kXPZH5DO0hwuEPReUXNR35cQLjjhFOf0ylhBOClaVJhMQOlrzlCT
eJ+J+KbEuEoUtRsHO7HbRDzoUKRRehABIpi3aS7t4mWyO46tBlxNyC4k4WbmR7dUqJwH0cALTC9n
jzXNF4Bpx4VoRtET4lRkJKzmzlESRLHItiKJ/7/ahAR0TeB/m8IjN/zR7ujN5udjYXB5SEvroSD6
0elSHvVox0Qr+rcu+x5BSaE/IruojHkxe3tBdkm6H///ZOBG0dg8R6WBHZwtyjIqfo6jukpsFHYP
xwUJqBKpsbjJrzJ5H32LbHnPJFXeg8JTnfT8CwSrS5H92Euh3GxScx88brcNL+977h9y11pDViiW
VRDKebkWoeaDsWnUrQy7Vb+yxnmwIkIsk046ZpytWTR9j4oKlx5qLucN1f0jpSYDs1JX7+edT8kI
YlKkHoQc1U8QXBIjOXgJyRY5J/zViwCYoUCkrKxIGPiBtYcdbEuNlDrtsJGCa77phZLt503upa6r
6Zo7pKVpM++XOdh99GAoiSEBV980XrGXTOX+oQpVh6TpodT3BrbfUgi9VnczI7vuQmeUDcnLMf/3
iPDJufcpIJfUQnXFeAtnuHTcnDbsrhgK6cESezoDI5mhCIkOmA9RwZoVvoX+3DMhHJxH0hSDhiiV
KBRlZSBxXJ7U4V49lUXaMqdDtAY4tPfHtuScRq9OLtYZDX2YjjsKlkngbq8D7HCZnrPlNhSqLQJq
4aEeCU8lEa+N6QEnomT2h6iKuGLD5S10fpYUrO0J97Es4knde/Tartjp7O3+rtBpBg++gOR78WOo
5ry8xJK/kbzt/B0Z6IsSQ2mgBo8Es9GtNUwKb63Rsu+T4rh4wNrFTFqwxmNazfhnxmJ3NPJSKVzZ
oHpz5cEUIZd7NJya6ZDvoHaowkWVQuZblBWpwO/05ms9WSO3wSlZ915iuArlqxSfMP3DmWjUKCCp
ZG5yHHdBnRXSmJnLFB1KBdAJ4No/gUnfjAQG+Ne1nQBWusmJbm5Cr007UTNZ76HLapAp/sB66+43
PThOzcje/N2zwiYIHoq51A2WPWSMQJIOlJpSkbQIZZhUyqcK2EYMztmYJga1AD8NrdR4gQTA7ANk
nJ1Kl9ySWUNMfA1Xx5oTOvO3yRQ/qE60J9oHNIvZ6xC2oFHq2S6M7zMpbSS7rsM/csA3QvrajbDN
Wcqq1HRbDqVx/VBK9NxTjujezCWxzQVOFs8H/ztmo67gl7jclAmj0G7D7UatHDKbZX+TEcH0ulBv
ehi1ejD3Kr+TLraqlUXAuwTqetwQ5oCqaU6NcseOVd52JLMDUdQR4r6iBgL8gn6JXL7xdu1xX7Uv
oZRJIiAMJ34qIOawLt/3NuBUPMJ5gZEZlfUxPR930VgKro03a4ueXTcMshPtUgkX0+JtZA3HenAT
hhVgjPwAkGr4WOAI5K33iU635EQMqKslong+JLzTCKUqyYLpf6d7zB1eVIPOH7RZUF/1VfCjRBp1
N8v9ryGHAAxo+is45QTgogagHooQ6zBhKSeImOvSe/4pqtvn5H1b3i4dixHY3Bvt8MRQ0AHynzTk
qbsqp4djBPwEezuynYW7dRTJmqCcWdBDll8fUK05F3Xo8T6J30Q+n7htP9pJl37h7PJzy8AiSEDd
eY4EOhx1SHs0kXFXrco9r2ugXo/Bc9aAbUM5RWR+Ffw1ZDb16v5s3yzdEUv4m2g+oV5HDn8HoMx+
mtp5Q26Q9E9fzw+cYB6VgABfduaKhb1kXmLC+kP+MGTZHBcy1XfTXsZqtfHxuxTloVg3b9Z+pvOR
UM+Jy+hYuTYGnOhxlqAfM48YHM6OLagSeIk/3bcnU46/JYMNRwZC/5xAPN+yLMht8SDIZFQauZnB
1FIcDpcdDGnSkdlPKTBz5yvZ6YH2mXur/abGo0Cjio4QVu46c9o1MFwuuKNYCxbpJvCWq1b8CHss
chTvBleNbN8K79mYcwxh2YXjDjFIQZ0k4EQO9n5n+7t9pIqbGcVm3PZ2frLvCOWpvPbgA0zWKSfM
gPON0uGEXW69I2hxSZ6vJB2EpknjUoCtI6HW+SOhTjjQ1/DiEqRjJfcecjD+iQveaFTB5wZTj4IR
eomDtEJl16QXQH7VwwvBkA4Q1VgM48E0lgLZwE4a6rjpDxUKZIklo2nw4DG2pvlcZk9sNEg6jQpQ
R64mxaHhqwOh195Bf2C3x35xJbdfBZqjKNQcfDfa/8Luq6OcbYtQzf22c9MrgWtK5Le4pNRQSwQU
EALak3rjlvPOWAeneP4zdzyBgqH1iVrn8TQe5xni4xw0wn1p1WOSsaxW3/LcAwrOHM942pBzYxVl
qGLLPsB3n9hwpgPaeb2AlXajU2flzrjTbXPXwwzlHO/N/4ENm4kAjdbgn9FeKjjwMbm/4GxyFHrh
cnMTnvZ7ABvZFstriNRCFqR5ik4K0mkbaR5I/m+dglC7xFV4JqHFbUlGyXJGObO1INpu2zgTf74d
HTbjLgdVyS1fLOI0HEUh5EKWBCzCc2kCt/3ANMHrRXTjxGxPGkuEND4gKZc5cfmlHIwYJmSjwgOj
9/ybIr8olMsS5tgazF2vgsNDblzo6/0WUnmBNwja65sCzfSKRs0zdsDyZmBo6QON6KjiV/3vHGTD
eg8l0fSbAzLe0b81IAj4w7UPVO3ho5Po3kpGcZjSjCCPTClEdBsgmkoBWURlM5GAYtCpLhm3GMSl
ftnSmKGKhljeWIKWP3ejheYwwU56EOOyDrv9B2JQ/LPkz8zHtcvAtpwRJWBsj7C1iFdgOLPKnkWZ
Qy/uvLlFBsrJiAtTJI4DDbPC03YA15FMVGK7oVGwxP6txTVDrP0jzuSDR1Sdy08Y68+YFxkoqUo7
XGMQx5+u1Xy8htbc97qdkGl+aTzE0peOdeZ1tZagLnsLilVfXg5TWIXvjtGKyBKNNbycqC5HyUBS
SkXdWrdyP13ph75FX6f0EF4oBw/cITZbhHWVk0bo6C3Tw5D/V2BgScgp7drV2Hxneg2EplyHdwOe
doEc+/JlEhzXudkFKibN3OcLQ/fVgkxPo3HnqJCOngsZihTA39nxINgZ0ycPM0pGVNBZPJ4/8rgB
jpysX6HrUhVRtryv7THck+WNDTe6vLNcCrNzhOs9CX5yUkplVBveyzbqRbh1VIDKHsaCF2BMJhc4
FZt83KB0gq7fhkre8JAqQFJ+/RAWZB3+zGs062DE3dqw3PeViiwsQPUuiQewF5CZrVVi7bB8PZkK
svu6777pX7mSBCHOAW29xveqPiaktFIeVzr4I02C3FNauvn2HqbYNPOQxwItV0J4pOkPb4N1kk41
M4xlQV81cinc8JzTXlJlD741Wte7tkeHUxG65bgy88cN7ryckMd73sml8hle6werdQcJ7R4KtTq+
66OrhhdHbTJP5qqw4MMBe4GRRZI/f6K5S97G/58ZCqBqV6xBi5CPydoLQuTyL8+IFWdbAF2LX22i
goMic8/NFNiCJt5tQBUsfvT+w7t0+ee0KbiNO4ihj/yxnPg2bYLH6tuLnCb5z81PDVMdLB4nbye8
14/149nlkL0uwmwdKc5T9HW1b3iq5dVlLGGLewjr7SshqYODcUYXPrDer+goVsiUuZ5cPyOzr+bG
qPtRAsWtG6jtEaRWdlr2OaZEN3BJ5p/M9b3fSJwRytljDIrIF/oFSomD8dd1wHpkbsYshlunD6L0
SKwZo3GUBkk0NjNFxksiBeld8UR4BWuYeFEjDNN1Ce2Xz8tGTEbgDtoS9MqEb3kIJP2Ys0ZRqmj3
O123q/6mrGNhWVhapSB8/zT8EQw7fCBIZKQWSx0SJuIWw5ohkY+qcWY9bNTwFbIPduyemrmm6bqL
B6d6+qSAdYFOs1wtnPpv8HchgOgVlUDlamAmAfB+gvbSEG2sA2eE3G2YVTEAAFpmIzqoH7QH+wsd
CID0s8CWFX0vwmiGhh1mCYEx+2Uj0xivJMhigb4UX2BOVa7OvnZ0nK/bhVvfODg9c5W+LHy05Xzu
eyIQUkNPqC58K7bncOPFHfhF90CXwnHoQUNTQ7xd3lu6nnlhV5Ce3pXLIHD/kl7aekmUx948m0Wd
sx23Fu32nlC/g3911pCdQqSsgCuknLItSoQiO5mTrGggdj7YxwUTXQhtgL46Scga59D+fYQFm+cE
VapzR3o5ktefFMNd8Dcy2G9kjM8JOwesuy69CyEamtbWn/FYLdyVJ3FLyYrM++mnLE5zEidJTNJL
vJvC9JQFC7UesO8RUwUj6NGG18s9uahEv4gNQUyTANwarmASh/0pkydLvWkSOV91CrQLeCXQDZP4
BcwSul7urPvRdr9bV+KJ3I3prwlm1xArR965vqaRaqXd5ZuMpsd+OwwVKSBioQojjGCwI7RIixqG
4H5gHaclSY9T0w6vfyQtl8yM73UDCifMKqgGL9+5/gl+/3vyu/WDi59DR6z3ev4V488vBlWaEzzN
ElMzPvEeb73mHFjlILOgKxk9OCbiDREiKKjedhFPDfwDnPCwL5WVYYOViCsGyZCAwkQL+H4CQZTa
pMc2WBFQDIwPpc2tFez+1A8TlM2orFuU641R5T17s90W5kKT0kHdh7xcscA8g0bxXg9hMyeWFe/j
gX2FfQzky9gHr8Hl/+WU5c2RwEfLzKEc9lr75IFE94g/ErjSS4XTQK0WVtzqLqM+aZEEZq0E/zQM
zDQZS4fdjXTWdbAI31oWbwSawVj3BYUY1jS66PJjDwpLgO3TIm4EsdiFdfCe2x7z9AqjSCtGWdYf
XbNi1xGTWQqq+QpQI2JNWCvgWXiGrxEh3xSL5bAwi2UAt6/Tn1HmpmYBAqcWi+Q8tjGM6xl6sTUZ
YX9tO0aZrbyZRscHqKuhccvl0gzSt/fessong0nhoF3/OhTTySE/y1Tky3NOuBYGU6MsOGdifjJ0
EUrUUHV3dRjDJPXgHMtbC/svgdyeCXKIq1c+9btsVFZeZHpflDxUvmmUcml5xOSgxo8S9lT6yQuZ
5oO8iNwZKNRleXRuUPn/MAur+zr1i4cQt9zW96r4W96sX7Lo+/NObsIhZrfe3XUIHO0sAZtn1tE/
uefVXpWGvdRiZN8voucLC8i94wzN8dSQrGD3+VuA84L3wPShVEeIsthnbovTCOtSNv8wONXTor4c
tVQ1lrRAZQqRD9khrg/AgzZjAzNncGqXy9w0KnDvGHicOBDfgq1axEx6vzfk08FVrqJi6FiU80bX
lLs1Q9U8WpPxpLx3sKV5XOVvqZ8i2Snklobtb44frKe54UmjHynOU07Nw0itPDec4NTUY6cYyuUp
+wusaA/8eFU91kSjIdEvpFYWcaasNOwsFb+T9ef6053qxeYxsgue2AAqhC9/+F6zMTd2YYxLR+e0
2AWPE3P3f8bPp2fPLBS8DnSBPuNLkbr9ZHccuxlePZrOpERalOICTqfFh/VslBD9jK+nt8Wum2et
4ajF6D/6yzsbBalkulRpQxT+bDCiyjMAVGrQ5CfwYYjMrBlmBHTNsd9BquRjJfPg4VDUMayLDVcn
xxzfbC6/XvJTBsqqbiHGKlgWNtKviVLlV1yFzS3kwxXXjDegzpIv/IBaj+cLkvM01YNDlbuQOKWe
z1hmoPbR98sU01X8IQVIFj3YGVl2K0+q19iR8rbicsEROEaB9HH8jY2rqpzbdPgfG1xgN4zx8Q48
BhRjb0l84tkOI4AoC19VMCcIO/E/Mv71Oq0NxEPLQqeGHgMNdxo05xZyAJuT0d1fjeri0W9VtOMW
PbeMm7C9WQwIc9oInWHAy46oTRVLWV5jZ6VThj4K+DUW6DiWxeoEiyN+P8IdHEZvhmyCNlmVbkjk
DRDu8SidtIcU2iM0O9OmbMirt9vzJeZu74wXrLSOmcBSCcCHETb0IPOvSI97iu/1+/AAkIsRbkof
YHbw1s9UJh6CKs3O8GOq1WDScuhpEo+0Qaqb6WNkpq4by6YJlFsBSppFH4V+0QeOzfYYeru9s/hI
laRLIA6Ie+ieAwXDO/qLVRxyncyTVAbO7qnVma+XNMPOgCLBBunCzdUV9Q1lv8qdW16DtPKQoHlv
8GzEfrjuYwMsh2S/c3MMYyg6elMtHQcBhchJe5C+ccRikDNS5c5sHcpuplNMSSrXkntbc+T9OC42
S6/fWCTj5nsq/arIr/lswPF4PcKqeef3xlq/+AfgPlGUvmByKQcc3yv0W1AlGlaEerHgmZDXtNnK
wXWtGBpDfVG8e0Qh6kexttuxAoX5VvX06h1H+0japJnlNp/IXlKgmr7TQc5OSToUp9HK06T9Aq6x
mT3IIqJRQRgEzV0rDUE89cBNjeSVRYeWaTp19eDAqfnR9Fa0uXD+6YnlWBcvvddnETOiPUUSeX+/
MMBvdGGIi8qr/n88tRB9ADwh6+ZNl4x/tjOiGDR0mcaNHjyB1Xovv1tFhzcvb39JJpez2x7l4Qhw
vSfBSZc0Xnuv9mb2hv371B6Fq3i4YmeVSjFl4cw9MF9NIhSrqKy67q2QaEa92BjDHTAAmDQu28dF
abPZ2kJRGthCBAayrKNerOTW4piOJRFniQIy0PiPN2DCk53TPsDaXDgGkpDrIgEj1rtcVV9MzbJh
WDby7Ft1XRY21QxaYQFOsvgdZuNnxjEV1FFGIqhLXZ9bavmcy7aI7DsFZ1VX7JYqyG9jypBaHlU/
Ozb77N9wwznFzGTLe9/IFKA7UnKbGZQFOnxUzS4c0a9rqDW9P31rUavNfL5oXA95sDCCiQSfsG2y
d3uap5sftCbcmsHxbud/Jn9pggUqAKrXXPO3WyfBDovad/lG6uOE54nzI2wIRQb984jgbjPBnKSM
T7Xq0mDKBl4dxIqH66RaJ4B951+GRc8S0CO9OsZPiaK45bpuBYLThONPBG0kL1lfU1nada1Vww5m
wXOhmvrA5qMwbyMImL9yu5aPyQIWrNaXi0BsTnxLN5Pq0eS+xGmtiz/qX2kdmtPl2bjvmmo4+JpG
v+plAsWSBo8ahttZ0Uh201rnkTVC+XQ33ZH+sCb3pvpv3NnO/coDcN0F2NQT8hLVuuRbRKN3igvT
wfF7GMyUd6IwVAWdb4MRH5U0Raa9QuA3ktmd3tpdTGaOleBbNd05kgCdJd5VvamjBR8SbZwehYQe
no3MQPjq40ALBgOD/bfU9owU4lewnnhf736Bg/jIn0l0o8kX6ju4I34HIuXlEJkyTzviPjCEEhyI
1aLrZVjoSuYWrwhXpN6PKoGy7XaUHvHiN94z09+HT54h/Sx7QlNFYfaPSBIJDbuHE6pBTiTNydDS
fbgHJZkfJRKeO2lmzYg0pAA8j982FYqIHqOLXY+BMM+38EWAS727fCMD35vJheEk+jNWa7lr0+h+
LjHM6Er5hrwdiRXhJYh9ou4e1r0tTRI9jcHnaZFC191pRpStWOjEB7cksPaMRTmTtHhsSTcUbfoJ
2+kmeWe3PA/t2ZHLeKOpVjGCnsQcrzVQlYFa7M96Cfn3a/9lzKpsBvrayctvC1MeVsrYw+Yp7NU+
PEE5X8s3D4mbZg/OBC2gNZ94dkvaZg4oVqdMSUqGyUFA1gls5Qu1K1q3V2fpK8ETLQ/Dxgp7CSB/
1/kWIsIa7QSCkd92pe5YHBnMdgHzm+e0nLyVQwuJNxs5Nvz7q5WYNvRpKc/Jj6HS1MtqXeamwhOn
SRYs0nXyJSVmHilzqu5DNbkxVySvR1dx7+trPkNoPaeO8QzprzwurXcsFXJ5REkmDSMY47/GJ46t
EEzIi9gY1msK4SPysE41Xf2CdHnMORlVz1LXng14oLKdG6i8MnOpJOrIoYfArKZNrAsQ8r7usSYK
czgi7a+MSjmYTJLhujdLdNi+9IELQB+3TM4BxtY6j+9nMmTVkWXQts3mXsQxrUDGN0oVj09qUxlb
ODF0P063x0yoyD8SL3AZEDcBsHD2sVaHdI9t2DtDKupMh/ZNlbcqp2+xBOBWun4gDQ7kN58aAEif
Y73L7MZ/UEfc0P7MuNUhybsPlMFKri6GhuaNd5Urxn26yYW1LQej2rGiZduXRY/JNBxTVW6glCZg
kpslc8HqRmjQPydVAEPt6YckfilyXUKbb25INDg2CunYXdLeg5OzsHtb+Yk828E3QS+y7EakN8Sz
2QSCHHeFROKPkVfAYIWbjiPefJsv5Xpnm/51ZL68K2FRkCn8xeQSFML6io8B0kzuFcf0ZxzG/RSw
x0LRATwbqg6oGuVEp6DbQwZWP1z/pAxzrVEA8U3NoMsT+G1RAm4VPF9A5n+XgjgGHME3LRgoGLve
0F6bFSP6t5Sn7xFJdaSz34hmfvYsD4ZY5+YKhOg3pPQYnePp8cdZUOFG/P80c9Eovyc4GQ44BuHA
CNWstsUTRUxYnb9WIWdKqpYzrw5t1/LG2IeNhcIkxLX2UYmVICaprU+TIe+cQdEJOrpR9I0HcYbs
FLmP/O8A+qxsLlwZaN9Xi2YZWvIIuFL0Dseg0mqRRKUr2oHMbxCn9Ga6CALACjZ3SWLn6x81Cjha
P9H18bzdUoyMWG9Qcwk6U9xM3yHb9AClleFXDUuRKSU8pT8Q3PtKn12ODGYCVIc/leqdVbJ3HDs2
FaE+vy8Yses6OXoHBh7ULMmm2TdxbYNUDP+U83rHR7NigNxrQb0Mld5r14xeyrELNFIcUyWMMUPT
4ANXRdQJC69AUbScW6MiCfKA6W01rMQNklM26UVKp51akfJXHtKra01H1alceoA5VSRBhsLFvSft
OwOx0TERw69xyhDWyfZFu14FpHTsdWk5Hy1jUBSrpr7D7aKwz5BcM7RssKfu8AXbg5CSZEsTc7vS
D8xKPSq3TyAPXAqstXXrq1yKc/14jrmq38vfQ94GzADJ+/wWf8wGxsxs/HI9x8IN4oxB5xYkHj8y
2MZOEIn3ZoQmEoiBfuVNcARrSEX7uiEtq9GR+x7vwJU5+9GfKAHXgmDqEkxA/4y2hJPLHAK8PZ8L
8bSgUYogfq50+G55v+8CwSlGf7j4gYzWdlFSMgdyFe9kWCoaU2T70Pv2I5jOuAGgaVHkDNB/Vw39
CwGutyznvudt2SsUqSaxyFH0qSnMKdFSKSQkoXUgQRtGB2MsA3pp8JCmyMAkdHqCwtz133fhkV9D
oldMc4RcTBRg3dm3Ck8G/ltWbi7l2btLw4CuvwLsAYTb29oMhoq19NL/7rvVs7pEvLBDLV9/2b4w
dx0pqIvwjj+owMaSVxNeZD3nW8L1UoN9wgdX8HcATag4rJKf8vpbuWilZU7ghJ8n2zMv9hFtM+eN
jDPRSD7OIQWBuubWLnUPewaNLFVgQrYyA01n0uRHfSQnt6Z7fgReumLVgyCS1MnN2+8CIIM0pC0g
qG7khVTDsUXI6PuEYJ8epEmj023pI4AaSEUgN5MUO5KiROsgMVnDaiCIO88ApxyyIaD5IJw9S/yk
Si60YDwHyM6/+9lnPmhymIpKD42wbAyLJhG5Aq8QUz98b9pqG0EnIt+hYOFMFqzx1beKMIYOSmPz
m7NcXSCSzYPkyI8nGrSKpPPaevs9h5VX+KA6lA4hnbKgkWNKXTHwhZud2mQz48r4ujJWcLHe0INr
y/bRabLjOJplyge0Hkut+G44+2uVLINH27Cec1ImQDNQjbNcqIsB/MAjlL8Su1dQYueZV8/sQT7d
/36O6pwpzY2GGK6VubPaD1vRA9O8sDiuyEHIGYKVya/OaleYHMG/thAPSRdpR8kA5WAXSLDqW3Qp
GSq96otog7EFRCC0XjfuSm9Tnn7erENIElNlBCwksGjwMtc3z5dI30uIo38ZcyLGHRnXlYlmavJC
9UFPqwFlmqOACAsgB/we66uBLyIzMPUh+BtpbrTPU4cNOWzNcaG1n96myI/0EFzun8hWBHAsm+Jv
1KSeILwqct7FK7fsgEsa9/sjxMb00l1NVs2dDpMHtAslnOo3AeC6Q35jGB991/yGOM+LKGDGcX5Q
xWB5DWeSYlGF45aocZa+9oTkxPPeCF6wFW1THye/TOCOOJmrdoxQ2WoxwBbF3DOMSUmMwIKiNwaI
kfrhyRnvxNd0Vj35ag+Gvi0uUVAMN8Vn67FsGWZqnvegL59X9+iRh8VMo51kZjKwe5jkyJwk2C5t
KU8V6A2w/u31YE3ZqVLt0VAVYbB74sRNG5yB9ih9C24+It55iDeK4RSCrfzLDFx0kJRppv2xbIxw
8FLGC7ckoU6LimrQLUYSo6nfhqAzkDqmhYsxjuI2Ryur7gvQycwR+jfbjJV0kV0UEhZVMe9H2fjl
3oJclYj/tAyh2BYyFeMrRGJZEmJoCOUiA3FEhbPfduhuclGvllssFhiaqj1pDkw/qXaOcdkYRFf2
8gOn5Na6Imb5YrFHNIGp5XBdqYpo5Pf5fQfxxt9wcpBzGmGeLE/sLhbfDZI5ww+F8wLR9QrIEleH
XfJfi5VYvit4BHqutdjnpwJo0CeazKyK2mUQ8OTfVP0UkOJi/oYTyrZw4YOmu4+EtiSwUnWF/w3R
yPl5jJaXdfuhMULxOiOpG6SoVHMh0e9DqA+UZh8DAfALC3ohnD8theXqDPUOxDJ2u8cyvCGSwB+Y
emHMuRMp9phu0I07a9ARifKyPvbHWF0my02R2qkPBZmsTjPbFejYiDt11Mz3XhEqrgAUXFhSSbc0
rFCBNH+VlK6O12/894q5AfqO0FD4hpV6mmFdJbwLpyPIMsPJe6HcAdDV+k+DEPOQemvEORsyjFVe
IDV0TG33K60UwL68muf+a1ujGmLoBXPPUnFTUq5IiUGYBDuxjqkAmqONMrhmNFnQDskxhEUExAMu
4kda/CLFeX/pvcmIDeiywefx6W/eVbMZKf7bTX6QRt2aVz3O5EejLC4qxIa9aafoeFME3V2R5OYn
YT954jNZpJb/xGiPnGxIxl6vzwqI4QvRyssiV4R1vMHt1VTt7qP4OAMUdu5CetvUVriLMYvFDdhO
FPiDGHkgw26Dz3l3hTIYIVaUIBjtH/hVGGGcPubHcAMm7ObM6EkLALkfUKtwO1ZM10KcvJ5DsEOl
RIYWkKZzRiIPgKFIqwXbVzS27anKB34x4A+Ewbu1jDqS9R0qXieyUT3HCFIVeO5HQbspS7JF1Ioo
fCk7VDuCFdS/Rv/LUTCJwirXN8BHIb+3iibQ0dFGxyGca7hffNoU00Ke5EsFaesVHKUaQ31hU5SQ
Y7f8sK1IMTR+VLXfujjOJBNPXQRoeEISdJ1ioS3fE1LBtfMjIwoWUm/6misS58qNbilqCkA5MWCk
jgMZIcEPG+RMUhEPX4rKL9oNWGKf315XMC0tWng8/2hyNfwWPaA2Rxc98YGmg57g16HO9WGWjCfL
7S1HdZVI/uTBYaGvWgrBnKqwzDg/rdSdhU/L2+wswYYG/UFI8aIF0VsSk8MnC8IeWmPaLePBYyYS
QwtGdGwCgE40Ewcp9Fu9I64GhRI6syvRjZwuhjeM6MaTIyveE9e+Hpsm2ZByVJ29NQTaaYiCgVf9
1yJyhPMZJ2wa/MpJ1sNV7KeepYzS/ClM0H/sUaQ8hCJY2Schs+Um0HKdX26QHqd7tx0LRS7VNazk
W3qAO+cl25AtpvMM6BXpXvyRQvYrwHyODSEPNKanlMVo76oA9cPVLT2v25b6yilWvtM/+d3ntda1
lXAVNDDX4M+30FTmQjVbFR4cFt12/7gNVBx4QUfsIuZaWR8hYh1h5h6OJutZel5zDz3JlN7x772w
wzewk1Fewyyws/iq2fojYEz2LQ2Jw7cYq6nEcY1fIGT8P3iyvdDvJYT1boVyhOagmc3gdaiVDZI5
K0MykYjk7QMek79rr5cO/7d/+MEzuQAkKLLq7b8J63H5Sab0NNVPHLwXS7iq0LCxOHhTRpqd+Kpd
E/zj/9KezE97urvYNNcCl+lqBGG5fSPN7c/Ehe79WpNSKyIK4uA7Q49Ep/jghd1Ab7LJ36zpTIiY
Z0nISljP6V2VHKunW5lfTbJeRThYp2OORSeRNnQluen5u69LkOqFK8qbQ/Kfph+z1xYXa6tYSnbB
sM0A9/NzfvFGOiKkZj01/4QMSU/JbHdTZzdBC3E2vCu/RdyhvDdaAAAcA0YBwU7kheu1NIsA3eAC
FOHDgmSt/92wq5mEFaaekTZa+HoeKtbFQcTmWXxLJeigL/xy0ZjfOXn7vyKFIrzSAk9gcHmwfqK6
ezVjRUVB2VKTWMnowDrtdkb0OSdT1B8cAWnbnbpu+cUDHs4Syd752Ys7x3SfPG0J2UaLhMlclL7e
kyTlrlQjz9LXVw56kYOaFHEQQU1RC5KT0a3iuQ8ssvrRm6vmzI2HhOaONQhRvJ55+7nOflYELY1b
V/qPEt5Ep5WV+S8VBgtsL1fyhTToSzQxgd20YRpUv8wFGmyQ293z54DHtgXbxAaEr0Er7GtiKhXn
JqGvO8vyqzw8yV+5YAAg0SBeAFX0FDK3ITgdHLZKOXtSTTqYqBrO/lC0/RZun/M5q1Mg97FVCpjR
rJGgLZ+gjnMHgRgqJj4ShmwqzQUl0SW5iRK7tg4yL/FaIgYHBAl1WW7dmmZoE01Os98fjvtZRYB2
4qIwPbdzYDN4j4+3pcobo9r89AMTzy2A4/OAiuGZXsLVFcK+eTI4St4IseOgRBHjvfUFu+fsYea/
e3HAShi7W4cYy1/d835S8uEVdNxhTqFiOgFiu9Uxar/ugFVqHNOIshopWGEannaaZrpx7mwGSWbG
KzKJr/b2PJK87Wvtfp9ojhB+mNVTFnvsG2ZhS565jsU2KuMjxjI0RNIZxDDkQ7CxrloOHROBmcZc
z0oLE3x6Jg2ETVBloQy/V4uY/SQDkFevlQyDHUGVnehjV4O5dTV7GXyRnw6Ywpo+99al2NThSP//
yT1lXAj+4jgVRNGheJJJTMq3dZh83jo4tDJjjX6JTNw8TuMYrV3pzHuiiLqIJ/XdupTgQzQi5BJb
5b1AYI5BaD2H/h0uoaz/elbxEmrjJhpSHhvvrNUjLlsWw97HCu3cQXtjvxEpwqnbdy9CQcjiZPv5
yXz0M7aPnNI268mQcnXxYwyXpc35hxi5V+zzib1jgYbTFVyXkfIHAqPpbztWfTgoddweNePvkTb6
qABoKvwgcBh8QCkdv6LtG1krCiKD/xmlL1eWkF9XoyIpF7Av4To+SAUkYjL95/ShU0nTNe1eXbCi
goD9f3/BEW2twl036TD7etanjAYlSbmnaXOiXh9uL/PjEtenTZvYHUehGkdWVPmgU7V4DD7ogOSw
On9cFgBV+lgaFjyaZlostY8Z4xbGwaIMwwBdjU0mAOf2CnlUt6nWKlkAKZru46W7YH6M1Oy0zBUm
hoidvCrDiGmBXuJAHiG+29ykfc5+NoB02dCY7QVbD0FY6sgl4/joEt8TKeUORq3QfpQBlyo1um3d
Mvcm3njIe8NGn9Qhreu57uv8C62koa87rjBv0IyBNuwMFK11AZihQ2nF5iyy4BVnZ6+UAIQFIxoH
cf3dFGBQ2D/xiZKRHxaYUticrXuosg4R9Gd/cz1fsochjxK2aPM+cRtBk3P0L5dpOSajI7/bIJuZ
3xQmyOGcsrUmy2J2zErM2WHVFXD5XvVOdZCOiR2W2ZWfRDauA/25IE3czAn9coF6fgrrK3rcFiIG
udwJ5c7YlfntuxPP2GiK+OmYh35L3LiJI57XbqFc4EqO6YAnPY34tdPFpzjKHms0DTHe5uzKKlCJ
WfXwFD+FNEkHq6ceYOqCnPYZRlmcTrosB5WhcVF0LPlRD/sYO25K0ZIGMBlbJMSlhYYdGcFIoRz1
m2B5UZJchyi0TbnVyC9wyoIu3qC7nVR3sLhw+Xp+ZEkLKPf0ZcyfadaZQDpewJdUyoaIG+Kd1moD
bAV7sj5wfdU3yd9aAbiUCZ0hbNVAVQCqqTx1F0TDXuKxcFNgYaDUiQjVOK1fnJesS08a4OGNGNae
V0T9y5l4578EDiqa+TDQdlbywxAhWCSGnmKK+6dzzQvh66XbWxldlt5NFr/gO/1IwkSz0XonPmgG
nSxq4GXRWyVSPe0DLNPKuX19mcsjVt+yHioeWP/9o/1fdFGbsiT/Kh702TilCowWbcf/NZilX2te
b2lIf7q8d8CK/Sd+MbTTCUaQHCiE1MGSeUmI9JDEkHLMaRau/iZI0eIuR4GoY8zoWtKRH09Zo7oX
0aTAY/Wg+8luSThYZWQy+W2oGDG9UVwEN0WesXZqu/LgyLo3Zx+FlzRg2H68mF+x17Q9a7sQUN9r
aNfWWw+Do81I19opRPWVxjZ4EP6jAA+seODOtEq33VBOjrgFs9tI91Ek20Sx7Wwz1BoN4Td6ovIj
fp0maJ7qJNoCvVPd76341wAPfQ2+WQzyJYFLawuQNF72FzWTUMTFSALNLfMnYasD0fH+iDaCs9bW
gLyu3gcA43fppoQukm5gu6Mn6QHfX/hksbrw4u84M2fks6pzZ9OLo2xomiVdHDB1MGw2Tw9O0p2m
+nafHvWpQBEcHVHbpfoybCebY6qN2eQ48kHlU4rJOujfUjkQpJI70SufTGKuVneh1hrwg9+D72uD
JkGT5iwN5mvUiubKsdnGrpCSDy5+/p6QA8+qKThIcg0dTHO8f7GOp3Rd6c8aEqI6kAAYU+Ndu5J8
GRXPtQ8yk+g4lgw40TXJuOfb3C7RZFRFiHN5gbQ7MMZwcesWdbtc84qC5TnW14RDmFybMQQ8W+Bi
7XkD+faWl4G3LODrXwhXxF+r275GAZviHQB2za8DJN25AodgXKUzZqMf/L9zVGUgVN1MNAN2jdMe
QvfDoEa3BHVgJNJDFo8SnYmAKg5ptJZC2COqMudiDL1y31hLApcC5mLI/V+0HHsMMqz//tzF6G9L
J+c5ThNdl8Bw/UXtSNoYs22ozRKaT9YYzkYMBCtObBvA4dlAxrHuN6ira0wz5/K605ZWAcJmuUMn
SU4v3BeZIqeHlj2yj8uQj0OmS0lwpozhreaKWDf882NrNfV+1kVd5sSOVEnGoIrdo8tlPzrghb9B
UBtTharml31Jq35ivY4JejgX9QnLaJtpB/058YKYJWB2S9yqXqMBVv+dueLTKdo7hwq01NQKD2i+
Vm7FEqR22/N+raUUcC1q+UNi8kbdMRvsSMuVc1OdtiVaCuBWp75PxPMz3Hr40Fj2VncK3P7x1xMc
PaNgRAOEvE4MIWsmrBM8JqFBUbfQ3IiJfNYnNdxmrIh9NipQkKNm4g/7wCNn82sAJFmyoK+V5r9c
IzeXOaeKuSmUbe6IfJed36feWanMdKCY/67VUyoaI980JOxLn2qc22C93DVQpKoWXGvTjnd/Udrp
zMoqt6w6c5TIHOLWaM+ZyxLMGF6VgNyjSWI6tbh3qGTQhG0cRHoYVhGEtIMLIOKguTHpCrwgD7pn
tTGpESaUw1dGxHZNZlwRPVjfkrcHirQlaXLqEd1ZUJU8vhfVxU9gm+p3CNJ+FAbPF7vI72OXwMgI
RkB/SSYvOxiR0Z2ZMDrZRs7LXISd2ATWMjBkWLJGtxt6hGx0MyjfIcBoC4CqDLGAifSmRKkmK0/E
DlR9HgAgzZWI7GtmARFU0z74ZkVPCrc/hVVhEBq3r33L7xPjUJtuM+My5KjEUgoAs7O+fHp6xRFv
daksLLwVV2quykfotKKO/j+QJeedpZycL+QWcXJBmdvI7cgaLDLaYCaz0G5b3pmJq5sI+Sci3iUG
8TjuON0nJuWd55898e14p9DRGEXsIRywiDJvmsOqbuby0YiVaHz0hMh0GLx71ZOyfc4jgTANtAWf
N9yL5R/c+bbf1Zj7KkWWrDahnwucf3mnFgPX02JmldNMiZ+33E+vXkvxjZyJjZ6p7pxHNv6tVMgo
tD46LvJNwC7TFHsQSmnm7zd+/E/KIrxMFlEA2W8Aveqy8tvuJzG2tUJ7FQ+xIy3Am/90U0c8QwdI
KHjtxoWdYq/qlkiS8VmOlAxbcYVuiKQpoNAGFdZYOjjZjQsfKytwRzT0plgmySlvRdHomVzpTORD
91MLBIJZG6mR9MLkHXghYg6NDTWNZKtg+jUo3PB82ES9oqCD2r5dm68c/Rhe0bJP1wmGU2AWnVOf
WHV0FePLOBQ8QiLfdGLu3LkbBNhDSbPcUuYc6Sq8tKyAceKgkgVjDjfa3WVLqswatPN0m209AG8r
DEf5cmi1DKHjmUJcjVTUZyHEt5W7svp+bqboD0ALR8m+q5RAwPvOBcI1NJ0+AqeP9MSChUJjDOpE
IFmPsJpu50KwV/yicJL1LB1QAfI13DtJl2RpqxTkmU+FA7LERlwZ5xLwxEAfAqeLLdlCz7CmFI5J
sxa/sj+ElegbAIZU5oiRa4o74t05dFHkmOhxeG5kUeHefXSTsueCf8PlYaRrPoTIQxSMUaMdFikl
7qJ1kWmIhXWWf1qUcBcG07syjjJpEyrujuWITKe3qSQoHwKb8UtGvLBG4Vyz9oImIcHdmRuQenNV
00pzB8qjV5FUo9RKhNYHi/qKEOyDPC+3x0uPT0nG4kX+XgpwqTGuGPCyfXoppxp8wW6DkLnuaEGF
/4wQPqG/J9tHZer9h3RsDTL5QFA7osaZIgZJTT776k0ySvVvq5GgQGUBotpBUqoEz0X/HT+FlTXE
lyBx3kJONv0p8psYsD69tyRMJUntUpX8AF9axnzJZG6wUZnXHWJp895B7lYvY6oErBnuyut6Vl92
wVMAHZilAy7JyTf6xnSkuSbzcJI+smRAaIsS2J65bWwqTYFn6PVMJN1kkqpWn5pRXXLpWBvxoSIM
tJ37nxBld54eFNGDNR1wQYZO+u7wS9Te2GV5Lsdk4BOhUBHegM7SCTZM+TVAD2DgUCOpGBMeUyGN
m4iNm9po/Zz4v6uJzbFCtHOoHBYZaRRBxoIgQD2EEBekwr5dLTiHs+BZhmO8GwXOvYk/u53aHngt
O28X3LSqOfk4xjY0Vt2YJlLcaIepICVB/S3964REvm2/1BRb33FeEIFjxaLqWMR95Sz8e5FuTB+r
eqU2ZUqzG6uVe64PN0YdfeoONwnQ4AgECdVvuRYkSUo1XvZzie5xecwjks5hSnc7JL/0Fgp1tKVy
BCZy1p5jkmaiJMO+q86UErLnSCcIXW8aAd59uE2Vuo9ij5em3X2ytzMFK0apSim32FQZYQQ1Ucgh
R2943qsRexI5OjHD3URG9J7e+zisF/qQBXkB3sFpzH1mwB/qYybqNAzJ+pxJCo5IAoKxbFwbb/9p
TDXAZSnkTJE0a6Vy2MbpZbDSq5bX9kybciQxoM5z6zAHcLDg7E/4pBMqL6AnUdbNReYCZwlCS/lH
TKagMjg9vPDrOApaqSF2hj0z3Md7obyRv0TljzOF6m0IU2J+S3n6/koBgg3Xzu7usnbEW+OcOAxs
7AGmpugwy0mb6Zpdi++ODmH3eS17/ZfPB3H3B5sLL+WUSV6P77X0oE73odnTHEn8ucKdVi4zBz0/
QMEFdOgTnXxj8Jnb9zqFGTshCEvEHAvieempAwtnkl9xrR6sSUP7QkHsBbGneSoG/mfrVvGAfRCD
7ItPPA2jtZn3XQEUKeMgsDAeg5ar5uCmI5AXdszk2vJG92PWbmZHtwWZFy7V48rT0kua5ex3dcjU
eePY8iRkrlmdSXgY7RaqGOBfve3KU3qD1Z9VBOdIzHxYQZpNBFHMw3uiomsQAQn/fmw7v0SbmmaC
CL3HkYfFA00uzeLRy8AE1CgTftV15jeewaI+Nixi9Dn9K7qsfv3vcxOHn1VaYPU15Y3oD56jIeR0
QkaFCrW77KBKQzgUldN9XLahtKhWR6tcKJ829+J07wCpbLvPA9XxDSxLmG1EiXX9E6Y0ZJdRcuPq
1vMYzlhUKkhoVGzOGYpbkELHcg6Ezg5/YyHZG566DZwTB/EE2JwxXW5Hn4QVPosGpoFMqcrPpHar
GcfrB9fFDy4RcGP7JtaaZcGjAgUP1zgvjaLL1uWRND6bAk5RZ8cy/+JKEIinBkYQ7W7tNY05i2PY
6/JHndKLVcYflsLhdC/oQioDj9X5kVmkBsg2ykiUfn6pQ0dHae2HbeqL/9KgDI5uyzzDN8ZHA4m0
K5oCaxlPhK75PU2UmaajEWm6npwp/MUX6LBA+HQRWS1bnZsRMZdxCkNOiKoD3tugBbrr2DSVq3Ko
1OmQM0yv7UVit88ll9Q6csXKpun5eUqoy3ABxgtrWrNF/j9xqmBI/eZOHDOXARP4TflGIPadQ15h
m6Iqmu7SkE4DsG2/S88TfGOEFA90NKpveWE0QpmAiDmUx7A/7fjbSkjy+tfuwRybTnHUpRNTAjTC
3newlKhVYSasMqjoVVBQWCJBMNGB5iHw1ygyvs0KeIweT1r1sp4Hup8XkAMImEVQDx7exsxX303U
WS7LKlE/CbiC3FbTWqBxKBSsOSx3kUkZjYkPP5Xs9l6poWsfqsAqoZ57AlU7hmaPiMvTcL5i1KpT
avubLetiO5PycSJfPt6L5I6to+PYWOExxIWRJcojxkXDslne9JmKy65NRqJryclUcqWc92e3PxmJ
BLGHNczyTPiGyJjGJtCkjcGu1HLi5eajX86U1mNLNcaRUbNLXaHnNvr9m0zmTYnA6E85TImp7EO3
OHT0cVkCa9ZOeBscdEWDqkOf9/YNjSyNScVZqgT0LC2/kSRZvgzBzxf+4hc/uCXW1mLAn3oWLxCr
qZg6U8/y6AY2g1mcUjmsdZoGuTQQ79vJ2rC3amP59FAGowdy1aF1+6D5LRrjG/8dA02Ed4fCgngE
GX5Gi4ZkER3+vILRsioeOSdeO2YisncWKp1QUmdFezLXpv53vhNPw3lLxwK6f3xHLtho1lkFC7+M
ukASCKnClRuqx+RftnwyRkIDvhVRBcSp6EOPdqLXjGxW94ZLsX3TbFqa1XifcciUZETDNgrrtgFN
cO60EEXt9jFCxy7LLJd86t8x6xALPdiE70sGgAVhSswB8Tc+fNGUf40m1NQ2dtESOxYtmg/u+8+C
n2UMBqedJPSssHBqJPkZ7VQaObTN/bF7wJgeiJnLYMYMlIGDh2qsluPeBdF4rhk0Xc4lXbWR7Lgl
yXM6vLeEUy7nICvhHXbDkKwv1bMTmMkyCTW8pmGULxeZU52bVD7sBVBJFDINTznik6ao/DOq4usN
Q6Mgq3UYiinb9tOrzTfBngMlISp1utBSxgvST/pHFjEoZYocqmKnrdoEpQug6W9FyfAKh7ijPaZy
sSmCZavcZ8aJb4RR9bplCA5Yj6JLAc/QQNR+RKkvSKT/HxwKCxyiFd5j88wsHp4/JWyEMj7c4OfJ
UpC0v4oJXa5d4ome+UBgYUMn4HSFg1PKzs5hXPqOIMBKdLTR5+qUK/9XI9WbglgsByLrkprh0orK
xgDGwCdNg0tXzHKEOcaY8tRuLKdI0anKJtYTe9jEtSaa8/vwzsF7owBMR6f0Dl0eyPofbySX8pfV
/B/B1/BvOkL7D9AenGq6cTJlhDu5uMtmrIZR11Rob4QtWrYoRsXDxc/aFr/s3/ukIEGFf+Ohw6qu
+gQQjar6P9V6IgUFRzBM55ifrHyPcSR4NkiG2IaSK62WtNPl4N+nfUNX3ioj7P2Km+YW/qnopv5l
7m1gjoEu33AyukYmH1cNLtlE08ayPJ2falqzUuM+8LRc+hFy34KBOuvDnaqQJSEWzqcwXvbdFaE6
yPPkt+kKSRf66iOn4iGOgfWfoOaHqkSEsUfVGOiAeFp2xgYE1VAuYjG5Wgkv0GA9mrygo0nM+uKk
I3iHWtPtO+j6w4xs2sqixwiMkq7AxBxdDmpjUHmNsQgQ15qYkoleuZdc1VHyMVHAr0ioV63BnnXS
lhmAcbV9nt4TWtg9qdUY++gumR1a6P9UTU4saSXm2UJsrKqDI7uNSkU3jNkWRC/eIBogBK8MJ3HK
g4MNp2+uADaIE5AxS0f9HtgqUGOBW+0YX/9grrqCM7qjs5NlkECHw/S23yK6rZwyEyT33mzBcG9C
FKjsxDhhSnj4a3ha3fUzj2zhtPF3Gt19vyo1S/CZ0nqCsfcC2fd7ANlyxdUDbt5G4w47Ibnn5B5L
ZKABRRB1ZDRLigbJli/J2+g/OwikJFYjydt4qgsoQZvg7c8GK9bUdIYUC1sIwNuOgJaSDu6Rbvp3
DxjDzzIeaH1K8DlmlO4GTYDBS12VwMskP3nLELl767OxpGhwcKUlWCbuBmAMAW7hpHYvBKfitJyf
f/CmERjyv9iG9ohF05xduJ80eh0plgRZJbqE9sFGWunufMDviOnSAmzahvSSX7ZIU7gf0InUx5f9
vvLsmIKy6bOP8CWL2fqYoO848J0TjZZQz4CPkB2lCwce1u9Daol91tuSo2OG1ukaqXpqZg0yisLo
N0BxjaNQ0kr1FNeW0W4cNgtafwEO1QuZ3sHv3ouSguM40/+rK654CnkJycdp/fUNTfGE78H0fCzH
ZmnWiTurcTMNPdX2JdkxSMzF1qxIBWvCAfK6TeOZuFu0Or0w8PqANecR3zN7JmivfjMLM09NlAqG
mPhjhgoMfGZQdtS6bViD+8wcw1prwa5ujJMr5zFcjeaCiiqqC2fFXTfbrr9sCieTRU75tJZbtj7y
ktJKnqe8HoVuEzTOg8tXjSfSwkfeONFte24XunjBTUee97tGqAh9MY1M/wxF3x5lw55upD9VD1XR
MHhvNCh6B1iTPIxRN+w2hlR+CqRfKN1ZoHjSiBw1zNOVALCIBJOP1wikEgIWEYNJ3Jg1SxM3dlbc
8OFZGRMY3UclMHYYeOcNtm7DkLXZlpx4XHQO3Oei3pZH0bla8XAqzutfXl/hWUYn0/u2Y6oGJRsS
qLL9ISElnmOFxDkZyDb60UhQboL2n3ACOiC6BA/JPBMCYWiJVAELfyvaye2vClFeDDlQEfRPO26A
oyMhbie8MhMdPVwa4WgKk+RUvCGNglYdRkNT/RUUAylR4ghIH2p8eETN06CDtDV1WpZNTDSgj1qK
D3Pbj2tCypOzFv9KVgQ0DgaqPVVYQVanMpZgA3eeErzq9qD7ajte/y+lFoL70oln8kBU+JM8ftY4
uIn+GFx3GvNMN4JvE0XniNyKSfUO27ePfjqWwIR1NGqysCuAZkfCX1/tuDlklc+JOTMzo8uqHvT7
RzKkDKouKpgY1MVxU4ZrRd/9kYTzsh9gkdbNlvz4LD/GgoVCgSAAZD8L9OVfOUt9vf2Q0JWjpL7J
89rIpAg/tJuC/WdmIkW+KWcnWqllOaWo0HAT25i/s4aW2fLYpEienMePjEyO2pQZ5ukNzAR801+l
Q0STnlWPGhGOVfXcv74RV/VpUNnbXYLT0QyYvWRngUlL8NzVBA7FO7HRAPliq0Okk9K8CZgSZORs
0l36u1sgc9x3hfykKa6WWeOLr9XvbxYLpvmCAa7J0X7KeZjrZJ5YfjHebP8Jt64kKYvLdjpuqWc4
0NBkTAIPtcDw4nEnT9uUFLGf9ltQTsjaezX7+PqO2c8nJEgCcTG2oFU2SigIqc+Sjg8dVvQ1ghX/
cTU+PiYZhjHGLk73Y5N29YqPZqHvWulMoHOxDdjF4ECrR2q9DnCThSgrq47IzkSlOFIKhfXVuOO6
+UX/+wYhuk+njZ9+9EcjSju1YURqYTT+7wcrGVWpFkSaIA109gCC3xx8DT9DM5RBfxI8Wdj3/Yu4
HD74Kbnyo6cSGyjMTAlU15amTe3zq4/vBz91cVeeRTSHKCtAVT4EU3qi+HDw3CrDjEiZdau0WUP3
JT3gxgjL6zc6bzBTEefngXDqOKfmfI4bNc5SbmOXdavKE/jbToaInPurmNQQARNDCI+pgWLOgLtX
GITLnPTABE0Q+osj2yT57VFbEUgdtKQlNxsAsnE5k3aImsyMS4pyT4ofbomYD5dVh8lj4uxiL7Ay
p2Uwl/ER5/oyeOL5RPVENMaqoowkajU8T9JdESkKQIBZ6VDOA04oF0StltEt9OpLI4iOelMHEruQ
3mJ4w2TENIw/pR91snIKMvM/4W1AHsvHhSANB+2zc6Jrp6cG8bWzb1oNpKkxd0ulai/WWE+Odjur
7jKQPe6e8GZowSmULZc4w6VF/P+rLUOeIOXpx5KfGm9kijRsIGl66v8WC5fjYv1XcDEGqbRbMUPy
HyIXzUCDf2VLlsRMViJe1BuGXCZC7ScSsswlQi/wevEMhC1tJXLh1MEkTnWMklqf4e2QCn41pImt
uh5rQhf/XLQAsK83iUk5VgVcRCrbHbg+0S43eez0tIn9u3ibv3IsxPzb2BUglmbbTdXrc3vcXqwr
msh6v0fdhiMERLwz2uUaNHa41TQeX5d0E69PfZg2U/4lIChz979gpTm31PSIa4gWHi4qgtoSJ+lY
z4ZEEU9ikV6vNsp6syB7jLpsJObKE4kbnpIIjF0pG2mQ/H7bIhEC6hBNWAM9UhyZQ/tUq7S68R9W
6ze4KGOgaLC3ex6qIvp7LgPrE8xMUpEIzwAPra0Q3jPjxXUgx6oRGhBUly+sr7CwXxVZH/H5M3ej
FrV0rJYXjXozRC/sBooGqsvOJM8hJrqfRVrRbsi/CZ6p5ZImavhj2bMChOMQ7uZ7twsLw+3JQmWU
nGbpY6jqtd+plVyP8THF6rSN//bcmE76GbDNjLjHjnnPO0rYyLOJpX/HFDBR3RLsBMspwHWt7zDG
qNYpOrQVx3mHvtMIASOYpI4hdQPdHqmvXnTJrIgIcWpzRAAvaKuf3x1Uk8ZpYEadIg3cfp+uv+Tm
Jk82SZ64JXbzr4s2/9AqdwcEH8C524rwrJe8pJavWfIHHlp9WAUsX6GVO1Q+Z4+EjxuwGKKW/f/u
qjIqsTA9QhuvJqiNLIgQqJWrjczrb5g0bel4uuYjOE3Cl7RbpKNsRHziO4cRZo0+s3i/20UPHfeS
KlgyWIT7LeuFeBKMVY9kW5mOP4p1G1ti9xdCkbqRz/VcCM0UF07E7pxTRALwinFHxRwnKOouZwOL
ys39Ed2GXsHMolyOV+dkArqzATbLZhVDUgdS/h3JRsFQmVBrmPPMBGQvf4y37rHTf8oLFz2UBspV
Lio+KfaYzLhx2I+bvz7KX7sg2KHb2k5Af2enrXzvk8AWANf70KYdIl62tnRTff5AHvsxYTZOjfeJ
Bz9oIcZZG1GicRR3zkef8zm+MT/kheJydWjlhoIG6cwtZmVqlTOslMhZd2N/NAMtGTCboanyVnjD
WlMSbBerKz1Sh5Uo7GDakHBzgyXNtoNALU1Hn6EWyQ4J9xmFyeEDEWNcIN7s5sce49dkZWjk7IZq
KYp4oMAOTkYKTgS4Ug5PoZeGkP+73g7KSUuwURKHPYNtzze6O7wAELLPmv5uVU73xh9Us8ZlV/jl
Y26MQsBTA5UawLNO14dAyTTt0r3XhfWlD6N1TV5neGTeO6MOMlBq38xddrJC0y1k5SMkGTr9ZbtI
uMmgiHOk5l9VJBU1CLJJmwqQ1cyfWpd9Ykf1/WcrUCdUQGr5ii8xvmA6CaPa7lXlvXK/bDHgcI7B
nieLsNL/CblX49x1s8zMFojd+e7MB1uEnAC8BKZ2ytf2hNyah2RHPmado+tD2RIQvsgjBpFUGLcZ
5UPOgMHXFeIMxApTkitx4bStJWg0XJf9AEm7DYINuYjUir6NIcGXTlREhLc70yOR7v/s7IXon3UJ
o/q91E4e/y0FE43BjMqF+vMkug1HoD3l9a7N+C0MpoG+JRGHUswcBHI1429tr34cQ9e3qr5+90fg
D9vT0MgWyB6Y04ED0pVQDLTM7R1X62LyBzgG42/NPCZdj3zjjUM2bn8F50jCfSlQLBEaDdiMYl3I
4Or0Vf6OGGiM6GL2XCD0IGEKcphrxM7Qx/mvRjM22bmPwgPB/cQnuFRB4zQlZR5Edxk7yIy6WGls
lU09ADaZa/otlYHOn+mwEy+y8rsYhUwf06uG3CJwP5hbEuKGUBezyUTgWnc9URNnewo2kqTcGFaR
NDPK9n9iTc0IKg6ttww+u8jZSuilHb7MI3z0FY+qem9/qS6/E8NUp86M5kBa/ay+76skuWRGO4YG
veCmCPAdj98rK8lmVxNtAoFbnRMUMu5ZVQFD6o0RmThtBBdvfEifX1l41VAL7Go6hUZwrHl/kPPV
wu47O7e4VO6xyPbSpOnP0J64h07PFosypJ63jVqp7HM4kTAgB1QiBt7Hv0qu69V4yWpNUGdoGQbD
fztvmw66WNYmUGdJUTn0x9qoTk8lplVFZt/KMy1L7xluisFugWmbtnimh981p7FS2CgkZswEe1S/
DVHE2WW9DUeKr+lfVCE409U1b8C00rSUf3gBfAmFvxJQal4sjl8LIKi39uZ4I/4qAbVqHersrexq
Pie2ZWzfebIGy2Fj4H+unJIwHZS42MG5ACOHBUjCOr4GymCm0NSp4JCkYyitN0mg/pVdF4uUSDpo
NxHDhSARTCJyMMDTXe7/ug9Mhd3oqNfjoyYyMjKhW3AV+uHZNgMdTKlYfRkoL/2Lvo1v0F0nMn3r
302eTbOBDR7C9v4pE+Cvs7g7EZ/aId1O+hq1uxYBUi7lhokrz0iYTvBAiC1YLl3jhtjtxFcA2ICL
P1Whj7KmnzpyvrFWZK71HOBO1MeERyMtINemfbp2q14Mwt3mbcbreRyw0xVMjIVwipWn1gcE1MuR
yeu+wRG47zVmT4xwTvwhMegVn/clu5bi212TpfxYYtebWbCwh6hpBkGXYeWGR4LcCn91RmgQInRf
bC9PC1fVRJ2uHYe23KVTKtJRNVqxvwuJaoY7llRjDhjGqIxGYbJP7LMvga7gcMkekbFEsnq2Btpr
QjxpPllCfccejoctk4ItLmZ5eW8Agb7SMnAJ+WU0NSiXBxZZQDL4nZRNI7sQqE3Gh+3WcjYK4PXp
RRsWr9cQSW9X7H+3XCYWCEh+QtmKCDcwLEPcOVnuKUjqBQmXSqyQulvuqSAQhXRACunqqOmiwg3m
iiNJaZbub8TRgRyew9Z3uR4958ngHlranlH012H0TWBIAnRvI4Oex0C2i659M1+/D2BdUk4Xya9T
6699aVtayKjWEaMuYr9kcy0HCd33KJ/+9fneXV8YX9FfZVfrBfVIpldA+JIjn/lSSYpZj//xhDxq
PUVMOi/MuXvOgGONRA4aVLUhuMjh9DIRDElQINZZv4dm0mAKM9UGmtKFH3+4ZgCQWILdd5No1+9A
LMYznoAyt6ZNS5Vz0xOsQ1rHy6msiJ5x3lOYvPJwiOUpxJZzNDUetWyyK1rDSjzCAmELUdjGI/VW
UgTAxJT8dTJhbb5fZ8Xpek9e4M3n6Vut84A9bP3XRLnbhN6ShiYrwpKfq89pDftY4xOpu5KCyaWD
X9dLbGTX1SmD6OVZSFiK5/65RJzL3hzfS9E4K/ERc9vUBqt3TorJc1W2MWUzXQV/bMl/umnMPt1y
U9/62/YikDO+Nuh1ExGIJl9G0RienID6/CPYAtPRwzyS18dnQIXsi8CCpPkE70cuJyhb6wI4pP0O
dFFa4LeDL4/08oFHIxwvryJaCGKINWal5XGoPb7/IaEWI9VC9mAnEJEKc8PLEjpC3Bo6FaAbhQkC
Z066YXsu/76mJO7QowZliBGg92XCfblaU35rsr4h6Auf3JP7yt4hG/x8zalmsdNP8RJXFU9ldUO3
nljWxaILwwzqFdgk4BFSBavzI0Mtxzq/nn5Fwatq5XluByCUSwF+F+/Tdef8bzJjUBC9A0bub7kZ
NzdGfXZ2JUd17zYzhh9bbitFZBk0h5WWo7RTzuzYwPSsJs2/NwgcwejFJtebo2cElFjgtWfS0jFc
esirLUb3Eig4DrYk1GFpNUuTofsfjf4CsJkRivL0qmdeewSppAYChDcxolY9msKYTgU+BYlqr+kQ
OLvMQ1vI06VVWEkId84aBC0jLs5PJ+tlyvjwtTA8JOPJp1+in1g6jKPWLhpry6l055R4nwMQzczd
Rotu4TFE6MLylBZumKcF1RH/BpuebgLwgAR4u0R4obPsxRLSo2ty7wWMVJgqKZiAc5seYOYhiGAC
WgydjvHFukD91zVj8ave7qvLXRX2uFwe+7Le7C0mgvwLNisLegBSf0qs7YH9ND3IUfVv+jVcnxR9
iUFc766dJ3MqfLP4G88ztzcuKg0fF9c18rT8CaGzsOtnnQ0O34tRPKsz/DQBcsHD/WANB3npnBu+
ie39RiYZxz7UJC68sY7Kip4L4ShSxpfYov53Hy0I7Fz8JeIsYsMzvLpkzOY2lLLfx6suBuAQHICZ
sTZJg5rrUkQF/k7elLX98VBBBDAfU6QDwjWjafM8IxLgqlvMTc67wGqgPu/qb80930Pf+T3Q8HFm
Z7QtKwSlfSeXGgio2piWctGTl8i73wxAjhRPo/7hiRd/vpwVWxjVEKkb3B244313EA08UlRHtFIc
5gktflSRQEoWKFai/dGfPlFA91M7fcpUANmTS6zAg7VHuJaXAgOytmt2jZS8MRxGcXjHnVmKbyYt
q0Js/v1r8W1uSJ6w87Qs5a0Rxoesd5hFfdo7V1k8hWFmx2mp2fw+lSHEaIyv+k4NRtdgYlB6+fXn
IhbBUBH9kKhH7WJqbnjMdN8WPVMXVKXZoOIw5dWIYayf4Q0ATA7kE5Wu0LGPwGlkohmnna/zArXc
ElRXurEmhStNCH0IKxFOaQKRS6cCBW9ezWnSMQ/6FmN/tXGpLTlQJz8PxLsob76kcQGeEPyUXhg6
IC+k/4ICoqQ9RXiCv8609CF2/bg5RamSVSNMRJYztqzUGRXTNrso7SXKlMn8Wk0FJjzG1BN3di6q
WvY+RYx43/bh7aDtfGbC+QeQKQTFV1vMSpsryA1kuwOrpDdyvhfuXX8vtTf3cke7MJMmkMnzVbY6
QwelNZPQDD66YCu/vf/Or8z9NrMu4sXko23gnaeL7Dxu3RcUsK2D9P5kNsncWXMIL9FXnkgvDXj8
Ru7tIW5si6rptYkPYvVby8KVwRbl3rOffwRe75nTbge9EN01/Sed2BKFJqOyqBdKE8fz1dRLGGag
RGaSWn79qtsUWpayfNR0ukLpoKd3g8W/UlaWPtYtcwLBGN+xsMj3hFF9iVmIRfGI/h06NWGFjZ3A
Q0GVTEGX9p4oeDqaaqaTTh2r0g3w1s2zqHGlRb+OUhWaK4hTGcH5sPM2YQ6ny1cmPIRIoeicr0a/
RKtnU5raSNyEdgTJinLHP1qOnvVoTqAcqufx46PJ0BQNFUTo9JUVQATDa4r1ToEpAYOFdAYB/xAK
rj83fsPMlv1VHYdCLUPPXVag7rozaW7iKLHCUEp3XDFbKcGju6VwNa5Czb47PJPW1bmB9feFYRqF
V12shYCtIFEdFEt7E/dKfUOAw7H0FjG9C+NZnibLbsuUnOH2iNuZcEbRT6GcyUhayD7Gl7qgkA7G
I9xnwSn++29pSxgaDmBK8zlg6jv3EfKFA/InGQiaHRzVUVZBJBaFaZcnX4MEi5Hs1mC4oADN2jtM
SdeZexeTlBlshz28BH/v2viEr1BrbpgqaNJRcMmUuFpheP0fLfBsYqDr+rPTW7ewqQ67Zl0m5Qhd
Db2XHzqikfb0cGOEqpMueZbf1xIdhVIaw9tnmfNCAcAmSa43evgrFlhJgftG6gAjehU0zZoMXV7y
OsmEkr1QoYlHieJw3vEG6xo1NF3067KSa8YQc422FkdlGe+k2w+0fyy4qSSO+dKnMrHqP+rjO6x6
nInlgwkFQvlva5f3/nhP20e+qCLYavCyxHK4JAPstJtgUifoWUYNk1lcgDrsKfV6kC5BzxDJHV/C
sLYtL4o8pq2mEAoaov95D/A/T4MvVXyafHdGXdU5r3rEcyldujBGOfFGcx8DzwZyUTDhQNaW+0jU
TQtJOhKb2BzW0zHzD2dXgSrBIyZ6vfVMbyVJPLyUbwgAGXxq6NCNU9fRoyX7oeT7HNXkKe21gfe6
oom1867YTQUlcXzG17kt+sPByegpA/oPHbYY1UzIqAqxThthLHnPU10B5vvGKXZ/rBI9DJMQIOXV
HmBvXY6wEUyR8I0b/lJo9OVtfyDtkuvYhdLcQT81VUAE/iE9qoetY7AR9O3dN6sb/1J9A8DzqK7b
6sL5Tt2nucr1qHbl4ekOd6sR/JMyM9lab3tufgreinUQDq3JqRCGWm0s1b4hctwAkBhKwz1VA+Zq
VrlED6OEbbiUzkhIlDEYaYWmbl7PWCRVcEVYwzcOeRT5DdkefwGt76F7FHI9muRRAKd1WBp/6Asb
fZyz5wO1cek3mFBgw0gT1UEmw904xPQUPbjzSHbBLSLTseoaPYjOlw/LbZIY32XSYLkeaPGca0bw
thMeB4UC1q0JxBITCBHEWsB3feUufrbETgDA+IkmgTiEtqnciEUD0zrBjWMKEu4yD76czBvn992x
ZJxfkIACHqJLeWrOGgpNaunj6Kdw2Z+ZGHTiqxg5Dc+TsCZR6z+iXKEfnVB4/tTgMebZV7Z3GH6q
96V2C9LoaBDcpsR6pzcI6K7MKe6WGGZdNzX8OHDERA+OOWUN8yul5cvLQLNhxIdsMxC1cQM1oi3l
m6vbp1Cn7iYBF8oVolqQiHNoGu131QQqno5wZHNO//zrrfn7kI6lQFGHz2i7GA9lV/FR9Fq8tJ4Y
C6ZYjmZYCjzu01mvqgWukKG3YK5hnrRMtDNAFkx3WBJJmbuXDE6bRnQKIw8hcFunFY3PSELnWdjy
Yxzz8WYUIMKjtA97wl2HScTlQeTQslHeCBfLxLIxbMdBelCo7EKYPb3GYby4eJK1CK37DkMOLpiW
Wms2fH75Fub4EEs7azPxZ2SSXaF15RQBi50bcrMXD4mlG83uTs/a5KKrxxAg1hu/HWsa67zEYPoz
Wc0srMc18rienf5rqXthwfuKP4PMlpYC/wsG53gCeGXCJ2wCPobv8m8Jdb+KZ675reN8F+n6MHD/
KJeiaM9Gfzk3hY7Gs5r5qPe/9zsbAU8NpKRMzWI3hWoLJiuNbnyWruibOJcn2Jzk8A9xhfreAwYv
FYdvDMpS5fwAWxiBoZtcBi2Yf3zVoisklYy9PvDcshycMIBVicn7zG5jR6xO1QZXSEl8A4CtIaVr
bGqk8PN4OykfxFUrFtslcXFZKA19y7Za1cCq4bTKIqoxii4bkwzl3oarqokusWqXxg9C3Oq/48hS
y+TvktYzaJJEiGem8xfakuzIUf2kazaw1IIIfAPQ5tp4ZEY+jzpCwO781fLJupJOEeDZfHlh2hsQ
2XI60SdDepMl5+oFn8zzH1C+0J9q4vjGQfS16LSFBRaTE1IkaYnHHReA/wGcNEN7xLxz2fdY9kNL
bLjUiGmEMCqbHUcYnC5kSmkfjLHQNRhNPCzfe6Rg4rJsYNaAGdpOJKbFaQpPRZEq1aGR+sQKWEMu
wXfPOWFy4AaFJQWjkzl7TbumowoAjh0XZUS4fS1fd0wWQa5VKicYxB5LP/PV9V+w2dr0iN61KBMR
9scJe3Fv8fngHEbcx1AGnPbUB5dafkgcosUUb80RHdGDagQyBBRYFcGzt4kvHSaE8zOd6Dsu+48l
OR0a6wh0OzNeMyJFr7FGPxcy9ucVCkviLYZ/hS9cYaMaws/PQJRctz9FfExfPSEQPQQfkqAKfFyn
By8B2JO55YomgXBcfK08XUmDIwLMxJ+pL5N8kNd8PFTKRsAAZ9avH0pYKqhhl40gtnoZkstNkHpl
baYu5zUgcd9I8kX3INQSdnmsjT+568jsoGFMY3s6rRvqtZxcD/DJgDDIXXmtSykycQz0xc9czwe0
US5Jyd7CdEfxSnc5wuW3A2MJw1umiBJXYFvIwEachSDU4O/k2IVGaxfS3cTahq+mGesH6nE+9zU0
KIIvLdQguwSQOzwZaiiEf/2ia4t1f+VbfVQcK3OZYGBkX7v8mH39yUeUVpHFJNjnsAkhWv0lUUCa
5TlDKqJcVRJwxpqOaJ4V8MsZayJcPVDe2Al5Xav5ze/jHshB/hB0yvHf1iXukTT9l10+Ttfm3SRy
J1fZTL0iiCU/wRShFN2jB2IptWTh5aqpE8gk8jtX4D/VkO/wnRehFFRyV5/B+5k32QGaBMFEaRBt
W2xu+8Jal7ul+e/beQXly7jezwHJUGnCFCSi6hca7VPrnpXVsVIMlBC5DKSHW0TZdzNQyF9iFev5
yeRR/3P1iVhoJzbs1h4TbzjmJry4dgNFcl2BFz3Q+hVBXu76WCW8WVepJB6shIOK/jUhnZ0IKpJ1
GTOycLEkheaBptJWujr6fCeEiQZpXeWad9bx9OzSo1GhGJAf5nwz6eLhK5LdSs4o8UcsEgPY95MA
+0WYGfUZWFT6IAc+3y6l1gD1AbegB3mgV2TSc2d0Za12dJxH+nxOPJJ6yw4CqdKnDvJDqmc1yqjl
v8U1ORQqN/DUKw2FgD2/ZeyJX1YiprBwZyBZ0qJTGGSTbHvU4YciiVcIxOsRV6Ul6RtQzNK/DiyU
PdJr+P9JGqjFJGlaenFEaFLAfKG/kU011/+MfnDKlZmgLZ1YJLFXBjEzh0iXlZ+TrDtqOLxyQe4S
G/dUToLL6OE77krH6dNUk2P0MGEl6bx224387ipXpPGhtev+LP0jHk8t+KDxcNGRdaTVQdosqKHt
rJbjZNPfhpJvJEtz5nq6R5Gyz0eLAYNvVaFhmiCOgEw3r2Fxf51st7izbF0nlFMgTKhlJghjayze
WVLDU/EO/rrxicZ7ay6/kxQUTT1It6SilaoLI/GWmo+paFc4dLMvB1U6Erq21DztOGoMUhFa6pYb
wUz/Wlm+OGl50QZ3hwLhghA/8SeH3pVgxu04MqMPr8MmaZciv1nhsR1HTES/t3CHR6SM7D2e08oG
vXIAa6MZ9wlIRRxy5lYXA/3yhXlwkFcLiTxjWPBAnjMwsn8LIFm5gLDaG7K11Putm7q2vCt7HteO
/PAD9E6vum90bjoDb46jPU6DubaQR++XGUOyg3p7Eo0RXNNkgqnshyr6YkCjkuQOTx1qUsVX5a69
dN3numRL9jtX/TwXKqCKGjE3QsS0Pk3igAok1SK/P04t1Sazb9WpircHd8vXVJJQcrKJYDEIR7ET
P9DE0YFafwPX+gTFxxIennNMKtnrHzBTEvyBovCsuoRgk0H9VcfjjDPNkBZgAtKymktoYiuPzKvx
iPLvgeR/uLQH/ojl2IUbGnWH3Nx07PJ9dvxAJd3iQxiuc+KXCxNn5unLoteWkriYZLNSmH+eVkxq
WPblHmQqCOQmppYzB8dkuz+a4crAUlASYVdV+OU0JOX/AReiwRlrMaEtcZFBlLgKDQjVdf5BBPeT
j8q/gkOcA3B0jStZ5+e4ZGp0UBQ0rCUed+EMIXRJG0Ga5XXltvylSiswaXrKTHIeA9qlG4Opk9UW
ha50NKA57RirxvwJ37L7OyyEW78sj9I6L3kv4EHDFTD/hsCC+jBeg8GLXLJCBZn/4SOLH3HLWp05
of6pR9uP7aW4nOPo86PutWh98bXEdNDxpsinWd9Y5+yjJ04TBhfPteLVZoRqOFxJ2eIRtK391Yr7
WZkBMP8znD+zUl7Esk9qrCrlxS4B7GQHRA3tEy5IMIuab3/lf46ds02q9iCt1rQPmzpVJ1ddpDa5
MvNCL53HTKBPZ2l0GxImpxnYTCgZyiiJy2xI/oTmPWwwoSNkLdt2qqtZrVIgoR/Da0xq6bdsFtgS
2tdxKiASgII47ZYpLFqhD9nePOyO9rFVnJeoA+geTrfkldatcUkxHzLX3Ud/ahGS+/bIntKZqGSz
10N8cFHvwI3CHb7Zn/znHwrRnZ0fFReFHP8S9EgxVaJAs7yOwZShdzYKfacA0w/MioPvT/DyDgDg
RQgjmmzmGWieLqcUFW9coWJIgBLUlJdrIlHSfgo4Fy3MPcI0ZwstlP0+r8H1alhoB2ShUeiq8jJq
fKen0/IMsyiJtjUWG4KmKbPBok3pn3goCQTrINUZLBRY9TjklhACoSa03qO3c2mnIU5+yZY6/RoP
OG9oyIHdYlvEjQQbVcjI9UqDTZFXxcyBPpGqQu6o793oN001cosuJcqz3KqMh5DQjDyDb7050jEU
ZVxbW6lvObtU42g67oCN22rfO4Ev4+2rCS7TsxA15F8z9cCEqJr/YycxqGMIUZ8HXWDWoXXNcxe2
t0Nm2yzwcOHUNVDCET+KVSwpNNPBdMmg7EaxOdkp+QX/2SOXqFE+HsBHsyVIn9RDL6CN4wLUBy2o
7j+EPUIkka1ko+qd0XH+y0ryF5GhBUP/bil6su/3UdJ0IefYg05oTSDqzjqKVS9oso51PFvf+5EF
jn07LR/+WRys9aXrcI5+il8YFvyCEYeP2m/y3igfla/VRHe5SVqaGOd65020vb02kL6thwQhEkEi
uLO5JoCOHe/8914MCkMS0hnAHeuU2/ulrhP+9blHsXWnkzJx+FoTPHDZcjzV7fsPQ0UWxu8ov16i
fBxjvwME2YZYr4jaes5VjeCg81FNU2D+O8zYUhsTCSHsOHSMI6pd29XcenrX8Tc1WhOwHfXWdDhz
ft2aMb8cUliMSNC0Tldkh5SO2Yaq6bVEjLIbqNgkxVNxFiVZUe459iFn0lvULqUOjztoW8V/3Z1X
43GfFbMf8d/Ho2noXssROygePDY6CwX5Z5qgCxl6dprSIcKJJRr4dXBkgUwA7ZM6CR0m03DwByln
4Kml49+OmalWezsBIJyKhtYi18UK2956IYwnCrCi2/U8ptZHLtGBr7fjYfjON+w/bA4Xq5JgTdv/
vfIUkLVpW2gafzhhWBGu+JW8NKiHdvWVENZOHtlPA0ooSavWGrDdSlbjf2a0q0Cy4CrlboADN6kS
t6dTfLrcrT77vCQpbesIuegcjTFGBN7zA+6CR1x0pAG+MLgXZhvmST2FJ9WfdNRnOgKZps2bjW5X
cYBXrLaZxuiKOCcq3hngHryZVWG9J5WzJFpSP9+uCaNcE2UGBjUx1WZ5Ij8Tx5+Y2yh6l5NoXm2j
QyzjtL5jKXE6cfF42S6RXnzN3Zn1MXgFF0oxXCXeP+1GtR0MfzSBON8EOgl/z0jt96u7JUrESdwU
PYtV1vCrHAfh0iQWkza2C2hYf137zqLycYy9fcBmJBJ9TkGD0lbxm7mriGVHkG1xzAOMbBslFG/4
f/aqgbKe/PCei9hwp+MYKljJCr8u5mUCIlyI/kRaziA3QS+eEv/z5aKwZ0ZXAde96Njt0a0AWzzv
UoKXvUz8Mq0YXuAfRiNjFjgFyyZkcx3xKbqbRVmiHX3jS6e1lRkJ9zChcyQCx6VX60Md8PCR+y4K
eR0vs1G9woGcCsrrLcyuKVXAtcBKiBx6Nq22WyOFc9Im3kLQUGbu/RAEAIghn8nGyToKkGjDf4ss
uRa9eKEy20kdBIXtE42QiHe5u0/i3NOgibs8zN6pt8zgTS1N0EuogCVS4ACCGKITSXFiR5RYz5+4
bTtQN9B5BKO9diXHPxBgZcwxvtoYIAtHqwVPl7tDCraILeYN1byIfxDCcBIHYTNAfvQUJ7/Iy1hr
u31vj+Eda6rxqqLbWzDswoZbY1UCuKca2AIfMq1GEHwbOIIum+hH2b4yzXQaH/yPM2IH4DmffLrZ
3Zyk4f0jeva8Cjb8qy0hj7M1YtOkalcLLUiMzftok8+U5aRH6HqUwELIgOHF4EcOe0TlrByjqnly
wZmOB3bYsyTolWOum4D4KUIZ84x53WF93oQb8d7oqmokdG0ySxaL3MK6+A7W3w6SuGoycV9Dj5Sy
xzc275mr1xgh3jD8y34ZTM4JK8oJIL4FVnKMlVEVpykSIf197ieHJl1J5CCjbonXaDaIlMJbG0Lb
qqrxcYTSKQtQJzVyQYZ9uZsJGRU5edsypBdEyUjsi4q4QL9x9KhsX3xv+A6R3C77DNhEaM7GqZIU
/JBxqiFla7uIUwq1RYV4UcmeNgMd7jtnnL2cmpvfITgGCtK2NlKboroZLQ1xkz78nDVlpT89DPfI
0mwU+v2FPw9LAk0V1p02pFY7TPRwbqGwjSFtjXiEIlqpABi4AbRkC7ec1TtMmrf5NUWMCDuoi5EL
KLoS+nAU60lItXkHRr+ihuzrgfC4yXFT79C+WjrqvXaS5sSbtVkDQaCWLwevpBymRSris1G33MdV
Wkgou9hyGYc90kGTkPti+9MnVl+Oa+Oc4aOBkbXmXWz7RbtjW7ZJvPfkbae7lzbO1h1CxMQSmmWl
k8T4Dd/bObtjAXRwUxx4UXKr6ZinDbToI8/UpgNGm44xyjw+VGVbLjckOjXRQf+96PsSZDmc+3J7
QxEfySx5OsSLWZM4LD9Fo7B+NHCVJ7JU5c4auh0m/hozXv8pXn/uC4VbhHmd+POCkKjtaryl9yu+
vcfv5YHkjthG5ozL0sD2b/H2OPpGBybIksGlsI/OwWy6hOVKbfkQkEgCrP01QGpFGbHKchq7gZlf
b6zFeNz26Fdo/GcEkbUSetMgKwir+46R6eGpT8OKGOr9SO1S/z8dg4/ydR75KDJdBmGMsV3bZQBm
D6aKRjsFo5VXy3cVqdeH5Z4vE9gvmpXnkTPmR6tkc/KHUQqO6YeaG5zGE27yQ0BkJ2nSZhzGNkYp
2q4432aIWm5hNvaNkFXkp2p03mcMJGUtCn3pL2RI0gWgSOU1xqCAheRjcasSE0XZEJ2NkUvqOzVf
gdwYjtpkP8T4OauySCK3bMC5iYuwcouiV8s3QITkVBOmgZU9oUiuaybGhIuzrFi1mMIFIu6x96bN
uyonkeMhdodwUB2SmdqdPzImbk7VLqifvNV86UmbsPgZvsOJSUsr9DNQmQU5cBpJP+yXRikaqzZS
jBTipEEZ/yc0S6dtSf8BOiUibNcUhLDGvX832tTUOjkh/zUv/Ei8WXjnSp7j+yZ2Qo68bK2/15x1
dXkxhJfzbE9pywBZ1vnLUB5x7wxNTbz5XW493E3AiqbXh5G15f+wduso7aq/kSCEP53W48ZIs1GD
BuPK6IxUaeUvFGDSNfLFuWiZYLKm9BQVadCLOwkfrNpMDGSUpE5w6M/RIYvygEbmrMrl3p3EMn2e
oMBdGLzQG4RQbkQil17AvG+poresziHhFKk4jAmHhE6aUF8OsCl5bov1RysBAvgoWstnJNZfbt6H
vHvpoiqBIWlYsNviOH7ISPGrDnCbz7COCaff+gP1BhezogM0lMPCM0AhzZzp+JMX+x6/9oDbCKXp
Bd+n292B51agBTO/DLchNwOFXdVvAmUABmO4vtjprdNJ2GU3VIOhuS8gUAm1mKOIJIDRzUcM5e+e
qwWFQ+No5dRSBJ0J8Jl75KSkIngTDtcZDA6EvH2dbHog6B6sqqeEETxIa0IxGYjNPxGbJ9mEE5ld
aOFouD29HPIiQTIziqTP8xE3allHyNe3CsfMHveyluWCbgyYV5paAmRCgGoxvae+m6iu1M242d0a
n+Y3qZhzGdULBrYZ4YuDsp3axf079aV91Fly4m1coMdZm+87IcBAWHFBWutMhCyaVxCHVcaL4wQy
+fqCoFxDiR43NsAKKT6wOIX2WOVKhWQAhV3xhDk7Y0XCwPowU9IHNKfvncjH+7d7eGDmB9WfTQjo
I5rq0O5b3cOvl6vA0HXFVYGrwzyFla0jGvk2Xh5iiLowdkUzzu4wUoYMrUdTe68MIDkcwyrNa7ut
hznuYg1WiTnNWGXWrj4vfM5W1CAIqS2ozwzOlcIrBdgGHt/Rp1vnqIAStFTmwgQEK8FeJyJNyZhf
PmOqyjZxSkQHKUNJnQC6uLp1bmOh3kBFBAPj2qPE0NYvk3kn+DaQ2TiQe66rkkbF3jXaSwPC8ZZM
CUXBZiFQjm2zK11HnySUgGvKHOMW7HAY/gxoV204NH9q9X+CuG1QMMAFXFK1Eg3B7ZGxJGe92qFd
MNdYUjnnsYC4yq3yh/QK/ha0dbgt6qabYgo6qVnRguTMYTb1fU9Ba3JInJgFXvysfN+gwgY0IVcv
iZbj2jj9G6j5G7JpdvdeR94304nGjQVU5uxWSLZjtVqLNh0t38YGV5Db4dopLjoYJa3pEOcdwyex
iGFYxHuxdc+ZLEo03XcZEY84Qz3HRpooOOm6nQ4Yw2QNtJL9yyjQEKQb/hYeK4M8Oiq07meMflby
O79BzZDcSEeuFj6kS0zoq5Te77xHV5hfoQOeQSabEUFQoCgNsfyROhLk9L9+xJ/rpIptYE8GH4OO
WUGBmf/YPiISbz794zC5i4uIwC1fV1i7K06inf0YOZV9iQLutwG3vPUzHxuXpzUVuItxonXm3ErB
qj5Iof9MeNEYP62v+s9frqacI1ErL8KgRIpoqdot2mYS4eBFwtq/yzxrjGmADhe6zqzh3YUQ82te
iYtc5qKVq03WfomTboIFvBoNKe8zVPgajkPFx8cGQ6EeF7doup754fOf6DKlnF2eVTF7Kqo3Ik6Z
zFjvLByqy3h7rQt8UJShYImNoQjxKaZ2Z90mub0buGwgEYiXeAQheFDnjcnBvZWftF4NJlbEsXxr
n4v8MEgm+EhQGHSEloZFSxNmRdWbSvJL77hIWIHVDm/BkKvBkg9xe6vivkFgqgnWTmzWOuY1a9Yo
5x/Ly+O7J2Fjlh+ZeZxYS0lv4PA2eTwFMAfRktGdAmcEizzLdGbNc/OSqwP4pL6ibWTD2Tlcl2D5
f824Azs6zOZodcACgKv7TmkPIoqxlI1imazeuTZzn+dpboIiUkfi14pLDg1Q7JZO6+lD0KZhUfPF
Hd/GT9c4/xALdgEnz5VmMVTAlhh/nw+KM5wqYlGiNAjzWuxWf40O100h16nAsi5nICIroouwYTRu
fyqdTUE9rYVBTGT0wvtveuCW5SijcjCd5/HPbZkFOoVtm3xB79dfQy6A3k1P8YI9dZW7CbKMGqm9
AP3Bls/oGdu3br/QdIlv3FZ/pAdidgiZu0I1l4EzSz1A2EnBFVAFrYu0AkGZ8NG1+pKMW9Wa2bop
rhI6SCqw+xx/KgVCsVOv1JIr2OyzDBuJzpr/v/Z2/9WdVsL+fteCRqG/RFX2zhaLCx28at1trqKW
L3SgeXdCXS/PtnnhuOciaKVBKvaXWXsR3pANYMbT3/ULxjzrMkbs4oZVonVk0aXlkWIklPfBkE5r
p7W2kjkUBUFh6aucB/IPnBGpBXdMkCxyJ/2SIyGFR0W5hjab4+zh2szdWtsUQ5ugUi0sBcbaPfJ7
pwN7/60K3oWOAspW2koOpg9aiyz7cv+9ro/UDiJagMnsQi2ZcOVkFtucn6E+XAKYqVLtFf1HR2o0
KEpWSX5p9qn4AQ1f01jDNBEHmxU1vSqbhJpPYcGHtdchlA763EUT4UevrRLhsDRC+EpxPnmcaX+S
wlOXLV1hUwIS8HY1ce8KAdiF3A24QGkGvijucNcrnq4x1577z2pvdCcRnobsQSxrs1e6fFolnFJA
YdjYtdaZ7Gw67c20TaABkq7zqrVgLCvUw4jeEgtD/EuDzUY9o0dy/bcvEk1OA/PnbdLaa6BeZUkB
U+Hrxw9tBf+O1JdNiGcMBHy+4myP4xfJgx7IWOvm45SQL43lbu35ZDGLlc0AJ7QT8LVoOXljTXyo
ICmDFhuWyu91QpvgtKCHl+HBoa30ksp8wOP7lfkyGQuv826G2IzvDrYnJqQ7lR/CY2mc//syXUuA
jZ1IeU28DIgZDzHAii/2xyCMdFOvKcPgqhup3eHduf3icdtgA7vl9jdNvfiIFh2n8RV7/RNcdTEN
S0NGAJRP9Yd537wZtmamzu02Q9QIoFdA+QN2GUaIkneUZQ/YIKejEv9THsmawyqRd6RSeRe7647z
Jg8FEGX9Tz57ffWy8sCOvpQ6IUpU83ESq2/8RBDKdgDmTAzf27jMcBgBgyqGxKzhvZWERfI8oG9r
hi+jWNB9YVT+J0+s6/a37/rEKQjQwOxJdwRf3vd1lT2ifL4Wlw/X7y1QxlFbRSu4oLlsdgqTsm4g
ExfRV8y10HFA3FQeUE91GgbS/7mceqTyOi6ZWhCDYj42EDjBs2bmQtRBiY1loiGxlBaRPJTl31FJ
ZpAekpD054JKJuPKLsqr/bzEtdd4SFRrkStBqmv9S30zB2JgqwpwLikyuWHpaDvU4ZpTdmdDbGhX
9nAMI8FYu9VKTMM3MVpv3oHnzvdzEkPAbmm23OOLYIxSpAwvmDQyyUzc7PPwCyGDa0K7nwwiQ6OV
lf+wjasqqf7ocXQIAJeLRI53PaFAshLAXaqWD+6h/zxhqs9CrsoMsqCC109WTRqOoNFgg3p0hTRd
UV7D5DmbceslK9yNZ5hdtIxCYpbHFuVcpXk8+wkGwG6EWVLZvvfwLEbLjNCZKUQQwoyl7GjY4xu3
V9K2SejU1w/9VCUa/RBFvfmb7j5IpzXmdWIXOuxWPVGt8Oi30845ht3y6SXoFf2AmA0A6Fl6KJqc
62v+IpGekXcl2s0qmT4N55+FdugGqt3IzrniAgx/vWRpfQ9Xpo0vfWld0XCP5Qh2z9Lw77pAdmFM
suVxuvTiGmJGUIwirWhtVeqYRmvqYJUDIo/ugSE2uE3F/vUsMZjxPbJiDwfqCFJ9UclHwkul/gg5
HS+vweWh1Mba6bT2EL0wkIC8MTScXto1SYYvnV8aEaazd3F5hfY57+dnwvvVWbQJ6hhiVDgD6Ife
pE7sCuxurIMa7ga3h/4H4gA8mjf9qgIUxs4RWjFPW7IZzVUNhCqarG17/CS/VDZoC85ZSR6vBvQ7
HFfXIqdD8vHwstTegNABzfwJgq1UibaIrVYXAGwNbSN+4hgM3YJ9N+uIb2uj3SKxvPe0JLgkRJXM
MRMaW79dEzdBChJgJOAk8jIGx2jRdOglj+fdAfUDhlGHNyWSv8uQVhJ42PsJjvNAw/HO5FaIkjrO
MyZ2t5EYn1zdKK8EpsEfNHxhZxY6f31lSNS1NT4PW4tfeoMfRc76fOOrNH4y3m250tvC7icr70s5
SF0nC91uT6fYoTxDQGJ0Zv0VTXDnS+XbdQZQZj3zsymrPUIi7W+Uzk9UqiYGfmI3vwY+I4KeT1hv
DfPVsjEvTIBSxOI4+2fFFkvCGDkOmfodb43JmvU/CtEr6mTuWcQtBnmLt47HlK8fX5m5ToO6TUbE
vvBvj0h80xTUdlch6uwMyCPUCU6/W3dhTmZMk819/Rx/s0cfUrWz7PjxBIWiNVcrme0li0oyP9DH
s1Ejop9lDQ0k/8FCOJOtADnNMx7ssN6glSBEGk7vTXfnwyZSFqxoszLK9k3xPkngr3RGerFz9EMS
B1Zyd3GTKagAjAlTf3M/Vw/QzBSjVRI3/1mckDrpNps/ezQhksBfDBcHOI9smR96sjXPnlf2xS1C
yGlYChHEEUyznE8uOIkz4KkpmrsduljHpH6gDz2W3e+7Z+1PBUoqSMV7qZMKCpE9laSJ4GumJ2sn
9/LWmCvMePFZbs8UB/9GOC13musbpXOA5QDqeqVTPj2rLzUqQCfbnOgiD2hKA70I/zvwFZ22hpHY
FRw9FOKgGAKOaGmg2iDZy9O28YGjqbj22R80OTLfUuw2UzmHCuycIawby8Wbk6IH/R0RxxrJ8NyS
KeWOFP3lfuU16e3lnbZSr/zoMKRn1kRVf0Lmr0k4oc6MUmqRe5mCDBsOxFI/btyIDDfhTXP2bMg7
Bs1j3yrXXr0CMtEeoGVqvTfrgj66XgBfA85CEaDhs4FZutP0nTgHvze21d7sr5G9T5qI7sogacDj
au/qgS69SisTETGl0YedkOXx6qCQumrgbKLSYg3SpvdrTTDNT+nik+loP9FHoydU6X0c8IzCCiq8
CEWRtf2oHeCb+FyuRYkFCAEeVkkNVKx2ICSRWWX6BW3AHrCRe4ifC5VPQWrF3g5K4Z7kIUW2QnPU
M623hkHPIrm/D0Gth1U+ZqDWr2qUn0PWahUZuqmyo32VyWcrehc2g3kxLHNnQfWVZl+ZUKKMqQ0D
yq4UBV3MBgCMNv4JsZpnrFpfcYZ0rNdKU3NZnTkg2CdcKI+M42qxCmKaOe27kYebFh5QSD8Zb2S4
MPzfpwXNHjlLFnsH4rb3udlDsreFyMALi9JQ6makh4XIjRpcDrAlE/xcwpTFrgXv3Ipsh7/YFQUg
vkTyRQSsUxXeS2Zeapk5SBDDsMWB5q9pdh+RFaubue7xmO1LEKoeGgBLwc6NWKzo1SoMxdnVtXgA
W3AxNIgpSkDKAmicqhwdxXmmb30BOfQT6NFzfSFXPlBhF6L7QZ1BZlNqnenJtt6yCqoy+5GOrWYT
bg7qzw6FH6bQlkVmLuFM/UUlYTrUT+o0AnsEljxHbj4iQ1kf/Xxd6I+fo8GSaXCAwhaeTZVgaW6U
ZpGQwwDk6jPTAjwRXK71zxYJ5iNPXDAAOZyE8Qy1HoPVfirXMJosvdX1YyjJNcL8QWnyY6CRpfpL
lKns28QX55hL3iaT58nO5XKSKBPU2TxsbY+924aP2gijvH39xE2wjOfFXpJ8W4MeOfI5itOzjibg
6QMYnn7t2oYF8jRxZOQlu2N04rFW/PdvYQluA4Y5SyESQ/FfwL0u1P45qM8NGpHGnjqdFaK/7qEj
H3hVZC8SlL/z5R0NUae2qyCPAPNA4X3yMvC5tFnq9SjCBEXIQ/uzh78LbFkwL53uLHfRCuae9V1d
UaIGNKRjMQ/IXBd/0MyJMt7ReAS5UEa26VmnTdnmlZhLpd86Xk4hojXHGiCcews26FvVD9NTHyZi
wn4hehg+92JCwVvpwagjw662bmJvksR6QI1HZzXCWWWl3NVhCW8MFQBMtHnDIzMc/U7mQk2I8DSI
Y3Hl7GSthh5UXWklt2vf67hD8CwG157BhqsV+YQMLdh3d7vMeXJfQPdsHOVhBTOg1k2cLrWnzTh3
QbXGxO/VfksUBhegDys6mtephOM2V7YLUlxbvgsSRFD3i/noWm4U5lLOudZjBrrLdRt8J/IK0HR2
EWMOmEpwivTnVrOUrnPeLtLNXvwalhgVoNSGCkhJm1cjoc3Ktf+QGVijG25NOtUKxGq5yq/AL6Zj
DxrXtZgNzEtMWVVcWaPFCPbpG4qA9X45YLCmq8NrAYHyeoDWZANX53dHbtcnHvw3Xr3qiNjMWdQZ
o9zZGkten85DGi7K4My8jqTg+kMUsnzVhByIaGxqNjh9Loh0i6zHGBqW99taJK5oStfvf21kEhch
yzizCozLy4QHaorVbq1hf1ZWPQyU+xxzoChzcdNhU2tvNsyPEPbKFwujbGu2YYMC6+GJ2WbOPckZ
m0EBBsip3j9k5cpSxjgc9WRQweY1ojHOa4XwHwdY+ffD+pdfb8QkMigY+LdSdPIRviYSggCJIz+1
Oa7ZKEnI4o/oa5bKCOdolGv9M5pVH59R2WO75AJ7SQ5emrXIk8faFRoG3bIw9vjGzHG+jeQxV4qK
fk6vEjfzg67tVJVhYLyOBBVx9p+kTYyEsA3hx57CQNQCxSZSxSN5esN1L46sxFgtdlQeFhOCyMre
9PTEtJ4tiUpDYysnbTxSEB61AcJCfOWTJACG13eJqJqJQcfYIFFyulSIGsVI8oAI4piyCdA40LlI
jp905ZHKDSA+gZhN3Mbffxolotpn3YYxcfaL7L6FvbvhTtVG8/VzJdZhIeGhCK7B8F3GhOBTohaK
9ugelU8135G7pk7SnF+yZZXd2+AmV6WqrB+yx9mHK4fa6ldj9RYGGhdETdMzaLe2dT0iBPjzf11V
Lxqcx4x2wrgFD6S7VdI5P12tddKu9sSwpGdBWiJ6rrOR4jkaP9YSldOISuPJF0MI9pdTcG9BmSEJ
37FT9NWKsK3jdu/cKm7ssFWCULDVz8XdXOAcqcGkbNlsl/k3UpxyDfQ+Fnjcjhq8Z5c2+WCsLrYq
2zNIBWSEWoQdw0+HbWxBEYJzEIDJzJcX52GdbHbuhIpCyJ8cFU3D77J02b/UUxyd20SNi+F2L/t9
4hmDeE777oSCaDdpuKuKHopKebMkLNKfDP7FQUimqcqgRJ2AuPgZo2EfGrbN7+PoL3+vI10W6Xau
bHt3P9fSeBVqlUOkHoKe0xhtMXwfgkY//QF9vQ7v6EyTs6yKX+b118yD+lmNQuLMHaXfSsx9ACpc
DAgMIY3cMMtB9+2VWyVNGgPjBg3qfSnmwshVwzUtxdIUKzv0ea6OtWgPCQ6d7OyQWc7JHLpbdOz1
suow1SUSxq06S0QiCQoCHWeczG+59ft3T9eVYOYywkN1FbDV1j+yB7JSl50D4foV9SsaZZXznrJd
SbGZ6q7tgeyt3WJNy2IvX18c+XTNZg3h+t0B9iZz5teNVlnTDPt2mGEpRqef9tKeA6pQAT8U8P8/
mPkzd6pbSxLHar8DwK/XWd1GW7QpEvWGxYQrSl0ZgSULfMHvKK2zwgomARULmz1iPAZ5oR+HGWVj
loQ06VhSUj963N1T3NUpArwx3TX8Ke4yhv4x9X702NKjqspdOqJDds2oQ3J18oHS4F7Pn/lWsu3B
D7qd0i/uZHZpBBHrtx76dd8/j7GpxNso82IiDZFU/kYPBVYXkPrbeFtewX22a0Em7rGkhQz4or0A
9uh99Rffxzcm9DbdkZNRmtJZI07kDW5WGJ6aycx5okpM7kWMwcf1asc5KC0UkIJEU1g53J0tsGW9
Cj/wAyW/oxyMbvXlZTXlqf8rVHqv6Z2yTDkD0eh7JhS2CqaKcaaCfkXem5MhOJHWQzsDCQmmJzLr
9ouLGvzK9kxE/EJMmkxhBhR8qgjtKO5rY90DWHPV4Z52iaqaXo1hqg27wjoKk1pHsA7/G+LZ98Hd
4yq7d66j+x/EkRDWUBorJw4LaRCLWtLyAWqqt1ycSNXOsmTL6D9ySl1qP0R5q4gjbA41bi+AMe2k
xhHm9mhI/vbvlszKIMWWml4jBfCzQZvo9hJg8KaGUM2mXYhU3jn6+BWDI8Ts3PGOTJQrdf/EVdqg
+VsoTypESpAD0n0ytMBgZCppr0bMnY8gcwUmPlq0cyhKlzdGZCEx92n0/Q/Tp2WLiKJPQJwdfA0r
zPER0ukIdu/NDPoGvqNCNuP49y8bR8LZmPk1rE7Aesm3OtRKOfB0OuGf2y+r3K5s284s/KRRKYiR
eajoCT9CvXrdOmM45Pd1l5NrM9w1ZAQ5YCd29hKsd8EuYmZtguo+6uYpl59eaWrIygKbD1xN7aBJ
qZstmsSHZ8x7URFLR1fyVVWP7sV/PW5BDWnM5c7B/dln0nRHMFyh607D2lvkj7KcB9wnKmwUJZaA
umZznG7AkA1NcXhQekm/bpae2v/URXpr8/9fJ2HprN7hH+rrz1RUMdTyrl4u0fJyXja78s+Gcixg
BW733aQBPbV/7FOwm3FbNIWmD7dh4B3K/FILqgW+qWsNE4EUBuhSUNzg/CzIut+wrUnu+ziSRjwt
8mgFTOpN6KIXJj7XzQfdGouPYzWF/9S0TZeshFuF7EA5SWcQ1Joy1NTndvl9Zoc4TE7BKcgYGGHX
6VArCHHnWXrY9rEeWAEpJflo0Oy1XcfCRMjpBpfYenoSSRyCBqtKeB3pH8WnIjjrzN/Li4UrAozN
rAXbxZaXSsEyqv5uS1TapCQBCGdpsNhWVwp6i7uXppFEG5jzawRFN0kVJVzO3F1pfW/xEWZMHxgG
6fgewG20RXnf0EpD38mFpgKdZ8mqOTkpnwQ86RylBUWYRR33AoXk4NcqY3fuEN16VdptEp8gEUI5
a/dksTuYF26laVFqxPWl9HLe/5SBCTkzdySQpMxYTT2afIa6bO4ogTx6T0MeFLDIBddoYFpOZflB
DVfOVyR2PfzlhgPvg2nTZRKWPuvn6N8GQumtHxKyzK2vBfUjWyZCS/d+Cmz2AVu4dnTYYhFSVeXo
ZlDY4bQd1FDTQz+2QZD20qhzGoLBn0U0A+RbumVU+FIrQZ0uDmBOupLj1ZwYP3ixUF6+D9JJkqMi
koiBbPV9HOjs7Ldh/h6WO1QRboBCyeeRNKmI2swPohaDg4f1H94zOC+Z2eEASlZQd3/ellbAGCAO
aTBt/E7MbT6BUqS/Cr9+4kGEWktBXk2baUHbM6BwIuksu/Q7pyC5D99mxPI+Y3bYC/WuFpn2siXl
sJT03WWRVD5n7+TEFYJj0JWRuJv4WwHPdj47dSXTkXv9ry0BO2MTsWf0NYj/tx5rmOo0fE5jSPDE
53bQdwK5O0zMivF9utGPohR/+KB9/QoVd4Iw7vK6tzvYYWpU5wgNXOTxStyemuroyVlCYHitT+IO
VGALHgic1K+v0HpXm8H96PRwJUX2vP8WoOEm7ju1TuBA2gpjbg5y0SgGDgZ97CwXf2vOys0axQ5w
5IvgZccH6dRp0xumtnWemK32aDac54UBs2qAXun7j2DXcm/djFyyCpAyWRvsylOSh71E1ySGaf8V
Dwif5kXqFXGIzo0TeVT2dLXS1xbREdPsfnoBxUHOS13Pn4pYH1Hv1yKfQJieGXhEXfO7MyU1AJ2B
keBZvgdWyFITI8GzkrD+8pKSwul7rvbICbOBFJ2/dShWlKE4TxS3+K8HpOA13X9W8+7OK7VyOFhk
zyIsH/8/O0R1Jtf9LL6f369wvIs6O7bw/QOpwIUMsSQoOvqvmDpzDFGIRYZTzEtXemNcOG0C+z7G
Vgv0kdWSfF5iIn7gCpgOC50+n5F55YUOTBZIEZWZA7kx6JLn4XiFw6kfevTgu5VB2EY6+Ub5rgYI
cPQP/IDkmaOcIdXnHu2lF8Zp8QRzcyZ5kRjTCoVzzFRgpExT0zqwuEVUldNe7O+1ZoWaNjCEv5SA
7c0zdL3AXHkdWn3IV/DP3Ml/UUbDt4XI7VWEBVu3xUo2K3NB7TdEKyZoTGRTNk2HU1u2e6sTGOzW
yOb/QUcYJ8mwiyalsgtkgbZa2lqq9IN1T+bGfoTHVQC4aA0JyFfYFx+Boiwm5vVYPuCGtZlX1i5O
meCCPqBEnfE4g50hSZG0k0XT7KgFc8k1tzc9+VuPD29hqW+CtNryn0cnnVuRE0DIHjIzYrjcuOQZ
Y71E85TuoIiknWeTRwnEHkm5F6BvF7yqkYq5rI5d8N8+QtvwJ0ZE35aTw3U5AwEMUKNUGLjhgZsr
Ee/lv+HcqftYAjMikU8D4M2a5Zf9Sue+zlZUXrjC3/6HxNjI3aAVAR/CYwVMihuUO3pkCmtW79m2
nkloBByOkVNbcKIGoihgPEKo6zc8tVP+Do2F7CJ8ZfXJG2qinm5ijrhy0d6Y/Llq9r5QRK4fLTZF
2D2OtzqdocbU1Wo3IpAfnb14OSzFG2BrPPq2aL0fpzyUAcR/Gv2885ukunq5GYLhfirP3wlJ0a9a
ZxuAYP8KFq/Kgf7rw1dwcs9ZcLmXs2i0/xcsJCl3uko8kj6e1mhsC6sM594j03e9CkUySGRaa4lV
+RYXRQacCURF3xWrOComslVK0ekUH3wFoakqWlPt1Dy8UssJ5+O4MlzBM9A5ZbA4Y9N8wPimaH6m
kxrFjMi+8Be0JIjDiM5IKV6oAzFBtLUSTDPsOdjBDppFbcg4Sl7cDX/U2U4e+cNGHSIyxnRvJuQE
mRjaT2+If+n0i5zpRRnk4eweJ3MtK61QIj3xHrmql790FTkvoF0vtcXHKrCeplJRfFAqCPlHB/zp
gm2jbb+uzFkNtHrKhWV0pfixZMyWVYmkK89mbi3iTd19lmmD2UXLeMze+WNwx/GsF9kx9pInF5BV
IL2E+GIEHZ/aGvcoMTIgZdlsnudoNjod2BNhtpyMljGVqj8cx/Iup/cXLRS1p1zzpGNRgdLGp2kb
ZOFdGL+LAjX/3jL7uE9kxynxnAeCxfnLyg9SFR+XvVtsNaulfKwsDMGQdXa86XEGAhpr1yjeM8FB
GyR8IEFLUrW7Z9Gh1wlQTBDjLjvW5e3jEs3+MS1GGYNUHgtbiisPyZDKrNN7ZBo8vQmTtcAhxJek
3Ir3Bdp8uoEm58mEoeFc43BAmhGWj5msYIjCMgbKruvZ2btpf8PQJ6MGcVGGxGD98tvcCAJz+AUa
JstA+rETCrH/GlNB95l9XfyfD9d4kWi8nDzNC0J10fpflWriAHnjYUJ2lhDTiSMQeKCzZKpM3iir
mlxDuLj7g8DoyMCJftssa8yAJHj5Zr+myG4RtCqlVTLMIP7DboHWTNlq0jjfRnPPyfV0RdUPJaCy
AJ2Yn5ECAMPg4bWbl1/GGioJDpktRruxVF8UsGaKIc6EHCM/0e1cqRhWiqmzdd5ewepkvNQ1v4C4
3i99y71/KW8y1rE5DxLEokn1C1WmmUHLk/RSBYUEmt5m3MP5F3PS47wDEZ0+4qHVtoIYYsgIc94M
4csERfzWIsTbkm2XIP7BTOVV63EMLYZd42IonL/230kyqXIPrmcMrHG+DczE6AXZrFb00NjCIYap
752OtUud/XlCnEiRRfFvj+AXtkA6FlCPfNo48Ihm+lhTxdZazY6IDnh2taZMfOdfdQ/J8yBXX4DU
SQqV5W8rTmIlf1JjUyquyrWkza+wu6sTS74Y2I3bS3zjN6YqMvw1y/JF7OLHqwVE28croEAB0FPM
XZvPrLTZWlQkX0BhVnjfpIuNaS9JTbqGa/vfNLqtENn46oiNpiQW5KF9e/1AxW8L9OaN1Wd+g5xU
BHKC/JmBsdccvRDIayYfTQhsV0fmORWQwzWYBfe1r0X2OwPBGnjOOh/S2PWZWXyFO/aCAHq6vk20
gwj0FQYOpkLilYSfibQTuimLdxn3lb5NP7KO68bwa2edKsoyCCNYllzNhsKfVXDBZIol1QnSBjKV
/jYYlgK/QQF6xKFokBXIy3qvhANK0mD7TNjyrdtSvZvVrzjBaQ4jjaVZHbie4fm23cVm4LyCBCoD
eaZvAleJnlvFLIbB8g+blo1zJgwYiKwBaoBS+Ks6m0DGUqNlACRh1z0FqTiFU9BjT9SMtAr66KVd
d7qRNO5GYip2bY9NX7Mvz8pNAQhwuXVlEiTRmgGtPt2+3UA9qf6w7lp5/uMDk4A0dF2Jl9JPIBSq
q2ys/HSRTMJYsNr3aDY/wMQ4ehfRC6KHvnHLYcdIFmj5E3rRIFYEw224dZ5/VfO7GbH8kJDFkubP
E8WIItbEK9Y6LeUPSSJddxGbFdNUVLkQyMqmYizkHTg+tWdT5763EDgwrso+Z6GshQKi4OTySHrH
X5ICIhq7KSUICEjWpbwWaTFRnalEvoL3D0ezgJqXyXPPR8KpxYEM0C5raAE9p6LOvAbiij9WA1jv
NBu8LOiBB296jH9eP+TPwyNq6F5G3oDyUdUq+WxEk+G0hxmQVqmBZhP0LQkrG+v0da2skyrfyP6O
+AmIc71qwTZbr1+dKzTwoaEE6QFNDNgjTNSuR4Bv9qo0/JxdTsuXIzQrSA47B0F4lC7ltFsMRVVx
URBCT2OZmsNmuXVDgialsXIQLm/3eD6M5QzTOZgS2tONXS1HE/9D+bbFkHhZqh30LlXmN1kBlJGY
T5ZA16XthUky4A28MSgbFbUQJguHo8mB16++phUFAl+OnLSt/9eLjFSy7wmPr3L1ZpwBuSJw+BhE
OBrvqd7bTcVZtLtKlAQ+4O19OuIwLMlXlrlSTj+WLQQv1DXIURP9mcgjubRI4ZMaRxJkbIDEpNuP
6keovcAS5z9f3/avCrvGwa5JcUgdpInobSlGIxcG2hV4BAfFAh/4MH60Stec5NUILSUY3pH0DbXg
TPN3RNNC4Pxmbf6d6VVc7MZJU7ozzzDNXSloVUgxSB01SRbZ5YWO8Ti5TeuXjmUor4x98664kiF/
gTUJziAzqDIfN3IyMmTvyYiLThgNmwDrfuaU8pysEyH2CltHJbp83xs1MWPcdJT8damkVqEyRKC1
YH/bN34lRJIB2OxpYjD+a186mFwrt3irLjMKF38z8O3W06pfldja8MmRWXUR6lJF/9+xaGuUqY2P
ZOHIL3RXbA8z2DjwpQeZBdSjS2tQG3/5BpWGv+aebT9yRZJp+duaBC6ncXHrI07+m6wCBVZnzQyZ
jRfVqPQwP+0Tc22qBOTjIx3j0B9EGjEfUwVElc0q1KGr/GbaAzp3X8wbE/f+jLLarqXMgGtT/RuF
Bxby5j+qU2iRIN85X6xRp7Cg0dI2cwM6jmqZF9UmuU5WZIjTbvXsI//3fNMjWk2NPEwt+LYXRiuh
J3ZXrHrnw3XkNxNiT+Cq/vvM8WclGkZtKnqkYocFqe6esCbdg/Wee6SkU9g08K9aKIKGBg1dz361
lJF1USvUYLYHtutb+78/6WidwENQxwIQ2JU8wITXic4lfpDrUSH548qUIdkc+miJcLOlFPD6qnN1
Sj0LIp+Xh+p41pQ9UvDda1NbmrvhEb6o4Av6BrJmrpXh95TLgmNf5LcjBG2NYtIO3mnTVHYdmSpE
8G9mdEHLGeKtwqfCt3WtXT87NGhNKCh6Qg6+oRdGvyFqYQsyXovyKr3gFx5V4z9sjTIV2jHOJILH
qEJcaRIFlytJb5YjJrMI0JyHW3uKBl8dpyudZPjAu+ABu2ZoU0TFA5Az8z3kUUuASYwFrTBufEos
hjQfUqCum0SK+WKjwPM1NpSgzHJEOue6h0SqMF2yHdcFiZZO/+N960LHok5ZnuATlLGOlCEwbts1
c7yLpNUX/n5pkXIZkvf7yC5/7CNOS3kjqrPPBVLPF8VDbdCy+RpPTNUOIUk/5Ayr2Y+7T5ylYXOb
6xSmxnoutlTi/nUlaXFzI46TMd5vNCO/2dPlRqkX6QeOJaTmmKEyWTKrj1rvPdIiXyYM6ztsVMUx
jE/txocponit90YrUl+Z8ymDY0mZs6+iXlzd0sKkwRJmRYWDRNu+it/1zntv4fTnJgfF5lidRCKl
n/LXql227rfEVxUjLATOFfyY24oNUoBk7qKevLR8fvwG1654VjkR/aIXhXtltoNcc+Pu9hMEhdx6
/55WWfIgFVojInat5/ZYscfu1TO4DUAQuLz0ctSyhlUKEDKenFNPGOjjyDoIpnpqFhQcxAckIfCg
jKasyzSHs9ZzfY2SNM1uSGz+khbidx/vymmVlCYbTmoftxhy56zqJ6kDRvlpPL+6CZIITNMVjGAe
GZOlCh26FpBqiRpFT0uuCXhBpBN17sj6ndwERpFfWXxRzq9LnpXcW+gZ7hDwsdJk+CmAKtu5AjPI
QBzbc0bTO7Ce/zLjTQQJXqPwWGh9NNQwcoIGXmX018uRL6KSO/BY7pUNxiwCXi5TkKbS/KeXD9k6
6qkaWjkCgasJZCjt/Ot/Cp7O6VaMn15fiSRDueHOSwTDUGKa3oKfBJo6kyfovZNddvG0pD+ZO6VZ
aC4z9+20OitFI+n9NvIessovJbKdV3FkJ+3THN3jA4/MHmyzZtIsXrnfq7IwrFG/TMXuYqyVB1bu
QTr+s6EpVsd8NioRZxLpsiNptn2wKgHarj5wopzZx03NzB7LpnH6iFoLCaidw99c1Bjw6rt3mFE3
3H6gjZ56EJBiGbYc5Yafp0y+dMO7EPka4SnZIqhqhet/OpesiP31NlK37Xf/66s6ScWc4e5qHHzi
zcy7nFPe7M9jCyGPJHJI6GNLrs+CLD/d8wzoOqtw71FXAFeuvZWJfwT7VZA3WJxWBkNLjdEICZjU
tvdEyWoTPAeprcQZftWOsV0dJmzpikOMmW1hEzQu4Z4Bngb/hHOZRxMEG55MgmW5k/tRp94dr0po
5mBoHpGyWuVw+pNS3Sr0+3cY9E4QxbD0mtFOYThgpd+PAb0HQyslusHd+xrb16+4gnLNp+V0rY35
FTYMrVxaSR0mVZEFlg2yYlDaS+VEpr+omvXku38WIMBKyg4ADDqmqw6SOV1lyuDOVzt/pAYDeNNE
aUpN62HWytXx+Y7YUz6arfEqZjGVIPoXs3CRSfFh+Go8eyZrASX87Y+wAXY9XnZjIgxXrYyghMg6
l5uQ5GEGr0uTNDcHWzzLbbVuxkpK/MSNBkX4caQZVCL0/xE4jEUAmAFpv2XOOg2HdXj/W/rsPA7z
aE/PrOTg/VntYyZvc5j5H0m3iWWyhVQ4LZL9Ozq7imLOcEdnGAIcqK+zP2gcnk7DkQgRJJ92SNDz
cvCsyp2fAtBGnf5D2sB3Vm46zhpgSRsZqJPuXSo38iDiD2932ofJrkn9N5ggJd4aUe/LH7hVX9v1
pwatKiR40g3LhL1AuK3o+u9tBN+fa5mB95JR+as89tA0vud7eKxXXM8M01U9cttS/0/V0f307aXs
7tDGwOpOfjJLSUwgG1fIHJN4Y/E/keGI8ewtv/o0BNQIMxHtVBFFUaDbCqcu293p0ZgTGHxmmAFe
2i6+Cre3mDI2MpBHLwZszUsmsJL8V+AMxKqPq5+AH69BBKvYukm6ojwxDIC0T4S48TjTCBfx6R9O
c8+svdGA8aA0qaYySyq6OQ4EL0QMHvbTbRxArxc7NGogR0eoDAQW8P6Y4SVPpYVOi3YQzsr2WOML
7mR+nkKCd6Cjt/EQICz3kiOrV4w22dkFeuU4fz9UpeqhrVDpMBZs3puWQwWA/zL5+MvjrNcKU8Ee
/J3rHenJvT0Qk8Elcl4MvjirS7piZEJ+49JuOzo34XZQYATT8H3IAAHUVsCRBGUWRTueiQWFBUS/
v7IJxjfy5q+xmOysdKNRmoCTbLvRpxn8/iS/pkI3Ild22gYizcu44ne6pYrlkAOO+DYG4Rs8+WWv
mFrXt2p2ULWvRoFHX0kPJGwof/7tkp/Z6jXgIORQQyrOHIkwHhNiupRA9/g4Jebosg6lWhegj8s+
BdIO39RzjJsd1JHobMUJadZbfuCm7LUWEhSQG8y7b5fQ961vqu8rZ6Yw1gZV6ojD4Ve9+gZCVX2q
rQli7+p14if2BL8OOMew4O8Lw0JcqVqiB5PmX4BdqhCsW5sLYFdqXZMg4u9kvpQuHqRFzhdtyP4A
Bmky4cWsPpKg473yl2mmzAXnNa626/jhwI2YwrkUeZB5Fr7UakgarQBA3HIqHEF28GnoYOEyoPs0
3cGvj/KQKdKHcgHw0sasvVDEsaqXMoQi+c1n4dDskg5GImbmxdH37lcGX/7lvT83NMyyF1bXwY6g
XygWZCl1zsjPV4QvdfPE/8b8d09aWVoalF07zHvs6txj/uZXG7ri9rfAGNJjozYUMh1YhPmANg86
nIJ33s1KZ8SHolC1Gwpqvj2eBSSi02DYQCLUfBACEuAkchZDSqEq9T61TfjD9HBnkHN7A/VKw8KL
ZPNvtcVMCSPulFlCu3Q+5MpusHxBmqGWYY7/7Ef879kOeDscmXdGDA3VgD9SafEMOHpQdQh2L48F
g9PGEvcfBO7g4B09+AyZSgxsHVqzKs9b0eHwYrhWwOSBCNYjQBRBJ+poQUdD0gb4mnB/XfEvWNcH
SZQFSbY3zhvzjnayr1m+DOxbj/HD3Cx//X/Cy2TFDuZP27pFI8pAIYpQWTP7nukbdl2t5tkdZljW
kTaZyWZ+0mZRQhBW09+yje93t7AriMLvZ9EfBfDnZ1+VArDS1sLVJYMvV2c6UZjT88QI/9Uw/pTW
GV0bOz/XzNgeJTnAVWxwjA4bevQNduNhDX26PAqY2fHM3RZKPoRZaBFICXFu0UNlEiolS7t1YV30
d9BQ3+Mz8xkN5/7I4wxwi/1VkM6W3stp6NnNi+67I6ig/7uWY2rCcF01us4XmTeN7j9h4/e2kdib
1Sdl9llu77gGZjWusMwIpR1PPCRWaPvRTcMXIkwbL7ShxntaJmBJhGmPHALgUAui+hLofSrwfWKp
Ks7ur8A6vwrM0C2pwPjPRRFyeOLHme4EhIHFNJDELnZkBH5We4ISWtbWtRcYOrW3oKtjUAEGfkv9
e0R5RMJmXafJ8m0HkBbf7J2sFsx8YOfvrv8WkaOf+bSrRFEv+PswZioNqZhSXdkxFLfWzteW7XmA
iMfwuNAGs427zc75Q2UpLhUSxSO6C/frLRsts2Lt37LCSIZS8RdfuhzwXa91MlNja/xpvN587IyI
bzA+qDINNjZTRtQ7NcTnvAsLt7SHE2IxM/C82fMOCDSHUSSgpfHLOoAZdFrhri1KK5ZBjwOV1cpm
aprD2tTdSJLp8EnbmgJDknDUjC6NuD+0P0je3RFL6XDZ8sYYeWKvNrN+sSZWG8SRS0BHj+v1t2Tw
hQX0qRzpEINgWet68qIEK10gfqN8ZPIc3NyfRvkeeexu7T1qSKCD0ju23VWj8LMBb1iA6nazDhVI
P8af/FUmANlD+MIgLu5QDqH3dqOdyUi+2ylas+1lR/eZjTEVYpji6dij3eOAlGC6DKaJK7sIVV+t
ce6SV1B5AiwqdEixCx4xQ+MAOZn0cEmOIKXKSOqKg/rB+RABN2aAbqA0toNkMqsMO9wammabOIyN
VDU6hnoDJUfqO8H3WA55JsFK3vJfEGHq6IHQBne4TkZDlmz7mxrptqIRDRck2k2fs4Leuq+gpOxJ
ts6vmBA9ez6xvMB9/9wY/zACD3so/d/njo6fp1sv/Tv0IQNphRaQiIeJjeLz4g4hKtdb4BVsDK5v
76FTchUnnMbewJDfMVMWb/hi90ZFKHnOTh/b4Df91t+xOVg5mjZo+UDNsNHGG/3c0baiqre1oXuu
MqIL/R2nq3m62i9WMPpvB70zYibPTKDVtl1qK+6NQjN4HJY7nI5HMarG+OFkABNoez49L5B0qEYj
kvGkUkBYPP5Onax9Jh7i7WqmGedbKqD6TNpO4FOQ9xLGRYM79xIqIoC3DG0XdYw3hMfmj8v05eX8
5ood2+AXXJUqTWnzRhRc48+jMfWTJaDsQFiltBXfaCuHCRPMjinDTDHyzAiNcLg+qF2FZ5Y769RC
5SgKcxri0TMkv0y6gumonQTtPD0KiXrT408/67KG5gpFXhyixHRAGJLaWCAYIBfplV7bBSaiVziy
Y1Q9upQS3AHzoIg+GGnzgborY3pC3piEgPUE7FMhCKzwc6roQDRju+tT0NRVmNtDa80UTJUxSiT3
RztQwOrgvEAbGXp6OXeo32ZDPv4hN6Qs1n7Xl8cEPtBQtQqLzpt/1gjOyPAUUqNue5DUAxukGszR
PkhjhsGBi+ihd2nRyBsLmMtLJZfs+P+dViHdwgESSvON1GujqOxXRQHvDsdUlYfJ/ZMNcYAYuRnH
Fys/+oyxEJFH+W6MngxcfL4ipZwYpfKnYHa4DMK//z6n/H6Zr5KOogwmKZTktdJpl2DKfhMfrI7z
arG+5WRLyzKmM8tx+1arkaorUX/i93psYmB/qGi2dt3aQx9QKvX+KCfhGxzg2WYSOfMi7urTE+FD
OoZhRv2f2nsa/zQvX3IO4dqFsXfpMyk0QQ3xK35rBpmRxWaY1Izi2GYNYGa2LVCzzO+1QSfgsheO
XMkF4njcT4oVfLOmAqeo9M5v0y1Q1D4wYghI76mx3g5RIcbPmSwIl98zTUvJGO+zYtfchMdU0+Hw
s7Z5eNJCbpdx2fxpw6zXOJvG5v3NYo2PZ9Ug5a40Lt37OXZ2pLzeiX+fWzSXfWtiFXfQpsMRqpfh
qfGvim2F7N5NcQq145uNPCGAZwjG3cS2lgxZMo9mppCEWl6q+aOWRGC6y46w5Ttj1IJ16uqQ1tEf
7q/F/tIMGxmkq+91W7MTjBFBUYOxB6nX9f1OzlC5GWH+tfB/pvchBx1CRICA9A5IOz1g11G4Svhy
aHTbB5cyJ+2UxlPzLRTXL/Wb1YB5Wk8P/ORg1s5uG5DMykzpAbu/uTWSjhorKXkYOi6R+kDHrAG/
TAcYjU3UTD3hkpOBrblqMjS29DHuz66wsPp1iYJ4SnEF8a0kCv6477j90oi6Fb/qWe4qVLAqQjK/
1J4Wd1kdaCrAqq1u4NPraVIn417NQ90yxaAPAVj5mL+8ikwYzcmwSFUwwPl3VI5VXCNqd1EXr9IY
Kh3i/8lgE9hDAKy755KyLNZOAEGqasNlPcjm7xFUbeq3PtmqVXB1WABjBwbwsqHuU5Z5UDhN8l9n
9UFKPbDROekG1Kw6ZLDEC6GcuG85nAxEVi9w9sGjoycvI1hBrGC4D9cJcRjpWI1So3w891lAsTi0
PQgzgaWXRqi2Tho5tfnedMluI1UE6yvhzCN3OglOQdqpMV81/bg8QrHA1/2LPxVRXZYypJLBg3pD
meZEVqPtD7BuN0Uu5/vDXdfOy7kQBndnjvQdVCYBaHp0k6OcxqBd0bTgKYWqfhqEtBD/lkkBgp8m
VnghURgSDq5RLdGvyWp/ddTKHmFUrZGqCXyWMBO59fOlIrqepfi3gGkfqeWYc/oNKzhJnHnoz3A1
RTon4azo21ZQBV+yCAFfHGNv3xgBWzvuEmuUDCwz+SZbc0YF5jlmOWz3yEYaR3+HbTqhy1D28DZ5
zEeTdc4ndgtUUyo6U8vE5HsXPMsgTlfWMRsDDYHRjt2f9qPOOaI3qDvWytIY3ms56tgOhRf/euBs
oPoSR7PcquPHJQv0obxiyNq1MSxDSDdblYVEK30B9j4qInReDFFmCr6WiRwVAYdXvVRPLl14+P/v
ZiiPRleeDJvuP7xI8mrXL1qSNIzM7/3IyYGI8XMVG/iWyBUgPF2L4BmW73UeLfxjvtD3cH0a5U3x
2MxpYOdOMUH/ZLNFEtQovn810j5yzNDj7qH7PPYeCTxTyYDej7Oh5ZV3WkZJaez6oGT5Jf0NXwgK
ZFSMTFhiAaT3UIJp/+H8IK0rWBuFEbAAyPJTZ11I2tP3EqF6PT4fubgSQpOK/6x25GS871D2Ua9I
wlVFP1pojMPsu+BdPVeymSvn5uR3gBxTgecC33up0ItNihqqY5GMkKfWLUrr0XyGtTZttyT4CwSF
oJa11oQ59SFzEE0IUMCRl0PJgqMEduiBPD6bSMBQLUA3z0MUrjm6hkk5JOlh/D69DRznI1C1tiWF
QrYhi0szYyV9DIHbpMmwoYi21Tkj/m66k6tsSw8nAFY+mXervFej6eo+UD3HHv78DZXS4h08Xegk
N72yrTRepkljq1D70m4Qgrx+YtPi1/aYUbdv9XBpRQ3Lan1KB/IWvTUYeixJ8XO3m/uzcfva+g8C
DTwY9SlbXVaf9zYKeDHbGBb+xMUHsohe6pgf1mG3JHnGLLOp1MH8rUfH0Gc1GrnbczV8H5yhL7xm
NVsqAeOmiEFJkvDq2caV2b2xjT6EhRzxPC5rVvOT3QYSzNoOJvv5I3eiIbKceND2HUvbefMzdiX9
o4bwPkA5J/wuwVoz7g+qfMJ0K4s/v3hRWvHDTAAjAgpwc91+wlGY870a/w65j0RKxgNURcr+TqnN
YKgiY/uldwD/WVENXXv1NTAS+mrcQHQM5sAIZs0W8JfnVR2rX2xVnJe5bdXLRRpcbQ8JoxdYcAtX
6xItSW+gn7l9YlWtn8zh1XiFaaKsE+0DLOQX/EkoA8cxpRC9fcfnRIt5s2qOJV67KJY4G/e5YR+e
JGaGZiH+Y3JNbkLwbahtQ6QlI3xnSGwMaVnUUQeJTOnsCqaaW4TY95+adqgB+1z4xHKwU1NpfDU8
aTZC9ry4V3aOYTsuPaIgHiRSoGLWo9Yd2jJqHu5yTyfkMP/IEt9MIMxPuu1EFHijidqlbiIRa91p
ODrMYdq18rlGwQKsUQquOcb07IiBFPOGEpHAerjqLklmsqtAsIeS6tgARN5Czy36xiP0BXs9W6e+
VACJTN+pqtySMVG9ZosMmkJi4KEbexsxJan55dOSg+a+CpwM4pV3Yw6ARPmZiFPMu326P+1mfZ9k
YzqPSteYnllhmFLOLGeXN4jf70QguCLQknJQNFR/720pE59PP9+iqNZjULutW8NXT2tiDNnC+9+Y
CWXIv1tv47sSvic7M2wf3y6OGTeEOTJZB/iwKyyOFFnjVMKS+9nVmDIJhvAETFRB/dwd8h9tQSCA
NNLYSCE/ALOflIu9PV2ZLxU3uupNyrMienI8ZW3wt61ezqGGO7uS/hIBkiQ0wJzcu9qPhKq0ogoh
tV25DK5uDUi4+lB2sfMLDyMHOoNrVcEoeIQ7EiLHFLpmOsV4yrq/3N9r+q+HLvKsySCiM4Qk3RYK
fSqT9ZOGqI9NOJh1wFsYlHmPy8Gz8+0tMrL4g26bC1PS5s7jWesp0mMSgYxi9EP2ha891MTMfojf
zTkUH5595uddCy//JxEaj61W/HQMM/J8jYl9OdZQdORDAVnrSNWZIXzqnYGvd91mB1eAsDMsFRFr
HnZSTrNvJShByKYWklnz+B+mnjl5J5aDhwK9xm5udncQ73lJNwO9Iqu7K/8MCLC6Cd8uhuZSToRW
GdlsaafvS/dJOG7g1v0hhcCSA+v3Wqd9OIlUuxGskztpdlq4uSPKu7/5boA2ZT+sdY78+fSj/77v
QGm5yUgVxun/Lx6dCJvWtEzt0uAol2vRbh4p5QLdYncaazZ8024jINvYubH15ePNVISrMd44Gsyx
OFnb95jKC1dK/dvxbFmvZPxhevxV8YqE3qXadRg7QLTDk29/valzo/HPTC5Dqndagrsy1ye8lDOq
oQDc84gOiMvjykPAaOL8fbwhhKgsQKreO3lox2BZujFILkUoxMgH1yklBUda18c9nzmye3tPVksh
U0M5bZr40C8jwMohvC7PD37ZKRMOM4dm+lAFiTXWYTWoo7ZRM/5Oxa2+rRID6kRXnkFao9O2U/l7
tJwvp2JdH/yWfVhL6DaoAiTVoDF04u9CLWM0pw3Sl7LVBiMCvwVK8z2fHM+nN+VpLHonbqVeYcds
G/dBv8ePodcukh8rNYRUy2PRvEdL4t9dVwt7S0PU4ahtWDbbYGw0rr8zPNNRjwF/b4IcfhisGbyq
8uiuV4oCHOwNBErWTkbV4W5BCfNWEuZDFAsnoaYAdvHEU9Ghc/Uom4GHBRhO7qpfCMsggSdqhCSS
XPe9P19ybDzZtMll9pSWe1a8PyPIsm4PxomUchNRA+bp8x+8KfcQdyW/CUN8uHpl1a3mwPMdXq3S
HcHRf8OvLLmrP11sn4uXrFsr8GICLkaQYJX48ZD+eK3zUtUiv5rnZY7J6Ua0KnlwZa23wLaxyeLH
xcPU4vnfYMpZVaiqqsYRTRww+FQFLofri2RRIqZlr3EBLxYzJOJdS3WlrlSHyk8Swfg0KsqTDcHl
qcFX1uKH0R6JuQAQDyH11/mF8cLeXZibZhxqErvf6s9MyS9egvr+cky1r2O78fJ23BDh3hLWP3Tw
/h5v2ne6rsL/ybAnDaVuV2PDCmC8B30gSIRlPzk7mvTgrUPUbMEHiJW2lFRNQDkVsO6UEjV9xkSK
q7nwMjZPiBPQ388pBUJcRWWYYuExZ1OaFpyNdpZ4I/2jUyHyKRVGrwJTDNaIr8kuKrDStSMjC/yR
6GZAoAtd95ev8NnC+XqYsfk255wi4bJdhKCDPuusDjJlbntajlVGUaR+9Av+Ofs6tnBMl7NC9AvZ
oN/56aXu9t+r/KyCLFI6f0WYph8G4UoQh/2cyBlSKlDYfLRST+0EhM/HteFAhB1oz8HtU5KTUFkU
7qRfRandD2gmvknh3e8Lu5gReg0yFqB8SdwpTS4z9Uh2XdVwWKce4YLoynT5lYrOCR1P7QzKQ0Yg
xu9H4U5z/DzmnBJ7XaSwbANbiE/ghuPrhr1IYBmr8Lp5BvtrWpXDzNNjhBQ9qEs1xE8Heh4tSIKE
FWXUHjDayyoVHTzi7l8rYA/vrAS+ijHOluSiIeXtc/3ocksZ6wBh/bUsG3gx79XkrYwAlPFsEA6P
4+DX4h6fU3uxWyPAuf1JBDNPaRDl5uUYehFv2iASII+5nBSPg5/t/ofKDiIcEwzVapInCMA4dKEF
Pn3kEGJzWlcpY559z2gAXUp1xr8JUlqf40yY09w6UBfWg8m/HCefAHghWTe1FduBa3MdqUk+/gzg
2EHsFRQYnhF02Mx2eyVhIxPZqSQCDOTz13R6kN9NaoyWqPTrk0GU786SqglqGBDM/YyDBfu9sY00
ztw5wrZcRXXBExgDHJf6O6fLiWWGPcmZDDMq3kkvrOrAR4UfwsFHOiqkhTkVNntWCMc/GnhTuZqX
HQ7TYbJ4rhZqgAF0/2OmLYpzVkfpFSe7KdmJ6H+1Fafx6BzBcEV+9EjsVoZ29Ju3C1L/weGVdpQq
PNalV2sThcKFj4F4vsWXWSEi8XgvTII7aDpEdpVD1cWGwlVO7Jm4H7Ab81XPF++qzuifmjsnlOy3
Pbn3PVUKe5+9GJ3ZUHvDayrGjFsRPBEkgqEIO9Bdp2zvHC4qXsBlc7lbZDstJP3D8DN8hO9BTEP0
s2HMCjWZdM1U9mWTT04QHQ6wgPNlciP+r9NFIz3lhoOxPuyGWdykh9f9vZAkQwIOEycBsFpsyG7G
sBv21eBmbPGe/Q12NDlZHCbyO9d16OFy6w2ude+Z28QZmaVdTjyiIUMcBiKeSxYx4MypXW1J2430
Ss0Bm678QxV5cZXl2IEZwyjK9KUPeGKYLgkUEHjQhuOQg0qG/yeRdExbSrT3QXpysfPiBPVnW490
ShjLEsE7F5dfNX43AplxCz3zw8sSk/6CX83MMd6OI4R3vwRv0ID9ebvcHZrcg9gT+gDLAXDnQcsa
f4bTaMoFa5tO9xOgQVSi3BBlNNbXJcwVwdQgzk3vQaxicanmRoR2tKt8Hy4ZRHG6+nbDNla6WmnU
Pnn40ApZ71yKtWDiO6C3SQ7TvAxSvH38an2hDOAoGPVw0UQDR5VxJlU/ehFyiH83i/sOLXVtZlGx
xqHiy6Wrt9shztq+pyZ5CtBUzk0HP0LcpMv0p+TwDMaA0yRYWceLWgBIU/QcfnXdsHqx4voFf9tI
SwjtP8mthNCddJWmtrh7Q0VJkxtJVG+PELWaqEGy1AXNv667H1eO1mLcl30VaTt64Pn39KaSKtqn
zosG6vCSal2jEzX+m72eEjC5AwsH7NxcUffdDU+H/gBfDm+5UEzknMy0cJKBmH6ASmOcd0XU9y/D
ZIo7cbh0RTVo6/6edjpA02s2nP4PsL5vE+3AWZV8GBjUl5YxR6+tpBbQZ0QZtpFIHpGCc95tH15s
ghiE3MYqtaRQVfsSHBhjxsdW/nOP8KFslsholVnBc1TsoIDzEvs3RZDPL7PU8VUhb0gCb2m5oHs4
hDqyOyfDUemb97REz75m8XMHtRmurZGoex+NtJEaVL1Gfdye5Dz7IX8YkC8BSS+SNW/scDzJNH/+
b5w2WpwRsOkmbZyrzqkBOjOWiRW87s0ALZKJpOR05xQ+lUCqA9PuFBpYzOBw78OI+gpcdxi9g9OT
IJAg1i1CjRJV7oY4YS0OnQogomsqN0VFwx17rWnI2Xn+ncRAu0hheOQQt9TGKXWMX4ZJF0GCukkg
pOpHxRjY9j44dftGVf4OTSVaxd3AmOmcQQQ+Uh2dyDXSsJZQU2234iD5ZMxkIzpgrE257FCsiNTT
OEcvo2CLTjRf8lyZhzPuu/nJZWDwhn65vqMzFFM03tEb19PcA+MvdjnxJJN/gt5O5ii7EoFZB0EG
KcZnqADm8IpuXWrIIlRoagu/OsYMfC6ABkPruhDJnbA/lnwZ1U7Tl3Rs8EF9MHZ/rQdwDednmCWF
/cUduHUqcJ3JRA1vOS9Gdg8OCKpSMJ+j8B1V3hfUx1mvKDs6H53giJXOG9hz3tVCgm7WCI/Mh3Bf
DdnbHSglAfOa+A8b15lPcBkSHDsa1QrHJhEyqlVG3NP45oP8FrISCH3FUpoY9vDFdIcu9XtsqPpD
FlY9eE53rXn5JWmHqWnWJA67cEJFVEnWjrY/73LsSQB0EMNP4yl+4pzz295Qqbr5ghAv/uTyxZ8n
WIzE+SDSirNfdRZDqEzXw/7txsqI46uHXlTagyk8S/O/qgAA71a4kryZS/X+OKZLERMM4uUc84//
HOvZuxrGhqwe73dXoJEOKBL+TKnv3CxpSGl5HAGcSle2xtjzdgw3zAVXG6pgZ41g87FhwpRnHyNJ
mn5th/4RJ9JFb6ByihjkWFaxPb/rpju84VC6Inm1Edsc3dXr5xuHMgm2gVEqHhz6R9K3To+6pbG2
6sqYgC7MBX7EPFgSRadCtYbLeQM1KDKwlFV95rY0uYOiMyxuzTGtFMqT9f/ZmN+G6xbGuJSUUdAt
HcJxS/wTt0oGKfxfUclqEnKrMakhZT68nuItMZ08bgwtuuI9+rgbJ4ZBDOqx1NHRrLx1ynjweRIH
lvGYxqR9pYsAI6Kk51wAJrm3EtBZulhK2TiVGkMBpKT3pjnLGRTh3Rtg0z8AMa9zLdlq/sktI5gW
TPAI6A7NPX/bVjfvwqWyD2woI2qer4i1sf3EHPH7WcRnwcEeA8Um7w6KJ2aGrFEDSzkQ45hX9jkU
0+p5J5uRneoOM5f5Go7nRoQ+tDB0U8xJ9j7VQwCDE/OfLvmxVExoBR/d63FS2VqrAmBekkW56wBC
m9JaqQCWUbtmAPWppzJcw+pwrd84F6PSRt8s/W0nWAP/lQm4HCv8FqB6+DzAm2HHwhEr2OejHuB5
yPKOXJdm4yMIqOsK3kFxidXd+InTD3jPUUJh1+3HmbRa2OVdz3+jxArjLpCbduczni0H8dwm26/1
f4nm/n6xQ5qKZxSdWbL+7FgHXw/h4DO46BfGqk+jJzVPhCnzlC/qMqkIi4QIkEXChCDUho05/dNl
Lvm/TGvdYVeNVchtrTKpVmgqVNlN0oqAm1x+kPzfKWjyHdofx0TnZLTE6R0SRCmcAs5q8qsmNLOq
a4d2A59pMK4mphWSAYqiUE7zFAAkRozyIzSDoCBOxHCoCZY4of6EWCYlyUIlKPDjKJQJGFV6+zmW
o4seLbi2UO5VgObVnpphtZyGWj+LvGAAz/m1hzOv0tgSZCISYSo+utjccZLOpdSoqJVE5xW2rE3H
J7nvX18njk33Hp0hmIswFqS5muFjl6VYuzmQs5dp2mdle7YVHYPkLj/kbGJBr3y0TNLkpXisEXf7
6LmLusTV75nURtwJO3Sq2PLt0LKEQJ5t2mKtDMWd2eaqfAFRUax9Hmomj9Bl3JN+QkVbEB1x0n3c
reJiqD/XrtIG4JE53UhbkLNzBTXE5/xjiQF5rnUC3vemUL3ehpXUEsMjNXGTGwzbN9o6YfrHZ3JA
ihdFtSJP9IxItJyOjlFpBtSS4/GSv3O2DR5O/BMQGkRJVwjgvb2EymmDfAaFXcc/VmbXsZg3QaYC
XaKfPUQeXcxCqxRTvLZR7aAgGU5snoGzsm8Mg4skgEzJMW9vQt3Aj6toVR7jXq5/gjUbwZFNsha7
O4aTVE+/VhZmCxjFwQOPut6WIijNjDJtuDM3VG9pCpGECGhR3Yp7ER+q3HbNQ7VIndQicWfKCAV6
VEEyVeXRdxbhRyvf9K0AKr7ZBwhcPaiWKELEhw0/Zom4ek4dBgl0hAP7iMG8BlTuYLyeXxFA+YNe
N/zCwzKGpUkG4AlmtS2BvSTKEjD0UPoQUT3lXoOdgWCajNFi54rAj4GDogWg73kvNpfK7/ryeqyA
DMbZPZAPlmxIHtTQ4bP7LxUTwfl6jY6PktnNIeQDGa1cJjjrWZABDryAVNaUPRsenArejF15ubeo
kfGcKIoIYcV4Aa1qNJoL0iLW1BbyHoo7AiG5V2uGdAll00r6pspDfqCNNdq7hlRgIhmuEbMJGyPn
qRydKScGvfg71ginbn8KgGc72sdY1AN+A7CRs1mnuUsQUzaJSp0UVfKAL8VAnykLVOOHk0M68SbW
yygB3DxHWLX2P2eH10EBSItMHqagYwRB7hy17IwFcLEJlfmGklzmNupEhGdz1Y2WyFBLdfjVqq8D
ChZpIaVvHVyxVH02GaQJx231xyTHFYH+IqctkSWlpwJwAjqAaCf5F5hV2wVAKZklMdTVMpDZA3F/
8tk2ED96zUefyePNqUYiXlCMdgDfYncSeZJi0N0WecmGSuk5Hms7OnWwO/24gaNqLh9OfI6IgIom
Fywufegdi6PRHEXKcyVMreHwdEeT6eKSJeqoIQ/G9pK26EjLR5Bt6Lt7sPirWLutfNrImQTIkG+e
NBJke1FbQsJTE8uIF4Gcl5Eeq4a5kyuhs0+gSg1fMqDwyKOcrOGf23WwrEtR52z7/U01td1tfIdr
BZqREOxFYsQl/Rr5TDjW5zpIYtNvRpFkQUqyvpVwR6x1GVLhoAy0nGGlvBTked3eqIxw4vhD4T2D
QV4r5yaj2sypB26Pc/TcLVrcf766IiEqPBEToz63K+NGPNIBe2mjMgZms0tJDlpuR7/rbKrFLtE4
5qqYpYaS3K4Quy6pRY23cs/nXSHII0hZdfVEvQ0QLWy3s24U+fF5htShqLyA3pVeVPwmG6XbfqJx
r/YqdURtmz5+Rv7YUIkRFW3vaXkANPRmpZgpa23MOoeNCKKm1s067YTS3TyUtmx+nFl0Oz8GmU/9
hM6C+b6KQrqCLgGXc5NZ8DpVeSIbZ5gp0SM9Raf5MY84C0nXo0mTC+BpB68Gz4KTPheXFzqNY8vs
20h5ux07nbU/Ib44Tphs0rYaRwprn0Rouyo7jp2ACyoJRzI+jJAfsYXhNN18QGR2MraJVElCrr4M
lc82O45MXV4iUyTrMw4ccNEJxnxncaG86S/o1huVZV+u34yHtIrImU2pTriyKnPwNynaD+VprEez
Vatvja++TElDQEiHt4Zpi/19x8F209XZ9l/xVSnnaxT7vM4eATh9rnl08RABv/1c9hWKJTIXuz6S
7FozDKnDZMIOrCudK8yheL4M4YNXicODdJ/skpx6dglGylzhao+DosOfEY+J+nczkxYnNyFDrYoN
IR2F3qwtkKIz+4OYN1FHtJySd/V3N1hKwO8zHCAK+UnTRdC4QqQxclMPEc6lSsF2Kyi1NWYinHKb
MafV3mxqHTYhDEqEIoYF1vacsjaDviXEzM5nMWNXVH/sIYgJnUsmS6vyjHlYEngaBIjSyQ/UekmG
DyF6jsYuk04RpsA1WhIFBXUN3AbXWE9S4kogfNAqLBocc9XAnS0H88z7A+fYXYROX8AAR7BPWfP3
dY7zwjJi7JUqHFE7ZP1Ll5U9UrlKxiuLEs4ogAXDEKPZ89SD6BlguPLG6hRKRkyF1i7ZaxIwr/jh
6eM9vMD6ZmZqvGujNSorI10MYE5W1gI9WuY9ztZL9Tu+Ir/0f5VrEAXccpv/nQTT43r6fXXL/CUh
HECNFC0yi8Outiic2KOobJ0BBvI6zw2lBEHOPKJKk0dudSWXN+wcyaLnoOcXsr32vmlwM2CHR9LY
5rlXcWdAhnJGKUuezFyIm509GvJQUZrrGLqpu3Wsowt//vsPy8+7OtAQKfPi9Ou7y23stz43RDcE
ajRsHoGJa9mA80ClYnJs9WyjUY/KiyVnGzJq8ydeVQGZZmrAws1Z7puVibV4muciTViGg3oPfuLH
uB4McSYNZbEczdsAQsOi9CouXc4/IwfNihfdoHybXUc1al7o9NAM6/c9yEolCb3YR+6EFZl2wVX4
76Z/IBXwgwzeF7eZQJGOWDrM6yOViyqAwt+VxThDoAGmd1XpstTOY7OlhRKFIEQUzh1EBPgAT89I
Z7UZnS5kHLsQ2PoOFZpssuOgTeitWjDfhQoJExa0EAKs3aZhrGwa1H9CdeiPIoN1lzy70+W/1jVO
3K2H64WL6f1vKl8nw9YBWb3QhNOHr9HuL+3FxTvMw35t0861/pfKysDSCVU46wKkiyjXuyo1FKUb
ZjvImm2TFmEeFNm8V57uu3po74R8RU+aQuv/VCJ7LA0OzF3EYENbvdJ705gBqnSDTeb8UQVLpW4E
BRCQbAsIFvF8s+dKuX5HZZknL/deY7rt0FZimNzTrolIDHa24emtna7AHVR23DI/gnEQEL9h3rlH
LaNWxaJhnFqaDvgPfmATsmyAn8QebUmTIOwZs3SPEY8J4MqVXu8UwTl6RVk8qjswphKAMNGRS7O2
lDTzDqx9bazFsrr3CI2qtRnYhh9yVHEFBepkcJjx7U4vKAXSqDYRBlLNXj7D26WDrc6oG97hG/jo
zWeye96/I4H8tQnhTwHUNAE3wQLxROMS0Df+NjYd9Aj2tTWLi2gEpO8xNw6YV16tsREZXO3asP3K
z1z1qCDrLp67YeMUoR2V7efxTFJYz1qDVo7xkRWkA18SYyi9KoDIkq35K800OXPHCQv90hhsopp7
hkZiFAUJ6/7ODIJX1JsjtoSdvfDP6s/EkHvCHLBjOvclcNBMg4/Ed4w58asvb5wrWrstJXGxXate
XJIfl5Qlke/mq3xQxC1+RtyNxO8M4S2m7XB6KlQpN/NbBp4x7x3YAZSS3S6o1GEF+Qi2zfZ5iGuB
pjuB8MLjaGuK7kGldI50rwnYWIijHDYjoRABF958spSG9RVt+/OAJ4t6R1O5uv+Jyi2zZ+qGEIy5
44OUuOIveUpa56xAzYlGKeyJFLa4ow9b1wK4drbjJz3B4DsE9Azn78cZdr/huvwIKYIOs71RFlqu
cMm4ywiNjFWofC+ECrwKlxbFl8h2qjUTf30CElbqdW2g1oFuhZfNX8Ao7RZ0chdZpgbD0FuBgJoI
pVHgR5o6v02ujN9dLD8groYPU6/vX8mrY23fX74rvJGlQBdVWUKO2r9yxLG1ZifWTnoaGh04CM6y
j9sN2JxL/32c6NCXIRtyQ2F2aTaSCSK+dqLKycq0xK/IQ8/Co+TvrBXOOoRRxtlsSXYiH5Fwd3ho
W7eKPEJZW7x9SyESBJ4P4hGJUZheNbUyeRKe0hP+lhqEyxPhevczBlRp0QS/5KLW4GtCrzBzfCG0
5Xxay/gREwjFq09884DizS73ga4ZQwR0Evwg+krI+wVKZLgqSOAyqzZB7jeJGTktPoXVlyCYafci
r3VpGMq0ZT0n2UCdwkeiyP8cAtLILQH2hKD3QmIETXM9XRdCNIr5KoD+9QE8Gk9R21RLiXhJzuMQ
v7Cu7l3Vq3spdNvxhE2OwVgT6fo0We+AEiiuQ8Nrbwm6mtvwoELXB1AQEBZpgyoJtBC+hN/NPKf9
wP7TsftXPvKOxMBxv7RU3qs8y5FF8kEoZth0rt0QaJgb2bse48+eWdQ0ODyLsEwboL7KUIzjknks
HFageZI9apVyX+TcR6B+/LUhsKgiituGmTR7GUC0yLqvKHBBKhpQrvd3HL/pg+aGrkO+J8LP4/xr
J/ew9cs3Xn1uLwBS4M3soRk52C3Xt5EmWhnRM+K1LCcAFQJ7xOBAu4V3Q+TQzagA9i8iFvGKGDg7
BIebVmBV6YZI9p7xZXE5bTvV/xQRYXX+3b+33m8BQGX354HuXlyYoikl/8qvrp3INTErUwoKSG9w
a6w3/YIULLney/vYSybdrwqbySqJea2oLqNR78w1hi4B8KRzKY/OSa5Y2TzaFDIHdH56mAUcFV5i
JYn8R6Lot6UyDHlZarujpj4NKfuj3RTJLM6TXHAsVuYSUlDCkI9ZbdoGzBwwsp4JrA979D7N9YSi
ov/nGF0fUveTfOvSmVq52X2vXvtWoNIRzm9mYPI8BxcYuv2TAfg/bzh8B1Crzt9FZTjLcSSX+0Ny
caVTepULy5S9ViF2cpkAaoTod4X7hgoTQN/moh21yzb4belDLOX2K36ntgUCibsWDY3HDFnunSDS
DSmo8HEh5KcZBBClQGTOwIFVcajT/rkXqmk9Usfk6Nbk4qw4mMJO1AOq3Pv4bRypOU/9j6QKDp/V
/YgL17rvQc5bco4n582AqjOJ95jqRdW61CnkdPsoKXhlMT2nCgbh4DX2Icc0A3xBBmQpYUuJLRMD
h9B2XYFc0nRbVGxogG9aeLEzLcoqLne+Dz+6UKVDUmdV5TgEk9ekj/SKb5I1vAjHGU7OL8q0z0VP
uB0ztUYWXKLxPZf3ix5M09xBVyiAeQ7pHZn5zYeC/xh1mHIeryYreT7cHwjND6ladT7A/+QcrNQ2
kOqkHtuQHu7GicxYsZJ9/CQNAhVyLsw5YpW82Ai2tJGn52/sc7VFg1WStRiXjP2vNLVCk3DtlrZU
l5mFQezvS+SellfvEHkUkGowGUjImLimvAUm9p1FoAUJfZ9sDvK48TRQ67MkBNek31jgXdwoKl3x
efD8fAXErz1AxBea+9oTFefyl/DKqTCavE5GcTQSI43YPxyKG3975UqJ3IHXfec/CyBorV5+eED7
Y8fnr+5wJEjy+N2rzIeVhAXXuNg0cRM9adD5+nJg2iCy0gUD0Uxac5KFTOd7E8F/qAuVNA7EZKvN
U9VVDKmlvHl3zaiPk+fHQ0jFcd1Hda1bEfr2hHm+NnfuyctIR/k0Alf2TXnM89znVfvU1Yx5cRim
8fsJLJFk51dEZWa9lB58dgrEL4ih7MuAzOGJVJyN4I4gCW1gT7aJwrOH2s7DcoTuEXz757BbxOrp
McBlIUfy3eYLXZjs702/XNJ3+d1Q/RjJBSs3wGykOgy4FuQttHgTKntSO1wyfh/y4hOLINLHbjLU
DDVSDU1UPcvgnfLYfnnszdzCybsakgjpeL8mEUX1/ne+vuAgjZTyHNP2QM+4arYaUD4sHs1XKi9Y
qj2GYGH7kPM6y0dpFHPLwtz4Bcf0VQKiF2dvjkMPEGDriDSkSICgBI/eNazAmYtS8zchdmnhjz5v
y+3e61i/O/9+wr7tfZRKWAMxaIJc4gbIDTyh4HIQXp/l3wLKhJw43f6ekx6Y8wxUroHeFSkh3grp
UvMDlDQcz9/Bi+CV6RrphRByFm3JJOEewgFRHEVJARLtXk89iZKuTMAwyKolhby4BdInzy23hUyX
2VXTyli11xbw3dQ3aJGo7QHuUXBzsZVUAxk8oSQsPO79+8DfI/mTsL+nNnm7hB8VMF9O9QtdiQ1p
+ubrjTtAV81QPSrsY5Sy+Gp0PRMA5mwYqvkKwAjEQVrXbSPc+TtjeJOLrZwpWmsJOf0zib3VrPQJ
L28UPMtlQ2iujExVkcnFvodJjVjxViOv2GXYi9ZnZzoZe295+npnR31KV2EtDzCxSqmBPLdheNPt
AQAPae/ditGgF0nn2IhT+dU0nrbtnHM6uiZc+eUwb8kZ8v4QehkWPQMfioavR2M7wqLWYIwGQCQZ
EyxksBrG3f88NwZCs5HFEqYGK0n6qF9dw9aZy98BBgh1FlIa//zzFUrjEczqlM27kOvqwpWLu/P0
EFNJ+QMth6nW2/dAKWreUfw3ZQON9QRT+FQXX6UwIUnfRei2lLteobzRqysg0GtGdo36jVJMYhr5
i5r3FfBEz/J8HPl4VHqmyZ+j49kgWe+Id57FB/BjwY58tvSNA6M/rKVB1MOCt2bmOrbIIUdiHz/e
7m5s61um2KMf/kq8RrCvNIDYm4Fvqgg19+RkQd5DrAUKDf/p2eMoRgWs7fOydXY/WuFXm8/bQ3Og
2WDH4DfO+3Ta4K3JY1UfH7ZU1cVrhU9czeOFoUhzcHZax48yi0NhsXbFMZUO7F90crhYikpiKd0+
D5/+QWYi0zNEqUmiKSKh2KBplOl1ZtuVlbZIhFBLKD6xgSMxoqZ3fdy9bMa99JpDoBqxaMMXkhCT
qoUNrjHkDc9H8hSE52RzaQhGqkSHCnR+xGtIC0Gf6ACdOzFmiz7u0Eaw9YfKBDyf2Ms7xK7d3OPA
V9yUZlEn9Rwbol8Ol6PfDWSDcTJDTesII4blrzC4JbUFDSHsRe9Ic+9SDAsOmLUSH1brvvKBkVkZ
bAL3xhvEtDf/OsBdY1wExCMJGUqUJIQO0wruvokFTfvLCK43jpSDIA7+2hnYH0/N1JRVxYIMjFAn
1yKA3HOoI/CKyNdAr1pzGrcncbyISQApiEiW52abyGk1cdcqM9AjHAEStMzV6+IcEeBenwOjQLZp
3RYSd2kkrtuwTOToq7BpB+58r7RPl8ZkBrY1YdTVFdj1RJOkcSrC3lVPx7Z8hUVGyW0Rvgd7Jpa8
ZLg4Lrk5aOtoatiWqnykNrRQmY0hszbIv3xbwz+Zvn9s2y6lBLCbLUpzwyygQo6me3vH7OJVUpBk
ysHU1L607fZIsvwx7rty53ivwrpZ3gnQKfUrZtuG3yIJFjC18yXOw0/BI0b2R/b6ioiF3bRQfJw1
CGwTVRr4jUuXcCTUIzi4Cxg8vhQDIkOxjQ5cwM4NKep81D93/wru7ZqQVxJzyvEb6oZzm/CSA1y8
mbBud9xnb5RPDCD+wKPki+EDVcD2rcBkuZ879Fvd4cBRDXszigfNbRJjN6QrNHg6Xx0/AGgnIGHZ
rIDt81yTb0p9BkmUhHWCQ9s5r84T2HjxCoDTqsOpahXXNcu5Xb/8sDEc7d32i/CsxQWBd5FcAAbc
bp4fQ+0LZ/NocdpSempQN7AtHEr125s09i/QD+ppFMpjSuntfXKKVhj8CMYuw0UHBpBimnPUCdvI
UnVlNISgeNfQwyX2PUPmpeSjSOpIX7Q7sUVqK7U1y4NKuNDDgB0djE/M5Mhizm6JTnqU01eqIilS
n91NqU3har4ssyO0BCyPSmyNGYOm5q9Lkbv3qeVvGK4T6qGGrlJ0XgjXY4/KbPRV8/6WcbV35xZ2
fLrYafmsJ7oqKysMyIVh2PLXHEI8kR+mM3npdxO+Ypu3bQhDnAr8lKkuSBX9WeD2CVXtNDz7Axri
fjzlGDMfo+Ul/FcT38afh4LDCa7Vp+l3tHNWd2cTg8hJ3zBcM52dz2M6fNl9UotTKIA+Y3bz0CpB
A5Q0QHs9bWNc96RfWGK2SNwCnzdZ+YGrIsDTJNSg/MT3hiSF5Q6S7QUEPrs09nLKyKya2pcE6HTM
5MqDNnxS1DaFw6ilBcW4vGiuzd4vJ5iSj0tL/Tszsebx1yFY04I5DpAJJ5DxCSE72qAGTesE4KJe
WXf+eLit3oaeLn+K1LedPLXzPLUxJNft0zzvT/rwzxWQB55eEyG/REYvsZTD/skRwXUL4vVP8Jfj
LqWNaLIZVGvL6xzRAvMAQu17KXiU+FgED4mZf5l0bR0vZJuA8BQX0WQqzvVOFaq1OyPpZUhY+vxT
wID6WU1MtMsZ6vh0bMkBIS3nhcaKbrlcZzwwWZjk45CDiAfrarrKeGXj2/szhK5SQr/2keAkz7h5
peMEfroa4Jm/zSbiVxTMwwGXYF+qhW5ww0BW9q4+SmGSX2mwKr/RhL0J557Lone8iO8EwoHhyYP6
UgUngD+UTLDwev8RVQ+XfyHIhp9uZ99msOE3HJYcdTSk8YclJI/KeKD6bRqR7Gb2jhJAyDe1yGGu
CVATONRr6cSwq0aW5uDaylMAQq+x0hSgqIezzCmoEPUZMTPSBWGg2w9upSZnfvvb/RNP/Jr1AZdf
+cwlRgXYqPvlJSmyEBt1YK82BtmvWzPkNj1M6zqNPbocME/XgG3SI2bYxcIn08SJaX1ob97G/VlG
Vmi8im3BXUWULi+RW/15NsMcmWm6qbifkw84K/mm2DgqcahG4U029urUUqTjo2Y7bLqClJZTegml
2bl7joyvkul08+qS0UnAvH7gCkImDPqZTTpelnbfldyBJyw8V2Sd6iztyvbh5scRD33+08dgfPpF
D4GRgMoCoZjpxQj/gRs9pJvwLLJPJ4JHISuMDdeS2Q0HZBN0F7PyhnMWf3aVfMt13fV2KfaJCObq
jZC2XL4vRDZA3X1RyuWxiyyV5ZHSGvro4ozVxc3uqk78ahu+85p4+NenErA/pXxtFVokNFs5T+Um
1nOdUwe2HqgMyJYXS8Akz5RCsjW9iS68L7ISmkLerZPqjILPutFcuOcxImZOdkVYqZRZdMlGXthq
Z3nPsIgTc2Ri8mRzxU4Tjdz0p7zAJSoRYMiWDO1h+J5fPUjvvY2sRcR4SDnKtMi3fWxmTZHz4wQ1
zNVsXfs1UNpoUz7aUWjdUVK59JqyV20iS0czjeD3dmL8z/1hMZ6kQMbpK+/GcyOjCDeVfChJ8JcP
PzpOMHiuZHzJz/pdjE0x9RczyyCbrvCqmOxDwYV3XoT7JbDTvgORUBcSafcJhcavl7FdaS5dl/On
ny89uBjxMbaFE+WpbK10n2ASUM9glgFAJUHBGb8H1hEUlb7FcQdTk97opwwsJsa9fZbnNBOnheo/
l676QhHP1+t3AZvvzDaDh8LJB4ddfcklqgroUQYlXMwIY2QmaB8YwFV95BYlr8XO0/N1xOBwS9AG
FvBAYlLS5xjeh+1jIsR4ShmFj8Kz8XCFFpU23zsf+G9VOcE53A+AkzmPVfdmFfqiD4DI/J3EzEqP
8LEYURG0UDBVv9X6QZAGlI5PYiFAM+oCXp/mChdv3VXQAofKoT9n3Z+v1He07pQ7xdGxBaF4M4PN
zeyQ8nVFP4D5Mnf+vSk5iBRvgV+hHG9dUKQBrRxkl3oJwNKNGaUOKBBdSxqc8yXscGMc3BdD8OOn
am+k/EQFSIrqIjnQ35iTvhruTm/GgrL3tYcx9eYjW3HbuhpgV+AXbBApc7m4w8MPeiujhSAvKD1d
G91J2e7ZE+l31uXzBSxV8bCWXmiGgBQWMZXPAA0e9WoIEXhjmo5DRa497jaALtw2KE+8L+ZcMSqG
9042dJt0urmCM/vETLfGuwhuhy/e0+TVkJ3isPAKGv7YoVP8j5z5wWr0xD1M/lfosqNZxa/YxG3A
rFwn5DeK3gM0mAh521KG7cHMlkyywqOum1zrrapoBbxUmoPk5Ax/ZnrHw+HqH+oSQGRyJgz+kD6r
99hFlSBSf7ndqFZ6XoGiJrYkJ4b0Dn2QX9L8RiUpSU9pPmQbNgjmRyQK6JsMz3RrStSOUGcKDx8i
kikpRZFxzacFyoV6Zvwkz/s56E5kGqIBhmSUPiiTB3Q/z49L8mEY0y6lnvEr/aOSSVyZGXuaJQmr
yI1A/tECmwRjRYYdpCytt2vo/xEyzjq31day/x13LKlCqdwVvDggiGuIYKMkN2bk9TOq0IZNs4TF
JF33TgCS/CsxYNa04XQtYSOmwA0CPqFFGhv0utODVQRc3Rwr+WuD2V78MYUOzO5+xdelfCBHHr3c
8ImRbe4PA7LGrEW3LFXoM8xMLMagD3wIc84cllkcLIelGwuM5e776L/kXL3QLH0s3e1NDjtOSGFV
Trr9ushs3G5bWDtl8QnlBsTt4+XATOw5B3HL8wBtkrCKhCeNRBx1xFYQEOWT8yaK3P94kAjgECSt
N5TVknn6jsRGKuU3mxPAbV9/dIZO2J2+y/3aZdEaGUA8UYUCxVctegy68WoMqnVS7XEKLQColY+W
bGeyu/juSA/3MI3p1GkEHvmFBTYPJjOvtPqu8182E0cTUIIGM92CsZT0gH8H+SVsl90jHvm02b/4
54q/xv33C6yMJFKebzSgKbHVgWyep1KssR520EkFfYsUfCru679d08LQJB9S1G9SbkpAmcTb+Gb8
ZQoBN7tXrKztBURJjN1i3K/1HNK5t9TKV3gcWRkX+BsDTbj55tB+i8Goi8LLvEQFGQaXCAUw4hRl
RZAUQ72/IKppZ18ao6qcPfxD6x4F/AsPpx2JhmbWWO3k7jehhwf1BEHJzhwUIk9EH7Dv9J2lrlS5
i1UxoJRtfceBlJe92ybiAVU8z6mRLYQ3sG2jiCGGCmJffwhcE+5ZLK8FVhsa6OsBVLmXfPAYxN0a
YaFjfS2z6axddJC2SfQVXp4ifS7csUHfS2oTHruzNo88jGYFtrRkf5mltUbVzcJKjaWSkleCYbME
39IfHG0OUUoYsDw/5qE+ldaQ/3tGZolTKI5Xy4p7eLkyYcDUkqY4lxgG6aymEUHSfM6ugClprrJM
D5JbnMRO+Xxi72X1Nv4ZM+oDsnwGfnl/FZ1ejKvfSgmyZcnb/nwrXgvKBaiF1VSNUOIVh3iQrN2C
sBDBPjeDSHU6YWHfEhOwfBTYOTVnab1oetsyeYRs6n0rV+96XYrKy2tGCCEz0gAVLCIEv3NV5qEF
uTwzDwDRGa+cw9kTyXlhI1/BbhCF8FZvPpWU7KfiS+d4ABw5eOgAzj6Ni49Vgwo17x7Ao5BAVc+m
byIxYXl6aMz//RzewbLejZfUn+Rc8p9/9DfSaSzNvht8HijBXDwIOQc7CjpnvZaolcYcdIdAVoSU
mnGLV1fGlcFHiOQBTgyctniU63hxgGq3Y9ZpqXW7C2uR55R6mxYngaqgpn9R2d0jraOFdL1TfCvM
CPWfyh3/eHMJ/FopbvIRspfjmDsOYUJLnQf+r5dLcPBkc8EGfVGUZ0bGJGQ9lfzLHj7da48GmUtT
hSyh8yjrWzu9wodFSOgHFy5F3KA3MwZV2tGB6Rs8HGMC0olqhSJ4cZAq7rL9si+QZmYyLcogsGS6
DxO68l+OhhzzSy36Z2lJgZiq51+cptugd+3jm6BVgISBdLieIimfrTwxnORvF9biNAcJQjvjOcUn
x0Aqin/L2EY9y6x3/VeYNaVxZTT/IJprASJjQ9fFvqbcJsZyhGkSYBGVAJmTMRyzHgZDdHqyRAdY
VVZ0/koGHj+DJv/dYTPQsLsodN00F0tXCpmdel9YBjAZ2j+r43jyAzKZHkTtA9sjQnoKJiKSoptb
2UFB0jY7KXZBCYz2CZh5dmX3Ce8ssbj/bMe2YlcRuxHwrPHb1/z/VmdqcCioOEzAPawv2kRIGTui
uQ8GAvZTfk6BP5Eq8STNBKzwsql1c2fFsFW9tx1wCq7hZFyugzPPrTIjQf/TWqzaq4liRg7phXUf
sFiLqrXcRuEIIxYk6HLq/ExsyhWwrd8iqAUgDLWMCDWe3yu6NV2P91qDk9Cshcdo+tfH2leKpsK0
seqr9sscy4rfzeJOwYq4grsL7ezjpqerJf6Ij9FaeOaeCJ/0V58CEHobeer+wZLbGzEztBNa5Z/4
j9DAXu2U2sB04P4JuK0+aY5yuaB/UISIoMgOGnZXbqbSwNvA8i68ngN9JgUlZU+G39skVpyjsp4t
Rf2psdbFqgXh9l2uLA3xt9ewmDcZCPYTVl2BayTha7IqlvKA5lWbgxPOjI9PTd37dGBJv92mL/ar
lNlR4HMhurtidH8M2AnWjiv58M34qfUso6roi5tL/mLzuZ227533gIZFUXO60m4lNvQu99PFrNj3
DgWpZLJ1HAKBpIX+61kA+osu6ocadq8UXH9w5QR6EZaEvrWbpyInCAGaKLSulaU31fm8/0m4tS6A
MqCVoFocI6qM7IHmJbc9efehQ6qzt4va6NOaAqp3yQcOdmDPk59DM/RzyhMlRbJrkGUcAg1fO1Jl
CbgM4cGHMKALSGXpExA/NCAlsuiR9xC10+2tM5tDFxHe3PzwqB2T0R0aQ6Nmx3nqC4N718EmuMfw
+8tlyc8E2GBBXOT3cG47CJwHDKa/HGYd8QBYY667kpJtUj3e2HdlILUkMkewISRXohfG/od9rtu3
rrQnV4awvqFDhLT+El66oyET4TIxbrGkqD6icH+jozwCWXoMe6SZtSNoYtbpW5FgkZP1HMBzfgS1
b5YIpc8DzpWHavxSQn7/PwIPO6UibTr1qJZMV51lfQj5sK91qufhrUF3VZGm+lBnV36Al2EoOGHO
bki0oizaEHRyTiB4LfuI+BA3c5KTcYU51IN8pItlTQd9b0GNj5xLclGgU5PmJrFDbrxRdQhxq2+G
ZQMZs2+KRUYv0uVIB1nZGdK0XwxM6D/7msxs4jchpCxsWkzMadP63n+jV/OETUT2dRdhTLLJE9g+
X1tqBAgVH7p7qU1cEgIdTsgt0W4zNTrk6DZFv6QiIe3J/vbM1mBoxJM3t3c6orMfFONo1A5olv/z
VAPX2y1RvW1oMPtccjyps4Cv31gZLXoHEiPHXdE/tUqKGWhN4uuoxNd1EwkROee3U+AzeogCHXxD
RyE+e6YfIGjiFvhDWcB/WB2RSxIXEI+zjQDBRt+zWOQaHNY2hnNOYMtQgGYv+tUyIsecTaHJmH00
2iqJYdCoOd8xxTu1cfl+V1bY6LDk0KTBYq2SF213jkelvHcwT61E3X6bisAfvHuWBvs3VtuEykOM
95+Kieq/tPEi2ea5BRoYL9gL64RoxcUw/X+Mp7hT3EyaQ6T/lBNHSef6mIsOFlDO2P7n7jHcqRAN
3jJSGHKvDPipAEBhZlKLl90ZrBuklz3ktrY4XmbmDum7u0aVmBx3UkSvWleHpDAzBWOkOzFbz1ka
EuWRLXS9u4BlwoYWk1BnbhXWMVcvKu03CVoSpgcmPSmGRTLj7TL5k8JekcNEAYY9fIC2Ia2O1/me
fW7qUfKVPuK8ErFAwk9soxsqMToTS312ubX9dTi3hvMUofEL57pYstNb7O30dpM+cBUOTFxgvIl4
hwBzReEzxgZgkumBKmuxSWzF14k0mJQV4c/eTC1aveYh+4luTWbVGFnTXOlZ4mKKzYqLb/d6aRMH
5Cz4Ax3TpYz2uoCgZu0eWTCmkm0GNwgPJlJupvNRSgMZr0woclDhOqMD+r0Ws9rK/wxdd8TIyTWT
oCvKwqPhWMk8YglA83fPpEr69XC3ik3HOXDYH+Mm+AV2dFm0dhU4pgBO+FpvrzHHAnkiIuVdmPT4
51wmoLcyPU/gq4gZ/Ri6wQBXnQoSS1R923Ue67jnkF43JMrzkunE94bkN7aL2UCkJqyPUHtzYh/i
B0j7QaiBnrDq3SnSc1StoICN2xusKxgqzEUj0vSF3WDJbwjG/h3KR92f9jrZZ8YHrIbH2B3h1/SU
uvFaIR9i+GkjMuF2zoyQYNKA48n3cHmw1uov2QwAdw0xrXOd2M21/W3yCoDh5H5VruMn/YSJJaTv
quP4e4x/QMtYj9c4kCa6/nefYIa/BGw7A3GFQLeFinZ3nL9i01E2V+J/l9eRNsLFfUb9MEOlrYva
hbYonWyRE52/Gd4HCIZ+sNTczg6QFPFPLRESjRmnXC0PDw5I5nV6ged6Oeey2/LQMo2k094LMDmd
K1flv57OkKSE3M06MRZiM3+nqe3snT5pYzmH+Rs2/tjkzWPj9EGgwJxBYEyelbxuwQYG3eD50C2n
UXKMQ7yF0KJPCUNOkdKG2aSNj0zRL5KHgYYpNW/lbRJSMgnzSqEgHkLY1A5/EhzB8OeZU6ua868U
ViaNR32EMh5OwFetSbvZi7gHz5/zYm1CAmA7uxNQVFjsvg5vJRCkBtnVCdHMExma1dW8G0+X6Ae5
QNL7wFWlrhlc6F6Kb+8uLEi1/TTOrpIfmhZvnPUrP12e1nhUhmE1mSX9Q6x/hKLMNSJSMSvArFPf
c6Z8jaGXYdJmUrhfMC3Smx2M3nCHx7VI5P1N3BuQY6TqFdDMKgxJP3Yf4tQ0wnQkhjnJY5yB3M+J
T2w2ZNPPFjwBKmmFMfZCGR1qsEOrJiKSK8H70jL7WWj+At8JUnWxDkSo1MPgw1IFlX3VgR+t26mc
w/Wq2r2egsASxA6jRzEiO7ofGzPQ/jFPsIghPh96tgACbErpgaXhlNARrVMGKtSWS/woJDwhml+l
nscMrQjgJM/7leZq2MmHf41lGoSqYBIsAno8XSOc8cemAUygYHM1MjZbSg26C2FHAcuTzew5zqCl
rm4+Cu2158z2szZNw7WOJcaAKXrkuydFRTW+V730jyBkzA+yW4sJJKIj+eVpAVatfvOa+i0KJjOO
rVsnfTb3TwhA9+nPyI3wqoUGB2M57JQNJw8lXwD/11X2mniadpXebxqkhlL3ze2OJUPNuBPAuVZd
Lb6cbuPZtyHwk5y02ahhu0ej1gOiij7462AcFLvKYdAOj/FRfbWaq6AkajXvwI/9Azl6Q/YMdmw1
hBJVE2oPn0WPbInocQYUffcpw8IyT8Z9rPHCqBENX7s6AtdIh1BuSimtKVikQMygp1YE8suMCToX
OPrMd2LaPqbBtOrVYEOJfw8MUz7UiVuZICGfaZQqavQ26rGvmruWb2Tdu8ui3PlAHd+MOIBUlz6f
yiYxvLqwyb0cuMDfUr2YfI5os4duWVwngR7ARE35Fl0DhYSw/Kq3QS8tXJqulvIiXaoqQPRpUMSu
5uQgA3ehos05jfscwiUmwsLucOpiocOg3yjJH/5Lc41zsjwAbYmJX2zxNOmf+/NqIcpvwG2KtbJV
6eaork88ds2oP4yzJj1OK4ots6PbxmfCBz/qJAMorvCHRoFZn7VSorK9ZFZQbjNXac/XuFF5lSWH
4ac47RnCTBqVa6HPP4CXdN/R9p6/E79T99YiPVJf3b17/zwm+GYR5c9gekGjqp29XbZx7DDfKT7V
HejIFbF3UJDm4/NKNlEX9UavJ0Qy5FwPrIyuHyzKJf2UWH43YyBwFVieH0t7JyRml7knyCmqnpHf
2tP/yYuv9VInvuMLu9jeFExQxNOpJIxFGO/Ic09rUkgZLbckzpEaaXVSL1qaGyBtPYy0wAA+s6g2
cJCnsGQSmDeBAjT7hFQm3uYR+ZC6Qi+PhOXXJej5/sOp/1CQDlxyWIiNLa9DcplewFArCcWVF4CG
ckqxYOQXe9r3DZ1bsb7i0HZD0aaASxRjODDDSSpt4FbuC5w449Nq7DTXGip4KRgOckOWvibO+eZb
ebalJnTYqH4xZwFADOG8wk722cHOCVIAlcNhka9588ZMmZQ1/loFUp1nU4BAoOOgmoC31EH4RonC
31pRE724AfIKmWlkfIGW4RHIy+o9Z4uYlkpMRbLmzcQcUizw+Pq6FDtSEjvvdcEE2qrqiA8pm4mi
wF1xDj3ym1iVRM8aNjllHOt/q+9IQJNwfQhYEZDY9TRAOfdjdoILLh/pKoLgSxApauYtwUXO8ebm
v1qDP+rzb5aumg2Vzj0RUVUhyVTbi3+KMxkZstEQWfN4afjPJiKBM3cj4+n6mQ5n2D0J2nHYBLHd
lWy79Q8Vnk8u2RoQVVmJ6Iz/+z1oe2jyiq4pmq1YWwd7oZOa6y3fRGRdr0eUZO0ikipLYl2y+GGO
cZIKGJmXlGLxaavmmrM5pqZM0j4GMfKmU4Ihmq/1IUNHleGutNa1vviN2B0VuYRix2JSyk7uGROG
EHzoTOr0m79Ybnze1mQAXCeZw1ntQyQKwlDNP7m7TBqhIdU5Y7XpjLcIH3qt08oP7+pp5gzhYO3i
8QjOwY7sqA4mf4CBg25HoF+9TTWelEaIojUVFy4URHH3d8XzHa4C362n1Rdj6Gf/3A9aTOxOWQXH
SUTIMqePXiHNLen01/0ADUmtL7Zr6Aa3nCLBioFJSfUma62Wy/XP2b2ZxwqKC9P7kufKf0O2XOg8
YRm1JCrI8sNHWnGTYkIoQ96wz1n8z3X987v8EwWNrBMb/Hr7IrtGAwfXQ/wLTjuGovX1L57kHvzr
jOvLCSb4BZD9k5ipLt/aVUi4o3GxQ5/XBuoc2MofFx8pTqd1pX/u379piafaS3QAb5i/fwbah0g7
VUiH5hsda7lVnn/UBaC5NMyX/dEhcGSrXq6BYNqZXgn7IqJlKWlFrmOa0IO0jNQmMh89vf/w/+nO
VrmT3SFtnUPo5dzLZYBcs5+qZ4+0Y6eBPRj629zL6GRNMJXGJtePyhL8r1KntUYVXbP3p/GaBl6F
9uB3oe6dklHHWodVGbnbdi/zPfGGkJF100lO7EyojmFroBwKW2niqYRMKpzPUxN5aGddv8+vzVQ4
KgQGYGeHkZxdqu+iRKbEoleD7VmMytKZzmtQCQvDmHhSwVGKtt3NeWk1bTnhBZ6oyKy1PTS2xAXY
Rs5c+qOHXlrgBElSIwK86SCRBS5654J3Aomw24/QnN+00h7u3QzKlURedf79Z7QVfBHIYi3Aavek
I63I0ZbICRAGbDCD9FbmfA+QWYiPEQCcPx6WCrKPxWmvLGA3cs0EslEfAhP3G49O1VHsR24/SsP0
wPCmW4fu/fPrYVB1I1s+wXfOWZhBt2uw4AEyclhwbGcxunaGHQ4UmcRaiBuW/XUg0bBZtt1LU/Zj
cIZtvmzDW5iGU05nL/JBPawYG4w18PSW3U/1OXVl3tDdsPrUozI9kgxwCLICdDOZL9j1Jv+tWBqy
TRO7FKI6YqRrqjHITPEcn4lJ8krlw5kzyOOnE4KPlk+COfklBR6SUChL58AbrYTC9fSUntjrjxSq
mMUZxov7MN5Z6CYcr2cuwORoIE1GwlXtUET83FQDsrDtIccChybVEs8/GD+dJUZTO4ctcbPcAVWT
IH6vkyQDsDJ//jdVVpF9Bz5cbFeC/VvHCPefx/dC9OOMeiMBCW+odnWKvj8dyzbikZkx6TrKAlUG
vXhQy5A9CDBubxiG9aN8gXjO5VmfU9Ka3cUIQNwVblX7RsIWGvyWMnlx3JLVKBdG2jiU62l5yPHy
EYQlw9W/wClRhMpM17joYP6ov40OTzHtYssMlbhOwTdcp4QukwsffdTq76l7ta17U8o21rq3BrRX
R0KSYZlrMwLVbUo00w81+d+/4DjpaHtZVjn8tWS3VARcHWLAvEYPVyn0rpPV1xvpek+FEE8oUoeW
Gf/Abfkfa4tYFxIwHZWz4oaLAzj/zISHgkMolbJRUoM/053iA5AR60eoaDhcu0ljp+9f/tgPPySj
KXER2Dgr0Edhdc0IC4AIKPKgMWrj2uYOzKBt/KOZQRiRxE/xZYzvFK646E0ji9n6nLHSuuez22ff
PZsHrbEPFgoY0UK4HS4MFmJMov0z54s2P7gq87jNJMulPaqfaEbNqGkDqL1reCnf2hO3RbYCRNFk
7PuO//tGWMHrsb6w3g4B2kvYYMloqSlfyvQhTq0yLgbWSzzqihw00ZT7ytlsfoPnoQavv0hkw8GS
Uc4Da2A6mEqIFPXhyPprSFlEoVq73yjXMjSDmYpyqo5xtt2hvkxdsXfU7DPEDKWE7yDc9jDZmrPl
D2cikjSIw1tTr6RLF45I3rbE1hyqLJA7jenCPi4iC7QrKxAfftYLdCjYCb0s7fDmClatDCvrCIki
+ZXp4QwXBMWWaycPjPXLNdfbAgjMbcfHizO0W4a+3QiI8nR/p8v8E6EpmbzUpcLpN+zijjlAiXfs
F6XOCoCOvfGsL/vbeSYVW8/A3TmakZyYPaLXzbEuOX+6CYwF8X5b/4MgPrv4YVr/1bTrnMrnFQFI
dNIh3ehDIDUQU3CGEPJVKg6Xv6RQt28v+LGuQ5udRNxLBHh2ACBaBlH9tDt4sAJhTjda7/oc9oAM
38WbpjDLE+hOuS8DTsIhfIY+IbSHNZVMs3Q2weOqI7aNXtP+GyC6cQhB4xSwFZ46ft+kVyn3WKog
nW5+Uh7Zkth35Zi30t3q9+K2b06OTrE/JSTcxCwE/oWQRNDobse9Ni8OaV8zbYc9mpM3q1VNbUbi
3NAYb4dO4uuFggihVIo+EuE0bI9C3SeVEqQlKrmmui9aTE9AeOpx0Hkwv4ZmXh4VEgDQoT3Acf/2
ThGKtbnwsE9FCmorUbTLqKWXcM+4A9iO2MhiezJiABnyVP9BB15CSVDZ+j5Jfxowj2ZqXGPDa6U1
7iKPLEVkOTEArWm7fHST/hYgt1qXOR19Vf9LX/ixD9FnDpBt12LY0W2OnXe2bqR6V2Pm5vyB9wTD
m9vdeAx/OuHuAT6Foc1FeaAADfgF4g0/WDFqI93t5iBi4bZUT7T/H0/dmHZf5vXioz+xsHBO0WOs
6iEgVelzK2M6s6pagBEAp0cld6Fpddl1zTKelUk0X0XQrVJWwBoGweDIZvvy3JdRkUbf7/LtZxT/
LZoLQ4Dci4nBgT69L7Ynxy6Rc6YLa+ilK0mcSCyY/PFMtzuMJ6W2Zz6o736aQ4bJlGLj/IiP+QQE
3e7ozyqNaNlkV3lo6tTAeaRwE+k5ZAXBI66gRpBajSsTuaGa7rDm46y+30niCgvnVfG09TfPG0aR
mkORvk4Halzet/mC9ZZ+2db6ST26DovjQpn4z3NLA9S3jsvNHuiETfgdkYJz4CG4D/6KouSmiNva
ubmYvosLa6DwlfXSo2KLEKV1IHuh6vYwrr8XFd1NhhgVxP/Yuxg/g7LKCtmEXpVD9tCkBLAXxXho
POU4dpuX3xqgd5VOH40lo8qjjBT+ddsTJOPosL7DIY+HTE5iP3mPbSthQdEIT/0HJR09nlJEmU5U
QAbFthCZmebg8envdobx8NMGB6BeTBVBqN28tzGtlHWKCwiFfXiGJsZuvPyFTdOsgW7uttdVPrl0
BGQS0OUtkscM5V/M90bcRsHCwq18hixkJhECvpCDCxxvOqpTWUWU+8UUGK69+wYYsdIL3QnOf8rG
riOUst6oYAiDXGzwBN29Mz0KaDzS7TsowjueDpaGhz/6+4Ay0l3c1I4qR0NRQ7eUdhOzo1oBDfv3
vWcR3QRMNcJ7jxL3tdAdVSJc3jQFeCfGUPrDT3ksCkBtso6jS+Uv6uvxMdZBKvezCtb3ejtJkx27
Q17EdZR/KmYkFN+J78xmNk4UZexJuO0w7FTldUsoz8blXx9MXihVPEMlewrAMPmJS1Pm7gUyMMAb
B8EMpZ+d4Hg+WsnngT518ey9pZ0vHgbSJhL/4+J2NNJb7UHGPIp6T5RNPsWpwrWr4Lcj3WugrvUD
v6RVTc5mM7GdtQLTPN0sVROQL4agXbzH6uxI5NLKr8BnvsWd3/qXXPRXkp4eED1v+kIj5kqOBKCR
K5iTGBVNdWb/iHYMCZwz+yWTU+6GRoiYNVAsb12ACI7SvqF/olOwPYs/WUXQLP67T1zlr7aiEDkC
lZIstIT6grBOyjlG/MyrK+BLgwspvLzbZnxaNWz+pmSwpsVadI95UnL5aCrYL7g/vYMkU/XUfn/S
JGLsCm55cRSXowuXt3oQtmJXDSX5KUASz11JU3cjm22Ao60w472yX3y9WZt8Jaa6aeMVmVmdk/d0
CUFO0fKrqLgb67noOhIw3fcGKQIrp8iW0t77+JnKN89odzXdjSQMk2sKTUI0F64yAqhZAJjXKcXq
3GBTD55Mm3nzJe1i6deC4Mlz/nQONGXFkJMk3+GdeJGhBQQ7he8Yp8W02eJ3vCBINa5aUHOrcTwm
qbbN1jOpl2ER/oauZrzEn7BZmKrw790IRvIn8uBZg+ZCDPpQtz5kdyjNYxUiZ2t4jOT3JRtS7gAc
9g2oVHARp9+0kipN2ELkvAUkkZNY2jZ0llHSFQrcO9Vg8di4aJQYyaMQfzsUQj1wI6ZPhwoMLx6r
dGzCQ1uJrXUTv1v2cuU7ucTW8tvJvLwkfbGReRc053GLj+nloS+tKJ1YQfbhglNt5cocPH1ezZHk
EP0Vf92jE6Wn+7XxOGxMNTuD0pZdNkN1D+K6AFyLpYqimaOJ5OWRLVdC9+OYynHmfNczUE7NrEJV
y43cY/+lIXJgRVtfSR/mzrW5NgD9gpHrNVlJgNSW3yvISv9ONuBAu8aQEXnZSyjQu6w2SXKZKyKJ
dC71dhK6GZpcmf8zkFZUQQaTTLS6EFeofX+TwwEeJ6CRE/DuvlqQLLIEkllg49MlQfDHBTDZ0W3Y
HiW+flLaTJCzJTsV1NdN1Z90g7ReeYLwjmC1Fvjt3SqQ0NicZA16wYFKe19UfqgTm8owzGgQ1q9A
wiO1YbL2mwVB7HBNoZCYD5qmUn5GJHrBbwPS2GtPFXDkKKZjzgfPKmUyJJGyj7XwCnzFHV4l46gP
SaLd5r5vOe72tRVFjKyEP0xxRlivilC78xKJUZiUAEb0r/lT/kCjjYNOBVJrzmU65IbZvMRH7OPw
bfBkwC4bGl6R+ddYn7f4rbso8kRkUgPlULiT2pw/pqOiKVgtjDIa++C0n/5MwAvfdmnbQ7eHSZAz
P6/DT7GTlM5G6yzhIVn3IPsqMefwIUQPC3br2ez1DbipuuiJxA+URmNMDWIL8g6AkBsDYumOVwng
t1FTxyJgWCA0VxrTYGC3AoXo3VAW2j3V6kNHCHmRMc3/ybqOQV4ai9GLDtWy4FlQdEX5IIiAXSZS
gigBFmf/WgKRDtwW7S8R5SE6S79EuMCHCrLq3ciTYUb8CM2BDf/GFkgX+ps2wxDNZ8/a3+huTLX4
eXam5vb8shEGVaC8t03wj6fPmZuPBY21PN7Kj8WAwdNcDB8ApFuu11Ukjtbubr2IFZogRzmopHPK
Rhqc6gQP7c90QkuyFmmzxOElXHrtpJ3d5asad9hsdUY+blkLWzMkKZshQ0QL8XumJOr3Tdq3/SR6
L3b3nkCsaJJJ7XklkAeppnozSjWrn9STHXOov2kkJO26TuquNUKMwU8fI7DJAxUfHk0gI4gB2Xt9
TJJ1jF9IPzCYzoYebqBVkBGKFGG1hsGpQveTjvPAqs2iuJRNoMGEK3IYlClk0hpBOIbivFN6XNSx
pmTNjwe0aDdCBg7ybCLVVwuTnQk3IF3sWmRy7S+VB0Eg3LyT0LGI7pycMK5g4g121rpGKa1A6Y0n
fg04bppBdmygOv1E1DyWC4qRl7KlTrZhwZSe1/+H3/yZEaohiQ/0NEFTIwXwcINwB9FdDYD1JYQy
/9gW16KGxHnbB/fMiKkDSEDDd8t2H0vDdvXzFIoyGEGZ/kSizUTkCnwAlU/SFsaqHl/Ic2Q90wOD
K/Mtm1wWS0MeoKvteMwhf+ESUFHpzqkFCDqP9anZRRPlVKrF2ajYzJoO5vU2y9XGOdsCJ9f9RKX+
tn2XSpDHP4uDNjhWibP8AXiK/omfM1lQ+Npbhbp0k1H0hMLtkRWsPC+z2safHniyg7cG+KIlvz23
6gb/HRbe1+0sTtuUZo+BKZYZh9MTGr3PD/38CCVbRbQV5uQU7WfLU3eJg88OyGFEWT12/3pBLtSI
E27O8zhCvSHlCIpaMcAkhXRCkMUPJc8xxnqx0Ya6XzRZF2ykUcZT7WnBeVN+7BvCGAGQ9vgNeUWA
+DblkYJIjG/+VqKSUpbJ6ulRP/gJvFv3JLvp8OjCUkwgtnYkTChQW/Yyl6g18mwYRvNagIjtEkIc
/qEUwF41waSxwWeNSrfP51IkOrvvNjiTdeV/t6vs4cWqIpqc/b2twVw41YSRVcixcMjhvHyLwxhR
OLK98pXXn46Cgq4NyF5fNS7U9ZR3d3B/W0yHW8Yud9555mEezFoFiL0wfjAhhKSdxq2TuMh3Gu+4
Zm81VMAGTpOczCUKuJIS0Brn0bnA0Z2eueGYRA9r5kPZJfib3/Aai4k6Yc+1czmwJwMa4e4rqysT
sbdxG7E4EcqajmJLrsmMLSOx8KYjOF98avAXYMJ6SPQFnouuzhZdNRQ4MvtH7NRFBT2y2Iwdc13j
tkGtxDR/4R8H9JuyYopq8W4dsd69osCxX1FefjN1GIq3SARQ6CA/n+ML+YE34iN7m3k4b4cx63qz
TN1vs7TzVU9/xdnKt5fHmR4+sKXsgjpwfI5ob0q8p1clGKhxWSub1jtFn62EGHbtHUnwWUR9hJGL
Y4VlN+KzVqi0TsF8DYBjtrLHmdvKz4qs39IPwNMzRk7t1rvXc81oq4sAC0ZIVukjNZegLMGVeyaU
6t377PJVQ314YgD94JvTplWTCokr9ndBzgIEaG7MHbTW5hBS3tygDJQD4yyWbLnvWXHnchYwJ6wa
VwvgOLwTHG3Tg3WlCjqUCYZqWT9WZ4Z0CPMtJeSUZRZ4+Rgb11dn7RFuWNiTDSZFRdUhxjEd7hb4
DOxxK6ONxe6lVOsXyCVuCEDMfTvaPyrtClCV+HHmW8Tp62U7AulKQiQ/iy/AgdFTA3D8PtAYv2zP
Oo0n8Baeezj72tUBK5sa9Awda3NjdoXy5WTVg9VSu4KIL3dWtxz1tgPqekAdPllLy6sOGyig4qaW
iz+hlFUyCZHOLr5WArJVlLmpypXMn+1RSZGeDNUL8MgDyzKKBM3BCrKQ7QkL9pw41jIH8pRJ+Oj3
qNB7k6PRFsZnud1I6jPzwFrW8VjZZDH8cIxuExTTpUBAXmG6wTZMwRUlbAlzLZ9WqxVboeAQ4S16
otXu6X43ETAWu6FodSRbX5k0cG7oTFflcI+ukeMda9zBe1mTd26vQZ3E2ModRNaXxTQ/ZkwmozXc
mza+L20KIjlha4SYA5JE6ONp7GJi8hVt1fCaT35vj5/qzH6r7mWtwm4t0zortlQitK7/QpmIkAen
uKkUb27gBJ2GRsFVeJhTdgQTkT/gQvSU8ZYyxdz/vu70+8dAH1xQZhZlGD3I4gz6gTLrcz9aWhl/
DjhQeyy5vczXrc4LOORXCi0UwECbjK4uC5miIgJrsMojYPnUM0/xkpHcV91uhay889+xNXMb1d4O
l5ty2/vvikAnuJr9pGM7ZgrvW2NgiccUAx1bhiy0Q+Zx8B77uTp5UnIm5gBG/NKoZN+v0pSP4twI
LKe3vNRyYsMocPTR+pqeNyZJgc2aK2kXLjB6ubHi2U5YHl1OGqc3WtD25rToY2d2TWK3VnRmChjC
vXMopvw9G/CVI6l+pM2M0UZ6ZG+8H3mvVnX5OrSQaH+3pc6d9qqiZbOnAnQrIBDKG5Rh0mZNQ4mI
VMpeumE1+Plr0lAbB9kyubp4eD2grjK0ujXsY3OFSbv/FEnggCW8uuRo3dd3s/ZZkpYn79BHe4GC
l2Smb6tAunrHcOrTAhbLeHrpi/eV+aCtI95dP5yZj7BE4j7RBGiyVKp+aN35H8k97OqoSN62JHSa
4YqNbhPdi9R4wJ9vNJMQc8tEje2XnAoQ87PoBbrHcIqE6twwcZHHw0vHdkU9uetWVEa/aoSAsznK
h34LtAUyGZSZbkp+6Rgovt+L6VhN7w6InhNr+acvmyy/HnWoMvItxlDg0wE5S4/oHjQwnKTEiZT9
s+lmYdMdEm4lb5u79LQA/f5mXYi6McD3VEKzLApuiFAXqIzpPotG2+3sSG1dgpX1BOHJx/QuU79S
XQ2iF3OyVc3sQPFKk71pz8ObKjZoXXF/R3I+Kxfkdts0cEJijMow1S34q4cI6LEqEvGScpopdqnZ
AXZLWWjyjXR7E5McY8hL+G0yUYXRyJ9QUuNmkXPVcy8FmeZAorr/CVedjkta5POpQb5p9s+RriNN
u/ZLfX40NQVI2u6ggw+QXZWUgAz/bsGR338IDMqoyvKIkO6eBFIUtzX9qn8P8DWMoYahGlyncQFK
Y3M7PQAPzTTAHOLba1m//OzTMOGpUghF/r7X5LJVPySwYWcXBv+GwqiV1dP4PoCW8vJPgH7Z580t
f423Pp76boO4pVoZ3Jq4VJGUGcSH7UxXWcjzzWpP8KWCJ9K0lA1tKuD3329J2qB7YHU1+FaiVLeH
iUz6fJfCWb2aiQqCLze7qVZuy3XcqLKkBzYxEp88ZDeO7H3QfMT4Jpi0ntBPr/eLIK4RAWEtHdsT
/QdR6ziNiVFdTOr0bqSckQkYcaEMaYITD2LmT3a0vv7P2DTTrA2Igx7AQAushjWDowf8nLmiR8RO
kUZnONzBMkebtfGVmn3mJDq6rcWOchEZ9iOaUZBBaEYc5K1/8c8Qam+vTbEOir3fQpRLMepH60Ft
kVOBSBecmofrC9diuHjzAg0/ZEObyVslH3UX/lTGJOELPd6xl7SxeTrU2pqw65TZqqUln40uG4qk
SJWddZMcS+Wv/XXtla4UbkpwTtjKZpi3G1Q2WdGYS54871HRq3/0/RgCYGV8BK6OtdJ4GQQbk93W
42weMLOeXqnTw0hZReq/8gWVh2wlT6yi57C0TM7J1KLQk2pDnlmAnS67y64OD9hsEY49ELoJLzjY
yvs5bZnHBAfuNGGABF4ef0F/NwVgi3nxvt6RmgJEPePLlnDm4KdaH+Wl8MqrVesx1WoO9IrR0Ikv
yTNeF3qieHg0TcTYWUFHzt3hGx4SL/Nhen0B/AcJwDl9Z+qzMxikjbgLJJHp0XHjvtu/VCIAH54R
TnKBhquVTAtMXXR304Sza0GLQ28L2aKpQ6nSxluyt3G+atxAheYt3U6w2/PkDqUI9qGZt69SOL2Z
LeWPH/0hUQfCtQWZgc7ZeoYHjQ4UhyjJIngk9Sr5NICdV2radkWlHumPB+0G6j9Fa2ivHS22+pnO
1XNi8wGdCWnpDi0d9FSo88Tryz74WlCc17z6TLCT3cOj/B3E6Tbu5mEdHh+TbzbNi8rVDL/brEi9
JvXVyI2RZP4uZneb4b00MIwLOFe1OHVzv1tpUZ25x/wpRpyif9DCrmRv07jfCQuEJOXnI9G/on3Q
/4tX2CGf9ZZBAlmDymEZkR1XZAnmyjmrmt1TmCjbj4U6rxy06vWjjystbvdn+/ZFacRIFb8XOEwf
mcyNRa4Qrd8rZE+75NT+uV351udzVGVL9eVW7MyWnIyZcUSwSZbJXhgeoDwzVIkxNzIhY7tCjliO
RimCXrauF2P9S4sAw178HeoAaZ6j06gp2WMBUuSqUCQbxcW2UIVe/uQjMr/SzpMeNPp6lESZCp6L
z1ILpvdIzazu+GVxeBjb5ajxKaaN6U62X+V+3dtTyZ/k7F3sLYzHITmFEIzmQMTujcl3E8Q+RjSV
il6stnkulsKvRPQ5lxlG3o8iJmXNJabgH+AN5lF1e6m6W1FNEPXlmLtZZ8aCTYOYFVOiVc+AKazk
SOW3IETfXdhhfCdMAem+CE4aDwo2pYnHTNtAPt2crR309wt7KrC9s4nnDz3vCkTc4KfyzhfodOim
NwilK23HzEj3aE/KgWKUnf191Ut1AP1mJWDSQAFmVRy6JQ3TAE11DEe5IIeaEnRYrX3AlNoieaOP
DbVG2xz7lHPDotX6Zp6RZvyLrT26ydgJSlKMXBwFvWxXfEka8ierMwHPGsOSkwiQQCuICoMUQUMl
o8ZN0EIPav9TMynBurZkmrBOAM4Tvkp7ptYInraU+DgMoonUPjdq6/7nPjm1OzrcdhYe/U/plU9T
AjJWqpApmA9gn1tcmzlxWdlBVzXUkQhhY00mzGX5NSdt6ebM4RVDRJRx/pdw+y6drK3H/FWyqXWj
TcxoxPb6oKq02IJ71ZsT3xIcksw6xj0n4+EgqzCsvb+Y7X5Heyd0p9f4R3dL10zcNwRPHPrcGQ8e
iXpw0mykegMCMpkSAqQ62SiNHK8iPZGis2LKCruOie3YK5U3esmZ+KoMrx6qN8VPbyh0V/pkjKS4
M4eviL1YR0XNaEJPb5tQD6wBgHM5Gp66MXs1HMTQVqpw6HhvsAHhl3sc1chUL01g7OzbWsJN89mw
LMUaX6Njf0DzYc2IVppz8YbegeizSuBDhyGjUBj2ueD+SMUClrJfvJPzkWHs2V1zkzCn7zkKXH17
AYwg1dtaXWCkeHv/JwbqS9z4mIMRJOrwi9ezdMbgA21eR9qjr0zHIKr0kPKzb21QZ9Do7qciRdiO
Eskofn7S/Cnf1oTw+ukpHQKW0AqYU0XZxV7pqCmIr1FV4bQzDiAtpVhRFkKayX+EkQgN3AxqXEoq
ylxJdxQee5e1diTMt8LqNt0ObvIXuKQd8h6SI/P0Vh/8nSnILmGO796TCJbCHQSWpY48vBc9Px21
pyt5GjU38P07zcWy+uUgG+vSW6hnvKs7OVkuIbF5j+DCzlut7H0u1WkEbwdereVWe6v6vkW8sgVf
rte2stVyyqucjTYqzlnpzMOP45voMfYoSAcM5ftXEStP/nL6rUzJQs3Wk1m+5r2eKB1mZyhmjWqB
iu4AMj312YWYDB/PEvrNWawAQkL9CI7rdPXVRIPMXhLOp8ae2RT69laxDvmI2xEDz1UXOnnvkYDk
/Mmpst5SECjooc+1HQnMio0b3QEBgs7hy8HQ56RIjuZalqoGheL8sQLrlOxRH0lZ9J+nnMtST57v
58w1lIm7ltD2/A1bMteE3BtCaDY0ouNoO3Rg+n/7PX5AYEf7vasuAJdVnf+AbQ2oAuqHu4AzD75T
qvTXXw/8NHcoJ3wmgVycuO4P9MtzAOMy/X/kzmLOvML81bVJV66x+7nhT3n0n7xQFrPQ7iUNNS8v
DXU93BVoxCL8R1RuLL92TAN4CAmVnYMa6qKtLzJDM3okYpJyJFW3UqZlXVWcPdBT95iHdweqzhwh
ORB7SK2gNYDJjirXMrO34nDOZzOK1vc1ldpEAHUnayYYAqYJ7m+qvRU5qSeSaLr0src7qgG68FVy
9xtpvMBRtQvSqBfX2O66EDBsWIZUFmSuxBvRWJTwK3lOp/9o/Y1BLrVhx2W+Y6kDl69lsLalmar1
plysmGtfdTueVpPueCDHhk/sXLWB01WCMVOXR3AAR8s0YUJSqa3I1nmaqeCYF4aLH4RJGUH/Sp4P
4ttbmNkq34gAId1dfL5D2+8kWIse6dXG/PICctp4OjnQjrpkghmcgkMKtxgCGFZ2GX5+2Ate7bAi
uy2eYCERmVKbFBUEqR4ohyZD+XRh4DqlM3r8F0ogxG4BNAvEu01Z4gxttRcrHTYitE0Nz7ZYS9Sa
z/EFS0v2XZODJoi2wcDEomDG1FxSuiMH/TRZndmdTmVHkNhm/JFftYGi8StAuhUWh0A2k+uMe7Zl
zEHmsP611AJRuUVBGH4sPKDxsd7AfiDahYO/NuSlQpLp/G99207KK3dYJvvHK3TH1Sn+ZeA938h1
xDAumrExPum89qFDqY2RyuImFSp9EfAH79KcKKqAyuYsqNAqFQ14Gv2MZreqmqFMeI9S+XosFefP
m1WG6V4HWK0IIv91C79ciEHCdnUEObeIXjDhpLupzjAAXTLjcOdl879uTpj5x9T4GJ33C9UdlZG2
Eaqj2r35LSfvYcLd3GAj6Unfl8YWULOPq28lhhfcbLlIlnp3JcxrpRDPrqyRRNi6SAkXcRjrzGBq
dn1+iB6wCfp7X27jy56md8gBnTSlrJPxtDs2qdPT0BW/JgKvREiQzoYRocBlVdHeEEF+V53PicMU
unn1u/l27dtU0VZ1tVkmv4wGnUg2pzu8b6GfYZKw+IGf/NMN4NtsqUoXVXqDzh4RRfipFqOwYQx2
3jSsGDrP3/to46/d7Qc5mJS2Q1YMdTdNqvuewNBCsaN1OjA0YVntUQqDVzba5D9UDRmDAFVIg8zw
zbFJwRZVcg/gc8Lfd5wDlxjKBZYTuI/0ir+vQaEQVFaxoB+gXH3go+bYfnAseavgQOGixkRKoEPV
xnql3yJY5Ie7pQkkXY98Sxkoz6r+p422vo15NHDxs5K3CbWXBCC7bUIxbLr/xeiFeqcvhl/osFzO
+pEy8IL5sQtGVuFUB15nQxrCt7G2Q8eedyO40F8X6Up/QRgY7wAQbyjfu1YAJnEwbuRCJLsmdmOt
EIXJH5atWAeRJm3VhJFI8wYWDwPECCeyIlVrdrEzDj6t5W5GHHW5x1tLYtXmptZ/0ARhsP4uojD7
ItRfR5PUrnQZnRMRVu3efKSPeI3YIH5XdZwdHusxLAefFVriH8Vox11EKktmZsvIgQeans105p9A
LLpDghpaz+04sIbg179yaqwTCuNWZsCqiPhvPtExqyIYmxr8QcSwJb3L/M9fkAQ8LB674WdEKTE8
LqL5CJMEJtnbgdBoNWnOK+d7NtYb6KXLMrvwXWR7lWfjj85FeNFtyyDQrYoBfWzGr9zJK2ttonem
AJTQYjHyrnDLDkVlnCfRHKM5nror9e9pCuZ4n5xl9DjfXGEy8Td5OAAgllznuZQnSupeUhXlKWGP
6zcRLs9xc4OResZU3xgYznk22yJquHm8HRtHMLPf4I6Tjc1VmqDLBz8BgDu4Y5xu7z/ecccWbnGK
3HBdFYwi8lPuRkddsyZeX6yRCWxSXu/3h6+LMCbEaK18iiGwNsasTgecLy3NqfMqgEkjaVovpBY0
3VF9tzLKCgnpfWr9lZcmYFbaPQYcFW0O6rkXrShU1JGc5JLoKzxWNzP+qmhXJD2jaCMwL70e1lv8
SMWx9zNeiU4L39XSezfPPvVd8au4fsj2R+sZ3va3z2AfPKB9wzjuaDszv6P8mJe5lXuekvJMEeXZ
9g04SidSRlZm9f/VgYhyEQX0zrA+ktTiwHlOuxRR4aYa1ggvcBuV8l0bBOr6y93/2KOJ7ooO21cm
dbe5CcagoJcbYLiD45nY/nGAhjK1gZMfLgcu4btxijEXMcay6KzGgjTmCo7AJQeXITlTjbnTY758
uZABBj/dCrTikxUonzPKGQq6gim7He7O+iuqkQJIYVTb+But7ffIiZejHsJNHQ36ofH7qbWlmLfS
WB9kxZpLqF3XpEkw2pKiCNf1GLW2/oWsVClmXSnGjhzWvvCey9Gunsb41Oj+9ILM51cwpGXPqP8b
/UqIYpsJ5xEo3N1eQ74GAF21KPfi5gJ90IuAIzcTEgNMXlJ3bSb56PUnM4Q27h3lC9MSlRerDMjm
tuWmnjjSo2e5W4KMcaOd8fCRFTbFkwlldAsaXikpS3FunzkukDIZNkoxJRskrLKFIAKUlQkEVf7Y
ilmf0XdN9vUQIZZiBlJaa/7Y6Lkcr4z9ifz+vs7qWGFme/CJskIRfmA02tqTv13Y180jOVBI4x7n
XlIixPzxtcCZN6S1d+ICeGnxEjkT2ZCe8UssgnjNy3JUJr7vQWPPHCfqza4edQC9eelfLR7B3nk+
S2BEgjXuQ+teU/uJSbHe7pSJPTkObdUJ/B1RAI+GWO9BedLKJiCo+x9udXPpwFIAI/SDs6UDoymF
pp6RDVqG+CVGYHA3Qg0xPQ1x18V00Je50h3nU9HmJpr3nTpsCU2goZ5tR42njNFrlPxmz/tIN+2u
A989vVRrJZsklCmP/O9R+HAWDTedSR/bHEMv9bjgK9SOpQd55Q799pFsUQkDotnapvI7JYsjT4Sb
oP7t1xT0N87H5lmDuM3yAgeOfCbvV6gij05s0iVXUpdbh68bx7MQLIJnNp3W3ICdEpTykrgFg7KX
iViHN46JFuTWk9FY/QFXczYhEBi/VfYF6JIqyQ8TdxCfEKh7bTcZM/OLkyXJg++zx7IXTBvSuvuv
akiPjFIcBqkqRAFve8C7NDmNZlSirrCJz9YGwiCTcNE+2LY0jCfjWtPvl05NYTey3reFTBa9qxuq
d5D6BIs0VXf+tr10hhiCnRHZuRv4htMGs1HviRf+mtGfLCtmw2g+YK7/78UJ2mQ61ieSeWeRjHVC
Evy3VqlRNfBVlccqRSdULmi2rfjHRkbRRBQwWDp9eWjPHaNOg57tp++u9W18x/Np8xV2IaoBw5L6
3X2DQQEX0dIGzY+hBTUHzPRxl/VFk0QrZQ2qKyagnnmCUSug6Fhph922EZOp9UxCItkVa7vmF9oq
y9Yjd3xsAEEqY46y8RpEyi8NCvh9KUD5pZ2b4BZ2oD22o4aEpp3yCJzFe0oL7mFlaPG9zFfcT4NY
AmfMH8ovzO/ve2zfOmt6fbK8+6D2HaaNs3hqQi2FJ7ZhXZll3OcOkUzJxs/nEOT7r+LUKW3QMXGA
PKvlPSFo5vKtQvSatgmORaLB0O6FYsDX/LjnUel8fycfDsSPB8FC49iUKoL8ztX3f8aEwfZNiRQm
hsn6S0/opiFsp6qJGQDbIhSEcEOwcMt3yN20OToc6d6xreh1FBHonLeiCHghnKWDWWkvIwsfN9tI
H+UWJsry/PYl2vZfhLVA3Nk3+0TG5FBKU8OrEOaQry3yFaZl9C7/CBpdIXU7AKSChl/3whzGb9v6
XL1MC8OUPIxUDKLQfcpkdWkY03qUsnlMf15eAW6gqKWkdCZChIUMELOsN0W/q0w7puidKnUTSeSc
AaORvBQb+mnybnjClJ6qXLy5uSFz4fraW00uQTBCS2K+i4apsAuB2giOflXlbc0QpcTYNHBMOBeK
MSoshbCRLfzqObPN1U0lExSKa2wiPIfWjDQDMAZsjCa5r+Va2akpcMxm0ebAGzvdcjhJXVeLDib2
vyEvxUXX6ZBSO937qOm9O0Vi6z9b+aIkgdDpOEFLfK964U9vXr7txhy2wjg41+5NYRzYEneJT7jf
ameV3XHX6adrOG5XLOdmcgYpyhOiqdg7Httvtw2KNL4ZGLOERWgd8IAMvOf9TqzXix5AkBfACN2Z
EOzR1AKcgYzHxp0p4Ruu9XhWXqdWIDxwIa2qpSYkRCgLRSzUB2dN9+Jt4BemMXmyZDFzqHAu03bt
CF/0pKipKIvkNTK5UDxLneqtrR3ZJxNJ63By0A0RemE2y3hxGJ3DM/K+iSzIQKDANUy7pSj8wzJ9
7cbc3YOg+sXlJsxkP69hmyOR/cP31CFk3m6ox2JUn/fd7myxhjQWgG9elBmObPMdCf4xNJXr6j95
BwvglKmwMURw8QvNKzEife6bng8TtFfNMV4kh+5lqTfx4lqoPGYv35rE9F0Q7WomA5oQtK5/sEJH
17q81nhpBUT1zWir/UzG4SiCX2lfVV4ZVc8rSFOFy+FZwi0c4VX7YZ2DXg4MDsnOMd/IOsjywB8v
ePQsDuO4Xk9zO3AhpkiYVh495bXWbh824u92N0h0hh/za87bHSQzooSXkb8HC8SB9HpEaSbFtr+T
HnndMK1oZS681yaKRM5h77k5E8JFR99zV+0832Q/84xH8zTDuGZtZUv5uobQ37iAkhY9KAJG8/Yw
iYw03WMCnIGvPioMwcb4Jq0f1ilKu6fQOvX6bzdQqNhZdICvDGKiiR8LzNH8wnPtkeh6NgVoWrHt
lYaASLjbdcqZQ9GVFvzskqzDQR1DK9tya/0Fjhvbj6WxId0wz2zPcyaVNuGu189xjl3UlyxidOhd
H1HZ3PFT6Pj6sh1GT3+Rg2GKT/eqsevSUaaEGIpQAq1uZ9umRxL4J/xDSD3XR46GNGeTcoqqd/rJ
HFHOhTUzY72iCZt1DMDnmuNIW56TlLm/QS6Iy1D54bmpgjYfDrUPcMvcQJHiQQer8tvpS0Ev/olr
ymlUlU3P/b81rasvh1paFN650bZskceoPXkMsKYcXc5JKHHeGRp98wPsFG6sFxkKaOswFR/+GkF4
RJoESEdSimm54mqPIZj5KLctGPkBYnbHGRAtPV0EtrWjshlwGdC2hYLK1awveQzMlldGhaEWaXfI
jMvLIZ93ulsc7q+NAej/l6AEELr4Ddw82V/KZsSLErFwv9mUtVF19MICQO74nrTH7KWnAoVk4XGy
2vLOOJTuyWxORGF1IvkO+OqOr74G8EPkqOWDV1SOqer2Dit/8zVC6VpphN3MBmzAWVH2i5zaCFyZ
xh+DbmDIGJkvat/i3DVkOc+tescaMXFDWeqbxmmXO/yqNptw+yUyGGXvpiK5QlT1E1iZInEUS7ZA
PVMqSYD0W9LdtNVxiwzzh40Ia/aP+E1c5iXg842Wvk3pnadiAgrrZIvj36iG/KrjJQdQFeVdS5SE
QUPwA2TqObeJdrMM7gqWszczAjb0SAjqH00cyOgTZ68zcn3vGCPxyGzdl4eT6owKdVtTpCq8W0Xr
zA1y9vu+eJlins2n3KI77UEGjmriccica9tq+hRF+YMjYG2LTxnLdFLV1QnT7r5JNjwJGLYsszoQ
8tsBGhvhGdJ6QAwrXF6EVeLIrwNYiIK8SwjPE7fqM8SxXF6SCjZKI5PNuxIaV7y267Mbek7GyTmr
vJoReGubx7OyKc2BIpXGSTn9BoaFfj/+xjYpHTGKMxuj7suLdbyQQMEw66LWreYYJF4Y7FRW4h9n
UnbrLxEZHnj7Gp+Za2C47L6ONJF3Fqe2n/DHuQWneDve9lTqeG70Ujr7xsfpCtWdVWQFl2HVf8GP
hICBQ+Gv70rn+G8EhTgsRIFSh0bG1caVALO9uajEsg+EECRo6Q5FKb6+ZTJPP0J9hf66V/JTovNC
p0Z+DYFxJIiXPevkB+bVNnxkbCRed3lsVGMV4Y0Magkq3UxDwRFPa2T2+fN9HZoWZypnjCG9bwbV
55J4pilsGF/ArBIuNzwv1D48uCRArQAyLHBAaCdnmTEj+jfNbb4m+vGREqq+g6dKKJjvb4Rgs69a
/8XwG9LDkISlaSdBbxUjsu0K9dBStVkmJMFXZEiO9NwpQep4twsoAFw9ee35BXxdCeML2vyN+Svn
G37WgAi5lDVnxqUvx2fGT0ulzMJ/7UhLElUAe7uJHkxNXwBGPCssTNAshfZwKHgvkGDRAzY490gl
4JzLQsf5LT1lug8oCfB0h99WOttN6tFWSxdncxhTqrLIKXg1lNIzfb4viBLmmxfw0LfiKLsGJQM5
MVhNO8pflOc/+bakFa7chEhdbTZSKHblSMJ1MQ22rw0vA6eXekQ/SX25241VuOgBk/ZB8Kdrf+at
gXZsamHx4wL5reNNAw5OC9GchNidb3Q+6a8OM23NCDjE4tYepe1gE0CJKKrKqW/4hk3tbKSmjgpQ
ml+WlW1hvwQdSr2SQdHoLt76qf/LUEIgwqnTXyNbre7mYwlreQkU/h7gg624Rct1yYi4tqtkuIpd
omXKINA2rSDp2cPfM2mFNOromKj+Qq3tItS8GM149Nx15zqeXGeM6OkG0ka6Fs7TJkbZ1j553mq6
VAsBiEqqv0pNk6mZkduLeWFT0wAm62591MBfW7wgwm0zyqqVv+9Wt8t7lrMd6y4zOy2QxD1vabQr
qWm8ppZuHSDDjn05nRi0skFmU8v2Ol4rCB4YqKrHF7sFrybnLX5yF0VqkZgFs/Gr2cyT23CXisYg
Rt76FAXp4HNKLm6JTmhQ4NzMhe1/CmjyT8hey4zpFh5gMhfgOty3PxaQ4Y4CLzfkFK5zKRW9lcZv
Tqw0RVVCQZ+ibyD84Yg2gWIAoWv9FULeYgz6jsSg+W3jLgviJq4MC7Wm08MSxJUD1/qYnJcP+ewX
z/u6jMGESMCvPHObTurxkM7y7YpmAkPEaz9k09uOvLnTIIPYQ4tC3P97F0smSuQrU3ilBDbTq1Wl
4Obo0sFLwk41UrySsNRvE3LyuJ0K5j/89ACArCq/6RqwDPkda5YkyUHk5f4m0tMtLPCtq205xUfl
v7lDPSaujLQqRZVjTGQaPbFLAyfDezDFbxNb0vL7KQYYXsqWlrxdiiIGeYBUaVn50CKHIKZdklkq
2x+m05rtNrpdi7wfbrdUBx/C3ClAyoTCDuat3m03wX5m1zzzqGelsnbaXipxm2OxffZ+CKg4XFsd
BHrblMmhlZXeIPCrweHzPWMDoeoFyCu/NOAGtuVe/ntOnsI4MJrS39sBImAx5XN4obyC5K4ye1T0
teCh1pl/QhCagczg5IE84MR2iW0oR/7M/kTN8xOT44DsEaufBx72QdRwdeDLu3C+SZNcaOP3K0ep
i0mIVYCzGLWJtaHUMnN4hPS0ggL+5WH0nEa+CD8Zs1P1hBPr1jCV3e/wCOFo1xDkHa8D5SdK+gYA
M15MMfZ4s7GXgViHhbEeuSpfQ+Hw3YnefKYb/SnKb7AdxbLRZrgCbrn2xyXSPu997sR57GwMfCmQ
0f1cy3q6lAugPrcv6sb9yivZzKMPRxGO6I2++DulmsDVtQk5MdVas/gUSon1Oz3IzVFMTz/f0VGi
swcIi19otDwedugYgo1mySJPh4SUr53B/CQpZgJNXYefQuc7KBjeeTyw+QmS5s8GMvB1k985mJHH
axJFnk9eR8M9Ewp+jZ+7lIfaOCRRI+V1ML+KhZJOKMcAqA96KiDGhQIYIncQmKq8hQWZg/1PsEn0
vSuIMNsKsKoeOzz5rk9sPrFqV00EFIvKxGWLNS/7aUDmrLIiGXXU8PLUs0Z2vIeLnPjuy3ynEs2x
xoaBm3Nqh4iB01J2ooN6JATgKQlD3RgF35dfVZfSWj8HS3BbpVNSvFz4XB0kCS9V6Dpl5X560Cvn
5A2/mWQPlJaTburwU9wBpk7lsFD98rfC1sXP0xVcvdNXzkx/EOxfcNEa1D6eCvz+tgaaN2QB5lCt
5vWrOxUZvYUB0PCur+hoJ0QJBAjRV62AMMqXk3pSycRB8FTjkKzKkFn9JkH/rLxSk55drjVDtVXB
4lKp0pVuN2GB1t4g9rhaod49YM/weLp+D/jRJ8XW8uBH5pkH9bfc4bhJIMHvzpMNBuqBKCDgUSuR
zuHxY0YB/wOC5oPWHRJReJlRom8R9teDARpFT1hqmdcxtPsHXlxloXll8uZHHCZ5TM0RqmBKKxWD
quA+YLEX3OiaCj3JejkiyVhshgO/pZk9HXnDIsaM5jldDF41K+Kx+ne7672HnqioRecuXq12VT0m
QjhIz7Vuam66GXAZUh2u2D2iSjO4amDifwiLOkUDNLS9/eQWgEYu33AjMOrqfOXoExbVoMGwvKsA
tjq2CfMqnS0mxy9o3cmhLcNNajnDXwIkVnZvmlp5xhkum/4hRRWQEBmwjQOUaw5e+AB8hjJYATyT
YkoYqN52EkR/vBWD8+/Z/jihWHSMP4naTBZVungjdnKcI3ybwt4H733lZWdGy5nfOA+PBjUBCks+
3pkCoGFpjmfYetxq13bw6QBxXKsYFIm4+aEyti4wt9Gu3wYIpzY3KUgzw9U2RPeIlARboSUxFTMB
A7IJIX8JG8aviIVBMeH88xq8/A0uLZC4L7iAqcoMBVVNn81qb5mhuTkSrWYC7FaqsbpNXQGipK+2
eoEjttw16ZTSTUR7+euccNZ9Je/pRv/k5bol3dozQzsqC9zItdfh3d4GqJewfVdRIzTuD/J9qlO2
TogseUbFLSWrCA47UCRMm1LNxY5rKVh7aEDPo6Tw+F32CANMzrIwDWSVl9QehyILKP5lg1FsOQoR
9N1Huh17d5GeFmDMQqBlD5cveeVM/ZA1yXGuyMnsQ+xjnYsRpcgfrbxQcXRWG3PPOv+uS4gu+qya
2M0RE/Nrz7K+nvJxzRdo+x3BuJvHiZfPrcl0WmhBVFkHcVOrIycU29EIg/p0tlFSA2r6SK6bjkKP
JX/tl/FaLAPzuMKt/NTLpscc8dJdWq3UBxcRzuZrH3/puggziX45BSJ7Ix/pDMOZkzATi8TnfTRD
X51ZNh2cQ5D8pX3qWG3LJBFNJZQ4BdCqK6JVmfiXBfi7TICViz3xmUQq/RyaDH9JH6PbEX7taCyA
g/pKnyurhLP0G/4/iBTqzFKZUYn4dlnWnJG21szFYJKXlMCPuD1U4IpmyYBqcaNbAIjuVaRYzmrP
nZTkjcqstcLi9e2oVBTLfU2qQnVwkM3JoShafiQSvnQpdOSidCHJ2uVKz1CPRnFe7pwxfO23PXP7
RmQlRd2QVwwvbmSA9+2FOxyduNsrSimXXGZ3JZo5PN6goEDkIY0UWCL6Qyz6w1bm1fjpj4pKwMHl
RY0rjsTDOgY3ShnRPjV2NF9OtorZfkHr7i1tfhdCczyAi2vEeKSPXKc6EcfETAU7OG8PpvqunWaX
YZ7OG+Lwv3oamaNHVWfQG+Yz2c1x3bvc4FzuSmTUUQVFOFwqs3cUZpJ+goKICpNQqPBB1TjHXr9f
RCstOPtW6lWIf6kYqocAp4HMmj8j2sA78sx+WxA7P4GUPlPWeK5MiimSIFdmNDEzmFXasr0j8CMZ
Z9EjdWESo0KxRxXkYW+ssXfUwPH0eoOy6dqZ4V91bJEYpS9VFP+41cjRHrfK9UDF6DVQvnYP3j07
5AOidMvxeyoosW5V2bAg9bmV+pUfGBrpBa0OcrNEXMgnSomB64txyZvAleduF+gdttrQ58R751vo
3E9hjFhVhGq1eulq2+KKHzA4GUdB9WicmxMossybduOoQMxZG/PLFhTAfCjaKaX9Ruimtl8BL4KQ
brgGG7mdJX8HZS3t2OFb8FMmVjcYpTSu5thu7ajy5Nojs5yGBFicAqUv8F+8vXkcI3DsoxrpB4Uc
R676OCIFlWkvuhnw9WLc7bQIDJoYP/MYkg2ze6i7M/PvvSVtZJK983LuXlTYoctOfGQrUB3HP2Eo
zuSjwwtMLezAjYD+mlgJc8QiF5aHdrk5M2Zg6vTEmIxvK0B1XnZOu11f1r68Fc1nWIVnp+z740Pm
cMxogR5pggJKE+CTjJk1LboS5j4KVNiBkodnIVhOeAjiAyOgJdtjjj9o6HzhrC3MJe57QCk9Oqog
FfBvD+J5SjysB4qRC6mQUshlN+LbxBvq7Tvh524ANnjST2pMpDQUV+t4VbkKWU7AXwzP+2cnoH7N
LVEcqFOxu0o99gUjjl/FKR2t6jA9azbgn1mWpvYPxdpzxYDgq7l4NAkSTfmaxU1waQPz+r583kiU
NeDE7XFgAbrInudQymXLpYold66dZIfpRtehRsrDwAE7Pb28fXh8FEFOP5aiZ0/hH/5qRasMrQep
ZzEqU1l12pGvqtNfAa1mkRV2tpPFQRCHE2DMPfSTwQw0nlBzXXhxL8xDnu9C324iJKaQScXT1dK2
jpHhGHSXi80HANfRPLTPTSGnOTATjPza5vvLS5mjdVZOTZHqFO0I42ecSR189AsiJqtXmNacVaSO
TUUdAWVYZqwbqLQuycpKDIYWh+x8OOl7MlCkkgoR4d796jfZWhNx6nAq+RIOl6iFU7d40pxnHQSr
DW0Pb1QWnlwe+rhEU2RL9pPQpH2pPIM/E5V3vgh2WrHr9vnqrYShIsF8UzYhAYzPrz2K7K2pUGdz
nB4220YdscxE42p7z/fMoD04cYFvh+VkHR6ikeHOjG6gGQ38Dgx4kTAJ6MJRUz6PSMtLjtyx+nNo
jc7/zbbVKsI0MRerX4HY/MjjMQdz0CZ5OZTKJVV5s98dGsEaWrnNrKCNXjkUwCh8B63aZoI0L+53
CLylacp9vMcD5pAvGLa+FyWnfQcQNE7kwnfpviIfIJqi8K2pgMiXf/3FgLwsy3UHS+ZkNyPMEGVs
hrdqp3Jw1F2UKBzQ2Kx7vsM3daIjT0VbN9VSISAmweBZwADvJliXGDE2I+QTWmMZHPhh6q61Xqf5
iMzMHQvHUpU2RmKP97xVQ2zYBnXRCQaaO8C4MKOYtmmds2UOKNDtOfZLdbKNjSZTC1HhqUNEj7od
nwgm2xOrB+TGslw3bKwm8SsdkUHZ6lpf529PfOlabX2JtHLMunGqPumfO9Y9RQM+piIXaD610uDj
P0xql1FPp4MV34MibdEznDBgpAAtfbxyWuCAD5h//0OEIS9pEkKq9jHKMd7cRH+IMA3LIOF3iG4m
la+7ZJtPbwC1SPCZI5hglTfRorIuYoKYDgX88NXurfIeET+eOZwFPL9DLuqE5meJ4ZjVeM0S7r6e
ahdT1OBg6U2B+xhj6EkXPdmc7ftobW5MM6jnuIFhkTPYSsjdG1cIU7E/6xIkCRGQS74IeTsoW+ZC
JB9zijR1No2l10Mp38iuu4YsKN4T26ZWYvudAzUjL8P5Ue1DEv126kYqEc1thvxqWwTUMJ3rPida
GTTyUOuDzLdyJmQTEihv31+/KrL/H3/emCckMZ2DAnDM2j7nYHByZ1U0BbieY9wEA12HSftVGR+d
3zmA9lL2fIfUTUKAuqaaM3xJoGiL+N8VUn76xD8B4QlTpAx/2lF7/hVePNv2BeVgVurke8pkzHlM
MdHqxkVl4sIIKvXk43hSURcDcFML6GnC9cuWa6pakmD3x7E/kZh2IBe6QLD5CfBFAh++A1ovyqdm
B/kciU75w3+tj9T+jmeY08ijPOUeUM3qrBRtw0ksgcRWUd4tzv1p2ooMPFYWc8n7IconLplZzxZE
EahK/M3MwSOETjnQA9bBT5uq0NblkWL8a3fR5E/jqy3XH4mtmQm7fXM/aE4TGuprxcsDMa+xkd3T
W0c8rHl2pTMhHJ3fgfIJKhZdrc14u7dv6uz8E0VtDx4HZEeYo9wXjP75uRLc9rIFvglCxWqhAKSy
1INuR1ag9NWTbkpByvmwHBAcBOZQbjlw2EmDMNAPQSTGnr+KqftiqocJqacLC2mMh2+dT9zv2YME
m1ybdkVtP+oDPQpxzjvfGlRvEcOWguEjiTOO79HG7o7LcnXaRakNU4IoeYyTO0Gg8B/FuLMHOdHE
A3OofqkZkfxnGSdTgZxP9cdZ9jFmi5J4Mp+DJtXEyMXsckkcYltNEL5H3TWY+TkyzY6xZLESXrls
7DLiX1rLWWQE4w0+sFFOty3BeA55Uoou6l3+dwZzGNKCFaGnHos7cnJiMTSLld87BbBKzhxu9ikG
DgintKLtFT9ZFvHgfeGht1J9MoYztAR60eOkG9jdN3hgIShD7lVK4VFdIBqg+akg5ogqr3hDV+Rz
LMv2PONz99F0ftgzv8+fMO5EkpZgaFdgMKPr71BCJaczZDM6AbamjQdDoA9bN2bgjS5JGMFjHNdy
HapLJEwoljWSKRvobarpG52Z9T61ZCuu7wxSadYDujDcwa57zsQnmBLdpadOO2gJhLNZewAw46jw
66P8EIH06hCMuljEaE4xYXl7DIewX/hsJwaVAg//wHh9TsDr7Ip25WqtICiT3HfYSTT8f5W6VO79
9+W2qSdqookcjniWPWnbH2mC+bfG5KZAQ13Xv80jAmI93a28M1yHiWAFwskF8+rrC+Fnym8/wZCV
CIntbLmc1hvubaDsDZOBkaSaNf0DjDyt0ewy+vUJ4i3726EWZAFeoBI7IIlLTzGX9Wkz2eg+p8sG
r0U+An+VPaDRZI5ExSFGIphmOI9RfyfoGVKk5p1r9JQkGjrZRpNmOUQDeWs/Y/dCyRzO5AZwrJkj
8C7ADV9MH7EvD2hpylAw8YfcebtiERU2lZae9S2m1OeUMIIhFKH7JizuSIYZUkrZcWaCvay9RRgY
Pf5fvqgRGAxQF4wov0OKd4EIEhNeVSpcBHkdn8FAA2tu6vN9iW9q5FO86T1ZFsZQ3CakPWyTmZdl
JVdohqozjJoFzM3evxLemfMUFaWkSHSmEkcHUL0YSJn3eFOm0re/qKXl2z6G2oxO1EkxZ35IXezW
8ZbHzjoSwGbp2SwvdxvabaO6YStytxqQmF/l/9DOGdqO9+cBf853dRywCpjz9j4fNFDVT9xrU/lz
sei8mnC59DWDVu+zBFYyeJWcEgRk8bWgF07QqiC74K5RCDc1qrtN0rrY82Cr0YSxXNISfvdXp6Tr
64xKqyMPZ+Ms9Y8s7ZOdkiaZiRnLERHBFi9QMjq8P+hLgRnIsGNQk4gJxAk28aLlFHH0QzE6yo5n
oYy5WlYxm4Y6AEDazggKX31iHXWzWC87iV4CsZsCs2u6OcAehqgcUstnAerHH7SLVrV0GS4j3qP4
H8Egj1JV2h3adhHV0ZR5y5jjAlf8FVFJIOW6R+X+3TRbgU5WUPxOXr8i/bygCMPhUWXXFWwHoKHC
wqgT1ws6q53ZeWvAR92+YY19QPdOAvz54pfPzuBLnV6h4tkuaGd7Zbkpa1WI9Lb0coqhCUdxoI6C
xx8wiP+RBV/moH+hhaVv64hcgXinEnmbRKZQKMg0xbZBNzJkNi3/p+N4S9gpgq8aPVBxfbPTUvWS
juc7F6CNAKi57G+zRtkv1vlor86KqMA2cpzZKcdjOaOrFWfvACISpKXxNlXgE3sOAVpAWPnEcv4+
UQjgusHOFVav7mwsdLLSSTtH3nl5lUq71Izx8nzDbgnu7P0csyaIvptVVOr1GZsgUrL793bFqOkH
DVwamMqXT62cuAsbWO6lFhkPvuA79q6faLN/zO9WTpyyQUpWNQr0jcFZJiy2zc7fWNt40dTar3Sm
R2SexX4XvYOS3qkGyq1072ozGVMRWOYf1j8BeY+aGg93Xxj1IkPeIyTGZ0poiCBYaehBqgBjQ9sd
N9n3Wloj3sd2He/EiWXbwOyfDTni3ef5hyKZd4UYybVrMl6NcnaHRF0P4qABU4TjOqdQrYwszjyQ
wEjUjjVdcEdp8a4zr7AFR3l6wixSWAklG5+fdLB84rHTuqp2RVdh6U/HtpANaXzI8Vri8ua4eTlu
u1f5f4TVyApTUZpHzdtUeh3I4HSvb7LMK8es1RUvVzudA29L5Sa/QQN6gKYFEp8xyKJCgI17B6hs
GVRLUqBcFElcRBj9C6w+SoB/J8mGwr8iIJ9OSSjem5Wnq5QZeFW88E9EzXZDFQCrrKShIB8SvsoT
BtjSxMZl5v8Qhvg8z6/iJI1BshR/viu7RpVV1nC82x4iiSn40uc7wOHBAUNik/BnAlCXOGpZPW4B
FNIMNIXTN3c32tlwss3SVSC1ovO5dt7cuAT/5lPRkjPazsV/bZS997obRiYJljQAYbyk2HwMTGbV
OxQRhWHVAFKNibrZ1zp166QHKeJ81lv/v2TpqDozV7AAL9RYh1rpsdmPO6Zr/qkaP/+8BsLfZFlt
kjfoo17NHokcF0L5aXYAVrIEYLgcasSjPMT8frAWk4g9BZ3LrVUB/niS7b/XDltA6uFBPy/NnSnQ
d+FHQolRGAE0yrQ7k4TBCna7gCZpsPLhyMxGJ+uGdLxN63kM2TKM4ymzYm8DkvFHb+StAId+UOrP
ffk2nCpTjuAhAJyE6HPykc0zpV+NsLbj1xIQnOX9fL2lX1oXGGlT4kaCSCYvSuTN4wA4cU6uzeYN
iziqQVIc7ZdYxmXwVJ1i1LpbZjQD6HMZ7Xak4WziXiRM5DXyfxosFbc5HPzsHfBZdieyD/Vk+756
xeptgB/1WH1OmC4tfGY2efuH5FeI++hsopTpWdtn5n6oAM702HeYQyIbk1yEPAH867CaqCS/zt8B
BcI3kBpYxj8V9TdMX3Odmlwe1xz5nGRp05q/Ht/uJr9XuzX7ZQMBL+ABKb5K0i7ywkHJ1iIHZ0yD
KHy0+e1fqCnd/rTHW+h0tNCJB8B9ZTdnc9tmNN7NRMg1k+2lGL65FX5UtPhinufh8K5t9PmYv1PS
VGQwtWslA1u/JdqYi5xCYYBZkeu3vqXup+a5Ipz9Q4g/+6/JYxLRa1RlGrblaHDRZ0qKdxiGGy3F
pvqYvNU7W3Yiprf6B++0RKlcr3oYfqKUO1QIYt4a55hDrc7axj13NrWG9mLHkeKClfzVfD84pTyp
Mc48MIxKcdWdWSXoDvEd1CHKUdar7JwKbawaDtypuG4nx0rBOZc+NlzcN8rXc8MFBYV7CsbrQ+02
JnGlsvuaOxUdHi3zzxENToRA7olF0uB8P60r4Gs1IjOYT9Dcbv0bfokEesE6g7j+5OpsddpyWrEm
nD92wbwS50BkulZMa/U/HD0UVuQt4PcxQkk4lSdOfyfYj2cXVeHpaYipyAQEzslqT7j8Kc46bPLP
8tuNz8eqr23ZVFFMnDYYYWy6XgDIqei6giFPOQ95l2F5TRGsBZE6Q7D1WKD7/h0tJ6aFi7McSQ3Q
IJMx364XozUmxIBetpfHnhErrrU7D31HvoiVsu/iH+Fec0/eRolAgvj7sPjoJAp6HIwS+Jil3PH4
SRXrViFbsTznWFdz9ieZz0XN4ofCTBGJa7sAr11u0Ugb5nIi3gmu6pta9am/X4FZ+Dd7dJrjgTBr
P6lOdpLQmZAC38NF/h4Ud7SpFl82PiZ3HaZFtOKOZOZ+mx44Be21K5YWmBsZUYsCov5wWwGM3cUy
CpVSYKT8ZkTeQ+NkoDd6ru1j6tKVm6ych4lv23FvCd8n+Ip10Y63wKsdeyFVlXDqcFECPvQaPRQX
INdRMO6P4yRLcEu/7bl3Twa+r6QXKq/Qza3WP1JigHqvrzSxpzMR3Bb2JDtObuY8ymeeaJivM1v9
0n/TVupFiMnwrJlQbB78vQBARannYeHjYT8KaaxheL8zjkFq0nBkIb6DF25oFHEPQyVB4hgQtvPw
0p+BwBxcVq6hmaEQwS3B8joKkBJiCi4x8Kwf6zc0usFXD78WKbGsXT37mLS8eHiwWzBWxIRxXWf/
NBQ4UGuMN0CgIqqN+mmZJioudOvHk4/4eZFkddW/kpvJUMpOvRC+QB7FujLwaXJ/umy33FZx4xk9
xGhpgjiTw4HSC4Al3Vjtkd3sUMIJxLdqT6E1qCB+g6YwB6ONwVJU9iEVHf1aN2ft3nVzvjMmL+8O
0reJ6Tdt38wqdavKmraxi2ltNI/sTZ7eqOedIkgQ+05jgcIfRnzNwkD+O6rFc/4YOuCfRTJ4RmIv
ht2Esa/VJOn5V0A99g/FiO79UhVkybUoMxCTqlPuVivsqZ20x0/2UoeTg6lgtvGwRB1XxYZEP6re
cptmkr1vVyyjbZyL1islmKDRUmi+HBVi9iwM4xqHHs1fPv+/n6RxSInKY0GiFoRLNkTuVHwBhBIK
zEqiQIkm36RbPRnjOZAHKr34BU8vMrUNYFOJJ42XDLFOuDsd3jn7jt2Q/C8luP8oXIIrUU0OkrNl
UPaXkwrQvoHBs+LMlbgPNMSEu4am5AXJoSm4EQuUTOSjPeQEYq4WkHryRaQ7RTHuzL2ls0MnFhru
fPOqTzuH2VYqes4gqzqJ4pZDF4OiUHN/Hhqy1Z+CSBLs5uaDiNld7Cqah+yXemDmjah/njeQhS5N
XDdQ25kKcOsE+KTHMmQ71uR6CxeEUPlDoyV1gIpf0qc7KKuFKS+DQ2jpBBJo5uRelLtleGD70nfR
fMjp5pGVXWdEu6msKAY0LeeaxPLTXsEOXzEmfA9pVxBmQ1gZVfsbqDPKu3lrYm6HduQLCYrMxy0u
axMTGH3pEvkUDIc3egdI7DpW+FdPRpTwEmnFC2GL5jERfGre2Ois2tIB+Qekh/YZ+ONBoAmwDiYR
8Y1sRF6s2lGLaSGXdg8uq5oIgpJszmRCbkJF7w4MUYk/qGGpbKWwqbCsIincVS+LJ2PTsRWB3MaG
UmkYmeWBcApapCtBp+XwSSzfyus9FyOBhuOu93HHKFCzTgpH+jY/zSr/LAsbFOECdoK3ltfXURsP
E/bBo2xFGa9mPuuyIoCjp4JfGHeyCNqYrNnwO5raLuy4/2E2uZyaKL64jZluN++C/UgsOqd1wDHZ
AGpIDqF6VUfjfC63Hmr0IhRWhf5jjI5FBD3or9snTUKHw7iBBW4J9hR7DbQGRT7RcET41cEqSkX+
X7wYXlftU6cW0moQOUrtZAYmGygoZniRpFJyP35sE2WNWpBx22MzchHJfuQGB3lShvPYoeDcVNhr
rTEK7m419brFsP7WInH5ZnUQhE6hQzt246sVQmldynMkjVlzfXrS8FtXs8zG3u4Qi60pJ/D0rRKZ
4J+ywbCEHbH3nPmeZSlp9439ZQJ6qBgdKasSD6BKuQgOLWZxxjkgNCQQoCo6bX3TFd8yUOflJ/W1
sqgfP9gDh5WeEJj6O0r7Scj4/wQ2VwlzMACKXfYqzjpXER9THues0dEujCl+BcmpmvJJdLzzWoyA
aqCyEus7Qj1ucAai96JCm6up5p+MQwqn0iMJigF2B7BR/9jlh6LCs3glt28FOz47aBLMZNbwig/P
U/KrQyvur6B0HtdPROW+19lwdqTHsfB053lZUYwS8lkVmgy0ejYwUJQlNqErVr+5TWFCRI9B6ndA
PWIrlzluBiQZ5wrQu6ga033tqMBuN3dc6rzaSKZ/QYqCt8OcQMWl3M7i/xVuFFz/Co44OgGNSske
kSMUFWo2fUjrTYnFVOBEoxDymbceL1D13398/48aT1N1hsasz/Ie0ScAfzRGFN1LceivTuL/q8I2
3+HNYLJIKp6+A2c1i8bhw8skg6fOK/dFdkgOI6E8xEhDrYzEnjoX9343GWUgrwxHMoJwjIid+bb1
doT7JlkW2JfRCkWXT8rgl/XlgdWn7EnsJXiHcheGnBFcuPdoHmJWmDc2KY20XxetwTKJM44CpXEb
+QHWf++221crbN6q/vW1XEeo+B5BjUNttf6wo5IecOYmMDbVW/z/xagvhNZUY0U6fZgicnlqxZla
msYZD5sKm8FKRVQWKYRth0xazLYzq1Pg77m0eob5dqViJiTcenaa6edVqaOBacW2keW6xTpuhHda
BbCp8uD23e/sJA75GUiqNF4FVfhq3KsCkGZslVtxeroHGeHOeDE+iXHh9C77ycOunfJpNp7eylc8
eFSgVEZ1DtTqzyz0KrxXSTuLpThzLkwP+ntGQpxwH6ouamMLCqPU/QCO91CIiTqETEXgz4oH9kAv
W5fYKMALztGjX6udg6fvpzpsWsTzsd7pujcVmkws9m2ZPqIHEaTnIZlaHaGh1JdLbuVkIeV/Q2hi
D3rxnzP03WtufW29pXAyMGQkcCLDbYgJepORIcTKkZ3PaUM0/bEtd6b6/91G80y/pHtluRiic0HQ
7ouWoOjPguT4tmgSmXl2sRPPTcChSCe47aPnQze1pe064A8wIwDoyLZMjAK+jb5n7lM9IhDXg04c
iG1lXKJLEi593BnCrobmhQ26Y7G5lKMh831U59NyMRtHDQnxK9N1QcZEIWN98FL5KkhLDgF+zEl9
vSIaolrpKCQvCoizhswe8RKLUWMvraFUg0ftFurFFErrzdYdVd0K0d5anDV9ppU1e5aoPew2pU7L
cRkYv+Fv+0nPaRJ1GpnqymFeOTLlJkEHjHxt5Ntrv6qZ4Z7rbbY4vqj9alq6kHYg1AaoBiYShyrw
MItuWXowDhmOXx75Nhp4I2YCZKZY/wDam2qCTJmDHW5XqI6zBORUv7oIySHtuTBTPD9p11C3O1bY
GNKG7+sEPC0KjuGnPxNrqgFHU5ArwM+0wNkzcINmbhrIXl3tC+fl5IUgVGMABNC0PPStdOFPSVmG
zUWIolDtkBE3tfXS2IIW8NtpN1VhapyfPEyBs84LJ2tr6o2S5TqMETuPU9u9yqhue4zbQTQnomZZ
7eX0QuJGXGVL8ycI1FWdOSFJuxLShCOCbbNQSpJtbUZFvWtqZQgeBO258S8nVk89aeZ31Nw4RCp6
pGc/00goCp6EvXbOq+DaDEyznl3pn3I92zS0dtGIWuXifL0xmVtVWqjNnAzcm11Aoh6seEFmVKlR
uHHgm3DbOM6on9WANCIS30um6jF2qDsQKZfu1NBrLlsochlVSgdnDrMWM7Hl5rqyG3l+hSIPz5Kt
J7lEQ4HfjgiUemwqEnYDAcU255DAAFLKvqvUTpTVhZeOX8uBypZ1HfmmXPtUgwdtb4enCq4O8r0A
beqjnTfbLheeU0S60RgwUdZSim5LpPD5tU64D+xwe2faX67cIEAum6087D/RryHv49fosMEvoUMY
P+2ZTp7DFxc21mUimfmKwAAs6Nt5A+AUHlZKjR0af3KOIe2YJn313Duo5ph5oeHYWoeSVoEMbUw6
5QuF4VFlx0iiudnpLksmmLDGovjgcS7K6+dTvNYlpSWbQgb6IkVPxFoha4nK27pJo4gXWa6HA1aw
YMcOhmOtsrFRy6qBaSGLx7YFDIjd2wn2Q22FJKAUbuQaVerrCpXTeR9bC1h382+HUkJxwm+CYxH8
iF0urVfltVkjHvIo/GocHdtvGkHrZJ8MBj2gNkkX3X5IaheFS0wQo1QuBi6Mx1P1PoaJRppAf6UM
Huim3Emfz8q+qtv7MlEA/xakajbJmDrh0SnnypsiNFX5GbQ8+BytuIu49s7GxMEx8rpnCOvg5fsV
6bPAsYoeXKI4tvgz+T3N8gjU0Z050Kh99gRk8eYhA5GGf5YXg44QUnU6yhgJ+z98mlXedkHk/3Rh
a71UDLW9Q74vCQo/cN2VZ+UmsrDxiiMkF1zIhUkc5VY3m78rac6w/bWzLSUBQkmzH9EeBzH+D0Gi
MTj/tDeIIRrShK1WFxliFVdEZzlQdgnHbupjSCfQOiF4cPl3QpgRp8EKnRoq1iWWa4OPqWiV5xC1
wUFoWOs9XWZbAwF2AnKPcbT0WtlWoPQeeiIEw6auOMghufcZYLL22ifDVJ69IujFhvZ20rrO/AEg
zjcYaUDumIEHNz8fEZF6PVl6ZesdS+X7iH4xto5qyQ+G1fAcWBh/tCe2bX9IOLeDRJErl/qDg+jv
Dq3bly6H6tYJ5rDkZYvQHFjCr2sM+/JrKjiXEy7ikrkeT3uux96/na53jRLt6+8OgaWwO0qpBMLb
o8Kuum2Vd2GAmaFM55HnFnrb5qlo/ml7MVES9ZJGQJIspSHpkmPv5ZzwfgE2zxrvBu5lJWi1yRu4
yftmILl/QXWZlwvJgMRLDkNDccu9Hl9WMIZs4U8Jre56KxX7wMDAyBWF5Y6M7ewWhsWXwopDOXm7
y8fj3+xqIaDQuRFRKxYIvLq2FGM1F9kamMViNKqfcqMRXDn01VipWTmdvKUq2eulnOIftMWtBBfe
2FrGGb+noBjI/w0shXBzWc7b5Z5LyF0TFRWm1xXghV65w4bFC6PJiHBTCKUJ3WhV3Hrcwlgn2kjh
5vFRLwEDxxhOM3L2KNJn/fUq30L8sDw+qXR82jlXpons3T5bd/qm5gOi6R78DB7uDdOq9FOmFYz6
qZ76hDFpDJV7gW2ms0iPfmajgMwSOFd5sTdCOxOwTabGkTau2jp5ftNszhzsTrqnYD6BppM+CluB
o/zmMYLiKBPcVXCx6wWfRwERJrokuP+A2v9Va3CcIR6ha3RZg0Wd2TzeMDXuRpDmn2/HvtJhHdXP
7tbckOi1gKysx1fIrhDKzT8E1NWMSjM4K3yOdB3Ug9SWqd47hkH4Y2kZ0DokgukZqc9Ks2YFQ+2h
bbyQt0NHqAcdQ5tUgG9kgABXbL01eizC24Kl5Nu41FZCvJfUMBkQHpcGmhYVxi5RfofhKzJEmaaw
ftt0vNUUCSJ+iJquoR//gZzCyu7Atim7YekJ70UFgVTWWnRlh8j9rK/8UCZli06PEkZtuWR5aod3
Rs8GOj7V2H39gmWAMLOU2gTeFyn/T7bHn3IuqvvwRIMVPs0LEx1d+Nn+LjbFAe5Ael48v9Q+rfLB
hM4sBL/oC4z7gXFUs+0Od/q2SQkO69lrP2dIuFYs17koI4f6GSX2YOdALIlM3qRpAnRH701RTZuO
vVrZbtXqbBk/+lr1kuuRctXX5Nuqu6+a4FvYL0ixCVGMo3MZ0alw+/GGuDZFZdxF8DYpaPbVKtLq
CFSBFle0eKjHZknIL5QtrMaPpcZkisDDMxDYfDMsOEk0C1YN/bmnkH/WxCgXunaOICxkSZT+mmuR
mqm9bFuw1Pa4sM1lrDdey3uSv3s78eHF3vzIGUvK/c7j2SUk+Woyh9izZa4BGZs2mKywblZKY1y6
7WeZfH3h0fIIlY93W2foTUEYekYLyB1pIdnZooe3Gf/Ef+YiTNgppzTzU0dotYz8y4x9gcbcg4vC
RKL6wpqpQPjN+vg7nOAB4w1m9E/MMua8l9TVjTqASXd5R8R5oUFTsofoDNgHxOyM2kIT6BiwDD/3
6NaZdjVxai06ofqjV0hcXuqGeL83eYxm0NSqqboBpHB82VetFFwIyjCJhsRtxenwKtQ54/L14oth
IxL3tu0iNvcd55FfpjR2oE8i5AB4Z0ox0T/pD7GvTBkkGMUIngVBXH+B+L5Sfh4jz6b9fN+S1J2V
I/Km31vepRgITc1Ms0BDXhc3oD35QicROh9HPw3oKr/8BtrGO+iLoabfM6RaJRAU989hGQafcJfn
tjnB6EBCJ3fuWDAjCjG65QJLop58W8bpPc5N8AYptJEMXW6BLgA9WzmL0YrblMa8CQlqszE3TEJX
ViAWNNtBfv7EDDeZuggqSocrg8bzlxxt0bXl7qIxCYqEccuSBAjflDBVZf9WVTFMSM+P6fcurKB4
1FplXHuCJtO6ivvUcsZYu4uP4zFzUXiusItCjLn+ZPCQqwyOmXuFZrI4WcThZtzSXkMYdgQcmGIn
6fxAKD4HkQYcsZ8najjo5HZ4g7OJO4PK2xdNkvG7XIqeHwWbKscnGSwm7awzHsNbA0maiA9J44v7
NfqQrUbkpb08oZE56rY41Tmoon3QOw+MPLK5sIoLZwJfw823Eij+PM6auOQK5QumCBHgNIOg6WYv
srOJjIu4YNPxK+8gMMqjY9/btFBWd/FZM9Peg1T3Tsf6+H7GbCmUQw/sYahvyuBXUeO5Bh+RrZMc
xp+v4lCdEqYZaF6oO6JSNZBRGqL+V0yQb2TlYVZ0+rNCpPLPGnPtT1GuwygFA2fpdTzmbuymjh4n
ta5XgxGGIJZgsF2jc++Ez4xUKJA6hnLph+ZL6VWNDHUbpuG8cvWBnYe7CxwaMm+gTi2rNaWP2Ocr
7G7Hkly4nwmVSOzgag0SXS6rJP4EL7agvO7Zrpj6NjYzkI+UyeGJn3sed6MOFCxEviEtXG1ZJ2Ya
DbMfIt3xnQ1aYeuGfWjbOCpQhAmTkfwYPv0x7SkJ/6J3qH41Ekjt8MWSh2oAfkdOTxkGYz7irsC2
46CLOE0QNZvQNTmL8offPjR+rEab1VH6dnwT5muE6gUEIyovMCvb40SrXqcazS78YR0S38/XlTWj
QgafH/zE0RHC5vSP+PQ9R5uDnOdnAz4tzfdmn1G5iWeKBrkvSTyB+t+y/YCUy/oEM+1QCUlVC80M
lI1fZ7VxRdrxlNrTtdzS7apkmgaM93IOtuMNLV+spY33BoJ3iGv9QrsIaGCcikVNUd7CfOEB16UT
h3qFeoXko57WBlADk+LqNqnc/+zj4WMiDpSA2sTp4I1lweLqVasuVsL1RDwb5yI/i6XVcdJwRqcR
xpViT2/T0RZ1isoUDutscbgS+gGNjjrq4pX1dAi8UAo1uFQkLl44jwdk4oJ+6AJeiQxsKyRqk4P5
jWfry5PsVnUQ8C0UVP+tu3lPfnOtVpWzI1MCTlEWEygAGoiL3Bf2XFQHhym2TrFpxMbtnKtO/Cef
OTGlhtTdT9moMiBj48ysZpfyIU2QzKum2I4sTBHwsnK3bilZ4wuqKY7hu2scanXTdIrkJuQqgAgT
c+NYrK6O945tAZPeYcWccVtDbTtZMQ55FvM6bugz34r3zBNr/gi7qtu6zS2fi53M87pvOK1IPM3n
PmR3FYirg2s9NxXsRSnKhPGpRVYfzMXkJbZ+MpE43BWH8kVLP5jE/TaecHxnvlcqp61lL7XF2IpU
5MDltXkAfAJdD42fzYTw7dJaRJnVLWRdMrGN8bzfa0qt0zoNi6ZAOGD9jDe3KJzi6U6MoFjc/pwP
lyk3vFOzDO0mve+wjCu61pi9ZRdzfFl9F+fCYUIURJEgIDJP21T4vvcfuahJ1XpIznJjXkuoJ35R
HMKmj0Yxv9lqUM4hYI69cFQxfvUsRjlur0gZrsggv6jAcv9omNkI/oEgGow6hn63/IB9DB+o2x7O
shvgzidBi4rtE5ZBpdqskjkMMkgm4eOOZhwUA4Z2WIKCCx6wRKpFS990hF9hbEoHpWuQmvbe7Fjh
OmTrwWINjlXrQvhdOuYcePQa/bR5X+FPTsWZssqRkqUKBkOdqyma9RJl+FbMKVOVkeaHWP7X/BO7
irm52zJMuyYW6Y+x3g8rN8SrHHA3d3j4GAoboi4Mvv2Xagb/FFOpqw7ggY4i5/veWEOl14SpAcZc
CzJTqjIili8J0l7xTH4lGAp/h0VSEey7n2GncyHLTqad+Q7+EyBDfWFYC34yJiN9/McMkMUD5NiC
IP6ECpeablUS2+mOxkhrwED0Dyr/So0pILBpzV9WQPPiy/nD9qJW3VYD57YomAohWBZIUH2TFDam
c+k1Euyag2D0fvFnmECD5nH/KAI//igwUBI0+Ry0GyUwGidOJUdJutxQ5l4RVtZKYtw7mUXrWvu2
bOT7yzvjkqhLx/u4tlTMFMzqMQO0pN1AIMw7zfDTkxsRrWJIiPsGXdmq87E9Z7/nBSFiO2L9qaR+
1nwBfLc1E0qj4DtybG5g/bd2ykngaRfJKl/5Mc0d5snZDEw9TNZ+T48XNg9RSNpk6x2RbNTQLm0P
os8y3PzKO20qSyJbSNKX2SGdmiW+YavHEiAgiQNHmHKMVw9hLxS9evjyLUL+rGGZa52k37ze7E5/
6/+JGLY9zqrPRlk7GwEEKRhm3r3xcJIXFrSQE0MORL9IwHQfLHwyKOoKQvxcQKV7Joh6Hx86J2iV
YiBLl7PbFGSYN2HfeQ9zJvU5l+Hh9NiZaqU3IKC8Z2Tkx8l0SEwAu4lE32NMeDE2+8AS6H7FeGM+
XiV4U3hh+0iC4klRJSZ6joxSLt0cEAQ28AHmdTkr6O1FuJxWcqjq2P78Np8zL5rIjLQhndRPm+AE
Z+cQhOlnQaA9yRH28R2YoxbYTg4uG0fVBvn8tb+gK+Zmk8cJiQggBdTYzR0fYW5+lRzwJ7zZrfeO
tGGexVGAT6+fQFGshwz1ZnvYCUqUp+mYwJvZtcX1dTXHHngKMFh9pk/KI76TcQ4uSvliRCjTSZm2
G0ihEEKhd1m8xK/BH7GG6Ag+E3yx3qSAgP2cYVuuGf52t5dso8LxabSI7DOuzrqnN4qYjgNHF52P
6S+sM++QHY0N1+z+mSjIvUoR2j4alRGwM6pvS7NF1Y5OF0ZxjskGjilrg9sCbKBkh8zsvUyS4DS4
ez/9ulyifbVyaekSzgnyogJmb4Ft+SeolDPf6Re49a8SII911fbWuToJvn/re4F2jH4fuB1wOLlh
c98yOOFFClHJF4XecBJKj2ZZGsRugM/aZz6CK+s6JYES+8qfTxFB/JpTNesasQfuTHYNynazZyz6
U/dnDMDEklDxFbve+PJWeT6LcHFeFhWGt4jisWEbe3m00t25I1Msq9WJxdJYhBm/UP+gAU+T++vD
5S+78GRv2pjKFbmqq36gnj3QmwsbfPuceh/hYO24xxDroHdvaNK/zCBR3PR8ADaqSDkAmZHMKPpH
uhVmzZbcdx5nkSZU3qInKHNqx4NVlovuHQY1HgxV+/koYQk8yFH+F4EEGrUOBV0gJJWNhyF9oMVX
Vm9ANa6S4eeI7XuztXEr2ilsuGximw64TirZApjxD965W6wixJFz9XSqwMF1SEWBb+CviJUEPchh
ZfAm+wSvW0aNy0ah5SKoaZT9VlcKWCa3k2tnZgyCQV1SIx44IYqh0kg8VAROp8qdg6dnGV9uu3ab
R0gof9VawsVKyAXFR1Rrm5Tk8LqLMCiI0BvVwHzfkkY6EF52oDefOp5WUC7ksjgVvTntDprMvYsu
EjjxfqpkESnswnQoD0vZjnfqgm7+j8c4kAIVvRQ1pU5Xfejdmu4bpzTI3DmOxTaS+bM5ndy/FCKj
0Zb08JcRO7yswZadNLbfr4bTXFbbLxhiCQj5aVoBsWbO4+0rAIL/nn0csCuA8cDokXt8YtNfWFL8
NUSVbm/lx8SxWKbIZLskQb+WbJOL7HoB5aQvSYR4DyiPg2jqkzU+7K4JRdYZvoxWgQaczvXkmzRX
s2H1DV1rOg0LuboyIrBzUXfgXNwkHqDUDibjlat4RIdjo59ZILTmCbEQKx7DGmzJwEs0AFP6ZaNv
QF4VGaECExsL0279G/jiyZ4qHvvYGSgYn6dtTU78cDsZiJtMxRlz7X752kwqD0f/kAxSIuFXxQr1
F4q/PJ3WG4FRU6AbEKoolXxypMoKCBr6jyUfS9xPWBZjRKIURLhtE/mtwW/prg1gmys3uay2OIfp
F0VigOywS9JDIJ6u4ZPK0qq83J36Fop1kTKB4bBYkTwkQcn0qYtqoHB5iie11aYK+JzF3xrVA8pD
E1MXNkBjfobvT/1kpy4daiyvHgVvO0cKN3YHDm3QyhSvjsA7Oc3dpkrTmfqEm5e+vvWD1WdtwUAH
w7PMJF+aGEXYGqowaEB08OkZ/AcQwG8jeO69ByoHVawPUARuS3B9oQtTP8geQwaK8Q4wZNmFtg/A
L4gVi8Hqh1JmpNLS5EotyZZgvB7maD+jHQI3WKIs9AHE57LPtjwjeU7yvs7ePGHbdNhYavlUhWSX
IBQS+622JoLUrHXonxlNurS32C8jezANAwRY96TMx40Js3MpzrwO4Wt65dvj2j6MI41YdLRfHer0
0Kg2RharUiRis+LhEsg0TlmYymMGSLaSlBztpQk470yHqG6WhoWDcuuvH/U+oaNr3XPo6QPQhhWN
c7gK6/842vk2ytXDc29lQDUdjKEGPY3ljASJxbHemiDu9Wo0FR5lWgDABoBkfHXid2fjap8Bw8H7
QtqFhZrFpQiUzEXHwAYnzQODNJo9H6mDdv/UBVeRJHjvqL6GZEDHPjs501q1u/UmZA6j1f3PWmSv
NXJDN3UylSmTEgxT1L1TKYzOw9MPsjoVGax9dkzik6xCelSryiCg80VRj4DGfk/4Qxny8+Ve0bXU
OF3uPgnBST/CJ5qWi+2HQ414vwM0v4GXZVdyA8TIYPtYfVxbkztlDgy8AS9cm81iVo6AurSsEIcU
t3LuT//rV1Y5ItYmNhPR7we4CweYnDXbTExGAW1+sfBqxELYW9cjHrAuQ/XnU+pd5V8iUBWbtWj0
NuE+KDlH2v7x4xMiGtGmWFXUZPVOt9/Rf1s8dKwd04MzynYe+nJ3hm6nXAwD+dNGrB/RyFnTKTO/
Ecl3JI0d8vnSna4hfLj3KIK2Ob+79yGxIWqHR/7moSMR57QUiZxDU5UGXetnji1rg5Tp7MgV+2/A
7CLuBhJ/E78gjjcoCWplQdK0ulZqA1AQQglw8hMAdueeyHfthu/cJVd22YuNoVfq8PGb+S5A1LON
cpiFhdDyTKKcb51DWcUgu/+6/lGZpourmmHlfQmbPCO0r24REw46MMWE5F8B5StfMsbl7Dn2SBqS
kQ0kDEtKalg/qB1UH0GSCX22Fs83Vd1glC13+b3doufVGnSSwnFyOWRE79Eb+3qFM77W2WrBpkZZ
Mch7UnFVRP+mUv2dZiwok8V4xAWQgNzgfPrFNJoteNBVjbz1pcKHD+X2HNBkZxnBZFU23Ik9Ib7g
KlRTDHXimG6HrYTAyOdhVgRZsn/TCqaLRuS7WnXLNVvUbyGUDEkgogLCwqIwvc8gJ9uaCAkPseoI
+OcDojo7+AKO1+tb7vyKV1xm0kCTlYaYV3UNdwhQNX0tUvwG+rQSMoozY9Dz5f+RZpXOnhPvqyM3
MiUnqR/l2U/jbsUCZl2WfF0GLUEP4qtFdO8nk6Shm+dC8MEJeE2GNEZ+MoyKZtFq/Zd2FaeDubOL
0hxim5ZJts/U+OT7NIZYDik8nnUt7BhS4aV8Cup0zFLyplyrLbgpMHpb+JFT+52slThYZGw8EN6a
remHp+e/UvpaoOvCuAQBHS731mIA1kd4qF0LvEToGaEQ+CZgpkAgAbrZNhwVb2PandG80K8kgMnE
c8rkXjDY/GiqCk98pNPL3liz5aQCLiiIWnFMXcQBekjbAOmyPYJ0JUZmL+zUOHoG79xOFF8pzseb
TNh9wp531dsSje/ClERBcDfSOmFJeUEezkfBV47iYg2AqCCWyAwcssj5Qf5NJNpfGBfD1uafeXQ5
PCjOsVbyCdhMZxx+tYraFHAMSnOzNGqngIO2RZdOczP9hKtzt0miAL5XJCRKEnwUPjtpNCvZeUVe
nIQgI4Ow3cPRF0nk/p0MqCAfaRqwTKFtT2sDjZFxnlZUy45eBmwJ1MMMOyN7w3KunId0jeoLsgv+
qPUbZpQh3EvNoNTcvM1wX0o22AaJGSf/83V3icdJsnUgR5zA742CHO8I7O6DRYGp6MoiNnlYv9Xa
Z0qwywUGpFQ1EuvQknqmk6NRD0TGuNmhbV+cCUTro8bGr+3jZ2vb5H7KgDXrrnkw2EpD6Ko/eS8O
JTyf9V4VBgSohhUflI649PUyPfiSbzRiCBRESdl1XUYzrSblMO7ccdC/YYeJI6MZVldeNX7LfiXL
PesjNN9WXb3PH3ZvSi3cyXi/+P79x7rCjqsD+Ff3S1SGkGCQdgm8RMW4bhBDONL0mYk81AhWhP+H
KeFIXgAJ2dE4V9SIaTga8aPlbStyhE2TpvV2gPDGYT5qoHa4+7AqKUDDbm/ePEaQpzw6GnHUhDdG
sAvCgNszE+wMYxkxG5lVsq54uJihU8peX5vmClgZXyvQXkjwV++gnhb6TrhP+GIqmibwfE9bnK1c
IP3MiKnacATXgVEw3Q1iMx1Cs36pKLbIU+kRkp9wbUf1cUT2romouEEEzAOdNcQsJQiU9TeAHlgK
xGyJ4/h3xTmF0xr/muuvh/UtTGkjGlEfACanQMlMkbVxZh5pbnuz/Yl2t+yhUc09NI45Jw+tp1nK
POHLvMCcntHsOo5ySHNBIdJOSF17CuoY0R172Vo7ljvZTBiYu4fPKAIQFO2P566EVlKKwGVCrKFx
oWWoQw6p/8ukGHpVUAktJdu3RAI4OmZ5p992fyrJtg8hXYSv2iGHyc21uwK6LtnS6EtJwVA060dr
2EF0GdkFmdV3SEuzub6ekI9nL2qqi+TzuBZ/COKNlxP9jniabFzdJHmCi7SWcZdVqLg/kNounUDW
xJhXJSyuDPAemYAxKCVkArlIj+5DAZBrV79Xn22Sjm4xknlq892oVmdHNow9kHUaW06yje4FjObw
qvab65Lc1EpZAIcT0ojE0/Swu5wJFr6YteyvKTzs/nOUBeygSFJ82bcOQEugm/ODE3chVa2rRN3P
CwsPav40GwfwQp117vI/r1s2ByE6ai+f9bAsoU/DQEN6SxnuUUn+38dh0TdfEtoixVCEeTxk7Bk1
uXJAyANQ52NH714rBOxwlfgntOmUIY81vdShb64cWL+48QfOHMskaSLrZyS47/P/mBO9GHxS+qJD
oKw1q7igc4yxOw4DGrkrI3BcZEqYoOT9qzUvHdYoDyWcx37Rwkd83ozK+nrw5z8u0OzaCNdiYZqy
AHJyfcKjM5caSK6TQ/Ose9tlL6wPvREDfsxZhslmbSiNy3978QRLMt1B9zI85xG+ClTjya9FXhut
Pn4eCpjQlMljRkYBf7GD32FZoPnPyKAL/ejQdvNwQLDS/f4Xd7ynU2BE88f15sI8fX4vJI1Yh1KR
p2+QGeryzh3Z33rXYcS81Ggdp05H9KfYKG7zWE/ksca9JH9MLuq7or6Iklt60tU7v91ejp77XElw
AYs9pOGVYFwPjyvFt+OV4zIx43hV7jjCwVhvKgdoEY9v2gFKiDL9Y+iHoardFYpcCSSaQXUY2GAx
48GHMqhy5HjK6K+qvASDdLtiexwwFrtCIKscUlugp3z4Kq6K04U6XXeQNDZ8r2SxN0xPdaKyZPfg
kVdXFmTReplfqqVwvLZper+O5GR00DKolvkrdh9tPDegkjiblwhyllN9XNmLfozdoifrBxD7QDdN
mJ/bcjRX4W6GpZreJ+q1K2r6IKzZRT2Ws92NPYz4gIyFr/agNyqi7CJ4WduEY0AAP8siWjdbk6Qh
ccYQ3hUclBoRBL6kM/lJBoBIXmRKgDdGxqNCjEg3WQAmPrPzh9h5IPOvLBnGHRDDwaJ3TCWXt0Kd
2Yk3klwG/CdlbixWXr0Tr6AVqetqc+mBWtMf5fm3b3VLz6OIFztxLPk2K7l1JhG8XxQj5IX02/ou
ilk4A09rF9pYNvvb0MVSh06RZpSq4x8iY7+uVPrwbaemoJc6tspVcsALFQJYG9Zlo5AttYxwtNOn
7Pjcewiz7GRR8w09OLePMqBaTN6+h7JpE7viFMXYxN8TWebMtB3ky7y4C8tz5MTkWTyQ6EjC3sVn
cuM3LIsCSiXTpoIL2ufizkssZyaNVkmDmqk8vx4g9kGlOmGOx6hnJB0srsK+OkhauBdAENRX5dUw
qeDCdTs+E/D6Vd6rUdf9tKsPSH/h+uhFsRS9/py21VC8U2ualImI3jlPOx5fYI1lgcBSPjepEpef
pPNY59uGXDSWkmNVbu6pY8Yl0JrSAsaTQ/SjKe7Od1yvePS6yH6OJji+uG62v5ub+UqGNGf3w/DP
JApo7qibrr4yIGDBlHja0RXVRhqifHLwUaLuo4LPPHbWAdKuOmWLH0rVKj9LyJ/utRnUx9Tgwmqu
X/Bql3EklGeKBqB1xMsvrVyrbRtLt5SHtk1u/VRoom0IYs0wanFmOnHkctvV+3p/WNgUgABaHOuL
opRi7GtY9QLGskk9W/iUCFEmR48MU1DZqzlCzj1D0p4U9pFl0tey/NE6ofcjqxTjRPUBhJRJ3bB5
eTxw4eR7Qsm12kvppBoWbB45m2kr4iD/tjY9BHWszLMUf9PrbZ6JqHZciQvoi7GyudpvTW1SRP5L
d8MW4t6ju8d0N7ZW8ugFbpdvVXoTvk8935WWCtuDS6pXFwUhzBiv8koiQGhjasV+LwIrIcsWyCJG
tnNJMjFHOLRdHsdTm8DCcij5i+wDY/TQyBxbq59Te+8E9vyszP/CLseXQ6Q/0VCU2j407FVMn7Tn
hTcgcSJERP3oR9GoR5gFkEzMkJaYt3/ni51g2fnWgkrrup/BdS8wVllvApXDYrZKHkhs0geBMAqf
owV4ZxcDNT7qvifiK6REjZZ3wfvfMM+3QG4ZnxKT9RUVLc6PZLIGrziHvq9c00sOFRno293b5pzy
UCuyK3IS078ebkJ8O1fB6f99nYsXpKdmuXE+Pz2FtoO9zjU1JEst3eEBIdoLdZfRMmwCMaiUZrVN
G9UbcfV7QJZYI3hiQZSCbgxxpi0f+EcWt8cVrFbjfD3k80ZT9A/i/uXWLkxf4X+3HPCoUdvA9l6A
lk7x1+K+kFaihZlHsGu+W7sE52PgwiZ+CUwUfSA7q4vtS4mfMU0yYqqR0ZWk+u4CgckQvrQNDsQ2
pISd/6eYbRT0PuDoyX+PFpqw348Tv3rLIA6m0CG5c5aVT9IvQeU1Qy7zGa2roVYfAqtULdmDXbkD
RykWdjF66USbuPERH2PNfJYbi62Y2BnX6lkCevVRtkLZeGNOS/NvBOizlQ3nvPHO1zJLhMozbYBY
Hxv3tYripZP1Ql33xw9WExrJr50Pv7D8RxjRj92h1ig9jBusC4dmVLsL5GDMSlP+TzIQ2W8K8UEF
vA1S9XpI7PPHMJcxTUDt9l/n3xRTqShpBxJO9S4PZn0ichj9FRRUF0j+Fxpsa13ON5EPH11nITtq
9DDJmY7dpkSJTgvllwu62wDHr37cDG+a9fJDmcyldI2tIFvCJE3BfgL/rOAYrNodZv1a10Nbx2O2
r4ZK9VONaLHSgArBraLJUJvP8lI35TH+e+w9AGRxOCcopJYp0ReFijrufSgkl7/7hxQgbE4QqGSU
FkgjBJyaedjCuoaYFMlkYC2cQVWBwBfuncrRzUAKyJ/7DQvMTT3LlgT24gA2/gbuTBgj0solWm75
9jLYgocomHjaID2EIIdSYmjUfukjvwIMWSOIpWTnsRvKZ0jmbBTXt5jkFuiW/qnMbkwfO2h/1fOm
uzsxFWdZ6HRzNAT8bHIXgwnVFsjjk5BIv67Pzu3yTGdneRRnsLi8ITwpmY617mOnAcYhQhxXD2vt
jfUqgW4OewpASiN4MXIVXzyk5i0amymxKhfsg040QuA0CYoHVESc2JakIFYnshsi1zmNu95Yi6/M
4xOQDtbR1akxeJudC3tILJWALe0GrAFJRrUj2hNQwXEsyf/Q4XzxulcTWqkKT+4PpqRfJVzWVi2i
9Yn0+NPUALy5gKjR1qBt8an3lTwr3gVVXxJiGbNQwFGnFSsvWx1a4fGHUcFxhsJyabisGOAwEPEj
0F/4QS8thja3bkjeBVlllvPKFTTW6CuW8lx73im1wECNRmXX86QX3JnURO6Xzmi8Ip4o9ptRKKZG
kGvSrrJwXPm0O1+9mcJFhcLM8bC1Em1ZPcPGR20ZR1O8LJ64E4YH5P19tJOKOUmq8oRtIeS3yoT2
IzxVQiIQ25dcEfcnPQbU416apVyLolPxnzG7laQfpFjZiT4WLBzhDnSGqU4NLIQzUNy4sFTrlfuh
eW5nCRaleZzCmR697huBxpXNB9B5PB3sdbQJu8r5OBEdEw4T+7NIr8qZse/quABi2fTsChjnlVV9
aFpRIAdE69uYcpNRp+6KxQEZVUnjL2qSTFL76cmHD8FyOx7azNyuZrXZP1CypQBWJcBpvVBSg4N3
7GGkyusX0McTjswGyL8ISlb277sHQ98LPFGfiKOFexCrQlkVU8u7SRHqkY2Erpb2yPK7QTl//5QI
PbM11POoymI2x3CgzzFAwOl01Y8PE/N06hSQKxWf8YxuMuTztkj/Qw4ckpafIh+dN5qmdmKZnFO0
dT6Sj+vmAXkilxJqMU6eCabdZJCqvQlc4d3NULhdxqz/uQ94cFLIsIlNjACPdoLNBvpFaRo76D6U
EkVWhy9I0CZ+EaDx1y+Ho3QgzLbhUB4OVkh/cCQ9CF2Me1OWQW9AUtgkpwkqQOtXF86a+lWEX91G
FpzEaioOHF7VZahz9j40DIz8I+DhZhejUhJvAv4KJ/zEByWUmGkUXIT6I8D7e93nfj0wnS2SVILX
LBI83wZ5ODnIA3p+6QPiI6YDa7qIXe11/ut6dyxQBsaa981RIS5BYFEf2uRD5dow1FdtoCXa4KnW
TO8TfVRjsAkTf9glnwal8waxK6ygp2oubfBybE9xluwRnOuNMRQqcInC2vg9S/LMU3/r6s7i4vcO
CcMmADqXxQKoO9EWcmG42826DMhvmdfbwI9lxdDd/t8Li6dGDVf4CeHb7+Obyh4vCldyR8ZtIrrs
oe7me985KL2TcEE0yD61ciqHKJFxSD+4PxX3E/FTgPyd0l5Ct+uN4damrYCzrfeoNYtMuU3tdYWi
UTmPrLiVgB6oCnno6ck9YIwc8sswVle0KKn9JG9mDzUtscIveZygMurQnFQAaQcVvyVpR2x6PU4P
rAGb1vmH8aA3+MnHMJIAz0X0cC1Sq6uTOoeVTT1hrCBwrUN5TDj32S+nX3Mnsn82WctxpLWfAph6
w8+GBDmWWDpyPzn4fq199lxlFkELgNxMhyMmVHqfHrFUfIpJqlQkB4JEZAfedNsWmZOPp6yOpIpb
ad/3kp989/Iv82Cy59a37YBdrAuIXdqH53VHQci7KHleFgnQlF0fu/2ArTVnC80J2KY4v081lxVT
uW6R2YeReB5WzQ+43OGLCdfzwQrCY5EygFRjNy098kXcZkJ6R5LfAS26ITst4goeR3wKqbGlytgK
LoctjgSGsNwT1lknZzyYxJB7M77pPvUyIzb7M7K/YJ79+xpBkFcWQNnsAI7cANZBpenU/wu1jTTf
1/YTTpVs85QdghVKhNKUdDe4t6e73wOkAEwWdgBMuhjP15t71scWQ7bwlFqdR6o0bd3UYB6cZjs1
se44OLdJ8SjYFPDGgaqR7pNoK5H2nos4aBm+nC2ueXrCHzbrR18wCgfmkLgTp8cBKx4KhavBFxb/
M6HWRFpwhn8OOyM26QpRn2Dpgm/nWNEqqkbe3UBZjyYx5pBiQ1xtza132NiKYCXVac41P7FipaIq
PFpx2dH7JD90KDpNgFEU1qYvwRAm/S4PJyzzFXO3bTfHFxNrQlohcNgw5LdElVSvqSURWDwTUNVs
2Rec9dZvwTOmvlUydcsl1URmR0LCMqDzDXKVAlBDFIJpF+unhnTVp+U49k4OUIAuwNp9cJHxa3qR
DnIovvuXxzDYxahURX22DWRO18OhJjWYfWJOOav9EPxNiw8Y2JUgL8RnSF02CcAWeYyBTip3r2ob
slNPAgd5tAm22eAqJ25Dtp8QlR1YyW4rN6D6W877ww0LJxwZOwUYXuniNa4drZJ+aMMg6LRF6wGl
UIa8s2h5+7+P9Z8wRog1rfqCoWeta8Gp55ezZZ4h7zfSq5zGT60ZpaeEOC6CJGq9WdODS6t8A21y
7LDSCtmmHIxBqS72VKPxvgsfiJCfnmeQWa4fZ/BEvFituSCF9AngiZH6iWO0lLa0NjEe3XuP3eDz
nJgDgOPXtrrTUNGkoUyFt/wdolRcHhTEuvjsRvpDOaHWBIKRAGGORu+d9AzyAi0E7XWsA0PAYdQ7
72OWljLV9xSWVUmBq5y1mWmpygMIe2XqMypoXfJI5e/JnSPCpttMbfs+6ry44whteBE5SWfzj7xl
pitQlm66T4j1FXHZ+LvMnXqJM2XmxZr9huQwd//Dn6pNJ9xZC3A7kmNgS+DVO3/GMX76hLVzs09E
m7dRXu83atKTCgujEadqxZMnBLU2SLUzoItfdkZWahtXAWRFY99HF3Ko9G4JNKhtqm3I/ziyvjvF
zZ+Hrnab8nEm5jOajJpkYJ0wy6j9CXbpTr2EdW4S5lVdTZH4T+LKa3IWR0nTCR/yc9egV8vpQZV7
ASZdS5KDcb4asG33byC8LN8LVumvfOVacogHwnvXaw2/kHcE50CnvOu8qPjxxx6uc1Ru18+2LWgz
2q/1Yetw1AjHbl/m4C+0vgOy12lU9oNiHua6KuVFRReWh11M+tjvyIJYNSL7RYfF01/RXhxPPJP8
J2pT9s369/lvQQ4iaKFHMTVbm53HQJwbEbFVRyTfJzznUYNLO0N6fg6diioX4d4BiDAVOhyS3/fR
L+UCsigug9pjlrG0LGqYQUuxF4wJ2Clzk04pOGvzAv2GIv8sPLckSUi3V4tvRvysEw3l6/O/Pg9T
/NF2WPvcYz9/+AyqZ+paY5NLCR2QkS8LCvXvYQqq7FV6kiR12PwZd+YFDgD0T4yLmjM84VQNxHag
/PQyba8iLy+lSmNfzJtktrAyMmSTGQ//e77VvhQj6OFRtHLIxfFHLIDqFbbQhvMjSmpllomm9Zr2
AcBRAdYS6xr8lDseZwPLpoIjVXcj2kvyCGOe84tEmnIE6+eQSUrjB861l7LNxvxq06I+dEi14mkw
g9s/BNrRYJCqc2t7+N4E4/pWIuUjl320jHVSRsXwSUN0iDr3SNitE7OB9yhxJ8eD1DdKb3iuJZq/
898DDyNLoyLNGmunGeUmFXdJ/v4mnd8Rk2XG1+GCm+TTZSaT15kckZIkzJUxRBTlJEiKLkf6UZF8
vfNy7Is64H65wOsCu/t1MIqDGCn2ZGCf2xpi1aUXLbKShWe1jhT2x/YzhT8V2xK0V5vAuIOH8Zo/
27z3b9n4CKc4wlURrbS5BTDoELM+8kq5Ivwryjhj1HkOLgPRu8wZDUV+DVkyeiq2iFMeARrHgFEx
Db2Fl6DcrqIQ5VtV+Zs/cbd+xKwhuJ4hf9bg6Kt9KUPfLWGVsd6ADrOFR8qQwK+TKKy13D60Rs1M
e+NggfjKf9Rg3ntkKR7szimGjyH1A5SMLo08vWKYr7UrCrKEFKQRWoP9uWLVHJ17XMOuN/QXsfhV
Z1zGPMXWjL1/nV9KUPFDKgTxUZHD6b5xFUTipF0yW40BEyy1s0MCcfS3f3a3OFllhDXtL7uDV+N6
iUrW/arzOQmsJbv3nB/hYQ8GXdONK5f4tNyIWkevhuT3yNM7Q7pXvfXr8Wan0d8r2RTpsTH0xh0H
ge4LOJv0pvQBogULwbPwmuElEczA48jA3qUM6S5WgC/Oe7P1HP9gSmOuSwSXlohYeBVL+s76y4Z4
15TIe+Pscy0EFEaBHOyipFoUYWGUHH0Y63l2tfumLxLaO4z/pRzV61GLU4Ka56TkN9KK8oQDHjJ3
kVLn0dSeshmy+cgh30fnR07McpkzUzoky6YR9fh1cHdrqXBxqAUPCYmjWdYm9/b4odtxZwZ1O9b4
Th5fVtjRyOFtz92PGn2uCCgWRASGSgpynQ90fduH4o8kCbuLU6AoHQhrd3uVt9LI++abkFji55fU
QwOCLrpHtS+2gb9d/TJzyNDsI96Zczv5Kqnl7+jiUE/7vlrKJX2my1Se7ActpEsxtbRMY+V3BabL
yBcD2UYNAWmvubbqVXDpV9A8B4MxcHIlTgg35ki+RRgC4RegymyQ/AvHuTrMjE2MF0GBh2ILhjC2
MC3OHQ95NH/1CH9XfVJfWYX87BORsNDmkhEZMK/ot3hXt24H6w+1jnTLE+PWGx01ccFMiiqHuADi
m3w+rI4Ygq8A0CQ3yzQ2zL9DUuQ3cbasnzayYPXeNUFuYL8BTer0jpj/liX/eqINF4W+I4/gGLZ0
fmEshrmj7ufiMbLcbLM85GKFbrrSahIwVazoSxi1sZzoXL5qLN+3UPgV8QGRMSFj/mMft29DFQIq
3Y6fJJTfcvD9dAankQMrh3UPsaORhiS9fwxqucV00PyysFgL83Jup4zs6lVCnBJjMrlMm9gXdoUC
EyDCkkKr6CnkwCfMwzgEZRg/nA/+FnDk/pG51YZRUwpmi+bOHJZP01dwFgTEDOP23PLdyEjDoBQu
7If58lDZD2lEyTYRoB87XUJEiS7BS+9+G6QXYwG2jtEywKVGCtlVoxFSq0CZXN59gMPcbmqagWyM
aj/nOzm3AyvbmBN/5KjbebY1tK4is1TbBBW/7eA9YhTnUJOfb8lnPncLa6Y7PIQ5Ed9WcqXwgZpr
SFgJtOcqCAWfr7Mb59X137nyn5RfBJ+cOFO3sB0e3Wi5UMTgttfIvOEgpSBrv5u4jj7yhJ2Ss3So
tXoUhu4Oi4Dv7sV6YQ/+QGWg2rq9HDmkr2PLYH+Dq4o+NoIYOt2uQDkE/C+MmtBe+Ft0e7se54Iw
+J6UtTofPJc6QGJcA0pZdtfxN6Z/Y6x16Q9JqmvE8IgnuDX5PEIeYKxnr3ggMRmnyJ3KqUg4IiqL
5nkdk/GZBROsgwDOmmysG3kWBupioJWrkgryEtmi69CDzJS4dzoGII1gUJJTgFQEFwgCWxD/Sqld
NexeQqLP5jQxOXSdCK26DZh/pp5HjTGA+GXI7VOjR2MzqfkmmPPGvtUSMcwI4SZ0KqzTgeGH4oLS
UlmblGajTOLZUO2HGUyhsPwYgMNA+tsk+0LhT57gxqaO7hMlScALFhc3PSGLeM/fhVD2AsQpM/Lq
fC3Szm90lfK53oYIWCmKXLJFvSHkXBMEbBYgJBhu1Mo1KVk9/ycVwkR3PKu6n6zbw1UjwCo5SKsM
BXVtKJAjspcgPYixRPwOJQkAKsrkQNqam+xb9h4beS8nkJ/VUpXoVuBGPJG4YO/9CTAbHBzUvKSI
//8fo/pAWMsfBpmZs10IOCrojr3jtqcfH/VBo7uDEwq8X7xH6cgfqatUS14SWoVF9vW8vUpcneTm
Icvu4PjaKOz+EXfj3xTE/jrCoj3MPNrLUgCiCutF/Xva4PzQL3Js809uG4eSrZKslMHjeA71nIVf
Ho64VsRVyGI+AP3AxxK+Lf8IrD+JmWevetC6eWiCGruLPCQmshzoeND/X2W3Y/DTNYIaJgc+jV+J
D807HtW4a1NHwl1PxqXkn6/VIgIyybS/PBMayAlunp1H7Eo1n076XAcoFo61oYHolaqO5jA19gkH
pHQxx+uHTjJEww2x6h5mz8kbn8xPh6phdi0RRl/A+P3Hfpbq/suKwb95uBDZ9iwnQtqkhK/CnKIn
4xOBZoVADH87goV1EbjqbiTX5Ax9qId91pomTqJIJzhDwMeWGAADp9uXjudXNvhY8AQNrfOggLIq
MQITc61iD68V6qlOhJtLTxKDOZcTlmLHHM/u66/Lkf5otLV/WCpdfgGVQXBa3uWRcaNUsMNJdUot
y3I5hRQ0ahimeElLIn9UAt0MUhi5Exd7Obllv+vbdf01ABOypmCX82EblanKHvHtZxhnEAZ8FxFM
Dpa/KMrk68upDOxvi7GaW/mrp5EG6D6dyra/jfLtgOGume41BmP0LOWjoZZXSm1Ylj6oHlqcpD+2
Zp6hDsN65pOcCJViFs2ERr3eR0bzAx5PlCh/IEkzCy0ZGna/DShLXO3+xrq5fRhAdCURt5Y8SQo/
cXJ3rj8GtJpYMTCA+c2S8cO7oxzzr3Z+1lbQKGi1NnnDRe9ZXS63v4xqRwe5Kr5FUMOXVVjR2nS4
D1d75gA+VPbSXZQ2wZ2z/4iqmhb4bTOzLxVArPuNrnPL57cStPNfC1HDpbybK8JPQdG7WOJeF+K5
fz2v+UEYuUpi+u28C52SjpVTdiQ/C+RlIxrXmi1sotkaLFfp/a6YEne1TkMDr8yE69lUzv3sjhq3
wm/Z8aDHTGHLZ8ovxgsYhDLZSLxr2X88WB30cIRUzbMdxvUt4DwM0/nvmuelfFB5XdV49HsnhHO7
NRgQfi9y1aUCD35jsjTE3x68634K0JFpD8k0abR0Suj8l/qia5Ckyulel+zMPOSA1g9aByni1S5A
ZzTllOFdMLfJbRnOOlzbZBbzw7bKO3LNN0Yn/9cM1jjMBErgtaWCJw7kOH3kmmndlvtv2YvkOms1
ahD4vKPr/lwvFfzTTLUFr+Mo2IUxXgdgaEMB1aIrdhQilCtWGEsUsjYYVqAcHUEuqFmiSYlPB0qw
JIQFrDZOissDBIib5EZSKPfoU5LPXHjr+Rf1E6CLrS6l+ry3w++WliOVmT53+4DQgsDBU0srNNLn
z6biYm2/0LZT9L98louXVgIMpr1EoTbk/DuX3eGHWBviQOGirMwGRMEYpbNUox/UREQpEQr2DcRW
zUtIc9OcF7VPZIMUJi8ejsq+9Wu5PNyzEOMTVR7hjKtu2pTx90hh9hKafMZzC/OT2hQsQzT/mzRa
VR/qCmVaLghdBO7kgvvQzksuLP6MSlLuWl6InXzyp6m/UtAXc86h2cDRkJy540HqCtaQx4X8jfni
TblFiukU3Zog8tl1pHDzRobmQeliV9lSvp5PGNnAzpdAB8z2+Ut8bDZWSojIrvswg/bsSoCerVI1
Gq/Gt5oOvvc0i8jcyIwXMB9O0CiJLua9JK3QuGA5VAgvlvIciXr5kQDXSiaZSfLj0tHStgC3mN4l
bnsu5lzQCgWaPguV8oyo7DIeU+C9pnAgebPW6gIpZOSloeyVLm4hc7JijgAGkO8/MD5EJ8iOmitG
ld7lhpTVqWnUhPuzewjnpPJpHldmPOpx397xZbTvquYmLMYSEYI11OEl/3/cbNsljD9zJylj0aR8
xDTDpwYoaPWG88a8LyqoICHQ8Mw/xIWzYIxkQKXX8g0vqjTd1n1pQz04mWiTS/RYreT+3cHteJHD
9dTJp2lnGb/pCqUWOlx836Yq9wbz/9i5IsDTV4dwXXEUbMK6s2q3WCaBhcAezqX1+I6u+FQi3lqd
fgt9LuOdOPuNbI/n0fd1pYtqg+4voBIH5ycWK4FcXp6leruIGeaA7ewH00yaxvtxPOSYBRKMyJT+
/xjIR8QYF8S0WiHY3mYyADAQ6Plk7EBCAezG8sbOCyhFxMtckvPMvCnVowosDRLgllf88CPRtnjV
UbO8Jrf1t5BWsbNIobEP2EhTNeOxL+3WDunR9o1vl3M+q9UkQIE7QcZc40z6sELKxz5FwHT+fPj5
YszzD+bTIeXR1hc3wtsZosJgmrKiMXRQbyqby9bqV8AxmUKdyunrGadpbbRw6NBEamAC2AYBYKkH
RgMmcvD/kh/ZNKKh2w11SPtM/oXz8E0tdBotyvlnjVuYPUh/dE++t8Lh6S46O2XmggiYMk9f1j+a
U/oEKiC2DRaMk5bDhJgR/MhTauvH4ITzvjnh0OceCSZpfdqiqeqN+336NJJSaLKgWh9eUkMF69Bg
IcKpx6Xh65NsiWeJ2e2Mofn2YDzn2vNSMgmcEu8oRZEEr3QM5R6me16j4tc7vPhdGa7s8aSyI5Q5
CFExuLdZVFiQZPL+NqwJqIwSvRKx2Lb0+/hxqtbbjsYbJYdFVSd15h+mgi8LVqz21L/r/JENhYn/
qAN7JgL0vEPnSkZdGh3rMXOf6a7JCUsG+nRsfYOEX1O/Hb7JOH8oWaMxxHhdxWspFHKdpxdIxvpm
z0SNiYs1v3DFgsDTMDACIs78p8Lyt4VDmHjzdJQ7MosIoTiwJjiIDPVIVdH/IL6xILok65mEeMJb
Ne6RLPHGJIpYdepxUCFjyXxtLKoYw8oFiXUzxsZSx3f/bkT5zuXM/6zV2F4nsLsrtsWktxzXxdQv
omNEYGhxnvcfNp+xjbfYcETH45JuSOOPM8YmyRPDvtr34fuZoIRyzxHy03TVRVlgHddNej0JIUL1
3ola/bWSzucE4a93Id+uDgUj30FC4Xr2+R2XMsAKvs7M8B7sp1S6F940ihEaAgcuJVnKuo7tOujG
qfrrpRkVWRklxqQCtcHnNWUNAA1rFJWEukcYyKYv9SRZrhX7Ir1JOdLI0vhJSFB1XMRhHgchcPar
t9ieEdp27lP0TCaCjPl6LU+hIfdi3FKHjWU6uzLHenvSQIBF4xmOolk1fCw8bXftR8T3diOyS2dj
b9EPy0HwxplcJc35Tx2KwANtUQN9IBC2AIkqiaH+XK6wkUZXKmzwFb5PLJixFAAa66IJLvYxUAS4
kALFa3eCFTACLsHSxEvyUQe+QQ3fpEpHU9AOK41qb1ntHUwoGYrP2cWS77O7SnSkU+s7PbpdQmeA
A2OKRNVHaiuBfvEUvOC1hkk/VFPrPFzAYyu2F0ua5SGOMWNwe1Run/By4HLu5QJ07AEed3F7ufrt
mlaxUQIxfWx/Ba4KgIvo0ym1HpL2u2RKrQqUdFR9zamP3K7qz1H6kl2vmgl3jto9TDeE/J0jMjRS
yNU8QQLwVALmdI1Gp25xflfu/DQsn385+rkR/KCzr3tPP6wPwhsi3u7uueE5PG1ONQ27PdURGiRq
7MGcDghd/dTm3J4QLkfNv9BS/erKekjN8kpMgrKEvW1E9bD5MlvNLoNedql4KnuNafacmWdk6Axn
VbWfkWn4QLGm8v0nGy2N7Mu2G2NVw/w0m1BoVpaq+Pm8LBc9BU0Er8DyAZW1ecmbSQ0S1vWwZ/2T
/ZYiAtTwYdn3IRpv7TQMpYWObkvhfC/QI2Rkc/vcoDWYD15JmtQYJIcRehvb3jFGEeHNOrVn1Ysp
f9ZtV8yXjriEbuG+udj0x0UUaiBTzFguHYT+JXMVcI1LbY7vqmhx5KaEvGi+3w5PX9xt9HLaxGX0
VMCjjv6tUYNpfvcEzf1XusKoZcrpW8vV6ixDs254FHEDrTHKUhhViepCSa1685QN4iFAsbNioPlN
WrLXNiViJhx6+kn4U1ek3mgMgOXp3Fp2MRiaMrOi2EI1txeI+kYt09LSYI49iUDcZ6+vNQ1yDFXl
WZ2M/PJe4fInrJqJjbV+mVGcVZ/q/cQmmmkFvOGZpQS0q9f3lG7+NGw4UkNJYN/7Dl3Aldi6KYP6
NEInpL8gD4bo7LDmtO6qeOPf4YnXa7vaIGhGBZYRTpWjvoIzFOUYILchwgZZO4eHgchX+otY6RXU
t/GQpiTySPn1Cai+rerkXI/YL98RJSvLaXkkpE+jqWHdFj8U1uXt3gYWybIJMVGulw6PTz0OISaW
9Q4P5KVLHSM/VfosINreXiBNelf3cB0tFQUUSP8AZy0PNIkppUVyd6ZmGPc+UgrDp0yyQDwa7qmj
rJs/TZy6eodUJRx3E2RG7wHodlNPQNogKXVVswqpOtd7C50bwolZTKJKw3hV5Txtsu8tvFoOfTS/
QtMObDC8aKUF7IEzRGCg/ANvwL3eOeHnh6igpYwdMHpJInpAfg7AxtcFKFlLnQT4rUrCB7bJGBY+
+JQLPYEIo2fGZI7mOe7EyBwhUdWE7safduZdmqbLF+LGUrEAK+5BLzhm/dXCacbELdU9nlf8bUIl
MK0/DZkVQDJU5D4qCL2sMEFpZ8df5dP27bQvHQthl455+GHga2l/37/4RFH6x7FF0q9/4kPTsL+W
qhPAQffT4l1gmN2yLEsNQVdcSDPdTFOeygb7nQaoKkyEIKB0yuqsSFxoFnyI9GibMaaBHkdX9bh5
dMpBJ/35V2JUpzrMR01fNH0Xb6FaUVsSJnSKC2ztmwuPPI38Dl/q/8wbTjmYpOqvzHF28RPGeEeV
F6pPb6STfEkt0OX9iw0nrdc3+KKI+MrZQN6LJYbTB79ONH4Wehc1WYqlM1zym17I6W+Y4gtCKlqK
GVlpMZ5jkjzuLQyIdPpdeqej9QhRvbe2/9iG82/rmm/OKhrzn10RWBXCtb0h0BjghQK4NFbmUKLG
TY/YnzjSoYVhJGVjnHmGzeIYZJYqRWV2hl3pAYkarXbMVgsoGl1rTJCOG4LnjBCf1ZzpChQt9OKW
keWyIdFTjGTfJsuSVUiR4Rzj0eUHfa3xcRkxyWbKZPNLHyDDV0faOvNcqwl0Qx5gnYX/uW/E8oZu
krrLEz6jOkAar93+bunB/F0s51gOWAINOdcctxlYFgWVIvWZjQBwgKyABhsXMDSIafKPpOdtRs2T
BoyRZaOBc6+Uzev5RMBeu19ZFM0vydlhY3gakktUjjbIYR+hJjOkvMDwfAYnHcsxBVO2Til6vY2s
QmuSS12z+pMyJgd72ywfTIdruxay1JglawA6mKPNjpXaoFqFrT+DLf7obK6P8N4gzCjw4Nm/a8x0
WA3Onq4LfDBWiJzVSozTq4K9Suuz0I8KP08XKDnq96vVClLCto5TGIxzMxJkpoyZYoBytCk37bfS
AW89DLQnnBZoqo5XA50G3gtpttHNhJLYd6WHs+o1k3XKg3i5wVQnhp9OOT7WaG/qib5w6EiTjLjY
tize8OjOPENFc6fuHYFvEWq/xJirpiRJH/NxQryNXBA3qhKG91xtdxga19aBcw730Ea6Jz1lRrom
Kggh8YzwY03+H1xkqbDImk7DuRrJZEfhW1ygIVZrEXo/87KKcn3rA4z8c4nWsP6liXpAtZ+T5inv
3hHF5QPD76x1fn9lA+dzNaAtOq/CtqWK8VccVZX41FkKPxAeLsqnYw2LNLNFVo22w8roXyGQIVQ7
O530NfoMu2KwT3+mEncXRyWxhiQyrAqdewG2DFZpVRXhmOV4jcNRoU97CGolZiSDRwOuPsb7KspS
r9pUqncXh+FG0vEHw26lQWvcGPrySgjKbzydpmvEAgdr2cJEZnxzqCq2YI0+lH+pkJ02HkH5RddE
Uck4+0ivk7QypVXT5p2tE4whcXj+7XHuTP0nO0MwOmmfbNTKcNdlUNDixN+mFWisC4K0gtavaKKt
ZVndf8zcrzot+A7LVoCZ7gq0DrBLZZisrLjo0pv0ONwrAZP511NVQ5rJdDFFFm9T5l3KelkXdt6j
bjihGbUcKT6p9+qmv3knc5pFCxXIYpWyR9SdzWMBOztKRl+KTERNaP0fru1odv0rfebnOH8AgPR/
chdN0cXuuqrnMdjVpaIQhMN4BqMLZ0cFH8yTySzv/UmNcszn1Q4FJeDR3jeAaQiuBNL9KX4b0jF3
ewEJSiZ8CKUrG+DQ29E26A9io1n5kmo0yXznOkzNiCVQ1Z0T64PeHEnTtUPxffloSG1uWfVzugRV
EpCffHb/lLelpnCCT3tt0THn9p7G5WgDZ/nHAfBCDDK6+mQiuCS5s6p6B3BXInyTbiklBLhRi1Kq
mg7JNJBhb8ErpcyVe4hqbbhpPU3JnbVD6m1GJCdhm2pCTQN5lMjQNLh0wEMn/hBjpBI59beAc0p4
mk3btRQEdL5lDPrRvVNjKewyw4KJDQYSoGe61XbUSFmc5OnPSN1q71GDF3rjsPj4e4M/P414Dgt8
iE6dHm0ZQ0sKlFLpkXnfc+sgIiNTakZG4bWJ/gc50fMxx7uK1x7uR8HrL8yZ6NY1sWxLWQtWhDQ2
4FQfe2DYpB56QEHJYCwPVKXPK/yOmJ1yJQff/BEc2jZxgOe17ea4yUvUYjwSLj4PxCKX1D6/z9Xv
/Nh9YGu2zmUKP/7wwwSmgI1bwyS48keOn4xu0/rp2krNB+ZiSuu7rKTeA8GAaUkLKKbb60Mz4Olv
gJolE6HFl+P+SO7s6UbQy7iq3W5m98X+QXRhXveXt8oDEnVwazrYsYR/ZkZDuqSZp7D/HTDnA3lZ
eYdMidqDmMM64IMHJBErBhrswOT6fktF+zykX7RpwzqvyIdX1lTzNqH64mMT57QujyO4HodNtNa+
v2+DLnwZc7fM43eHDl+ppZ6PFs2a8pZLoGVWyxs9E6gx3Y9AFztOcr0GMrDLkXdMLnSzc7l7r8kv
2Jq6fJL6rSsacsUqI0b83xNQ6+8m6VLVlN/t7sO2UOwJTaNKmwtSl30LBWZeFJ4vDUQyI96KKW3K
+TKmI/Gq4G8F1bMUiC/yMoSSBEmqEXJM0cykp/+2EIkkXxd0PEX3ITcgbPs8lZm5HKuSObGlMSY2
pH/dcbGGnfhVvdoNhwQW4eVWpuWIfZgh7Obzy3EtBLWKw6/zl9fCVIg5/J/XHf+j/TrWNX0juZEr
tUcQh64TCTak1fp3IaOoAg1BQJKYolvEb+6M3fjASVgFvve2HYjao2xemQB5EdYoyBvZAV4AYUII
A5iwVKhXqh9ASv2liKBT3lUIOd6l0SzKYKP+RaHG6m0yB1mJawaDo82e9eP5mIjC+HFhtmx4mvfR
ct4zf+Zc5rKldff7xNO3SDz1qPOH33ZYH9YKTzPrAwN/JzzaQtBeB8NsKPIPnBA3PX5PYN74mKRv
/nlbaz20FNWlpeINvc6G/L2oLxdYNuSQqOJtrgTADJZU3ARFxnq7UpaH/Vg5Ha3VYu4PvdzwG02f
2NTbdUaFRk3PdvjU09c0H8Lrp1pJRlIePDXDd3QCQK8VLAsoMcXvGvS8ZMeCGWMSCq17aDhSV/oj
Nl0yYBxUyNAjLbuRIXd5UjV1Hu59JsJ3Q8gFblz31Jxgrt2TUJofCShJINrlL60n1ZNr1+kmU47S
xamBoRSyimY3SLETeM2BZe/dPlrp7HL7Camlmj1mKZHSHTa4VZ6u2j2iWeuBTp+fuJNXjIxwQ0yQ
6V43x2iizYGADBwUc5rQVnP4q9NfwMlEDAw5T8QMsiE4patCiFqNe/7jGaa3hql1DdA+32wdPyjV
e+rp4KzxXJsVgVNIq3MG18C1pePeTMjnivdz16OPp7LDCtcvVV9pffhCk24wGkJTufyEc2aOGzBC
yZUFvE2ZImM3dB1BVCYJx9F32SYzlnrQYdltI2rVI7Qr74uaXW6A4JArlv35nkpuoFx7xYFpwcIl
8+wMLJAFpjqvd7ymX0Dm04u+O+fHCVj/+jWxtzlS9Cj3A323NonEBaFk2jlzQXlRn5rpsIHi76fN
NUcchvQ/NpOAKCgj1qcOCiN2NYhjnC9xKN/lFKXAF6mR+foG2FTKKdztkrLbqoVhkZsr+sILsIC+
hxgJZrZQA2dzy/J1NAgd9/4yRt+qpTYhP3+tsNL+hX693aSAUfaZ1i3+crk1VYIuKpWCgkMLsZ36
Fp7m91wmBEXtH46PmdnSG3sayMHq5p8eS9JjhgJ2ikg5lMx2IY76TciUNehw5WtlBDYI/9Ay4RDH
qG2OnQAvf6Usq8bTQiXJ9xr5NgrN96uEvmSJqVvoddHBl1gLqpw0ON+cPSrocdKZ+MqPFDh8G/IL
5KRGVOQSU38XjZVaDYFiurny/cTZ49pLAdPDyZhksGtJrgFcVq/Pm5Dqiv8G1NP9B5YpSDlzJI9Y
3y9ydYmPYSsDd0EJYqB8M0VIUuBmgJJA3FxtHKhIlto0uMTR+B8kZZ3OBlm572pj/Hp/w/fCtnmg
ZgBCMLg77ytwPH8bpulK/vwi37CiJDL7PF1Xx7FB8qcxTr9wGTe1ROf/qXr1xajk8rj6/2rcovvb
Znk8ahMpvfeZcNQLuSWTHAVDjggYgToAUCYCM9L0U+S/FKPVgsfXFvwYTPdRyuuFn3B0BJ1TNet2
xobxmD7saXEVBKiNhNpYYybotJB+pe65hYpet9BRkNYb6V+c7JIvyin/HCK78xbJ+rYyDlFfNJEH
lj2kbSrh524pv7OTIdPYOW0ZF11bfoiM5HfuGXOfzD+O4pA2KEJG47M9kClTe1Wppm/Lx15+bPGU
rU7t9qhv8QMizLqrdsvAjdtJjkWRe9BNRGC3UpMB6shZQUDIK3Bx18JRQsKOt+5+Op15qpWP4rgG
RdQ1CQf7+sw/RvL8dTp/UEhh113XAHimsNxFuQn13O/a7UBmVz7m7BDl7mfIKRk9DC5UngXEyTL4
k9568ifGi/KmtySM2Xstmc9ZtofIhFQyH5FbGt+Pb8uKkUiIapXWshTLqoN6S/QF2OPJpXoayQ94
49s9i6iVwDLJwWMo/p8LQnlKabUFjMnRi71LvmcwCGqcoe9XvSjTnJuU0XiA5VvxMusgKAmMYbv/
RrY6qMUtv0qLMfYEnfuX4NTRFjJPXU5idegZcZCub6eMzTwkVvNuYNAtzTTq7nkZ76nBCUqwsjuV
lMKJmbnirkBYhTwrIrRo8ZP68WeTiudw/JDgWe1ewr1U4+Ah6V8JU2eSoG1TR2xYzEIZvnwUI21T
jt/0KEANIsZ7++4lXsBMPEOOrlpZPNSNPl+DYb0h2PSUwGJ1slxiwYMTuLJRsKKD2NQp7H0NHxbx
Vz3c5N+LxQF8wQIAvlpAP+b/UdNEJaoA65z3rziuYGgctDnZS+JZf96PL3kM4icuf+y9Mmvta4JV
QH7lMcJIxQHoHfs0I7JQ5zKAXRA7bF1IfwvvksXZvLhpsAgXuPcL08U0mJUOX+WGw2WYXdA8o0q3
zfmwKlqsOSUjnBN1IOYmhsl/fkW89giwvbNe2DEcPYo4Z8RkNfXt8aQ78lSxOFl6x7IyCp/7lfyy
jf0coUtEIg31rWxWE1+Pm8x6Qemb434b7pugUVpILT47lKnElhIhzUc/eGFEQGTSPFfpktsfZIBO
CRfNTqUC5EB3xnffGHi7s6pWT3g1xKjTg7B9N6oYuK0ao2+BO9+flmHGn1zYNwRIcxvScLAIX1Fl
FkDKRUyrlkVA8CpBppEeSvQUxGOuq/9Q0T+xK0uJNZh/39L+/q3zmJvRr3fqNdoByGkSN0GGq5Pu
nEAarXxdUd+zxCwAM/FtthJkUuG2s8awttXonlTYFFNANUK1VO/e/d/zodokQYrhjgkfGiB7CO01
HeJIQtESOoAB6lkwoYxKLffe3Gcc32/DeNSn5hJVbt5Yhc0PNUNmveacaI4vFkaZAcbpERrYBkUc
+1m8+23cDYF+qMshD1txc5EhJzTTRBgn9SgveTcGvpnUG5Mh8v0HdzjsrusrqQPwNaOLlSmNp2Yw
fhLfRasGMk/YT8CSujYuws2H+wLB5gF9Z4XDBx6JcreLNteb1KKwI+p2a9A/ckhslv6H8/f9rNBV
Pp+KMwEvGyPcoyRkcs1Rsml2kCsYSqrk4w+zRe1eNm+iLGa2Qvz4e4aYPgUz/2XgvVHM7TBIBwTc
9H/8Akm7f7uQIcH/So8ur+S3zef0E3/LzV/PNjm2QhmjjPaxnPcsS3mymGYqxW3CiT4RIYRwbiQ+
CRdqwmAI8yeMNKPqP9CV0358lcDOo3XNcuuKJvr6Ib4RlvDLeSwKsXGWJmVyk/FATjUQ+vRu8Mek
FOReFXO5qBYkhCw32ivAu6u3sxtRVNXeXxyveZ8awOa1t+Q2a+LNoR/uk+5h2BcAZfn/wooL+hA1
Q7fDqIxj6bzmJnIK2TxukYnp+nOUBgqcsScsTtul9SYZwgCVg3TekFC0rTAygvjNXMsLjET28R8D
0LiHjxOEpBxdk49BTluPiDw72im5cOOaqBz2zbydEQ0zVJpiFpaUtOQot2hnSWIpysL2k/gE103B
wxAvNyibAeLDTp69P7+SVsgjN3vDi16S8ZCNKjn9oUMG8RZxY6ZGUpfCtf8bMultjhuc3oo1ZrIh
yLPWlkSDnKvvA4x/fdHuwQxW7q2PasbGlu+8SLvoeMM70CAyLmrgsd4Peen/nYjeHrIoRBDghpSK
X5OP14eXJK4VfFl6oos1YUMzI67IxKcnbBBT/ZminLhOYv/5gH4O7yzAJLjtNOtmcS9rfSKUe0hi
nE+lMI1tmLbtL0sBfqxiQXZktpRHUUvZSGfeUwSzgImoRwec24Sy0YYZopjG0wc4X3Xai4OZMccc
0l3ATBLy9dlSYiH+YrlaMuq66OuIbBTVdGz0iwBYMXlRCrTTPM33aH1LX2RD9Vaici9D7p/eXel5
/EREIAjVYjV97gSGb2/CWB9NNJPjRi2LzHPDuc5Z15Hp7ZQBI8whxxPzgAOQ0vUcCoXRYHceKVaB
hPaRBS2EF8xz5aN5Aw57XS5s+5b/zYcpJk0OeGXIO05zEjJ5ReWbbU04QtjtqDGqFVpURkZLtgzs
5t7V9K9p6FeJTtG5FTe7dx/izYzFZwHd8YAxKVSI2g1+lssWusDFs3ByFqKgg5/+UH9CwoOhUDhp
J6sw0sNa/lHhlSDodVY1f36Ciz1EAYOp0YpdZIR2UwQNZIyc+pT5HrO+JVcPc7xnvWd6YOyB3tDF
pSVxuPUNj+8+9MJmqMkEVHKetCpIDiGsX63387x4B1Um4KL5hjN48q1XDdBTNQOZMKSGBOhXk1Kw
6ed8DNdCJqzCge1lL6oOV1VaLAjQa0XVHq/ivSMotFJLBJ+aAHLhEJzeb2QQP/t/bFhodnaRy/Ln
R5CDwGczgiyGQNX/UNLHEpcmLBN2LFeBtsu+YaSbVAcXZg6GJa3g5nCt8SLZrm0ff4+sQPK9mBKW
g1e9/imsR8dWp32lTzCP3QEw5tYDBVdpESa4/+iqKwwuYaAfiYBWjWcPOGCiTxWeeGvgJsqkQGVM
gsP+HNSf9j/F7IXSmjlNT1saA2hxuunUdbrN6j6hS8oKybaVx5pSMtx6azN5JwC2orzJGCLcMXH9
3NLP95J0tle6TN6JcrsF774J9NnVsAWu4/Vs/9f660vMuNm24BDYlAPCOK40wMSDzjYWl/prWGUU
GJrmhoFBaTGuD9Nd79IhzH7DHkgdJGb03BZmj1uXZnRleHLsxKVVDYkwYMh2n8kZEJ/wesnPN9HQ
O64DnNwCIRLXKj7bY93+lY5dFquwo+poDsKMDkmeIt/8fzOSBY+9PyYjD2dgK+GHlvXC58RnkWLl
oqkVriGriVZhipyDBVI2ZgZ0lO5XxWWXNCbzDS/WgaQNYszJreMaSu0q5mgGi0crTkYticutU6iT
2FvqTKxtn2ncuJm8m/00+FZwFS/rKFk+MErAAVu6dhDqSueIAGax3ikkkPiBrley07tDI0ovZ7OE
tfmQgvHiYplr4kaU4IqPqwodMiUe+kFKJR9l5MGLUTnZlvViJYUXnLV+sLb36FDUJ5v14Wos1pzF
ShENL2Z4awM73CBOvL/Gr+xAvftw6n73Tt3HJOom12M6oInXUGLOuQqI/iPVfYJuz9eu2NXHfWWJ
/PPOIrUemYvR3Grq+elObEUFtYXgZrlYjaRmvKb+iGGYf0EbbqubqDV7tzSg3eCESQMbHMfsvxtY
alU4BCPz3oMulTGqQCPWNZXKISC3LtKQk5HeOtvbH5lMF1eFZqG96WDQAf1F854tYvjY21LYlgfo
RPGWB7et70Iege/Bb6IfIfuWCrg2UMjpWlKsBRzFutMEPQ0uspbF0PlJqmaydh4ntc61wKK+Shss
WPvMZvrTn1UH9F/OU9YrHkg+XFID7EnoQRk88luqNQAYp2h0QHK+7FMsTxFHXrf2o9jTrhXe3r6y
XR+Rmo76ON1eAvQJdH1n4yzaNFTWAQ8LrB+RiYNGORAeUuQm/6vICkkh6FM0POBBSKbdEl46/LxX
I5XfAoCKPtNibOM0x9oov6VFwy2hj0ULdHf/iI0rnoBctuNkMQ+3NAaesfjSZAtL4ZGK/h0rnV5c
Ds3eSWauLWlC8lBiFxty7YX2FK86d7BZf7sYVWrIZGAiAZR+W/ipL+sbjGnO9XWBx1jBG5mS8W69
0oHShysaJMFE77R7Ba17gIRw+0X4H3RHtaqlFuQqTLZ2m1pt9EIWPugCvWkF/sSrfrzQ5JVlb9G3
/dVFeQKKrmJns90g82oDO8vStXIZHzZuv6ONNKFxKqLnSBA2r6NL0DsSW4sHgKRB8+t9Qi04NEwr
6JZc7Q5xdECJQ7Tl9dwsSd020d9spl80Rp1x9Wd4Zg/MYymV4uK+hTJOGc8MqVD+J10PeKBiayvI
7+LsgoGciA3vxylzgnHbUyhTuTUnMBK02d4gQkCd+MCpQNtbEtIYxWonsd+tJoPxMmTRWE/8IrJI
WcRIj/zRYzh5vj/DHz92p5qwSQDRR3OSVTiliIlUZbCO9XotSXjYttyWJHWT1MOBIujAPzLIN/wf
XIULVNpxZRLsdypT5yD3K3pnONUeMfJUIUtEDrg6Kl3O3pOBr99kru8A7fj0bEv6NGZICOqLK2mQ
+RjIvUW42xBNFE7r3L+u6diIO1NK1rhl1ClPoXrCgGa27GsuViuRUcPYpYtTtAU3uebOFtlPs7Nd
iqjxjps4oyUGx+GV3ZQyx1mx9h18TQFkl+3SkBjxbbZVle5LWWqtStQbT7F3njPPi/d+4oxy3a7O
9p40zX2+dIR9ZrST6/2cuPS7xO8N6sKb2oEYtWFgTW0pkrDq4GFygRj21QiZ78d4SLuFXm2R4GKR
3CngJDqiPqdrmeJGiYGkt3A/2ueHJQ/b3oQSWmlBTF+dA91DMxmXRaGkAIFHYN/zpZRPD4mMTxF5
m6G1tVBdzqqGFV5vCreJULZcrPmWXsaFf3DoR8uB1mU2tTP+6op5ZFpfYAGW0jsaE9Yy8HS60WVg
A08ts40O1123EZwesYVwpVjDDDYqazDwrV36GZ76NNyHJZAiYLqdOEBvOonmxalCieJ+3tI+IrRI
H8XxaOVnXDLUxSLrxwOnDfAOx/qzHbYhAm8iwPkEa/e3gBQE3o+1e4f/EZctw6AcXBR/IxAIN3Pd
1EBLSz+rsbmcecWaEF15kbvKq9zrosiJwwKQd5R0Bmk34ZerB1dc79+MB7yVZvrQuzYUs2huk434
LtJBLxIRjoBW7oHy/IQx8La7+S2D7fw2HsYSP4vlJZdXkN3audCGPgRF9EOcmeEtNdQ6KCeqSN+P
rffRnHcQOPJLJIFbVIFq3y3jZitYxcmSj8FUnKFBubW9i0ACEAV0W7qwi5OM1QSNtpd+TIrqH+Nf
itI+FdzDV46NOC5YOnphzXOD74Ahn1lca4D+OLKAnjnKfu9pyyr27MSmv73JlDujGMaBT7ZKq3cf
2NFrHesOIqpfVIvjP7OWblYV50fjA11qxODPqHk9/2LhW9CiXqmLwJNnf2licXfG4yRZ3/0lABcJ
qJZbVbYMxNY9DrsciohEHHuMzoNcdeUwHTcyY4yJa+NcB/6yJRT3KoagGLPeB8dNohH31ONRE7bc
sGljHKxujHXDPGiAbiAjnNY1hIW3/I2NfRVQbPjFVlK74kgoOvi0c6hRgZs+9y6i0+MB4M7tgyA3
nw2ZIVoyidUDekroV6uFX6JtyfykxzxF+C7OBD6fAljDN/rzLrfaoKh+xWTOaeHdqSbUk7btixZl
dZNG4oNv+BGnOc0qy8wkQyfzRth17rb6mW277sQzy99W0uT10KOVwdr4CkX6l4euVKpMHwLX8Xq6
R+T2oRSszAVZ3tZWrNAN3wI03eNnVw5hglKG9UCqxGOqfxW/LmfrHdY+qXl0oYT6BIyX3m8l1pqV
7PbeZjh8zRNqM7XRrpCRi1aZn1prqCs2wKcv8O2XL4+OekGqzapAYL8r6XmZlSg7MeHB/IMJyk4F
nl9RVifrdrQStbdM6BP90KgLDiS504f2A0MeXWjGPOBT9zjFmeXWs2tcpnsyu95EXQZr/Uuo7UUs
qatIwVTQiZ0DTTIOKoGA7Ux2A9e5qCcvNab+xANw1p/ReKy9V81I7ylXwke5Kvk13sa/eU81eyNU
ancPE4It6sIWYFU7CNTqt9FAVhoXvxGoeOqcXIHBLQI0lXYRc+PTGjWujcuxDNw5ZBxAdPepHktZ
hEQPUYB8j3dI2gaJcvgnJvB2/N05tuNJCAuzZBs3xwNjwIzdR38Qn8Uz21vAyOUoleXFnQi0GKWE
GsItwhu8i4MLMukRg+l3WyZuRVc7xHIArjtDKoeSzbVntn+5mBS2Upg6jMvVt+sLxbgTlsdL2N2y
t+kXWVM2j6JI4//1pQCfT38tki4E3xZHiMsaScmPEr/5UZFch5DUHIkZ4RrxYcgEarjkLXcrl3jW
Gf1YKjOhKpkt8lgJ8tyyKKJs3QZTYF8PJ9HPh60J4bHFQ6ARYHCjWYDa9tBTCoydqr7ybV1pnvQB
BtQ1zoBs4N6SKPMVK8zrAhn/UTNySBJ2/pDKGuLO6q2tV92hbO2+oE3YKo6NA7TlZw7Kw6q7JGVG
cu6fkZ8JXRXwK4yMzCxzHzYzetPGbZHJVgPr++1nH2gicOrfoD/+t9naQl91wLN3MbOWmCuydwW8
341UyhIDLey/b818X4rVdtkLy39cE8CXyxdFQnD1tyOpimueNEi9oCxkuSv2UzC9/AVZDzTq/xUt
BfsS+Mzf2pnhdFUHXggYB5zpkkPJQPOI1MOvhB+LxNohNGJpc9q6DWZ0L68Fka3BwTpWLvMkrO+9
LprJdlsaXIvgilvaI6t9GebN+sVRdEbGoHRZjb2MVXThWK9F0IvDmzW9pBkSoTuPbaJxn6pHQ6OX
82KUhBRt7sxpDuzfWs5HCxshUs1LK+5Cbr26eXISUpz21KE4rUODlbX9/yk7SxLw2nnMLAid5Dqh
EIUKud7PqgG6humO2XVWheC/XESpWH7fmQ6spOJnCiHmysYCZ3WZt6kHHlxJKgIez4qn0Z7FpyQ5
U9AbIFyHMnPGino7MijGUnCZPvffOZes/3/L4puhWeenTOGnLGJdAx5cr6rT3NY7EXJNQzi488C5
xmKHP94dGP3e/5QVfXktVNpgTNKxk0+cph7h4Lnjbrpm9g2SrpbkQOeN2MCDSHLhTprqLMjqs+9R
z/T+VeSR+81ZlKdtbSKmocBsvCI38Npq9nimqs1QhMf46b6xe1SLCXvZRotQaIxv0+36teVdbxGf
Mmba5lsZwvjEicHZGp4rYzQPKmV98UvweZVlXNIjceLIV/WylHJIrGUx85vV3hdb5e7vlMimf9M8
h8cXIFC5P9rSH8ulcjGYBlVqAUke9ulWZDiotylj4QEKXcTsaxzTI1Mi8YUSQpIxQOzyPKeJXvqq
JrXcpnmGBc1IxZrzgdP+iqnoqrFGSSVq0zlYhvdtKNrYVlX0cRDO3A1et84loTKm9zy8M92YDlLK
mW1ub8yV3fieOGidFpwZTq1swCaTCkw1YFmfbUPF3eoYBufUa8+k92Bex/fAieXJ10GM8FUrVExO
kXQyeIPtIhisYyKsB2ff06sBAtBDFfsFo9mMaZkfDQeIgBDUCljwRqJdW+2pOwhc9hZuTwAlj4+z
Gv5ZVY5R7NQpbcSZpEkFMtDzYV88auC9BKqKjlxoZOGpqU+pIUeJx8uGAhibQlqhmHHjuZBe131H
DBsOL59E5fx4vh7F4nrqY0pY5XHpodE6sczNKpiju5pT3slHqrwpQTJIjGWjGRbDaCTkcCcmJjJS
4Vrxr28uksdUrfoP03c2w44SCU42VjSePjD7hL4gJtWOD62IsBexLi/CsoGQSR08p6F77zkYDkQf
oue11GA75sALhTDQWkcTaXcsRO46J5P/JM2TCGy9vTwf3Iqmm1kCAeopj8fWrlxsUC5zZ72UXu1T
gG4EpOZWwctENMK04MNrZs3EGt15w+sgl/okVKXvXHRYaAKkOnrEwEQOBMUnY09Qjpl1xRWWbjue
wA89nd4/R6a5oWz8y1mysRu/7mvJ76XSD9bkFcRDS2VCv1LJGAXyhx3s3HBqztANd2Or7UFCrUek
pbBka16S6DJse+vG8BNTETfqcQmeMs8NH4VvScReZZcB3Z3dRFNai9faafENoYN3ptqHc/6CC1K6
6qEBwI7s5S0Y66nfMl94Z3B3uyL0B3N3+usWfvUwQ39wZTJlDO2qxmv0cF5ciUK8CSrdXxVgtk7S
rgXgw6CqHFYiXVxZCyQIcCrPVo7gZgA6VddZ/D6lkE1Mv2+ixCjFl3CZJuVBU6Zbkc6ZspzYv0Em
94rfkdIzD71ciEEp6bkgsumglNKM0ECx/iO7+HHeSIR2aTN9BREdA4CmMMz2r0T7/+laad6mgYTo
MRK/GGG8rKOMlEmq9Mqko+ul7i0ZwQDFfK1ke31fm0UbfMKfbYI0lanmiHv1LMOMJZD14YA7cl4s
yL8QFX6hGdVmvBw8agrnir2NSnXAVGoRzJT+jb6+e/a7YiaDGRz3z7PCB7EurF+ja+OQmqRUKV+X
0HxTvqZiWBlMThJtbaPS1udIeHMqoSQl1ydM5nfXZt1zl1vWhEuq/BNdR/uR43aZ5XeDdVuJcnux
n4LoxJY3d6p4d/jMJk7Ebf7vp+3DXyugnJ9LVl3lFtnFVxXS6dD5VgDZDASrvFebrdo1gsjvhRA8
Gsl91okHpogSyMjFUm5T80J9uqY3Jp/KHpcir8X4gzRsyMJO2Vm+dHPTXn0GFY64LRy0wSu1I/3Q
NeynidMlMUY+QP8pGi35EySdwkEWEh+8i+dcEEVhpGsJkaWyhLHnmC+kIjYfx6wRgsSsMd1PRJ7Z
vRmkCDJn0dofCmULN9qOgVpqVae/ibryUD0nM+G2KHLNa3awFfcJpkGZbChvHp8+u9ldtVBz+SVn
dBRVSU2ADtDGiMoDuQAZDsxtT4snacUuDwXntVQt0Ycupn12xudvprFghUW5aS3pEl+SU8bURJ6j
Vnn4by84592cSUpmggc/OKY8tXbqubitfM3aGswch1y2fOi+k7eGJekHzp1hj19eL+0zwQwH6qnw
7bhY/avOD548SihRcYkFov0ImhT5sZ0/ZW+oM415xHuBagtTbcrmROVgFBpNyAN6+go4ZvCqXiLg
P3b6MbwBRw49qNu0KrG9YRt03RTx1WT2TlcOKAvcZDTASd9eCTtyIEGwvohYWXHnoF4oivXKMuoS
Yq4L2F8bdgMRTYwpij/pkTWRZwMNrwf6SbgPZCtWF6OS/HUkwIqYFLrdhAlRaJNtR80D7it+894E
jZi5uLfuPkdwVQ0Y+OaZpYvv1GXQ2s5Npg7oP3fpUccEvovfP08MxKMOjdKGQ1u9XPc1w1QhcNkg
UopIyaAjABufyD/m5Sav139S9z62aAItNU/VwNN16/znKjVrMM91k8aawyI40N+0Faw5VnsxVl0T
s0TeyMBbAG1QalsUoK09muacHH0ywkn4TYOVCwTiPihdhA962W/phLPdyvMbQOfyInQSNaBeAZKF
GqddDqDTMQ3+IayvTcaxE2rmXaY8e99Htwq+BA+Z3kCFlOu20jKg+ruffwLXcsoxVBQ1gR1S0VFJ
x5PCbyBEp9lYAVwlDry6qM46+IuSVlcvl9z/vFd4BbXqUh94UK08CO+TB/mIOAbgwJriJ/ONyozQ
VxKC0Sv9RsGA0SfS6mOynJ8f9wylo8F8NQIryJNp74e1XuE9xzQTXUGnbgoUwFOQjjaI/Zco19Ig
MqmDPtyEexgi6LZH0SaHNlRmCMVZ4KeH/WEYtwF3uQf9vGsIAwu3l3sB9ULlPwTublCeZysDJ+uW
S9WZY6Jaw6Nfs62dFI1BCzpUaNn0V002urB1K0nbrpOx+w8rXNAag899PgwsiLVrJL4sufbtPoiX
MjGTkfy9kk/6n2XCpYFc8U0meJbK/7rmGoji3OFSyLznp5zlRv3JT8oVm8EGuBC9C6I5qB1Z+j4m
D8RY4/qvgvpA88eZFoUVypfwurJu1++9mkeE6HM3dQERqNHylN8TPgDEhOGNPo+WQzXl6c4DvORW
FwW1xKKsC7sMIlAdVkeFbPUYEMKcgboQLBawUUP8TE2Uksyf38n5UjVEJPKChdkRX3J08lG9bd74
4JXjp+aljqg6gOgRRgZvdb1gt/XSIexS5j9IxwPoCflL7uezL3FwGqaNrg9YLDTi7joruQv4CkBm
mQ6Vg/WjVqLENU+6zuMWHuSvCXw4kwlvivwXnbVoCzmfej5OryhOkLDPU/Di2/JEopuiqiFg9+ti
4Syh4Ise7fKSGUyiLaVhH1YjNoP3Eald8gfJSuESpig2P+IQbYZN0zKktDBvrH+Ofqslb7KrRLml
XCSDarsyKoHF9dZxIbe2JV3vGOJlRbn1hhJFh+DBMBo+xOdPHxypVie2r3OxDsVqez0htYIfVhSl
CgKe7DqMiYDGssLn8B7MIrITDFuiN5Z8jX1UBdxwLYapDUIm95Vy8Tl6rBpKhppbwGebbCifKVOz
MKjOwgfNkHxSCSOo/lRhXjZyjPBHMETUeBDonTS80jq2XSqa8DO4y6i2g7LzekGvf60EaHl3Y86J
TC8PXYfv1x4kEkW/DDyzD1NE1kHQGqB/EsIRnLzHlgUee0gYR1yEH3WMe0Eb20OWR4Zi73X7Rqia
8WLcu4lZr1NcM5Cr4EpMBwx2FSum1GpuijQjWX0h++3Pj1R0VhyAIrranlkxHBm+SFDaRyEvj0/K
ZHZcLipuF/T6wSN0s9fEsZKhYUh2Bd3bdDkPsjJvs6kaOqeGzSdIB4NJOUeIPwI/NF8Yr1vn4xVV
Gold4g+2xQGDEhPh6gzyBgi9AkxzL2sl+ZouPJPHg0EvUrDhtlTXblJnMFGl/T7ubcfpw27kLeWJ
NIJDbeJbESx4ZIXNExE0XEJ2L1EOGryVV92JHwrEIx/dKvakm9sml4kjZsHzjCe28DE4jkC33Pz6
O/5JC649/g3ZFwohbggWXFm3z6ocoHc6Szk5pzoKw/O6CYlqwkLTnXg/8zbprLzzGe/WsYn8G0y7
n1ngX3u/uNUBc+mKlmxvOvVhAaaFDkg1AH8VSD/j/zVbdGuaMESMqXiIuKZb1g9NKfpEc/qDyA7q
xXGT8xmlBAXyoe9LC+rVSxDK5RZ0gyO7ATEos0GoCINezVmm2koc50ptH+cxnMk16XgIU6Poh0eu
mN98O38Sw5UKlmAZeLmXeaQdAKxsMywKmizy75ppnzC1bi93Z1eOgGKzsJxQ9XcwjKOkLIkz2ldi
wj+jWtOT4gKO38nUakO8ApY2mTgP/SoB+WGRSw/MTgIhKBdqn3uWKN8T9olztyBWtg0CDggNKTHS
NUkHB2QYW2uNJO/WM5loKt5shVSiJtXaI7LNKEXA+fqlqcsbfOKozsPiG59mcCDwokkixEizmIkp
wCh39qAfZJi4HFMiU6s8o0sRp8abUce9VT4KrXQki9GIpg/RSn09337DavSN3Ym1qEp/W5Js9rJd
rmfTgiScCGnWIO8uP7PHsDgyH35G4X8pfHZHOf5p544dcOWfNJBcD4F94oMGtzx5ZwI0eDol47pP
u+MWZUZpiSF5N63Oze+enNqzaqe9ulAcS1eKZQ4HK6Ii6bLTaAtlg5FLwUNtcL12X6bdlNGYDm/k
6OmFYx+44WScEAoCvFuJ1dpmcIpGglRapl1ATOiqAHdTBQFzncyyAHq82lP4G7evFO99FNLjijrB
NPhBnG/CDWeB91QDQjOdzJTG13EgkWOGpUrFk4EQNBsWXjNprxRxB/+hGLkTSk3+Cldkx5BRK6W3
uwyKCtGMxp4iN/GlWCtssvlSaUSCSawDHs4j0tWVnaiYeJZtgSyMFMTS/H18yX6uartSpuQlb1s7
Vlv5YgOn7oQAcCk6Bw6g3L0kS2SRAidU3pZYgcqLcbc9jxlS4axKSAJKUh78MUNxXWfNY0y2Bo3f
QCG4oR0Vv7kl8wjshphaVEK6f4YMsRLh0vBfIqag7A+h7sjN00lcZ5JZ6JlHJUwfpFayVuHFlMYh
GXFRn6k/IykTCdCAtznm5QHfoWSndeLh6bkvkEu5pdiDgS0Nz2k0l4ZlZHsR/z3Siv4cDBTp5wkO
HLmAAng3LwGjflDa89VQRp8OFPLfwGHyI+gRx+6lXwvXENNwoaHKTgae48pldkKm+j5suX98kym1
+Y1y/7ZoxVBjzChxuF7oZvnoXLTXmQ8UxwanKGACbojBZW9f/dlSUNLkWaYJPoCxSl1je2vi291I
QZJjrAPxaGA7byTPvF9giY/qU1qt7jn8ZI4CdAwR54HNnKYZ1kb1gIbUjl36rTF8ztXh5GuUBUSh
WETfsTk5NBWpVDK2K6gEpzfH0/Zp2WFVFaPATnE+IGhguXCnvinHD17CHH1ofsAe95vRH9RKlcAH
sRtEeSBVvtkLZiwxPVojyILOdwk+2aguK5Zp+XZncO7Didkx+qJIs9l9InQMO1nAdVSsVBPu9HZk
SPKxg6OE/HfGUw8KweRilRuzGY4A9blv+TtmT33JZvPVBbrmRiBOZBVgl10aI7Z0oHIJW5++KYya
Czq7L+0wGBZ9hAjFr1O0530Yk9vKewixd59t/SO2CXIxWpwTfxfbtSGa71GYrvjuZyFSKfqMnXzZ
oM7BDDCuDdBW7KTApVD4BE9Yv7KPqlVOJIeQlLNikkqaqVYXNhE1LZp61jwsR8wSG9x/FmvAIoRs
slwT8Pl3OfpaBsQf2MUpeg+ZCstUbbtf0cdZueqJKAH5Dk2dyTpXkEAo1uSNvTR6zKhrnORmPBJR
SAHQitQTdJJE+wTrwkLVbarAbhQ5+7ocjbu8XIh6ZmRBitj6GE0Y0SORWu7pUkasLgsJYFhWMhQV
yypScdo+hcotSXlJKzys9cJoos69LxU/pkhZshEqaiDxWs+64llKZs8NSSZ2oVmuWgZLViZz4Bh1
t0pWXO6P7QvmHNV74kuZ5F+G3KaHVtQkuyC/oTYWaNcpnUTuXvyxDD1hiGMMW9ScZIJqSx27jdRj
9SLR8U+rkEis6oGUx2vXtgvHZy1QxAF2KoRkH53Z/ZZYpLwB7d9rGigdY4YenwDNAWicNCMN5u/D
5ZGQdQzxMpwEtT3RhiywtXt5etYRMA7HSsx2RAUQcNkbxTpHh0xBeyotSbDsDG5HMgsp/SeOhLdm
xLKULPsgxFKs6TfWMkwrPifjd7hDAqTC+C/sjx+CIk1FnPw1ZQFk24T06u9x1v8R1eJppRHLViG/
tVTio+YtAuP9/mDA1LfXwVNw3TqvkgZeeIbXVY2dMGEP8nfo7MCm3fe+sQxLkWuQfxVXDuH1EMBA
pWAQknPL+6mW4f1kngdfH+lvmZUEDeHZNIqBO3FHkkNbEyaMTGhVC/IxUiUElXMx6scZd/e2Oc2b
+eywOLER4LOGdDYJaVITyMRF0iX+ygPo6YbJc7ISYaH0TIdwPdWKP/7+z/vtOZFKg0/+ior+9ym5
7z1SV/k37dQ2e0RAIyUunlHjfkpfyUYMpr6TslZEBLJprJGcFzw6ZyBgVG4N2agnl+BXlU1GUthB
t2swxSckUdawaAlMXtPABYiOzdOtFoLg2Tvc4nch6TgyEyYBwOTRp/uNDK/OWYzJPnkCzK36J2Br
TN8VOiqrko8eJw9nIxgnmM+oww35lawwK6O6dC0gdo9cueIrNCqejGb1kOo06AEPz3VV5B3Jejjg
74DckL5LJ/GCHz6WXGDkl8hNrN8n/13m4WcYgaKWhzELj9mEax205IszpbtCtMKF3lZaojQWImaa
Amks/MOwK2+V7AZcjS2Vf81tZD4XrJ7cRXfvbH03ZAIPGvoQUD2zlnMxB3Hu3CEaIxMfyDV6oEzu
VI4IEvUrTGHvYYUFpXW4k8xvXW12MBQPZTUwaoR79Y+FrwzfCUl/BcPiXhtetmTjzLiBDGUi+MG0
QScpLqUbsL7NhQsz1D/n0qdyFxaCHPB+/6q/OBerQuc1jnx/FRaMQzdqUHWB/7om55k4h61fFm37
tWQyQUT0/7+NCAmGk1xyNMls8zgxpwxAG7YrODPEKnp3rLJl+8cLvPaAxvfst/7QWHQ7ZMdAtRwe
OZOufJFjp6CJfHqAzLmPERlhuGPCACMASaj3gJLtoV5nPENu+35nSWqLehFZQvnlaGRGQhtNYzNO
VFoiBuH2QsbtX1E7sjHh5c/mQqhCar8IGQtPRHi+SulRSRvz7mw+RTtstSmpnuW8qkUUEE9HglbL
8LgjTmtfNb56GLHNKiikDD6CEHNwZHiSD2ywWCdlCghIRPUXYobc6AyiuDjMjtcmFlSU29Z5AJW2
YjQifsI+E3ZjRpxOds+/pIolQ/hWo0i7+cctPd0fTiajiOtOL/rEYuSJ/Ik8V8SUMV1V3BQmDpx3
C0g8MT35eeABoqxe5uuRZ1bOwakoy3ci9+48XIdNZk3cIf3OjsT5FHN1NKGh4OoMTAPgS8hr/FCV
Odm2Js+HGmBwiiS5zTYXZ5WeI8C47Pmg0v3SH3WeN/NpHIXrYQPqfn0ye+dFl5F7vz4EPj7QJfhr
dY491HOLSDKQiLYZ1LGwTefyfBx1+cwxVSOxJrNuvXK2sGVFCb+C2QERoWN5ElJ7EA47MzRo3wzP
6H+9satBftQO4gy8B3YblWDdicsC8Y81XBpxjUMbVGsiShlh+EA4QS5QxnH6fcYC+Hzrlk9vCYUf
2w43/hUYq6wzK+1+4fGWPUOmaAC6rGFSlx16C/DOIgKlUJXmy3TdZasXDcIXq+4106dm6Bhmyccm
M6IbQjQQCaBxc5OjSI+hzvYJIfuPo+w8tbVi05ydkEdnYmEV56lDyLySSsz0hBn9G55CPus72HuQ
S0xyIseeBaJPZ+JeL7fGAn4Q1/g6LX1nP+J7FCg9L28mKb8NK+pJNDXd3GQf65mwlu4p/RzLM+BJ
SBE8leeWjiWKkqCz8O1QX57bCR/5b1YYXL85Fm+OYSSoJ3pXC3FPiyzLPuTqpXVSZdd+XbiCjTng
l5PVsXDMOwwOetnDoN1sTu7ROn802nJ2cEWNYssyIR8Qhb+Hu0nv/TZMctA+kJTAgz4eP72+8b85
FO+OhINAAtGYbkFMol43vLxnOLLYAqQmuD+GEdrcuDdRkdBQ703IGlNn87zpSs7hKlSIkFYfMwIW
XbTjXBrA+ILBBA0tQYvaawmtj0UtVpOjIMohsd77H88Z6Wj8lJjenJqSAp3Ha3Xa5ePGBcuF86gQ
P1Yaj4zQ4sR0uHlX1tPRB0PQvDAjc4X3dNQlN5nQ48iKG6zksSSN6FyEXcQ5oy4/kaIn3c6SVi7b
VNif7+PaJz/Al/LeHm2SKIFjTv6Ojtjbj+bz183rP64r2aK7IIpRKugbu9/0rdJqN+7KvKMAhV/A
AjDYRbh7trAKoCGHfwZOvLQW97Ca275HpuQMJ8jzlO8ulGMyv6A71FfMU5FBefOjCiPcnXtuGMQJ
bAMnKu+5SaVHlyK4HEqPY0fFkQCfPyw1X0uLS+LwEzYpQgLYdIm7+FbQWLiU8htWem0Z6J/4HYYz
JW5Ablw2hPTI7kiVxaeOfo0ISIU6Qe41NJmdO31oTPDwb6q4+cLNTQpC//SVXbXrnXBGkC5trWfk
8rvCnbtVGPzpaL//M21jPzfXvc3bzCUY9b+s9Yrt/gwb2LaIrpXhi3qGm7TiVqmjIz33acsB+8Kx
Nc/5xvn6I2j+gw6vim+EuxWOI9U1YBhVpXlS6ZNdDC0BY6VOih+ece1ugbQjKeVuRY7/hB6CuHzD
QSzwMZVMr4EgiAtFhzBlLGpZoen6lxjzDI6zot9435dSiym+TCSrhYeNnrEnlRBbwpX9m7CqESp/
vpMI7xiloqUH2ddjUrYG6XouhMHmwxF1M6agRA9F8q3mdc/WSwyVhvu2cqNk0YleGAfT1ItDpUK/
1yQajJs+uK2hSOywgO3oUN9R7GmadkBc47aOJpkq4kUslkNAELfYJAsyyPnck1kiMYVu2nO46lin
ZkBOVICRlFULIgfgAViVx8MqYDf5aigteRyzryKx9lJzRlnZuW2LiHIsEENugFmv0BCSX2+gYxih
dO7fVuRc7Xcv3ymXwNgt/tXFgmaqIz+Z87xTbQ3ErRDpNEptLGkgm2Oevx2BngHaW1vPu+iRKXlr
IRAz3YASg7UIou1Yj3W7dsGZVdLgCNM5+eAL9ZREkMHpZJ2pSdLN1qGnCqanEXcdAJagxyBrXeHT
zvYXrqyvMiSq0q1bqdNQBX8p+Efp8oLG6SFkxFFd3J+HXhIKQ1THMvQ/pmaj8DX9FwaPe/jZC0M4
dHr03x4LyKfqEo0d+BRmzqJWUHx2FB2Tq53/gFMRDaSCIDA3RfNPkw9BdY6M6O8pmmpPa+RDOYAz
wZmDO6Q2cJxYBd/DC3q23BvYRqCI6n7m1he4KrqyW9+qP4NffbZlkElc6qJLMOTrfmGF7ic4OUZX
v3mtUP0OoZanzFVwPdFcNvc7uEOSsRtHWjMcyDrqI00JJgoZ1rZrrRjI9Qi5WtSz8ZN2rK/BGVt7
F6DS88ZJopF+EVca5r0keMXJOkVHcv+3vkbxMB+nt9W/0KRbvNr2BQ0E7Kc/0YsZawCi7aIs6VX4
MOcnjMjpI/cWhkSYadlNgMQed2aLoD+inWrkq2EeSMmvizFoGftzfeu3ViRWX9aBsU4fUzNDp2Dh
RjO8brxZyq2YTDrh+b2fUD9rv0fj31mAzFxDQmpEqmHmsEAuqTOnI7T4cAQ/3X5TBJRPUIRTQHBA
RsaE2ZjHUuJkJfffW/c7YpkjOwMsl7tTr0+13ybahce+rAB0FMcRIevi2rsZXmkCz4iArM8DmqBJ
LjnpN0O++UHGcIkcNz+QPmDoZgBsVd6rVylJsYvlBCOhAEHAwV69ZliZQ8n9Y6qmLrH6a5JFF7Fp
4hiBAK2n9+fZICLSGDTOjuWNJ7wKZqxF6UC+74vBKL2UvirJ8NO7+9r4fOJwSOn9O/ai1gVq48Zm
E2lQTW4uH6bCGDt9Di7GIBnMi7h+jzEZDpkN4QVGPVMgA4YX+Ih4MBCEhRennz63f+DKjY7CtR5u
pEXS866Gllw474c1CzZ37J/N9zgKGQm9BnjZecYQjNU5k3BccGxqJ8+VbN3/qR1+dmOiAkP2mbjp
dfhxGTE6FzKrlI08Q9uWRwYPBY9BWTosJ36Lf4K/V8td8nBwvcLOHvDbhpdLj64x+HZX9ALX/gKw
JCgqoZL1kzSLGbuZky7OdTrIiPjkOuw/0Xr0s6PYs6InHJ0/CYCMDfwfXcbpKsiHVQPqNwPGb7+u
+qEDkhMVo+SUeDFKrKolWYTVCHTSvkiowz8KbIZiKKRkc9/TyEIX7yk+E1LmzjWTJFNPP1vTPz05
L3IAVULZ+Tg/9/mAG+5hFswzZOqdP2MIb175APZhAtsl6YJXAKkrEA8osIUDj+NeKKN5wp8mM07y
e+e/aXkJLITvuVqB6oDr7iF09UG7NPfVIU5bSoVH0eezf537osLe7JVuxo5IwwfUc6k3xq7wwGgC
45U4Jv9hZEQIRQDr1d6QhnDOEyFYlFCVOZmFBoNMdiHpTR6JOXKUemwCWYvzmxUsiRX/ogRyhlbK
o98mRCxDUXFpyUj6ikghZCITE3tsPHmgRZ06nZ8lDg0BsDub72Xc+5H6raGBxClhNgm5rq7dgeCN
CD93haXad8WSSUs9LxKVYjMOCSI91j0N8W/zodlIlTjhHrAeShUbdoLVRfwhf5F40oUhi1CLmPAi
a4y719VRsFbysGqVTTniqAQ8jEAtmo4fz30OeNphn6BM5npBwPXCaYVRc+F5n8O2f+Q8Kp4fvyhv
qo+ibXXqRG3l3Q1Q1EAuDoqJ87RWPbW9ANsWCOGGAjfQon4uQLHO2PZew1lBq0VrKlpFesMuaja7
uyKKO9G/uZ7d3YsPJHR9qpXwBlNk6oNRPP1weOQg1dLOIbcKHR906JI9bDNw0gm0xpdEHLndHvKf
WvRu3CMhOEOYFjyUCO7G+vfV3kplZ+fLEEO0+K5P8QRAo6utC+EARkRoUFyS+d0nizJ0+tjSqZi2
c5oP2QlpDg7WoJGaWAkg+pBMx+M2xdpDxZ8hPV2sxIEg1+gwAoauvcqnwvy6f5EsMk+Ee13AexK/
3pYtFo5lmkkVg8mN+wpBytBaG46p1JgXOV0VXDNu94MYLWRuWykFclhgslh0Kjj4yepgSOTnOB0J
0gd2lPEZpGCKIFi74/AInEKguK/uZ1wI0H+ZbIRIk60lM3fR+GkyXvrrSIGN/dKyC3eOLraEkqDL
nH7vZ3CmpfylUeLEhsGPj6tKR9Tbwn5ENsEpeAk9DAu/frMGs1NPu+JnUj0nngZRDEEXXajrX3mP
xQLJHEXAdof9IZ8j3pphrvLDxANQ0I/6AxtNS6khyAgrj9Ag7A+glTPf8NBEkg87PwuezXr2ey6O
KLwwuzKJWRnYyrqGdPvxi8fRhTgEoCQp/vi33BKVDB+XhkykRGkGG8parLu6JcW6LiPbWiO8ySPh
zIXH+ZM/vxBvjX+NRxPCSipYUMk2hGyqeCutFzF53s15T5E4PMPkgZo1/LjIO+v4umOpfevPk69b
mzjL5NTO5u+y4YrZCzJtHlW+TK/zjUoTrRvSEyvn7sxN7maKUYWINiq4qpow3JsSVN51JEHdbtF9
UuuX6CNWexZFgFP+bjv1zo3kzcGkPoapg3O6mNfzFoXx5r70GCevLPcEqvwmoCqWXczTuHFQ1Et6
zvf9ZLXCqmJYP+q1vmaQsNwOCpa0JuJmoHydXYO/TG2ixu7Xf/bSLYRnXqjl6G6gi582qPgPFt8z
ODx9zk5XthREQZ0TB4ckFzg+tTyKKgyCHeGXLOgTMiTK46tupIa1Ejc15AAdjG0MXdBfZObv1Dob
59FsczAW0SWNNNQHnsRz+YwL1DBcHkxQKJhmvhwSyLmBWStCVQdmOwKGKDar2l2izjFYC19PHLni
+iWxDmJ2A4ukmegYke6ObxADobgrOcx+ZiCfbj1nyAFSRIhmaNNVV3Y4geJ2NPlPd4FwwmgZKxTm
9SJYzv57in8TOmT7E0RG/YEKsSJ+G489exuz/uRawOLWQbuDQCTsOKCdXD4Q+SbUfeUyME10UW0m
ubF3hbnBRWH9D2en1DXEBQII43jb30SX4MA874icAzQErfXYaSHOEFq4t5trnmK+svVfj/u3zxmC
Bl1CusADJVgYlk2WpXghuOZf7e4t8FsqB0snzOtutr3ncuIepi1/i7heT2S5xSatIx+QCMDJJBhL
Ge/MI0sYQ879vAHZ9wvhHwooBFy+kkNnBkeOZg9QirBzg0+5XIxYW75sWlfFN7wNhHbcY8vgWxaI
x1OG44JD9PjZDrgCJlRHlnHw4IhQehYdG1inkUqlcIMcY3MjxHqLz6J1Z0WRc0S3yAnMjf/VuOrE
cGqh4la6tTpfdT38swxtcn5Q3RZax3S6sNz3RopH5SBcecirpW8uxfdws68HkGBz4Dd1lSKNQPUO
b5rAMtfSGyg7XrfrlIQVhXJxVpXUU4OSZAWvtFrJvKTshZeQXfQYYKrsP+BHCJkCu9jetdHVZDSz
xQPO7dtr45NAtnuQIfhTyqKce3zGJgj442DrZvjDqDFfzRGOdcebOAvGLFnVilJEezlcI/ujfQnw
z1VeTvjwfGInNzOa6+nfuzlPg+rtOxj167iX8G5U+lBdCLcfz8GhHG4rY8gs1nqH1flpaaxtQVXW
Zvj+FOS7YokPfArgebdikAVIRxPwjlME7cjqBI5MeClecDMMv0qifPodHYr4H8mnN0VxOHN5ynWi
e0pX/O1t1uOmXJeyjjAyLSFVGNWEfHP5UfvCPTMlN5b1zK2GRy913Zoie+28wGZe7nmoUWMjUWeK
IlJTm4kRPIfOV8mTh52R3WPDKZ1jhWVDFxxYjwiXOMk0LhWy0mw63c9A4aWNrG1SMZV5HrnJN/bV
Xh4Dl1nxV8DGJx99EMMF6NU0yQFoL7+GKCgMrSuge1vHhMUNwCqvBJteWn9y7fZWDbK1G7CoLUY5
RHZNYHayJ70L4Y8A55WL6reRWphfqOb5SoX8vGHZXp1hYEZUIGMoNmuV1xewvHUykmGP/yWN2Cqy
gT8KcG/3PiUoN5cturDVtRETYWwyrXud8AyVXGVd2nxLCeNT66bjIWfi+MrMicySsBa3Zn7hyoFb
yX5fpcy4AdV55qUq+dt0KSd5Fs3thZCSrUGVmGbyLBhm63Zxs+QIYLFmu8n2UTc9gh7zV/FbxoTf
rCfPc+LjKFrCO5acw+caKOGaRKZD6Oj9untcNi7T1pk8Z1O6XvuJFNiVPgWBHyY6GV2uXVED+gh/
VvfR5QvJSqYSYxBCO0JMMEzVptwwyDCiTeHMRHkgVul4NVtDMuS16zUiGEczETnZVpYbKdvavgtP
NI6wDPRbvJZP0LIXRYDHvkLZp7rHNj6782qYJVXHqwT3r79j6/EZ8nJipeMgxWjcYlKB2pQxYu3s
FtdJOkVb6UTZSk5mlH65vprm8wV6MPd65hRDgnA0aMTY5PzS66jYhS77IgFKo71ryI7FCrlslVoG
kD+fRkNliw+2vyhEeNuk+Gfq3h1yZGJtsL3vNgNwucC8LjdNMXuBsCv+TKx4gQsgkqan/fTbhVr1
whQ2KCFcol9hFHqvy8MoICbfe98l99VBIAiAH8o2u1xTB83N/fyEOCQvj5BHfxFP/l/8jkJXf9MF
oo1GOVrk/pxdLtaA1GpXEGmqneP0rzh4srZ94foVXL7jOJJ7yDccxVffEQP0n7uWtUHjPsnb5vwB
F2Ekq41iJ+Rdz5/1CmRjcgDzSwCF4Zbknk284Sa+7Hqac9I8i4G4Q33B1HWXJdPE96L0R85rcops
fCK8ITCn6fSBFS0o7NzN1vwv1qXgmsIMkuZL4b6U+0rxKlrksDGE8a7ZgHJ4Axglmi5IctBEOnT6
l3r+FJen5tgkERwA4YMpDe6AOhg7O46ptXEqoInvWRT0AlSe9CTRz3sdduTKEO/ISZlrHG7JesIk
TQH0vuTRo1cnnlnPk81qWbO9I+tAaw5sUi5p0UDxvh3DMkp0OoDD2hVTQ4xho0FvSl+bAu/s32fL
8//U3kM08QjLZDXCGwdgenBM7b+h9Y2xrNa7NIZ0HbPKs6HQ4zKjyV0KEm/GWz7k1HWKva5UThUc
P6DFb9JB7JXKW8Y/Z/qlcymH2BgyfAKWvhtzPMLZZyBaw7RJthroXhXiIzmWXqDE2/QxHkqw6QGk
DZ4qJIfrhGt4lWWOhN7J7rtKdaH4Lqe2m53V5JhwuHcYZBvDz6sI7Q+h3m0RlGB8ddU+QITjDx+F
qh568BXjJe7DDECsNyfv6Qut1aF2fA6UEjH/nEDJesoN15ZPGQUZUwzL1ecFV+FKmSjPbglWtAEb
gt7F/2USoytHhzoOi1FFL1FBzZHHevSG0OuYnR8wXSgrR+7+isHRe6qz8hmVZb7Wm1SSp9X4ZDXN
wp3BhpvIkuLeQNyIpoMgukhWAz9L2Evak+I0VrPTinXYZHYJcD9jd0hspMnaTK1PmRybUEWM4++K
Kor7pTkpJX93cqqbP6rCeLg2Fe7TCIrwupg8V5rIzQuZv2fnd+wW1il9tmzyYgNKwlN593weGm67
aB+1UB0l+gfCDK0fyIwDc/cKn4kHU4R1u6BNo7lfkJR65RkiQ5fgZIA4oF6c8mm9JXmtyh7kZyGh
CcgG+PEQ0v6hKBFNDanQgC5kC0y749PbktOSHknBwVGATX40TQbX4yg3E3Y4g3aMMNAKFykJ666e
1J7JfQmeI7gftysuYbsM2INgQYm+omyAWmXTelVT7hLHdeKBg/U4mFazhvW7mwXV9ClnahXRRInP
rSzKFlQJnULJj5jdf023Q4G1V3bT8HcF9hgWH1jFcb3WOqLjCJeBSlkXEwALM2FnxDdlNulJrWPR
vB5yzQAn/jxvfqvyGxDMdgCyryV1pa1vlllaxC2GFJlqIu5dQJyhpxvNvbI2tvAtzsLJ4B4ithJ7
eEFG1lWAeyP9b5DGdVibZ4aTxwSk8HRxxevIORk/aJTDJTSY9IoxlW2tkAkqsjlCvAMEYa6RNw4r
H/Nzo/FjSknqTCMIxpm498zV16fXaNspyWdCEEf1OGxy18YbQEfHhaKTY0Nw19UraRWLuRWgnyP2
CPlzdZ6Gm6mW7oo8agz3o5/Fd7SZ00qF7okxbtKjf0kEM641D54lTRDYjORo9XAYNkqeZ0gUTq9+
GuAZhNCSrGD4Ezk2JKpj0vlWzp1aTJbapIMbV26Hqi6taQNEYjIOfMpUb0S25n11NpRhsp/s7zHq
aO97Nn+QDk0eaMtySoFB20ych83N6UbVGOSsBX4OKHTQiAw51avxEeyTsPzcRaw/aoEBHMyJFqYh
mSkoXGuHWbGnHASTnaaKuGlXR6T99Pi55xgtyA3Lz9kb2NrzxqjbQ3yqM8oWXJ9M8c11txr9ZntA
K030Esuo7bJp/zpXQtmGXftltyWNDS6fm91ai1mTR8UqmigySxpMFVgurbjjFZqnJD7yph5are0z
ycyE+t1BW4/IyiiuYGLbAsPbwRSqMCa7hXozZXEu5RSC7LuZEe9kE97ljFA2HteTBU/9S3iqPO9v
9lGwXG2zfS18AMRtb24mOqu32fATvRPyfe6dZdo2ZH/waPj5z6p+cSB97ykVGULXLyULqEnNXDby
j3oAqAXH4KdJUYjd0dK0rHJnxCdMpYdmokh70Al0Tfepyov2E5s5kiDqZPuOEXGqpp5i2X827JTI
gKaRr20soZFKeaNUf/X6qjPlQUR5zrrMFGOsol51Crh5H6WfazCW8L7zIXfTgkUFMOE4XfUAyLcL
o6iEeWQadxPk06zVW1oh0tDYFAdUEdAUV1U1YKWc2te39XvoabwVPmgZe8a8CvOV67Wwaxw09OD2
WCKPHjFCVmM74om7+GzQSsblmimuB3goEi4KHAV9pqqYHbji1kJjUQN+xv3YagLWxU8/nxbaUpBZ
i1hhaImQiiBP3vtSjnuEQ7Ru0ToWneEdUsNW/4zkjZLbTzNYgdHIjkfzTy+FZWBSEWldcG6u7W++
yrjym4b6af981pShedHW/HwsEs7SEiVXB2AAOkqJf5fX0yq0IHv85Qcn/M1t5c/tzP2ym9DNhgic
fZapOxqNf3GQc/AHxDGwAXS9ymtdj694nfKLVm9s8VFdYy2T0PV/X8L2/AvT/ehtrYFo4ZRlM59E
MUL/2ZQ9I6psq9684aY+UpZAQzkLX/h9gNC2318/YJJS8GAEPEVH6z6PY69/TypMTgzYkJRREkMQ
bSS5rpcjiggN8kt93yjXMKrU1oPP4TEt9tJMKHDgPNv2VcCs8BMWRWT+N/nsRW04cVJSIM3EMeZh
eqSCVHZBRxLvnmy5bWMv9qVXEk6+AWs9jYoMnLAMEZfizGDLICdRdXZv6xv2D9pqZVEOPnJmov1g
380g53aOoxMuBikZLZAC5H+qUTABWXJiL9FkItUAQuknKpFkfD3VbW2exb0m/kNdNItKxeCxXIMT
YnvdHzQ4xHIFNEdCXSaw2yglRumybdS8OSgW78xVyKMCiXuIztu51cdW7ADAao+pL81UAO2A2Rxb
YJ2s2yAzl4Y+Dq+9mjNdVXFngU9RLJm2tqH0p4hr4Vqe2Gx72GsuyY6o/w+QGy67o5yMduCCzyYW
cip8wjfslceHUJn3F0l2BY5oLTQpvd1+sYSQmQMy/6+wvpvA5VxpY+r+uwf55mhm/KtJNYlvzCyj
Q7OjJ/2XlwA7IDWmT2bDqA/ac8TeppPNwoQ4QTGzSHvIDn1OLt5OsRPJZQiwiFb4UlB+5VEdl8pV
xOs10nnGfjdR8IGzRUixr2MlTbxBXC0XAm/EOZ3LaQ8yLD+DRTe4YJ7RiBU+93keo12zJmy2+z3D
nEg5hsoxxg4vvu7ZpEyKT/HpLleQeRZK6IeayvJgvwrqLLNL+UO4zCU/tUYd7BWObvgVoI3H1k38
YxwVYWfwcvEJTR43pQpYHAOZ6CuG4qOLCZYr3CYQYrY/BUw9CMJ2l3ucAYDdkl0A9z//UJ88uBu6
c3HtuJK709G7JvUHke2N3uZANyGFjQlyMNcjkZTz58LPq+DmkWUsMaya8z9UvVqu03ArgvYu5oIl
jLO8uTm7mBvEpnut3wEXEt1RHPaZDGhxbuibA/+3swm1gIZDVqDyulQPlhJLYwQqaFtSAni8IXWI
AGy28EZ2y/HhZ81hw/LwZlqG7sQh1T3sNsvIIzUHKKOCXVaMzsatC7J1d1xZiLDGtchdVL/VatK/
oDO0Zy/0lSA8k4Zze2zTYoCLIGwhcexSwguFgKoWrXL5ZuQFHLv4HiUPusjuJ4AAoVWGNM1NctOD
5OlX72WTgeztDACOwLm1DytukqF2ihrqrhDMRmphK0XovBPD0a93tdGngDiT4z8gnMHfXdgefBNp
AwUwZ30H4zz6848yzVanLf4iDOCZOTzMTo6nqARxORqDO1lTt6AXshk/+PmHKQm64vWEHtoY9Ver
mmR258oHKIDtT8GuNjEeptRSUVNOCHcttUMS8JTBhr7Bkk3VDwiftwrp1VwHEPbAroAILyr/LMSf
b/Z5xJY4iOMVgNGrXeVSotc5lJXXwvmW5N8zsmU0krtUG+8KCQtJsGs0qepo2paOsZJtAgER91Lk
CRWZ8BE+wKbslJ58j97wj2sDWUxVXz3GZozvLZPWkQeYhltW2UsxmZB1u/KCO1bsgMisR4Z7K8ln
R0lnoGu6xHkgwznMqUcZWNcp6zQMv9tjIUp5vV0LfPcIHle0TbDFIuOLTcu35Nr/ej41hLj4Nfwc
5Xsz/GdIZH6nHv0GWiqiyiMRFw49KxNHDD3sHwuFuDmPvPIWjDsqoHR9ik4FUv8/Z/p+WG/g1Fzv
2aoDfRJwbO8NBUlpFwXr5FTwGrLsPOgA0xEeKIMfkiHk5WeSFM87YmHK7cWg9Rr85Pp0FCO/pJJK
0gf5XGW/lFQaoP27Qv53g3TESpedgQ2mbgf4uuRVVuBoAJ8yOif7XFLY189c8V7iWdsrFITxO9aN
/w56ReuREwImqJl509eOySpO3imFJmRiS+qw+/k/cleLws8qtOQEQD+RG75iqtGga5CPq/uAx9fr
+I7/dZXB2/LZ55fRQwM5uN3OyUw/feGbuXxgZE+8BG9337CjxmCFDi27jRCWxdWeYBlA6NLia6nF
ZxWeu0r+EZCPonDDLzPLiPeP30dL32H2be69NceVtCl7DjH7oCCG/V0BUv2EdQygspxhFbs5tu8Q
TMeOlB2nVBT5TYQSf4Aug+Dk27byjwqgYVn8BGB8eKGfClx/fzrttDSWn3fOFeL9W9DaVv2H6bFP
Hzdr+4/bXtlsAhtqPh9CXYuCGK99ldZO1iSxeSv2eHEN2KNQDOmspjM5+54MsJ7LetAqr9t3uxuo
IOVCGvAdF+CyTzeiUhXpv9Wkla1SMCem1DKENfZfYUyTIjzC5eu98p91v7o1grmb+gmVUWCAunhw
TfMQWn1nmtMCS4qMQc6Tn/VUUznmk4IzFFE6j7Eu8zI97UG01OHb6DOtcSxFHls8YQARel7NlguY
uZ1UVnqOqOXFoymqnMPG6zAjYeJ2K5neqVjp8vvhYWQG0F+8RcTWTfQHamdwh4bAwdDR028M12PY
XvQ8OnwVAKbl0HiEdni9lZM33UToZn88xZSiWY7OfGW1RlO2njWVWWdFoSuCSFz6qxdR9R4H9D2g
av1qbUIjDMstTB1Ex4freXVlH3rLevc5Sk9CXfU+CQdmXMx7egbDmCYLeNVS4phACP+Y/LinfvME
k9ztUZ6LwsW6rB7qT38xxyLS6zeVDb7lHA1X14z5N2tHUB5RzAxgGGJMQVRziMtbjSSriVrbJKC8
bmTVIesFXwq+fAeGAzaTgmzoyarBVwclzC5Nd4tk+J1BBvN3V5mxJTJifDM+BqTrfAMiDnKMf/mt
ppjoqnYKA+fJIL9J/7gcITUOS93DUunUU6Vd3hEW6vN2HSkU4gjPu4BDz6mWxrlVwRzHb6sB/NBJ
NaVVdjZjegqdPjlkFe7KQHFCp5mar1IKg8kD/Qjnc5EHFtIzfHE1hbK7BWpJoeMLS4ZOzrRXdjfO
DPe9NZQLbZhCoIwdxbLqe00jQny7Ii1HwDm4/AO/4QVtybQkat9ji2JCfjeEMFzcCDzYYBuC3tOy
m+/UFutmt5WxmcYkv3+gK0AenLqbr1uNTo0cpmxXCovT05UKUWjtGbS0EiJZmBJ3gLe16ACxrXiu
O7lUUWsIbVqhtg2vCBieAgYbXru7mWdY4oYs841QfRwSZk4Fow2TcKJmG0EQPmGt7y2Wn1EQgLZh
wh4CjlduNbdZUdmCLf/tsV5V5cIJaQB0C0SiwO6wkXvSVbhEl4zYTZ13kTTuHFoXsr83dpYISLXy
82Gvy4n694WuLN7Jk/wcZALYOzqnUFpy5chS9A62JLWebZiIG0AhyZWXe5N11KR6uRvkBCkP67aT
XmAIbByTlG7Q8fYi7qWhEmOFILJ/ZuvEek0lp884ZnDQrbfV8YKzSIDkxtINb0ujnIHXacAyVegH
RcN0wC7/AIwNNFhsPdPhqPSCCjBmn510BT9dbP5jLPjSEWFq66/RwtEpfHncqiO8nFU1Dsa7x3VY
8g/lJ4+jqhPxaZHUhCAFk7WL/LsCDibjuJwB423kA38xmqG7eB0nooLUxn0jFBWtw3nrPe7pHnPV
NEevcS8phDllBCkHL1wFbNqsNEhihvoIHZSbA6IHXDTmjBg7T0MWCiVqDZC2S1HKATSw0VqFGtcF
n39nsJSbF53XdN4BB1A+qsc2c+6kWmnr4o7ax8LJOIJL8FWJcxbUy7cclh8O8n/+36HY1MUT6cjy
+zhfxLYCYjbPIfX69GA6zmJjjrmVjLKrJrwseqv46R10S6oDehKEoYdPZAWdGFdz1nd3dgch8e82
zi3sPt9IDkcPitRY1zSFi5U+7q1ZGSySs4x3wrGFljcJjS9gcaO3roiJkxa3JbebFWBdOnETK8+o
r6NcFBbmNaTzRGDHe5+LnGWZzhv6RuyGgl2ipid7h3RIFzOIE204V3EmsEagFloI9tCIE6BWswLI
PhKa0Gs2z/9RHukDOYSw7I0oUK/aNxIaZfGs7iPsVoHaTTjgFYw6o5ThKSf/6Mm7YvFpdohVd8v8
7aHLzYckicJXrQpiyJDSuDm0X98roIFns0SBB4P0UDsJHJGUd0Chtpokl/cQ0PUt1mvnEQVeoHZz
CpqR+yCmZlpi4LMyMOCMAWhN6nHG7gXh5W6M5E2jd3Y/Kmz6QPn8Oyf+pWqHp7gNubHUKjurpryc
YWb6P8s7UrXwAcAfOWG2t04WfLm7kR6tzejxoIGRbQiZwoD2wIAd/1DnoneZg12FFbxWAIE8pIwf
3aA0EaMfqhvMm+a1W+Y96VmhXNeZbvjs14Wu/tfWzEcVzHp1etzb6RlvHb8Ac/yeNGlxU2+H3CYq
qMNOGW8E/itTzzsbfQnbD66YDwji9gmliGax9avuhaqujthehejtLY8hPLUYD7EilUasQZtXmUem
c/qlJlzv+TzPPghCAzhZlPutAK8kM2PPNcEBJ3ATpKaqb2xLBgolV9wgeSMH57FuDsl2dKrRgd5n
fsfQ9JSaBHnNBep3/R9dfa8+uqPrhcWV7XUJT2euNkCjfNC8mjbSvB0Rfrvw6jg6LQfSqLI8QxcY
H1nQRwHPsWJMF7enuDe/nHnwoX2HXYYiKT6u06rUDgKYB3u96cT0QUEBnE24pFML0QwYPeBmdSGi
jnArwzGElmKUeLY3Xr1QXz8mUouXIaYzsayTJ1kfD8KJEnp2n5NDTi2slMtR9pJ5uJN9nrmSZm2+
TwiODeHit9KkCLha0DBmFFGW0M67QiU9BBD/z8wBbu7HSJZCdnd9UmVoUyRln5YvfJpYMOj1Qr4M
cgHVKFbS0DySGP1Vt/fyq46aeNuO8h53LH+yUS1v6Zni1LwWnu72pqlFUiyxm+2fkRr6WD3IIoWO
u+PLIMiJ0jTAqAfOuuWgsvNnxqPrCmzlHBQs4gaotjw6D5q3NUOLaTUwu4kcFN0wiHVgPAYFqPOB
ECp3Am4Ab8lKpwjQ4WpJX16ifxWYBJFoWCTgipW4WDnVPDwRjhngju/ClK+J2WifRn3TRFnJ/4lH
suQe1eG0RqALZaaoaZ2Zh6PjbBmgXuNj638sBTQgcUk/dUrzcSKGCTTiOV76O5mNtGePB12cMjnK
6DZdzEFAtVPYAvMLVmVMdR1znpwJe38U1bVzIvcLEGV8VI04Irf8ahF/fp5ko2+RETWAR22kCn63
m5ZRCqVkk7PvdJRbzVxG+hLcwDXSKELd0+1VbVRSI80QAENtDCPVhtDUvpRawyArZjha9jIOa4a7
yhLkAEAaB/nQaWoLLmgtA6Ihx4tAjRWcXzWVNNKZRZdr9hhLB8RBgsouseRGFADjjTMR640eUxpO
E3d8+NpL7lJJ8sQuGm7QUnf2gWv8GvlUcTmL76gn1xt9Ph2ZL7vUxH7yU53V+fiyuRAW4Aj7GohZ
kOYgRl2gJLuarFOnpLnlB1KF/RqUXi9E7jehPiT12xPFMHwbocZSKlemfULc8Y4ufALlZD6jCN3r
fCWjioorIvIhH1VMF/SsTcINmT+YRB20zFg+Zmyc7Wpfltf7mSsYKsIZubtgrTnaAurhvQOUhFPK
UZGfpGbUObtl1dLGVbAR67Uj2X756TsPPk87Y2cDanCgD/KldV75QxPSF1FL0qHrHLwg1WHJbHWA
UxvJKmwIwd3L8VKqkbVMaWe47LHfU2Kpv/MM/WtAE9wivc9i+Ejhbb9F6CK41PbkcABsY4JO6LSy
biSyvV/TrvZIXQhJRwBGRy4x72O/kdhEMnzDHZcIgjjGeMvRPuf22yqKxz5yAH/tRjID0R9p4LTw
kSfeN68yB98X3040p2mZrjQ7bGYUiIy1J4IojTyz7VbVmN8sC7b7k40cABIoo7h6pUS3jKVtRD+p
J/xRUw4CCug0G9uksoaCETZ1lpwivYyuDAc7w0zR0VT4Clo/0E4UmxPqC1zu902M2U9ditbOehpl
TJE3DE3+pYYwdYK+LTovqfxN2FmC++uX4FpyJc6FzIBRu3iHNn/yATfHOK4PUcLBqaQ1r3uBIjz/
PRN/LcNwUkw+hZX0jxtg+0RazfcSthsM0Afc+MRMLZZXZApba6Sd8anXlD6p13fbWEY6b1Ri++lM
pP82BDEy6akPJu0VjOB2y72FqF9QM0nTDVAz4WLaksr4VVL6mrQvRw+swZ2a3CvI/z+YLzKgkqHQ
PvTDO73ZyP3rrum0Y59WDo2DopTbw8kfbnqoVXg5FFS90z5jQlC4TsFfAe7kbmUSXAHa2tThmPiB
1vwQ112iydF6WA6/MghJmgd6FCVbsK7TD+oHCowc8uGtsSg9WVTu3c6vjBySZznoJv7tlMwwZpxO
b/xPRzFL26UX6/OI3EFHkSh932bZm16Ckwou6Lc++JFYcFzw/X+ord9CVmig1Pk39ZqLdDyIQB2M
R7kXCoDOhyHqWLogPHsYbLx0Om8w8PevyowEvnuaCupga/8voDT7CCxElS0aFKaYJgTKTE7fEDZ6
uJzxdDqAAkjy2bkBVIgUH1xtLNj4Pe6D0lliZogLPnG/VQ1DNkruCh89fLJ3WkWNOd2yRm7kpHxq
WHDGO4dXQGtrkJnRYx133XDzNcLzqjbJ+ciN6NYvPglZG8+q1ZG8vrFQlhdaJtSm+u/0YO+ZwsXn
LOT8tM8AgR/xcOLC15FBhswEtONkSFSNcJHDzfOnWjEvgt24Q2HMNyb6szLd0WGD6Sk2BU1MSPSZ
8Qy0HwUwaK/WFfZk0iGxaaYadV6j+s2Ghhd94rsFC5QZdYIyXA6b4G7n9jwEps+nWERxLmdgVqA0
RG5dKwlkwEUtaqXAktvZPfHXB36lbDAJyqH8mbTONW4adgEbBEG0IGISxuubIUtStTB26hJ2CfKZ
D8ywJzcTBN2Ud9bZbyJJs96tSiGkER+qEAmnWXLqWks+omXhzKRWZMw1ofxtPIsnimwK25QtBw89
mjq9JiUfBi9grQ5yBu/FTmimKYxfyjzvUORgeG59N9i2u79TSjfTLbNH/Hjjr3mxOvL8w/CoHRiU
D4Ah2jEjoyWKNl6/1nFZzrQxyp9mPk5FHryc58GPN96ezNkfxotg0M0oc54zrsiMofm0aD0dzVBG
obO/bYOHo+CHmuPcWInUlwwSXV/33wiSg+nm0XIEPwF00MqGG+xh6tuWy9vZehyx0F7XRzljfSTb
+I4mGsEt9D+1sAQZQChYwykoS6UsCfwzPaa2IIy49RmzQiTfxrDa2ynw3U2p69MzkTbpN2B4ohbl
H9MG/pW1l7/REp/3khH+BeAiWqCvxhuZ7TkhxrR95ZdV1k6f8tJOdytB/y/BuEC/F0yAdkaja0+t
S2IIDL+bu3z0ksfslwRIU0wqb3jGbFRBbzTDuj1KGVrLaGkCe1ghLX+3QrSk7CSrYt0ziw9YV+3/
khxqmi21AGP1Oyuoxy9e9rpREHjZQ9qv7ZXpJHXMQGlCfjxaeU81N3wJAusF5w71X0PSSilm1eam
J+WTGTCt4f8DAuRbtgaXRjfhPN0FGY3TV49KmRdO61fqoO0EgJb38glXEJLUSB6MuT9Q2FbigIIJ
lkl7ZKZ5qk3C1tOrU5vBQxF6aicJjh7ROmpjQHMWx/sl809fW0Q+FVzuYv0gVmOiVyGpRbwh+uFu
qJXApTolXAdNOs8JwxujiLExQVTlbdMVg3O/MhK0PQQ1cdIKTkQfRSEwu67qP6oyVqMAmc4FdeNY
4yNVM+LVGwQn1zBQuwTChR4eRZC8XqaShKLqnRkaKSPdPr0RzclkyULOhAS4kihaKhnIEJ1m/pVU
5DXsPZWD1dQHGAOSqz2MfgOZw7tlp4WkjtdboPtUR86xsXb9CtKtrvsPxIDoF4Umn/KzmBbUyHFy
8DLBluRRiCuDVmRZnWaKGdCoa1L7uK1BTms2evXnAG/7N+jZ9gdUewd1JYL7yRQa82Hcan6DHOc4
5HUwT0sG7DgeGnwZftyW54srUihlic2/Ub4EthSmSJLkxfDOofTryz2X0QnER4fhLwXjH/XjmJUW
1cMq+qHg2y8oOFSIZ9MNxcKpjSOzlmyXpNu6U7HKWDu+2uE99E//Z7DKSgpHVIt9mZUhCSN63H66
jWDfxdJsn/LEoegB+nsrMrWD/DQplFK10nZmw91vA3ZPSNUimpbsNDR8CUdYuTy+zS2Y+oM0saKN
E74q4hPanDyTcBHFOO9avg2zZlmS5MM9YxiUDNNgPTjROHQU1yoUSYCbBPhirek8cE5uxM4rXoUe
awjwx8hsd+Rcy5uAfM7Ixsf/e6a4JU1iRKtoUemA0DFJiw9WlawsOorPMJsgUPQ0qITK3xgM7GWL
ZSiyUtNgTX6F0MwRvrJByxsTF9rwcBS77jFtQJJnLxHbQDOze4AyjK61dIXrBWxjYW7mpk9vPRak
QTm4xaJaOQZstb3DmHHYIjivzcdmoqTA3zlRVM/i1brB+55TsOhLp+RoHWeIxsb2Dx0qZelpR6Nn
K++Ru3KAqA41IgahuTLlS6C8C7lqlnPQCyvOUbYCkjcvgEbWorMQa6tkQvLLYmer3rsAzOa/QAzB
VwsNAd1aDYCQGs3QC28MeufRi7I971Eu+zNWok+ygxMtF8JSQJ5Sc7oTFQFMvnCDhR+tIPjqiwQG
OBlf+K+Am0j3GHOqp+FuyxAIaq9PzSxjFrkDi3v1BHVKiBzv5PFzicwQ3pkMa1q6YQyhzdzU7kFA
aAd7yM/6UTzZy0dMdbNc1Hpl7RHIw1/jRMkJ9Gpw7hphw1zDAnwzds2m7INaOpHi5z27my5B4Esa
WAb8A4SoivcrxS0iuLfK1Q0jsDEK4T/QcBWN2961ghKFz9b1IjOZWHYhkfYe92i0b2s54LjU7LTQ
9K26g7jjLWVP9+fVLXkWBI8hZCh19rga0fMHIMW7nOYBiBxmzzHXF9KefEiwL7PU2Prv8WjZ1+zJ
vImjX5IeUqPzA4sFQ3wg8EmfCHVnXjZlHjH4aIbER3WrsOWUYYvgw8nhko4r0/yEzzZDdiXmvBu1
DTe8XXXYWU7NCsZVH4ZgpburajRNuYdiQKjaRVhmEpetCffiIM7J47RpObZ48OPT0mayB/KWRVMd
XI6ZbgN9VW/PjrjxITv8dktsa90qxEbeoxUCaH/dw9A9gtRg5jH9ilbroSjsLtvRJ0YcsCc1vjWw
doTjcQAZl4iz1dnxhUFU9dwHE6MBNJsfsQYoIuYXwTLxp3cVYkT+a+Zfn1rJLEcHBzP1nCQakAU2
FjHZOKpAotD8cSYqzSVbB7HmFpZDjc8q4kFMs/SqFYaWNNGKSXOgWm3t7KtaN76m4Jnwlgye8/3v
4/6/LrBcFPi6EBJul8+NYkFI1XX1z56ZZ0buIluAcVTe9GoNvQt7e+iUcRO16faGOubeIfHTUMrT
k4rBfe2c+pgbzYyMDI72hIrHkX/c6xZEjhEGqnIgHIqUOjJq17gh4MRfD7S3MwxuaiXok2mclIMM
TsVyUn6RuQJgIfAwoXeiuJwGfAAHYFu17cx6i/UAtuQjhZa3wC8e+lSIK7YG3BJ6C60YJiZLn9RH
u7H6GR3wTZYHJj7PpBOvsVq601ATSYnFTaTzHvtz+fdWoL62eyyOtqq5tOY5OPzfKBkH9SCypv0y
gyTdCaRsFIeqqRvlofPcQG8yjjPgQ5U4tJoMuc4ht4ejD5W4VWP3jxiRpwMSI78cnkEXhfs3k0TK
gB5+WPV3jIGRpkyKdNdqfhsCnxjBnEHRMzUtSWPwvR17XkoWkZx8MDXJ1OlUJsyv0c0D+TavXNy7
gnrV2Y9xpZQOSCv2Pe5aQdPNT3/7CJ0UG3VzcfLGaOH4VTH2X5dPYLZ+DdvMhxh2Hhw3mQXvHiCV
0FOj0x7lQ6i/7KSaoIMudXn+yMtKQcYh8/seqeqi5Ghab4UmlskBDL/mt3myXJYIK6srghecGnuR
iA+IpkKrmVKXxVhBdKeAu5rUTMURWMGJAQObNCU/V2vsWq7R2Zzx0EE1SO2w4gSXGI/AFBaKPZDC
wrkLhuTVDkY+d++sEwXOfabypzw3EPaB5vMVbUKdkjXACYxJNg2BiPaMcgcf08wEoXxVExSL1CRG
fdYb1jE/j8b4aDoPjdkeg0cPOb8QJ4Cw272N0HruBhe1Z8dRq+d9Snki449yfFFU17wcwTvlr/0s
+kvF7GtWjhcF0NHG4Za2vTkgqZ+kDN5gBP2e8TIcnVgaSbHWfmmnqKNLYIj/VW4o4xAryt5W3FDZ
MizQnohd1vg2Ly3OCpU/OhPd+536OEh2cIMLGmTkeWXfKDks7L5q08zRXFzwl4HRXmRIsPWjDJwg
lLxFiB0joUQivvkZsMeewUN47BwAoq96ziY/iCykc5f3N7jfX2yhZDJIacBhcEgMAENQHGgM93Ff
pc3N6sqY5KTsUG0csg+QL7OWQC35FSCHKiAkp0yglf41YdnkZdrwOKqFIG6C5G3K6bQpnd+JdjWO
WkbSncbUT8hqheICXAMxAVFP4X4UtdDIZUlWJa55+omJTZ0V6A0pt3MDlkLPMclPF6Et6hU+ODwz
AM6/hc/kadLAfLATVzzAOax6vVNqWuyQZSBKpka3iz8a86TYf08I+N8ZOxCIU9VtJEWeEQ3Ou8YA
GLIFMa4L04YMdaXxFHWLWj7fUxoYpV8QM0OnpUqsCgRgwg1Pgj+NwBSrg//EYlAYUxuGbVCh67vJ
iEhajEEv4zXT8T0XvbezSJENNK+n+jny+OJcRVm5WA/9Cg/JLCfi0UAG3DM4Ep26hUS9TeF86hB7
AkdF3UyFYoanZ99gP/UQVRbiDkZBbEsZbH/DEskx6SdxbVCaeI+FcsSTGImRFUdukn7ir4hg/yuT
+IEuuxNS5s7JYx9NHvyry1QYmlYoXemxkDWTFrgJqQcN5VmwazwqWN5BGxD8oWLsTmNhDz2xIRvb
jjOuvIxsOr3lVmFMQR3CQPrV+fwSGI6slKWTQ9PeMFSrY123mdiXkWyL07I5kwBZqBlRmJdALtuF
FD++x1JgUhCXDzCKMVc4GlWsdxQXYtJWlTzthJ73RReKFYq38HJmmNmcgG6iJI1S4auDTiaItGvq
D+b+CUOT4S2XNZy8fYkkP9LWzfcE+VdvDAXU/Ui5erQkPPFnpTbVny0RSYuUQctTb4geiN/krprP
Ucr99KeFV5CVRe9yvSYKMoymt2ae4r39uhGMtVv0WYBTb/PLwYAk9J6m8x8TQPI3uAssKdP/hnHj
VrdIKdocaRvrTnxNZKgg4YSrjZPhGso4Fmq+pOv1/aILUqw7votmBwcUd4pKtv5s5bU/HYQfuQ7U
JFelBkppIuHKPugylfwrN77N3T68CoBDm9t1ZXZXmVyFBBD7kOCF3ZBtRQQw0n5KuIGDd9NBrfnH
4UlU6x/Kw6RDTjCjyKQ3zcFcqO+2mhPIjrKWHNfycJqIyWhuELVXlOYinAoNMM9WwBJ4Uv3hpxKS
8zXr6wTXI0MdTxDb+xYgJtvW+//EQe/QgFwwmnjF3YwQbDW1Zw95YlSFEzcz3Se52dGfZ2uWdZU9
mxwWWXa77N7bzv31wlN1/WuEPYvDLplZ+1GAvStCCEFkYcBnNKhPRd6OzhYqkEjKUp+QW3zvq09T
gSxra/3TUcUdvb1nw4a6RLKaI3xGCtC6NgWZOQXbsSSNB97H2jVQM5nCLRqPAxFtYzdaNNi8Ch7c
pWg8xpGophpbzqPnLCdDaknL7K4knvzyYqPwmujmDq/gCJo9Fzkvz8PRHEk1fjWqeCdggDCs+pl5
WLwZZv3ZXPXSAt3KpQT+PWSNxtKCewnWuFgtqseRftc99cSMTI2nn0kOcLrmh7tWXBHhqan4G6UV
DEDa45rxbX35XVXhBWbAyqB6+GoI+wBp4z+Igf6Q6QifImjqBuGrVKx7OrmiREvOOFJej/DZTzTu
X1CCsolhEjc29RsNHkjsrJmDTbgztywM/BQnCd60RkXLpvs5E7N/qJ8ExB6P3s6OH5BWCtf7fzTA
IZGzqBHeNntevueR6iKKLP9/3np1++Xp+TtePUxYLFCa9WWwv9dWGw3ccSG/+KXwg58MNaU5i02i
qmik00pU4fu6volslMhmR41DTTGFkhFzJf9sshj7U9BXRqTNF7HgilvdPHg6SpmZfesHKz0j8yy1
Cd7ful+3TGdZSY7XOTAvwcHQ77j4UnvHljp6tT9OGrxz2GbMmtCFsX9ZnvK8t3fJGQaeWIyxsVL1
cryxqJ13+/MKmrHdGMlrl8qzV5z9IFb4EXS/1/8kuEhryuGGHtLHSIRINLwXyC2qlophpiWkoAey
WOGEbykabzi0Aelposv59zh0eDRzke9pqDZXBy7r6w36kVwlGDbN9mTzt/beM2fANaWY7zPbVvow
8hdWCv/ZCs5Kifg0KJlZPwDJzYpBj08SrvDlyzoSx+HOSIgzYX6rJu5BxO8pFd4a9wpysC+AJUeP
tEhUf3fcuBJDD61zxuBzmQF3AwqwYAMMrZvqob7QMbsIQH6Ag07OvJKxGtlCrB/WdSRav6QgyzBC
ketno7uZBq0mKq7ecvpchTaD04ePn6OjJtJlhfMlErD8FWdhv0IYJyCuQ+5VUuf3MChP2km2mTS4
nV8gJPPVwVMXqHWbPEKdpKHopAV1bJEsv8oeCvivbj1dAT8rl0EwNN9V5FATEX/fOFipX/Pn0nhx
QxD2XEhBt4f9T0RtcVN5xeUg+uG06HD6EOSaojlh2eMJir2FIJ5moXVenCtuUwF63xo/s1jcUN3K
afw+eLOroXV/c5zVA48PiqyWOVIxaFCcVGpkB3MyjgTj52scBg9Lys59jGoQa1dAf+ToT1KrYnQq
MDO1XtaiIQ64DtPlU0RZPwARmttKpiGb1IFTRrmxGSiO4N7I6YpoQplE87laflx5ezL7btnPbg01
kxjMAuwrD/+U4AHiO1WKQDp4Q4UxxtNy/smhBym4qQDo5qSwu2dXC+9irHOtPsegj156ChP5oBLp
19K2fn6CWpP7CfAOmp3lY9pxX7Ano6hZN07faF/xRrH6q6YKepSCwC0y2ztk32EypL1ABMyI64gv
dFa8yLbRYXOGUnLBwBYyuA3/2ifgwTlUYs64bki3fOCphhpFq5gCZ2mBrQ3fG4+AupKZdWdyDi9H
Iwu1OJFkAbmm+lMr34+Zw+oCMud30axl/Cb4H6rlFE0IYPqANxE6kQrZJFWwB1RFD3LecWGXPLsk
81ops1XVkQcRKkkqKMmXBL36kdu/73wlv5d+URUamVBJm2iCetkc5PDrrxdpwpj1ETHoryQRbNk3
2e7fUWicN5DOwlK5CcRIzoXUOqbb/TrEvf3r7kWHS4rOCHVYPGGc1naPgL22DBNNSY/6wUiTBWbj
YM8czPDMlcn+oNJJQP/PeSev8CWiow38pHYD+4qUZozopZUM+joH8p5DWX7MgAsgrWHtUGUj/hLN
/4nkWgvfmwuLhxnt4sdHlwgpAJw41qJUEjnEnCvr+dUowqSaViRnsP7Wdz+3rxuLZ3EJcFBMBpbq
oxHM+Y9r9u+gi/SM8gXW+gO1CToaprEUYSnv3J+4j7kbRwod1PMbTm2Ks4twAv6YYy1ntuOn0awJ
rHKBVRTRTXroYhxesvUg+C73KYSwOJ0e399EdNfxU0B8oLWnic/kN6DZe0rYPYNDX/4/Eme8BHSQ
yksEwJ0b2NuzEs1gPHu/iqmXFHpZOp5ZUsFHg4IvDxXdjDCjrp5bIKoEdRCtR4Ylghog9RMRneo9
L08dM6UpZKM9u2uH8K4Xk1k2/FnCQUeF587ElYQ3Ct3/i6qHA1EdYD6VXTGKa7/yGG4sgClN0hv6
IplCK4snD2BmB3ITtf0E54omU4FFnSn3zxbQieyVSSbjpkowhZyQlgQnJ7Z9Gr/8XFWpX9MXB6qX
XiNkM2aUAe3mbpXXrEDarr9nJunh6FMMVzenVAaZthZou0tpLBBXQsA25G3Sxz6/ShZzV8+nHxTj
1+mwDRbtbBRQdpGKpcHBoNshg89RxvnAuVgaejH6ZBXnrXSIequv28Eu3Cad8RNKSWpFP8vxsXia
DLh3/LHjJjz5q+FU4nfwgPVbwWHqYzUkI9FwatwNoRvD7ZdM1PLJ8uVPvwvTd1sIWwYcIcQkAsAd
u7wrW6XXVbisE7marP588+GwApYFTHtBqTUW32/cZgnU3YWL2IxoRw3uGGG78sWm45QFmSxNcWjN
i8b4vVLY0GNjfzE/Wmk0swMdvVN/J8AgKB6KfyemGIkmSz1FG1WH3VoNdasFUGDCaTzjBNj45aQj
8ILajCqwVLIPlbQqVc0B+k2tBjg4Lb0V5ROMp8L/AFl8/aN+fUlhBCibqqnyWZTBasxnR94POAfL
OxHPdJFD4ZsCUpXz1aBZZwFNeYowez4oSzfAaz6wqTmLTtNjFkxA/bZQ3manQm5Tx7bNsGiUwy4S
1hqDbu8zv8vjDPenD5aVuJyn2WyuGx5NioeeUz+9ADXAPvgFO8EMzMwIG4fokJeAGykDEsYk7K1A
BpcztvBPn2u3c/t0sKb9iBdFYKNEa8AjpFF/NMGaiEizmLYPJMR4O4746+gwc1cRAMOraYmM9Ner
iJSGiWYPtbmZyH5oE9jWNunbzipZsS6NFuvJHlOvo5TD0IcGp2I5biMKdip7WXCFSkkP4O8mO8dZ
GR++Kljd5D40hKfWGQ7jIZBTSyFvy+j0SKByq1FXvPb1eyTu89S/4hCtbzwW5iCZZBlhcUiwY1qd
FQ+MPMSKSUodMB0SlXY41xVfoIXHWTpjrwSk2MVy6X5kmPl1hrcndG0iJ4FK4bzp0d0jRizXdz9k
vTxXsSoFjKbR5scTV0kt55L0O2lKm9AFwnEh7G8DhSkeNazT4n2WfRuoNLug5z/yRMok5XbvMJrW
1E3Ev8O+Jzcn6tFnOrTT8ruR/YcMUyjKVQs8q5tyVC2S2s2x/SqqBI6/9Q57nvDprAqFtqgOtxTD
4KJMFSvBRmaCt426rPMbori13CeMw2fJNvvLQBvUAHvU2/NjWRNAqo0bM8CpNM9ZPQS4mpPi0LAz
kUMpox4KqVIq+rNpS4xTVZV34ok2Xn8108oK3RDMIxMnSbD6uEdlSpJ/o+nTx6flOzyvfZWVq1K1
tCSVSbUcQQrssa+IE2tQg/2Mee7/R8DaUpSy05pBekv9CBUNgxyX6B9RWidf6/2JCs6k/GE6Ermf
mnheV0H9Ew2SIwNo0k+8QqdENraZ9+R2Nn6LjdCCfJHjzkvh9F2n7ZyY7bL2ZUPZBGPTIYUGYGvm
O6xf+wnJwO3noByRfMa9aXldiIFPo6qwVc0pGcoyfD0GSyWi97wcm221/T5PorsBr5P+uejt2/jl
oaVDDYkWjWh3cF/qekEciJrygmaoMh/1c3qssjnijcpoLViGCAdoMd9Rn1Zx+d8tKj8ECXvzx3VQ
r0rf+7WpMFkQ7muolsK9UddPNaRhZKFvfsE8yqF2K0EQJxkBrpvGWqD36wn1iHqgXs+SN3Kh8fc0
6h1asjF9hpqNMN5YYgeDEyrOvUP4YA7vO9Vr2KvKGC9wbX2Zp6OOZSm7Qr+FsI38uteLzzYToUg4
c0fsk0E9C79hWJStsMLeGroq62hLpEjn+asm/taZb2FNxYivxO4nl+UIUnnIOQW7Fll4IUTh70ij
9d3iVgINYXEC2hMA0Ekmw9JrUmu3dWP5F9BrHepirYF7EVDUD47EpAKTz8AwzEA4PEqj5u7+fIYr
keCh8QAVCkAPo2u92yF7iNV0rkr2Mp7nDdqs3O1TTqQfUwLzz/jR3cHSEf4rpAwM/rYj8jWbHAJ1
ErU8nT+rmHvuS3SgrupZey17po2vWlLLeDxrUT+RmHhB2V7m376+DEjW7J+yooDVFlHJ/KTqzBQx
m7yv0oAg3b8jV2zNB3IarxPEP0adjUK+lbh4Tez4ONiDF3V1GtLaaDXCAaTvxwYiBTT2KKN4B6nL
jbvIznSalWUKIL+dkAbuL5a+/WbFJ2D/Roj+HVyElGIfk+5tVjZj5R8e5bBbjBAPgjEbn16BwCxj
wAGVKNuj72Z72npYierxMWxbsmISftSdSyHrgu7x8rKZyqJ3FYJfX0kN0+yfAEjlz52fHvmjT812
I+HOOAIBkxGTKuUwbC+TnDHMpuqt0e69BxcY5QZReg6z+27pcDIGg3HzknoacNse55wx7Sy9yQor
hXvu67wmxGWPNCZjl6MOE21Z47C0Fg+5qa9YvuTWUijBLB7p8iimfdT4x3ARaS9mtY7QTddDfr6h
Wx2a7Id1eiPHhZ/q+4ir/HHyiySdXvxXi4fyrzKQk5s+Eora0kjEKzr/M1GRjIUKY27TVFiPqUqa
NGygbTpxSWLtBuYltAd+Co5rhlXS//DlqZFX0LRq6+CLcq3GimvH3XPnLs5rWDlwT76IH2bhBRUS
IOGSn3gzY7llLkvb72nZ1DyAjIHjud59eo1w7/dJ7wG0atJY9DZJXvqN8EoQfKnhBUgvJrVM/8AQ
3QBUOiPHmT2gsI9awUsgBcwZ1slWc/khMlq9NpVMEfjcf7860fxkBiSy+vKmT0d+KmIDFm+jm71X
8CUn4BVQx+2fc+jzfObUCwCHEAfOOezooqvbq04MMKCo4GOOcU5jh/DSErJ7gsJgRotoYTI7wyq7
oPsaMnSsdCWr3LThkhdgmWUBupujzfCql0rT1CMrYnGSQes9LIv8ZEg08R6fPZHr7zSwNDSSiuWS
fP0hWeGS4aOd3rDlU3iQurfDqBYE63gUufbLmoByOUHYYIwlE3ANfh9UiUdM8J13vXMj6V+WPu9r
7LiCBjxzVX0Dcx7ceJxXyy9BpIyhJyAyvv5JXkLwipLFBKn6sU0QbNaMWdLqmGoUVRIioaqixhIP
YXBLibS4g2KyKy85B+ez+eTkuSBdnNjNhv3IYV0XIFWryW2vThKCcU37HgHeLEmMQJpHySEGvX/X
ARO1AjpCXFsRA18vv+8orEwxOsGBX6+o+BqSBXMXuybrByNewmrI3JZJXnHGtFnWf6mWIFUo0CsR
BoVBXi8vQnOBI88KUbciVUuBYM21hWCC0VHHAdy2SINytcY4D+QBPIdQd7Zt/oZYQYqwkh+7GbLr
t9eIVP/OwGmdnKrIV6XLex9O4UYD54WNdxEEFlEWBHR9H4SjmBmQxU6vlBsIjHVGIJZUp1s8LcDw
f6LhDVrgxZQw8WO2YY2Hze0VnVyOWB+tOQJAP9jE2PmQ0zvC9WPP883g1zVdS77i71+MeApqWTQd
FdJjXcUXelykCVyDsABLkF0BRWi+xu7xZGdkaSOQu6rB9x1Xirp8RvgzzNEl7yRMgfPUkNR1DXM4
k5yZMP4aMY4Q6LUfLiEHKWrfUt3Mi3sJi+izsSZjQMViyPHnrSg1Cbu1sr6oryxcWgbvukgYmoKB
etNWcYrBBk3i4juXl7mJZKZ8Hy6k0IOa3FFy6wJCRKLJfwdcGoHwMifWfKq1rt1JK+iL8GZbaJC5
/vm7eCI1sBox+CDgd8SBx8oFZ3XkU0c3+ec6Bn7SlyIrHpOy1dCrKqw96gmOpDF81ve0sNNYacMq
oxSsw8iEEO9k/EtrViU6z6dQNlUei4/y3iMyUUR1bNaXV8GZ0djKt5LzmGbcM9wtYp3g9RiJ2WD1
sPIZ1y6RLy/SgE9Qr3/ZaM0Ffcs0P2iL3QcdaTygVHutIg0O5e20akrq1zu7mb8NlvxQ5w+Gpq3t
NojW+jGcGgzseSVldhjYbV68Exy2KSrZ1qK53ZEqu5aBTBdzSmK7o/jeAf3mtSKWn1rwM50V44zN
PUf4aHTojeZlNW9u9gYXKA4vW9hbr2H9GaMo1rioJNyWZJjDQWIjNAVNInNaPxuCRsACzJOKSvSi
fRK9vQoSYrbeRfd2q2iIo50M8+oPHqkeQbHqC5psX2esLc+hRDquVIZEVQkZFN6fG40seSABbaIn
4qCNHpzvaFY0f/ZleEx5120moCZtz7u6SkDQ9zpBztGfaYTn57ffqo3ImOzDr2gX042oFzcd6O/4
Yv7M/lp7/tEppCifRk5OBsR7stx1W1UZlFzkLJP1Z8hSc/mAuNj+wd1EzEr0Fw5kaNQQze5lSbom
YAS92E2B2EsbZxM/0Tm90poHqVadQMkoEZ3mYXUiUWkPBkFiTHcmJfzRWc23p+0FOw6R2sQDZXA/
xcmHWu8rnpZXuCDgGBObNkL96nX3Q4RxPhKP/IjKTDlim6AQNkzI24DMW17hITlYwIVOaVeilc2B
wRRJeO/U2Fwy+GAVRek5JHOIURp23BF579vRKTVWcNhvQBFM2K75d2YBZjZFduoX3fL0jycGJOLs
ZS0kh6m9ZSHt+/xrW6yNjKGtO0suNdBWR2cwiT8kkUJTPBwBvM2ixCD5o6Upf8f0glLR6zAVbevQ
dPHXuUS1aYRA57bhwWNqJIpaXCv13aczVma6wCP00K/6QhSFbNYaDVwM9vDs8RR4+DKuRArgeLQs
sQ4ZEC3tekVMIp1Hi9aetFUyK4y2fz6KqnvX//qDrioJ+i+h0S6sboFJW5qPS3Vjg42PSHGzDj8l
sXFdyfvXnJGuInyEZ8Ol726B2QDdIBBbDsUlFpIoXxPBFfnIXAlkZPyMK2YBAsrb+c6QqjSA4+Bi
7LLxQz3QYxE+J65LgYDSQ9MQm2i6sypA0QlYL1/JW5xssu2GGHHKee8lgUtMGqjj+sr2yPXWha2n
3X6HgU5+p1fLpLPswD5H+rJxyDOisQoz5E+RYstnxUGz43eUT6bi6SM7v2ODTCNoxqV7oTYUdxmv
QQ/uMU+bcZzXXQAnH2/Zh39VOjYLHsHP0aeG82js/ut58F6V3kbF8DffUkOHTlkTnNenY8i5hoUR
wSskwBZW0fDEQtsYc2lKvEmLMMafdjUud6GMo6MMn27F02YFUXL8KAQ7rcEU9LHy/XbgcIaPYMyA
gShmrEh73iFi9VWkk3+1smQ8fPeUd8hPnSe66kAb7qTyCoIXgGgSNwOF+fMnXOEoc4g8KbfH04vc
rzLSajFtj4Z9+r2DQ+6GW9ek/5rmAaLy9kQm1DMjtTj+lYs1G7cMJh00GxbQ1Y3nUNVLpTfubmQ9
MjUhqID5FOHlC+juKj7HRmsaM06wRaHKUji6MsPfqNlYfEH4Q081h8FOSj3Pe3uBJI1K6PiMqv0S
ejcnY0hAj1ghf2dvyrZP5w78pn6Sq0rvFIS+FeBCqIIADc5om9CF89qHeHxhr9Pb468WaFWjdcLa
TF+JKzVyMOr/HuLxi4ucBbSjwbvf6DCppzBdqMzRNmxDFtzIfXNPEgaHGVeglSn4dpYqk3dDOwIf
kNdbzH/r66QYrKwoobr7076qVB2wcABrIOJj192nIbIfTKVjEJ9I/jFBBgQzJHbsHH/1zGqfA7nY
y7rs6l5pNUVpP7SbrUrHV6GCaoxqRemaHFy5Ji5Ry8m9nRuPZwi98idZlcjo07WWL5oFDRY9XAus
tF5ly2vBDXnlVHdTy7IiuXKFfbqUtGy1DutB7828CkcQH7co1TnSX7OCtSOUG0WKbd3N11khh1NY
0G2s2u3EyeqlSfxSwqpEiN+Am3276FoOERVFFFG7CXF3FHG33SS0sTnpOrDUga9+6F4QFIDbpAQ0
YaWep349phl/bCgErrWoepu91FV/OPqTt2FOQma8uUVRzgv+6+a2s+z+Nc/lMK3ceYhJgpr7hAJv
B/zwjixaFlW4OAe9cZeiTHNKfXlj1YHAyAYU9ShWPrGOVG3QIcXtZ78wCTzxbm4H+4EjVZSt+x/s
pfbQC64JfQNSZgZOUDzyEn1cy7RBhv5vt5v+gCzHu+HpcBcBkHod56wDvDA8K9Vd7XfTeun/dBs0
xo4sLi8Tdz3pNwm53h+mMLTKXyII+93kfZu5dksDQPxKTPClg/25ctyHnpY1mdyqPBJ/OjXSwO7X
210qJfedNkGXbdGg8DorAn1Rqh4fN8UCSR5jJKsK6N9r3MZdjdNSAExEGXDcBiD1hx25JKHQ1D24
pftPMLp89X9yt8SB7DpZ6499Rcl1wb1FzGd4dyUIkM/uMaov79hslI+rmVwu/UzwGLeIA325NdpG
GdsjlIxJKVsbaV4k/r+zoO0qk5KO9sXrVP+P5lLRub7EuvcgVGZWvVTlefaIWgDtqvH/b836lKGf
gcHpgJVV+pdaMwJURoR3RyfyzkHR2dO6WMmKErE0KqJPVSVSzwPuSqH9uyV07nPMf6H84Ve1CHqZ
A7HM382I5QDXOpF5cwrMc2WKf1YM4K83+PxrnCu/noY7A1R3fVRkDqFR3MdoqdhmgAh6hQuHBLca
TCv58/Qlwhm8cpigsL8vw7v/5t2U7oFH0LtKJNN3nXoHYHNBD6UbuqALyc5tbFeHcM/aRyyXNq0G
4C938DZphzro4ZPTz3aVxTZdaMwXZNzfZBjmPeZRBIdVeRcO6NK4AveKJwGp7J8OY5setHN+wXlX
m8GV7QGe40+LHZ5WuGhzjS3vFr4JrNtW1zuXr5WqyqBRqK/BSVQvHQL9jN1HZ5CgbMZ7UlsRb2nH
T7g1oAJjt+tc+hMpBkxyJulkm7ZGhz225QMevfV7nJVQcBIIHozhZoMWpFn1eiIk7ZN6SWO+6t+d
LP9BJ8PtgmxAWxljzTo9QVYLoU2r8qQGbw6zKyNfQX2siyCzaJ6BZtV9/vmxMrK0CWnMPVMQB3lo
L/eUCSQiFfCr9MQNR6rr+JFAWjf0PhMSL/8znC/DApbpp9oxaEfaJ9up6tvYitD+izAYRL+8wzR8
a/LhnMuzXZ2wfEF+wQ7qogHhqjMVAsQFgJmYyGYLPLWBkErLgRCNunyDabWs0i7jQDXUYzKYawW+
TdQeBEboCUz2CDa4sCDS7l1Rz9Wx6KBp3HgD9+gJO7FcOQ3K2LuHBtY2z8Nmi8yE5ofJ4D70ntiC
3+wlSShRoutdUtoZZ0/GXohaL6kuNapohRWtVU691WeeQjNxUQBJ75XAk7/TCpMLmhnFIDeC0HG1
D4s+/6UjL4Z4GuwckCu7GeR5PW1gwyC0HzI5jDKDJFdS5s2WLRvsTPUmEqc730vahYOr8lbaUYbZ
pebDwKnk8bElRq73//wXE0GtECDNgCHCntbxtUHGrKMB3/tTwj8KxqRtBHam/1Usn7EnFV3rw0tl
SMS8J4+zfe7gy5YqWVDtKRL8jMgcgPAC/Arefqc8rJH3Wym1HeSLGh+wTnide0T31nUFsSw/HCD1
cx6+86Z79ozGpxF8h20ZNEgKxc53QyHx/nGOdpfZjOpG37dOsm10o9W7BL4gootrqz1m0cMENZPb
y1Y/OgAdqil01I8d+gLmQqEGJTQfm3mqhOuvqzMLBC9srcHuyOnJZpxff1wWtwFo/GRRYHFd6ifQ
JEne1lVUXIE+4DWEOM0qfFf1Id8+M9vdGKwj8M02pNQ7dikFE6K+lWCL2qeU/HoA3/VjRQ1Zb4vG
jxp/XFfWSnqpU8DECVgu6/MkFG8np1C15JhpKXwb5wG6RRwU5JqbbfKYej50200xiKuiLZB8M1Zd
mu7nVJ3vi8zCAKeYYsVryEOhojqBFsorl5/Gcd7xzVy8efKyNoyg8+AwOgkc+x6NCImwZNMNZ2W0
Mj1BlHsIZZWC00qsKGJU4NtiWGHLmmWZA36k2CNOwnoiOy8kbX8yaPGE7R8MRDcTMQ/9+CfHIL6R
Sh3Sgbuc5hlXfpg3q8iqQzzazs1yAnNCKdPhD1ErYUmqRy9e9Ksnn2JLcK/D8uZYownwFXfKLdib
4XMyIjqEaj2WOlFZEez3uxRqTFSeKcAIaNdl4vZSZV5hIhXFNgJb9zpGSYgSffXJBcqSTmRs+flq
S+hJYwLTjDPMwfFxnLsT9Zsn2WnKEfS/ZrgQML7Hx7M8t12fGs9XXn1P0gRaPAx0a/guF+aFccMK
1WWz3XEECj+vL1bYq37IaLPX8ar1/8S5aFYRN6gbLenBXIGFZdQae2LxGZ6vOmuvdr43dpAzD0Bz
x2kPIImNav4GZ0CSf4Tv+bP1FANUVvyZdkSat6atsIqRN0A5eoc69K8WeOEvqtcq8TzPBFxJGWyQ
6tPknz2HLxiVKFdMwhzN9ucXkEkd0WdT0K9+QrgadAFPim+FCOVgW2R3wu2fXB0Zg1LUEzQvQbX4
l2BHpYmb4huqqlJFwLXVjBTj/G5mauFsCrPT/5jGaoiRiUZsMxmEngDpHqgw7ue5Cu2+4XoTtifz
tPoX2nynzYhR4YNPkKOAWtgWb1swpTCkkRn7wpq9+c0617UFY2mfODAY50xjM+PvPQ3uszN+96FV
pcBBjbRtbCMUWapP6b2+RQT9/KuwffhsLcDZEtUzo4jmuI8Q2eiQMj+IfaBKrmGLU/4RqHBjsGR6
JRrv/0hpuIebCeqRk6SkeStwZR7jHvDK4StahWxn2XdaYszI9ddAYXdG528nCY0LPrHp744gpPR3
ZQQHB6xOhqBZ1dKbcigvvWRWHamueP3btOCD9RpwJActfJvDjf4Jj3hKXICfWson85+0Go3cU22Z
PXY8PRYf90Nk137ykF5eEFRLiDDFGTzhOoiDH2jBrwwkI8Kjk9ymmbWLY0YImfcBSqM7a6t5QURl
+/iGfqrdG4QETaUTezow8oajXARSfMP8Rprjnh8AAx1JEGyHWjjmhevMZP2navW/0j4OYbkalodm
rekrcxmkAiFozIB8cXHb8EhkgU5Hfonv41e/kFcrf4YxoQlWYWZ8cP70zCpPqa55hO/YOaA87T+o
iabJjwmYtqfzaVsS5cjaN45+foLnPqbhcBH5rC7F+fgG8DqxgpQ5rrE3zdhk8X0uV8J4+46Dazs4
AuRFh2RxgNXBavbWojHOrUJiZ/Aq9jaLI3DZPUeTeKr1r2emQk+338JAP/i7mcWNYtA206BpRdO5
G9R5l8c3MWxMkrF8c6180ofzum04PZ6czTYnRAReVMwB0K02x0YihfidlYOAg84KQkuZylg0OhAO
+QynOY59083tMvOaxHqxOsj2SWX5gFokPZRdLh+vja9SFCIC8psfcHMgEIWnI/qR/sd6Oi/4W4IZ
rWKbLO2Kr07ruxbgXLi5Msc4ZpnCyi9HgrZ0fxKhEmkg3nYIjY/Xyd8HG7/hI7p0qncbmb8Lixpc
E7qD+t+P9mVGU5zkuk9Rq1Q1HzEcRWrxON1IntTb8pb0yZPgzALwDegv+u8SZW6oDQ3RC1xQvLFD
PWSJYUzE6lTxJ1TvdF6vN9NohoLcJfKRzqLxU8ADGRDEBaj76v4IEK5Eql4AsH1qJVjIrBKmDpk7
hGKTnYQRJmF3RstaTpAIAjSSQm6GuLmCt5TlP96L0Tm6oskhkKyabCkC4EVi8+Qt3fDbtcDRI4DS
uE8CNst9hyJgt2RjMdY4HZQtdmNfXq21GneVFsWPKuaJ0gaVzn6psCKqKzE7vyQxsWf3EMmsvg8R
s5ZqW/EUQFM4AlJB4nRyQ9GbMuXFJGQ11vWIObQBiC6BUzgmKwjPG0Te4fCpch4+NmYyXgp8oBib
L1h/AFQLT8q9AiA/jUARYoLRjAKOKK0Ic7zqp2f7u6cof6rJ8R3uHfUF4F4tzWj7ckyP/Z3yzMhl
lke1WYOsKwcjVRsSQV1xmT179wsSgwrFlSRCTHt1at1m9WHAbAEOOFsIy5ROI151d7uX5CdNJFbO
P/6OE+NRC8AGpsJ7nx9mCyXsx71HOb5CA1LWECW+E3YhpOC0pfTnj54oITQptvLgA9tr3tA8dlQP
rIuJRdzo0ffreNAqZbKKm44Sts2j+RoHzESf8e/ZK+p1nStxuyF2XGWG5rZMXr1RLfClwodGT2TK
N8IukeOY8Shpq92+nGqtDYLPKOGp6KX/3nHDro12YJ8+HM9lQK6mx2OhUifiCQs2nMyscbqiQ1Ak
OC4S+L+o+WVs4hvBN/950yZv6wPvEVsniupNL116PY3T+koVYvqbpnegvffjlwW6HMIMWEYYoXgw
Or51mfZWezAL8fqOPp9uAdgwSyKjPYx42c3v/qiTjTmDHHxMM6gPMI0gIdVKNn945OXu/d3UCpzK
881an/9pWkdE/TJwp3Tq9uMNHLxaWlXYXiOruuPF0bD3wpR7sBCowcL5m+3R8mJLDeXm00gHv8q0
WaTrlMcmASAlwop6waoMmTSzH9uq/zD2U4m7EHWG2EG7lsv95/9fAv+StvRR+v/Wg4LjExn/w/Lm
lWVaH/Z7OOSE5YqfjD2dXYIOb5NdW29uv6dDsjojK9aGFr417V1K2BJ7dc8OlfTq2ugmyyloY0Me
UHgAFHTSEDx4OZM9WrXI6X5sW7jeBv9dmImwnMMTgJaRTTvT9jU2DEk1bnchjJtYIJxMKpeif/yc
gFXDrweXQSHAjRxlDxhJwGsSuJkOU4vBkMEcogLAHCqbbajc64wV4Psqdq5Z6P60VhES0mSG0btW
0JRHsqlfziZifYoPVPP5Ug/CadnKB6hOnWFgqxosvMJImpnHSUo9fkJ2SXttWkUHdd5dXPbxjWRa
KP/u+Kp/RA4qMlwAXIo47uU6IVS1PtUNI3zyGmZQfbMY//+9N5WxR0xpAYHXoPF1mQPtD1f+oR6P
ICGWQ/hKP3zfKhomoy754tkA9McFCl+hrWFiOf1AzSA+NXxUutWHjNm853V52oQFaspJje1WeaSU
boO/AFpzHXmwkKsqZzj95IFqa+8gfWOND3fXnIem4FnrcGHBnRJmG/hRscfVbRbxUc2djVp8Ev5W
umXQIGaAr0WoEa3yLSVQ9KzoIt7+oZoXsB4J1UZxzoNHTKJ7OyD4bLq0jmc77DQ1t1tBGmGlmC5T
hiGm9tejKGaCgBGyPHc4wB0a0QHu9vWA9Q13zbdGMZQtujqi+8gjFIPZf5edjulBGbvlx+CPqSwV
icnrjjqURjXrxQLy7G7s5BS0S4odwfy77s0deM9dDes6J/DsSX3U71yOwOdYMh5rI0UQvxOgYzCw
T9GpsAkPhxtcN6xcbo9aBXx4lApmYFcWtBkyWvui0sPPsg6Gk9cfWMnTlXICWW0vJg9EByuQboqm
eetPFmFoIc27T2wOZGtgytizv6JwYrY/P2Zw0DZp+DcLcWLnvrqGtUQlURcu8IpxxMBKqxh0fCta
5eTWBedLMWLvnAWz1fzNS1ptpxjb/wTECJYl4FFUzdSbnJQllZB8oRqaAunKZ65XHsF72DtBPlIl
tqAAFFLVDzwMqEo2eJm4ICMLapaF2IlomYmItKBmYua1Et3vKwB6szLlHkJX37KvS/BJO5T4Lbjq
i+eUof71e40GN4Ii3kWqn6KQUscu3K9+0nyYG+Bi87fYNXHRFMAFDSDGxTDv3SM4Mgy4qeSnHqvJ
I1dQXC1gHD50xT7H9dA6r4LUogJsjWHfq3qdlE+tTty/430CMGDWVyuuKemEFvCLNq0LDVz63UNP
swd5ME/qAhjQQJG2sUNSsq0pVhAhrCHoN4P1e2bO0uuk3cFrUVOYaOZByvZ1FUH2GRYVAEXhqWPc
wkFz9SQpWbSFFXwhtB4s8mjd25ZgFFfBlzUHUS4yUS7vjV93ryCJeBkBrNc71uLykodbsRnUqVga
h4VtS+Ij/hQJqW95AmPtpUmc35YktA5ow7N/7D8MNZRKcRBA9AohoOJcLVRbEHHgv2QMgz82b9W7
x1dPddcdC9C5CXcVYVjM64ts0g/K4lM1NmXpUOu1CDc9+9mAlb9/WlUPm5RPn4yqidBAIc6Wgrpm
BRc02Ks7H1k5yQsEi2xWo4iihlom0CS290LmTIBm7yiWcMn0ORsrFK/C48ktqOJWwwGZ/1mf6mNh
I4w2AcfwlOzsezbR75TyxSFrSjwUpkwqp1NDNP59TB0Jm/VsULnaR2kwesDdsOz4QYtZ0GRzyNWg
xGyaV/EXLAdl9tP06fbdtcGOK1PXzvPT1S28dFiYKGrf4Xvo8UDgCuRmOcROOFCPN+jmFF5mU5ST
qbE36b67vOH0Tpjg3orgECIhShL8cLJ1Rsl4D1EUOHbkotb/n/iYx1v8ipt8az3FdJTnfrkHF1gW
4VCJVGfS4U5uslCmQ/tO/fvt6LjS58d2Lgi1gJxUGq7BORkPW2GQcq520mKSVoaie+2M7ZD+eTFF
RImmlMeLD9E7HZkC5A5yEa7OFwRjpYZHmlLtAlfXLZ/FOVb4nPKqfMaUzVYXS3qT+9Ku8fhUMU1a
UXBydNLHFB/LLB2/jJC3v/KJI0ACTexVNXaxwkciGKcSuog9EjCdHy/4xKAtbb+QVP9rGntIYiSI
21iJcScwKKYdxfrJqDX0NeQfdUQuyaodutH94TYS7v3R7J7eAHW2COhYSNbls28059YPvDoJ06tV
iZAiFzC60gKMCnvRUEzTqbuV9y6Cnf8GT09vLSnDwqtdpAitB2pr8IZ10bUSzDY6BeVKFgxIcmxK
3lZwVEPJcZlBP1UsA1WULzhh1EfpvBZlmDb7yw55G5t6t4r10GoELpM/hz00kYw65ABTbzvG61Un
t2ma39mEZ+ornCk+aaI3qMW/Jp99J3oIHswrUSROKokU0NAf2ZiSx23/S2W1d2cMeAAFwanZ1VUW
dqzcPYdkvGeP4HKbAJBNjA9jYnkoBAHThBHJSvIOmGwYTi/P7Sfox8oYb4a/xgW4V6et7YbcjO1E
CurdMK6sO3wC0lpCivf+gOScz1yLWzTQQ3npC+6AsdDCp0VKEm4BYP0jgYQ04EbHJvtX++2GSbow
g3hrw6EbrbttBAFFX+fPOykB6t5EaBr5bqw9Me1l/Q89hHj9bdVnREkyOWFVyIxl7QQQp59Av0IM
/M0NDFhGkaNzRaKeMTd8tV1dv+XdN4hlfRTlrQmPbjVOar6dTXOKDLr5sA13pHC6xigFjGc5L8sk
6p0LDuX57EHVi+0p25h8NDSHh9lvTd8RmTdYDJ6XXmBzzU+q+BVA4I6X9VGJ8FSn8Qh2zDiJBZFs
U+HrF/lwb2/XZTQ7UOkaC+yrJSOc3OF8hInRz185jLQxy3Ct996YPWt8nINXxN6ZwkOCFVSSqurN
3mwmhTPKTZbWHle58JSwayd1TEvdoChQ/5vKG5lcGyDUJ0LayJlaBxXMCkkHMi/+fwSrokP3zOPr
EuWuypzZPZbxDxQRyRSuNxfOs4QKo8QhLh9aHSuJfZys61EwZofymesUGAMq5Av2+5cWhMeX5iUt
Z9Tr9FQXXErVs80Cro05iE51h5wBFXpJmaa97MfpgF3CawOm1fdDQPqdtq1RXVhYe/EfWPWVbz2N
/qdDlQzA4aN0DmXH6zzzgTI6OHGAQ26352WgOt4HCoH0oLC4h2KEVFRdhdkgIt/iGMhvxde7BFVK
k3+efNnLMjaFZMdlO9ZCs0ROCriLdXKRnYxoHZkZ1CKTMoSMqBujWJ+ArwU9zNcvznmBrpe1rFSb
E4QOIYpGmaPa0OyjbJAbR57f1riEKohoKDAPq7vJDl/n8eQ43LYHqNr+glVn9hX+J1D8zl2wl8Sg
b9evr5yFSMwK/8MGzqrhIDvHdumc3DThvRQzvgnYNOFAaEBqc435l+gIv+iuRcTBdelGwFxGUszy
4jGraCjZiKirqeHxJCMzoDlrFTh3S4DlzPEtZGrSGXyl3+AAazJnkGk9HF4NS68zkVn0HDvGWMLD
qoZETh4ixGUZa1v4dhk6yzgjlK6UAbMh0LCFlF2DXG6LW+Aht0tZ3n/tTfQXG8qTKD6NJyHRswDp
KUKNIANYLMJss9mksI86E3gRw2KBU5owGtU8191HbIga5DfikQRNNU+M77I2fVllc+/D4sbtsVhG
dHAPWh7LfxXhrlpcrVFXmNq9S54Njf4fDoTpnNwreYh2sNfldw0pcL+576SYuOPans+eFtjEo8wT
hhS+2bf1oqyGhBNvv45owFfXxQHXvh7dtzw1qchhHse0EWtVwtwAjspmloTD/3rjxTvV33eeXrXM
Igh4vuwIwMy/DsjK4wwX5zfoo9VEFdGwhZUupigjTEi8RsZPRx6pABtGlQPDQaCc/nzUkpfs0uZM
ZEhEiUCI7zUEnsvFXkyFLcZzZmTXnGYYGdU+QCwK9oqDZp6+QdwgdbxSgYhvzUnGXKUIs8Fs/9BX
x1aHKIxiXNpc/URhRu6v50+x8IOHRXqOYH4Xuwr0tDyGEjvqXI90QoRyN6SSndY7wizAJgsbDcAu
ogNX0EIvX1c7XMTTckxZRAvb/zCINlsphqQ50IUvwtIHkKoLNYxhvSE7FoDl4vs8NpPyABxX6zyy
Ewq1VpED+vyYwzZOjrQPwDza756mjCNrPn1uokmF+zT2Z/4Aa33Sfrcaz62UB9UXbzWwPeS78ed9
I2Zx77NajUnq9yqqpe0AkANPG7F7LZIovqpc+WmSy2H7xL8NU4nYNFsEZ92fligRvD1ZrXJzoOL7
ww/qXxYvLajbbCzUEkxDoy3A5Jv5VmChyqfptT1DcV7S6O0DSMFxQAFuMcb/yRIMlPjqYDXMZVWH
e0TDCTt4fjxydjxBi7fCKX1Sm2mFw7RAnLlV59oatKkdsAwVBgZcC3qxUxt9L31ce0/s7vbdjzv9
gxmx51boDI1YV3mFx0JWfTiTIZ7PMJlmW331raVhc4YBS7IypdNFcGCxidN88kBFezDHlo63K/OL
8MhIVyEPZVYIp2C9kPAf4CmxhIrJIGCJTUYZ4luhf3HigXv+577my/IYrGffDf2MttQTgKRAw/Lq
90j8h0pUY6dfo2/n62WEL5i+8KvhEPBd8zddjbv4SwEWTaH5YcNYUYmogGLkO90mMGVYETmak8ot
SypcJtL+6VEVpAqOJLykvYV531hS7jsnylxwQqIqgRqDt+AH2C1hXhYyWed+e2XiFggaF2G/iSEN
/nqTK0jvE34SFRJv/h0w65KCsL+NOB/gIvp/87hsdboNUL/6CC1lqKTlpHZEX5GRyVbB4JCdsyHz
7PkKQWTibHnBwBl1TAJfO7lhYn1YSbRDq2Ce1JwkaakvnyEegD784fB97PA/02RMj1APx2Lt2HpO
ME+wdm3V/1kKB63wDsmf7E9jSjBBErS++kHiqEg//NqgjM0HS5wa57b+R+ZKAVR2iDfgSasGiqi8
OCt2/XX8wKrIKwVldiwS97t8ZRYAdwNII5g1Lzx2MOMf1nF/6mgPIjIoXsKl2UPL6kFV8lmgKRQq
FI5YM0PQFdvxtdM58aktD3O8mazOqdb4/33ZwkpH5lb2+RA+2sSuLvi2xMGLMxELeHT4LQ2foo13
LFYYgQO6aWejHvOJdZwekPfCMNxZlIrbbGt+lM88QD5YkrExW29KV7PurKP+enAE43CixERvoUSi
K5ebd+nY9ho586ESGpRNLpwF3GtMb1vdVl4PLtp58EN5atwgDHUR0W7Sf8AIPe4cMblvg0EulegW
oKdYVQ/Y8CQUcgZXLn9/LfqyqURBmbVn+2wJMYLUEw5pcSghrYXRmRKzfRxJlKJSPvD9oF+VJnQB
ifWsWptZb5meHvyHMTlpmRIbMUYAx6QjBTNiZV+i4iJG1XjvK5Ye+2Pm76gPNIzFXjpup6RGKdiv
SAXIo684On/jm67uBcnhZ/In1/epjXUM6dGJuO3ZUVhPVOwAmPp0sk6CvxMZ8bL00ImxhVE8nTd6
dC/Ojkhik2YVan0Swv3di8O4Gth8bwGMvylPLF9GGYzZyUyMt2P8KG9bQ2aJ7gomJ8mi1uM6mdAR
lqBFcldKfjI6ZKtmrtpK9+aRKsZBvTqH9PtMUamjE0YAZD0uFNVA5Ef8InZ5Pxbub50TxbGEzH6k
uaE71weg69MzhWyvgpARDOsY2WYnQQY4Bb8hqW3hMaGMuwsyShlLX64elgRfImTxq4dNvxKPhccY
q6HquUT3y3iuBKsuoy/C9eaPf5UaPtkc9D5v9XV+8jhX7bMAhNjpCJkeyA/zIayE7lYaUk7sldPg
uPS/giaL+bnw58Po9V11spu3X3ZslIk19l50NnkjcG5QXNxLq4XIW/KOpa0aQruoh/KiFsqq2rfZ
zU0TmjAfJOLKBOwgR24WibivvVzbDtKgHH3IefPvMmLC5zo230QJbnkuVTG/omGBAhBH78LKz8FO
gFgcqQBgH1g4ORnGIgQhRPy8NJgW8LJx7smWjX0NwbuVBYBeLByeUbTWe6EkPDDrP0zlFgYWTUT+
BQz2myIWekREcPYE9EJwd+VOvzw8OPp2kJriy2fGt91pnsZYOGIlsAg9s5kNFCdeMdC+H8oJAIwt
Z4SE543bP3uOqCdo5CJvIPCd8SSBo/XKkyRMj9uPCDyq/BxuecKNAC5a7Bn9iL1UdPxEGek3Yvcg
D3leMNcG9vuDWCzXU/f6FzeHpxkA7cg8Mhrvt84hL8LJjQWYxF21hoFvfCcOCBptdj9E2xgtM9C9
USfEAP/QDf/bgby/YN/BR2XZP8MLNCvmcTAnRiRYlcWTkI+UMZ+Yg4Wwj7jAcC2q4svnK1Bmly5R
JVdnJCqtJZH8ecPb+Fn+AH/XdnZ0azzj0snTreLozThsQ8JOYuiY47wD9NYKVxFnv1uOLAHk94Mz
PssiY07zk5XMYtpKOJC+jOmSvmhzgIJEgDxz6lljFB1oRiKc2SNbnzFMOs/cejUfFbBMg2WRQPb7
u8Zfm17Kf6wWtiO13YqP8iVu6HKoYQ7vni3laYYLJrYvGf1a2Nv7BD4D/hhjhldUSkaY8aUVuuQ0
GB5BattmnIfz/q7KmBhLWcy27g6wajkMU2XuVfsE6hjalIT3Ngxmzm5K3AsLQjzZb5nn2T2bk1Zi
ZlnhVc/69yZ7W2dj7BW1ToW4FOoKdXr4CBU8kzJILHk14ZZHaEaB7JKCRqknjiQZT+StGl7AWCuO
2xI0ppxDho56XLNXA/gv6ja3um3OCHvJXe6AGoCiqCzwjH2W9zI+KkHBi0KVYccANRc/ac9nEpfa
wzGW0BoBaTaW9ykCCQWJxT2dSwDV65nL5SOWIcMhlRh6Z7swxhsYL9DM+C7Vva2AFqKzB2kPDU8Z
jV7vW80eTY+pjmlKVJc9uzYsZd9eEr/vL73oF1AaBWKVhlkjjc0UYp+rpYzsOC9i/lPg/lgu4j6J
18qlmRKNttjpjir+pSSvZDp0Q6hkvDKxyZJufBjhGjCS8vnogVj8KZOjtDpHNMvYoFqdr5j3A5gn
NxFd7QCpSlh3ISQC3RrR8ozCtf8ldb8d29dPnEsilw/HR7wqN/1E67XKavKLV/YVrymjzzx/iwTE
OUcbHRfbUHlkIr7Z/HF4TCQIShg7/SJl++s8O1WEftu9Tu/L/oNZhT4CXmSES3XYrq3KfF1WSIS7
w6er2APmE9t0JUnAaRO6sOGnHdY+XCSdDGKO4qd+arT71BnuPb91rvnvhdUO7s3IusvcgujDRpOx
ViGGfPgBXUYk5WD4NwRuTBOklZtepu1BibOVJNZ1at3Aa07dXc5uBTA/AS1ZtHOxERqAd7b7KpMQ
A8rnChuJYiV1wTbrkSMtrjklm0jyilwOdfmgPBPOLpgweTlgFoEFg91HsNwL1fzBwM2AHT05xCSb
CJX1bJxjzQnk3ERgOsNLocNwSLqaTGnrU7xGCfWlCYPIrbXRcar0n8+sIObUwhu0VUmEmKFGIYEa
ae8A1O6m9DTh01AJGVe0afWcVnzUIzQhGDeIn5fcqWsVB/NEdhCUVh9HSHnSYgUqjLE5AakZ4Vd4
uQjsY1OenDKBUQ8vSm85EVen3vOhCAQc4J6U3Ui2YhICEalYcBu1v7Evzlhd1lrrf/HW6PWb9Ee7
+L2VD9Mz6CZtlHwgwKxUsvtnI+iIk8P+spPpXwSyUx4/wEq+/3A0N+RPQzzDiQJ5XP/AmIDrKeYK
NnBFMdSil84Q37OPW3v20CvJ4jndTj60Djl6MBxvafHkhATu95McR1sCVxp8BSBlq5QPGqemK1qB
N8U8uWP3Rs4tXVV6vjtbSi5imA6xCxwBwj6desBP1b7aBPWIvC2vX73lpPZxtiSFx9wWe/7ZjNva
exbpx6DAUR2Et22QuX1s0q9Z6/eiVjfFihUjml5uw6g0wvtOQL1Kj7Y8d7l8534/5arxcvVBwVtN
t0vQ1X0jHMMVdCgo6xpmtl/bZ5sCX47n3OWaOW0Er4iHi0v0WA8dWKBr9xn87u40C7ihTn0vujxQ
wCC1HH8itqWp6HumWm6GWBDZjDKsPoLA6zRUiLup+qNgkSxo9PgLsAGSBfVj9Zp+4Y4G9e4n1/0W
iMvWxt1QvsmjO9kp5htwrnyi+l0vpPbuwbC7a6iCGbHo6SKq/je4FaBgfzn3QpcZjxitQCHJUWT0
M1x9y4h+V/9eQeZsMLi0R8sCRWr9LimHuHOMZL0/+2+sdacbEZBWv7NAg30mi+z5W0MQTD7e5nAm
2bunZ9kYEFi7e6f67EV4vIDC/09vK9tbY7IxNbDd0BE3Qjj44aWjgHuw3axz9eyxZDE6AfvLRVJS
Xp9y4y3EKzhHsj+Z6VTavrV/Q2zKk0342GpHMGtdmBy2xNa3eS8h9HWp2Z79vMpoQYIEz6TWBe5L
9AkbitSZJj2Y0aR0aG4rtsrvYQh+v6mQ98U+qdiOa1c+rbciBOIlHyfCOsntQmQRPhjLczkvhHY0
yjalZ2yugTRZRita4mAfa+V+9UEHu3gy9yqxS8hdOGbnR1va2EewFb5E5tQoLL925zoVaqia9yvP
cYunV+iMKClFTDYonKSo4SfhmKWZB1B9dMKh8C0k5NeCccBfVLuzfgmuEX88CSAAYfZ+FKtb5UYJ
2xP+yfrcZzOz9z+xJZOSYYRvus+3JTrsyyl2NkEaPdqJw0ym+xOv+bhRY4PaurQ378NWzzSnRNiJ
ayG80rsvoKKu22PLj4JXhuc7KSAppTpI6cHz6ZfQCZKW1QU2WYD1uH+evObFvdoJ2Ruw0eFGza9S
CXfgkEnz1UK9t4KoujScSdHaxPP2RldsmZIVUH+aiuPqULE3iH5c+KktAA4GtUUlY1+BGqUHf3IY
x/an+oM8jKtLuo/DeOoircMj1vnx8xeps2lEpZAusb5sXXoJiS3wJNDyGhTORepwMoNRK0mUqiuL
xiE+n00dUK0TyUiPKm2Ous8C5/h4NgPKpwK7Zdvl4+H5gqWhaAGe8XWgHJ6IN9JJWCmgnfAFBgiq
YN595HO90kjwu5Vs3kbMSVm5x/Zv7rugLuiZdDsjQkFx3e+E5bTsWInAcoJ/ZthIv7GFK4tJ/Q1q
BlS/LSXm47xa98NCfBflAtuvafQ+O56jeacHrC/wTxZZzev8kHbslpGlYJwS+huAQnUjEMTM6rIn
hNFNZ/yEAxPQZMv/GAFlShETcz7nVpmpYw1UHsva2KqQb7gOz+tu0KHCyxJf6v3Ya5mmmT7L17gK
waB+nb5HZk8YKryAgulIQrg+0054e/VY4DKCcoCEOi0vno1DQgvXpPDOQgX5u/tPGgtZi6Ukkdk2
uQzpaV4W1AH6vl2Z0q6SMyct8GbG2zu/Yxj+y/0g6BwQE7IRvgp95u9sosl8dXisIF9lnFUpIl7v
irraDNOy/dJBedDtmJ8Cgtui9zIFkKNktrgfyk02XPp5O24L5zlAY2K5Qd2uMUO9O+rnmdY4OfRQ
qtz4rMh4YOnERJ+5NHeFAM9achMi8nIKKetqMILTOn+OQuUmKyxn2qetljvehFMR4zkEd1IWfPGk
EkVOxc+mG46ON/bC1rVTqSIw+pV3nqt1zWf17H2xo1LuxTAvU87RSZmrmow7j8+wOtfA9Hn65lUq
Om6d8dKqTCxwcsgg3QUEKsKoJxvg1RFZIc/skfoFHMfRmqqGFgco4sGm29OR0MEuylHjfcATWj3I
6T4PcscYX0o7fMPYWDsfS1RE6XZ8EvWenL247jj9Ccj5Fttk7pBOeAm13bjtmpLpNBpYrw/rM40Z
Jigh4wkRX+DmZYddG9QK/kZvfMtMT9LRPGoUhm2h00jWJtjOgdDjX4cFYhRSFvxlc0IevRfNKc4K
FEdW1YROO4i05EACaX/xNX/gFy/mfArfy6yEdwwZ6QoWbLwk5vlzrHVZkV2Ky0Tyhgnl8O7DTkOm
JS35bw+d3LlBRaNeQkDM7QOrgGJZgP5bRRaZbu06SQV5zT77SwshwkjS4cOOKOiSo0xlyORsdK/Z
OZD3HU0bViIM4TsJKp3u0CzM7wFfKvgSDWlR/ACVhSvb1hLrc2TcsXluvWzGiMCM6LAOReXL/OJg
hPz9xQkO7FCZhgM0A6EcRHDfDBo8NWU1GfYYK9+BcMQPZzMNWQWVrYP9U00FwKVwfxzViRGi9eVc
0LR+llJkXQ7nz+CLTXjK/6ntCBcaeUgyEgOehDkavBG3Iz546b762106WkLWZmuvdN8YQ2WSDZTM
b/4bJUF71i/XDQct4ZOoL6AOZfSH3I2w/8pGCbg1IlLnitk20whmSpiQ5NWjzzVx7R8Qf8kWZ9qV
FPQ2evyKTdvBlt5j195SnLfLIrtlZu3+BKbQuEUs7hbHH8MagH+LlVEO/bbjl/liH61THEd+b9lR
guK+0ojjc+9Kxss4rK5KIxgOk3/sjY6gmS28fv9sMewWwXz5jnuwZHynVnYsPqAaoh+bqFPpgCum
wFqne4MGb5n6QR0tW8qei+/Vj5lApm59VzmOfKWSeXU2I5YhKHWFkWN28X2zyx82EcHSn78qNvuM
0JSxEdKv2q4fpEobSxoYVRPheqaEsCpF6CahWdAuzyS90hTHUF9ScLX1KoJlKiMRagxMzrmbAE1S
4T6iGyKXARSlGnfQwoFkKWN66iFv6bB22j2gbgPti3+oBiwsIxvqBfIj9uOPMPmTTo6pW6INMToR
RRs6v6qXAnVqxGgZU2J+SKN5mWv4A9kzPnyHbyjDtsDn488IMdDnaJlCs5A3N1IVjugwrU7uPbfX
NZUAgVRauz20o9+cjXq4dnGaeNf2DV6qn2FduEQsNHQjdrcY0CrXdC95vVGnrAEKSst9Razl0IjG
ofhjFtRaWEMmiqZx/sC49ShQau82UGrtusGPYqJUscskhfsIkHsVdxDdPa/omudYzJjo0dIHHyRQ
RKqcdyTWWWXzmm49btAyfACHuFP2NzZidO/LSYi5hSz37Upf7bgFAAoeX6tYv5HTsOcbOa4mQM4l
tcagkEG9WBgC2yrTiltHOBL89MQKmtEUr/ssnhy/lodrYwK26Sui5i0wlPFn8pmPQEFsl+xlYaMa
vQL3j6/Dw44HeyRVShfE4K+afYaojFEzfHL07A4rpgoMoK0PNzESVdINT72bv8mfAGD15idJjtUH
n8uxb1eHUJLr7NDcueAxp9HCi31LMrJqMgwwCRDlmi63jeppOmYM+wIPGxYKXc9fzvXVFJg/jQqp
Smr8TZvoDeBLLRMLpzudGCOZmpAyKh/3NAEoT01V5v5drupaH3/9/3z6qdq9uvQnLrwJG1LVqWSG
12tG8Ov2zYp5ldDEhPrcvon+GfNkAz/sGdehR+QKH1vYHFN2FkNHnoYMnqqx4H+b/Skzx7XHaI/3
f9ofndivIVuKQ0KUURIwlFyLx4Z7DN7R0NT3QkFQqwjdcRVwLAGK/3e/Ht20i6iHLdiGkB6N1zcz
AiIi9OyA5kIgh9I46yHUKtGrTlyjqSJfoF+bAUZbTANXnXuv8C5hMTIBV9LiTj2aB/awH4sUFIqt
S++68DMdGtCpOg6e0anqNfHBbdD+/y2xb3iuWMIokWeCiewnywiq2IGdMcN2CSuHgHcLM86C25al
vGBXnHo/WKZ1Ikz6chG162JYS1FmB+9EPWwQM64TLRyVYfNY2aWaDueD8fO9flmmTF/H8ZkTr7N0
KDJzi3pFT80ynObhXXf2A61xIr+6fOzxOaAJ14E4i3x6szK0BviUxzPAwzBoF0Sr4B+xviVJ83Hm
5PVofE5C6JxsXYwg7AkCecyODNzmDuDf41GJpSSPCOp+ceyYO+rZ7S7QSEVqW0UMkCoaNHgOy3vB
d3BBbimg+caZCsosKwxqlj+2ntT6G5WBrlU1GUyp5NDKX0SKKNQhT9y5ieuJwNHL3u03jvdrBfM5
FqQtC3XXY2+op/12GbXGYqGLqF5CUmn8BjSAB0gIeHZ3UKzRkIGASoKcHo0thXukmxJQftRdGQhH
nOw86D9AV33L1M6hxqNl+zgSXkO8g8VN0ZbeKQzCtD9vD+MH4nZfbKQwaB5LSHF+3LIy8xlHMUnr
5zXFJqZTRhRxgnSZMosqVX+PZnbMN9NpGdh6DdA6VHjDqC2iiobuZdq0ucuXD/KC3uhuWDwKXR1K
mmLf4G319KtgcBk4qCm3aROOsQ0ymkv3iy+BCfgiUJq7aXRVN3rFbSpIbctZ4skPP6szcnjwf6XS
vPu1YolZwsw1CNIFmAZpBk5MDdK4Hz5oRqd0SavPubbECbEklBx1tD/JLk+1ztOvDT9Yq0W2Rpi8
W0z1LzypG6B9J8dEDRKT/j1KzGVhWqGvMsgZGGEZYxdtQ3UaBklMCKJ+bfvH8ksoDoWU//ATBMsC
D2lQp/vpB/siP0K62QxijRF/o/4S03wW23oVe2ZXEdD+Joq6dVUVA+wxT4WC40FcglN6jr9vXy4J
JBWPH3jxQz/S4e2HdgZqZABOx6EQrGvxahaYlL+5MBYAyg22RQPuI6HJftOLYIDn8cDAMUxKZHi1
vBkT3LTrj06wbWs100ieL1rQNgRXizJSeFSFJpftuFhWqsY0L9s2quEAvn4r2Dg4VPCHnBHTzGwP
Dm1FRmlKJ1+cAq5+BC4wq4ynhi42I5Oc+p4KE4fr4/kYwq2kFQwUnC+NCQpg6j21J+tzF7vzNOc2
rxrQcBA+juVEkLoXtABqgJzYuJXos+r16kkHo5b79qVkiqPdtJYVqKRFvwQ0fnIw5ivn/MNxPL71
YXhjcWVsWk7KOLpee1uGYL8Y4M0+5Ozog3zuciiYm1jJ87drRYo6SG6+hWl05z0dljQ9t2skzOf/
I+v4sT2QbAiFcuImfy/LOd1lIo0EivtAO2xbjT1YsR92Ie4H/A4Xqd3uYJdM8X8JVDABriv/hdst
Ih/jy0XlL71V2LMwvJ7Ecmkzzo7nMcMlYb5kl3SgqDYNgtOl1D8eK5rMs8+VaMTUeUDKmNKBGnIk
OHpgpHpK4tIzHqOfrVMtX2+B8+wc3isUGXLQvWavXqSwbPtau303Ij8ObvXUx1TRgvA4t0qNrCN2
5DG9ZrMtcXsp7f5xT/c5/CkAtVijtYm6D2LKxOn4O62ZKqXN+55b/aVl+wuKZ6VH8uWuEMPyckhd
ZXGN7HJV+sNWZdIvGTKRwZ3jRhRN83LNIB/dzLMeXB9Twn+LIL0FoGiBsxUll7k8fmGQ9Pvucjwp
aJN+bDPEGuhiQDGn/kZhzZvH2pzN9h9YLQiZh46rXIHdnyXsAecXtO3BuUj4vZ8yJ8n68fornLwk
FYZL89f2PF8C1hgyxUZAXdcukgJdjCtEk/GUUAxIyDreUqRpk6N1v9OMIRZMufLxC81hlLLCm17u
nkQDVf5cORG5N6ZtfCU//eHrqlel851g8AyQ1ghIq2gX8DWCXVJv/6hmtTz5DmaMPHO8Q/CFdxh5
/jdZA9GppvUyPpviHPfts35kenjMsS809zTEmygki7Ibi/4VhMb7nlrJeZPhDITPGM4PE36lShXi
478ytHDUvy/relYAGmXTwwbEV7XUl8PtFxDgqz0tJu+2q3imC1jEDB1psCz1aVa2qH6X9phgMNIL
RaYxar/Syx5wl0nmOPyD3ElsobSs1hTXfQmB3Ai8xNggPaI0v8smGnEWMM/aFfiT+7Mv9g1LitCV
5RmNqCa4uIW2oKLVraVILsTToGmcXDmMfAc3f4K9G8KcXf6N4g5dfFnzivPwfUL2JO1PRz5rEI+7
frD9C5Cw0bKA+j/iKux64hjJJvACvEcMUgh7I2cuoGSBLG7feAjtqARhM1POAL/I59u8JQGJB0tF
czr0nrbxtRF3ASiBaKw5B1lgjPH3zCnGtM+iIMYe4RpBBlXNEo37jamXMn+PP6Bw51iUZStC29hn
8MqbsstorWKAZvrKOBHlSQVqN5zkqcCay3V8Y0EMLXOnLEd43NPonZJjOAF15Q8qGKe6f4A4R8UZ
yOOob7R4Q4U54wHWmuB2AUhW3Xxet/SLfdmomM1ubrEzp7jMyFG9BznSWoMUAwVDnm6RZPpwqYQ4
xWRbwdGxbGTewnVL3ol6ZtLiPiwFhMAQMmVzvGZvtCHEeSe/s9dUYIU0Jmr7mkHr0BUV/EtwBk0Q
LFjhDj0936DecTf8lStP/gqdx02o+7kn9Jh+IlBBWqdqENcEImcs00Ghi3fOMEjD1NXfYUQNZJFw
0vWf1V0pTlUkf7PVK1qRwkY1Jen9aqSB/3BWiCTbYC34LKYviM99z2S5t4R/hkSqnR6pbW8GGZTW
EtKqwb7d4RqWKWgXFkSWzdlcG4ga52cn9t8i1Ban1fEieUF0FKB2UAudQ1rpFRPRJeUwqus1tJ4/
zi1e8bQUn960Zp8MiJUi7jl7Cn2adwzyh7wHbZbjDKPJbXuyM22ehovqM3cnLImUJFe3jNs2q3ka
SGHgNksuQswJ9kL3zoMEUwO/y//0mRSswFQteKdnx1djuui9GeNsyssGThkse/zhA6/hq+Y7RRUw
9qNQ70uhHiz98njeJZLyGx2Lu2bB0FEqNVAw/SsEzhZS/yrCi43uGCWVfJiUJak79EdT9m8qxWaU
v7bY4rFLrJqHKA1QSWTfusPeUIw5T5WLct7ihmItx9oYJjc00ye5KM86y+dMuoWp31ofaDwdVMQO
VxFX9q7vVcbR7bitrU8Gl1aLqFIMFLQ5CzMs6LoGLLH9AtT5QSj7K0QhSjih58VcBkglpCzKd03+
Jo7DmEytOxbCMwY8eHlEO79xXEDYXYXpY/XEkwdxFAKiRlC5WsWhAq495y9YKAJPc7ZEgLaQhrKy
PHmEaS+e6YkUBM5lO0DNRIq90zOv9n7LuPTPdWtCE5miOO3kOK9gWFzPiChYHxD9xArPhaWoc9b1
bKa10IiFJjT2/Au/jFcSj0EFn4WPKyYnmVEUz/4ZvoMrDkn+ZGvOyucSG9XnPgBMCkUcTgRlwxzX
+XJ8cRbEFL4ZDkgwrwAVuzV1x3/PafuEwbd9sqD9TYw6imbFpUva2oUHhBfqb/bx8O3nbxgkAaeq
WlvXNb85wUXyUDFLRfDVpk25MoGxV7iw1zqin3BJa0WFIjyqEvoxbcNz+kdWrrTLo35uN/A0Qdh2
FFA4PIyYo5z0wEzrLnCSNuD1HMswWDW429SzWr5/TfWl0xZLMyZ09w0/y3ZxA3aXVXEbciykh9uY
rHGA3EORA7Q51GVTviXAWrVhOruVepUNGGw8C4RsqTn7/SPKSV+Pg529jUVEbVXyrmjcZBo2QyWH
EbuzPCf5FrUR8TcTKSSF+QGFX8WENwIjZNkG0Iv7hVv/9UabWWVN1EHKrIXpBM7V4c2i6rBbYMHk
lEdzQQ/TMk805z0ZqCJlsc3ZpxvLkJ3TBo+GCxVFSm4quYKIMKcpss3nmO7EtPPr83UsIlA2DM4V
HeAfdAbnoIa/bh8yYldNehR7giXvXXjEXq2dUgUMVeRRPECVeefeYqtsfAVnbglV/YvSCrrShTAW
U/+iGX+elxGJQ9tIZNQh8qanhkvHPXVw/auHXF24ls20CoWwKJcYmtM/1+gtpdOLFpox9Ey81A4M
ZOU2i0Rk0kbPukZzZ2GYvPKGZzZb04zbQC7d9uIGXs8RRsoGwOwZgmXBABj7vOu86ijLV4Dbbiw2
LTMidJdlKRHgTZhBOThT46VcqSUpeArMylA345vpoFLJgnxJfqnr/hxPqsFu0Bhyhvwohg5XH4do
zWFaAV60akr+e5N8s0eBtoeGP347pmVTmi29xeocQqc5S3tp6BQtQOW3Wzxa4mcgJyBxdY9GDWSp
zMtZIQVFYPD7d29/8N+i+RshcWR5+TZwniLSMuu5jTA3skw8VAdQHM14LjNC3+fiG48vw6i8GRwz
jLvut+kYHuTgnv4e2v2NVsUfZANxsnv+7ma6SuG8+x1H5oA3HWe6KHWfR0XQyP1K94SBfTT+R2ey
Rd4++AyNUK6ol8FewlIUfmkvWwTJjrz5LdA0Pp0Tn+wVCqK2J1q14ng+zxMnHKVU+wJUSALGruvc
n/j7/5J2LOeA5hj7esh+NpTABMqBUQDQV+0Y//Td7SVykpr51MB4g3eh/+IVHMo+M38CJU8X8xTF
69fO/8iTou76UjZi/NrE2jSiGI9fRqB8a8Lvd8Vs+TIo2wUSEOm7hYU06uEHT4c/mXyCjJOAND+t
56F1JSVnpp4Od8ZVEO/t3b/ox6rWcRx/0rVgBh5nPEkVuaeRftXaVLkmYvmKIn5lCraPj05jsAtJ
HMFV5iVqB5pA1nG0bjW2uBf9Ns2KUmZ1cSD5V0BIdH4ZQfW6wbx8lMWebV4PndqO85/bKnSDAyTY
OOTyvVEqF5PCmmKkO9BCSk16VNT/PvxsCvAGGS5lpvq/BTn1toGRJyZB/dKtJcNOdnoofp+qs6Ld
ejypofCdYrk74254N2Qk+QHrVPzXhbyBIRvHk07dUCu+mhK9RvFAocwaOagdbjTfyO4p//kdwZhb
N/sB0/cQeQuGoit16FaEZ5uA9kW352cWyYPr4FykkljbkYWEQHwIaNPfLQ1sOdYqOiwhsdzl33P6
cObIdeSpevfj2F+9SwZ/AGzrnMEE6kgMIL0nEMtBiq+QTTAakA5KHfpsDNb7rEsPPi/GpDU4tIxc
3shg0VpvEYKFDdhhzKJJK6mKhcvAt85VdAxFm6Lwmd2oX6aNhCa7osRam3xoSwrKXTO765cfv77g
Oo6mtwKl4hE/NlLO+8SxzmmJtGUNt3JgW6NM+pxRbpwK3LgtFw2QhVexUgqfvlNqxjAckK0lb0CV
ALwbwtBlnf7l8UVnwqjiKRVBVF6fZSYyHhuv9B1iuluu4D18u0lUDx0GmNT0GNjLZWB+JhwfuFUL
Gr8MqNl4MNVhRJgs81YcER2TawCjnliCRE3MPmU07T2DsXlaMUbOZWFlrPrLVKX+4ijKkSHN7Fjh
oFe1ZYlFxGVvbL1GLSdXPxcUToobQGveb2/A0giOYyaEj+Iq7k27YxUDbSpHC4wpdOQhi9BLZpOd
mYyafRnuSf0jJS9gtMjBYbcPDIZJd4j4hwRVspoW00Zb8+YVeoWB4OCBVdvMinvqFoz1k+JgMdHj
91fNWTz+gZmRU6mEC6Xr0VUjyPxTNaTLL7kCqr6LSSpffCGxVMi1EqdgXGpz9LGvIouuXm4xiJ/c
1Rbbd/XEjeMnQMGz60V7WuUSKT4liQ2aHS+9hiENDx36oNGgCm8/5dRMXBf7znWN/s1iEXdfV8G7
hZPZpX5WByz6caD8Xo75IXQLUInKXD8fvtrY33ou072HUdshoqLKSMq/rBTr5R9ENgtmM65UfS/s
oVHaSdogW0c+CFX90oA2L16yQ+dpvSiBSOqZ+0cjyocIUp7TJNAB0OTqg9yQ1PKo9iQDAdpdhOxE
fLBM8Puc7wF9brrP6+ykeZ0q/aXtt+4Nwn+7Lt7hgr3oEAr90P19/4aNL0jYUtPQx9gtEtivd3bN
5t4jJ9xYQhdIj+/KXiCAnsT/8XEW+Rh4FKhZyiQO6LjddliNHc7TIKpMBuuf19hBeg0SB8J7AuMe
IF8sXpJ4hVIi2z/kG3b3KAjR4b7zOC0yE2g5g+IxHQgu3JJ3G1EB/d7S7542YuQnPqnSx9+mny0D
8mI27hNMFPap8Ip2R4PBvyXsnRH8V0cZTAv0ZOv8KlzekQ+kWap0Zjy+694Q/oGa58ldPFxvuor9
jOIANAevrz2kXv2wmC9GghFL/14OAKjJpovR5PVVNT6fIpXHfrEesN0dNm6ye3tuLMKoDZDU7MWc
kZ0+cvr/hw0odA0De4espXb0n1+INpqBLMfgY7YfvtA7VgnAqUbRijGF7mR0V9sd/iKlrJ0WblKj
j+ZHJNE6yelKu6rukQDzuCCkyUSjF5PI8kc1+cqhOI1awvVcU0aV3WVpxxOEPnHllgKEi76tP1U6
yLxHoLY8Z+QDSvEALCoaEO3ds1S9aEIh0T3qlje4cowYZmyBYwg4E+JiAt682QO3dtcrc0zGJk7J
EGPE1ybsainpzIqZ40NRnSngcpC5T+W2z6gH/0J3yajdD+lN0BOe1SCP2/q2DpOof9u2z+ONv9xH
yLH12uJLkdQ0rNelyM1WdemJdG6xDZ0f13/EREyNJlKEqV2iA23Ud9RiXD8midZ6gH2QqH2c2ow5
G6KlUBFQoWXUDGolKT54a7rwos15Kwf9m+3SzCz+QCeExwd760gLjAxuGKCe5OVSrqfXQtxM4o+E
LBml1Uy8XiwGHcDyWkXOPNSQayDuicb0R0Ku1Qsg06vGqfbAJM14SvvGPb7bHMVfebIrKUguzbF7
Xhb3Knn+nvlvXoJH7DH4WHifRE5TzEYJOIVpzLMqfvItjhNoyMbJkRO4DgiAs2QBSN2+qXn3QqAt
WgKhb0/qzz0vVoeqrpxu8Ae5qMZbVQJ57ou6R5jfj1Ke76/pWO1sZ2MxBCmF4Q3HI/gQr89GlqCO
3sQVHgDJdAFi4+4J8GuSHK4WXimTnoCVdl7m5nm1fuM6MULKXlDOegQIqhxY4CqSbjP2d2i+8l4b
0jdpmkYWY0X61+DHqD6zWBn50ngqWRw0HFO/aiFPwKn2DH0bh6ofPejL2FdQgMhnww1KczKNT9b+
H8DN876zcRi/acEh4feJ5rK9fGKjAAX4OzZvvcRq7ZXpwNIrOeyw66QxRcRMc+1n6P1Q15JwS4Mb
CEcSPMUaaBEhn5a4ShOdjxAuMq2mHylltnWNO+wcVx5zkt7yWC/i+JPdib56g1glK3206o5rEB3b
1wZzJ1/asxtIMOYQ1/VpNs9bHf9Jnca8WRkyAQzenuPSFkeK8M68ck3ZELm6w2FZbvTJDTRG+nfm
FtVezn6EXXuswhrdwE3gRDu2CZWrioFdXwh92VFrNKR0fXq17pUb2qb7VS0rlDSM47jL+c+CtIO4
QHB+PokODPmfbPoknyqzHdI+A8876zDqT5SM9mG6iLPt7A2J4KhLGXq967vZbXoanmCB/DHwPmP+
tCYkYOihvx8LFYHOBTnpM7S237J9eEwV+6LCsnkFd++cVIONrKfrsAB7S/M1SX4FKrY0bnhlpB+X
wsQuAHO8HV4SVFzJfzwrb0bYDtmixYU5pvymufvHgJohZ9eXcH5lmbUcpGU4l5HU5bc/PqtDJ0J/
cllicWjtHejKX4glg/kiBdkvErIZFbGgOd3e3VqUK0mpxeCy1VYX8aRX8ImupM3qRz2caGGwJty5
8VMyDe8HfQCapyCbYENJusnu9tSND3hA9y4N6uX2WGZQz91I3em2Vrs2PCQ+oyO5lb5Hx7kPpYhi
jFsY3ifXCgirCrb83jqRjdDloQUWz/NEGf3jza8TcSIVu9qIzOg7jlUS9v4EBW5NOTIh/2Hn+ZhK
LUh/OMeRhdphVjV3TDuoSvTvqBIRysmeRU46JjmHQA9PlgcZ0/xgvMc5iMWV88NXnNTprdGC844F
f2H4azWvFOa+m9W/B5tYZduvMl1q3+XoqQ9MIehp8zdYx541CCzNqREnXgtrBQNJB5uyJFRNmASS
0yeN+f7JE6EamW3hYddqyYaYFK9MRcqKdRTre1bq1bxt2BcUYW+4gLYYxj85EyD2HlUFta5YHXPA
5gUa0+lBxyDxvkynrVd1Z/Bt0nZY99VWUVorbC9MJpFhvZzIhtDhZriKTIv8FeX10HeLDcR6XQWa
c0MFxPw4lhsmGLCOXasiIXwF76P18sVBeDk+1iBmrJjcKcFoQ/KXjnq1r4vYgkaXG1R42QVMyShR
C/6egewl8JjIDFLmLQOM1KF0xMJ722Cv23boGsY4dbBiNSQVwAtebS9iV7St5Cni6cywF1HQybid
vT5RDvlFa+xgxcFewE00UwVSE8mlj6RagsOEepQvHqQlJL5Ib//rbndtGQmbpNUzLKEMUjFx9mro
4p9vcR260/bpLq+jtiypZCsTjdboe27Wqsa8h5YbVvfz5LyYxV/HduXxaMhbmb6s1k6lrWwIJPFO
PmZUikrhYl7QADgPwAIMbebJMna+lCJCuaVPJEbWPvtHiZ3bYq1OXO6I9QNL6yF/7yYRbKEbJuFM
x+dCHdtsn60On1zBYbqMDORaDsNv7ozjdKtQmFuerv1E8Abtk0DL7au2jkyOgCggJFlJIMWS83/s
UnHialJ/J1JiIZzkgn6KKSM8z3AtIZyU8ypCU3q7bFFBozhAYXs//mzzuWR/qD6OQK/aHLIZZsWF
SjcCDGoRMGl8h//w0YjVT2Kczx9fbuheeW3220p8DzsTwE2n2fFWEjgasXe1dTQ4Uxr6Af9srDjD
LcV0xDYwg1yUJoWAb2tEogLlZ140V3/faGEABkayN/a+Y0fPHujV2N/yG6iTClbMOSA+g2uhWGDa
bYAOvPKC2TOmDMTQt2nr6EAQTvNvaRyT7agmtLTcNfpKVA9Sw/8G26OY6IWTqZFr7rxlnSRTh8sO
VOg+oT3yFqPuH8lqh2jUu97JIGIV1Nk9uHUK4PUqA6wwBDLMqqit/aBU4qEcJa+4SsmfyhD0uANu
NkyZBeCPSyqTvIThlG2b5FkhT2EV8ktYE12e6gyJunmjeh0ph+B/nZYfSDOmrerD7gw1eSHQRNv0
76tAOkOxiMpPnV4INI4A4oP/wwBkzLN6zmAovn6sJsxgpS4ERmY1EGYsrIY/SN+7PyFM9zl74X1+
8odeEXiOyfli27jcwOf+6KzYwmIQENx5pZmrGdwe4vYjmB6DcbTLIfCJo9++OU1IbWqyfG0QqHJd
UFjLHGD2sUeMCpuQ8ewOFnnRXmTMDp9sOpx3M96bciYb+e9Onfr7gFdYu4wjE3fuR/+Xb21h/mpa
6fALKZx38rnd0fheA5kcCsKuj5h1HEUzvVukoWaj1PAZqjinpoNQ1OmugZV6M+luU3E0Z0QFpHEz
YKU+oECp72Bm2thrIS9qaRn/UH37Z9jYY6KZQ2TXRpTc3wqxqx47EPuPBvAFJN1ToH6RfdT/iR7m
KKUKslDLwcEnlApWXvnvd/kANqXD0i7Eo46hjcRaSRJK1e4+5MkjwGsbzHjx356+JGBzWowACr91
mkKQrhDyVwDHbd0MhRRkk36rOHpjZi2dloOjc75Rx3RfJ4f+t6xXD/YNykNtyr7CLWT6BokRNuHz
8w5IqQ7NGtLigXRrTcCmBsITWOEP5eH4PCVH8+xx/HgVF62FpnXzpwv2ivFtLmA36ABiBT9rmiBO
NyYsM62SlR1PYbAvFf/spE5UpFoC/vLPQwiVJE9SWTn+6d4QSjqcrvJyya3VE6Pf5LoWuQvSuQkL
DKVt/OkmWR+eFyqVdNRXpsebGHF6ZPOB4Rm/b/YQTIwImbqJNJHUdoLdVDBfL/kK14YxpXt5tblM
JYnFL13pCbJoo8egDh8LQ5/OnCBUs2aD+7knyMuH3HtAKmNhljJXkHbTj2KMBQ5hBDsWjMSaUVxB
36WRnBByLbCFv2gZjZIxnxSbMeSQUTGfxyifei6H7DPLP3zamPUhKtBPe1n83q6oCEzobezybqBk
3GaaDbFjgnA96CPcsal/qCyamudaGvWebmdXAfacWiSb7RrwzyddP1rho6+KNa0xrdyoam0XEUt1
7kqn549+B67hkgswfKU34Kev29vsvZHff8hofmxCpFyXeGrk6O6OsXeNiUIhqt3lUVq4fdTKVhTn
xaudX3FLco48P6fVIMOpFRSs9hs6GZfmUBEPi05USn3mkwJm0MN+QAnj0wiQMb5r7sNMXCpwm5Pj
+MXz8ZtT5uelo0vG/9AHaOtgEXck/ptsTNhsTlfwOch+i0bVBPkUgT5hZ0Z+chDOPPMn5HDBPNXw
mHqJO9rJw3gguBfSIt50R3Sr95MdgNgCSTqx9mqKP0o+0WuH8e1Y9JJrzy/90y3G5yJuPJr0NX/s
QRr4c+zgwtgI6mbG8V7s5LU9ONJX2tS/sDn+QmYtTFdkQYR7x39WP2wQepzXwzbN5FkvU/4oNNTH
bEf53m9rmSFxwdgUAil/CqPJVLP3Zw2Eovr0qSo4zc/QDOU43qcMjy12bhVJues6VaGq4zXdRfeI
xtOcDb8v4pQFwXcjKATuvmQWqBTFx0I7Az60lDXlptghk7exhLL7+XX7nrDS4jVdvMen78XAF8Ll
q6yozsU+uYRNhLdBe3JjBhbaVqJHFqMe44Kv1I1VLX0FDW0UlIaJ5dFTpe8ylC3Px6oS1iJG1aY7
z39aQEMYKoDTYXbSd3j6o9JJNVbvcyYqhtc0XidmLKIYKdbn7hCc1fBvMJvYuTEnumxCdqqDsesW
8AJRz6XJweB1n8o5gB/9PU/SHkigqalujlF5wYBzDvVLG2rtRnTNeBV8/thGX3Uq74+vtq7OJqZH
I2ABLbZ+PZYbDf4mNRXzv5CAAA7KPPYD53tlzBArT3uJnIPXw79ls1eZLUfO+iN0rcllmWfVNTMX
X5ACdox8E32hCR7bpqJjbosCnAMF6hwo3KzLGcTQrKYX3eUbPDgTwpJ+FBLwdpJSyJ8jkutk0GFb
OIxGuXGQjPKmiw+/B2d3tds/fvcSZk/N0N1j/fIN6KP/kwyImEn65NLBtkBUOKkskV2Eoh112Iy3
bF0/5mDzLtDwh97fx1e57AegD9xouzMSUika2gl/2USHHkRERJDYbMwpeka1BlKeO0JzEl+UHX8i
aj2Rq3GeAaZpmMWH9e3eG72OriKjz8j4HDPprLjQH1SX8dpJjZ6mr5JDzDCrGuOl6jfSXHSpt3Ba
LeNGmm7TXVXl+JH0RHMOw2O+al9LFLQwrlgARlZhQorILkYj1uJUn//oEjJo/5tWKQZyVgUXH7KR
vORKbJmCKNh0aJaX7FpR0XHnbBZJHxMLqO8KXQGnPAsusm9TwSALPNPw8RgPfufIPRjd27EPkpZb
QouvchvVTEnyjnC/7rTa9VB5MYIZGk2i2mOl+i0tgFT/1ntx/i6REqXrF2hm+RN/rcR9SjkmcHgS
JRhXIU6x2aRUS3ZRK+/nqZIlV93BAsy8B7n1+65n3oruqh4n9nzr5xJktK8zvWuapy7h13v+nPFl
qA9EZXhAIQQhXgnNDwDQaL68yls0/KDXImER/rpQw1ZRmx/4KlBEaPCyPG0C0HCo4seQuJl+EMrS
A0Y4QQSBnRE1yPH5i2Yyvp6cYqKplsEIxFHnfYbErrf2RA65bCLwZeXo0VBXW4BD8iLSHbEfsEis
thZ9/s/lAq2R8hqUbYfgtqQWML1GcZDp0A07SCOmtNABaescLenmJaW3dNd5LSRza+sw9RGaBoML
rfJjBttCEdZhluT5IKYImP4q2n1Z6/PoeSrqa/wcOuFGfWuPD6qbXaICRL+xjjS0I1f4y2cCh+Cx
gok6WF/WW7mj43CnoDgf9241YKmrremTiOuXVJWnKkMgpPpbKnb3f7BEd0gIdCXM75LVqYJg/aGE
oAT2ClxsEmFrvrRxbFGcN/DH5rBR/GIqp1N3E+3USfeL23vtD7QGs2ndTOzu5JtVusP8C/a7vu5B
pANkYrZb+KGMnE3YrehE4INXFzB4HVQRDtyvmekllvGwey3QY5v1jszrifSXLF4qwuKZl05TxFcW
5hvgLsMd4HeBDCp6ALXlx0CJ6Vig8Zclaqr6Rf8HonQcM9uMNeAgBu2WOVLaBOftO+n9XGUBfzvI
g3o56EKnIuGjJis6kyxvwfm2FRFAFj5XIsyFvfiBPoJZzd8DAmm9zkwpluICdBNwxsFW9ktvptaB
+fCtB7SFDDFl0ogKdaldQ21AjXigAeaotwMKCVcslJksqrvxjJejEuVV6glaCeaQQA9Os5UsnEzE
tJ+pH21/Wb2fbh8MUbEl4h55+g425US4XxEvH5lYs93Erg0RKFf7yNrtZyTI8GdmDForzEtf/rqJ
Lby210hVQzCkfgjYxW+o1XU3+JqVPkwnfleLl+SBL5HckvgoCrClvm40FvkIU8Z4pglnqEQmgeLF
k+Q1JNJpyyahyO1H0Xu6uRKw3b66GJ38ZwCmwtL5hu6I7A3xEsfCh8Cy/KdZqzdgWiAqv6YKd9eQ
m0c8v0q0ykIr5tSLUp32/ZP8pwuOD6hNvGd7I3mHeeoK+fdsdNjVnJ81DGfQpsx8rFKyrlnLS0lD
rT3TgvBrrBKU22R0vdLSc2A3Fsh/zAiRt1M1XOKqwyFkqC3ltdhuCMAcQJXzxnWNfftVPr9Rf+Vq
WgzVSW2XzZSmLUIjZVeolpOY4ylphq1gSOk7vMPKqxgswoS4wf5q0Cs+D5KH5OXlBvVmnXPJ0xcV
aDs4KF4qeNod8yyaVmT0qIkOE5qaOEL6JPimlxKNat5wHSGhiTuv48zsjd9bw0bylF5nGnRhbQsP
6mGD2GieILlQb/KS33OdUEYDm4xm4HPf5w0wxhIAJ7zWD8nhtRPXxe0nDAqGYnQ/sHY8zMi3nQmm
El7wcNwcWq8AmWPyvuAUqoimN7Hi4p4ak2HtxCzGmQdtZKzaNEV0wtt6d9jjacEUpE7Ixn8ekHsO
50klR6GXeZpPNcG8Is8kcEuh3nkblXz5AsZKwH1Npi8L2cf9HiBYrOCbbSLwvllU1+7h8He1lMfs
vPCDVpkQ9Ixs01K517pk0/OzB6mLEfzEAmx1+uhccKLw56AqEHYDd6QPfjlB/A4SKNtvUrRDYFyE
UGbZt+KbJKfo+C5UsparVrnqtG1WsfqSHQoprdgMzQwfdkJUTwZfJTatwTyHfG7O3bZXzo7K30R8
SYMCQpnRiYDHx+FXmexj8dvkovPwXx5yvTdJaGVtmYK+rraOlMneLiL7QE+9P+PlHvaGtiVUS6Ac
fZswn3WmutPrqhNl90w3c1CJLZHdqW8hD9aiMGPJ57IxRB7Pf821vIlSpMmRDbiQwknhHIbUIesa
kEQvcVFIiU20J735OXOU6Lw4lmFh7/etrsl5pgJ4rDGj2aj22YSnmuBUUeKFc4OtdbYeSVn5y5Z5
ihMjPascoLT38GRDvg5nWnhX9Z2NQYcydrZqMjCtzpGq10phvZ2z3F+8PfVk4SukCiJufOfvA10X
EYi+6likL+r35E+2xgSU5r9bEB1kyilD5aBXHQ3yNrTZRfcXcLN8cocBe1pH0tBvyAOtOjyN8B/K
m2nncWychnnf3O5KnWQH9JO5HJggS2nKnwa5TU1ebpcaN26gqPV6S+iIooGWtuntdaejuqlDTyXX
91nzIiDfA8T+eEb2hktL6+sn/hVghg80oNTqu/PNDTShzcP7kE+aFzQEia/GblPwTVjvhYvzxj22
l0KxwocByPL9zpXAkmRQpKs5w0ijOjT9XtTIUt3X7rpun13ENo3HvkifoGJgAkYf4aop05yyzRhB
a0H+NDu8sqQd29nEVcPpu+HJZJ4vg6cXVZ65Eepyd80YHDMDC5T9nYaD1SdT56+s+lycpT6blH5i
QxMDTbNUlXfEuhk1fi8VH9Wgf3qV5FMizxTdGYJE4+cKpx6ckqZO5/eUB8jjIdoEAtfwigZSxZsW
PoEqumMnjJGC4bJVSFGnYdfBg2xL8pxs+TYsihltAA0gUgu/YpZ9MpBgVmcxaZaX7V4FspeAG3nB
bCVFBrpkSwbF/IMWumc2vl5hEyemGy+G2laROmvvPlo2JtDlT4J69GlCDRut2jGspEHXewlbQIsS
G+ZqOsgshNPhE+jW2FwtTFsejyMb64ub+2BXCN5RjmjYhcRUP+c1zBz7BvjSzEnGVDES644N1Vfk
JeUWo2HjYioMn15qzo7FfAWfcmi2XyK2KXZ1inc9U4MPUb6m2Y6HNeSuACABNwf9Tf4IVrQInUYB
R+X6GrscHqmxh+5euPkKuiHHdvNyYDu2nYTcZTU2yIQXo1IuhT40dtoZmawrjlM9OLHAWjiWPqkd
oFGb6ri7qW91uaK6uh0vmy3NVpjea4g04Ooc3oZ/q4e3YVQPxToLy44Fh1+2UAnv4ed2wenb9i5l
uI2lRYifdDY1RfFk3WeHeohBa6/pRNiJfrHMzabBfwMTu/46FcG6pJUiMTG8NjbVZLgZiDjdlAPY
puRJJsm5Of+a43uP25eaxXZmDKZY3HL0YEuhwgweYwIOTRk4Hx/obHSDM0NW7MQJpX+5oKhLnvBw
M5dA+Ab7K2Ug07mWOekwMAsFhLLq0PWqo70St0X10UwODIwPoGLLBqi9hbbZMY7+WZ/SQE5W3yxQ
jqOlADuw+Z6HeOLVe/0VDq+xF1vd/WKVotWs+xK6ByHeIFDd+44vKUjcgx7Z4wjB94Va5yKk9TNa
zXW3C0jCoh/XiAG8IglohuW9iShpgUia1FSXIMY3SETyqo6cWt+YkLB1v0IeMQlyBNtmxxZH9Cm+
/IXlu7kIfjpALwCDX1jmjJUXHsyiw1Nc9bI1xrZIX4+gUY3yx2zvtzd7hQyC8KXvx99ATR0ldGol
KhxF6HdoH4NS/LXNRtDw1BtRzJZIY3gE+JkPb0UiA9afH+KRonRkHJqJ2Wo+xzdHI9Ut9Yxp0hB6
xbRNNptkr/gnZijbcAKhlOgnQRjBpxar8SuScurNCQQ5j+zpz5HAyUQOrTqSGYFO+XPEmo1VLNky
5oPNlS+bf7UTvR33Gviz+i7szG0YndPH4r2jWx3A+vkp59Qs0h6ajQQMZTgcq3b341dzZESgtKEH
g/wLowT2xzcvsTpMs2zMyJSzzrLogU8UQZAuC70hcov8XbRDCpTLYEJg2njoccZS6TiDUs2veilG
t2k41n0k9PtQb4o5R1xx1B8ym9MdK35ZnwG+rbRUmjOSPO7+S4AM8I/cKwA/dC7d3H7+MZ6/Apy9
woV0kEYmKmB8NG62GTjrVUkyxJf0IhxgKkCwt6vyINhvMo26Lag20OB2a7dH/Q0qmj+h6gESeS5V
w2Ub5eLrg/PmIj/c1RDypo1+VlCq1Jz9+R1QqWpDQpVlgXoGcs3oLkv/o87D8PlPmEkJsrhwEGgx
9FEV7mcFBij/dPYT8tL8AOldd49ayCurTk43dkz2fPpr//K9NJa5G95icSZEcR65f4ho40r9banB
E1I1tXRpD4VVEJixPHqxwxms8FqXxuwksySr8EiZgVSknT8Wdb/SoSU1MWUc8r6HM4XwDz5CdL/3
5K57Ht0yZsYfaQ0Qcy0CBw5PPvNrke803ZfsAJSk8k0fnAZiX9K5yTa1itsDUiOarAFLSDgPDBra
LZnKtdZZgqSsPH6VUJCnrjJjBgxSIQPw9H3JIzu7eOW9uIEBVej8QLn8g3tScKTNHrztW+CFvIln
F1Y/5gZOqPagAq75iUj8oR/MNZNN7HZz0O4tip6J3As0JF0+nmRRC5UJynG7937xrfTzGvfzzyGN
2orzvP9jJOmu0Bl7iMprmWJ5tnPSdzB/wm27/3548BgadvVX5RW18CEuHh1IjRY9eLwt59470JqD
rhiaNIuFSEciF+fjPtM2YiFEJG7qxYjUsJ02MHBvMKUX7oy/U780keEiTLtgZlHaAYh/iZ1Uy1sx
uko5ihT/2i3kcPifq3H7XRx936hLqrD2IL6EHJfU8dnqFm4uASHAZ4E6HmQe+T3XISDxl0b28ssL
VjH3jV+4seGeyQT2h+ayaDad+9T4uD9FkRWyGpct1eOZBreKMqxm8fSVgvVLlfC8r4zj9kUEfghQ
FUB9zJoU5d1SduPQoFIfzpdQA3I6rqyAMqmPpDW7NPyCE3U7E34B41BPycEDl7jKsSC/LwgDdLI2
GZB22wslgO3KYeZINX2DgUR6NcMpyRlcF4JycS70fwFuZV2Wr5quHOUq4u1tSj6lvY17wckYTAcn
oS8HWb7qCn0oM11saB7uz/rNkIWiWeuF7zeKHT1KtHRPVoS7RUXI/198/aiArW5KtZCfhI2yIzcO
k/MQ4c9tQfGwnSgLGPu/rDGekN+pRDmAxJexlXpJVgoKPQVjQxv7N1mENkvh0aMwHRARH+APTa7N
+Dqr3w7Y3uAPcnAgk2n4cEJEb82plWltzymLMHft8Encp0/+LhaMEFi4dM1+nHpUUwRK3sDD4qNV
k6UWtJ6OcD9syJ4x2/7mxyy6rN/XGui+AChw07Vk+KEE3IeUWp6+FKX4uRBsPO2/zagfHav8Sxnm
1b5AO+6bhZBqTppXC3CSDEcvkbFO521L/bZu4Ut8m5ZxfSA1pDAcuooJZRRiN0i5QV5yeNmUYmHT
rHxrp4UblcnIQ7oZ1AZw54v0guyH6tCc593AZjNvxIJxCEdNKuUkzSkKonTnLWtTCv0HaLyuCX2u
LWQ/ujbMOWe7xSwk+qk85SbDH8pzUQAnxJNnBS9UN8imi9yxriXptu8+bfdMAyn/e+Nj/g8ghCLD
AqmhVcbzqGdmxELuRcfIF8LcbhEOGisdEGdufj1Zxf/yksQk8djb22byjFzDUTW27aOhCkd5Bqaj
2mCr7bmQX6hBJgdFoFctwOYkbJ3jtreZ04/btJrPoYNhue94+buSxBx3U8qOUCIfMCavcT+6h4hS
y5lbUymMxZ5hBnZcTBdjFrySRl37mWyhNFzdzP/RKdKESY2UER9tpPTt49WenDUEeRRTqKWy2I2m
PbTN0wtrWq0Fy+8eRikAkqvmQFq8SBonN9cDkpNZ3pSGqc3ZJiLXohsrQmyLN7DbfMz5eG2O1ZvQ
q4mczS1csKBJ5DGDMlTFQHPWUTvfJfiL4G0xAwuGRHj0qu9DGvBgfiSJ6BM8KhZKIgNyzyMGUW9G
yf9VJf36jgg3q0Eb7hZvJok0JFdtHmpJG0hlUoY1cHk72kHdpbq2xmCWlVAcfYBibS50Pia+SUiq
9CPczGukWh9HAOcU5UwgAmTJ44JRQaTUp2geWg6iTxDOtwY7MBvMHXnDrWGkzfUntvXGxsd3WtEJ
bqlzAzpNdY2+E07+3Xmia09zgnBr9zGJv4fOgPzK1mx+36ZjljLSRWYMpyA2RQ6HSzCECuApDhfE
/kcR35ZeT4WKWLNcId+I7py+yn6kdt41AFMUqKfSYrgH4RFqOTSqhYKEkEGRfG8cSV9DeVevqP+1
8ubyrydl2C2tqpSC5ISq91ldL6uvo3YrQpF6IM1C7sQr60q/bfYQWrPxuGrLilGqWcGzOnRxVTI2
OvqPWDRCrkOrIFjU2gBdJH2mcYxCYmAA9Frva+o45jQgt3+gb/PNs/rrUqkHPK9xZYVwb5tQwrFe
X8lSBnq842YWXiYXJz3ZggFEqZIKtP17CYbGRJkJs3BngxpUtZP6xC55QwF6y80GESNtopgkUB+m
cfZLsGV24SLVoGHFjT8EadHMHao7GKx57d4in3uetZjYiVbexCt1/JxtfEkomRRHfWR2CtoXO7Up
zLKHLZSrH1rLoG5nd0ZtIUYPpP4Igdvw5X3jZ4hk6xzcGX2em5S910/T+PcCKvYwbETivOI3+KJi
HmXspkGaW8AYNZezSkv2A9kbhPhgB2P7+5XqKy+SU8/K3tBeL17uIuPeh7mRMZnFRCR4sSIyFis2
WrmPpzrtaTQk6NfjpMpa+JcsaGEc0xQLV35F5i0RGuasePjR3JcW4PpyZ5z6SrrJ0ldixB8zzX7C
pt3KBtuVZXRkxfFUETPIfIjoMdWQ4fw4O49gZvJKVi8FYtJ7tyV/EtIL/mCXaMXiUp7o1KhhExcH
1gXlVweTrdHjr4nInckbNdMK9RKVPAIpfAiM6Wj14ZWdjYwwSzIc1TO58cFv8MzCu63MKNXBC2ta
K/wecbKaxVREmQL9A+9qcAQdpTyKfL9B/NrA3hv9IQicN0YDYkUKxxSBCIxM3Dippu8S2TCIN/Pg
ohGVnet+iwlYjz2y6gzr+A/9cwv5hyF7ZVHDbyee5Vl2Dcbczw4GTdyFDslPqD6WIEtjk8fs/tXC
NPUJaW1l8EMpQEYxVSegd5y5fyX7uHgtRnliUhAdraVq1cEFNDGztTuqK1Emx7AFW5YsR2oa4/ub
gNe4THZpHEoxgNnO06OhjgQCvvjzeikQOn1DOWE2iIqHqPHTU7248mihLtgtEP3JEzQpBv/hRueK
T1FypGf5zFBlRIyLysxecoC5VnZ9MDir9FJXVnenRsGPWh91clgNUiarhWqnx335vfN0AnAZEHTr
sXofn2yjyPRbA1JvEENgcTTFGeLo77d12BcXu5Yh8XmqxoQyYzysKB7xooL1WZbkycF2Y6KA+LTu
GOi/h0m0n7NaVj92QBRDbjQtGDyj8eNUNZ6MyXE2RgzTXGotkRYhSGo66CbLJ77x+CbjWeN7TNmw
g5vbXBoZMjMdrRllqv9u2MuvAQmGvRxE6BiGbq3Tqu2q88QzOktEpgLjr92IBFSFAahOSq3pXN3E
B8bEs/20GqZU25Pe4jNocYCjtosFWLUEnNwZbIswZERKazktAlWclVV6PKkHZKzAkZX5IZ36SDEp
29Q6aaAtxJuIrIc3Jb1ReBngN7uxb3Npy00d8MZhXTwpIYxt6lGVGQKnvLaaXwWHNnUNAmWae/Tk
al9ajXSVKIkDJDfC22P6ma8bACyo+45xGg5g9BeVaijHW0tDNDNEYYzj7gkZaFS7EdyhQvQM4R63
V4Or6+21JgFRKAw31pN2KIId0sH3WWrPd6FSgonaxRuFde17c9Ae5eksvvUdOEDwx3TD72WwkfXq
81coQ5pCj1iD5IaDG1pZDZ1kunr7ID6up7e/275Ccdq+rJgrhoQ41qw/AdU9hQa0bXmixyT6D2BI
O6ROnB9XwOjb3thWAlXyvvrqLNI46MocRJUDl3HnUrzt3YJPWVmUxpeKgFQ41zdk5dQe7x4wxA/i
dg6xzPpIYZU/K6cuX0XWq5l21qKglKoWv7X70ONwn2DNy9PFx9WW68g/tOYbqbYLhfIayx1BBJ3n
RC6Lgk3vmo1izPeDs5+qQtJ+B5j9apjNgxk6s/QT2GhhlNGG/AFvT1KIJ7dBRShzDAlq0T9gLTA7
gNhoWe0pkFWR+PmTgY70/SfsRtzNi0XEtw9D8W4t7MopDl4euVX6fvbe1Dbr6dQXmShgq3GMPKkU
TLiHPsad6MZ2k49QTCmAIJEt09tWYVDV5QB+TNEJILVLOuXd1vACUy5zcP5Q/CAxlAHjZPfEvSTx
3gkAfGRKcwCv1pLRAvEdWlSxYN/uQcRHDewTZyf4LbQLt1f+lGmmmHj2oJ2sspO/NR12M5k3s+HY
LrArWfSs855jJzPQbvZOQVjuyeAGgTzlwesJl+fRwCmDZZHazcsCcmZTuFKlCkoTJNrid5dTQd9N
8TJJ/C5y+ZJLujcY4froHiyHr+lUzoUMkZwpZTPPa4YFiWH3XPGBBuHFLc6//NmQbIYzyYhAf4iW
oQy3IHlst4YAY3r6FDAYjKpV5oT+9b242vTDU0fmrIjy5Fq9im7WBu0VeiwaBnr8fUcWVw0t6Y0B
vxWrfflqNccqL0TfVfklx4APrR8OZn4J8mMmPdL9bmX9VvKNitWGptt+0tvT48OyazreaZbEs5x9
YolXayAt6f19OVIGAu5wog0VAvapWnctbiZnP3vYXSWrHQEbuu+QxkIRREVrLOFU8fY5jVji/cdL
HMYxFxfzix5ISZu1DJ0g59ITY6Llx3LYKKc/fRfJJRUcsDMmAY9HqqvJ0JWOc0An1oV++J7NN1MC
SU2dJRxZ75zpTn89Elf+XoEgypn1We1s94jAgTbrp42Cht6j65wKws1KmEzUizXBEXFJ/z0QUNz7
JzgaJRVhAJjrpMugbstyJj+7Kd6RDs/PSwAXu9+ACOsh6fx96dX4msZb/0xOBKZk0LN7O5occMsG
9g3zCNYI9bQY4UwcCOXvVfDLJeyW2XCilGnGqQiLwwsOkeqsXL4bVIxGcZ/R1qJKFriNFa6R4iDD
tScrSYyZgr7q+M7Cm4TYa7J9p8zFpgMgi41RMdTbBdYuCQryo70xmi0c7VO74N1iwwRbEEGsbs5K
WzSm7vOIuXiYs/wHWPNgKswy55FyQqTuQ88LPI2RzA5DefbAuRDowqB9l3ue8hWvKOFmGBb5H1t7
e4Dswen7gAYO2V7x3FPf2GqQlZlt7Awp6Dcyf0A09zAlhCFnlGvRCmsJKn7nrBsyoARfwHqdl7ug
RDxkuelglNChRE8fUWQcnxYPg5YdAy4ifLoK5sEP5a0LavafmbLgjTgbQO25N7Ouf+q6YaUGSMq2
VrEzA0TgIH1QxQLbjEcpr0gHrfQIKNWjrruKhkdu/4upNoKGwMB2SFCDKS7Ia8ZHN6KYCIczixSv
9kjuzd1r5mVAdqVYzpHgSywKlPoAgT/zZCkjDmzwFpNTz/aNmNSftkuPcgczTGUpwSCpUr+uZzLD
h+4j+CcZu+nYWB2ScNfF8NpcrmiD7mkXB4GQqgLiweuhUu9SiVyOfGJGQtTolAh982O602yAVbPZ
FUlWIhF6exoCTB3Z0i27L25FjdYuZEw85uLL40S0MzePt6+jKLaJGYITmcddPJA+hszLm5z1ZSt6
SGenyTK4dMs5Q+NZkRfrAVziqd7n0hQVOOvqh7VX4RZzUiP02EfN4/TeORE6jF+5aucpe7Zf5Prj
9QGiTGNUqNST94bZWt4xvDAT4YrhLtMpg+xR/F+jn/+vOkCCEO82p7FEZrZUIuWNbAqHur1sGrPP
LXHJjIQM94s9uDO2sK22lRqnZXV3qFyOAap4aPVqr2H57sjWXsOKygZ1nxgqxQ9cIZMY/1ksPQts
uCI52417fPgmxP6ajyRqCBXNOCleLufrfm7k8uY+RZwH51sK3z7H8a+VxmMrkp+Jr2dpIlGcW7Bm
m/oXjrd8I1Jk3mNQpXABYaYGrnyaxetg781iwUD0VkKYrhsRjHLulp+dobXV4FiskQ3Q/NydmEkh
oOx4BISuEFHSqiFqeb6HcZW/tMAdn7IhvW6C2/81sEfgCfVS6Nhrqn02+OX5arAC8CP+CIFozy9V
1krFPkaH1GYVe1ZJ54eecT3NEQ7/qT9tlnZlTshuk3dEGAIWdyTBWp0smCkzP1NYfX5hUk2PngCJ
xTKMn/bMMPcFFN1X8pyhCj4bbxzHibuo9UnYvKJD9bMeiXoN1rINzS/jRBs/4l6mNNp6AXnGrBMu
gZfHe3YgygsOu4vMb1TCAm6lH+bmGQg7aOBxep+ybB5vaQQkCVdOHzTMPUiq3i3eUgtdOy3V1YCB
sUlh3P1MZ0kms08vKT+gzAuGYoJ5wYgNaGoj3YQlgWu4wMQCDXE5p5+Nb7KrmIcKbNhWoJ8SqvgL
JEApysnd6R/2r8hkGobZzoblDaiC0L59lA7MFB8iUBypkj39rIxseaCchd2D7hVbGbxtJ0SMpuk+
CmeBqskbk8U55kU1bQh8GQktHUVv7GVcSZ6BtNEdEKpEnUG+Zq7nA4Nqhu2XnGqxaSBadq8ClH0m
xMALqCMYaNQDfdH9pDJ6nRRi7s1LOnd1rlFPE7s9JYEsSqCoOklq5xDcRrPb/DLOlTRmFMXpPZx6
PMsKjfhmwlu1QtTh++q6sHOKq5m6ckCv81wms7LtksN1/IODcUdCf1OlUTD7DpIxYHAAFnyIYyAK
XrFXvsmm36JmacUJxmWE3TgXYcT1VHNLoTm1j1SKVYoRGeQI2lBihN9doCuYRbF2Wc3x6LHVG7NY
iiac9pnQ0W+VsqPylzq1mM96u2hNdzZKGaUnfLYdig0h48HTqAPdVVuQclxZnpY3O3Jqk5F1mzf8
pteTXdWXjNhlurbhaRIOHJOVisIDC0Nj5uyben9cT74XKQbsZTlujQ40s8q3TfezoU9f3IUHOUoT
1uWr/IYpg/Pb6sVnLIbJ4ubKflYkFX+5msC4MFBvDfKN48nBOpZwlzoC+vBPK39orNwF4P22w2zq
5yZ5rwCSKOh5Sk5BU+PwY8aDgscdCpkYgdShBrVsTeC1lHm0IUoANlY8XyVsE66l+XCVbcGdyXqM
xubpwQs3NUUXsHl4KGk8J20Q0YuwVNgpVbpoTiUiZUDX6PpRaX1uNEQdp+La9q9Rl0Ng3pu6xpFp
dL2gPGwohZWLBWkF0DtUKT6FK9E+fZ7gtfTFrZAtlzTnmzNJSMe5pkGOAya6JYXVtv7Im+J0oh1M
O8QlB0VNmuMpTILfpTsXKVaVb1hozwoxoY7EjzaACVdDY5pwZPej1U4aMRz5pU5A2au8rI/DlfvE
FeJiWwIhw9+3gzAAC2PAzC3SyfjAnF6p09laTFZqoKWFB5ypDYJ8cP2jAphaxbAqti6jBMvo/LWV
hW18dhwlUw38WYRwA3zRsYNjqBFbur8ak8oewxAV1lPYsA/KD8uXMCqccVTmp1jHVBcSTogy5Q97
3SGqMO88CWpzS4OopUuK7S6w82DYwsx5N/rLlwgQWYI0rXAa4rWBe02ba/o4oMxozuNIJ3yDrAs7
NKzGBMwMbJlHRgW8YI6UEEGmr06Tlc4vemA33n5ozWHc8YyT5JO0UVgBlBY93BLC6C+yZ4FcNsxY
ZH+M7VazAzvsn4b3yTfKbxVF4s/pd6NjIVYm1/DTniCoFqAVGkp7/aaJNJECjDucvFOrfpSj7vAL
3KcOq6vukdKAt312WSPzv8257fw2vwizqrSh8df84J09a0POlc9g0YNwY67EGrAUkm9u58dRMjMi
/mXGS6jQB6SiTA7N3D0oABh5/zf7z1D2GYF4EZFPc8kchVqY2ubNKS8ju5nQ89Q3qRmfY4rfsBpc
SRl0u+/TM7IBQr6NY5MSA7uKV3BwimGGYg3cRjEAa9wYfoK4mOMaiACic4nKJppHXU15X2vso6LR
O8ju7iqv0ZLyroUiQZCTjcHAYCPkCF2F1lDWUrlqOTfZNicDksTBtXq8jaWwY7kLZtuonhjlyDAd
5ILQDqGV4IzYReOBs9vi6wJ+jjPX3EygZAqKNTDehEVUG+73LAwjTppZO2owNsHwqKZlndhB3p44
9vSPY+LZ4G2e0isFwXUzlzdXXrGt83xPT09HdF89oQFpi5y56m0w1Y1FVeD/PVtZp3YGGFrEidyQ
2DIaKJoEqpKfKPv6ZRUyaWcqTYI6a86AEqdAMyb3zE+ruYCTy8xstmXn7qIWI/9sxiaF9GZa0O4c
LrMLupcE1loKk1cOgWRqs9yVKACQSgHhUSnt9KO5ZlkXW0uk9NNosao7HNCiB+KS9Of/1CISKV1H
flid5GD4HJLlhex2tQIXm4Y0VY7/yTltLT4r8UGF7k01vqxWrMd5NFNscDbouE4Qc4RxsP0WKcZJ
FJTU6gjTftAuzNCNQDBqo0TENkUe3scz70yaXvTU/HpwN7ujY12BXdV28ZrVvWexwp3pA72OZdeK
Kqyw+tmKppWyuR3ZBGV2kZQXqlIsEVcB2+3T6xziK3ewlkxVZkwoiuxwYi4NQT8kGkCmtUbevlYR
ow2MzZgU2fEAef+Kg23qIkWPIQ7O8RVAR/JCVz0TRugNSPdjhQHaQqagcm0L+iK9xAF2vpuwsYxm
aeb82SBwAwVqEZo2sYi+FNm9pCgG5oQR8EaelG7+jv5xfbSI1NoRY8lkKMJywU9vLKG+qk9DCh8h
AZwnQHJvuCa2q0jHRQVvNUSbN7JdTQMQsAiT6r8+Cuo9t9Gjhh8jOSjYMpaa5Fimp2Eat0/KdmWn
HkSGVdV2kjLgNlGfJUAOGBHlMT0tXxjCbRuSa0Q5ZFMVbgX74ptD1VcdQNy2y97SjefYM9uJB8GP
2sYvIhI0C8fCcTz3ZFi8wDLbahH0u61u3td1hbIdo2CTu5vU7QPo+RxVVx9MRJk11/+xWLW/gO7e
mLwBavA3WkT4DNwYe10hWK0KouMFhkNufFfLCHNrVKx3L3fzwD5C4impQyxwvbfF7CUtJcVjilrn
anKibrz6DfUr7ms+nCG5uveITm4A8DHl9BFgHvCJU7CsvBzcImSCyxp1VRyjHmzE2RlIKrrIUhIp
9EOuWpKLKw4CBRGMDhToRs1DH+NXQsEc5HeOXMULkyeXK8ilq/Q3dHDQcl6jauh0XF3DJJ/grN0X
gH+0UdcGQY1VQqVEhKCsVexwcaUZOOEoRSQ7MllE0ajuh2JXgsbn1I3wGT9HHoXUbGSQzvaXt1ft
OXvHO1HC9avCGj8XqIwEn+iBQdtwCWdella9JAW4Vv1v/8L1qlT2ns6bpF3S6DQwx1hN2j3HccYy
bkoQ1q3A4DEss5EQQq1xJRoroD28j4C/ujpxdLcL5PRSiqhgO1zekOH9NCxDsY/U+Pb77UemNkQo
Rv3t38IGQ9tzf+BZwapOKQ0ES72zrL6gJNahlydrP55dBiY3L6LI2IhayrQCa600//oJ11MZimgl
dm5hYHLJhs7IXhTiRJZ6HxQocKx64/ddyJ/DLju2o2YEt1pBDvZMWKk1XZ+JyYuhep9eU9s1+iK/
578SD1odDKyQ44sc4SZyGldciUAqXIO7nR98Nk0Dx+HBc3npW/t7kwqsN/26AwQm4WImJFEXK4PN
35gNhaIN/o+GVw1r21H0e5fVyQTBjE7DG1ykQoQfryzKS96mvZEZ3h3wQlMbFTyU3WOJnBNfOj3C
psVf4LlsRYy5M9m4RZdJZtkyHrV6tMu/3VLieeNdWLrXBws3DL/QyC3Xjl/ipcUwBhaBvtt126vB
b4jCkrXfTNwTR2pL0wBrsK9UA+QO0njn2K3mvhK0+YBb13CyLfibBI7bnl+VuWUNIc8K7fOEXX9C
4eg1HZ+DSID3XmIMRWcoaO4llCVFiaEIp7Zs9VHBRUPXprLLinnpmjmqiVu+jjjIJuyVXb+EL5pf
N1Ri/l3o5DkPaacnjFsx7TOeG2nZ00B+GJcT9q2ybrNZohtITxWIp1LHHHKiIxwDr2LQnX3cxhh7
uJWSiv1/P1xjJIOQXxIvN9SS1Xs+2RoUxr/dyFIOFITkcn9tY/7tHKEYyCxa6yhCQ/PeCyH31VcB
gc5NVDtsxvQ7nK/Lj3dhkvefrPuzu5SnLPZjTOZcUF47V0vOb5VdhxDfkKeMjo8QnDK5urcxQ/gZ
iXe8PeESZJ7fbzp3avNFpMKODxGCbU87xMrykingHZpHQi/w5BWIZudtCyCKYlS73dKkUo0Aor89
C7rMXbol4fs+R/V0qx7z3hfkw1wIOzaRx0VwvD3caRcXnU374gExQyzJKbKa75O9L0P0NUCKAE9r
ZKRlackcVsFhihkGX5YMKIDoARriubEtGZdqZMPGVOmvfHfCGA9UP6npnpkMY34FRqRibTD5Ky3r
9GqvmZIm4DEYc2TMhhbkJDW3E8EtiezR9dicpcyPtPCKsXJvgu/6budFgRUr22iuz2GH9OunueSw
eEKLSGTBxNTQwvJEk8w6g6KvzoH7QwkZVu4GqztaASGxeaU665nhwebOHlBhBsyrzBjeXr4lPeYr
eEP2ZYlEuESk009PvRGlrZDM0OfY6Eu8vjgLrIKgwrlgVShhXyvZAB1/T/6VJ4bp16f1j5tOhEs4
ZLYWoIjVHQrrkFl6TaaIgzbxaC5MMvIIX1W767pNJ1aPlUDk6i15LHssMMsuoxUZXEwleD3jjeiJ
aQH+KH/6VVp/3+biMQIoqK9mVPs4gs7cNyxp+G35TLJT1U+MqXc8wmL3B7jc+3slXQm00QiyZLd1
fLTf68TNWXPLz2S313nGyDsTQG/v++7+XCxCxEv6R6YPLDr86dazCG+XT/FnKOOTD8mGohB6/bE/
eDPr8im4eYxglkQNRaxPlO5O7EGRuWNu9aRj8+qibiqpKDXaHpOiem2R5RY7n+doCgAMpQllF+ZT
EOGO42orS5J8AarYxf58kMg6dFAwabnDyeoIp60O2oYQkqPvE7B+Y/a+Br9iJcnlKF/HUp+5cs1U
l8avQdUw3H2FsFtnmk5y9MG4x/k8rCdsfg3rnqYQX4G1q2oUQzwrts23LGK0keX44YrVJsyOYCd3
qOGWHhvrv2nmXv775DIAkLolzbf853J1L0yOXQkm9MtoilFrKW760LqMW18k53thtAyGYW70wX1y
R1rgOHNbBxHV1SfkBGExzC4jh1/jfOfB8n3uNVEqfXRjJO4miD8csDsSA+knRHClo90Wv038R73S
dO1HGW5ScWLyz1vqGtPgIsonX8CXF8Y/yYI2I5LrfAOT3G95Q1H0S1Xnk73kpE8TZVQOQe1NKCGv
UHO0VOkXD7r9RecU7wUB39OG7F8XYrr6Uw/KEAg2Q+4fQJzPY6Cb/qqmIZP/w3xmNbaDPX7GotqN
JWZUEk3IjnM5mbqfN+IEf+l79raB/+m8uOupFKML+AZc2gfBOffv+Z5KEWRXEUsb9ssJYJyCDmDe
Oqe8DaLcQqaQrQk08SN54MJzWKntd4McSPigjb2624h458R+aZfqv2l+ZCpwANF/6CbnRkjLoKgm
priXh7SsGMu4Y4D9V1U5DtsImxJtUJyuqzyfaRThZ0DHBULMVIUNvLm/dA+zVXnJHiUKdhczQRnx
6JST7K6C+Nop4VLGS2KPBio7KwyzUhTrsgEpie3edEr31hKmxl9E4t0eWsq8e3sZjefR51XYvUlk
l5SLjlSneBAEScZcaupHAOxy6VPC8Yp0/DLvpV9Ol0xA4pzKi9EgyYfANtDSMP4aLJIR6JG+W3wI
CbRb36H/LnnoWEiLq8UB0vQYih476MNF1g6JmOHUL49VpkTX9x3ULVP/9kMIZFzH//afx7sW1GGN
a+9ToDfaTBYURV/gwGatyy95Z4uFirN0etsIp7B3AoQWgPIQ19/MAq0m11S/hzcxg08gXGuxRvqG
TujnJ4HqjAeu343/U/0uEmhxASDihz+a/u39YA4AzHz0Ix4rpPUo1h/Cjt52XmigjGNdKwspE+HH
ZAPpdagfdGfGmdflgYxi5zvaus8uaWNnxTpCQIdlYat8k5ifEFtD+xkREtbvMNLol9/SC7m2dBHv
W28ckVVINeX5ni5Nfs4q/57VCCkaUs05FwmbJJ8X4MbCO+5jynt/ULUIH1CrgflsYuANhKmY0YyZ
gU15/eq9oELaLgrfESPHLd4YpssOSMSX7WZp6oiAnU3WWMK0WEQDH3Mv4eiLx9w2FmZw+vmsxSYh
BMCKqaEIBeINH3ADi9nn4FGQyifrh1qxJ/rGNoZVJXQWgw3EK7f+IEzzDVu7jGPFyZbkYSpfLCZV
boDMXElkLgI0jGhrz8UODmAsHGaksuQYUA+w8DFbJuSSCEUYa5OgG3axdgQJ/ST352/5xTG2ySFJ
qR3suY81ebqSWBaVo7CDQkF6NOIXRMVQFQQYAlInv58AgTElRQt5hRCfbBjz4/zYPDWU19OcFJtM
vKxEnbR5LUFN1XhC47WBMj1TK9m6WQp704wDx0gHwzULsTgOGvCEnql8n/gHQ/8b/n8yE5kEwY6M
QaQ8wX+H/p1bnFq5vVYNMIx9fr7D9LA3AapEYBACLSo4XRRkniWLv18fisWSpmhpAjMRh45yzdqm
UJvCkyhZ1AqmaRrp9FQ6gdyMnqoHK9DpF87gpZ9hLSIkDquugNB2f3mTejYqIivhDtSl6P7dWCnT
Z9o0+ZZKn67rAfYOwA9kXIkK9VDZ+472dMMYHWge36hZ2nqJSSw93/ujtTCzrRuIuN0T2LvOrS4B
0nd0gGxB9ekM6bKZLns/CqpumLKVieij8nKmjMqFrp2T5uowe6BsaZ7PHTxjZys1n93xUOHCtGwS
ZDYB6Sf3gpa073ZSAUaT3IwAMqKNDrjY8+fHHVSKWr11HuYxPnYh9ZzYE9G1Vl0NEuPFFxArSD6N
6vWgy8kAm+XkA7GRNqhSVk78U18bpXgxfJWkklVEcNSAJAkvAVeoU/y2Mch2sb1Wa3kCRtelMB3u
A5+riFdDL7FjDfLYI9HV6iUEDKUsRfKRmitaU76gvaa013WzcOeWkW2rH3iWPdR+KQeC5EgiMjI/
BW0BTu1HdKlWucB5VDFSAmAJnsECRwQ2jxP3oXQKlNJhzKm6oZukfa7kl1uj+xG0iD0v96elbtDB
ad91Urbjdfiqa7Y/7Sh0BWUFSeINA0SP8icWgjhEsrQbjiTCH2cvcdUzzV93Jb2diP98F/kzJ6C+
CYwoXV6LQi9J4HA9ZCp7Ob6lRhFpGd8u85cAVSlFt3+KO0DF162Rc6MLtlbR7w5srhqxfUSGNjiV
yagaQplEsCA8Oq+lC/OjFqgISHyt8jVqLdgcnEpbAGfBlwD65uIDsZ4md6hAptSPrX7QZ9prAIg/
FYNnCSNtGn91+Gs6aX2CV+FcADa+TIwl6h33MQPSNNniz4ANOuj6O3Hm9vyhF1a9RSTHnLWFqyoC
tTq1yb5wnMF6L4oAyw1PZWSW3fHQgmeOmEdIjWNp+z1ThkMFjzK+lFJXgCzRiUdj7oK7UeJxK20T
ZV+cjpTd7xlOMHOj5iwO2I86hW9DphIRtIiHAZV+yJ96+c29RhDBIdw16MSMrd95LMyjTnew4Mvg
9rRPZoqUeK6Nsyd10kjR/PV2uIm3Rjs7GklGvNIsgDRgm0ohA105AuU/cpvjoFNcaCzI34Ng+j+g
vo3QjAa+vK8Coml3gqx4F2noaCIESHP0zvxXjfAFop/v82tdVmm2MtZnhXPqZcKlJHa0aZlKwvvC
eYeqMsqAVhF4SZumthBW0aL2xZC4GNW9QVahmlkp3qr76/aE3aib8tcbx7zE7YoIeP2eE2EqKlXl
AFIRiARKiF7xu+B6RcUl7mBo9bgVyvzLXphQ0VWqgT/CFC8y/DWnNmA+HN+An4WM88pMf7K0Xdaq
QCv5mUdxB/VTDJ9SP9Mv7EjT9OKmo4lSllN3ZtgNEBr/Ga2IaIDDXQU1fp7aBJ06bkfHxKP3lMkh
Ria3oxV3wsEjiiZGZr1uolU7kNYQ/yIAH8E4imj/OD9YPUxtOppx7myYI//5X6tXPTEwaChmRzSU
3cJFgyfQen+JRXeuweVujHPTaKsx01sYCZAz41IvO7pwKFUihSp9/M1s7AgdS+qdjVHYf/XBDeix
NVae/Z4fcB0DNinl5pUR9pb+YXD882MLooVVMv4YNX/ktuvAL1fLB0nqvFb1JQjgfu/r5jfAGQcG
4NcbWo+2pF+LO9tF6bveQYcQDTFkstV80sbuwQ3yRvuPnD+kHzSrLN4HZq0zC+MUuhTP+tb4FGQE
7g0H8ziuYiLwMf8XEsD+407BmTIBLViRUs/7dTlKgoS8awi+sOHlqQelNp77MMmqb5tZjpTacuZ1
2j4ip1KkO2KNOylQMTFnq9PV4jWTI9endiwXC4mrmThrV/TpObngpguKXKD6K/8dLLka/t3KTdAX
yOGlAuK9fPwcYeQPsX2Y6/6EcnDjl0D4I+EuOHsIsfkF77kiPZmUH/D2pJS2rFn1i/Ba+gamryYd
LsNA2kptduftBE6+n+9IexgfPONBqkAEcfVPgbDsGwLtxrItYrir0CPN4neEHkD5REUZCOwtOZ2x
RxDIqzuiv/Wc2HZy5rT3J1MTvDkfFly4sosaAjdbuYc2Krwx8zMIOOFO0ajfs9ZoBR6ECgIhBGHm
pFM6Rl7yEE6pvpH697t0ukuNf3xRGuOS4uUKI7/2VrxtPjjNBgUlmm/oQKwq63zV0hSdIpqck9AM
5ZoB0wwEdVuT59/hRj7cTDzWOwjNJ17eXnFxsnPILfaZOoaBE6uZsEfVYeTPZTJxu7KKIpvIBdJs
yOIO1zxIdZxsFrsZaH/JcpyMAbBBHowk7s70SodCWvJBOTpTTgDfE+L+y/4xdsYfldysL+M9uHtm
WlYycbvTf+erlSiwDQRZ2fKyfG/Y5Lt+6afgSRUOFd0MfwBqyL8RuaSpCpPrEPm1XB5RxFxoPj6A
us1IcplAh1NuWh6HPqPb8NjRy5pYtgSOj/m9RESUnZA8iHyH3h3fAQHItR44AKfGhWFHZg7CT7Ab
fIGRr/u2EGueXNODW5rB4dFUoKuU1ykEMtQhQqfXRe03b64FBRHFpYuQncWmQNvfrntPN/peVA+x
XMuz5I+A5tu4tysW+AcAAnXIJQ/NtvJSijf3DOchO4uCM6VdCqZBfh3Dx+q5x+60Qz6apk2+QU73
iz450W3rgGJi1Pqt2cl+GhX8HDNGBjs8LPLfEoAGUR8W8XLYmQSOcAZ+IpKzUHptLLhYRSqHOIWH
k41sqCiPowQIZRsp0w4qDfcmEBrNvtd6jmEkuNKy5wf1cmMost3SOvu7gdttsyhsamewtiieWWuw
YBDDkhM2mGYOSR1FYC5oWLUMn9FZUUEeB47glHkD8g/tRHDvgdp7+Gn3diK1022LR+goKOVI5/A5
H1+C8kdycTImtrAz4q9I/A9DpVcDoaDLQw3pM8uo0zzosrqq5zFOWoORkDvGum61C8ak279hac+X
b0W0Zv1B/g3QAHOt3KkZAKAqTE+I4jd+iWKsU/8wZEM7yU68xyTxCFi/2R9Fs3WpPDjmglEdwQ8e
QCKQcXTbBYqQ0jTYWqy7zFu+OpSF+eD00jWK71ri2awiBgKXOn/4PAHCgcc6yD2PpIpJa7pgb/Uf
LGoEHX6oOqcIo6tPAI8HofxMFyiiN+jAbJ7IslOkASv15x/4N84YoqEb8o39554mIx57woNfP6dE
17bn/L93yZfc6MgktbS/NDCsDBARR+sNyKoYrA0ocbHu24gea1zbfJe4nAKMoTORrJhAO2q1YuKz
uI0qJJUMwfLV5mx7pFMuclOSVcaaiDFOnVS9xP3hQ5JQN6xn0sReNYyxWN+DA9RdnjLr9twmC7++
YBEQINWz33dhwCDkiHccw07bEKpHDs8r70uS87lL8RBVDLVaLkVf13B9Ictr8vbTl/ZJPPQyxX54
lsCBiNSNZy0LvqBUj4oi8ywksAv/UHuYF3UCumXE/qN7ECJ3UK6hkvUlKRvx9+NSSq2YLjnvxUQ5
ht49ux+qkKv9PqWX6v47gXf30tJBb9HsuDHXzeTjHnLnNH4q9Lv3YL7FsshvYND9yGBg0+vINzax
uuE6MPWAsT5+9GVU7IFoEn+DHfHH6xrLP6oYi1tRqTh4vLIB7Z9jBJHPtVp8xI/VjzEos+MnIs+e
lgq/2tXg0AGJjedZqLxIwxxaDl0ceTLrILTJNtLQvpHRPRt4ITd6cz7/nYOpxbKyqaJwuSJyI4DP
vCL8/Qs/kl6I1HkvE9Wk/hXG/PTo2v746QojTuUf3xUq+SI7mLlQKyupuVkZX6ECCOMiAPkG2S85
OlXFgsjzCNnYJy0Ukgc13eiPxI9jfzrqLozZ2J04mHpas+likADGJT4UBLiBm8SKLoOwB1V+Xb70
fwGDvkQy3jYv0GFWGD5lYJ2U+HVMiVZRvDrrnAeyngQ2JG1Gt3PabGOQpQHaQmZL29wHl3HBVT5g
lRX8waRP9LVC8BKjaUmuV8dFLgd0a7m24SAvVQ7nzhisB+d2tw8dqAYlrudVlcqo1d9W8/VY9mIa
8gT0G91yyFlORRPa7np9U2ow8lQsScFmDb9wWPZIk2BuoF7jbJ5cH5OORVt1TIaldYklqJIJxwBA
Uu5AoFargShIRQeybxQOto8cRT44LNhGvr0vt+NHhnVvkplR9VKUPpiOpnxGuTuoXpgs5gWvs6HI
udvNzQ1k95/BvNxNkumUkIy5MdnY4WUjSGgNAql8RDuIc3En+1tM2f96VMIGcsAvSnbRk8b6w6px
YtU7jzrBSN3ClJfZar5108jtyr9sCb/InHytR0azuWahx6NNovOKs+mZnCxTJddMFZ3V+XvFI4wy
3lvr2rx6B4sWFMbn85stIkHhoJJmP7QrLk3aCM21iRS5RM5MrU4WQI9tR/TGV+VLlAIRcDSxU/IL
hjMf7oGoxolFPfV5gB+t8mVtGrMBL/6/GZi/LRBOOzAsL3Fs9IJi/yewgA6uXqfZ/n2gCA4BuEVj
v3Er2b20+l9dLzlrrZ6LxEbq5dIrF7l46TT00E190hQG4jBBeUWyNBrdA+flntY25JAoq7GmdvfX
rt67uH5L/r4DabKzsklR+CbP88cuR1JI/r0ggO3Nl8LtybuV3TNXmw92xE8/0Mt0Ws8L0DU4qajD
jhiVZawgy4bU3heIsGBGzhoSEz+NVUd2o9af0Hs0vGIw6cX+yT2aa7hcZgynsXINvxqIlBX3XPyy
A9q/huHigVMziIfGp5h0l+sjWn/axfF08jD2U7UO49pYLudkrxQWk3BkWJhtSkYZibr6qfwoqrtf
oSWm+CpTr0ccBGRAq231W6MVbM6fVKfSMsBzjXR6akJR+2jm2mURc6yuiN3XC9YyxJfse88ejlju
SuHsqtaADciNvoVr6S5EQEGrPRZJgmKelDgBuTAND9QSBqCSYvEYQIGt45AijtlTT5vAvhJ5Tq8Y
Pvmfad0t/hxiymapGclHK47mGwjxPyd5KRqBCoTeWwCVxCODNBDUcnjR09FXDbCF0aZYznjzfeRc
muYtHDh/vEV6NR3wmwvphK1GX5l6ySBp0WtzaL+20fLSjY2C/8F5Kb8E64NaVSDXbLGhAQdm3ppI
fdDaTczIg6GN0bgGO2nluXtOV6J9i+gC5g4fVK4PN/vsIwZd2AEnGeJ8jPO3jk4ejnzRZfspaUYX
50Yz/AEPo1PgRhcJOyXcTjhohniH3tSf7RQO1Z3QcAYpZ47Tx8p5K9iTNqPPByecVnJ0j0r6iRas
w0ic8JBuoO/HvbRWuDEvSpdR0WB18DKxE1Qjk+rChfVrXXu2qXAnmQOrq568BVxmj//Lp8X+Vcmx
I4Bl8cdJSdpfTLPdgti1o8p+HswuUtrfXPuo7aRAWC1xZuaCGfMJoCu5H3/YCErwzzCplIMY8YDX
dU2i9bsyvwW4bjtFB8SeiBu16VKGq5DMCP9NLMZsnmDH1HN/31NtT6hFiuQWH2+in81M1k3HpfSr
gBGkxE6flor8v3/LpixkSvZsyifQjLU3ZRgE7ewv5H9nPZ+QHDawIQ/BvjiC6o9xUc8AS4PrysW/
nffTYcBYe73QI+xWJaYylLNRpHPfXY6YHd4jO60GWPJKuO0aWpNMLEXb9YiYfN1dYNpDENo6U2wc
1LLwqMxGHcvlLHEHVB9sRXTwe9slThYN11sTXQn+rbvE656b6RtbR/WxV9XJ7Iazt25ZM1b9KoDi
u7F6TGl+e5Zvbp3f47ktMvLKPCDqBx3GwidEnK2aopSl5EJ4JbDKcWoYFwlnQFlGb1cDXvkGRbAQ
Bgnb3DnP2/3FKBSCgVWRkwzNBuRJJOFECcxZxVZe14g51aPc0rgcFsfzA2RPPacmsr1MhC2As9sb
LzeR5QrEXb+CkXRYo2NkQVHHwhLqA5jzlE5sajuy4ANLluuTpD6fhhq4RNitDRyH3jMb+pKmuGLF
sGEU3fi9zjQip+aicMYyizpm//izqt5M5vS9BC8tnODm6LB7qFVXP8IgDnAI5auX9/EW92DCtARJ
LhOUKVVXaRRgkVhnYrGrQaBHppC2Ab+cUZR46+gaG2rVj5P0JuWVRWU9iLw7NPmy3a06VRr8bhfU
+Skp1mzHi2AtK47m2lm0chgAt5IIs2bNracVbB8khMBxFz0l+XW4lbHM/JCa07oKvadgJ5Hw+whH
F8ukpAC0g0sHG1MUGrCN4h07Get7q5DhQdgxXgA7vtnri/JyVWs8oBjasfale8/52wdmIrT6uKPk
W6QuTMvpUPO+ALrEJbDLHnNTlQ5N8F5xmFUCNbwvjyL7UCgxwq8RjTbBffZefHf88yEggDXLCCkD
7nvpPMVpf2WEhOSXMrDBqP1Gv8F5n5q/SjIxBGf7rak83jnR1bE0rYYkgTm4ksgX2HFaA9vf87/P
s/XAbr7OLFisopF9k5+wgqOPdoVdrO5DvCcrLC9+u3h6eiPi5DwuXUuWKN+KmBXsI/vcUzCCzXrw
h1wOjJFwSrWl9xAsZ7tXXk1bC9yRLgFcYWX6GRgPd8gSzFUQByHXQ11KfVDsmBgRFLyMjByiVK+9
y7iaEYyaaP/Pfas9BfsktyqXHvl5Hg92Bo/luqA/RooKLsPm8szrMl56yEN0RvtJeM1kZYyMhUlV
FHTfYO6RH7WqsrrZw88mbKZwVC/X+K8eCiHdN4Nebml60Ds7omKk/YGEhiks6mVhlckHEF+xofTW
Rb5HhGcFhw+GsES+mRVQZQMdiMHWzE8Nmb5xlBxilrVM+DravrMFMxRtyNN+LDwxECz5GvmLUEwH
y55jkDPvcFwDimmeGhhRKThGsoEUAhl95ugdaApoZIRpDhneRsN/GJFikzafkr7qvpP9OGCy5fE8
S3b5Z6IO2Mwjfh8Lgk8NrHkP+ryuEd6vu7C5KKlezSvFIZznzEGLaINWZdMp1LQ3JHWSrNRtM747
dMmAbaVwLVDE9gJJenoh+yofJgv+StIN3fgZbBW2dG3BE0CF5rpv/wtsE1SdCAh6OG1LO4RDzhOL
U5j80KQvSIS8Ol1eXRFDr7ujTtS52BmX4CSvuJYApbtVAK9/J4YVJ3pFQy7nUUtX3MiC8/pPze6e
+XuQWMzWrL7w8QaPPOJGPXVgRjtUQdpMp+g+5WYAVG8KAYSjbXshzpLKPeT0R+QsEORhQG+21+9B
H1uv8FqOYFrnN4gaZZY7wiotQkHrXjjASEUa5drnYh3rB7ZJzR20wzX7IUw222yhe+f82Pgazocl
/Ju/lX6/JjlYv0aBrgByVGGOvyeX6a58nSAp2A4ugNdJ+5tS5IiDwXgoT3E9Oh2N80bP1KWmJy7u
IV74PEuAy4fsTlLRMRFL/fIf2lZjbOUmJLZ5R33+HoMaagylZR0wlSQT33hEm8KMTv7ZBOj1HAfW
HE9gcwreDj6a6nVo60XqAkWn+36TOWVWOkP9Dqwple3yPQgUhbQB13OWYr/bY/xJIVs9M2DnH5+U
MovqIQmCR80fN7NUF9FcUwMtoS+s4+9ovJozy+tjv2W9EL6zKY/OYHr8mEjz/K9EhvSRJC62MwsO
t1x3u0w+f96byIWM387V25JaO1X2t+Zi+qsmc4Ji3eiHNk4n5jLdXtHuWww0PoW37ZSjJ58Ue+Lh
2FUylc2FD5Ey9Qxf1PU9WBlJfdKFvkVjs8YT0sD757BlXhyBKC77C0zJfdnYCBkoyOq2MYWd91md
+Cfa1l/7aeR4JkmYmH7MECq0zWTqWJUzcxr5XW3HOPj3i21KZKqchqxJXMq9PITgDG6tTcRi8mPC
Ad4iXECqeOWyQnW2NrkoFYd3zqhdS1M3LPbqGcBTiRvQr0ArMay3TkKq9XUN5la/FEqvpbzdDlTK
VxCsbBltNqUbgA/fcIBSnoGVEzczNmFixhU5tGp8wwi9j2TNezwh+F1F256NDwdClBNuPbey+cWt
qhhqawfyI6ytDkoVOhbyBQT79yVAVtccYopcPPtDLh/nsUSKiE94REwp9xrxWuzw35caVPrILYxr
lKPVIJhuDVJPmovdAdp2kRNchI36a9VCdyXLQ7zG2ZE5NZQBLM5Wg9kpvNHFWu0TIv2FSFkKiVmC
4mvFksDbYkoPhUAMqvIpt9tQ2E2WIAgRIgxhcDlQFaLv6Vmgm2QW5Wbq5T6A6NE8+M+IH10JV/oe
Qp4FT8HMV3vNkT8DflIEF9MBBcJ/Ch5Tr9wh87SBq1pJgjKSGK+QCOJZslod6889y0xLKvxdlrT4
WzNIiNC4Qz3EoY4Nmvxy0MEcgWrEAAshFuhbnGyW/A8m0InJJbOKQydrjd3aVs+Kf5KMRjg2hVPC
0fnUbn/EqtkYOAr9AS4uaq4z1d8h+YJaykQgnH8QjpZANbJ4qmTL0mn9wI8tWQvkJv21Zh7n+Msi
Zyn+GhkomteJZ/3vjfq5faGoKRp6kqOo8qRYcAOztyGS9LTqGI3o5pQtXnXofg+QCvNRMUp1K/Ku
oXHTjJIDONT8mn0fx2zuLFi2sb7IOHG1hiB9rxm/B6sSyX5nex2SUPUJgPaLupf91o1BGhEBTh36
fBcYFUZ1mLH/rWuXCZuosHpxk9Axg7QZNsy8+h9bTNGDi3IoQyf6WYeT/3d3TUd71foUCQ1XmM5J
wDW1jP4hqBxb6bbR0THOqcOVoqaW++uoWy70KzqYbBp96TKKngULPEwrluLASXvAw4mi4uo3K+0Z
leE5jUW+gr9+cll0kzbvZbTsO9A/3zDGKEfxtP4Tm7cbVhi0za+U+LuBWwxJrMRH4fLHgy06SlEE
w8US4Ts3wUoqyHCQt32on73w92XllQwfCbHM0VWhAZC0NsWWcosj5ne9n5i5b5CpSpbY53Y5YduW
2hXdhFVdAMfGlJY6POtEcJiTvfgesTCD3qgjim7pSDJrrWHs+qdo7gyNvV4xyMXE2113ibEKeFYf
+NscW65CYbSGgzf3cnXwxfBi++1COGfpYwFGps5jVH0M8DxMwzfWkp8brSXIMoAv/bQ2KIjXiv1A
41rn0prt7vFpPIpIafCP3vWNoCC/fGkEo+J00/5qtEuVhryfNuBWNM7497/gadsVWAzUOQ7Wex6f
QkjvvywPe+8cVMRvCJYr5sKZmLpQ+PjKo9OqVgaPPrw98jSigkPsA+Bl2f1yKnhTDDtfPXSFb4o3
anF0+d5qClB0xoQ3dQp194psUxxUTzDF/zvTruIIr4spDpljjdhNKqmEFuKFe2uM4rUngn6zNRSX
LfPKeW0JunTCrrGQ5Z+ol20w7H/mfuDDOYvNg6auWOuDu0VUguggCVYGHNgcpDLhV5+1qkDbqcFq
vv6H2kc34Yc3StJaCWU/EyIek3vjXGxvHojZ0nf0fpKWAo8JlBLO6EldTc6zewWerCSdCpOCpT7t
rJBcDv/5/mTQMF0vp19rQrplyJHPXP1a+X7Zg1Uza9CJ3+XihXha5mfiXrwnL8ma7aWjPhB+AmVz
dXgMmM3G5EeyqhxXocEgLH/Vj5ONmGGtBZzaG54n5AGFTGmZey3izVYVHbUjH6r3qlk5seUo1pXG
w4xMjdKiwYpjIIvsVjAxAHJZZ9hOxOpHRwYs0Ss5gMAoyLHKT/XyzCnxHq97l5zN0qG0wacaHxe8
VJ1iAISEutTFDvOuqWbZOEO7yi3m++XY3T8tyqjdMNDUZl72aX26VDKWziaXgb2c4Jvmdz4I+f0e
ni7TA/IfaS70PvBDeVDWzGHwsAr4gxp09MWNs5VfYkVrnFpickW2BOxYy/fFO+vj3FbQJX8RDey9
hHBVRa+ficwe/hsB6OGNkKjcXhAPgFijY01Ebs3cG70uojwKlMPtU/y6iuSwSQxqw48L9bkg6g2A
AgEZbzY6SwuE9buLaxGJu82OiF8M7aRafL4Dos0EcCpHf4LOFq3/WHPuQBNid0ivHQuW3WU2IKs+
AqSkPDxSo0sMqGg7kYOZJIfQlso9QeDxsFhJk12+fHPORyUnL8dCXdlQADN+YGy31IAPkA2/zu43
zLwgIZH3Sjwkbz9OS8028Z0gtK5FTsRLrq+8Q+LM6BRzrRhPoHEnXGsO7O4JADAOgl508c4kzyKc
bibhmXPLqVvU9edtZsi9ugFzNPXKb8pq48gsGrX9iRfAhcuM8V63zdo35mspVYeEhoHvRNzfrRfs
g299MqCMbYlyokSuuQRcAHatl/dFuTTgx6ScAqIi/NRdlFMXdDucIQgxHrH8Zw3aiZ0UcSJJaQv2
jaxeNM6mKGK94AKB0qz63g1HOml5vw3VyxtrAIEtvHfbDaFUCj14FcIDfCFLXx1/Cqt3skYq1mSv
pcpatD5oPNJOSgv9/GWikEvMqpUQ8Kt5d27oKZ1fsjR5nGr0YxTuV0QQ9HD+QYAlbOVg+6/be8rO
7hl5JXolF/m0qPFQ03jUO0Pz1THg3q91ub6lOKn0/4KLHp82BhCCPclVLukNfvVI4Lj6XWfWvDrA
lJuXXFnGPLYvAyxNRU55c/N1p74oO4t/7jTRAXpY1TUes2cNa6XzLvjiRJAKHWGSyVoJNRInDs8s
B1Xg43uzWLFhK9wT5W3Y7gHUjP4QLGzPujeiGMkcZ/ascdAPu8ECXAYzaIMQKQ2lTXCSAZ0mH/ST
nhBLCCaQrSdUTHfrXIJQQ/OjhRGhkfo1YBtGsRHB0+zlW8zNde2gImBnYK2YABBHy47BCeTrEeJI
MgE7EasIfqbsPLCJgT6fxDALnq4gqen7HtI4QF4PI722tgT4nreQtkHy/uj3nQpkZ7zaVN21ZWLt
64x4rd55La01aalQlJDLCwxwrUDSQMnetsaglglUx3McweS6P6eCHl/enVAMhVX0vpMVyf5hPOFQ
3r9EssN15W210q0FbR6dUa4l3UiOQlMZ24J+ZO3cPiU7yNRQQdxshfbj8UoWoLHk0JrT5nUlyYCh
SazUEJZWdxyyBGJBv3+wllOzCD1wgUk6Wzza9LYycS98G+M99gMPUxRcXbNoNCL3eDGp1MxOqZFX
dGfpN8Xil+3TWWXcBqWgilmpEmfmQLH4MXZbfvGkrn6pK5XIjJCqi/FencYUl4nf8rg/i3F3z3E1
Q2eZCZt3quxhAHCZZwtVR7Y/U8eHj+38eussVhOEVtCIb0skM/RbPgUNhPKteU7S2+1HIDU9CAFT
pcOS2ihbrbByXSQdLoNDe9zipM+ys+kQO2CaxQCHUkYV4nQwlpE8wMiFgMFGL8Ii0iwEHl6aVgFB
HbEhBeNhL/JQhFdK1/And20abynk84g1Iaq/VMVjiKqaqRm35X6IsW4uehhtB4kt2C4xTOTxDPBI
ugXPQYyDiCyXz3jRWK/uFyOuZzmeTCH1Tt82t3urtOdOhDmQzuLepg5obq/YJFcwRqAO4Ff1g7cG
qFK0lgHVxptftjhCT1D/9UCNbHIizH7OQofOU0xA4a+VPX9HpCAgJVSyAQNlbQizjH0HqLa3aWL3
XOGczQe4CGjw3cgmKCFM5kU1FQWg5YM59xZ76xqIJMfOdX759Y8wPcjlJyYGk+ZeJOz+Mwrghddl
yBQTEN4F+7a+pHPTx1yqXu6NolpxTzLsYI9OGotxnZDb8YFVxg/+u84/DxTMnO4NDzKh9ApEN61e
7DiaeHJ93FWjLJI+NRtS39Wy84BPEzZO5/DJtGMyGqlkyIFYHL5iSgYt6M4G6O8aiHuF7cGCn/Mf
7qddxCLlgwKT1v/s9Q+BH/AyunPhNQV+M1Egk8wkKtJMDFLSW47/6V0Myr/ejOT5oN+Iso19KD5v
6rQSnuVzrdInc5vT/j3EiDMFd/HN3WF+K8BfvPCAlFa380x5Mz5QSjpNMc8C0sQGeFqLBqXROg0P
tlTGWqp/EtIKXHFAGsWdME7wETuV6mwQy0G+7ragdBlwB8R2L/JrLjanRNl3/HKv3kGb9Ak4QWyh
LTqhibCDIVy2M2Kk8m57ZlOv5yOD7YoM1sjInmhK/0xsKOv3yHQINAanWhjAdPadf0P0QswonyuI
lhCx/2RssvZEa3iRL5odC2El2v6LQ2TTXDgWAVGhLLe6FgKb4F6G4PkbzotmoeCIQNgAdPLMPdr7
0Qhse3/L2rXVxCZWY2Myvoo+uIEDuysqfI9JX76dKRhcMmviliDZG9GXWFbXm3skGHSAyOJbK1Wt
Id3IG6UhN9ePHfXQ5FyB9btf0HG8HGKXz8PO82JMh9IX33ujzWcu5hG8Lp7V8eDcnMOtYAqoQrGw
emvZjTmiYUD3s2lxW/P75BPxdQ7NBCIwWeFEzI6hbDkMD2tmlA1tZD6yWmXF2DSG/OoZZAupIQW6
kEs+bCJjmz/J8hVv104thT6F47/7H7Vpb6wKhF3DVYQIpbwjVIGPYnNtd+j/9c208Z+8cGVQA8jj
d2HZtgygoBssfbKzCc8gp+/GiI1VCmtW8Z/ubOoGBcwb0fISo3BLTCcgM15PFpAgaZPGk7LetKKi
Cbuigb4B6p94OjbLTKq02cZiDjfdDur6vZ4spfje2NTt/lEoEdMOh8tjZqPjS4RagViMaNfomwXW
KDM8+/qLw0UtEHA9Asay2qQcMsvxllUBBQeEj9zc7M//v5F6HRHYtStzWUQSSA69GuX3uiqtspVT
swsxfkg3TJm0yyRjU9SQr656C3sQOIPey67H9Woyv4U6ak4PkCQ2uWDsoe0AZbcmaKOkAjOm7XLp
Uw6Vql/Is2w57sRnRVnsJbH74g8KP0vxgSgLX8RJrxzZbBQtWX8STJqJlpswCxOWZHEHtzl8Ygv5
VIgjrzy+FVBMJ7mBSXDUwPYsgrhPUEBTSujeyRbTlABK67iXsjjW4PFQa4TXxHcJfISTNfpTay3n
D8FUzlubSnWmy5LdTGnZTFP3Q8JFYDcyFW9/bWJr055qBIr4ieLr/xUu7FmDf2k8dtiudJ7JNw/T
mKWFLCj143HALMIWeS08mO/L9MUiaHZgOJedC0ILX8YOLHRyhCrYDTV0sKKMnNLCeWb/J1jwDiZl
1euKs/QlakFxajDxk61m+x15A42yfYBblezbOwsPowfWlFaMwm4Srndr1a3xQXoV04aByJC03fXU
/uW74/fKjEqfiGjw03CS/OIJiMUhhSG+fl02PD9xv/s8MuWVWm733+MveNtwxfE/BxAma5NB0UIk
EtDTn3FBApxAWX3RrydSAOYcczL41X2VpzY3g957+A5igRtD+a7rSII8+ugnupg/EJ4N5T53eYTK
LUgwGIQ9ywz00NbWlk+rxIwuYUQutfBafihnIkOGyDofLJemKguBSR7YHLh6b8PUSEk34KXREYi2
gDD7Hg8wSvaWQA6sp6itV2+us/sssMR0a2xtbRlh7Ubs7jnMX1hryXzRJdwMi7R22x2HMk2ZGhYs
3jY7Dqgv1dmfgH2NlVuLq2p2xENL/Z04Ya6cvm/ncpk1FVCcFNLZN4+KsrQPUYAYd1M+fhFpFEgl
YbkUlHOxL/sOZDz4vnzMsMtAB6klZK88mky18zxBQmgjwTJ8ALjHpg/nF8zCydJGcb4H3uicHMp0
1wgDBTMCFzIxb8JNYBDqhuZ52bmJZZxug+qVgD9XWaeHzhJoHazfFngoAmfZPf8am78vC35n7LXN
jkKM/22tYQ7n1kJleVejWqJGz8CZg0Crct0P3nI2eTQnJQUkbCpM9JBiYpZVw2n6YvZoTxI4aQEj
JMoQ+SuPj55vV32POy6AasFMq++/2JES6LVE5GqNczy6Ubn04y6j6QfW3TeMnbFn/u6yyAwbo9XD
i+qXr4P3l9RDWaGXjSyOXO4VY+a+Iwbl8CeWs0joeUGrWMwJPKl5ekGppUuzlo1FZ7IdcIXxwbqD
S0Sja/pTHiJ4ubCtGh7eqkXbbZTmHMjJxXCuc7KMI5fHN69wW+Xa+SdzfNVUIYuHTywW5wBsYrsZ
YKH2hkHpTrqbc9f2QYrmaz+gEt/QN2mp2exT1mIuV9VfYir5FcSUryFylDo3rJ8MkgqYO5iFYcK7
32zI+aSLD94nCiy7a8t/TSAu+jdcUvQCFjZOdtNSeZ1svcBtDwxLIyX19XUjEPhBjb/WFSD5xBdH
54NK242fuJW/WR6SDjkK8oV+OhS3zibB5jI8c+JaL1qd10rRpoxAKsjrPxUuB0XON6Zmhn97+8dO
cRwZeoIIxBVi+FGJ0qBvFPKKIds9kDv0koIsoybwDMigWDXGKLJ6CzCMzOaxBIQ5qRQO2llXPip1
asmlIYuJXLsroxWLtN58QPSuwYvd8USWUWxcmjTe47fpwX9ZrSE43eMg0Rtxqs3WLVZHB44du6sF
uv85jQH+w/eppTI0U0GON3fgxESOsRvPauyqPZ8ZjXQd0ZsKOyHgRO5rKEI/W53Lvkm5LT0yN2qu
L/4yDwEaIymKFEggQVJak9FNPjz+f3BSf+C/f/hp9idTauu50mjO2iyP20XJct40eTfmquVDvVfi
YCaTZ58IxtjzcD+If0NSA3Cdani99COJsWiLfD1RePKuCkDVPF+tZPlV/ydv5G//QHkWiKyT26t+
YHxiC6BleJ7uhFWBu4XgSn/LXeG95N4xlRmmirILMrFa5dEeLKSrmB3tEK1snZ6100PFt78zG1g1
JDrnohBF2sXlKHogMeS/RbOgaIxHXq6KEgbFMh0YFhcUER0/FN88sGuM1aXnDMQX0GDBPxtRxWxH
3XVC1S73+H6gOcrdJil7dZ3+Rnk7i8keeMo+/A9HuUkitXFniU2f63Q03mRuAEmML2g6wfzM4w8I
F7P22DgWut7607lYc/OryuOetMcsfyEUz116j+bUK3i/pu+rHNpRt9QM5Nk9r2XTlJtiEtCnargG
5FspFZ/JC98y3TQ/DqwFWCmSBFirmphB03gw2diF0golH5MGNdXK/rZxEhSsB/x4fJNuldc9s+rz
0UlLq45N/JyySC5rpZBqp4TQid1GzMxOiKu3zrE92945w90ZsMhoQ5mZkz9UAs3mJKSh3dfKpNQU
a6xFlm++MLLD+R4o6dBO/3eBdwAa2LoaUzhoTXSctDxTFff27HXU7HO79KkCMD/YIk/NhpKzfGJL
lHwETKjfLtu/QnZHXUlW8lw9tdxvW5LkoDF175OzAGiy41jtMX7jjw4gRAmbWqQY+9+9edMNon3g
+I55ZNo7g96QVNJScRaMPYq7xiLMW17cit9o2J7hhMlgKj49viKLcA3l8oYlTz3Hs8KuXlbGx6+J
JmoHsQYCllRzxRBBZfl7YAabW9SHYxx9kP9VIaemXgcMXM9LwGRzFB9YLbjsOyS8XMFlpZXX7Of6
I7zEyc3K3jbVVTJw4haEh39b0l0kpuRjbbbN7FXaCF4pOG9pOiB2S8UmiD7WlWUOUu+qqjI4tokj
dvnL3EV7deMpZkmKpig4HlUiBGSzrrXduLy3XB9u4gTe4xAHUEzTEHgf2ExNPrl99pbk7Hk9Su2e
QrKnzg9Syvb/fTHB8mDzunVbbNYMcrTsknsJjkzCPmPfGr1BN+BE//S1YFFxuqKQ5KYcg9BZ77pU
wQtocT/+87XYvCMfgs7bIpLRsHMFCCREgt57iYOvuTNGl4oWFL3loc3JhQ/lTV9Y9sPRPR6zGi1O
W4poEReLQN9jvF6MoK/df8mS0Jg4UI8h/vIfwsD5KJirv+OT6w250S3Uc0RyPk5ghOf3PVpWHSHD
1yaSqsX9KaXx5rHpfLarzbKtGkOn3so4Tn2qbpWy/R9oc7zskvPgdBC5yVTLk2KR/SiTrwTgC69T
sUQvj3Z7teqaB+irHZooSj2bAfhg8OgOpNdAdj9hkMyHxXJ8IcMZG+8ppbHcaTrTJljfNIrvX+cF
bwHl3eCBfmjAUq3/bnf91/TEY8yKChcs/MChCO/aPN5Jmw48tYZxWhTok2nV1WqepJFZDo5NjXRD
Xd912Nm8D29OzxTTVs/9aaie7o22gJEJBQAQdJtnR1tHsGyG2GaHlhaEkD5iQi1YA1giIo8QYG+9
qHvdGVohVhvWM4OzUV8c6dVBoVjqR9wUb9+wQqqJfHC26RkHqdVxkxz0jHjT1IVf2XTBIzeKEqvd
cc21Ig3gEhAKlN2UPk5aj7AVqde66kGpjkOhsgMHkp86UcEXcTmYBkydv7YgFzpodRX2GZc7WBD7
8MhsJ8kOhihqR64RZ9qolQU1FPRlEC/ZbYO2N9Km5rEfM53DNqBfsBHADZZP58bA7bkoIFVGVVLn
Ua6TUHjbfu7C6VcSmQEcN1NhN2qj0OClkrLrWHkaWiaElmW0K9koIq/WMe5kSFIf1+U8op1e3wAp
qQ6NCrRggD77chdF4pnNOHOYmOLn019doxkKsrEQVQLPDowXSTg/zEqhDaxcev2Ld785AA8DET2/
8sRhEDq64hU3wSemOsVWnXiEFl7SzJmRVi7u7ojM0vBzljthuFJGexgP2W6yPNHpoea5sydMKkV+
CH9sHDfsnssWHtMGFZ8Jet9yA4ZICw4idT0XMDvuXtnloa1kGy/0e7HdurhlPbeRtTZecSzseA8p
0gp1jYCzSfecnqHm4bhC79rWtmtdNwOIgax3my7l7OrCGUlKFEwwuwSx2/a/dMZ/A1tc3suxD9la
7nh8UlgOrDbSpy6OUqPzxcO5g8vgnYg+LXA6l3C30Cl6iLr6G//SGVnKsHxf6vAdCkZMPmUzTRMN
Lv/pePRhaqUxwxPMaPQTcj9P0XKBazcmEHLxPpNhxuIRR7kkxz/pSsnob8zWDyoanaUbjg9AutIW
fCPBrhK4VjEoXMiGjVbRIcnay0qQurr9w13UlkVPF1L+G9puFEZvzrYhFJhB0B0k8ZsN5/ErV0xl
r+RqEU4WSRguC5y/A1wR+Lupi6obSAQFsHkBuHumtRr7LNLJNLriNOopg0k3g8auxIsRYLv9/Q4/
Ncgpf9vBazs5uHSidSHGdQPivse+hLsTHfdXJKHiwMltyYTADzi+vjc9TslDz4L5XdDKHDn2nW01
BEJ+6NbtIbnuxPdFEFR9VHy8aFImwen6WBlfqKUXqEviXXYRlzqO20EGLrfn0qztYR6q58L6HAEz
dHqMCdHsOYVMOfkoO5F4Kq7d8tWYSdQ69Vh2uyYE3Nj+Rru1BuzjS/1lqpRZ9kAYJioB2EFKNwz5
wCOoV7uG1vTuICWZT9D8JmWyWnmOnlv1hCroaRO1Iu7J++zMGuWgX2+fpWykx5AWT+s01TRq9oBI
j2qQYs7s4OmT/0RRHqRDF0+dZ/vTmkp5kQgPEFKP8UM8k3n1xMnmRNwkzxqg1ZoWjAmTy/kEX4uw
a2MW7tTBXuYEcTM3/0IZfGhwQxoi3muCADXnQkWOSJI28BvuYgI/Tbi7rE4DZheJLxJjJH4DEQGu
rkP2dOocCdwYy5mYpGKJkIc1HQm3M4YXHbt0EfxE9ZY50J2vfbVFADgmzzQLe5YhFy7idz21Fm7o
8h/GkyX4dZtrOigvQVn+r9OKVCz4ID+7ceAcgrbAbUFVAe1xVJ8m89XPmZhPlkRrlTf3I+B9B8ea
OFC0rtaBhZVUBRlBLRQ9+CZbaq45lzChS83P7AkEc5sTgGOIuVpvePaW6m/KRSXtjSKWHuJAkZbk
r/ztUUfbs2H3t8gzIZj7HuuGEJQbBcDKFBnTCE0zU+vgyzzIMYNsX1G5CEfEo1PdCE6vKUYy1FMi
QWPpcdiBGtF5fgQmXqAwheBcCooCev28vk+PZb9xU3uTvyRqXo8AMpxVbjqnrWTL7PSRt4BI382u
t8BTQ6sV56Yuxu2E0ZXUKeohmBg++wxd6fOUvu3P3+5X7GRIHScpLOwvcdDR0h/CiTbYIc8SRaH4
s2FSkbH+91IPtuilbVq1FXWEW3jke+RShUcAYtfYejxdzZY/gPKsf8PZ+yQEIzEqhJ+pzO/VxsY2
9hBfKjswc47cB0xoNF2Up2QcPhA4de7k+NdANCNMOmHvE9BQ8P3gV9g7BeoLaTwMa0Vo+krzL3EK
R/MWgwVN9ppo4EjniUZ4YPTof0JE06TsreakH5Rdylv/rEDUkiKWYBgktFMQ8yMurinElB1D35wy
U3gyatmxcr0uQTEZE+Zipm/+BFbRXswweknf5lXj/1NgX1KVvQ0ljqnaxavnrHvOCvHR9kXUnK5n
6bh09wm++x6aY1Bit4AxwVVm59zjHHi/YP2RcsIX0eKC7iB8kyELTTHSomTOGfKWP6N+dIEa8lHA
NTxlFwHUK7dQuoROxl8aydrXQkVwM9yrISlg9Kn2kgVvI1lCcgNwHH9gbAxkUVQ0+LHuUN1N5smW
uDWKtydB+yHIUwPMb6GrSuuNeQULX1/5jjTn1h18X6Z0wGSyieaQiCN43wF1/GADXO4Qj+3AIUmI
Gh8fil5c9HRWbd2h8sBbqUEWCo6TkJ4zssXDXFPsfr1/77br9zm9nqmkZvz6NjKUdXyYE60uNcai
3ObLxyWCLObUnBH21NS0WnICzwkncKL3TOWO3K5MQXmkpwkbVpTHQw57kyjZsL33AX8xIGLwybeS
kW+8CdNawyAIKtNN/DN5K/4TALN2r0C0yYgrwaUs7P1HtLsL+oBETywpF/HaalIhVxiOFAd/oPUT
MeU2ffkkJ4kjxKYQ2cd0RN35FkbzwIsmmaH5lDdMRfnyL9Zfsn51mb4dyHUc/2neUv09S/78UA89
oF7F0TE6QvCfVwAEzYhbWdfg/fX1EibAa3lbpdTUy159ZGrBxwsMmrLDMHWED8Fz00oqdEeCm4ud
zRidycb2ZqnDH8vQmqLx+vHLvrsI6dO0iWFo/bieREsQbf61rGWsEVrs63pMIJcgYXwDVI9lIAjR
zVMizRdEfdY1B8JSrHX7eaxLYB0Kb6FaDdvHc4n4WL61k77W5196u+Jan5fN5d7HSExO5rzDYIf7
T+HdYg00JvgUtpTiWXo1FXFlETE8dz0oo59+UF0HSPC+LmZGnp4wbI0Vh2DEcY5wLMsdN9riQ5x6
TuCG1G6lDqCZ526PRfrWzDpfyTPi4xEY7vzdBBVMBvbQDCvYzLbHAivdHT2mJDUfFs7wtx1tQhnE
WkOjmcMCg92ju9I/ulfuGXjh6CXKrDNtTTJZ1wwNGHMWjsWZFN0iclOHsEr5COqTlk4OcHJPCPCf
9R5ks7665OErBgqtoAaYkUqnpwvN7Gza/K0eXfBfNz7pryaOoKEVd+OeF2/JTKUXK+nQ0vnph1rO
3xCfmY7WNK2LMNYyiW0Vktn5IOAf4Kow1qwDM0UDJLU4NqC0DZBI3QR8uN5KLzDfUcMMzPqBaH1w
v8CGKe0h7ASOaWGDCoqky702hw6dgcFd7tzkx4kakvf+/Sfpi0Jc6x/FzMJ/Asw2s7bjXT8QirC6
44G5szlrlbXOdC2CdN86pJBe7jBIkzxaAOG9TYlxC8p86y6PEKRBXvqhDavR22xDypYANZ17pQBW
FvD+iOAaM0eD72QJ5xKcD1mV2hwR0kmM0RubUHNEAogmPkTm0DZwXd9DCKcGP/Sq26jiL79azlgO
fUFi1JE8zG6Vya4TfjBblKRD/jgko4pAIJwF7nfAFMlPgPlbcjFewV/RJwpyAFinym79evQac+R+
SRvefQ5yA7oSuFBDt6Et1uWb9FFTHh23n83CpJiBfaGCbrYVII1WIBJlAYQTBXVwnDQUbUqpMLDG
3c2YMZSaU8WD1t4bJHa3ZE7flsqNGjvgcGz2VFE9CW+jNeBcuDL9IJZ2BL/wGTBo+LGCDOi7LfCT
1/5rkj1taBHUfNOH+Uiun6Lp68s+wXVOZscaSfa0MEf17v1mzUjwHyBofkKrDl/ycq5Pmq7yFvrY
X/jEdFjHw+i1eaHhhVlQ9Hkq5p30Nw9R+kknmobNu7sm87Z8vgjl4smKjMmn8bPJBI4VIjytij6i
g3qqOO+CKJ/m2LDByrxnvoJ5r+kWLxzr73hmaQTu5zmb5fYERtk0+/SoGEOSl3T7xiMyr5989VLf
O1tKCzrV34sdEQgJVDoxIXae/ts61VjUG13HDv2tagMoyk+jjgUZdMsiw+78+wKB55sKuFV7w/kC
Q+kN5SSDD9wjL8dZWz3H1ppekuf9ay5Kjie97rcTAz6imvrpP5BWDomjfl6KuPTpesJePR3dPg9I
9Va1f6JLaVGSRYthVcnWZ2bgsJLmg14Q+irvLU2u0XjADZGjoUaMnYH1MYCjD71KrcuROODvj0zk
jogy9JQwzMrkARIPrsovhxsu4Q7/Y25noNcbCogpFd/sM9ir4iQNofqumbgwRKYhg0aD1qFgrf25
gfWH1X7yGQdOX/VkBSghKUwhlDVZ8ggMnxntEU+SIzobFCgpjgMEhJVdY6kcGBGUMtWGrbnC223G
nSrLfv2NxwdRjoyqdB0KBqOUbNMe3F688sRPgjwZ+/+3z9VTXj0+N2qABaaZR2ihXybLTO4AXIth
zbW0Il3Nm6vyYqrz27VhyqTpOj4a7Np3+n23jhbr3TeBmJX68E6HHS5/S5g4diPyy4jE3IRWqFHB
I6Sx3NW5R/TsDkzH4Ov3X7Akh9kjae/qtGNTYUGHfc/BWAM2KEbbsefcU8H8U8rABgpLT8GSxSz2
B2chQWTcY0rm7Rn1dLwMlJiCKHxvGDoQ37f+lMgTL7aejt0lm3DBiR4ZMoFEt9u1VTiPxb2pTxN0
ef8CzhX6iKOQgAxxuHASzIyAbtBNXzbmI1RGJjFqfwXO07ENd2OSeNmppwIDSMzyyH6N8F5YhdpQ
ApmURpGTj7qYkaN3PNtZz6aIEOqsRqSpA9T7NrfDmhOddXK8F3+Eq29ylN5vFZV6WaSxoPxsfrKX
MXxTsXDfJGljy+ZpaSoRrtuZrNP31Yba4kml0fmudm6b0LAxA3R556B03NYxZiklKJ2IhjM+PGwH
BTuazWUfobOZVOhjIk3rsa18CY8tB3OvkkQD4oBrOZ1T+Y1y1pL6xAcQ46XokLNlRa+hNKn1dA3z
CAA3nGconuiICon8E79Vo/c+nc+rSW8dfEt/E6GT13uvPBJgK3Y+K4rN7n+xTRykhO1yGQgilIKT
sD8A2V1mu+cl5fhkDKsCNt49gXWCMr/ABGv+BwtSnYNgRYXZJpg9xjyImBEUfP6BNo9sp9C0TiL9
NphwKW9dSnv0kUqmHMrC2M1nqqj3O5O8KzgQCDJf1EhBC7mXubSK7jMYgXaO27tP+TxQZN0/ehk+
qU379yfPfAC9M3ApVQcaNJDL4688DlQuELnC2MdDeucGdL9dlur8FUQU+ptzFoacgQXylZgzeftD
5CAAi8LEfl5gMVTCLEuSFjg/CP3g2qxAyqVqQwm0MDLKR4ddDcSzcyje3623M9Jf9ZKfeoZTTB3T
yW99PcLXJs3AzwAId7VfupCABqdhf6Ci7bj5AxQKgC54Bev26/xK2BZYe3qWuppUP808k+1X2u/s
TwnA5NkNZMaq4Upi+4yoUJLZJk3qCHVQx/zD4Ll670zvYzWeJCvKFdp63SqRfandIcrDIfpFq1f6
6+4roMmnUgm58WOwtg7+3y96g0Yc1GOmtKq8b5YRnhewfrhgfIqJZ8YrzP1Q3BwzOfB0CWhX4wrc
7LjXBUNjWKQmUIjjmGUjjTFoNnczVHT/KwWxyHZtZEUTLOqLegGskzO8ztsUvfwnpunz7F2inkA8
DvXwqBvx+nM9KytR8aG17m5CrtDczUXB5/q2lorQklQ4SlppRbDWlAxubL/Ow2gpOoO7f5KVZZ4D
Cb8Eu+VBxRI3fxDQUig7zsBAnjOdcGcbdOap8kcMeKdEuzf4Zkyzb2ocYaQtRj+JTYQgA081MQ55
jLt6YQCYGBoUxsku4CcWqsWTac5MHv2d5racV/lbElXZW1ANd/t/YLjr+oDMv/wW1liCbPkH51hq
IiaB4NVg2GkBArYCgb3sMUXVLFMoDU30EQJDDaQGSzJ1CUjhq6Cm1+CpHLiWnlDtuS0M5E16HA5R
YU4KxwZsWqk/JxRvMI0CfPhQqvuvJq8lz+bxrmpgB6nbAU7BTiXjWC9o0jJm1ovw4DQICZVZKC8B
9PyFg2moZN5tyOQPeumqWu1Bomy9S5LvAbLvOIklWhMG+qK+DFJ7KnmqADI0FBSkIBC2bhzMxtiK
NoraUrqRuNKvtqMv4oW45YnAZHJkuZ0hi4Sj2WEd7cSPB4P8Drvi8KzqG68Odg75zP2SJMfSLnWM
8QUVKggNXBSUVyqyCKiq2yYKqi8/ciqpxMBLAW6Di8NwwDnYy4w8M3rpyKpBjT2SMJMnmFHAe+gL
boymwbPMdCCY2MdmGt7Gl4X5R/lwoRu/0L7CjakEKFn0viUa0h22osK2t77sxflBOyZSY8g+q/3D
7OnvFz8StB1B44N+yteHhpidxCLrCZUQhHh7VNnZ0CCyxYecHpcWzINllqVBYWEY/9o7JOIJKKLD
WoaRn0gv+Rr8tq4r3f+ec53/59XQs53vOPEUB3jmnkb2iealupVJIct0IOCgFQW7SKXBa8+q026K
pa7gFwAU6jMwlDQXDeRsabYn0UbKMyvJWoeptrycm/n42VQyRGF2Ka5UnzbPyXhWDM/JiEChjU82
+0hPG+DxH5GJXccXKuBQaNBEbq7fH4z7oATRFpyhrr6SWraieTRJiTJHXBwg/Wquvd/cHTiBPGu6
HaKO75TUhlvmk/93G/sJtWCVDVQ/FIhEOzKNa7IPZEgKwhzprKO6mdIlqxno5YIpXDFntP4P2uBa
TYAKV2gayxU79uZaCwtq49T5V32fJ2+Pd8dceeCJa315wHN0PEtRMpGA0Z6tnsZVlRaYeLzFNAk3
yxACJ8GKzABePm08NP2jYx9KIVWd97Va+FdS9JO5ZUi1yJyoRY3pKCxNQHOk67RAajBucUWVKQWg
0oOszCkNdHBWeGQ/vPobxZNm2mzl+0ERZWrD8sgVbcVx53SHjE620NxBwohfD/0QIuEAWBoI37+n
Vzbp3Zr1hMPjiKWJ1aBmeZegV/Xq8htdMSHqc72gXjwBpXKtxWWF39Kbg/UplPjxGmBjL0NMQBG0
0MU4iXgTQ+BDAFBny8KGl9wEeD0XE+BvKWBO2GKMBnD1oTaOyOInsKQuikHC/zlovPeXW4Gia2PR
X83jnwgftbPRjbOAt2LeSv9dTQ0mf7wMPgFQdH62pCBwJ7OziMA8GHkQ4yrT06bSnmH1IYX5Ghjz
r0WfvkmBiYTTpkir4oBBpwZ75Mx8fbmiDUBf1wQloeB5hb09UjHIL2tsvAU7l9fDkEGvIaQYFGMM
6+F8hFMxZKtiO/HRlQjaFQ7vfPUghRJ2b7qexKBzSvf6jJ7xKEk6aU8u1EZFe3nAS5d9Er2is6tK
nEnkiV0m8WGLrZwKTPa4qBVNoonkzwHTHeEUzv1A/isXHGZrqE1esZGzcwFJKy2g9DIEQNnbhLkL
sVaaAWDA9Ltwu5n5gK0nP2x3Fu/3yYBH+/FIJXDtFub7sibDcvyAgRVD9gPLFZiCoVBf5eIBuBkn
RdBEXtLPLq9G25A8VoxuYFKB2vBxbtK1Tun+9dnQEW5WO3p4bLx1dI+ynKjITUr9OjSmUsoE/omR
ZWrZsojTwmAYrfC/z0UcBFrWKYJs/34WvN3UPArDI53hmH8Pg0c+l8sykwMM1KCRHAjfXtbrgLy5
DJ5s05memyj/24ArGNsYkwDRBRIJyMFnsOGNASYo22AN1wTq9aG0XHjgdjDIGDpS8mfW3hbueNAP
KI4D2pr8R2JKvUaqNHz4wGzw5A9vhYzjkn2vIaoygmeuVdTpcIniOoATwJhq75kK7Uxd1wJpGGWQ
9644xh7m/8pD3tdsoMqIurliRJIhx9ZfbmqK63ORnZzfUcwznNTrco4hPZpLA8eVrHXm61/sJIg3
TMQtAihuwVIexWSoqBDpuSCf9R7B2rqTLJki154v7nZLPWrRrYl9+nCIVXMLDJvOqoUqoV7IFS1P
CJUyuxM8p43TlnFVI6GpRIPspUl1MIOjWDoW7gzWoJ6QQ5t9tbaFXjGHv129oxfGSv5u/Yk8JjIR
PNJoquShQtT6RHk5IYyZRhBYAnnCBYAUh8fUBhCIsvUNF0C+Vr3dIDikqon4A61JsyZsFActFyPM
hbNdKyh2K0XXmJ6iIrjvw0Q+Ng0EgXHdl7pgXhAME6DXE9LIDiZOZrUTlmpIiwsOeZnpmfxNjeZX
UgEcx6OELRg0/BLnETE2v7VZr7Ij+iVBkjgR0k4yNzcpaPq2OxsG4Cuf+IxcCBwPP6UqyQ1kJCwi
+XpoJ4UwInoTzJ0fl3ArROu+/lFsWw0tH64jq66kV/iOVBU0L0tkC8UueSIxYoJYMujoqno0G56r
my+ra1k1MsKkRKzrC1puTPIqkpxpkApfp6cHEYVzf8aBFjqF0a/5YGM34oSau0BGImxupfrVCes7
gYIxuZrAFtCnbS4Y4gpKJkOvIRwwbgfPLbDEY6DhRQ339ZGafg7l2Y/F3oOzv3Y/MUpyZVngw1J6
/qEtosU44vhVxNcFQdz6nFXnurIJ7H74+svVYc7x9zjaeTGMnZFjUwX6g2xJ4RqzL+YTsOwZvgDK
pyDprPpMLQiGEYs/AMRrBqz4KOvIgYQI9XkBoiXZDc1dK7Z/wImVT2MDVjza5TEH+wLovjQrtuca
XFlRInTEBzie/unCSq+UZ7+7ipwh/xs5+cCaqJCK/p1pEeAQ8IG/yDnfLt6IV+SMAOfVBqVmWlvf
oWAKSoE5xhRieQITAuDTDNdrbwYY/41Yo+njx3htXLI30k3jxFbbNOUBqqbNq1+mBcH2mFU7uHtP
1OMsjYlFzEoUR8KgvcmUOAo8Jb0kJiAkQBTE9zO9ox5E9UXuwyJ7ojfC2uH+EMUDJfHEPu0Gx2Jk
eOO2tbLj8X34818i7FTs31TAHPqYZWwj6sfugCDGZwR8wB/ELYFMjcRZycMfHigg+wLaHci1Zr+i
tmEUYzSOEuDufMjTvo9L/dRLJzJv6cfMxoTbMHFT/q5JwguUkFEqup8wU4lbey5BF3vEdseCk4PP
RGCgEaDF3uv8o3ilyJRpP72p6isahyjrf6YsNokpqdFTFaxL1bjHv6k2bIt4PR/jSBklc1nqM1Uk
PyABagZA+eV8BgEnlBHYQqW/Sjrj1ulB89BgB9u8GUHoUkaOLtxcGTrRLSyGfZ4KjoRWgCQ8BmDN
cjKzNxa6OFbwdDX1jaK/Sabk1Z/yZAfaa7y5khkqq4mJlICgpoPzLPn19nZKdUnkgGkX7bTPRmpq
nkYCUdm654X2sz6KeSUtxsqEvbus3ffsYwkqx/t8XSWedR4vy2sFU9cacex1c+XLx3ooY1iSAAg+
h2BBRKRZW+oD9hvtBpfEKkhlYH3jNUnhOMHODR62nFNG2n/FHiobUwsohr2aXiErRGcB+Juv1aYK
xr5A3xkO+0FCjghHzuCoKyCVqoDNpneVIjmKYnXuxEMjsooTUfqTn5b38iYbr7oq8Xe620mrlna7
zWodn+34ocTqlDkFy5HZvW5dfD9kLj62CW/Cp+120FGLdnpPzgeRHasWeIgUUEMJYpWILwsy2JkF
anHSlKGPxMTKgFB+gr20jQ30f1jln/4P9a1aAopi47dBQVbLkkcWui+/gfmFxdOK6WCehi3zP75R
eOALpOFciFvDHjVj+NW+vxfmiaGA0VNqtn82rdiw1huR1P+rXrNl9eTn32pv8VsP+O5PVi8vD+0j
MkzgeHRIvD+ADAZ+QvCPGT8zr+MmHhtLtaGGmsOkV6xO+4tMC4Dav20Wedj5H32v+uay1vMftHP0
tLw1Xn1Uk7DdpTbZBN06zKFLmzL+uprUTULW2Q67ParnCPvpi3zRl2ZWlBN0hcHU1dpfyzP0e0pN
k3RQXZRHNuERRJ/VKaAr2qIo/HmQdTF+FJ08PhJM9ENwD0+rNyEty/Zu3Bg7NO9BBUMOkalnJOlK
Vhll3Ji9upW0Hb1m3vdiDEY1X/7p1A0Mjtdj1jNLm8OkH+DllaM/EH7mekQ9n3ra5UYiQ297QENg
jjOu7D0eWYQj4k/yerdZpaXHpDM+f14U2ZAtiE9IA0ROoTF5MeINAavtBgFEP3CRW+nDLhT0aQir
5bzivanm/SknCsZAsLe0aHByyUVcmW+2XNj8mORZcIA4AYDxOgqNrx63PTWVEwDn//aQk6DU/5BC
12OcS3JwhetDhfhVGQmsQsjlfrgxNnDaHBxDggsNxsUa5mFsmeOAii/2wTy2NeiGFt2788Yb/PXq
y2VszusBn82LEL4F3QMr7ZFxBlkcnUgK8c6sRUGF6eL6t4K8AeGSQTtF8/pvvDyq7AmbOs5Q+n/k
k8KX+oRNF8XPJd8yHyzh3v7oxrugT1IA1QIZWJ59dQ2ijCTWoF1twZF03IdmeLFKuKsbceIvEqKo
6KHchLqoSvAwcoYVk7FFAKf1Yt/EdraPEiN+L0B2xyI25NmeXVeooNMpen3i0C2E4RqRlg/e/aq9
OKUnS08KpEm1dtDkCQSuO879MdWD4mcpzsGlNf0DRgSmQ60nzKDl99F5JYqoWreRnnBOZMs2N7GC
3hDGPIVngxeh8OjuISeQzS14uBTXm0NXM5zDHbEVB7j3zqmVKFJk9rJfems5n9BLqIAhVkjJXUV2
BXOkFo/NzMxzhLVHGsv0l3YFINR1B49YBbVaYvDGVvBllCE7Ash0FVG8KCBJi8EhRfEyTMaKxVig
+sKC9ErjYEfUzMUwtlg2PrStyIckq7+1RpBNJP8lXX2eih3yZlexEWV5zXCpbLECK2SwFQp7rHWb
DLBaDUqB+xEvHRrL7wCQcob/NTXtLtLrDxm6AYb5O6Ak6wFz6og3wpOWKbHnz8DUGFlKqtUCumpm
kL7v0MztetQ2up7C32U0Z2ewWAKW5Q5fFVZjnO8BiAp3fqD5g+VBZAh88tITYlPIyKH0On5kf0Lk
u89xaVrQ4Zy1fPSmaf3T4wV97T0vhgmG5WY33DutcXThDYhqYKcUPKZFiF2FmgYd6kMxAlZvGlO3
C5y9hqTWonWj66YrJbhGe7eiEVyiGxjdvEyEbXCgGtF/KROjYWC82bcIfc6GKKzxX/I48tM9C0et
U47NFghWpjifNnBd0w7wLP0kvm5rexEAMdKED+6/h2PDlaSe01gz3Msy4lqOpGd6bn6eE/XMw6uE
yR0xt+bdxX4L/ykcr9D7Tymls0wya76i6SmeKLpE1KpLJTLmdNdpMWyx23hAJHgD5e01780C1rv3
wmHunahSWqno3Ec1o/SGSrAAeJp1g86+hNckW+nnN+lg9AuZJFT0jUZrQGoOqtUpidcs8s5iKXow
gYKmnf+4s70hrgg/ZqrCy13bItPth6W7M/q2/0b8mi5LRAzTPVi72zCgpp7ojsfXeA5oix/dQhc8
v8gVr0Jiy/uzFynJFHK02lIPXiSU2mnEQDprs2qa5Uepbo2dpytEEJHM9EJEd7BH/CtvL9l6k94x
nSmn0hOoSatxmYWkDJGky9svddweqp7pDGQGgn9NgoNDRAOyhClFUpCZKXBJbAnQnf8WGTSs9Gff
EfBl5YQX5eV9tibgL/uMxeSJ4Qr7sZ1KT1eFpB4im9M1iZe/2ec81xPfSYwInfgo4sDaIvH/JFXF
5guEBGCtRuHzYm2QOnhpzg5QDfkAiWJmydzlUc+32NceoLeMR56eRhsDA+wU5BCdlyLQsAGSVszI
4bv5Tvv8VXGZt13gIccbvOpM6L3y6Ygol4ENJ8yqvIhhYsL9T/XeO15DAeba14WlHy1prvi2fp5U
uzzsIRHiKKcle/HokheDHN+9WBsrce55GcDC8OLry45BZW/pmhUiSXS5jt3kwS43SQbfr5+VOa7b
/eyIzbQB0t2pY24GFnxTZfG2HkdC5LNTJA2OAh7jl1dEGlytE1duOa6sHkAzJR0X/4fD1k/o7AK/
6Z3yjZuDvfFMcxm1q2EYY0l9lsKPuovzJrP03D0NfcQtcH7VFX+mBjJeeXzenT2TMnRkZ3q+xWtk
p/HA3nU4eZxU3aSXc8oaMIXTVh5KsUTNjgSx48Z6vXVd/tADgP294UDNjjOzS1EhTG+aqpfBheVx
frDzFbS7Kb8b52aZHjz2ZWJGlbggJkQS6Q/CQxWQtwcA4WeDNDu8HnHoKwtME/B9Sv6vMxJf50rP
EgdCBOyYkPbtlOOE/tPgtu1WCnKEx9cFeCkS0kmM8t3sSsGbS5EAFtCCp/gjfeSJTYBE6z8b5BPy
obpu+OOjJZgX/RooW+6PDVwdahP2pmm2CawaxffQWUasuSfiCPHIUW9azttzTqoG42LddMi7GgA1
T7ckPUwpRtqLowR4I9YnATjs7Yo3kRif7E5gKdSN2tATT4/qwCc5hm11qHRsNoBh1ORBSWUDVN7x
YXX0klzy2Qn7TFVazZ/t3PIjrYxyDVwEWrQtPvp3Qp9ILlKOrNnd/7PP0zC1DUoFlceJyED1GGQW
z9/WkJ1qIYtECnI7SqAUsBNNJhrZGGqMLhgiWDUU70FHhxpTsz5MeNiBVC8Jmlib5bSZl+QwZLDN
KQvSFdFg6/WBKPIeR02i1jLasqvjFkDFL37YqgDLghbaEiODqtNPLPW4omtQxSLzEgsgABKG3rAn
DF139S9848u/BND3l9sTwD66OItgZM4Csf8bSWpjjlTJwtcjNVBi/5jIe6RiXjuAd1PlIef5h8BW
qjg6lFCbB2HQnHF0h+8BU7jNhqt06lK9ElCotEGQgZ1rjKju8TQWILnASA+OvPSRQ2vyy9EuQpBf
LoEuMHgkdrH3Ii0YKVqqh1eDKH6iZLOt/pKTQmFjBVnOiMfHlImo2WsbfBp+mVqu2UhmMiQn/xFc
rKqXNYmBXgtCmw8WrfYxts3oY6vNSJKHxNw0XnqnVDIOoFod0aFZsLnwr6qp5NNnu9aKKmBqrrmn
tDFVqavO/1+KJ3li0L/+pxBO1wS4D6fzpE+kynPrMXYjh3/Pg/70G2InJ1SA5R35DTBtvORgrL+I
NGGq+EXBA0Ydyta9LZygDsJqSiZzwfXOpj38NVHP6yKeZQsbaUkl9bPokVBuGMNJbFqvWBwD8I1u
hN3mUFEnU9LpZkR5/QOuqz1Lqab0Wh7tljdkhXKHQKPYr3IttcWVYp3Hf06ddFrzqSGpQ1NiavwB
FWpPeDgb60aqbUNLZ4nHZA6aA9rGu/Miycqfw+MKuTjE1lBjT/XJQcZibs/v7CT2jkJub66OToXQ
59RK+JzFVRur2oy09gF7+MkhSdXo4KP201M+J0Yb3Qm12emctzMGhIVcVDPwU7mSpPY0KB/nMU7L
Z+7gSBBY1sTcpuxUzc/aST+oMPAiercr4FYvEFZDOh+o0SFN9WTBaAmmKabiBlEob4ATehrejkym
YXg+gRg9pcDRaAHsUzMaAb2Qce7SAbPQ+0C/3hp9gmnn6AGsoiaOWIz/EhvvPx1TqNMEhGrbpjYF
VEnl3R20Y7qcT8bb5t4qAa8rBpKBo4ZqsKqMYDh6bR8ey4eMyJgBCmIrQHIjrWXZG9k1650Z9xWH
s5UOjWDizs1PQ0p5c11NejJKA3Fa2x4HkS/UgPeCStt2wZC6jz0rGfvBpaaVUkZA/c35Fn0tsxm3
8IdezM8Q37t9X69x/x1Ew/PORbBF+045OWNZezsXRY6VncU2q1CCr6DKgSfur9fFQ/aJCk4RdWTG
Kvkv8lsgfGAG25XuYDmIMCDe0ZTh6+y/fm7hBwjHCq92cVJzzU+4dSUQ8/5qnT3BfAcoLuU3dZco
jAzyOCz5YxKGRpvFna6BY0wh+PpoapTtVVDQOlOkGRpauuqyyBE+bl8Tv48yKwCeg4ajZHcgfMHs
9c9qL4LTFszZkaYMiv3WbjEvC7dUD/o8EA2KLKou8YNXM09lQqaiz8WlPX2g+w8eYge1cfV+A717
ExbXecjYVES6Nz011mfUsqaxMbpg/fnUoSHYZK91JfbJJuzxrGPDwQYYeQIgHZvdbt0iqkpDK398
XHe1/D6Iptl1sbR4cmADPxVMGL95K10RyEYACJG8a/7sHz+1RUZWBWPD5sDEqvc4J9O3VP1rTbuX
5HcbMxsR5IYIrCNhsibpgcBB6SdXgBthNmZIc7aGIwFIldrcdp/zvA6Nd2T6OKelb4vtD07UIjTP
/Go/Wxjix1S4iEVPBpUbIROMZHV3o9poDLtXZ2afD70DrXoRL+0DMUpKH5a+iO19FA6eGe5zLkbX
GVkKMWHEwL8itUpZrdTkBTZU6cKe5DJ0IyH4yyVY7aw0U3d0RJCoQ7+0ixZZU0BbPsR355OVcihZ
MILlrrZNlyJg8Uns+Knn3x+z+3VtQ109qXLKCgKyquaL/pW60lw+VRvEIgnwRwjIpjhN6Buq96Yz
gN2Eaa2nlrnZqYLjWqET+11c1sUOEQdoI4+QTgsd8u84W2lJDjXxYKX5l/wEbOXg0Neb6nw35t87
nTZgXtDXvAKP7UY4Y8FZV4J0410+AbFa3ExY5nm6yw282SSh6FYfCScVw7xywShi1nMzarKZM+8x
fr01XrQ6P+5Czs/ULaaNQ0g2mXppQUtDXEG1flUsHIYkZ4tHgpO8N5miwW/Jth6Xhi7m+5wvq6gL
kmOYhDlIzw83pv9ifNUjgf457FSw5SR0t+7TBA9vG44aARUzNYZoUXUOBow5lzGey2ZJI+5ScXhz
RCL21+GfEF/GxM0+AGpFqVkkfRGrrqiEVq6cB8Ep8ossP+aKJmSEsIMF+7LU1o0XSXJL1QNs/iGD
hOxjolId5ZhC/KShikZs/8Cj4OqRujWKfD4mzIHehgwvQ7IQewwk1G33eYH+czUpjU4ga8gn2P8o
foVL24LHKJk0jNrwqVHcQYvJaeK+h8uREMKwpPPCl43xSCWceezE6EGiQNhTwD7+n+0/Uq6caWBr
lEqMmTSVA4x6tNvQ/UwG+WIlhHlTmlawZGLSx6xO7nCj0oviw5DL1YH5RHpWfZN/95TxFQeJm58l
AisVu2EdNvv4LHx9L1J6g7FH1TYRspfrBY6M/Hmmzv3sOpVFZVpNpUrQdCHmhwd3EruI3f/8Knvf
NSMI/MsADb2Iv3g+1kkYUs3WCIxDTtS6T1cHnCydf243XPh9z9F7UnHbQn5okQHC8vURBnh8tWIt
gx73NZ7EVyVMy/GoWGPy97xZd2/zAUvHhp+I26DyFMdxwbjUPz7JV7326+hkhtaYOxesnU3LCIct
sQTbc4momwzpOUF8bb609VQUHIXijw1NvZnDoTOZ7INzlFLNFscTLXzTILE2+Fv/p67Cp4mex/Fa
nbW/4zObi1V2ojGsPMSjO1kjHdAsmniwT69BzSU74tvnTgCg9VoIvTC7AdMTY7VsRLhNXZTpqaA1
t2b8rrIe9vWoQWYpBxvudk+sOm497/5bB1srjqfIxwxRK5nsySYeb1Nbmqbv/8JupDzBfPTdrWYP
ZSEDMdqQoORk/7caduE7g/DwInEbDs+beBAMKlLAN+f/yV2lzd5NDbtnl7K8vc0GQROyVXkgVVaJ
LFBumwmGj3gwJZGFI07JHjh/1YtBlqFkSdZatkXIOnVXhAA/cxSRjY+06L1Eueug+uWZqPHLIXdX
XwOLZ5BYMv6c7X4i/LfWi8SJHTEu5pnCj+OH64E2i5ZJT0jUWTvikmEP45zAhyGt/KVDS4SMMHWt
4cy5Kc/hDh+VFD7kxqRol3f2r2FV0ma/2dberpjXr+UzRsmtlfNxzi5a+DDGoHdPTHc7BuK1DzZu
IU5xlCaXRR8m8dK1wsrwiTBGZJayeyH//betmyMiT0LT76jAPedJyR3R/hqv/jtwgVAlVa5Pge7q
Bjim/4DxPTF2E/hDG7Gq1bPdS08X1c0JNdd/mxuv2alj+ZIl14Kn6GWFOLMY4WP9FhIP5wXEUqMc
DCHr4F3iN6a9v59pzmPX2zY74pwNkK6sLhQT7uj9Y99dil/ns+2TEUJ93n3FTTpHDWOFuyQQo4YZ
qVjQT0WWzAfK3R7/qqb5Ko9T2V9D5mkYpujf2hfl/4nFk2pZLXyINfweh0lLprFfVJg0aFJQyvxc
vr59lLdo0Di7UPKEMVWRNy2IREsrYX3XiMsp/FdftK3ey31B/IITNHAsuNu8ARNxoLXIvS4kyGld
sqDgHnbrQ39XVFV82E875BT0UNRYdGcYiggQs2ozmzv2LNAZLcPezHa3yZuz7JuCC/S2gLUrkr6G
5sdFMqo+EmyDNIjQ1djt/qF9jlS5eHTa2U2+1YiFYVNw75ei//vqjUU95d2OHnnDQ3NDvPoXGyOc
C4TM/CE16EgdcNMceTuGObRyWdhSXvDm3x1zKavKZy8CAfs6GtlaGFMEd9y+EGrwRSxCvpcVGNpm
b/FPT3al0xBt1wnF646h1YzcbeSi0Olz35w5f+lIJZk9MIbD6EBI37u2s0Cr917Tm9j3LWJaA5VA
yrkeiignbqnjeVgccOi7Hm7Qn+C95b9D+AkQe0vzNLvOv2GBlJNHF2ORQ2cYz0Rsd2cZkgvRW4nZ
hr+9trKcMg4PHC+fJq9cXFsu1X0r3rGEXmTMWxJDMyQAGN/MOR2t+wGB+0zrAGsMj5H9v62YNW/i
5UjVK0iZ1lSjVAgYbcHUc2vG/WKg2cRwuh6RpuALW2gt3vCVE7hD+WUPVFtoHzHGETeCSSV1X/i1
Q2riCQraSQUIcAYa/hBoznMmxlhzvulGhpfeJuMSuQTY/i8iIoopjPQn1pcy5jive0qULGB9HjUM
2M7lWYN9OptbTXjWdJL6g3yu+j6VrRisDl3sJ2w5IrB8fo96XordcX3MWou50POSdxt8aVNZvaSB
zpc3S7MTvZAXhUt9t3L40mNLsaTx2DRKnIug2+DjP0mDZ+kCqr7wX3SORuMFLYcfdFEB26a3snkb
O22PTXythhe1N4pocQkESijCuU2VcxDV2CtsS7FLhSHrLst9bpYB2kt4Ng18UISFH4W/ouUZMgsN
CgSOdoQb5Ee9M7+WW31lgMCenGMzgO+0nNPIq9h5dQ5HeqdwxRickhDyEQSR3b/1L53kWK5KRevH
duDDNaUwrufUZrZ0MZgsvS53zC7i64lmkKU/ylkF4Xgf7Lei8+IYC4RjBnDSVy3PG26cHeW0eY4M
r7gGDUA4MJfq8yBdmEpO+ekIiBbm9/ISNo0IkD3gSQWxXOl1vPCVe2NwYPAXxlZ/EBhnVVl1Iidl
UCFHAtbptyh5jIPTXyzcLADCnzFA/d4HoVrteA6Aokx3WfIWo4NaCLXiqHE4ff5CIJzdNePj+gEk
wB2SRsiqIoD9GCf1SCZ6YKr9DllNSyFqDO7+qwrenAi+NVO8W7NusujlBAn9+pcLsEemLLEjG6Sb
tLVMm06mb6HH3qVNDIkIO9/qe/6uITGehNhOIk1Boap2x0l9FSP4x/78n4DoryYr7Qty7X4DgiLX
CIxJ6b55riHtuOKAkcrlDODkz3UJg/MrLubhhUckcRys3W3AAh7m2pluuoZ0BKeywFvaEkepa1L2
1PI0rXVhIwUV6epBmXZ7cYfJYihUX+pa+d7v3t/uVzKKf8nWfoULj64ysmpn8HEX8pJzr2bHErTD
tNJt3SMXvus60lj34UVRNhblt2inlRM7Kim020m2yuEDHR4yz3yZlwqHW1VUUaBL3krhOX8aVr4M
8+sxFgGqsbGm8PAafEq/Zvd8kJjBkVuVKNwMU9hbGlixO4+hlSnVP46NXD+The762qRT8Yt6rchW
L+RUCvi3Y5cXdRHIONMQNeckPK6JDAfFLCo0SmQgbg25YE1DXwU/0gyq/dtM1kCW5/UWWfuesD6h
aWxv7CXgfQzb8czvvQdEpHa0TLwGBYvbtGbxyJxANgSJEm3ehVY31ZBxH+OtJ+Y9VYIP31+CDZxG
N90SKaFKH8Vm0SjJVg2jvvAyLQgcyxSxdEecKP1S1LmkACGyhYl/BAGZL4NYFfid1N4dAuboHisE
uuiPbYdp03dYYufiWgKU1m8+HbOQE4hkat3s8OFfz9eEze0xy8rVo1Mq5B20PmLgRUgGpBrHRHur
gUTDrP15loVUjC7C3QliOqwS38HJh4dkQguAD3Na292pd76nc0i4QR+yfffzVg4E+iJ6LV0/dKEC
FT8TqB9xuf+lgWIrqxoW+k0ZqVwlSllFVHT8fSmODLrA0H7pdid0QibomLXmU/qUg+bsuIVn+k4K
fj/j3om7fJhNJBhwS6zH+1mWmlaUwIth2dBNnNUft6EvExI6FxDOO/efjqw7h5DXHZYZPaUSvbiE
CS451urJiMe8mXYWrV5QL0v1RwUtv4muagsUqXs1uyDM2eD5ddwqmqtGxDL7MBds0TK6FaCyEnKS
KsCOyn/qJhRjbJHvrLvOoUNK6RrFIGRA20ayHmyYS73DS+PaBqw2o5Ycbf8Bsvy6vO2GniuWMOIf
N3pesClZvFvKzULT9rUy2KJ45fYvcdCHYPXTFOVmiqLY7HfVreK7JqIXY/xcxn3qd1QwB2FU8PtF
QgVZ6CAFZTalaN8oYm3w3ceLOQLLQdQ1YRl1i0Hye8pmsSLaAS/ezQbRRrdO4svZ16yLYCSXixyG
dzscFEfCNdMteVgm1RRRQOrMLEx22ZmsjjTiUYkODbpnGzAkBVSItwyR2zFUXWxZCN+rzToRmlmn
wxL9NGdwZ9VrZCrqdvwk7oGNka13SvutqetbqeP0mUyTjX9ncGQVRIBCPsd8Y+apXUIKTpmkULGS
Vh9DwE+dY1L1ypghAhFwzO2/SDCP/2fmx3VqmQWMQ+qnzPsXYymIandHIEuBKx0ZNJxJvLE2CLyR
YvJjTy98QFDULAvebEI1yst6QFxFHHHyljPSReJboKYjBn8Ebao6wzQQDQiH1mfY+Vy6ZP8XJaxA
0ja9ARkZjyqQ4//Tw5WtiVgB8QxL/UMa78fhUXD1Ur1o8AumXUYQtOERHyPkXzgpP0h3KGwNIfdq
p8Jx9hLcVBSQdTVKPqNEmPL818bKWs0qfwOR8B/wnt3dYhay4MZFFnCm/diYQlqCENyn4rk2xmRq
+S95SOTEMx89YYc5Dx2T1lN3y2vLf6EWvn4OFaaQU16bZUeLO3i+5SbbHS0rx3Pzak24qboVIMNk
hMu8kgR6qhZegF5f5i6ZUDpGYeph5XGD1KCVYbft/KKegzGLG5BBTdCBi2Tl6DbfNZ/PYaYF99MH
P//ZlJVdkDRROYQWZRKGWQYOl/Aqyk7g2mBUmCtQrwOLNclmZ2p1QdOKn0cpIVkQ+ETPYdcq64/o
Wg3GUVZp6vlO2lfp55RW6mzT4AkTeNEPtWDd8RkOxA9WRjSgbq1mxs+bEnPkzxYLbKWpZUZMU2+F
Q+OeDsWB9Pol21Z62XGN64yOUCOWML3E3oahHDNVJlalPOEWTLFdsPz+jghLpnqnKskigcVNC72Z
Bqxwq8UDZbeC+6gYsHYQMpVac5WHFeNAFzYinckaejJRb8+WKItiq1/Yxi1TZA03RYRI3CJtR2zh
afcKwa3uzeAmuH6Vs0bjsLtFpQtuEhdyaNLx/A41aSR9QIZwOgFP+jOINLsEICel/MdV38gH11LH
gu9JKNdpfqn8XP2YD3qmg6WUSHg2H264W9vJ3/fh+GClyRrHS797U3lUbjjK//vttuE1T1el+JgW
nZ2B6ae/KUNjFr/O+9UMof/D3wNfX2PKarjMW1RSWe0e/gxyi3eXhlGzqrMCpYFYzlJHCSzjv044
3d5S3GIryYauMsXKuebSWc0Zl/EnBkbOILlnQ+36HNtxzPQSB1wgyAYRcun82ZrQ6k4VgWsu8qjD
Z90XW+X6JLU7RnMTFRFdwXFyeycwofJfV3bljS6IJH9x8gcHl0243e6NLxrpqeCwofxEMqjzZurY
/99OaQvPkoRFVZ5mA9XewE0zRoBsEeU7WUDdqKN5RkSHbMHV3U56NgBhfU4GtzBNjKb8+Z7YQAor
Hx5X414B24S5fqf1EMUAlsy62tyHR0bm+TZlx0M/TDH1IQNdYocLWJ1fzqgHyyl8UXCjZukOHUGE
DSgQ6tC2bPmwzUggDDfq0kCE5JY+++uf0qWGMsk7dGdmvnC8KufbZkb6OyzMlETNP4dD2UBQ/g73
yDUZDiPah4onXUOy6X6+PZJ7N9FNN7Rfeimu/mw/ME+CuuLTOAXqZfy3XoJcQNBusQOSuF2//AlO
lcKMHowt3QGhzEY29fTuf1+TcKga1vgOh68V/QH+3wd4v1wvmgB9qAQoDa7WqF0xS4efUA1slU7R
7gYyzbfgyD23anOsclV5p+uhRPPfJvGCpwsI/mRSWVzptebbQ2eWgmBLmulXdosDDQhl+bM7jC57
z3+XKIMi3Y0u1eP22Qt2yIhQmiCKQWqeD0dfbMwDNvk2+PkW0CV3nQUvSI3k7r6c7Ir+EfdoVl3V
9Q61rVlMMkMLjk/TFwOBXmMr0lHAiipny6U9vvxAWbYYBeHH7gpklHOZq2dp87g5YS6JwHzTpSFm
gACMltFlRb/U9yxen1JgWl9jJo7WkTmvopVsJ1CpfreUFRl76dq/7riHrkjUI2IH1rcEVSG2oqeQ
ENe76Ku+OJSv+enRPVxQAqt3RvwC0hz0j0zYReEzvpKJ+TNzgCND0J6UCZUNng9V/KpOyjQ3SJ5k
N7oAm10TuKcPndazFfIspq/iwro+Xyy8jKOZM7Kv0EBhi/Qr0YqVg8u51MLuOtv5QLqQTlQK5XwN
2I66YfZS4gU0n6vb5vg1ep41Jl0R0XnaDKdH5hksFSyITsX70sLftFTAfoOKvb5fbRL27nfI2JBA
e2+f+e3RVuzm2KvGZQEzypMjHXnM3+/MiOmddh62I7wx0hoTOWjL6Es7PaeNU50Own6tVAmqwJ1P
wWyfw12LQnSmNfP1grkeJ2PIHx3us9BTFsnUcEF+AfDXyQmxRH+TTi47RQZId/OJo6123owQL4f9
lawdWr5V6Hsi43A3z/nD4mBmxc/HV8Anp6KYjgrR180H0AugbN2XBsX0GXR7eJm30owQYbWpRjqI
j6sSzZUjYF/llIfEYS2o1kD5XHJ/aXHRgX6zBlZahtWgzhF4k0NBGM2RQOM2oHMZg4CxvKEgwvHO
YmSz1l5MJL/72eQOI6Z2c7JVVUQtTcSEvqqpe3/ekWfsUBwH2NOKFSjygBmpb89gPOkF3gmMV3L9
x3X9DQAXMkKQdBA5lFBp46CuxpGWFga6cfyJMxD+TkAcjV3OvrlTHFldszqJ9vul5FE2yTwj0s2O
jsoVIej6VG7CSZ+UdmIUiaaUeUtDbFkJkQUd2NHIlPlmjahotssVaR1mR8YIG+85EQ0LOMGy1JXC
OW1ccHhoVSWdzCBgL2kkVQANK4iojn00T4QTiIu1M5jubXvfv8d1p/8N3bq/QzA+vILx/SWTs3g2
DY76cNHJ7HaYiN+G4JWi4sbP0X1MsLF5vwB8WzIJaiQmCxvvEh5pSPfRZtQ9XmggNjJuoJOF6LMT
03TCmJ6lXnNuJ+Hq/LnK5gjCjO57Z92iZwwISKtnw2JaBn23Gju3AXE+4ORSKtjGzes1TzzCuKEQ
b+tQJVgQ8ViDxSdquQ2fnZN0AiepU3D5WgFNpgCnbqCJMPmiyL1CpK0jgJ0Mut0g2Wurx+V2AJ/A
PIJhgcJpXmV9YtTzCoay3c5zyaSirE5ztkTwjEdU0JTsj1mHK0MnDjFs55ap6ZPXlGtuv2p5UAzV
/KAIqqdY78kOwmfFgYpMFMsLU+yv3N7QRMSiRtepCNePq8sJjo6Ao6psMVxDEYxgsxvjN8dm5vQl
coRk5iSh2/ZPhYWdbPH5JzQw156Vq1y00k8HlxNwEMrz8QspqQJ3FZa8lHvG26S5QZ7RH7pX4l+S
FYbhHST9AX1/ZWUWOUP9/1xp5TsXsIARyqfbhhtPZqYqxH2c6kP2g0atmyKQrztfNmGcbDweNxJ8
Um6PAdzakl8nQNQ3e5QKnnk6/LuWYcagwjcdNn2MLBpo5cpkr9YrvcLbbom2AorkNVe+Dc21t9py
uWevfLiRy1AOQ1cK+7GPMmVoUAdLOFh9JqY88amaWjFCFZJSwGZxjAUJJKjURQh/gJh1OMSFqv6R
yHLrt8VJxldXgFaJUBQc1ncVFUyOefmSplyo5ZpM8ZAL4s9L2ZSC1rkvIseqkMG9GKmE0BKjasT8
FKYSGvnMkPmup/tMzWrxI18Qo9f4VYNSC1l7oFFtTkV5o9kOQPRrtKc7fSA6vNqgK8Y44R1jTnZY
gC/lxQ0+K8NaQWvMRRPxHgMRiwClM4kdEYwrcfmJPV6odjFo/U08XYuBTa+4DLxaJ7daQO525RXu
zX2fDC4/WMECDBQhXgDOS2o5sQbCUk2YkJm7GurI9QVf+OrAamQHf43SzQmLeGkv/5abKmmfKJuT
aoCDtTlM6cUSoznvF2pJBo4VZPQVJr42CH+hR+DzgtVlj5OONXzirASENP6CTzqjCXJJQnb2G6lM
XgGs7wyGzW5IxnHIdh4imuWrHWvMmHgRvO5Cg03/f70OjwbG3nEPEx2Yep+158/yxd5bTErqpEqv
csWL6spCtjfg0RVICTcd3ID/IQg3HwMtqWG2jUwrh3yiCTjxu6OROktI6wsU1o+oVEEUEWKQIUXq
jKs/W5TvoTr0xKlm015+NDgShiKWB2QidIIpCrY6DlS3MsHX02X1PzPs7Qn1cJoOAffti6HwzFWE
IiMcgGF82tu70HczNV3Yf4lYTQmrAPOOMcFOGBOVx9RoaW0Clwd7njvqhKqCTUInyqn8YihAB7UR
r3/GdS84cq/N1PO3KJIlf9oDm8wIFHeukQzEmL9i/7cGJKstA2aHo2eyIaEBw7nGtihmmhIWhu76
ieMKOHOwo2k85hDM03HGTRdxhzJw3pE7fibkaxfJWPSwJPmUXVR9KYBLttLD3sR8SAwxfxSnQxw8
zg7Jxcg71b5h+Ps8t+xQ7H7L2K6/zYTcKksHBOg8tAPkbTS48N5kP0ejYqBcgxAYiEgphQTPeP59
Q4TFP8vO8hSwZ1wbRchX7uG9D0LS4Mcnh+uR+jeHRBb7vM72ATyvsvHZJGGK/PedmYFiH+ou7fxx
gBX9WmCH8UW16x7wfv4ZHNpO3dzphiWQyjLYhkkO2Xzm/YbA2SAlqFrA44PJu7o88T4qEeaf1BYC
cK+lcIq0gJIlXh5l/9YF9eB/6NIsYXkSSvlX4hwrk6mF9AD+Ip4Fa640cnduPuQUVGJB2Y2Wvjmt
Sfrn3AGhMEwsVZI9haGSd36XQ1xoW5WUYLZtdl6QN3hnstfpOmiQTgsUC1HhCWmmogGOzcsi+bLV
ivoclMZGriE5ubEzmzSvvNEWsBjhCn41Xf14C5PRuPM4rfuzc5jgycqunfrg88cDHWmokVsrqMdZ
sNQMRmWUGJxd/XptNpaKWHxxWGID4A1vA2d27ZlWM5n+6icIBbqap4GGh4dfMLiWSi/V9XAQ9aG1
Yo6UzLY2H+1t3k9VZjNidk3RFKdBmcancL7zwwpiVUfO14/iQj8u14r+bg86yg1v9F2U/we5E2iX
MsKZ+fIkqZf2QOAQOS8BfcJQCMbXpMR6VXcKZm9RXGhpkSJ23Ng4pJ9WCN7sFhYWbZ8nHCWh0tVy
351aFaFzH4U21XeF/MQIHZQOnJ6Dwm1lUvYNljNY2GOFfmc5G+Jp/YeEXuW8CF4Pea0IO2kVMvAl
gMVajIOWmcBxU/sGgcg7qAQmiKHcywIbBmi9d21xZq/D1aF0bw9iBJoXtFDpOJ0FROjfPoXu95u1
J18nopDq3iUIgo79pEKSBZUgJ5NQeo07Fx64qJGsOspEH6pRtifAVBAZpAY52oENq7pqucfejXbp
KzjqE64zq0rLfhcP7JFTMBFjaHlJ7iAcSPaLcnGcWPEzNFPbe8Hjf1KB/WiEeDhk+h52380ZpoiD
M1tY/hElkWVF9T0CfP08G02yfkxPgDfaZ4vf/vkpY+h0UEfD0qYdKbIg58BAsZbh2hXMBC3r2bX/
veF0t0ZeoBgVnz78oxC4Y2qir4rBEhSP5xeRASKPW3GgCH4ie3fpIJTLgTLBnRNkqN6nTBeYzotX
hGs+EBIdvDTNnS5LmMl/4hnd81fBSXSRePAhC4W0AXsdivoGWFBIgrMvo7zikZol2rRFqf7QUli8
SEXfojL9p9vc8GSJCVald5MudNEMQXa/R/DiIQxpyGrdPnLMTu82wSpGMArfUu7uLsUO8tvy+/vf
v87ic3aS/JvoLn63CP2yJAD9e1Inu9m4TM44qTobMM6Nye9mpBk4mkOstqRQQIp6wCYLdbCi06Ha
6wSNxTfKhnx0NvVDIG0EHpWXxVQm5hsAefwdNjJwWXoVgftR4ghlJPaVYll5YEuBbJKnKr1qzhxw
SmWWQtWcc53lf8NvJUE7VD9BRiKNYQaeAvSkP7ztHSfJlGYqBiY2qBKrqb+btqGaaf56hwrAy62p
ExNdTlVpNkXUG6+s/f2E/mBy4MsOYMHGSxnZRSJRQLv28ADjwsMLZQjsf2PUAFj1mn5AtmjRQQcv
UP/7aa+yTVLOOPWYRv3vy+gqjY1mMOVAYyf4fG1fNAWYTV8PAgvR+591vFFEUwAqpLZRTrWJ3Lps
A6Zrox901YNkuf355IXIneF+tIlfY3NBmce8QNk7Q3YKQsHlnHwHiD1FgYpNr2B3iQ99zwneTkBZ
rTcrS8spaL5kZtuhCuYokiMdtiP+3w/Bn0U+zUWDTtmbEE8o0vqG9R+/daaGw0qGhf2bWWx2OCq2
KRo9T+lNjioy9YVVnqED0oOF5eOIK7hVew1otAcjyuiWC9oHtz2JqbN5SHJ+M1Cl0BjzpJrriCB6
Qe2L6coEQDU10fHAB1ThS9Yws3PcLTvHNp5PorxLEaAVZtkOhuKfDPUlJM1v+1KZaFZu0UUkBCF4
bQOWa2YSdnz4l5RXg4Uw65sNUQA4GxrYmiWuDDcKBPTAupCZtCWQgHoXgxvpMw9feyhPlpP5Ua7t
HGw43D9yjDo6+55etDpv0qcynR3KWysSPu6GpSENHc5ka6/bAuCXve+hzEabqO315g7Dk9Uhh6es
3lDTQHnRVZ/LXkqmEtWs4daYMsK4VMz4wqHed/z1DRy2eOzsgDfEvbnyOl4JkBgFH98BGARxafPI
zVSvS4XmhmZNgTL2DDLzdusX9A9TD/CKg225nMjUMGtFXkV3U0lJUdo6ziW0eQPwC7i4yLnWxBPN
Z85UEeLgYaGwaQ1C0+wyBvAeE6kvjWiMy0m6EU2wPA2FBHXWcMzW1GdMM8zdBCGou1vSQ3VWoU3T
/kDcx+0YFsUl+kBeDCwV/mXO69vAJh9R0elN1ASXnYr508T7vqqlqBhcDaWa/n3p53T3AtH4bp63
VTK0ljYN3bBwTg1VFBOWK1Wg2L7KBImgNLl0R4lt+8QZ/qKGApJFcwOulbwCpPwCPJSi5XPY2nMI
QTg0vY/TdBKcqaYb8i9tAX66yTRQ/6GRJVScoTzJkNAgIkTJt3VeycFF/lKvMxBNLnsRF3GqEDn7
pTJn4nZ/mCnYKvMjmKBpp/Ai8NzJuHSMu8Vmjsf9ARrHDzoK4sHAJ+oKaUV3ZhElvo/st2uBC4Sy
aLB02SB/uBSjx8ulpZJu61Au1/9t6I0FcPZZtLat7HLk2+Gi+x0bsk56fyxgVdxrq6CaqCsL8QXt
IOa+XTdJ0Q5bWnLvvRZChXrK3KHdWOJfzjsbhCymgSI4zsKfr7Pw6Ps6SBkqOTuKzlckVsAM3PYV
PVspKnrh1A7Fci6BdY2W+RoDblkgkUCFzrohHIzy393TrlVEuOoBpysFwjQoEJFXZSagjZ8Qb436
+Pzxd3nSXcRCO1HYxPv9MFfEL+r3ZMzWCwkAuUoXihO6mjnWENb3Hegk/s+QH8tYck0I0ftD7pVk
uvd8BKtlsZn01+UZl10KrbyVRG83vkuyDZdhDD+qJRymyujZ+dRFDt2D3zX67nGEukzVSQgciAWK
XYDWyB3SD79DCDk15cLTGWRm5vNMTMUZQrfgKrgBQv8woZRYodfx1XseubETMX5EWPDmSrehSEHa
xSZzfpCdHiJQv+cKhsn+ajWSLWqodG6EqhpLE5zku3tmXSLIsiG7QyfgJYcSQX2mec7kyWoDS0Kv
tpUr9QtBoIlx7sUgf0uiCZUwN1/bQEUQpYBXFodSaKF8+95fhmUw9/mbPT0IY1JPN+Xp8Ckswfkt
PyJdFYUT49PJRxtzRuhxgzMss5fN2+Toesby6hWuCSdWy6lHgRQZUNVhDPpY4E7MDpN4rAbf9Wdi
ZMm7y53QSLDFlu/VJZMGfPSB1VFP/xLayOj12WuDyw4y+hNSp8lUl9XH9MxDet8RewMV3e9m8+kL
ijsURuvvbGHhgsx0seJ2ZJhPXmSkootxmJ2OLmlVJFR3Lf3EDeNlCYP8SuFu17L12Mh8T/0EOkrM
U3cHkO2nBpfpm7bK6JrVrr7hoti+b1tijAyqm8mmo+oLBb6j9fc3Mw+UppvxB6CB/B2Kd2qzZgde
RtR0aeKmUw/k8VUFJ6yR/yEiWVW4WeKtmuPelMqK+4tDfA16OxZoawAY0H8UKxyhMSxexsAn8iTh
zpyKOY6Gjks5fq1LIsMOIbOYTK4rfdgCQn9jNNVUIuWe/UxzXokEg8hJKj4NDDt4OUloFitKKLVp
prcVzvatwQLYfgPw/RNsIMqa2vu0N5m9SNQ7Nnxx1SUJhsZUavEI2zMUVqN3OtLmx1+NsTcHlM79
Uktkd/zgR18dJ0zI8MmWiiq/1966q+PJou0VPVOSLDnFDJcctZEaoYWGJOMVqp1Rvo+xp4e0/O4o
d4I4aeydhQwWQjGINxqQk1zec5CO3vyreakLhJvh19TwDwRfY/aSjmaDB7BH3FcvM40mWV3uu6sV
DLatTKp+bJSD6mfYiC+Of6w3qwUKRh9xvfSUegQz45EKJ2iJvw+S0pf1s/dPXlMzPjEKNtNAvBiu
qOevML//CuCFrql2tdTf1IF0Bpzd6rn5T7oa9RRb91MAlUqxYNdkBoQG0eoQ3S3H1F++/qg2xRPb
VIWVxcTzC6s1u0kOPOnxCPJA/I6D+1FLVwqUW4rVzMFwYJCddQsr3HMoiLFQ+TDPGjrP73T9lweO
SSI5Q1Y739Y0/RXt1ticWHrZcrlGQIqvWx0JStIdxN3KkztjUU4reZcf8KazWPXKuVs9qlJmblHk
HMG8pUSV6ncclaQdcii1im5gHUCmLNVWOnk7GB2NtfM+YN2+OkC6lRT6KhlB4SILJchlq387qTNG
fBAwOfi+sDnovcGsRPwCbfmCH5nBjUrBRHd35htLv7KPovlsiaKpLP11uvH2qxqcHd/5PRdQxeA3
Nlhrk4Vnd50dXIH+XCvFB8ufmLpPOSofVxt+1UctBo2uX5gpFSo0F5c8qYR+r9EwlA/Cxt3OmKli
s97L5yOQb3D219SNs/Vw6EJOhxzoN1VTWhqIP9pIpU0PRLgX2qXteS8PfEFsnKj4P+APYlSp5Xio
rmRZwC3VP263vVklLNzWQvfW5LnG7DnuP6tKlaFE9O2UVyO/W/sN05vXnb/zLJXiboiY48RfX1Nq
Zy26PtlhzvngEzSN45mqRRM2IE8tLGNDmfYVW5NAvOTDmUOvjikebnbhM4UNGymp6LzXj3VBbK+r
uzb4Gbr6kSEmnYgocghwUsCnkceRmgpjySKVpgnSoALzjp2NuKvxMcdURSjm5ouwRccZinvsMaux
HxTyeDnQk61LtX8HFfN7NQmhdzGw+kPDVpC1BYaJcWOMUKBgGtocMc9iHkEtnECAuqRU2se7D8V8
no0Y8U3FbQg86RkQnqiZoJ3Z7TLH/AGTYvCXdJd80XABO7PvRGTwRFvN7UUMog5AjnZaVtpI3NCB
c5zVjSOrmgDlGnFZx89YJvSXTaeeECahYYddxD+kTFmNTt/4G2IrHJkv4Sfgdq2n+xyn3flMDCM6
7myfj3fllLWzWHJDpATWGIZjgdbXdP29XA8OSi5rtvuWCcuAdDkH4ea/fL8JQbNPROyxoxd1HulY
wzIsR6A9ArMA1gjRh1AIRlometZ8+vD7YbDs0ABE/1RIs6uelFeBjTGjRXTiYX5gu9aL6kotRCVB
vTSOt4mar8DJIr3262pkbYsJXNXL7fsl7ye/lb0GpyaMzE5abyZwec2/nkjSG/1KVAeiiAz2YSk/
d40JA1kCm1tgwWe1bukAfVi0yH+7Z0w+2ptCW+KjYcTmqGx73bnaC7TaHnTtlIcS4RiqMvKYhmWs
pMCGkel3674lc80Sp2Z5okaMCTLA78xYLLcU/Vfy7MUguc/wMWvHnsZuffwbzw9RTrHd1JH1rC4J
C72dJZTbxE1hCBdUnZeQDG7tJcatuEqEWcvWWjfhbRzmyOuhUuZ59zVB88tTsb61iaYGrPhrJn37
l+eEt6fA30WD53Jnf9KsFy88Bj+BvRQANiVSCSuj+F8ynLkGCgc0aS986ZCRcU1Q29CwHaLBLBsq
VKrNF0bm6WFsHw/YB/1kCqrka7ujGwZU+e4H8g9Fui1O2CE4tkze5mFHDj9clU/SLBr6p1sg13mk
ADs0daM2qQc64s//Mzl9dDla+n3W7pY3wZCGf4zYSXti51sWgEXR37lfKkPJYC3vWBBeo2m5se1Z
fkA5jt1fGTk/sUj9KtYlYqjGGVZiIqMUpYCDS6zk7l8X0m5ZDkjNS9bbQpmosWyHQH21Of5HIxdy
UCF1yqPw69GOXuvy8j7WTVnJ1GvCJXWbrfr6Tw8UkKJDtsc2rYhhmZIeMXINl2fg7Cf17xF+M2CD
WFLjZfYnxU6r37/kC+dUuhcK/iREEGkNY1aykkplCtS4wIJDqZ6qdou4LlsN8I83MNKiAH/NSQre
JrHLs5lE8/bYfZ0pJpgA5OP6Kh+S/jZ4rLhRjNgIwK+RvSPI235dn/pJ9r++sDVgphvr8khtUbYk
tMoRxxb9hcZWeWVIFNFnkGS5HuydwshDrhy4KkeqM2aHGFTlAGgTVchRXmcs0rsH/He3bfC5Dris
2uq/Aw1tauP6BnXSBnKHQhb2L87STISv4D6s6H+r8D5mCNnTIdcVFe0CymRaJIl86VWoe5xu+lDt
boZBI3//UV3gUAiUBcXkuofzRgn5193qAIhoKCOi46GhgZ8rcry8KUJYkEd48tjCNKEe+zCo2KCJ
qxcmlg2fyLtBFQ4dBQf8IdhCjr6/cgsitRw4hYiZ5jzOoxP/hZ6pNNKqGsPECrByA2RajhcPQTvy
Uapx8gruDZdKxP0nZv55gzWSSht8zkrr79hPq8/96wsnkMzBglPJGJnekPaobMbLTiGXD7cvEZIO
GdpACU5LbKTyol3PorHMLb6bubX8qbn43zo3z6VLnsZaNqBStW5oCsMCyvnFLX0pjSGr9IXYWeLw
cdLATYAXs38vztv6tIb834AueUyzrboaY0mmEIlZJKswHBOnwpYDNaNl/M5UoEhakwr/Xz4nM6bT
OejdrkejthkceXGLUEDDE5G8En/607JVmRYIvUagNxV7zv7IChSsSGbivIuTnCaJoBgsGghsXprE
eu03K4VBJCeXbBDCaWh2XmBV9nSS6LxeThPspOrfF+icm6upewGCrod03Cylm6tO8Z764YSqmVZh
gD5Blt4BQyINmniavTvQG1uTYqFMstUDodlCoGHMkYom52u8LYbvumGehUb1lJenLOB5D0hiRHIm
ZErhq8AdRnuvFmy+nl1EJAu2D4hNe0DvJfTXpnihX1E3YuCgFulz11qseuQMTRQbdt4FMeQMe3fI
L/4JKIW7Vv8hi8gHHJFq3dGKTuzQrOoem/OY+JXZofD1nGWP7HVTyYTHHgg8qZxX3XN2gbj5PdHt
ladnpzQAa8rMOEvGGn4tnR3Arw5OWoe1D1QIsitpOLdTSIozhYY2RD/i62JEt/AMWwMWWmc8Y+7N
FhHst28EJQvgBITx73XtYPvDpfWMSM89t1vm5Fh3DAvRZmmQwa9ABsLa6sn8PEt0J7s4kxm0/VQZ
pxH6LmehCUBxXOR+Gc6CaQwy68Ul2AP1UJO423ik3NLgWlW+N9ZLpwQa+mhuRyDbSDbrkxODNabV
EdH1cN1xuj2ubnTW6tSiA/s5hP9npeqWphgGpAhzkI8oD2j3takJk1Ja3ROK8K7ponnmE+P+hj/Y
ntHXD1YeCtZ2yedoOb4GeR2Y/ps0c330jZ3f7mWyFWHGolcQvbFgtFt0b6wKgfD3ptKsAalAmrQD
YAvc/sE8C62A1xCU2s25XDAOkBhTs3SmDjvJJwHVsBUipRo8J+s6Mxi0SKlyZBqhuFUdHdQCORBq
AzKCZJ2gmGJHoMvBmFq6j3dRTjwVAnnh63RHAhhsF8yVMbp5tmYXxnkW7r2Bmo1doclIECjFZEa5
7lsDQbsPLiR2/YGWOTwi7BFgzgkoozqeVWwQsNnJ1LeeeK5t1cAYxY4P6SUrvDF/OE3l8Cjy+r1x
BJZes09E7uRazcdydO0sW6gf6yvaQyQo44Yng5v4TsvAi/y0RlruHDRcYqZKwHL29u1mcdz3lV9M
ikX2m6mS07PGhddzgRr/B4EKs5avYDl/a37G1pDE/V0D061/k+QT64u3jeKMS7cIGpam9Y+M9TvW
63NTO0o+Q/PEbPqE3Pk8JUNdOYf7UEjjPV7fhaIy6VY718iZ3/BGHQ5zVs6niHl9Ici8kGbuOdJt
e2cBGMpMmNIsJReokwrj8biOrdgw1w70J44fnBJEYW4Iht4tKhgECf2h7YJk7cU9lvPGqTM7X3Wj
nodDWrIzK+0Isokokb/fNGeGZE7irXtyvVAjh/MPN2ry1jD4Dbny09e4AhBh/aOyb21NSR4sqbRk
FhpB0zsNwbaV1U8b4iXTrhPBzNADFKdJ7DaQQ9pn+AaX+dvR8Cs/XG/E1euLOzU1ZOcJHglXP3R7
lldUsgHxlgxNJpGfOiKR1j4QyNiWGhvriDkAEdAw99dnaFt1dtGCt8X5pOgpVK5yLtRJ6QgaBRKT
sOl1OyIrnFBawrkz4Q3EKBdljmLBqzM2X/y5DJKAgjT8NemHO9gpkfrJTALQblhvGOY2Z/gIyQXV
Aq27FJhAQMhMlL/apj6aIdHb9PpBgby6RT9j2Pebw6kojMfYsDG85RKJfgUUyhVoEhdZP76QttZ2
4CoL7K2r6gY/3C3ViRurA1U2G3M8ClHZzYnMio/f0kMgxcscXuJseme4HuPF5ytx+ifOKuS+oEqo
0KN3V4yadcESyOnJ07h1ij5R/8Y/xpQ9lCRZWaOlsDDBl/ZbOw8/ScBC5lDQ44Szl7/xHmJoHKxa
vRcIigBOBe7ClzThpCYCGz26iMB86zvDi013XABI6mZ6X/C/TCAdT4hNXKOIEd54kjhHw9keCHc3
9s6fLUqU4ZjnbpdSFKc5mCzPUZ2kby7tZw+8LbtSTu02D6bXJuN75jn5UtfNDgUDdPKUQdxgqm9V
Hl2Jkc2WS9Wha4kEakvKxKBScBRoZ/FCA5Xx6ydhkYYxEFXxPMR9NjZxTzNOZlbhhxFqyUC3bmIM
i3GaB08S/tw/TxX2SFJ1tppG016wURCU+aicRVY/RxdQMQbkW8GfyY7AcViFjR2D802LoE+TiIEI
4Ncua3s3Vw6KaH17nC/DZonuH7SzHNhwKyPPYJ5+GdJk3SKtMvGHvnQ/TfpSf10mE3EHXBIibE9U
qJH/gEzHVT+a1KA5pamisra7vr6rsC7awazELvOsy04j8uXQtrs/NiqgY4DfehidIgOGR9PENqU8
t6vzpcdiPdI5c6C7guQwjVi+qQyhEJaKPPBcQZcGH5JFlG+jo0CPqsnHvn/WcK17w1YdzzibP8VC
NamGorxHArVhgYdgVuOPPUxVUDwJaw4S1tnq5YRVQ6XTS1VDRqepQTnObXB71P9fQwlVG40GaAno
JtsCJOtu8BQ8EUQXAtQ5QY0mU1FzSwoWAZFzNre0gyozc2ubly6uRFAVF4VQcunMDPwUeLoVvgcx
/cNZmg1JLijzuyxh1YdFH2t/TN+fCzc9bBPu+lZxA6L0Fm/SUEdMu+mwPIj7XyaM8aGWx6Owh4kt
sN8K/maY5WXvB3k8boszn24FMkTyliL0ZhLXnGe8hIuK6l+H5MAWdWvdsEzJEsoggnylZYfMXzIF
MoF9C/5lQx8DoF2g3OeRLQy76xUyPA4WtXAZzkQc5MesTUT3W44CJehtPvg7EDAWf/nXaOBWuzXk
eTmAAChUNLnmBYgBVqUT9UurXIhuzJYKIQ0JnaDd3zCgaW80o6ZjhnefZV8bOFS9CPUyfKMAz3Fs
Z3Me3jOTj9guRiBEfAOq/AcemG4mP0e3EXEr56wqGoUjHXkUH2EkoYDTscmnLwZpDiyT7Kj11yUc
QBaM9MeGw7GZEIyoNJfGX1SzTcjLcC+rGvuRtfFEY3KysdG9XXwWG68Skvc5wF8sxBzGJ81Q8Zqn
bIul0JK/2o/4zmCwfnukAVd7AhXqO97a5HHkBH7+lBzHHb4nB0fYlx4DeywZZJv4uGVwj90CHBRu
Mq9Ws7XU3itUc5ScSnBfSG5zydwjgAQ+GADNVMVzq0YdQIsXFg328qt5WUWvocn3VFePDs6BL6yi
qVMO0UI6hjpw25g/9noky23OqrPY3Xp36yID7PZC2rsj/DCIWBXfmstGUZFDagVvX3rLwc7AnPMg
x05xwiAhFJNbvpoQOjndszUWCopUl5GqYOuuyPrXztiDJoOZ6ai5l2NoxpRsV0ML61Mm1NFceR49
KdTTmG9zFbg9yUKXcPL+IO2MWVwGvGvCIqg9+ntf6Ey9SXsZY8gwN7AgybhlN7CnpotUY4UQQCAF
CvI7z8LED7ic4t6+9HJQ3iuF5GA/qyKcswceS5Q8ZF/TWI37gA/u+5X8DHoyG/oKsMVgbkcaWscS
6IQq+uuaVGIXga1Tju9PH0LjwdWJyedG2YmU7pgPeCtPFy4uAU/C0fTjUuBHOiLHsJvGkQiex9NE
bOSe1zF2C8r4Q4+ms9ZYku1XD+vm+jlI1n5IroSh47Z3KKVrhvoIBzMlWIxhJ4xabcHBMCShBYXh
148Rn733C3Yb3eugQbHReynE2GklaT3LoCNzPg/r0mFhxGbN0vf91CJcEGc2UC8CFtK8TKBmAMVn
3RtQ2bCQesaYKbFeMgh4SMNvS8Q2U0LHeKvzKej8/rJ0xkL6BWEW+wSck8A/htGN5C2Oaet6qIUI
JiKxTO9wqSR0anKSt3aTX5VReRxfxqlBtzJyhU+y23ZP6zvJey+eoPqGcMiuKApajoIZZv4OO9TA
QmBEXMBUWBES+XEV5ZJu5k0clzrqg00ZQ+BR/ghQ8XsBmbs4g6x2SZBY5+9Pg+AiG0Z4arP9XjXR
nHX/RPl7mliPIbWq2lfS/x736w+kKv/waxgzr4aw3ZLACOPvxrRK3/Q8u3RsHMTmvigbFiR3H/Do
ft1tm5n24MVqcdCSxGWvLwVgwSqwSBCms6kBNf4un8MiMFPOiQaubiKmXl0lxyX4bRuj3o2U60Li
QXYBZKdSLdK7WwGLjpgrYFYbMZ3Fz8KM8L7AXksCLKunT+Mv4g9Waxj4SlcAr5ofkO/4YSuoOK6m
dYCQ5ez/tE/1MHSb0J4Pm0Vy/s47ieQVpGynfWcRkHJt26kZbQhoRuUdoUvlHmxhxPlTqs5+ZmjB
wVvGiRiByjTMipFm8/OGsdO6UNcx3Fjrn9y1zsiWwryvl4ApoUBm7n/vLNYAZu8sMuwo9a1VeYrD
iJmwbpfEKzzTQgFVZ/NhWogWTWJgOdUuLmZdpaeZjwzko5bvEWVi+co3wPCIx1B5+o5OgqQdyOdK
zNTCbKGwPuyjNPa3Fnpvo+6rH7dgW70w94pLcmX+To8l8hkvxCxppvUaIdO5pBERJEnVjr/Kft1Z
TXGuyaQE2wFFUWcd1hPeDN2XSbX15khkRNPO8oO04HPHgqferYyO4NMeyI4230D66xKSAEeIh7mu
OLMwscuh4uNqNjFlTXFWLRFrBNuaL5s3zsroNPqrjE/wkDhn04LJsVBqP5KdF7Y48NXXv4ISSsQa
M1k5vzJ5cdBmFIeHX86KqdZasn+aWrJyCxD+KVYNl2COW1dWsJjVXF1RXvkU9NeOYd6nnR7xgNmX
hxza63wUnGjIZ+t0aCYgy+30UmS4yLIiOiRpe5m8kyTzpSdyVAfSkwt7vyzgV98Z4k77u3iAK/TY
ZUkcgy3a1aFFS2qRkpV81BOKqYomPv7wI5/1AIwh17VfnzJjeYCOI4B2yc3JYwVhvahC50d7XBqz
IM8h7CZiBttvqgJIdSc5/QZ/NkJDUtinsn10nKxrGjCQkLV1doXhi2yUhttwRpI3K18vrJW8XUXr
1jWpR35/KRckGgnVjL7CofmIiuW4jK4auemrhrxzIxSVHhjVEdhJhbfwUdxtKyHuAk+3ePea96oe
JCtoROdamnuhUNA/ijP3VzkGYK6jQ7vk1K6W2bJua4xUpSo3+Fh/eGW8UPAy7vFTd6qrBm4xaAED
abDdU5bD4iXMB+NRY0wpTWakdKV8RTDcnRIASDndn1cjSDJyQHYEYR96WNmyebnkQusmfUSLK+Ai
6VVlCBVxjRMZ5f7+vxw29SesLzkZImzCy2F9H70gWHWVqTofpev+/j7kpbEsutiiHc5kzyfKmmyW
Lx7yx0L0flnzYZvYWzRHe3BbTGF4B63PbIa0/YQWoBniilJ9aIwb4xr5q31App7YILcbTTW51ah0
jv9UuvcXzdA4tSO12ZjkNzBPWeGpOGT0NdlQ/7PMcuvLJjRFP4Sr1xIvSawBemrp1QR6advNnn9A
aBO6BxSoA3IRYjo/2B9E5q/XL4hsBeiXh30CxWtZu6FPxa5AyeqpmKlHhOACYc4bM25FsriJz4JJ
181xn24lXOF8ff8Ns71wnjTnM6NOTJN02P+xHrGLi8FjPBIqNvYti1dcNDW/TKuNe/N8qnFR2r+x
/E7sme3mkRazY+O/riEFoMRE7rF/L61+N0Ip20mluDiYIhunnok7TUjpnOyEagYIDwx67cHA9K/3
D5xwm9PwG1EY1i8T5BIsZeGJrDpB2cQWUGAfNn/W3c1EshVqeeSnNsVs7Xg2Lv0S6p509nmALIW5
0Qg/1mquoCCBUzSBsetGGB154MleKGZSFYvrs1Lngq+tSbSZXagaOgPylm0p5t6iQ2AxjwPjSXZD
sfaYaZPnDHnHOhhAI1jj3PtLKN+27A0Woi24eKCiabN8pMtUJlRXqXCuyJw5fsJt6f4L+sSsfUQA
564LMo6vIb9GbBiQIVUae2pGroAXyOO2LPsFPDKB8dAQtiaLSO0EWhhxOsTPoSeLoRUw9Jgq27gy
8MIcCLtdooJlrXoxUtvQG7G+CINYvOSNZOeoAUPh0Z1/SlLCcEegA3S51GsjwthAOomU77AqN9P2
86N0hTe6A3M55deuxPaYOytt+LvU67BjRZyrTmXU0wqrR9mUIBuWq1a1rF9r0kSFpb/yTHMAt0sA
piio/jbfFPqny3ZB35S0S7My+fcNvW8vw7GX8nPAFMUsFWwbhTzpN0S+CsZ2D0bnIjFuYdRwn8LU
vl01wGTiNORoCLwwbi1YwrNJKF0bx90gS1Znt9kWyWtWIaQoMx6Cx/+3XnTO80HAQcPSmBWXFEu/
+RkJMrScE0EhAzAQCDqH44ieoobRIiqzZE//kh47gdXrSEVef1V1dyJwFow4cHb0v5ipATJq4BL4
TwI/fbAat3mw5po+mXuAI2ESJZf7T/S8Fb6nuG9513rTdUazN/lKABzV2N69ySgYqRI3wDZSNmzE
FrAV52mq4/QLq4pqsgFf570wb72LJqhAGA1ij+Tt7Bf4vxGiEIR4LCSLge3GGpuwKIXxzIS+DPTI
ZIEMvZ6bIMSwTHjGOW685k/db0GXYqdXd7tTnR/bcut+1R4e//d0ryKb0Dpdlh4oinOlz8CqpGL2
SIEfwSuHliNWBGC2ROGIO2qilp3Ez2DbDOhxnMAUOJmqdrXpvO7sR+vYW/3GT72XgA8ztJBTrW93
wvO6DEgDnpUFIoZMFigiPZoSESikk5qaHz630c1XB3x+6ZSZW1mCzrAtOn+noZnXR5LoB2GKe2u4
OtZ/2tm4oD3elrxBD0/kQUiI7TvwyhiV1YpFJJRB9QnM9XYicT0LXa8UnaRq6kKnSE5LeCR/kHER
UvCqH0fd17DUqLrzVMG7tXAUBS2w6nb0w6nCaRr5ndTgxvhXIRouORDdRT2rumuPEHQDr68/uH7a
NIIyXCmmZZVKW3F13fao502xhd4weW54FyXXwlPpPO8kVWKR4Vb78O0oypMhB+Z6XI0tSRZYMbTI
W2Ux0+4Z1F8ywCFaJvWhki2ffFPBbLsHsWhIGSxwOhn0oxqjP8lPzyPJYxLV2ukJdfd5TObTVlW7
IKVHT/UN8Ot6SejVzPoUOgjbb0O4bfuucPinJwrZG7i04MKJzeQMy7qexPtbhbXRG28rAx0FLkIH
ENx3+XsjGcsNi07G0FjcT5rbhedeQHuxf+FdWWE6pmYU+EBqCCoV8bS6MFHcqb97i3cH+uX5wLpZ
UEhETB2roCU1RlsXd/fuDVqpkUtDrhlAVkKf3G+MzEgCDsLl/dRlRnYHNdSKkme6+oadYsOG2ZT9
vH2nI0X3z7x3sM9/P7wE624vss1oNdFId56c+0djOalLetyNrKq7d5xok57V+P/vpighuxprimgS
GfxhBoWgaL/8qJZVGh/FUdLBnk63iIZypDsJQqCOsLj1jDCKB/l0P8xoE4htSJYH8gX6LCprlRdt
KN039zZaT4WT4azQ6IphOuBWwlGfbsa+2XWMx5v8Uxtcu+KR9eRYu3lcTglae0lMbkn4BCg7L2T4
a+IcK9bFSSi4qXbiWsi7wV45o3Ft1lHXXoXBeDOplAlN/ZtAeZtGVzwgEuk9NVS76NUEdBgdKTSD
ZdMjQHqhTalIJWDuCgrnoShRtpbmdyQK6XbCClHWPG9VzI+2FZLGv9o6t+CQicVYk21iSLKqq1c0
xy+0TeYO5MjJ7c/YuRf6z3QH6Y05ttksLzQSTnyri81DQaQKaW9sgWee7Cc3T4BEm+5J6ZOZlVfL
tF+/5262Rue207h22gBvSbGctKAtB5kczeXu93sBz7f1kFA42yi/Hmaoib0Rk7MbpPa9VHxRvKO5
yKaeK/NxTNI5rQ+F2tRdxDh2Jx5/XU8bbav8hMJFZ38TZAnA4z7jcazCg76FyCe97wHCmV1kihKE
sso2W6IC4dhVOY0/L/j/QLYVbGWQ2WF4qSsmFefWxhTFp7sgs7F8CC0Z5B/OQUa96ybinaeCszJG
B+JxO4TjR3XW2j4D05HI0ZZaot/gt+52jgr0SR50dnU8Gxt1CZ6CjLcJr0PfpLjGbMwTA4B+HCYM
yMGCTknabLNkIpYXOC8s9k8tggTeKbdELbCGIvI4aNR3YZWikX5IYHPS3/fcbB0FpDXQ8ca6ukHl
7clytEPKUITHCi4mSwei03SRobm7IW/OvGIxv4kSc7DtmwJbKxdYiO2qWVHRLfgOf9RBxt6Z12rN
q7vhc3r2v4MGS3i9lb8wJ6uxM7Hb5BguKUqS25KMdXjB6v7QsRaLeFjR/f7WX24jZpiz6BVHmLSA
ypQHjJAgb4IY86MtW3DrusJfjALDvz2mvJ5/e/rB61LB754VUC3NiWIPBnuQVHDVY6P8r7brxNZ4
RWuAnDUqVCgL2alveVK/GCay1VRmuNvDq2mTLq+ZBSRWYR8GjSs4rj5ScZWmcNZUr4E59s7Ce03l
kyakd1bBR9zqifdt5AkTwLHQTceXWn3H/EbA+xCU8VB/rMKKAjdNQDOmnVRRVnwQvUVDzj0pLPfq
xik7WvtcUL9BGb8KMBamndL/woqpCzQc5bCXPLpJZXnsfRv2LN1hFC8PvP2pfTPW0bI27HHQsOGc
0wOuiXKQBQUvMd531iPh8bxJPanJmfDf5umGUMGSz1t7jSc4aRXdfF9hvJXJYWX6rFvs28vIum9M
mZyiZKUXIrjvNiChn85CgKRQrieAZtGdG7aiEZKRzHx5YqEDLCzt5D0uY3Kr6IR2mY09T4GN3Aw5
sI/7ElEfFzZED1wWRXoRu5qK4lsWYd3WN+Yt6pNjW7Fwm+p7JKTZ1RZeZv1bomj/B2WbzeXn7DNI
eLSx60NhE5pf7MgcDBp9Fo+weYivH2JZwkLvfYnY62Nv+Np8l/bXMkU2+VEJM31Mu8RKy66CzTRd
QiDjQ/aEziMFqDVw2X2lSbE9OOZHGMWm32Pf/DeIvBXwcrKlm7QWvGLPyLilTMWNR+H25Zi/Z71a
0t2VAlOCESQvd07NEmLUPJGUlmvlw8ylOdUNw/390OTXIzAB6x1I9OdqJzo1zB/QL0TCwYLXpUL/
Ds+YUNBRWvh8vIg6iN8uVTahxMjPHpTr1kgo89vZYvG1hOEIbcj5w3g4d/ST5nC7CuEH1B+4CsK/
Zjz9F7Ttvfz0MX2UjhgjisnlqIkGbn6DoMAA50WIbFroWfMUx16wgdB2dF3NtLeN9dCbV1vltjfN
Lc/YUUNHcTo9YtQrhTPVSeDQltR0hTAVIz0H20CDmOu6KrLjhxEwEap+u15zJIokFtStaFOP7V6T
RaUVOtHRrg6/NMdv83c/rxAHlX9mLaGbA29MIneZmwDX3y12bdkrRjAigYPOCpjkHDx0C/SLYK0m
RLQSUcQjVeVPF6T7hupf/oo0ZscEeXAmbZKXVLo84Rhnyr53D+v6nHbKROmF4OxSqiyhUJfX7R57
AS6TE9jGhQwgZupbVRbTD2nIRX/TbHsE079JRysv6c4W2HlihShA9/0bEAYmb1nvXTdpimq47LWV
ljkO1N4acfWZWZVjQ8e2mYdGWx0GIa5kwBKOajWKX9UYtTgAI6cI2gi7SaNgDWnrfFdgKf+Wh6Ew
ZxumUHYhzE9eHyejwwo7SnZcXTc/64N0rikBG0Xd051+d/watp1UH1uMpEBOpf2ouHnypxpJ39aR
d3XKkiart2BagV9dj5uVRnB1tp3zajNl4hya9+GfXkB+HZGArtj6sGwajVSJ/XP1FyxdU+ee3qUa
cSwEENdAgeoxHQG7F1WNKDimszpGMx3Pl9WM5EZjqyNGUDqExu/NKiq2DG1xY9+qnA6DZ12JreO5
5rCWB6gT/VgpzW9qg5hDgG5n134xkqDkp+z20NWS3iipea5RLQWgv3Cj9z3eHcnX8CkGGIIMyNCr
E64Xt0PoG3KRr3DTKGG13mYKyQ2X6LqH4lUhgj3+BlGbvgb5ZFeOf4VKYTmqboiW+G5tfGbOS4gQ
ARDVvaOE532naTvCiYEe28JZIY/CvYL05HFSfFG+/ZfNfTDBgAhDG2OwdTtmIVkAAYFjwy9e6D7t
3JhxMWZrgSJKLhQoyRLOq1NgxO8f0vkaslZ354e1zQ4mTuonz60cKz6WMoWW0HKGdgeIudHX0H8O
VBBgmv7g7En6Sb8HoGA495P9KeOKpy3pPoCranTQdv3MMCw7dkqtHz3cw76XsK3e8vdNXxy+YQ5F
AGACxKdKKS8+tJ2fyNP2Z+MWYRZ8wMvGLNBo9e4ybMggHEeGjCYOHbt6GiLwDj/abbJThO+7H9u5
fLSHcUkON1cL8EJMgo9nLFvcLB5NQXbD8Cbbns3chnF6B2sfmmWXJIV5l/GlAgs5y6rSmeiN/dnQ
yEsnFtFdo9BUeFsLFDpTjiJ2iGGO1XmExUEIG1S6na4s2mRmQzLxpvU1PvtNtwmixJ+QjsFPd6sL
nkjMRli2Q+CF2Oscvq2G7kYoDK2ZiItJsqRLJA38aXEbE1mWnFL6Yol8haP3yyWfBDkbiyVGnOt2
GeBwH6fwk8jGRT5CMp+zjTyvdfM07JNoKbwZvd7JaIjhRaP6sQTxpBgTwwqB4h1Ecastvkp5cbdu
2uVxG7W3A4gqksHpBjOk8wWfLNpLh3D9/OKC4WpZ87dKndQMaPRAhDHpFc7uUS4Pb8/E9WeBFsCb
n7kTh/tC9qe/7G0FhjCywlUWFfkyDo5yldWjMg0H2rd39S4zkT7YIRn/X4Sa1LcWu2d7PdiSd943
jlULZC152gQUj6jEmmp37E3C4bw7i+XHwtvGEhgJq3IhpjXWhhiDZUMdH+tzSA4P/HcN+YIsRwzA
kvhM9M0Jr0GZ8Xmuo13JSnVeFrfrvddsYz7IafYCeP1zaKXj41vOKXhjQzd84o97onJIOMVlH+Zh
hTC8YfycSBdYxJgpKs5zjvZL6AueEzZkBqO7iOE7hxY4KumVRMReQSz/2hr2Xzw0lPZg095sDdsw
fJoiF4EJLl//ThpQVt8mrIL6/NOG7P3LxgHen2SWhYH8BrLw/mSkMaYTBslyv2nQWSeKvn2XxDS/
95AHu49lN9J03+KK/LcxaDJ4vUZLybJ6oGHQYlTuP08CwWccxro9pFe5Q35xjhKTmFxeqSiD0cMG
G+Y2D3Is8eE6y5PCRD0iU/iE9wJXBsvyqP3G2V4Ndc9uFR3Te12qSpI93X1kM6Bo7eTNUaIQ0Efj
eJEG1z6UA+uCIs1XDIN/QzQO5SbjR7p1URc0Z3x1Hxc1H6J2G6r4NiFUZbrCR1I/9eHxDi6NBurj
ZLC0+FhA6vqFD1Mi1O9i//xLwkWWv7269vby9K85dBG0lQZDr5tdP69KquXavGBeJZe/5Bm9IdYX
f7WdypdHrJ/Q4C7CtoStdmwcW5x5rsYeCTCoAP9yo1U1kKx/J07QdVjlpjdAq4klpIhPTZ7+bboy
v4WUSUwbQHym9rMU0TXwb5IWnXBRWxQynidKhfGlBfKpEJXQb2UTS6BHQZZyHqVjajl8pgPhStsW
OZyE9+vGhhXPONuzabS/zhLhVbT5DV1gyC/rlbyK2aaPUNbXUHnAzTrCyw1KbwbFKuD04iMt+MV7
gFA1C8O/fnLj+MGfQ3p59NoPtEjAW33/rTQPNQSGP1D8HA2WcO/G9oeMBp7Mu/Q6SboQbE5Ywtxi
HcHtvrRQ4UJZPD8RAtsyDhIC9ldUf8U015gX9m5EuzRHoGCM3zjobSo3IPBe30bLSMSNvy6ATKA9
06ZR7pPQeYgDuwqka7varqmJt6T+2X25A4gdpx08QLwmar+Ccn3KRUlQwFrs4qtNoeZ6Y93O6NHC
ZlPnDxluJowcK63UT3TZi+VR4a6NXJKuI8ISdAwOt8O8YCgE+1Fqhfe+5HPObbCwHsNgBcJ+guDP
3EVTYzVhCTk+tljU7hiFrY8y9toC75Wry4LVNEhhgVMS7O2GUfuN2YPom3RLU30/cF55kA6CARoS
xUyvpbZ2uBzEU2g7FiFcdTUfD9cijtxoHZxPlLA1C/iW2CQmP25AdsRL/3D6e4N5br6Zsqmr7R4z
pec9UA1IUjYtRDGdCMFivvpvcnG1f7S3AHn2sVDvtA4TpiP4o3E5wXqO4vJY1RwL4ONtNtxAcqbq
SN9KZagZujTQi4OTdEvPiWVeFLhE+bh+5PxApxHUttmHanlX8ripT0fqnsPzWF3O7ls154l2y66n
ohIB0oY1m57AjnwtnrNJcrxM05kBVapiWQjblpgxnpVdHm91OP6/4MHQoAi3mNhxHzETSQCkObns
1DpdnEj9on+BQHxtIHEpTmEVBxXDz+PxTrMeBXFv6qMEjGyJ8LMaMisw8cWeaft8vnbw+zQLFNec
AFnzHm74mcswOW5E7qCLa1DcEInWLKN8KTh7mSOrd2g3b0mz85JXamUGz/YBXatHw+ukmYZlH9ZV
sO9bmVlG6RjUhT/WE/Tzbi02Kn14kynSyPig1VdJkwLt4UMxXD0eU5PbmV1SVfWDZ6v6zNNtLAW7
z//ydmJo4AHp135So0m415x2U1pfTESFBjbzH4RWAczXlEifU5sQb0zLbgjPVkkaNI67JOc4Fxeg
86uslPq1jioqILEgL+wZ9HyljGGsGDffNW5QwAxaFiwSzz3zDs7VUiJPqpSftSzPLIdTbAT+Gu/l
SPjTh3HeVH+rhYq/g1lRDyCKbfSFhi+dPHOHbZgafmSl5BP3gP6WD045mYKhgx+875iKec8BAi7H
LV0YIMnJnsURC3pQDNOoJRj0Ci8rLneEGgaw2P3jkqWXKddFpEEEtw3nGqlPgPxpGq47Cvt0kVjx
wf4dZB//KCZ5LPDyGMncF15a+cB5pAjOJqJTVnOVhvcWWQ+3I+VkIhgaSlQ+JAsGbr11Rgr0LgFR
61EH0OgHC9aA8ueTvdNVSiERLcqIBIFPEuS05CDH0rRo4hrQlCl63sbK2Cl0bDHsk3p2AWtbwq/f
J3vYIMPhgD1TBYC9XfS33u/wclE58PaI5EwRR516+0AgpFkOh3BaNYLGNMlFk9kh5th1crbKvdX8
uGgwQVbpRrJ9w4e37rG86QSpOgMT7civnQDye5a8n1X1vewRw8NJudRjYeYns0foJse0Ic6HrUX+
7TWOWY6hnHXHcwkICeq9sAisr2EMAtuZrPhx6K21Ps8CGHpUWbW0pVUGlQjGB5lGqRsrO+bHt3nR
gqovxCULse8bygeu+TXV+wJesctegYmQQsqSgKh5jKkC48lnTVcMTeEli5q2C+GGl5P4p8bzqr4k
LKnb9NQ4e4ARskSWYJ2VvFtdfSfBjWtg7wca9U3EVo8/itim7yWRPztzdCly/nJRDhmqrXTEvuML
iIOk4imlOoVSq1m3bGaRIR0DuQcH/af2MmDxVHbRRaVAqmI3VAqp8OdkLZQKECS3bMki0mcc6xXY
Z4oRuFKTh9y/Gb1hjUZK1s/jonlVIvht5o7D8GPBMvyVVqp1L/HWdDsIKFBszxRdnEDSzn9CaURo
whKYT8H+NyTU6d+68A5YO7odREOP5nJ9cBspODvi4cxuIYm+1zKdInJIyrhsa2muPblf5opwkW1j
AzsKlTshSwQD22NdXWO60FTkfAq/7/07SWBBarlfw2DSUVMKAvjxlkf4EH1FN8DpCMPEbdVwEH8I
cksZRXEzUUyCODLZevv5vetZRjr27yAPjdx0CHImPKHZTCf9QraxYTY3CU8EQG9hchVZkRSa+jHJ
lwQ+eApCw24EbDb9fVntsczFVqq0hvzWr2L9mpdI+wVogLt5Y+mqNgSjvi9IHRkfOaPBBfqcjH7p
H8SNalkFX2Afv19XNiT4dqQRtUjTYAERlPiCVy82/N63zugEBb36y6qj9HoftT2RILME6y2/FwE4
dz9MrYQEehsVvQ+V+dnyC91E14igJZdZkxgudXXfLlHqgvmjfuSkWziQKn3exNfKduiwvBbty1cu
SSbc2thZIwLH9xg9O4BUnOVuUvS8XVOGIahPdtByW6oip6li+lubfxiHhsovPRNR3LdCI5P6GG9k
EAdIm2n+095xbLysKIS4hmRxGQ4wLdiLsrnnlbPs68NnGxoFbo/c09ZVywRSmcf27JupIRNyZxLl
pEjx/ufS0uGsgwtlOP/FwfBWi1unS3tkB8gNtbao/DcTKBzufPSorC3O9DNC8fdFGxdfhyj1JBQc
x8FhVgFpbPn4zLmWAo7Vdhr7HsNp89wkLK/8ChxI6lGHIVc+N0f5nkLVHkMt5uEOd8l0bplt96MV
Zj7vKmA3LWRW1IutglFqpjanins32QugOnyX95SLB1b9t/u1bnvlIq6mwpe4dO3MLpS5OVAa+GG+
TxniV6xjXGXdTlm17GEdSz0jB5VhO0mkZ4flveRGP3EzTj1IRigluzbJ85DnhzWgF98dVbZ0xGrP
OYNtLNXVbXecRxHhoTEwsNpxTjC69qcwhwWhvHpbIBRULlrhrDtmbEVfE9wd9iTdCv7sRBQOpapi
Hz9CC/jvMQx6x0c6UJNekbHH1G2mi7jf/K1t6j2LskinOg1QX8zp1NsQhvrrnyHsKB3sfWn+EDZ5
QnCJW8LMomUlPye4BQBqJqyBvj/92QISoh1VSlwXK20Wt7bc08+VnXQIDlP/wjzQ3fWultZX4eVv
XcHA3LuWeakTjFlN0rrALkBveEtjkTDs1duxnkO91wHw+6HfzbLirqSDTfx+bW4jezilHy40Mbrw
8TM6nZx1WlucVj1/8aqy8fsNyra/4hM248/83jDjRNuVlbAxBeKwCT0mRPZm4KPwQS6of9EYOaLb
ofxuel1SYeEkbQVesvazHf0p7edAVgO6NavAuDinx5mj/2BakSzOXA0LfRckWkTodOaM3e8+0sIQ
UG6PHVXWOwvyITx3iexGIzWhkOOqSIZgvpObwjt0DXj+ukKTrOrGLtUFdNKj4DCT97931TCkk7jg
2tczOqQkSdg3IoUWHsBqeAyJ9MDgJg3sABnKHuyyQ9rf4yFQhhwJj4w8aEwuOqVkELcSDcJnvf5F
qoHVVt75XfjclVgW5lQqix8E9KKtepRVxa5146BPtn4EU8Loy4yq5HF1gtreA7uiuw655mclmykU
G60dD6+TJgG/huCcEKeLF3BpXs+L1/duOgTqnMvAomZorNEOTzk6qatl0Phy7pKbGo7Dm5rsqJMw
P32zIb8I4L9RzDoERrCLaeqQySNNVe/0G5TJoLZ9YBtPFu/EEfQ5HIoGa48k0mmpugIYvP5Mg2/M
SQBvy1y7BfoiHiEyYmDOYjomi/TWoUX5WgbiQcp6np3+M059yJfTTHhZqYVQdVMDOENnbcreGFYs
GUVXvNtH7LUDpfmJO2+9/x35QxF5dLZgO81wRfx6pOjZzEVxF7Nf3k8rxGM+es2ExveLMsBOhbOd
70ICLaveV3fOAA3Nw0gDWp2b3SMjM0Huqby0dqJlxwsGUVdph8T1v24cskCYj0NuoHchZmnQ3YsL
e2pSh1P2tj3b1s2R+VjOvF95WPEu5g3iUSPj51UYAu9VaUexdhhteTJNQuBHBSStVQl7N5VjG8zh
+qKCqhVWW8YQA2z4uLnGHWtAT3JJnJ1sLpeDtcjcBOyjDnmw27JBlJ6RamVXvKVsPr1E7NyX3pEF
0En3LjqIqq+ijHTeSacB2hMn0lDNOb4E9haxoAnqdpW61JB+X0Eu+tcG2CzW0oJ8wKYGaASyjoQ0
ezlZQRoZ5FDIs4/GJ2MGPmUqYbtO62xM05wtvhaLoOpgH9zzg8yxD92046VTLFqenPNEcXkdbV8C
ATXLKPt2SDOzNPy3HiVaKj61aKOodee2/yCxzIcgIXs3jhppggc8dOhYyg8I9QSLQ17MnY0eEB3i
8vUDfm5T9uXrrbYho9vv16KDoh6P3k5IY1NiL2YthML1yDEjMYxEcm8844mDnPOKv8gDJhb8HhbS
yyFFsxFvMfu9ITABMqk+omqODsvnOEBtSv6GpLItjd7zKIqy7lSUp5gZNQxcdO2X7PFGFGyV9Pkt
jxx6rMDR80llNJkvNbXw1zyy6AQS6uc8LSnjOYTGrtF54j9l25LuySu57wa7iib87CTWQYNuDrJR
vmeIbQJTQIxNNbgRPOsdwhl+9hdYKsj66B7VgP+2xorOHmTeHwyl2QAIzSYQW9COXFfl49M7/pMK
On+r+bWcX3XtOKrFENaPl6NM00+LZ60Y9r6Cohfiq/IcyHL/6ve42ult4BWjL8ZNneqj4z/16ma1
JN0XzOjMK9Mj/FgqdCVTBA8b3FlRw6oNmGFxQz8ocYzE7UnO/FqFJSB3oVFhhAS8qqYKrQk9hvKT
vKl8gTcKo0Hp5tEjyWo1hAFNeZm/dpMIhfnZAHIQbWLOWp2hbJ+UMC4Q6A3zswoo1Y/xgl1hd+IL
25b7w3qmCZ0FU6ZLEfhV6PR2k5IlMv1NX1RJUxKHXgN3IFQkpx7E6R8rYme0HWQR3yukT4/Js1Q2
u/4VX8nEVF037Xs/hL12dIyzfkjlzRRqyPPtNSAywBn25AG7csmHkFibETbHWVOzutDqukJFBLlE
quy5BBJuUb/BbE2i/RVpomzaBIZZ/LN2XQSIYfhZVoE3SW/oXsfbCYYrKS0JYXMse7syQPQJjgjg
puR1QYN1Try9gQJnsW7daAHaGp+5OY82M5bBIko2/9F9cgmZPCF856jp9Gfv2YtINGiUJ8nETQXO
FbIXPZtMGSnqkMi1RLNDJql/YndCXAN/KYTK40+XwpHhaziUjmExsGlx5H7BIPNoWogT2WXM+aT0
MSrFDpxvfw2xpvvvllaVkicFu4/ixorWpDfqIFEMU3PJf0+c1a/Qn2nclcSAK5CwWia19W7P34Hp
D9vy15jgsGH2/HSD/nUA8uAbV9/duzWstQ+/CDclofbRuLVvH8Ey+LeYVP3Cw+YgDFDkrzO5+qM2
oaqqkPM4RMFo+xduxaNuNSGxqSKjugnlIBKNA6YjUHwZczeAH+TIZeT3Uvw5l/ZFMlbU/p9LD398
vSiPRr2a0t8m591xs+CmJF81TsEa8TvDiGzuawN+J6l3Ls8hdeanpCriDVqPRojO10ZUtBb0lQ0p
0Q+bM/zN71fd68ztTM3JG8BrqYnIoOFTQsgywVPaTsNdpuZKJzTLNMk4ds7uc41imk3raGz06w3D
z+cB7b5slVcgOagMaIdiE7moAFa6YTw/igtfEviKLsnvkVUZRaL5RZ7zk94/Zbr/jz8uU9wxDSvP
gi9Z7mPzfc6qcko5SgeloUiuG1cdJZ4eLl/ROkxjTA4LrLxJEbR5CxkAjupn2XNZvZhBfsqNI7hq
5O1/AL8j1DqK+U5YQPzvBKLbYJo4jT7K5+s6Lu7B7b/IHOsGVL62QlNy/X1Vb5+c+CgB8n3dFJt4
RK/GdGeJ3FCwrY96arCBcK1+Qg8jTRcKECZ6IOBw6DTE2rg/fSkIOAXp09EVRPomxr8fnrlmyBji
R9Ho210OxPeWO9eZdcir7lvlKfRexY1+AMQiNCw0irJh98AsHrEWLkgOc+Fzw3wwehA8SV0iI+OR
Tzw9akR9B1Xt4ZZrhE6f8sZdDl/9W4R6CrFarGaHOdqytztW/9esZuimG8fJ8WcC15NTfZxyAvl/
V+qJp+n1AwtQgiApgtq/rsMEuAZxXb1cXNorYbR3KWRL0bL6s6+vppmLSWT/frw09CyVYF48iJDx
Hxm7kS5nSNFU2eEUQ+8NM+mldi/qNiv/KVFBw+m/bDAI33osNDRHbP5x4/cbRNSVqFzjBAW6f/bx
mrUUsVkJWjtPNGd+rkdDPZsgQy74FDg1QxKh0GpcjsAlnZ8YfmFDaPX8a/hcbUZW9WoMRpnqBj/D
o/HqoZM+XMYkjskWxb95SHLCgSP+7iTtw/GW+P8q19LE9Apw6tUXpuJ2rNSOWlaRZvHmULxB+ta3
3nWfqn6YM4Kh94qD4WmEgRXYbWKiOZkq3MZdjvV6t/3TrkN/cyUALzAZxcCAzaNIjRVmNSm6IxLa
wOSJhIe/sx1RWAesvNVtTGRiv2ES1mBZRfHG+Tdre6rW361mAkdVI6qR7iMIq3U7uRIYnLMiVQfC
YL6ApV7imbatE8DkwDeYLJ1cZDQa5S06HnaD2WjgrraerEqfaw2NDQDa3COJIcDazw7sFDPkVMYz
k8MP1I8FGON00VC4ELXvmF4x4deosS+Zop258iW4z6mQofH/joCR0UzwhAUtqHWnFNcZccTb7dur
WVUpejxVAp7C1vtndvqc88n7VmW9D0WJxJYo+43tGerQXEwqtkNmiPIksPcLsjCLaQ1HwNtpxNu6
HyoSjkjQGnBlk6fiU17VEF9ImjEwvSSrPtha/pYULX1CCA6Ntp7me2WaxtxB+MwYSLynasZL0hDL
q9qSxH5hSsfQrAaJyohZKgC+3KoyKI5zuSo78OEjfDDdtP8bQg5niyUEGOXoLnF2yT6JdiYw7tZF
Q5/1LxXusjUwLqvVtGd6/owpfJc3OIMz/mIeTMh5Ayr6cOkAUJp/1cAV/nD6Zspen9pzuoo9iv/C
EZPgImW3ZPYT+Pg6nuuNycOG7VkCfk5V/ds+LJBhXAy1AO9SXj+Ap8PqU8k7wa3uMNgb6Qzy8Kwq
uveXNfkK33VSpiZbpVZSG4PzWE1pip161l9LViPtoFLLLpg/XWLlIqX1dIcxU0fRzHesAnMIwbZA
gzeqGNTD4x98xOpb59guFPpuQdud1UjQjdRKYIUoUhiTl6UMvrDy9XuoLMYwmyjMODBjj6TWvwRk
wNP8KMazkxEFrOgjutRkqhufXMYN7xSAlSQ5QCFi07ndkYeRV8bvczr/AyJ/TwHcSCxk4isFm3iR
oKGPmZ/2JQ8B9/mvdloY8VpYpocIrVBNraiGr+3imd9ZiiJlOaLJzQxXqia/x/gZCkWYZlUh4pAO
NzkctZtIL0/idX9O9i6uFiK2Dje6FtCLCZcVbp8h+qOaaz5BDutEtvvqQ3wftDuWlRY3Enh2gvN3
Mo0o6NiZh/VxHDEkTEJJb0rsKo3wqhVHjP2C+NgP/ywHdOO+8q64D3VMdU/lXVSsPES9Tpq7T6BV
AzvwiC4oNb35T85PwNdSGbOUthYrzmfklHUKc59eQnm9+XFdMBvfBJhnknJyIti9qpWbANfFDOKJ
ktFFkm+fs9zaDf92rlBfmxxocB4zgOU2QFTnfdCGImAsqNl++75mMRpbSG5Kr5pJS4q6EFSq0ifb
ouBkSsBVTbiXCXdxYsoEXa0fa/Fg9Chj0nOqvxT1BWD64w9PtwJffratQk/l6bwkT/5oFu5oXUHC
ncO+Ya0iOcXFddWWSFU9dRTWuZf6hDpB5O0l1G9LrBB8aG44npSmrWN2JdXT1zPy5lknbp8DEe/g
TU//Eje6ncjnlAro8ZRuzUGqFyVfKdWnL4ilMZ5gL2ZvMpZIxdPebA9XU4JOY5eHKLY4qnHEsSR3
UHaBp28Q8Io5o2bka4B38tjWUiK12DCGRndJwF3SYvE9Ahjr7JBSqhhd4wd667gFP/xBcgB7vg9s
q7sBg6PDBqFSk9WMPa2W9X5iy1oQjOQ3G2fLMp/CJRqeIwHR32vlYrk1RaocFH1qx8hokfiWC+RF
nKQ3TtahCVDubC0O9KvNbfl2s24GjZdeaPlivkU9HeuN1JD4tU8HbvrNikzPSqNA2x4XGnq+hG4y
+i6WId75F9Fa5HqqemvkRdeasMSbdntShEbGjyO8y8nx4OM+j0UP+we1qAq3ednwP4qmxrZgzNEw
koixPCwxGb0CUw+zgMKqbL3Y9JtRgeWb0rWUixpf/frtIf1oUW8s8XChkzcNTNirlnFwb6NDaDYU
dbClIOWyvVwHxsbIb4k7pNrsTVxEpNh1G6qOMdIbOg1vouJxhobZJTDMGSUL9/6XkNQ876T9Wub0
wGY8x3IXGSHyISkvKRH/9tg2QVwv6OLy8FYAoopaH9u2hReGFrBOOchMbgHzLWSmrxfl69/6X8Le
lQd7EeIum3ixXZMv18wugKz/DP15DMJe48M7Pco23x7NqzZdo0re5Mih4qxL1olw62PVZuDmChzE
0mTLs7IHhfXDQEvAH/J7cbQj2G9kZkSZOP89bZRm9CGBXd9SxTjb+0e/u8Q0eGbhtICOUCFSJWcR
W9+CcGCS+WAWlp8ieLaaqSbBMumdqUuKit8deap0hh4xUCgrK3YeCJJi6zUWWx9XhdAm8sySl/2K
zq9aX2zv2LhSN0qOGK1VZ7l3clf8/pqzCMxuzsBt13QwsGTKrzH1eOfB1pF30G4a/Vx3y090xVQP
zI7ghEYpYgQgxEPGm6UG99X+S929ITOg4KpDttzke4dQLquftVOcsZWjdQhWXGVJd2DZBC0X7rlE
w4RXBjAlJMiM5kWdcsi6MgN0yBWPNeSytB3YZ+pgiFDuU7TcZm8XIKn13ADkRFXT7H4k+XDSdE7v
VrKzqqb4pznI732AYA/4KB1CTatWV92UnsHqLDMn4U8Xw6M760YtPuwtKv7rAXl4nZr5lS0b0kJw
4l73B3hHrQfptCd+tWKgHnHvOyhKHettaBKifEPkqscOjV0EZjR2oEBCNQAIlYps5nAR+8Wi11xA
Rk30wh4EwGnLOQ1Ja6CINMk/dKCYE1QpIwEYpSqsaNNA/xNPYBq+4FbjXF4hrmUrWSlo4gxSkKCj
YvfR1OSWHrWk3DqpUrkBeZV0MNWkg3TirMA+2GAGgq1kt9IZEMUnh41YdWkIKchIRDYasOpXel4H
sU4a9+6F79dQf8jGziJ/YEEDbyRTqW2pa1RoMl6wC4xhqXw291+3UfU/yX2vl2HhkbplidFHYvXw
eU37bPIguLpqqq9+jkRFHEW+JGen4guKB1Cxc2kT6phTaw+GQzAjCQHG5XEcRDHk2xDpOVFc5/Nu
IVrE5NIbQej9GlRrSfwEsfvI4sNlUV/C8StJMz4Lcy/yIbmxtzeeA2OJTa4jSRye13H4494kmVcs
NvdBp1WavaVy6Zmh0i66xpkx8o5J5cVE/iw+8mAqbqCfJdlVaMiCgSyE+dfdGsMGYe8l8tFanr3I
d8AFCfu+uzu+PTPELN3BfNvWbm2MLsQIP3yzh7BID8o7/JbFlXyiKNdxxNgHfKN4mcewbOJqzmya
YmYk1E/I2QV5LFnf9FIYhbGi6V3QiA+oqS3UpBTVAEC8o7deQgTuAIc4hUFrazaAgj4xiBa/5Nfk
UOFjy3/5K+X8lxQvNolUs+DGwpUAitC7u8JNc0uQy6mgc2mLsEb1vzIHovYZuE+U3fkDdcyX45eY
oRl28zhpeKHAqTZkk2yZwh5RPNxZIHHUPZjzJqk43OOuMGQ2ndWu9Xemj5lid3cHBzkkuSsSkJVG
U1I9PkX9DHSkdWRi4RLWVfXwIDJNGzh0VYD9mZCDbRgamLBkRVHWsNS5BqajLpl6d/rWr8PblcbH
+WeBWtiWpoPAddG8/YjH5EwWu3izSEQAoI3uh2i/Dv6vk8muEHMb1uuos4IEGlAUG9p0q163rmhq
fqp/VOnbWkFNuupcn6NqgYLGzxRAByY2sEXE9MVrDFakNaxMh4Nw+InVHsxboaH8xp/pwVojWd5K
IMmcslP1YI5xff1rG/eWHJHIrnCJa4H/CXL3AjaitHCVzRAYyCTLjjJIyqnJBxRht5LOeKmtOEal
cFi5qTHgZB6CcEDTTn38rsumLLlKJtLl2hLLO+GaTO7RDCJOA0SClwdD4dbAEKpOOFj2v28na5qa
iOEwPd0eVT+Oq7UkQVtEYkzmQi58fpqfKCsMaK75ssZIRx73fNh6lE8z1C6HhCFPBgu1dstE6Gu2
/xWAvaGAtLIAK8HNGwy4wf7J6hdrp+wIsChtPzBFbrU3cnA5z6tmmaOpi9WM+dPNU/W9IT2v79JK
m+CP8ePegSaWEN1nIlDMW6bl6oGz/a4bj9EbQhtNLozXgvB+9t2Wh5PVVXMb68OQrTL6IHXWXIf+
pYVnJbYLMK5xFjX6vojtPAU5alZZcUFMPuKFv2e0WzuKmwj0f2CUfdmJX5MnMkVN5bA+ORNECHNq
v8uH2RgdnNNsG4/sevMcqzQ46bWXYly9MqzGDQJ5ULsioXxY407N179TSYbGwUCFxDv7vURy3Exi
AF8ndca/U328z6n8TGnoSiAsG9P+Fz8gDMlPKPtMtGMwjcbVsXZiIQkyBfqiz7yTz+mlzp6cVJUU
acbLDPNsendHpTOWCEmbUrRiwoWW5t80BiFr2ren/HQbwuE50D11Pd2h+w53uvYnkz+VhFV2sv1Z
Q0EMR+WxEK+M+7FB6YOMcRcnQesXe79pMANRW6u137m1auaNWfykX5+ZSaR/IPuWG7xP2DLRRaJS
dsiBwZhtZJ/B4PNePcO1elGQYgUpFIjxfeqOnKgNzK1txrHJ2l6YWrl+Gs1h+LVKhjy9Q3BYl0uv
YzcVxyTx0xXgP6YTEn4xnU3Dd/c43htP+kXwbGzxC0kL5APvpv2aiAohZtvGpWGiZ5t+TjPhg5ED
uDoKUIlLinlElOxdDJbxtBK8bHmmPe7UmdFWjb+EC069GyhlsCIjvjyxN17zRQ9bHaPkG1oSZfsq
KOq5u857/oABOhC22gCTxJrH44YIP4LntlQb9/YuhH8m6Vc4wteE4fVnggTgnqkZFdHetd0zVn4/
P1M0NwMkbDYC0gEV4LvBfP0N1CvLssseUlhfki4HZaLgVbkAIoIz9oCIZ+GHI1/xLbZmImwNf3BR
PNAw2K1RSN6czoVejwNvufF6NOEp1m2yvKus9MfJJIyQGP+g7/MaMQuHsZPZBA/rkHwhq2dekPar
SxrbhWhvpxZ5o9dtHfjEz9kyHB9bDDOt2swIcbISnM1yjH77GgVIJ+lMd8O6wFYn8G663r6LktqR
yStliux+tsZe3iFFjVlZxMJaq1Jh1CkWvFdZLvWdctrEVWFtV49Ml2BTTPAOfBYcAEqeD3Y1IQ/K
x/yl/1OjzNoaAiLWhsI5dTF/p8IKtvtqq1y+vqwrsyfK7yQMV8BpuBrSBzs5Xv1G+tA37uXJ4vMI
hjMMgNTo21Jtdp4MQvtVp6GqivM3L+Vl33eogPa9KGfMFj9uTOZX+Y+JNomJuz4ycGPBW/uX39Y6
815ctcMkbKncXGj+3RENJAqfoC3KoIL60xTYV1eONJEO4YHljG0R4bjpCW5PMVx2aFTb5osS1F6i
tzEI3KjpFr7otIfGyxX6h+/uhQIxASk+AwWk7F27KhFNEeESNJgkmpeLLVXWpynZKo1GDyrXWU4K
w6VYuaCXE07uptUes4nfVfIOOX2lE7xkNccuer/N6kYMkV6AABnGbuaAPA0o8R6TD298MxWAJOdV
YzeeiK0QMFmpXx8UYvQfHV6U2Pjaq45cC9K7BCYW/qKYOl65QfUulY+SbcMd2L1On/R6iO0tByA2
gFuceD1F40mlopfw8nKsD1vWW9k+TtP4oLojkUzWCyIHfjxqLN5+8dj5TheIRuBZSO1bsLTW+1PH
6TqGFgHhXE1pK5xQS4h2RyZNmwHOr2S2BH/8Ip9pbrLYzceRcsZsNqpR8ii/vdrdBI/TFx8ZML5b
FVrbsL4sOer4qB0PVeIywogwZqmoCjKJaEP6PdokeUQAQzu4a1C4fY/7iUwpHGkTpN7ushpGqqt+
yN6Hr521q3QmRrn3LPrTY28QgjAZ00aHSoSYVlMoCTA8AnEUn3oF1gxiNcmTE2WLz78JZv9Nubif
xENn+EcamHTwyAb2VvVgRK9pKmgbhUeTp9yHyoXJbylF9tXuaQhV3++gRbaVSLSCj5dA5X4sz9n/
Vw4+/YtYxM3DQDxa2E7MEsVEZyhL4g8cijrbS5BNEwDhOhAp7AESbKOOmyxznbWf0xdFrAVaS8Yi
2+ig7ff++N/7zEPbO/R7Forx+WSB3xZURmZTA3CFGYPwDCjtWKXsgv2JHbGKxTbqC3DHjP1AM7LN
hSniwukeZsHzLY5wrntrMZfbtiV19Y+3nG46PBuyxCRcFGvCCOM1+X4TlJa0DAp89u0dlls7vWIY
3nT7h8ESMCgFWZc8KRmkUBRE3wtNDejjqBX3nyOWFMT4z3F0/BHS4SVRF+oOje1svjaiE0ET+DSB
1MUtS0wpAX+Su9kD1aDfnREQEpUONA2VtNfUGooY59rjoGQf+Ta1Z+FrGOrr6RvmeCIGQ1km9TLZ
K62viGOR4Fbt6JnU5c2lUX/kMY0heIvgzr5Crlg/gRSVn/x5y/+6Mey0koXMW1DWtFnw7F+xNNYE
xSZvFMrSToMhBACu/6WrI37kVKge+n219QFXJskt9d+7NeWQMvikql9UoXjJMvxOANNadevgZdT5
aOjj6G0IRRGvuQCZiYiCKwrRMXXmQZdnMbbPPfnGv+spym0OImtwaGOxp21IMG8JB/9IeHUuxSeJ
QQKKBQOlqmy26DMebNFqfx9gYk2sIfRhLW9Ur12Ss17EBMEZXfmT9tkf6K+HJ3ctLkTWNN9/gqq2
D30RY1xHVOVmxdmYZpYRQ2soPu06zWCWnTbqenh+mRABxcmB110Wwy2jT2Wz9gzpx2XJEhIHQVhG
Cj0S6+YrhI+CMAthu/VWAZL2ccGhuAFf9l8PRziiBtpnFbgKSAbleCqBhrSxpHTeYLEoSHgEmAIe
e1vvpqle9hYPJ+mjBWzVmaJ269q+3ORPR9xZyik5rMVCScxjgbRmV7yWAjRz4EeIKg4QCjZha+oA
36rnKzLV4HOIsFXBpRa99rb/85PqLJSmZYeZ8io3QoKsmYxOEuZjvhCZHMaVpZTrd/m/l0F0uzYm
2Xy3vKz0dFJATwFNEjjJ5RKM87jpyQHyxdegAXBSHbN0FtVckNXshV6X8ozMkhXnOPeTHZgawsSn
WSmNxc5BF3cyzFALbkYL3Hz1Zgzj4FL5WpEo22anCAuESg+zIo+av3H8ukUva0ThNts7kQy2vCf3
uR4sVu4AgOD17kRF2YHpFOyZmcrahfFrTrx9vr1/5/29ovvunMWXl61Q44dTw45Igwxz6aLDJIpq
3SlcnOGgUjylUJZwy+ND90qLaFIWZOOhkdEQUTLhZpuXlx0KcuSZFuud70O7uUOSvInZOuo+0lkz
JdImn7P300+UNF5WZquUIklaahiyUNvizoUS/XanYKe9jWJpQYUYgF0jKd3exMZRg4qL4K394D2B
nO7veh/SM9lMtAFumkRX13F5xVgeUac6hsai/aGpLNJaLxBG5WRoa08qv6BAkHgGk7qojsYedcgf
pSdm8zY/6rE6xifN99p3mMAlAFISzyox68RMeO0+mgMw/afZbwwf+kgGefHLUrvaqXDq9k1v0HwY
Y9eouXaU7HPhpxAmRoR9XlGYdeinRIS9K+y5IQyX4PSviU22PDBgfkuduACTxZPPV9cQWDYwEGnD
Zp0ggWRjBrmg0pFab4MxaiQnLiyXi5aqow3n0dxL/vMOlYFsomIfQdxHMogRGtM6qeWIDUKKMc+S
F4+BjY4rrevjrPzDXjNr3hQdC5bY/qxYOvThDIM62HOYUAow3ziatE3Fz+l2HOShYlKpcOiqr1gk
yBvYyzTxSfBZ9Glo+Sry38LFBIQHwN+mQFSu0LwQsjwbHss3fOBlCa3dRYQRyFhjJgWFQlt9u4lO
0+9APMsj/lKbShBF62edNC3PonXZwlPoaQalFc1wYf+kyQP/kKz8wzMu3sSq8o125An/DZXp1dNr
cWibMGVal3UIBU3qSvcdvBogSLvgHZrsJIO/4ZLyvDvPfk7cA573vpEmzSftSJ1bxOFyBPUHrf17
CSviS/1F0vCnMihv1OwDMdzTiG99rYyFnwnaEp0fzlf39bwC3GAjcHEBqkJcPpKO9T3Gx38dFIln
uFk1n7rViXeSsFIMhnORPRUCvSh50ncBR3bDnXxRGGDEs7WYRhF5dv1E9RuU+QGaonRZG3tMAXn9
bnRg41xgkI0BBwQo8X+DWvGUixeOqy5mEtmsbFuzufaQlJRU5vx33DxJ8FBf1AkSIm1cp/KIrq7z
DaL/D2woH6F/KA3UHtdDyQOolYuuZVbf3tuHGlJ4MG1cvfHEexdTiB78PnMSHcsdVoZ2N+aRapOg
KXDxD5gcyGAXAgalvag98AfXDOK7YKDevapKhgNycPZLxSlcEeNebqLMWOfGqpv//V+GoU/inUao
ykJZ3bKHOxZCYD0bocrPCKJaUB/PHWRU3HAwJrbNFv3a4B/zkktpl2AM7s5ZwMN8uziN6emZF6vX
Jf18BmMVA37kNcZyXvZO6i/kPvnp/snJwjguydpxr2DnPRy9bzWxKKB2jtVm+GaxQg31/U0YwyBr
3SIAJL2TMt8xHFK8lmcH8f/HUqz/mi/f14BlDMN0SmqPMSbMnYrCylny8DzDSbZYvw8oP65qOe6F
2LFGWh+9JZERP27PqD5c6zvLkUTbDdcH+hKLYbqVUss6Gjms7+0Hfh8NhDjkNx7dv6FJrnIByIWl
pOkW4MoNL9AfemqKXMCeBJomiG39C/FuhJEdjZaZpof3nKNUh+Pn9FDJHKbTTKKuGhMhGKHVUC+O
FZiOzAJebMAT9ddv/5sEzQGXODhg1CAfZcxzMoOm7NEfXtm4yEjHf+kYL90nWOaEVlNrAAAv+Eaq
IcL2AS6iCtg1vJFctLpk5O5J9ujRol99Hzg1Qhc1zayYr55Rd6tq1x/qAjNsm4aFMU0gSs2ewTGM
+5k5ur0Trqx97rqT2eTyYX/HwlKnKbn4QhfHN8fcpNlUTV0iLfwCozTp1h3H+ZIPA1LP7hAQMwnA
tU4ZyURO7Rbvx38/8iDWAo4GwXPu6spVzZ4MzqotI5D6NV+rULvT2L07LiVIxDQYzdQtrUoUjeKb
RlSWv84N3QwrhG91u6k+JweTRmKYVPRV0ApZxapqA//YTJM1EqeOWownFs91jgKupsTvr+5o4Wb0
dINJmg3RXAzImoeQtgiYKsPFZT3bNpl8g8Op91MozJW5p50arYI/tBuz89OKLSjeslOgxFuIMlw9
w2hiOQOSYrZHtzkN2LLVOUv0z9cwNdUqocVjDcxFwfdbZ9Av2hdMjzjQDwmV1h+OZ30bFrKr16gp
+CCkJDe+F62GCh5X1rMUcflWfdQek42dwd0Ni4+WemQy14BciqUue2sLywcB2GZfN4r2jLjqza3X
WJZvy0oxU2MaU9bs/uiMZouLqfcSbLGARH2l45TDpJb/8eDzCet25/1yDVN4iJvnqXicnr7sgvJa
QVy7TOWm4CmYPl7KxJPaeSVBq6tTib5Nj2X5M/WHLCD4PX1zFoYKuVKs+tK2qKdAZMjo4hFmsI6B
ut5g+lUnqcyCOCuRrBWgD5nFT/NrlbudqnzF+z0jv5rYoeqv/8Ewfx/C0N+9se1Mo0Qvw9zCEPaZ
1n1ylOq+boxU7yJxVwk8qV6vWGesbggEB0VaDsGXJHZMVWPr9t/5VLomRGNfNoBAc2IL19jidMDa
L3vhJT9fDtRgMO0/PMmaOTcSX9DoEwE65XHJtfMkpOj7zvD/Y1iyXRwJW7IDK7ogUvDGYGT/tkXW
ToLT+WUadEm1bGje7RA0thD+VuKOm33ptdAF21JRrig6xT9sOcdQfvUUP0n3xmPmK66x5kfQDjAG
SladiD6Ybm6VlW/mZagJEvN7QOY9slqbAq0sJyng3YLO5mk68rdars3flBcXeqb1CtrSYlLDc3dz
HxJG6qsqUbEeBkhImgE1uHNK0drQGORos+kgPb4NesPMCMpM2FWf3IflCoy4erv9Z9BKK56CAKyL
7DdRooHoIq87QBSYBz/+k7LWLRpnjLX+ChdNXDHcvuzCtlGCuSmCjaK38k0S+BNA7+qAtypAAy61
zIVYpcmMRxxf5y9zhiwZxJKYtNV2TEhZl3nYCfAlJTd/bCQ7kYx0naR2KV3VNEIxBfW7SqQl3vka
o7GBI6EbHGAlMrJnpy1PWMZnKd8ym31FLFR5q5teTC8QRpgWwHqc1QgbgUE4sgnwUbltCsNCD/1/
mzNozedxxeEe1RVb4I6BWwWP5y6YJhI00S5KBwotk8N9qnepl+Mom7Qmp8Uu5aVOqQ9toUoppUjx
jDDQbKy17tLj4UORB2dqNezgHy6//vHqAQzrZPQThu0NP1V15yJZhQHPsx/0JGcXmQRDQ4F8itv5
tmhU7dG6If7TcPDJ/JKQXt+6ljR/aVZk7ABG01oPqtJo2dTPjmTVcs7i0tVAslwnHs4GOg5u2GRE
7JP0I4eZv4+186ZR5T2l7U9njmE/T4Zq9xUeYA9Xj8HbXZvPVQUULB4gwwzFMcFQRqbPgeS7bpEi
/taGTd1rYUfFAk/wc9bEkCapeWDEhoB0DnECLm3Fpj781s7tv66PheZ3Q9SZi4UGd5UONZYqRZU8
v68CWWkd+VqonsvnwH+BBp6jnbwP6wI8A68Z+VMrMr/GIUSzYGsncb8O/G1Yh8MeAn/tlhqS14kD
OVU1Tfy4GS6NWfWFma2EGjTd8Vn6J4ZkTy4qeTAgYzEqvO7SuP4/6H040feIj8xep2YlhIqFuGHD
XlcH8NuFVhmc4iQxmq9VD07NAOrGDG9lPFAWnk3U+GJqTK1xxx1UJs9PsLXCxBWmo9ZQOSJK9/P6
ATiu4P/oYcLjc9WrGIm+tB/WYSB3Fb63Ri3S8ybNzQ7uO0WqNpvlSSHp0gEBCVDYksAndfkWL1kj
m3ivTU3OnddEOEnbuZFCpnQj4o9RIHslYzPFvxK/FzJ8FuJRdupGR8lx01N4sN9JrKT5Fr+Hl2yW
D3D7XSmytdFGduH098L+OQLfyBeGIq3yzn/fMQ7Kruc0wwCDqDGaZDDD6psdHR/9MRRj+S59haNX
5SyKJ8Tz8kwWt00GyScKoFo5QA+L5mz3EbuQNwzSGHbvsoDEyv84JJUziEZURU6RTxE9h3yG6At1
rDorJG7kE3smXz5KDF04u8vbohRZOgRFMi2MPI8KyOQFczLA8ISsHsiDrMGiiAlji1JYabRfkV59
CKnayoJKYFyCuZzu+ZCxJuzyGCZxwGpaIYZZT9lXh0vztDkn2BZfR7up0ZOA2qbM59oFIIL3w33F
TFeZklP3jF66b26nhAUV72pUNyPjKALaQ1ObAMG22/zb/K0wLK5i7A7JaWWfEuyoTmV5wZcy4VAx
lDRx4ssdouls7MVIOt4k+Kg8WBPkqdSAQdG79+krtSAx1YZi19lcHMDttnMsS4G9hWVqY3OyoDT7
7VALk31mfsQ0viXRdXMgn34eOEOd8LeZyo6fLco1fq4dqSJilylXV18kNn+hyB4sgW3GO2+i3Bnc
1GJD2dFaCIy5L//Gl6Qt/xvQ6gxGRxRgp7NRiA9rGSMXsqZyAv0Wv621nJCGSH4GEAxxZy/3s7eP
0qic9X7d7eAhq+mmZNEKU/RK0qDB9UWgP8v/xGyBkTVU1TIoTso22yMqJq/4O0V7Cph1x5ezg8Xo
hVQHf1rAx4arPYGyeWZlyinBD76dvnBgvl4A4+4hl0Fv5ZQUrC8oT7grqHqpWcBOlkMaqH4GbTrj
nR0V/VhhnrFNB0yeZn3R5q42H/PswICbKnIRYlqCchVH/IUDPIL0m1yigaV0/NAUHJhvqIQFYCNa
gzXNzCPcNZEFs7xGpQMSFdDzmIq+iD0rhyChhuAVS/QyLLwoQnC5pUAA9nxFxnkSwcKQJsCrqAjc
cZ5sevtuZz64L7ujcwG7oe0lYaca0why5QZndHcwLMfUSapq+5iCgytTbtWh8U71HsPiAbdD7i58
XWkGgwM9zZlzWcALdWLL0WeOol6xE/ZoGxbxYqSMotLtor9C1VLpw5boD3UpuFIdcyXzDvjCUHWV
BSw8p4BjTGNbA/MJpGJQ7kPfSNtER4EKBFgVSHwvJD7mpnMu482RM5bdk02qQkQwK9bgQm2pXYE7
fsOKUP3nABII8h2d2113D56Ccem7MEyH24Zp5F1NPzZ2Cch0GEH/JgJf5RUJDluV+y9cULgQbSbi
RcqKT2+WObcZcUsN5rIAIXUAe3rPyOnNDNkc/RIJ5uxQw0kizWfM8GpJmRppqSaPO4iNNqYp23pf
XsiD7NG42kH5NMq8dyiCTMYwKb7AzUkZAaWgsKznfXcHnGOTfJ+riUr6vO84q6VpG6SUWo1P1rZs
hMlJIhPkxKfO9wAyI1Wo1kXdfLmS1PEqx5aw4qGYdCvFNGXSXzo+lz9G0qMtU77QZH4WbRxrdfp0
uNsUajwlT+pQvum5LgtF885CGkWCs8gTQ5eSiDu9ihhHOXs5me6Kwr8PalNeRXNDpca+W9itK3DI
ydQuMpwsFhpPKgivLZ/QluIGIPbz1wtjYUa0M/XHqryIGW+6AkcnMod9uRn5KsCFujiyapSGi8OJ
8vIJGLW+pwIWYkAGdsiIRSmSQ9VjfrlEOaechIxajz7qJPiejR5P826a54iKsVvvBdYGCe73TxAS
fAfKhQMHXlU04MkfWHWtfmmRwqTYaxPdYmIl4SbmnDss/x9yr64lfee4+b8liRp8Q9/Su9byR7OK
TU2orcx8f9xLMNBuNln0g6uzoD4+nLkdWDAj53yIFxtIEzu5gTEfTtbZ3ir0ZMhP0gm0vB1fal9e
bvWDGJtjXjoiNsPDXPEzH41TAyqrlgJGUKZJIVtjNUD/AUMYROiRAiqAHHU2c+xg5DQY9rxyl6SB
KlLaHMfONaJQLIDJw2ZU2jVO7B2MdJ8xt1mWT1LNHgI5cFmLNdPnuJGZgnXlXYz0l8iHemaWT8yH
zSCq8znm7xI+cIvmsF6pRYnbwUYei4CWAozz2cLZlrPNFbg0R6OGhpawXkpRb6Y70wfxTrdNTvOU
ZqC7WxNmdTF2OLn4ESDTpTHqBRqgbSBwmTosQmwSXWaSzT6Q2BV0xx3ReDhu5CXnTDUjBglmdjZP
PBRSYkme4ij62nLrYneonMpiE2l/2HCEVQOvRQp29s1BaVnS98wJiz/iZ4TsgZ69tKNK/KVZ8BoQ
NGizNboltdXFuwrYgMOS3MzQYhDjMjAVZ2ekmMmXyu0+jc8lvikVy8z8aSu3yw+FIoUP022qNKez
VntFd2wZYs4R+2CXfIzv92qJL2pQm+QojaHk6gb55hUJwfzFbXGZ09oXLcVBMa+if/sTpN6v76Jp
Y7BXhuYd/+J48ebUZHxY5gLbb2gpEw02U2MP6qNOJDBTYlb5rUim3W0bmeZLrR/rTbOOTf3VY+Oz
1gjDpHFW/meXHikSeYrxx02/NbcNH86+KLATCzMlytu84UQdis+th/EaRRAUUPYm4vfK6qqHzEzs
b5XIal3BVk0ktZSt2tIxFb7ZKvvZImEgacyB3oIiImkSl1p0g1XdZ6iRMhYoECUdkCeocM79cfAJ
qNUw7w4VFus6A7AkQg/9PlheEd/0/zKfkiJkPlriWAGLAOh93lG3zDSsB/h/Kxvz/hZDjc/gkPbO
O3qVqjP4uE/VVsJg4jSXATZDwZrYac183Ts7fPaUrGOfcBH9mOW5DN3ey4oTxbHUu0lcX1N3CU+e
Yv43lsD9SVTHHdScXVW354TofoyqPAOoiFmpSXjTwsko88QYvM4oxR520TYmD9aDKO5xpjE/0yN5
yNvEH1/29V/r8XwVxrTzGtadJ+jOlnt0/9NNxk2Bb9pOAegIws0rO26qFMoJpaMzRwr7F6la5/cG
73fqFCN5QGw0XBwbFDf8gXmBjxURswPeAhBxI44Mc60oNLyS1oonza9ZOyIPMfuLlKYCD+wFh+Jl
5b0wtRt3KystNoRnfZLLw0CLVeQv4phMMS1HtoKrMLJ+K6v28FLSaFWltlmB2GKUMQB0oqh7ai74
7Q29Bf9u+rQtLN8DBhF8kZBtEDF2zkUt5WuXY4Mc+zfRI7swosCvWM2yJdRuV4m/K2PD5cnwXJb3
cpjYBQZvm21fE0le/0VzDY6H9nKQM+WCN/3JfG0LeISqt1h8NeooaWpoWVxEwFhu9kX1EMmTQwNE
imah+MJ7t0UURqsa+5WEaeHGrdcz6rINP77KrKA8Iv12Nwk5QYmK4Pz630srN9f9XHYbldNi72El
pyE4b1R8/ASMRCZYhNLJ8KCDFgg5WqXHGIJAcSjAPtteKCnsUzFN75H62qJns4usJJwOgbXdicEe
Jchp531H1fHNNN47Ljwd84f8KsILWPk6wJIqMF4+pnqxHB1s5wSzYePZ5cZi5WZz/OZr+U37VyyO
Du/ZvLe2W3HapBGiIXlnZDM1IHvdypDIAMGo203zIw29/ero7EdRhDs5J0Hlm2/satIJwYyP3OTc
h5LHQ4Qu+RVM0e+uST4Y/YwhimP7VXy0OOgL0tiBxNk5B9ZbMn4Thb7xdVX2PBuLKJTRGNe9qdRn
a2ZFzS76nKABRiR4w0iAaQGabYQksIqMgeIo0B+inrFZz/VS+8QSQ5w67raUrSghxcAC/aeOilXl
bQGG1VkzTzA6Dw18DwLiL8sOTXZQe5YM0m3cHQfJo2/wJwzNoSn2Wm1/CFl6bdjdawX9sGUcVTEE
l63wcty0AfHY2KeDr3he/3LGgME2wbqMFtoIJ7nHscCXOeDRbs116AnF9NjKwUS0zTiW2W0BCp2e
G8idovi3EjUeyq2rUXemcLaD+u6AnaRu16wdIZEfp1r1bxY1prsXPksDV01hxJY1e9b29wVfd/Vj
q9XmAgeHjFXKYH8Mo8IkjSHNO6NfgFKLOJabDaOS0+GRBCL61hxXehCUo4W/R6udwrjBRirvoX34
sPuLOiWtwb/20bY/9kGSSP0WxomvUY6PD5TCKOH5VWBrjOiES22rQb8XT7h4sySbducI0407Yk3c
bJnvJ9uYI6aR88Mdc1qNdcqfkASCN6myT1kJxwYc/JOzwLg8kzCTMSzlVkN70BTWdBTg/TH+o5SN
C2orVSY/oz+Q/Mtfc+EBdgcZmfiqTR1qo1veZtk8ieytRY50kPtF4xfQjyuQzQYs0H9fSS5LhfPF
CUMrw+v5qqR6x5uzCCrSfhwg1ZE5Q7wuVU0vh1FSeFQ2Onqdgbnl6ddsKqTazmIic6WvKK7m2bmG
vRoHXR6yvWz0Z/mffnumlB//jae6ZIV7olf3hKWJ2nquO5Pb4c6ED0uy8dMYM7W7o1F8sDrsPaag
JNeX9T1+R/uOxKZdntnF5rDS3fn0H0S7o7ElwGrPd9HXIp8fWQoeVGXt/cxC/RY3ko9d5Wh3dGnL
4fNc6OOiW2LYzJe+n1NTXUYY7kunjsecieHfKuuEWTPNsGVtVHjid0WtdOzqeQQLVyUDEvS3bgF8
YNBJhr04jcOTyi4NPuzzJDAByUCaiqupvCDOk2F91fsidDbNdqbehPbCuC+Z4HwU5MhHdTsYvJfI
Rf0CjWhjzKxyLu3hBOdGhRGcZYIo0dF41pblqBMbxO2gASvs7rjlhV3YGO7c9PEsyV5G1kIKeYrj
AmaAvmnZRBLN+Kdx7z8V3Uaywnb/G29UtHVXWkfjIrGpTEik6dW3+I0x15mQRIUHx1+9xjrQJP47
RMz3OYeyoUEw33PqIsDHNhkxmSiqNrzylYtQbGAnyHFBQpBw4IeBTgGe6pX5KsB3ZuMNIWRMzenH
Am7UoFN/4JNol54sqR+t7HrMiAZdnM9i0E2lGp9OSzOplqB7ibVRDDoD3YDd5qzF+JPWLmOlr3sD
qSXiVwXBXE+UPC7HCaGiwMRh/TzcAOs9axeYucPmMvuPeABDkYHvv32kfRjz7It1ZPJjEAEowYoS
TszKjN0MaCcmkN5Ko5A/TW9ujsl8XytT/+DLLl6h84vwiL2dFJUJW0KASnwJkpMuB5dBjcH3L8Mx
IjEj0Colb5FJeNkjprMmY8dXMoZuH8m7w167quIZmDsh9vBG8wbbhJyGjMBdUIgb7TDXG6qU25MY
l5zbhIqku9EpjvRP8vh3c85riM/HgCbQLZDYVSMBcSTiShwUoEDqpmZeIYVzUy40elb4Z+/+OpzI
Be9W+DkoNuwvUllFwTCnnl5u6PfUKZXH8TXxQNe2D+6c33PMh4y7UVvpHhhoh4cRHyNMMHJSz3dh
txZarfiXT+khyBHVAk8zGS7gMplMudyR6b1m1SdhFzPU01i3te9WPwyqqe8ToLqTeO4KAIi6JI+Y
7C8LzX9SswPJasqNtgJJJ0zuFVrgqyRLMxR6GjpHcz2UN8BdQmeHt4V94a4g4/7fYKPdxv8sSqvN
IdnU9WWaN6jpt46Xz090ykaTBjP6vio3hYDPtM+/tXJVSOqdGj7LhRwboF6qocQkFxqusql3QvTE
+ap/mPFERGE4ro+mavR7gme+FZeNvPS2N8pLnTFGIzcVxx25PBtVjpam43dOFaHsd1oWVlWf1C34
wJ8nJebhEoRAAPwYml4BbkdVkJuWTHUDWBnMSFALqqIMUhTuPaqoJyGxc6HqAgHH22lc7uCJX4Og
O1BJgPgg+Uagtz4O4bZAMBUAii+t2PBQQPSRs7AWpw+gu9OUDqVD7xtMDSs93LajPY1zHQIWH6dR
PxH6vI2K3nP9sQiIYvYOIHrvysR4+asFga4tB3FulnRjaD4AUWAgH2hp2DWVd790fqLYai3FqPK3
mlcvO5WAq+txHNOz+m6pAgfLjccJr2qA3/afvvsbc5uW26fGdjRTbwXmYmDzUN22WeppIHU5p1ax
g4zbbAb+FFKXbqxK/4XsiE0Llms5wUZetZiCRigu6maC/hdX5xWYFuOffdj49j0TmMej0Xp1/9eL
VzQ81h7ZDV09FF0w3ccaW7T7G47FEBi5ASwA/dCBZ+gE9wGAdYnpgygJ9sH0xjZZVhTYXSXjdFL0
afO8v0J2STAzMH/iWhauh/UXwaLx3GYOw+BPDD5kMWVN+EWUZUX6Zlw2tkEhiDQcmrcLDMDcTwqm
y1HJnY+YJLj0iK5jJ1M2Dmtvb9XnDC79l/ZSzCOBO4gwEH6uUP+bqR5LLejfENltBo2znfZdQlK7
eXiHcJZ4zGLl+h9yZub1b9E3TP1/kGtdasw5IIKmT8nLwFcepM0baZPLvcoZ1nD47XeUXyCOb64K
ON35T5mZAmRnrJM1i4m3Lrmxc/Fmwv3RZx4LLJzkOQD9ko+ELO67PyDTYExzxYWtFgRxjlmLHI09
NA2TgV2Ltsj+iY843T7OUC+/t1RSLsAgJ67aCYKUoLkxdTAcwUBMIyE3slJIctHydoTp9o5K4ee7
+bZ4nJ1feZh8Tp3jek0j7Km1lHoufJUTk7368fj3DFvn1sA4yqU2WiDAyEvHigxDNgvz1j5BCC4E
Vmwa6az6HL6Vz59h9Bs0AykYaH/C4/L+/sOyEQPAcOTPx8veR9VWcIZ9tmyzFnw+OXBqUeKvBVqt
8ouP3QAhtz7UvWgD6oxCObbTwFYrd7+dW1gsXrJ7CzCWiA6vY1QGD0ZH4Gz1OEwnlzYnAEp2xT4O
JeQWSCbV9SIeP19P3F6cu/A3U9J6G38joLVsN8O3ZkgdxRxG7gHSuOliHACPREZtYcNfz8h0aYXv
1+85ypavj5kV3e/EIV1T6D8nbHJ7IiAqbceJ0Rrnssz/5+QOJ1sl3iHtOO3mKQ+7+PZ4UXez0g5H
UJ65yAWAgSz4aXeWD+x4zs2NL7uw6mgoOZcIWLspT41qdaHsCChpvxuqgSoz33yCQ5+OqCR+CYt8
db18GcN1SlbRBvtHzJFxDUnwi/0M2yEVrowIzEFIT9ZBglMdOH5lWUSGBHRoprI15ygwAcE4DJ++
lQD6Va+8TEXm1vmBnCKGv16HhYHtY574MPt34Tou+aaIZKe9AMVHqTkpoTLuUrkJfQ4LUfYVRvUV
wY4fORSch6X30TaOlK/tufJHznStH5U6WuLK4VK7I0IuQgnWcMmw6EWOaS6S2HZ30ADc9RO63wQ1
Olk7nYsmC6B/YT142EE9eRT4Qpf8bh7iVsRQ5rEThjCpuMlLTfaemRTHc6bUelrm5Do4dURmAOYb
TIB13nFlefaycRuPPsm2045V0hOxod9f+G90302PywxXTlWnvfiZ/dYHCJwgcYiK2sv66hI1p44n
hFDxoJXRQPnTzhqxBpzkv1JBf8WtxTlg+x6jKKzu7nQp14GqJHa1B5v/ezfTR9CeMVBrz9Fj3s3J
QV8vRayxCUw0MpLkvo1qRHt0skxwr3eVMIeK5DFpQ4mNlbMFrIwCI7iY+YFxmWeWYhzxs8bmyQUA
jJgh8AZ43Ifg/fGaHA/6qz+5gDQSWHJn4STk6lbb8mNRjcy8Brerm+YQpt3ph7KYrxMTiLhA5zm2
s0KY9QOBDvt5sW3DL+NMmz99cTEXnlcEM9danQimZ+EQoe0Oq5+NAgtfk3PNJQBAJBPDDrRsSwoo
RqJlKCVPdbXAoF+3XgV2fNKt/EL1GU0l+HUElWGjvUL0ljsm/hD9j/ooRl48sapuwHfN9jlhyeaV
q9XU04FPJkO5Xwa8FF85pGu6KZz9E7O49c9BtZj/F3zyeOxj5/9M73fPs0CU/7WqQmeTom/8a3nr
JN2phca1FqksxNMQDAyZp4ogGXe+wFjhflF1AG56ocs+NwqMSd6aR5b5oYoqdVYOHRelY4pyp9cL
iv7ZZrYcZIjchqZxy9Qs3MKNujLkUiIyr3TcYWRPfL9qNDBIzpF829zMPuA3owiRZq55ChhrH8Dw
3ZhlSEctAyAbSA6H65lyuMPY2es/Q2t/Nrivu8Cigsmm6cdrIXTZTbX4eBzz0Z5iXhaWqGkuw56P
B29hxog1lenbJaIXc9kp+y5JwwvtX8vGWcecFz9pv7CO+N60ACSZ99/cTnGIz14eUckJz+2/cYGS
mlQaWkPTg04FaA3K7+6duBESInNLU+mY6hxF94jXi6iNA/Vagd7MIB/FNmtw3Wcm379SzytnGcxP
Fd6ToU30eS/c1xkH7l7Vu9b6+YUWx9G8zv5OqxcpcrBT+9/cEP+IYBe20Fag9DysnwTplw44wz3q
fgEbcPYCbA5eZogg6pPph34lE2DO0Hg6foQlFiH9ByQg5hMgL+itOaZhEQmWrBoiuEirHJubGCTM
27Jfvfuf7JzasSjmqLr6oMtKTtya6gWi7yHaSLkH++Wpzd+GRiHf9Grff/pr5jxsAZ5jb8zpbrjm
f7PwjC+d/4y/Fq/Hd35jqU+btpiVZJmCcVtvIiWVMDSzIALiuUK05dODKa9LoR70BEifDf+MH516
BXG1NVoIpA1KKu5KSQC3R9bMfZfr4jFXDVQFpxDBCO2pdDnORfxs+fu8wvC52OMYUjMQc3Py64/k
Qa0fVawwbqLxK1Zyhk8XHkukUTAjNOhXFoS9KjsABzBsdqdpIn8XrhefLLvDNd9763fXXoYfBhqV
LKhTbgx3iWUVTsNQtJScg+8n4vEMkSSklMdcBbrG62P7u9eN4dFFQCkX9AWVzKRjaYIl51mJ+ooF
eDr4SObQ47EI1eJ2KZAoGN4RxHBFSEIQXV34tNel0QJJVMD8vW6gh3kWLKXmp1NmifUOuev0D0PX
yxYDsjQjuAppmKDKv779nPCHUVVPhQxoXXJkejivcpiSxWBSV8hFrpPnJMMjWcabR1LqC69Ka/xm
QBRchQWSW3aytVheq29GbRMmUlr+dLssFGi+j36Xgn2gUgvpTIZvAeBfkike2nkAeIIh1HQrITLw
XKDD1p9uH9VQvbMLDOOdGZScVkTCZDUpPRnarQ4ujC6HSo1KG/m1f8yTGdvzonifh7GuLCWdGiQz
DOo5JfiR5aOpWVsa0ql5Q8/O7J9epkrCTEf3WROa4ghq5QZgZh6F3PiVjiVQnLFXfy3mcKODWyn1
GwDu0oO2ZoQo82Ik14v0P8BbfzzUIcUWmodMPLERzBVO5WlURxVMFkEmyCS7T1z/8UkteKe57Hjf
jdbDXh12OsCGvwLTe1Bv+oKJVue7wA19Mql1yZFbtRCYlUQeH+j2vnL1vi07vmg9m7GpA6erBADF
YCo9pgxG8iFkkxDirYnlygOXx2sHSlfvMRq4cohBT0/DkHN6OVSJJ1p0Jbf9YeDKMg2TXUnKOQDO
XCKpzvhFjBBhF1pFHkpwVh5eW0vqX3tpnxEQR3akWKalNZYE8rVtwL5AOD4zoN4wkakjigx76ccf
GLg/madx65bZHi8jqek+2Gt2skcVoGlO3YalrfcXCLSzyZ4etpm1Xa+nxtTISvHy0L9zugjs4pmG
TkPNFEbrnyBLdwv6zUModIcDOo+brSdXR5lS+XYG+ovZil/qzkj8IyTwK+WVNi/+to6NA/CGe38X
9S/+Y1PDgYzGFtOflJSac1yBpX1pV0ZTWNaxhrQZjh1KHvQyYA/lfKY/otjooPt6u69CAZmDs2uX
Lw1CCuFDT/dmRySqi+hco4DPe0VNyPxn+SB3WqDu+TeNm8U0dCkOWrfgIB1zd4QcEFQzlcaYFHhQ
omcGGiESElzG2hJ4CA7XuOsVnZVyI3/AZwD/xkb3Sp46tH3G0r8glMI76LCExdErwq65zTs7qa5T
FKw1QFockgGRJK44HB5FtzWBIPPa8qpvAU/lzcGgvkfAsZKnYa+lo/pJdHVFAVGTfQTOSfKu9X8R
i0Wko65t2fhAmDtsGXX15tcQFzDtr7lLsuQ/Foem0IIWNDGBZ23+bAcslIikCtRopQy3clZZ7vPQ
USloqxB3Ys6WucfiB2w5cfma/z5CWbsEo4e56WUZtyuBPvFOE0vWTAImKKPc3pAScrNBVCgm3FFH
+b8QCWcEmQXYGaUp2nLVu87Is532OozfnauxQm6gX6yEI2mU4qOFEJ3b1rK2nt0+RnASwkpYGGr6
FmIDx0q1wIkyqj89Y7K8bkMn4vtzT885+y9gMDiKRx1Aqvo9prFpsRPvaHd5C9xGjIu8QhmJ4ItA
OuNshEgPAhhZVbEej9NSdUv/2OLLKRinlmYGIfkJfgfnX8UPenh2x0RgBLvungDM1bQxU4QaROfm
ymHv97mrOmbD3EF1EiPdDh79I+5+ucs0j5hft5jvmquWFenm8qxA5Eylzx7wRzqC3cjr2Qko4g0B
sDnc9gk++aUnHOFoDQCfv6XanfMrWJP2AV3P4fas/xbjZm8sHvF6Qp6bI+mxKb61CaMxh8KQUFgE
LGXimGvmjR0FC6/QDH7fPjJCzwVuaqfbq+yWv2h+uWoxL+WnfOF6ZxsNQk9IhxBkWoxy2UbWoynW
R5pp8bUHH5cL8MU/PU4h1BNXn90j2d6747d7ud9lVb7ZtHZOEai0yJ9LEuvMg4Hx1t+JypDY9Etj
vAHgsyWUNCs5jbCKl/DqxsbTeH5iLY7PZ4g0jIAdW+LmHCHgh3iBxnCOe8TLou/0pL5nBVy3Xg3k
EFPKPqIfCY3e1pyyupFN2nueQP3wfYprGnM/bwD0gi4CY9AJ2iNgML4OOaq6gkcJis5f3aif4h6G
RGVvbohbPpN+sNFJ6l3JGYHeVcQHrBeP4hCcFqm5nkSzHKhIjGCeMZej76rKyqaUqTSd1+JmOO5p
TQ3uP+mjiNBTX5J6UbGxU9c8R13oJyFWi7ydcJ1kui+3UVL83cqu8Z3dU2Zxz0dc8SudPn7LRqbZ
UAxOyqV4XPj6w6zY2VDix2dBu7+/9n6NmGVmu9ZimjWelYDrAP4TqhHis5QCkj2mIrZm7Ey9U87T
lKhpvsWBFtyMvmZ/V/8dsW90P+9auvQ+7vcYoEurLKDK7ilzynW3cd6yyn4lxhfptf/4kHsnVnTf
YoSqzzAxVcOtFfJFKBy2M0losSmbeA4gDGAWV1JQ2lFqRQpHRm8ULWArE1IpL7BUfsMlp8FrHVoE
T/mpBD51p5jrwJ00NZfN0Qu41NVf7gd23WOF9v2YhLu0zUp9yM1MpNQH4L6TpIPA07rrnQZHFTSs
5TRFe3GN427Nb5ZIExFHyanpLa8gApKloRezKs+HemSluJgZB7SoFvhDiohHd3JUHG2+ZBcA4vpK
3TrXWMLgSN/K7f57IMXcqjiOTzIrGDzpGGShmXx3eHqN47fwuIZnhNdTfenCiB6eTlClcoQAClEp
eJ3oH4KC9Ds9bx8tUP3EuD8jT7V4TNGh3b6gU/CNUTgNNhIV/GSHGq+7Bq29gGJd7yc6tVxcOgVH
p/Bn1cz4p+/YN2UHwO1dQlE9fhHau6D11s0iQviwCgnroWMRTt+97skN4DsGFEYhsQq+lbCMmFuX
M4CdeAejbN5RWN0nCW2Ane/QTMB9xkClQXq+oii8XNWrivTzns14gPxUzHo+awoQEMjo3uopDItG
a4P3pjN4OKOWBty9q8mnB5VkgRg4fas/1/PqJACU9fWgZakL7QHnbo6VUbqd7BXdgGmGQeB/BkIU
VXc/2r85GRl2vm1dRxf4vQGdQoQLs5DK4PolYLmcvnsUB4xaGPWuR2gOt2aZF1zY64/kJowMoNpw
sGfRFHKuG0vADlF2zzyno1kvDdCcBUYxKkIgQFKdDbayApTD3s+3Ni0c+RpT4BUUhNFsevqcwFNJ
XrUiYAj514Eb/TjGMWZltLm2eqI429KOyy/frqj2sUMvm3qAfIRvPJyQltOV4BDr978WSA+RInZA
Kqh8WkIaEF4+UYZ0DI8+xn1qZnat41Nkae9jubZrxvv9jEPuqPPz/G81s9FRkhAZ7eWi+g5CxPuh
ikoChdIACGk+zdZDuKlJKyuIf3D1LQuquVAeSExxf8KU/+9gwajLf4flSkXVefGr2/sJ2vFueWP8
yt1dPqBdqzghoFMrCalyrXWLKHuMkLJQxHDRI90SYNqYG5hglO/T6ryhuVm8bWflqedLBKsNnNkV
4zZYmXKmvWqp89okguhCr7F+PQ0AYnAh/Z3gaLMF92SmXANb629RAd7/NKA0gGa09VwfffkJ+5om
rKu2V6OlVCFDySrU0hENgtea7bWYgeMbmYLwu3fXBvZEEKC8BaZ/LYTsKvmZYKNs6F9amybRefqk
5OrVC45DqMMIF3364/w2OuSZV0Xaco62iOIiQH69VFXLLyTUDMOzNMw3kVHw2J1oADEqgxEvrd6Z
dX9IBj/gUZs+krr2KdhlE5xX+mCqxGM1/LKfz7M4TkFWcOFrsK/oPDHtnakhw8VksWv3soZwB6HU
GeDs4bztQWAFJeZ9IvfEbZjvHhjtVPwoQYigapQ3FhDwejZc7J854+UIK5+2WlTjYKrFV/ZU62rq
jv9j8fTAZ1Yhc4C9oFuzhKj4Uk4nt9XOh6jARk8SQuif7/mrnxMklxNQLmat5zuQouLu5ml0RaWp
0EHYxPj/zbfF0Vg07ZF99CNuIIltND+VBidGNbnVrBbaBRzNAk3KIBzu9m84BeA72HZnUjyXxR9Z
MZhrBoU2E/g8RUYmChp/V36D8wXuWKd1UYZ1gfLgIOa/Qw6P3xj/ygU9943/c2drgCp0+MHSJyoH
SK/hzOGwtkE5ZZAI4QRO7tXU7Rwx/ugi7lVBGF/oDenwLJzv1G4aqCJfjR8F0NgcQ1NaZTkxefGJ
FYpSdCydxrRT9mDm1gMUTh5mhk6u1EWJJCkIQpoQwcmeduZ24gLHHURStXHgAcXDERXUBl9KtNbN
4PfNHZ3S+u4ZpLxCfpKiemnCBRBilrDKxYsIgh9tuUf4L83SCfyAOl1XT1nC9wpx/RgJxXrGi1O7
HPyu5XxPVVl9gGpCBLLFcoxSMaDvtWKYzubfcWzSi29oAK0iFc7JIwnxy8t9CQ34Yr57j2RraPG5
CR41K2UY7b+GaM+7QecCQsQUmISad67cPKwUWGPvKuQDtDgsDQDLIEPghRAqoHORWMMyvC+NXtYm
uXdHTV/IHfRMQlLu0d3Lu40ECJsJajHE4ztHuypt9wt38zU4ASexkSXpLmtYplpSr4c8azVEwi2z
Wo0atakbEn4a9klNOXFLIV+qXc9CvpNeAXBsRsAVp5cf/TA4nQmFLfVdfhn16QlkAqPEO1iRJV8l
v2hFusUINmO95ZxXv6DrD1jHMJZXMlh0tHgXGrx5wL8aSJmrLu08Sv6fk9ZFxQsKgdZ0oCdrT4AO
HUGz8+rJrfpVSpUnFOpf6I/pf5YklgacXKyShJxreSKAyDG9oR/PkaJAQjflDmmDMl+sRg9YkV5F
tsPw5wUVWhD4mqxactmKpi6S6AZ5cror6uWU9SBdHpuwXbV8adKGQPwX8fjkF1wbNHOwWAkxRqnX
McQChwzkG/vPLKAOaWkjpZlbKEfjl5IFqjyvpWcHkqBlumCbqE04bbiTaWUv/XJg3Kr+oy9eeWJc
iPV/w9YdkhlFVtpEZ0moVOOeL5oaM6FUIvHqYo80o0Vb85KTYTNJzrJRr0voGbr9y7HIjmiWCM/G
PN5DUs5OKsjst9LOk84aADMyk76j9H9RrYERkiKmIf+dvaR3QpKkgaaE++St+JSgYPTtmxFMXLHU
hIkgEjS5N2k0agCZeFuMt1GQiT6cNlZUowzhEC+A8VK1ENJx7+h2NwEibPO5RRiqBqR+jpQ9FyS8
CX1bgbDpAEveT9wG5RQG2jh+J9KVzknuYzFgHbfPkDLtH/t1pw9tFAf77zA2i66/5bNvNGNJxZNf
nfLukT68Ps8lJjtIBrhOPSvqtSm53iVKXQr/9ckzEeOuz/tou0QLraNDmCrWq9g+P4A8S4+vUJ8n
4snzMlNOy9LhanG3WomHxr5z2AYnEVYAPbr+sLXJ3fzUNHCYRBBqQoioZjljrBqP51uxfb4VDqLH
KUa4NhUTZ9FwQDLE6RWB2Wrk7bvaW2XWueUKEMC19jiSdiuimWF0IJAI/5d5ChgChxaS4AsV4njz
/TUFDkdzokdawr9W18eG7cxn7QNBP8+uWGY3whUaaNxKHU9X8YIPFa+wEiuUx99NfSWGLAAF16MJ
O9r1ay5rxikeYRy4e+XxzeYYnMbtFmLyWNR4dJ4ZzsYeaRLaRBVzGa39n4I52g9+0UMDZ7I66B0z
ByOCAy3wg8o1wMaGBZtLpoQSu896VYPHZmeDdxV8pnG9tJtoiqDVPwG7smKgMdA6+fMqnWp6u418
hkNu75toO07bmaddQXqUhFUUysNLraXnofa448KNjJ0Du319SOqIxUku0xVKqLfrcj0RiNS3DhIh
gWmTm38Cai4oCuNOruakRNd9rMYyFfNiEn5MDRfkG0p0AJ/SiMzI+8UPzwGHb3ox1Qvx7OrmdaNe
7izHXICywFU9Vxo6wPSV7m9QOxjCbu+rkgkAc5II0vTledcM0LpQ7it5h4vFFtmfxWRUsfksP14U
3d1Fp5gVFR9X6KHHjPDERocB7HYJxyMXlXZ/sXYHtEkOV2N+rmIsFJoxWYiwiLwCqkX9lmclnIAQ
HZw2rxk4Dt5QTWr4tGX8/BNNimpyZixbDbp1X+jYMBKibH2fG5chuN2VGISvaUK4wXsvZ1snY/O4
jCYZXNVJr9100gG/L1vyfm26VAKxwlgvTs//aENi5ijndhChVPSWzE5lwfNcZghZsoQFeQXD+d9p
Yw5yMnQjYei3FlNtJkkRocFUtN0wFPS9tI3F9kct9pIuZgQ7QxiG1UKQgH0e/sOWtddIk2G0pi36
thS90NJ9SjDbP4LBy8u2+pJZZDh83GljJEwnuGBne1MjR0Hs8HRs0Vf+aGkF7Mt9mljU6WkC0bL8
BgW0u4AwQ3di45c+4S52paVLD+YIDYQWI6LKUJYNTMXmtn8ADw1N5ZLYRJwdJKw2vAwPSbk9JkO3
FaS7Oeq79gHYe0o/nBhEzjlu8erOiKVgAzcKaFqsoy1FK50K8QZcOrHRBdkoNNXBRNlt/u7v2rdt
QqKGEzsNoQw6rVKuaRWFKs+OeFTaSLnwYWWFJ4CSvBJyv4zmg8m2bmR2Rmce1nURaY/5IHcqJpJA
QrfaRG2USjhbdNpLetOSgulKprabPLANz2iadNqrhmTIpOSLlSltHMsxe1iy3NbeV1Q3bzs+e8Pv
mRH1e532AYIpDqKqwy94NLi7MYPAEArCBK8htAZNmHBZO/lJxal8BFzxwyqBLIVi0lr6Rn/fruAc
mE2upOrRje3KqeUC6OdIMVGc/WqTFVB9Gkc/HnReiRLRh7C/ThJ6H0NHWjAi61JOFWRH1G5FBWMR
tBoZjk5Nem4X4V1WEqrBlKJzUgdxhf2/1a170kTZImWaEkAOfDLsxSvQs+0gnFtauEvh4KBtDFlc
ZVldoESU15e+BMcO5jZGRV2e7rvyG1JKSEkHmy5LbCqYCVt8V73D4UGPqJXCRD5/5U+qlzoADHeJ
k+CTwvIUhHC4Svuznte2HcXeglozyrTgocO131rPudsEBldmoUMutt2qkZvXXPiqvd3WGPTcEDRk
eJBqbdZkeoIM/1GBRerBOl5tfGGGcIlHPfJMtkoLDBxKtvWA9kyeEEZ6aao+9ODS53srF0bk9Wwk
sA82xF5qEyYNn9Tu0jKIlwqIfoeMsP1M5/4/8rdCMpuwZiqHEdpoPWpyDYxw38AOL7hGGSasTLyF
W9zbfMje/wwl7uN6e+bG/twrqwXekMtzQDAfwCYl1HFez0A6HIx5OkUz96sLQaeOpPdWs8rpONEE
dP1aIysLOucJcsll/SjCMYqrafFjEwmsezqytg4jfyzd7UgMGE90ke9H/xDRR8f2kY7Kev/lYCLG
WlJSnR9D7cxdcPMJpksuXcVpxhj3bmw8RLsk9jooP5nCPRBBLVZ1SZ9hhkWA8nJCV3E3Tbrm5+fQ
mHqxbJwCaL9KgziOVAjIdTvudIxK5TrngD5J8++hQKTbrzO1cmIq++wjPP6VRSLMWY1m1YSgwwDq
nTytaJ9giEMbjUrDCEmur4FCT3OWRXd1D7neoFL4CBRP96kVoeikB/SaHBHmL2uNUAmMCjq/65fN
XkdZDHBLsDPDqNXcs/T47s5M4Eb7eIDXfI6msy5vjPJutGPC8xon1IuZ/45011EqdZ075C8tpsgT
GntPOtZwRwrYpTk5h2goId1RSktKVymr3Eym1qL0WeaZdIP9TWKSV4RwvTR7G/y8IispUntryzqd
ELWW/feuDeodFf79qYngZkswHdNZZ84lrJ831Iu262JaVIN/NRU6TxkCSd6GFnD8Fr1NABUGTQYT
s5sYjF4/25lk7+WHLMGBzjRvsNIe3W4nEwQWMlj8aso3ekZxKPpkGRhsYgylydzR142KCOQSWAve
SeHhpail46bCA23mzHWsIodmMVQFcS3KCQuaDAzaSnNxNFlcMghHtkLdl2gCEknjB2UlcrMmBzdj
6HCc5YPsn5bxWeUh4Mz43Vovj3BHy7vet3sf7GlruYeavQSQ/j3M9HnK5/TFw5BMQUM+TJ3JYing
AlMmJg2pPpmy0hXTowJPqYy88zmBI53aIaLpkYS8UdjQqbunl0RY3cZPVf79u+nDb+HBcHZNFT80
mIvlxLBhmHM8svmmBjUcSo8qqqQZX7zaHUOO7cmRQ7KKp+OegI+tI55CSTC06lpbsvI6126yOrAL
+mxynCoG+T7DdOk3iawGLm4N5xaFOCaNUELLJe3OL153mDzL8brzur662qMocVgy1/PBvXlqv8Nt
kWOkiLUbMAPaB1uO/rKTXKRzpPsU7YTXeOzafQZ2gAwfDmv5OPOn/PXwMTJb8FNe7AWviklQ4iI4
DL7Ud/OZRuY6BzZ+COfNVhwiO49CpbwvFWNnrtt2VI47sPFy+rRlNeXUKgHzKB+ktevA5CJHp4p4
XCxxRb9ET6mZn2e9W8NQjhRaOzsOOWBV4EJAYhvHUuZXwVN5+HWHiVC6v4+442VmDHjIoe+GHB1m
nd67fmJeVH8SSsTDvO9yqTYEbbINDaogfeqlXNgAikj/ThxSCB1WisuVFrWQ+6/tFuphoNX8UQOJ
c0AHBEa1Uz+uFCJTLGYnS+n2M1EqZ29DRQgvOXLbxkGzBHXDXBFPFlSBLtxsmGBDGXo1t7PrO2L0
okWAoYsB+fQiNNBmBuzZDs79A3vDzjsaTRjji5YnroYqvJiM+BG8Zf9QlqSnVi1TNCQOE8ofRhSd
iciAjYCYMkVhqUCbIhjRonoxZzmctlP08xaLc89yTtpfgqtm8BvyJx38Op1ciPddn8I8k0xHY2Aa
y2njXAxpAwtADeuKZyoWrfaWqwImiMb7ylTD2i0+LT5p7o4BIPE9u8ARrkDZrTAivs/bcVFW1qyJ
PrZMin+bpBkTMDI8rPdDxP+bnW3SZzsuwlXAZCDo7g8XIxKQ/qPhg6uucyXha/ObuAWgZNkr3uei
qaU+2OaLCHcLQtPCGJGZHFwjae5sgHVpcANhnX3PICVFq500L65GngKpMHVPkHYnQQMvCdzk/fL8
h9sWSJQcDBIa25M4IFRkMLR6JcGRE750X0m2bz83Ot5pVxEHdGzq7x4IUriP4l0FhB5jYEuTgtv2
Z9QS2t4vwXJjQqvyvgXpeBCOZtQOcDx292U4ok5fO4ZGKZXPG3q1QcotFre5x0a2y7XLlMMZUahF
pCH62lFnOdzYmv9e7/UBLspSqTPuMCBo903YA0jpxGKgAnYV6m0i18XlNDYvzhoORmQYPul6iDGl
4iECgMgdZZRP5MzPGiw5Ti6ufESWHzz5L6ZeHENGFRuXHt7k+v+Jrwq8kI6q1R13QeXp75AOTPPN
A3JsfKiQyJ/IlFRAFC5jbT1tWsLj13Gm53Whpi3GIAXnduuj0vq69VJ9YtOS+y64MzqunzJ36Tge
qzrBS1+AsI6w2vK/CpPdaVJb355Hi+yx0gUNjDoqMNOwFgoHydp2l/+ZPj1bgSY9PPA2LCj+o15f
MM4BFsosPQ77wSGafZXj1sO82zDSB92kUzm1cPhkvU/azbWez+OFOlXlTEnRntYml7INZuH6fMG9
L9/HP60mSzwMd3ziKohOCVLNIaozCeSAmtWxh3Uemkr8MSgOXAvF2zPb8E9B8R41Cbo1m3ci6IK1
I4H6kczmhDIK9gveGf3jl+aWJa7TpvWcruj8xR83UUPXs+oCHgcUkYfan/OuMBO30kSYX9S98nuE
TboAPelhokJbhsyY9dmBmsV24w0Aok1xQsZkKozRv459hnCKUHu5qhyy+0h0lwr5PJ68MZt/dFHs
PCc0deoF6cEGmowUvr2cWtlTj1g/GLK3B8zP4GI3xJw6DuagzuRY7WOcMYu0XSn8bkA+oFj+30kg
oC6nwr1MckLFtsKvfAGd3+7nHZhQf5cQRpZu8XkqTifww/7+as6K01QusobJtVGNncbTbyMhGnoI
Lz7IqlCF6OHatp9yJPVhD3bM3hj9PhQUDtg70pzqvKPKAqJfha3CWpXAveAQK4qyJV8+Q91JrbDL
TWUmVFelpQ6McJCxQPnpyXSpqiZlofft/UxbC0uJTxzobIfsiihjSAlq+14F12xlez9MUhhyUuES
8pzWYx1djN1J/Tw8ruwBINwUfvy3vLnQpAJ2EruIu44LIzEGt29HhjK8a1cAoxgGhC7jlL+uixIN
RoNbJnaV9gaHXCkutov/fl79sSemQu0zE8wFWyxfQJvdhXpItIXyTo0+31WYmlFY2j1Mx79KS2yp
EI+BkAy2AB1mu5LjussmQx24un7ylovvR6FLYU78+YKtEzXLSkrYH5adKrRCRQVmDdyTcx2YCxux
yCb+v7ow7QxzLpJxv5VFIhXibeF/ZJxjHyPiwjYEVjYO/9sfgkwGhdMniAJGpfAlrsbpQ32M+8zN
0UShpKgLfkVsnyCnsCfD+ct+Q2HTFMZZonn9q98tNnHFwWfWMmvV0FANVDa1nDvz4SWgZbqL07vW
slOikrlJNju3uSDiAtbQHABX0kLRGBnKZXz9vWVZ3VCa68llU56eaaK1CeN9Zq3P8DY211Jr6h02
qZEufeUNiTwwlpBvHjpgLPn77JbTwyVLgVBBXiJz2V3d3A4qoCBCldA0DfDVXlShmx0vD4jz9q7q
7bA+LMuWztC8ZW9QTe3tDVhMFJ9U48PUTa1qKKEya+1/E+6MjWK+rt0EYzBMSBSfJi/m2rPQhhsV
CEf0f9YpfAoim9LUmLeoj/8UKuKUnzcDkfPKH6dRgTdyJe0lt1FiQRZ6vXd0pKpk1QEfD8UYWQBi
dN32yho7HYuoDIFdZOMT5U2O5UzOYA8I/CUeaI8ZNXoKToroOBtJP2MFCd0XLjzdYRkfuQk+a/pN
LocUElnPFCJQNJPS3+U3z8ktO/hZ8LPLl9CicM+HKJNV2ITkSMb2OJ199g0v3s+IGTof5zBg0tfC
NQJanrGYLpmnMworxjf03uc7GQSgs/vt0Q2sfPze1Dd4ciEaWiyfPnqgNOX9/1rpvxKUeXLtY8AW
yNu+ATRWPaUYgK2laW5gpu2dY1FPprCVQE+UPSDcnxL/1IaGT6p1vmlB0mgHjtTGdvGAP7F8vxfd
8aNO27pUs5HATbcpuzN6BthzY2hU4T7vWheyByvB4UK7Wn6PbXD1D3/+75z+4OsLv5V51+g+scqB
lXl/Kk0Yqo/lo8pn9l00CASDEZ+tgohwj7aIkkNoOkTeVOAsQCHdq7nzkC6YbB6964AzItsbpJr+
exul1Gcn5l4XSwqKIfVtgyvkmzqJx3KXLxjffQ8gAhOsO8cogS3v9P8mJkXK5fUrXdF+anmQqlyh
/hf1PXPGwOrKhAps7xFm5shipAwLTnF2tbqTO5IQD2+QdhTwRcfvhx2wUlxULvlCn9Z5iQZWdlq7
w0Hwsgk2tSmbgyAl5dvLjen8YXItw8E785VjcOQp3FkhM9MZ5Dlv/hvwJzqKbDcfdJGAvpyACBm0
VMyiXlBPkJXkpiV7OP69WLxieLNU6OJMj3hOzJf+qpbaSqJC/9YjBXA0H36+LO361lR6MUN3TiA/
vBirRBMudmVzVLnJ1GAvy2oreusE0fVOaDLZ3l6Y0Z96cRuhPX8c3DPu1rBXYau5947sED/Tz8do
jde/YJs/J3MvBT4At9LbbYpK0NzpS8a7eop5WgdMMjkvbiAauqNn6vgJu46ISXIDcUkZOODopPwF
HQyPk7nzdudiHtEVoNGZZyupSt2DrI0gRYuNQpRvKgHKULm1kqRstwzS4IL605l4vaAT9BvOTqOy
plajvdfhJ1DxFvKE5AeZI27pNDuWDCm8JXHzm7VjuHoLdDwJxX+ez6kmmIqtlnzAok4b/jApIF1c
2U4pdyjJ7vsTh+EkGTxXrRoLj+xCa+OcH+I3CfumT74WiprNW4dDFI32Py4RaARh7M2bEIdz6Nii
xn9Jy96m8vW0xI+Oob4xop1H13luHoAkciOuJUuRk5TehrzU1r04yRcRnjy/3bXvaHRnZcqAcGOy
2t5EpmnaGE6bCvC2XdYNXNAfH0sWHr+ggGciCi411qkXaJ04iV/6YdtRaMNw/5q/4535rQJ9CMOu
j+lTx8WxmZFWApE8jpGjsY0RpQqXM6n+M184fteiTQrCREPkZ7yR8EGa90Pp/bNlyWVz4hFpDEPw
3pboaJlQT+jVVonqJmaJ4jN6oiv4hNy/eri38y3wooeh5synwwNcrIzj30R5Y1oK88ByeRsynZv7
YNLbAcWdCGnEuU7SUplIEYsWq1QbHatyCfh+4t8NauZ6KRqSLjKakrUpDut/ybTkQ/vtRhF9DxIz
txYT5VL81d74n9JwWEONMy+r9ck+gY1v77Dqd8OkQa1NWt52xijOD7vMfpbGSUcaFh1Hexse9IQp
l9Fb9vKeGb3SWDf1Id1NoNuEa26k9+k25gqqZjH5EIHAK3sjfPi6L4cz0FEo08ryve6jxrLXX7xN
vOkF6MpUsUAnbXXrK8eSZvkTOxc8k2Zt4BAAo77AtBTd00NzmRGkaMGA3zjzKX4KG8jXII8JYkq2
k/n8Kh1zhD87qOjKWZ+uJk97pKxZlxPA3G8TJgoAqGuJuwTpyQoLo7hj0ie42yUB1xLmaC+PLn21
SX47FiSCVv3tp63btOSEQmDPe/Fe0vWNd4nF3WwC1kdtPhHNXmK9hMOfyEmsVMABGLRypGE9agqz
iNDifIwbd2oc3L3KQGWn9Vnj3wbjRvJYZ8XiizKFDmswmJSvhpb6E+kwadirv35Bm/fbfBOqeh37
KLms5jZbbWEmoVmETq+/Ho2ttWmddvfwa+q9boiCt8FCZKr4jPf98dF+HZZFmzUBX6Zh6CQ9j6ez
SlDKU5y/b4bLRB5QFUl3+xsW//DPgwtzW56MieqSJOHBZ+RL/Z2471zTcT6AyntC8qFKLjOkXBQ5
TYq3qLiBuvHdUtQ88YdfQ87gH+3XHvJe8+GyYwC5iGmvZ96XrS6QBiF0P8Tjk6Ik/XgKw5yLOFiu
rxDDrnmAZY/iC/UeYHkUJU5lPYCf25yqKS9XN5zwXLpFVWa0AGDx3EKSQiw78DxvZPOuAr01FPSF
XWsGR61NaqdLwJxbYZ5+ms6Jzoe09VVDvcKBnJTFQDNA1Lp2R4SUHn24ZESjJI5pZQzuo8fRYkzV
XOzZSfPlrytOOafytVUok3mU/JnGiZ667Edm2dDCRkf+M6AqlxgJJWwT9Jqg2rr0t5Md5jTYEYbv
dmsHRDvG/zx2owB7AVK68KbCTDmW/PT8v+8J/HsmKUImNLZtpFXunliFmma38Wbefaur+j4e8ema
8lseRXQJD2/HFgrghAbB/QajqI+v3PZ4JQCQSQB2PK7sTnL89frHgm7BLSgbFOPEKAYGirzYjEFS
Di6uUwE/6WeqM0qhZaLc+DZVKTbLMRm+xcEiv3krGyPpzA+X2b1qRUjc/lTKQ+X+FqIaMj4jafFd
N52p/m3Rkm0oLh0wGvsfgJChPPPv/v7QIMZhOLRdOyhrOexTj4/r4EqDiQ/aYhmteSaaDbyv6nhJ
bUiR1Rn60g6xJjkQPdaHfDhhXX353kapishewC0fTYZOVC0ob7pjVrn8h4UFza80IAtwmwmKUAVC
0KgSEuMC/l0qzfl8inMhH0xN/s3sM7qrnpTdHUZgce+LHc7OQA2l4pSJq/1v3cfL1XkTX0ISgans
iAKLur4LyilFlnz9Hf7u8N2X3TDZw4TbR/hLvkpAaNNh9I5zOwFopRqNyXFR7Kr574Xe2+7R8LuQ
UTaPy8Q9M0k1PJd1OE4jG9b+/ouX4+Hbfg2GL7oXbtVSoV0mbGiqmwQDer7qDRyc4gpPQRuLxNn+
0SFKGHeAUYS8D8cTIk3CSYgdIHz9mYVgfv90o2wWwo4+YWht5gZk8utFxFFRTGWV4xyvgjhfxWqw
6orOFQMYUlit4XgkMpPyZXFeQFff+UYNTZp9iCdFotB3BvhzJiXO9s6r8pkWieFXKCd7i+ntYJDu
8P6cENtU+9rXrAGY8hrHfb9x6ltONF1TnSR2kX9g401wUcqCOXZSy1MctbGX/o73uMCkPMepX7AJ
PNYo4LDFLWr7geLH/P9YS7JLvScxA3yrBFMRFQzbo92VCk5tnn8XPq2qr221KAkXrYbXQKFOeJn+
99V9lHkY7YznvenKHciC8ZvT8azs4evVIhI6m5Jm2XFR/8Onj+YcxMRzd2xerlbW9J7TT2S2405e
B/LSkUu9j68puhBrbKxxpzUTFYEpr856xyxE6z3TZXMcLv0v+H0u1k0Mx4p5KgxYxRp7z4FdLN9W
cI+tyByWCAkT+VZd9kQU6ReLk7jJXM0gQV4vZVO8EAk2j7FhLaZYoBHjUqJ8mmwhcO3HtbH1I1/h
IJry0LXEqMvAXOC2gsM6Um77ci/r8TVb1TRQlSirxPag88VYXAF+736jD3/i78Eoe/JwLOHWR7tt
Ug2ymWF2l87kx2i9KE5y/xzEijVmFHpranZ49o0HK6pX9WClWAnaBJIbOfy9dKGLcAlpeYdMye+W
dVbrF6egnRGhX7DIqoz1OaJCDSiqbxXagbIRJZgv9G6wxpxC5HjDXx6V4DQi8n+uj/hrymTbbL0o
8cLsW/89UIw+DJm9YqNmGDPCWLnvr8TMnkEcnTPso0WyTRvmOe6RzKv/EvDUk1vD+T9TecLZq/LN
8L6NdysnYkRMz6BIaEIoEeM93gPpH5TTrFja1ER4AkrhY2XdIiZU89Duaw4BUQ8S8535jguwui4m
H2inNWyZQfV+ofDqKVgSt7B41JQdXu6dhW5DLEec7AE6ONdNjaLTKfNaDYrUcBFfTSiG6ZdeASBm
/C6yGQIWDqkWu6Y6OJJc+tnTScqcFcksfttsFS9S/PVuu/fueFDwbGNnxM2FOB9X1Ur/Le77Ru31
S7YUtsc0dRJe/3+7ZGHtwUO2ezRkk3TJb5hKwe4z93I1uS2DdtmKz7rZZUoROoymiMJni9rxEHnc
0hsEHsFyOUu5p9R8q0UQDY79s5d4+ryPVuhoa/6xd1Pq66kAhXoSf3p6mGE7rQ1t2eKy/nnObOzx
ttXxQ/wBpF2KPGV7+MZs3Q9N+0qN5qFP6grjPhaYhzZnkxI8aFSw2G2RIaRh7uDbNSSpA2fV+J4H
NOD+4RQgqA1kSajz5kDaBydpFEUf0pDQ1iPuljnX0ZVH6P9q5ac1+Kn5G39sNKr5qGrzQllVbyJb
DS5VYz73HzIrKFC6Mj7/JcJh8oaBw5GCZgvRfa2t79a5tPWvDY+7OYC86emL6e64KlppPZKai9wv
xhu4RnRQXLsECtNZVPPI3xFL0+ejjCdJ0JN0QIUb93j+QQj6ugLWzMKm3TcEFh64oxoUlVJxwpSb
i5wXWPxzAShchMhHKmwDa6y2g/pySb3o/gpXPV9vaIluxJrFvJdwSETxxjk9mgQbpMoKRTzUB+/Y
KOSVdJ+jcecy1KjmIxYuNku7fLGug73CCJCu9i+kSQ+LDh4KXt+vbTR5aoWHExY0x0RjGzT52Ccj
xa66sMzUAJSCBQZ5eFz9Dehz92xxnusZ6erN8At3Q+buo5qSiEwirg5HN+lr8zC/2kaMBrYPVNCV
jobnYmEHpLwPucODZeEE2IN+MWLruFcMlz1L8ErDOovpnNJu0wq6bcq013GdMNTuPvuwPEfHXPvt
qjQ0/+RTQUCXEoMAzdMqmY2INN5V6QuK5F7fmF9cohM+Lzbzk2WWbee9YM9ToMJKpT6MI4YmLkQi
56ZXx2jMeeGqjp0rqio/Lg5VloyvWua3AxmyHl42o9mDLc7gSGg3siXPRNYA7gSAYHiGzBfu0iJj
3+8xemCCwrOi9SPYdvpbfRcdlsDKoVOSQ3U+0MnDt+fuhvpkNZCDFbXuvlZhnFz7FnBTRwtRDN5Q
5A7f+Ib2rxxAQ+kR+oMK/4JjaUaGpRwN3u6WlfnRTsl/tmLzBG7sMsCRyumbXGL1y6rMEOHVETX+
AZVHmcrWCrxTYEzZ88HwvI0E8hZijOnosEE5IYfNd9ksY5qgUGlmWo2UfkXNmmFl8i36n+MZy26a
WaWJcVLo/FJz1/CUCvVlfzBxMbHbn7NA8b4dd+F+j1umqDFKGEWG7k79NmOK6FehTJHFR30land8
J8+8n6XrAxyEL39qBzdGyVoRit6asTjiVZkYJP331VGS72/pqhHe/sAuVk2JDLBvpEYU2yKfFT04
kMUAkCkHQVlgNTl1h2oE5NM+CJuATd3KAOulkrw9JBdwY9SYe00jU5pl3vczcK4AewRwFpOd7sVg
Acuy+NILq8Aez7dLRgffZqlTd0BzlnbVo88iz7liQH0CJ5AbvsBCamL9NVQy3qSXgaYEK4aXqUtY
CkA9Dfm50lngCrUmOTNvvQ60XCIWV7B4z4NsWt6eamK+FHwuN3HjslALtg2xhomHC3r8RRWOygZ5
U5XJ1wq5zQ2LPXFbGWeYMFjSvT4mPjcCuxSyuFjajxqY1OmiWl3Ki5eF63pfFaXumRkhcAjstH0U
WcH3syjE0vXk+Y9n+qhpJG5wJ3avyPIgKGjIOX093TQsQA4kGR8sE1r9sgAhtUh63JyWgSuYf7ov
StVJZDvlHi1XI1HqQx/9gZf1W/gwAp/qx1OlwhpiAJcsc1tz/3zJH+JYPFmNzWaQxBOsqxiISRz6
uKTbza9Dp6UzPuxw8pPeWe3mePURx1TtMrp3PEmzGjQo7gfPJAFYROm/CScPBJEM4lMDIZ01zybF
CZD1FPw9j9sLJnJ+UmRJp7SxydYKoLBHj1wHBH3UazW9rxb0D5j4gQifPrwWNZyutCL1ut2l+l0G
IXaGx3PboV9CPWtAmPCUWuZ7rAxTfwe3pNHroJSZrVPgcilO0I7fXuHx+GP4OhgZl/irVO6HgIcj
bDA2IvKOSXvLvPqjWWBxjnEe/dD+bd/fHHLz5iUQYEPxJYiH2wizA+DXra5W8SHCdVn2LFmU5YvN
fYJVpwT96qmNv8Hy6gU1soRyQnV9i272+eMp24Z/lMiQ59xH+vCt0Uw8rDeKNWDvr6SRT6+6PxO1
xx4PdfrMC5UuRLITaaHJ+LFohkmq/7Yuwz8CiNrdqyUjtrVQAptat/dMNK2QRpJEiku1qvBObvsH
tyYuIVE+WxJW//YlCXV1z3A36HI5KUg8sGZzFGTU9Q6gmXKrqnAMybB80WB2YakU6TKdkI7VNWfM
sIYLJ1Y8PoMbroKYDTHMGY4PZWgCIDVmJxjx4I0SJufs5Zu11Au1y6stSasq3QbVC0KOMacNX1Xs
ONCqCf2TcSmtfs/lnuUAaAtE1csTNNHYWCt2hX5v5ZXe4svTOY1SkN+sCShVDHKZOu4veGehjSb1
eLj/Jo74XzwtGe4FzcMEEMZVGMThPz4LiPntG3/KmRbQdRrDdK9beXcPk8CnmwpDA07aQTDlYXEv
YyzYX7zAUr4Nlc3NADm67OzZGSLaxGvW2EXixVQgxJ8pfim+xwY+D+N+JuSKPXd3/oX/v+ZA9nFR
RRI5GawDFYAbDkzvKjSwf999Epoh9OcsM51GO5LHw//SU5IumAxbhRSUlq4UsUI3avc+jpS7xrAM
Gc+YUCLgD4jY2C0sziK/73uKyohIqH3p2CnJT54KAFtouj4DuAn/yNxRFXn8nBK4dUpfq+lAVKRZ
de6gWVOymxNLkAFUfDugygS7hGqJj1hej/wgmhS/CDfqeLQCVt4Klv+Qh5hY28PnTcbkebDrPYXg
06jlRbtYHPPpcg+tVF4BxI/jc8aqiH7XFmmyO9G0recw0IFdU1vKqqB5Sn8hvRguVwgCwkpxfWpt
HxZvJQvxNd3QlHrh0MdZW4W2fhJijsGJThfpE8hj++t5AnltUYzYdKqoaTje8lFKonpfMl0u2f8f
bYqB1vremZqf5kF9gTglhtnE2omlmYl3/9+vJ6zJOi7ClumViFa2LuFc7WPOjnzlEAo+cZqX1pa2
q02DCdS22ws7gG30pn9169zNo/vNfRIYPpmcphOuJ1ZQY6oX0pjFwS5nUQs06KooglBBAky45J8B
3jHbdMhEbytNUdEz+9X+7ybwCe8OTl6L/5H0sVmgH+KyoX1UJkA4ArOJF5TBCO/DYm/niL4JEXO+
Oaa5naploWbdI+8yhfWEmQr6uVg5yVdR0VhM0YlofEfHTlPlLsS+PIUSsdw7D9byioMV8P2FauNc
+u1Fy2Y9u1QmY4LkUV1sHVfnTj5Ya+s9xMsyqKalgEmaEE88rc3ArdLlciv47RcGLac/TzWVD46z
tQowkj55hSnIoaITgj+F6ci9ay0TEogpJxBcDNRISxWV+UO7Dye2oYjOTtDr3emgKoAcJjq20t6s
WXg7mNdj5NlcWVKCjyL+bb9xFiz++pghFz1Xiyu8cWFKYC7oXLK5vPl67mpiVTcSdjdM+JLporot
2bqJhCq/3PLa+psvm1XzMDskqazo5hYy+ygPZYqTrUbveZeTEyL1djE8EF4Cme4fTbh1bGY+GsDQ
nKKW0nG9wftnx5+KKqg24PVrB6FvZz/h6QI0s088seqmTrHoJFMg3ySWI65D2NGHC6yWaSArXgEi
10pHHmu5toi3zGyH5ZfcKBEQEc+EPBWhwCVhISRcB68e8DXtDA2gzdTSDHiBGkSy6VKIgms1pRVD
fZ8fSNohsUnKFugksnhHT8SSP1MJFTRDvmBjnuybcJT7Qlo8fyh+rENvxUEF/7YCorlgoMUZjBFB
t/5Jjc5//Wg+ZWt3Dsu13ohM7s039QcI6j4ml2+t5J7ml6v7TesPtPEjoVVoEIQKOppjmAdcIpuM
BH9eevCks01NDsc6ojJuSRXO0UEUwCAks05qZI//JUvkhhyS9EkmFjpbA/9928XFufM9Wt5Koflc
qo0zo/2m/lZHHcgy17xQ8L5ZLOiBz5MJLC3Y04v4dG+GDDhfp30O4ZAZK1H0UJvrNOKdFAGEea3i
hVLkIZRtyXdUGgBGNSBfCyLp4t+hwsl3MU/8CqBANUSHKLK8/4HBbGtpqiFDuJmiCVTqSLl34ebB
1GGIXqud69Wl1quKvaas15Kqf+3UUk4GxqOS1EGcWQo1OxK2+qUI2V7a6OjOWdZFS3i9aY6qpTxB
EryAsq6ZhIp4sbDxssIMVNP1PYYv9sFNLU8imvWNhxfuBtIiVEl6rQKfqBBtRb6/Y55/YF9f6p1b
NuL3NDRW5Kxx4dzYuVDSCoBCVVrhUN09D95HAZt5869FEZNH1zHGCAnY67bCTps7XX7+dHT14UqH
PkX269sW4SmZ1fGfd+OT4DCN9PCGGqcToucAg3oro40ppvrkjUCrSkZ1eSkURPp5s70Qx8bgDT3T
BtgU2awQqTZQfxgU5SI594Q8ZhxLFF1vEIXdPL+yAdBLpYVbny6+8Dbn1UqU2WC+MqouaXF4ynE5
gHWFXbe/HiFXS47Ih356IGTzbowkprpdexFtsaL7xxOLPIDsB9bd3/8IArHSSEKhqM+uk4Z0P/oB
AmnsPwfubWnqnngHrwWanEoZA3KWAkTHrF3FE9lnmOX0TCfVx7JhCLJuD+HChSZ8QItJwqbITo1P
zUdqDn66KMlUHpkbGmYQT3uA5/d8ZYx4kRBAxNU6kepRy7MPHJxpibPUyWdLzKNxYCl9e1lGjgio
/xb3p5bTAToDi7Xgzuy7z3CsvglE3dibOzK6wkTLiVFS8kMBaJV96dkrMzsxsnQAhfmWULxevban
OJKaUHoVk7qKIRXDe2bDuX/BOqOz/YPGhtndALrakNv+JQKTJKaUefYOUBQ0z2TBw1aUCaL1FlO+
ZKI4wZ2+oTrjEMEQ5qEkPmg9tofcLbbA/f7VSP7b+5/zLxy5PQIz9qTpAsgnWezEsmaNh/ZokRho
O5JZrvmlGAr3ACOnXDHKw5XczUNIBB6FBMKuFl8TSjKY0UsaCRS555K153+e7VaeDqZJwSG1CJxe
qZnqs1T2mfeiXmhro/dYXxi+2Azyut5Ip2uIcFC2+0wX8+QBQWh++uCp2ectHB7fcM9CQcJruuJo
CMzETf7ShI+NPaqnqRpVKB458xcimkXs/rBAODiOBKIp+KaQt8CVGTWQvW0j1kFcarm8W4X9yM3f
HQdDGz6jq+7a8P4lnDEZIx+myEfGbuwcb39SAJb1ZKbihLJv/o1J4ZPxR0i61wmBUONEl4B2rou0
a5SAQ8tGHSWl0nn+/5CulohGqquFRrBEESkn1gHTdDrCdJVgoYAEobrkaVHEsMLn4FC4TmIusYdp
iOYSfnMpy94CNza/ulrGirGGadP900iotxZMRKRFLpkh9YEuUJ61KQR47I7TUOW1hy0nYP0Uygii
9ywnmetDQdmiX7wsFYC78KwpsS1GE7fCIx1N9ym6urHyj0gHflAol2YdjXiZS1d+UuozNJGyNSbI
J8IxLn8OYAq4dxhTixxcqI0+5Rj/1yX3Uo+FhhszwRmbcn81BMH8OqGD5y63m/kkS/2HZ6kwcbpE
CMt799g1wDRxFtrBFgIHS8myBSnOmAZSPH9OQw+xKWy9ScsPNfjax+pxNPlVXKtFmNljU0zNtdEM
7JBL8QFDPSJAx+aOQs8+PmBNxU3GsEYLLtKP/my3akzFKwzr6XxD4CUURHHlJF/1p1Inr10snBOh
WargpEfmOgG3Io9MGnnlUwpW5yGyf5WipNyXIa2E2pnq5Ra7Tvvsh64Sama6A5PHDPd7BYz/xB4j
je/ji54OejSHIT6HGj8QBA1pEaIOqfprb5BKZtA9Di5TI8nGDCFR46TV/9joK7JfB8fkUBVSSyE5
xHy07Mn/eBgW4818WLdXrX/PElpfAbI5yFT+77RiTq/13ssviRAf+nEfBXydPofcUVvmcnmWJ66J
x5IXu0DxJlGAWUHC64fHMrKTp2Lu9g8obdInq3zdemgN6TmKFtM1n9BZcP9ls8bN7cK123M1Vb1j
EfOY02B/mCmCJKYRnCVvS+cvJECcgs8aI+ZtC9lM9sL9xSSeME1Y70dws0ZHPAYnTPnkLIIgrrMY
9jf0vTImXS/NXeYobcBglIBuP5o/MrP/ixNHloogQ9AS0y2kgdqpWZ+4sXRD/uXMQIenAs3MzGvY
+ZGrsS6Qnu4C/0Ysj/dk7oF5YjNqSWrHmWOMY6AV4NquFGEF3GJpPkJyNHt4sEs4ESgyz/7L7Xrk
aUjVfPSNXRlVrzTtYYqYnGv9qsM+txohqvYZsvIK5OH67WWpyZG90+vEOYiPrrJKqNn32j0CGECc
MlsNI8yjMe/CT+tu4zSZLJ6er8/iEgd/PSDxMqQBuZ8gw1BEsxOP37v5RBqhsg6zmLbozko4aueh
CmkVXG0M9NGi/ZJ2YhatGb1k0CnZbRcmN6DEX2V1qa4BYAZlTK/9TbKdTbIw/T45487881DG/Kwp
0U3L5wNHgUuM/06TB1JxKo/3CtEVoMx5vDGGJbRUEKdt3/otiJw3zuuO9R1+eM70kpHF9tx1Z5DL
Yj8dTKrVpGAlZL2YD26H4geBWLKdyPRcZ8WcAZyW3lOFCd8MxqTkU7TcBisSBidv0V3t3FQYC+mn
IqKDWNs9MRHIK8LQqmv8o2/VvbYXY+T1+LNb//4VHQ/i5Me7F02UCvl0Ohg0hfqXCICPrLmogoBQ
AZhqotIocleje0M+I/zTbNGUxFdCAsIcNWc0tI7BfNDUZDQdsAvHElvD9SMlKKUjXuEX9iTlND4a
APkRhSqDvAu5FkHqyL708TxdmE7RQ0nW/uhGICHCid0PiYsHmpZ1EymzUUu96zzX9wRegOBWG8Jm
ZezgsooqDY+SnUm+V2BBInujwau18unB3ctOCG6yZYBf0ggE6mnrUcMLvCsB45YbNAfawo6rqBBl
wxOMHuLBP34AsbWNmglPLnRf0FchzTaXhQjBezsM7ILz3srgqICG/zSdOWnfidZ2YWphbWzjbRgZ
aJU7NEWKL89TDZFc/jn0TyetTMkXlWayUebBsDFDc5wYUjkkIE/ztohK/3Nq45Y9fwwo1/zI2bQZ
Ut5X2LvDp6/KE8oEPFJcs64CtSp3vRUDk2vIH5yDo0Dw/FjSZrpge/3/QHevy5SFZXVPUSmTGzLX
KZAl/Jzuc8PL0+ZIgySc6q+pxA52BYMI2ifBWAD/JXDBFMzqh/x/ODrpX0hOAWPy9fO6zvBUxQzj
7q+Hf3B9ZLBwgXyDATJiigiIAvgvibG6o8a4yaNX4vIZivulxsZqsqANHaDjjXeFgjZpYP5r2kc3
9Iv/FQoFlT9kovecBoKiK+iTyhjkvysAT8XypxW2HwEkEZmoY/nLnvQEg/av/QpuaGpOBdHR6ypQ
u24Fz5oRfRlha4EMafy8RIB+oybZer/DJB3jEIA6p2GiEebQdocR/7nLlT4gR6QMLr9MIeH0lAQ6
Thba+HxIK8W1mmN1VaPJtmDSPvPb+3sEnL9U2Oa+D/gO87mlZ8Pnchdpj2idBH4wD/7i8Z5ATpMI
w/FKl50M3tR8dvVIGwmLXv5RmbBzSZfzxKni1IhxSvI8nYKhrnLb6MOftx/1IGoPl9H8972U8/d5
QR7MWqaIwJjKNMG8N5f7oZlj3f/mrZ/ZTlHUACun089HjR/MsGgnKesM5poYhngujMmy12GDvGZ5
hML/mw/92hdRHV2trGXdzuac5oFHPBTm7I/cLOGoUcTC8WplH5w6ZLhCPLYZihLJ5XCv+EASkIo7
bPq85w/epXFeROLWVRMvQ1/+JhhNi/BpcFQLIY4lUw1Gv0iumHPlQ0RvqhuvLiwtQI4mqWRAn9u4
Bgw3PYEMBLfCMw6s/yXPhwyi+PkqmGcEu+Xle4eK4iob3mEiZe7bjzbLy2/JwS9uHDiDFk58tn7y
v+z1UKhNbErst2TrzftJRksTvnHDDkG28QLEnnOtphVM1pLm6/n0O8ROJw16VLf5LV/M8j2JmzOb
MpHiWs4JIUYFSQNczoi5RXhIkCwksF3nrXwOS2DopcL5crr0Crkbrz32HnrPokpuP0D0apqqLdo/
oUnCLFo9jyAguk4KNHq/JjOo9dGypqcyHRN8uXBeuDRvexjcdPHTK7TjteYtdVU3u8CX8vB8mnVs
wPAimyfQkCF1YyDqTT0AUYk7+PfVe6/ib/lprEe09VEJ55ARPHm/mcSQ+cDqTSjX8ppG0Dej21S5
nFR0dtW7RYm0pPJsb9ho8fouNACpZ20W//fdy8ReOQZoto28l61EKrWThD+WepMd52Iy4XnbWAFA
srbkdOtla8+AJ0zaHUAhJeNnSelgF1ZCaUnIBuE4mLDPDKbucqiUYtW2zFqxy1NPvxcIRLB2geMF
ic0TkAOuNAkk6Of3xb4NFIJ1Yqli30POLWwdv+2gkkzjJLMP0L6DSHxL1l+WGaurqfxu8Nypn30V
PXpFZHbwS8S0FYfQSjUUYnPPfITbLKRz0LrOSqeEbMp3Z7Zu8ZwAHtk/3Hhec9G2KPHNJHZ9MjqA
0iwWzVNoKlHS7qjU3oJ0GZ99drwYUe9/Mx0w4g8OYdH/oRwbJHq1AfZ5tnveonj+0OzeiUSdOVAI
IDkt8ZmHlER0LtFVvWUGK3W27oIzNApCvgxUgP8hzUBBVzmdb8t931u/3hZlzVnCHXu2ht5oVhwy
dNK4FJrjNIN05jI5nubwyoiBIHpQazfyupJ7qZKeukV/4cKE08aTeEGfPMtX3Zz+jpHssZz2ohWO
lRGOlUodRVWZjjElVuLhn3i7lYfaFLe+nB88Olw3o8oE/LGixrXZCyZKTtB2aHjagBoDEE6j1ivE
If0IZqtB9vj+6Z1qrGSCaHwgalBVhrjrCNtmlHb92nGirktJT4KKp1kFhN2TcWrGw5fHigFniKgn
FGHn5aYmBVFqEUZYw0Y4irCK3HuTYMhQ8gZ4yu2XpjdbHQujRvdiIV5TjQ5DNdCzK+/r1ctP9uOj
uiRYoWHnDnD2faIjKrz4JWcwvBxRFmrpe8Fh5nTEwwixhERmfOsxvdLrlAa06gqejhHzQRc/D5BM
Nili2KQRBPD7A5AVgrazga6xX8173pYOBfQw9vs4GH0NCjr//IsHqpNiv/Ddv28J3Juc2y8NMlOi
Vgg8AM2ofvJSTx4Su5AG8h+aNluJzeQ/W3MsRRYoNnxdNqQoeswr0TuThOQTT9cG7rqfZr49thQC
klJJKn6earuxL6PckiD/cdTKOiVaIuKOIxDbXWl1scAQLZJv2ULYXiJJZrmeBPNdIybFQAQ5R6om
nkYhxEOBnUSV6U/3JIxDHuf7xrH4vToNN8UeSPBGNFz5sCtI8XCdOfALF57a8ADbn6KrWejlc0Pz
eCjT56BRL5X5vgJVZrIStrE8/t+VoIAHGCed3EwRPkZRP7Md41pKbrieLeb4XHidEj9xrpBzG2iY
8u3WMfibgusveRh10mOE9xxaueJQUE+yAZsWptKpWGBLLl+o9EVUX+QQb8bV3bRWSjXu3dg7JIDQ
D41RDRbDYRpYSOzthhb5gIOR/lwQeUgbLYSSSqvQIiC4InRNe3rmDhHh93GmAYIWJQTw7bV29+er
bB5MbRYc+audEgodYkywhiwCi4efa04Yx0cKCmodoRddXjMQ4p0PruGppho7gLbbxy0PBk2W7UqF
L6IWNdiXcxVUqP7b2h9UBKlq3F9zxtLGJNOkdRACwoRjO5EhjLQoOd1xtNQT9kHANz3JnOPhwac/
aTrdHHmR7mFoJdhMMOiAcdNNCss3Kwl1otygFPaZNyNOOIo2CxGhXddMMoquJdmvhETWa9zHrEfd
zD0hWR6nw88fJMksIjuGBqHF13bPSjBnKdHEqJRxJo72UgUrwAlZNIlJFoaw8OPY49Wv9xh4Cm7/
TYLKF37Sd7PBEYc1eDHVWeeyZ2n7JQ/ZGBOkavbwJvcLlXNzl52IVIFGxKJ15mdSnqm6hEYi1zRa
IDHFdrz3YoljbxVnlep/qnbdM3lDGsoi3IljDN5HqSAOuJsfd9NnNPqU9kbzY0vHFYJ9k6/kvKLO
kUWzc5PcvXxDIbe4TXen/j6r9qO9NLL91kdk4Iuj6nhoBzJ+WcQ4aVcLyVWEl0oaM2D8QXDeSKRB
rFTF+3hShx+1+aWQv9Qsx1AgzipN8egvF46kOaGM3AR2UNaGrQB/8VeYOaEO96VEZx+4F1h2ZAI/
mbkVuRcqBZe/rP5kD69gdbQrAfhaMiQVqVWhvwSbxU1hTdF2U0N/0DpvU8ii6MlvrE+e1n67y+Fz
Zkq9EWy7uArtyWKz8K5I4TWGjECxIv6H0fDlJLwMHCXuzheVIkq1piIJNJP1vUSQeG+efpZnRqgy
e695w0VeCMvAtYKrgAuCv0N/NDNu5OAJor8LPBR+bgpzmqmLwJNFbiqq8+bZxmN/OPGY4tol40iL
gz6tGDa5sJ9Fkn8kZaaD7qq0WDaTt9GWn0cU9WsbIcjOmDqq3kuua6ZCBUxUObgvvk9D2Js5VwB8
kOuco1wO4D4cr+lNKVPm75l7Ndv0JhQ1REkEysuJAlW8wghZ18EVUKbmc4daavkt44T1vxsJF78E
uKDPybmyS2Zjdcqi1+wwJSiaqpjmQAo2HTxdnlMUtISeHBNnnh/8S0sSykgf2Z/1e+P7kdtDlcYJ
mgo0ZkVCSbU2BCUEW0bi5XPyZcQesrCy10E8bEIAkVgFlqIwKyO1NvuL2Zekmt1prJpunGFWkhlh
YAzc+7D1HZJRjOb6x2XY4wJej6RVStLojOGFJpPxLTd9GKuUoSCDmeWG6PZkuvbWutEDVeqkwUaG
iLxdrEcfj0v6L58I4NVuUMKxNWuFoMImpJnintDjhcu4jGKR1RC7Dum1390r0AvIdU0aueIFA+Sr
+Rc6+hgi91g7ApTzbZVD0mkFV+1qdlBEdzK+Ihxz+adOjuo+ncKqOftAzwUbHYSivUjhWDyQRbOx
rqbsE9XVQKtgG4grqawrMlTuHD+k1VqYavniFpJSkhPHL2mdAHWA7D1nxJrx69bLIWIGd7ow9A+M
ngSm9PqXJkLUSEkiMvgTnzdYPurAAr/KxV+DGVSf8E/S9LwZc78Yzv2H0YCyw4ohdiTATQXCjprF
nQEXjwR0O6GOIid3272fYyoo0xNWBxIhNOVqluaUh1mrZRAmOp0svkpBYe0RiIGbbL7r3OVez7DG
uI5/fTak8Ip1844jRifpV4vu2lXagHF+r4NlcdTc3acereRj45lhYZI6KsRZVY+9jlKHH0XXUj70
BRQX7ulJ2+iKdimewtFbxX+ODJwSIEADGdX1Ou+C7rVBxYhS8reUBe5kflz8fXEySSe2w6D2MBMh
yhV9bKEhm/HfTiHjj8sf2jkBGxfSZwI/8m2o0+O9JMvq1bOyAxXENq0J8tCZPyVKyIY45aLJQ67y
hp3ji8vUQEHGicfpqWuSd/Fi6RbiFcTXIBzdf8nD0dP70BLxndK7MolP1G+MSK802aJeZpIUqOez
wn/OScDeHnymfjZTz+T0Hvo/LuhokyKcFxKV7/UviOFhl4UBiMSxX+1j6dwnkeW9MlzXgLFRV95N
my5ueuwbiHfEuZYmCXQ9Zjt6VnmqWNVZgt+fFmmUHmAmzH+9HjDPwRVwgruHqFxaMwJVeef7Jpxt
YQHcAbBqV1g0izb0W8I15G1MrpHL1nsvz3q6shugIwXoCUfbDhgNYBnF7wJAfQbaOb/u9swvRfQP
oziI6mlfQrv5YU6eLj/FsdHn2DF7ud2qViDLtrMxgGEHZWjNWVmOY8+/vOZMqZP93sz3Lgd/b+C0
F3Qa1ciW/pLPj2mGmkN/W8w/44dtTahUJXcLLk7d3jhC2Mdg3DY7ZTnVTmjSfuA4Rm/ZrLzev9oI
oqnLVHlZpWRx5dNv1ZjyNmbdbX9ueP4ERQvX8Lqg14W2IeP0H77dpG+kTUUSxIgTgtNT3t9hNpLB
nr7XIb+ahJiASdyVSnmXLWLfo43FSOSvAodrsnag+911hLcUWVTgdngWDKv7UzLJ75+2f63aEcSj
v9o3oYkwwh9nTSMFSSGLUSQGH38jsNJ1tQewMDb98/p6JU7peFajB31zrPR+kDpibdGtogbrMAGC
NRW1ppvSxK2XWAWcaaq3qjpsXr4uLrREePhO2/DsNOcs8dB25msFozct71SLFJB4PH48rlw3C5Ic
fmoZSh6jWs7RjSKlQoOnb6Qz76njuog5jniSG/A7OQ9iHyKL3pRRFXjG6LHNJbMXtFDkik6lwYR6
OeKv9ONjHzcn86KgVYEz9kfWGoB8Il8UoKY8oU6pMSh+UxqB5zdEZ2E0uwE7ruTI3XIfMJjpEMAi
xjOavmrj049XX6IqEcYnSB7nivGvH1eeoZ0hQZDEx3Uc8t6uJhTzmCYoauK58Xlh0pCFxcuME9iE
4MPEsbTwS48ANHT0uD2n9kbmC6aG88veljUkprlDeMw1r2g1iAGE5UR3sdmFu5uUvYdPEekU1HuN
S1fqY2tbbX4oS/QPHe56nRO1HHdkJHFTGxA/Of9Un72c5/HABfDCYbSFioWx4qfTaisG6zpLzbTp
TiUav41OYRyIwJxwTkbW120kqW395n/ecZQAegtNGgbrwgoe9Ns6eM/tQ1D+SiwzPTx0oOmP8UwY
lIWuNKc1hnmk7RPBu57qgCe2rJptIll/JTlqyOxINs0c7vlFgM+U33/rDchwIw6Kzcv6JYatz8Wp
NBgh2/Ne+99Xaghw6Ww3Aqs29b+I7WXMsP4T7BVbVTPb/qmMr8Ng6xI/iJ4sMgVc8grWrge0Y4L0
2J/AgPrpMSAcMwF2hDPZt85HkUS5xkjTSBL7XNfRBeHSwCt4+gFv726pdgHPOP50ZpjFojzh4ibo
5pp31jA9Od2qVmCEnYkEfOQrxfSTq6fYV5r45Ui/GcKjcyjN5OR7ZuYWcAd40tb2c5lDecbgeUcB
gqan4pbCYaUsIOKpgx4/nN14nqH5UIWB1O3HUCMucnAlCrXVroM4BIRO94NAirEv6RD6CzswB/BS
jiDMTtIlDzKStOr67TtzWVtkqlH4AqGdIF/mmj4/9CFQNJLprDeCKnTJfM4GjGDgP36VilWsSvlX
oTE7UTcypPndQrRSvnR92T5pfLD5X+i3BHhLHAM5X8vPB+AlUXAbuHYg/bOqwA77bqpbwSU92jId
MnzmroooXmqGvtn9YeFTQqtVIPFAr4fJh/27cswqDyeEkCWvseDyLjWgI3xHNyMRUdcIc3+7EIf4
CtPH4rK38vSJXWb+U6O8hnhBoQwC2yflsAbX+TkElMD5OxqJqvhtmhyO3z5mCg/qDsB53Sxy1G1E
t9lOjuhf4tlwoK/4cwahJnrrYX+fjlQxixu6vyCUmmmlcnRjDuZezRRo8utg6kDM/w2X+nCg9qqb
qZVBjAhxc61+vDJvOzHX6q99uAvqP3xS56lBDdfV8XAPkr60Gikqx4wL+XExOMNHK4dvg1z9TQo9
wEMl1dzvJ6Q26Fj/A8If1FwT/2+ksvR15Nok+RsL0rjUUWpfMcotHKuYMLaHjgCfMAXtRS3VyNt5
PNBHZ5J+BOL1NwqP7jKPNh5KZFVV8CZ0erTQASHCCazMT3IS6e2KipaXlMnueP091dRVZZS4J2Z/
TCxpYd/DhhSQBN59TbECt/oSBC895zV+x39G4bb63Zuetl34pVIErmJtedpLN2Mf0qzgpPyTWWpK
YTT9UUXCdFYTEnyk/8Yce6DLavS9YMAe6uoaC3EgGl4mppau3bMWndzQkzvD7nPoeZICX4/dmd6y
zdDgNQCy0tFEX138fguILGwm28im8EPyHVrSuDp3YfQbEofW+diiZjVL9v2IESf2ssIwFUNx0CaU
HrFXMLQ5Cr2ZHlwtmOt6nA3RZ6P36BI4KJIepdIKY5ptuRfv9p9gtudvjeI4yFYXjnALuKdeVj34
abe8hCnzaYUDJ/042BewfRrNrXsoChSQ204CZm3IKT7170Npgw5BQTSYyt77eng3ESAnrDHmRoTS
qM5imY7EMjTqlvju8ILAcRMpM5Eti/2lOVNA+BAmLq+WduEE7SoIPlcriGlmkS/O0riKawtSNifL
VOW9pPw7UtIItozp2GcNHJB+FaGY1BV+sRz+jVPxFsFEmrPavUMM/IhXQSRWV8sjOnpzYtTI+UhZ
SAQfJvAYGaGP7T+LkM7Ld3Syk5dSfZViusGllsArm8g+19XCtPrNH5q5uwQEhGUwPWOfBEoxWtH7
Lw5waHcLJ922XvoRKTmmLqBZYBIfXzzrex+JrT4v27FzCC6C9WHxM6pX0/9C+K+kFBjdFvKo6taJ
KABRadpjhJspWA3kKfcLKQAc3DYbmJiAvr8XA6xCWu1mZ9tuPe6AvAh1Yk3EgUy/8LFtaJSiC4Wz
u+E2G46ni14rRs+F/UrW9PqvEeTxw4Ws92CeInHKeBhfOejN7WauJLS1j4NXa8TnN4+ZYsTVNsMZ
+wyiGH8W+68iPFKiozv+LonkyzcmLXNLBpGO6s5gW31+LWRBh85qBGGdeM8u0aqlg0S3Cok1IE82
obpsLQSU2lQcM1MwEdtDqNkXbE8v/pBdwnkwa/TgAd9u/N+b+FD8MnlO9+A1eL+BRPyfyTmknhuv
H+bPR2cKOV10Hi8nnZEhZAWA9auNF+izLi4yXXWkv62G/7sfaOv9pdjhRTHGedYk1H9y0Z3QEvEh
sXShIKvFzZHo/X9HiZv6faHsV5lAS5qQxTERVEgMw8IlXo39COQI/LoEef4WK48pLp80TikdAWS1
QLcp29Ty9fzma6IfangdpG/cMWaAObU64tu15MBrh5/RbewcQ5oidkRKgmX0F3rGOIVujhOi70oB
QwtKpfMKTXcoLCyRI5uBevvNfe+QNsbwMSdhqLLm/6lK7qJcwBfydIeTVd5mzmk2OrI29QyEHFzg
TptDXFxL883+ClmD4WaNEr2Alaz8DH/LORwyYmrAMWLEF2uPD0+3lgnlcm9mjeURUn2rGb9JBejX
DSO1gin+IU0WkMXi06UCX7pE0kQnJpj/Nq4qxCbB216ZLtE7mPc0dU1i41EwbIfDa4TRPAJtJGU+
yOMCEO1JqX+jsRbdzjlEN5D8SLpAy0PukAuo9SlCFqDv34syQAUKJP0JngzmEEk4xCbT36R8et2W
6LkE/H2wT2+3TnxmK1ZVSJCnF+Prpr5xIZT7XqTiloUeNY7nwIlvaSndPq6RyzI4pGmeK6ZP0otm
6H0q3F+I8+WBnFl6mplMJRzn9tlRBF1vJ5MHNEG7ge6zckgYX5+L5Xtvw8yNj63lbpYJgXL6Dr5h
gC3hOcCyPxqaXvF2/su8pGHWlu0TkZvcwaIabbbg9E5qDrCWmPt9KAlpG4bnfV1cKHtUy34I4ZxN
FbgTnrJUmAIHa1Au/GH5qhf7wLwkKmgFz3SIJadNAQViCZ2PjcLtkfUVNMrmwHZCFtaE6Frgru6z
xsurTkdxzebbnx0WoOI38miHHrBNfIu0CTfV46XfTbpo68CXJRrRZviYb1sQVRDvqILePmf2D5yE
5hh56I74iHXExsKR3en/BDZNVEerTrHXhbs3oCHAB0htvQ6FxKqFYeegTKOz/gROl27QzMvtMXL3
Rl+yLKRa9B8FRK7VeQ88VDvh7j1tDid+0pQ5C5XFYDd+NDi2meM6Qa3t+teCDowZpVP1hMNWZ9L6
m7UebmUb5Pbe/9bRNk91j9Xft9NPsMSAxDpAOnM196i3cgPe+k1/Zt6LVHpeGJ3zgXl01vMkQBUr
vLKvv/Wdx2bpwfe8Rdd2XZ6VeRF5nV13C5SDyM3+ejvd4r8a1ZkJBInkn8poaxrbw7swdtmEY0fn
5dZDtzEHkIx2pwg9ajolBcGwWlf3suNeJxt5yPMmRjxa7diBMEErHeJAKbd8zGsCgnZXq880TpAf
yAszvm2ICEyCMnKNuEP02Rvu00xXGBQmfXVtq8I+Pz0fs23CYPgLrWq9q8eO3b7UOFbn+Ed2r9UQ
2PzbXkFpThRzWnCvmGpVKYy4+dgXoPa0n2JQGnXKkSea8h38SJUFfyvwOrKOeYUt9DzoEBXzAxO5
FpbGFZlX6M7ssj+CcfGc7S5vMqBejEqhlb5UcZvlG2M2z/AYCtbMjHAAWwrKMGl71lGDCBPk9xUL
CTgRsDWx+KILke/qeEh0F+v5HMfYXKtNts8KH0cElNkcK/VB/tCc0msUN1HqaNSPwtpY3Yq3hhCv
k34f8kNKN9O1EwvO2vrHTsPk78hCMbfHLwLi53zyqlSnimF+BIoppJH31jegqnglY33zCRdZlFCZ
/G6vIRlFUi72gdDBrb+bjlLpr4QyDRflZbWlKa2EgNvw44B58fNgZhqq7BMTzO/LK1Utlvs3j0y5
KTf3DVsQnTKHYnpghqPcp7WjfkzJbhOU24g95kVp7layXQJ1GO7rbIOviywI37gwcb3yI/MLd9kZ
9hWh7zkGhN18Eyhjroi0Am7PtEqYqD/Av5pVsNMTgdeHeUREhcIqZF083D7cxGAnrH0lirCJwSQY
wNLfMfn9LI2zrGQ6BbwJbg+yAbAAORxT0PgO8NfgNmpVfGg3FnobPqv+DL3LglkNus2k/765XArs
KJ0j2QEAzQb1MUjtoxlKMO6euvIydgJVPAnxGGKg9hl31VJfoN5Bm6Em7J1lDw07uIAS3JV+Lgcj
A/mMn3m/7mGdmWC/Q+ZV9o8Ch64Cb0r3Q1UWQugA3Baj0Ww6+Yt4dvch7nRgSi1c/kkolYU0bkAc
3rL2ehCcn9ofF0Fpe/0Bvew1+VUP+UMtZ20RkrQN4Sd+MJ5OGPmiS7JqBPe43kriaLpgfykXZabR
mfWhL5wC5Edy6fM2o8O71oPrJnjQAY0sOOENagoo5SnwzS987EUaqXcsB4gJ6ja5xvjoMDYeloOw
NEncTU3kYUPdlqcOUIaOpfoJYion875j2PlFQ0tB4XtLCPCGbg1PLQFejM9vplGVWDo8sIgzHHrz
7EiY0kzdzYksfJ4PmmJOYL4p8jOG29qVcoCkKyXbT1/jrngbcbqwfL7LWoz6sF9Ta/kaqrM3EH46
IEiv4y/AZGe0P1+PDJbSM7i9PggRqpDAJ/MFTn17xfgnDnOy99MCcfZvOTryigSeyTun61KDxppE
DQV7BF9kEWPFpaIJK7ibPxFCFQQGefbAQUjdohxO+pbVCfREqLxU7AI5V7Rlgp5PAqplyqcletDu
hGt5ZACfoA+CAd8j509qrw2KgxZmX5a5v30NHW8YdSpXcdsu4GZZrD+I4VPrsBkBASKkxJcXv+yi
8vJ4E1tzUptqTZJy6Qcs9nLO0MwZbL5YuwiQdY/EQQf8ekoGBmgaJGDZUOkjf/fUQEI44gA+s51k
/ykVjIPfcSHR3zSnTclEQror6qGm6nJVMRDuU61kYyzjAW6kWEy6gbNEvn7SP977IIMWthyzMSao
QSpAfeYKIzDgKCjB2uCuxFmASYpcR2zEKcqub/CirjU3Ml+WVo1ulsLxmgZpYOgr8AMLsAGkCvcB
DlGg6rA1ElxrSl7cU8bNy34WpBB/jHJsi5kvW6cJpftsitHbpkQCIrYlJVJbRWVt2xIC3/Oa0RI5
TZ8agUNQf/XWjKJ8PHaIe283of0J6l75Hpc0JkONVlmUWVCRfkR6bLWhcQZT8ACoIQaIZ9slYxie
ty1jmsnbJQ2s+XNCS73z9jbThQ0mcb9vYVV9Rsd5QQGsSU6wSsgWmfkLm2oqIRSpUKEGgQhAT2hW
axYsRf16Nr/NuAeXEWypvipk+dpyc/VrdLyZGVlrgSSs8CCrgCXNKGc+Pnr/SCebLkGVJ++3Kv0Z
M7HxGZtsM8DAfPxscYEkXdCrvyEKxF2nGtH0Vjcyu8KY3q7sRHKfIhkm+v1P7ffM9AH7MVRRAKLz
L/UzMDZNawtWXwWeUAf/03vIEgRf0Rn46qfxcUvLgyXd5wUwlsDbhdXHNCkpg08i5NVg1G9n7SWU
+3ZHjJ9OI4aCJ/uDpTMOSbDzm2FVcRpHZofWE2B1RGHy/u6LduuJA7GIjAHfWyHdL92lKQGWtiEq
HNVWm3bae+75LS6xXIuGWoz7lVcawky6CeBX7YW2bpLU1DaGq1in1iudsEHuKxqdtgrsnvsEdNYm
OCw1Zh+cpmK0xVWSnNUSVVgFx8ldEmvm365m6iWbbV79J62xGA77qN1bnZyzUwl3QqhUMXFcvpeD
I5rm6cciQEXGA0EKJWpTGhqLp32XGBDm1KXz7n7fBnxUoYunOtSQ+bgBJG6fYiOw0kWvBKw+EXDQ
JEW+hO98mxfsJp0UQEOZadpUCOV/jbuyJLoT83fZ4nVIfBrHrvLhvkfe8hxrWcFwguhuv5ZiaSUW
bwU41NzBqhedoP7NV+UVBXN9GCVldCKeeqK1zhT/WDVwxX00tUYeqk+9fu/phR6FGgg1JXEbb0HT
nuXRc78HJ3yVlVf4gD4u54IXCFWU7B/eUczV1le2tKv1iera4mJ7sB7rFqGOrogTKhSscdMhs+CN
QX4gsYbYRwS2JCRhNbbunHQqNMg9cVrxZjiszjIXPbFwUIj9umurDouAqScmkoI/R8Zfr/G1vgFn
CNQeb+5DWqedl0ZSg9bl+i5KNznGQ+eTCChXQzUI9HR5L1w/QP0FmsOJa5i0xaJPz5SXTtrk6+A0
2gKh4itTS4mNQfO3hGxxaRiVewrzgbnOAdupOYuyRqUNgEvnHqF+036JHpbtpRi1/D0AErEx7Dye
HigxVI7ACzJR90S4hNRHLdj6a05GTwqwy0PWxmIGjFcOVQXIFptTRkSw1zwXDKPdvUHkLCSWtfRA
SNgcus/iAtRWb+hAcODZ6JspWA8KlVudaGDwGLk3bCJKOgXcfwc29mOZ7qE9ZQA/kOQe94b9DpfT
yJ30Y4vfiepzT83tKt98Ctk+3yW46rQb481yf7kIr8qpsS1CuwgGTWIygKmGdrOuuS9f5ghLY/sK
FTW7V5HMt82jmZFOCehvNQ1K4fkO9dt4yQ1XzSN7MitpvejPURNbtLrHMUsVtm0yYcFPkgM2Z+6k
I5Qm+rCt67aVxNyjKDOnnAuew99Ckvsr5WOUTqFaDeIpRq0QrqkLmE2F/rPPxgsW8dG/OMhiTxGp
YOMKQG21gnLpzkUX5JbWqAlC82JI3RLgV0fl7m7pwcDnS7QZ0EFKN1I8zDSjvs/sXnBejZM7NTiH
wZZ/9aW9ggcZttNc51fbyTDgaRDCJzGdbCprJu5F5241wNC7i7ru5TixJ6JU8oH3JX9YhX0yIbxI
b5gEOAfHEuKKESre6LQ5gqDMA89gWcn6K08V04vLl10J+MWkjgNMokahM1B1sPznHOdlHTjRk1PN
XYRUwGlD9BwCDvJASnKv/EZF6ZNiadZgTv9/9p3On8fiXExwDCs+Dk7q0SKF71Gskp1wv+fQZwZD
zeSKo0iu15vEwwXyf/sFIGC/Tyj14btLS0xQDyMg9xnFFci+EAjZaDjgJdKzqQA3um17RB2RiDDc
vDclXOlX7YTjJJvGa1izSGe4j5kJc72TLIHb1K2ygzQlJZJr2cZkeFf6KFuZgdRLcQF0KT070UEJ
2IXf1lqrtw2f+g9YIf3rm38dOzSzFDAfe4Nz5Dj07LnPY8OVU9P7+LgBRsPmxZItphMZKdCfwlCH
sqIYaWNO5G2Ij231siZIi7j93Z4K7TFFnEjy22XlEW8wol5DHu67hBBDQbgV5TM8L3ufnm81nRBk
2j6PhYpT7+cAi7IojPSc35oBDLf7Pr23TcTzEj0njqJ4E+aoSRquiPg5ZVvuwAzuhnjvz9UZ0dZ6
K+8k51SgvsuFY1Ll7xmF7oeDiu6T557r3iria3YDNcpE8IR22EWuqtnZuzYRAwNF0sD8vObGu40Z
xzBFMcq1p6S/PJ4A+1U1sanhMNMWVg8h+IU2TKsYbiyIm7od4btgcQIW23YDUJSwJyFVqm09aMPW
B8Ldf5YS5ih65mZfRwlMV0VeTKgeEuzo6pXpI7Ir/NcyEAVjk+JwhqI2gXYe3Ea29ga7dtIjnSO/
jjYIi/Y1zQFRqqtgfl9GDaShK/+t7ngjdNMY4qqJJMMduYhFM+yPyqsyqPdw2N3zmuTrm1f7ZMDo
oGXqyOLUCkfVI4F9n/WFrZfCIoDvYSs8tbNc9T/hwVlxJlM34D2vlt9Rr6Rh4nkToOe5d8vaZ4RS
cBiFp06aBlhAXrwSnHFS04npp72eOLatUM9zohCX5L2cX2o4FS2OVC8F6AKy6hlkpUdDmmKcvpb6
46VO/1msQS2MlIZFRFyP5KQ12hFUsdDbXyn45R2OHuQJuOJ953VkEQeN+T/l5F/5cspycncJ9ENG
4IlDtClZ67M9YrLa5DyegEz3KvUEOIo3RcBAruqpFLsj50cxy45ctWVWmT3YtS/NsMKe+XRRDu01
fvBloNwqsSz5yWg2duhhY4gIRVShoMPzwIsSuyHeNTNMB3OxAA+56VDxXY6qvUkjwKPYawgmyLd5
apFA1fixOSi7d5VTn1lX1oCIdEnZMthje8Xb0OpCKlOl66dFJUBSKMNV6s5QzKoV31uukC35+8BD
v5v8gEvfF5CdE66AHTKJimHvx48NWfB8evybpV+lg7gAxn85rUuKwkbUf1zzDeqkkV/7pslbaavE
ImSk93O33Agm/my8LsAjdbsW3E0aGVzgvMH2hmKbFLX9ZQeL1wtaoC8JUxxorUyjpM/WFwOAE30c
9BrIHsvo6E3ZsBbVoN8SBbgpBTMXVEdc7Q8KC7GpuXyvvx3mDn4eB45TOmsIavxhUy8r5ATMTa56
IM9uZ3yrpDxjurzXHjwG+1/dgFJiAIo0pOrGC8XMujtwGfXqq1csMjtlmqTL7a4vbYzwy9Q3euzy
26HkpdGXUFmKDlIM5Ndiqk8UC31BbVzMktofruen0fBTW4fZ/bSgw6HIe6j8CrsoeyTw2S8jDPw0
JJeajbQUSZDP2x6TrfC7QR8ZQO0vKfqlNNqBCVDQcSHsofQDwHWr4ZsK/ASulKrENMeRODxM95Uj
QG8eYfF4zxRC97euZtMkObzwMOJYw5MKzGHELeok76+DU4Mb+5xcV6wP6TQ5X5QQs8IbuIEm/dUo
Ie5tmSiLMacX7kGzkvEgGJD7MdO71q8HQ21jd/zy5K9BbYRSea0xIGhRHytpaPKTFjVmQVocMh56
EyV5mXMfAp6cf+hywyS6k2Zgdv9DQ2GJ+gcRNBy2Le6uV8b7uZLqZ5FmMdvqRlE3axfBbU19jqXd
dwx0eeTnG93O071UUlic4BXKCI4lcKd1p9HmOKf8BlHkHc8FctAdyAErBMUQcNGRT7dUu4ski2rA
W3tbciO8pAkSXv1dLfy8ikihKlxHOIZRFvYnMfDiq9jpbRpd0vHDUtffbljkaNrNA68FAXtdl14q
sECdff6kp3tc0KUm+NV64PhKC8MbY8a5sT9DWiX/uzSVtAmHSbRW6/TaEh33rlvt0LPp1DosFLCs
RaP0TnoSW7DtJCpaTTUeliG/2tYyeF4ttGxShzwBHRGHmf9Q2EzaiMkR11ud7MNdtRL7TmYjeySN
+9k2SOAVpaF0jeCKmFarD5K4im45oEgkW8UKFGBrPa2ipN9d1F+1nBNyFnz31sfQTVDcIsdSGW5B
i/C+rUCnnfPQ+/Y7XGFxMiAsJU+Te0TPigm+ncdSl9YK28Rfk73urqwFaz3LJg8A6X2HMTSTqFwt
4NVJ3i6jjJASvRpzrmEw/kQ20PgXX8uKS4dbrI4mgkAxWcv3k9fHahySUIybQPJNTHwYiT/BkOq1
MQDPyOcp3S+PyOdMSjzPbKPhT/tI3mHnZAq5vwP000qnjMTNzWdFIej9zzMXvW2xPQVYh7omkt3V
kvZueHd0wKQbnLxpJzE2ESTuxa24tEyLwsmEuVOgCq7lkPd9XT75tDrp/uzfy0mi7wEg1qkBzY37
gyUFlGKUhlhTEhCnQ3dNZKPTeThEr4fyQ9QuKOXsmC/AK1E9VEWUN3uxrVurXst5xP2lfBkNUQUk
rtVi1g3JWk2Tf8XdCgnKPomMgNkMzXFOIhd1VzRWWvcneUxbbDcmYfYwg2LWgo8i4c0JAw5w0QRL
9umRqQkz3U84lXtcSo957JBcEwhJzOnB5L4m1FgPaDHostxhtnkx4htw5f1NCqnqdpD68NXdcBFp
J8UeROvObLYrg/QUobDj+EoQxzl4KUskSr69sS6uIBUeyFLKRTte0SVoXzMMtm1/8z/exit//4Un
efaW65x7Knd/t1Vb9hb1UP6YRLiAUgU7NXtSriPu7KLSj+ky/dV/adzkDBrUZssWX41/rz1LodUJ
Y2xX8A3WNUzQ7hGdbdrifUiSE/N1595RFOTLdzyLDS7hyWqJHrorPQlnPdBtiJDeQvqog4Ojr4Xz
tvpZIBZUHJKAdZAcvejGsoHbvC8dT0/hh1WFS9zC9dhbsFkfnojMT9gjXxGEOwU8Ba0UDuKhcHeh
wmpLFzMhighyCokbeV9onSNZ6R6yHWNStT2pqZzYp24dQ9o+p8yl65MqcL5hY7owZENAHOIEF6Qx
Kx/l0/ijEY6RlNE0tzf4cOf4Dq4zZ31l9S6JJ8BuS6thEPeRBxpd2E83SLCmDe/QnV7g+OiQcd7W
66REatCAIkIF/PMMNyE2H4ohe99g1EArcOy2iJ2qUzMz3inAQjMSXsbCHFjBwb4kV5OZalF2Gtof
rwAuRE+3DjKf4KhVNxKOlD1Jq/Zdtiv78lg9KEm33Y6iDbgtfq2GHg7LEIQVGg+bHCl6nSp5aY0y
O4xFWhGOvsVG38hH6AluZvNb2vakJNAfAbg4EzBZSeyPs5jgY98s6QHhIqe6YDll+tLudSBnpBIU
oZuGyShJMMNxOF2aNIOhnItgOspk9Dlq23RGp2bnYIJqP0S8HXrDpozY0NDfi+hdjGmOVocF/heR
Gs96Ho4moT65ix+FOTdLvF+I++wjMc/th1O6YoVu/Cfif3Xg+mp2AcNU2bxbzQrIygPHGs79Wjc+
qa5mr7frKSXaD4mjNKDgnAxFdGhZMUwaw6VcQR48yGIQjOsg5Ij8ePXRi4UFPbfgREq1WakzG4fN
yL/HM58pi+WVzOhXDgKFyaGlR9ujZ+EoEPE2g7S6Jxv03EtyY9swWkvVtfY/OYzEx8tRyX45z2Fb
/tZnS+yRbLNVw1Lk0uG2HfOIiUA4e6Ln7NP5rb3Xsw97in4vO5DGrx3rRngUjLJNC4HZd6bhwkwi
7J/ldRjcVUppkDQljtzzh0VqtCmQ5aieE3VDgkiHSmDtluoRSgAqBwvg81oC3vCyqBbHC1cwjvQQ
iq7I4AJZJljeF3QnThAcTFKCXkE66qhepJwIaOanoiHqpALeJOEsAKKko0Z6VDE7vdO8ziVtCn+m
QxdFVICr5r6BS90hTjQNRtFWQ+MQMhyE4dgxNJMxq5+9btPWKJMDIzua+XsehOMmc1rnwrmMiI+L
rmtEYXBG2HmsehFuhhgymsQA/OV9w8IAEXxW6OamETWnn7IAd2yNct65LlOIRl4BNg5JIDC69KIo
4D97JPmJSYTpK5XOd2m9qlA2Ot5l8ot6ll8M+s6YAsD8H6BrVNEC+6Rj1l4B9JR6qXMnsarowGMI
B4xuGuLLrZRr/zvTu+ew1sBSjoXqzLXALcSSfyBcWqpS6IY8GIU4saGuOZaJRpBVz47ythl0ZoQR
OZoVw+0yylcdTi6DAiAUti16QXULHMbd3NAdumaGvkZ7/JYaPIpYcYwAqr1dSTrgMQSe/Ao6cNGR
Op+1dfxIyA2ApJsQI/Ai5R4VhXP6iRDsxMPIoQcNMrp/jS4H30sTv9OYp7zeS0msT+k/5Ah8RAks
L/dRnoirFC4PlkQ3srJLZzsjLNXt/43eMIVgVnXJ2g+TxDBkTwP6DM0mxPNjvHJ9hrsw3ZGCVvlw
ARxV4sb+mBEf9rq/KZvdbtUrx70mVdvY9Z6OeKdj6kxC/lcLFn79X0T7cAZEZ4WvhqmHp66P3O4s
Zikw64moxCGK+DNYVvVWN7N4HcoSLdnuIJ4KOUpsYjp5JIK7EOnssCxXAYbaId0DU8eSm0IneyU0
1a9MFWfHZIJA13a+s8Q3+Wb7W0Oni9lTHrGr8WzMr5K0k4Lr15G1aHk8KZ+nqiJlWi8497hBx9Sx
uW3stjzrkHLsJc/BThTidKaBTgpN7TZ3fIoxrOXpWH6vHf3iZuwfi3kn2jLl0/W2gMdjblNNmtjU
4Z2aCs99Vq7vNbM1FIEoXfiEAnoAGESwsuAfkiEYm2y9EDNjuMG/WkZOGRFChaBEQW25AB8Di4t2
FvyzbbicpNp8rKI6zmwLrE56ZuHDTRDGXB07gqmlP40vUfE4uE0h9or8I4pG0D9sCg9AcXC0t4GQ
3HInnPHfpUB0hcb8BQuSg3pjyDOj2LJSGWkM/cGiw5Kl11qScZ+h8oUuam0CPK+y54Z76KnHOA78
KM5DWwNFp76kENnND07DgcDLzwlFj4yf4IhOg/lrTeTlO4HO/19FktMSt1XBWd+rye+tbsR/8SdA
z9SbEC46wR4IjQr3NJE9tmyzpk36PfqYX17ss09jmB+khPN7Bk0sSVwPcMkKZNKWMOKrPHdlB5Ld
wghgXB5/+29PkbQXJsVn3COuYIAtj+/M0S4PVt8oWIUdpnwzBjsdte/MAhPfQgXNuhtZAGYx49x2
L6T10rlx0vtIDPoMQdQEDINTzaPysOtl7LyeXgelFJzYOELEn5rP+2uFMCeMvB2AJ61ZNO4tdPxb
w/B4EYgM8aDNWfS3CmzMRipTyx6CqRDiuxV3hOQ7y2XnVc/4k0/ypOZ2vLlXeUfAbWqzyleguFxW
0sSjlVQtEzWXxKMjlKMqI6Xy30Nu10DPjdWP30ZeStqTuEshqJipjJgCkhgYfK7x4zD0r9sdrAsf
BFuGQa4UpLuDtAkiSrM4or/OOsZToue9z++rfdOvX2YJyPVd65KQgE4ZLhe6kaLx0Yc/gG65VGnh
7+ZZNRoxrmuEUC6ZyobuIRnAJcZzLITpercKiuyxwlgaee0rkHDx2fmb0CJkdL06T0ZxO8/TMUKo
6BgFRhGcD1HibjNnwqonASmEOIZVCEzRvzz56YcYzJAATTdxSXgSgFDpnTo9HA+onLJ9WZ6qnx6n
S8aHpl6+QwkE62iGpWMpJzuD/915aV5rH7caTsJS6EfGAHLZluOCQIbSnUkG9iLte9I1dq8gkNYO
JR+fD8ZRbCp76a2Z0ECrshANhEjb//L0d/kdYX95cMz3mC3ovTMqNRt1H+LqJfgt3DUoCKxtJKUH
bscwI2R1Q/nP19CWEsrW7iU4rAo2OKg2RLfyGYUMkL2F5iIDuhlxntpn2h+zCeU22XXlTByaO/NP
/fY3u6H7qXnC+CsAcENU8jVlJ0PZqNwD2cI514pZg/Z0MCBn17/OJXOfpYTfJKdLMyMN3QFeyVc1
TUZ+RNvcuFRxApuQ6PtuCMpbnc03Rh7/xkrKWhjEfnAts8+9K7UmeyQqJlwfxRpxjp1SlMPzz3uI
fM/NcckJIewWLxNqSyCUgNky0VHcaeAzIn1Ip/rFEfCpRBqoTjX2du+Ms5wnKDgQDihHgrJvd6w7
WIRvd8qe5Jk6EfsyCLMu4Y+XbT6YY6m3DVTunH01O+kF4YFd66rfJiDT4LumZt8SR2u1tdxGaTQ2
N+jm73uW4Yd09KEeC22hFzl929tPAVn4QvTW8joQq78nbvGRDozKQKHBwrUmfDBKHUED37wYnsX0
yn3MSsMepUpSXXHgLqYKNl1OSvE2WVsUOtVoVuMm4DNTcHLQlgaGUpljt9cJX6/nviYu9kJDKrpg
FmWmHMlYS//Keoh7ygft1to61vvsoBez2umFxbPaQLitd5D4MLa5sKTn0fOgOZfdi8oQfXzo2Mh9
zgr3JkyQW3nLjjyxkqxkbkcg16lMxe+DeGtRcU0PPHt2mg2mFimQlD8x1T3JkGDaIa3C6QQYdVPr
QBtNybt5XVUMi6Oln/xAhKe4UP+XLv9+FVxNONE6Z4o5O+m7Y6dzYVGxbASbBrNPlUVUxQUGkXck
abjNqB9jFkEDtVIyehOlgK2Bkx6jZC8BMXr1/MPPMD/5iGFx29vNF05jmd8eEa4dLTB9327emvfk
L3z0b2KZxbAxYj4iNQP4hQLU9cjPBEavTHF2S/gjyhiUXzeSkOyL/jqD2trWQJW0AGNImSMBEco5
x3n13votleMmbzyloNJ3StAznnfsW+LQZmQsYApMFZD15937MtaOwqNgJqmW1jsuR2otKk6lR+0m
k/tOCSdXekl67wgI+o1lBdU0L8AgRz6cy6pzyqTHT96wulhiu+9xXEnfYFsFNv8QQBrH0wnMrkxb
Y4jDy59/E1pT8IVwcYd+z8vQHL3VqLrqgs7B9AZrsMKhBmTqgMYRfXJt5skztOInGsNrTuqEhdqV
kVQdsDkqnzORZh+E5Epbv9nqfIEYgtNc+z4MSr/SYYYRMD/dSIW/IFmnECNWSiHIRrV7tws4Yo1s
Fdj3zoSbMxW3D46BuIDaFDjvzVjkw0nWVW3uUKO4t9oUY6KeiC2jIJAGQCzVHAeKsAWINial5bbS
BNKDPhITf+zBKm3AUzK+GB9C1CJ/3RG09zd1o9l62ZQwt7Wtph2Xp/tY/jjFGYLWI4R2E5wzN+HP
m4PTmKazGbJwjUpAVWouA7updUCZYJLkStPgjo4L1WojC9VeJgR6knoC7ZK8Noon/yW0OlHq6G/e
YNvZA003lDez5fI39q5s8NXsIlK62VR+Tr8QnuPJkefIbzvn2AmequprKfdI1vciK5el+pMMNU/5
avLW1nd4bODmPbSmEyWMI69iWGDdVKf+hLHzuS6MmJzYRNjgSWWXXDBHJmxKEDCve5DhNrKUzJSj
NK3LcLbLpUYYvnjfmfH3k1q1dYAhaW1pmtv/cH8gdIE0c2VCXSjPYLO1J5OMKqUJWH6/ZXxsiBxQ
P6wZCTed4PhZGbuiTE2U/Eojv3tTWl4rMY4CvHNFUFUg2M5tBe8FnNM9G+n2zOyAkD+KqefEQwjE
9SPaXlNe/GWioToXTustH4KoJN6iLn42eoYsK1dmrxgDBYjSVmzUJ9KhQO/EW10fzfnpWmte7lkW
sa1qDB0iYuzTPCqFJrIC7jB0aOFyh/rk2E6rVWFXP4uNsPBAjs/JAYwBJPOkdz36x/p5ZAkGReAa
Ul5gtc7NP4GykKH/13pRWwc85MZXiqUGI9cE1myvRJ7K1PsIwyhTtquZUW08Dqd+lD/57nymYXlA
HZah5g13eQNryPlup2hsNK9/ZjuuxJn1OUePxG1vOj6fJSbK5MAubImm46aw7ttmtL/E6EzatYyD
+Nfk2fAtbKY6xHjWsGAJXZqvpjNtOOXHuj6M7cYKXhNrfTY/sW/9aWhqL8Up1PKAhmpq1mgQqH3C
d6mkY5ero7j+T2h0RGYmh2gZmvGWLBvFafBiTROMnrXTa6wBUzsjfpUklmYiZPhwA7xdN6vdLw5+
L784Klg99frQ/2mYxA0F1FItvOvK2R+ZL6+5eOA+N4DzsQ/HDoTD7g3qbXIcRcGdX209yYLW9bHg
zNJUIUj0n9I7XsoftmAWSFtWnRY2GF1/rMHO8hcmaPPEIu+4cA/bfY+d1oAvvAO4Vna5fzeFVTwd
KVyBkpLR+u1e2KYY7nlkui5xhjLDZXSVYdp/0JqDvFd9wAIgMfLQOZd882D28wkE0ieOtM4IE+p9
db2495F1P+S+e1bqwN6oNib82ktVnPa3t60IkiNfed50PPHaSvs6LRqKyo/axxgUf1DzhMDsnlWe
wwFzMmh36PMtHK6Bejb1+ZJk4aZtT30S/AVsRu9KxJonc+cumnwEbcXOlWhObqRvj24yXTd7lDdt
Oc0l+w6o1AtTg3CB9wAiwo/vTVToSp5n0zrWTfAZ0kFUNxj0tmVNPEXqG5EIs1JYbJpS0FIwCy7B
mK9vSl3fYkxaZUHPalOooVElNZhrFyuf/MARRZjBSFVOEUVUxSVVpbQy/FKIZTdhuSiyxOJQWoT/
PD16tQKPYU5a+hzNe2cQvvigzueSQa3TkuoUy2nx3OyW903ZOSNJARyjMGJL6pDUPQ1S6iz6HBqS
Hs5iDxgYXIacnRkuanw53J7k+qViw7rEza9sctBunjWizQdNo8nBswKgF1XxEmZVRuze+F3hlxEZ
NUQsIU0qPpILGJVEYtI6ido5qbMWeW9AIou5Vq6e+0E9wQDCVXURsW5Rj+4Uhs76/2eBvcQWIwlZ
JCjmR3KxOkyI90gGlM2nELcTQ7zN1E34HMa4XTi1GUHMg9rpUwU+ZV3XkvpG7ocZWLWNhX3ywroh
AMOEAzYqyJOmz7NrVrIo4UbLeTXvEUf5332qxeCBSEf65VhZMU/PNvUiQeW5ey15NKcgJSeiHuMe
9PfhwS5/Ddh48I1+BrGIft8DdnaFpctgk6prD7Pyvw1kfZaDP+BE6RLRC4X7FyubEHnm/WewQH8C
uCoXIaydKU9hLlBefsP34h420idKAKBqS1nSjJOG7GmQqLW4c+dAmUZx59UjnS5e9PpL1i/2x6O7
RRFCr784pEV8LvHIz5ZtgFkfTqGiftdHDIsS/vgg3/Z2BDod7Q5lRIZPL26C8vUY+EfGFzXG6oAx
Bp6poKAWQVWS87O34a4xBTbfiN70bjbO8C8rUcNE/ErLni02NPe2n10RQIrFMMKtiCw0WdhaWHlp
MI2LwEj4w8GFNekINwLCKKo5j0EC/4X7Skl6+xKBJDQAnvF1TzUO1bE3uxZNrWB2xOxFmU/zLYkx
dooYXomvIMCuZRWO/JmrCa+ilT2w3sDf0HjGmSV/4/5J5D2QVDvtqc55Dvj4coB7oUvqYMWN9cwf
W1xrTHF07kJLegGnY18MqNS3D3HYx6+qjW1fAWV5IDOx4OAi5iiR62+7KxOqqmX339qPMJ17nvhx
hqMFUIu3kS0OBk7OESMSI3IN3Tj7jZTWSz4ObnVhaJv7WrnDBo4p/vvLmzLtqLNQxiaalOfAmplq
MK0UrAm9awtZWorAeup6ahElqfmi/eqZeDGWo2wiAtSUitu9i3hICmNluTj/+n8HOQLC3K6gyhdq
QCaseatVkWz0pjacxy/fbI26/GIC96LXTj1Y1HTWvrhPZzPaXq7XgslExMqlUIHsAIUr71MtVpJO
xY2uKsGa2uCVdXM8xbTE/Mg26nVgCZNeEenWPqAKgxuK3/kI33fR8+LWx6hSMzKDNV6DAnCgstrA
4t/uGCqpIPlBPasYBWEvAPmuulW+jgooT6OMyEZa4qAhYgUvS0zAAp6HW3VCgPRRXLX0pVYcRVWr
WRBFlYiVRCo3ziwhbUMFxMpwLyUmHf7ZdnWxr4yaa/gWrxxFunqgoYNl8xYOpaa6R9z8zaIow0e1
v/4S7H5w9hn0rug4YreFrUVwGcmuiBoEIMhjEzOqG60gmTVEdE4qis25XqWscvul/QBzkd0FLUJ/
uEZdyiRb+rVOgBYLXti42yBU0oglB9RjEUOTfuN+MaARxihfZTNACQ+qWCnfNpEmGQ43e0f5rivu
BAiQMgTh8j+U2gI6uPx12Cvwk+DjDRykJcgM/75a4ZZmpJp8Vyz9HFUsT8EO05ljXTut9+9bgl/U
g6epXhsuOa2b8WSL0dNOwGser+w3qH3gBwVvcYvF3xFqiOLaBWBCKQ8TmWgNsSgINBmtYR8WHsRE
FxAZvKtEGHMf+v3vwj0QxLB1pAckq9IXeDW2gM/1Tf9TjnrnGLWkU6PqXL+rlqxcDuIn3kivwUAO
TZBlZ/kQRvFK0fkaGnGE7B/u05+jbxP1g8xFGwcGmiPqfdpjMr1TiJcVmXrdMTdEGODiI1yA6BFD
FJw8hlf60W6kRdOnjPHTqQRSR2RWFtdwt4NYjCq5mA3/VnALrO+vQP3UZnEE2D58GodRgYqqmgeb
RaKmj2ppcOEkbmk3oufvyzn/AXHyjqV4TwQGwJW8Y41lZ8wzAFRftmdyNJkDk3xCFj/QcnXFgc52
Vs1ebj67ieaANVpJJg1tMH0GrW9/0dR+3+/BzbT/jW1A4VPYeOyUyXB23BzckffNO9Nnp6gXIGZD
v2IoHqYCrwGd8XRW7nLuJwwPAtMQxjij6in+aCyTi44Vvs9/JTAyoqr+QHRvBkeK7xan8mvUalVM
hdCek4bIyl2pI7d7Ugia4FQ6scsHxUP/pUn2JgQPAmmNi46va+N2DRkZwC5D/Z1ROt9LOqs43wi0
kdN5fss/5usBsTdeWeRynghMD3GSr2wdueex750ml/bykE8ve4QsvHCUO0mlqWvfmlonP2wMAW2r
MbXmhPnJXtHVulZNntC87kElztlKokYIjC8DyCY8kb8v2V5FwDCh+NkI0W/DdhQ3eo/I1Gy3/JXl
qXk5uJtcJWjBbxAr0zNT4gcVE9tJcOlcFzMziYCyYn6hKcMA8Uh3Y4qF61/Y6CKJbhWvsu/BU/lJ
Ipk+W4ey2zInJrKthV2XrGua5nB3dODVXA15vzLMbKHSJC43gsaO96B4n950Na9wnFu50JO0Tta1
qNTFXSFrMMzpOm00bC9uGym7tdYkqNDSiUfYh6GrPzN3fBD0g7sTj42+1jfh4vEvrNf/Z+H7DLPh
TofYU1LSHJjEF4QwIQMMMTNGOtio3G7KjqpShH7yNu16KebZiGdlx5WIyNSOqjIOppF745aYBCAI
t3/OuDfMI+5Lz2TrylAUmqu91Ry/DtRbMejlRQkBnCN4xI2+rst3v9wovrBMnK38CJHrMzD7fGRI
h1WCQO9MM6hjZBjnMIdQinvCR1D+qIhMBDX+zZsRLNe/rQURu35BQRG8KL8V6bNdzhBk44B8TY59
mxRKQSjSIkX2lyoaZsen6RbIiqEqgw/U6cES1SJpzNOv+c6my9V1S2qNbLnkTXEmyjtHcNi7hTs7
fwoDTnHLNSdHxJY842oNmGzuVhRS8d0GgGVo/mJcmr0uYmnm/UpoqkTq10qNPuArKIXt3MTYEKQC
JwY/4YXvZLSiF1FzMTOpVlhu+81KCFK8exOP1NFzaORCjKcz2kcmx3iAgfkJGbkh0P+B3FXsMivh
wWIRYP7mmH/UA+5wy9hKzW8YIQeft2RTBdDy1MwJOqiauZ+FtKhzPvQuO5xRjOmDHIKEkXJKHCV6
eypae7adaQA1FzeOVf46cns3Nw1o5OKuYtcmunR6YKfSSPulErFgLhHEOpvz2GLPu750odnGxVsK
CyUgTsg9aGxTL8PD50PqLPxZ3jgXt0CGYx+VRlQKQOa8sWriz/YvVYLw/qBkdT7qiSwRedy4wNdB
gxrytQTSiHrZKTPZ5DInrFpHTFBfu7kotHGx7fRx81tx/0usUjDTAVQSMryF2GbizSsv+xcGfw1Z
mMe1YSfiieV+RzA50eSlyCIO5Od38BJugQew45Ze6pZTpHME9eLnePLB1OjG1HcCsebksvL7LAJI
SDm3CvU5uFhcLQe1ldugASXEs3m6X+MPhReQHSV3UZy9Ov9gOxbREBoGWFQ4D4NtLumiiui+nk65
bjnBLywm7FElo3M4Ws8EnrkFpzQ7zcGht8QQtK3wtQS2M/N3Hlz3PgCMCM0LJ4+nTrPFPGRFI84v
5ErEbl4n3RBEdb+PTQML7tDpRc/o/yuIzKywqaRjKdoPxwyWjMZLtdPDyxsCX8BVRT1xhJQ9MW/S
AjJykLWDbyTOA8UgYJ8p/pw0ZIvnF8Rcnc1mNwADNYuHE6VC+FwJp1+i9Qkosd02lg8nB7mG6nsR
i11ofWGdz9aRFPlyhVanHZCN/hy4GGW1wehmgM1A3+egsWU7TnlQwRBzzOQ/2yJRcaJWIPDMDu8B
fMzZTw3JyrTMbXoNLbT6n9ruwGv9xalVKeLPpXzhgf07MRTH96XfAyGiujGlwVr/oHDxkBf6WOLg
/PJ8UACmGX7bTMiEgdhMQTRvULScsGu+0CndDfilo6Re3lvEH4QS/EVOI/8AfpODkQ9sIgyJwFEt
SkQDoz0RFBjK21L3hkysZ8FQlyRnT5qEygHHXu3JamZ3O1N73/X/2bDubBThA4wytTMa4298H6a2
1QkmlKK3lIP4jvc59UgeZB6ksPMwyMuJUVuIP3ZRKGKp2c6HvIi8ZP3qy2PbvzH017qSmbA86c3a
Zw2wjYyvJ5a1t/7xQVGlVPrn0jWBbwecMC0JEQX0xM7ckLNxZCPRWggCLcYhRthaycEOuuvLWvzw
cJauEA2J0BSgI4GM25Bj+WX3x1apqU7DT13Cdf+Tb7RmNmsRO/U2GwlQ0hk79i7/wJgBybcoYQ5a
j/zrKtLF4+Yc9QcTnt0U3Y+inXL4pGneowko3Eo9lHPYy4KEMVeHv5VeJtcKJEUxSurnRgerYB5Y
ZK2YXHThftJMK1nUr/p75bEByOMUw6cHz5GJxDQEQFlURlREffaIt5dHZhYMkfUMz+5Nx/UupsU0
OzwdVszaOVqj1MzIKvkit4agTqvFpBVMkFVjmdwJvFQXLFNKT4COowuDrM/YNEbn7PgwbH9IxXo8
SXEwiEyoMMcFT9V7yGIIGcEIh+vZMPdkdOj47AEfxl4VRSGXq94uZZ+W4mi0JqZWRA+MNBj46DeU
v/k0HS0dOt+Vfss50wfXnkPwqcHPp8vpZurhPblaTXiW1uEGjK+ht9/YbdEScq2hiMFPrdN3h16A
EU66UOyj1tqnFiiFUcemgOTgyy9RTgTPg739x7npS7X84IPSh350RsBGMizO4Movf9L/rYTPn4ln
IeXudN/CvAeF89pbtRkDfel955EWnJtLYNBEr3Aeja0iyKqJJYpUTYcqIJULAvLTZcftQVKKJDOZ
+1ITS3Q1mvknCrg+FX7o7pFDapuGy0DYBW1mTdPK4aWTquqNxLWjPzVd6Qjv/lE/m/PjbReWjHKI
ekvvWKcu9DauZMJEHpFJrbINm7/ji0sW5GV+DS25ORFLbGB562R3VvMGROA871EBdrLsUt70jRte
mhzfecm4e4W4/I4qTIA4Ty1EOaDTck1w4nOyL0As/SJr0lMOvFrT537/+bvDGGbEQu9fvY/GSv72
SWAd8SOHzpgUUhkP+N063yWEU5mnPVOt4HTZd2HjQYvltEr4ghqsigXZMyqXrgWw+Ge30gGPFIhM
ZGSQocn+SnRGIG4uvz1Hfz9PyvIiALp+y8GCEZhkd3jlvGNdWQ+lYlrj+t6u0ZtaoyUQ0XMtiM1R
KsvuAoYQh4xrJtcOkaXxVH/aOFMNT04mN8qUgekWsdO3yE9FTdDASxbHvTSKqCipcI0r5hE+wpBF
K/Xiem25NOXPq8MppD4BsmALzY9tnyo2pdOPUr5tot5yo+YpiV7VfzJAHDOQemArBU5idw0MyB5e
Cd7y29rCQk6LmHXQwEo4CBdz0gEzDXDfi/7xA4qJBjbM+NW73pkAf5borK1DiWSz4ZclR8bG7xGL
PiCgUKvo00TK4qGpIcGtWmg9LFnz5kkUZfJ6nyCX7JA5taQQf5VqmGCcZRII/X+sEDJDeG0/9Za+
a1gOuFIQDHXhU8ePsXmiwT8h02nMuyrfqmgt8EJz9349z9IcfhI4jN1AKdLcF5EAiPKBR1MOqOSN
VR/WCg6ZExk8iCOnCnr96SQWbTlcy3FL5XejQF8xfp0rrtAcbSnHyQ2iw05YuxKPn5j00R+6/Xr4
c5gkCT64d0Z7OUNQ8Mryvl9nwjN60QBq5ZnPrKSOUto+RupHvPBus08z6JL5IaBViphaRh8Kjy3Z
6katJyYuJk6IpV5tQb0FFZlvKuYtvJCP8ykzEJWblSolpmFE7fo/WcLxehOiV2my6quXXPaCqCrN
QPPNTMC0lBshRnsFF6IE9UUOEvFNGbJQqImjhqV4RFFMiF8tuyS2mABi6YsGXRA4CUhokdWHomfJ
PQfXIUETrL3A/LaCne5jyDQ0qcLFj67BZlCJcchAnxTrBKTTZbV2Dvu987SsRBd5/Ilvnxy46G2R
dax1P9tI9M6GdO8veI+4OOVQWd3E4+GRS9iobVgIhVZhmfGFFp6kXiaEe96+iVxpGicE551OZpu1
xgnjdsTHhO6TowXpF8gI8BQNP+p5jU4ukAdZcjwYr9wt2q0ygAK21+MiYL2Ls1uJA1RCSfUcJeZk
1mqsEE0bBH629rH/j6yRPCPX20qsP8m6RNWSgldC0sva3hMc0ctaNgIrwT74pfKvrQf5HvehQpG2
qOwIQQ9iLy9oOXwzVro/AcF5OWoyhIkTIsCLN4kxTOF1BhGxtdRvAFfqAmwlHwc7/9DaK2NAxkyR
/MVMqeAyBLpItlIRk1SY3Y0UHESE+yg5uzBmeHX/HtmDbvYKW1bJ+JdqVoM9gbNA9PplP+hnEVv1
tXn9m1J2HH0mJYcHUaPwgSRCVFVS4n2hxG98FgtC4CPOCXHw1uW4TGd8tR8IAb7cF10ifuq5+1W5
KofHPmOANJwEZZ7eqUyyW+H5KwScs2jZPbUirxOOO/gSpnF6Y+eBTjviNmU4TK1gJKAZjd6lSMTl
ThGfqvYODp4fk99ErrzwEy+hCYAjrgf/yVAsf52sJDVr30IpOqCUntNAlow2TxibgCrtOMa3HGRe
fmpPErtMaPyM+RGi9U29AVojwuwLXXxRcv78aEXc4VBvgupzNJAvf14EqmWE3udVOKTgMit2Cync
09Sb0H0I1zVQFdipXfD3NTVxWvRvBR5nTab5Fa7pDSh9BEj0N6fSqUHleG2G2n0+5SJ/G5JIqrms
83ZiFWgT484yOQ4edx3m4Swk9vMZzTtoHasWeDRpn7XOkLClSwVc+FQ6jCueqXEyJjmQfLNaZDB+
aDL3x/z9TBW/w8ekl5XkkjczFdTTEnD9vjeRCPLyLwk/H0w/JWy8UVpWqt143sULiwu2xERPmw7e
xIuutzML4KOdNMn4omnxeZ0am0Cs9Nnqr3biAXSUdX6g96xGFwLCMY1yuk4Ca1eG9cyd2StaA2X4
9TBiUW0tlVYn0blnEiygjC2xdM52GXCbmPQAwRzLI1Bcn5QW9QQLlzFMAB00OM4RiRe80mJOjxVI
Je8MwE2Sg0Z0TGJ2qWdEoynBROIBKaSu291iyRqOilTR9Fk876CN1i0ptzBI0QQoiodsnOD2NIY+
JQ5z1gsTNwPIKhUu8haJYAovjyLwv2v1hVWv4KANaeWJCMyYQdOaGowShMW8I7i6x6plZBfPtNwu
/stKVQl2cHvXxX2W+0ABDV96QmL884pOiYpMjxcdm8cScG8/dPC8T57a2pyPpKU6xRosrmUuDj7S
jRkp72/b3SO6db7Rg01ZaZthWgVGhLgUBQwZWbD9KP6If4Q1iNNtZTMHiFUxowOC+Y2T9F/Ayltd
lzLBfIO80hvPBwchb7YVvC4f9abGWR6/ZSgmh8VrkejRyL4rh/kczSgSgfXqOA6R+8fx099WsJpo
8FoCFB6INxHf+yTVWhcUoe1OaSZ6vJhqtq/56R2gNZDxJ0ZgIQEKGMsCeFqpc6LyqNnuOhgngn/t
afqac10fG3oOyzvlgDiPs8SFLicpXWj456+SclIsOkwY0MiP4y6ONgf8tNABkV/oUvkoDsbYtgIZ
y9ycmc++oqE7XqhyGTz8BLfcssCU4GKbmueqHdyu2ojIVApbxQrZucLypAWaZNzkE3RLW5NIgma9
P5aUUkD2h7YpfzKL7YKeca33p8Q+qNlNqiWxgqtgj70d445gKhtocjBtSlZXbQgoWffrlnAMnwnh
1j8buEjbXE8LULPcXURgnc4mYa9mBPaqRx+rar91uP88X+lLrvc7reAa/6yKtIv2Zk8atYhVNxxM
5nANjnRv2w/Umjn3efaOrfgE28OQdo5Y46EST8iP8/3VM7IIGm01FwMxp0qyvF326CAXEpxy6DDk
V51CtUHCaHPrKIvWnWZHKfSygncHn27+jcbAmjfTnEM7UMKC5QyMugVqe6o78yt22LzZ+c5vpAHB
NPytouHSWOdrRZRk7CoRojCu5bMAsGo9/CTmkCg5WyUOgOCPtuBCNG4kGSoQ8jyOGMv1sL1zQLcS
57aO3tOwZG7C5ecDnAmf2rvYYTEF7eoQ+kehkN4aRoxQKD4oognLnLv4XoFi2PrxtD79XcY0MhXf
jRihgn8TiuJDM/iMD82fzXFgJTOPsIt0D2NUKBLW/GFYeOdh+oSl1pUc6ka2uyoI9hRDmHHZqq+C
nz+cwVEOV+6P95aFCcB8JCL/B0ErEvZ76cPjgsInFdpe5eyLU3ewYcISad1x6W+fCHz2RHR0PiLB
UU/BAQtmZfxNJjBi9t5ioyHtMDtttcvOEMBxplhAmWJm5lf6PlKhvUvd7besqV5lvaY1X/IAV3cl
CwUCZ/7OMCPVaZytiSMG9Ynmx34W+WCTdi0NsfLFD+UAWn6W1LlKF0KkxJh5SCuYPCQUXhmEpAiJ
SNZPkwDuR4w53UlCEzLjfz/QzONmBIBvGJMfJENLMJpBjvoFY1omRO5oQa6jMnick9hnhMPPicxg
Se28zQOEBuNo7YS6vGzk6GfaG7ipZYk0sSuw7UdeouA94U/TWlM40Iqosamv9RjDv4mEJOBxA81N
FcRYdR1hT7Mbj/iLtMw3ItWpwLyc3GBttVzzNp1P1MiPrDjZs7Oz+owQWPPwrFZu4VdQ3UJsW6kY
7Vb38wSbVCPZSSfQy5409yFlX71rCP9k9KPrXIrYmZuG7VZQT1qydycn9xMroT0WhQ1JhaZ7zcBF
aAgZkSZ444ghz2ZHodIcSoLIB/gIPIlKDHYULj51WVXhk+bjX3PPYZ61WCt4fIilajnP2xdjUS29
8XrtGMiOkFXGIwXUFyG+oNmB8ja2whK4qB6ZSArQP9RBna77lqrlIDLLExI5U3SJinPtdsw0/g9D
HXw/S1hdTqYkQrShQoOo/cBAc4vhqwQ+TYhh2rR4aX/cH5FR8kjDgcNVVCjSUuviDJNHINy5r8MC
NDG8M9q2LJxhc7cQzZdqqS3tnn+IYkbAXWWdz3P10Bu9XIYIUXnJmSIBMfxMCZ2CHz/aS4FtKuW+
ZWP5+H5tWy3s9co3uHA5s9eFNHpoHDIxwsgUKmcw0Ii31z0x/8smUeh2y3vsFL1ZWdcUcu3n2n5d
y9yW5gwztFYQdaED8b+byojYPDaclvWjNWJ+Hc+s1dhFX6DBUzZS4i1kd9wlr2tYcw+42cKvPA9b
R8rMGfxuK1Wex9LCvKuJFGzY6iZqOhGNQULiA3n9CfIZyKtDp4mIkWPSA31kIVjCAPYzAiwDn91U
nebS/Yt6th654e5GCPE17uP7X6rU6kJ7zunRw4+sqTuztD+xvuBM39TPm8LjAqYWVoVSf8AHJopg
zkuFjcwNU1s8wyh3G/dnt0ogGsv+E4lxD7rws09hfOFTng9iSRTyAzjkthYYFcw5bQcyrPSVIq5l
Bl2Q552F03b5tiAk9ERUi57PFaMUVdkIgZ7R9b8yuhJ7ZoVNlpVd8b0ftEW4B/xWNelxUUkzOJwQ
/wSx/9HT83+605wf+TJHDdZwIKLcXrU1iXL0cqYqUehpU3/So0L2R2ct0Apdwe2LoRyoB8JWAh7Y
ZCLqztLNRHsXJdzZKRzKjG5CF1XPjBRSXdVo7ZJpz40yZCtycChyzVKvJAKKYrCn1jOW/Z+WMBA+
8WIDE1LQswYakAB1DUPLJoDOdNLdI9iWX4Quh6v8q9bmX+RnVu/19ZFQE0QKwQz3peftVYBNeaAI
txLyME/iwvQ8byjf+DD2/yk6On9SCDUryaWzPnMDH5MsMiIBMiPQzp8eNvunqFb2M+g3Mb/3WfpZ
6aUpJlBoNNaaBnBWufr4Rvxl8im0/FYbmh4qZNqB6ngDhGbOMU4cwYoEB+ymC4b9j0yST48ShhdW
bFixp7mXMkxAruyJp0Xj3+2jR3BNMr2vekONXpOQ6qbtN2olDIBabFXk2rbcdN4BUmvr1smLQg6V
iu57qypMgmTUc7T3UNSQrMPLwjhLhBgxo2S09ZJ5HmRcNeAe5dCP2KidZi/U3LkbIja8siUkyyTD
i0tzqFKe3IIi5eZkwsLERNP/pCiHcnADVgcHo9JYbYejGPDR6zh9oQadkd9K55htg0N+z2WYSruo
oPuV+CDIH8At6LqZp2qWm3Rr6SmBg5+mM7LavweO6LYvDI6pRaPwcsM/R/4WXQaxwCYE5VZPGPG1
V9J8zQURWt4tvTfv+7ufxxSwNZ7s9FxzBu6mdWIZEYm/WOxZxRUjoIrAix+hTsogPRGzozb5zbEU
tQdmBexHqv4UO91R57zwMQ/oSeqjx1hHj7C8DkucdTI6vE0lY21d9iByL0ianESTnIfU/dNVzQ/u
gnNWc0rr+6vjX1jZswA9a0yx3LF1xMXliACvX/rrWqIBzh/i+B+Rwxsu0F6rZ5rmwi24z2EE8CY6
JGfaYUnzWo3B8DOd+R6tRGSMvA2485KwSsDdvePIU/D/P8wKEmEFF50qchHprjgFtSKz2G4fXFQM
IadrFX7YHOUaYNKEGv3ykxW0NECbIdVGs9etB56Gey3Lz24PnHJ7YgUTSkIjbyiMJT3/+rrMFx6B
uzIxW7vrmK0Ccf6Dhkie2BS+1T8Oqjg3ibZIWk4tQwtFkTsq82z6zQB2NQOGpvDMTK62VT1hEhvc
zwxcKue5T/FV/rf+/HJhg2xuXM+pKYoGLC/VX08uqxGdh0gBD8E7MmhCTQBw0s1h2NbYHt3kuyTl
nBb6wY/6G+yO9tUbF0VCYtl72xAo1BLXmAAgLfw/L4l4tejgUvgnszP8mnTS5IkzTHIQQ1mSFY2i
27F0WyYOIetWRRADE+AMrPQNUANzc8VUvvD5bMPNKHxNLlJjeQTjXA0jwN2wwCld4oRRtPkg9dBt
/Mpc3g3/1MsJPJb8sFzXFmGqUIhqCQiJ1VRjb0D463wd25SHiBDtvY3Q1hDCRC0fUAUlQiQQt05/
Q1YuUIaJt3izmLtCn8A+eTFKMV3+P3kEOmR4f9PJnCEuhZafbfFmfm2FiZR7S77ZvXp6X6J0NilT
4/vxeox7TFHCCMjh3IoHq0/dBv1HkOeS/ZaV0cR15xpzlXEWpTISlPK60lAKRNUZaJxA1F/ParBL
yEWeBVIV1T+kut19AawPNo60yp6yztfwCUMrYUXRyQwUfAg4/h49nFjc/WJh32IcQfd/VLikI1Eb
HnPFvEyLAi/6oiFUh65r/EWuTvyzqpu3LhSudzH4nO8ErOkjs8j5Pw5Y1EbRExLYrUbWFFzyHZFk
OxCCG8uPujVo/+oagnioPYvaaEVRFjGxLST7vBx2kmx/y0NXAxnSspIuI6LWtWkk6XVhD6X+I+0i
7tGPlFXz775ubp0DqZIQvULOWToOo+AdBbvKVpGn7TogsQ2HWPvxDMPUcON6Yn5kZrLl6IMmPJ1f
Ob0O4BA9e0DPcOrilp0eXGtLho7lqQgN/yzT8ItRHsh4vvBMZLYbA8X/fM+awXVQNHhkOSxxR47z
Sy5QGHaqkbr15Rqhzxb5XKHZ7jlzpMtggWrjIkqXL0TNYl6U25HrgYkqsUaAX7IFZHeyuawhLddn
3SqTTe9UNg2PE+yyiqhI5Sc8fMpph3E5RL3uQjVzzP4tcFFa88GgfPlsmfd6sKAquAmm/iWd08Ip
kdCcrn0fjCKrcYPrsVXYZV0BA1QzykOVnSCsnx7rbiaJyufzfU6CySygr8B4bdP7rRoPmUQ7h7fq
83e6YlfVAocYxOyQlhjGNls+JoARmHVdGoZ6ggskThiaIaFMeLmj0/KGWURrJq9XAwuBWv1Sxhqd
0lYJDOBgdEBdXGqaApFqxX3qZt6+HMVY50/pJl3aJhGbSjgUJVIUIvbOu7Si//96MtHfDu689pCo
0OCAyYbqXC9G1Ot2F+DhNzKrQmCjrWcSvAtr+/39YjrfaWyn1xFAXylMHKOJ2IRWsWG+JBc7XoRZ
ItIs/scaUvi4s5oGg46CEt5/HuiC0HHAOCmEMeO/6QlS5plYo2yGkKN6/O1Q4ov4MmwNVDnr9p+j
jF+GnjG6lrIuN43fKGFFjmoxZ5dbhvVvq5S2NkWSbYQHLXQT/Cpmm9Usx1V+NKA6YXGly2Z9C0pl
nMtZ+kdQ8SdPSNDy32gDLIl08/mMHyRVlPjSwx0mHo4IFmRae78f2hBJvLSawzJ4RAHEvLIMVQ19
VMdRRxo8b2r1FMF9t3KTrN1x9gZ5ycuphoaslrysnFEKyzP5g2Alu8kq95DUzSWncoamiINjvdFq
ebRtpdgUHddlE+m3tlUhApwRMNxxHPHlMYCx9ieQE0o1xNEg/nkAeRwHIxjuoDjHZkUAvwGbQJHY
9inV+bRkzpXhsWATmv3In0NfSi0zYaC2+dt3TGjEuECtLXkrsRx6lc9ILTuCi4WXPCd9zZ1YB/Fw
AQvvFTmx+u7eN0jUxac9SxTDRD8nafws81scBAouPaaAmr8kY4hrvcXp6RwhaWugibd2VhfSZT+F
WcL2Q1UU6awIesxGsq50fXCBlXPH0gkhf0xwGu46QV+41XSnBA3VHVGB5PEmMjjVj3r1TSY4Zwdy
RtBdtebFAumqxSJvJ29cjteBdE3NlMQV7/8CICszHHlRoGdmxvj7ReK5NdOr2oMNUlPq2v84g0Yx
ImYgcSIKoFGpz0FHN7t1mLMs8AnnXJm50Rwm+KxAnxzxCp6yLUYkB2b58cXhgQqLuiVzJvIsawdp
WnRw42Q8oqqpVtVv0V7QyEOzrrZ6CInMT6lsBng/7VkqQyKXO2BwbptzU2bhMWqFoANJMAPbm2KR
OEfycKDB0PbAt0jr9V6IXAvYIT4EYi6xlmQiUJh27vxGeshsn0sqBDyoYFYpMVU19HWKvT4vRuss
lkn4pX8/iyfO8izFJ+DLre9XfnoAoV1sJb869kW+GJ7+jqzGNHwVYNmSRmfd/XTyxv4/dfGaM2FD
CcIEGtUsBsmUmbOngUz7+lD3K2xsg6hnS4f+gaMAibCuMBzhT/pB9ZNua/NvsEN5C9CRBZ3TsZQC
emB/escwNNTzdCzkA3U+dTxPB/LmpwvMTw1Q56ETAbhvzxgmXBhTAYHgfxNvlvwnJcbpAsqeQfSs
DoM+d1SROQxnw1mLJUDDkTGoDNyfYZxlLv30xfnH342wxtf4Mr3SpNm1bhVfmXMJgUGVh/yuWCtF
s7Ea+moih57YK8soYBvfVpAgYjVyJUsrrwQbxOM3nVwnyCVS/5ZtLMy6hDNf+N62CahoSfYsTLei
MSF9t1d7eALTqaA8cvrFGqWMbOYoMyObqV7UKMKvoSsPH04tBiuS+2eticuE12Y9sPZPA/6GxKG7
n+wOSkVZzKdo72bE/TpRILOAF2eQEdro5coF3hHRdyTkCnylZUkv76LZ/5JsPM4AXU2E8RYllo2m
mzN8CQ5Ao1uT5ndeXuyq4eokzTpeOvbZvibFfoEph20Ye5tzOeTA34SbeWZMVycOky9RNJaB5zVe
eaKeoGQrb2jg2/00kfrGoYN9yXXD9YGqC/gFvLSwpk/Qcf+dre0rpnyzRK1DjdCNYG7JWzvIew6F
kSvmB38XQkWkEE8fUdyj9NmEB9eY0bY+sUE5ftUWxlAUoDpPL3jLN6sXdlLm7082GRuuZzu8iBeb
a7+XQWB6uvc59g0IryJQ24GE1kSqHHOZwAHqJ5ENxKeLHtwChyQwFi4z0+rFnTDSI02tavdF89vo
bMAQgImyTruPowFMT48Rh0Wo3mJ8TRTaje/qMdUbSrRJFdpnVzYXNWOQUMWFUCjK+sj5iXLAn2LJ
iD0NpBbSQdOnCaKzm0FXuDNzptYAobq3ZD1pV8C2IFlqYEwmcz3lNwbsLksIJHinU95lG3Skwsjh
g5M+EUnWeL5QLjTRtUTGa8ifiVoGNRo77G/eb/njb5vF/TkSNf9bY1oz+djfa5w4A4vNivr1x/Yh
kRnx3Xe7H1Gl0Rybrfg8I/lM+RHKTbmD4vBJAWKvFFlZ/ZkqWTbGovX3rObB6uFGbdofZEGHZqx4
8ywyC2+83LWN1PI6gfdkYoBQBLtFENRSIWmQWYKwV38e856/Kf6ZRVca0zdbVwsfnFU8JM321beo
g2uwrFgj32gaDaMiFXcZG4V3wAqLAIqxIkx2qa2pHcBnY/zWW+bWypw86U1G2SaGhtxxEOBuoEmo
OCUyNLQiUT+9ae1QBWSCPhqkZ4PLsfK6NCZ5Ux2fFgTLxdnwdCey+C74pNerPp47CUCon2ctRmLJ
qfSfqaEq7XtvuE3rTrB+Z1QGhrNQzC4iGsuEBrHb9fq4QSpS9UIPodJh8/A5MFH8G+ERHf/Jw44Y
OidA4SGJgAHsUlfNb4rRW9J6jMpdHu79PWfYJsTSpjkm5GJxTg1NKRM19KGf6oPly2O5h1N8eRp6
uOgufC7x2gt+3tlef/K01qJFtMVXSgxMPapBu+YKZ40/gB29dbM2q/YbefyeN2d0ZoI+GmNMBayF
9pY1oy/jJey8SSXueFoETam5B+wE170lGCvZikBckGNQV9LZH0wnuWkrkENVdc0lxOkBd00hw4j5
EBmxOO11b4c+lzRIvn+mdhPbY+YVQA5Z0OBIhYXGJ1kgqMxoloxowqKHfyB9Gsm5a6AtNgW0slDP
TFcuWv+NfX9VPXgV0YX8Z7KufT47tKET6nvulwBLFVu6Mcjb3awoK5utaAnw3hZQy/r2XmrWokhI
D9Ik63VRUgenuMix4aX5h5OMxHwcEnnb5BUnvTGygChqTW2S6bMgd+yGRUDkCEgONrHFVf0RR+XE
tRA6jMINzEN9UqmFW5MkuXxr/edaDStGAQWdd4eM9vHfUBX5++c1ugbbP3pjvclarA4FY75aXk39
rydVpq60hVgHvyrnMM9bPF0R199XPh9nMkhrR8CaWfX1P5x2Fl+NJXqmngYT2y9yMzdyU+327b9O
QkXjqjuCTFaAAev0WXjyWREtuYCl34TgfGJXywOcGrCkrFlpVtTIj3NNtI0GoUjNP8P8qspo+QXW
JixBWVWkfshUlYvy7VOIP1ZhaIdqSzzVyBFag7P4/rI8ugG4eyZYHWm39pT/YBnlfLbnJVSClpyL
asn+mkUCFyeWWq7dko0UJWEMNS+v/Yt+fy+NJJhHeeFvG+1L1FdkSwe8ghMyE7AL82XT++pB/ZNz
Cg5dZUo/lMWTowrFK8Qx8MVeqI1uXiTCFwFDIfqIH1r/fwb+/4+EVH3QIErLr9fbIcwlE52ZEnq0
FNl/Dw9zS4r1z/8EbioHE4vyvCRoG4ebx88Ormgya5oNkG/EMiFpnFiyZd8NdypRPCI3T2he7SMQ
lpCEzWOsZ1UQpVOM0pyDiFXZrxcSnc1HWvy8R5kSLepY8Pv7XyZ3n1iOyV5PFJBdkLZYOsWMEZDf
sQt+FmFa4qpjv75ntGn6XsJkkkB1QVgdlBokpYkNCU+zNZ0+dSXEDFd9IUzmHmEmA8W0yJgWFX9O
UpLrVLiIl7WmmCRtOpctm9Kog7+C+2Tv97DtuI0ZgnWP9lMtf1rbT3qBECHvYtN3ydEdbo1RXDlq
rJJUg/0j5FClTrF5Z1WtFgWL+BJVePQo0SS1Ph7zpOfIy8QD7+nXQ1eXOP08L2dT2fsC8MXlx87l
zzCT1M93rSES+LQdGQNvC53G3CaHecsx+fzLNLTgnwUqzO4QGVs1xto4ta0bR+13tWKiYI1mm3NU
CzEhwGS/1osNLH/GSdW2RB6HvEXvjxLEfpYH+GX+2Mi9Z+kdfJK1nOUhp9TNYfAIunoLre47hvg0
aambHEQ5DA96Miha0isr/A6SXPLQHzfRrfkzYOYDoU/Dpg9UdvOD585dKb5nT5S0rmQdUGWm5ZN2
2GWkHzrqiCUrPcuQD/Rozq8VLZ4CGArav3EAHXznCitq6YuOR3JDF4ZGW2X/lB3qXbJ4Rm3Ide5A
jrCQ+G6sXkro3oFVzWRTo+2EFj7FkdCg++Ms52CeXUwWLuND9dSN7SdCFdpFrR9r6czvgOfYLTf+
i/oAdlAnVNZYXjEYKKvSyl2C6Uan0JcsZ0bM4Xugjt2GTEAXec8ykFcnXTf1GUfVyCsnEaH7IbN2
2ioHfNVnrV7Vhd9D17NtVtPnZOEo1j0OiAKQDHrH02rJxo1SPkl3wmJK1jhgGm66OVbv5XlJ7HGb
evR4ERHDikK28ooSid5jqv1vZoOxTwSrbb81stqrwu089C/kqtKklSyDtNApf15JyFVK1nllPMOQ
sH2gDACiufh54XzxLFELIWk/joNNsTc0PWlBMSZMrtMzkrm5pADZYYHW3b88u7ib5zbPnYSpFdoY
APg3dVc8d6nim4LFr3lxrXn7+ldTlFtMdIEfQf9Ymlsp1ECcWM1MvSgk+onATBjcw59vKeWc9r70
W05oxrJcbahn5Po57e4wsA9QoKkDZvAbIJNeknv/rFNs3iRpo+EY/HovHEG9oWYroUtkBxjxlZbA
wHYNgRYyGQjv9YbtOnK7SwLa5DY9qEYkqS8LkeVZ/ufKa+ElsDHzW54m7DPthhC+6pho01J+Lqsx
j4W0iN0Z5ySbbPYQM3cRyLE9PobD1iUP1MSAG5d+uMQYyHerTOfUoHpUSlZN1o/rYbpHF1WF6WiE
THiC9vcbKQ93ULJ+CHVLe2KMq2Tjlul0/rKrwB9l8Ynj4ZhQAZfMdTpRMs/s4cCqXReJ8sfcx9Wc
jBk2EOI5OqmGuWnNApG9Uq/JTGqD9eg9eSw3K9Qv3IqBFBOydi1RZvhkZwHojpK2RJCDE0arqlZV
prNhKmjoOC9hA+aAaXhtEuX9IgF0amSDItXSmS4OFWTw7Nv8R2Q6B9AuVAiTTba/Srcml4ForXnj
Qv4CIkHSebRIxsVMBOfi5oPQ7awsDxxMo3ITImBLro3hNdcBroEqqhlSZ91Snylc/kA422sh5n6i
CW8gjCOePNPfD2l9Ga5pSe/0ykhh4SIFMd4O4l5Xiyl2hWdktVrR71wOD9SYZs24E4G+krBxVlXJ
pJCrb3XugtMOhYSV9xjxznTfxfCeVnTrloDQYM7gIAcPC8QNex1G9+BfFKV+YLZe3YaPNtoCBi9p
NapOw2yWrr8blNSwozwCWDcBkZf0yGHocWw/oJB2jbhnC9yEzBGHZyKzHcsWZvy0dLG2lRSQiRtn
GDK11RAyKBEWMp5zboGxnqfJFQMC99+76UBh+7Ut0MsFuzN75U8P7XgBWcJ26x9pSdeVvDN6NFBF
EWYpzFcv8Ov+b0bzW04W50tn3nWaZFTecXIt1Sd7PQpRZStGHCOEJM7sOnSHeXHJIcJsoujFE2a2
sG2v6d1e5NMGsXWhfmDrrkBWnYPyhbm7r/qFWi/Fca2yxz+ktXGu8O+cZ5RGYcXXfb2y5axRMd+8
MlxPGNV1BZUIjZWNmP22vxUifWLRaErQc1CCHzNV/chnVfi6qMU7cjUkLhUbin+j9npUl//cmfzW
1rq+wyPVXqA+vtzMDkUEDTX9myKPB9uUgdygh0aLZsTwqRjAClCjojeS+5lgU36Y7UV2aU6OIYY4
jQWJBsmq0dqK7mjMIzhmYkQF1uITyiC2iSyldgXXcg6zVgyETAWAXHYCw28RKO+jD5MdPt9ALXK+
4Vt9lLrd3CJJpeT4XvJEccWMdRafELhTAlsPyWP7Id3NoEbj1zSlb3aT0ZVHUR2iP0e8r4wNG2yL
goeU9XC58rSPAohnbI2P82NS7gGHLscCA8lfD9nBowfDQZk5irAJ6E9+VkqFN/wKXLDkfg9xyKWH
jGyz8lTdarjFpOTOJQrabkbX7e5S9HXMX8/ZbvAPbWspQI1ykvDnQNNoFj79gz060wk45ansx3Xi
b47FUmPAbz88m71rABX8ke9NY4mWt4YLPB9qMcZDhCPmZ7sBUmEIcIBtv0CDkXK0Mh4Dc2OatToP
brE2Wyd/bUEMeSUB4bG3PisTR6K5Va3Bb5SdTJGlT+sJidr7AUBCS6M3mS1rM11l5Z/11Ds12axh
SVZt5ZtucRtZzZGxU9JpW1p12oPVbbnIP0L/he2sr9ht6/XsnKz+rBHiPCNpw75MeZXKMxrgSN97
0DP23w86ukw/AKqKVaMKR+81sQp590zZVtvSPTKpJBlApHCKhUt1EHhle5IIaq/VENAIYc3Nd/9a
JWbjur/htusK6Wv15gWorj3TlwCxPm6h8QHCFsNyVDiOcDcEBtUPH17+6pNHfR2mgVH4RYscJX9G
eczOBpTXzm66IgDUFVgcx8Jh5DHNR77C4xkDlbx9d9ZLdfM0UgNJxaulTOJnPhXf5bRgI9zcbnEF
zER0fQG8/r/0p9AQ9i0K3KTxO9/QLObeYhfZ9KdFUbMEmQODC/7+f9fcvh/MBjZ7urKOvvn/vmXC
9wbf+JQf303+JD22kx/dl3Duwx5ZjOdppko4QgsMW0COn9o8VDuvaxniiYzSMr8zcOyo110DGzo0
VeVgpIU38h7CvjLvhlAIobMeAsOwI+wRr4FSmdlpQauF84EhOukfTN1QkR9Cp8HSG7E6ZyX8mFGo
KKRlYgjDc1vRWmq5fJr7n9By1PU8cnQmSMuQ4nD/MXsBR/HEEDsJC/I6kKWNR23ZP71mPI92YjXI
wlcp54VmgyXw8RU/XUedzqxlJnZsbJGntm9SkePBzAh38oEF1S/wtN3lFOAYV0gIznNm9DXpzzbR
FQJ9yDQTsJXH5E4YdarD7RHot0KmWhmAoQcvSKhoiSTZzXbUH8Te4y92SttaVAOm4NX0W0QkqYVJ
tZ/Po8o7bx/c+gP52SGXVikyG/Gt8o/xbdVM690bKEZcO8swsxXSUEcjXVeJhnSRCMHZJRQGClQ3
DvkWx7/i1B2M0OVZQTFPJnSpFuYJaPYcaitvBVXMLG6iWzvk7Az7ogb9U2hICeLTJvQXvSG5YgCo
1wgvjqhNNJBQgLVl24bMeo/b/UNL55mvBVG61bUG7B3FRi6EpiKOaGbc59FEPqpcAFuFMtGeKgvd
f9FtpILuSSVSAYfAJIwG9RMR5rU9tAYeZP3Z4hGNC33r8BA1UgVjJ/hjh1rBDRQ0itfghIdszrge
9jbvNHc6DWJFgKWQN9HOHCxsPu6YTrCH3CYEU2CPCPkAwdFInH2KmaHclNOonT9blqqZ8QEiz0BJ
DJEXtFKcrrCa85T4XI+NWvaBr6HbdMlIAcn6AdFiM01ye2uBmnYJii9PdVxrIwCo8g8A5HVo4rPf
n+NiLOM/VPk974GslNqoyQK4nPWX9/KNaYFytmqL+wxdcGF2NyHwvPrZ0VQ5fgEYv54jgcBpoExP
5Hqq7Ge9gr4k5pBAfx6oeUwHTgrl7BB2RARTniOvbwVOmKzukUSVonwpvXqBGeN/vAdnXFWVM/7B
n8CHmB5qF2T/H1dv9o/9X2MvjKEKbbtmrzgc393Oa2Kkd3/zGpU/RTV0bOEm7u1/KbNbwq/DB5Rw
H6RdpwpLflSxbSo98Dp062JKWn12pNBJOfx6T67uuojEMn8QLTufypRMhS3rJ93+Ber9HuhM0Df8
WkZwhK5w5OLhvq+rQ6CDWUoTTdIa2I7R4de+o4zH62/YN+NiFP8t+l19bUgNlScPKIaX+NiRIjqH
xdwGAM2i6MiDFpBFjZ4hJj+vKppehT7jvfGXQVZmssHJi9d8gCYIq4nqhMucl3/nB7Ztdk2Fc6Gh
wXCnQthnQu2shuU5z2aw+CnF7lpH0YEbw+fNLZY8LkRjBR0u/W0qiOMe0rXCt801KgCdI+T+CK+T
CVuETbeq46aPxWysbjCkAJr737CxajsqO4E0XWVu6op+8dinrLG74VFhBLdAjAwTYGQhkzwvpgw3
OPQKCacu+0JcRiEu3fDzc1zri354x2FAqQONc0bK/bHyiu2yHrKaKnjJ3K77YL0H5lIG3r0n+YAv
1HdpXWSdT+LDeA01YIK5hlNUra8jIzwrhtJNl9dTguipuWzlFDuo2vPZiPsoliIGp7kwJ7E5HXH2
JS88/7o8/MAFHVYu/PVgNNv45+qAawktyyU/YZK73+0CYQKDtYDFRFbB9ZtLh+xqCc8/GEJiROAW
lwGf4YAb7nCZIH8NxpjbrAMNkVWQasBwTHBxQjVuFzq/zv4GZUYwc4WeMJrRGhVFxV9hMhsMtsic
hVgn60aEMf3KvuF6bPR84mGRymdl2/97gTDint6BwqY46PaddKyBNKH23CPwQ35SVynhoel7j4tC
43cLyZ8/3kbj3K2QW2uin5Gl6otf1Cvo9ZMEXTU2t/EDFQ3lY/WGNnB1EGZut14slfy9FM4sL3ES
99SYlWQRqhQ3Wa48zkmkZbRBBTOo/J7XizCIzyJXX9Kx/cXvLSKMYfCOIHz1d8Drf9WcTpzRMGAX
L1yCo7so/y40I4jPQmxZdSpUxOLoBPhWkpozIDsXaLj75YOk68DQhpjCd6wl/3TU20Zpn0mpwWwx
y2iAHOryfdUkzN1/gCh05eJuNB0B//Fjc3drzdAztrbzRrBccm+lWhkAOyW0f0HDARM/sCOtHWp3
WSYgR5uw+30o1/EdX7PFjkBbexJYrhOuPWo9djNRimAEBwgcRIXiXl9h/K+v3j+rZOULNzOfDu7l
PqIobGWiZNJJm0dzd5MMjV104ylLC3Ovw+1W3bBVtug1SfKNPgygwtTjUwcM/uU94vT9XmzIxKAi
QfdI3cJw4mN5TyJKx/1NU0rft2fPqkDWRcqxnWau3w4x57Baz4kHyYRqTM0GqYZg8lC87VUwlS7d
6D/8nXQFwMjy/fdz+GI2zjm3hyPo0pwyoVP9GotNSQf5SgTS7jR6Z6c2ME/qPbxvJbBny/21qTEo
w1qeESbno6cdHCwI3tDqt9/9Fn2NYG6ndQVnO70pr4W5LxgbUrWJ88rtScyZANoMLdqOckxYNC9e
/zYRRhyHaAdTYMsyMr6rl4gymIvQWPTBZxhc1V2d17y8ke2IWrvIO8GIKZvOW6OuPxc5PiHorC6o
TFWu/7BtoGoRpEdhWzfpA+/kNNXxVycCuoXhzE/B1+nUNK5J16KEJXqPCdlmnfCaJVFtiu4nQf+W
cgolXnpoFHz+Sq6tocejcb1FET0acex1MT+DykYQcWGr+y3FlC6U0208hsPEvsZwyKfekEwHy+Q4
WJSeH3qoHzQJdR2WvM0+T9Ao+9Q6bY27dVNYcsf8Fgt2ePIVwUd21rijeIMTllkq1OMJT2jiTHEz
S/qQTKGZq6Ii7hmGKWGCRj/3XbWaN93RqGWH7mx5FQxqDbe3xMK76vaBd5reirksvA7obdL6ePme
gSAXHoLYZOeMvjkEGZOKIIvQ890fNYLEITE7+TQvp5o3Cr7YBiisGKxWc1JlBGIyBZCNZNgN+d/Q
gVHZC5ie5ReYBzjelARVJmP6GS7v/iSlBL7Ckp6xvMT+yL9ktqaeqyWlILpkHVMRKGgUrP8opT2P
rYel32UGj/AZLod6Ww+Z0how1lVoFkoB24YnJ5+uyTc4d4p5/r7Uj3Rh0K0uMLsr/RJ0ddSMxXI0
G4jYfgQzXo39zevedG/+fJXTc8S+YPuXCn8cIH5Lm1OzrhnEn03cjoHUrUVMPx3VoSlmcXxSMFK6
INJt65kFwazgDG1Ph8ayfa1k06Axrmq3l+ZHiQ+R53j9KZB2Usy19bNF0vAARf2WuPJYlbFu1Bm4
mr3oEeauLFRpHM94KdOCT6iCZvn3qu5eRj+AqhJ6ifFovlGeItMrokiwEXTbxKG3WgwMkWvv+4Nc
S9ZGC5HUi+JiAIH5W94EA8v2DqRshFUYgMSK160CVd/chbnW3/wkl8VUH1a7tL9P6Et4fpm+hdfi
/EgC1V2UeYMz+Sb/EGXVa4JQfP/j2m7Eba1x6Rs774cmgV1G+rshBMnOJLidv4TMadrqSULdXQJr
sgzlR/ZVRBO1rWERXBwQBI4BIdmRdZ1v59P1sjE7QfoD8dpr7NwXC02RWD/mzt0LnfY9Ffj/up2m
E9e9vq/JfxBxMRcOcdBWy00WO7K8joH3hQwEmRVAhVNfU6lQZjAHhVj2yf19WlX53KHTt6bzFXv2
TlJd1+IkkskOD0XxmZxqppN1JKXQPyGHWmZYEC8ijAef87MM/kIgDWoAOEzTo4r7JdEqQcCuv60q
DS6ZLJZNu4RJSypq4WPFR4bCy0bdBMrhI9ch+J73qRNvQqTSqFBsoPCWNk59/nkjbpTeu3kTScqJ
2lMsqDPWFywJytEkqx8H5QHr/HGioCS+9c9Hxoxkp+TTo3n1szRXQzJ45mDYvDu6wamVdCJUx55M
5iHFaaxd0fBvnh+G2qQcwLagu+/tX2fOWw9atXR1cmaz8z+lvOOgViKZ7GB20f5V4rf3aoA4C1zq
fNm9RyI/Aa7Ddr+EU9Y6FGlHInCQuCK5Id02NO2hWQADi9Tz0XRXRopC4pt+McdOnC7z9vX/aA4M
PoQP6ceV97A7Mry08xZdVmesi5ZrSKqZkuxjd/P3g63pn/gjhu7K4ToNy5vTXmRMEwxCmKV6axPH
aanI3Xibdbf63FYomuVpoctkmOoIr4ZioZ4uN21CmSyNBMjKrX9hlhmcayzYedcnMfa85tYQ2aJk
MSJUIM0+kzEyPoXunMQl5NWOoi7egV2rVtdGVMxvdK6+OS+l4RdMHQGu4QGuZ20QD1nc9/C0ex4d
rJAtz6gwNZ7IViJ7bU/wuGpZowAgDMoQNaJ7EyKLMDhYqdDNbQncOIqbS3Tlo+re4m7W2cixnBAa
uKH3R1BOWv3TdPuGKwhtmDWFhbsnh/0UMq0cj6e4XSFQj0Cd9qBnCZ9fXAE/D8NbzTPXX1mjsRp6
3P+mZmE5AxsqRKGN6ceFZQbVF/cHRLGHDLEO+VcZ7U3rt6Z5QpdcSHQ2nGR//E/qZcCYXBBwZyDa
HUCv24r1tSLuySy7E89ilLKKUJEW3PbjK1Nbx5gazyXPb/JJRYEMToxOpJsiOwBJUQNxvIlcP9Bx
3UwOEVYCn3H5zjBg2K7e1c9Jxfhd93icAxLMNCrU31Z0gBZ9w7qRtJHZfUFQ18g9ss/eFD1eK4vr
cdC+FXNiQcyGht3qhkyA6ezL/JdtvatSbu5HBwe9iApObsN/Hk24eZs4yvoyCYpf9BXWkWLsYquu
i88hEZQCinZD0t2rgbLg7sZvsWdglTj9PX706iUtFkF1U2tTrprbbZ7RA8qMJUNciEX/MNAL7DaL
IoyMm33Awe/q2lxIV12mlWaIUFKOB/JuFcspDn7JbQYBnpngOxXI0CYv78bfOIY0POfCI8VP5y4j
SnsRtB57coyYFKu6Bb5EMtiHn8CfkAy+hu9utIFMxNPX745c+aKsCS7WJh2PD5fy9FEs7EyL58M5
gtfXNS599ueHBUSLnkDEWuynTNrtpfxn6qY/V3K1P7ZxGSsWoKMmmoaE3PATjnAmePnWkxf//2iw
eDOXGRzMm60BCdyCSZ9oYxAFTxLCrvOaK4VYWYopWOB2SvltASSrebYAIXkn5r8JcQU2Ce47eZrV
NS4Zi34yHVHEp26kMk679dCaCfw8dwGuyknHRHAKg9k+YXCSxaHhe3sKJLPs5SSsAXkdVBOUZuOG
tOq6G6Vf1oV9pU/rEVYQI/jsN/9s2iAX8wYDcEY0FoPbCjZpMrpO6q57BCgFeYRk8YTaSIzQ0bas
/ngJYqXM5sJQpeZFf52VXLRBe4os/E1heZ1p7v0/DSzvz49i+s0e2qmkSOY/PFh5WqPyhztjym2b
FzTNM8KwNiVkLf78vF7VLoBjiY36x8WVcfKaZRvL95cHgbfc4NWGcNc0p7TVSO5xe/sbWUFm++/3
N/ovcx07orJsMBB/oIZyeRubcpYXuaB2S1CCuuaLrIBnUK/9kquzSOux4/ZKs5rxxipWUCVNw114
id3F+mrNk0hHeW3w3ntFtCwg5pyXrCWTb48ILDW7+wPJqV4kiCpYtWe5jCy9JFQoUVTO9RzhgTe/
EiTXULT82444TjrLQNIZAajUTeCcLRCBABiN+HxXEIa8AKRNWUw/j8IZabndgUikAA6iJMCko3vY
RoGnslwrMJXKF65eaC2JFUf/tHsckgpmHKfZdVXd8RaMVc0xci4Rch67FLNHN34u4Ee7DuTuLBAT
rKWwGzqXnxfEpXghdKnyHImPOXDaSpv8IcoWtdweUa+KJtxiZmce1sgeGovVHYxAZ1QvcUEYHbWk
+SD1hHy18QSgOaAaSFEti2cSg5EjmYhx37pPe6v9aPSWirX+lMCL6FgUuf9sadAw1mNVodfLaTQ+
rlVj1bykVDyjgqoSMyjT3/aJs7lrtgdG3NRRpVYQAgt/VR6nbRGBdVYzQv4/IY6kOKZScnU1WqOr
ONGLjoYD0yUXX14d6eoAfo8WxEPSac/QY64zZR84Zg3aajHgUAtS6oplE6jYF16KjnDUrKbK8A4l
C5MbwmZU1G/QB/bZZ+x6QyzGozrX51IaJOU6xK3dXj8jIc1WGEvKIvlgS6a7Ij4Cjx6Swgs4e8BT
1CCPCbNbhNQmPgQWFZhS7L7Prug0fi686X+4lE7rhfh1bUfcQ0G9J01baHBCPmC90kxZogH886QF
gLCtCLTvQKDIPEAibLlgq0ILsojmLtqDbhixWzAfoQVJPQpHw+sdKlKyRsZNQnKU+VDbsGi+xqQH
F7gKBJvR2NF+3mz1ApbNBsupYcbddFSSj9AGGj4wGkxoaiaB60i6aBCbAMSrez8UiytUr3Nhx3mx
0xBxHW1qGarGP9w/mAjjtZ2wzK8w1e7HBu5IiNLebeIKacIwM+i7sRrj8w8jhWgIg4AYhCPGOTPd
dZMM0PdeIUMTrSfX9Zu5cZVcQ/+mCinGopRN79UbHRA7+gXnOYE/Z0OLrZPOtjmJnLa7gbel994F
8dDj4ifqL+scjfJBWHQPaFyn4WALihN1o5l4z6zNe3fnL1m2xE3XXxlsEoCCvMkmqaIlNiEKY1eP
ZKKORhD0XphHPhRAHHpqkcZsURqVksNnKsjDoy1Hjtn3RBIn1Mc2Pi8EYqc46qZHmM3tngtVyc00
tCqabPUOENGjeVbFc4f1nHpUvMmKEhizC2l7xszutarw/nwKFu8dVAT4JLJ4mADrLD1TSC787dNh
/6OdteTLzMgblLxW4jgQ9TzxBvc24YkaY7qU0YQBdp7XYcVPxZWfKN9yVo6vwyKvUmhXQ0xkl7l3
nccCP30/pHKY9ADWEGEbmq0woJ/ijrbMUIoTSewvsYq4WxRI14QmGKi30KkXpVAThajjeZuQ4bZq
WSoJ+fgbQ82p5k55czp3v+cSg0F7rY6pEZn6v0xYEd0T3xy3rn1Nz0IU4VFPBlKlM/rY9YkYNDVT
6herIBE7B1NYWLEEV1vlfYKkVLkvlT7UXRUZDwqGhPkasy+patf9RklF+uBfQLS8WoLbbGQxzoCb
+Yd5XRyaN8GyvxlI/lboyGG2bRV6/LGIlMqpZDXbH+SPdfZdf7w+gCmZnkZp8u0tGfjBbMTC9iCS
5xI4CU4wdv+DoXXv6ehWvLAcci/ugFmot6eRB4tbXJ0IRt9ZtFzasEOMBXtavip7CBYaaxdGbRlR
wX+rjEMRbmONPWEqPzUrINTnjWGleX3Paf/wUeabWKbKYY79DPdj9AYEML7ZgujChBGaFGycs2Gt
4VQLMUDXcJqMQWduOVFPrDtL3NYI1JaqEx/RMIZ+6kyuVMOKGO7pZZUAbn9VZ4vUE+W7X0hw+Xq+
BcZ+3qC3GFr/YB/aOfDK1mg0T1KZs2XXOlgEEYkeIkrjHiX7dzVbmK2RKUXnWJ3f8GZBD5AQ4vOS
stVhJyv9MVj/4eu81L/0keSK5q8Auvf6yxWEMNEOg8KCRNDMAON8idJYLslbrysLaKjXP3qQpUAO
ZtJqtS++QtxUYC0wMlbMQkpWWNnXQPGoVveAhI3WNLQu7JW/pFhIr1ftw0upDYfsfMKGMiPo8DfX
QO1h2TR+Mvzd/sMoxyZhV/vVbTEb7Ld7NRiOIVTcidC/HkcOKAG09slbyaLRTKsKsSgjqIvx9nb/
EMm5vz+eVGFDn9iTMgz7sbBYyeEt66L80l/xjBnuavjZhu7zV18fdOKJthuITvc/WdTKAvCzHhBk
qFPCYa+VnkE4GcIBXt6hDj6RVphFHvt5y4mMqgDpKBMsggsRUgwqpgEsuDUJ0OuDWsBV6j7tWUtL
395Uw6ySKcoMNQApGwxsQgSBD3/YfslNuej+5bBC3CSBPhpxQX4bEVpXPemlY15RNu+Anj7Zdb9q
4dukL3GcA/qfAMp45j6XnCrzRlkYBwla74vVpcDuEaz53dUlq+SaFYFep0VQCpmmEvrHQ2hXRaRY
ZSLhb1aN26W47YI5aiSgoEG6z1oXVk1TR2emAeFbo8y8ci7r1AgkgfQJ3fqz5FXWNSYqab2EIyXT
oJ3/ebHWeDUrwi6Y9aWvteZvNsPdYGMUi+DOf04xurgW6briZWgxtDkPeRK4lAUYOgTWV0vTJYxN
LaWHcJGxhAGMmMeGSOfHPB636X2sruuuB2wfibqPAcyRZUopwQyYUArvpdW3DMZIHhJ4nyCmTj4K
8RSTpqwqWy9TuZRfQZAe0Hua0Tt/VWGJ1JdUE2dWiYZkZ+cqroaPLed4UtzGVlz9g+q5Slhx/zDP
XW66Kiqs/qF0ICmjeKuYO95Uiouv6WHuh4C5AnL+FlXWqih/Wjwe+trxhj4DdKY2N1GNL9zSahtO
kpFODllgMFW/YAnGaZII49l2GIW4xQhkuplVFfsAoj3Sa+CUFeInPt+xVUfls27QTseSq6y6lXE8
u7VUuemrNtJw8dut+8UV2Tn+Oh9FmMAjjREW4OKue06I2ys3IetVJ1ns3WMVA+L/X01j8h7vc4g4
U7RHqLXJ3OxHAQQ9LRhv6adHv5yQPqREOjdcC9c0T8dhrv3wG9Ow+I7evu4tGv3K5eWbGDVhlFw6
Mj/ErCgue77Zbh9amzEPuJZ2DXWoeBU8C/hYp8I2ZzSxUmFw69fSZc8J0N4k8Cwcs3cj7VilhhzA
D+4l6xTKFxGmDbO0WQjrJn0ScRINV9UF9SzKPMKq834cHFNdbMnwExrmIolfbusJTI89Pgg+S74u
3mewDFnZr8z31lQUm4TdByRthDRTHvPn0cXAc7dmkdhl5FHltLQb3HjAgurmgz0QX39XmipS+Zxu
tSwkOtKH/gOb1vQ3fIaA0NL7xJLGrebQQ04EkSI9TDmvBpaKyIICuVZ8MsdPxVI0TRBY/ZcJNiKd
JoVoAS69QA+yVXKz+IeEqFv+WTgAWTQfELHR/JkB9fSSiXyaQ8ejrRUfasriJikj9+WYgEpAULdt
F7guFLwBDZ7RcgajjSX5RmT9WzMF3y89DQlm+Uha8FMEbAjL8oji2/6OvSFqJL8AnOR4d/u9/ezC
Z7tUco3hTkEqOHxODK7ToFD/7dCw/2ETWGoaUcRaBe5svfGHoBYqAXvDna4DzJ7PCmKaOKIrTbAi
Tr65+TXY1Wt8huEm4u9mwv+yfl8s/efoHFMNXqSNmjpjRqhDMY3eb3QBHpPXwx/Z6zWGVV1ENueH
nIqEhIYUqO9kGQMkzxJdcZ9igZzaZPC/55D7c35Socf92nYeRGdEr2Q6IoI5aQhfASMWxRVTq7ZJ
tyzUMNPq5EHa4UzUuNHBmoKPWjh9eaKObDlUO/DbSEN+jD7o0QKtsuAKNI9WKyhZfD2VDSfhDzKO
URKRJ3tAhHtCwP9tO6WZXnMLxipVv+v0ND7QvaSbuX19X5CuTpGN9Os0EWp34LhJOMkUWglvWFKR
MV9B8zaMeulSWzVSBLnBZ/WW+uMI518VXA1hOqVt3B1/TxS1lrQDEOvTZB11kzZD+RX3o62edmKT
fCMVpr1pJBd5afL9d+9SGwcXWgsErzcRVwfwSR8OidXGMTqxmxCQN3UaN3XyXmKSIPOvyRVWrfA5
6vnAIIfnFxEagTLRcdn//3+XzrqkcnNQmck5yXmWOr/B+wYazIXNmHmaWElajR9aybg7if4KgXEx
+GMmku7x4TZEcZQbWfO7wqY270aB7BTfd1mBTiEKWjMAEjzqmIWoEi+KqT+AW/IFwwO9ktkglcDg
JulIa0Rk8zOh8kr84lV2ilut7J6KpC3gCYscsCIzuzaCiw6jxn+pEA40j0UCB4H5Yd2Az0yjn0XI
tuS2NSMvjlCI7gN2mie79AULsKtY5u/d5cE2EKWxUX0veqV689BtB8jq1OpCmGN866xKQ+Pz4SmB
ywmI4kPU8UqhAG5qaIt1VHm5AC6K/JJCjz+8VOypOMhxakUtsmJd3oEYAlvFFBk229Sm0hr1oZDW
aOl3MBYVtNkeBTMH/GpQj8wtoK5/9LqRVCjzQ48Iqz8vcmI1vM6bMODLX/m2CT2d0gV1BkWBHnd0
p8BDMZ7pIdDWEQEvU8LkDwUqkSoDl15oD8BnqM+Rq0j+1LCX0wf1BT/6i4NdRDzWXuNJ5d+HPSHw
zK9jw5BArerAyUQfRY77lKd+aSaocovwj0mxt1qjizidrDACUKSqGdjnS3mnctX/GfT8bPptWenC
zZ6vaSQftLND5UFnI+hEzWLfzaGRoPp6I2eYI7nWn1Zil0i8deVsKY3t88RBf2AB2AWtyRs1/ow3
qRHLaNcSUHjLFOY9RJK2YReoYNPTNRlq+kjR8vWGlkWhkpG/vgH4DobvS6l9S8xhSzqeKbYCl2A1
8jSQKoyi4hzLepMwfkAKRpIfQeqwLaanJ82wK9S2B1uz2JtEfFak/5Ox9CXBDAY18uTnsOIO5WAW
MLUIvxkTiyyilkWnJKp4QWL7WjNY97mDtgkSXrtehnyaAikDwATqd8uqg9EdQtAuxxeLeneYm9XJ
BKLHVYCqhfWhq696SETABj/zFadmGk13FAMXFCPHjLb22+YZ3irHSEfmTQX8O+HxF5PrwwY7Daz5
W5cIrNOnF6JgEiWfyWbZ1qb7YlvonlWOTAGOnTdawFmo6ZNG2sjWfUQnieLrIRGeU5hUEPB7DtgX
JaS6Jw1R5nwpjwn56FRU+h3s9woMfoQCFsM8EuSf0rDpFp332FrhE5fAgWL2KkLIci1CdPLGo7o8
RUYmyt/RQUqNxKdN4pOmkxhyuMDPBO17WI0X+aRnA4DhepPag/Z7GnPHd23hfzvd8snFNxE8NfgY
VjEkE/+irFd2SLiF7yI0jbbeVIvIbKPQTmH6YjGAH+agxduKRG19m5Hwh8K/0xUmBtFTt8M+XAyr
W2W8H68kn1jASnc6QeJ85QB3+fKQDZFtp69hyFLkMLuZZsfBEud+7a3vzWmUQSmgHFPIVHWlsbHW
tYA0w/FxMaBkIxD5mECrsanvLALhpuEbmkH+wxIDq8x4gXWQXr8aUmLu5j3KkmDZEEM4nmnoYsVT
2JHvEejQxVzBZqAaxZ6dKJOjogFOtJR5+59dGVSMvt1Ogu28DcxeJoMyQROhG5nbWI0My3K6ewWT
V2t1u3HPhy9xITvo7uCgK6S7HuXIBkMIkoqVWUyANLNdWym/DC+ZfhpcfGXKGHcMXiuDjAw0fiLj
g0iVanbuhgq2blgf2xHHhjy5rpJ3KTSfHZQAi8ipwma+1ILHUehd7eUvj6IoUd+lbzID6zafc6vl
T+PCqLWkXwBAn3xoecA5vEjunBwfzMeW/xUt9vBczOSPi/pwWtg252vwwOvwjAve72idcxTeiVQo
xojcI71Tdt44FViIExOnTAkkgAaDNGyers3veeDal0ul29bHG+p/xXydmxAQPiVAsakMlKnleFTt
GvWJ5uITXR6eEGBcbXdy/UTUWBGbEaT3/jNsRfZVq8lR/qzqpZrlcbzkbcqakem7f0oY1U1SKuaD
nVGtVoOjKGIWXkKW6/W4Acaklw4WbRJ9l1jAR/DubiCsFj7lZdAMOzejRjC47mxMvbpwwzSqz4xK
G0HWSJ192LbUwRrvEfFIxMawOa1v6kOY4ejpJox8lw+E/mx+EW4lB0nz/+1SRRLa/DlDhdAiTiJc
w1A9nD8hbSGRbdCRaapbc3SeYAgpwig8sy9A4yYh+72XtUf5tm3VdvMhkVYZZnrv2XKQH5Xh/sIt
X31oKS8Ldzx/OnewAKxBlap/RPiU6YorsRw3o2M+mLXv1zho9N9YUAIlMWSNhvHuqXYjM0ZgnYc1
Lvk9QVh1jQXF//5Enoc3AW2WlTwZ1MHFXnGzi0jb2yHGfFKhZUJ66EfCvop+ZjhW38fMD+pHBj8t
Sx8hjC0X3KQjeii3fKnHFVvyuZptabnDSN0XkE54SrjiFwqTFhIvERP2qSuWN+o/Wn7Xb4EcnkS1
C4PFVCCYNtllr5ush2oUCHWDjz9CArMF3MCDD3s+amTqfxmLrECQ0j4g1T2FxEk40eaEoDtNMObf
4rWXbeFifHNcV6a6/ZXERF3lD1jI9G8f/jleZy6XfhFmKeqBzaTdfDx2GDwVZ6vm1hHzz6CfkFIf
VkqdTDf5Q6xFv5pCNPq2sAZas/tE3Z/tKYdA1NA+S5K+nbZFhM1WLZKQn+ZfWpsitGDjqtDz9EY3
qty49YRI3ogrGwIeTmdF3rnqzOETLa3YAmEhT42+Hl2etEnuuLtd5hymppPBlI2cT6zXGA4Zoiuw
CYqhpHQH6F2nkKNn8qmBqyKfhl+RV3KKugiFshcHDJIPOfwKWjcevbnnbovuQ2XepJYE04UeHo12
cuNQ3K2zHYBXzi73BP7phO/pCUG46ctZfbCsKrRUjeEyhrFn8mpuk40d5VcWbRigF+3mH9lqntUI
NEQSM6ETr6FbC9T9mty8uUbrW5YxwCmFMfyH6VO20IwdCIR7fgit+O2Yl2JPdBJKQ+Xklj3jdric
jXT9owIMZHF00uGwS9U9Bkct5cZGWSDFTCAMuzxPwHzSV5ybNZDDxCp+jALtATJLDR2k9XjajSbB
KSY0c2ymZLMnbo8MFq+GIPuObsSlXvKfQh9bvNb8EweLo13atJ2kL1/CB7XkvEU/oerHU1ldZxaQ
txvTaLbq4Fu1qkV7wWT/Eeogus1g0WsMzOg6tAEnPw3VKjNZcwQKThr8ihsDW++HVDJNJqwqzx+h
q5D5/rc7vv2odFQYisDQGund8jvygifG2ZrTXjJnCyE+R7EQ6Oh7O91kUS99AbgKQzuPaXrTpSVC
b/znQIqO+yUqFMgA61k/qniq1JqJqRfKw/ki+59DwRD6VwiQJU56iActdvXFud6I+iGY+wQ/4IyY
Y8EhDIjmjZkIGHLk2k0/JtrKOip8N9TC5I+hgZ/B5+94FlWm3A9H7aj5ubtcPIQ+yCaUg4oX+fEy
8N+k2iLXhfn0uou6PweqRBhlzt3exQl+yGMpcMEkmsJk77dHwcaAv9botPrlhVd8fW0h+sGQKMvq
TKRdshgWpObn547r4OAPYkJky2NhOcWBICTcR7LoGyhbRlTp/GrsWiGdYTc0H1xDt4sU/pCQdYtG
lC74s579tPS0+DspeJDzUsCm0vCgen/QvkInzIPdAIAjAhnCD2bu75iZbTkYKIjP6QR/Y+GVkXWu
jNWbkNXqyGri8bbHt+wse1J0BLv0CaKxuF+z2TbA3DhGKJ0J0lHNbbqXXpVtXUlkA1xlkFeE32o5
0J9jBbSsY9ZrzjOI83xymySXbTWyNa3ntr7U3lgsHWn0k9UQDh/c5bNEFN4DKXWTCFOgrtwuUaGS
EEAVH4+X2aWOfNI+fzN1b9hxmOhK2rT+Iv0tspI4TDZXEg6w8iHnuEAp1j6CAWy5D/YlmiCQ/15O
5I5Em8UkP2mYW07zCeBzEnYovkl/0AsH4XagLjT4JjmTx+96f/mcsJtNWrrFUozqicxVhrnJUAzy
KBelmd52t64JLwYhDnkSD0JnnC+uct2cN1slBbFdLP7hOjH6pCJ2kAY4axpgtC4XofPPqBTjGRbv
TI+initvuawA/yLsoA0uxRoObt/zvxBD4nYJw/tCmFo9BBxB2iJSBEiUpsOd2eUPH4xTaAgFD/6k
1qUlVMSE8BWd6aa4eswHh4ouH71oicQCJgJb/2EZiz51so9wfenDfpT0nHpxD/oV+rsFci3AHdf6
CRURgL6NXzXnVPiSkAi1i+lW04jxsT66ItgSNByLA4lOjh/d2s64LPRxDwaTkEm74o5diaNNka4R
HTVf6PYlQ3FIjiCQ5yx7RU177iZh7sHNDuU6jt5rGVLZPGziP6ICkTrd5eNiYSX799xIHv76ZLJU
Cc6QdF6nqnuSYo3qMgKu8LX58BZdPdgX/dQTNOEZ0K3D+uBT7ulgUW2g6YeViAs/GnmzRoBy5xSb
4Bk9jBfbTscUSVb+cyezcVr90pOpsVhRCHEE1B/iNI+nbH8waVzQtxXnqm+ZOrSxpGXxIizZd+V8
nkjDuSJa+GyrRjeEC0tBgwQqzNWYDIop+Xe2EQwkqxgheAotcbXudsAdwGgOR7QK6CfPy++rJxlP
L98rP5N5lnwTVJReVLu9GYeccRCJTO10dPPWYwNbVUo1496lfH0zd38KkzLimGR3xOocKM5WQMBP
cfW+7dHaTtjn1ylHIKZoJzwD8lpfw9S5IIWzXSvoGJ/8BKQdNvHAJb1AaMWlOxNoy27xX/ZebvvB
8sM8uflT15cKMwHxLmOW1lSyRzheTCoBpXtWNloAKMhrZd0VXucfmY9ZPOv8Br2fChnc/NEPnvam
Oebb3ds2CbmxMr2KzGpVQy/1+FlAbJqxM6KVzpnvR+mVH06OLi8+gM2Rkc+9RYXQ6CFlEY0cVnKa
ZhVkFv1/PwUoXLPOoqEYkKpGy8Y2BrlBZBQYtJfXNqV2U/roz/ZCZBhbG0FWLojgHUc+x01z1mys
qMUCIuQWkZ+oKqBZE3q+GK7rL0AAejPoSVI0AucweQeROV4fYYVCAJMvN8O4/1rX0fNl5X0arq/m
fBPRwGsDtxb+FEN7emoGPOabWjQVkiNRTeXl1mrEFAN2J5rEnkGZhHb0SxcyaQIRH69SXObRnf2Z
oN7bElUVa6A+Ea+AQFFCkgy9b6PNN74sMhixHXrn0jsgZeVEG4JgaWtUwiBw1sCKU7IXBfbTnCMT
cyyJ0hXak4MfUCEjHGsn0cgJJa165Qnz6b3DeLQ8rZ7z/CZ0a9tCoP9M3KhqqB/pTNRWCCy9vkNU
QMgEBeygs8he8PFhVZQo2sd628c5MvIFggC6eReQeZjjXBRgEjhmD2pgoCpffIOO9weN/b9apbIo
y9hhn9XnH+jjXS02ZgV0NCmZhVZS3KWYwd+rLhYgJpDGTylhf4loNp1tyTbKu/QUh1STXl6qktcE
UKKPuk2Md/x+MENonBakvbMyWcrSgvcGMWbpFA+o9zm5l9+dQB3ibhNopM1QMpsna2zDTZ7MnwuR
4g9z4SmsmPxLqStFEADZoe1/92LFTgeveW7mF8HswRcDFQAe1Ghnl7IT/HlRGfeu4v5sDJ5sVh8r
yCC64Zsvu6MSS6vSr97vtiJkTDzDKf2p7YF66a906rnFJXe0qxF42oWpI4ouXIxYjqVLehHFcMqG
EFK1LMXQ7dHrZuOxXnvG317zr72rtg/336AAv9bN0xOWXySH1ZAb9PKc1t1db+sA+ctef/Nsj0td
AXRg0opPaDZcRtRWbicFGlmHflP9FX2sxafUBqz4ZTQliE9kRQ0CicuYbLwPUIH1+4yPArbuskYp
E9WV79Xi8ikSMivcD7Jbw2+nt8EWT9B8yp/K+LXE8izm+A9QGyeH02nbVZ66x9QQZWRe7W5zUc9u
DzgBQGfiuL1hAfnHw9xh6OtzwBGXPxPTHXlMXwjSquhgwEzIG3vCehISn+w5g3BN3pstxoWM7PE8
+YA4m1nmLuL2ZsX0oihjinmCNkKaRZ1GdIlE1HWfDibR3675AOpG0mQrlAM2LBBqi3/Nvs8BFtT1
JFyQ4jdOv0PmvnRVHEPq18J3xH+62kKrABKNsd/a9l8h9g1HpA30ERBs6llP5ErI/yI4oBalc9pz
msQLrayOmWLFfnthSRqK6SGfw5CXt3I/naT+GVWiZQFGkFOrnlwdwYEKhSGdg1mUsuIcwT6stY2Z
bvRES4IZTT+MKtQ9yuqSOrvb6Hy65/y6RlptUgvR7XMS071eaJ6ePk3ImwxqIFHH6oXSN0okBmxb
0IkXf7D7Ad34UxqZTybCq7R0H35G0dgRTgdgy2pX1kCNgOf3jHAUaJK0gAAQsCyPVgJZ+UiPgmhu
NN1/9hV9bZVReDrgq+aFOIloibLmn+359+hOzE139D5n8Nmh7xn4uIzFbOMetemi8BlAYUak8Z8H
C4dOJrEiMA4jkn8q9KIUt+bGx/Igau7+AstG9XK6cAcDI+Xgt/3GWhTeOZd20P5V1di363W1ycsj
AiCyiF23yvIVFZyuqMvwUjzsgdeost8v8twtbb9bc6fppZy/6VkcONeXRlVi5751nJIE0hh/xioI
BBvF/0SLYr2HqKGaC6DBXEnPqwgiGD+Sr7cFcI2R/Nth+jeEqU21WcviH+rIk6lIfzLTcLkmCaPE
q8Vrg5MpPBqm9RYW3b8luJ1u09n7w2/w1vsQydfjHsIf0An/Nrf2jVgP9al/YfPTLiRvPy5Gr+cb
66FZApd9N9iZSxbXP+HqwKqsUqKqoFbvC2tJuBWybeW2k6oNeB8onmuK1AhfVqrJ4m6O69XXuUro
0gVe0wMZcfgZbrUDEqykqv9E2zH1Nn/BGqBEhtsPeEpqp+W/yrHIVXCKoXPOyecmB14nAGzLkKWS
HPw1bOTkuCMKxyvAStXmok7pFIWjoLP1VBv362nFP7lO0Z6S/6rb2F1fLcf3UWtwLNYZNfGoHztx
mJUO/jR4BtTVl2SOgwXaFwFh/s8SETY2CLnVrVYJfLF+ZASv3yTO/my3ExKOxcqzhKj5otMve4M6
mS6rhhC7D8Tbc6Uz2Nyr+Fy7CXoPQkigbLawFhxL5ayOjggd/fb+3QIjSgzX7yjCJPVKRMKB39VS
0gf9XikkLxhC8I56A4f9fZ9FdODlZUlLkVKqGuAP0KTJOaBEF32scxz6ryGI1+zIg22pDRN5mMc2
414Tbgvw8ZG59AfrCmGe6SjYsRlhRsC+Pit1M3bWuNLT+g+sZ/EIBRtmkYfajl7QyDY5Fj0XKNMT
R9GEUB4xonrQJxoGn+AWqf6uxVP0dbG1OewRaKgNBFRsKzZtxdYNYYaVGkpm5HHgxRi1M428fIMU
KzsNFWeWCJwC+5rqBdNfx5ntb1mKpT33HhUSWqNMD/LwVW/k0+0CcFaq899JuIdpE7PO8cHjFfA8
OToi8znTtPVldcHju4mRnfxRabWQMfEj2S3+Soz8pjevNQ+JCSYwoiSGubznyJlBQnglOWpW4PIP
YVtTtEg9D64TwY+FapdTgH9Z76GIBTLvI2+qYUSGe4K0obm4hmJL2r/UBQAuw3ZyjgLHJDKofwF2
rNjUPaQOYvmp5DDx2bphop0B1rJMMGZPTRL+FKVx2h2tGOfaLXqSeqxmbFDfNYSH3Hxz3cNX5TYW
HA/xN7PTj9rJIfjL3gnGssEEhMYfKJG9WJwHbXC//Uevm9IUAdmN2ZtBot+H9UNb/IyWbL3fPqET
qcI7JQbe4IrBxNbV0AEGT7Sjljyo4c3chNU9SOIReFu9t5xAZYGUeXM6GqsnaQKWUITEHO24OeXM
3qDkSKBWmCFhl+xGEP4k6E9DyxzdodaPxxVa15FbN5XyhSRUDNZh+VNdvzuO3sQERLvzI2JxpjOh
4hiK2q63DxV2NyKhwQ/NRlBZXRGIrWizhbQXMIY+i5XBl7vx22mR9Dwen7mEKOEYpU3FAWrpdFzj
4CNkPgiLRnM90L1aQCFq+Uc8zzxfcSZ5pn7rTxreZTO+v7TS4wMa9VmC4c1/p5s3WT9KHRDscOGD
WndMpfS2kjdz7V2es5tRJqfxyBUuxHft/OJPFyefgKNXb9zfuQPkPHuCxNmD2VtTQh0bwBHseodg
xHY4+SNRMItokZ+d7KntJHL6hiA7UFaGOXfoPJqNfCd4vXZtO3LeQOuaEwcizVp2E/tW2mWkuFDh
bgiryPfCIB3ceH/vlSv0c770GAbsqoHvQI6uFHie3B5RxFz0UrUckW3SdwbXMQIp1NPd1WjzbbBe
fC1YVcFVWvkiB8ZJterpUBQQWfd+wWLg307dnN3Hs3DjDQ65y0eHRxNeba4qNMskG65OkePoIjHX
whOP8Z2IhwLNtS+Lv4OQ+FpLsP6UX0ui/3WspXMbjYyZy5eqKHwlC56v7aW5chXRUgdwawcGg9j/
apXVTBZM2X9G87VhEceS7chdCnKDT/Rjj2LWlv8P1mrl3Q4jLYHLLvhhY7Cf5ulUW6SZCKGLFc1O
zGvpBTr++I9hHkC1hw0PqYtWxwINc6QepPyIJobGeIJnu2qyBg5IbeMXSEo504H/4DEXgDB89kpQ
MUTxcM48lb+l04zS/N133KggNaCbbrveSSoV3scdWFuO1cXcu0IK6u4GsFt9Aqu4aRnPhiD2Z3LK
S42HrcWbWEDwvoYIAsmEawuPyaBczTUtT71OAsYsC+egRB/RUwIeKRh0oGMbkymB0ULNA7X2KqnT
7HV+SPwYqPFMCXerwQb9xbk+d9oOlTCbfHo1aUupbjp5JWpS3k+jwttFomAQv+bw205kygftfz0C
IJ1Om65mTIWGmiv/zP+FwxOsj6A8bU1d/xA9FqvLxbDSAa9VoAiLfCcel1l+YPRiMo3jr7i4xQZW
B5MvAKKlsJuEU3Eocf+4/bo6eZ2hfhsHZOH7kS3zskwFETLzto+DddNaGyGM/1mXbPo3+Non9oPB
VR4ZioSZJutzM4JpK+ek8pB6ES+2RfrfVhBjCAUBoxqGdtDXIx2cCunjsL4O+Gg2DBZEA7kLV/AD
E6bMTvNO4W/7gHO/kJpeUqmK65ItR3c2b7/tbKFWNeRNrvPMnGbVXqe/PzAakVZNlPKcG5HgxRt8
hz8XXB1+Ycyl4ZXnt0RWXQzb7WYMt2njOzo3Dw2VDeBpsbm1SVA4ehl34ROebQFM2oyuJAPqApJk
cdrYOKnj/Ri5YnDEJ5KTJyY71utWdJHHtqrN3lRYcIBKLVTML1pEl+M43/kGXTSvI0E/5bxUMFo5
SGs1QTCg0XxbQOhhM0JMUO36OJuwHFvAyYne7fckN1ev7LN+90uAlUOMLzKK/B/JEWXr3tljwftX
7rE7Wx2unbpJ40NQ72xQmne22sJB5IskPRcvtKtuwvuOjLLJ8KBT9aFyG4pNFQnGptlv5fZMzejo
tNs1mn2CVg68ORXQWUADZ01uojkxTvWLuEJGuotr4mVekM9TIeePST88HQZRoFTf5PiKRXUSGzte
mF/4/nSwyGj1kCIqfnuHNeCgROw5nbZfs93oUCkVYBcv8IpjXvrAQhOK38AO5d8xf1itNL0DpE0f
HD6ROi0qE8st6CYUUv3235h5NbYHDpbPm4BT60zJ5RgRmFzGhsr6n85vS89UWRUtG5hWUb1jsUkh
RyPMUgcZXch+uiJzdMmKZo6pB0A/7Xd4mazLty2depUOYKNSWtLjgXm6IMifPOtQsHc8sbDXsmhi
bsnbc3pwUPZpqvW+041qdYY//f4UTtl80a6OM+S64D2UPrJC7hfrNbCbga6pM3MeM01bP7dIh4ZN
21fes8t9DzmlNJti8Ya0pVOvrVq6Mx2ZAKCobQ4vtoxQVsiz2b/IjJhDmEjNSpI0ptDDqjrP297Z
Hr/SMOv2J769KCPZMy1FyO6VXE4kmMJAIU8Wjn4/abmvnTZrapquIOUSMxrZ6TxR9PuZYIslpTtS
u1foDihH9aGMeuONWLt+371Idu717og8Rz5GTofHXyY222Il7eCRl74tqhEEWDA7szmo4/cJwm4v
H1u7nnJW1IAkovQFTrWoa6y0zaq0gDPDJ/aDd6woFNfyvq7WiNFC/xyiSLE4gXIT7GTc1P9y0Efx
msRCIsMwuHOyOZbSwBDJ0eX//8KQu0u/yYwgBWsX/N7U6ze/k2GzjTpB2Kk4VdVYtt9GSYj7Hlhm
E8+qhF91kTBnOqpxUl2y4nelXELIqWff9EIyn69ozaDV7PgkAeqGcyjnHjsCGxPR9ow2KM8eEIul
wbkYSgw997bxOqeV5xrqgobK/q+54ofICFs7hzSAdDWyrw6AuD5XTbFnHbKUaNjiGLvbufo7039e
RBScmj7zV6WckNHJvJ4V3fqulIuRvePP6KwcK9KCWBGK83LWEKlGYh2EL3FwEKGYPYQYn7bYtC4m
rZvBbplyyllQL7poI4IH991F1pV5U0SHrgg44E+L58sJYBFcBkCDI9wWJSFoTsBFnhMvZDBUxDNd
bxxAnhC+2mLY16DHRosxdyxk/g9XTQIRaEFvxAEBNxlVOL/5y7v2MbzVgj9v/rqggdUqrP2qF4aH
TIL9i03Ncm081ygh/OSTVbHhUcUUe8yxm4/HfkkFyUoEQEnfaiHCmHsKAYamFq/LRaYaa/i+zYoO
aPgtvITjC1NJwFAti+Y/Lxywkqfl/SGoVfP3t2qxUwo3HAZJyN0QKjevTSjBUb2GxTgwODFKCR59
rMUDWTp3CD1BMUMKZAo9wFxUKCIepRSZimeoa5wAAb8Phc0a83yzSorBoh0NwQgJWVXOSFBIeCUL
T4P/BCdnKYNNr4aDZR4rkl/rXTryF82zdyPF6pfxaSLegcTNJV7cutcfI8+J2B7g/T+7wyHVlAUC
qvsRjEaqdq9S3ULAYrM0ed47oW+EVmdQo/MAOHMhBEi8T3nlQBcXc+bW7JaypoVqMfEcFvwlf5cT
sGn3xJ1eX/HvIWlVPfEZ84HZkVjP2ntA8IUxV10rICXjzdWCXMt/+U1FQviyagnYFQbh0C+i2dvY
CqvNznBrGnksTccp7sdU2fgzym2v/nHkzf7Y7emAhSXbGlnDCnZ1xDOdOsMYaAZyRXygLnogr2gw
rA2UQzrujEIppWxGrL4uUvDo5i8MzX+SJjr/aKMFGQZrSI97jZ+0Ff4pEjiBLU7dMbg3Euvl4TKL
JLdfFuzul/JzVAUMnsTvKcQEEXfdS26wdryGvNLAy1FMYmV5UY6tkoXMam1DSDv4FwTJwjRU+mJj
oBz+tRDFlwsKN83aRboiF9HLkAOTsw9VqBcpbNnbJuJKGNsdgfYk25mwjKmf4mpEatDqbOzUBwYQ
21UzkYiOhLduVdaRT3yu7iPCLLcDuCvK4iN9BSZACioqPDuFhcScw4kxpApRDZcXwOZccLHos0jc
Yt4pRj1EjT9/Z8ChiZzRw8vibwtSxclra+viq/IB1g5w/6zXTI6PmO8yQSt2Bf7A0jR+IvQ1VoYT
ruIl4el+CN8D+surX3s6cby1n+PqocC/Xykul9IRLmxPt4Rom547O++RD+E8wU44+exBIDbg0+03
4eFVaiSvElDoK7bt3tz1mth+9QkIidU6U0qhdwrPhPMBi0seNaBpLLFYsu4BgHV43dWyq6smCgXY
Vb2Hf/GVN/drkAsJC2yI2IrLUCbII5FCUV8PpuLSbBjF94gikuJdxi65SmDjnnTwKh8MW0JtWUFo
QkUy4dA6Kv+4ChXOZpM/HdBZMREGEyhi3QtwPyVSyp/0w/kFiyOmL51O2n6u54ZP7NjGgmHpseRM
mXcGFjc6TXB/RWgMcJnysq4Iq7MTupHwLiXtEjuCbtLgo4Q6d2ZtHVfEgbhJhQsNY0AHe+SWcEWE
WwxXf4I3rFWvW6JLailldTbAT4PQKbeQfSB34oavEldoB4Uct4dkI/4dCAiXPwCj9ttKvuZLAKBw
ZGxqHev4RwHLAt972FDiXH2s23ul5ldQgkQogqwkMGFst7PmUi0fMUna+VY34l7QENcFlAtK+yiy
Q5DPZzCGEUetXJs9cHoAc5s5we4etO+fkvt6ATCLqFw5YpaPPmyPqqMskw7vqpVxEj6G4093c/Sx
KX4zYmTEWIR/FwVuJxB7HiQZr+hP4pQNwww3L4rxbQgxDyeodBbySm+/2kylkEfeCUEhZezimLh2
eX+3iub7jOghBIppjyVLCHcQT8eCfwXm8h9h3R8W8T2e65Y2Bp1OeDwajqVE3plc2qBAuRX3SMFs
xs0VD9OGAX29tt83KEom9eR/5hjDoTiM6qbQB860YUrdC7SAzMS+CIEHM8SUrT1Mil+VTVwrKYIX
bdHFaQzNjSgd/OePc4M4OzlzSutTaOv7PPh4rwKJUcgUrDjPS+Dte0xew54fOKjRpTj8mSxK76QK
r4Z/Eg+pTOJOW30KgXWEzoxuVfLZULKn/BHvPY/BElyL7af43awWAZ7pUvuLRbdwkTU2ElSuJJts
SBP0YhzlYwUWoy3ozi7J0CD9lC9eAlkN1h9MvctwHE+6hQ7mUAgbhmXoMTq7eamWZ/6hsRLI6RwB
lWzss7b2xM2XYW8VZ1gGisLq2SKXHEEMkVwrRySbKcMyAYadLoqjTRLixDPcu93D1RmWAkVlU4fg
9douAlhmd2ydJrvMp7eY8eLkZ9InGEuDuDZAJtx0rOkJoNYE2HWiUAy3e23oNi5IsEOyejEUCt81
qqB2WL0HVYx/jCrNXo1uhZLimgTHgy2Md7/Bs6DOHTDw88a1XKHLnqi7Or5py7C7ydJUC7tDUiws
mxQRM3dtZy3EDUNSe6kBFmLy+GUzekhcFMqWapui/T0qzqRaluUlwRQtS0pszkeWbCuxphhp4zzK
L0AQowRdpU5kY9vd+jTD+7YECgrRSVC8nnrJNdIes/lUgursrr8IcJEIvvuM2q73HiaKA0O5HHSg
kqtPb7u2bCdWsu57dBKPBQ2GthOAPDPdwdP1BnmE1telnbJY787/yEDbMNImrdm3TaOuRYmlls3a
Fz0vqiKjvv6sC97dWD2NxGvSFIPF91UmRtRdUEWzmuq+PYi6uP90UgTrOUGNpmS+O9PMVH14xleR
Ba01TI6ZFFpuhqOI8h87Ap0DbfXYV9oR5qreCuQ67NdNBLMkn+0ndNpTFYaDDDHJsbCtg0J6NKt2
5EH+egLS9srI2ewy37MbcZElp/sXP7/wfNfaCF1Pjayghm2vs7C1WJTTuQ/FhdPEHhg3RsTxBlqS
LauBq69eTl7Rz3EDgK2uI3xDtIJJf5kACgEqfkdiRxF55Ji7kLOXv7XDPcaYPp9OY4uLkMNS+ZOF
fz4xgNlMKSLQ3/QCNVjCi3dL9nwwWFHB1Qwd9uTfDJUhhNTRrpUck/TOVojahgi/trlLbqQSW320
uK7JBMs73o6pgg5BHaaL+7jzjjdeKiO96OxEh5PWEuIU+lDKp5mcfqsWwn28p/gT5ukPMhl9tCQL
5FQZ52aTwQ65Yimdvl8+O4I8Fem8h7Zb7DgGJxF67PP3CV5TlGVpfSzwjDYVtLjjYRxs4W1OOxjy
nt2joIWMK75iEZL5uOCVHuqpjriKptgEvbzv0xUN+OdRDrGbL7VPsAHD6YN77uvL2v7uh61iaz6F
o+WmALtl7y5N7a4vRi6UOTTMHPEYSZFaOrpMGO0aCspe4BwOjCGRR52oFi69Ru2iE2B2z8yul4ls
4RSNK8tMJ0RphK/QCzHmyyUolwA/2K4HzY9zQFD0wXikmngJ8E7VHTHEuRV1rzH5t+rcvKb3L7Ri
3TM2yFZjE4kg81RCahwaWDL9WnH+La+uz5udgZMJ/MFOvoUan4D3QK9nyXOV1TKVzYwfpIdF13rx
1oDeG4QyvIGoIUpYmhrIlWkMGTQDrcb7uvSHB5n3dFeYajQoUEk0xMqATo5nHprxLQLPC3fePtPI
3v/1AV2UFkjmOZdSQIUrQPHKiMELZvPS/IEAkzVuJxPvRIwKb2YopvX1It7a/VW9cS7kGNUcsBe8
GUf0q7qtXeeb0o17nQ+hYcXQSnZaktHiJajEtFsiu10SlKjtGK5BvLG2hwSg6Py664oDnt7s9N1T
Qa9uUe2QqowVDLQXV+kB+08xxC6ro0Tzu1Wu99SAcoA8wtwMqVlGWVLsdTPgmLYP2f4mEq2e2EWW
cYiqJ4SEaxX9bxEHLfTbCFFFdKt2fwSVf7o8ASEeNrtIjwxt9TPMTQxgFwPEpJQSt2LOGZH+xaOY
KFes2KD2D/LEWoslZzzonStfZ4ZzhCOQbhcZQxzkyFsIN0AA+tM+4qPG678Ek/eRmgc8O83Eazmi
kUXMKaz7Li4gOuzLSi3S6bsO3lSfkfN7rtB2YnzJyKsS/USdKnBU5mKgyK8VW7aUDTvNlcWuHKJx
7ya6c9z6yQBpcsMHMcyu9jotzqFc326To7JQ5CG4hFOOQwGGRA/hxoqUod3sjOylWq0qJ4HH5DSr
rPiBY3hyDeIje+bjGlA+2v2Td7dSvKiUVvJW32YsERF6pfFo6rIGgoYL0Yve34Prx+JRZzKOy9kQ
3R/QRMEafygz2ZHj4n8Mw1ocToV4YkKQe2gGMVNrMo4He5AynOVTB43sEunCB/E3gvDDFYUDIW2H
sV8crq3UicCXXQ7YKwRZ6OQaBCxe6ItofS9vNQe7nR+vCKmMewoi/XkuQfj/fbonVntGlnTBCliF
a6hBZWl7LbCi42GwDaN+sb+hDG795+5XHwRN1KMRl7stv60Cak/5N7RjHEjdhMeAjmnMALwFJw14
LFRncVmvr/+pS/LWODd76SLPyoeAPSrqNBYtqoFVM6uzHUWxBMs9a1PLJohA2CBkY0K5Q48ZiXjy
NwkJ0ITCXfG1WQAYiK0cCgkaOef88BWoZwZ83g8VUAo4PuWPuCWwErXdxkPMgQZyoK1Rcpvg74qe
En6GkZhHvW7JfQ4w0uyZCrTOjiwHKQll0MSLi38NzbGsS5PqMyUk4NINFE9FpiASLIOxtUvSuUUD
e6lUik9QXsJllASpEgGp8eu7dP7juQRGnoXo9wrZqTkNj/FfeE67tQbdmee25gu/+jVNW/daa9dd
jcEWtlioe0NlSrylZrrLtKUpaKK4ZOuDISNDkvd4IunOkysGtnt4eayBy5NdCN9Mem3o/RTsZU6L
pWjlbz5s6GdRzmIH9tSHMUc296VuBS7oKCz/HNNHu3SsT6iK+dRsqQ18bindS8KYqMxxQDmB7ga/
J0/qeYZVlvsbKmcIWQku7YncbhNnnBjY4D65Enr/u3UwIR1kzUU4S2ykOLavY7VaQf57poaNVKkq
ABQIx357m6PBG+dUkNRIzTNLGOFJNbw6zMpI0dqTmjk9YzQRbfOOCn0aQVBABCP8aoMh/QW7HFN/
j3YhrVVr+lLo/rBysyOKBDvZtlAQ6fLHEZaZ8UGH9lrOcGPuhyJLoSnDCfJ2bIi6cCLV32EVx9Yv
BalhJwjTwR0aKWTZOHnTTj0HUxBKZe3FAN71kCcmy6wvXWOMEW+RbY5Q1CJqwS2ghnQGKmyFGlQk
9tuYYjI6F1lrqQto6OATGKSyj3ys+7vYazgNAHV693kKmv65mP0QeaEcczNg6589kJM0uVpRObJ7
mHqggKU6rtwyMaxqvOUeNK1OSl3stcp36bd1WludXPd2lemKcYMlEMubP1P+G3NeUY8SUiuHaPfj
lgewOPpLHtZu1uyVGzV2nz+zJ/lU4Ir8EXT+WaP/Lv9dOnVmrYKDtxPgVY1fkBe56ViMHXcHRHi0
C/YtrHZq7g7GsI5gYB2aURqAtA6QjQIWjyKkXhvb1Lxjj19VPCMj7jNs5yFdF9Y+/JvnYVxSsomJ
02SPb1bL2YpL+MnY0zonpoUpdMj/fl0ZnIndzQ0ciUU8mSeoHP3WyELsQOySK8n0Q9qwRbczhLEz
v2x/MyNk7uuUmi2XydoBiU6CT9bs6KBUwWwt+px1NYgp8HM/op4SAafg6Cd1iH9XsEiXid4ZSYj8
ggcmkw9f0B3rQ792jM+/LlBNSjgV/aTJXjuxBDDxJ9N0AYhO7rRnxDbnlQJjLKTEet0KZWBBkgPB
rTbCdkMDeYfLXhaXOzAUIhDh8S50XJN8fC4EoH2l4MN3Mp3VP+f3qKxF3Vq7QMOE6EVcTHYmNimW
MsN5HQb/bESSmDIIw6f+CYjdsg6Sb3YHNz3H2D9C+pkAjNGejyI3IVcAV2FdicfdhtrXU8RNFjMZ
mLQIR3NA6Pw2GcZXa8Defs1n29EnTaM9+sQaZEv5UkU5GxNooeXW4D4YjMWDeXWXkxL/DwovgVGI
jo9Myr7SopAGnXbn0EeJtvcI8A85kLUIoeYZRHsyrsA2/azbwkwO5L4FdqySbu+u5We6j43XIuZY
BR93PSlwa+Sdno1hoSC0Dv7cOTRa6pJqYNNuP/PkTxFNB0A+PObbq1CBmAhtBwxZEYO8Hp3UZa73
c9wfLhGXn8nVZ2S2yEAJt296NpDADIAy0I+T0E2NdjEZ6nApQZPWoRZ+X4gNRHjF915Tz0wc5qUa
rxQ+so2HNOeZm1mAUpba8A/DnAiQV7X3IC69Kh21Nzmv9qeoV5rQbcINtS/CGgm3zps7kTvgq6Gt
LOsSLDsEdiV9ceMyaXtqZCv2nsbyoQ7E2/eGAtoUWsWt72KqgTR6NfdBy+3hULLzPX1x7TjRt85A
YMk5U8GzqUFQ+7EBfY0geuoPG5j8zsDtPQxilUW0tRY/xi+4RcXnKT9WI8bLjBxwg1MpFxF1MCC1
cP8Lqqnhn5YWGH7iD/IhCQLmscydGgae+lwkNn/sZ6YXeexx/4wvz2mca9u2YDVyXzBJC17yxmcw
LdQXGsPvY2z8bDnR/vCvE+mv94u1wV/CCKO7u1M6nvg7iv/ZEHVidamE1oSQG5+zDsJ4UnfiZr8C
sbT1daxiPFyn4xnTaQQeA3rAnMVewyXgOvIvj5wY9MVQLQWxZwZ05ugN601odFqbZDvE7dzQJOGm
B1ZQHEpwCKI/PFGNBFUe207nwrNVOolr/T6A4fDMm5tdjkyjxzqKtGtVtR5MRxIY+swZWh1egMA8
W0e6q3vI8na8ZYAAkifhfOXkLzNul18PiHUvVjWtpr2f69VKw80RlWfd2MzId+e6OQ05UywW8aLP
ceuC6HsRucHvof2ryxD187UC4nrqpeSrGeRxfRlYpfmBn0Lb52KuZ2BY2NuLiBFfSABG0K0Qbzpg
MQleOeyAXqH6xACUc+sEDcqaadUfoeOKrwg4PCSZ5VyNmCr9I382+2ROijHhRdKj4g4xqvubA8CZ
xwcDQdqvty527APK7PvHUbZDxXcKpnHIPXVlbuGjOfLrUt04JBjuAf0QTXU7ri+VeEFKYPPPtjKn
sVed2KLPNiJ0GIb3R6Wod76stqiy+PKy4K5U5DBG8Nl8Y4KyS1rT/fAcae3BxOSXEW4H/Zgj01as
7UbHxQoxF5xXdGXdR2I3fmlZsn2Qj9v6g0TMslV6qXsSkeYItBGkRa346jojNVMMysqJjdsrWaQA
zHEUM8nkV8Ib8BgvjPmZxdgCT/z/D39vsThWO45mBQ0hNNBsPkY/ODQRarKF3mzEMxmESDntk/ht
vkcIFZI6RAmKrMnULPWKb/1Y3nV9gBUM/j7v6j49J6NuXRsp5cyEX2wD54pY6WwmI1OyvxXZZsD+
orug/Km6v//jqOB1x78wbwp6LaH5qXkmDQtN9YEHhJQ/2AR1WdNJrdsH7J6jFqN9OLThMpKYmKaj
tOphTiK+G7Ob7HLgdwL3dEb35K+SGxQ02RmlCMJ7C6RmOQagYgwZ1tvdDr9RlkfU0p/2QE50iDNl
TYRwEPPvBU2v6lkotolW9HCCu3i9HvNJ8iMqtsfvHLO5K1J6AmfcVwrmKVIGW3h/uqfUPZ0xug9V
/TUmNLkwFHdhYsnxubRF0xFAc9Uun5qav4Q0DG0MG9GV0jSS3FAEwy3ms6ZjD4b9QS++ptJhBKny
zd/5uh7/wIyd10jnLEUuk8jLXaiLsZ6/tr1VaxfbFxSk/u0YGNp1cSRULdHoGqhCqY+t4rRl6aIg
WxaEBtgDMZw2q2UPM852DvLk+lfa11meDEmOFvdji9M/oSpMF9ur/GxlZadz4zKL2chlkf8KBgZf
YYQAsZVh8KOkoGrlcfI5Y2xbIrxFOUV2eGeFeBo+ayvxK0+ajPVLiMY+kDhJX+RtsRQoYlhVjGZs
kiuh+2tFZjyu5QBcIkre3z1L+pQq2uQr+h0luiyOLuqom1NePFcCwcqVfnykYsZ9nbiCu1W6/7mM
Q7QzxWNomSJv1VOwOlL5NI3BueY3urWORhjs2T4t+neW47Nog4pIUXC7f2yvcrIhCf5/jEKfiYrM
HjWbxi0Dps4Kn/CXWbWd6xJzbFjS28zFtDjIfAB+H/5gNk69sv/JUx7H+eooiWHokVilcsJq6/at
92uFg+PgdnCcb7DJFwSLOkVo4ZOkyuO5kYxvzIo6UkIyY0IoWMAe/ESm2lPbWVkEYpCFgZ4Xfbyk
Ephn3lBhwOtFOGHw5xGm4991bqdad4iRIlKwSAbfMEWXftu6U/Lrzne/Ug2uFCWrwj+8HnUh4myZ
XXznpikABNTnIJFTQDFmiVdOCjWhlE9fOseebmGebD7MrHFnW++yjzH56ZyVkvGyrSCtJ7+Pp3Fj
/v8AFRyKSbMfpvdb6YN+YnhhPcEkcKzKxgNnzx8YtULojZHHcyVa08hP2YD/01j+RFHV0UfCKdy4
QwWwAzuths6WouUpfRCcJ3C/zALc1T9aQcMyLe2Hx14cP2ApJuiquynDYiYDw4RsZfuqrFwTCcqU
vs3bSKp2nioUeKixPx/NcN586u/+I4eiCUP1Ag4zW1TadfK/HVz3egRmMlhnp6E7HTu1GAytpgOe
oC1dWRz3ml07RSjRxGGV44pJvYOufVAiZSw2vEj2eTt0wE3gxbtWHZ8Eh5zy9P+Fx1lXbfboXvbe
/sm7hQQp37UmZ1FGyGbws8kHFEnYst8LP7sYlOlpqKk+FfwmQvOPkctse6Ch955x6A6g2ihX/V4q
3DP6l2W4Ct5yvKif9s/hWVofSUnMXuYN3V+/VzGNakSSrWxRB2xALEanBzv6xZdz6BXIWdCjjno8
zhGUdYfX0+4prJ4q4PnnvLuFbUUVwIe9ea+rlNXDGnFEb5Xz5L/JoTNSAMvjFvkqbJxA4rGTgCQA
EBN0VnIlxx+Y6mbN63M0suEyGpdggC3aHFwTx+oChy5k51VkYRs32JIY/EfscLbxojWDGDny0wPW
ZQIgQjtzkSCmhIxTYnTBn8U3PycwEbYLFPg5L0SI6uUeBjZ8EZrQTHEJWKmfYekeKRMWbY6aJzbc
6kGBmQNCntMQ1grm1GmCKmP55RLf2bM08eWcVp7lvuh09Rxg3fWcwCGUQNomLCjweLN95B82O9zF
eab/pylGth34IaKdGVBIp6MWYPmcCMCsiYMieefJUFBklwy/Su4UDIlsX08RDr81CiXp3k1EQbWb
dQGzicU4SCqM9e87pxh0JBz0/+uyQEe30ebE2CYl058CToblsu/jByH1BtxIwcDcqk5VprPqwV0z
mdKLKf/XuTcsXADuiJcb+I8KahsfdEp9wEXFsbUk9jGqYwizXpTaYdPG0/vaieI07KO6ux+zsfXb
WtMCMezo9+jFTR+BeaQNUwLO3uMmAiCcC/V98a0g0VNI4WMXEY4GleGFO/Q0/cAenyxYmRvioKQT
Hx3sELhq8agzQcX0E3H3MRDDky9IvJIGOK7AX4FkQci+8YS2daKRvLXFTr8GeXMc7ZzJ9Zud6XMx
Pn1oNeRN6S2tCOOY9pR2qbsApo2/OIAJztnssHD5gMqAHRBkLJXlgZeZQ8E7nZli4NIX3CCaH5eZ
lpmjP7y1Ze4DNIKopKPZ9Pg7gNcVBYr+YkbsHjIeg1Z7sripFCc6Em2fC80rEF5SyE7zaniq/TF/
GjjH2C5n1o+M+cCBQ9GI+vmKMHmYKJ6R3oQR3ciLt80EtK60gOMCISyFu8opFawedEZURl3ovfuL
imuXEqW0A6fxwA9NPpnfemI3k96O4ntPvydVjbxSdgnX/RB+vvTnJTr2T3nyb1tsO73M7kRbKrVT
YN0izGmO7CD37G7Ny3DtXphPs0Gmu8d7DDc9QQQpbsWOC9EbnMTJSDrgLsKegd5rkVvVHtyVLvPi
p5dhVaT1hQWenYzTT3afAWTeO2klz3pjxZ0IXJK+iW9aQXBSuF0VG8vn7qjPcD+PzT2aVtrtnRKj
0WToF0kbpagqpkAy4NKMINm8ajjqeoSCzVyUka5FslixXQyS5Dc7TxA3SKl2QaVl6tuUhTJlIoXB
Wf+45GQjiV7o01VD2xBeKVN0V6anNFGhEL+5Jkw4bBD7yzikrrEGucmkOTd5mqygr+mAeY+DFugc
xnp/OoNkcnIvvXipEhYWIzJPsSjaez/Uh6SUJPJjdvtfuK92vi3/vK3X8xQNVCj5NuIthkJ9JGQ0
zK/UbppIgXAXbEcyP4z1YiNrXOX9c771yGiHIWd98XQCvMmiY+KBqu8apGTOfy4gpPuNn7lH9P/R
UmcN8EMcgYw8aUrfL8QmUtZCeiOo0GbDCW5REfvyS5VK6KJPVS+IiZfaixchRJcKh48DEU4IA43K
FHXYwscDmkIzijtrq7UEq+bsM8ULYNba1hiRvMaTZxtgqNhbw/wdQt3LjOiblTlQmL108SgMBJZx
TwwFgQgSOwvONNUZHk69BfH1OmqQrWHeHX1M4jcQg2ssY60VzCsP8TBocsmxgojFBMgvcPUwOU7c
YPxfDhWHgAwizg0vq0ffMBiQKL3WgK/ClLNzKkhgzs1Tk0fQGd2pxw8HcD0faHMwpfESEYw2QNHL
tjgPFDh0L5dzLVu0Yz8F6QG8Fxqhi5i6inuoa/FSX7CGgwa0vwpSntugD0l1f4SB4t9hbv0Mg4F1
Si/lB+7tqbZCfR0N2nGZVpr99nJxSpPWJv6e5SJVaey7+R+NdG1k8rnG2GItlXXCzbNf2SnZTWnl
25FtHILcY/9YMYjvYug8an9BVl29b4GEw5ndYz9dTm7eVMiiOu04ijuiZHnr/76yEDGWtJK8vOln
HPOSBZRIbPPt6cB/50oPhLbE53yYADdTda66eXFKdzX7XNk8/1qoqJfIu9nGR/Hut3Zo60ispGQR
miA9JnrLk4d1pbj/rYBNxbwzX14fveIDfzFBq+x695miGl+td+4liVdtkbccjJ9S9tI5bB7FUAR1
dJkGDYLNsPR9Ejc5PLKHanrmR0u3ABFzFZq6IC4//9L1YQbzuzH7dtrYjrTHcED3YuSn7TPj916u
iaPojiIPtLVk2OfDhIQln13TJ2k7ylBQxyBk8pys+bscSNQHlAALu6oQJcp+yNWSha5QPGsI8Lni
9VBfLP3Rn+TaXIl4Q/XD0lbcE29qoRxqTiva6ygRwa7p91LdK45smF3zCe3KeYt6ZJs1Q2VS9MyO
Th69yx1ri3cnw6UcIM68TdTTWzSnVjEUb4jUUnQ6OBPtR4Qt34FwMnSkMo/NgbwznvqR2cACpQSI
Yb8T+4iMWTNYLM9lJZxo32ItNxKTMFzdbnVOzN4hVe1SDWD7piywCbIWZ4fv2/FpbE6wvaN+9bLa
z9iXAaXtVPoMRxVtwEbl4z/esu2PAhJRzjFnttDVhVVeI62vAoFkxLLTmUPUKYlhMgbm8oFg1eOn
YBQg2pQk3FpYYLMIC/pNBPghIsUMAE42uDT8xWAT/3HdOlLN80EFRbBxzjYgawZ11bIaHrdgrpMx
uUunQgi4fEQX9k0NgmRBKfoTt0cckCNuQPpWHmYtTDDAmbuU4m7WRiXhxLSZrSPh9niHCkslup9l
rq54x2maud5E3TU1sNya/VM7zZMJge2nzy+1orlL4AFOd5I0JEt9lhJICG7CGslCsCvkq2OjtYaf
OiLPHVfCJGBU0Gu0xRk11KSp9flR1ZvMT/0Ndrp9kFFGskgatwiSooP0YQPVOC0TGm5+FHS5kUji
Va4iHpyr19okMDBKJLNXwAS8zV9r2vV2A+mPYyeldPsiogxpXbQMFiSZHQgEjAcZBDAcAtKgUZml
GS9fYLswzDYM6q2uwpWy/RijgJ5zQxHKbtIWJDz8c53oNsF/dy/7Y1e6Ag0fhnjRHfM1k5gJLQ3c
cEWPILwD7U1WyUwrQaBZRPnr2fF4RlFLMR8WZDUPHeYRzJm/ro2u/81+AZliWreQ+YOWv9Ekq3/S
efH0K5I9LQWPq7UVgV4k0TRPtGy0FkCQqst+lOlBDcnucCS6GVfp83KG9ewQjKQ4NUCPpK42kgFw
KP0suGabUGHY9pOHbEsVwqy+8i6p5Jc64U/R0rCk7465NdMJvUsXRc52hlTPWVdaZBdw9kMQXd10
HM9goqKUKFQ55/4al2R3a4MntnyBAabqIwV0zSQSa7KsifDG9/iJM54EW0C4a76PiQ6b+MhIRiP8
PaIj70EZNsCQwMbY+AeiJpPIA+cClJXkKszyjQOFVIm1cwsH0dicYXn4gOu8shZBG6XiRH4+cpUa
ZyasBk64wBOAITvrMSYHZc+3tnaVfRQQrqr8BO9mjLwdlrK4t8eA5mB5HgGMid7tZyt5zdHHQPxM
ZNELQNCf9WGjcoVtakBJCDnIGLaP+IjoYbb3yb4rIEwFBhdlbAVchPBXOFeUc0G5SFAwkXDDL9x0
OQosA5twcEQ6C5QjeCiOExlHvpKjS32kDcu3TGHqxop1Ju3RkjGHqN9wBEsonkwGn06fmNrMU3aK
Sz+stur9ZykoISSl7ztb9v2Z/qYOpu38B8HV1iK1RZfS+qEN0c5e7qTbBPPL8bpaM9Nn5OyIO8JE
7wSRr9+CC7G7Vkgf4fcg6WisBEChwcUjSrXt0JesqtQ//NuPeE5X03nTH3S8lRwTMeouNGEGDNdV
aoud8ZpHE4qs17IGbGV1B2q5s4NYNmUPW/dIhNr7lmLsPD77zFoaNwapVOdWkZm+CdFxcMZ40wN2
rujYvAwVDrn0eVauIGUJytBWFzn+Sk9KdVPI2G3XknHmuoiYH98cIG4FcHMujBzHmcies81tuqR0
tlgDbCIzA11P9L5tk0GloQlA1gtkkvJF/pfY3Sdh1tWWmsL2dxBq44dethQp4A09bT/xFoK3X99h
5/dT3yKdmBrmonZ4HW8z/we8Ijdkz3ENm/qIfMjcR9ABIC7G8EEt6nrPk0ZqEWnbJ2IQPa3otfzN
ZD0VY30T1hhnhAyRkD3dr6q+vIGahK8j6xwGW/ABjhflG8d+sTA6UfG5i9xvNG/vSLqYBADKNJzE
fdozk82bi3JxoJTK84IVHyVdjcs0xpFYB7+QxtEmhqukPCRkvW3gme7IibN+TBl6/dVi51s4338O
pyz6ufiQF3jN1JP1QVs1Uzo6RjCRrswFbJDLmhgFcjzRXVliTl0G5x0MqSqH6zhI1C310sTe5ztZ
2FZKXG1NUgUNJXJbCIHul8niDV32Qvzcn3gkMzovsjEyHPuyvgEzOanKrKrYRyZNFua6Q+6H4WSS
Nqe4nk8s8SdjrdnGgWI/FBqmelSkZ8Koc4/8a2qd9jMu24UiJaivYKub5tvOWCAMsBK5GpjKdqwA
amARcALteTlZyI4NzP0z++UGwyvEvwqKmdhoQ9+jJivxRpmDFm/xlCFrZpO5e7lZ0g61hqb4dmf4
GOK6lFqNq3RKOO7xwNBlJL8jm6x38a7bzkoUzyC0yjxwFGehqL5T7J13ac8kawera4YGUuniziri
+IxsMpx1O+IX2sBgvQ085knR7ET/lbDa2ZG5tMLi/4p3XY5mfJe4eaUQKmNkmC6r/wZew9DjvFtM
J0HSXhkyTH23QVYUdYy9QUs8RIpJBj1F38sl5zvNIShvx7WM6ypGKsy3iOGfRRhFXkY6Xta24hHJ
XOzgNCIyoHk0Ixaa8UtHWQ/MkKSYA8cB3ejNWUCIqOVUARIprmKhuO+u/s1PzpL6orLeECLtrMzY
4ysYwoqDR7ZhgtAoxrzlmulzyTjhAch3drSmQ17JA1MQ+Tki/y38I9JjvjFf22JXGRl1IIxx7gbH
dyiGkRvlPC5S7/mTetldACQV5HguDPaQU7QJcbORxhhK4/pM985ET8UH6DQhyYisx2XRB7ya7pmA
x22+fHYalwdbEWc4dKNEWSMJDvkG3SgmWFQxGWuJ9kHZBI42w6I5CgVUZapvuXXaFklO0cR91kIx
3XieZmSbhCMpogqWM8O0BlW3sOQZBMnG3o1NMx0pkzaSnAici8MB9cQTcQJgrNXstJN1nuQ4KttS
6OMKzf5aTFTD3HHFLY1j/0tDy4YsZ8fdmGLSuT/M9WzBviR/nookQD6Twe3rFUH86AJPa/oILdNe
MIyMUeRkbtnQHK3JwPsAClAfWju8H8+gm5IVNxqtmYkbrEl7UAoQI6hEHgjqCcm1ozvEZQ/CoFdw
bmK8ilYRGUsdSI+Z61JhvHO6ZLIrEQalnvsbEv4/PeyK6VVsZP/Y45+JsxoF1zpSAIV3Z0ylbAki
DZSw/47X7FJ8tCz++A0Utjf4Sj1O21movznpX/cKdQkR9axdcy/5AXrHmLqqa37tGidohyHzppHk
mqTj7+V0k+sIB+KdVNFnEOAUnVah+9oGpIDMc4hSlEVfZ/D4Yf7yRxhNvBEKEaJYwfy2/Pork8Uf
dgRIjTZvX4ktR3Lbpw34MlIYLDWxXme5SYAgcSSMFR8n9Rh9pyuZYwEQ6urcw4MxtBDEAEF/lYcb
8n32cqJx0M72XRJcZmSP3mJbu5ZyLdAgqdkhziOajuQR1gwaki42NuMKJ8D8zEE4bmm3nXQdieIB
srw6jipQkGv77ddmDniM/bcgyEy07lC2a1i9h5NT20y4hSRZNJOKXmvAHHfsTa9un48K6icYqzjh
8YTnn/aekV9F6vJp0pAk9ak1iYJ8HS3l3EoOIP1vmIHv2qq4z1aoUNc0dQmvUJxrxQe/lzM8rAS3
lEcoPSS6uBDM0kkTh0W6ZmDmsXpArGTOY7Apz3GwDeyTNUszidemS3WjM36sAa+w26sTNQjM9yBT
rSyxHqh+8WgaahmqPeVHXUUBJntKubSRUswj7YMmhO73B+/7BfH0tce+IE3hJ/EyINCevMesXCbK
t7hZtm3jSc/juiAIny0oaM6o/0uU8EJ6G1kJmDRtDrh58T68pTWE58YzZqDnvqHJEsRkTU0slmeM
R/+zAz7aLuEc7MuB+f7iZZrMLwdLzmvwifgPMwBORzmTBySPxct54b1kKRFOo8aeQzqWjDiBrgUI
Udh3jzAJZyqnuzebmaRGGJZ+clkKxAsSoSRT2QytfYMVRtVYdubChl9ArMWpS5kkgi33Vjw7Ik/j
/t2ULoxgc6zfGsiZ6BqPcuQhejqdBauAqLAKUC0jYlzQbPjvoBGcXzzzr/tAt11Z/wraXa29TAa8
pvP6m+YGkNdSaqjKCVaA3j2puTBj/qiEoZHVpovVgxUX0wjZO3M5oUDHIzi15tftZYAUT1r3VSu4
3o6uwY611iF7ZcwymH+hZgEiHwpaOsrl9WhGCvF3tHYsgDJ48GRYpuzYSA+6SahW9B26h66HUY1E
SsdmjL2j/AnCeRHW9sn1ZpZdyymMxYndGi2Hnxx2acK641Mx/ZLOJ2SJQcBzE8smryrofxkeSz0w
Wnu3ipDQFhHOZEVEWv1bnMiOTREI7d3d7xa+HfTKV3T+agaJ+v899fy6yHqFtJ/hpzAQ7qgWea96
NzaeNJ6RBnBd2quni4/I3ZnnBv2i5hx+Vt7ITH1yA0Z+xfJPWbaAp+ANS9kBcme7oyJSHiC0NOL/
FuTzsu2DhNwOIwVe7fW2A5UEy7Y875jzbg/iuk1eY2hOxUxRkl6f9jLok2T5JXuyUsZkq06vrGcq
PKUCwX3mWp9kA01Yb1YEaQdTJRHUY20ctRTENkJG0hpOP2WdUHJL37rma5n8yirB9G2OjGMBNoeY
gxF+/t/rDfWSErwR+Rq2BHuNDj52WgIeV2iPleh41EDua4VPRzq9jAhix/BYAI8QcEJKXlBYi60i
Aym58CUGahSnPigjOG9fXLxin7h4k/8Iry2F4wUuOGWdCIlkxxH9DcItgPw+XRQlhYQhtvG9bLLm
0C+ZSod+FGOO8TIPZZCuueZxWlZ+4RyQ6gt00JxRWroUugQSgVmWDFjNR8OWjjhGUul2RcG6WaLI
EsdZnOrQ7mh6F59VqVULNLuf515QplLrUirMvEU7PUetI/0er8Qz8SzdhV6hLZIZhH9xEetrONqM
zPHEv82iSHkD4xsKYG5nLWZygIZHa88vpDlRStHed7m513m28PhT9fyUELH+1sOrJnO9Dqq0rLKy
LsY28y56raqKjJhNfN+un2moSckPl0xmFScqhC7rY7ovfdbrB2ZREJB47kLwGiOEw++XR3L2n6ah
BuvT2V/3FGqNvvi2+n6v4nhlJsbgDM1GianYdVILIt4I9z9l/zcP7bp2u+of8XYlv6mW47rJAeHb
IPPvVKcXE7oouVgTZPNPw7Z3VWuvFG5LqDi+5a8sqbmR34yar9BHX8+7e4LiEEUW7SfNFccz5AA1
Az9Hg+1RQnGfJtrN/TYVSjxmf6p1ZQrKkN3JAsCPC2r8LKk1CupqmT7hXVU9uLOKufnGuCpMOB5/
BIlJtyPFoQYmSAPQZW0DJ84KxWWEcJyqpaCmqVvCyZeuS5NzDNWPnamkTbial0dXWb85iFSPHvfl
XGNGv34HNRgi0aRPWfTduO4e+MrY//ElQNT9G4YcVM4ycKrz4mK41Y0VRfqVock8Mh01h+2LBoUK
MFUUnkv/PZM66kM3CpY2OtZQZ4Mws9PBODrV3CKPMgLtEFeN4fdCA9AIqqprMaqeGWyhsvn7fm00
2mpGDGffeDOOOVFXsCvzfiqFNxN4J3FozxVb5HAVJKPxSoQ1ZeQpJ3caLINLJRvN+ZiOGzvJ8XaX
LXZP3s13XeMeHETCrMMg2gUqbR18NqQFF2tOlEEm4HmLSE4mAPqXNc7bvW8F7kw2fQfPjGBk0X2n
9ZYlu+v7KJq+vmOBCwlD+oNP37AyTzoIesEDi333m0rXR6MRLMYSllmeGuoqzqdWWo+YCM0FGSi9
AdFOgEgfa7vpbHkoepTC9lwLuyZrvhCF2ihKcD2bdD1HGcioJ9vnTPNjCNlwaVKuIHJPxbhvne+K
loM+Jd+UF0XttH+PnUP2ZXUGRVWZvj4eGeQ4YTVGvoNGWyArtbPzWkAV0Mu4fjjI5L2orqqwwJzf
Ige3JzbqmG/Ns3wL/QgdKRmhjhKBlpqfUCbwj0GoON+6sytH13pT/BtFzdZeQtD1yfaiwRBE5QbF
OXKz4qlnQE3GDHL2dNIEC93VVlvoA9SDF3slY9eN3O/ck5A2dKEP/SeAHr2KjXk6uycw9QNz9liE
2EfK0XVrbbgtM5WeforWtDQHcDuxSmm6/54xIG3e4/j6GhZgbsajPj8wabPZU56G7nkSik0hbvGM
EVToMv05Jowcmnj+tTPwKLXnWDa5J3D8FVyYqhpn2y7jOPUQiqNcFi5oBoLxgd7SdEANypo6dEcL
B9ecD9k4Mr9YKloOUYRHha0tH/fAC/SQl3OG9Q6PBXicrmoxvX3Oj3AvAgjxvrkFX1gsrCHipgFq
4KSIelMPpVkb4tqBfiaTOi47hS6nNpyTVFOk8BeAV7wnMhWQ1gIaMWVRTTYYyzn1ARYCLl6QSN9g
l9O270G6RDfJPH2H8uFTfgonkgy/bnLi8h2cddOXdGxVhjhii3g8Sc3sxTLg46oML+Dj01I3+t5d
uHrl16KP99mY3pSbRYzKsCt6Hyl+wu3mdZ6HdhyYYVaGqVZ8D/UgeOGV43v07hMaOCkCgRo08N+g
GomCFc5dyTh5BVI9NZJAJe8DuB6mEyMGya+q7YOkvfUoFFzHP/a9lrF1O8iY8WzWkGUaW5ChbccM
dIMhKcmVO4GRUniIw6RJJvhVgQXusvBYBDqm7oNbCQXknz5rJGIYzcEa28lJoZvu0vBdIAZKI3tW
WJ8LfQOHikhGoHsPpHQJ7P3noBmqp1xK0nk9cwvFHbD9IsVmXuPhmw0OmR6OCRmGS6k+9YBWXTQt
YhUrWbASKFw9av2ZxvyqDj2K89Asrbn61Vh/AANTabEv/AMhnID1Eezyu7ZAs2MZqkoQSxmdJpJT
jNOQdMUCZ/KxKixwQ5lpYpYFzVw2lfFbBGczpxOm1BTluGPS+2LLLvgWWX7/10JhBGT1fguSyRd8
o2uPgYfGw6q5QvgzorVOyehjDnXUTJoCvFanJ+Mcynp717AYc1mjcP4Ua2pK/oMx28zEGBWw2b3N
u5H6QqlNJpDoO8rMmo8Y5ohN/H0/hfXetpvvrkW805ji6/oRuOUyS07M5IVK0UNlJn1L4XRAXig/
xrWqipwlO6hi+Hm3sJSx6sHElYDPZ415lfhR5quqwMu/OzsI7Zdn7ZYL3XAnUu3mMuLzVjHTMO79
hrk0s2IbCzWR+LC6kOAcOGl3XFxOKPieNkNQJzw1vySKrIbHgSF++hqtQYsGg6e4MuZkOs/eGphq
jvOWk2l3Ijv7Mk8R0/mSy2Of9qv83hDPGhjomONihXvj3WtPK7w3dkWFOS0F89qeJKSb7PJHoRBa
5y7Mw0KsmhaC+gPC6UxDQSZvljcMt4Z5wGSC+oM1bAfK2PC37m2eke5YsB3w7swHm0k5sJed2ROi
5Xlu1CPZnACRaRJtpFqdM3vLNCEji4gLjYsZ/CpTwhrEgjCvSM3qR5TurWYeasqV4AOp9NJie+EW
mVrUniDxK62jreKIUvOGkvFSNIFKM3ALFqPZIuIY4vKtX47klXheKPGsNB6SDznvKHWMgZGNcULu
xAtS315rEYj32CR9m5bp5zxQtEygzPmVF5xIk/kwsR3IiWqteyCzLkMXHEFO5Mgn6JFtEymswapm
yGu3DlmE1QDjBcaHAl2p/xSg0omSpTUiKorTEY4r5PMHTfILA1sfwvIu7XqmTjTNUzumLJRnNXm8
IKRMQnmYZ5//NTkoZppyxjlmFTl+RnMlxblOjnkuCNc/75yH22k78IdgQWHhyx+bTL3MbaZAdHCy
yIH5W7TXUSBXmtA/yC6P8t+xj+WyuyKPAaZo1jKLCLeBhsAGXXE4J3sA4JY9iLWg1IHp0jYU+VZ2
s4gKe0/CJXwHMBYw6uL8iz0LdUnDGdSqFv9n/h8V5baOHGDwR0rKYMwJedH3aH9ePw4tZDbYmmRd
MnNpGZ5ISd3SuqqbeQdUoghHy34YSiK90+fp9HEMFq09M4mlZts6dCS4HZHdRVO/v8dPNK/i8OAB
+PEy6JdVnvDvGWa6aWMlwbgOhB+ybWqtGdrj8zneB5+1Eu1wU6L0A9vS0/YmBefbEh1Vh66YT2Xy
oj6376OVxIDb2rVXLiuAlMc03qQWUuumR8L1nGUAHtr5vNW8X/Z0Zm6lmKKlyAcpMtrAzRah3xR8
4fzq1oMUau6OXSqAHF3gPzXn/xDlIittXrnsGoTzEMogAmerIcYucaXfSE3DG5dt6RlR4c++UgNX
gONm0vBFR5JdGl2J6odRVPpKFkRhILBidVbxtp6WrXI46KlcvcbT+9MCWyQ33brDDuQzo/pJi3SY
SL35HOtDGm0M0SyCRk4tdZcuu3bDpd9L/Vny8iMS9UQQC5wMlGyBBlttVHE2JvkotFtjkuPyzeeH
bXts6bAKUOCfxxH//DzIuKWhbol1Rzh1gVkVNWGKoENZc1/ekyLMIdmyBzY1KR7nhkFHqnIBsV6g
cT442YWl/NlHnuPcmtYhF87wy7Bhsi0PZCKa14qnRXm9a7bjgFxwdpRYOEmihyL/5yje5oUgE6fn
eG9773utZ/hG8n5H52yNn95ni1EWmmm/Sjr5IPNytEqDvFfIwXSyINv1SfOY+eVRBHS2GeDkAvKE
qjS8z8XM6qGPD0uOmGbxRldOxCQ2/fxd0uRJsVG/WHzp/hg2BiWUvxoMaR9yCgUpC1d1lzSCJ+Y4
8KAj7PfcDTuO1zw40mmvVttQK2PmbDPLYqKGoagHW/q4OK8zE6qHCH/TqXeyV/LXvxhVRjLgZzqI
D2E10igdIundeiWcQj3xjkauMMLO0By7BOjXd5182LhyWz/OJoqdPAB9IuPWb6UeHJfsZdFnI0Is
iT5iyrQul3U3F3zDi9C5M04MWz7iX13SokSdGGq3S40x+5iBYv2AwzMMOnsjwzzGu3t3dP0itpye
h04p2Or1WYfFN6GTy1ShieCrHADct3VH1fa7sjop22xQpB71doE2fkTkwiDO/iiYZc/GW7OuQmab
vOI1myKqIE3WFoWrpGMky0cwC0FWODfK0fv7IwFxCVlyLLIUWvp3paOHPpSmGuDA5cGC2WY9zo1O
5ZJcjdSwtXMtpoXZEHZIBcisPIV0srrWxfhmMt15NPFTZlOQ5hoK3rP673c3ekom1dEXQ6i6frl9
xfbwRzB0JNX48jWMmiqoHQN5xoPboON94eSzg2bQtGsRzhPZsqSQAVHzhvDOYHn6ReW1mdq8SQfL
gzBTkVXV3mtftN7cUCWhEDO56+HXoiWIrFp8KihrdoLlb1hS07xahmfLhOidKDW6UeKxZ4FaA5bU
7w1RvklZdp7+Biexy7eabV7W7Swatj88564sml7TwpUTeAKdGPZ1KnZ2ic6MzIlBiE/DeU+rH/Q1
MOIcgm8jPu+0Lanhs71Ee2f2tOMhqnWu+J3qvFONqaEO/iX/TpUP1P4Mg1YcfHIp88/SyGnUTAe9
U+OH9M7FVvZ68woYI21GUsBJ3yuCn+tlWxX6nXvxVv3NLNnLl+2JAxTgrhQoQ6pPRAbpkYALcebx
t9G65ZkenYQdwa4hw7c9hnnupwUSXmRRSIvNbj9/qhmz+DdCQVL6QgnCd9EZ4OGsumFJ8fyQ2ZBC
ueU/QCeJWxhLCLVsOw8jYychDvaf54V5UEeTVRGpuuWzeIVJ6qdaJQAQy2ET8mva0I8ITTbjoomZ
Q1RF1zUvo3c/rRfNaA5qsVwINH0iBhrAPbc8Bx4inEN+NIar5m3HUIVVG4ShWnGEEbQhwNgun6s6
9bgpIOu/E+p3Ct5GdvKg7iawMQ1gnDZIArobmNIw8GA9MmKk/wOaOoWh4xHoVxYlfo2rwq+4U8cz
w+AElI+YafyX6t5/PAZyFOQ4roA5+fUBPdSymGGyCEZ983o5E0N31HHX1VBcr2U4oxoEbNN7IDka
k2Wc5c7gNXk5hr8dnnAIY9K5sDS9Qr86mW1SFfi/7Gx74pL9US6q8F107Y1O2Nptc5F9Iyl13S8f
0JutcLzLd8jL5u41paYXBDQT4WNcAk+ULYwoakoMMeJjYt1i8A/9qbVvuZsMfOxQSXkDs+q0OF3p
MmzCVsJ1dx5njpNoGgBEgltd/NKddqvVuPPlQMWq6brseIp1EjScy7mHdUceYggJyweMxqdA7W5I
UxwUFhfFKJ2NMv1r64UusrQdIw7QCygnI6ejuKTBXJcl+qTpiSNhnlvXfyCwGx+xHKHXqqLd1NVI
+T4g2hE/4eB8DoGaxL17PrsevfWG/FDiuaNYiE9vO6sFkXjY1MsBKDzX5X8b2xjCNYduM82C/US+
1DQO6Oabr7soWRxkPrdPK5mqqKVSh/2/n8jASk07VbTHJHCw2T2KVPfNZt13jx48Lh9smDaKMAL5
gGIMRD3D73ca6uJIqt9wPzO2avdcC6VJKw+yGkAiHEb7iXqnF13eW99CSxqnZftvk7XmlD+e0YRE
LkCRZGdcCOOJIlwXEOQDdGYW/8DlIJrqxjLQgVEBPpUghto8hWKqrdaQsXfOB35vqzXDvDGOquoa
xIA7ylPVEURWXnIvoRhqQH4BGnv8U69syNoVeCZXI4uiKz4NImMpxOGIsjHrCYVuJ4BadQbcbnde
FqZnNLHha83kH+yjTO3uxd9HRLpJxA8sVSwzkxMO9z/p3wKwBLNhurLXlGRy/nyJ3jKH+Hmsobvs
IkgdQTr2+0uEthKl008I+w36+6xNdaALpOGyss9qWEm4I6335zqUjSnRjXTxSQkxM8/0IWSZlE7x
R5NV1NrJDDYibB5DlOnmKOmR1rphpiacusqbt2QSBJxXnJcBtdpbe6/vpHNVL4nxBRpcbpmlqkpo
s5MnSmg6ir0Vq1vaMXfPhqL6rm90c9lukwyrUpibljlyZMJokoZbEjh4VoyxL5F5AaWCa9MrUF73
VbNNNGe8mk0JJyVRXKKAxgxR8eawZ1EWH5nVXrzg+X5wprN/4SFNEq2CHjXDL7J8xIEd/sWgNYaa
4DNZzm9Q1TJqE2gXrFdO82sIwq6vfQrycFrlH94uPqrsmehAS9QB0RHLh6lwTbQIc5jUmQ+pMiqg
m6FtbNJTs3sXAT2ZcsXCnhIDGcWSm2ltuc9ZCtspUm3HCtlyvvyp1Jg0ZM17of8Qr1HumStfbAY+
4Oa6MVgyF8roUHpAtg+gU/n78NPglRJ9wyDC2lwcrpSY1OMAseJziUtjZ4jc/X84zsAuOVEGKoVs
x2wvMLcQwsuHIDEDM4jZn3kJTXSimFxdsdGHjLgVQm6LJ2kUTO9gsYTSE3EXO/g5rL0k17dA/pn2
GE6ifprIUPmDMNUC4NOXDn47Hahzg6CEs7cC/d36UqGXHB6wGp2O7BZLhhk7zt2olmvrm8xpOrFu
rwdGmIjiTTpTuanfE+QmTRGri1Os5HAVUufoZWwOHrzKh4mq4N0F8KeyCmmNEPFUU8o1D3dK6a2Q
eI60v3/NbjfJchpN4LoC/mQO9h1C84n1LrYUwd9my07wy1LtHpxBrVlWz+XOcppo1H/x2JaYRmX6
xDYJO65Zya1qjDKuW1xciBjTQXQtGNZ5eWtbo92B3JvlV9jhpfHOB+9TDpDPO0pmkFO0mI7Ykl7W
paNw/t7MdPFAXaifotgCTgoXXHw7I6HnkVlFxj3BtIp9zd6PKxZxsMu6y/xng8VXeXv3WKGetxlm
CJI1VVkqP4A+nUEpKnN7JnXFWq/3tmvlm30TJj01xFEx+qrfitr2I40UXI9Sb0pr76avI+u0kW0k
yXCBRv6TENx9n5e9XLiCOPxFwKQw4Hjug0sBW3anaqhoe0o+mHzXEjpkORpOzIZxLi2rdyjuTZJj
4u9TYH9XDTZ4ZW0FpxBiYPrjyXYIvEagb8QVD/MwW6wdBKatvOrCrNulJWxDPDswW+5LgNbrs/fI
MYgsdQGeJ+6yZquWxHXde45IZN9GUldfFtSksq9D0QLtNiwnm2h+ohta4TewKBSLi9X4qhVoF5IL
yP0Mo3Cvt4ke9Pa2WoDHEaGnbcvC0xDP/ljoK8g4VpSrTmr1sodDifit+OIyxx7C6HIc+xIFnhrS
a9tkeY+2Mt3MLW53PJxBDc1vuo7gWlK4M7H9H30ceiluH5aD76Oc5CoWPpbhDtyRaL0rUjThUwGw
HSkrLnm5jVs2NE35idwQqKEFo8tUIV+RFjDcqgkC5y+zJJI/5IAH39ilqtMUCypc3Li5EViv5GrV
XCAYtGYMtdbWVkC4y/2dulirtFit4377J98t0tLL055bnEUk/A38mqpe25uRQFS6cjc8arGHwb1L
8W3lu0ybT2WepqcovlDt9Sp4HRj0EYX9fjx25tBvE9L2l/xee950Hvw/KYo5cn50CSW7ZSO9y5oY
8MT5oQ61IF4U+LZC5xY+ebvGjQoZncJhgApUjKIn3BC1Itso77rqhwZauzMVBwa0DlXPvHIQIUSv
ztIWKx+UjLpeU6JmYcD8GBEqhCKYd+0++LGyHjZGRC5MbJPVQf/KSNfvyVxA/C+Q8XJICzKAGJGo
N3P5ylESzbTeuKC1IeGtA0lnEeryk3ZbNznb5Pv4Ko8f1JEH6bXT2vPTkU9Hszj8Tz8faAqzbd7r
AsdlKFsy6oS2+fjMoQyw9rmK6X9ecT8YZGHfKqS0QVwd+b6pYZmDph91o7uCNXHCuNOiLD3G0rgb
y1cl2Uf/YtCUY/FRTjtaza0ApP5YR48OiGm6aIifraQjaF2vXr5oQ3fZo3DCjKU7uq1Kr+gzSSNF
WrtTyFE/blTeP/bNsM791utfnI+dKvvR9TA78Ghq3uOiXnqPGPFoCy2NQ3l9vX4K5jVAzJFRogEB
R1didGzR7Et6gXgH6E/DVEYOkeJjlq/ji7dobHZx7DfiYEvnWymQRc5+DFmIo0pgLtEzSrMK5H2j
sW7vPQmLdqFYl9A8hWEKGtp/C2BUeWwLiayFNbma2ZiLqpMd3NNjg6mbLB/ZuhzroMjHduMI6tr2
zZsLTtR2jU1IrboDXvB8sxqU9jH5U7+J6VQJmr5f4XExywMqnMEt/jA7a3MBK/UV+1rVEhL8YCHH
+rs129huVsmIgZqKQh4NLoUsml4WAI/I7M3Iw4a1oyGNdKR9+6pOpM+hiIJHN3aTeSNxie580lp0
kDAjm5MCpRAdgTe3Oz0WblAo4YTRM1m7eo2ol21OkC8nhzxdoIMQmxZBO2up9WBfFDMEIYtBki1n
jTauEcyAnz0Vl7jpE5XkBQbq2Tr4tHLwCAWtyeYO8H3t9btQOGDnvOhzpkIws9/q4WE1p4aY8LWr
cOQOD/R1MDNHBzdWKCS+63QJSUCu0/FgLOkkfvyDGHAOH5Y/ORfPwByUwt0VgJtbSXtplVkUysOy
jOFbo32Oa1+XJ5RAogu1RtenFcY7qBpgbAqr45p3+b9edxOfJH3odHxC5bIPx8dC13O5ZtuD1ZtY
JSLSv0cS3PcdVgQyOnz9NBMfsiNefpT11bvMzGNFJgT7IynWSdOxIGfT5kzNeUz8v+YOkOaM0vPh
x5i+6ltf26cY3tb/Tx397eZrbbD9fFSGi6HFgi/XtrTuJDqPvskyTCQQunFwD5lb2vR0vgjj70nE
lq7tS+PKF2yYDjrqdxkFD0JNbw2+ABY+wcVG3WfkMYP4dz4vVM9j/u3ipJ/N77ZNUd6CgGhyzLWJ
k6PRoj338TgD+pt8nD2LEOs8cEKh4fIx48bB3UjBxCtkd/TeHDDZFQfREJmdS9IWBVhYXKiGDLS1
3LsaQmoXFX7kJ7Kzq+w15vOWY3iGDlJiHXE6D9jOtLk6BPBbEE134Q1cj79L2KShF6RbcIlratCJ
BpsKvltAX1pi4vWnpnSbPu4BYC0WzdQwTH5eatoccYRSrC6c6xpU+hcBcoAPbe2nySlSRpQlWgcM
WLfTq4F5vAa26GiXG9HX6TS4lZqecWlOWtCt+aJ8iOGmOm336b9pmass3CB65RMmViq+8ss36GiA
KqdvEKBy/VIadj+jMUlN76p0BokgafVgG4arG+4w7ex07pROYSPC26YhAEOGxBHysx3KKdPBmrAe
AFexNxwL9TTs5PxfSPHeCZrvtz4gNHM6xeui9R7Q1/N1/oj6TTmJEMWuzVW+LWWxBU6z345DFB9J
h8HoEV3uPyBCYnboEaIIR/HN7fQIGJj+pm7qeg2FLRtF//Nw+xEWn+rFCN+5qTYF4Btcx5V/fL4q
rFVGmydMRy4mn93+Kx/hCnV/hplUD+/gxqxM6E0BwnK3mS/B/gJx9/fcocRi8174nAawZrEaj/0Z
9Hf+XGVARIM4N0Ul2hTA0NfwJjySou16+0UYR7x2D/SQnMS9Kqv+OxF7IqZA3puyerEjilzUFAZ3
ITSS3QbK+qrbgZxL7pJVWXsaDhO4EDMTrai10VApAhOWTCJ9tHpTB3lkyh1clDVJAqMpWAmt9F6A
MsrKPLilNNeoU5n5Fh2Hhvs+cwc01SaQw4gUhNDkLsO9VAjonKzVmbQ8ZFdLJ/afbuk3uDrlTYLg
rRL770LAWEJ/1vnC78GgaHdoJSdK1aFnNKhiH8V1UrWYUnBNUKRsffj7AUJ06a+e5mz2pHwTvFdB
QZHCSTI/8B6hV79XFXEFxtzZV8P4HSEUD3db1poGU4c46E6tjpm2rkOJjFbwiyLfDuw0aEmKXfJM
XbbrSQFdVuzD666u59aNi7nbkW1oDW8yyMYH27Jv9SZpdmKZJxVWoaJJON0Snxg8QHiKeHqnGJOj
dHrj8nN5G0HHrPfS/6D3SiBEj42ZjdUmy1Ifwaw43NWA1UfNBYaqD2lDDyCjfvCdy1L//03n7291
PeHLptJQHnGspOz/Fq1bz5GQpQOGQGB9lORIjL7mJfgKPmLn6uTCTW7UV9doer3lxj/WYewPcHeQ
Eo7TtiOBJa6I6/5XN1sVlfpYG/p1nZ2b1+nivH/3cjMEAU0cn6nsoiKzF4VbsXTL2+CLCamdM81f
5P853JycXpFL403Yu7MAKpdnFScQrdrcdnUETzyvhX3Ud5+Uub9nvpp6TDGSd/lgxMu/9fKeN2Kp
KMbolUALW/PZANhZe7CXEjVYoDHFzzZiQgBPd9711VnBIuXlVuFHqlMtzLkTJI6HFr3y4JkVcuUe
dyG3VlmVWkGWeGTdopeFJqjgBDjkfOXZJrmy6jHPY2+pfuua3KZH2seeKsIir+UWTC8VajdTyDMv
gZfDMd/+ajL+KQSskv4B63WReahGZHx3X8dxQfXbVLzYW4J79q3WI0TMaT+amy2nko5n/rHzk8C3
Wlbg18JBO1DXqtk/1FE2goZtbGx6vPnly5BL39Yt7pd4DrUs9cIjudQDQKdkZ4hT+FaAG7h6A06c
4mfn0DhbkxCMAjMSX1B7S+hR2x8UOvXSYhwBBmpwo2G2CJ0+QP5IcxxFKS9HoKOrJiXhT1C7UnpM
NKOD+fWs8ZViNlUrjIMw7AiitQpLffEhUC+1g3Jm+HOYEHWrGBCKm3oWN1KCHl5g3SWh933HjXX7
QeZ/qsi4gK2KM2w/a66m7GZbjfiYY4v7g19Qheh10XAejBG4NuyBXTzeGWr+2iQ0YWk66NhxSTfn
PvPbo5DUl0ATKp69f/MZDynoxMoRYhLg03TZnrNgXfvQNHwJWa1+CwYyXzGZAsKgZM53wG90QXPq
T2KSM9/GrGUnuXfs51Hnk7iN8brG2iUBm5WW+HFNinlDcyefkGQ5ythE7o4/zbBFRe5x3WJ2AhYC
IjfISUT0PJP9sSQBVQqu9QA4Kzqmjmiw6bm4b43+O5dsO4Owe4YwpI+kSdupYa/RiXpWudAFtbWE
wfj53epRnEpAQ4oHXETe6F0kIVaruDS+ZeIW9GLqqMrngZU+8Nt/qDZSYXmvuQW2q0qRTkRdmR2G
9K/ZZTbE4yuMUzSGRQgdRWXX/HGpGTlIW4wH+qpEuXXNVt8gHWpbr1H7RqRNn4cYCDrKm79Jhy2f
I6V2awpgDuVzk1KF9okWzi5NTKjJiWZmu7CJPak0JQTVvRujMrjlKSaOHlRZ0zxGrPRuFcUS62Rl
5lhMcWIINWMYNe5+eDkhsaVPQcvcG3xFRfdv0heNnEVkuuhBN8Iz/KGGBKXH5U7/HJ2GlEuzIWsb
EPa31we+XuHDx4UduxmNQNeM+ghNvaD/G130UFaVssTmnQoffjLwxxKkzQnAwIBGHPSbHMD0lSKF
sWoj+NTQ3MDE2DbRuhz5y5rU6xxW7UZgtApGyCpRmGq0kTKQD7mpjtd72pOo6Z1DXL9OZumpPwut
JWX9//XUgjgJrqRr85CyhPqnlxe/Vfuw0R2BQtwecar8ZgNNpiTFywcBWjl6aC+YAZK41O/GYUR8
gjo2VUDsubgCYnU8ek8pWloxz72WelcMOGRNOvZGG6Z/QXnTCaSrg+OCGfN3H7kBpJPCnA+IvRd6
qo82FAIwnX4eGYMgTVZg6Cc7YL78fxDj0JRVyfJi897hwKc9IMP5zAV4Cjz+gSgyRFDJQpGaKSRm
gX0aIq/klRKProB4cXfHVvGWTZPzcG26wIU+MMPToink2Nci/wz4YkE0a9BOsS18EovB6TCAgKur
YbHhqkREf6vgX4uG9IqOIKmBn6G6xrYluQk0UcB+VHd41SXp4MFIYdW1bY05Hk8+6Cv08cg/J9LB
M/jZr2speYpluB/i3uFsgQ6EzjPjEVjzNIRS/HaA/9w9zRc/kPMMx86ayfAfPSrq2gfOzUc2AMN8
BNf5iYtVf4X6rpXpSvf32hLov7rlwjf6BKbkmUNmec/9mi56aErdVlKPx2jrvqX46pwsjbn2fS5b
CBawZfybo39aQYu75VAoDm9GaOWzjpt1CGRIv4XEtc1IynFFRblD4XQJxDJKFYSbpt+LRjel0Aab
aWoKa3cu7uOcVBfcS9cPFzDHoEKpQG1snnLNOfwGik3gVIJ7nMgY/88vcIpc3jZIhk7PG5lAk0Xx
W4RSfUcqx28OL5bfGn7A/8CdneVsFGXVmPhuNZHn4lZBMY0eWj5jH73XMl/3K24DM/yND8aOlTN2
YshIlqO0GSERAc+4jUd+8qjUSrPtVDihSbRW9PPUi2dpMftG2rl5yLroxPq2yCFDb9alKxtcNlgV
FZD3QHuCQMm77loT2awvk5ASMAT53cdEc7VwCKm2YQVM4o+lvR7V7MH6OQLmy9jyM4YgBptMx0MT
yZ9yeL+ki77SFgZWbV2ZEDMs2Hgddv8DeqKqooX+eA7eNiWPeBLUclLzlahsx0s6nr66XmYgpcVs
9Yr+nr+h7prHkDUxXGmjOuunMcqc7OCBu3HcGXyu4K/QPPtUULIrfhQ33UaD4Fse0acSP0kN08JJ
bgqLZcjhJSE8ztMxigQIDWxCzcX3uP5K6TVdHdYV3RB5VUEGnENeMCmKNCZiyUIBdoG5U5RXLLnq
vf3kzgeXKrItP/LHSmU1qq6qAy3pq65e/qBBtl5zXd9zm+RokyF150kyacn1T2WGAiaErQFW53X2
4URQ98asIWN1+DtOg3GYCVunBaAhAGxY1i9Y2hejhWeE/riFPISBPkqeRVo8FBZNzGoowCg9WYpV
3oKz3gopvjfNynQxQiBbf0n+oAfegVq4t7WWfZtE0URrcaMIht00lK8qcblRP9gfBijRBWtPPceV
M1zyL0ZxJ6hjfyTpIVVOggB0kUVMyValamubxGI8YdueJI9CNXAjllC8/feWauwAx4RPorWQ+No4
3xL+Z7IxTfnUIurPkEXV0cF2A6NS0/Fu4MNu61g007BtREEHycyErRQEqZ+ofD028HOMllzYFfa+
A634I2JQLWBRwnkReJrEq6AT9RNEAiWi2waO0wL5ioVooAviLKwMAIfSlnednnDS4+t0rRg8f0+f
xokNY/7zdxrnpX9ZblKAvGwi6PJgyH62CYs7VzfdvGLtzVWjfyNb9gJcWUlZVDi707DjCdNgHfpH
cMAN1Ebt4kUr1DAqHMfCKMhZkAFy/sFUEovWpLud/Su3pVugwrknSTHcH/MZNIFEvJBsq7idbKRY
ZRzEO+BYpxjP4sdP3EtnsAvA/lQqmUt6SVovbqGDAZRHInHe46hBZy7LVKVHHpD9lNEJlvSP7ypu
j5SFOVE1uHWMb/NeMhJTYCQcmeQr7vbvoXML8mSm3tjcVVAxYbhJWpHynl+3/BJbTYyrNWPp5wZw
eOkRfndwxgCKxe3dEign4UX5BE91qEJvXDMLXT4JXw5cWENLHRdw6MBYxS7wpFIbulZZTwyQGkug
NitdTYhQHI5eq5hhYzeR0JEWxd0Dkybw/PwPf0rufkGW9cHX++IgAkMy1GI2FELYzGHH9UH0Lsqj
ho1J3GWVhChuY+ykgeU9+FYEv6uvy3cwtRjJY25UgEvztdmdwH5N4yAzhR1oKaX1/KqO+ify+6qy
o/TcBm7n/8trg4QDrZucmdWnSo7MCvWTYz+WhmF+mYLr9pOU+ixHIb0WtEiDA1wdncozhC/WpWxs
KvVm9LxIl/iwClnfT6Vp/hIfUwqRZo4Gm4X2iqVkju0Yu52hZBSNASoDqMxRTtEq1IDAZ1A00NJd
/zxnp10xPXnYT1AnGE4JgfJGmWmr72bbU/9Mhc9PlmRZgc+tRyCHfgmloQBG7xpjl3A72DKwSHau
eqlKQ+KphhueY9xbGM43yrQJfF6IT6lWm76ofvCrBt2aNI5C3Ym8uCcPaGK29EY3cA9t+4bVDEvi
1AKT2eraflGEny/qXVSgvpIsEq/mEA6iu29c7ZeMF7lKDfhT8ifboaHu9/HAq3ThbIaAbectBLDz
H6wGXEAD8I8D6d6W+3vy0K0gSNdZO17mJ28TzhC2Rtodpd/I6vOQw3BqWNSNDmaSHSw9yVNmSsly
xsmHS/FEaJFsIMLW/ZgXZg+8pWbBOCN0LJsa/YJjCJtweSbnHxERxC1VX5WSxD+FUVBXkY41RINU
wH4inCLblHe/PYaA/+fTJZbmv7fpkkuIKXRt5sQWjoWzmTrLEdYliwVDXcGRapl94gVe/UNIsG8K
tEv2X4MBqLoY6iIW0PY6vZcjVePoyvkHAumw6ydT+0oOVqTevdxwsmm3Wxw/UyQmxWxUHyK0/Pjj
2gmddof+zGlp5xcERWO+vBZAtaxe/bQDclJRQziY2sf6cZW2caIDMuL3wrM+cKnyv1cV7AI+Rlah
ljizWDkqiZxBK8IOsOZTH2Qcgy0pGeKauNj3cCniJcn2NYlVSlk5WOljU7nr/BXt8QANuPccIWUm
TSQve9Kd35gEanjTYP0eligKsDuHa/5MqLN9FNcGNLd5ccb4s8q0UA5AxjWVnT7aTuv8QjrV2P8O
IKniAUaEMaB3IgZjxYGdfmRXTn3gcmK5GhgdJ5zTARJ2MOocHeoMXM4LPzMlD3I/dixOPRn0MDDM
TuMSsWeU7NzG2qeLXJ9Zgp8YRFol80TA/bgn4fvdavXa/nm5nqbdU2/GviHR68bywnKpMMncYgvO
+ZKCeP/lKmhMz5hVm6o1ALddWyHv3yxoQNP4y491uBV7Xl28QciXdtb3EktrtmSAR/YbjpRHFqD2
R53zl4GzE/5DnJSqZCE8Ml96hMSH1hlm6hlgrBhK0AkwHTI4ERUOZbCjsgvviMjjNsiJxjNfsMKI
61muRiwb61lOK2Bdcg5LvSyxywZoa4sU+hZTSQ1ruxc2DRYqIt32ewHSRk6QAs4zGcgJlRet/hlY
CC4Ej2BdTwkLTocogm65gvR/GRphdxc5+iR3GDGXTJ/nO+BbVe2rk02RVp4Ou1LmKMEShX3HuKvu
F4jjxqtAoeMUDih6L9UTJhCAAHeKnPmOmwJO6PBILkCdJeOerztfyXwTlMXyZkbRTJIwTbwhEzoc
7dRqocJLiahMhsHs/skoNodmbDaXsxwOeZ3Y1NAkZH00TCnSvLicz2cB8c3BljSE5dT0dFdjiztB
2PYs0hpvHdBSKm7G93zOFqZMbQC7nPtGehR7q5ERHmpUmPGTJxDqu8v5pvEAzTXkcKkEKqOUYUTx
fVcD0aiIExH7elWmNpLI+6MGVNsIEafc8Ryyisz+iA5OUT6H7H0Kx44nPSt/eP7/yDSf4HaWZpUz
hst5Hvqk7Kn8kpGsJoK+oJN2F4Ky9M19c+TLUNW5JIrEcZOVFCOPJmaHMnC2aR0/T2Or+2BB2CS4
v0tAPQoYgAJxpAbD06WvQpbg6vsBP3v30ADY4mNoer9knsPco26rSJtHnPO/fgM1TZL44dZpoVrv
0GmaeIGZfiYRH+IZIG/5xoOFNlReXDc/L3F7SHYEM9/JHXHeq4XY663vtEdYu7vPYrHumOO0ZetC
rA6q/jYeMN941hSF9/rsIxQttVYOR9VmVlROSpAXBsgEgtC9ib5CJQ6eX8RqyHxLaHsVuAoupYoS
mQOppFnHKWQ7W7ZNLkx9Ke03PYDR2qX15/5Bwh7lwkEjdUSijN3xsdQOAlR9dXxocEG90D0+uWd8
Q0wZonfiQz0OvuD5pkYKQ8xhdMTohk9Yqa5EtTnOjlVxNgHpCfki9kQLYhaM8LQMZ0uEKCVUZVkc
7xRNAKwNEETeOcmsDFB6y7xm6gs2VPZ0GUTdP+l3hrkjPNzOTwIE55BufQ1OxdNbk614dmpT+NqA
fw1PxrJC5mguuYIS+U2pZo03QIGwv1Hz0d4JXiQCIzxYavgepApH1EPPS68iyDBwkOgd6XWDzIKo
ZpC34MHLptsn+1y1KI5LWfBhHA0AY/jUGH7fHg+3+fNbX9LvFFNVFnCsbRjr3jwfiMl9WcWhBA5y
5FQMgMqgboG8Qa0u7HXLipbUF/CImtJRHwbVXk3VMhzbp1oxfI419b/or5wVs3JT99CCCm9o6cKT
4FMHJoavnmn3QKo5QFLMLoBKMXExky4lRWtE2qeUt+v3sU2O6HsnaqSayyjATnhkeexVD3ljI9Eo
B84+GNViPpXT5b/nAhXB5L6CFPeRbBKMdljYiGuX85xv2ApuPUcH5zCYxH+orB+8iPKpkkpI8HH8
TwG2wpeAfOsFdqdRg8eynlBpZLeg1j1U1KjPZjoMqV4bpLpiN5j0Uzyle8FuDwHfOdSLc28idqMN
waCbuMwJE/6zSHsfTZeN2ZtYgA0kh+qiw25SbYe7MevNNfsVu32ziq19+hnV/MJkwIAGsyFqFrKG
hwqomgTy4kgwJ1X+38gPuBifwHf6377DyP1r4Ux7r8MXnOtKj5t2f81DJyFIcEeBDc1ZRT/6D+FA
Hhkv3IGT/gFoJotRZV5lLPSKGD/jNTw1Q2VBf9U1dYACvsiIW1xF/3ATLMiZmoe+Sg+JNbBJuUi5
fxWu5Z7B8Q1E09uCvPM5fKAzWTXXjRejT+bufhsm+0ucjLEFnRaYTZN57hHqE4/4pObXcrXImVM6
VOSFbnLwRnpAnICMP3bk58d9jRW/KmgRXu8kWZGFKMNRbymZAm2fjgOEqSzOvISIDdSIPMSiqgYJ
gYuT3LniT1xxMK8XO3BSMAiVnmY/H/b5YXMPuaqTRCLgTQcRIPPtytCZpupyTb360OTlgKMFqPG6
NXRjaQT1YnX/j3pnsUEpvDutVlQ+VYTPaNg3BaHUj/hdFrufeUZ53dHPfsm6Xy84XXfDuGxqlr4w
J9gkTWQ93Fw82RXa4tFeucDTUNSZ184ZIBn7+Bao1ya8g3b9NOsJfN52hsE4pn2Vb8xL9jCHfrm4
RP3bo+XaBWxJd3lVeJFcs7rSKmMjX8vcr0OTqBhvkDCm4tIXLxo227saJyJFKnrKfIB+z1x0sUVI
rc22GTj/ylU6EDQh+VQ2K/kL7B3E9W8HmUKgfSlR7U2CigcHIjQ2jbJL66t0rWGGI3UT0IojjrGU
174BfoV7+QJJir2YF6DBO31oP3STQe/L449go60PDJwvfX3tYJWJeC11bYOFq7tQzJmdoded+bp3
RLDMcuk4w1jkYi9vimCYpAFOZKfs6SifzvcSw7B6Fw48BkOf8soVbq+jN/g7XajiBMvknsRO5zIV
Y8bByCOJJDA/zA+sKl21Eg3JyVsB1dWanGaVLrrKm2onGBbfLgF50OUqNBQwnZ5Uym13+t4zh4pY
H7ohvbuUr9yeqpPSqkDYML45gXEGxpouY/7AKfv/xLpvz5+SE3xGRuzb8NGAxS79Ozc8eGThJgNF
svfoJm7uIl3NLTt6aj146QWVA9ydWkQ7ZTiu16dmdxB1LTrH1GMdglIWeatmWuPc/qnKXKvNukDp
2utMT9xAtAE7VT6sYXr/qM8vY6hY9A94CPV3q/54Intsga6w0jRWoEB1Lk4n4kSsLDGuwbVdaa03
fuu8JUxpIKeUtKDVNq326TUhS0k2cs/dF5jRwtu8nW6svIPDhS9a3wnOaTTTZ7kfqOqN6DmhQBC6
vUBuPbyJBrWHBRZ1MJA/wesQOB9GPENzKMn9zaslCl8nVW4tTnsZEAY+Ym69+0xffq2BP19Plq1C
x92Isicg5CP4hgjju399jMaMk4OYIi+MjC6gAj+u1HRzjUQdAX8cZFuaCKQUxL4t8jIqmm44Cyxk
jJbdZpk6c9gUN0qFPC5jncb0Ovg8dGqQNfyMUFqIDSNmNhU8+10/3rPQbXjFO03ty25wgU+T9ckc
Vmn7kZvVHHA7G7QyjrdYqlBr9D5VITG4mNIJ6SijhzabEyDY/2vsZCLYmA/tzMoNfiqgkbPP/HVt
zwP6cFdHign+JQ3eEkQm3CPOqCcnFitV6t0s/n2SdLho6WGGOR6PEggO9C+rUyAycDIlrFWh5Jn/
NkxMP1D/GczEXx0pu4kABoYxkI7FfpnlwFuXAt93tmEhWD7lBxpwA1o1ImDgocfa4/EshPr3EgkF
mHwxemOuZe4Dnhxhjgg9QntUFgyK0CV3CSuhtyF6Wt8WvYlWJt52S12xiRItMBGDbyQQndVf1ZLs
PZFawfyMVgycMSPY2W7FcKmBDXk4CqMArkaUhXN8KdPb6Wu0CLwhRW++YssACMnwhAaCHePX/7/r
8Kk9YLGWAtUwyuX63TbRZEyH0+TlOXNm8gh0DL2Ju1qRaoGBrSFw3wRni6UduDljChZ3It4oG5Rv
/6qNHvF7zC3tB6JIZbCduJHZjLyVekosuTMTErG6SnrCBld9fAl7ewg/T7W5exabo0bM8Boo5HoB
GEVGkGwxCcvWZ4B3FA+cDHOxjbNJ1Is7KlwrlBn3b9sVsZeEDvs6QIYv1UHFaRFFxpullILWev+4
gdjc6IbN3VrLWlS3wz96l/Chez7c1nyKUBFgsl3UCGgG7nPRTNhL77QVWlc4WSFjR51UBu34Pbqi
uMi9sZKwGg+oYv2l4+nWK6Hj1mFoP/UW7BM/YLnhnukloNXQWjg6pIeP4CjjP0DWa1xHBK9Nz4nI
3K59oieDUDquVdEJ977jjV10xGjeKGo5jdIAfKABWyeCFs428TV0051ZLHFMAOBnfb7c8XKb7ooG
oyxaR+HmxXpdNcH/i/MFJYCy2wMXSKMRcZw3L3BY4vS0tcUCBwise99wv3KGv9UVBQ0DgISdYgqv
2ir7IWI6HXZNnM/f/GWjONIuCym3GCgN1bUbjyHF9eHTD04dOd7b42O5YEG+xFGksvPa1ufBJCSK
Fd14NSEKAuw4wdRkNn9OmZkLVacxv6sb53idCiMNx0GDh6z2CwalTpMP4lB5jvI9VroqeGM4SrBT
VaUupJ7aXsupJt/DaiVOGCx0rlJxAvc+AhxJR8Z8tt5LL+M50YhW2iRCtWiaQxwInHyB23UOsmKk
WUzoxGJ2MncoxyOf/FuWmE0+zAyIkVjFxtGaavxNnfeIoWrBQeN82ISzUkjIxUL6rmgbQ3W7reio
TWqqeSeDCBvR3J1QZ+1FZoVuDHbzbUutMMJfaQ51DXvCD0MMXqEhdg==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity divider32s is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  dividend :  in std_logic_vector(31 downto 0);
  divisor :  in std_logic_vector(31 downto 0);
  quotient :  out std_logic_vector(31 downto 0));
end divider32s;
architecture beh of divider32s is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~integer_division.divider32s\
port(
  clk: in std_logic;
  rstn: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  dividend : in std_logic_vector(31 downto 0);
  divisor : in std_logic_vector(31 downto 0);
  quotient : out std_logic_vector(31 downto 0));
end component;
begin
GND_s32: GND
port map (
  G => GND_0);
VCC_s32: VCC
port map (
  V => VCC_0);
GSR_59: GSR
port map (
  GSRI => VCC_0);
integer_division_inst: \~integer_division.divider32s\
port map(
  clk => clk,
  rstn => rstn,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  dividend(31 downto 0) => dividend(31 downto 0),
  divisor(31 downto 0) => divisor(31 downto 0),
  quotient(31 downto 0) => quotient(31 downto 0));
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Wed Feb 14 11:12:16 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPDIV/data/FP_Div.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPDIV/data/FP_Div_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
EFUG+X8nNHSIgjIlzgDQ3j/skN88IcqlJ6BIZrSnfwmzV7CqyrusBOSvt16L3Jw/fR/t2u6LkI1K
7VpHiWQNinnjZcmpns5D+RSyKHs91+dATlxx8nZUz1UEEpM4i0tEVAsrj0i8SP9c3SOhOSWvwqn3
5QNlX2K0XOXlUg29vdKJO/unK4IW+dX3RqEBWceMqiA7i/te4pTQLyldvP0Tkth+Ba5d3b90D+ml
fhZ31mPbor7CO/U3BZB8FF5G2OdYAx8ToEbWrItjdf7KBQ7zbvjSp57SjQ6fY3xdkb7tAqGSPAG+
ZU61o/rkdWdonBxQGaGXc2fV5RuLzGv+ilY7Gg==

`protect encoding=(enctype="base64", line_length=76, bytes=983168)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
hLClCAymVIcrtSJsyDrGJl07sFm53+zd5+XCbzpWvmijE2pqPUx5d61U9LdyvDqyjF/vwntRkiC8
ETUO2LhU3ORouuE6c9SBQNEpHv8oFnr39Xg9Csfac6jRTdfEAw05+vkrw8dr6WFMZTAr5MYlyBQp
qFzRodjd+4AB3gdvxIbtWkGrHZc37RqH9PQT/N3HNcNd6q9fAd97eIBfGeKN7z2n+1DO2SckB+0M
VbbEskATBBJpV3/SP2kpEXsTygk9o2yXjmqkpPufI1dDmvVsmQZCVypevrG4k/WC/9FF5iwidYv6
+sQm1Vl7SXoru/Yh85CxiUDydzG+Xv4yQkZJjwSk2q02nqVXh3jP/gpRkSOgil2PGC0kxef95rmL
pMBn4TAwuGcGIQ7YIkCoDU5pSWSJU+12a/o4cxW1inpmbRbNwZcAO5x9ozeuEAuS7z+eiw02DRKA
X/gBxHThUfn7Rq+Zq3DMKlg5iJv/hQg6q7Jh6gMhFyKbkj54IBtkK5mpDLhyQ7a6xZduaKHJzFDC
pVJQgTLdN1nuvqYBZzcEAYwdfWP7y8Nbe41fYHLsYQX9giG9CaQi3lFI8+ZP319/jTqM+BFv/jRH
b+E0PivzKt7GNVTQYCzi/sDgzI46T5/yso1GhNlsutYayQPvUd7yrcWyMWU4fbW+C9numdtBdIwR
kH6Vca0i0Oh+wc1CL0SmA+rX2WbKmbAQbeqVgJTB//YOmkh4Ri1BuD6KNYcb+OEkHWqkSioKAGgH
DiHPhDNADGv9sKg6KgKm7lMQ4Shq7xve+nq+k+h6hlluwvvhbho7NK3MUvVBPYvXtCZinuxIPRkm
SuTv2+5cQ7UhsfMbfaWiGdgZIwlKN8xMseVZ9QsEIAuLbTEFIEc5r508fgVQaAuUx4d+usO8ad2m
QprCKnH03k427ihr7GOtnHd42l50zfVxru6Qa8umAhr98eyYiKf19T9kbHoRKFBqfMatdX6j2GVZ
a5nLtMq+BLTtW4b/zN8t8FbnviF5/W1k/4LbazrenShR9vtPC9e7JU7DbvNOm3viFrBweu3Zl/Ly
zxrKo1srj8hrHIB3Zrjhnd1/x/gDextUx28EX9sABjbsfdabVKsGX7JPZKOxIRDgw59Ux9Mqmw5F
eMH3fI3bUMeKgiNJmCcb5SQoEVxzI/dvYCJndOATLjOqnMYx5fPXl0FhsNtIzQ69WcAUX6D+rbxo
6rQf9JDNMaKgj+pCZ+8YeaiKv1HBoG8fHPWb+yCIbat4j72rrPRYvTNu3rng1jeKtpscXKs/9j/k
dRP6jnP2IFAm0+eLcjBfdshgxyrz2W+8IfwJ3Z8k5KpKRl5yz0B1BtXgY1t7ye2zLgmH9ZPm0v+N
GFiUBOvcPBdl081a0KxQW4ahxoD//4gP33jPR/ZoseVoF6xwnpTkipUUegMkPSp0YO8qjBx1flDw
N6rB66nWZv29oRmQ0S5MdFq1xazBuzStlHc+Q64wlY3xKFHHoT7fLD8+qDCm5SQbt26xIuAKZlqj
Ct7Ew2M6uUqT1eYgOEW208DR5nad5VLrx5Zmxzdsn/7cr6XpV2DYSPvM0D0H335loNns+mDazNg4
pwMss8eTTuO3p9Mv9pcFFDMxvED4UhPRDPflQ2TydlwJUQFJ5KNeEpFHNgBbGL4MskkwSFg3T5WM
iblBhfXm40ZG1DVXvuq1hc1BMAolcvbwg+P2fVZlLH/irxgXUuGxAo1bWt8V7vUhK9zb5SV/Vxm+
WbUvxjkKBEadty3Sem5ZcGA1xU6AF7yWp86vX242ux9S11zkrzXS9WW5kmDEifHI3aLpdXn91W5K
5tTLFw7LPvLgZ1eIMFhCp0ePogJBNlm5oNhz4NnEdOwI9yXyx+d5Yikxuc2foJxk0XLoShODVsXB
kQNM25TW4klOjIcKQOoSj25KFog2916OSjFf+Z03vHP/hrpKB7iol1kPsuSN3NdTDGaj1GobhmKS
MbcpzyeIm71OfKfwsQhPTDuYRcRiYbxkJSuFkPnQT7g4c5kCcF85s8gVkG0vG+894bbKiYuKRTar
rc1Gs8hxjP1mtJ1G6II5q0HL38t03HPUnsYrtB4y8ecoD8xEvTgE7Lbky3wPog6X4OXQINjHW7+G
qyKEObAq7ewab7UlfmhgjR+GraqyYNOLQFjho9Lg+VHj87Y9Fb3reWwaoj3APqvbPjVlJVOHXXz0
lbkU66R/q6IqYq8TsF5DRirSV/+iw8A3FTVbMO425L59IAozHt5CMLC5y/j8yJvNkWKhLpBMCPnq
BLcP1OYjhxM8MuIZnO2vja+PNkoR7npo07g344OBkBoKE/H0u29BsL2bZv31qzSEVNf9jqwe8plJ
URJ/raWyK2zK1ic5TEtqgNrP31l/kDg9vkoObCd8i/uVQ1hcxdpQUImnS2qOaKq6/nMWzPueJx13
ap1GXRWhcvAyM6Pyws2AVzmyN43XxhkJ/6USsWANXsb7KalOqVCWllGsWQmbtYy8VYYlH4xbGCAB
oZlzXBxXF358xPc7ticIUhqpXYkLpXRdXYFZX3fdig3eNdiU2j7XawebglW9qcmjOPHwWigAm6IG
gbc+Jttbd+yAQul4Nvv5sNEl61rPY0k3dGroX7l/Vjm0z33ZTpiQWZjZ/QjU7PfA4p5af5GM9lNW
6XRGkSaOM7q7/YXeGjfPOJmvKeFYqnAr4UlmzqbWfTu+F9BUExp+mjraICieyD9YY6cAcMfKvmUg
Wf+HoW/kxDP/Tq+7LlIIkEStMnNupYznpiezmXYFY7or8AEOQBxvfKT3GKF81uInBwjVq6XV2znZ
ItF4CqkTcDkYnf/EGAUlM5ujSt4RH1AsotI8CKi6vlBrZTc8nwSPd7Ifg4nCSfPmDMIA/z9CD8R4
zJHkKKQiwuU45TsxBZcincQHRIqsdBvOhUScEtlY636IdWRVelcY+HPpvgGzLeeivOmt9RctVtLr
KQaqDHq9QHPyHRZOLNi30GAlk8uUjkZ2JFItnajwrPiGoMq3jP3KTkfSvc7ahR0oX+42/Y2N4/sb
4bJN3OdLKv3L8yRw8NSoN8ai/In/PwGZkwNe8XKmgEIua0y7waZtvzchL1cnQQht8YB2ZgM5Q6p2
jcAdCHZoEWQa5h7mzTBE1knAG8dJl/ipRDZZu+vWjSqQZhigTzHQ3LzT3vpoQ4qipXduDTgLB/y4
tuVvoe7MIG7HSMSSR+/0yNuAtSD62Eds1roiK8umlIOcLppbzdaUSvextmtg+ggMUvofOoDomnl0
lwwYnZ7ZGUZPVjmmqEZ8Q/Hhh2nYgWocNglvhONI39GSOm4s9Tmi7aXnMgwmmN7PSbrLz2LqHMQF
DbVeBX2BBFcBsTC6GghRc+RWg+ebVKVEE3X71oYFqdhqy0rrxQWM6ifSwxLCV38LbvHTzVEpllEr
Dg36ULXtZTigNve04GX/iU0+fZ45YwyWDsTus2sWIxBTEFVxKGXxBUIQ3Iaq+GN+16oyzOU99yG9
YWxap+nBiud4Y/ml15L32tJprdxTomlsIqR88f36wPNIgeFa3IPt51TBccLwj4aOhT2Vg3Lz+QwP
5R3UnKe8lAOERpnaPKrhMJRnf+24Xgszry+IIpWnGIGHeViL1yY+JeZUerbEZdSNUTIEPpZJ5j5B
ysB5dgJfYQ4BMKwQBtxRRMDTpLZfiD6lkWJnOY5vmZ5B3erN2735zkCjm1UnK4EvQv31pQ0ZJIPH
4zv7dbG5qsZzBIVfgPw7Dq1xOEzsSpHGsU+sjOOGNw0gPejNB/BTz8RXZObjjbS0itN3F3Z/4D3s
3coPTUvLWX3lyPOnVmj2hLQI7GdMu4EeLNjJUwNToRq/pfALCiXTQbhwrTFgPanteD/nCfkrVyHJ
jFKoO50yVUyUGoOrBjbAZFv7JLEkYRsb4OEBBdJOHDp6NRm5og6KSDrhoMAjqUMpCpz4YHZneqNf
ZKdGoikW9JCWAoOcSYiu39ZojSQzr/hLDvAt+DOjwhr9JOLLdjujMQfQQYADlfV6H19d9sare2D5
fSKtVFyoWMhRmGgiYz/Xg+HqiFzLhCYfIO+SB5uMkh7GmLUcISBI4l5Cra43+4nnm57zzK0AZUap
aNY+k30yoX0U6NQMnkmD7CZ/bGfHMEMWIzNLh7aRaERVb4CuAhjv8jBxqU7ZEdNXCUa8F9yYbQ8C
Mwqu0O3DMClcMcuqHLwrdiH8VNHKI0dyU9Saz85ozcgiXGtUq4Uq41zIWS8ti5AW19n500RLyrqC
6ZCY2ZtnazZBZ+voIo37FPwOaGT7/T071Nfn0Zv78WaQS3lns6lrdzqcFzdGjcmpYGR/lyCqSCc1
JfEaoqA7QJ5bnOMyN0OwIvPs3tr7JVFKi+h8la0L9eaS/fVgrufFtWw+9pWnXOTm7WGbMe47RDsM
JlG2tPTxTjpD3aR4FQfAxaIQpQMaThNjfnOJlRqqKzcTXaZD2nsDLc20Ug2SAJf2M4SWlnpjXfDd
HOwmwZYgKO12Z+Kymdd/glTFo9HTXivXMmIeTVWCMKEAEEpy3rBePdZLt9GkQZRPRifB/SpV4qM1
iC4leTMgn/P3jG3OuinBGwtwYO0KyLwta+QdGVB/Nd78vvgH9UxklWo87pNxKPs5OtCjW0Y/sEVW
3iibh8fi82WrwZk7zqA94amnMO2/KtwRrl/UGh9inOxvo6cWDRldXpt5NsqmMN+Z8XKpbYPwBn4i
0OPI2tAdxl4ondAbytnRqPVLXpBZ7GIbTyd1tKY9EZBGO9NDjYzMZqTOUTFNURallepxbM6q2CLc
R4OcPQnvXMRsrDAxiuY97HUuWlHX0FVAcZYjh9CXZpWY7zzeaECMPgnxzynIIaFWWPl4UaHNBI/C
hDP5YRWDmgDkbtSAFgD+Rf8BdVTCkOvIsLbkB2W+sPIQhdp8AeBmuYzpmjbD53nDFhHZXWZy4mJH
csklWC6B0Kwr3FZB9iV5h9AXahYQGR/4bE3pLspt9DgwChpDhOOCbfTBvpCvF9jMXJZnc6e3WI3C
7/ev0FmzSh7HaY+ByG62OFu4PbYCqNRvaj6KX6M2fliVnIr4ih7FzuMagt2299+k8NPQfr835WMZ
6OaBADPhKw90OV3eKDJ8poJoeiLYJcEIWobteWz6nGv/VI921aaQFHRMA8U6HngGGrTiT8Z7ko/3
mvYygZ+ye9LXaNQNhsdGBaOjKDZ95tPX5YE4dhfAJcrbLDghi1jwI53n1NWl8CHPYkguo8Xux5pc
aMMuFpR1NZhTpSUcPIeJAKCkAWts+EewppYPLyBcjZUz28AhZJ0E/PVYCBqEfbbvHV2avTec889e
tWUMR0pjKcORxZ3d3wZeX0JgEIosh8ijTBSSKKQH68Ir/pp3RPIxn4I6UTMpHA0AZJXKxIVdqqm/
vluJp/Ghkr+PhWY3y7+mOwWtzZw9xtVy43IIfGAjQ6kC0AOlZk4oBDaIml1Ec3COOOtsvbelIcBY
/INSCpx+KB0EkrgvR1nmwuAlJURxvp7oaIHg/XkiWIJdKRDAcEgWp6/j3K3e/AjTA83WheNc2ZBQ
eQHl5Q8BOjH9b+wLopesHnd0KNyA2lyOYdV74CwbOLe0sx9MkPIXFtcAi5HyBu+MwXZ6KSJcijju
KiPCeUlyQR+gyDvVcK/GPTH/w/en12jfrtcLzbo/FOk4eKDXzsrHe39npldkRV2YSuNdWkNhLJzm
bJRBSi9W+s1kYxfsuSIdXpPqKr+SkSwFnFvbec4hwE2TmDrqfTFTIU0C+MAe31UcNUnqSFHPG5Pg
aLtEk9FGC/ZRgYUEmez7ZitXIHSQmTerw0uD+hxdO3FjpTZNNxkmsolgqsbgkScozkssQRNnLXL3
HcGLsHoEM8mDLjnuzO8WN8FQdgzXa9e9ouE6hfgv9wTMVEEZ0plGO5owq8boG8zyfavbU1VEHdrV
HYa0llAoJKPsMdNnKc2ugXN9jl53eGMriHYYi9oE9hn+UCfwlCvhvb+kt6GYLjPCA0C4TiP9Gfwm
ZiWc5DyN0s2mTPtP1jxZCCTA1aVgOvwpVQ9A20H+4Uxc+9QxiMSTWCbdH9O+jx5Si6wKnZEe18vU
jFQEsl53lKea+PSoq6AmH1B64ozwdmvznmRAqdKNueG63lka0bgWawD4SyYIBfpLT5NR5RVrEx1z
C7UQLvgDkP3hTe75couQ0J4/2BkvDRC9aH9YRGmdjxtKK10nYOsUSx7do2jRRL1s7tcPKZk1M8H1
UPUG4U1iEjpxJMnAfgfA8EdyWRBPz0Nn2ryufh/syxt59RGVdw3aXnvMFrzgm4n7c7g0uQwBxY8r
8AP4ya2Z1xMsY6nfKsVkMw1QhDbwSqfB0+GriZsw65vIXMuMzbttqkZFqRersWFvh6J0mmBeqx35
SMUzInnPQVWaDQQT2XS6WKKZImgJL206kaa+bpO1kJttIgVSNa+DtPIxSKjL/GH0se7PTsYFd3I8
pPWkrSM3JBe20KL7VggFjVGcEWOQt2V9/rLo67GU53XpYq9P8Fa1G41i+l7EOWJTapfOTwoatK8x
KTimlp9CbGsVi7XCP9li1w4LyjoYx2akZBD1nVFMa8YKjeLXtEDocwBylzojpmx3J8YFQT5TJ9dZ
jFBaoUwfnreOztcZlIeFuDV94/Q7YwsZor2aqHhRNBvgffxK7p6STeWR+a3JXxL9DmJfwQPQbjBF
mTI4VqjmqcO5YrGtftHH+eWPOJLDE1B4+5IfAYV0KSDCeZFoRC6lcWMyjwUy2dIGlFfHr4e6Fdyy
i3fKkB8uKcp0pWl67qt+HdlnfmGt7kqfJ5FwjUOdC/NPlmk0b7qbd4VVMP8AqWnCAQZZ8sz+oBCC
yDH8ONtcS/iCQH50Ja4L18inebsJBkniFJ28yTlBqyBrG7rp/FsZqCBpcCOIRx2LYcOVhQ8Guow1
kpjLp6zB45JdBbayK3PwTuGItC1affMj/Vxmk0JmDXdAFZ2i7yFSnkXEMEhKA0OFnTWo6eDNrkwc
8iYeEIYN0gcGZjK7UFl05dw/mph1aoelHwBgWNIJC0BuUNlAwXroIGQlsQ7yT09HRQ4aYNOXld+c
o/7a85oIgG6oD9YCLM+48VWbGqpyA5k+oLESsXnUBp4BfAh4C1a8etM1lC6Ao7Oqr4q4yzsDR3Fd
m96QEFWx2xjiRFUFpdeKgWG8ifAmdjjtdiZukVR7DcecyAlgg3ae4cp2IhqtGakw05kdTJObA0uO
6kom4YT4IhHpA74AGhBNIRWfv+Bxts22jiSx/mrBFmcteROHrR4BDUxC1Hl66aZEqNsNGTW3NFO3
sAmHPvaPgDc827Adi2Il1La4yci+fYJKunG8eiPYdzxtuMQSUQ6gAO3lNfr1E/HG6bIiXEcQqbUv
xl9esXJZs+xAiG8DHrhSNU76kVrLXOCTfqW5M1nIzFrKolw32n0oKwfnoohfMRxyavp91GV+B0ra
1eu5sxqanDDZJVrsUOiRGFg7WUihhyJdEgFQFxK9InWA8Jv1Hlip+LA9tQGsBA2YOCi+cBa5cXMX
KWqRXbeMIcvuOK2OZlxDMLzbS8RyhDS7/effyZP6ql4RjH3ZMT0WRxZ2f5xScJBw9zlbA0QXAk1a
OSxTLEAjMtoDmPksT4h3nbtTI4RxCoMyYWj0s8QN3CUIgAZzCiwKXR4FOwjIQvSTUkisDCfCJEPv
bVNjQeBfcyebzM6aisIWSe3a3aeN7nQmqRTOKAfZTWUIU9EUZ8XVxB/La2b7pfMZxnJlj28fOtEr
yo07RxJ2i8bA201XaWXllrgncgS1W29PTcERK+JQEQfh//WsRnB+WdRqQYswLDTBex9TT/PFtSBZ
lQ0RVeFw0EP7PAX2XGr/xi7WkLz5JhjxiPBHFfPnQxqWYUlnef2c+TXg6ZbcwioOQgjhhCR0J6zp
TfST7lH++ig/Co8w2FdDYG7qGl4Vv1iY8lHsd3Surp9c3QC6mpjHT06WsjWroPHmaYb19yV9nAXy
I2kc0HGg8YIAsGpzjOVQ74eqTeKwgT+uSXZj/7cA1IrV591PG1hLLsNdswpdtkV0poyNF3NnfoJT
xAFsDmaW8TIi+PB2YNpNAbbOcV+y1TvXiW++X+cljSoqSrBbjmTCD4OjZwzdWwWFdtwFRiWKtsqG
NsISPNu6D8vl/PluvpmPEhYdSZ+thVZyPA8vPe/0bmd1K1A6wUUeqHnxABYi697ezC5uhwIQkBUP
m+FZiv4OlKjRSDInserHMAY6QEcm2PNakhyCmghBkaJLy3qvQqDTVJkdbcMnIXYkq1yAyseQ+iAJ
Kn4+LZVegIM4BV2Fdur884V9NlpthBy8dYxnTEMW3utBRbypvhFlBv0fuJghKNgc7F5Xc5TcDV2n
gvwYY7YV7fw2OvSgBUW20JD9zewN1/eAYXFGCdA0zfi5mtmYgVrTqe+dSRne8/gz2SS9Y4rjPkVQ
2+rZ93mepTsU9FCP0RSQ4UXAgJ6efzFTYAP87QGRFmH6ADxyg9PTW+77PyN4HaayVUiHoSSqsfG7
Ba0C8g/xUQoHkO8z6RgHgJrJrtw41r+qpBvbVMXwwT/QTvoBpWX7btDeDlEPi7Z5lhs/eIzoWLhq
PnsHCTke0prpooymWBnyaa2l6LBucuxycw78lYQWG0GhBu9SxmLzWTUmkm4KL32Vb3TaywHc1sTo
r5niS/J6macP4RIY22UgyvJ31t0503TGiimuvEUU2tf79wMC6DZ1i1zd+wsIGbIlo1UMvp1+nyXd
LUJnKzyEIanLMGt3UF0p/f4Jjhf1h0kI2E1qzb7tiYve7waa4X3r+haEABC53UBhkADGTtD22Yl/
qblZIg5H6pjrdkixisCI1WVyuoxpHuyjZre/MLs7c2ULd6dlZh7EYOMz1IZd5d+Z/5cy6V9Nk3G7
s7wWfJDVL+qLto2FMiv/SPxUaHzf59m4iSbGWqMeKuCSVpQAkmT/qg81KiqsWdKGTM6inGvjWBXE
sKz1F/AGfmrKoG4EdEzpCrkT0OTiwrzdEzf1+2JYJP/7T+Tkxdhyo2BIq6JO7O/bemiFPnmrbNoD
CJjZGyv8MEhF1YeSqKL1TBb5t4arqbc5v/HvBYptqBZXqgBEJRH7OTlEOK0Re/ymvQUZ9NjBohrn
7dS+s6FWXH4eHBO6sm2HVjymTf66ay8s8eeOQfGguexfH07IfTv/BtpRurG/DuMrT+0DyxXLIksb
Pk8jAMVl1EVdO7Jzua8+RZ2/Q1W2jn/sR5g0RCkEaHEAeo4zsqcDSD+akDkZEyeEYb+tuuCjHeXJ
4lNFdL0RVoTly0U+z2Yl/SLgdPsHpNU2iJnp32zlJHKbObS2ouq+02SEYhgPshVV+Q+eFdZ3N08C
5FvoMI+++uE2LTv6zKOy3QGj5k+4C5iPEldsgteQcAxMdl5iKxjjEcinnTw0u0tGx87nwJH3nkYM
KJJMlFWUQWhEvHavX1wJ4nV3TKd1u0FmJxKMWSsmf/vivVHzo+vlQyEKfcfRvsDgyrOXHQ8ylvpd
T9ZHsG8MmjXGOxCPVQZgaiXQ3WNxm/wKtTK1wSn9IUBI22DqAsgMAV9p89pHEsNTE3LfBVUQdcM9
6vJavsLX6ldOMOo8qB1YbVJUgTYg19Ndpm/PUygdSyK4RKTk16pfOUxXv0jwna8BOzuO3l8Nxuyy
31LUuDtMP6254a2r42jphl885BGhuwrSc4fXufVPW75jj1bGgTbPHqfrRgpleS9KChYB6/f493IZ
d8YkZbEZK3lIP/9AoyI+5by4Wmj5U1b4VCiQYqYHX/MCe345Udm2BYssZcmBISe64YjEi63fXDHB
zMu+lwbM/BTS19hnUzdSU/F10MlQwKv3EkDAsFdS9q3063CErZDCrI4O/Q0ZnpiBgC26zT0j1YSM
NWPGuKsf9xbFmfu46aKryq1BOiit5SOYKvO0J8PYZxbsfvwegZGQdRvT1HdnIM27bsm13+vlflab
B+9P1TKuK1Zac+8wSvwnieecQjWhymmsVjEDvhcyjjBHCDur8ESBQ5Lff+hHSoYdMCvB6WRCLsic
RucOqBPT42xH6vS21fFMGIhTChVDWyu7ChVWbro4ESumkZ7N9Gew9dZlpW+UNMJ4g+UJI2AMxaUX
FYb+W69rw9qxWyCyjazw6DLBI211XFz+ieAdfQT6yrNC71RRnKy82L58UlJzy/Z9Qj+sSXQ/Dk1j
2xoz6JDQ+d/u5JmPYACtwObj/7a/HsswzQCuQ8TYK2XJrTI2zWs2kvtinXyB92UFREdy/B1Ol0tN
ImOiLok82UWZCTR42hKmzsT1NPDm33S4haqbhsfhn61efj/m4rz2Sg2cpwvJsrCdTNUboTnu+z4u
G1Cc7ebozlndteMfe/GOJB5XtdPZqnB5SB9hsTeUAOgQCrroFpbJEDS/jcWHmPsr1JSxWtwi8Atg
9pegGz6l67x1zUBAEibGZk0h1DKl8FHdLz0q5Pc/YrJuPUbC/a6HlcEyXCAYuRMudv2jmqLgq5eg
dwWgomnYGEfU/QR2eAGEmHiIMhlUqCmho3+ER2Kz7unWPzxTm6/XYw+BIIazz9jf4YR2xl6KzL4n
eF4bsHkmAcxLR9cfmlvYVsKMcWMmSI9/zgMJXk0m/J7q0AxD5D+Y/9s4Jfwtw2oUt/Sl/xsf4rWd
9UFom4CSNVdgSgoTOmBXuLF/l9BepewiaByqmE+PbS/F2IDEBBwEW1PoD9H80ztsVr8fcgtElL1O
KC8VlpQVdmguugR9a4bfo8K/BaMtIrWSQEyySD398hAcjqqyPvpyubBCwbjXwQ3NkShhc6zAW0+T
alyOVe5Op1Wq85QiNOlfX/XmHzwufqQWAM1rDOsqRo3WloeayYmSuf13lbF8iMbHAFObdk/BHWZb
TQkMTkeWMRBBViAXihPAnrvE/6geKNLwGgcIU4i9hyb2lixjx0lnUo+KjtO+QKNI88xkxgd4FKHV
WrTUm+EnXLHtUaATSf3asFFpphNOBCtA6blnUaqg3X9LJZoKD3WSkXYVBscBv0U2joHfFmAbErfU
bJPGKfwO1Xl7K/QQ6NDo/ia73QWTGdRsEjCZfflU4FWOtAUc/VVJNB6nPc4+Tj6xyXyT9FCg9KwA
5BrRvviJJwtPEFiqBGmihYuKfxK1nXo6sCXKh93CaIytYhsTPILzyxPQIZUbuK39w7DH3TW5YdWq
vjCt3RIBaBGhUV8PQ/Z2yuwGjRJJeEicVDtFPxWEBgJCBoOetqaeTv/3Up8n8WDR83+oY05FMCaT
yvLKEv8QKnb70rBTWUn3fe7goE/oJZmvkO5TGotDpxRzzJkOKt1Ur9NjwRiiTg2OIshLEVAgdYHc
JpfVFwMDCvlisINNQ333ycxnyAKlhQ9rL5pHhl7pfyjq9byoJROAxINN7jrFes72hwxqR8oT94p4
rvYz2fmSKaHcBWXd7vhbGz641yFq6qceEBydqJKQVtfiQUNZ50X52LQVTsoOd5/+MbRATfE3FJgK
Bm7v//g8mTF6w5pbgtg72cH79kIz+Pkvw46AvFn/X9WMlm+0JjvGgNWuUEwXocHhCQWngWyRHRP9
Ds45NFFA8UoR2eSU5t0sX81muDuFYbRqfdqdtl6kEix7e7tX4wO83ODGyF+qUgn9lYOG4sGvV+4J
UCqmgt3qXGcjW6CyeF00FVPZpCFuAjrB59UrqVlgX27hi9I7JJMrc7LjE3CbeqUmsM3uH2BUTzIn
QjUEV0cMPLnKkr1pGpUjNgbYYuiROxQbcbN84Kg+GCyyYZCDF0+O6LCIKBrK96Jg6joHUZ4ns+IO
ObHGDo7G4RRiNKnG/SVeEBjvAjr2I4TGiCPX8W5CpZHZr0qpFYkLJm3T98ndHtHff0aT2Y3aKK7I
deIiWlO1mZ/TC0rljpyH/+mma1j0H2TcMPcRiahk2xzQuAbDhg8Hxs4Ulg9cFXurWtVDqoHNW+wy
+tiaYo/YR6cUfhTcX2ACUg9p2EpuM/Js4JIAtCh7UAfqdlbPenHsSMYnpBxPIWnM1I6cj+MWwv0T
pynBfMH8pZOBe8Sv70XNDQ/X0cZXsfjzQAkPRDCSDfDTHn+WY73byCNPhBei1AXqsBv8V/UhOlNV
xjyjbW6fzsG2enpCjk4K5A+Uxu4gNl3NSVtXNolTXB32OBo/O7MYcMrZw+DRFOHx9GtTWxPASUq0
/cw4sqNRUqJHoUSEFaOHeTs2Ddhq5Ss0/Mt5ac2OF2n7kyJRrt1156S24V3mgPnj1m5W32Gq82k5
OW/LtoVun8L/CepElkVAPwvkke5zNQUvexQLkOw7UDJpUHdeBcXnf6onne6QUA7cEGqJwvsTpjWK
b1yfSXIr0ueghTaGZsLL7h/osi1wrxm23gIRud2xFDMFVfxd1YUl3XJxpkIf+uhFmJM7LFu43bFX
S+uvUm4FCLAHKEHC9pKh5R5x8//2gBrbIDhsz5EB29dmAhtip43ze97imSHRo7fj5mNTpWMQ74cx
J4eIuHIxt+vcwaP72DwIOLEGa13abRZcMc+V30UFwYlD96bibZCZlVF0nBA6GgO5bfe0YI0D+gGm
+82+Dm2Q2cKS0rX0ay9SQazFo/HFFRIBHH/bMzA0T7YvDrctHGhRZTkVPaNj/GDvwDNbSIZakKsR
4JR5t6QH/JWeWR4K/oV62BQzMknURoSngMFKzVu1gfhS1yjLG4h7q0GX/4NEVFZKRAahCF8sxITN
jVKIfq2bLQFFFE86MuvTr9nQiNx+U4dMCwS8KTJfGbzzNybcjquaaLzqcAGgBQE23/j2jCvUrA/C
F/+Vb0h9IYihNxlu3CcBEJhOm+8tuA4bDyg6NpmpXsS1BkBip9sndU3O3Ufk5mkisll3Co+qeBL7
GYoInXCQFu9dInreek5THEO7lT1B6tYedjtce0q87n03ubZfg3wNdr7XZVK0Lflr1zkFWY1RUzIz
xnZhisYr1B/s+uzFKU5F5xDDg5dNrN8n/3kOTQpaqJtldC+idUawe4mEF6+pR+ftT4IVRnfL+HUW
d7dasWzTmDM4lkmyNN/p4vF9KYxniY0xL790cF1JGRyKOwPHKXNvEEAaj05x0O/hiX15hjpSGH4P
i9qk81lo+fhqw99T+XLmvMzNDcbmPd3IhfDFsUce6lwjQhxs7AQhN0nYE1xQ+LQKDr9xs7O+yONg
6zdysq53tJf3NA9uYc2M9DRAQZbeVg6mt6g+Yn4A3JppqTTthioe7X+faWF62ItFcntl1CrnFkY5
P0reBow5TCSFsJP1kDn+60xToe+GRS54WrPllzjTldCiAmHJdeljF7eWNEpSJY599nuwCtynlDlc
TBZhykWuOBBkX6fl9BVlx2AGG2qqvLK7ldWj11zk4yNdkxy0I/NDQa6TuM6URFpe3qs5jGE6o0It
tBQdgHdZH7ke5z0PIpfDJYudbIL70h4zvdiKWgE4NjnHpkS2zeL9XLjbNJOAuKCbTVwIgOcJ3mfX
+d36iCqzk6HEm2JDzA3kZlIW6D6U63aBOUm5eEzcSHxPPQmS8k/AVZmd2CYMAJywwSJD0ad5MGIS
dygVEBEQvuSFN9JFYfI9ySWIf8Fev0QS/VZnkx+hMOK4wKLaqO9NmeWD8RpWBiJpGC5GUaIZMicU
bfrcCT3Ak2LBO/1cMqcPyEjIbnTEVXG5O2t80zMbxBK3kAzgn6L4Y3QPe6S5tli47lYLZVKShcwl
hyvX4sWhC4vKJNhQ3Y2CeVWnABbtMndi3HBQgoYR/VSKVIm//2q3ZpTjEazf5T+lYSwgHSopOkYo
ZGyK8cuFwJCXHSOwOoz9J0/TbdPbLRs7BDcwmOhWyerJnGHZwa9fdC+S3P4JUCTKdKUBeJHEzNzD
jW+v+d9hUXtxTJImG738Gv3Qd243Jz2RVEMjhjOGCSpkefJdNOMUe8e23SDo0vkaEXXh3e8aMNAu
ptXIHCVidlIQis6we/eiD4bo7j4fxovmn7pgfTVcglliOzXZpZe1liEPyTiAPxgKCtejP9iIfvHw
9QXRztQj6PTMD1JZFQKZR76nTwTGX7aYZIEsN5cf5RmEO2WzMnB0UbCRQcvzzzgzlgCghzSjqSz2
4jSPIx8v9LURwZzTf3YPonY+May3l3SHZ6sCBKzsb8RiRWy7Qq5Cxn2qr65dDJNhRNdKvgiKiSCa
oDQZ8Gcw0Mcbobzq4b4UJOgJMG8b2xPCKYovhpdlKwc82Ccvxoz5OZO976RsAXK/+EpfRC1GeDab
pk1AVnxyR8WNbAvU1xtHXAILJQdFGVIdaVWf5VSnKAkZYK4pJrjFuQ8vT8X+aLqjIG9qQNzlf+oJ
1R24Tk6fNaDsiBF2OKddwysdH+xtzRvB+kagXHSN7HydZYnkmmYsai/ACnpaC/FuLvHAZQ/qrgHt
M65Cf5hWHqU9r8+wdWbiSEkn+aYV+/CYqoHVRFC1TScMBudlXGnYnnI+zljsU5eeVmEqrATeTMLJ
g5+Eeg9NRDCUsM0HDIczdYOAnl/xcS5pGORRRu4tGHlrq/RIRhfUX/Dlu9tgw9SBUG1AlPPWhYRT
wxnelzco1CWaWrlMybZ7b+xNmKaQ4TNiJLwsGQfK8GpLGdCO1WMLAH25BV+pssKT8821v6ZkkF+e
NQrYKCwDICQ5kcMcwNn5dnNAUiJncmmilinir5zs8Kc93Q5ZFkgaXo1QJP/AjUVksGoxoAOKjouf
caPa2oduF4Hw/cWvxG+SasjvuBR8PPhcdim0UEnVt2xPSzqm7bDuf28GrEtCCypMq6+HfUW0D6cm
C4VMa1GlYFGev3S3f8zlGC5akDdccahwzUF3F/oP9HGH4KcopJWotBM9SVM8g9JpGtUDRHs0/uBA
VII1EK4Qsti2Ak0RPumdUTiV9p6gINNLe1NS8obNQRzTqEGIo8rza5wY3MiAt/FptHIk2eJJcToE
6NJOyIOaYgdRZnzjHftQkgYVUoPS3NEDBKJYWaqISSXjdGrpcJwbLYWgXLxK7ZlPJPaGZ5w5dVo7
23VZSWdicsKNdsBv4MBIyojC02SuJeM9NQUxu4RMz3sH/NHSmNmRu3WGlAPJpE9WRorSTRaqIe/l
w8KZeibxoLemXmDbJw34zhihDo3Gb/fEbTpDxE2i3QG92Ult0JgWpCtqIbvDosU9hivqXgrbqhWR
2/+MjDidJoF6ZP6NAoPl4SuT0tm+HCjGazvwRBqPopXrtmwvFoSDCaIEPNmO4mycivdK0zYz6cpt
SMzRxl2oylZvlxgHeaI1mFbHYSLSZ+ehYLM9CrAgZuYRQ/GkI9LWfj41JuIMYu5hNSrVQQLtk5yZ
8QM+X4rUY9b1IAnS0vcqplhGsQTjNbTwkjORyINsrVg0wxt74Z9SZfPm8udbf0mqi5RA2I3qkSD+
iKPfh3KVnU8eWa6B58nrRJSKDAryJ+IcOGDqh5x6oKcqvbupxVKEcz50v/RTxWnPwDr6qTmJN+/H
A+xobyiGrOecUA+ThESO7hS4urnO7BR0CuVGdH4JInO4miiviIw/Z6al3tfRybESZM6j+jbDB3CU
KYs84enIaAF3P/3H0C4kWABn/M++tHlSvP0l5S2Z/2WmCOSfMM0MhgGWrAD1vrP0yvOdembr8Erw
XZsPvyxf/kZBLen3BmQkSrC6v6+XBD9QCn9Nk+XbKvdC/Tsp1td6I/1TNbnx/tmB6eBhT8gSpYt8
Yab2bXY0Se/A9qY+VPDw91k+tJleyykUAdMrXytaLmS3Mk7BVb7ghU2sgfsuT1ZH+z+pxnp4Wcib
VL2LpZ2G2lB6x/kYHF1RRnVW9HJDxfbgRUW8cRPiOIFYrkvTCnCipIzCFV2UClAHLUZFFbkGnQMM
nS44Ah4wSZmH75Qz0Sfed3y5ULPBzcDnbctQkTAJbijgY3cPAAeZ86ACmg7Ms9eR3zri3euWURE+
FVF5J01j4KDfGQN1l9RplP2eRUTuoSaUk5FYU7Lu2SmBonGjfZvnGsSR8Cv8dqFKw/ZQhazbA49o
ApX6HU+mGT1DgOeCLXcImhRHmUocfDm9Rlm0ZYDYl6Fhkm6zSv84374smRoar8UYisAh6ykULlr1
XTlJ57jLyh+ZYNl+ir1LrHPgxutGT5KekogyLWaAcrLoOYJPqB6l6NPdLxwJraUGy/oLAwhRsp6J
wtgcZinnJ1Gz8l9KJInAjpVZ7thKxDM6Cd0O+u7Q8v9ysuMtwdNFW6RugTAaC9VWCAAMtJJFGa9z
qgbjYQuswypblS4gIQx+Z92rimZFz0H7z//bI87uUGFN3A22uN/X64ziNnHB0Ec1MYp2aVMWwDrr
LObwHvtEjJT2SfEbDPiGt8OG3S/S/wOYEENmr4qEuUFWS1FyJxSxFl2fK2mTtGGv4gtEXd12pP6G
P6bE21oofHlbHQthMlTDmQ/qrnKMWRlp9grvjHr1sPuL4QTdtQve5rMMVkdgXPVuUyKWDHaolP2N
Qufdl6d3hgVfYoozo14rAZIiBP85WBW58R0zcbXCv6jLbCuUpR+hJk2oSw2ySvUWZHFcEk/V+xMA
fAcjr9SQ9xaFjxU3OhlTJDK0PRTrQ0TuTHMqAGsiVeyA6EKuQxKdfc1O7zAiwoGeTlXvQ37YEDMz
yrBovHaYL2lOOyENyxHtVTZUJOIb2HFyARit1AM/4logdX9ZO3pRbUfgBMwVZBExZ9JgZ/A6D03M
agcWC7EUQgqAbFDJFRHPPT+dN827y17aufheBPf7OdkWM3j7/p1lMcw8Z/9o5IFdG9xtC5s+01l9
FBG6J/BRJBTvbA/jPV2xMVk71KO0x6iN/MCvr3FpevX3DdrDZtzXZ0B3YF8eW7L92V+4e3MkOxoB
g/7RuS3pSPJUFz8/L3nAd1TwvR6BGaDHCk0cuvWjfZ0PsDgV/ro7EUAMJOecYBhuO75eoDhuWDa7
BOjYlY3R8k76yoYBpKPo9daevbUDQwmW+R1p9aoRsXims10AxFtO1ppJok10lHEi9Fka982UMQj6
b/60VL/p/p61WUlHRNWYnylxIwEhg0nZ8ZdLde9NlwIlCqe6ne2SLzUaIqdVyWHoHAWDe1o4LEmT
BjR7TYoWk43bKPG58PAl8aqooRzHgV3R1JlY57wEozTPmqBmpQbCwQ1CGA4SEWUX1H4pOTJKqyVR
ZxrqVhLlefAKhUDoR9RFWgYKxomFzo6o1iCSnxVlTzLSa852P1gy03m3WBun+xMM0qLdFMyAwYP5
6fua4+XBC8H3tofqisiXhvAU47Gxg56bAJ/d8zoaEbzzdKzlXnwSviVH76On9cc/SSbzHw1NGUS6
y/nRUYkN3ApbyWdi+9PsiqcEoKSp5gxNkan49AfktWd63dTCdux4kdk9/JN2i9XXmR6YI2e3VLDa
9O2M+EdEhrwacHQ6igQH740Jl8xOAUuLXWTF80dbdkqamHbOLnvpyLsSbLhugjGILPJVCe0kq618
+73dEPGZ+oRo6XcbOPUUoKDYra6uOnTLNCLvQkZ4HpUeJVRD5ZsNaM0kyUYoO1o36J1H1OwVLSzd
h58mkl+SS/klc5oOzQKqUvDLsCa+t6PzPWesMrMP1J+dQsiVHEq+AOtEMJ3/fJ47q6Aac8iXCxcY
h0kAlwMoRY5I+kDmmjBfQeGsUVFpImda+KhTjmSn5yG6WG57p6dD81R8Lnk/OlvWHDZMlfSmmOLs
64aOdWfT9nBH7LvkAmT88EasuPex1BcWwIX6DlnH1Q396ozgVQe7IjTxG85DP3LC27OZ7F1wspMC
oiYhpx9XwkPc0pzjZUvDYjRCTBpOE2X7DBr9T5lviRCqzKVBLnJJlfBaxSuIvwvZ8GMst36tnfZQ
FTZhTn/0Vm/NG+jCeCJe66Dz/DP6R61PqcLZ11FT60A1mpYpQuoxHHT3uA5KJBDXUUdSBBISv1d5
HyrDhgO8jdQ09qgnPiNOi6ICAqeY8mncE2BlGZ7PZi2U2XhFR/cMyDSF4aIVJ4jeueCNx6Rneq4z
0nqzPGbsK9HVC+cjTBdQWnXkfFHQ2X9Soy4KbXo9C2qI5+dNJ5dWPZzWPLEhL89HmT8bebns/F0K
5Erw3AFN7qwYDqW4y+1s/jf1Xn2azaa4tAABGIyyTxq8TEoigBa/0FhaJTgqBDw92pEDE0HMoe9U
CxQYVfJ+6zO2br9AH73hJMsGF6gCchaeFRho7NMivJYiYDsd1d8M/h6TCmVNuhTvyvQ02G3bZJHF
y4RSGGGi8fUZK3+c4r/64H7z3MCG9gyiMsevTm6tFy4a4wfortMpY8USLPmcnphw8GFkrI1DMQrN
WV6BqGtaAV84Z/P5MIlcWn4Zr6TxjEflafVRQK+CnuG9r9m0yE9pNaxzWpM5upbZ+uopGze7jO5W
gtATcLN5oJ4cTK9eGWreSssjWi9rEp2kenNMiqaW5jSLciy3idhxIMK+MCjzK4PjoiZbwfh322Bg
qhmUdoyzeaY+pnetqXYPmQgcm/JBLT1olfPnw81TGZ3a7y7ak+pjTKjHECGMfIJ9kr1CxPrhwiOJ
L8WX/k14dQIthiLMMTQiOEFCKWqeYh9TfI8LDRSXvkCsET/Ap1y8/wgd5zzZXwFgXbYRKPZDQFEg
Zi1fGXYOqoKhiJLJPyRq/7QtDs/h00W1BBuCHjpaJiEI8s/YFOkr3IyDXjZYa/85vOBuP6t53r4Y
g9LGXQzXPKoLixIUz+VcNK9APOYpAYmGxudp16d5Nw9K5PbcU3Z2/HGt8F2Vk5YMUeJnzhTTX3hO
Q5Kk1qP+eJ2Iy4Gmf7zL0HNEGm5kFfy8oQ1wiLjJ67nvoTuEe0vYhDlSrCiuHI5CVEnoUxWqYZWA
6r/M8azwUtb9iDHucjzQTVtR27qxVlimaIhgWlt99T1wLrCiG8IPMIDkRw3RZgLiDAMwa1srT1mD
bOCM1wjx3Ne18nzCQ/8yJ3CVBCwZElOnSQuTSTyArCvh6ly8yKTfgGF799LGoBD0qx6Fnccm+A3L
gU9PqVeCdrs56t+AJ6GZTJOFR04jbZCUA1QsV371qCA36ijR3bfX5rf8E4o4tZekmIy1IJ3xb9KU
frkXlWjXouheGPdHt1zqQdEKfCL0XmpFxjjEc36Nsy183erGgDBnPs8MtdIHoO8HMpdbhBhMLmU7
IuqsXBB4GcL5VV4MyNkeewPka7Awyk9nXGimrBTOv8yNCO+Od5bjMuWr8ZAN3J5ibM1xoPfousHi
r6J+1nhK/ZzDJDtzlqY3GGpOccRRJfq+FDJiN0O1MdbhVyUx+Ic0/e+D6oJDRhaqDLEC9hHwsG2b
x5rYyhhqAfsTKwYBgfy33HxuXTSJ1T681jJXvU4o4axS87hgMOZ6zYJvOrmN0LY4jWWUnX+wd79w
okJIDLouUgkaN6D0PTiZtwzZlXl7NrIEaywOZiHCurI7u3h77ox4ImVH0DFGGB6TkqvBDky+3ZL6
Z7mWcMY15ujvhxbOKMSp7CWbtotIplPzQcXI48wwsWc4Fwp5PCxNTY/1QMBM8rM+77tyk7+/CnAL
Uq6W7w/mXC8pQdE22vdSOtamcRxVPm53qTKCdm5tdWnb404+PVpLN7Dl5F6ony5hZkn77Dl5hQMx
uFkDUxeLDMN9ZL+AFR4v8zkTbkv+Gqlr+uVsJ9+qw5gasvDlD29AkS0cw9KEOwep2WJj6v7chR14
lOnfY0q7R4shAJCZWEqDFL7Pvs7OvGRuLM9Jqy4v8kvhOf1fgSyclMFPJ9cDVK9FGsHNZlVh05Yj
0Zf6x1slBc0vxYDkGyA+k1RvDN3WOCHmnhAFa4NC65zym6G/1S8Vd/8zfidMT+TrpRt7LvFcFBXx
jvLpBj8XBZysU8ds5vbkVCxdsvZGJz3Dxz6LInIOjmS57R4rcq44ueHbJA1im/Qqu/MkxKA/xfCT
m/nyHA7hYdR251ogsIzqL26UWxq1IoXtTS8aH2W5H3V9sv6/8B1SCAEqKsMEf4TUVcqN0SmAvJSB
dFaETOSzQO80FO1+TogufCFpk4SOYaQn0LvElE6pvqNYiUBKlWj0ZwxUKyBH6IgODZJucmkF2eUW
zBg0OnJ3WLC1J640SAPBelXhH44uQNu9Q6fmV+7MykbOhsHBA3+CXl/ISsjIqjYgQmDKmAtunYDM
GHRfSmpda/huSkUezLE8Z3RNY1hLOx0D4GF2oqDqJgH6vY+0iWmcinvwGBCxkH6Z/877vxX1QzSn
t4kL62iw1FX8Ll6aQsKZsVy1WPs1yCkOwe9rSBbzJflLpaK0Bik4RSMul57RkFT6Jr76U9wc/rvC
Vky5dSZTbFUB4uROPl6HelLbSskyoeGKuYb/IpTNyzgc3oSp4rMPEnWp3T1Bi1/9d6JW0GgPfCo9
XzstPnogvb33GwIbblAxXTIpIlnf6q1Poxa5rRYjsxJQLZqbF7fV+szOmdAcXwj5qQawGTRBCPNj
N3SGAI84+fJtvTgMu7ZU115JHVBmxzngMmWb3RGE2rP5YsWD61DS7mf+5wQwqykdMvDKh18ECY/F
eIHlyb+toNWO7/Dgl6pGIdOYwfUkd3AdDAsj9gRT22jo613XNRlLKqFNGRrkyV49mUPSejXDhbwR
PYzoNGhH+wv9L/DD4gvZiLmbjIIdWiPSUPw47JB///AcYV4bHZXxpjb97cQYehx4LHpUIyklVWNE
py/Hj7kVGKT+EIEBiJK4NbgVJyGUpHe1Bubelue09XPbtg9PaGhB7i/D34eNkmHaIDod9ydUFhWi
FsPlaK8ZByoXhOHApi2gkrs8JOnTDLTwQV8UHSgHc17BbgDXFuidHDBAlsqdEUzc9sVWYF2MN0tX
u2yrffbu5Cbh50D5YjmV9zw9Nz9QzsLksaIfogHcaz98iXCMzWS1DzN3AJ6gIvNYCUg4WNwqbZ9s
ZqknZ4lE027HidhmXFevQHD5lPDuwSuGQMAgYU9drKYLHieIMQCuOV3QORg5pceIhjMOd2ArOnWp
S8VkJKT5Mw+Qc6A7vzzMsQKBrcNy+KF6lXXXO3bg38S5YCzdVYBRNw9QGyiwFErPZ4GkTcVWTH04
aSO3IT4Y8TradgCLb5zYEs8V9dmA3rXgwQYIlsUqgn316qKQ5Y5QB9QbvGihmvNCrHvyFtY7WTX/
RTkedGPt/lnGjY4dC9nCs2LE+mg5EvmE6Y2+aDQsoDN1BKMNTVAMrkU26NIUjqYBrg63GxDE/pZL
jdLL2TY+Pt5+h3FDV0WUJxCK+8E1RDe55ioetmfRfCbQu1zwv3ethzfwtGnfrWbA2ijZbG2Xuo7w
hRbQkGhJ9owVgi8J45zG7nYYTwisKCzbgD4V7YkUgBi00SFvLnrpFs/Q+TnGkP9pmr0kQLaW45BH
z5nmww1j8tg4fVvPxt+KDbPqWD7cwKL09EYzJKYErD7KNj+yppvHVsz8hLSiwtSRAKTxGlWIibmX
QuIWnAJqfqQUFmTYlw012bUrqflQqIUkZC6dRIFm/O87oTkF6nb/9qqqnhO0ype/u7vMQDIKFtdG
+4hyftW1NLAd2tS5/BDP/Gs4W+pNaoTzJrm3uBP6XC6UWRsrHrwt37t3wF3WkEdHtYb/npYuqvBt
exlCiFspER1BEk9AwWHAlfXliMijFUrb/WSIIHMeX2K9360RDzgBWYUCii7jM/OVQEjqevQdTBFs
0fiNkfQ6qrJ86YsNDF3mB2+VQG2yCLSvGk95lvl5qky5tGmDrAYSA/eKr09BtHqFFRcITLG3pQbX
QXDNUlJUtbKqyqLbk5aKfLQKjAeKkgNTJ8uDeGCxYiXLVbE4mQFDV9w9ohpWX+qqxEswfz7+0lQ5
pcxY15SSb7c4t3cHa/XCMX60SZCndMfD7ZV+YqRWBvzcUKcrEm/92rCGnMO49ocxON0fuMzAXeUi
RJfjK9/jBgAsYeImnMb5lAyAsp37654ZDmsI6mxfshBPNnQjOxvWM9MAMpFYTeeT2xRQWYs94X/t
PVEJzoYpbfAVR0XU3TfK0eW2fTwnWNFaicN7G11PmQsYcUfWfefU7EQkAJqGzt4JH8EPSxr/fzyR
n7UAeFmp1Zyd1aGQ+8IuesJj9oD3KXhW0n3VIwqyx5w6YmWUtFjE6tAKjkDgzap+uS/wTVi0ePWr
SGkmOmQq00ijd0wUnBlJohw444b/dKBCMA+ZO5nQSEZpw0hgBV+kTyBqk6wVU/Pain492HKrOgY5
354YiVDC3dCpgyrL/QngNHD1fV17WXiTxaWzdMY4CrRBUGI/6D6kFG5G4nOR9lgnuUk09etRIPEC
B3yT5ZMfOIkyzj41t67xpnHDrNirOzkAvpgmM21EXE2YGb5cX3ynXwpiAGqFHaXhI61XPhGrEP8Y
5uBulAhNTo8494BtMra8Mb8nC9MwcBrsxRUFuy8ydx08gUdr6S3prZY5i5msYS6UEYVCObiCU/zr
eQGVnCBNaipWvjGJH90ZLy8MIc//C1dUPUZASDc0RODDKe4/CNsPD4CBJNyno3lgvpvRzEpZjWsf
lste/3x6elPRV7fJN1GtG7K2KWYbQjcPPQoQ6JJf96cRL2c885gznIvXLxDJij2558HqRDnf30P+
3aOpu/WIBe0rdlgB0mDkaxpwuXsM9OY9orcXSV2grYcA5kZnEr7O48cU5XXApYKhAsTbqy8aYEjs
asyQAdBPfRUX8YkZXIHooxArXML2owtjOC/lLN6fZ71JLP8W/x8eGezG89h6swu04qVdMShQwzwE
pzPFSoXDjsZxrPhIJCSOvIippV6s5refPr4U2cdf9+7LJLGcA2bpEoZ54M8m6DeCF0Khq+1f+05D
ZdInXUjHsWJjxpf8cS5udY2Y4ge+yHSwOj4oispzx3dRzpwu0vEi1evHEjw3sRiuVUBQYl7RYRs/
7g2mJokDIgucsn+aJ8HeaDquBoPns1cKJENXrQ+4Kx4gVXqA3Yshfmw4GkPjW74JVMmJwjQy0ejx
oV358c4Gh/48CVYX6iLj2wiPpbfmCPlUpl6bjHIGpC2KcAQrLKr+Pyy91OH23m4zN3PSwE4+7etD
nuynIKn8VE5Du+bvDupKIvxHBrIK0RUGzou2gjNSkX1q1NsIx0aIV9pqIlcqtwwg3RB6umuq9vcI
u4LKJ92R3w/U2lglzw1mZllhOHpJQSRSSpTCs+oNTYNcF7uJF3bRlaEPRqocqVHwxLNgdIzxFlWg
XgLikkl9VU2s+IaHVsh/qXRtn3SOCyO5ouWgMRyzOJ5CrSgaGhZfZAVd5HVvedCHfXhAfCqJ3duW
i5PIlJqeXEPe99eH1Hw1Y5EPe42VU3LARglvElrIbS1D3NATuRAjpbFC0LkBnjYV1bIyGf21yueH
oUH4AfEUaHak+jyU3Y11cuvyc62X11EeDACPPg/fQAkdd8KDy2HnFrMVf3MsgZwfH01azU6uMCXk
MyUJRcSDC5X4/nm4yDVQitXW0kWTE+tev8lhbjr2ap92bg3nXzUSrWchiSQ0ix9Uwf7Bk7U7rmcv
oBLSRlqCzRj9IHyCIKgLzkBJDObi8l42F1QxuZFIBLmc7yO6TXNv6CiXra2I2VfMXKHJPQTFiy+o
IOhTNLm4SCIw+0R2dR3WkRGasBORH8ErfNkiQnEs/a+AR+oMpJvpJWzi1PBrwMXDZTlR4ClA64SV
B8EQenbnCSODoiksa0c/dwMAqaaMYmbyzIXa0XuMZFWLv6gpFM5jDoYAlvHsXsq26UJ0nb3y6bXe
sbl2dhp06SbQ8mHdQXvSsSQTiaTnUmIJ8xH5+8VfaWeeruEFMLdQufHLjGTZ6XxWDnZ02ND+0q3V
+c8Z7QacuW53N0G8EBfTXj2docKVAFz+Z2qy09ez9t2a6Hhe947GEjDX/lQ+6gYuu3vc0RO8wu+4
gNO2ljlZUmyFHCjOMyqOxoFsJtp13g1hwrPc+C9pPTMr3IK3CFlAZ7q99p/IrYY4MO5GPBDWXt1l
A/IJOrkQik3gqWmyiDnlErZdehRPlTHRlfp+zNuXg6D8XgV5usGTYci/Aoearjah9Syrih299WBx
zzcEn2wijpo26+sRgvqLOpxImcxRvu+43cPY2x3SseGKsqsGIN3AL6t+slZF3MX4izSAxpENeI1l
4woZ6hUZvaY8G8fyICjNZ/WWrQJ1bJ6JbbLXzig80qHm3Z77YJBkBFE2FAt6C2WOVynBoM5aa4xe
tr0GkfAYAyp0QVRomAAYuiadwTLCcXCAGwhCHDvGXWoG2EUYmz8zpn7lFqNAkqQMpdrckVSgQ28Z
PJ/+d4PEm7IrvW/jsZrxCWavQFAO/vjw5zj9dqr4z93xdRLj33epLIv5CWZovwwUFS7zialYxs1s
EvQ5c8iXX4jgLzlLmG076I7Bs17tNVIs8JFiuPWjBpn+N7usbdYwd2RlzvLPqkYGxnpGXc+HHyx7
uhhXwNCLKj0ZMieF+S+fpjgeY20h8z2w54aydP8ks0P0o7dAmoEcrx34SL1nNAI7pbTJgRgy7pQ6
ajrrVTO7KAED/LfcsnYS1Nnqc7wfUrA0dRG2s3zLiQyoYjvdhCRg97/YcFdBmoWlj1ET0XOCQ320
Jx8JLHMmk5jIZiOJJJwCSVEudLz5pBzHvRf14PW1eZQJMVA/Rl6HtMRB8XwAg/PFePbyw2NM+K5H
wr4J06clXW5Y+LDRW4W8g8DHDX1OU72t7fn1BJTPFSm2r6/hqn3FSwgmt2QomHurWUHG/fdTMDyB
fwGeF94C9Md6PZl4qHk4CVpr6AGFMSbRlqS4DcizlCFuxayFyqvT9c0xjqUeW5UuQ/UPN/HuX72u
NNQ8/P+GSsKE6d/1dRk6ik7sAEuX2HHWFtQ+Zn7cunaylXLhjPHTv43D5vB7X1SfoJlRWA7aOR/A
TYV6AFLIMor2NOavuBpQfiSohbCuRdQ3RK6We/LJfIEz4vTJYvr1SHtTSIvX+P4qVYOcREK0GKjw
X4kZsiP+NZO6ZfK90C0MICnCZ31BpkrgFRaNi6v7GJghgVwgECPXx1TTzRW2UXXPBKabpONtNKOl
QgufL9r5RwXi198GCZBt78zuBxoQnAQLC2O6s2Y7rLRSzdgU79limbCKo8GiUlDf0Mwt854YwdAo
IZJM/Qew8LBIQOnnDKv8hpRXS3SmSZUXQeicHYfh9qqTRQO8ZY8DW8/9uqhrYzWdbycJlAMuN2LF
Cm/MkjVTMXpwSJH0zg1ZT6vM6APq2T2vl+mgCongBPO4tEbV7WesGkJzY7pzqiRhzoFeEK4hOMMT
b/APL8qL0XeQHhk17dYjSan4SUx0C8yyDH9IbCv+4fp3zQaTvGTLjjiOq6yYHRvMsyAAQh+7oIlq
0cTObs0Tu2HTugbrezC7aS1J/5hid2xmQJK5uMlHrgdK71uhA1PVZcoFTaf1ncXTxbeEffiSxc5w
oMsFC9+RQhEqP1QlwjQ1eRZw/9IbBkLH7S+cVx5BpowED2+gEiY4q6x1edf44tRrjdB5kSjF/Ph0
fE58DRCJs29VU6bUzYsdeNZFvOKixyBi6cO6zY4l9jUlA3ckEOaBh99ngxETBhM7J+L0sZmCApz3
idDwazBZ8vDwA0gXMlOWkzglEYSa/Rgb5YvQI4d/O8pC+CR3uITkD95bYb5hj2B8shwN0epQJ/mS
jqzSOnNp7Nl1J8nzIrVdfwcpBJaBJBoMr4eJvhqdOwJNJzUTjAng/3WvXXZUZnbTIgYEkhOWb/NM
ThVxq5yhqr8GrhTHjMGkzVUomUsuVZxxEf/16pQRRnIcJCEciVpw1Dxs6wfEl4oDKCI/4AFwg23s
G7zpGxK+oy73r5EEXStukbiTXJLGxxLSRdJfvPj7IH/NiJkEy/LDCgmkndwbdk3BblSh6ZNKELh9
SfHKjEzkwJIUZw0Tl5kwMG4gFPpwCSkYoSLjY1GO5yt8FBDtiI/AGWjSi73jiStrQILUY1gqo7Uw
7LukEIAWL80suJ0iFbI0EbLfed1wWuSpCnpWLxEhwaljakQg4z+5qDZEH47FkIi4rvpewueV3YrQ
/1vPP0rClicL5+dPKQWWlDO//13KhUFMFaMJoZeCMlhY8pBf5BJJmbDj76xi5kvVvVZ6lJokfMWf
qlRJ9a5RNs9P32LQ+6K9/ctBco15H5H/bwOu7cgiavUSSO/CLWOX+B8VFBafrYigMIccYmS/Qapv
jMXgf3uW6P3j5ZelZJJJ7EBotfYVooS9d88dgGdA+FvKlGsE3qR7ZDM6odnQaLeDi8GNunhjbftX
uRUqnZgcNmO2zcPSF9Z5nYnMVAgspD3N+RBgEkY09pv1FOdNBTyafdwxeUsN9bBrq6kBc3hLfUaR
kuOGtFRFLwxEz+L6dKBVm/Lkn6kjfmZkEDj7sA9sQOsdAQMqfXEt0s/GSUTFWcNu4EPINfWwL9F6
6NZ7fcZSvqQEQnhAzt9OpmwnRmlvCi7LnuvsR6GWyIKOPo+v6quN42cESeZaGmamBF14oFsO+eWS
JovPxk5IcwqTXLtZ4CVZciU4TTTW3t96Olv0VjKo2aIEz3GfToiQKsL8ocqGNF0BFCdNu53Nxofd
vPKvGuHPHms9RtVN92IuKOgaWQejir4UWfMxRA9qhrtgiItsaqVKjApyJFCNfvlzVzMyDNeTInSP
M15M4/tbBcRl1WPhqvyyCUwPSnBXoJXWC1Q7eTM7KgtmQYlVw7DIrDlG2HSOdSUOMKmWbQuLHihF
lkuR3Kq29eC0IgGJuPpLt4xk8qyPysXnEXePPJwbHw7MrwQ61xyfdB1geLSLfcS84ggdswQRT3E9
fTTMGNolf35o71Fl6dpjttB11/gfIZR+Ss1aPIiW70N6i4t9HZ6vx4m3F5aG7K59wkVHKHL/GkHN
3k4gusbaW3zeXSCSlDHuhrE6fnHlRsPwnnRkBxBGL6aJHyWS11Gmf2+aI5DP7hRrPM98cDdzqfbY
6/V2UcckpAy6HunNG2iH9iRixDEBDMGtvvGS8uFQNXaYcLAmbNg0N24dturTMAYA1PfxwZJFE029
kv+xHIq6XROVlwXk4s7/Y/W6bmZLqThwt8PZp71F8cEABvgBNZwd5Qb93EUM5L2g680cwSK+oMv4
Fl3XXWKKJxrzJFYve5XdHUphCWnF0LbpF4WWSR1J3De5QU7Qs2YkJAxsaf9rmnTK5zgY7lwG0cJD
mQdKea8eMow0pMZe2/D5a6i9vs5onofT4kkTDfOYOqcnpxt3CuF88slmRbvfmtgyR0hN1JtekfrY
s9sUr9CQIuhdapkSb23Jz71a0bH7C9DLEq+SCzYDhFIGbpnJAetEOKnOY+cQZU6IalL2gdWj3Xj8
cOCESdUAfpKUyZ0vMFEnu+8qHLCVzD5YPg9I6HkfrYperWUyMd9aHg73ExX97xU0uSmD+ot8PwkM
PmTcVNJ8Qm3tzT0m1v8aIxZWODKPh7xWfCJZVM7+gMtnVdvQxNkAzCK5GL7CviQLfCOe/JkHFX/a
9CQlnI4dqfXQFHvvdrmIEbS/v0/9QORY4MnJI1idXIK4W5T+GBymk+OGgcLVZITkVcoz7IPB/8B9
uvJz9DbLXcpy5yu58SiBWEA01esK0Fq1BQ0CHRgtQnkCxxd8KNBd9HV8/EWVwYB37OOfNMFCFcpo
ryP9avWoVLytR5BDp6A4B3jl+g58sMHR0xVrMCx2tkJCvDg/azGz7R2foeoIDA3/nWk2KmEI5i8g
ibjWuXLqjXgTszxLaRR4a034h+2m3TJLEwFAl9F3fSNcDQPjgch7z/2mqqMunFEJO5UGYMdg7nTl
LrEvieWi9+HsHEYgmM2NEjsaSRGO4a+gk+a8MYr+zMh9ucyAgef/tPTiWrzz//oUSEb2bYaU4aso
H1uRN2orJoQVFWNuccxY0bsCSQaBjPgNUX6XU0K/1g2oCCvskZ1mLE4iJTyjw0bUsPvFCXI9pY1j
ucAwDeWYUApmWBOSBgaSSV5TxJfUTYj5Lxc//JCyE548pX+SOq64csdzh8C+OzipqjkabFeHF3+I
9ymG4dscNwO6NXOlGQS/r/Nq0TKLCXvlH7ZAo1lB2hykraBmJwkrvvOZBAsPgA/XDdhBw6Al1XMP
z4QGeHQH8THFb6IGyYWDClNzpRrnyJbzA5QFrqznd3YxFu/EylHE8pyeD1Ztw9oLwQFbBLCu+Ejm
nQMlwq6cwX4du2R4KfyybBGSY5WsbJRio1fFwrosJHqx7O9fMijGsSxW1InzBREH/9flLfvFtZ7+
EKSSU4RjR6xdhRjJRPYWCrKRUaFvbfF6pqJiaQI2/gba6KKMReJWjIehpNMn71c6BwsNVXQykrpj
VBbhLra7XFuoIQ7QLNT/yZdKpnhlLZgyBeuBTB33+cpFd0PWO8AqVPnn9/SMeavkryxlHL7SdUIX
E8HGrgIEAX1sTflmM/sDDNalW2IXfxblYy1YwAldDP4xP8vaa8H0pNG0faX+w94CMhmcphddJ2Pv
XPuunS4QhHDN+3Q2RB/O51YuLBX8aLJtSH1BKNCLfXKYr///2Gxj7UIV50+3gsKp795GbkywYedl
RC7WXL3JhcY6TBT4HpKHN32dA57USV8yldTg5Czwq9ZBE5nMjXB+BN6Heaz563putU+y5tK/o8ux
Lk5LlCn6lGFPcTqeOdiCsz0YXQ0RZf5uE0p1QOLXEbAgL43d0sCyB2cFXNudvq9CqrDiXJ+Rit4q
I8CLSo7ITr6SRwd4yVBInvQF90yR4ByonwuzwJbD+u3oxPzYhSc8Oj1vgZ0RaNyJdEoS/eS/7TKO
dn3SPCaRjnFvVvvPCtXCBc/18hh5T3ODdkSmRcCCA2mh9PE4yelUn/OlgQIhHWm3jzelXumZMVUY
mE09uKTsZyk7u+k2ljJqLPecMsdPjGJtjHS6DENJcYrZZG8V77QUKdpg2vWd+uAlx2Q9r8yZhqXi
/P57ChLYvMCnuGf3z//YgY4L2x4SSWUoeUzqqWZ4kBlRnYbDCL9qmiP6wC3wHCAos4+vcJVja5R/
Iz+NMaiFqaq5+RIPjrBSR2N3M0nTco0+F69EDMBwluKQ+9UxToNyqCvk7v6Pi7XPWWwak6iR/NoX
CdFbCYI2/lxcAKeyQoJQp8XTaknxzQUnyG7gemewN05TRByet8l8KBHI9IebuvOV81AxCu6LoY0J
M8jE24Ilm4/mngmGRv4GZdyWkYTbmT060mvqdvJJUFeHyNCj1RRNBR6bLYcOqlPAixjwkz4Fshpf
qSJ5RJUxEa4fl3NRHon7rnGXF/LlkTOSU3/4pCYc5BNInR1dbXeDb9pc68otIsGT22q4tkbCgGix
c5s27fd6xuIAF/ZH5L7fj8wIwFe3+3Vxb9FjVnGGsVpJjfFoiPYF3Ne1lHMAXnUvZdJaJW5n6nX9
XOEgqObtN/BH3xJRNOK2gC0jDVEVkYFYW8mGmN7DQbj2GBgu9/CEnpNejc+1C8OhcESokJZIzFZh
Po/oeHC1usyvT/aExZwadLL8IyVKIG+fB5NFKogRT+aEClimgR2wdR2Z/zvJL2GpKz1MRZKXP11S
TITl2cQ5jBt/tH5S2CDYAsUW22JXfDK6xIKh57nt29rJBvSS0/tt498qHPGSFx0g0HrTAd4QgEFe
sjYI5nL8x6bB3PmxDfSOcQ0bmmrvxrLiux9Ijp9tVf2WJHxHHE7ATF4gkRWIJYkep7pEShuFZHRI
SFr78PXt5FwhtXxGy7OdI/M6U/QC/lxAFPqsFgIHnch9iUNrVbdSfYZrb3lEk8ZYwjTHSRND6eVB
Nd3S2ssIMFdGVAeuwYiJOMkJILGmrLWBPeeZfV7XRf1SSUnvSlUINWfVNCmCrPqNVVAUIt5bhmAj
TWXzVNqHmA36YbDi7DT0lDDEIBvnoMtLMtF6OGWgKetLIrOw579ig+L4Qo6a1z2AhONuhoNqO2bO
MKuOe0DTfv09R+Jb4oLXTEsNCDiBnOC49vjqj6axhMrs0Xtb+9CSk+8irCPwc9GKzwpVnFY2/nQ/
K/pM30VKZ1ljjXET0YTL1zZ8ZUVHj7drAcFfWHYzaunukb2ddG8Wa2PwtYoYaenewYo3ZKMpys15
NtvwoP1TwrGYu6X1LzRtyjD+UVKSopCiEXC020EvlUFbyJGfC3ylX73lRhC9JMz6RNmCZkZfCfk2
zJ/O89wC3oVbkeoF0GvSEkFTVN99On0Fq/T54E3WTz1TNx2FkcmhpqDMcURbPiUPWEMJhq+maUeA
VgwaA4MZm5D2hBdCYXKlpEVCQdSIV7sXmw6xG3mRYerJoCk6GcGmyimKFBTDT0iIHRgyw/ARSYSA
4X97NUk9YDVKB3OKjAfSjzxG/y7ntONpBkHg2lGHYQwRVsQAYClIUK+qeMczpROvJSTiaNVE6Oli
CDOOVMjDiOGg1v0mnsodUOjcjyjAO4ef5LBwitHgYDvnwOry4QbDaN6lDjzAgzKci6DrI5S7ThPa
jspJi2oBLgH8M+gKkNzYqiMzyHudErQW2U8dPA5FVKAqA9TOAYogwRstcRqDL8O1zj9QDC6a3VKg
f2a/eKIxMrY5bP99HYJZBL4klZnZsnQ9k7relgQMBPJy7g+nyMmFSIQGpQQRI5bCArFaVPb7EHQg
zfGN+u5YGoSMIC+7mpXfL5SoL0c0pdpU84nl1NpZAkvhShKTUsjZuoGkdXXeEFa/Ixp2ziyNan40
VwYfH0UvdKiDarmCtXdIg/ivP9T74ox9ZX2/4DOxVlxKQWU5tVRpVsa4oQdwQG7usSgEtrcHUMRh
FWoLBaPZt3HoeqZ+diY4kMl9FgIlW1lRMJHJgmNIulR53ZDHl+PHo3hEUzN+I240hwvnxa+mCAT1
vZ/UzXGwiJEaFVBjSEm89nWiPeMc9ueH7C+boIo0WCo5Q6snZjj2BWqYdEnB/+c4KRrfTTl9rJAl
u0Drjd9EnBnLEzIEIQihKMKbMZ0COYTogeyTUJ9TImS2SMm8Nu0si41YZh8GTJ+7KT/tBM3I1KUe
Ls50hBuhRv+eIWZAV39wBfiQsDqjAqjdmi6BcyzBRrtSaSmwZ7opSn+6FAZlCFwNihQF924YnsA9
HR1+m5Ej6JgYePmTf0gM/s+3wHhn6ZHxwuQIGfyJQVNy4YpjJcD7XVgTX/3b2i0N6CX1c9Rj8m+N
pIqQLzoMAb8PlUmgFQh3VPZz+PErLi1cfiA8GiEOy/zKePZlQrZq43vDKDYneC+vcujPdcX76mmS
HE9rjSZzcQVuv87kdLwtawbIPM3TZliS27oF/09D475zv7rEVvODAMykO9Dc3rphhiqSVSRyF88+
xh16kA0t/v1vmAtdkHeGBqxJgBxWAuuKaEVhsxC4sULnhdkGgQkyc9jSbJyVfeTG05f45ZGca3EG
cjgQCXDPry41itVmGtkTxjaM9+ZU1OzmbLwfNJtBMVNpgkb4INkLtVnui5nN06IVKgudplMwchgP
laTpO2OmkbaCBRPCmZbtaXwhgT4ITuuPUs884rPiueYminMS9PDicp7bVscbNdCDw1ZuJc0foDLv
RDD7IFUqGTmfwnKGsr688AEMCh9FjKi0kQwAWOn495iTeqVqceN59td4sSF3U9M2Dc87uqPiduUr
4BOTNDjd5uHCrEk0w8fhY7jvJkxYO6n5M4klctlZBbRPOiwav6i3Ii3du6NxVx+AbZRD89RuRHGX
cvFIIksUF+Rd0oBtIEaeJryvL5KdNHHlWCCqnwrP8rGtduV9lJLtVW8lr1sFr1kxMbfpTG3oPmZ+
Uv1QYwab11DFy7yCTLLxIoQdf3+k7oAZnUt6h/H1ybcVG/btnnH8i4nWBUJdmaEx6SeNXlM7n1Yu
qZciBs9gLzzd5RRW0nyJgXGj9nSXZzyTL89FEhGJYeRmC+/SamBghjsvvA2uHsgzisG2iiUp3HxN
mwJaeNwkY4+gdejsxO8ttIS8ujn3pTkTDhdQbvk7tYDahu44OeqUEGQBTVZrzjNix77IFeZq3jpN
kkvaxoxbiKKvapsidpNOgzRJxvLZUF89NzpOBPvqTe65OE957OnITQIgcA1eOmofU0hevXDoxmZU
vvu5qWbZxvOdaOZ+DQhuDmExuSTNlckUMmir0+XveYOFw0LoWDtPpYksccESnk8sjOCj2wZC1UhQ
ywx/as73xGwxvi+ZiHCoD6mgMyQ/EIwQw/i2M5T47x81cgRAJDvI2C38+v3CIO5iNUOGQtgAF3rX
tCOoT6b7pY2PAqhMzLeCTy4hXtrd6O+kJTGXcqt8HDKuee+ooKQse2NFJ4na9Ly4NF8RE7T0fqlU
+RNHGyV/rDENjf0sHcKVj2k1zEePucrNx4zv4YZM2kBP0kFEJesKw/yWZaeNoC2NzkOxRGaG39Qu
tikj11lTZr0MAOZahjraH9CenshpDUpfDLqrB+GUBXLIPokDVVZOIgINIB26zUNWizcJi4dwUIDi
hh9+KcOJSFo/jhyQo+KbM/HmExCsaAUkE76hXqE9/sRmtPDX2wMwdYd9LUwknCPLC6olEGBW8ar7
nixw0pWvZcEFB6fNMl1bSXE1Mv3+No0hbPhg3SegOZEazQIqaOmSuPpCxN8hy6xA7ORscRuAhuiS
QKPMIDgAoNAzzhNWlPNED+KVLqtx2CC8YYQFuFKVnGsxFyekKkPeNvTCDR+3rO2XzxipMsVyEZ15
ecDcgdRyjSI3M3d4rz4v3tDfLekUWN3mPFu9HickEexBMZa+ZyFunfAsbYgNOsfcaIfOqjdDRNh2
kzmT717MxWL3xepcDPo9Beukngq35Hb0C256EYOa2jhPazsnX580X1teOkFVGvAPci7+NlfYi2KS
DfB7pv8e9PFQhTq7PMGS3lQzSgefcMbjlHXP3QNZ13Ia5Wn7/+Dk5WZKitelw57ZXyUP1VkqNclL
Gpd5V+N60L4HrwMfa+r2O3v3xjjych/xx/7PfXbG1/DKTZ2+7XTGoPj7wA/ctp05jRwL3ruYF+2h
swQknBxyVqDkItX/LLkmGZ9RhQdQcNeO5UKTyi5k0vZ9q2lDFTZ1jkTv7N1S5TrPvTHMzGpTvneE
SX8brMq2QW9N4/f7V5aodzwOQUaV4oDz8TIVlj18R267F2TpVyuvM/7R9l8KAUtrmex39CD8DTIk
7ASuqKy5hGAXD4gL9XBjaKSB+gedUQB7O4mskqMdaUt5MFgg1zyovetHQqGgb/Fp7FupCxye8N+e
VRtTrdwVhA1LwgUTvMZIYwJwh0uYHOfXn0ActadYijSysocw3EsqaK6hvFXc7vWdsKZVpJBMNZqe
hYMSuueBUb1NmzWMNtxBuyShVDAe0ku0FocHXG3OQ5C6bS7Y3pwhBbIcCR+bG5KaxE7PJ/sgO1xJ
4x1roIiWeMroTsAuMQ1hsYqGaWNqgAgmcS68BWfeVjNFI1sjxhwJh1DRLaGkNRWY3YDGi7j1Loo5
896BmSCLRE6MwtHQSEw40WVHPu6dmfXJJiQalL9Q0epa9iovL85IqU9k8jPLzYiegW7Iy7MeCwVk
X+8KsxPLPN/RPZ7GurdEtvdzPwi3Xg2FQsQEkrd2YOzu34iSH2aQbqMBuD0Eny6DzZwvvqHRITDv
zPv70O6riwZQ14uSD226tScGOakqIYNliIGOJtmFHAkI4sNnW8MW9GJnjtnBVmvvbrNKnEEkKoye
okaA1tih/0ui09FR5vch1ix92xx5CKImEXVQ5qj1+8Ll0XHYTaGy8bVKiE+s2NYgRc4QR5TSfcqc
vuWc15AH+wnWnBgMHMhennMqrK5S2MN86vp4ztwayzOeb7t+FJJ+dQ5xtrldnqezIYvx9MdpfIqz
9VpCZ7YmAoR/aylwC+N6gLxVrj+UAB+91OUS+//47AYX67eWYI5PBRtsZ3//zuAdIIsDnpV7Nq0j
GXAMrGXYLL2gcLBU3u06poq2nASoRea2iHWhPUxBB0rxe7KzO8CswjSvpmK68sE8R3dH3TqYMHxl
UDw6Ue3WUnE9FL6d2VeIbzSYzaWUGWmxiKb6CSkMH09Lvj3hNUM1uzOHcEncsQb8RGQ4f6LCGcgW
rXsKGM3iFYkTpheG//eqd5G1LFS8sQDwcqE1ecC6dOqeoriDA9rQOA5VjnixkaBh7Z5ZjQiAGpam
Xiw+KCh8vuBYTJEFgsjQcRhWeRAgJ3Ply0rh+FhQG5kFGiR88aS0hzNy/tQvivnFKUn33ShM34oQ
tHQus67yxQZgiNZgKMMqAVbx8YP6GgvkLYjwSQ4PRPtpZVe1Sf4s9E4Qu41hMVyu8xLFaWp5Rae+
QC+YQgy1+Q8ICoVdsxMzKF4fiUfawd7kckgsyrTEGe9CZEJj8bVF+EWJCNotND83B4GJfQT1ZsNq
ek2oDz1yLiO9UtptLTjfj7MBLGR3WEvjmnX47b/XltX87NvT0K5PN2Ba4e0qMIpfh6Oq02aNNVcV
+x6gwp4xcLd5Vog+nEgdkx/MlBVUrCjK2LURf/vhrd6lotKnjsIDlanaBQ9pYghFJFFUJnFVwuQm
DT/vBZuJ8qPu2kkT+8o70KUA7gsTgJrWtIalGq3+RP1Zfy7xUOlmjhjqh96NPi9lBsBdPd7qyrsy
webmtvMEqO+gGDJdmb3+TZFgeZKfw2jPu2k7qXkW1b7fPAzX84B1t+GuLkQx9LO/i3i8QGiOZ3iJ
mOoi/O6Wgpb18Q4cAEvs9ikm+2CiDCSPUI/dJ2C/g/mCSN2V8eMD4BaEOV6Va68jDPTu8ZAgLuU3
QPTJv+gWp6mZxO9Wz6Pf59O/aD/QPduWJuzFjGq2cKJbrAR6brkoisolMwW/mEOIAdkiafghxa3o
xG1tgx4HkPOUS+V8UggHOeM7hW5JNLVyQw3I820f9tvEXMHroBE4Z3fUMuu0XFl5NV2NZ5EHhSN7
rfmpPmZAM4Xf4MZEdlGLhSdF+DkZyxSzjqSMyP1OohKSDlDXEgnKz7cidUuVPPV0iF6Nf0PvZ0wZ
LrsNUdZEzGNyIHENKFruC3qK8RzCIJw/NJB3zdJTNWhYf+dyg/u0Qz8cccRMumOcQNbNgl1QbLnx
7kK9ke8wECY5eFlpgZUfp/a84Y5WhiM9xWf6NKLBrGIMMHg0UI160HdWUgUSOZm9iA6cgmaUm3tN
L1i/c///ef5GXu2fxvv6UHfihX8vOT8CupJGAvi7L34G/Gje7kpk+rge4iR8fIY5+cqUUHbglV5k
V2aokUW3bvN7npgI/m4a+xI/6ojk7gQVgKkdYJKfjwI3tV+/nUvy1qVyJmZCcFzSVFBHc+SMgrk4
+MPC4THXmtYj8Uzu3Tnnr8CZu5O6tGgD8X98PbxkvFaP4/hgPEdRjoSR5Bmd+efEhuqafxLBH8KI
cDyE0u8XLejqSmEZ8uRlLlKJ7Noazb2n9yPNL7isz+1wRbLmiLaxfNEA3v0XbNcl75VL1UAFSigB
LvNpI1RoN71ziI4rRDZlrLv9HNW74mMX4GekhHq2NjhjdKrwa7D3Hhv8AGc9+tJRSzU5ESxf0H8+
cCorrzHY+8qL7kpBk/iH8QdIM8fPkkaXzFnfNdjqnj8ohQmoHaqHbHvdFc0gCPMKWjQv/FvNH1y5
tpTgPslCshbUEDaGlHCVX2etzropw24hyOTBUfn8kOAIkeX3H7rddHitfa51RpVHHEZBU81wuhdv
PmWEZMDAksTYnUgn+tPR8l9VOGQ3cgsXwSSJO2OuzdHRbBP/4372ZN8zS2PxTHZGXkBxjDsRO0Q1
iyKSMEYFkszAUks8ew6sLoX0P/zzjlBOQuZwpC81TWh97gLMmoBDG6B5uV0D86V+J4iNyXFOKzBb
wHfppESXIbDqo1BQDgukKRbofB+U2dlD5jTFGzpYEajr/N6dO103KwT5z+eC4U9cwf5bPvfx9eMf
Gt/oWtd/P7sBd26Dbk3l8yr2GE6bt6VRT1WsYsklHtofl4zuYlayjL6lMmrKuwVGPfdbNHN4SsiM
Mg+8USny8j6PRIurBmzCrtcEnH1g6Z0biChnPpNxQfRjODzajB8scccZqpqPINK6IqTcdXK4HZPn
o6nOPUgRCAvxzx7GFD7xN/4vXIqApUpUIdfCHNJ2jaOPLCUU6B3tgHF1RgnW6YzKpZOpKwjqn8a8
wNpx7qYcO1Nhlx9sYGKrAwGwOK9T8LnAQhuSohFRSIGrsnyrFl4KDGp/ghT7GeWY9JPHhKxSYz/L
kCNSMKaCwimL/+7podaupbs5Ny28KPcegh9D9VhsA9gKMNkNaH3CE9zNqw69CcjUcld3hZWW4sPN
2wW/myBJMN5CpQkKA8CeVLsCt5ZIBI6yDZlPnsBrMGgIhlcIJ44y1Cxwhn/WPJ2JOMmgzx7b4uXA
dSrlVFRThwSNJWesGqAPCUtPOk6BiG4GFS36HP0KwAFDTpQUp6oeMDy6dnPicpyd3u/LVC4tedb3
ID4v/ONudfgVQrYaaOev7h+MsGwef6YU/a7fSImHDe8hhddm3ZYJC8NXGetyfcjj4JnmTmm/3TYw
Ief28LIqPIh00gSSCP2YkfSXcXF8izt+HOk9mz1RKPo4VzqRhjBs23t1oRr0nZ2tgiojwFeFunc4
YW81WHzXKIJHn6qWYfGmISGUgjCRFGeFYkBsYezz8LcuFb4ryRdpEPM6lPwTfWh09A1vW3jdTMTb
qt6+nteOvCp+4Txp7HShdVKxPtkr7fOchUkWr8RSusc5ESAkyxZpNwS9+RSgJpgcuEAlrxvcaX2C
KsPS0CgMOhhVPpasXAA9hIyFHpRiJacqQtYJpIBIadZ8GEKalstDhyaflNTg1XWa6SsPGy2wCsJZ
3tWT7+PtiQ4xY5afl6EFFc2oaKFD3/mqaui5aXoRKZ1pwO4tH0VQaCx0ux7pHY+XymQ9RJCmkMZD
UMXIJSEqG8xXK6DKQByxJmSYRdFVKG8thi1UkaGQc2PHT6jAovDQGfbrG2ghKNwig/H7qUHXdClS
X7D4bQt7EDU76a5sZTVm4h8CjsqXErUIovkg61dl8xuo7qieexXGzeePJfL3x3yE71KMMOOFtWQ0
bITjLBBUmBanqhwSH74nmId+s7hlxjbOr/WgGrxFY9sex+PnQERmrk6WnnO4bc4uTd51GH4VN6Qt
jKxEJszt1mFniCRgxyOtQ/fyk12Kg3fIrx/8MmnofLPrkX6D2ZCNPDi92s6KkrGnh2YCaCLRflyq
ETamYacbimCnjBz90XG4nEMdGVyDfTyTpgn78gU/1Mb9Hlf+F3EcNT72gqwnsAMM7E07B3z/FRwx
ghwh/0jZYmbyS1QxJL1IvZdSopGyso3Qrx7h+/EDuuFUeIXDuTsu9SJbw1ZTKZ2xEKlpBM0CPtbQ
DRnpVyHErkdjhHj46vtPLkqx3AsRnQsS07QtmXNSAmEKoHzDR74eh3YokSFV5AzpK92SObdns6JT
yq/2En4/9rDvQ8lUoEM3nqC4ykxeG9w0iECnnsFJKso1loOzsEWsp7O/4t0RLZeCqPdtML/+HJpE
OuKrE1aho4kwi3cFXSW8MEhMrYTdwYF7nJMsBIh4p7JBL3h7RlmixFy1C35rFiEtzyy59Ip8gxwt
vsY82OJJQg3GOIn8P8pD7uX//LiEPo0BegpC8dDqpqp0Kp4K86FWyjEJ7A1tSWo8Dbdk2sS2SM8c
ma9jPRHeWKAHe09TTCeRKchZxoF3C0Cm8pnYxh6Q7b0M1UO15Ztd3aQJlbUSNpq46gSwj+e7J1ma
d0PFnY7yy8Ljekssw4lVCkexLzvRDME3ZRl1SeaJt7roRM0JhkycUNloclivdT2ECGpCMKGD+9Jr
7EoMSpoHPQ//008F4krW7pwmgzF0E74oKH4VVRa5PQIPYikJLkPBGlwq/M4Y/tXkhfKbn/FMcume
jtYBG95BgEd3npkSRo5VMBSqErqYD/OzCg+2DzvfZi7BgijbScjSZDtSKZzkMhMmyl7QQcmEqBCz
8mb1IIbvcBzI7awjxTSdrDG1FxZZKuHEHKEJrNRvZHFNI3jTIfN+daJD6/Sach3H0CYkQiCxQFdl
1RFYiGCtisx6eRbsJqnvP7RQ9CqdTeJZuQNnyAVx6Mk/oc5gYZKTOVJZWFWoHX36aJhtOgh3gels
QuOuKg3lhUjiNMqzTI7zYJOBchKYSoJTaL/AYZdjbp/IX2TgcLL3Nmd7t7SSsZxTQ51Vj4fIIWQK
Dm4ikf8ucgCatPU2DU7lxsmrw7SnDvmtSIQ0lhPYFTQsg6bQgUUFEPu0VWdhKtqAiwY/ZLFZQtf5
0FiCFgjPxcVcGxGjLyzQ79wfJa4iBO/2Vbd5S0ne64vZpJhXJs42dPp8ieUEILXLk3/g+HWpb2yn
Q+IFu0ZHMcO9Td4kIq7bv/YIsGpGPpFUp/Rw9/IKnY0uZLvzoKv0tXeK9IOfYG9g6wFz9IEzcKoT
y4gwqj2zCHB3QsUSYo1e7zXeFbOAKWbfzrFZgOc0But3PUFL5T7nCf/axzbadpg2RBxQ9ntJ4fPe
c3R5z5W71l7+fK9ahL9BwTYLms89fXkeDlxGmscJ07uuGqkDSoWY4ifDo+ectSvYqmK9mGFXI+Bv
EHxBgOs+ocpDTj39UQlXKAC/xIuxOfWph50xjy9R55SZ4pIr9WWL4/F2apwOkCoz2CWLxnyp/xax
TD5ATFHgkWG6D8h858vFOP38IBeZQEgjfVieQmbPFyXyY5/iGQnFanaX74yv31z92CcC0oumJgdH
jhhNWUGxA7aiJSG4cIKkpCKXCjPfbstaWG1fs0Pa9V8HGi9x2FzfncFfdjQa13eb0E4q/Y/4o6jp
dPTF81RbroVdJeJKS+frYt+OY52bc+ln2OQEnZ6Da1s8VaKCWJkC9TNFc2PqkBpt34KDS7YN+Zfy
rZJOWgse08E3B4Bbzz7DHmc6GfNadCL8pwAc0D+2bj83o88EJMsTSOjwfFIVrWXbMtYntFoea8qL
hweg46RlsUT6JLg9ipVafWGGCLDBDxJrD2F0Dip4FSCimqTBMuzdfXfv+H7ycHs7cqNlUhDX5Gbn
XYxbCHDbZX54YHhYx5jp+wA+PK2n087iJPoDS4jpkrqGMeZw3Mx0cAFeA7Uf5MquAbFizA9rTqW1
D0oFec27o5cNVZYmt40L9bQ30oi9xZxTjVKmelbXeo4cUkFvtO0CIx4OuHt4nsi+2d74uRcgObXC
iDL06N2+3UA/VlFqIi4iIigOiIGFYgZUKLVVsj0l+S7ChIOqHyLTSZUmRv5kH6hjB1Dpy0568mh4
y9sUj6WzaUyJN8jaO5EWSu9AqT/XDpjJDED4/bw+dfdXqyjc5+yusT1m96GU7BLHjAf98/81TQhH
Ak8Sli0MJLEzo2f/UDsoneUaW6WhFTjEBtT6s0qxM0v4N1Ly9hxzgipCSEofNpVRQn/EmhDhXi1r
OjewzO1AEO0uKljV32eepTfbjHp58XtEWXok+JYw96acUDhMsHbYZiezGhhIoaZ9X5niySvl0hMV
n5VnbBgRjMpOHq5UkL0ok8S6pUArTHWtZeRUZidzitgNUPM57Flg0rOrwKfrCTkmvQEyAp0Aa/14
NTYbhHLrpr60hddP60NCeaDTpY9YbsY0SknPN/SRhOsP4Mw/4TxnRb3MVyAmoKif1+pyPUFT5knD
D7xO3xu6VKDcDKs5iF7wNNpvmMBxwgjpgFsXuKxNj9cqHOD9GhQAcZ+piEw/UikhsCC3TYMj5HTJ
28yrMUNx0o98lpCAq3STwgSXUhAf0acZcvEwcSn4PIRPnf62RMNO1fceFOhpkQADk9FFkP0j/uOg
mYIU7pjQwluh9lm2eZtkqyshZTlbZOZiygoof4tLLMKUf/MFRLOX4b1FgvtoNFBZd5tqkxABbBhN
7IctVRbBjlM9rLqRmtPxlclEBBV4EwPQhxodGBrDiTSUlADlcqK+jIHPTlX7bK6BCWjwtjKcQO3B
ThTg8j8De6uMtefTF2kkB2PPOGGcgP+3GJvZ7Ibn+C+oU63+1cQd1/G2WK55e7zIuNNYILhdv71m
lLOe9zIihpWYzfeB6+6pHQlwhuMnOfNILl7lLo7PFEkbq91EEpzzScdWgTWfbY/J4L59B+ia05ks
Ub4T5ksaHBwpa6ou9ia+3hfwkcMufNEM/3m+uPLDxnr+5lrq6XpIY+GXOUuPStnjcYEjN1N7Dh6P
/ihFF4IJNAH4IoPX1+ONvVglt0fRpc3D+IAWygBzW66JTSzAlALEgnPIx4Nm1fPfFWwzdPiC2vKp
f8jzM/sY+VzaY1rakZFd0budCy7yqIoS9u50Gjzu+a9ejPjPkgc03dBAPPiwegj/Rz9usqCm0Wzr
JIdJF8JG7CSxgw904wahx/pVVHf29ajG/AW5/3sk/9r1OEbU7mkUJkb+HnmCZXq37zRK9Qb+KDG+
7XkfXZBCptUTBVnhnfBiZOMgg+fjvpSiAsCOTe/2zmO8UlPpViomv7uhF5hcw33GhJp7f9AVgQZc
PALNdf0ChaZTbu1xY/Msu0b/uygZNQFAPN77KuTMoIgU5dJ/XeAY+YJNgmAozvMyu4nYxvBMNnFi
CaqEmgJSPa/JOjYB+Zaa6AVnDlTVzc+nNfi2QeYvIFiap7cEFtgavuiVjm6f/MfWGm1b9/Y0A/E4
OP0aPWARgsRkDFYy9CpP8NsmjZcT/uscRq0mt7IAEZJGW14RX8/ChnOV7mjImmx/jKrcOryAltLt
6NElUrxanJs4RlY95wz3ZA9MCFsWJvemAgDE78DpCw0nitAEF++yaCyK25AIFH2Jzi99CFp94K7e
RWRAID9M2pBo9z1NiCnU7UjTkvQP9aZktKJR10KAhZKx0FBFm8ly2OaiP7leJ9VslMFzbr952xPY
PJcuGm7Do++S4pZbHjvCFWPUi804SM2UfaFa7F0lgx8nEmmiXwQ8I3BHdJKwvosItlXzxL5U20fM
cw+nHgBIe8MW1ghacFfCleibfTOc3ObjDXQXSHIPU7oqKZsFTdOjXdc1f1MKMeIfslSrXPHFAzH+
MNLd+c5A62AooxSoMYc2Iw0r6f1Z/+PT0oTySFz2DOGXrzd3durKU0rJCxzLJbyW3Jf5yj45e/9f
QPjMkjWdHyvSB7Z49cY66635bXCsY+ZqtWCfdRhzBgf7QP/fSIGcQSqWaKpbxm5rRBOEkBUDOTzV
Bbmgwkb++GMsGa8aNb960R/AimNki1stF+qUdl7uwXOv7uz/5KHVIAt/Jl2YUFe96wNv0J/laYJE
bRXlA/l1NbJ4SzBpiqD0u1SZChLvwZUosypL0d051U+x/AsH/231v1jUmAh3Q48HFKmEBFeLHL7P
A1LOjx8ZGEsmJy0UrWRh/adN7ndbx/2gfTiqRrysgxD50muZXr13HZOMcxbPItrLUSQTYBZDOwv7
t0ZARSg+yQuglsZwyUopas5azJCwOjfgRgT2GJ2ThevCk6DqMEpGRS4jBzkwfWpBZg0xDq/sVk5R
gGAtlfb6/LKhHz/9wrh/YAqQ8TrBt4PSFahhwF2j/Ua3gQ2egOrWp+1cC+L9PX4Tggf9wcK/ps0C
z5rkffAqID3znCHZv1eWT3exRGIuw8NWISXUoRxCEMFAZKr/ZdZyI7PML/hGHspaLkWPSG2VHK7e
HW6hVAPbxuGg4vwsl860dT/k7H7PjXHbOO866CT7qePDrg0v4VJkfZbUdM+9jppCScIHCTqapHLZ
Gb6TAzmchlfYsamR7lClXk0yWUXmy+/3wr4mATtzVADtXX7k7Nev6TudhEwKR9jz24JOtEsl5dhg
n3RferNrNazHAYnUFqjWEm4gcZXeoLC5+DmAf61AMWzj+SLVRsRO9PVjPvjs7qUcU7ffgAR8Aqad
xmb977t4oub65Iq+yvlcEZyjHHRbQu+svh0vTF7TAb7rr7erGUoo2SbwFrzxBnX70GHUKs0khs3G
r/uYY9HKaBMyJZAFaPjZ7YALwkn8gGRHuIHzEbP7ALEkj4lop46LzmPsN4mG57MCmlyhx5G9b62b
jmKmXsVBGA0jDMvI9j6WD2aHOflcSyXNNQ8KlDpOFpt8YK2BCmMYQG9DDaw8fRuhihbHq0Vckck2
zKfYy7kbKHxFYJNnTeUJdAFNlnCzJ7ISYWy7fnHMOaHjSCYBrpSdQJvWl+2qPktvjDrR86MljT/L
hxZh18PsH4wyGPmMF5gK5GNjoDDYTLnTAEv9lGHuk7m9AZNhmrIkly4Cx9FVIjg3mj8Uuj5354VP
rFrWQji/A1l5MU+1FgX+dAQeVT2mc+jI18gJ2v7eBOCrTKxcXXcKrNEVcAZJIuhZ5ythTcCC7vKe
rTHjFblyxLPIp0vqrjSW+w5PefDVRF3601heyMFwFDj7YhB+vBrB9+51yh88hE4Z8A6SjNRDVK77
zOfxyyi6dS93ZAcYX+XUvzx0/WjIONUGA/D5jY6htL9lwayIRnu9Hnelb3kqo3D/y+2S6cUq03kw
/mXohuUn/B65unphHIP6/W8jMfgwVit0WeoKchNcrrmYElXdzK00oEeCXY0hv8ieSO49LFueJVDF
xMjkrWkWztX1b+IaSTxW/37Ngnt8dAqgD5YxmCppIvGepyZOxEKleJF1sZ0O2mrPPMoU+HFRml8/
Ct6C+bcqLP7juhiLeD2SjWP/FsTWVgoo5ST5BVXjlhWu6eJ1WLPblNoKs6FUbbcZrVXZ/3saWym5
YwU++1hmYsdrrbB7gY16NTmbMQkBhrV+l301SmMhnZVxztlKfXm2+kUAP4bynLaTJpWA7iEKshbS
UdSzeGVDyS0G8maKHli26E1iKDld3e2eXanTw8nulixcV0RB3LP60TmHImd0fuyo7zA74diWA6ud
EP1dXLql4tReQFyZt+gkdF39DbS7uss1rouaSaHM8HJg7Pw4p8AR0MXAVsF+k97z6ZQXibt2VKvE
MQEHGBqtqqFPe5QR4j2KmomzoIxGyLw5YlJDD7oXiIvZ3HRdhP6mTWaAcQ0bItRXNWZrQkn72VRp
VMloNQyjGiLB7yNqku3MwaTOgYYtPzn2H3Ud/nfQFuiFaETeyOmJt+dPBxOScUEhnc7xKq453Xn8
txUf+Urhe+mydKzkf0VQWlL6PAA2A+OUyd4bCjqKhWeAJ9DmY/EAnQeCYy2AlDZ1+EwTsxkLKgmP
Ve1MASyDtRYSh7UDUKQOFdiunuukYW1rnQO2L/EUVUhzlY/Fjwd+/sEeX27hcl4zOyhTYFXN8ZvV
bN70jUTVyW1zVS+g+Ve8sy3+NPH7DFg5CfZCcSWwjh3zDhQmkzBztpxn/UitXjyO/l1e+zwyqPel
3mRvHk+E3hj1ASeUfxIOCoFv3dQNkajhdKPcTr2XfLwagfob4JCtTmXy4CajuULeTl8mSbOSKbRE
LbZbccKd/gqX8IpnC64tdf2oJICdmMnE/0lpmPolKnNUjIqj83/+yncQ2FUWy1rF1r+ztoBw+qBK
mXRl21z1ynGpV8UFToOYHtEIDcZq0jd/UjI0Fj7QZO7a8Odk3hXEafX6caK0g2KhtjU5WG5AE3ch
zRdY9QJ8sZWR/Vpp/3bojR24KQT3846T8ZWArAR7esulx5A3RuX0+qLbAqHJfAPdxmZCbSFBPrqg
hOhP95OdJVJY7Xw/kzpX/5N3BpD5nu2byLdq0Vomjri4YvzSozSTrA3smQmeGTc0x/l188nmFQ7M
r+3bo6k0sH+N+dfMDZolszP4rZfoe9gPwoxX9EHTHhFvK6pslaaESA+wmyoGKPQ3SQuOFqZdnePE
SSLx7kNsmWbXl33o6J4Viwp5hDPjluf1H1ElMYGw0C/AvJnWOq7SEgnJFvxiapgtdurfWXT6Nm5R
oQ6NoIBP2mkxbZtNIB22hj/iqrJTSs4wzmOvg1AhClxfJtf0Ix+FJkWwiYHOt5iYG3nyk3X2L/ap
5wcERkxz5wtGmf6B9J+DKg0cqxAEf09W8aZsxch1FjCV/Xzsr6+jN/mFfxDsgFhCcH4VhhtNTMwL
jVdsorZkS5WwmDcwFGs7iscFS6OJh6cs8oyv1kbS/PAyHjB+Z/B2MCvI/9brnho+izUiVtX74CTK
3Km5GDT/PL2xkkJODjC1DvB3NLV6TZKkcCalyoxepCTVQeiE/g8jTKDNEIzm1+w+j8vTLlrtBJTO
abDwdQviv3I6e+ypHhg5mhD3fLStMr9TXMUpkvR2bRWPCxknhlLXiUp59QVXd/QSTYD2fnKpYzLH
YJgP80TXPT+XQVHf+0H8pXNacJaNnndZoYiZ9V9cs8Qu7VYcr1+Vd5BM3QLfOf1ZS11wiv15mlK4
lhW2FML1m+vpJVtrzNwQWYvZU40xfFwQlx9TvPyVmcB0nLVZ0eP+nz5v4UgzM73qiXnitRkgSvYy
z7O64lQxiPdTxPTYCqsvm2tVvf9n8mX1gpqXkIAirHrh2qvP6MMggarf/o4C6jPUHg8GxXWFOetV
xaH0V/gLIKwu3FDH0I63ck6EFZaVWYYFxFOCpCZlLqWQ2vWzskf1Tmw6kVcWZGkdY3z1tA/cJsRU
SVThbQX/Ni2LGgdwx1AHb3Vuv5fPVKO0OmMZPw31KG5ZfaXPCCTy0mcp9rmcWr9IRntXDJ5pp6bt
T/nWnnn4Q+8gcbMuGeviAFyb4AMjk9DxFnq04eS0ZXechZhmWMKZUwD6wURpfjdFL/7qI4KaNvD1
nt447Wnn6EA34XSKwx2Q4CdBUe4OgzfGeZcC4P3iXLrULODVDDhWm8cdG+rc1EubrCOpINDFI6mJ
gcjbkl6RZUIRWdEoBi9paESENfrddc6EcyhulmwJP8xzuNzljDnxLvmPXFbPmy772tc9jDN1z/r9
TEFrW2rlu6YqTK+Cz+ZlwZKimHNy9n2tV4fLzPV2PKq1W9tcpqGkh2IQFB+SoYDewNgfkMdLGxsT
dHfoMAYhgsnacJxIv8KpozJEhIuO4JprWWHT1QCMFQWSDlMee1+HI+PDrZjh2laN51OGPAx18/Sh
/gtGHAvpu8oUW/FGDwkAx0t4zxH73e3j9bctslsjIy9qwFHfyOdG/va3S+KxX2GA2giuREipp+2l
O9S79hU8z/f0TYYg8ZDsG5jCJ6zZ5Dce8kqspm5ZwYP01u5gvKZ80kXt6pFFWICQBEZqxrgEP3Ng
zo48OiP5yKtprLNPWljOqHvkbrK2HJmeUBEZIn7k4//gOk65D7pvHfxNtK+Nn0QmW0oSzqix4Wcv
uGw95Jm3sRMF6f4omKqCwP3e8l0paXB9D5CPd34Etja4GWqmDiOTDKbU1Dou/gfbFq49tPyuV5VC
ko/oM6apVXR3QNslboql16tUQNYD0YIBZRiPxlWP2zzOJ7SOsDDjWhVzCIrj25RSTITDA3GLJ+Iy
3DKLh8tjoJ5gL5sLtr74JZZ0XmU6Y2+9Yh7ZaZc66UWee4bkCC/aGVThFYBPJIt2a/9J7Li7kVuZ
CcWKlMvKmABoStDM+FdfcCKHUejQXZpAE0cwfmCjNpvCeq1Te9n7KP8gxyermI9TODLq+zwKr9NU
Hl6I2sigGLU0dkYuxQkEuiyy/x4er6H56tuRF/DrUhQf5Zy4PQ1m7yXpA46BugvWuhLP/BbRZdST
Ly/zp5QaCfI+YrOZ/PTMaRjaR/jDn93qm4vx4OYznR1PrNCBZf8J3A0LIyoG43/5VzUIHX//OTAI
jqmIaOK1EMgCdCEMl2s6zmwVs0CSrXuDf3nlPLlJSedofoww+nCZ5fDDkr7t2hjiHyPY/2XNITm/
fKzJlvcsFGRgpS3KHYO6mRA+M1BLwC0yBGtAOFu9kM0f5RI1stwK+vC6JR33isyc5vMOyrM/TA2H
z133ovNbFwtnRQ+tGCk/2838THIFSBpG2UDxIQu9HBRtlszzWd0AztaJqNNscOWw3PdxjmlGaVvw
78x8N/oaA8pDMDWpL9kfVmo0cxgKBHe2CbkNoD2YtyIRWQ8aRd39b3R7IygqnMOmUOAjwnAJx3Tq
RKuHzfnJFWpMAtzlv0pv+Bo2IozwGxSvgoxMjlf2/XjK24ZMLK0gfTg/cu5eX+/l9KM81Hctsidv
Sp5HQ3lRj8BlMin/7E+GBfLbM43Kw8Uehe5eIvqJ9JKqM6ki4qe4iHFb9LVXCCEymKS/1SVToFic
0pQFeNa57YkSZFMIIH0P2k8Gxvx0sjP22FJvmPpFFEzW6UyHTX9iGtTbQ8KlF5aJhbpMIyOH8C8H
6MZBDk89UDObLR4Ww5I1z5qqr9xUutoyRC0FcZf9hCzvKC2iPCDcIxrOrVtK+3/xSRCp/TUs7OTB
ZWxdABkbBUVBWlhiJGaWyXdsbmyqQxp9a5EFx2sEoMXlOa1hyMNgyfUovPu9oho7hUgNVRL9AYX3
k1M+dzRZCVp/6nfMIOH0MEgE7Jowze/K9O0JgqHdUmVxIa7HzIRQ3opBgI6AzTO7LxZZofcXEFMK
O5X8dCVSh2WF9yXjG3i5HiJH8HAdhyi883m45h0PmBtiGFuovmWaSRWL7nWjMMDok6kYnKjMoF9v
vWdU8nqC4bPtXGh/p+VSEyjOS8Ci8ZqATcCoyeKHMuOoSMXIguMccz/dv9LUYTaebgOStAKARbz2
PpfjxrDfzQLB6kotyI/mpxgZq8D+GIDy1DwKI12DZPNu3QuWtDB+1qZXNkI+e/WOmyMaV6pS5v4f
J0kXoM8o8A58mfPh82PmFGvAjUcmVAgGzHwP/dSRYA9jzm75418ZTwC1+F9hLhQ49GSQbLwKrV6W
e2d8Gpu3Xujf8kJL7+RZh381WGUdlWKwxKNUVlc/2tbpCYEWIB3yqH86ck0hjtxQ+OSamgwBpqz3
3Rn6Wzfkiw8Yq49mv19JIIhCyRd5mV3JzRvCOlCtx3DUdECbfBIBL8CLA2ZJSA31z9FyFfIbJqCi
7L8+8YDsj794fHOc1386bo/hOE9ymOqdOTX9C1S2/65SqJYU4WHBUCT6ERJHj1PRriUWqE6FT1dm
bXCDVCR6SLXwDRckT45FBxZp/vgs+qcNYE9EDb9g+/09BbaB8vo7wqdi9yAcT4Ux1OtRoHVyZEFv
jRi6nqLaiOvwGIj9U3HRBhDsgfYGzpRQgjBR6UbzyqscrbU/ERrRJmc5zFEVNIf5AHLUjYk0fWT8
rbY/Mry6EVUcR4m0NA2YxitSm7q/IhLwxE7aPxR4ZsxQvqy+6DarFJ5nYX7HplhRexanAoJg3MJq
kMeql5xCyTRu1p3IdAqn3gqcr3zOilOjTyWPEvjHFNEO3MqwL2kxaH2aNurCHsQ4H0cOhSQ2lTXS
BEn1ll4U3O86VAvR6NzyB61fWceJ49mf7DDcel3cupVbDyv1GiJkJ8GQ2jdGIJqwuL80ZIehBI6W
Tk6xiC0krit3WAUcQTg2Qkss7VYtfOuqipD94britSDqPG0Tm5EaOWmVcUltTATxjFmcyeRo8WzC
1Yhs08t6LrWTwy5LMsQkTVmGwwRHWcMiBM7y1C/Tf8Is/tHubkIBCYTuWn/nQCfsh64oa72L3Pxh
/yScgOJzBVbKie3AZBox7+UbiuPqB6zD26VHg7h9r3iLi4ksWdrIhon4HXyLpsFpFPMsC8rIzHmW
aX0BU4XNqcNU1WSV7sIXj59dFtlHeyVNTuX/Ix9PVY7v6j0x6QRlc2NUOLjJAJbbueRD54wvekZa
JZQejhS2BMunuEGCe4/LK5A7fnpHAel4QNishx0sb+5Tdrcc+pADaSehSOz0Ckc02yB2rCKuGzqx
SCVGYuY2dq6W4fDqoNZKA0byznSYQQo2Qf/T6WNz9wv3lmmNc2wzhevxZMkziICjsJycduQUv3oh
JzOen7+0BtxhqfLxBcCYFalE7Y1eDE/bOnoy2WtQ5eg3b6gxwAKzu/kJFTSOwPttvW2A0etEVxNj
Pozoe7+lUQwjxCswKuRG0uISr4NLOGnvQi07eq0Acg/Vtem0fUk/iRcLXE5Tk7SIJ1RPf4fN0I47
DuuLKQvosIm2G0X1xptOUHf8U6cVqw3ezXoaBIC7qc3x8KPT+nfMqUqwJFeZwjPthgeVJptIqIhY
5joWllcsSLKZ/DOsR9QavmY2SXulw/0BraOQW1VcRbjKiollQmxfkZ1Olp+yZ8vCJsleCihkza6S
I423kvflU2JVE13odpGFOQGzdGNgdMuFpXiglR5wlnyaCVNBYWLJl8MaZp5rjq3+QCgtVeLQ/mPq
Jgb83WVEAo/7M6a9sTa2BIPZMDIrGNI4GbhAUa/ILihZHPOEzrl1XbjS3VxrSZNL0hjv66KCiEDE
Zp9wdH0AttlbSGe7h1mOLB7N3U0htRcZ5hQ1q5tBgU0QnMlUZlDoqjQvsNDtPvNwPaUOM7LH2BDX
g9749FoetaTvytm5+ykCw5lSA1A0wMOyx9oQRALRaVeIW3kkw69Jt60Cq8AHHdoxz6Ff/3uB6S24
NF2cw347ecPBV3i6aYNj85VfAmC8lm23cXZrKGayHXCtBvqwZPEV2ZkhqDhKDTMLUbCwD9dpK5pP
sPgwRnyTVKyXzNPznEdNiE1OiNIsOt8U/VUFNKyxns6qQa769fbh/zpmC5slg4lxaWaDh/RTdWC3
14PmW2XmyiyOsdtqTbbwWhcP7NipYLlTiPynaR/WNMvIrz9YrwVVP0qsESJ9+Muhml9JgrEx9fLl
cmFwQAZAzOLyQyp+cOd3U3+WYIJ/FHilTYbNxEKszyEgVYv8+1Jo8wH8VDMs0HhCunaiUfLQOHtz
RgSm/htIRWsEKrBlpjsZUUcnaZw8idtNXOCeh+HzVhXm393K3QSGUzn/aQ2OImDhkQEZVlBy0jpF
NxSRLOs6fU73ICMo12S/sbCIGxJE+XIMWXN5W4M709bKEoYG6mo9tO+JRmY1KYTxXexjojKsBTDp
NWRqeE6DfEw5mNy6tt1Xx5YKwk8xie6twvZPTE4rglOuSpJo8SjbzCIdNvQBQ4VlupNlzBAABWiX
i/JFxAJkVEp27hcWBSFWyr3KDEKJz5/X5xe5h7DFLPG3LZ2Vy0oybF3yDOui3raJ5GRxZrMwZ8kl
FaeKVuq25Cb5ScaEZ+mxdroxWv5IUp7+IVTrNHarWw7nMnIFyryPLBJVCAtRWgxigj0QxHBmz1Nr
YpT5Rnkol6MP5EKgM62FflaswVnwqb7HDNuw1uSztf2IiDIfklGdf8u0DUpniclE2FV7+InFWFsF
Y9efpy1IydpYHlfJ2c9s+2XtuqNpKOnb+H401Ptm1PdZT06HIxoNi3enYt5l5QvwKwPHhEPwX6JS
T/Ll7G1uUjinvFw2WTgxc6PIi+xefSnyqNiZJbWUPf+Dj5aWQ060dUHGuXPmCQxSV4C7uufg4jjH
aptZ+Sr/vLrCs55tLbpHQGKq8S3lS2LWEUpQwrSrqN6FLfbdHm0trp7p9dT4fH7Ye5FL0xG/cZPe
gH3z084RmMRLfSuXfuWJA/NNJ9TENiLEJFwvB4akGwbdjaGxfYnJkPMpj9aYPcYp/tZNnaaI9q5g
JdB42emaMkY1cz4uJWOVXj0jpX/fVS77kuk0ItFANfVL8QavsQUE5S+q1fV1jKDYVOpPt8XirgCT
CXyK9EF0wuHhny88MFkAlON5DzE0PQ7MkQ864/490oMtBT6p8WGz49wCUGe3xAnjbKw7H+joxHoH
mz9YsPyhAdAAHfnN1SKbKtRhy0Z43RoKAGeeF7iqmWg8pEBwDDsVisT8X6QAt7DXo7D3Qw3jB21z
3eVimF/vdLKydeJ8l1ZlbFgO1EpNMMOZVbexT473EkIBP9fJheDXr5miZwKL3Dn3fk3nf4x78OCK
v0HzNaUP5r5Im03RuZHkFvBfcKFQ1EhJT7J1mFcWEnhhqbOBBtSZOUQA+KcmnIClZTcC7Gy53fSO
mPQj+ONzl7I+cYccPcZvrhLof36t/6DL9wMwodqj0IYr6E7Eleg+RAc7yRfpRKYyZS1OQXE84bId
7euxtcIfR6NevQP0LRAc2t7vPzc00TxYB/nnyrdqnamqVXr6rKWnr4U6ueQ6d6fzThHhi7J5NaEL
ISyilNIpgp9La9eoDS9pa6rggFI8Gd76lAUXq4r7YcRRmdHWjLAV4QI0XqAcBwgMk3iOanu4ziWp
31WmTKiDmmu2xN/vM/l0EsUDhph2ONDHoE+s7EEFfI24JARFDTlkMFRsvPOd9rFHatp8I09V5kCK
c69YuwRV9Nla+uDpHEGHoo4cKngZ66OodcPiW8wOhr3uIQyHJhppHCazr0yNhDTFn5WSFzhGT8Nx
AuNhmxWjdilQa1MvP/7iwuKGD2febETqpXYPd4Emb62/z08GXwxY/ftzUVyo7R1819QDmkPRnJT9
ypHQ84yB5queJbefc4/7F1txmOmA0yHkK2S95QbbdUmb3I1USoBxV5ri5SyK3NdpWEfwX6wwIaX+
l4A1LyPaWG4zzTuy3OZmdN96RP1wv3ScUG1/x6VfB1qt6/GaGh0gdFbb9pRGdzglZfYtA5ArJYDs
pD2FlVCSpdJACXo3So6XqfC1vfNmVX17qmDl5Ry0cFB3B1xchjdwOJTbLBJd17IW3CBSf0tU7LPP
Rp+E2u1Pl3GGa+qqAj8SgcpfN+86YC1DjZwPSBdThk8KL/u8IptfhC17CYbwxkOe6D+EStuVPhlk
7Bn6qxM7LhJ0C4K8U7zgnvEqVGev+aEjNdi7W15s+A+KULZsaOVLG783ZJIRuXDYHWhc/zIkhLNV
hbGXda1utOcong3pCIi3wil7uDZpnpU9chq+q4ndITopMS8JKdHCgmJVMuyYKIBWG0kTTXZ/O6cL
izvxbYZ8kds9eaucA8H8u22ogC0khYhCEru84YHLNboTJpUmWbGuaj9+C5+TbM4NErWXMPJdDCWU
vUToHAoIyOFMD768Z20OFGedNgWCfmw78rCWKLsUbJ3SEjH18u8bS2cw0uAivkVRQo79IHJ+QzXl
hOHL2BsgmqDUWnqrFXx8Jc9F/cUOyOTVRhje45JEv1bG8Uygyy6nvaSq+4VlLw2X9VQdJiBsjUhA
OQLLZZHXscnydtaLRz7bZviLWL2mxF1u82VTAusEw2fjpadj/jeaohHRWCGTVgu8pUOKf66C9jJJ
2rVJeE15W6PcD+QSd/ARj2sUwLtVK1/dD38xmcFk35oEBLtO231aHeolVpgrl4bzOpj1s+QmT61z
SvwzTzb8H1rrhCSxPiTOs8TvvO+Lz1Na49amknyrypi5IX1yHoGIYI/6vkxP4h/HuBSUvGAJB4IZ
bWRsqItgCwfSN9NKt/5VVEMpyG/pvhEhhmgDdQ5ssyV1fZ5c36mzRhTi+w4kzQ3v6eD4lFFrDJFs
AhaVzuIbIhcGdz0IkDHqcTyFYn3ARvcKept38TbS4sDeV/Et96Gf1rzoUxiZrsR8NVhcP1EwcSxa
cqcNIB0lJVH7s3stzIFOfS/IabrPKhWN7fnOjQnfJ2XuXw+cfO5hdAb8eeyL86gGdZf87ht0uZ9f
x1Ehl/cJFScM0phqVqj/Vi0EGYNKfjCQdlXbLYpm4WzDz8VbXHYW3f75dIpsKzgX6eYiA56pMhTk
Fs+X6M5RX7J/UKJ56wToo3OlJ6RpAwsfwaH8GaSTepNxnBVkKgw3EvpAwKfO9viIt6Zo067j6Dr2
+VGaPTNoUBjEdy1fazNF/0d8EfWSbbJ2ZJsYlJsq7W5RUvCziqA+yuiDjB4mqUa4FLr6I6STFvy9
mkI5OYvoaAvGCM88KgNKYllgtWQ2sVKE+97y9cAfsefTaDRKYpPgOb/EtPVxfRXPUaVxVg8ZqCdP
JeFeBd7Bu0IWZ7+uLGEcBJ5BDy7AplydUYkbjyGdYPl3tMoZ3P/A4L7+EoDVYD538+DeCeT21VtH
vGmJ6s4GvnxdKDwsTS1k1A4RDsnEimcLs3nfT3fEQRjica29zYOd7WOuwWukM4TxmJw45d55eT78
0H7ifjfS6ccc6OEgjdgY2SUzzkpUcXBBt7SpwPWKWf1QOjHf9PIwnBBr66pkbZAoYO4OlNUK89Q1
wh5ZKa2ggbC2/36FAugpBz+Z9QhX3RGNAksA9COygWJJ8MK6JCY8ZS+UvG+GZfLwKHldUavUZQsz
UPcXYG1hI4AVml4Bugeb42pqO53iyOVJumbUf2H1ByfSMMvIFr2Y+gh//j4iMovmV6797p93Xdxc
E7pDycMlTYrvM9msltx6u8VkIkrkOJH4OyrQ6D20MIRuVEYiOQNYp9Ti/hD5c+OSVS/N1VL5tfQx
wi+gDtRh7kALUVUu4Czf7dvfYyQ3Ux+ruhogB1rz+pNPLF5iwTv9QGi2+c8wZ/ew0IAzl+mSx7IH
08LF901esLwhXHAj9jlhJYV/2kq55MWO707sWYhiRyNQS9+n6rxejpcQk5BYMswBjjHkVk7xI/u0
4H7OfO7SNIu1mJuNF6xSS1/9PQPSM+b4y7EqOGWJAqHSq/sI8PS5vBkArH0sH+8BieeXeHihiFkl
ivQlodLlZMybdCyosCHC895/JyFnB+cAEtuShjxmL7UfDYKJb1OZPda596YGQ6w8Azx/8dEfS8C6
dC5B5lCDLl5R701NwpBPzrsnZWCU1NPc8bomJHQgAiFYGqy0sdEUbpvDhUOVNaiihlBLgU9SwTOP
bYOUwnb8ZlRRwhYJRVR5zrLw5hpo9PA1pnuRyTLd0rHh3jKvNHSDIl+MA2ez+uei6HJV0ENubq0B
gNbwykVboFNv6eUnSIdvWNhmPAmUa1gUCEFPlzL44kBaLSeO/fdbljIgchH856egAp2GRyHr7FXv
B5S/1a4JcCe9AeT3NkrXnAmMFc00nxZC37Iv4qTwNGq+fR024RMZz2bbTe5CGkTNvkqSf/VBjZka
UvG4dBtrgv6QEPBZ9YyPI09J1YsLlRE7GcEui3lWk8oKo2cPNW5u+k5YH5yzxQN7VRNtrv54aQXp
pcMo2Zj1jNiFlEkfiwDPUZUaXhmQjgCwp5ptwpSR0XahqJ+xgzmAURLIGqmFKPvSqau1b4xV/BZj
wnwb7eCuHZQx0i4s5LRBRWmjy4C37RVon70Ga0wDo4gdAu9SpefjhVisuC97lGmoHSv3HsOp8gfo
vGm+U3882JZVMCJvB2oV15p+pkB1I4dwJgWnhwcBvHyl6kAsxfcaxS6cdpFPOF+bOvOgteSp0UZT
d4y6+Lz6BdKVBdzGY20I2Jc/Kert8TGQm49F3sUon/U5m9x6yNfMDWOmljltCKKkc4j9mtmt86mT
SJMG7t4wRFzIHhMrHpchqE+XbCIdMElXFUqIGANmnyJcxYgoC6I77uRZgAgQM8tbV3164zhjyDJ9
5c9/dHM8AXdZhGbkuVmplLjoZLg4j32B8p5r7HZRhDS9483LhiZE1OGtD1t5njUhDulZIWOlJv/d
EopXvta76ZJVxO0EYxkhY7ugq8YvkgHK/iqvOrv4sZOKjJovpWOfdq6wS54GKt6955Jx6uZI0gob
NAn3htD2OYotpXF2yesczypWPcKdlgl0F8khQMrNQw98l6y7X58lACK6mw+u2i8zG270cZtW8SJf
N+w+J+vuy/7kAWSwcjLxvicOZO3aQHhvGslURTQOF7k6flJvgyZhyN6M3/7f0rLVnXPELG2p2cLZ
3SxX7PARRS+qYihWf9B5N3A+CuQR9ZmHqMrYG/Gkzk6kgpgsb8prTZmobtiY5wa0hOsCAFLcHdg3
EW1qdmfZqndwKew5JR2Q6ovbKvD76mDDTD0fTceT//qlTjHO1jB7G1culy2K/dCOZOn+EGQ814UV
sgknJtVI96afjlS36NQnW2zAs79KPlgfIroF7xiffNLXQC8OJ+q0cJWJ3yrmoc/CT6enQJ8ehNs2
h3pAuQLrCIw17yQLoOCO/NHJuGihQdc+BJCbVL5lP5kQp1H/gCvU6eVfOrTmqq7vPXNLOfS9CLQb
WOVAT63tcZE3et1lJtGTufMGIgFhU4gdW7UCV+B2ImqkcjvSNznng08V44Gz+gtNwuqo70SeZVN5
I0ECfHEn5ZG5ZA9IoFpCq3KpRvLK8Iy6VjRc4+yZxSit2QuGGX5N7j4aHw8xKShsB40N5CE2jtVJ
OelNpDOhFVDU4gH46KpcaeV8dXD0qZY+2bH5W4cBtdd1DLdUN+hkuk0NKpmcGLzKN/Z5ZWlv1ApZ
AtgXT5GWTTXkG3tzUomFRLD74X84/nqpGRCH54QxGA1IAoX94EJzTxYwZlHL0Ip7MpJ2uQR+3Dee
Cd+KlSkTYyi7Z7D7Wya1Q/0iFcAIm5BxQZXtOD5e/e6f7i6sl/9E9PqgvrL8rois8OVQC+dij/Uh
uzTPJ04nr38WJbL0vxGlFXeRIoRnaa9qa6stbBpyFpBZ30DlT0dADLkC05y7o8NULBMgJx+YG31D
OdroPhrNQxKIqcj02v9sWRm/uOYL881qV9sMzSQaupzAa4jLhv9qzjeqRFGpD9XnAxuCMDtLzfGY
MzOilR/NYoOQiglEZVrrrJsuuKUY5FY3gD7exqNlDV+rAhGD2ZAzRkICwJTkfQgcqrjh1WFqoroy
Gp/NBJXBcJjQkHSXJ/vMIR+LO/K2wEWKF3a4O7T9chl+VhTHm8Iv0RAdKzXVd4YKdOs8JHdK0TYD
TAgdAijbB+OlT7eAuNsyjkvTCP1hO4XaBL3u86pS/93mtdyIUfks/ACRWt6eFrhNe7zfh1cVYQxJ
+MZYyld7AC4TpR3IoKAI/Y2zwQMocnYtdropIixH4e9BPJdq1px8HIN9SfaocEjshf9ss6nfU9N1
UlvNw2mBBrfAF90CWmar7IvrGEzxIiGGayNlzdwg9HyZNrvhTPRJcby/8H/rM+NPqgdpOCw9QDUt
dvNmPzUCSLDBDXfqUaofrLIw7EpKQcz96Ra2DoccqVhiozZhCa3cgjSwT3EQ14nzb8hoE/U4aCw7
opzXp4vWRK3MgQpLO9JBrE8wOp2t1UvRMQUhN8b9n5mwTDaEZwn3NCb7j1Q35XkAZ3px43tsoBcL
liSjPgfjDeOImIVp6oz/KnTT5I7lgfErLFDikfd0hidDuGdwWfk64/s/NnY4d8y2HNQa7vOD+kU+
RYj+Qfgf8CJipyVZou44vfwlG+Y345OA6BATc9u5PcDKwvF3MYQdWuWbrX79WeKEZWqLuWDRQGHX
aaGe+7rWkVbZYGtQhx9NYMlr0q/tBzXZ7m5be86pyB6wng85SqMcSraed9lde4nyKrin/vtFf41J
fQnjM9nLc9kcdbNVr/n+cUQ/rUxjz3/BMa3cA+nFedVHpWOlytIxFfDvL4pZ3knKNKf3dUTg8wuJ
gKBZ7eaaRROD9uTLZQKfq1cX5Wd/Cq0PhrKMUS+bjUznh+Q8zdMkS+hUtPakm3UE4jLc1xnRbHPn
P0xXHVLnbFCZ4xXORn1pDLvXwCiQh1LwIRewE5xBGvr9IyPXt71zzuorxU8GW7jZhd2CcZ+QLugU
8Ho2JxiSbqDTVsMUueeP1M3bh2+20GuGx5sIC6UoRtlmuNuWukCkzXr+808Jl456pjzLI/G4rqxX
5eZTBlXNFzLmDqMEuxzhTug2V4ys1zrW9pdRADblBxQOAMVvWCuldTegKlS0MQpyGGa8L6usTw8r
dN6cIPRkPiKiALql86GkbFInTX0Kixw+KFcTVf0T58bQkxJeNSZusL1Ra8D+COSXgVqOsfG4v8u9
MV4ORaF7zlh7Cis2sIZzLVa6+fw1HPuXeHppbHZ1dei9A2qpm3+aW8/hrHPmYzHRzh6XhH/B3TyK
gSbB6jqmR3AN6ufQvMW1XwuIsvB61YNtwajXc/GHk5oK/x1k2SyT1okkVJag8q/ELVxY7uxPmbil
BAcGQv/FgfcvbFR+k/Fasvgm3MEzd1WHn42a4pgYbJx+BHcZNiTdVhoT01P6vvmXhMNblUFRVwZ7
DNIWQglyXvKeWMB+r1rArCTMVRTyhEtPHMrfpmDEbdwacJqlCUm2qRRAHTtO7J04AnkZAqXfPQNt
8KRW3AcobsE3L6OCZP6AzQX7O1vA1iePBpftSP1c+EqvBaKIKwZm+xXW57Rjy5y1JY/rYZrab0Nc
chfZARrkVl8XIUsdHcBFeIIYPrSFDjPN0JVDcjB8yOwQFTpcNrpN7xCYAWcLccWVQw1upkmRj/yS
UBPHEVOhOqZKuzlkiudW81N8bneA5vUbADGZhVKbP0mvmOusp79dP898lE7nMVc7uTNQBNTa8dl7
hM+6zzOcSniLjvR0EbBrmbjV2aIM6dZ/O5+gfamrljS2f7YLWrnDcoyy3VaeGzMubasyGe6kjVih
ytuOBoigBCVEkZeOes85d/fj24eFAiOE/qLFgBDQCxYwG5IkxaYjkfm2WCSNxjyk8RgOQNAREJ1/
++uVwoOuF7adTNtfhk0uCQN17/kcJ5gm+WHgIsS29UdtsZ7cfFcMXp8TJyWWaBkI7OxbA1m+ucDq
mXKFb4z67CkM8BoiW/YIIWh0j7g00433GMkijzTqyGhehFkviauXSRcqxq5ObdmbMqaOJ8Zpp39/
nDwGjZZRG0Kq/gn+7C46aBi4SEREHjMDWyLx0ADtb10JOYb7W3FgwSKbLdmF6E4MbiFtn7wtsky2
MXS2eYff7Dp7U8hpfs0dtzywj/iix4QlEZPdEx0uUjvxIlfDhN02D2+mpjwKQHT4vaUd0DmZ+vKe
dswfF5Hxs+Ejz7bnJ28Ug+9N/6I4llPWKfYOThMQ7+gRhZwPy7MvUEC4YQkecFpqCTJlOsC/bGBS
6ohFSJwpDrIOaweX/kX05wjJiBseX4n1wOIdiyTZ6ikw60KA79GxwsjZ2spO/pWMlhxBdCfjDziT
+8RUYG2Y2nns5Pnggak9/hwnWUWa8gZjeow6asARl0x8qskgKxjS7ApmKG0sDXwB3dxrHRvFkAr1
r5U2coc7H5UH6bL4hfeqA/QOGX9ATStaGioX4w9f1jbO5AOY12b7wjpnzGkiZtCb6Dy9Peet8MFC
YgPC6JF4lrmp3nLPOAMsJ7aDacNfXUCOF2yA24uXFPB7nNGlNVod585IH5stcGQ7gd44YdkVFPf+
kJwdvVfTVgdlxNsJLXXmdJiqIGX6FA1j0pz3505HPEHCy8kGkwgjDssXwwuaBEFG74yzxgT4et15
q3bNypO4yP5BzcI+XVJ2zy8eq85wuLWlHzkceKeXIQK+rC9fyAmyUpdfCn0z+Nb3y9bhfbZdf3Eg
In/z9B6PgssqGZY5Vn9BKyKaTWT3kj1pPWOrzLYKcbEwiyJMf0hsiWzW66e7zSknIHjngowcM0VH
dZ1y4JumVq7Psw+gy+30Ro965wVF1VMaNy3Awa37uk/4QnLBM/OJRDwqaxIoLmIygydDVhxoreB1
Qhd+Ji+0SFndadG/o4ZPGZB6k7hq9VyDq30OXLaZMVFVmk+vbZ0uoS3buYvZtfpqKvOK3ZDYvWFj
AO6D21VJTIdHJoXpHY7NZdUEUKCtvWKrMjEj/HGnwQzdox5wLJD2rtwNnCqvXxhvyhB6nQBBpEMQ
A3jqSG4D5l1vnLyLQaabhrYVcjCBjBoiQwScKHskyEpt5jB8xgqsZ51a+sglWiavBczildi3TJ5N
jFncuX30GG7BvwMsEDQfQ3zAR/FH/NP5QMP0a526He54NZ/lyN49igL/Z/OtqwaIXj/uFJYgxia7
JWZ7G6n6bSlidU6GLxV7UGYPHIPoRF/piL7zq3yA0hgQClCNgw7oHfdHBsR2rep4BIZZRPjaW8Iq
S/Pu/rnBetvbaOaJln1C8GizoW9PsFt9xHL1DqvAdBdKqx2fy8gUvPz1yp82p4ONlUz5Kx7cKh7r
pIVZNSxEbO2/EaaW6LUtg2Wyn7T3zF9cCoosYkSK9SuAqJN2uYpTCH0Ue4HR/xtXxCBcob034V+z
hNFOB6blE08srMRNC8whN0kXL4eXtEf2RdcL1LIJ5XAWr4idVQ43D1UWr2/V7cyWEzRZR55E9FcZ
015hMKp5KDSfJP62D9uD+oQ8Pd5Oyoy14cNDHqd5mzHZm/ED2IujrHSIIhRdL/v0i2LQ2CpB2bpL
S1OuU+rs1R4orGdcMD/CC+YeYGCGM4UGom9Wc7p7gUIFP6MlZoBlS5W1QSVy5h2ORijjlu6Pkfd/
CywUuslL6DVdnuXHZLRHBLGjKiNFhnMti8y5SUoS9Wye9NZ8zIeGxbSS5bd/4xpPmLrcJ+s9uppT
9PVbp0qZNvnR7n8niIskLhaXMk14J/SRJksKWDZoJG67thomjRcEf7822TbZqgLjRZw/MFXWWevi
eNJMv6wwZY/jxOgJZk1zQWI/+Q4IB6ziXANM5I9j7WWB7cr7K4INzAV5tfeMLBzmoGXKtco8JO6G
QeDkgl1syHuvVW9af7wwUXVJdJR8IOLKJDX26IZUfdy7PGx7cO7AKHPXnX+Fo4lW69sC3SBSUS6c
QJ/vXkkEnoYsd5G/0IhkSPGJHiN3w+rIPyZSNDjemrQXXUYvkY4kJkYz4ayN6iHtOovJ7NDDXEYr
KvgUCLJwek9MkAawUv9gTLlkZMl5dexvE7tN8kTFVt+hFWv8FsSW8ISCrwSnnDRFhG1N3c5+etjq
mxVMWi0gIqEsxa3ukZnUbuQsA/wo5WgxoKqO8pUxlmtd2X70BrUOECLLXfFlfmVF/UdSrWd/pbhr
Ca8WGTC4s3v1BWG7Y5+LsKGOL8lXkJu7USTxyU/B0hlOLdlaJfkjy8ldEXZmp13Pfqhb56J5xbL3
nR2AratC/H8hM4lN5kCTDxc9y4gjJwTVdC2Zpd/O6QtHrvEnQEVH8xmZSP0Y6vtRoSVvtSMCZyEs
vkuQW9ZETUaIP6qRuMY+NG/WT9rtdvE1PZdk8v1dDUkZiKEwqFYWHgc7cFJg1CwNBsMhBPXrRj16
CxA1ILsINVPp3skP/DbMtv1ar7bfyMDiTfKO6GAGqKu2kL0shjBlMCnVq5oBMcdgqSW4soQViFs0
Uly0Stt8SCMsooN49hFK6jRtrqUjmJhBlCLRD7fKlnWvM/rSqhJ1Q1tyTyYMgB311Ez9foSlBwcL
nSYgQdkw417vEqhOvcW0RT6Lc8q/ZJqYAstYxHLHpLQYXQI92rJXlDhwhzuOjNvdhVhBeLyw+xQk
nQR/gIIQ6ZxABMa1UNDYETVCDk8XKDLDrwTkaOzvFRQPp/Tcst6ZGxZMvvksSPq/D1ugsMhPH2zu
bAumyVV40X50Rhxf2ijxS9amNXD7M+jdx3O0tnV3CzyB3bdcT/rDkOXZE8AUy3f4jI9FgZ4XakyS
iYR6VXMApFoSXbTlheNJ4GbWgdSQtkCS9E9ogRYpCACC0/lsAkYo0lqdBYEk09tH4PCv0FXZKBOm
BtAXJFOZMA/+LO5DOpY+6V8ReSD2luXNpA0MmbXhT5YdOXnVV3FOilJNRQOq+djwQDHkkmx2tciF
50lLxxbu9B1opNZSJ1SieJ0d20A7kKsAk+fSKahjAJgNPH0NQOQJuU0zeDb+yshirkr6aU+5ymf5
HQcS4ts6Fm7Hs3LyhgjWJG6dhAJ8UGFrrltxrbiFFfSAolzpYxREHE4LLVYnWSvLObm0fUYs6jLG
7UOMJnL+m6fPWosLs9y0eLb4j9G3T8qnz1y3c7Dh2Q369wkJi3mJEjV4Jtq3t/QoR6ty9liqQaQ3
zKiJAGNfwYixICAbhhYEal04R3UO4sxR0hpGZp77G1m5Ci++RaEblmkjqZbkGpCpBdHwkCjDgmjf
G12kUCVqSq73fca8Q491dmJlQTf1Dnpv4dDCcsP3ABrSUl3aOEUfyg0S6MkCnmb+UI/2ciQssm/H
gdbFykZq9sHjAHKd/pRHO/VBY4kR82SGp934++DIJuAs8UP/UjQCcXqEc+hhL8vgiZkjJ4bHUTH9
TFwY7KRH9rGnYn2u/WvPBTIkf80jhgZLfW48hj7PFWztd6ozB30xQPNzeGvXqneXxtBq0JxDpcuR
jzwTmoQu1N/RlA/PcY+1/Rru7hlu4i7T1vS5+xhHGKf/WWS6Bq7k7gglqP2rMry6XDNAhSk9vwsP
BHCpaDH7nmzIHBqEcojtYV7dzewQr0s3J4c4BCPTEHZblqvXPRvJnLG47Q8BBzML2pPAp45YQAak
L/rGqeOVZtWY/dnXxx7M9dwWVJ2MrOqAF+HhvyFGa/In+oiSsb/RZZRorIJkj5nJjmO3qhBp7d2f
4X3n+Z2mzHksJ/+gifYG1y3Okw9BmKsz4tmC23qoNLw/T/rq+4hdgaMX4OroBMsVlMofQNd+BiJx
pGENLfYh+ScgDAxUK6MwhjV9xBIzOulGSFrVoaZf94WvgZr7KDZeH54yPG/rrTWmBJ1rVaWoDSot
6iW9Zufwpic2K2Sv9Zx1VNT/bl84R6oQjis1wQymaeLGjavgmyff3jBjxW4MUmdhqHkdN04nDQBm
y95jxfAVv+3bBU+HFNvEfCm6Zs/iPwd1Q2ZBXxByyMrDhdGUUD4+YyNTA1pVhbczceBlwsM4//NA
klhZ3ogeYuGoWJhimPptO2aKmloBcel08oqPaJU0ChFxk19fSB+t6In94fAFHhecleIFljUqnYfL
J0YsANJ9lnimnIEygAbhBZ5Us5Iu8304FRZVBpaGe8zIBTGboAYOLl2XzWRQBxfIBXYIn0hTlP2G
ASRFXSRykx3uyitK7QrmJe9+ZBA/i8eTsdJwn/iGfbWQBjCgYLFhKqn4ONntR9HBEQ5K8RQ/tbhM
owPcShSNrwcJc31PStG59iVZch+r3DBrosYBygO9l/KJh3VZi3CzwzBnpgnAgDDe4tOC1c7H5Low
Ceunxr4WnMzp1Eam3TUo0y6poaDqETdmYcUE5pHONjMmeFb1gkcDt5uKBdmfptjopZNrV566mCzm
P+dKAlaaE6ZzT1nXUtWStMwYgUsHgvMfK2P7o8FJBcsYteVZPOdHFd/uBIRM9A3qSw1qYEqH43cF
dVylxPPMVPF+3Vqk0S1QOsWfJ6QyuqzFp2bwJtLXqUMCaKP0hGXc5CKzV1jdn/KQ7ad6XzTUWX0D
D5XkX7DLCXFBulE/Hb58Hztbc/wmidqHYUmjXrHJ+yXwcD/NsluYYx9eE/fpUOTVt8g1GvSbhbKM
S5e9S16fWLAmoCZt/zwGOWBvpRfmreO7ncxd2Tqs52qNLmy5aivAV2Bagh3susVMLbkaaOyc1VoT
QntAtn4hUYTZNHlJS1XUyYgnaHTyWHhAz+RcVCEQB1oYFNZfsfMq+yqPTqmnmmmaH78mpPwBLG9N
qqcFnsx+RxQCyIVRRYI4t+sHNev2aE5usRyrhVL5OqC99Tts0j2LVZnslxr+UHw3aju3OQlm06Cl
PypUU9lEbGW/1RPxeD2pTmgJwN/ZU+Gt9fZh3jfBqUzs4l08ohUdD1Pmsq1sjNp7EVuZoi7iYr2a
5PKUvtd5DkTz4NwY4fF0cc9/o2TT2K1IfwO9L7sGTuA5LSv2+Tm9T1+nAsoH1x/m7Qj34KN5APE1
n5jwMJQ5uYW/5rrrTCMb5h3ezR29jhjmUTvlo27IytPP2bIuhZ3Ul3bNIrbEa8uuUy2nxD+tY05R
EJ8jmhqg/KRb84UMjkTwC3DuXhgZ51ljJb+lvyVYvkhkcpMX8JH53e3r/fEqhm+4i2X9CvsDHwVl
tRhNbnRJItFFMeVQMklm+S2k3ockmFOjDaVBwZcFPwdIvdG7tJWNPKRg7EEe9Ehx6Athe2Bob4uG
wDghXARcvFH1gmzXOsVlJUV7fKZ5pbjOAW99olu+gLMl5yymzQyk6Es459HVc+Lh1J161MPXvIQ1
TxQws0hYQZ3GiglaqQkyvGLGU2++J957y99Vd1EoILpFFV4MIAjYRqxoCPJJ3tN5oHXieB0vP9/8
5c6TG0BPOrfKd3uwtMUXCqskJ8XK01p01yGPXysS1VXmTRPoEoOqyeqbfF0hGBtElGCEW9d/RiHf
Hf7eMcY/dX5A2U9xyRo8QwLi6Q2+JzxLLQQuKYTmXwyFVbUJwAF/b3NNm5F3xDBiMf117jXdni66
pwUZaYG9bgr7fWkxocSk1DFpkrdHxiP///q57U5oOBehQfp6VXMzGQpx44lhCdLauWKErUA8hBT3
CDsA0qpJOinQO1q6uxwr/dJnS1QMf+mcHKBy+K9oL079M3ZKppRHZf4Dm4DTBLHnn2HNQeznFOj7
kQWWIb0yALBtWfpbRJaI+VreYTaVW6a8v7zW34j4GCKQi7kc4gYp1dGB1UisEalObw4lcrCOb73b
4jZijSSSPF2xLPn084Vw/0qRur0+xS45Y4X842bww4CDy7t+CQZPuSBbsIAlLq9gd8X6HYPe4KNm
ywBUpcDvpYflOZSNv+Y3LPImRXmxkhV5EcUScrXjmxJzqpMce6RzN5lq8nOmwAUfRTZIeL5kHbAG
ktx07hwYKfDUkSkOn0490FUnBrdUS/ski1SZ8wjJHYBdD2GlyxZpwhkgEgTarfS8qfyx3YRfBVzS
N64eLrmqcUin/W7fKuoxRqV1flmJqv9WtV12jfSTnKZ7y7Y9XKkz8iybsshI3EuksJIS7cHUBgY1
xlbhMzUBqDR3tCk7Yh2g3XDgO/ufHZX3KfsN0V9OAXBSKQxtgDBLOzFedm2kP+nLy4K5bGI+PKm7
IVpVIze9k7abPV1bYROqJOMOpON7B3rVxhsgt3h4UtlPPO6B2bZdfDUKheg5Ea8g4Su1LpS0A5TH
tBpO5wI8akk+Ya+DAdtZxLPn9aohvtWqJSkK1DzY7Umy0PKLX5aGIbRokPXvhmSvNXa2vzteNG1u
E+5603Vcg9eO5gJ6BewfR9rPNN8+E+l8sra46F2nBj0QtGT9A+HRUYBNiCeyk4KWCnyxhxd0ZQqn
918Knf2tXzuG0EHpGY/7sN2eXdmpamtpJkYBU+Pqdbm3OLYjpUGUbWuSK5cSbtdokAkTZd17+1F2
kZD3vuk/8IwHKyVhRIDIiZuom0kyIXSUpFroFCRK1MaBSadMzOEl3L27dxA4qF248RX05KFLEuQk
BVScIK4ZIv53wlpjXLnlOpUJy8bSHt191GRaPvP7nKTz5OgYP4IywyUMjTQizLIudcC+FShhfFgF
K3wzvxiIUQmdCMm7btwwjuI0bN7Houc9jwK9tMXDZO5FWfz+tOOeQl34EzITHERqcttGuwc+tHlx
OxmkEt0qe6D/YSAs+leNP/iuKZDxSSVVY1gP7Lcoy4D/8r7vZYTJcpXayZWZSTAOArzU/VQwnYW/
tqtds0VVRu0ZtyjvHH6Vnlk7hHOxOuwcUqOqeEmc8O6OUNGSiCar17btD8QDI7FeiJdO5Lvg6brW
yHt5/H1dbtUaOUx1pDlFhFORcXi3CXmwA/91hUdmnmbnS7fPq702ZDi8zEaWlxs7lTnnWrZ1/ixB
cYvH1x9UzbH1jDMWrltvqfxaml96LmlPxaznpg0jmJxoCeabqVHZ97/vcST9L5t2A51faJ4iXYgz
50EYC0oLG0kbhXj7JqBeXoE8pQuqpMnv0w+hdwXVzaDCi7TIjvLHbBgzgHqg4hTOtcJyooAKhPOE
c/7g9pTfEs017z85dwj8FNZG72PnC4VL9orlLg08Ua/i0xSMjuMhGx4lBw8ZFRT8fkmWcBgJnsYk
HzIsE6/FLCze+PmX6DSoyKuMfcZ/b/+BRY9VbqS0jJXSh3Lq0IyiT5WDL8nKD3JqcpIxSOYXg66j
YKvYb0PilzEZ0ewL3YY0iyCvBN7dnzdZ72VnV1XkX4X3gIUtAco1bDDBtFSAZtN99RbD1bJAMQpn
n5UwTzotE6Ivy/m9lWbFYC0q1TS6y3OmtYr88kUzv6nW5kmVUvkBrTSRAETni4ztiuBy6EVof4/m
0E9my/EBvdnxYmPDAClyK8tfYRalN60GE9as50zqQiM7PCrXTiybJRtI2apEAJRXZmZH8wNjhG5E
Vbk1DH743b6VNgVxcRmMFfFCfbLG71WjFTXE5Hx6MqdppB9/41UGFlKnbyvSTzewJRltZMNnR7YH
+2zg1bTz0d1tIPQkzWhqVJOCSq0gCLPW6mg47FPGmQBYfMSTd+eF5U0vQfeUMm+E5xr+Hi5HvgyX
6gcnqQg9oyB9YYqCcRZHP3vlEngV4eXGikvkCjrjgvtlj3TgXUjVEK8XxbLf+27knLxvWK6kYmy4
dU4ub6NLCBYMUPSukhK5EOCuGJ7yIQ+8dSXPPO/SN73WO+hZJhztOzV4zeQG2S5o/o7qxy7tCrgN
XAATAzUm3xMxDgz5La74KmYi3Mws0oRz49YvbfhAxfi4O9dkDeQZplZHeenrKB0EOBlpu5W1y3X3
4kh6n+BvW+50YE1JdzYjDIQRaJjQiIIb976RIpzLuaR60hzczdFGjdP7p5zkwaeOsrSpEmMAdobo
7ish23fdMmek3qEfPLRODRlyO9gvf6CTFNBI7i/GgDPYGu3fXGDR2g9TO4wUNIn0/V3Ze2XzkqQr
T0FXLGpVsp1LAVbr42Mxzj+z8WpBOYFMlv5Ts0bLUNyUnAubjS72Ixh9Cikv6CcqjcY3SzRrLQro
D+ADRfTAP4AQJ724hjXAY31Vs7JSFy05c3cJ7Pv5M6Nwygf2EkHhqnVWlkH4uNRnwH32jIAHOK1V
J4E1zABwAKZFTk7nCAQGHMYg9sXKSlhY3EyHuW1RZKxpXjLJwUVp22k4FqyGqxSarbAGccqQRhTP
rrAMc0c0KZs5Ewrqo1Xe85O6QKnuduxxexSWAUB3Fy5T9eVRdrkOhaKxumHoBZ32qJyM4CRPm1BB
2X+AkE8favWeJ+63ntvoAzP7A7h7fbs3AdOmSix8K9e4Y2vdxMwiJtZtopoGbv5NXTpX5EQdm+6E
Z+u7nXNsVyAtsSrLIBAjxBLy/yf6pBxKa9muxotp4F2oV+NnRRDs3Ih72cLXaStOtFzlwsytc3wp
YN1rY6QLksLzOabEeGSQI9FiNkVLn7EwkK4ldT3Hv4etI20lISW55+2IXoSRMKmbFziYoMVBx+g+
3GClljkuTkAtBVBu4Zy14ZcuA6aCx6fBZV9HtRQGzNveanffpDPo69VItXjaUbugpagpHRa8SKgi
3/ogM/dT4tTrOg7MtUBSULdo7kcxaAKJgRWAcNhSYLDxlSqU8ooXt6U0s3JmiYwcq/BVQ9GJMUZF
r1wd+nODSotpcrVHLcrU4w7Q52nAL2lFEF49umIIsyyd8aB1fg16fYd3WfjRRAvEMcUk8lq+F8Tr
/a0osbdMFwiLEpj6o+GG8S9bKL678DElwRBYlRZziADDHtxrF0mk2MxGbJHQbh63aWwJSgoSdvyI
Bi4tJ68CcMqCraIyNCPEIG2icOcNC+1/32+NNygOY6TrSvQMjDw4jofrSDG1SIxutaXXYS5gxmLe
E9lZqEDWYFVWNFezW9sdITzLYHZDOkGGvkW0KX7StBod/dsBGzUFBvEwvb3l711DlnOAYrKuwpkX
w6PvGYjj1FyrlDl2Thjob2v9MZM6xruCaoWg5ZDCPe9EV/g0yRGL/2Cp5G6jjinjqgEW38Ppfk5A
BhxDT5OJyRKY4/fApdSw48x6bIUjK0MgDiOmi5mBy62rW33m+k5a3gaWQdH2uBIqtECRwYoB2Cx0
xIXZdXQl2pcfaPMPN8/LF3wpNQ/ddA+gB00d95b6SSstcKQTLR6aq0dn8jMz7Ni+vSyC34t4XOtp
27PVMBqzgm00sddOKUI1OUc3+uA2SDaMsx4O3s8W8ZuY8+KF437FFPoG85O3cEAMsDWlcF+q4rDq
3XovmsKtaalTUDJO/IhkyeLkGxgPefB1GVU/yh63LhVGCB7h7QqSGJjVhIh2g9wEFEU/b3EVnBTF
uGA3AEfQf7jsbvHhIVNyV1EQK+iUmzVLzfgNlxYjER1jNsZRt1JR4uylkJwpPLOMd7tU3ygyMTM3
LB8J1wvUl8yvl+sysTmnPduBlO2S0zoBFwH+QQAk2kwUOLkJ8FJOCIKsnReK/lthe6bngc6WYFKL
izPvXiFZHMl71yV/Y83ePj8JDbsNQ6DovyRzkLOPbqWmfEDt0DHWyE6Q3/2VbDqHeu4QLaOuGFwA
IEn6PNzeHylZap2X95tAKV47Ih13yjAJTt8UQ6FpcD/BsW06ISNJvskcBrRh0kdS18ezs6Tjy5ui
fIG0//aAgEsWv90P4iZQB49GGPSccbvs8Xhw4j592VT3di2uu46DuCJH8EKnhdtVl8XjxRjynNK/
NY3WyIUxihjlyORa10VCErLCDz3kvl6hdZPOgC04tNCLgVkCadrI3o2fUpA7ofArtyhsDn1g1bFg
Fqu6xdbwSfgKdTJaGOFfupF3nck6so17ObldmzDukhitnz1LPM5/j9qTehRRdrbdYdaE6zKYVyss
Hm2rm2L3HvJqGLLEMDiThHt7vrPFCX4I+5tqz7i4RJvcwMQOOUCJon+YuwOYZaM8R/OFcoZy/RHy
7qzvX6yLCDVih3exbZW1dofK0hNWKnNDvG1vf1ngS/r0cBUxQuMtV7M/aMeZXBZsyF6CnSzxjJFf
6TThUvIQpUs51XhQhhmKPF5hVNjLh1nfHC+5xAZ7CWuWULw1YjEzy87rkXYQ4V57QQzh0WZi5g25
CLMQ7hSQoFuopYquAQLGpb39TlxVmxEc0vFakIyuRTuJGURFqcTlNQvjZftcgPgx1P2udErOzzbU
PTfy73+5ZALB4cGt+WI+x2ZSlPMuoLkYY/AxXCsIZ2o/dB8p7/yL0EY++gpjnftT6wfwciF+1q57
bA4JYBML7B7aE9iTfN59lgGk4iGfA36KOeZlA5e5BNAdB7FozTCq/39XfKhlhEfEPx8ZLzv2J69S
LUQ7EXdKFLZSeVLF9qg9qloImbJJJ53mUndDniLBv8WtnC9eZrNjGvBWhZBVZGYrk6NUHPWFGdel
TMKjh2N0rsfgTAtlRUKTtz7CZ/o0RUBjY5f90ETjuhT5hvxMuHBmmUbzJR00eWqyuw1m6SO77hw7
q07SNP5s9gUIH86YysjzQaxoXdeBgHb05lxtFCgM6I4BvHSYMbRRJCcDwkHWoHXm96QRINrOlYKk
GHYViShae6XgGxe6w6Uk4m0GxrDUMLFN59tIBRWNgv4CUJUW5lyK/TH40C49PgqCknGAX+69nyPo
qn5gq9woRM3pNcvAAw7Z766aYPwC/e1tihOVLBetpLxvA4jCR1DPAWmiQQ+kC8Ra6mwiNH2uwDTQ
Idwf9rXM2WCpnkv2SqcVXBYkwdzYK0ASfcwicRge4L6AxZc5n79npKaN+WvWW/fmPzNe8pkK1BPq
7VW438f0b77kZXbXXsZq8iN++fLC+EHWJZm0bJNfmWMqv47eTBJ8Gsh38SM7WMniictKiRSXcPIe
OmhuKExC41Li8cC88JmRFodbqPpJrknkMxayEwXkaO58lGAFjqOAA0SbtJx4nuvJf6YAoaYKa1Cz
KVCpY0lYjkpHQVbNn/f+mt1JOA1wT6evdr+0YnZ+Bn/8GpKcDeo5a/crEaSBBpunXwfMfQ4ILwq8
4xEP3BDv5v0YbovJ1VEcj8qDw0pqtM4TfnQzdw4d234djtg0kzHGy76TUpG6AFV/GHArrfFbPurQ
IZIx2CY+JSCq6dAVQQ6R89JeRXS4t6jzDUnb5oWjdXYBHfDa3apx9yjZZp12ZCowD3snj/yqfNad
PMJDflTRbmk6rg4cl8kvT6VMpwqDGoMgn+nYats534DW/wHAh5XwJUInpz1svL+z2HqJo1yGxtBo
KTFoJN4zyrSuc36h6ZVGLMHhr9mQD9ypWhXWWPS1Gp0NfPGiurnYudibAQrhmJis2DqzrFmxaj5b
FxPoa/uo8ocH1BzxD0PSEBb9O2gQ66kF6DYq5PICXwlE6mKzsPbKlkgtluoTtaNfcU1w/bH2zQPC
k1EF4657RBYyvst4dzdVwqOxZXVHhd0/b0Kirf6EiVZxzH3BcJsu7XsWKywvfB18/j4MDSseP4ir
pAIFZDz7ZdLJ3eZaQNllS84MmcZEBAU1WtSv/EKx+ACvtZMTNfwSVG17unX+Je2aVvS1ycm3XPx4
QA+8S2DLgqPgVBLXMkoOermc89j6+8KJCUNljqd10VEefKZb9B0MU55SPpUaNwWlcswXUIhsygyW
k12V3VbJw1ck/cUawaaBQ8E4sVdOdaq9fqlMmwtNBtx0srCdbE+JIAq99pMKjF6bG1LIjJNgwf9N
T4zKqujWDhq658EOruShSD2/kcTpBjUn029Sj/Gkd9AtHGG0RxukBwouguPQ3m9RSq+rKXWNebFM
iMjMEiX8qStokBznAUyYyPj2QQ4cQQ0EgXXvYPzXZbotBj4Uz9Y42aDK2PhDjKGW2XiqIE5nY04N
yF79UjKWHHXmC5PTOw/MyOrYhE9lauotSXf2F4aDW8EyQjuXr17+h/TF6wF2vCWSeQBc6ZIvp6KX
/vb/TbL688tNS0T7wVUr5xIXaPWO6nIWJH7/vRbMehRjSMXQ7TC+Xm6QZvy78pabjO9Vni7wd3ap
2t0WPMLEWtai5ApJ+dBVDK7V5CMkYKSktgCiMpw42h9+5X44DvQU5cadCq+7U2lONj9MqWIv1VPk
B8xAkpjGYoKzPbQR7dSTr+M15eNAAHcBWkHCq6DZxUftfUgWOGzYBaqbY4jau2Uj7+lm0yTAPLay
xa/DNcuueKJc9wpjKRQAC7+WxGozO+F4DyMH0hr23a0f5s8rYbwUPBqaI7+BUBW73UQIFaSMTKRu
r/kFYmDLgiNDSIwh5q8IiBwVzaDJhYj6c5kTmgbHmb3193Ti+k6frGXpsXJmzDv6SVfqLLIKxOQv
aVuI40vts9VCVnmMfQ8XuaK3TXbl7KOm0lLShnryaJnBGriP3NgKIdsLYn90nGB3dEXyCYX+U9lp
ntjgZocjKpPF8ehRAncfr9q8njbWveY62J61A50/tn5VSm/VPf4914DAT7GN3AuIAY3ArTdMGKbe
GrpGVUNBhJik6+G70D17Bq3h80DM+QRXRTE12paLBvo0/FZEKxYPeopUw/3fMZ8Y47xH0AkfsJIp
G8UQZb9yVaf98h1pCMpSdXCNTvZwkKRlPQrBTGqZwsujYqWygdpa42AUvBh3iaBsicnW4AncPJZd
tGW1Pc0X9tTIeRy7HhIDE/0DvfCwxWrQK4oLPVMOCfDRAn636FUwFEVKDVeIxO5frSPpWj6o4ioq
CyvZwaTbo58Tu7a2TgSRsW2AnjO9DXfLS3qlE+Hy9YKj/s0+G6duo3sX8OYjKu3u49ZsQGmHt/Wi
jRBXjWSi7ZAsJnEPw2GU6oEe3d2DbBav8f4uqTLl9eBX4IMlrX7moqPrvcXrOl0zPti4sT6kTfUG
+7/qQsCvAaIKYxKtFJoVMZcbvjFQ0vaxKfFqo9mc5IeDy8ZrtJo3GPnKUQVr5pCeF7VbqyfbiI4j
WbQdar6WzlEXTCds8JCsQyGpeJj6BdDNNLqFX2OW2JqPzjmJEgj7G9UiZScAd/hwJj+tZaMbuA2Z
xYw2mcxEK46fgfth0hhbVJRDHacYB4mG2hLazI2OPOyAID8x9uV9KYzFJBp+K0dKtZGHZZDlzpiz
GC+DSa8duYckPyFbDoJh58F+Ave3UCOgEHpRLtnLMRphR6m/cQaPiocjzbe19cLMe17V7kVSvP30
f9yuql1Bo+FOMo4HBF5oZJp7MwXpS37jet5nUirqDIAaKs9DPmevvlyrySE8dIXDlSwsDmcT1ka8
dzKcYtW+3HQdGGGqAZEn9uR+1LQjYu6Rfuv+xW5txE3KfGrGq1g/VDKres7ubXl5UW99ksrUD+VG
ha0MR77oWZUtB0wxfo0MPF4g6/Zo0KLtp5r8LMGHLQACjjCzln/JrOGJFAbMsMuHeIME2OUZgyiN
1QysWQg9eDXzb5MPVQ3HHevXcnUduLdRPxAQTHjqAq70KVEJBmtEKGDiq5WfYunTuPLeSg96JkOI
SG2sxvbrrbA2G710oSatyjJeMBXnDyoSWPMz/Xd8X1Z6qjGWbfGlSGVDz3G3/hg7KW3o+XQ8/6Ur
WTOjryYUy5i+7GJjuEI423Ym7Tg599akV0wWXYELxEphCL+FIxoBDTGBzS7Ryu/hJWxk0WJnvXvB
//dA1g0CBlZ5/Tb+3bPlwidPSm/isk09TOq5DOgZqHRIEKu/DBUQM9fbghQibWeENeRXP6rRsfAf
FqZdzq2j9X8A8HxeYIoG1E5m9M739bPeI+6MYbOEKzSO6Ou6CfgzZpUFuMJYpweap+xMhpVfpN4t
uki3mDTfxknY0xyd8B41LfZUdevE6c1ehtFHFfkq/vtLyjH1dpvUe4oAfXELQIrQvJiS3xNyayBB
o8WuiWKbGzHcliSBuGABafTzlpbf8FWp4S9VNmHasgtRaCGxV99cQSrt7ut2Q30BHwc4+9466uPd
gvsEjLTcXgtazSx1r3Xa+FJl4D9E9YsaEDnOBGWnbnudAageYsJhm8mVsC/8j+7MBZjaMS+kK0ZZ
7nsqvDuioA2c1ac9sD1+unq3yRaIjJVC+NCXX/Eg2XayQKmyp9LSfLhrQ6Ow2H9YPc5HCurRuQvl
GSIUxqk4mm9SqSUc7IMXrfh71rRnSVZBjK2Gk17YArjkd3BQ5xhtKHoiE/ydPwK0umt0R0kRplxu
vpLXp6ZSQX6y/3T2HL48ysiFwEXpRF6C6W87EzmfbQHhmCAtakT0oxV9cyiy4MWSCpObbBvaUnrH
sYAxYIr3O/Rpc1GZBXMgfjAV7LogjTytQNsUEnTZNpgSD3gGnqoZz8Ex/pEArpEGnnwQxswj3rtO
seYGCmYePzj5RazgZx5uJXh8ki7JRKnj+IMJpyRKgYHXvwDOWebyM4CMS+sbpMASLBvGTuE9Vdfc
blKw7eA8B++v0ztqqaKFbZq+oF6+kQNUjO5T1+0VDjmGe+2RT3GK7We9XccmqBfRirsRwIKQXL91
eL70BsrorT8299ocq2VCXqDZWPpYLs7v076Qi63EbhKA3dxULRut1sLmjPgyGjIUuvVa6HPWr89i
HpFK1SgwxJu6PP0AdKkBDAfr449LiRIWZo0KyclB9hG0jbn9bWOJc0/fvGvjEdkqZ4wtseW0YthM
uxdULcaGwx2+Q5sG2DcI+brzCfXfKGCcI0RF5DWsV2M+mI8j3x458CoUXJARByfd1n49knoyEP51
jY18q3lQH0s25gFkwRVSCs0uOpyXK225DsG/IBATXnvhzi3Iyt5yVsZn1x/6dVJWQutoftUBbTp9
YCE5TVvqkUqtGdt1ZE5fqDG+LU54feua7hdAaMS6z0bjtC+mLuFwXP0Ba6a1tR0jCwG+bDEiIAdd
B4lpfJmFZGgaNxglp6ZRTwC3VE8nPQCgg/LCZNzn16KoCDP0mNOWuAj5TjnUl/tP6Bg8qaXBrV8Q
/cp5xH9MbdzHT5DNs0g1dsdr+sYEIVe2XwVaNrSAQQYDdXEB//90pM8jfWKn9kOg7FBhwZ6H1n8x
NsZ8G5Gegkwea1egAh2IOO6Z36fIPLL5C7N63KRiPEggqqFcDmH47T2K6d2cgMHPn5NCkN+p/ZIM
FMI0g1hm22IGhvnReSzCsKnvaA6ijLWDgFy55kltAo9/m9CR9EAfsgjU5M0NxFY/5ewRt638fp5Y
TsWyDy+cBJX9sVTBi71tF+1kWvhLpUNsEgLv4IDXQTcN8BrzfNeMCQUa8pq9HY1zhVJVmYBFrno8
F5YBOHWbgO+8WRWbczXuTBbMvKz79Jwn0UH/jFjtFpLqHMbhwFiz2ewNriu+vzQB4xhoZMx+BrDI
Maca/XH8/tuatId5VZDlSpPbVuNAWwXDYMplFUgHoPFQw3isTsfaN7LyhI58HLvKDD8DfMgM0JVv
knpOojiEq01qxffRKYHoHcTBB1rdVgYUzymIhQWqRSt0WVzuZrrVUIVraP8moZuPRm44Z7ror+Kb
zhFNdC3fKJ7PRj9lsfdzLOgCSqyHeAXOQieZDOlXp1rOMX3+qHwEbxEwspn8Pjp7M6iUOvzxLyVB
V7q6Vcp91RcAzWz5BvSAEU2aiwiXFLv3sXhkcsb1MO5V1DGDGe2roLNu3hbWUGl4TT6EoaIBcMvv
8RpQTZgxVDnD/ZyWywnB+PfNkiNYH5xXXei38smXiQGUBIUr5jlmhY74twZG5CQEAH4+4slAZLBw
3VS7F47m1tmumppNqerwCfZYEMqh6t8rkgnUVxt2x8JBW1VgUHrm4ZOf1WUTQKzwdPrm61YFByVn
l05UrECy++njZHCxymBpgui1gy9OMkliq9NyBjMvd3aUjsLPYFNMhukQaFtQy4hKAyJlH9rns5vC
rPHr6uj+OCmW9Fl9j4XFK1v6gwhQdyatS/baXUs/SFZ+N2ApVZURZQaVQjyLe/Pm6phV3H37Kmdf
rUrwyK1BRPx7j+6b3SmUrM/J2ui8t8sQORdtYATSJ+1nLX+EdYnd2c5lm6CTpGYOj3Pt0AHmaLDH
zpBV49kSzvB55BFXA2+uAgMF8foFBfjWjw7vGNAPR04DHgCSwyN/U5TpZ0/wEk7RNSuz+Tc/MR72
m6w8hTHgzzgJY3bWhh79Lraom70fxsVICr8YgJyTl6C8OEJPB1q5qTdFtBiisBQx2J8oooLDoWUl
RYURl7q0IrqAqo/sSm/cVZqDtLc/1EqI++Jgb1F1ztz8Uz6qw85VqYkZ+z8uS+LN6AyNGoGhcfW9
Sda0bDIQkRRrf9WQba9UtdsJ4FVSNUweXWZ4x9S6otZiqhc5sEC6M+vpbiU5I7upDebMQvhs3JJF
+wxjY0kCsZUTMPRc7fi1OB1FEDLXGbjPdXQ9cToogQ65utfjfWhm0Ce28+tf+B/gIS/rNa8+jna5
Rx25vJzlBlPZnXro47Rq9HH/anOqz+DkrH0hroX2SqTWzMd3sTz2TVI0Vp03JDvgX/nzcg9DrUIj
EPDBe2TS2/OH0/unfhq4oKQFVUnNkstUqqdUzMc+rOFBOKs4M1JAP0sp2q3pT4Dyd7geZ3zjBLTd
jJiCw4cDSK8lV6bkoTWeJNpxAp5UG6+OpmZD9wphz7q4/FhftWBacnrRu/rGjQV6ZnShT3s6ohJ1
zfVUC8V5rT0CUdSd6rkKLqtBF9QufPIMGL8NcD7VUIU7hdMal67FyYtXyyTe4T4iocWVpovpmhwU
dyt7T9daS8IH3owJaKk8mqrkWhxTbgwT0MA4doOAUFpRxxYpxzScFGoxRSeLX2+Pa8p4HVvycOXw
+QCDFMbuCV1eyYFJzRo+95q4i595NrCBJW3QfMKGCgBznO+IWWOFx2aUmcGwKQdBqxPFkMe153nJ
QwCA4fDMeOQxHcgsFMLg3eld2Mp4ATCHjGg81JMVIDOzA65bbh7M/OjpWmBG0ie1qyr0TEapmy1n
TEAuAh8p3Og8vTaziqB+TkLfKA3njQbmK1AWOmiUpf6CJ/kKUQQ65vT5TfcQqdISnFTL0tmoh+3l
eO7vI5U4GgeQh9iScbNoHgVKbOvBxPlfppZbEajoMCTlW03+r+OSLYUhqgVbxUgzGzkYcDoRyV4t
kkW+AaMKL06tOWIrPrNFemhnq0enhwpYS95hZRakhKxb3+jaFc7nd0F91Mcnyi8BzP8ru5xQYsZH
c8QFmCcBV+bSZUV7oyJ9xJmJmHBtkdxBVRYeMkhrPyTKOYlPCLhVIWraGOgXdzQC5uhOmJuOX7xJ
DCktYBmggWxRfi310xnsI1jePE8/yuMdLwCTr/CfHmade9/b/csU6cve+0f93ktl0v5MCFlLOlMA
jpuTrzE+11KiDMYSgcSS++4o0bFfp3G4h3vT+b6EqS4SASwe++xbHnqxGA0BXA6uAIH64S/6XxXi
MFh2Mllto8363ILD4OWiE2B3wUuEoyqVeSn9Xs2eVV6z/TIsa+AbpqVfh4HQtfXc214d2Qnw5l8o
QM7CzjBXx3r+nJ6WK2rroKKHnGwC0YCLszMFcNtleEyigkEybV60UohzFBhdgolT2nVkliGDHt8x
k+4JNiq9gpHo4eCg9Am7yZDTi45VJBGAyRIGaYBVWXEZa8tEYfxL1/6axRP1thZSnjodNGPr0JmV
NYAPGuU9nWq9vhN3zqvp/xuWG8XZm+QG+pBJkbIt30kr9kGEz9mcOnf0AhkRIR2kXUTyNMxRMJb7
Tr6K9tw2KeT2DRNfqqE/eaIlbD58E+/CVv9ot+zYX6o76+PF3au4Nei2bHIWIFDGqL85+o+O51rt
3+yOIoq5yhJBkFdKZVDZ/7dSn3JD6ZvKClZx56AY1c40MkIRb4PR8DvHpAtWfm/bd1MjGbShIlYS
1Gh6HZVghNqHkIANG2fOdFM3JlXyQyQsby+iWvUbrq5jZbPm3K/Sbe7cXQDqwONy8fAdWOccgqv4
8A3VUQL/UU50csJb7Ekjq1Uqj0ueS45tHiaRyQHuteZNK+nC2DzZvKl5ObdEVZAPFUfJOQLou8tn
8QAKeaIQJKzaFBcg9ROwdIhBkyBeb7RyEyFYWOt7ZNi9bOUsuOusloSrmpM4GGBnzFDci32UD8Ci
bC5VixaA9UCG92r+yrMDObLR/9j4mBIZezPx08sgmbRI+iTYAiFAQDQuR3orItgEIuPN8a4p8OGI
Jd6Yau9xuNCAyLwR84R+APJfm/xmlaisaDB7CFWGUHNpfdgT0PjTHQmeTzDO+5x0JMKBOJTcn/gW
HnSkq+4Uk1FbjNzlr/7ZdngNMYkCFaTKpqInPpQjS8NW4s18THx0cVArTGac+WHCxGZgdLcl4B5g
GpGZqxVAN05K5VyPVIu9JxiLULw3azYbBLxBntz1Hjb9kXOK7ZN8w1Pn1SteB3XOFVccChP/vUST
II0XXiJCnk22Q5AAMTjIY8B+u6A3dUFD+dtHNYHp4RQu9dkJ1Iv26Rgg5sQETqTqCgyOp6v7sUyz
KhP9fdQ67vw+rV4ku8c771CO9mzWg3si5s7Oqfb0XV1CVufmpEigv6U9HeXJF6+ACM1owKgk++Vn
js6Bqh3zj7QKvuvYOWypAG2IlSkNWirz6m1TEWe2fQP18O1FtYdUR7UiepmsMZ0qBK7W+1j9zcYj
YgZR+39Rgs2UxHCHckzHI9AeTgLoWDcKIrXU1+mLZvnt3BcH3cUOgg+NHKZzJxdWRkAxb5LoSViW
o+bl2H3af4fkF4rcvKoCrSyzU0hPwAKfuAQG+nJRI91w2V1LKncCskhLNwmbx8Cq7FgxpOD7Rc8G
pXtzY7LgdLJTS+IEy5hP9RJOj13xdVPN4xQi/9c99+BTayl4aN5TBGCtOflojCIUf0U7TNkAXhvQ
uaionM7EEkKQcpmVq+HptB01Pkz9orV1mc7B8KqXsxy6rtmcdXF+T+V+oQVZVv1iYMkvkPbFKTK/
cjLRgWLI6cINKWa+D9Ja57zQ4Ut6/KwfqCWQBOYUOjfy+96WmDyzKxhmuxCDlwxIyQxm9bivDIJ5
I+4UX5TatS4wa/Nf+NcoJR7TzT+IiuyJyTb6RP0bW67gusQlgNfTvuv+5JejmV1cbawnYAxBNmVi
I2++Pd2ZnZnH529I8p0Pk0MLE8fmHGc6jtcYa+8WMHPwg4qmEvEvxUxQotlfXZYnEuhyOxCZ/DZB
5G3xY605Ix+IZhbujO6rci+zEkW2ZDHVBDsVLxEHZwkZki7XcADkwpkUu9+vhli+svkknNZam86X
dTwhDkCBA8KyTY8R4UfOeX3BMar6IZaHM1oU1vNp6U7RrGM1F6MGNCKqM3mqZPY8VVv0J6twd7yC
B52nAwrlL6ogt/+kGjw6xYCZqLHti1BH2bzWMbetMrYmgiobHC3lJpuAjg6pCwhi+XtRxVdEFWaE
iz9HS3DHjhbbvGt1GrnZ2mwdL4cEe3Rxd+X54m4BzUc0JEXkwgmXICIi/aVo9bWPGZy95lxt9nyA
ZgRaJnU/tRhirnyFoTodNKLzxgsIUs9ozhCNlMWNPswO8ZGRhYI4vgwMr3p6ea4UqcZu3KwkqaMz
KjIKPQLd7b3um1u+L9DRFodKOvJcaoIqMz/+gnNgXLJosd+uMAK8WUlhAN1hjLjlIfLpc40Fuogj
Sq2Yk9VEto9IFfy81lg3G4XyqFPAPOLxkg3yr2Ku0YHtRBnGgYtSCBYq+GjMzddv59o5tna4xNS9
1WCEhug/5Cvgv/pE00yvX4jAJ8qrN8RTLsO9P4SmY2XGx3fYItinjwxYhsVjjo942smGsqOuZcCD
U1YII0m40uha7Obwf1eiCzXHupoJhAPnaJGmtBejrFGH/5b2b241QQN12oMafQwdLD+90maxuM7E
8F45/WiKxXfNud/tvAv/WU/Sns4Q1mMxqxQn/M072pJTGAKbF4eQT5Qr5V1/QTzeJbkMMGIjuMHS
jYCdwHloNbtrOJ7xCBnCzU5NrMimZNAMXVhgPnnrVS+rckqlZBTAOT2LlmF+kBSyEZtIMbulAJYx
H7HXkZDsj5hAF9D+FLACvmXMI9tej0XPwWfVR3EEfMuqA1F6KQKeks3QlvmDoDBaYzbnmVMGcoUt
YZNAQSO2F72CTN+Y60ZSdQPUsHjZl4aytOWYpLJFWxTUy7DpTjqVALCMiiUqEpJGjSms9KGAX/ym
SG/5Dnye0uiH+BdG8/JCffzgu5hBbvdS0kt/JsATzU7h8Izpa1LtXD2AiGalf8lARxzTgIgCuUU7
viO6JvrbkVBFP2pdp+LcEvzcWoz2ghx/y+TphCgrjw+4SyMZ0+wSruhfHw92necMZ4fgTN6szhUe
8QRHNzDFxhDB5NhZTjwzVn2R/Nwq0EX9CNs1G89DR3Ldj2vU1giM0SgthrplqRLEmDS6tIN3qNHz
7U0tFRD+qeBSu/vExJKmGdcqsPDkJbXyFH+yH3XqNmcnvz7y5bJpg6QKACpg4b8iC/Gw4/GAI7hR
rZQZOGLDFY8M1Uz/z/3wbWQa6DY0WsSIJnTG/VEFiyxfoIcH0HIT03Mxzd+bnUNTUymc85WSsxLM
N6S9+0jlRnXlrlusa8TBa9iCQhjwsfyifFeXZrOJpzcz12yScmBYtSlnox/0PApCCEZEP7pkHova
KBfBQzLsXMXTBDCzuryqko0JcAU9X5rhhhHb50zcc+8b2Rb/C8WoE3sksYU63xvlVa1SAM492mQk
8E5QxalAqOGlmN1GKh98Nxyfv+/ytdtHGxstuc/b9a0q18lZHv3ZArnv8+xjH7u5Zuwa4lz8CAmR
reUJFlLw6CgxQrtXnFK9Dg5LQN2dJCLDWtDDgi/ktBWcxjcx99g7YLsn9nKR4trWfMXHzpPO2cXI
5k6c9XkLLwIbbncTJSfueiJqykNEKnC5vyYpT1j0DfRavrJZHxOA/dBEeIUa4aHR3N8FMCAZ/F/Y
g4aMhAhyylghukEk+c6aNjXwdFhPKJl8qZkaFVzfrM0CKrXObRnMXRR9Smx7ujJkXjtKrTZ4FSX4
cwCPTSzcPLtxqj7vIKwdvcqSbdIkSwihR0GdMaGS66o449HwPpIQ+eaB2z40A0TtQK64vcNqeua/
7y4RFtczwM7pEAi3RvhZgs06KeZ294/lgmJSndiIvwsInjdv0WTbyBWIO0KzJGaS7gsvkuhUHRIu
GEUpUKiYTXY0qZFERkAbAg+56CjdBGQEV7viFxsp8PAhADvDQbIEcwEfynEWrCqa8rTm/8bscXMb
3M7lqSZc6mrfFQ0Vw4koGGSomBAD2ezCa0ixF2mr55IKOJxxpLAa3nKVzvFb5MtgzatgBinhKmx4
23BmoNqNmpAkJXJTO9SYPrvbt3oz77+gX8xIoh4T5KU1/lpPRNAk8+dy+p5ZNPW6K8cS9D42s9Mw
JlKCNzqQybPNe9E24bLKjlPa00zT87HBnvXoPL+YD1sVzIlGaJXzQmD5RzuZRS32D1GxQ2XiB22E
o2AoDH7wHP30DOfXmeIlQTWqz0aLq4CThp8o2ZTKcjLq6SQeSs3kyj4hI5JHUt1X+hU7VtMQHkoh
n/pdTltr2N9UIfQq1gocTJW0rcDZeopidf9vwzEJZQERjAFsLrHMcmh5mr4GlUJb9oIYuH9EAGo6
MsBmNF++ga8yexU94aJey3SMEKBc8c7Etw/wSSEHO9LKP6/1WAo0WUZkMfMKJV4C6tFm8HMPSgPp
fELwD8BuBIc7ZenW9WyOdTeviBax/CEUi4iltqeSqn+eUQ/OD48fqtEWRUVFdZiaYovaJY2aYbDN
iJs/zaz9uhxEZ+9XhUXWUroazcnh5frlDurfT2Z/4tMXgX/pasp0xhL7sBc1oPQnSlxoE05bpuCD
6meN4JeFMDr71jqzLpuMDBBpNQq2U3jpiQl5AyLYI0YZkcJzRjWj2NMbmL/F/Z9AR9WSBmp1d1jr
fvd0jDaS/etcCKM5Ivcml3t8/D/6gdFs9KVELrJLgBeBBjc8EoXMHYuloFVGgesUxnRPbGU8WrLd
kmmWENcsakCwqxIOhMDfe0praqc3CmFf+QIbOk2fToQdT3HDP/6nz8ODL/KdshQ05ff7+NeU05Ke
73EQxeJehbhTtTIXE2jzsQSSkd9pFRDkHQ06RXrk/CLVk19qUkuS2bN3eagqIxSXgyAsmsUuICdB
P9LV1Z3bvm+OVhDyxS6Ln8wfrJha54C9UGUxg+cjmXHxUj45yirIQwZ7i8/t9nbMTWrLxVwJc8m5
ZMpv60SuQ8/qdj91sf3EEgT+nc3Zi6JGqBPWYgPosbf7snLGo4c9meITbDCt1y+mxIwJwvB437bt
3fpgJLbJRbuHHA76bsp3aq6EFlfPY7jp+ruiOLE+YVLA6ezBxw1MpX3MJCbU7UpZhEsg+qnSEz9e
IbX2Wy5wHJkp91rZYczKSW6OVwObv4DwGWEqqNKLT/BgXyrtlOwoVNhy9FELvyAo5Gi0ISQ2FI9N
2IYki8MtaI4LOfcPw72ik/onBzSH4VS5gqNHm/aOWJfZEWGn7puNhnqw/9/Ri9tem3hd76jtc/IR
KNEvf/Dk+i8hMHUhZoHIuH30Tr8XeswAXhUe/vJwcRryYnu71HNJmaQz5romAKZw/MJCJZiurYvb
ZEP3/L540FBbdovc2BLHtsbsq2ebdZONNLeqSocnZPtOc/PpGB9yQO/A0feWWAWMwncAwh/0AqeP
clNyvdhTJdLBL6ayxzazXcp4OjoxKUF3cGxDQZiFUDLA/dnWpyB4bwEbt0dLHIfRMuIRSi9CLdO5
W5L0esTsUqNC/X7RsAC6zEk8jtEME3V5EdtHVYGJTocLScZKENIW8gWuLCshQSgiJatVuqj+pGYo
KdFQL/L3zqUyc7i6dg0y6BlSJhrknUBUGSg9N219nY6H2JHWJ/dXz2h67o97eEG7/uFBn2q8ZJgJ
dRzVTVwuSZJfX11WVPv22Gt3JOwjHeUSNrHA80rUrJ+COzV1r50TF/Ccfzzn33BnD2P2t8DEcS0R
m5WQCrinVNOU23ECLhSXBn1UDYj9zQDEY743FxEiYjB5j7XZPZsOddzMe1tCap6FDpprT67tV56P
LZ2VRmkdRP6qWXo4pgVEWRY7xOWHAYynUJHX2O2J8sGEZ/o4M9L3dm33X4mjNJE3VT+lbdQibxS1
XXsR46phMt4p+MdDM6lHQKQg1ksZp52l/NSorjP4u5lEMauP+kkNtYDkrRx735AOpqheSZBydqDI
F3VNtmJE8Y+jquX88s9uKLAR44W5Cq0h8dv/0Pcrab8liqIoc9+WSwlYrmXKu2DMNCGDJC/PEzW/
8GDFxy+6rwU7uQKStlWTwT72fsGPy1klYra22HflAIZeOOnA8SonP5Rib1M+vBy4BXf+txSsAghV
Pbr4Va58ms4gi1KIjBJckD1B9jzeSl8uqURk140BMt1mP3tfnrkVcWEKqiMfNFcNLZYPT1LqpHgX
7r2R6IjzWHL1PGVgM+MuWH2H1nQPRoIPAe30bN6gYCHqMoq9gT2ZoGkF11iOvF4ICQ6czzGH3tkn
nyf8NaG0CqSlVOxnBfpaSxPmCf+iw3axr//OfqjZy8H2PijeqreEDH6m8H4f0hChUhfDbqH7/MQ0
9GgHT761Dj/wRhAiQET8hwVIRpmnIMCqXNPqTCnc3C7Wx2KgdJrEaTDQmBIygUCQmEWAN4LsV+eV
AJDxjf22CNdhnejoPmj2/HppBJD1pqq0CG1135Iu602uXVsUnT3RaacRoYaJ65q6mupfjcWUaYOC
YPTu0GOJt2WW8q3+nh42IbIO+UgnfSI8ILYz9sn1Y/KRz1mF9f/4stSPLepWwDd+ABtHrpNBjs7m
5oPKKZmQk/exk6JyF7NY/7j6wCjBnPZZufii/+HcyxrpzOPDs3BM2JnIRQM9iY6Vp1Vmghl0C5EJ
PpW2+H2Uoq+YrdMBngmeRFPRBmABQtT097YQuRUmaJvVRUTILW/sOtkbMVpi3OLPg//KUFieA9Gg
UIUHGvWztiJTvfjBPk8S5rmem3wrsxbIet1osrUqj4UYprLCPj9MMrjhto9gpD5hIxfHLQMEB5oi
CVrJQIF0LNi/thChWJGAPntmT2oyphS8glYOAWtWTFGhK1QDsyimCR+dTiF00Uk4YkVCqSuJCi++
JvlQUOG+H7SKLV5/cKm0fQ4xKqMwOraDKX5zIktJpGoQQYNOA9ZYRCcxlmXnLp9JoqT3sQiaPbIu
GE6pdzDUCEGiiLjwgpgGg6M8kB0PGdGu/v1C+LPoIltJveQlP1JSQSGpARWm+mrKTrfSTNhoVKlY
9dzfJYwqUtVIKWP0Ra8CcRBjmVyXgwcNJe/ukfqxTHDKR+BcwHLr4WRn74DUfYnK6qAoz5JlORLa
e/5UlVEzSMDufPXQ2ZeLZpb+e7Onh/UO0PvWzVPWLefzD0+Xsr72N0CFxHMPqkMzRn0+ckXCZeID
l7MrRorQRPTv5fwnwkj8MsaZTV+AG31l5p/T8qU7InZQoffmWMpGkarXyi5iQyrh8BCgPYE0Cv7W
dHfqByI2X22fsEAMf3dRWo4SpELYXJyvUFvmDaRpo2QZcYUEneCgIv91PfIvUVc2s6puQDEyzNTK
cUKLbZkpSe4HoWXnN/yflyPKWJwDmUXzLGJrw0fhpzsNUr0zk7i9NXHui7SOzQ00+PdAfKK+SZIL
Fai97/t6nd+d1ZIe1esllnGDhFsPCF/XGWvVoZbMXkoKCokFJ1H3v7dfknXFC0DyIVtQybtd5TIo
sVoxuypfzmBTD1O57IMq9HHT1d4UypcfrknE4DG3F6mfhAjij2eqyOs+h57/ZyA3SwKQ5iaXLm4G
6CAg03zd+y2HhfFlcsg55QVUPWCWVN5w2xXGGTEPA2r2y6S6gYhu911awXCo+q/5/FWam9havuEb
4Gka/Dtl8FkUCpyHezbgUMeNQM95r/JT1EMMEUtSPrpjbugMNI0WMcMzK1o5ujrU6se5xci2Oz+H
8V30ab7V3lJUowSTjpeMq0gPA0x8mNgvC78s2bJvKRHlC2GGQcDrlFFNNIjvZxWmEqGuvOlfKNPS
NXQ0+V91VKS1eiW7hKs5Y6WzQkI17XQlYPrAq69LL88ij4rmy2rUtjl8Q44NmSi78P6PT35a1ON8
q7Bq7XROdLlQhH0Y8s3oIlzkEuGXmYqNmlKJXNvM4P+O6q6P4895lTCqoFS8maGgUAlIWjv3rz8H
H3kdqkQhhIiQ/KDjPpvhLwjchb9GmQWis1XK7/Mm9jQ+vmsAM+NRLBUtmBFTuSPgHFpP+BBrTXkh
RJWM4Pz+yvonkbg7ljJKKcAzJsfMmZQmErtUoNUfcn9tk8IxNhRZoqqRikn3uldZpXguCGZvsXVu
EIwRYstVsx7bqEQUP0EasTNjjlQSfVVuLYm3EwQUA8UtSNHuuadxB4GZlzSMw38+d2rzyxEXnIS3
lKcClpYgnae9nKpuSHDPypUm6bdNFVdnHf+0Bu3cVYatJ+cWLHyS+nUs2jz3g8Qy+und/2vzZF1u
c4eUrPtC1Kx7lthLDHHhCoYWtwQvrkj+yZ+xSsDlnL2jC7lULOsU8CFtjjajtHlQPALGwCzEdYoy
yEwGjUR9mcSxzPGwYAWTtc1XldBwn9YG27Ld+7bN4CPCyQ4oQ2Te9WDouVUj5uegfQ4FSCjQ9t7R
DcxPJ5cGdW4O1u9mCFy3isK7dWQueAwTSbzKl7DNNdzH+hc2L9wZRj9281BotHLsqe4QY92DgBnK
ZS91Zcqsiu60xzO8Bl6pNIH+6Jz3+Hm2mUKvpw6wiqIICiVrvxk2xCadYLoGHfBqoBrOCBXBVlHx
5gyxVfS1SljlE2o4u521V1KdoK9lTD1qqVIvdep1DykaB1dfBlspc8qUv3CdVEMq86wrqpC+Ml49
ns9bkWVfJAcp3D9nM0M0td9nVF1mwkEcZwpb2wHGnUjOzxASj8MMckjcW00zLwUi+pnv0qh/TNey
2VvA+fcF8HYByMOd8b9kChfCrpQeWvpqyQy7YZXqJ8VQf7FanMmI81aYrjcgKQoOuvYMlHQ0gm0D
5l5QPoqKAbgVDQv+TXole0Ym+a8pFNrOmaw8PY7r+egDldlF+C58doyd2d018KjrWymV7Wo9nPTj
+Qd0erlX214EI/RX1H01dpyfFv0bFxtyy9d/ytF3XBOvMOjFalgxh0kXSbyEvjnz5evarywSA+BX
rP0CokKbiha0AQY6m6EPShrnw71ZOKo9IDtw2M0D0YRmYfPJzuMMsUEAK9btOpW+lZUejDRskH69
Iz7xjsnUhE7Ltm7EtuvN/EiNThgYARWrmrvIWOG7zHa/Sw+mCOmoPbdvXsPHT1JAU++DFS128RZh
gMUb7xA7Gsa8lIF1iB8K5NAvBEux1YKxeBZV19URUEyTutlJtUN3qHgAlslrW5Tw5phekK4BPW53
YGWFey+u0AHIV1hxD0VzpPDEJghtQnimX9cPxMbL5JBYwilYE54/o75yJu538XluepN4YGcRVQul
omiOPetrEHEYqOdA62D04ZY6e54FSnmNBzVGrKdinn9CtYfPnOI6dFkQ4HapWiCKSWVF0gCda17q
8Mw4ifVFCP+qQXeCyPg8N+CINayxE0UcmtBDeA47GaVnZqCzPldDdNIMTCHMY4ggyxsJLnLF9clf
VY5f0QC99F8/1e+PwPeIz1BPIvJVYmT9fMBiYMcZ8pv19XQ9vqdSPDpAAJk0tw3poJhxTMGBISdb
/XODtD461rOg8m5Uks86q2unCOx4LCDmhppi90ffYk8OK4F797SIhOa0iNm+FK8+4jvuZR2h3L0v
chXp8WtcgChnJFCVJHsyoC7lHbVzlwI0ahS76cl2OMNTnViMBWg5JIvLgJOaoR/HevYrnBEnEVQN
c+SrdsJFushenqWjDEQn1B4JyruDggzpBP6zWX+msNVEmxQq5SnMmhT+wDb/9oTXfA6cIve2bH4i
WNgFqCHVPUAyV+7N5BzyOQRcEW8NkegXg2JYacRLE2qy0/s+KQ8voJ8/3+5b3/kyB0m02e5zX4ta
ZF0sMlX6gOk0kZapxo6sPJ9uCYIltYNwrf8AUzuhGFxg4LiGtilEkajuSlSvhrOkIGg2jxM8tu/F
brSmIJDJRiM7mRXgMbAdui9/I54e0+b8H5hFPS9xOKuvHaYUThtyNmPbwXqpXFQge5rzBAhL4UJO
Gx1ZreGZO5Ryt2uKcdj1nCZ2fdezUY8YTYgCbvhK4LgPpgaYAYappMDDjwiIaG8SeoOp1VLKsUle
OL+9XKsRMKMsDGYyQQK411iO9/a3+2kGqpfLwyWYo4IT8jdefs2nXnHOkHxfOeQpByaiOJZxh6z3
4+HXB2cRjATwmiTUIrfLB2xWVYzHLX5k+3Gj5Lu/1qgeBk2Gp1dSL+sPkZRRys9Gl0u+FPLZTNgQ
gVATMvHLX49AviiGWfVwIF+FJ9L5waiaCoQ+nmYO2ThezBLYATZnCniQerE65c4gH60LZ3xpSmPu
t2zURNgmM9EMk4hkZ8tkrsmpcnjO/NxuKjB9UZuBxVxLIXEKmEeZGbWLwlxflGcdcUelm8+XcATl
6A9Mm0W4tKOqHl5qfqgAP39OemwR2m/p9c15T2ql63o8eKgEwbJeysZ7dJ4+OVg4sQCCq0UK/V+X
AQzh7xnwdV7qL5a6pImyc8pBHj/ve3KvxJvsM/qDK3/HbCGdPJH/ofb67hzD7mFDj3w4Ic/iu8sp
enxPtdiyAkTwwUtDuS9iCKLuJp+j9Hbjnuny3TQlNIF5vTRL0ChmriaYkLTppyxxwzXcsLBm+quI
pqnyRXKrZfyanGad1bOE071vD3CxfVYZOflE6UefLAV2UwGGR0ELQrIzaWAz5295X2QEDX/X2Z5b
r4tKArV1UneR9xk8fuO/u+z+4Ti2uaLb8WrWaivzHeQXiI36Wda6atEi991pEDR5+DmLKRkdHgXR
xYQL6VuEFqYTKrPneZRz9LcFRBh5wAVaty55NxF0F8Kx0yA8Gu1mT/3i0yyMMUTgj48CmChwumMx
/1hJ0u5vtj1KK4acmULhP2Nise0aDi6q7YPH3EPvk46Pmdcl4ER9dIdobS4tknrmNoOpXlk1DBXv
L2+hkP0L+tucT8UgV5PR6VyaiML9HRuFUNQqD6R/u1avQuLukSmnJTuV4OphQoy4oUSp2OinGI7j
62xxCYfttx5UvCNy3kVUh94/RwmmtKGCRI73XmfrU5WvRQ9e0eOcu5AWD7aBmNgcVvkslEkDkIrK
z9heIXLCSuqbBFWYBqA+rJvGmHkQvL9WJMLi3vaYoBHqZ0kP2RAEv+tcofrrYxuMjv8J9lg+awxI
9kSjxVmd4rVQ6jqqSHoou7S5CxqvuhCQJTFh0XPAwnOrntWcw7w8d+8vawkGgX9KMM1S6FS8eEHm
WeC/QVGaskh9tZtThlj5FdjI0cvwvMbojd+sXAx/k6DlICJ84Zyv0N5+8ipMTBGV+mfh2GyZbKrQ
WS8KAObWQcrfiee/I+GktujY+F6gO92El+zPG90LvsbSN8TerUJoSVRMfH8bUt6/pwts2BjQVGMW
5+7qNYvc35FmiFBfdHLtQpC6iZhtM4dOQ8Jx58MLueAQ9YzER/4rcuj9zLKj4GvyeFJfqSk7ZkL8
EXOOw/hj5OmHpEynvxFbiPBQQSWxaLDE+0wAVgNEn3DWLrZFM2qQZBF18c23BJfwcBh0h+YH2JDZ
m9KFPVAseGO5RGTR3euN87ujAlAhiOkoydmaeWWT9W29p59PSL8DhOUgkixp60/OHJdmudCT7gCw
52Y4i0Czh4oFst133sQoCq8Ewt8h4gIlq/aXSUIH/+vhXdmgANu+erN0+dWXhG10dlosp8CTgyIP
qM9/IWHTME8gg/yXappbywSRh/HVpWGAsk5IY+o0RaYBF1grCuRx8xAZ4HQ+ygua9BVLDxREFknz
RfFcOYyo+TQFUxDvkSczGwkE7qktm+RGLfTGTqJ2ppUoniouGtajvEfO+s+k7DQpthA8ac9LqmeV
YpUm2qbW1CN5hSOmgPpgbdEbC3YK2TBbJxxO3n3X8kS+9tx1G27C3rmT84/z5xDvbbJuQhxa9Eoc
k46Kf2dZ+FYnHyFdrvv6N+3njKONx4zP3fDLLHolFr+nU6ae/Qzncgicfw3FbubO34pZDizD4EE+
EboqybYc9+H/NDL5yiV3q1XefCHmjh4o6OB3QotqkraXweunq1YapX6yjxSIuNnsptZgWgetu3y4
Mar4KVdw9FfglWChkx+7dSoJ06mLSOxwO+Z7FulZL4vab++pMM/qVvIbeSC56G1SFfgLBX/7w5Rh
++4flJd64UtBMIVk34coHbRT7u8vuSaECgMl9MIw1E+SV3SlPneXFPxT8Q+FsthbWhq7A4sXqk4b
C2+nYQOoc+eLr+fz15evgXkbr2zafIq2mGnbASEu+j7as67/EPvRq8CoAqCaIWxzuBU3k3LogsyI
qvhRqQGUZTexKt4K5tT4ahNvSindl8nsD2tzk3OpyGeOtEf+PwQwHebg3pKClLQR7HFd6wj/tScF
s2Ia7pq7VYfYNvVVNQhjYTZYf8+RocHScZVd8S/uYTs2mfR4HzVfsBoIbeOsPFCLbIDBMfd57ZqI
VTyFCwxVmyAavE56tredQZTkLeWmUq9OYEKWw/ZjppI9nHPD108ZSAa8gzGkQBvArxUp7iVqJDwr
5LgDi0CIEyCHln/6UETBwEvyXrPyb3loUN5CU0pv8Gsruk1TC4t51MoaPSRQ/Vg332LhXjTbpGeC
vYXCGHbRzAgZ6uv4Y+Zb4Rt89vc2qGoyD0bxZ88JBP1auoha/ZvhZ0XsyAo7THazFg9liicfZ4mM
tCYGrYxjVEHGfUYMKJnmEAvuS7bDGGbAH3SyizP3ALDKZXdYCPWkaBEH1w+qmazqDkP029JkDqOm
53vVlH+UkSb9auZV96jLW/caiVcGwbXl6TcWBjaPNZvHkTdZqNzfmFNSxmv9w2S6S37Mcp3hqpj9
6KuxXjri4OzqBHeT2KPpEtOh8Q5lvT2wM9QvNFp5sF4VEIkEw+Po7CaKi2WjZgXFlNEnHTErnrSP
TTiybUZu5ldHQpXrcDMwUQ9dhrCqG2qEb+v9DMQEg5ctcQOov4pYPPe5czldbOi65O41RQ9NFV+x
B2YhG6taaY0KA1/f3iI+YST7mpuyqMXYU4ZuaLK7w9KMvm2cDSnYdhEtmFHEJyR0J+v1byucu4MF
/zySzqPbkUfZ1n3Z+B2HkbWVM3Zvsja406K2SkUzSPqOX3/Jj6PT/yrLeB8MKv98Wns2RxSMHNfW
8aX5bA68qbPbIKqW2VGYyKPL7rLRHZQBwE2idZW5oD8NfDNATVo6ofzvryv8JFBWYghMEznsFkga
+CLsZWl5PdEnSf7gmKo7C55Ac3KcwHjEa+S4U0hmC095QEqLeZV3x+ffzronFyBVm1sbJbTZaFBv
bj+3KTBMIm0Pc7d6A9TU69auOqAEe6V98SvhhMtXEF2FeMRl/wM9KgshFp28iuQWjIEJRokti5+o
DWRee3A3HLt+N/uzR/kWWfSt0pLaMKgpWLj1fw7X4uqb2nKD/kF0FkBOcDZcZ/3NP4PHYUIQ4X9s
PCK0ILI/k3dV4YD1foWqqPypS3ObHQpyf4Rvqr9fwT1x46k5G7PvVK/A7tSgBeB9+xW8cZrz7kpe
IkqUwbbyeOBItsZaxgP8BdAb43aat0fjsda5n4U5IU6r3TWitM5oua5SlV3gNpUuE1YNHYA56BuH
D+YYLUpxlAuJM0SDauOyabVuJPruNagpYXv1Hskx4Rx5nhf9RysIbaEBopBJ8bZ0YMUBNAD9QWoy
1cZH49h4V2oLN81oMJ7a5snhCHAUzPgYwu0uPoUjlPVqa2v8vKNBmNYOmzj2B+SBRsO1tN611ZLd
ftNjSA4lZhACyPrcvc//dC8oLlIUbUyr55kQY/OTfSXZlBVP9mdhJhnKuH367lecT9uMDhr5UIbQ
qagUhF1tHwTK5E4UzBXf/2ZuAaah6+O3ydyndyujyHWU9ATrzCgELFFbW5Fz50o52s/ua1UasW8c
8Q+e5P29tssSXSVwD+7tW3WdcPAjtxamQoW0FKYL65PE7/5YwoeHjuo4bNwMiIRO+T97Y6/0TLI3
WOQxY68HsQHK2BBcD6rUe3rMxugIIcKwrynKfS2A4aJEUmdX9Wrr3iYvLXLNHxWdv+433y77EccV
fElIJQ6wVe0K5hlBjbLMZf3QfDmzNWHCEXPryRMpqBZnDtoMPlSKkYO0vKCEz5qBDAM1DUifnXDD
MG2f5b2N4OKlyDKLbGTGyJWAQZOBgV1zNNdB7HZddf4/ORtiLZdSqMQJNaPPyyyRy6JKXh15bVsV
FFuRINuTTApb6P0GlA4rfacSpGyr62yo76kTg/xVoTabANJCqC8R0TQKfgmqeeLotM0v7i8T0Vce
ku7IvHjoRuO0vklCIDEtY8EykuZJU5VBYv9ewR/AIHQ0mD7s1xUENLzm3uW+V9Ef1ZRXqsmPpKUB
ax33LJbJCguesp+l2TQuqksxJA0lQA3M74MUtuf1+8GltYfPfw8EQgpXgA8vT5Wl7z/Laxg+6TJT
oD8t1qH5LEPm6pfeT08+QpGEgWTwoK+ilEFoPcWJ6jjhnpzEnEihMBpb+TwFbpDO+9x/HCG2gjid
k/MUlJ7iuh2oZUnriTTdsWH1uGS6ac3XGnt8I8/Ii67o2vhaYGCijJtbYWmaw7Ix6gX5BvUKUlF5
JY4Dry4cscGYc3Vg+v7kDGgR/GN1PmFklsQq0azQRC9IMk69O/I+xJCybgqEQFz2FgQZXt4YqI88
NUOaK2AYfsXwdbLtZ6NG2vq+0hsfky1OJmdyLTzv5AuLy7jz7c0tKgj4LWPK1onCHhbl8974o6jQ
LOYGrGTZAprK8YzrtuvKOcPT9NSpLXoMmM+qN953bxAK52k3QfR0sTZrxR8t2gMqcSjddFgcH5gj
8yBH+5yw9HLOHGJFOAqbRg+NbHQz5jKJ0FpAeTVGMTUbSt8HaaLG98kYGdk3TVje+rH+D8gU2UIC
PPlinPr/d44N0OBgA155BLNXEO5/MigwKLRzQ1bWCFZvl/P1nC2YOxm6iVMp1CpmJTU8iyBTnsUP
PoGUg5KYbwStM9Tl/nPMd3YE23C978zroAeoBG9Yyd0OPQ13AjsiMmOwyjyH0+LNFZzYc40N1G8v
hQtTQX3fwp39E6FHKDpanOoO3x4/PFMeX8KbCc9it599qM6TQFrahYMHxGRJDpD1Rf9LSH5jJpkB
UobQ9mrNcVfIaSIn2Oo9etXnQv0Ubu19yg3T0MdC2kjpUomlB0lAgS6Y4iqS4Ydi/r0nqQJRvkfB
jVVMB4UUCU6ppUEvPlqMZc9mY6S+N026CuosmDGE89CNq6Ok8T3jbsWvbikcz5ec4qPDX9zLkvNJ
Hj3iwH/fPGCU457ziSnbcO9+fLu/nPqz+5MMuvLgYBVTVkKVdeiX/VkHjMyHSwM9Yzc1crXx1ar3
zyy2JRGt/Xk+SQ5m4eTAU4+M6/WCyrXA0vjkqOQiJ7D9PqMGHg5w3VAu/0IZogJ6pYn3ItIsnYo8
zThUjc41ecMZxJ/T6Un/5G7pe44m6M0iVAellOJ7Z280PEp2I1wt450gmWy01R/CdH5i7BHhck2o
4X8NFD9U3/9TNlQ8Z/Y4JlGrh/sXP1ddCl65GspombILoQ3kM7rx1rUS6JbaIBhjGwIP35rEjEJy
NiNgouiU+OS/U9pSId2zYhYeAyhXM/ov3sorz866hQL/LKjAr71G+qUNDDwV4LSJndQaQ2Om1sD0
rMIjmWygcqS3K3tjQLC2WoVGmMb0tFdOqFYrfUnIaLt+j4QgMqrKlvwhs4Z+jZY88W3/pkTKgQjd
NVeA6x9CGapQulN/pFdcxlsZxJjg5nP0SAk2wrex8hY9IQy2cimI+IopToRGdnWEct3Oa5h9YPrB
zo5l3dnvASGSW26RNCNZOFsWlUidEJg4vUA3epNH8IVvAfJdBK43SuYtppnovO4rJ1ErLmm5Dlle
smEyxfYql9MxOCSZ7FkzqGhTYInFyrkFL+mFRPChNL3z2i2I5N7AoJUsKpkvghMSZDk5t+plsdpm
7xUEejrlL2Zn2yyWnNI5GHstAK5sfi991MMWfmkPytG4jQRxB3OSA3633qNbqBmhonXqRErJWtTN
tspZRJbbEHgnVUmrnZ0IToFvaKUBIVC9fAkjUt8vB5EebbqQg/qTveQ34QToP04shxjlBn79Ceoj
xLJc9MBQiwdabUMJLJu87rqa56sJC2ESByAuOXycDWW2QHyNywloIMbQStcmF+ZjgpVXQKOn4BVH
M08HpsYbDZyBg1uFm3lgeEwptXX7rbPgM9ib0ZglZJ4jri/37MrUnec8wtMPlOsbyojKRS/fy2Ag
MD9AGI0jKxhOKyVnqOjb1t59M8UbGoacGSshCOsyMeTvzBuhJ5XkuVcj/Jv6gRYI1V7EIB14/UDB
p3qwmnBSRmkQloXsR/lK+3go2xOsDX/ZeBLdWXrCvx3pBvL3S6tGq5dTOq2naao0aAO/e0fy7UWX
NPtITOOaRV5zqcODOfulbxqeZ7mMZsTyTe/Tjtj/X2/p3gwN/rWpLJnanskhYPJsh0UEtIsGArMX
9r4W1qMF2LNvcnIjKTsqHirwdOK017f4kAIf+7Kyu8fJd3BwkIm2yKOM7OGt4VXXd8QxdEIsDDI6
heQKFxESmevMGjUbjDC5bKAc7YdzOExotqK43jZqiOjjpldra/qj+8q5dGVl3GbipRFyfP0w9aub
GrL1zMsHr8F2fAjydCYFgH3Ke9UiUABEio5+6vovgdzOaGD6Wsw6h0EgMs5jtPDEch7Kn6v8v6rj
k/nzKotj8Cs1TGv1iw+JNXN7ucoWxCSWu9FlmrJMADEQVljc8To/WFjljTBFLn03s07KIHMyLztb
PFlhDuTRVFBKLIP1rY8i5f++3q298LN2rzA5Z/IUv4X7jY6tlxRFJ8TvWtpMfAbgTiCThpG9iZpH
DXJLe9QdmBTZwWfr6xXBQw+n5raQGncQbtuJ3ybblbO1Yfo0CYM+AZdX/xckYXXMxrgd5480H60Q
Kjm2IeymAe/53/OsaMRPUbfAZqK9BaNr3t7Jh4Hy7Yas2Wv6t3hvPmNzhh139NsyifErn8U/lpvM
/lMEFlC8vVQ7coiBPChEA7WGcJOiJrRk4vWnCdLwdfbZ+0i/U7dVauaufVFohmAa3VVaClmXxzvl
62eztatS2Uw2sRJTwprEBJHQ9QtwxFh+DBD2WwkDs9HhB9f0p1aIrbxtZzHburvt7hCFL5qzGXgY
N3rr/dixFYB7a3iJO8HdRTR+15umq9GkpwodHLkIBe6IbC3jRqtRK71+R/q+KK6F36qnn6q+bdNJ
i5DMe8diraVa0/aNtEOB+Oim7MU5nLCYp2l9eKivQ6aGEwMEKqxtv4IAw27m6ieQFAPQeDn1fzzr
WfAH2HkH69a8Jw1buRIIXul1mEHjXe0/IWCSWsN3haVmd/GHRw1gOVI8WQldKzQwK51UVEAb/I54
OS1YqbmH5e1jlW2Rg64LlRZHn8hylKOEleF7dJoT7ZoyQcyF8YFEjbGodY5qUrbbZ1lBCayXh+7V
4KpbP9ehHK+jY4cJ6qdoW7OABv7IIaRNSmj0xk1FYCFszKg8mw9kB5SIt+mKb76Ueck91ayc0bt3
v9EdJsoeb0SDDdRuN5OPIv8xGT0f9TD5Sy2V2UO7R9SSFaAG5fXFk50yMWM5iJUBpTtfA6/9SqeP
ScNjBy2tTsa3cNJCBrHAAIL5ZSzF4jl7aaMbA1oI/6c+ZOu2QUtrffcafp7uhOWbu950cywWCHc2
wVGS17fkr6ds2Qb5l0A4Fu1Nsyrmqsk5pBA7m6yxOIwSxerlk1yeJDv8J+oDDfcxuJn4M/rKOg2W
om6pWbUglEsOH9HwbGdArOCCRkGuZv5ykF187HEwKKOLAfAArWlEno+ZTSLvpbiX4h72b6kfnrxp
w9xTYyPaWpS3T3zVMe3shsyHkW1fWYQDjrin+yDAfIS44GfdIiAXjC4SJbI4yKcz3CQakkZ3MXOw
H0flLDN+HL4LWYrQSCCqziKq8tjgEj4wVpItxz994eO4vGnz+K3lDt/Qnt7WCwTbSfdCe7bbEIso
+Uvl1iIQ/hKGLBD41RZ6KUTTBg5mjIRWmDiuzU7BM/O7L9GMcCWPC3tMNd9L51tMAtzQT9XiJHby
g+CuX8neAxUU2U9dRBJBZ492HqJGXm042KRQtaGLc8Idfzw8mLGeTLFm/nRmtewIX3dU/TdW1cvv
1f03Sl+87TSSzHqE5IBK2H7GcvCamrdjG09263o3SeCQLnnGpS8q3PwGLxY+N0zakseD/BsX09ok
3bP4B2eDkxHfCdDGSvM4Ozeu9i9lB7fBz2g7ZJQEygS9nICbIWxE0ncbKUFlyvraJHz26/m3y/2c
8x2wWLk2ySqUou34WaDbd2+hv1jbfXqOWFhJHUjf244ymiUhD/mLeZB5dWngQEMaR3v9KsyIQU+t
MamT1v0RHDQDvrTb76s0wistQ7E0AXENj5c5lzEkx7PubdmDrmxmxOw/ZhVeNBXQeHD3SqlxTt4f
JtOUAmPZHx3Hiud6HQbr9ByShTL+TxnU0Z97pXeS25r1fKKJaSwd5GWGNNegyJp8OfaW/okxxT2I
V5yJ67W/N+aQY4Ho9DwZsiS9jFp3igebSkvqi34D1Wo80PLjqO2125INrP8oQf7w96ym6qJcc5Ql
Z4KOtSY7jto4m4yos+E6XAMqusaHzg02eLjt/hfbSgH0xv5KAQ8Iu2mK+KWBLbyOumU1DOA13Fci
ygCWgrkKvvOFICTJDdCuBjaZdv+J8I4FYNubl1F+HXnkEpItznNFu15ziZDegRi8hou1XFQX0f75
Hmqc6Zcilxi+O6WmmVmEe+gHF2Nk13A4Lkq3dLNAWTNWLoN9spsGLTCBRmOdF1QrsbNWf9YDrouZ
hMsr7vG+1IVGD0QwMZnKcRK6hK0plL92+MrhUFYZFw6GyP+lrOxmT1dfNbSWWblgwKTv8Sj+zAo9
s04ceSeMsodHdo3GBRLT2tZEo0IWvAwzsLgDb3xjxaOvuqyCVhbvzSB04CxVOKJDOF9eJqKNpV4s
X7Nt+06KsIbUZYBNjhRlZ9dROucbEF6kk/Nw9dtCPxno1T8MgEl8XHpVWni8dBqzJMxdIon090ka
ziTmZJLz5fZQ5ugwKXByoGHqVV6FWfNjzxHoAaosX9VdahvLpwykIJqtC9+Te56Wv4L0MaeoROjW
QQ8b1Tc+67Iq0ia1AwM8wHGMmBSlfA4p5LnkA3mDcYgwwjVyp1swGJGs2WPI1xpx4xBcVmJ8oFyy
WfE3KlUccvwjkXJYC2/fzHp6qejFGbZcWy7sAxTmjVyDC9FqutjWLv2Ftbw8NEYAsUnAfftvsoKD
XsvbZ5APWIh68MEdY3yHvH+vhNGzlJ26a92d6L1WuF2+MWgjXds4lN4ZFKB/5PeCEC9TdzkHUFkb
eHAXdDRtgr47vdKIWke9e/3WWMermdmY5xAkGh/XXHU94jHoumdXHeOVxq6FZlOjgeLq73S5juRk
jtSVszr/RXmXD6lpgATlBmVHAjXKvjlD1ywNVH5Z0C9PCozjCtQsHyGOWUlEgPT4TBaHtHKCXel7
lSuJlsFdy/kLKG/yuIaizosn7jtwWyFQQOi/hqJ3AWiVGEfHm7Zafjl6t6azfcJJdTe8EcdPexhs
JbV8yX7g1dLAcPVzx/Ac00PlBykVa5CopHsWdChqPvblS07YFN+zb5/2ZDt9ALcX6oDC1Qatp7nC
gcZx7m8Ekly8K89OpXGYf8fGsrhro0fIVtwKq2ezgZjGq1GgZCx1JmM7ydoO7HNk8Wf3iuvnoJ3b
4Ebe5t5VcB00LDZDEOLs/7cJOO+uibDQBrqmiZ8+C6qvbgJ/bdodetj5NcflMk700H47iCmFqTyr
l7L9wBuU7qYjP5SN9sO+gmqunADKz7bL8bDmq4xHIJ1fAHXH7qcP6ozWpJx+AB7PKeOdpaeqKsBQ
eywTUR5G9ZyM/bVvh0gOg/dV1RM/bDgNWmvpCWYTlSNEiDRjtmioeYW459Y++LI7ZtfodWDnbhu7
vrvGZ+PlQJjyQ+KI8c3uloT/emzKbaJ8bxWQ4FyPkXTZ2x3dBSWLE/poitovnn2brmirhNEpZ0Qv
ZctoZg4bxWy9rCcUTEtTOrhTt/CJf+DCUeAm2gkRAlZHf134v7Tl0Cz75CvrGlp2siqEkoUzE0YB
aR022cVNjJl9YLuReNXZOoE7wAzR0sdV9JhlQoEhJYrmbv7Y8NCFtyDTOqvRn6tChPA4xg0HR5qH
EfR6eiJcA5Hq+hTf6SyBJVS5ZLnLNjqtr90QALTPPMgAyMMONc9bGN+hR0baDXYf1G2A32jUh689
hNnwszIRCuuiOQVu2zE5mJIXKYGald/hpSDxFG/gUVCAzG4qncVBTKQzzwauwssKAhIUISgiQlgS
n/osdykLlAeHGRjQiwnpzIMxfNQf8sKIhODVR/F/0gmjS+EBtfzgr1ZiE8hwkyq8asTnu27tG0pU
/a2GS0riosqtvYqjHYi2yMLZpH/XAMvR/rOIasEBggDvamaZPnuGgYNTtc6ImEp+XQkyM5WXPDmk
4qiDsJ3WcCht9oUrMSLZtXy51GunsmPuYKSkaX+6mhh/QvchlcCOt3kYsSuGiXCZ2T7BAe7MqLBS
t3efQE/Aa2KFhjpVIEkw0ISy3wCQKFYn7xO1GXLDnx953tHsPCz3AIpQrppByAqtWyowv9k4sjCF
ArQfbtMcyg7DSw3TIP69xVgXtWwhicHBXhF9LloKIs2CD3dbGPexM1Ayg9UKIG8QZQEQcpIpEg/G
erFd9k+cRfof+d5YLtwE7xdSZoQCJTGu4NEQm7O6GfaWVXhHtdTvms23fSpvmPZCzIEPhut5RLEP
8imtKqi5yxm9P9x2IoKoywsAU3BmpaKQT8RJwTelRkklb/TTqdgk7xgs78AvpeYF1qegYMH1BTZP
6o+16Xeso1qMNl00SyGaUFp4yvZPq2c2enLdpVLNfkqNR37CCQ8EL+fcT80kYVml3kxivWMIuduj
bkhIdBxESoum3tQ7tytWkcNn5w/zh3WUKDqxzKq0DwnNQrIzLGTX9SOJvjmofvsniT5gbb6Z4bBw
CUPW9cPOUHuHq5X5JsUOCx1KV5yDaZUMRl+1UHJ9AqA6Lhbk+wzILMs1EC8j38IjHtWweOcO1/o2
IIUdk2FasZ9AtQk9e6t/K6FeAP5PTB7IpLEATCjRG3oFJV43nXkzGI/JyIA8Sg5KgE8+KPrsDNEj
seLsBmyAsuX64SroQZBBiWgTIm4pGzKCJzsKa4hEoLQEbmTpTvIIy7rNtXxZLZbxSgcgLDVt5OhY
euuKlFQ9EABCz5jvlIswJD4rDtCauxQQ0LqctgQ/uY5rOFznbz3PuY7NlLj+begrQOnq7b6tVmj2
befOyHAZQIoWYeHF4NX7sDE01h7JQv1vafncLuofjdoPcumfum0Ci/19maFXivB4WFPLiuDOPybY
IbcYzLIG4sGeWclJ/ebqsEZHvXLqmO6/AAKJjSMUGRyNBL/GMBUiYB1x+EkDPnD08v821aBvWjUP
KICLr5uYPenhHWXJZJrLQ8KPq/VrKfopaFg7N304HIDMC3UFk3L/HeBdPnEJGEFF2G8NImiEe7pj
/i7SxCn6vhXDJo/9bqdJEhsvFfitcYfE4SRmuPec9Orn5qeyZkT/fBovqCYe8gKRQ3RY0to2ioFm
AzSC4SPPjJbvpneQyQ26lP5GKjVgMqQyNGrwlCV/DHcr/k0njxZLekxRrtTc/HOpTTE9v/Zfs729
BBJV3L4xh8wuNiUvsQ2gdFwPbO5G51TEo9mPkW/UiMlSi7nqMCNH3mtptwhbD2pOn4FwHwfnJiZA
mUVxoWwoHJBtoAUdUmIcPZNmOvJM8q0HmEXuVohuhwAoyiRga1KlQCizWoHZ0Yvay5WBgw9rIbZY
IJfHsId4fMQYkUvLoRcCIE62YaUDYKmR7Gi8e8z8MsEaIOv2U4CnfyypeedQKpEjsfVTfh/fX32O
rPEW83eFhJq2X/MV8uvhFKJx3XlFQIkq5Fm/9E1y73vJgd36u9ULiw8pkZwD+86RmEVGFBIua9Eq
B98hcc4AfmY0kogCkPqgV+6WugdBIRQ33mTE7hBHkF/HYCbaWBbfSdiLl0qtDVMEP7/eww7bROgc
689YL8ojOLCJLKxo8q7sN9WAcJHdt86bWSvAfw6Tlgr0HaUginTzHWZh0b5pGGY10xR2b8g0hfnJ
faQIXnHgDbW/c9iqh/QSqtchyQHxk2ApWDVAbvgafmln6cgB2upA6VCC3oP5nSZUoXB9tG6KsXu6
WNReIOVrst/YKEqTpkwWtagb1JgF32OG6xkwQyiEa1gDzbH308bWT4O2Q3yV2viI1ITv2XfSEt/n
Vd3DyCWXveeHOP1gcsN5dztddYU4tuEqW/ElviMongx0KUykZP6TJ8EySt2LIu8y0tBVKqWSJjAx
67PJFL4QrA8te7ReoWZUBt/LuJQZrB0H6LzaKir03muaIhd4YttpwWAvmXLT/8LHSFxCJfOgVKgy
isZM/sVLL/tPoFGLETaGWFMyEHtD2+gBdGihnjxPAfMC2C96BAF/CxMCAtLHIXObuzlglF9AW8ds
OtkR84YVQgkYL0aPJXB9eXOpPuiIXx221945U356HPNMO0Ir6ycNVYVlIgwNDeyuOo5K92JVhdsb
RHxYDF3V0mXK86x940Ewm5j6t9nYcF6K+qHBFPUH+Oy7MJEzEKzrXBMIPZdTItsIEH8Re5H7vCP2
mQyIFwqFqEke7/xrjinh4lG5yFrUVu9uSwOqwR9oXsN9ntUZSeb1PGX3D34YpghLodezV90l3hQC
C0cc6vI3xBFiZyfcZhAGJjoLUt5KAuUkPiOiAYczdhl7VQk1KMdtNM2oFtxfgC9n4Z6nQXafY651
F/1aHUcVT0+y7REqbKxhGoyh5t4RJDRieKH0LRvSGXC8geh+I9TS1oyE7K9YyvgtswC/bOHxoHk4
mJcyt2FK3tSBZbn58TzJGRwd5zVifYFQBnOxhVBX3AG8uDgK9o0xFDTzYfGSx0FzL+aWoXA5ZmC6
fuUYGJwyFVNWmNtQTvFs4kP0xBTB5Z2NmWRxLz+/RDR2g9imxFA5QVxFEvHaKvvO+Qr1d1FaEc9c
tYZ+EX9rUj9rRSHFhYnlbnYRGQh9VEntvNox8+I9JvM/lfYbxfMhm5mHoDuFLf9rEwGTK/26zzob
k07hrry+nbMidNqKLG2DMeHBWFTWCHqBFGRUz0JzuZxfMkNxJ+hMer83KEgxLCEOF5jHPs2NK/IW
s5qD4eOBJsdXBiTj3ni/IFNq53/9Sy5Xi6pYZfHSviOAFrXjqCmx54WfmmCW4EGUykuS8iFRtXbn
fpnY3T0Q5xEUf6NTff4lH5G0GyTnz/CIOZqqekI1xBho6ABLu1dV2E3feP8oHMVIAn5aaBnYtomg
jz9yy33U3yq7yeQ/mzYGlEf+LgWMvf+92NxujWKJEI9XN+ZYgBhJBuggH4xx5D/euh0w78XHVPDY
AfhKTUpXqzi2ByB9TpimSrlqssg0zbZ/Hl3TUew1RwFtogDixNgr1Nb7nKjCcCD8d/9aJTM6N0de
uBd8VGgyPUyFPSksZ4tTnyiXh0CesEyp+V+E0T5r/PyXaK8ueeLpNDQl7VcPnBQJTQwP2lnqjmkg
2gLdqX3tE2pTY7zF09QJdWJnCkj9/dwyUdiv5FhNcl8wGAUVfN0DWuG8bBsudS/VDRu48NSHRpVw
kZU8FPmgg3W5mNPD0CI5hUtWqzuPwEIiEOa6ZMqYK5jXn7iHkcg7N57KMYWaCd+JAt+axZxqYp2t
hoixeG4ZVZ7khE7UpwViRJwh+PU4jeD7WYtz8WlgjFabyKaUzinq2tgwChns9kKCFffqOZzOfb14
XoW/OUIFOyczd5mk1sFeCU1Waa5zMHOquQXKbY9uGsnKGX3XOmIkrAEe00xiOQPHyGJ0BAGgKU1r
O1pYN+kHecgksOIwScFkUDTc0uJUoEzjtapqD6QUU3tw3dRM2GH1NAnm0QmpoQroZ0957D7CkiRH
OwpnHpKFqEi1ILXeeAqR7orH22JTYTzgYfw1x50Rq1mkusVYENGg6EieNymdBpOr6k35YhBHERir
fSrYrPlU6GFA19APA5b85MpTFjg7TiLsuipHFQ25lH2aqbiiNH7rQvdGlbRMALfRkbVjycRFusUH
l9XpYim0yPPzEFyH+Q1AJgwSVJBNgsJTfFlu7lkSd0ZgFEndnGs0EZMYhiEKDQPZ70aTRGnQEIfW
9DnX4wP4ngnadPhSqcER7OUwydaWdj3DdeUBX9j8bSGphLIs7qXUQjPuGJCY99EcS4uNbuf9YVfX
dn4wwrf0+4vG0ggledp8JwEoxKtDUhpM3EqjNqM9D75J0CwroNN6S9ILQ0LFjbwfXuPqjZJeC4gD
RU53dBLb/apVSEDkZtCTIfXFihvXZTlj7nxE7rUP3A97QTlZnuJukr6nVEnr9tOkfQKqRAt5IBdz
KfsM4UDRzovobDdOHHOThtkjCMAnE2u+5zvRUy8Tjq/c1R0duCkjzeiZSHaUe2whTAgyfyPm7+95
FPlqGkL8snfFp6Om/Vobh9t3Sc6Fd22WV9ypwHExFxn1uOhDoGtabNprIR3FZzdyALba85t5zogQ
qWuySRnUMPV8rTn45U+ArLnqKsjUvkTeEWmPXnug4S50gS0D0XC8lgmx1njvVyJIDreLaTuigo8K
HzprMYz84cQTbFbJM8fSD/4yX0VHb29gxm+7DyK5+5ABpQArQqSpf26fJe3yrwvokxghSfFvg6xS
KcgTB8Ye3M23PqGlGpXdXgN+kp6tRKPnH0SFp2HQ7g2P0tGrr4QrILGwLD4SG7jqfDKImBRh+q77
dBbELDebjBRyo1T+OyLBN1tQB5wbwyEJSABlRAoGZpHK2VQ0mjXPs2eDXQ35BvhU3ClQpIujWYZR
DB2M0SWJGfxALlfkgVUnFZFARFHnPQxIfAeUatMF2+f3spujTJoG5++8IVDA1egVuG18BcKHFbMN
oEhnKPg98yfv57/iwQX1Y7sXOdbwUo/16CHMbgyVFr6ui26mpoBr9O0aV1NHtMu3UVeTdQZMHVNy
pyU/b/qhJV7WA+h8BpSVDSLl/jfjEvsEmZxpRZKcQcUhFqM+LKcXuWNHAory+8xg8JPrInyXday0
zR0Hk5BGRZQIMtcKtzlrMIDaENZ4kC6pfK7pdwDDsJeotZTOgYi4cc+8Z/3MrtPVXHTiE1fzNJIh
gCXyUj3iYSUr7Jf+p0CzcbPiRL4O2Iy+vJHXq1ygB2962VCiWY0lDU36JK5GkDeKpJV1XxFDZCPn
G6etJ4Dbj08kgXFAejtDXl9a7IIxrmePFcsIMYYU4/AnXfwFacQ7a14vRFBl3u4yd1JZAKIwOIpX
ebx1Dp0K/3Q9BYMt9ETq2AADNsISrBGt3uKpoTXS+OMcs1Pv5KBsiGjYzPlpNUGN43UBLRjWGEIz
jvRWA8+ZoTZ5c834RvSSt/AbAlLcnjX8gmWGwl5kR24IQts650plQ44HrFHwVmTg9WetWWIy3HcV
CH/D/Cjq8W1ckbhp6OGEv5/N7xC+VHHygMKw+HtXVk7uau0oOBrZa5A463Qvie6NB9E3C/OiRTak
XAN9RXJWH6DhVohfeQl0cp8ovO7FwJNToqtw0+b/qQPHjk/rMRPDrDo/2uokgO9mgX2stRXlERIz
D1DmMa7AJc29Hs1kgEwwX7YnF+F3OCW1NQYpnfe2KEkB1cMbM6e8Q8v63Ra2/eW9zF9Bf03w0AWi
ealyPxBRDHZMCTzu1tcbWRIXTqXEHQZ79VGWzI0DTG2+61xnX+9sND2RK03oede0NLSBo0B0rtG7
zrAlinH/vd33DSeD0s+9e7pjfukZZk7jd9ooO15tWTulWOGPZ0s0nIQtQl9MT8U48ITssvwIGTUd
IWTTEnwmQk4UVJm7CoMjFARiuTlS+r9XPtWe7dDft6raHlr27BE1KejO4MEEU+/dYw1pC9cRaPzQ
0fSmOS9euMi2fhfjGlvmCihTVBrq5QsKl4YBKv+xaj6/q75/UMIQP1qS6hbCAZNmbQJz9WzZ5UF6
irzHbEWAd0oD9gnlVF82W+1fWHR7KNZwO7McnNodv940IusVGFzmTVEs1d4qxWIdc1QaL/10XA32
kFV8hOp9pgUtjDaIHmOl8micwZxjSF8H4G46yEE9Yvl7/26k8093DF+qPMwdWNR2qY/HtVPkIzTl
82yZ7sqxZ+JNvvKxV1u7IVNtsSx6dumsn0mymJDITu36i82hCBj58e5MJUJM3fCdJNlC//HpstLE
4bLCtWw7xsCinZY7dOJGQ+0Cqp5O5nBOd1Khi2246a7XSQmGBaBeyJBhYQ3kzsEpLDogvoEIXwPc
w+T8E1EnpfYZqOSbZz1Bd/soHK9KxWhhZY0Nq9vzxq60ZptlZGLgrckYPLlECoqIS4FKsxvnf8He
4Dwx/oe+Ir1uxkjibpsCkgeW5n/fE8YknKltafvS1Ypc5DTj248ukrbAkRqgBZfpdBJ0FpPtdOI/
M4+WnicI88xCnECBnB1CVNpw4TCvZYdl78x1UDUyeBWBmRyFP50J9lxo9Py80qT6NsR2tU02FWyL
eetu04qBAM2VZSkP2zUdUun2TNw9zmBkgfPHd9gPFLDyNRAdD419JYs1BPZgUs7PJpSONzAN1/El
eB4suXmGbjrSv1NQfy27JcXHZIVgrxlWlRxF0kcu7+NAF/UxKKXFh5CytPh1R38s2YoupiDo6DTr
52SCib3OQpdcnlaZxIbBm5VD4cO8XT0GdD5ecIAxFX28wCSlc/pcDp8z3U+6EGNkWcvsMGcsF4w6
zUIRHrvggxiVbe4GQFK4A8DBnufBvUrA1rlRqy88I9PN/FA27t8qyrl1Otj/1JXB2c9/ANpOEcdT
wkR78AFS21o4Crvj9d2Odx0AOyoiVl2NlHWsW/yuaqIDVzgPmxBKRMFbIEcNuUNi6n2dYMST3rKU
0qJq9ea/50gfEtdB4953fxyf1gn1zt5os6RAytW971meP2nORiljXINeh4k22cwArcLhTC1xj0Li
49RUaIAbaaICue4xNoaexnU4/pH8vemIB3Dn4l2SojjF3SqdOWEKyJnzZcQ3wzLbmCAhePN/vJ95
ncUL9kk2gRsJb3MIsjzyru6RW07BHaidXd7qNUazs+RU3MpIyltJeq4mTS7GnZA2vu/bEjvgCf5d
a9m52YCPJ0x9y+p4UEG9/SrJ1ZmPIHizXGeftmWi3XRP9Tu9K09uC88INNEhg1gdHoF4PqAn4gOK
WSLrnYxc+LcVGcMd4dTqDO3VwClLlk9wv847RcoNAAe6fwTZz66ajGIfGv74OkLJI6kLqcoXiUXb
n2hGj7N96/x/gQ5q4jK48tYpAYUkkEi+oBGFiIa9o4tuE22IUNMf3itCk4mj23PNkiW/kYMwoqnE
sFKrI3k1sc6ChuChhHsK3nklaTVejBP92sZjm8yJTTUlctCJfMW2csl06xI2wYAASeJ3meafgXTX
pW2oIO8fdjDzM4KQNAxX/wo8n2m+OURSGCHJnGpECuA8RI/aBLvPP8nE4b1tMbzll9O6Y8JwMgMl
PztRToR4Ko7z2Qr9Jnn+uVA48tjBaQx0+frsiejjOD1sIyk2h4alcaivXiwvnshfjQfPgOrawvxi
96BdnckusrRD3Jd9p0+/UpVEdFvr704Lo9xI/CMYqR2SjrwNNItK+mqnOCpBMoVFJaMo1WVcD3sx
QVNGt33Bm7goCR75ZQ9NWAf0l1Pu8RxEtTjjOU4WYc9vyWispR19/WC6CUMeg2kFkfWlI7D+EI3a
iHE7ahko7GrAp3cQOd3mO7/pdSgEfVsiz9OiZp/peQSU522MIotTBKRruLMNQBW/G2kHWrBFySm3
DCrXEER8ZJa4lEVK2aNpbFLBeDv6x7JY83lcg3CzCNC5wzkO88HlRTCf+Xviq29zuwWs9l9mveSb
KmdtrLxSE0SFH+7AAMfxLRtq/GWkUoFn0o2Bcv+D6sHIiYGetrka9wlCetTyZ2iRNnKSnKDavc13
hubX1k84zKW/bcJ595O/7lHJxZ7cZpgZTQnLYoWrJ/zeWoVLQD1FMdkpiax1+/Px9b/CYJ++z5qp
nNtPShyhCBd/Xgm75ryBKJos4GY0FC6QNvkdks6VeoOlCHXbC4QeeDSujiuDU760eY4yk3cpqY2p
VwZ27XzkbJR+4GWFCXBbXZ9Bdvkb6J/3enitq0vVputm/UibWE03qUshqZvwChzr2z2Zwv+/Rqdu
AD9hpco57o8N/wy2kK6+WOmsqWPLF9Zw2dApTeIpfJ2Le4cdqKcWuyKlj5U0aXlDuon465/bm9Pq
N19AsXSlwb5SGOuIdNud7qU2LD2rqNa1f7nuWJ2NZwYx0dQD3qnDuJglbdaatpr5YWN3uDzqJTQM
vX8oh3I2KSPXSFkKlIsJXaJ30Jyi4e6apapObOWnoAb+BgE3hn1+178Vzljiz2IO26dgU5qYayyP
ulmvHfEy+wwLRtVypRLUcXXok2E5DkKFBVND6KRhwaS+Oa+Ud+KTaR2LTrtfQvAU4qdhIRU1ZwQP
ru430pCTvnVif7fXN0L9lk6C0vQ98+avyMO6u4yC+DINl3zPdJM2PWzZe0rzi12DqJDuNtKdc5e2
g/uGFBhICN3ddy0QxRxEhuUpZF9KSLmHk48zFrVJmI9QvKXxpp1MCbX9uKPzE9Dcnd9LmOqF0QtL
DYQUue4MfxU5Vj3UeOt/JJV0E7GAG7hN9zwK+R70j3vMwii/PKr4Xux1EOlJ6ntpUN4DO1NKWE7h
RS1nKEtdWolRH9YXeklHWaYGrnlhKzmDGr9FZmFn9m8j+C8Z2edJHL1//Gur1Y0RfAmDVunIlU2M
G6zlgR78/7Y9lWqhMPVLy0c8jbRSDaphidbrlxcMgyV0Fh7Z5U1blmf8aYMuEaUy2QGxg1ldzoAu
edp43LQddGcW+WJ4xz1b+5xW5/FQjGoq3vlJHJdpna3Lt9bpbJpuUjiX9nEbyF/iNu4hXlV+D3ae
49JGo/2wzGDi5tEK16hi49ikEcjIWYxOEcCBzIqK2yJtLU4yDild5FD2sa0EmXtriEMKQaJHZtMT
8n/pqsP6rez9s0/lxQNthcOYFWjdQfHVknRrVnV2PAOTI8NVfwoamgWJI5WkmsOBNVDWothCtEoR
+DBlLtrjEUUKBTs5YqbEvGzRxCVhd194qwUJpiYXeGtH1JCRTjfmD58aWN3ZCNF5zcMjDAU+WlLh
u7fk5HOcmZY2xS9k437KBFFy6mb3JtQjpUFJoRYHAh2dbO6EETn4YiKBxy/b3rWBLDrG8KxHbuI2
QVTG+I/b6XFwr3w8VikqUph9At5eoZMCfhFO/zEuD9F+n1Eq5hNlFYmeqDA6Od1n3O+2/v7Wnd4h
kWDmKwNr+yeGwCtl5qwkcJ/Bzm47laoeaitRT0Em6kdtH+cFYaHygeP16/kkpuu2mhNGFp939maR
TB3OzHQ0WbUxXRNm5LmOIElVC1QF943ZUPWckxf1vHk01rdakByupAXTlCnQjCntxg/QD8cOXRoJ
uE60qpz+u9efedKK7IDxgjKscBYq3Xd+KzYFxTH2NrKTl8ovvR58yRE4v6ZC8eirGNvBPQ1Loinl
zi5tZbR1WEXbO16CUw3ZBlZPstp+XEPuiAgiQ1zrKP8fpD0RU9/bP8P2+cx8hAueOu0T04G2FC5L
XotY4F17qFNEy1rfettUi7cd1hQ+fdSqwdh1vh80rZENCkuZIDJPJhLx7LNbNPdhMLgSKh02TmVU
iGFPt2kRRf7uBx0SBfOZQfEVXfCwZBLssEqSxLiNCXEpypDN3DRS030GQ4OGCQkCcqS88U3Eyg6+
hsPx2i7apKnOv9wcJyGt+9EgpQm0V6V447n3ZYZQ787BYWAAqcJT9U3p/tuUPnBPooQ87BOqVdbl
H5DdtylzQ/HZasTpyezuJi7fx6DK5oL11iVK/L+ifOhPLJ40DBKmPBIr/6+oMLg6nFXNVqEeS/sS
zDrtGrHwrq2abvFR3HsUsl9qSoA8q7emIK/wYhthMgIARucqhobqMpgTlvm/KmHheZbw8BAmTjIx
0cLtIYrcLfVffoxDDB/LZD5nXngI5KkxWDgzq52sHEIFI05i8eSC1nbFXe20veqy4/1AbhfkfPYK
F1bNtLJKmQKMfO56QMX8C41kacNnIWFfvrWIakjv0iq1C6u8PLQuibSTjfElo8kiRXhk4mONEEkE
Wrt4ujtbVJA95+eWpIFXQMeBXIdLxGOu7H44/EQNCcXiZMp7GnSMAkNOzLBovbn/yfeAPJtyv4kk
baoYt9+Gue4gYvKyMh4SFqn7u+aiE7XFqhIlTw6uMsgbUhjmzOSt1m9em+bg+R79Q4Rw4qry4OJ8
ijOLs/uNiL7CqheE3pOt9oHUEUrWRi6alfpmyfY30dO2Ew85Rt5k683dmKcjiAkWQyPgDuKC5Fuo
EKUYceqBf/mjUNm12xUFtgk6bZilYWcDJ/gY5oK+gz4WCti/uUITUcF4/7rWKz6OLEogSBMQnIEl
wHD3hdhgZERL78aQhNTRkGTk+1Egvr7WT7lnTeNtATEllD1CHukXQr7e25ayGdTrzca0wigvcApX
7krJpxGflB9OapbkiL3q7izpzPPxILS55CZ0aUSiioOInttpB4VrsNEhE8MrLKu7c1Lgmb2QfbkO
eu+B5QsedXpHPkynZXTwjz46nE0AqB+qttYk4If2TywFhYujnMp8WZfZANklPAzpMM5Pv0UFrqEc
1awRUdNNeTPILfWsGc4go8Odozl7ttgvDk6Y5qiGIO/BKZ9DI9/VgGhcWoL4FW4ehv9fd1B5Hep1
2FkqtBj/bTLi8XnGmxr6lhRGuIlP30yDl7dTlyjXTMq5jE9q16ImJm7Irgqu7zRI1vTpxtUbXDGM
M9ZjojUHdvn8o/boj49LkMits4bqoXfvtS2flUL3LBG93z+sJ9N8xSOky01BLHCtW8eVxM1ujDzy
4K6qx7QXduAADUPVJGVQanpmiuENd6I2h7QrWwwy+u5fXVM/bwPiJ+OEuwmnCcASCXJBmoX8AXQ7
5nfY1W+v1ZkUT+yZn7x7WpeoWuQ1DjVboys7Y0wau/t4W8cvHn4zoIsTyENhdCX92U932JNufRJ+
5oz6L1dkOu20s7ed/ODGsbFGSVDND1bCFCSfzdzF5D764DQkKiPOt5CWt3NjXLnBQ02DawWxw3ni
2P6eaj++03shPPWeyfVhOjdRgRjXge3eBWmX7/rwoTN+RWX2dVLFsa+YuSYlUdzdBXZ6Fl+lNxaC
26WddtIwH4mC1AYScNnhwxvScJg51yB8L/VN52YsrMuAwECrry7P8D3QE+bjYHv2HJKen+kUkmfO
fGWx5OMxPTpNki7MdEGA+WB2oHdtQ8T1OKi/squMnkHzWCMdHgwKaLqr/OZ8bb58ouMLgtCU+y6z
gErU9/qOYfuGcqOGcw7yDAZ+HHukI7QrXzMq5WKhLhfpc6dV1UplTa78wA0xzfRZ/4CQXJoUfoSw
50phTiUlXT16gsIYLZnWsqEG8nqcgMLcxDx+ObM8WwrNNf8YkSPf4kE6e8V+1GoG2JMaGsXmDM+y
vI4kL3whaTRvuFCpQYKDBa3989+AZ+lpHKvlvE1AheFK29YMBh7B9z+/TdNd9I8qvL9TKStjEVaZ
CDOFJ6BcNK8SU4Wi0Frd4s8xby8ofM/YW/Lt/CcHS8Fi+WMF1M4ZoLhxC2Fl1jhxpYTkMoI2QZ9f
70bbMcIf0LkbqS4lExdYysfNsW5VddL5vaaK8MGIc7NAdrJqybTQnJooWUA4agd79lZKD22wr2yI
BFTU4eGfAeNvezZlfekyoAcQWMxxmkwzb6qJ2AYsdkshm0D8oKphcwcHxEwGusYwual52jZDX8en
xnyrMtKy/ophDNnA6xb++Ak8l3k4lKWH5jmrDJC2tolO0xtREmHzJkRIz71SyEieeMixs7O4Tyci
6h9oOOHej1hRZVLc9RoNcRWXw5/Ix+HYiZXYKnQ2O5IVQsfiSz4kRyFIKl9JKasuoWvtYJbBrbG5
w2fdjySrRk7Klakftazb9JwmWfmuPs74fy5EmX/cUnR1AVz7xmRe6ewZBEGkr8P8AJZxuYSVATOb
lkaiMCNAUiloHXfrO5Yftsw1QdmjFn1VwbTN9LAhHOgBvpI1sxtkJxx6aULjyKvpJAtemNZ5bVGo
Z/o06uirks1wELzqWWQwVclb8d/fUx7ZnHFrIn4mMxIwCLUTeskBAIoMXiYBPIuHPh3CUMb/Wad5
m5ySXbTJEbDxNsdznAdHDMrO+t9ujMwusiT0Df0TaeDz+CuBNDtLU+ZyPyEqdiQVq5K/A10qTrmn
/UUKZSqvEBmA7Ww0B4FxSKVggPjTzSrDSVKVk8PFUYvKDKAnaWBaNRjUpqDEGH+4x9Xi2ozSZXGR
SphSBEkQeVql1gk7P4lCbbd/7g1TTG4soUAZO1g9uw+BDY2V57SXDc1J2/kxOBnNwx0eHUwKEM0Y
lT7NfCnnGBxj0iidEkLzBAGjPgkrIgn9iUBl4O40NQmP37xmimWhCAoe+5DKs8jVt1DLqbd9Nksj
Vu2eq79zvVfbLZw7v9UF6rM/LKRdt3DYgLJ4fqDYlfUt17gFY1wRZJ+oWOCuuIvma85Ghri0/hjQ
mqm5VHJMi+p6OSTPQ5Nh5qSGFdkyjThH5Yc956doLN+noeCE9WKajASfixZtgg1VPxRiZwJU+ybI
3C7yM4uKFAG+o47YgT4OKYjeyjurC2uNMQEYl4TPBlqwBShULdBrHLOwbLMLFE/fuRnun8VsDTkr
gnarTFfWaMaZEfCjMhiQ5FUO9mFDaUdZaQu+bvISohAKf50OJWprd2kvx+ujf1NV094uaGotAQ0Y
udMMuU9DdWl3Owqa/uMbL2gGFNuw2ereEEs5w/rW1zUf2RUs5Kzco5Yi9o6FqKXxPtt89HRhQgrk
ujyQYPxwo5d66Va9558L/qFcFFC2WgsSECFLpc/ZzzVTo5hQ2VPdS9Px5C/2BxXdrk9bWSk//qab
GSZF2H+aw5VTsQp2sJzEZc7RPQLyZMJAzb7WwQ1s7EAUf2Ss+/UJmkKQ5tfVuImo/immM/Z2QsPX
jzEPeNW+C9jbbspA/Oci88c77c7GXdOdOv7RdGRPxNNNt8luVs3HiPXvxVHfQpmH+W5c7UFQ7STP
heOJ0gMcntJESX8C0f9Gmd0WVgWaFIUzXLt+9sh7nCB8QvRgaKUgtASHk0MYOLL2CnZMhVa8ueyS
X6xdjJISiG2RdBMKrGQMRzmh78DwBd3EadBCasnzztDBnl72s4QQPKAR9uaeHIAOQeIMF8OIpZ6i
9PryCkjugOWUZTyk8NYzXrKk3UrxHjNArAup4zP/cK3OkQtBRFcnURvnFRN/6kF+MY5i/f/mrwmI
Jp5Z/Hq6DrBxvI8a1pvIB7nDdsPhmvCuF7OSlVo/H8DDaVM+ciueeIS+m7AJIKmmK98DHldVC2oJ
RFtAS11DeZMF+D5oA8Q4QBSCx9GOM9YM/SbWEefP44Ki8UL9caMjjzAGPgUNopskL+Kp6tqPJ9To
Ymix4Azc7H59R3WD/k0Ts+w6q9KxFmgtZsNJk50MtwGP/TAEHBJg8wClvR6goHZRsaH9V+9jrdT0
M0gbJ3m5bYXN8ehmf7LXXDfQa6r/VIh9HjZ9w65/agsRtpa90lYxXNBLxvk8ZpyWRMJheA+Y+IFG
HtD8m3Hi1Z5FZFPhustzol+F6SAN3HdoAz63bdilYw0H4SzcxR/ZZXBqhnkfTxgU5oPhqGj2INoG
cFE11oBPQXzeMnNHFLSsdph/K7cwPfResLDZ4sdKWJRRP8fJxdEDwO4bY6N1I3LFD3fleZYTmpHv
DO1p8RLLDtUcZt+QCnShEDO+Lrgiv1GjgpHiRw5H27iKbHVpytv1rss/p34BbPARQ/VNXtW8vLve
c3fEzxPh7is6s7vsQ00H8nxpTxxFDWY5YqYZQkZGY0pQXodSNpD5P6pnXgq7W/ZBEmcdQ/kFfeqA
xEIQB4rbsRrvt2Aqy9zC6EitIcV507pPFIzl7uSjErikzj4G77BAYMMhQrLpZqtu5MyL4IHXXVhA
GFEIX6KGuhEku11Sewi76334mpmUfNV9nXumdT6jM3Fx+L65WF/5+mxXYQn25b6q09DiEIh106oM
KPbPmiRmZVsQ0Uyyis7IHQ0orm9UOLF+XzVhnT4WS//Wjx2B2/cAYqXB6RSJPgsys+IfoeXMALct
rlGk0+Cpi6pk0By2STbcaSCkecpaFb/Eyp8hD0yZNyh4J/d/2O2IE0wCsNzhDKsh4fbBd0Wyb1Y/
ckx5sXezWjEWF8x65jtG2G5wbl8Olan/NTXWxTb2FnyGdT4MSEJ71WjiF/4YX/VXUqYDO40pSdu9
1eQLkF0EMdqostTrTZmmJ2Y9RkRlBrqEW9M2vIxbbiIlrHePxcPGS60RyGWIBz+N3QNWjdD7vkg/
IpeYWMFBn6v7Mr+WjDbriwJqOMpP5LlbuOV4ewehTD22AhuP5SG8bhpYgYuPQ2Qh6+2nK2kegsmA
w0B/B+i2cWULcZEHsXRIFEQ0tGAhGCGy29e0x/opoDIs4vDVBtj/u0AF4llT67YgZ9P1Zvg1figW
2Rcdwm7/T0KigcFFyGaUn+Lk1/Ur8PwKwEIAVQTI3LP4Pv2cY9EHzsev521kpfWgGskOtlKnpCrz
uGDTIWFp457ASKm5lfLOD9TzeMtAco0wOJmA9hR3B2J6W+n+yPNI4DtAlZf6Zcihz4Etg6y/sTaA
MhRLVxoC4xR0F4jYtXbM/TysTbMCRIK0ro/EwyNmUdo2365kHAphrROQQoQs9hEAgmFUaEcHLOYS
uCJal/qhIJbjm4+jnGhjg+gtxIAe+FDkSkn432qgPZ3hfukDR2A6dzfRlh6ac19KHtyNwyN3jgIe
V3jynggu9uHG3nNGhdeTGTeiPr6hoh6q1Yqzdg4KJ28s9WzmPlQUy+87BprphByc08rdnAaKUAQF
6B3b+8vlsRTR029KWcIjVFzK0FUDWlhAAdmJqXrNJhURAktohVvAuaUslg9S19fufCFaSch7vg7t
kzUQ/VNRQ2WkDO7aJ6qa0iomD9fbheCbP1pdOTRTXS2mxxX8fgUPa0fIjpBPMdDWHyHB9DOpxoqh
7zkMHt+7lE/50QCKzC7V/81yq+JD/VmwWbsgm2YR0Zl23+OdKjCwp+8vNeZCdlZUeDuEm4+pczRa
Gq4a1qLsjjZmxRHGmEQp/Eb1FuwBjLKGE1n6iyIYYyMjqq5nza8g9BF+u9x21Ut/VQnRGWFXCm47
r3r+e5GigevfRU12vr5g6qaR+Y1UNM9E6aB13UsZ1ys4vTEipXLoNdyKAkXdZI61BBMZ8uOwvzXu
uP8knILca8jHa28LnX6aMCvP74+eDA6RtOfVh6T4dtE0X649fVPjqYkUW09CDnA63A5g2EvR1UTg
0cM9Gv7Emw3o9+/7G0NZ7GeGXS8lyMJH9Iu9RInJx0UfbXAD0oeEfrxOTrwmVBNvGaJST9K5sSLQ
iQJOXYlnWg6G4JBZKdgtiAVc53aMc0ybyvCKQaymhalndttyLw7w+hnGLXKgQ2V5RIzAgD6kxg1H
k7RC8v1JXyWc19+c+up9EKBX+QWLzHM+L9qA3Cr47fGQs7b4VeguQkJEkhB8gDQIrxyUs7uFeJVs
tW2ECV6XcFcYrP2dJPGXejiiq/0zkUatzBGFQD/b4rDLvOTOdxCDUqUtQnVvfvVcTOu8vlmRZ/OA
jkTX2QYtyUkfC4QdST8emcRMbDF6SW8OKfIleX6SWlz5CqwFpNzj8wNTPBvRGi96/fEhUp9unitD
ie/iY9fvA87XODL+jtlcIt16EDiAQYsKgHHtMB2kcS3Jp1tZrC/k0hBFLvZjRLdbVx7Xggh3yaY+
mWpRNSDR+l8PnFHrxWR1KUOtJwjHh2DhS1GD12/YwWrajmOn610GO78tp/V/ZA4akPFV/1ozkyE4
Hc6r5CECu033y4DBUjFRIxxAz5qHMIbgco5LLZDA1oUbqFPEHofD5GXewFYQcxwkay38KgXqtHE0
XJ2IAiY+pF822Iv1xYDutD90fRkBnpUjKHC4O3vOKOQ+9bfgibWN9+xVngEkguZIfD82k7nTPUzs
ScnjF1tnQbug4NyYOCJC8iCD6aATR3/+/1StcbPRq9s4l7seADyW5tDuf31JC9PbjlZGl7+X+s8Y
A/QNDwvT6dl4SX/HEGhE+9ss9/WxxtWRBSEg5z/l6DVPaVdDVy2jEOUiNZkHgWawTFKFOLUbjI4d
PN9C8yxDYEWsgu/X6dr2R2YbbRTNdvhfBw5EZMdilhOAQPxiOPKiYRBhWs64wUveDXJkwX4vzWJt
tNR+Sv7K6ByU5VK8VcHThBnXI59+zTRcpJ7Q2jYE91ERJp3RbhIoMNSNEVo7+5fG9ycIQ5w/g2qe
p2S/lQ53gv154WFBVg2ZZ6rW0IrBErvoTrvoU5po0ucR/jlU3ygofUAwPfnQGNlW/xA+/iMoCl3R
A0EeNqEKe9f+oXyfpu7pUHUtomFO1d0EHHvy9q/+BJHjWQMBNNIs/OyhgmjTfG8O5EN/2MTnkYn9
ZEu5pai87gbE70fdzgb805PnfnM6AOXT0CR06QqA3gBQnQEVpnQehqtPGxLaSRT57N6TDHyhSsfj
WRq9qhlpVVm3133fMbPxuypfHK1QVDcj9oquoS1j4rT20EvopNnt74Kjkmqy/sN+O4bDd1QtzD+u
OOhSCiCuBfVbhARQ4LOxD/1o4hxJ2AJSkutjJ97DnV0tFBgcea0lFhk07N4OptJ9RnF21/0yzCl4
7vbglBwYUUBGGuZnDgXemMTiFtZ6f/DjC1QzUMRD3IWUa7AOR/3oDahGoxM3r8bN+kIqsan8Nkqy
4sC7BG+NgLM8itfxUzuN8gZJ3C+HreGsbUTnGsJTx3dWDUp7B09xkQjrcN3qOsx0owCA/rZqp2Sv
5zSK4y8T7Dhw2NgVNo4HBs4XCmIgqVJSbHgYlFYp29OOhQG5hEvpYog7Oq+1aFt1TB9m+z1nxjE6
rLSA/gZHCIU91Wy59Vi/HQ4+5qyO6INeX/rlsAi/O4KfsGTFrVgphkNkz/Bt7ZiDZWYxbmyvr8t8
EjbQrqFW2uTOJr114Rzx4mxxiWv7xfLau7J9vWsC9tXejbjfKYvFFjdN/xgnllD/4cHrQ6xkeKIV
ig8ecONhTIOV7v4j1vUccvW48tBxjfOjSNE0xUQZWy0DP+kJjJ08yixoXZkjpcu3Ly38riMiVtXf
ej4eN6QevTNSfoHSkuvC6DaFxiEHyUqaklVvpxacJlqGPxseF42NmUC+u2tlLA2H4hhWqVkAXHTs
E/X020Kz0sNVfsDk6usTqBtUM9miJXsj5SwLfJq5JXfGMGKZCRWYmzGucqFfeZeozkPcGeBQcxHR
5kyGOR16a1HE1Qltm5qcHJDNRlEfL+RVb4+oqdQmg9JmSuihSMoYVL60S+jysBDtgpK3kXAp/7K9
+8a7NNghSLjqLMtCP3Pr7RnBPWHAYW6hdG4FirK0uu1Uvg3Jdgl/tzXuATJrkGnbAweyoCjNgGhN
l6Jbmcp3e9PPhHJ2B7zkWtSc+NqtpId3UFFUYS1S3kd/jGETztJyPTRQ8gL9lHD6Ts7mxw1dYsRY
4XZEXEIRZiuHpvNB+KHnx0kqTfxelFIU1o9rM54D5FaqhffA+1EylBLOrQ6QBjKQAXwu1Op9v111
+0oanGEqY9MzAUp09RuZ4yiIA0OJY7SDdFLY2Is5vXjTQVOyxE58mDrv9fuWwVcdc+rH13g/4T8y
6HrG366vgBLyvEoF162Faeua18MuxJonWLsZUsu8jv1S/9XxFIeOBNfWYFx9IxoYI3J9Grw2BpqH
bYpSIw8aFei7eT3L8ec+sFRFfikcgpUHr1jf9gBFd/GdFH6WC3skMSYy/Nv50m7H5mjVFIqMBT8X
0zDoii0fTe6NgDDO/fJdtSd+UsNqFQqRfmwperSUubqFAxky7JLjySfvw9aOZVo0aFTDUcD/WHT3
ZtN4nA2R0GMoU3XyA7olDP5/8lFq9yVrkIL7DyAnLIZz4+BLOCX4rXhJEwr1ZEOWxgeUUGfwx2gD
HblfINU3A2M4UiH1rsQYEYe49cUoWp3fgfTLP04byunyMOdUeAr24+TSSpw5X3ykqyt7JXU7oCDB
5dff1gVhUDQLa2JTqBtp0Iazy3s4b3fraP2rpprCfyfEIu3HCjcaOXUZa4FbsDS+xR+QDPXUYvkt
iqp4vVde7Nppe20YTuGICXODpvaYu5tJUI0seR1y4LZCy1u2HgnDB2p5fq9fXoh1yHVyDZusWpCI
8cMESVHLg+KYSt4VRYnQz5Fl1FIG/lHQeYnVUC/1XQlIVrXZJCpv5bFcZZlrVPbmravjUPSCfVm6
4VksN67o4+PFqnP6AWUC/zmegFWabL1egMOmDLdeUOyKCNZVKnsU62/ZdXLN7quRM7UMn+Q8vX/T
LsMcICvTU5J88H33Z/DWCNGHEny/X8n7xRWvvcsDVdtHD+2EcsenCo/9mnMYyLNuVi5bYrTnKaRh
bgWbI9WfPrS5z25VvZLD8vtFdiHPnk25FUIKK0znGccA5k9iizixYFh64s+VxjwHGOnjA7GZtavN
JH0WqZR8v1Kj4sYnB69LsIRo1FrEGisgaePpigEQk5M6RB7d/XSEoRHlR8kxX4FigNHPQMO4Vudm
jp7z7SMIruqoPggbBLQ6mrk39G2J021MQTNUyeAGr56D8NosHp3uTxFuIWVFhPvUqcVkR0v296VC
O8H+klwjBpyqDUzJKYglqDrzJ7al16SfSD8S4elFGiwJ7Z0UPNXJlrIJCayych4ZQLoOgIIm3rxD
woCyVcqyc1P5C4Jz40iwB8RDX5sODZkYP/SwwMDV2DGen5y+3DB6htf/PhKsEGazMhixS5wMZyBr
/0hWSPBWAvsPyDAOa33dtmo9OLxTSuLgkkyoe2xM7OfL9hrSbYkW+hFFRCAi6QMTBFbnbWo+Z09P
aaFV2wosUN7WPmnrZelzclyqMfuXzvwNOjhnfJ1l9l0aWvQhGevlFBYi/cnwYCKVdzxnPdE+SFpu
HpyXrtz17WO7bnG9y15FUZSf4lEL63559hzIVQ1v7QkkvqwqRkiVruIoSUEnIDa/zhwR6+Aon98F
MH9W/HzZIRDKQoaNAVqcPzAEBFTxohJfzi2ycfYkqA47H2Vhd/uEhsIN8GvxX6enrFaamwy9r2bL
VleS4jhf86DVWP9wIZsgdYhCjmD0uyr1MW9ozFVERXWTEGgwDjsjWFrPwrCX5FtJazc6/LDC6kh+
lDTuB7WZBdNORCws3JGXuM6rOValElI+/qUn0W5tGIqTQpg5jUTAIHbj/5ij0pgZGdZX1OG43H6c
hwWMfIEFxj1E+lQdrJQFk5P/0s2IW+uyDANZGr2qJ8U5p8ja8SIVWsZl2UYmKb/ak413f7dWnifK
qzWER0MoK0/rheOClVDsq22Iahc56jvCL0Kr5UqYWkpvoXKbcAfnCsWnmCCo5Li1YEsO0roOsLxX
6pwluK5yFYWxnN7ujYlsVH+KKSNQafUYpVB9gvzUNzGVRyh4Olo4brSVLLFBzr5X8GhLo5ucE9bG
P/34lNcXOUHTfwoUC0us0sWpX+bbaflIlu/giwk8BysmCgtwP3JC4KeIvSHHrIp9/rhj+wY+9ol/
AhC9EZXaZu4jvYFeDyiI/+JmbtdAX8J81z+8exFPy8QfpA9pGD5sLHkZFjeTMH9CblEek1Nwv6Kf
CW9FZ7AWIAvHxyyRBj6F+PrFVqJG9xIYy4zDxnXKvtEHwdT+70pK7WnJQ2ubBvVbwXGesxaIZSYF
ueqvRHSeRj/Ip7sNBWesbI7ZTrqK8gTO7YSHy1xwljr0ZUmsdB2NbCLL9eu3ny1jmMGkAh+JauDP
I8BYi8nsRkaobVZSSuJuFa0LrkCda73SfsUa8bDYGaD/eghjAmLoa557bWTOOnczsGnbU+gCqlyU
Y+KfoRp7CZy1JFxVTRh4pR+5plv3/MZuMQRxBfGXS3fptlTHsHt08ehAHz+th23L5lcW1fkdDzQe
+AyVC6oEv264Wgn+hDBVpjaz3i+1KjRVTdSH/gPjTUtnAwAfGyemNI2KTGRxZtcoNzDDOdfC5s37
K5hZBrdmctZ3Zx5EHAg2VV24dMYb/RUngA9LlzzOsU1WaLXQU+E/qH1vc270e7FTBAjURnJQ+m3o
7dXlc76XCEYYq/2duJt38C6Dbr3v+kRu0+73Bp8ht53lQLLU55KAM4l7wuT7MpO8RDSoUvm4FV4b
zLwyQmzawaAcyjOdfzqxv+aPUs5k5f5wkhNIno6wdaTJdUiFo7U9+gqDYtEkP581c9IHeAsmD8Ip
eygpLqZffuQ+xjrV4QSCZ1n51uMeNq2sbSwCum6l0ADpOFeMiHoxxmoCO15IaUFGxEO3L8zPwLXe
ulauotWQ5WYsZkh5izCQ0Jp4csvxy2KnvKJhI24Pr3q4+UhjS48PTFonO6DAz9GmYLaK6NSwUB50
unzS+lwncabSbf4BMYgj1VtgGkTAFhuT/ITdUvNpJ+y2lwYRszE/mStQCyG1/OcAM7Yfr0wvPfBn
9PwTGLnX8gEpnBVu6hc8txgTp6FdSwRu2uOM7iI6eMJamqAHiMvc6cyy4yJrvLRHOWFz59cZzxfv
06kCKiZwtRfzIRJp14LyS/Pq80oz4cGVjkbjPCOGy9J84o7BeFGgv/UxxcU4Xofw946edvmitjKt
H/TbIYK0GYFrUDZTsj/fj9yKMa0JAlctAFG4nzMnc26PYV9EPDhHli3mUVSvoK5H7KFxPR+bGf6m
TF1N2mToci5PjvaOBVvFNmCxjI3SuGX++jv18ZTcEVaMmIdYLfiKHPz4qIsasqLkEUitco3qEZEa
GnWtbDCzMkQW5HeA1lK1OcQ4fALbyrOMGo/01UXsPq7oiBjN06GSJhKTehUBlRCMhJQZItIyzh6z
OGQ1M0vTGnODIEi8ZJQ4fQcd36rsoEqJ2ULpys5I3gpmY6Q0nWiY9s5cL0r8TyzY9wJOgh60vZwR
o/3n5Yq9g7kQlMoXblS8P8bM3mCvaXCaTFAVrGZS2ZBIRfvGyHAC5OCtKTpEdE4zC/qG762G61uc
b3qLHcUztahCZhnhX29AyhW3QjLrddWuLNnjJd38GgHcvJw7tQhLdEXjN8BklwRmbmzkrEPMvj2u
ab6MtC+AuQL2OTHJKE5zjxjfQ0ywybwxrk1UvcpiyB17nz4iKgOrkPa+iCVL5+y/U7gUQSPLokgl
m/jgsiEpozMuF57H+/tduXc19UTuB90eTPwjtMh21WBjRLWq/ttLgFe2i8dLhC9JJKOl/DPncczn
TiBCFxYocpe3xdcJhHqnsL71u+VVn1HOdkepsVIeftYIRgOXxp16iIVYRrSctnXRkxpiIOsCl9pn
P3anNiBbgJYM94+1AnS7OhSRdmrl4bwva8MAyhOBgFhJsPQ/Nv/ULffeM2x/GerW8ID+PBX2jxzX
Rww+mBIGDGql5sRa2oHgXedD6jw5RQvaO8wc63PUsm8a/3OQ61QGq9TDyA8+j05EDw1p7KAF/bzH
GA80QldyVYLdGEcYfYQgre4gJT0oglKF5CAxqhz8wcrg4CYw40jdrAUQWOWkRsYqJY/fUqYWtsTd
FLUspzcMoBrPSqIMEUVS0gcymXFwZguCXX/N/LsmgkioQGxhbO6Wj/SEAbcJykZPRDVN557HO/ef
RO5qcCZkuKo+NfpeRV04RpBAWD2cYs7DCwpq9l6vWA8PHiL1BGIRREpeK5q/KkbBLdBWJKB/MOMM
xXnxWTPgZcCH6jfC53BZzZc9SxjkvfQ8Objspuu4DV7DbD6y71GfZeRStLM+Otd60Pz1B9foXGDF
UMTqpn4q8cZz3zvF8eo+sf/qaAjcNk8WYOuznDk56SuM2tnvlsl4NZpO8WcBPHGjjISYqLqCsXb7
MvLkWfXRlWoOXM1tLPaqpKrOA/ZVOGdlsXHtZ3NV8ep6STQh2q7Lu2oyckgAH2Tru1WjhiiZC97G
Rh0y4dHlWiTBicDgyHDRQtmLqlQYlXWtCM8TxUQk+XTrS46efma+teYYRcvdaYSsOMbhvRdZm00c
B2cfyG9qkohABc7VYUp01NbT3E8Nddp57+zc9VbE3FIk3BcUhF0LzWaaiVRxapTPENhjEc7w50HR
xcyEtN7NQ/0wALux0pml1N9f++xDT+8A8kB6TxoKPNRlq7Hkh++8XZElIqSbQsdbK6i7ed5T7qv4
VamWMFLwQwwBDgux/BsJNNUzPBgbOlvFD9tOX4Li1Mcg2Uprbo0sYenYKClJZ15A8RJKiY2KBWtw
p1bmqRnqodpqWoia9XFykyJINtoVgP1L83lsFiIdPdO7PoDDPmx92DPE0OwGAe+42zGJAzJiTwf4
SJwtqjik4OMg2JCjSltTHUynUhiBcwkX/BQl1Cmh4YqfTsNdTMiW3/5UNF+kVw77MKlzsHLumdBA
twlgOYBKZUcfFQQPSYLTFbwuCcp1NlgmFVNWsrHktII3vO5iWQRWHk04AqWMiY3LmMZcoOCnrt0v
8D0cAWb0ZjNP61EEoG84GYVj6zE5JuCNoleC6ri6XgThU2erMubDQoFy+QtsNRKvcDxkNvm6FJOP
TXdIQ3tyCF2P/8ueBNEFKREOiUTkyvuaZwdnkThp9lDfNNOc2OwiPZoQK8M7ZOvvDUSIhrEeyuWU
eisAmrH8CHhIy1KSBCY+2fsyV1t6pRq6/rdgawh4LuYMkf4kTgQLP/43QJocRWRp5FFzdCBB0is9
B85AfWOvKRyo6SC+QA4fYeSrdh/Z3AEw19kg1/A8tTPFQmR7r8RG6ViWzUjTcrscku1T7TUNDgAV
j0Veup6GQQjETQvrXYsYkQtrNmZsGx+L3Iz+w2vX0CGKL/fd1xU2OvSXvbOxzOo5lWJaw81Az+wS
n/T2VxnNHEX7nCWx6Sn73szSqoCEZIk/SIfDHRm6mUSOih2+uqSyXxgIStPOuiMM4Hq+LFNyky7b
ZWKC+ZCGgEBMXHf7xZ3sLRBaVnfEaYfSQnnLkFzaiyEJP9dcxGcFPYu7DV5v2RudaM9P1A6krs81
ZLerKk6WYr+xF28rCY/jMAoFIsF2r/HVeMsWO6ZICYTTsScwJLKaSprSW2HzibDqbY3WjvKZTRXC
I820XzAk4glhZX7Z46t3KWJhkla/wPvDlH7LRd18IPe3lR1FqXwTz423c7KWA4UeiOU24knqCebD
obMw318laxPxtZSiAE1edlHRRmKJLQtKbTCka744Tqd459Qo8vq+NEjyPbOqOe0TdEwJougjTNE6
VU5RE890rsvr2Hejk2VUKktn/Dqz+qIxrHmyQLSw/RJ8GY/GcQ+QfTbM7UN9tdYSpETGrK4IWA4t
hETbvjg61DGj8RZv9tzBb6B285rSYdSDBenudVHcHSPqwEPEM/VPPkEEVqyTcyfOi5BOHA2D+w3F
Bv91YRKHhzJA7rNtHgzU3cgt0tdSAXM3SxNon+I2SIJR6Xffm64eWf4elUlW/Y5ydzuN0fDPZ8aO
m1Y9dqxuDHW+MHFpVVkHiv932sq2ZtTDekXM089KjZsKU31892a+r3mDL96GNSShHRE9UEfs3eUC
L2XE/U+d+PxUgBrZfDo9PVUX9adJyFTICEVtLaxjdFl142gDUyvxSCqX0GbzWVRJntefaRLulHoV
3ZQpnB9jMvbd7AMga/RbXHszllvc7ho+Yr/R77o3shXfWwbqrSrrATrwXxmStdRLnTPZSsXCR13B
VgQLFa2/i7wFY8NnpjgyRrINofy+PHgHPJgvnFtwFFrtWW5Uz8k4vpnAlWzkQdlcLGbD6WSff4M7
uAtDkSrpgk9ejngfzDeqRKF+41fMwP00dpYsfn+udtzZzY/7fqa0zTa6LpjqhtVD+6KXT4KgwDTL
xeyB2ie4p5IhVNvB6c/DLQA70FD6gTvS8EjY1Ll8I2LWo3Z+GJD/DDnc2jqi+oGLaE2wRNZBMSLT
jkw5Rw8jiKMQ9cYxm29RepOFrr51XT0TNASRHrNloSxgsyv64+zmKL4JUfV6RHJMNIuCxmB+1xwV
Qb5f/UTvDRD+4w56sG+/GHvz/OxK+w3x9I/lPdHOoEh7Ja8j8Z5nMgN6RkI+AshvtTn58nby04lJ
+0KEgEnE99eiwsOHZ6PVwyHYBDq8utgpxBDYU5RfYEtcoANpT74qd2Svwv0jbCRaerhcnezt3sYn
WxaMRjwNl/wO8O4Nvhd5o9sYtDMgUAEDz6X/iigP2EXkBTLzoVmUOveZF3LD7e+6pal0i3BY/XR5
UEZ1DcrhDLtBcdjJBq2G2SoqPBlDiaqCG8YW+5tVEhdbrnn+S969H+6HeAqGdaadLMiSIwCk3uOr
UsiEiFRXTsAvwBdk3BYU/NqZ2giLwCuaKv40CyskkuKmMHpWUkaBqtydqRrl/HmwczlAlN+qUrAh
rEHXmseFwPFoy3Uh9h1r3P+S0mSazdscGu+17P2aobDgBWaYNB+yWaPowqm3UoJfdmgtXRzudggf
dGDZr5bSa/Np+bIM6eXcaF2FkBSfXfNcI1G4RHfG5HSsfvA56GQoRcuZ7gygUZ07+Df3sNLINS49
0l6rEdGii//FHw5/YoJaoFDekhkKVH/utYT0E4tRl6v4nna38abO6eZDWZza284Xp/UYqME9/icX
lczeajhXsKdrVY+zyHPM0Y520Ciw4uNuS6UxgrqOCFF1tLQbra/pzuukxo2ceevhbj2Y5UlCxu41
npyDyh+Wzf4DtmVzNFZWj0y8LpKem1creNiirVnABjHvhkN3B534klMqENyBzH8bNPzeRk0bTAQo
quHEHYDQT8GpSN7bNVlK2pyQM7/s9zoFrqZUD5bYMLPRshBGU5NBEDzMU/K50dvGCLG2cbYwsbw4
kgiu7KlsyHRVNAYWKhCl2mip/wGkRO4aKIFShU66P831L7UFGiFkcds7JjNxQJOwzFvkz8PtTs8l
zb1YrrF7WcIt1RKuDmx6TlqSQYGOVBCM/XM2zddJU8NyJ+oH2q1GpfNC0J7Y26nxmOA30esEYPJu
60++kyYGNwWNS7PiHoiUKAodG2AM4mk7gIW5o5Em28OjLTjbh5uaWve21+zLToaV+Gs7rbjT89fY
Hb90/K7k3EckDzfTNtAQLUmHDC4MPIHl1jnSWuxhnx5IAzbVsflC6HLfnfuLDVTCXfwId78bGsPB
1Kf0hNvP7ltTg3IVmoLbYdNpRUzR2RVxmJUBBYMpn3wt+3ia9wVsoumY/Hf3lJ8TfnWQ0q2rMFJf
9i7My3KkCCC+7obFN9Lui+Chd9RjBmvt8CqDH6QweQgB9VUdCpM2OAbJ4/8sH64aCOzd4wvyxZWP
b1nW0EfqXhE6lpmleWs20wBO67NLbqluxd3MU3+9yD8wzcJ30Mg2jTRko9roHw/ZP0Ch9m70OWcx
nhaIed6oi7P6Ye2MNBk80aH7x8DzlpkrCKQhmX9yamicI1Co3BUuvqxG40LFmdD8EV08+jY2LNai
jcfh0+h33YNuZ53OkcuQsC6685g7wvEenr5s5yYAjv8Tlp4PwACnGtLg8GdlvKf/R6hFZOM1ZQZm
ELUM816jjlNQoVUwWZmu/I0JsQ5LsvcHvknatbrYwbyuiU2hmeDowEqxXSonr92Nmd874OXUNnZp
5tmHGDzEV/ZkmSGgJVs4E0BxoKlpPFjIsVgQB7VlLYC2djcFPkQxO53HDePkilSqPjnULMBAVGIc
3PVuWr/zQGmJR+LSC3xJVP77pAs9eM4Y1hHpwLDwJ01EH+Pn/IQ8QsChBZLoz7Yb2gRuY7cvoBnF
ape600cQHjxZKx9tbr30J2FfRgUnyTnWOGxfM70Yaa2TfklAw6ycb9CQ3K4x5XlJwX/j34SN10yV
gCJvN4DkCcmV/wap41w7IWKWA1uZEKzHruA6FTlN1UJhsE+gAG06PB7TRh4o1oe2OxciympBG4yq
WdtxHG6OKeHkmWdsA8UctLpcoSY4CL9hv0UkhXQFlQUcM2JuoDSqfofgCYtsx8NG8by+Zx6Z5LV2
9z3XjTL13tn1A+/v3Z1vHkxodn4LwIGW20V0/x96OAGOleLxkxB3yFtCm2aJAbwXElEnXlPD4Zf1
2njghwz5scxeWikQEQZZ3mdRbr2Kvap/bEN/fNouvVFQeXZTmKuDaKoKsocw0wmd7aX1CMaUjfTN
h7r0S4hBFh39Fl63RcpaG7sMPn1IOUQxnOobHPQDj7PLn/RM2t8nBHj8+j8dSjG2YwEUHSsXTNWu
77JdQmc0KOoizH0cRSZJhyobsCkaXjDzSvUG/tiRYpjC8kxHKYTI3Xifzr2Bb4iVZoy3HGxXYPTr
ZJ49tWQly/Hk0AV2OnZd020eDJBDlnBTUoRS8neGMv2WfGuqb62ZdXLWzhAK4SrPIZbo6XcmFFTV
3J0QCkjVnJcM4Khgjbyv2BPu1KaYsp5TipuH5Ogr3/tNb3X6yfnyJkTjJ4tez+WbsGkrEGJ5+Iat
NmJOohAInYQRxURZ/iHBXDgt8wWhUzSnvp4KiN5FyOYKitEt7c4xeeOw+L1cbkw2AyeU2hHuDj09
+ASuTZs1HASHH7UpC30UG1S2i6vM1e0k3RK0eyAoDP+oloUNZcoAm003EEYRq/atSXs5GgFb6vy/
voSf4i28/tGIY0nSBb/3Pv3tapsaaihs8mADEnnxKaKd4SQfh1rJMeLCJ22Rucf1hJAy2olquEck
OlgYkFhYvL3iF5GPxwnZWHcl/Ffmw/hP7XvIxj3f8n6DGlabYEFFqQsjMfRwynHoyl+GlptQrLaZ
sztfqiRSyT39DMFBLaELlRHsTLud5eMJZ93xZLgPLKzgau5+1tYg33jpFDzfeLrFbHLKQ2GS7uuE
rA5q/dx3mC4B2yY4vBkLanLFz69zHMMOojiELrFe1k3xkOkOWtJ7XfGCe362/oEnpG3mesTKx9Xn
bUtPk9Z9WpizKEP2fVdLzoQonwwzZXmhUhG5cfGRXR5sTWBeSPXwu2zECdGQmV81/+lPDHWPzStJ
BXuhyVnW9ritGh9dBsZ8833m992plH8bm6h3j/E1MLamENVd3XX1y0+/FQvKKhrsBw69ERfuJ6Y+
W4BU5mB4oTGmsz0MJtp/IsfRtGovSEul1PZ4dpU0xoJVnaQ6Ukd4GUDCPVdQ+5jLtvkVAOx5krPp
bpMYYgAbyGvT0A2HmfTa6LK+aRr7OK/qy5AzqZcaePDSyx0RgJPRcnaFmYIyOgzKYsjanV2fcheC
UjKk+KZDFbVpiwBp7Ywqxm8tgXFenLVA3Ti38lUkDzqPMrHY5vjelaqQExnVj3QQ8SFNueqWoz0i
DrSkyTmnJLLIPsr/aGpX9nZClMLfb6zxqLLWuYv1Zl96/HiEgFNR/oNKgjCVGhyCRhhH3xUMTQ+n
pbNzpS+n+9ny8VuLd0Yw4YziZvwOBPm2Wo+taS3wumyzGy32Pa/Yd8EnsWmdw1hh0TpVL4Ga5IUo
u+qOAzndXVF1hKkpt/frm7pnMMvNLJ2gura/vNb8qMjf2Hkl9Xw+kYUXzfaizbnodS2h2qeFEv99
9MucCkXkte6G+E0qoVrgfuFE1UwELxK0kwWdtV1G+x4KQh8p8G0Q0fTL9svy8Rq3C2kC9I3eQvOp
/OYdhdvLwifaW1yglcP0baSkJRpcqvkD6WLYcW/mD1lg4h+QEy8d+iWCCF7Qkord+j/7MATkqY3/
xEmaBUaMU8q6em+3Xw+Zfd/ehiBOAnpCLEi/dMe3x9jTNcnn1WGw+7HfYwtOqOvZLe519prnyCub
LwkHmlZrfptV3GA9RXBkLHc7U18gneqz/ou+KNEOG8SWEGHw+SUbkWJ/MGXNySOibReWt2EebqT9
rMcjnuLBGMBSlY0wy0C3K3QJvHhQVugzr4rX7rVlJDzdy+X+Q4Z7HfCeHzi8ZyYFQhE7Y5kVvrg3
FuhCAsnvn/AUiR6sM90BBSvNy7gq1cZe0HgkNLGKrX5wpy7788IcJTtXoMW3lEOd8SJTbBLiWMYZ
sEMEJPrgMwp63sA1HtdxipDsce9XPXpoqATY2aWFTZZhMLYdGBe4xwh20t1NlsZ9wL2t2uBP6eVK
2UxhVP/b7OIp+iWvY4wNfmBcrhJhpITffZdq2RNatemLBdgwzQjlNFhANlJhCfXRlHPzDT7kStmH
mQ78kvzezgwq5nO5EDxX4Xzcs+Qc3dMWj4lU2u/C+LITYMaV/BhKUrH09Rvj8PssD/VONy//0Afd
eHAwFH/ymWrLtAJwM7wq9mV14osH+XogFJZEYpWGuOpwT5qWzQMbtwq/TOpSsBfBFZF64+0ECxog
4kIQlC33BH53+kOyQXrrkQ3zEGSac6Z9a3ty0/2NAvGWeO7xKQY7pb5Q0JzUY8Jiik5LN3VkeLP1
ug7E460khMpVVbykVJyYt4v0arovBJewd0SppHJoMJjaYI5Cs/e7tIauWo2uxC2DV1NssVxTCP+2
V7+cRm+pHh519r1tfbBBKGlRhXCeASIBs4L+w0oCFSMQbFravi0SlL093cLo5snA7ET+VMru6a8C
ieCu3MgVEgtg1r/gyq4qVVgNx4+UpMLjuTTO1HeLxCephTHRHr+NQ5nuf/hOpQrPR6p8utMTuSV4
8qmEfO7VCOER9AOn1gIO2hhhPPqGL7uuWMK5RyV7aHW23iD1LGx9qJln9Fg4D1Z36Z3pc3u+Ybix
x+T9qgQa094saVKnVb/cRw/CxGycwkd0nGL183EbN/afToF+RBO4pwjSqZvV7oncm8c/oITPPSGW
aC7T3FKlGzCGQSLmCENxPzQuOAD0Diotj5v6UATD7tmqZ6MoVcUItyfCDveFjoRoX1flkCuI5G0v
q/l5CgLrVQwhFrun877lvA1KK4i5YMgc0S9YgGD+t51Oi432w6hMw3GqKywCfp5WI7sbok03gLzT
byk2bnRvVWKzK+C2phGYzrH3V8KDjgWrnwskz10nThrUZfRiPHIXN3Jz9AeTI5K9sBwGn5VJjKHg
MIHNre2GcmvBW8CaNsS9IZnx6xRXGw3D/Pe10XnbelDFdcWyDwbSt3Jl4dTDRcsifbIkgvIYx5TS
Njc+HiT7rH5AIPMoohivdWKd9PhOFoUaJp8owl+rbq6MJPsEgvKq0PfB8CVUxdh04Ai863f5C3ZR
8dJ0rTX3qV3nCi3D7gGTMbrNvT+iu9LsXD0MbgkpC/hDvCq8qb4N9Z+f+ssnRLTZfLKbA/KUycM8
AEorYDyI/6ZdURcNv/K/b5xrrc30Ry1DHjxxiY/hqSh2HY2vfICp55SUR497qadWS/x9xzXFux5o
4omK9SOAlPURpQboubUd0+nmM3tjUKQ65LKb/W9eDoucLZmRnu/u0uhIG8bxR95Ed8NTmM8J1ErF
FjKta/mMiXBAZMgZQhMO+qJ44EmSHBYyu/jq3DZfJqvkqOXHOZ5UggfZeer/eSUp0L5dD2eR0hYb
98qBa8h/4MNABmu6UXewRDRitDN0v+wcbeqvI1BOQ2Yyd5v+6NBKe+GQp1F569Lf9DMQjc/9tkFq
TGyNMVgrbJbFv6k+BrkDkUv7IK/jYy2UIuGu3XdRI2MfnUIXRBhm43MDtEI0O/k0OPr41NBVGSYH
taZBlGllBF0H8BdsyG2kMVBKKjC8nl4aUVedUQEC9e5+e7P78g7SicpZZfFSY5t1u/qeFr3KqnCD
BVMr2pzU99aptnI2KDd3hLuHIprfOh7yqJfUiO48UPaiGrROiRE9otqZF1S5fQr4RVkuJtT3zaHc
jkGyFqt+MzG5giFyyw8GfkxPhiwcESliWxPOi0lDVPojgEt95qKROmznfZMEDRXeB5/W5NxBnrju
9t4QVMxkioLyiuQiNwNK5KFHhfZJR+nzLMoNDyo+jXKidb4DN4s+C00KEBnHc6HR0MZunRyiqF37
qzZ64lo5Rlo9x/iVswLsEcQgVhNgOVvdMJ3X03bj+EuQAdiCWPu+9y5+nHqEGRkXjmb68QKR5Xwn
REFa4rX6p+RCat0tth6HpCDI28b0kacvUfo4utssFhqf/7FUhQwR27TlXbfrCtZAnPjVhgxK3IXf
0Q10auUu49rKD918O7qGdKVHAwyAyQLm2LEglKw/f6wwX9LHNjYPbNW+SGpA57+9/TkUMEFB2Rut
jfZ+NvQq8CMVLu4qG7sihW9dUeGmgbIXiye+zAAhMakBHsnuHWcRfAvH+S3mx0No5AGXDlaljFTE
zW8TqDnFLuPrQf52/2hilode/UO05Tp6gjF3TOf2hy0nb8AmmgSBIGi1ZOuoeHIKSuvbrSXpJSdD
zAoGA+njPryAyY17FhfN8+PyCYuWzpCNTYMo4rb38NFd3yu87JdaBtWGgUPi41Oe3TivGubQXN8N
tc2UJ/91Fuchjb7HjPLgIxF6W7+1aQbRgKSI19GMwnrm1Enc8/p9xK/veTMBEWTYzV3sHoZ82xRg
bOycVi9hYqPAIliSA0TQbk2aBAhedJaQ6rF1FsSp+Yq5XQV/Zab/rbZbitJAR20Xp0e5ZOWdyFco
5ItSGvYsxied5fT6kNnocmUbTHLDIjih9i1AFDV1V3bi91HQ1E7PKjk395sGTl+gwdaQn0QH+ZQH
972D8epzkudU2BsIs7nWr0gqzNyk7D9d3NE3Bbq414msZLqpElk//i1fzp5/qRhISDlyLg2rIyyZ
cFRv4BVMOl7iOzavB1dEIFMGGbDInXRx7tlF5V/cEl87qoJpof09z+Sw0q69vRbgXghFWc5Y2gwk
tLpobdKrdhT03q1FXnf7eUEHnNUB9t+Ao+GaQuX9KRMzQIVdZaZLdGXolvM3yB3Be/O5Ycp99qoc
4MFFF47bluoN1ID85LxVYKT1cipHoPNmk1bJv8mAzqvvd4kYk4Lcaorq9T1wN8cjzSWk/mYV2XNE
jZuwRWuIw8t9DnCnZzMiDZLBa1SpyS2m6HtPu33X+ARlhuMssCMM9oj7H0jY2QJ2NGZWRWYMVNVX
oEVzBBahU10IV9FVc/g5N6nkGEfGGk9AbDfyoxJUC8UStnkBhLDu4fh5DiGcXzteFccieJiPKhCD
OPIVSBRkFqfwTZHN6+8tCY/bWw/y1CTgVCBZgO1MkJFobjnmMyKb/y2uuD8sSoHASOd6Y52ikrsu
fuMVdlf70hgbHZLVz/0daTwOEayq6PkeDZxwu/IPx3V2ciauFkjvCrGEQTLLK1rXopJcph64iBHh
oYn8/NQLWCajb55x7ar4AFi45PmW+sBFOT3myoA5OQ9m9QMkjl8kDNIKem8OCHbvvSmgrscPWaHx
eszsUIvhZnfP35CqN9RneHrgT7/PSleErivLCLd1pANc7bXvgatvXrFqWoeSwOibvDaZo9ZdkUXs
q6Q/R+4a+Axk9BQBZgh0aaFWaXX9Vo29o3ElVOO14/46YLyoc1f0j9N3dgIwOdi1zCL4eR7gkSfj
2uL7J2g3Fx04H3TbHbsDlvRTl68OBr7TutC9W1w+oHluNkvmJSa4DmGOroA8hvFD2v4OGmdDrNye
V3LoPTNua8EuQ+zPr1wLdDk4Bm2wlUQEJPjdhRJBWOfmT2yXYOuHtlQFXk/VfDiZIpHhSRKHjzLc
ZOJM03y8KXV0PkEONOSRkgSMIAUJYp47XGHSy6J80uaamJFSamldxSiuZtzl7Ecvd2qvUbsWddA/
YixKd8BonN5karw4Ojn56F5hsHE3MTZoRCEJgRtDZc5VMgoMEzN5YuhbB2fWSSro0nKtr+Wzwg0R
xFmkh1DXBJyoB4pApH2QnRet0DznjDuHP9zhbme6GiKN6op7OHFaxT1uj29z6AcP5OhurXX50XKf
75XXZW6lgkIMUXlBi5wBw8ULjy70JLGmrrbCjsKSOIyH+1/rEWdZjB5PLtD3T4vwEWeHgvS5qB4c
OPJbOA7533aPBvm3C+DZRXfnQoZvGstPcrMXm9JrePz4fT87deNopKZpSyFFib8WMLWRwW5K7Fxd
YtEArjUlNuVTm4hKhoboM9wgWt924Onw+B7HIuiQ50+SdrjJ9cFeOyxcC37X1L56rNxC9uBQHHfu
cbmRcIWQ+hNmjmklOOucJPpKlL7fWQGLdH7pAlKj00vlsKbZPnuPl912r5VrfUca9aHZEKQhRkfR
ot9HfycEQbuirJM53hYgcl0urs5sEf76M3tuBwgVP5kqC10bTlnv2iYJcnJnWW6oxXpLbrJtbXqe
6KIFMb6b3mhdU4mgPVrrI0X72O8+f3sGRFag3CWyowDBvw19uwJROhwBQ+ha/JEWHpyTggGfJRVg
4I2gB2Xfqi6ucC+ufBKV8ARhafk+FqFO22tO67P3O+WL4nAaVxP/FnPgi5AmrnYJ5sRKC9/BZTGW
OmYYtQe4tGiY0/78cRuEHcDS4Pzmh+j29Aw21UlsgwHKq+3w0GccqfRPS8RYr2AvC2K3Xw1Bh9iK
gwDQZZ3FRUUx7SYyxYsumYP2hG+sV2Bv8GaXYCX2DpZQFTF802nOGr4LZOXHDFYX3mzZcutDE8ek
KZ4JX1aVGV81MA3yejDI2VemTl2kV7LSfyfH1DBIt6faSjV0gU/kvyvQS+mq4q3uuVI1nPBhMHNR
I2HG3vxN6A3uJQHdGazceyBRhUsURW9b6pH6Iqmmh/vZh/L5X/PDVmFOwpbqm8JKBO1T/DjFnpc6
/KCMhXJDa3oXhOO8M1O9Zi94ED4sk48smaL8VsKxnhY9j987aDZL+Ls4FFvkfVCSzE1j5Jdpf42i
ui9VcYcSnq8qdbL6zJSeW70qB4UNpJHbeI1z/yT2xuhtB63YrlhoDAUBDVhMbJsImufdADqhL6bJ
g1kk5xnWb/4G9cviYdSkfx9g/4xRwGq2V8y3OphcsewnSe4jAgcoZnjsUtoe1BTBLofLPsBoYD7W
+sgwO4Qb0Cltf6XSVKrK7yO3/c3QUL1UEzi2p6Zpd52I4QyPRIOmAR5Gax568RcdeX2pnTh0do59
LVGAXtkCOe9KlE0wGAhYRYcnJobDBEO6MNPvSfrq+pICI8zU49SFI2DIHpPV4tbZ0RpyiG0ZzrXf
ubZsYfq/Zw0KwarPIoN2gURG8DlbcFim2uuLYaGChpLGVSeNx7z2Y5lJg2O8Ldc8BJXDIDeJ7CLw
fBI1lChr+tUIedlFApdObxBlVI8frmgS3iqDcjYlAKwmo+f+ciys171kozwdbRCgE2wfQwBIK0R3
kpwjT2fMVj6UxcuWhYLQ7cwkEpWmJDP9dpUGQbgX3U3JGwj5ZhzTfQ9UQWRYen6t+0eyOTFvAjfo
5Kl4S06c6rJLQO+seH5Ihk/pr+KKVQeivqFcX44FB8vU7hl0oDaNSJoUFlX9qdeQC5kJV6LpTUQh
IGgcQHD/dtVXUNs7PzbFStAsXLi4F4i+5SuAwJfZfXd+3Wl6SX/DmQN8b/BVihXk8Blx+niPFnWx
Vl2qjwqhDBITd2f2GDm2LURxp7Cpiw1o3xCkMq99J1/wcDvGzgnKFihdm4dA/j6ODthjhkaKT6wk
/dhSGHQqdtd1zii5mTl6gXRWgC14b/4tVyRPm1s12Ce8P7oxA2wHjatf7GvxRh/C1/2Q3vI8eUYp
jTNZNM8lLl2O+z3/VmFMsqb7HfX/6irui8kr8QSDDIobH0bQKicccXbbdr9yduehyCVuhjqYZry3
cGgNJKHXzQahUae7RMNhXaaBAZOtPdIN3RoriBN+DP0IeNAzArsm0KMrprpuyFxQZF3l4NLuEdZ6
P0yy/1x1lQNzxHkn27+AYPRXRTYYR0iJdcPDXYoz4MBoI8M0hNkFT0LI9abVKT8iD6MMGQUgoyAT
jUwkAJ/OHWK4agciRMB9olqQ/cDsurZc1Wy7WQt739EVTqz9X5+KJDfr2BgshOPFXisQdJ1tW31d
NAUdIOLv4SYkzxNzgChiTtqPnZV5JSGEbGaQMdL+4fzRd2/stDF1stsQxIe70EKOs7ktqo02DikY
jAM0Zpm7JUueuFKsHffGsHSjE5ve+OZlEbmvzMhMVXXbcGBIYmybbbTZLV++ezcYLjP6KdYn38eH
UiszisheSp8bvexAQEqvzmSPWJfjS2nFysUmywGsElgNwF61MfPar3/csxNFnwH2mtoLf77Q7xBJ
5iN4OhbbLUtAAMaMt2ptCUcb4BsmrIvPb/eJyUFsmY9U08yJz6vsf8TSspH+KmYN32tKV2Bw5af+
2HsXMmEbi5zhYf1/CkiYS7eoc5U1lh3EKqTtNARzxsRYPlH+wSrW6AO0k6QaD0WYyPP48rMLGfXP
Fa6vvGzm7MjFe08ktEKY8MINZTUH0jOBbKW+GF7ktFa/hRrddn3pgc1Pn1H1hrC3D+zR1hckuyfc
NIBq3PwN7/QqlQaRG1ns7Im7iAJvRSwnM2ZtB9j87LokgQB9PQfWpe7+U8wSet5+Q750Asho5Q3c
G790P4+UARdsSxTWuY8J80OZ/R0t2RuH1zAcpZsU3M1RO6REqX01pyWC/Nr4g9+OGJY4hmIdWmqT
KrIrWPsrSxLQHZegk6bp8RM+ZmKJ0PC4ei/78nGJr8oAFMsv/QPpaiC6GXcFj4dAi8w+nuY74xNR
OCGQuaNQj8Pi7DF3TbTqBwP1K8syVMIqJvdIlgsmC2f031SqApyC25RDV0DRnuU47ei2C23Assv5
FD0tm4gQY/ChpHg62UxWPgE0IH4kecwm37b7OC/5yIyB4cIzlrb4nGnRMhh+zLfFkEuUZil+GadG
wUyR5aY/ZWdZJwK4gcqfum9shTvSqGeZAE8k2kB/sx0R49iShEU95o2+PgexxlsPBumaOdO8WwkI
DD2c2aoq/ifxA1rVB8tRsLJWmRQ10CxG1XcIef4XVEKMq7IVruM8twUCZ3CaS2Zfi1Eq5w0tN8bx
miPJ7MzKkjGsNarzjVBj1tfQRL7vLzvnQw3Q14zPU1XJrDU9e/lV/fYBEY3zRLwM8NgDL0db69wC
bx25WMQdsxJYdAkAXYha+qIat3ldFcB+nBC5ta1Xc2nW0Q7G/hsf9suqkLN3xd2nqZqh4pd2AIQf
VmOVH/GVApsychmBYTDkMZujANh+8IOPI4ghiV62gC2PIrpNlmKGDGkHA96/pYx1mY6MdedIvyGQ
YE9vkqem/SJnpI7uAlydHYjg6pLeNigLDawzLctbsX3qIR1Wi6/68PoBcE+S/ehKDtgQBbobe8aF
kWGGSZDtacsfg5uLeYg13LaV6iOKPI3PTdU5iA8x4xnY+6bTi523nCrgGxeUg39A0F2pEOcVm7CY
fX4GTxPc5S6W5OiZ6XqggJfvdk4vkt82KQ0sDlVMzSlDuSMCEwMltSwGZl52t0AQNdWJ36fHDxmz
87RAfngiDnis+mxgeYTN0Ex41O5r+DUH7D6PcS4UnSTeP38euxDpYKS3+KGsy8Tzcq6itkGDgRdy
5rhjJ28xzbvqLATPQGnwX1sB3YgdkbqBKoNXLSfjs/YIn+kbffAvoTOstioftLaH+MtPOy7m0JrH
p9iSShyCOzoFdzvZ5rUhX2B0IBbZ6S7qvAKZxmHqWO6RALfMYLrXpd/fzgIsLurpoDQgfOhboImy
S/w5VPLTmHi2iR9uYQM2ihd3j0xypQDeJTjW6f8H2gsDm1YYNEpdQQhsNy+Fo4KmpqpB1oLpy3DF
B7cjRH5z4EnzlAxIA01B0n8K8uXhKeEabGMPKL1DTBz3kchweKMX3rKMEfAxlaIgMn25tX1bHY42
j8DdGiXG1ixRGjTLlsqHRRZ22UzBMUbksf/2eXxi85zWpcRzkaS05sKKqz1ULhmwTgXhLfPJ0JJE
mn9XNVcBRs1qRfF3Ss6ByEYIYyHwfZx01ubni077rNVkwEYi/i/3SAJRPCSlCePhlgL9WdppGqtY
4/5S5h7Y5GeHJxnUqIQmvGNA5FqMRJAlZ990Rhm1tqhCvO7X/ImPMRZpxlIZAuDaaETCQxyQg4li
zBMuff8qLdDsCi2GPzjhpiVz5e0ybRF7MAfDbohSry/aC0lYakr4gKvCr5UdJFGKgyVZv5YvvbpU
rI5e+BC4q0p5d7AJYIB71n1ipHC9hT+4H5/i00hyVI2ZM6oRoKZljzMzr1SUNoUijuNKVbLoLLcZ
x0KGiUOp9QnvsNd27GrYLl4k5vCQRQBkvyfeplvE8oxWF6zdZVNEfjBOxrEgRGBhs8IITp4fmINW
WqY/ZRTqAoAhz0Q+NLPzMW05vJyAiBPGxz0l7ljKAO6HVIh8KzvV9itvzyv9F9srsjcdgM6y+NkP
guF0KP1ON03zrD8D4CBwKik3oi302aRV/c/0b31UQtcSD9QtCkQbE1zRZ69s583iKRgI1GJbcxsA
bp5Jp4jf77LuqF1r9sZddsddjoIb1Uoa+IOM3Lwo3TCrtXHRKr7TFkb1Ty1v7P/ZE6yU2ztJjclC
95zPu36fubFH1saPIB6nyXvQGHI9DNHXttE0btrpiccbTGy5GyJbRE3vIhqm1jClJRuHrR+GUoD2
7/qkgJY/qwfk+KMmoy1C8wQ/Y9rud3tun0EEdjIPiCFRb1htO6IMzhR5NQ/Eq70q5TVMAp+v7q0S
SaAnKEOE5NnL9AWshD8WeZQVgFbKrHjNjdxQv4SoNPTGPFOX0S/rYWSrW2oGpt6yhLKYv61m8Ebn
ZbRbQRUufbLmws9ra9QyRMVGQF+eWBpwbcuKaSX31TgTUGgwC/NYxKYS7wq90jH+hTSMo7ycquzt
taXZ48A3qLt6VwUAp6f9+c+oziTStgauaeLEY7qWc7MOKk74l7eA+X47YMIysqEVQbvBkOmTn8h4
wAhcSNGEpFuY7N+WMuT5JwLFJE6OOQ2i9q/W5r+tF6PzuTrj/u1K2wEF3/usYN1vJDswEfSNNnjg
GcmCQ+dTU/QHjx0ich2qKSIEZ5QM8/kkaNPhdAaAvjrivRsFoadei7VinLlZMdxQd3A4ebGhACFE
0rSCXt1djxIR6NdJ2vnuyJwa4+BV2l12ujblNjNRyF1EF30v63/QRe2Fr2zj2vU0zqNxfIdR9E/J
yzWZb7xX6MnTVmxsWdtLI+s41+VAAB/4M1XYORlZ5BG5rbFjKX3ptSGoYRRem1TNpddO9d+BHjKq
xJDWmlhnERaix2OoIHRGcuhF9iH+sme2yGy3Tf2a1EVa5SAoq95A073D/bbjmBD8QwjM1nciolSb
Mehst3T0MguD6sPs0/hw/0HMDGOan305w9jjnlF33tFQ0A1BL4DRJ88rLMzT9vV9KT0qCmh2HHwe
2ffBUuyNRpsEgkLQv+j3Uzw1TNL2oFjO3nMekFguACakfjsfIYbvLqZeQNRvtXMBUNm6yWE4JYCK
JvXYXtlcWA3dcZdPI4aTSfc3XWDb++L0KkzklK/itlnSe+KIlvO4fUKs8GOvgApVMixJYNu1g8KH
4y0irvotgiL9EpdRPcDGWKSAQi4Qrz53xDaEt8zQnU4xtYprJFvwAQ8xm3e7u7mRt3UdSehVDRj/
8cFdhM2yU6notl1pRRCh8MhlSCjms1n1VRyomWJn2az+kr4KT6T+nckq+lp0aBlScR+mxxYBbWHt
LYdAkr0ix8iRtBhkvEn8zF7iJJsezIG/hMsRxq/JMvE/DCF+X8r4NALJb7gAhO3chbAcdbkdOk6Q
Kdu0Ln0B75bI9tkS1nrdk4f8VDQ5PVBQgld6eoD26fNDqcdMb5WGFit/7DRxfrz2Ll7AsZgLiPEO
d+OVH8i3+9gUQ517AL7ca6UdG+BrFKk6U0Bq+RrhypQoLPQ2nqsh6py2cAVwnnK+UuBO/YpAkgX1
PUCDaUEKiPJdDBCs57AOVryVxHmasHNB7fP14fhwp/i87V+Z1ETBwbXuK8qk7NUGXODkJtOBaQD+
oLzOeRmvRroRyw0m17rjhaygZBbvwx4MJdbjFl68ty6krsPISIqyFya+iwS7W+UrI6tM83qNMzf7
WVFsYg5LvXcHHZfE/3krwKxYrMDYG5SyUj87FQdt3fpIfBkRDAwfJYMhbsIl/1qSLbRgnRkEoJWY
FmSWqiXP6jfQLMA1eyVFEsNgaG0P7GrcV0i8v8sBmP4Di+vSWhIELfoNmL30XWqDv+cOu0ylE+Eh
rC7EBLf9vAQ7CRu9hFGY4cxuptiKlgUBeWZJdXaA45dHxZqjk/Cg7brQYP5pF7gNOYk+C44cI7vQ
kV69dXHmHG8TRaqxo7ve89wKosqXcnaGPE5unEJtv6YoPs084DuRFMGI8F8wZx5ZlPsJzYg2Ll0l
cyEMOgbi7WGqrTh4YWvqP5h5hjj5gDLZpCbs3dWF7TaNw1lF9ZifGH9QOUXDqcdLlRwa6wMOVVfa
h90hODrwtt4QSDOQZqf8iIzh3foIlw9QG2gTxUjNpmLLuUqsGLapLLgqjqj4X0Oe42hQf7mTRzdv
j+JEmnyd7+d09Sxs4ewPW3cNow0sW0Uzr6a2n26oFxDZ3q2VZ6dX2kRT4TXD+Ne7NWaSYpui5BD2
oC2z1yV6QcXs3Y9k64efW2YZ2T2xyyNOvYURU9FIYV+VtJ9Xf8AEakQLYWWPAcr9GZcIQOShI9Eg
KEYfjeK0vz9KXeF6i+60RsrdRUDQ3yG2vygDy2KKPW8FFEES26Am/lMCDrQgrzfYNI3jDoPQWBWf
n3L+OK2CGH7zVOyS/QlG0sKVL/x19sCnXzgpKqJrrUCdip0LIv6qVK8TuMCHTrKCujInsVJwq9GC
IfhresGxHHZAQ0eSsaYKTjYkAntccIAF8GLLN8H/+ovjA+yfuO4vMkykDxtQEANizjrlnMTVtUjU
qy09AXB+AFfSjj8nboRQGY3httS37ZIto7JTv2CokXxBdyBH8j5/wPI+PIXyK/odiVn8YbyDhl5X
vlN/yARXXHJWDyQM5LIq6Ql+Zp/crNWB8Gj03s/+yMrZjtjEbgUQUJBZwXCHcoqfxLXNhRWYcR90
wbtQ7ua00+nxHyVbtsfG6vmnZTZbmy0VqvI0bZJA3jGAF7VRN3NXNm0PJXk9+5diygrt9aCTKu3U
wpSmkJEaFjeLyyiID/+PuqCOnzDJZ/kDaccorEwU07SqrZUGY41vZwkzscFzWAxZbF9KWG4nmk+2
bNVm1Ode3qExGYRv4uLdxu11DF23U1qYgUi5BcfRmFKpwMuLHOKclZf9hn8wbH8N1T7EyiypGZY9
YKRF2kKpfWMe/EDsEIx4r7JLog7OvTY0x+9Wpjfbefivdo/ndGoQDgaW1S90CrT4NkXdDHhOE4i+
8RCohQ1sD3iZ4ev0DsQbomcdAk7AIeD+h9TjM8PPXIhnbwsYAWP+RLSgH2rCqeeH/o/NWweZupK/
Wu3QYIIY3h2XNgtBPWXu8cGNBMFo+cjpEmTYYiBYD6A3kun+JwDfV7Yzo8RWlGura2uvMiUDvNb9
Mf6u0H1BQ1poJexYQX9YGyFT05eO/Esqp5t47juLQdxFEq7SOBwYJLiL6asx6EKI3GE29Qy1SKQo
cd3rKgvT7fQG1zxUhuOhJIhSV68v2dlnEOc/W8rz22502vagnZaRIgi775AZbZy3Jjpqjl7Wge/Y
2KG0TRaHXPG/EpLqM0T6nsG3x5ueBazuS8J0ZSh4M4xcg3sv6QRUUUkw+OhOV3uqDbaHeU5nfs+d
OQutKjS2M5hVJH2KKLXzJDLT+Ctj2NAgcetIprV9IoD9fXYCBDks3wp503H0cXGJRxnKFVKucAgb
M9EZYV2jRRQ/viUO/1MElq0R5ewDfPh86X+jr6NVMwuCj0cnBAJJVo1Ldxw+FvV82p2XPcjmPVQQ
YBrhlavLmRFJ08xXQq2ZtVK0Z6qzGHjOYd5wtSGoH3gzFwPaMPBbRuNxXx5dZtXL/eHpf4tf59L3
arCSHEVTiDrwUiLhoepUKd3FkYxkyW+QCVHyzsuLxUcgZ4mVRLna9KgFLj0iQ9mT9GHomlyiiJXw
Ni4FByHlkeHzhRLWT3pPUGPMMcwYwHah6LBp7WYlke35jPcbICnNs0p0m5FCrYM/JpQGaQx1QwD5
g3z05BeDSdNUaAnR7K3puJaRHOIYWrqp1UKiKHtvs3eRCp14COuwNvV1jSFp4ZYbrbnQv6rlW1Th
sr5R7Y/ZwBtxdAbZm+bLS/y0M4M1xdUsIugvibaot27Qh2wV1TwkYSXk5W65NbQuRmp+cJQI5gOD
L2KTyA0AI5bhIIeU4j9gukztigN8Hq5Vby9hTBgB9boA3M6rNMrSlsKPy5iFa0VJGJAQbXYjE8qe
T/yZxIQ0FwhJ5dS53YJdEbn/mFx3H8so9wzPJQuNF5wmaclZauUECT07F3gyerbtLr3EPXnleeC7
pRcaUaVAJL25QxyV4VjDH7JVPIEv4hnuiMgTQ2xir1IIIAFyFNShpNrFbdGfL7xaKP6oafgiOVV8
DZjy0XTNS79I3k58BjiBFkA2Z4k6Mrv2fxwI4cvBmJ9145Xk7GtjCZkzia4vAvYnUIWodj/RnWCg
8z7BSatYPJP5ACgMPpgzhLAf+ROfrQHEjqyx3yN9KMY3vgnZoot5HRlZkx1HRdar8RQsJYfSxUwR
T7hTSu+eeCrsQuJknesPxV/01ET1/6857NeyGaxKl2xuWjNlwt/ho3+nyLJ67R4xSfSCbcFmskQ2
IZGPTBNnj4/iaHardSHg7iQEWFSsfX1XCuaMziXvZ+1aDopM2NIDPtpBsjbq68TNtJYBwjfnD6bj
yu1ENwK6dIpP7SpGkOj14m03C/jb5lg1EnFMUDt+GDcc/gGp3wZnT78WXlGdfJFiZhY7psY+wGyd
+fxPPniMoU16Yx4EjbaBUiB4Ywz1Qgnp/K9nQ9KHUrAEv+xyvoe6Bxnoz/UQ1Ki6XQWj0Yu1fa2t
Bo+zGQvVGGj18rnizQ1TzQjPmqG03j9HwjciSft7Tqroeo3M4B1ijVE8lxjUhnaf8ahyxsZiq7Cd
ZloGh4COQPvDExBAh9myhXpu5zcI4q1cY7AFlLt3+BQ+LrE9rrkLJnRRqVZVGG5c6sYiz/c3Gh+O
Wh5bbKsfd4ggNAMgm9+CnVe9U2U3u9j7hBTb2uWwqYTUfjvHzPmas8gus2NK71CGwko9DqKwMLDu
5EiUEC3tutoip6WsWB6VXVjLcjQ2ou0LWxN5kumUGohlUZlKJjgIggPKac765ffk/y/zbrdb+idg
868dDqfH9X03xKavXxIv/xPsJB13RHJUZpYCwdZNB+BY6H637Ll5Z//uo+SI1+JG1g3EgNDRxYHK
WLgnlEVJrnS3OHZ1Tsy5W1nWnw1vMsGdw961IqmUyun1Wazvzuvt9NoafBvHSfrQbsk9ZyO4fi+6
AR7M/IGgPaEjudZU9vb7mJhX8mXlcZFVuQpCxp7gQxuGGtzy11hVg9Sp27vVd7SpdVuc0CbtF3ju
+gnbLdWpW4sLALRr+XKHFQjdT5Q0psDV00UBzDN8W4UQ6IpH2t2w2kL6vYiUFNhndaCy45Yt3JXW
WAcK54GoQjJPxHXlPQ01d+lQPA5Z1p+ua5AvGERc8CmsDqK4w2j5ZxwzqVm5aeBN0WhvO+bYkMC+
YalHc0wPWJ1EHjTxO5JhawH4RxbJDj4EYkwzf6GWkG4VhWq1PtZJ6cjMBG6Gp/wx3FoMJpvObkCx
/CtKMN2UL3L5iVXBae+jXdReTpTusufKR14V4Xwk6Nm376bywYl1/6yxFXWXAKxpsVKSRNJXkCoc
NDCozyzBaCQH76szAZdXi0m+FDxaQEJPHy9dKMrPo2kNyfF+7TofJnG8LNiOGVmc6hRouz/omuv8
0b/PzYROkCcDTlJkkdEG94GkCuXTZx+HBi9kykeQr1Rn3oNUkLQNlelXvjIVbkUuYIf9j2ICGNTm
RFLWhyWYJMmAkerAygwneQfAHjh2/+HFAa3AkBn6RXJJ7bUNE52DUxW8wwH/jYCB2F9L5ObnUj8T
eVRjgkwBoqKvJl/wdG0mLeWlwy0fyOUCzCzYMXpUdmBFqePtkRou4i/eGR/hnqasXuVdvZbssVO4
CjzRzW1CZws28uWpff6goU5Qu96iYa8syEkNOc4A8WdWkB7AFbUsO6xdFd7JfJMsSh6zmUbfal6t
TVrzUpfwWPqUgb2nRBj93Ix9f9xnfcXiUtygPmQe7j28IdM97A/pteWwk/x5py7v3fSAKEJEma89
Kh5wYwe9u99kBb4t4kdEJvB8bE80sTsAaScEZ3mog/RverbKGlmhybVXQEvQFJZzcd6pWwjJWfb+
wW1Qmw8j0xR1fl/Ybt/Aws/sSSOVLzbPRHIvHJGMR/ngkPHu2D4KGnEjiL5OO0A7LNwe8cdmeNL0
nDKVjo2lj5965+Mg6akOM4VpD+nF6ptc0nSwIG1ZwYmlyL8n+PEj+1QbglkewldfLvfWxRacwkm3
s/hVVKWtPNDM6zf3UJZbBv4bS6FtZqTzVtOyTFD1Rl0cD9JPFzkuENF7gu2If5iGzO2lnV2KLtJh
ng95WSIq1HNe+dm2/Rqmr+j5B9FmlX2p9L8S3CROoF8Mc0GyNB6ajLnSQQw9vSGrR7Nppmk3yFw0
4AAC1Cq5yOQZR81f2fEHyAsfyD6Etgd1Z+r94k1Xwc/jTrjyqyUHX1gyG/MWcfbIuyh0M9YalroJ
GGV0EnKUbBDUGnucdNLdDIPbipXgbMfaIwmn2YK33u0Ba6TunFmG6T9pEJ1we/DY98e2R//rVzP2
gxhmpfF4qycDtIGy35mDGqqZoNGvxjop4RP428bMAnFHmZvMQfU4/AZa92Zl04eZtG066wRVCnOB
rnzwrJvuQ6njApVaA9okvrVWNI5N44KAUJqyEukqAdkmQ8uIEsVAf2OX0ob2DsQjbQgqw31NqA/o
40hRCFHq045QzqCDCdBIwN2zaLJuym7KBbVXRyzjtc0othUuMBdq93SfahNRmK1/0z7BbRGmL4bx
RkAEKXBZf7OfReAAOT31Vlls6sXStxgjdyglnBrAcuugy5dHr4YIbhhMJyJr5ObZ1STGgD24SoLu
DYlFbsniiF9qbulKTBG1MLCLLVRFw5brpAGalx66Exukv7OHxhYbOPB0f4DgiDtfsd72j20BVcvi
rnHr/140L90MX5Oih+oaS4o3IpPvpm8tgP9mg6BxrxhowuugSuoeSV1y6DGeWoUdmJftlV6csE8K
bvMCZdHXPEIyxyp0jD1bMJwXsSSk1YVCkoZP9MrTuEmE0cXVXz49jM1LE48IFXZ/6Q7jDhrLYEhu
FKDAkqT7usEMSTp5sIeaZDgfYICHCdBNUKSqTPqeGyV9eb3NTEH1cx8qsrLDgEoJTU+BqwYUohH0
WsnILv5tmFRpffQqbfY2+avTyl52AEzR4qsgompfkHoZ28k7TvJ8cheIY9dgDOAiKqiTACHV4Bfa
BS2IjgoXY0GNd9Hkrid3lnrUb0AheS9iN5ooTta1SAVmzf7cIU4Q7OL+JJtz/SjEnifUWR1ujXwI
JzsMKevUdkevA6DBbdkz++s+t6hc+x8I0yhj5NrPsJIj68mm3A5WXldoeO3tS508S/A8AsMsVbex
HVuK2aoHVUe4s777SoSolyDL3FkINBhC4PZC+/f5gYzjiogpYgfT+mt9P9BJvHAtHgu+P+Qgz6sO
PIVgxG5ifVQtJAtdo5qwN525dCm8o1pGgUY1bmfK8+U6xoCdqnfASAMVthD7+RoCjykRrr6K6Al1
bxqYtzm9inGLPDAChGm0ShCTJUxS7+2xNP6aForKVlWxIGCkr1vCq1oV1QBYdfk/sdpQfFSFukMA
FGrKejWS5DfXsiQLsdspv9n/ONgnnT5MWx99oZyenSVSyM7DIWEwOhl1Wf74MpdURfnHfVwn0dZj
28LGx+VYbmilb37SkfR5gBJCT+Yr8vG+LsCiJn+u3/DqcJjRRbf9evXNVh7b2o32b2RkMWIPA0Ur
w4SN5itYnibGYQwq16JlcpGzmJ7RCsTe3VHILmKIkfpPgIhzAeoXYZp3U5QE2Vdk4M6POs/eAeEp
DpX9qiKHVEivmTvu0thNcNYZJ70V7N6Lr8uq53p8+Y0m/7pmPNPXc2lm/ImUhz81FeRIFOdh3osp
JWX1JCpj/I7s4WxOw+7LgdyYYXSvi4PSz77EqI6lqvgF4Unc8ZPEDn0PJCf5eMTaMm6UEN3K0yeA
tG3k9UoDTatY9BMdBPJ6dj++XyKurj53BwueZsU6DbzvURkspu+yv3yeOoPOIst+L3SEFH/tgJkF
cJH+vNOKe2k+ZHD7Y4b+xAYuZhsD8m/mOpWEE3qPZBWSBtMNynySHtRDYMp6hq7Sbu/65ZzuvOjk
3/6rBO/demBneSJqTIR7QfyAcMOE4/X4pVtU35eOfnM7TIoN4iEhSOS0CEz02cTPsOAESEiDcZYn
P8o1XQnTzWZLv+nZwiagf3DFrTHSb6uyinrr3/+RFvacv91k0BlYb+0aboXT1Q3LYG/fK0DFHyzH
BG/eDDwXudkNB7Uq6rJnGg162t4QZgqr5bqfghjjduPpNEOHrDbUB02NXHgx0QU47Du6LAoFz2+k
4RA/+/tD50hdSzUTK/RWppQweLD3A33kA9xKCC3ysKrVNH2/JvNU56XK010sUowr4suPdB/hYy+7
S52vfkckezxChxC8QIoPaoy0DwuAIdG/ZbpsWZj1qJ3HEm+UiNO+3bMfqwOTLX5NxbUdVgWq0GpS
pJWpzAgHiYqiLqd5DuOIbNMV2bWLrYocn9+rzOmaf4pZyJQuf+FOCdbZ3BnkISfmwb27V3Df6bTe
dw7QNDtaa41vlW948P4WhuKYPIBf6Dp4hhipjlW0WKSieu8MhCIASLzE/Gpf9zUKH7VwFuor3lPn
0lDLuAbLCRpTzyhOqNMO4npMANcYAAnR3NP/ZY4S4Dv850qoNhqDgecYGc9fE1SoH8/DvKvgeWvP
UEkALji5ylxtsDRiKMtKUTsAb33L7veu4QlYEtY/l42cN4fwT8LIuLQnQ7Ah4iUa/R02xU79DTz6
d/YESVak7K8fsipBZO6gfLeks2I2JZmrFcuXksfldPMoWSqascGXlvIMucymh2Oq1blXOCGqNEI8
FQRnObHYyCuIahEZs1Dpwk90FyyIS9/ouoHd/VBuOVSuEBPdgcvQScwi8Sk8moawUH/+mtTBvWO/
xnDi9sZTOtNTffLqce23PNwqbaYytkNEpuukXK2r05WU1BG9WouM74CcKQWkST3axb4+hrgCuGZo
oEJFNF0pz2AtXeLwBxSekr4Za1fnuUUJ3fn70zwCSZ0xylzzXt3JQ4v1si/r0QXNKCrZoGjzt7Jj
obcD8vB4XiPP6sJsE7Jm14HrBMMkwHrmHPgcvxziJ08QidGqFSfYMxN3qrJRBtNrAMEIbDFyZOZN
WDhVGlWt674ZAHV7v3VgXjaGCCrMGCvB1bDm+vt73WJp1fhRj2LVsGsXGbJ/06ll2ciy8UD0YzcM
WM1gyme91z6FYXqSvGv+KFNko5QeJVivLGGoSmWWaWY+tT18+j7YbyN5RXupQqLoA075Sakz2oK4
RRYlPsuILyymLh712HVIrCHUGrAa6QTt4yNZzzYjK+gpnQnvFm9rup1E/WdJ3bbKpaKwhnG3wa6o
84RnKyKsKThQSqC5iKCHoMR2oVCW7x/CsgOniFVg4oSNsrgjChFY9Kp/f1VmB+fqc7ECyXWoWzPX
DhXOtHe6aYAYWG98zPxdj70rKLk2So1JcGwwVmvy2XBWV7SQMTt87xar0JGnDP619UxU54tBXqXj
7njy6u8BI5GOnzwj9wogD6hoTB41xh+hOOClqEX2clxQk7DQ/ilY4hxboitRGxKJLAZIiblch62S
IAJTLyos8WQwM5uckHQc9FDqJyPmpAN2B7y/2MeqLkHABddhKmHav7kdX7FR6VoEsR3k3aWRiI3e
xdLhYbcTYNMow+uM7/TR3eJYiDKlxRjQEFmRiVey8chtU9CqWbIpM+L8RVcR2yWF/aPnZeGCGuPl
lumCcZzEMWyrHVdPHcUZjBFLQD5p91V7DoGq2Xeudbyd6alzfW271J32yVVdTbegzZPhphozBuix
eL0mioJr6Bg28Uq1IX1vXC/0C+iqhQ7YoaIbgRHdGvUN01NqCOuy5/eVkT9Awggq3LqBtkEptaJP
R0r3FL6J1JhSGBirtEQv8SNK7R9gSorWrXmL/YGnENEUuPFciM6gLoIc5TxljPPxLKuWgQr/0Xxu
mq3uUBwnBHDrK3jfxKW3k0j1UTFOYd8+ojwCj8fFDaR8TXsKq7KKA2gHd3yXHHWzxukDSYbpwm8I
b4iVnCaNMfWtT1q5yE1wkpUvbb1C7+WwWica4OvrzmvBIYLZg7taXMkEfJxZL/iA9bpK/eVYEay9
QEoU1PkepLgMuQ/mcqCA379PvIpEXTvPS2x9ZGlg1tnyuF+QNVk1+ss8WgRSbSBabZY5pJPxYA4+
qgBV/Q1uOQT12kb8/OrdKXf0oxA9yJuzvBvYypcUpvhR072M5rleaB2nolm1GE9cVgF0m9XEDcku
jUdyYhj/ouzHeSXj1fHDkoUfpGu9CX7pSeVICFXt87WIvpH5WkkWryYlnQdJJFIuj2cSjfzNbYdj
1uPmu+DqoXiwWoBpXZ5LicxloLFMDrYLNp4PkYei4Sxyau5LYV94cinuTIkI2vO5jMbFX53ngxY1
aMzK9oUvCuitYxUljsRHCiWRHj3DJCGgrwhJ8j0pH3qp4ACbexhan4NbXuG8g4c2obL89MJs2gEc
v6qZ7AeNn5JJRipK5zAMbpJP2UFzKaEuMXAJsFz7txoCFTXXhVbdgzwcOYcHKEQcVp1YpME3qZyb
6e1ksafDDgPzUgQDoRZNo+tHsxEs0yhAtEsnipyk8M8r3xmj5A5JIFC9kDiq3WElkMidqZQHM770
HA54PAf8l+4rlaJsHWG8Mwa+0zqI+n18bRMBtdsDtEes6eek4B+MS1ZZfwM2USPHfofYQMLveCBa
5G1EwUA/naOg/WHuTG+cX98yf1IN7h4SRLnrSrUZutfYwXkf7ueSerXbpPJJd5OcDtryxMoLKNo1
NcfIvnY74XGAoGpxpdAdl/vKp36KZBCUxxlMaB2i8tD/8J5zKLXninrUAkwWloeQUWSLOJZYDLXL
kcRK2RbRiLQrWXiVhrHyBpu2bkhmt1PjN2Cqnl3F+HtLxpvUTetvAKl0+yRiB0z8FS0TQ6JrARnM
4ajUI681ksMKWztHdIRLPA9rI/IOnYI98lkYE6uo22ZzWpthPZGkt9DL4vtkbSgvKT4q1m8sCgP8
EgkE3OdxJmwp2Ol/ZsUaKC6OTUTmYRsp6SsSjbjOlAhtTdvzJz1ZLxFHLxCZocCXgKy+frn5u5Ca
YrofmMzZol/3TDRaVhvMywsSVK1KXE9oPIbAubAVowOBMHDrr7hjSgVfocgoNyTs35ZeLzlGU6Em
ZdNwAsXUN3qCbFB15Gw0O0sZL8/T1UL4Hq9pyfK6c/6+cwnQ+HLw52rhTDeiEpZrvnoUuubq5+pQ
fuYW7fYkwU0wA0yU8bBfWglmqfd8+KchUUWVnvgtW9otDwV7a68hwbcv6Ppbf5IoOix8va4x2i9I
Gm5Nlpd2AqEz5RjY6kKye4FKpZKLoHEG3mayYnkpkdnwFrz9X1zfViNu+6HREPBOeNToxgjLxkrS
ryGjQcOTPUe1VOPX/LCo8C3zYoh0KrkebSgI9PrHx3rUDveV4dwc2C74ZvuSgIDSEGSo7bIKwMw3
Q+sS4vQcM8aOMTBG/dpkwV7COa4gViLT3KXHOXz6gec4SZTGiMrM8OceNVz+ibA3iOX1ecxtPbmO
gn0y0HPsYA9meJrzyjs78s97UyaJgFnlTHkU/G5tIKo3IhBQkKC7411FGyf7Q75NjslyHo5ewfKl
1WbQ3NRCFqcMqFmytLMwyxQ2TGHSc65YgxVfw4VT9zA4xao5e3cj/55sRY9ycYFhjjhpCNM6IygO
vcSOwa19seVNXSkOrjhsq02B5qwgbHEmLFnwVRL0jQw3I+jbyQbdmhEMgo7MqFT5JUJQvHRYgN2S
UBAgUx2ocMmc/q+5jwMhB+vL7+VshiWWsn+BzAX/vSMlRYPO77suMkqV+yDD3UY2Qmexr6b5XMWt
d5cCNywqg2/7l4VWtmmB2qpYUorA4D/+VdV9lh5vDaRrUktp0STtvmG8hYpkXyjYDHaZ6Q+skwtI
l29Ll9zpwQuzMOZ90oFkBvnGCwwj7kRgtP0OxI9sfQxSNNzU9KVwtPTlfIKY/9i+rSH6/hOzv3ne
EltVm7LKvf5FOuP0UCltJO+s3JfTTBG482Yi9RoWG6LJOrAsGX5UcNVAgoCjw08FCEf3W1zgbeJH
JXth7q2uVm72ngGjPAOBbbLBj+yAFRVFf5UuMgzkKX0SVUp6INNiDemk9XReTOCEr2FP353G6s1k
Jps1nNrWHpv7QMS3n5l7YHvbFZdMVaygC4XUuk14Vw7LaD5OA4L2VvkGStT2Y6nzWgSb4qHDJX5g
vCP5RTxEMPx3z4VPHVuVpSUGRLSIi5KPECjefHNT7zZMkdclQfBstbtRSqylMbxBasO+qas6bZon
zdZvMwUO5BcCGlDyiiXaiPHmUNn310GBEocoFs7CRfCbfMQYcU/P0IVjMzQ1nr0buKa/VFRnCN0r
07L0d9p8fz1myro/pETS96VxL7+55l0D1tUbPFLM+lSSK7LNPh7bYhCm4OdNnrtMDwFgt9K217N9
SP7NOPBQIhOE4kBhfFTvX5aNGeY+zFmwAEPtALwD0TwPcUN2BHSpZddwGmepm/uXCHwkJClCRsq4
WLmrTGmjby2x7IJJkio4p+6e+BgeMdmdIdVsC+kWwSE7veSM7P6ImUoYnNxoBWSJBh2mJtoz2sdW
WrbBueeJo7Dt/zrMb2VBGBJi/oR28YTuS/fDF535Vxn2afIBgbXWfI4aXm5P6aqQxd710Ez7XdUq
7uq4NlvW5/lg8T8JpT0PCtac76PHm5dBsWKR6w/51j/j8XTfWhrDl2jn5ynoUh8y68vCkDUVzqhb
uknn5dieg9Bh7wo32f20UWzlmE94xvaNSBmegufpfbhbbmWLjXqF/pWtG0brwmq2cLOo5vkojPmn
lZ0zQWdT60o5L2rflK7AUvucxN90t+98ROC763Lp+bdL76XwQluyAXJfzQrtfmWfieF23l3P0VkI
jYkPF/r6aNygc439i8rF5cMDCI00afmsm/3HPVPcnNEMv6DHjce7JM/wyvGTmVIJZfxqb7YIFOEw
eR632BFpxm0kSe6t8mOx5sopv3nxdBOL+bXCafb++PjnTjRbra4U7el44hul2A8hLPXh6lv/v2CZ
J+CZqCk081bzSnQU6O8yiVYOItFH2zTfKr9CRhYUKGX+3bD9hsYAlsojfJOpLuBcb6gzcZfR7KFb
2nZ8DnMNZM32SVDaq6tOL8fOv/fr8jXEZxTQDuTU0u25/3BbyOaj5rhOJDOQcfbQIx6su3kc0E25
Gfwv1+67uXEQO6oqzx1OI2VC3TmoiPO2yzrINFEcxzzHlBFeCikJ4mkxCjyC4I5p4Yi1yGx7D5cV
iM7KKD9ydgND3YeRDpRJxdkbCLnHnkomykNJJq+qcWNWAe3s94f6v37TMdq6TI6sfDDqjiHX/zNL
LhCcXuGlknHnN37c1HcpkZempQdb4J+cIXqJWlg6vgd0vQqlj+e/o4WNz74mAyj1Qep2txVWlwk0
vQHi5V0J00d4Xsh7lqvYZrQT6yqujtkcZfHJ9IwRyEDqR4HzYSnaF0fCmn1EzU8NUbfSkckjCLO+
UlWXuCWK2IKvhYYEGIAehg7l5Gy+FML2vPuYihLWbaZe6YCQOLTxrXepPCl3m1COpwwJlaaJGyM/
4hpNW4Dnn5s2BOCp7swhDMuWbGKMLasnMshbhVY2+qdVqZQi7b2Bu/Bgfa2qYAbz2/cPpCo5bzRS
hyu8nGUYzoSab5t1kCnU7Zh5h81/Aai8AEchf9d8q/ZXJ70V1qrEYLQ80hw+PVxXWOf0shOn26m4
gkLJ+GxCJYsll9LbyhMAfMXrcsWl1ayFxSDWsrppq0sDQGe7iUH+1vUtuR+t0TPxa1HD6nRJFoVG
PRW6O7h4PU89sOhB+ejzNuihJ4mJ4oGJyXJO97NrmrJOkWejDC7sssdY66VuNN8bIjXJAysS+OdW
Rdcr5FTBOUZ61mdcQqRO3+Uq/g+4EmDek87ne8Q197upTYRHIgjlc+BZrzorRmLHBKbxUVpyybcT
8MIuOoJ0bgVl9WK7zogsxwALx3m1MSE2zTZtf5zq7RYYrryVFWObGXkj4DlorzUCtHyt2gBZtnN0
hHfvEuC2++ZqOljvS7ZC/neBAPeQ9AVXxzpUW4Kl4w8ZGXQUNnrJ+YGncdwcIHf3ru3zg69Jc2tf
t3AciXlBLujunVxBFL0pI/JC9oMGVNCqQwGCmZ5NUi49uvAR+OSyuIlWukGK3MUuvyUahqNXzjxG
mdaHoLfRmFPKUo8QEXpYDIW9MXEr2Wd0yickgKNt9vYcZoN42xHJ5vO2eZWC1ewKvO84cTUcYO56
b7XuRi9du8GU/f/H4MFbztST53xCRbAppCGTlctZZ/FgN53m2OBLtZbHvVpfYErUxjed9oTYAN0e
gqP23imRo3YrNk2VqgOpKNt8gaeD+Rj8SkODeG140t9eTzNG+RgtloZnaujW+U8uOu4hCLrtqoL9
4vCmQyMX1RB/bOkotFP+vkTFOHpPUVMYb11HAD4LUZgWOif6SUKL8mB35Lk2yXya4TIBqM3CrNLr
pdJEmGAvfKNVL0x4i4DVLK+wfivW9y+eYww/+hKp4FXlnhi7fBu++AyIplm2OregJbFDDXwf251h
8H0Dry4mpun/RhAPHALqegAzuRNRTlOqkKZEJlqwZdpD3OGhq3Vl1Rf8iSNASuOOqzb/C0/btJ5G
t6ROohHpBYRTYjRQ2lTmm2LmMo5o/G35w3q/BFyOh5uODBTlfjNmmDHqSx1tSQLsWT+U1sst6VZP
Jp/tSJ0jQjPg7LF8crtb35O1xzpTGn9Gmg9yq+owi9JqIZlb5fZBJYVIHaL+zAqXmHOmZddl93+n
20UlL9SNxnGeigQVTQ5d4GBPdwxG1hWQ7Jf+vZfR4yfP1/D+r2HW/LIzsvRnWVjmODqPCC8kp5oG
IB8CxejlHWCJ1mc9reqd+1q3TwyBiK1t6nNFIO5Yh35gUrKf4us+L5FzrxLF1vEtuo5dYuE9hvmJ
ET7wP0cshLoX3r63OzLo0RDvcP1GEx3bGdT/8w/EsoYp33zRR+S0cLTtbqejN4wacWO7DdJqtebZ
cGwk442yJ9PqHteHMtTH9n2PgbSMP2zpKpWFXIA5Bh/6qW55tz50n0ZQXYrl9pJOXwBvmD5yUdDG
D1ThbAihk8WAqn6ZKeHtbp325hNTPWGZF/P0PCiiiCIlNV0uhUQWWHLo+ykQgYD3RskIrzKxfegY
AFjmn1RpnyFodWrw8zCIe9Il6P8EjoQOkwnmSaJlPqMyek8UfpRdwwmKfffGO/KM82SXZfM21QgR
/F9PHzJl7VKwh0XI4CNLtjT+LMkg55pckdR/fP4Ua6JdZfrw7Ir1TJcYPhQuCY82iU+pEVsYctqo
lxMx0mQEx+n48vOQebqK8Kzt+hjl8jpakMhkpiuYXP4pfzcumk7JZJRgqsRNYqvXI3cWSza07BW/
BSxUib17AXnbnGIEF9qVwk/4nTxmpPd/UkfrZyZ5S91Xa5nHFN7LOZUCfZzMXUDKk0bmezalC200
hi/9rxmNO+02MRFZf3YQ6qn681AzjtVhrUsiizHYnm7Y6PlUi3jRnKUdZVC1yD21agxTNmuYZEjx
0gw+GR3KvELVVHWIASJrKBIHXXLq4y26+INIpGWkxGJfoHDvcNV/6+ogJjajb75X+0AQLo5+7sNd
sX04TB7ykmtkYiX3Lk8QGk0BXIyzpmJ+n6n2GDdjxgIXZQCIDpPVezz96UzY+U7v2atkpuKKdyjF
CqlNpZHOSvfRVQx+A3PZplsJkkLcI/5Z53faeEr8OWCfLQuNYhak0BdPN95CM9eGZqZrujzY4oug
9MwqLd5PntgPV4cLU0KjhhkkPkgP4gl1SnUMIXycvg1HNP5+LbKsqvFQsYloyl+uHANRpb6RyCh8
XanRmvGqqWCxic2jAuKR18jMLrz0D5DVOXWlh1Rv7IiznWp93QE8SwSZEKihhG41FyqdBlrRAvkc
kn6Sgh5cUcR6KSvDlnPPQMUNVtzI0LcZPbWgO+OnYvbU7QtBmS6sSN2K91ScjUY3F34v4q8zx/kY
6If9D6flQoxT1O7Y/dpzEpE60+zc6RziG6gGcMoeOm7J8k8xj2IH4Qa3PU6gweJ+P/5dMLEOl7w9
TBgqGleyKxqs/hf5/BgreaFebZoNO4YeGDLt0NPLb3eicSKmFYqMvjfWGolqtpL+mXc9CnX1RzRu
amTaFncSTJLf+AxeWIyUyqYkGRXoTzdt4nIUb0cdNREiKdvxjZoMW8iy9BAB6pwHHV6mLZG3eyn9
uioBi2ZDb4IV0lL1ov1/41DjUrbxOzMqCmwFxWPe/tAsRMHwsMDZebGzZBM2jlUWyXkblzI4POvb
H8Gw0sBc3R7YE6/MGFGcjl7+06jkdIleGqeQCxmIhv1Zbfq86iU/8j1HaZx8di7X6wyuaRzkSZCq
Z5NSx2pB4/3+gUhx7S5gXA/WZuF960yD9G1ZzaFJivo9HImuuH8LjwmF8myYip9SwAmu5W8PzN2c
mpcnrOyWNOi3+eGybWlkjp6M7OD5/i8TAoEYg34VTqxIbtQ3QYu5OW2CiiQpoij4Fxhq6pSo+m0p
b8Mfnio8BZctES/wctcLNy1wZvq88Lwl+NKPxp0k2gVhq2hLSG5RWACsv6uWsfkH/YyCU4ymJfjP
/+Tmym/n2jpuwDwV665dHxbm/VJvQKA77rYtYPia3zbmvshjUTwZPXIq8upngNJb1XlIo6LxcPIt
L3zLd8WnvXRW1FujedG3i8M+VpcHuYp8/40tRWAjDDBnBBjMoumzh9j8pDBFUSxdgASUrh+07dfq
Tcmtw+Niw+sYQEvwqb+U6JtAFD9Gt0rE7BxexPc8vv1/SaFTv42yg2YCAtxuahLjXXlb8sNBmyeZ
fQr7wZ/6kktdYBwpN3/Kko3qd1dFYx5EcOWv5geLZXUq3YmFiM3LrBDenWGZP4OKimd2SJ34tRP8
XMMHndC/Osv5A+x34zG/GoTiUMzdUF/bWjZncjmIfQnPfsBrNgRHIJlbn+tJWK38jNKOHN/Dro9z
tAjOfad7bwZkN7JzIvpRGPMFvj10Wy9X7gKqi8vnj5boCeeEL1ommsvRHxCgAyGQV8o2VG7oy+bj
3CGoBMcUFxqf4t9oAn+yhNWk0lHvcMcgvaZawG9sVZaW28tBLVoHMhphplDU1L0IEN0tbbqDQ9uf
UJKCphng6W9ZIdN2gDHYXIQF5fGdszqcF9f/8V+n2LMXOV8wBQXgueDGoYcAYZ7Wf20u/Ix3YMJS
qlnZD06Z1e6cI60ZFr84Voav+kPa2TEROyo9NnTGY4kZffJQt+pKxUIL6DTczYxYlRLQ0E3piyYI
N03u1w01jsqZNA0Dshk7HZuJcoZe70Fuw5aRynxgDDqmgYa089unWXLNS9GtIjH9nEZKozWxVKjh
m4bjXimyGOdxHRgpfB5wOiQxksAErMmGEzqFp/dW7yDg3yIsMWt9Z1rODMFkYEqVeDo7hINCsILF
ZMPHJXh2qkBH75Bpau8iPfqvHZq/xSYSe+3OnlcsV94yWF4SezrAg/Wqh50Wt9Jm+LcPWjGJHqo+
0Air6COlsUrI3bfg5jlaoLeuvYFLqktqRovH5rqZBJ8AUQHj4AzafgmBkpTbMM4LGc7IXxjVS9yB
Of+kkwyej+I0dxZofuTI6eQqrOfj0e0VJRXdP6vvrid4HV19tJBRTBOMO0qiFGsId+P1IZNbcDZZ
gkJlTAIusFuEmOoXzo9tgGqK58P8iV4AmJDJKvJN2gx2baDOZvLyUwNCw8qWKz+9Wn5iQkzZ/23j
WR5n9R36xQ+ISTuZfPzoNDDk/1jH0alDDy5PT/7ieSNcJ5nfp/er7UsAcWMxsvuZB95GEJ2C9DUL
dg7DbUUZ4/9ofcVc07XaK5OPogWLqSTWZqkeH8kalKre4G5irDoZn64XzPFYVSa3LbBH79qUWQqR
q+LngY2xX35N5yWj8oLD9dw2E7ZuwJKwLVZLhENucm5JONcKZpvkx7O903ktbPMmR/R/WfY2cuhm
h93jczfnSzyPHL3SfodBNh5+k42rbW7Mj0m1BZFeE7+6hkRS1fKrY5NkFk9FgDmEyBqBgpRlZdwU
p47TyHHIahYQBlxZbaLggX4YQJ7h2GQBUMxS7e1WGNR82Tv2s+MR6nlZukFFbXj/qh/MtnDiBQkE
p7VIcow2mwX9oQ5o2KmiLEmeZ5GAnjRaUG3nhfZwUZXhLpIrFog/91zpQyAEbhlSiALE/lGpMnNv
DwfxzwJcXfv0JryOdV4Dq2EKSjQH/iQA4Kf4EikSVxReTzKFzEcV8o6sDv3JRrewtdoQRhaf7Jvi
V2A9WQ0u5RgIluPwAPaxDg1knXS9UZJNHjOmheG9gF5EPXL/dst0mogPqCLW/JY5kQGvTIhoeUJK
FekDZEX6Jkdu3sXNpObuc16AVY3KJB70dUra9GyAkLXLeoIi5N/KycuXo7LYsVUUfkmd5uxxrIaz
o+vmMHtO5nbmNCF7V+naUxv5pTLk+vVCFiZxpFaMrhOc4IfjFqo7kwKc8WA9BPte9xjrU0FkrF+9
ZlpVRchZJxZ0gifwx4tRDptgr2PLqf5yAXERj7HDIglPCuQ5ICVk0pjlFEk2RHEiccLb1BLOnwq9
JRxxj+PCGjNFeLg8ahVBcBOXwjPl0nwa4escV32YKU2IcvrV+sn9NhdwCupbeEAXR/Ky4j5JE5Mc
+sADcbpPrl3LvL5Miulg+D6Pf+kyLpCDp8jr27e22OQH61L60uXmjc9KGfeiaxcKiauGFY3U7V31
Dta8n1GQspU9PSUVa8SZQj73fp2T46c4lCsGsz5EGfxYowXua9X98ouv+VH5PmuxLBG/18wp+6Gy
yIINFsRDh/wdpT8gExDUh0nWuzb9fDCcLNMdVT5dI4jhXFO7YOK0EJN9/QZFON/5JaYOg4p3FAzy
Uzm1/+HreuTGaxSYPawKF2IMegp6deGskN6xd3VTc3te66FUSoivvVMhK4/G6j5PvmEk5rpYuMAm
2c92tM1Xb465t7iRI/XEWJEwS3clADWVfbOcdggxujMGmvqCiYmYLgSgEeHiACIUqSj+UbFOtWo8
I2J3KhannBHu8eSGv7Q0lzKK9XtC0eN/91YKQgLAOvqQ3FAi1LEc+GYBD2sUfmOUxF16GimrJLKi
TZXpWm84+dpmlv0iEKS7w76OjUdHgyvWhvDprkagTcLVzTFhdeXDxv+K8FV8iqK+VPCFWNhCyJWp
fXUCrvJ8cC69ZnqgvemeUyURWNLbuJPXWnClO2WzGDtuTRyZNTHz5H9sVzSKKbsnfxvk6t1ZarK6
zt8ROU68AzyboSxwQ2wCi+fgvUKXZ7th4+X3bXyKbeKCbxpUiYe7RoqCqlTjWFdDnZj1pYN5Hy0R
iJR9rCAmjKBLixn9C921/NgPZthvutTLfHx6zkTQw00Ul5Xz6VW3BGPlXHcqaim23O/dDozQgQPB
QkdEX7LSOVk6I/pfQWCrDrsYz9e0wcecBUjPnE5mtV+m4b+pn/8UQIlKvlQX1ADwK65SFFmO4GGi
xt7y1cD9tHr55vWPwWv6tqm82ScBjLEuZ5IHykN4dyw2BpHg7Y1gCESY425POjDtaY7obIUinsrf
nKpRCMlZRElqXhHB1ZWx9qHaLOClMad36y3ktG7dO2F8pmiI3nf9hhUPR80yfimAL5mJAvaTTgvh
YSEgstyt9/XQM7Zx23zypREMnduxtshoyG4D4czUZngxwFkwG43aH2DPqY1CyBU1LudqvmOwH6Ih
xzIx2WI2GtUemi+YbwhbX7jszseQ27YAKfKJ0vOrPSYwb/mvXSWKiSSqpo5HMCeQQkv97iqiH5T/
F3gDOw/b+Bb2mLBguPYeETFhM6rPd+yZ3B1gB9rp5I2Nczi9nS3bioJi1KwLWlm0rLpi/Gjj2TTv
Ti+pIFL00f62r+Yv7p9eR3m1btOB7NwsTd8/Ze7IPbbYhtGfFbLtwbtuSvDO1GVnUb8jqAsv/OEs
3ba220cI6sGzQVokZX/cDJ6x6lITftIFE+vNY2Ui8UQpJZwu0bGbfgEgO4i61O03yTQb2aAJ4Ihx
iJI7hfuxS0wFmF5ahq7WeMoTvycYRPqxbwNHO3Ok5g9aUlyHrfNROMCCj7Daez2j0SkDHJ7m1LMU
Yj19AZbbdfvOFFgweA+0Lys4Xq8XaiO5tsBDfQ2ht3BbZaGdjiVNNNkHRautc3SSwFvYLggHQetv
Qiz+nIH9+qjAlNJwkL+zKLOWhWpJX8ZptNUmtpM0v8vmEwXU5hdsbe8F3u6TDkR61rHyDrb0zowa
aaTVuO09Z6yDuPBSiEklQsJmr6g7oKLSDoj5qWBRnQFGnuzyXzVKwgqY4LAs4pphO0rsHLWHJEhj
zq5IJMUwx+0p8dWw4yL6KvrrZZ/1iYjBKoU3oK6lYxIKhwt5Ubyntc7rCfhNGQvZ15jjEYWkRlhM
WyujFoBAno4mc/tCuqkB46H/gLs0jRC+zYWR2I1T/Km2Ef22QvvceOUBgKG3gmNECqdFuhY7M+am
3JobJKt9UX+NF1Ub7oZ8FTYA/0JCcPm2qwAZCZFo2LvqEe4S6InF2QKGN21O5yIPAioVxVKDFX/f
nejsWOOJfImbH8W0pfQy2d+Ouu9mIxKMErMqUSk+LZa9q9W+PMTxKCyE63zRAR3mdCgKK0+JEOBE
TcmW85MYdiN63G+jE39LR1OYvtKxauEyEUsB1a//RmM8W5xexPhxJEe2y6pswPYrXLk5q7bOHp5m
riyzmo2QTW+VXxTJxObIukAan1qt/Tz6oiCzTIsN+Ll0QiBm5oLCuLiYOaM/CpncoIgKneaC7EdX
caSSSw5iMLw+IGjd9Xch1H+zQ5zJnVvZzW00N47DHwsM1YdOON7QRJY5Wq4ZeIFWMzWrYqqn4BCv
tU+exjHWEFg/Lr4ML8qQeQS37CGupYcDKBdFdK/VcoBfQoyZxQoFEDoC4JJ4TN3kSUVGhfwGVFs6
DvnjqaQ63oGNvPLkWXgalVvEenQC0qoY1qU67ZjuFhOakaEZOicpnvwW2gquXaQ2vab3HVOJfGeQ
LmUwoyyzXkTlOAXMyxmIyEkuKr5o/Ys4xt2kxg7V4jlvYleIs6VyLP9nVigcQqoIXP5ixEuHfHh9
YPePpf8cvNhY9E4hpAYECIx6tPn1m8pIsBjtSWbeuuShQoH5qX+miXGK0uEKanyyXAO9QDd35I7K
3JZz3DEND6P52irZQizz6mRJh9YVa4gKgTKXvTkuyijVwiwI/B/nRX572f95JJtkOZhXhL8dQccm
MXaM5t3irXpPC35/5lxf4cL/9LMOpbMORXYIV1nza+NoSWBk1/qDO/MW7KASceltsi/WgFNYNxn2
YsnDjHZ7umCoCpz1WS25eABOf/lsJkuLtpbV5QJCheHFtVg4xPSyTa4NIYz0dUYNMP36CECC8CpU
ImzNYmT+5FCligwgRjzQuDBQ754nY7+FUGx1o7rQRmtd29DJ9+wiGmZgGMeKUppi979SQ0QqwgvS
f4yC4CBJn8sWAam25Ql3tZ8WgiNRgd3UKlypEHwuhdKsgFjoZcVjalnBNLIYcGXMx3JOVw/3Cywv
w2LbsZZtrXJ/PCXUDnxvvnEuo+8mq+2ec2V6TiIR+svezJAIJ480GtxLdDO3gnFcswPbK30e3AqA
BDu+VMw8ljcCvksWznWHUiJRgQ/2b3Eu9l11T4BfcEikNJEO35wm/31DhTDkAVt74OX+dbO7mroJ
gM10D4hqUR0YtUmAzjBPfVf3xvQrWTn8syf+as2eQErXaJskhxysLv44U8opI5+jLe5t5c/cCt+l
vozZ+bGHeRDsp3WeCWG8Si5M3NCGckmKMV+0qkD2dX+qj+RI+lbtkn/FqTn+D1JKN950qYh3aSEp
IdPzjCSkmVt/46//ifvr+qcebm+yqRjmlJdtr8pV9Lh2Ve06xVFLOUC/PYPXeTfLAeHLj6zYBQia
QjMdpcRlfWyNCCJzASPMMy3aBQSZV74OgQfoWm0qTAyExxfItjXoFhITneWfinPt/fQcVgGkcDRn
nr2TZDbcv4dXwJRXq6I/rKOi4g9AvlgdTu3X1kCYvEgEImRt6o4Kct1klSXENJU//nO6JKyl9ZBz
NiqPT869IwEitNfh2jUqJgsZd1E2FxQtEdYfH9vQBClyO29lhjrhKbUbAQstcUt63PPrv+13VOw/
FBCRxGoryYXHkubU18e610zIYvKE99hQxOZlfQtzmPGVZxNHWNAOJw0yyYGlD9MRXlCVOsRZZ3yR
3OPu5Q13ABRQ4h5qRo0SlFhRe53jgvkQfWTy8WrjprVhlwx49djdFrj5h5PSBsp/LNrcybSJiPSp
V4icQOTJ47NwzO6Nmtbcbs8+lRJaxFF+54MezXPFroUiu8H0injtuIQu2wPS+SmCYC6AOygc8Ft6
D8SRcaL223kahH8NHPw5qR8wQdDLMPiwUGAivJeQiiPOO/kcotAMH1+cyYOhhhG0eRdtJvxCnTn/
6SdYtv7b/yLVAyANplkpoTvOiPGmD3KDZ3/axELyfMCztQnmsvmy1+12TaZv33k/QMLtpqKBVbX5
nRDT2SEaOwZyC1KD7teoWQCozmfuMCQnOVLljmJhMYiC5kUALT+UkPjw0uIzYoMPT/qyFY4hNFxv
CWck9TbzLfk+QHQqPorz0rWbAMJTx6gV8TMbqDhPN4c6vmb06Ydom0bGCE/iqh3HmyNgaXbUTfv4
6cUJ2zkL4gqrTG87ZzFe/LkbnEKS7g8tSktF+/UWRcC6nIoAbF9z/WROd/KF56mvB8x9KqywleZl
twKXzSzg8za0WQMMKjG7Tbdr6LJPtNMpI/J11BwLEMyLLvm9sEZqcf6xxL3KbXA1pDVmLYxVImDR
bh80EoFnm/NlQH24eDHaqXtdZnb6hCnXUlZ5FYiLKvuq55Vq3uxWhaEAFi1e0KsMwbxxl3qW4607
m67Kh1Iwfd3Is+Ml9lp43fSR8H32/3zdXejVHLxdttVL+kVliF/Yjz+eDmTck4SGqXHlg76vLN29
PSmKpzCMTKKxsaiG+sIParufqs/fKHccdn8DAm1zP8xiH8iKVBRrMg5pIZsyLgchIOJoaHsAA8zG
Xnqp5AewjBsTfxOT1HVYsbsAcOv5k0cCZeVYIbBN4FV0/XiBZPNDTx+0RQI7Pn1Tp82ryAtmNnms
QTz6WoyJDODW17NU74hGTzKovnLCXtOzXGqv0kNk27UmJfyty46HGwzZGgg4y8dTQ9drb+MyUXQz
dt9U6vW0DI7OA/JKC7XwkJoKYdRBqn9hlu1E3LAuX70k8QfaoNX2utorHsjGjV+fo7TjEqMb4/PL
U5OWDfr/MjlHofzjcbcgP8hi2nAo+chX/J6R9b9YRoImgLS+0+Y3PfLb7SPSHIDH2r4Y5T96+RJ4
DlXoNgm48078AtZOFshUl+zXf1U4S3JGFqZomrGBVOvrh6J2tNbqLUY7FLmsI4s78+w1vhjedQmg
rv+1h9ukZ1oKzdMro1Kt7I22sYBtrmUIfvqE9R687o4UdMI6up28P9TzNjcYHXmr6nkZpL8a3Q0S
8GULroyt1dkAlyucVheamE6Tr7ytxl7ZZBWfkhfpMrNVCqpvQLZZwBVeml1rMl539+ySgM1puz41
zMAPh2xB9cceolHxdeza3airCtSHKre4DjjGRLQt+2aDX7cqqiEmvv2KuBYeiKLql7gjhLrDGBGr
fiNsX4CLkzIX4/0PF4zWKTk/TU1YuHsKpwkup3gv2HC7qQGdqYc5Qc7rcCB5NJsfseJN+cjFYmBw
pk6saSPfcHA+cLIyK/j9YQUtLDR9YC0BHWd1lXtm93qc27wF659YVUPe8cMdVBDEMR7rZgD/zOUH
uL8M07J7dj6+uNB0frv+xHm2tdLxbM6SLsj7C1RaxMHU8q58LnEfZelVcLNqFTm9nCo9sSbV24t9
j5CiSgkonxHO5wvlISaF4EGfgF0w0+co048Xc8W2UjcSl5zZQ9RsFip133MmfMKkM43FsKA37Y+g
dX9HbG3KTxq8kVhBemNRhsGd7elaR9P917KfA5zCn8mOw+tpuSivNTbY0SyXUuFL+5T+uf3t/oeo
LtSZCkchTAGkdIsGMKJZtx7NgtrKUO7F/g8GWwgtWu51f0hb/HPCyWnO2WK+sejZwSHKogJw2RF0
yTzw962YgGZzXc4ClQIPeCZlBBMvlik5V9FHxNImoHIkNTsHIgXzP2M66+i+CzruOT7PIN5UnPWj
FcH32c60hQbM5ISK3VL4xjghnzFDezuGGzlcQfM4xVoH8EB+86owttADlrEtR2auI9LUv1cG6QYc
WzD370jODNLUvgAO69Uaqx/3egzzWtGxHJTRtw1j8fb5x6LQTugBDR/OZFM2kw6Pq+k19p/QCq/C
qur4kREqx4GIZtTBZVEWOi7Q0pl8JDBcklHDQhDe2hjPMnDqYTa8Oc8Ccw4vXejUpdPa0Um9AECF
qGkCZ4f9G0lwVGBbFHAx6ulqEfnR/vX1+m88VtVqI3trOh9LVn61wJtEMuGfl1mdPyvcz3UQ7pdh
B4r5QPolLExLg4WQa7TEyZ5rfkjeQEAnyVyC8K6Oix1/dMyhOqeg5i83tBaK7J3LF0cqfVYkE5RJ
AO5dP2GhEHq0vgYQtTYJSuYKXGXGQVfyiW8z22/fhFNrBwCpyMsGV+wtP74dlc/QArrTK2dkQHjH
3s6ZmQ1uUCeWOgdmaY40zLogSyWP7f72gjQ8iX88nSlSJ7EbpnBT8sqCPANHnBCVvPVOM99iIuMs
O1AaIetHr9Iih6p9QtW8Sc1AT5w3qHuAArFkZW5kHyAajhHf6dg3hljHMSZgYJlC1GN0+icoox8s
dBiGPDz4I9l1SjYrJAGta3l6yPsV/9rWjGKNlnFDEa5R7uDYKFLPhym/h3O753Q+15ac/jPSmRkA
E7T3rGMHXua45jjc+FIBeZ4TQ1GOYCp64Wolwa8aCRKU3xtF+bGVqffmG2hhn4EiGQoE/AYYpslZ
RFZ0XWGvuoZ+EFSK1AX6SFGQFsxaXiuBiS+j7W5wd4Geb8ZF6ulf5akxHMY6MJv06QCaex4g/Pxd
VSDgqIhR5ggy5X4N8sLwmYANVVZcadBe5mTNYJt9TxjFldpUf96DwFEAfn4/D+Ffx2k83yjKj0St
s4A5CKwZxa4lerLfXrgrZP8hzy2+fHbTiNm+nwbKDcnY8mdcq29RXZ6DUtLqDDO2G4uyaR7tnLpu
Ewsq2RKfpflnN+dng400YrqPsHoV8NmgK4RdXTInFroB/TGymONSgMGH+ik9HiC21NnvxRgk6smn
zTnqb+v7B9OPul4l3YqRXH4jQLE7f2MHLuH2LS/KCi/dweMi+FZOQoXdl8hS2SxZqfWpj7eIoQQV
Cl08QeGEqd5Vyici7JmHZu56Vzs2PqxcZdMGX/NgrNUWegjL/Xv9gpSaglio3mA9y3rXEVlS5rvM
Xh3ROl1JIDQkF6GXP33am4poA0lN/bH+fxbByIe/oBhJoe00+hUhrHwNQmV7F9JHLoN+hieRYrtq
5Fh71H/iQZBMr0wZNZWMxqogc4AZKmJ52ULyilnddguVkshtqRW8m9fmGBBFYiBovONmvNbTxpK3
40Zpcmm8r+dZBkbvhchHzQuQK4zesAhFOJkgfojccvE2WyW162aCT9qpsHZEZBt+ptv2hNUhH5Z6
Tl6JU2yvQKL74sMrPb5DCQsRKgN0WXlYVZN72n/x5SRuGzw3aAr1CffGDUHK3Lw4jib4Kfjp/4D5
vYzzdFlPh8pfsOGOjWo3a7aEcIZtVZzUiGNVQb7AbKeCw99qPigKZjKxNGwu5B+H+e5M53wg0GzB
rKqZeFC4DyDzQflnrY+JY73K1M8UvAdqjry4X0drjLSaCO6yLd0ddOUUpJQgh2BO0yD/78/4KnpY
sSvNT3v4B98d4bw8bQqyhrZsXD/SX97xdkqCJthDzWibMZn/DkHl0/KoyMNGoXI1jQ2cr0a64j44
f7o7nBFiU5PzizaYE0kVEFPmP0Sd7MuJbEcRXB7TSVPxMYchFsW6oGCTnhhttEruBZRwXScK/DqF
pJQm7W8dWRvsUd+knSuwg5QsMt+p7PshbWNq5xiIfIwEZy6BAyT6Jqf9SDgpilnRclu3BdzQjEHe
MjGDuZGKQ0VTZa+8k/UxYzYhck74PzmoglCASc6MRDumA5717pNAHDG5ppQ2yuBwe5hjfbTxOvvq
djjNtbwoCEkXzOsdo99At6ZM47Vlq9ZGS9WDPmIFuQWQizdsFrP1UVApMpk6vgITEyCaWAeNXxx/
x6BZ2iH7Wf/waivIhUbGOc/A7rFg6SHhswFBCidaFpJ2Xjf9ai2RjZaa+BoErbQgag3d8tQ1gw75
sr7ghFSZ+ErO0NqlB83/u8ata4N/Sk6m51st/ttd85t13jZ2Lcjz0eGH3c/Y0QFXDNK2OCIh+oFJ
UM2ADNu4MIgVbk2pZHj+wqcf9bvnjTDRbAw7LWwnGj4a9f8zw4P4e64ADDhLGJ9SUkHmPp+ACafC
FYKGmGzcayi1pKQJWY//bMNTx5vCE4saczkJS+4m1v4FoJaWoD7KazgPrao8wRw7NojRh6aza8Zw
wwD40Xs0zS8RXrRemz6SsAShlm33TbgDZV7OmnSQo/rhIlYbJAz1tBH5YzuCT1eL/VtVzl81CZgd
gpeYkrBxJxvjXBbcKk7xeBcKEyqCzUBS2H3LRzbcCdjp8lA/0ori++GXxYsAjmFujAdFdjmnsuf2
gXJTyh0X1oIzv0wJ6gWw8WVV9/Lt635rZK1WB5e/x3mUhBeLa8OFWwcP4DPx7xehFV55ut8trst6
H4ltS7g9/sQOe0KtpKttco20eQpInYX5MOJJ/SuwZbASpvRedKRt7KDhcUJ35NYj5uiqmGKB3N7E
I/cpFSDrsOwH6bnIZ47TgZ3pSPVjwFzFODfomyGGXaymr+2D01fS7MBd3u/a3bSY3QtTyFh2UwSc
xqXrHMLcVdad3PK2XHpfUm4dV3BqcBGapuURgca4Yls273wUGMqcq/Rj7JAysaTANG5EweKn0eIW
UU3ddKYl0V1fwDx2dS3s4jtjTPfcDNkaCrxW5I8PIr6uDc6bvxIz4gwBFtrPB1HpUGb/gIhXHJso
eKCJZ3o6uY6WgMQElVqgbgOV+fcB0REzjc0dmzfT9lGbpC/ABBP14rcn1cVXw3bJ8dGWXETE999K
eJZKV9qDqRkJWG5FKSuavC92OI1+Umb7bTF1gcIWchtWzWlmHxtcWWaSbfql19XtlBUKvZsmOQO9
xoOWO8B1MVMVDIEhkTeU5Xx07GYUdkQabS/FD1UdEq4L+YaPla7px7c8BGNnTl+i5sBBvchJKL6J
7ThNLXfrXkdKtEr1CxJWkFfV+QU/ikL8NdTA+SVpcrQx89NpYsY8E9xVmcX2k2e7j+9M3JCvFfK+
AgGGqVNjwU0TS3PDWViiJrw4vBdytmu/hzge1WTEH5z2qrj890faT0YONBKSpFkYwttYSpTQqemw
2d2wYqB5t+S5nMhY/PCwk25HO0zA49x0p/ic59CIty+kTE/m7HtZZzApfiZmn/lB+sbXhqQiQM99
aAckj+bNO3kJwMBN1EfKZr+s2K3V8rqhnm2zoeBurwOa8DcSV9epq/HMoUVFfoFDgplt5PxFBmHz
Yx8wXXF0s8Sacz4OZSdm0Ux+2G310MPdv6KtlK0UrJSWKRROMej8Ho1in7hDRCuvAIyi/lhEGmVr
25+1k+bTnnFAJ5yD0yC2OjOt6DniPtYL3FeZXouARJuo3dFJWag6kHidp4TXKDHCnvNtyoaQWJNF
5GxxxPcBDQ89HOLf2ZpEFHYVS6oXurTwWKyP652vQ7D7woBlTwwetNu52Dq/JmkD1o57E8KMUKQ0
y6Z5je6UCmxW2Wz9m5yzjav0pHtGD3oyNyT3rLejx0zbxuywk07xQWrkJViA2Dmc1zqkMtHjV6Bv
miBDevibhhMB8+flR+rYjnD2VEO2MTWRMFyin/9oT42R2CczR/ft6Y/GXLuPfqGHz1d1t79fF7+D
y4Ap38j5YSZ62+5hE/JOmM5KtnpACd2qSuhSZTkkAecnlmsSpiyhZrP/ppiv2WfBvx3X9z9q3EUR
V/CB9wRoNBLG0BAk19fyRzYvC2O78+bZUV/P9p6/AKQ/sLPylGFyiXBodzn/aI65t7RJ92//Mm1j
5RqQRLnJqAZxZRoLdummCWSchQq8BFcFEvqzExXu5djr5QTYE9WOuMSzIX90hOWD+0xpiJPp6z8I
EibGOWwFgCZudOCo/+fOWbrSGT+wfbjOtQFnZY8KE28bztkHJqfmtM79DTKNqpacuA3ftndwKKF8
OvKZmEu/uz0+HFFUkDLf3gK1HViOK5xoJSGnK0vaqLpHd0QEjYur/gn+5gret8HAefn2qQee2lX6
nndj0EYvTy0cvQR8hlOcgsw/IkjLInKaM8SE6g1nbAA7YmqwJ/QCGtoPzmscTJrhlepOx3ljKCn7
35+UBpgfJ2jDTZtibourJZNlX7QU8WAAYEUR4fkjBmWej4K555a+O13vOS36jC6HTH/BEa2R6Cdn
Eg9WYBa2XnnvwM+Th2A9QIXXEfy/ZBJcydzZaqn5X6BPC7e1UhmO2LrC3MqzOejCRQmR2YO3JV6i
u5Ul4MGe+dFChqastwi9yXhZs4O3YBJp5XniwJEf/MnuHDEX+hvW25SpGD4MheqE4inDpcsigIsy
xYCfYRFjbneWA19a5X0+l2ywqLwqIe4AzdFSoVeq+qed+kfdvXtzkekXIaQAn5oyLsAFhNtxRv/n
E6Sti9hR+/lBM/xLLbN0kRymen85a2ubrwubnhLBE9iZRPYYhNmicJ1nFz3r2dzh++3DVuDtAdaK
ToN/FY2m4sdbOiGamOmlYTomk1ds6EiKkrulrNOzs/E/BsnXADTKizl/g+I+ghl5FYZNOGuWpVJI
a6FM1k9SzKp3XrXMbPhe/mRbILGlfbAJ/8Mg1T/dK+RPafD7P4haDqM0H9QBGVcPUF53BShddCV6
XTKHeUzqRofKK0zxJqpC4Mk5voFVJw1PP+OveMeKf9nVB18+PELMuFVTQXLjBaOf5lk2Y5cz8KZ5
eee0CpqJ3/S97TNhgftBvcy47MrOjq1+vkpV9kOHH/4htBYztuYvYJ2JshgLPPMnOSjPIygapv6r
LOcDe+Yxwzevf+3Gr6x/l/r55/vNkVU9NJCeKNtE8mo3kThkSPQXkHgT9rFvd3YOmE2oQk4UbC/q
UVaygt5dFL35X+SwM9Z6NQQi+y38woL+1NzfqstSy5S9Q4fz9Q1MC5NfrSXBvYt6STrtkz4ODPAK
f488zfShdf/g0WJc6MUsTEueNmRCdvb/Kh0j1F30s2j9UlKUYSwbRiFdaZkTAKzVptM7+jhRdKbS
sx5aLvXrUfYo6hJwo2aFN/RugY38eIhuhhH1WWudiLZvPl7ojf9fNJYDot/ChsNFstrNv4J3cA9r
QN0fQqwweIEaHFRvEqT82ZEjoDa078gTyO/lI+PkeC7RnvIcdW7qmM621NZ/dGNljdFLeiHQ9BBr
ey0OgOqjjuIEu5nkgg8ugfEc49EsQIUYsnBpBY0xKum390dJcRhbu3nbAZWEumZH4D0fpJzCcukv
zdS1OB/iteh6fw7nhvjnkGkOS0Afhgyso6K/WViIYoUdkj/tJU3GfxZtYtUsHaNrKEj7IotyfVtI
BLmjiOzl0Lz2J/eWudUw3tPA6ZADmhLhuqZQl5TFzL1qDkLCEzU/I4DEhGExI355Zcvn4LucyJIV
VCqPNZlpcrkT938TpZx2XIn/Vd0psQRd7Y7s69V1QadcHkVJHK/rlxEeBaGD1bgAGjzWmBlFEiQ9
mc+5bKs1bREJrOOliKud9oyKqWNk/+LxdU90Dh+DLIpM9I82kY6GsXFmrg5cggRs9/94UfHpvyRF
W/RZv8L3dxxFeWkv9BWG3dZuhCnmQpXiMMPNhAEOmJ4zJAKHUNrJJsUWabNUfXdZwma/2epR9L6F
5ioW2qAusnCEu87OSyT5C+m9db1k5fx5aJ5/XAJh55u+c1DKNRjT57zizYg6ZqkESs4S87jGEuV/
6sLVRus2XTK8xfv+rTfWhzhuGWrIVIpE079sYCxuC1yCHGNTHud/QQLMm4PCGfw4wi1901APX03o
JAVFsVoCVbAjjTZd2kQjRZgqWGucc3Dv2vcTzBqHoknBvhddedLFHP9isojD66PR9myLxwh5twJy
3mdUY5cyTiiCbqRHWUt4tPqk7Cei6ojOVUQPP3qNmOaZsU/NKA3k9Y3BZ82M+vmk/m+iR34walrW
uK6BHZiHP45h+mHqA10aRS17/qvzCOQoZY0jw515+IxPIoVyL/GqVZgiYS2cenI6717XCHHdG/Iy
MRL7PrdiHzCaEmIKASBBrKA183QiCdt1URg0iEo0pi81KfefHPT51rDPNg1Au5+6WDQPCFrtv+iU
lb8m/2ZTVzINR/G4vYQDYGtcpK8GvOU/l63ig4IfTm7uPJFDwCfVl45KatQ5gyFLEpfyNxfZdAbB
ZhSBUdtnEmSkBs9A5aafR5Eufce05wOA3etg8Abe9qhNwsCJ5QQeo1WUPK+9oQLzNYO0fpX11lqC
76UYhv5DTSSvT9d++xVOMURw9MRrvP1pTOWF8Wosc/tTi6zyoj7bAJnSqy8CAYKJOsyZnPyA2GOf
hmV8AM1WIZ3u9hcuH5CTwFkMr4JU6f0rc1bFyWFQjR5BfCHq500t0u5BFNJI9U7AH8l4+0updr29
mkSg5+7I7msOrNy+H62pnY0S71fW+uJLuq/5qkC62WKfHsxgRhgoT7Ho/ongMN/vZ/HoqbtU7fOY
ecA1c/WeQX3uW9MSZDwdug3iWJVpsU7IFA2skESm6R3I6UjuDQqP0tznB1ttv+xaU/5bpzVci198
H3cZGV6B7TKnO5ajhIgLThNj42qkZIKDvs06KLz1N4pJGCIt6KQQCQkAa02Ydg4dUJhonEtdw3i9
XexnGvdVbZB3Lcr7lbtBF4tREHnCOQ+6JCFUfd4IZ73EwJAVKr7HSVC9nqDQn92lUdKDj6G5Bp1L
zTjW2fCNfppdByJ1Gz99ew6d0bQmPsQdDkDtAR8ZQxMpK6L0IJteRr4FUjI+j8yUJn1mlJ3Sf/KF
56/yvlGGQ139ACFBEo2UO+gZUyt53WNpOFenO74zvS07AcY48Xb4soHrWlO8ZWG+dkYcSi7oBTp+
U2UZUwUha5zx7dabU3+SAEDocMPspcK1MCv97AAb1yNRNAX0ygJS5s8UwiAk/gxop+d4T3kGIqv5
Pd9q7+MDUPINoNTWwPphZbwUD2oF17+qVtBD+LDpLwxomLWsaJPjvS37y6D+JoR7PrKmhb3CfidY
hmWvnIaivt5cy0RR6jJXf9B7w8+G4rBTkg62827X5sk3Bbuq/xb8/yVXzcY9F/jNbTdkUSnQhhga
qZXyEDdcFjGXb+VVAuak4RlmFHKy6dFcVSy3Wk7qqMHi5ku/U/9EjjZ9Jxzns2FaTHbHzCWhvoHj
Ela6r6UMXhAvuCVoffxGATa0Y5EemWtM4WMbVovlHu0pJYa8UEvInkWc3qraLdNnw3g755RgGluX
uPpwfFNU3KwbcCnRUQEq/QHAC07rlvYJ3cW3tYkFh3G3EdB56St5Msl/l9xv41ud1TTJX67eRSTC
NDo/jCeR1AefiCRMGRApgF97VsLKJ5SQGrgVN/8+1pt9A+S/lClIjXa/Ch+me91NH7ie8ZCCJ0Tj
vZm6rAW8/CqsIMw0ma5ALLtFPO3JSIFTHm15EwAadX76KB+cs1LA8O50xs07jK9QIpRGUJ3tJgJw
KoaJljN/tG5Vh1fRsrCXrJ5AHYsXVW2y1FVLpKkkjvrYyf54yOGQjEASvPKidV2LYGz4uhWezxrZ
kCcaFGaflPNCGCXjuQ6MqlN8UIJtsxAa05U9ig6QiIBJK0J1XvjK+mkjSxr25NHuVUnn6g/BZipR
8YGMrwmic+K+D1pE4cKRlAxgcnEUDHbwV8tT7JUWlVtw11VDpxBtVSiSu66VGOvxUe0f5cNs6NXk
MfOH430Am/M4O3IautEbxEffbMmC9uwRgLL5rBpH2E4nCVvqdYm4BA7OLpBA7rW2Pb9lON+Ixf9r
EndnEAa7dt3BwUlgNNgSZj5u+ejnrxe+jz76Gpw5hQun4kVTb8Jl14RPSLm00TAj+gKjb5EG3B97
DH0MIY/3V9z9CcQKfZbqvi1dmw6HeAqtteomd6jT9zS0JGyuSPW8rQNiePUSRfLd4WGl8iGIKgkO
47brV2dLBVwriGIivkwGrvUV0vgUFrbkbMlddznhWOandLmF1fGx1p1P/j5lkOpvnwnRMLJiRE31
g/PHtdFuMcHfLkgwNmvOXuKjBcbe3lkzSaYW7KU3V3XS8fky8bGN213VmUcU/+RFrpaeiTw8CxXn
HJu02bzMxRORVNppzzghV1SLrMMAQkUDLr9WykGpd9nDpB0NIiUYeGqCsS0+LsDDTMx7LkRR5+Je
20r4rBW1IDwQSJP0zqGV9X6MhiSmmAj1H6Pf4rSM9Tk7O6dHAPdkaLDsSROmPKA8DwvbdmYFSQY2
2q0dPvx9VX5lAg70XXpqOMMRNd3L3hPc3Vru3ZaucoX+lOMpZiynwg8TYz6SSonXELE+b4qSeVJB
mJHmgxgKmZvi40mcrYU5RCh3rlEiKHVAHCTNO/P07fH+eZAl0u4sCb0Ij4wjAA7XvDjmtGL2Lqiz
kNe2h5/s74F8m/J4uF3b7rdKW6mc/T6naPHKfbBoijnzqdCytMrjDcL/+P0oNax5pl+Qtxtp/V/y
S+yqXRtEB9Z1wIg5U0fwU95MFUEzuAOYSfRbn4sVSo4UCuYns8L/dUNnm6iUOg+aPqSGOLJ9DsOw
kmahol6VZCEKoeP1iHIkL0lxLrJwdAzkZHZAbIrQwrQyEe1YJUAk4togs7T2BaHTjbaoc5eulcER
nm9jRj5IRrR4yOF6szOMCYr3ghrFW+dYBTcfysPdtJwfIk/5v/bd06Uwy02ED2eY3cCHcItvDsI0
pjN3K5n6wdazX8FKqKPfZ7Fm/yaGfi+1ozvPKVq8vpJTLKTNsIzchlW5Slxui9sQg2/pEsI3lA1M
Iv/TmuYAwiWh9RcKO6NP/pj/gofwMmgCn918mKxVMizaJIiEwSxJXL4WAw+ad217Y3AflJLdFQtn
y/xn/EYXXG/yKPdO+4TlSrFItPxK6Fj6SnZ4hFYgxm2cAvnmJGDUP26H27D22GIJd4hTdoXVveAE
GmUAT+/6J4iL2ccqgth+UW+msZjmqJ78ZOwVuFTpFOJlgZcpeZLVdftno3kjZa7kl0+1XNNuGQyB
YRt9EoISKbc0ilDs2q2ea4HBYHgaJ7Quctu0m2+/akItobTRZX3QaA8DnD8uFQgadIsY9tNlJlxl
jEkZu5LN6C7opEl0TNfgNAv5JJ2UiYvpmNeI85TBRHKt56hzvOpIxszTimlct8zRVcOgn9up+vBY
6aGBIJNtg+4W/VgKSlto1ZjJ0r32zGGTPPDhNdrhJU543/KjR69wU9CeiGMqdF+Mlc2huU9yPTSx
qO3CxjiPPViwtjqqNSlQlynkpyessUzxy1Fg171PrVofvapJliDaEITq2MZ56gNYcWd4RyLt+Mfo
ghGR/XExa5q5gzLeO80LiXVrrw1o9iwY8dhImDnNQ8Njt1T8Dt7wWGgxavcOEkh/RKOzMtmy731i
OG+pHiURcM6bGGufif2l4bWP2pkMl0bH1qf2qWwzopOBiEkYS9m5RJnGIVeVaq+AgkOc+RH6e9ER
NoDmlGj9lanMdDY3dO1vUb8HwrYmctYN0XMJTXzNKBs5n1nwqCyHTzOMEiQjkTSHgn8j/uv8xYEX
ibzleWQuCwux0va8VUzqQum/wW2fvCIXE5GMHi+VcOniT3cmJGJr/zV8xlaOqSW+TBGJYC59dsR+
CRj2BugudKi4dflChudhHJOmG3u2msfvYGck7fN63R0r7sP1OTlhkdlLCpQ7iXuUI5jiaaqvvBe/
sdNc4VNXYDgMqy638x1U89y9B6iq2ydHOl0nS579w9pItdcpsClEy636el+ZVD9ztBj+/uQAW20m
rt6ozbX9ljE7J/TQR3KpIQBVNsHClIwF2xME3Oex/p4Lt52wjtf15kVgMzsrCpRy02fa8DXyYZaE
Os7LNmVjAY4wpyGeslTS7NqKBv9XKN4shlnbUE7SgfsbWVYTiT5WT4gvvOsbGJsklKA8VqpG2s/Z
3i/CDYpWKH5/v508rVTdE5fWvM1BSKR6CbIyyVxvmsL9q/gRZ8i56Ym0NgolAY8vH9If4AXBZ9If
uHkIQ1e/cfI1e0HozpzMJzKyJdwxTZ+mR4yhLiLZKiPCu53OQ8QYAJQGq9qu9nJHzKtCSajnXRK/
Ayxma2zJKoE0WwG1AL6tRFrnFYwxA8klNI2G8/UQ3Mz8dZSA/0Vn+t86FfBPvbFC9TKdEnwyjWvX
JT9PXTVSpOZ45QiDPj3pgc4/xBz/w882oCRDGN26iFqVXjgDHra4w4R6WvLTniUugAPEGVRxPbB0
axQ0nGhq6QZ+Mp800nfd/u5q8cRKCXUTghTWJ7Za8JbsazOBzcopNa7xMicC3yqcpyyNmY1EgTBC
t7vkTRHA6+xUAirUJJN5gYdVSlM/WHximQ5wiWhTn9siK15tZfWBb6+d4i5Y9Gn3zg8TCBTxHQgb
uYk0WjpiRSNbDPMQtRInAvweB5YBCkqhAsLikVsSw6zUQNnZzAO1zREvm1FneOx/KjaZSLyCEQfJ
RE7mBV3fg7iZCX7WGrLJ8dUPgcDpLczolXqqvxqjMvqRE7Obo/crrXZlOaafKgSTpSrDjqbMApzO
6lQhszbCgWiUiWtJGI/wPaf5BZJlhC/drk73fcklAtX97/w37M8IEdDPAUvAcdAvVdPIAagFVRY3
OrXM9NhPurXPANVioOha5rLRykWgjl4P0YyzMT8sVqRy2AEMKDXGk3iirv/1sk5uY41hb0WebnDd
7uCypAcxo4nc75Jt+Ou3FcOepfcDj8IVIGO2Zsu1D31jJoP0hLnMc1fS3b6MvjyuNFeDWuOU9sdq
6DlzHzxLjKkrMGQT7C5qgc/YkUXIty0IcZkHknxUdeo9ZydBiG4zX+416k4aDSwRxXkd5UlL5fSs
dUBGcJsTjjFkzV5KZBuYWH7axjonuNhVS0PhlS+6xI2RmkZXn2NM1MRqOdvgcKBkgZvlE9gh1Pu6
cU+0sv2SrNV+c0xO283gj/B78wjZJX4tHL03KdiPgZIkNkHkn1GBDYzN3ZvtxZIukgA6eP4Mmlx0
e3RqXlAAeCjVOut/KlGYrBxyfu4y4VMKXL5QUBv5ehcPv1cUpupyZuQ7V3YLGvtiJgeqH8LvMCib
xdL4uFuvZY9Z8tUv9WyIDlnK57xxwjJ/jXjk/bnbqlrbHXImM8jIVqz1V3QLp69/CfcqX3u6i8dW
7xeARYCsxyuP7lEra2sIqIodEwE4VHOjqZw5iR7iKoVIjYA9mqgwRfIsCllZQM6IzPB3yWP/SNnH
VqT3iD5Mczy8il8frTVeXDorq/A/C+ZIW9GGPPWy1O3Jd6b94gJi6SpQ366IFRNvy5abK4bgKUvu
7HIsMzLOp/+nDrXO27fCOs3IbH5GFFOo1NgHJCIfSPijheFDNSkiyCBGtkRTxDeXLM7VGUIdoJlI
zga/LPV8f/ULkd0TICbKcb8DcdAJcDcW4k+W0xStCAAzMWxhW4KJJtHreeuyWvt3FB7Cs0A9+wyw
Zu/v4V1C+QT/zJQVRVbIzxzRKs9XNdGA7KYLY14XxzfbWir5QpQf1CgoAHtwYC9c/VzhvJco/7vE
BOmdPWl+439BInT8gamu8ooqrsr6RD1TcBTxnQjc4JyTsVHIbC7UwYNSuveyq9JgKubWPKTxnXBo
TKyVoqZyPLCb7TWzxxC9wb6t+y/kYqimWaJAAf8u0lJLVwimrfL92Qa9x6xlLR64Cq0IHtsEhGYI
oWVViC9hL/QLGEg3XFEornhhARTarNwo2Z4p2SOPXlX8ZF0dCRZUqMh8De/9iH3V13uqTbH4dIr2
MQ8fIWEd+aLq0s7+bkSBd3IbjMBrkCneAUwsqLRH8kWoIo07YPF2OZY/WKmWEENWf2fmLajlwW9B
mdSknY1w4rlsdqMR/vXPIy+UMEmroqjkyOIOLB+XHhh/oiinPNi0zzOPe7v0WPwb8z37y5bgCzUr
k48hlBzFhOHnZ4/t/+ueHZ1SfAHLenjB05tLkK0MQ4DEBLBkzEiuTi5E+lYuuPZ1Q3LMCwMM+C74
ZH/ObhSaUiPiqtOr6MmlegSsqAJQoVRx5gz0OUNcbSMIrmKiJdEs9UvC2sLqLBtgUNvhjgsIC9Ne
9lgWFBfdTttIePjcQP6UecZQfRy0Us7d7WpZjPDAGmSGzycJfMS0rjI7+r42OTlsQrHPBbQAZ01O
+EsN3BL82Q0lk3+Qwfa6QUBnacdMPbdqS6aL2P1dlCh5pZ8EhuhUQTXkRgAez2H6auyyGZDe1xDx
5z4ume6jIYXC0lM0OS7rdq0UKc3VlrtWOm31ihveZvvB8KzYBYf9qZJmIYsvSqOuw9Q7cRjkg/JA
TulLe0H1VnwpynfaZEMIRn6DiWdez8G6KFJJXoSh5PssGrYI+oTywSkhLw9GvWE4bybvMQV0xHHt
uMsm3EOLgjhP8xL3A5xssQ/cctQrdZaQ9EQRO1OqeEsW3GNFeQ0Us+1+TSkEvf0A2WNOVsLf12aT
0uQh3o9CtwE8w14dtfwzpxor/9He7VVkwwAe8exv0I+4TFT2Q69ABukqAlu8FNaRrWMmIGZ0TqMB
zUnkqU/2BctOv7W/Bn17q9YD3M1RA+OUHGkkYtFOhs+hi/JDi9dJGZsghbOGMoDvm7ulvuOgJyh2
3sr+MO72dl+SlwHmf/dWcJnBQfmwZxJpil1mhcLm/aR2/PX6AKwAXUfL1RflU8Nv2oai9dRVA9g9
ska2R2YRgPHnJIgJD6geVIdlJK2JNsh3P0H/4MuMosZep1zpk9gQR5mdQtfHjo8Pob6irfOzXtS7
ZWm3h1fhgPd31DlohIYsAZ3uQPNvcxmiF9GbLIFkurcj7f/4ESdSDSF6ZD3oF8vFHn1LEzWwnHJC
52qi9PE986waaKrFsoIPhoBFk7pGSEjIphSrD+7xJeQk/nk1lnEt8dbbjFANgz87R5/8o4jIdZYT
96bgMGKxKafs5iU5w+s7vV7WcHbAgIm7RhU1qkDijgHL34W2KBB1BII+2JYh79y2gsufXZKzh5zx
LkiJHzZ0i3X7xqENDvt+U8bxzsqmrI1HAuTvzp2WNBPLWJcd/ry3m4PyZGpeW+sYfRM+eeLNI5Xs
1W+ML7rMNGbUlXnDlWd0cX9hbPsKrDXhaK8jLwOlReK7Q6HHJBl5+3cxz0SH8ZzS/8c8STfeU2/e
GKcAMFfb6/9/2NaomDGyI/j7PbAiS4tTCNgizjSVpdYwZ2O1y+3zIo+HNwQOYRE38EOf61yG/tcl
7sy0xgI1ekJ6DLT5FdYMUy7ktKkQ6oOe6OBxMlNqC8GqoYXWOZDctxS6sJgX6V7VOomO51moolzG
ncvp3CtIpdAoEJ+Kzl45lfoEGlHFbRlcLbEfwhxtoUhaBJF3xfLvNo3rSEkR74/jX+I5JZjAh2TD
dUBa4GdT7qLjcSTklgej1KVtUlHpkAmdhm7QFdMUgh7+4VvuyofdXw9w7DxBXyLkBw9Dj1GYpxqh
fD6m6uQd1sAnoxcQtGc5EMlo4fDHwP+1eLwscF8viIOQ1qPfF5DnWdW0JZNU42QUCm6ujdb14G+S
kfRk+fDNyuNkfiZTbVY0+iyNVrm1n7zx5GDjiNtQO80CItTHY1Y77mnP9k/u3GhnrU6pxHCgiq8U
DHQSRfJpnWJY9DwdbQ7kL1OH8rwh/qpCh/lNQcrq/ljRngFz0PPNLFYgTgBi8ogHOzQ7rY0aY9gN
EyQkmi3zVpOsDsMTEhERa2LcPZ4s7/lW3jITMAgHDM7YHlw+dpUZ/BT3QtPOZAfFWdKxeB3ozrwM
DXL/e1YR6Zqqe4gaWvkFwLmSs2eSx/xLlvwahpom/X5AljrMCvWyLlFIA5Pu/KyZzy79oNYA/6yB
XqPvhbe/VfUN2aCxd3iguhrG38tjEzJbNunSxvPGVpNJnt/vahJP/c49lOS5G4g8IrYjgJL9DEjc
MuqKadpasuDL/leLbuypNzBQRn4L50Mivvzqzo6VqKGefWiCQ/0Pwhyive3p+A6dgC/xaUGgNh3o
6h92+oTnGvzEdlJbnZoslZIWQkEqyIS0RU429T65yud8E4rb0dLXIls88Tqt0yRLslV+EDf7wz8l
dU1klRZzgpbENXW9ny6DITBf+J8VYxEJwcfDnmBZD/46DI4LMW3/WXZNhrQ+REBhQg9hwdZD0OT5
b+zvZDDdzheQDtDZ83aKWVhBSm6xthtn6zhwxijYP8gaUrfwMbluijNxNxteS/X7ENQs+wKWEgyl
iYR9TWod4nTC3gzuOsj6ZRK2zgZi3V3ZK3M7R2+IuZCl8WsVVVscRCGRzRRKAoOLTPiI/OPpOD6m
LF/aGjH2MvjlO+A/syuJ+YJlB3tzqV5PyFzaHw8ekXZLBaRLkdBQ83sQxJ8A9ov13OxCTRWQW3Wo
ifa3pLjlfKf/WUDIgy23QwKcFiR9FKIa1S4mmBaKNR2lnjxhWqoTdnA6VHHYmRvff/3QrCqxmKpG
CZebgfU3ZxZ8pcTftKZh5sazswy802fb+k2JHHT46g6cOdEJBGlHIRwd9JXXtDhN/smWBNN/nx3b
ZQ9m2CtaFFv5arrKZRlnRmlb/Pgjfh0lYaS2tXc6kDMsauLY4zIhYffCjE2rRD/9BYIcZG9EQ1dd
biOOHkl0ruUHUXi19x7REfKqGXmKrrCaDctmVcAVsePHhknCF6zuKypgszYLkuyB2cg6yEIo2l8e
4CDsuhDZPPt2VwVo8/WMi1yFgpnVA5MzAVexm7B87bv9Ye3KCI5+nmJigUm1vbqDIJJvlYH2su98
APa7OPP9h2hPXrNndLF5EOezGbF2p3SQmvVBuE8SelQgkgoY3YTfZOn3YwVLs3J8T34BnWELNuwm
10a8c9CNsMqZbdXkNviXhKxav7NBQcF+kAOvWe7rzBHBWBkqQTZhc5CRLJaYpSLcO1l6Lz2O8ZuT
PcR55Sxy5tb0gaR/t0aAuOeobOGo8RSYvAUai81t8xv5iNbqfxpB9tGNCQ9MLHf6yemTHeWtKLQf
/2l8CZ0tWx1Xqav6VlEyGdRIelVsknqLMVmoV5lOPb+cC7PG7zxSVoj513EwwFmgbEKt9a9nHP1e
2F4LeizSk6AFNwylq1V8H1Ky5WvWJAK2lsufeyNev9+sAyff3l04z4eisHgFdE2h4eYHithKei2K
ET8i7ZHm2DsCqrqXt7GZSfrUns9I8mHu03+HuTVOr1+p/C//lxwQeCGmfOLHU/BZzaLjodx0GTUx
RA3oszSXMlLSJo6i/Y6dM00AFhL0rS5wBOwgnUR264czwKoKHvHBGW4GnVcGVjS6PycMNZMQr9kz
3LSSYEYIAWsqA7UGeukIJcrAsFjcvHaW/iGyIC7xe8C0QFewh+tyG8nKqeNMf+uEd1yYJricBZNZ
2YJkY42UcfyAQ60/uMxyaJOOMc9hB0VBfuxFdZaG4hlPLEOE99e0IAv+3rQPA5wpbOovFXMvOFsZ
f6TS9L2Mogh/+Q02tY0v17aof98lK3HrjU8nfgXAZguf8mPhffkF1hpvL7ZQ8GPA6aD1JPNm1Vpa
Kb8p5rj6mecHJn7XVDicFZmWg/pVUk/mHsEkd8jvqr1QMymcPBcOxL5mfV5yF8IKigFGgAXwV9//
uMbwGfldIUX3gIytXTL8WWlHt4oJ1Vkeong03+XIsJNW3GRKvauDwCR/OklO2QYotfxdfRF1PRrC
yw82vgupEz1jYJl0Wor34ORF2fLIe8y0PhCr5oXJFTRvrW0KeVxvnHuwOnip3z1xROe5sLRijwsq
i4EbBHbXJYgjgbtpqnRGEzWBio/4TLtH/XP+fK92VC5nu1leL1ZRPK/XGYO7Q7qPDm403o/2UUeh
dXiIjN90WvXszu4ZCPAeXW6aIllBw3uCRWkJsqIIJcgNQfWf1ijAzPxHhXuhQesad6H1/rX+jP1d
e+c3tU87fMw7m3zpDSGad8mOanMKDgEeXJ7wC3XXLGzFu5qUGsyOn5DSW9GRl0F8CbPdLcUjU5DP
HC+5+Nij71Hh3Ek7QQR9vXcPfwL6SSDZoLIe/NkGE7YvIrzOZvzGD/pXzSyYXf/QTEkpHjcz1IZ7
xseGX8A48FhxS/YK5rGODus8T2QND4g1MXPJCXaS7HnbKPfAjxRcfWRYnyS43854tXrPjhOApCRu
VeN0iZ2MZRlShAhoMty2NpZJuqZ4wtEUXeOTFMwFnbsZSqb+AvQPGddw7XBnnU+RvwG/+TIyNiW+
uLr9+yMinlZFrz6NgVrbDyf7+S2jNWNKP9bfFyxTwKGCgnUerDcgz3MKb09VncjQt550+KOqw08X
Xpj/W66UGWHaqGVG8qhFWLFzM0Kp61tIBQNvRw8X2cxgr/m14QX3xLvwpDtovVYG+WMPWGogryGw
+nF5pOAHGm4NnObu5J0gxCGQyMytxX3SEKegXwKBQmHxnZetIBi/lc93S7lP/4nOD4O2zfy6xxnV
nvb/lt+gShF/ajm+QsdwbZs9MDLlB0vcyzn7S87dDfMAztWauywDCjfjD945BXI+TU1I8oglvsMi
g6p3fWcaLgioXKYVtepEvBbVyzr94l0PGCuaCPGpKVonoHirfW4bkpK4iXU4JXLUI6CNwBEtoUP3
iYbVsPcmVqZ6kGMwTaAACx4kgg+MplURV7KHWJhchBHUNQNcbLj5g1THO4NzRVfREOt0GhVokKqG
nhDo17UB0eCv/Tp3w7ZRFvAXOMXxIQkWVk/w13OppEPpZNYog4gaymTtKW9TJcgZYWw++H3n5kUO
HJZCY6RERDklDVTO2Vr/SCH7mdr4kbghTPBu0MmwH0dLFXpR5jB1T3LB6cJ3G0B/i9YKGKkrLgyC
LJmzRcc6sNvN19lrObF3LEwNWkJ/txJLSNFny+D+8UL/Cd+y1lyejXfYjmLJxVIYuv3RucjRbhoU
U/jHBely4MPjYeB0KKZwgDiGG7AnoydY0kJioIx3eFTqnFxn8+usasrCa9FpBaaLUp1CS1Nm+5xR
ofR1Y+evXu3SOhzcz54AQxhDLWu9795xxN7JhYQAl4UDpm1DtY6ZqzHOflIq73XeaIcQe/O7V/D+
lr9xDLrI0frKYx5VTlsTb/PKpZLkcpR7c41YdhuYHeKd3qhjmkI7UIqKxJoLyU3xhsRdmHZbZysN
sn6+cyH0SQt/S+xeqwrjARQd7FIOOgrkt1t55S/WUY3cWdE0mQ0vWBv+pTjmKJ1dB8oLMwmXB4rR
eSP6K8pjThz+ynee/mBgvyYX8ogbB7haRX+Cx8WkerSwX6XVQNd6hpA+TiPFdKKMmJ0I3JmzWYun
9FQhd38b6boUZ0BRhx3YdfIqAleVgmYcaFmLMvqKooUpG0d4p3ikATWzMFwQBnvmOLFy74Io64sn
IMj6l1IJH2Ij4KU9KmdYSRZffGCNpD7crC3LDumIXhZkP6sNqUZyqvLyYsmSIVi6svw9354p9sYT
Y3thwcSXwltYaaxkMk17tmeBS9H3TOUMbDxNnHVaithycfhAztVoQHVTjMldTQf9qeQPT8IX3e6C
FGCIBiMDMeOylHrbcsHyij5xyav/hMvTgPA2d4yF/mwUALmhVyukegviPuveuuCwQG63vz0ZVbAu
d9u5vP6xx1U03GbAWEIwdWGCUMzPDIMOwjuVmmJHIQxGYq45duSAFyjBQTbnQt0rldeCaO0iaPCY
x+dcye/2stbd3izNYh3F1ByhLWB6LC92V07JmEIvcMN5oJvIAfDRIzLrvyQnot+9C5dtofZHw82r
4bgKLad6F8OVo8VSdpSnH2tF4SFeyKsj674JLr5WJAftrOqRaF6yz7zESb2xzFlg0tS2ONA84Dmf
dttUAiQ4SKNT30xpITb2+4jbp2IwubNxDwkKL95+y5/qIVTBD1P13WCcEM1kynhu99w5PAcxud8+
+QlaDRJ5VXMh98mcPYEVHNrbemN8bsPws39CiXo8b6p/6bKBA8OufJH6ZDJOCVDLuvJgcnqKHpZG
LbNDggDcsa2TIVUPVjFAV3xaJsDg/Sg6XfGqZ4wwi/2PoCp0CkSm61lANlRwbKsN8Jk0UOymzejg
s5ePltDQ+gmuUTKIgz4gYc87jO9w6ZeIf2ZgZaSJLovW6iJ7TpaCagsP7qXMkGB2ZxEZk3FWxmUp
dvD8v32Ddn03+PpW038RHku+oi1tISTYADt3mK+Yo0g5nsl4pU0+D9Z2u78pzkBDf+9PqefXDDy0
iNIXDhNQXS2CGYlNK7vzN+oc6JjW8ZwvROMaAK3xBql5MM/sVvWuEpog0+NTjmFstRraNVpgyVYN
wmjqtrqUIlAgI62mhdsUUnZ+0u9FhgFS7xP9+UhHM1FDgev+bQJEF9kYaOaYSsupoV0MLh9vg5ft
jGjF42ScJJ2uyhCavc/M5rVqFpv4RXNxefmpF1rw63IDQlaWzUhfqHt1E4d7hnsErR1WjiOICafh
shwtZAYTtlYFstyDDxF366E+lcRAeWIA0mqG9v5ZG2WnHt5mtRu6lm8TpvlEmsOQDI2zoN+Rc+C7
0QXR+HBbuC/OJqzrGRBl002fcZdf77Ca8hC2avTUGllXHGkJ2iss2xvGsJSAdBIbDU7rnXzf4Lfu
ILpAurEwwEhM5Gb5j4ueFXIjgwoprYzzUkWp9XgtJiht0rwtz9T2I0/R0cRkx8VFg6FN14tJ6fXf
A3uIyOiIDn4VJKlClqfq3/LuVI9ZduvwwY0lYysJ3qNb//Mr6XQU0NFEHuGw7wGqJmmh69f7G2Xz
DpDYZL6fmqMB4ZOOn7+5+Rc6FHXY9/hZIO78XkXHS6wVuATrL3SXEjkKnNr5p8SqTo6BeDByQBsi
ixeea0WT9rlIx0tAHZZ8MFbP2oaSJw+e1lwutD5nKQr/HnV0qx3zE85Ilncp/4wt9UlxTWGuO/2J
NpYAJX7U4ydlYSms+oCFGdMMBYIFHwVCIJqfCo8+4lJqZfGib5c79Xj62UPn7YiM8WlH/HyenFtk
0gFlgq4vUkF8Lx88WwPVB6YWcGWTvKnE+Hn7QxVv1/WySICU+uExymkGjz50mUevFQahes05IMgF
OCwIGIlZj3JJq8hAPLGzJD9Hwo7YKw17sg6ym45Sy94bffq6qes5Lvg76qYyFoWfRfRVzJb9MhXs
LtHiexjeTJAJ1N8gx0f7J+w9iwLbppEVkeMtiJ2fP/4nUpLiwUseE2cISHkunUZ6Wh1CPZW5JyV4
GtNCSo4bNM3Ww8YV6RV71rYnPRalj6slosDTw1cLZjM7szcIlY8AUZCH0gfZ4i0a9VcHw7N3xsQo
1HgM3f3FJ2jl8ZxrhOH2nSyyE+9PnNJsBONUhBGxuUU00wHOVTQmlk/DWHzQ9/zfesJdUo+T53Kx
MyYO3omJb9myMbmX992QGKV4obe8wTjTxGJ7Uv/aPI2ZJo8PMHYFog16TEeBrNS4lqnlcniWxSRK
wLgU+74wrLg4cTePO9WVhAQw7jJgJYe+20l0fGbFafwV0rMVaID9PZIFmq9tMzLQo1sVOE+lxOgo
A1ORQz5Lux4QzZ4mu0VeHahe2QXqc0sq9sSzND3xgBZJRyi0Jym+nd+rX1rbnJ3wg25RS8LZ+aLK
n0Bf6iWCPtETolpHj/6UcyR+R/Sux5+GUnbw/cTgGrXl6YhbedU51SBsPgtchUcX2oAFEvRrnF7Q
IQJrOxU/Mr4VyeL2IPhnkekCUKbJ+7bZNWKmBWG0NJeAjCQS0INFj6l82KrkUxfqWhj+ndqioNhi
u404RDjs909e6Z8fIsttoe7gTqT2kIhFj+CXuERB/rDN2O2+4JipUP8qO4g4lrIH+56Jzf5c0Z74
drIWhVmUqx5bxnLclsLJdflCVxcewJyBNrhorg725KjZWK/EInLu9kYeaWTRg07PjArm01VwkiOT
O07PwPxjbNY4CiBBuinbeCHXdmqYuUyeFyzWyuysy8rxrxUw9Nm0kptUDnkPwWdUdVlonde4PoWl
gXjoYhLKc+SWIDGDg6P4uk6XXodFM3uHj2SUi1SfFyUWvFE2SLupa7lsdlff+VxBA3dHqoFrVy0X
ZG3CByv2JHzI+hGDfYyRaxmzMP2TG7Ag4nlCE5xynNeBCIHetaVb7l2+LyBTToCxGlJnDd5ZJt4Q
JpNSGym0YUlux3NfT4UZ3uaDs9SikFahSdLh9Bcous3TUOFftStbdRC4SLO35gFZEtGaZl+37TPc
qee7MzjXqrtEySYdb7rNFdCdYE6IMaRJCtd6mayZy2UQoq3Cl8QJkfLgay945JhYQTrHkAWf7QEx
nEWxfr6QGKdTOL2CByl2/Qc0oy2kI9vzNsqyC6WfMBT4VF4iCmJB/b2GELx9GlDnYzN/vYNVnVwX
k8Peh94OLEzsJ1u76aJ/3cRonLt1WvC+LmdttglpSvM/KG+R5ZQX433pccMkXN6/uwD/uw/8LeUr
Vbjoql/ZRojNa76atBtLEBXbJTU8edGJ/CeOT4+LBLyV4cf4PYsbDDWvrjZWwqXzsupqE0LZA6TI
A3C/LnRaB3HOvfYDdWIIMlRc//UTlfzOtB/5Dw2CkZTRXUsOqWUGnbtbtO0cWU9VdzQrznZbZ6+g
5mKLizlMKGpBnMmdbbZntp1KF4OPE1w67jO+RKjcT6Pwga+eWBoyvGgSvFWO2xgOV8WdyMNG1rpF
RBRP/L5mUTF0VGzaxew81FGFheRqLftijOnhivRQ8yti/ytQmmKUNH4eCkaLaqtKWMY+EqK8M6yY
CtGD5go0B4z1+og+KEUGRxjo/O60RZU6wGocQ0d2lYIy7W3NCJ1768bHdMEYYQhq9xQG9cGY8hDy
TTAakzTw7ZUFvuvGPzIG1SUV5eyLqnbdGtzeW8yEQGpV8bMq3PCABxCRMbi+GqPtTUF9atJXJuYq
8N+IQ3fS+Rrt19Ls8VpKu3PCrAZs6tAjn75+bqZvOysuTG7qufXSW81Hl2Ivr9UBH7uvIBj2+vCY
X6abhJxTTjHMEeCrPxwgnHHLNcdQYTPxq5EUbkKZ6kjvv2InwHQDXXh5PAEEdXE7nE8FS5vHgn7E
HFFtPt5NsfZrDInAh5m1yk95uEiPx4Zj0AVjzOmdiajzD9mrXsKWVZJphcMaJIVckCHMkB+kY1Y3
xJImLF/3aHyIMP7FYyV2RYmmEoKJiAkGjnEY1z7AgjY3gQAHEbujlAQOwP9JAL7uvf9+8G/2rzZp
0ZcCIQwxflrOu7fMI5ENXDmCUAZcO84ITKL7+zqg2G58LuJNtzzVu/LM0oWoO6LRyyzykxRI13m6
5sSlKMTkChiUXtFSAvprU29HLlYxphgGexF5Sa+id0Aw1yD8qrUDBcpHyqfM7CnIApNEwiNwbJe7
bYtAgu9SeIhYqq1kaC4G93fYp6Si5rSFRKLGXCPKLFQQzemvdeXYsuXwrBSs7OiVyfWpU5poNPFV
CdVNW4E5nMK94nUZCt7rMOjasrwuP+AiHOBL3X/fvCoZHh30UTYw+Df/HjjpsMUp++mPOVILZmaf
i0IIvVZC9a23vfIxVLCe+/uYO+lWXLndLFJfVv8q9hZIJrJnnxK5YrOYudHDML4MKb4tFdeyFzvQ
VCPI77nxNEO1lPuNTVdc23xYBUrs6wHolEYl+CZQzN4WRPPCqrfND9GrChgM/dJ+Uh7geqhRsp+y
YylJbQEPJmePnFb214POMmx3ZEj2uxH+H7zrnZkiff2wzBbevEm2c6IewxVdyK3463LBEqQwttYg
OL5JwNrUSeQY+8fOCveu5U39RZaLsRBZopuQpz5ZivtwcoiY1WAI8L1Vi1uvh0hQCdxotY1XhAQv
4xe//NO01v7PLXGnfRizxgSQb6gDQOfKL5jK+E6elQ3Z7LOlnkkM8LZHn1l0Bt6mJq7sINpHzbSu
RrvwmhsrbcGcE+fkBqxzufETYl4ZS6bCTL/XO0UyYQBlSuCqwEytZ/tZLsoXqRV8n8YpFtMYEF0X
hoHNt773I/n4xFySQGvkstgq2PWDhocLudVhaNIFmghrgl2lyHfXQG2wgZVnUp+Mw8f+Ur556yWK
BtUe3lh1od9mfsJuNrehRLrDM4PKIX+jy1fWcW9qbXeqeTpT64ETXMSHJkd15WdAMIx6gHGTSOat
kcI/qXdigl4LONKfk2D8cJ+6MP18E7PEno3tONRAr4DIOvy9CztaSgg+zZ2AyGXtcGrJftLKuzAZ
uwv80jm8PVJxAVogrjbqvr1xBXxwi2vI67z/gD50kVipyum0fSkARVfgmzGA7hfyEhGbb5iKdJJ1
SNlPp0s1ZpDnR75lx7PpcUIsF8oL1Z4cR9wWu6qm5nAI/U5b3jmWps78bHxAUh7QUb1mhJpLHp32
GPQwxzz5HrwfSJTrTQuD8xTfQuGU43VOImPePHuJVi2O3M5ojPXRnd1sbG1Yj45iQUSi5G5XOpYe
PZeKqsU5nxLqQGlgAn/8+ZnpnDQfzX9llBGKNad/tISf53oVvuHIkkkVUOhkcdROWIJ2T2GN8tLL
qIbpNXKvDCRNjwXJyLVg/D+Fxw3j+PJ9uwUAQoKxJ3p0obq8hnF5Jtp4re+We+9XcKr437ktDrZk
ofvxqCFFtSNdGAMxgGdv19C4ZQaPxzdf/TwgOp1h7b5HQOZNwqorwrOVImmF3EbT34eeyP4SmiNg
QyJ4rEdjrQWTBiMVuZgBj++u6PvXCeru/tlfKqqlq79y6iYg8oarOUg+qZgpSYMHaPCzL18ReEDh
GTjbFIwmpYk3g8cUC+2998nxg+E8YUshODBQQ0yYrodrbNn5/gGLY7WzEqn8BRDnRMgm2x9Oulr2
txdb6GjrGsTAB9xDNzQe0GeX+k8kImYpz/DLapqyhNHnAN7E/1/XllIQVz6Oh06X9s64ru2pC8rn
bMrnvYXqOxddar8Jl9nYq/NU3DOyPPgFazldPh3jlBNOd2ZS+o5qZND4XlkZe0uN652KNI6nLux9
AZDtC370qIf6+3P0GKXXcmro5fqV5PpZjYHaZzDFMnhP0nH3ptaSdzmhiKEH4lzgI/AeFLijmHDd
xG8bf09Rt6oY1ISSep7QFLH3BdbpVPXVyBRQbWV8Mby22uozvXSDRPB9G1KM9kVLCK8VNCBrhm7/
gkkUNtKne2PgMAdHkXDfuUhKtLbhDyKI/o0bdJi6q6XdIr+rtzIm9G+oJCJAHBrS7y4fbde0H/X3
J23QRDw9rQ6DaoosGsX/7T63Ri9UVHAwhfc0vwcz3Por02rfcL/jI8OmKJO3hwb56/K90mkANoyy
hg0GzNfYI0dQDnAezOZeV0xNZ2E73mTxm4dfZ6cQy3Om0GWcMZdLlQv3qYQw7mY3tSLtOfWK7LXx
TOKsyQe9MqNBNTmc6WyuE3cFSAVSQ9bCLpgC5wwrFUpwRSoPnh3k7n8XghwBIZ6VH8HnP5lhbtLZ
6It7BXDZdWpy2NICuSQVXOfqcds+WiiBxnwChNMClFRsuasjrwDKDc6aIbuDkOE59lmA7oRkrIK1
IUfZbSykrK0JQXElD/IU2Iq7TtrDHL9o6ZRBmUceMWFnL9rS6s2//4xwaoGKeEj9EaG4Q52XDsu6
ZGXsDxki9RVtlwaP6k9izDymeRSmDDD6ZtT4Hzs4DaP+xImrSgG/4TZzH0GF4jVeQNxM8Y+tmzMf
JxDmyM6K//kFtHIjwJ+NqUBevoeXIS5QimK2xswu0lnQSxcpr1wRUUqCGJR9aYK3egkLdEaTaJ0x
lNaSI+N/OVmxoDLqeFG22xHxqu0cu0yZAQpdAnLmjXBQKa/J9MipJM6tZ4TSrgChBSr6iOQrKZ9B
afoWqiWXaPoTuUgW6TUNzQEHpUTtSRv2q56xIO4D+9/R6SGRDjMKdSR2Vr5OurMgQO3FbwegFIYv
k5jaqKzfjCbp5eCFVIEa4zMn28PzB5nARKn5CK1HjdwXh1QbHCyJ8c+k5liBZ1+g41ZO5K1pGl6J
La+G2e7/hsmasQ32z/i67bNemKizB+mZV9oRKIVfXGE3AvQoqxg7ObNPHA5lvwzKMEMs3kKmUd/u
CnrCYvwDi2+op7iR6Wsh/U6tImAsdvSaloXm3U1uiXxjTIwi96M5FwmRkaC7CwYMNBmcbzm5ILRK
f1QxOkJU06poGKK5l6499hRTmIvwrRcxeKcATJF0b7pVwx1nKVxlzPHMOPCIWMEgC0q6hhHXDi+1
Qe/RAD1LEsV/4GmQwMXrR+bBZ5oayvlaDOqH6w9sPNdIbY/hER4VY6kwjw74/HdhOs2+YR7jfcug
62tke788K5ZC3wVnl4s/dbNEvazd5EuFf1RewNRDnL1jtl/QKyE7OC0EQayNXr2aP9WPyzP+CDvN
cNd05I3Py6XfplpUoqQ2hkKuJ+cuSd7RLmhoi8PdgLuzOUzyo42ank8PFnxF5czTg5xUyAqkkZV6
Pq2HXOinH2EGWoTsVsu1Ic+iBnLpCd6lkXmLw+Dr9thc+zjhe4+643Wccea1bX/yH4zJpdElbcc/
PVLeEx7XdYr/Aewq5w7XV08EpBsnmQzjv4nnUI9YWyEDHq/NjvElGTdWPWbGHc6wIew5lo1ONcDf
Tc0BHYt9nHwOcyc0xB01rXh6ZZVMisyHComSyVwX11S+tEdr+p4Rb80Wj+NhnyCFRoAnzbogAOpI
fWiehq2ks457P7adLLwIUTcAieDyXly4gD781hcA2DM6WGorrH0SmfY0Ta9bFaEDL1fgyj05LcPc
hpwAZq5HbdepxCSF8LouZPsKOT2H6KrIM/2sUxxZFYj9ac+1n+iBYpS9P5yWu675uK8q5tC7RLlj
z3XdtaSEnsxWQ0xPfp/DHOMPxwLAMkCE10XLsfgUoHUm/smnaf5cruMEuZ1KiSENsbRjqFLqTV1v
AD01I2fjF4efakqwkj6uFv950oRDJnx7u50WaiAUQPFborFgqllJKCEOvVjnLIUC1cy/MUqP+SHE
iU6AO1Pld1zoI9+iA3UqS/qIRTmRfwnVCMn9clhyGYY6ORcdelyF/szQJhCRAi0CmwkiDKhfAsvI
nDMTEBAgJEHkhMmD7cLiz/qN7ygwRFZ458oVspJiq9CjADWpFLJoFL0e+/8tREP1O4lrIOz9RdTH
VuQzdv2znej41HP5SJWqNNDSzBppRfJcx5AazzM7l2/ilfAZZcQXftyasvqR3ahc4CR+oFBGNJfP
+BhW2WsEFfobvYLuhOLVTMPWM5hwTtlhRQwPlYeRjuXR5TqhUSVgU8mPbxqWxG97TLddklesYy6Z
NFuFryoiM3FTkbfUkJtO2axLTylYUY1FoGbtLOKDbamlGBicX8N8gfMpNbPX99skaxLcu33jyCnb
B9XAL2E/tz4OW+E0l16HH1am+6V3w1A7MzmDQ53c7GP001G1Pp9zKqjDezz+KE3ZK7LDP91cShdO
+SBHIkCDD323y4V3jQwxZF+4a7nQ83+z0lYyHWMi98nutBMNbgcndqSeH+wHp/uJQqtULJwq7Uso
bXtfI6fZPFdC/0fSwXnPr+91T6eRKlV++XMVcHRFMS0eDBEeDWHmobj0xAUqVHRmb/2+XsC1YuCF
xwGTtPT58t5K9MFLVPO2W1CrdqroDpELpSddqtegIAKncZo082TguTyXxs0dF/G4fltwneuQjR79
g6Fktfyy1uVeqwgUze8lVM8891XV4etzzhOlaMvdTvOXkyL6ACvkC7I3BlTr0KfGNNSlcWAIkg3o
NrxxXEG2FBs8VrdM85clUEiaoKNzQ46/tfZPJF/nZnj88ERVAb9ldfYp/snY77LzQq/jtxhvgYTw
KpJqwYWx7pg1+R9HVbkSJm19kwTyjcHybHQuAESBorBAmYMa7HzJ2WHIn4KyRayVLPCpjdSYX43O
7dBf/+EbTWVLWCP2DupBTTwCTQ+NymKINUL/yVs3l2/tvZLIriFauVQ2ZutfHCVKnVhl7T5EjeIN
W7B5JeETjAHWG2pQFDEFihBUJUcKmcEvMw3kH29WZwhqxTENcsItKRYko+HlS729dE6FH7UiH0gs
WLh1eeXh+LLL42ijf8mChvvj64J0wEtfHCPiyDUANdS/N5kMf1ABD9peE5q4HddSNYNJbZeNoEZ7
01TZsXsvcneVaGYLLTmiU/o3/CBRln8lLc2XgGlzCvzrq1QO/lfJ/ENO6qrpkYbNGaoQag5pBxon
faS3t1lQv5nrP6Ihu7cKLDM/ZnMeQPiWkbWPWJ/XK3E6kCy2vVPL3tRJOoBalJ/I1zULzf9OeB4E
o8Od3QXorftm5RV45O55qDn9BjQva5pQqPdJOfbp6OgafNVsx1kY7nsmL2Mi362JzPyP+jt8ENzv
1L2nJjEsXG4jnpAgoa9tF8Hy8dhWVDC/6EfAJvY+4TNfpdj8Yk535v5Is6VLvlS/KHQalJ5WtfvW
ERd2IXYKreYcps+wb/X6EnyCXB8iChNo7hdk00BrYUe0ctdAnLwaZsMcwm1Mry9B8PtvjSx3RWnt
3KaU3TenyP7vuHzfueKyUh8ZHpKfT2wRc3CDQuMCkD+AwOx5zic5vg6UBLNialeJnSKcftuj8Lhk
/YSYdNNi8Evx3NjDMCFWRlAh3sYkA8Tv6uoiEf4MfBTxxJWhNm3Tztm42qkyMqt590Qbi1VXuKa1
oRQSoNjeGVQgp+4e/uDnrBJNWQQ9J6GC8hKc6xdjEc/RGyTa9OKoP6xb/ugM/M3tn6Nuk0drIern
u67c5wQd7Nbz75yojSepByiydRvC1GRaiCq9YOEVuxWwXU9cZGXNchXPqhgBwBEgXSRi4/Nc+03Q
HNJus++jOBFPDBMJHjlKFtkhGf4SRCjbq8O8h8Xa76MTVvIX1NjrhmN+M0WqlgsxSRH7bi6rRuju
JxS+qoBUBizZffVCpRkGgmQA674SfXdDpmlUMUgkFxjyamYecU9ZVc6IwnyZT+T0qE7LpMQVCVAT
jewMzi92Qx2xig3RC96v5BdHy6fV9QMt7svdXnxMb5pmr+EN2JXwu+Ci50dhr9+wYTH15rcy8Bjw
vWCPUgZvCPZkXNzOlAjVsLOhWIRylqUPvjpCVBWRK3mOtnGJ06Snozhop+Tu0cjAiKEbfYoHQz5q
aJ38fnFQoYSxDOY1RjIojd4lA1TYt0NFTrwVtcLy2buQp3axcfLJmU5dq8kkbv+QlnTGmicrO5Sf
oMhDVWH7Ho1/v2BqO7Gs/o1gN6dMkjUFnmkDQp5MuzEXKl3l++4VIoCgMFMs08DQes7aCmKqEmk/
VIZ3a8R2a8bxZ7AGqUFjCBaGhkVctH6Jozx7lbhpQSqHoqyRlMorU0oxQXmHCoLh6za82joKmCAv
MTYNcAxCU1VW47TGqUaIc3+ObdU8qyhKqCSlvVvPrb5OQltpmuiX3Sig83bsmltBTnkdZz9lsRA+
YrG0xw5FzMgVqwD1SWobWKt2bfubo4KzJLdeGnXyCStnL9PZA8scdQ3TRvXWX/h3Rau/+72fYhQF
/psPCdvz4tvzPU5Xlmvxk0qELxawZ8/0RoAtfcIegSThpRT5X0pESmemVKb3slJtrMgshQKbNty2
bkkc/fxCewp9+TqQJysyE5puFBEP8zM0jG8OigRnbIyEa+OwxMJPuenTIaaMxjL4kjIWEdttpcfJ
3ckD21LlDk+w/Ch26mLAJXAKHBIZG1AqLcPilRjDuoA39Q+gxCb0Mwb8nEOiokl/pZx27tTS2Im8
NuNbNQN/yY0aHz+efz/5clMwTXUZTgFn17Ia2w1nDBp17lJcdOHN7Q2tPKMEw46vGa9b/RJK3sQ9
KdevrQsxyFGdgWR2wd6Fifyz44lRyeFsrO/n04rOE0PjO2kbcQuM6UdQPPtGpVuMZvQTnV+nmOU7
f66gnpLA5R1SVH5cVWOHL5hKXLfcTpv0Qyo0OepMR6uXeFmB6uikC5PrrRXK9F4HGkxsi9Njd261
OVfAtp2UdpDUYeqbMYGEXhjtLYajE4Cf+MDv97qJlCWdgvwPwgm5psl8PXLTZ29GcxjkdM1bOSMC
Geyw4gAiqVccmW4fKLnBEUghvIGE1cHFDDaCSy0sZRIs0nk69/qXxMI6YFuwUcbmeOXYjYqw5zk3
gUcNjx2WdNWABeLJfyfe7V+xDNni9SdC32So2g9CWuaGCvawAaSaV7KBh6oNwjFFB50HYU14xklv
3wAiOts8WQMR/5bG03WwFPMEHVQYnxFGG/jkX/20oVuGgJrMYApTP+igv9wUu+9EO38knirQ1VDB
0udOwz6sdb5GTL38IFUw0Y6QKix7V3D49p9xvkWyozgRXnJeA4jVHyGw98J/UmIJGbq+FJOq7BUb
3hK1VoNK5hUCujf0p6QUubkG5HzeunwZmrKR8pHyFgO1/RdVn3GkeSP8pEHDjYAgFPzOYJtxRbZY
FjC2JeYfUc42+uSLzfJeBTCorumaQybYyMN/b46HfPwJRkSwgeTPTKlxvlkDCyE7Ld39+P6A+8BX
xwdrfgB3cIdqagY/xKaQQon5iwKMaxB9TTLdGO1Kz38sGYrl0dCJT4O2hqqMwxHJspBZAjEruc/C
ZrnE5De6cBmXgw31qfxtSpOK54/gqPC7Lkmdz7Zv9WNgSUU+5+JJ5er5xRdvsa4vYHN+CU+G8fa5
/8BBTiVCyUQm0jUm4OKTeSzTKFs1K4LoW/wLVuiDlDL3RcxjcBgYnaf/m0jCeHKPeS30PuN27fo7
osvYWl+wzRL9i83YgkraBo8ncZ/QNZ7WVTNKGqttfIh/sil259TbaBjoCHYsaKNTrZNDf03kcBr2
ni9UHEaGH3MWGt3O8WZoPeeVdOIrRfohZ8W0lGfMuATLuL+rqnZAhg9GmZZyQsNmgckL0moZxLL6
zF3VzL/ssaHf/dcNsPyBmhqOIIEbat6ICrNWABQ6TgenagubszD+n18EaT+gPAcSOAkC72Na0rux
eZ8dVFYb+ZGNHL0gew9DP5qvE+lc/1QmC96Z4riF523LrSdsagm7zXGW5sJ5cXsbuFCCuxsREY8y
rL80Wu8zURiOuNMVtFmLizB04QfD2wuO75ebQqBvhi+i4KhCAI8t9ZanrUoIQqFB1PqGzAvOv846
cFZjGiy696vve/yhoKq4qxaoTflzxm3NDji/w96MJRt86i0lXnavm4WnP5iEYYq2K7X2lUVWsCoD
szBCLBBgmQBgwC2Kmq0oSNSFAtgvhCQusndHI6LJfOAw86sh0QGGdjBkTGFoBRsAGdKeGWzHJ+vG
yK5TDwC21eKLdpdxUFllxMD5VZjJCWiVAmit0pnxHtmun5LKw/3Stui5fuVZpumq4HVyd8ydzCyS
CNJlNNMp4bon+wQ8AxFeZr41o1XwRzqnckcwm4kaYY7oUXlSim+kYpTiHQRqwz8XJfyVOc7GccaO
QNZuIoEm6p+3bHJ9Xl1BuNEDs3MCuhib/M97JEEOdII7Kc8SbpvKD2QqqHAw5cAOwGCQasFsvLab
4PYXGSmTv+PJHJO0WuRW1n5HSr8g0mzgWZfoviyz9Z/itJvzLvFwDvrGwyr6AoCRIO4KPh0Za9C9
54H0uNDawIlo/k6pFbFvAisZ5qbDj2l/wljQNMMjVqHQ0QZUVgM4WxOEcleMmfquTSodxovd4Fxa
Oc44LP+JYiH+6FtPfQWmmn8RWF1xY/DPSHUyYgl0BUALXb7WH9Xd7EwVI6tT829O+JsvcKN0zChY
ly0tC/B0F8dgGdZRc2oDHc5+VCKENHWY3UZUzRO3nUXM3mPImkH7oabn9kKnANKTAacjkH2H1D1+
Pij2fqxEO6ahfGGsIS1kvPbn62S2WrRE4kgltA34vyo1YLuBqnjjiVb2MFzeAmHF+hJNRc0agYxE
QXca8puUaFnUiIoGNue794jX+g1Zr6rKlbS0OswFcXbyMy9hQMgWtgqTClxTSscYgnIw9AoPHpcp
kOBLoWJTx2XZ3VPlj5zVpoBznScBkBbzYlUZXAwbbKNwN1BTIJwuq5NGWlKi85000jFJVCC8iwoY
BCzWEzQ4lN1WvEoG/EyFhcPOMjQO5hoal1aojMOlLou88+u6ijp0L9aKvNdp5FHNikAUz4rKNCaa
0qu4ploJkw2aQSQ4ME5l4F4hwUcF1gWDtxY0bNHxfdloSb8frr2SP/TzbGYx/xgwgn1ASXGpk5LQ
jUCUttcCr3qmNIsA4vCQLJFA0xjJHMWiKNezBuqtuE3HU0YJDnjQOt6OIXrzF89ibeuqgj5eRmct
mvvs7P/u2FI+LkYoryiPTgwfWTMJEGiBlGEcLY+9Z1L9kq4wU5E7Izo6aBS4uzt4R4m6wcRvinlP
u7yiNIHGfB2b3eLYJcWR7R0ZGDdcaYSf9iCxvVJ/b1UQe8edewVHEtwzk0xDxmxjZ9WDDdeM2Ufk
ZkdJKdYs5pJ7Krrk4+34uVQrpuud5MFWGVUZYqdxqfgQAXZaqEA3zDKkjIi6SqFpcIjqxJN1fFVY
tMwVx9JKhUNxAV+LcPrSG31SRF6vuwBH0xbdNW3mo8JGHrjBBTTb8dYdw+idbrqdyF/bdXy0JHqw
rDvu47pqfpQnYvd9G0uBqcyIGCSez2qnaVFY9217cvlQYX9WRHi+0nXGgxYDoLIXAg3A5GVAchox
4kpXfCwMrCaGVM6FlSW8JU1+ywdI/2crYJIMySlXtCoeThkFdmyOCDAAiIY65ARbZCTyaYKpUk6a
vYeJt3tmkhEvkp33KuDykDvNfAvCC4v+dEFIAL21E1lldSZeduCv9kw6EM4P5/B4uGUEywiDcRhC
eHZm1OKAq+bEbCpy+6lACBOT1aZmbS00bXpA73Pz7OyaMcYVleoChpx++RCdJf3wHupjce3p1CgB
L0+6q1N8A1koJg9MktevgWxetjYz36qd5pKsxwIW0vpzPfguLlERGQtFwbaTk833nQ7Z8Qt5Vwri
cl+kRByUSa5U1ffnPq6ZmPAwd2OBktYlN0o9Q24U5aST+pREyFpDeeZRS9QZXL+5ZTq/uh/MJCnR
QMNZUrPy+jnEcq/Ji6mBxii8I4PzWq8phPFLaDRJpZV5Fw62ao9XOi9GuQdncf3Wfb2PlLCfSGgA
/8+EQ3mcQE9lfpAgBlgVA7DLu/Ri0i1oamjkqzh/FoQmfTVygcrS1lQyif4TDREG9tRs/tFpEdBc
KSLtMlsaZlPPDtFnk4ycBvQ/Iu6+ucCxN2dSmDiifW/1hqQOcRea9NiD7QLPRwL1pdnckdxSvCat
8uCAJxVCNzU7gnG73bNRv7fSaO/MGMuwQG6pJUULRWDW+7gGNS4lVF4PT5d+sQ2y6PdE/HpO3yWg
SEhYJXsoVDmJIajD2CCYZfL9mKCvCY367YzhUAgIEYe6pXkITLsoiPloDhmxwbKP0WAuGii6NU10
WmQ9JJuT3oOiEn1OgvDsXmfvPHTbTBtUzEwCpTLLr9+rG53+LPR2L1LxmDheOKzvyccrtcx9rbOD
1Ko3WSBvbM7/K+uxk01EJ1GPu5F/EYuEUmy10e3BnGfBe5JENLQ2ej9LNBQ9bg4KGX2CNtFAeJT5
KIQNlWv2XSqLK5fOHIHN4SvCXTijHrRWvDI8eNd8rIbkrFAdecm4Hlz3LFTk6dlKExnwUV80tVWM
BCk3p3vqoMJgYnTPCa4iRK9tYICyP4NbRIgvxl4KExaUtH97svvYFeKRxccZlxpquOqx3OHyCc/6
Jv15597prO0a32+4AGqSUKQD0FlOnDCXKWjfYIwm5KbsOwmYv+pETcwjQ9fR/+gg67ee9xHW21H1
90TdF50SnHjfob7t4vTvC/LK9k/BA8RY3aoN/nAW64u37rrFY+D1OSstZV0lXj57n38YYPpYtwWD
tFOZ/bPsYbeZoXtD0xvIYfHRxoJmABGIwx0Qp44xLIeFFpxjEDNdARVGQw7+lm08aiNHj3Gm8I2N
4J+AWhmTDstg+D7I2q8jz0JWJMX4FrR9n9pal29waqYlb1cj9xKFR9KpW3btLSekvtaP+UDQrAcD
yyVt0kNfvuD3KFsQhBATg8NVYM8jFTDDbZHebMRwWv+OS5U3R0aFzapxyRaYGWdgBK8K7s2NZxo1
wAY/+KAjtNjOpDTUJQ095UcJ/25TmB6fatOAzkU+T6FZZnDezfqm5x5TG/PlFPzP9OkelU8wy1FH
gHU2u4LV/dPNixYLjpJfl/rKBW9sq+wwgUIA1265zoiARaet8tXCzNEDaL5cZKbiXUwriYMWEJo+
OsGqx/4Rmuk3BQo8dzdoWGyQWGcvLJsnf3p9ecyMtWnrfPtb4ab8ByNaVdYv8xhQp9GMr7X2mwCo
5TIphgPGNgOsS4d7JtTxRs04y328ExNq9Wtki9W8UWErXLxEieAx9jzT1aB5RwZTVtjrvoKaryxR
tmpwBpkXDNN+FFs3SfwJc/zWW9J32wKAOrf1OGzCHEgI7QHcSxw3oQ7+EkknxhdbGdgxvd+788QK
5uqt9QTck21/DaqoHehwR8TN8jz7wTWTJGyk1Fivp2iShOOa5QEbT454MxTTkCCoBW2UJHouVZIj
YhsK+TKpn4x6N6CPz6u5TbcDJZxHH8eFtt5YLgNLNv3NchIFPhtXA+sQgwlPkox60hPC9hKe88JP
NjncBVA16qpUqgLvfTc8B6/Q14a6fjlxPJ6wMc1effc4w34nC2znJnMQhmaEXRVRm12mDYttiTEj
Q6gC++Rqg5u6ihBcl/hRXxMYKyZI1IPwZmEX5KdGowaM9Oc1/1Ti3fsEEt1aogVYTAareXQCL38Y
XWOkIZz/vFiXrMoK6eXwF6mhHqWlAw7whykFAUQG6vB3z2Lfy7gxnk49/urktYk9LfhfoyP+2ELu
nuKBqWSjWjgRpfVm9w9VLaWdKjhEnGBSOQntANfkgGP0mUar4BVPMSJo71gRtNH6bfcltp74RTPp
GlUYBzUxZ6FPQ0ArPg69VIeev95zgezW/ZjlzPXnv9vCOLsT32Wx5JW/Wn2bUpYelNgyAzF1q3A3
DeNjZpkh+SZmRK2PwKz7p7x/kIQ1Fz5EDZkbgu7mUysUbozGAHYR2m1j2uzkCjkQL1KIcXZBSLoV
iCiHrmXMU806CtiTq8vysFahyosSbEI0xBscbPXHDkNH3lh/An/XxgLnu19nBwMhJSz9EQmV6vwC
grIJg0kKNt20ovYYDGTrqZZFpFfmc0p7vaf4jDCymL7tCZiVnzjC90i9x7GNDsyONNm+V0EGMhkT
p7Lb3DRPiPBanWhvAkIDByxt0aQ6bai3Aks0EfSuav9cK+3PBS/vi1LloJqQVYy4aI9lbCQSA9or
CPPQQWOymEP+o8SSVB8msPBWNiXazLCxuUl8jDi3YcDW3YpIOxPp+DsQ1F0Kemy/BBi16JuzqVg1
eEN2QJ8mW7Jtmd1DtixiugQLR2jXKBCzP+Ehi3q4QyAqVWSykFmtQS5wCPXeKunpx27+mGVQKwyD
eHg60O+ypTL0tTf2OFTa7k/zN9A/CJ02tlN/m3zlrLbjoD18D0zC01ibgYoXAWwXk7Oi8I0d1Rc/
Z+Uc3hUDEmttJc97AnfUyzCEtKqAj5JDXORA0PrukSGJLJWPzrxz5a8MPvJ0wRcgdbQvI5YxuvTE
sMJUb7oigwQrygiwVUVCJtRo4WwfEiE6SoCbuvviOhHojeNV5GFNE2jpetaMdrH0MxVucg1AdOrC
vr938uRsEVh+JIKw5/cyxG/kSxewe5+4kV1UcVp0dj7+RTOK/jSrJcJh+1yh8mrkoCL1LVGb1eDD
k2qpyJtCRkVLh9eC/WTJQcFYFc62OAHFSXm/WwaiO9eRpGDklvmaVElU22rdcvdKA7/bTrvcUFfU
XUEzGs66XkEUMZzJI80dJzP9kjwj/jSlFlUc7CpGVVGLR375tp89ud19aosZVxgjS0V/JZ2KhxpE
ar35MJEpr3XxmB5lnekiAphPVyhfcvRM1g5Cp7iEQJicjMEHyjWd06z2Jmdcs2VF5X3d3RESNEzn
Im/+O+IPtowMilyn9XrXAGz9BaCyFpKhHWvG1H8p29ke+MU+QF/KB+hPxOFZugGo2a+3U2b7xDtf
7WU/DRIqW9ihjAZ2Wp/6oteNKLIQuRVMEkZcYevHti922X3Bw26PV4EK/wCm1voey9JN5/BFQthp
dsJSkolr2Qk1PnzXut2KminR/QhIBcpsTqloGv9YsteT14/4KwJfwjfiuXUJS1mvnUbPEv8sR4iu
jYt++FcXKhm1tyrQw1KkonVTcR9GFBkBvYnRQipnOv8dP9WmDWOSk1lWy8/2QDD4LHGdWgVC4CKv
w7Ecq3Fw0gDc4/wzDFhlMDVcCbLbPMCDAFtK3AjsOMMVvvT46YoEJiUKg3ixt4KMT5ci80q5CpZB
qPXOBNm+9EZO5PdZNVyYc69ZscQkmTPMkEY7n3U99/2JL/gOZeGnFwN5dz1/uwFpchej+NDbkp2v
RKWNCW3GX9/Lstvp/rVCLOWzzah/3B5l6M/vKinKbX/J7EWEXPc6xEjt3HBwBOjkF/MZ3OfGDvvM
T2+jarw9CDvV/ekZlcNPIXCQpSzKhGM9HsBiSpAkRmkQ+EHEFUOVxowf07Pv+NEqfjGTr6rqM/g2
XW13QvpvEXi9IB85ehUfZtRqjKoV7kA6eU9UPR+nJQe3Ugm0VoI3l8V27dV6YXn6aeGGjfVbi6ap
umP8P6VA1dgbzosDSq3y9fQ4ZpwN/M3YTg7Xa25jh/wQAxmYM2aYkd+WKfVobgygTS2ROuepkrFc
LI4a16NgYXzm2/M+HYMp9c2rlDP6tPqrVKd28BozWR3ZIumzEuffLmRLnoT4T+lqRaDkZM3liecd
lHbVN5/j0MgE8pP1DcGGdPI9nLxRrD0g8tWDgm1Mbw3C30CobIyVDjwz/cTJV8auRqVfNVXjGIKr
fYNRrvrNm6K3YmtNBhXmGRQqSoi18/loVity4edlBPjbffuy2Su8GxycQy02gfn6Tz77TXBcBZps
r01QQrofMlKHtYUgpELzbgEBkwXLYzfDab1v3AudHKp1fVtqyDvcwuGc54CYJLLTMyzW/A452Vhq
jDqFhjrindbaxKFpb5RGcUpS7ib8Lb0MXAfVGOcwXm0IYLfzyqE8hEA32pbR0fIdnG6/6xYoY7GL
3U820SQVYL/71iiECNgeILAvFsOwNX0K/YsZ8N1IiH//3b5IjWVMkk7SdIZjO4WYqG144n/vK8RK
DHG+SPxwzyJuwGGDlH+Ux+67epVeCodlEOdOb1HcSOqscN/Do9jhQ7vkbv02IKol0jOByes/bcAR
3DwY/gWw/Fmi95uPM2Dfzj0MkG9vsRxiAvncZvs05/AdEMnUISb5cq5Ts3+rgETytX+xXzGwQElZ
E/MtPBUdvaHPdgGx1276E7V62FxyZ1wNw8QNbtrEAM6ngYf94aap3PJUxkjIG8RFlne8uzyP36eh
dh0G+dpYUAdNJnsXk1ASypnz+nKck8xNJqXkCA8YOjpIDnErDasZ+A/VLjVY3Hl2ZqVEOsCQJU/i
hlg2LgFuVxqtko3G0Bmqa74lkKKDMeOzWSLxMYsbnlqQs6Pfg8UqsQd1YrFlKbY+XB+b85TLZXmy
YH5/KL42TSvuzhVH61GTQqf9NLylp+j8c5Vo1/t9xQ0pG0ENCWRokUYeAk87OhULFA1XsOymv/6K
Wp78pF0Cl9IiKCAF4oDaz16sIsOg99ZoEOXQ3LA7O7HlpI4gqnHeD5St3Dl0jiNkkma4BTAHr6/i
a5F2Etv2EDv+5PMjnsVSQRst/VBmFZGlFEgm+ZcpoKUf3AAA1Teuo4zfGKVk4DH8CetQdlfF4mCd
Sq9suptasFtT8/pGEoOs33xQWNfTTh0pZdbBnfIuCw+XDKYIEyATRAxkIKJuHo9nVgXv6wO9zIvO
MqGE7niWoxkSVpByCXwlVW/Cv1gNzXqObrBGWGYbkbF7kW1Ca933sEn7judA/DuhiPB4h/81UGdD
afUlxNiXvNaFVA5ZojR33bBQHgDXVmP9ajQ/mOTsudd4USoLvN2GaVCAE+qVQubGdZzBEKvUyYpu
/X+Y8BLB7YZev0pNmXCTFvK1Vft0tVUbUq4RVLucUX83BtGmaaHck1sOYN40w/M/ldB+7eR7tji+
eUbVYLoAb9oCU2EkrbPVE8IaVp4x9cnXNqrrv4KiPv2tJychtkhuCU0yvCCbulxLjwEXGQEhEX92
s0/F+J5/qeQzz8Ixm89Q+V2QG4pKGb2l+5/HMI54Fiv3X64G7d3qyYP8RIfTC0hCTkmZcRTZbVAW
7v/soK1HhlKJjRw2F+yhN8QUPcTcZl/ZB/vUcB/2tqMsuOjziiNO3EvQA8eL2cbiYmkBvBwUglXh
fKEhf1aEBNx2th2BJcTbKk6VNJcGXFyZugHMpTXs5gc2P1XlxFVTYD6Ch7KqKy2KQzwI5TJnEr6x
Z/80JPft+MpryK/jWxV/yhue8tQDMODvOkOtS9K32G5nmSLiqnTleIj/mGsOBzukj9sgoJ7zXuYY
BB5YTjDNruZwiJvXkP5QIHbXdlOx/33v1QNRpuJZkHEbhKDpd1KTAV9i9Q1Jw3dD31QL9bjZz/hH
GnHcYgTqH1If+OjQT7AfOy1XgFecM8ayYyA5/YEH11Kg/VrCV0USNrDHLcw/oG2BCczJYOKmhNTZ
TUudQbNfUpW/CTl7LziVt9NtFAFjmDa4qlINqlWBLAstdSx7yuQaprR2fzUUKczF3Y3rhUp7b7qR
szRIlMGc+iGLSsMDGuOryQVmV5dPDFOMnyBIjkC+Y3t6VUcEfGNhR2iJH3touVKWvAfXsN+5s82B
HDhzRhEZfM6j06uEAIXy43ZxBcPxfE4AONk+20C6qGxmrGgijMVnRmPDeWkTknabbxR1nONM+XDg
LvEeEfeca8HVbKaTeTO7MKm+W1zCa1ExRYU0dSfdTMWPROgwdLhx72q3lXZQo3iDbH31UrW75DNa
/I7qbUW779dtX63ZsogRLqLsS6tZk0L8JuZKzVUD3lCOjiYnOcC/9jvYGojQ8Yvm7iNavYb7cWoa
rwB0mjTC2dLUAFNsMt4IVBahG6BUheZXDb/Sid2KXHq19Qg/qQSMrmyV15m9zMyIqjB8t0ukAnG9
X8RkYEc0jDbbd4OPhae/9Em4q2aGV3F6wW2uZcaw0QhqlgPnpMRWwxm3P4lvbol9+Ri8vO3HFT/5
eD3tYKQTW00omESyYhIQNVuPdwL3YPRFAlr/Tj1cOp6wXzAP/2ThzaFjVwEWDyGGWDLEGZMzuTU9
d1wiD9l6st18JGpZbhPd4gMxMJwFUI/r77qxAF/JqOH9/xxrt56fNHV3TcL7MCjgnoFGdyCQq9BJ
E4qnh1epebCH8jqvY88JgEIjA4fB4hp21XXEwNcpXW7agcSWLNGm5LApPS8H+CLgebEtv2U2WX6p
y1h3DQvod7OW/xJM3WDarb9N99l6fHKqJL2XJyFaN0xahaL5lht5jSMStRoNwdJZHtpZuH+dct8H
ZQs+S93a+4mqRk22cNhLfY95Sqq5VGd20poD2H+uo9x5A1oUtPlT1bDrPuff/pfrhohX0KesuJRY
JBP2eJwhEXS3egfINlhoWubNGFTxG/ZcCOFj49A4cQ0mvX0x6YdK133GNz3v69Ze5WwIZNscLgpR
eJnrIO651/1TgccSWFaYEVuiMMqmn5Vy2RlJ8al+4RwAGOQJC5Zqg4k5X1inlmpF13bASvK8mwsm
jCYDcFznNjmECs9rUlvsvVcmf38p1QYWUmYxNSurKnfDNSFhjdZ2VHsBoF9+On+gSZUL34P5FNaJ
0WTvIRecvCAu9lk6MkeUSXDbbjyqdkuv+suoclt7NIpalCziMH34n9t+aBpm+dOpxgXtq92Y4u44
I9bRPOX0U7SnqxPMRv36KPD2Ic8R0xU4hEXPh2xXt8x17SE+iGGM1vZ7XOm8NsUkWI1p9RTCT04h
HDH0JPwmMaxwaenccE/1FoKJr4AO3BwqPpq3Nv5GfnDByGponppSMoZR8He53VQBghTiWu1Q7Xtt
s+/ncGwsveorVjYLxpzPA9TIG7fv4ZBjVdkRlOriZsTGZoaXv+5RKTv1A99Wzk8/zG48GbAvsC1E
mvRiC2MVVTWpFVfRx1tvtu60uAJSkXR4OufG03pyScbyZ2EuoP3tYGAIzupRNgyZoYm2RngKpHRP
BIheO1vP+wrJIlPy3AAeovCIr17pX3KYXJgk6G9t2igd1VxITpwH3g22FSbFP0y9ezj7GHPdtnqI
8Ez4zTaUkiFEwjYPTh9nPwhVXqHkH9chXN3Zo+WJTeVjA8H+Ai26DZu0hO+Ttjf8XKHVKfB5c2UR
nz1dzG1mbzvPuLNCSRKtkm3h9iVtRD8bP22byrlpQHIQGsCi9bShcaSITcbG0XI9eypRBcaOoZZi
UIhnzOBH73jkWuPJQnXioDiTt19MLsGclZVDmY67YSQIgy7V5gU0n8vgBpg1Gn3U30c7cQs6dOOK
cmdtHXxZjN4+Q9efDMrFJi84z2GhZbVgcBmHMnw4OpD5VdFY01w26ev5KFZmopValckJN8ogJnJR
p9Bw5S/lHHsEd+YdjDJidHiV5TVmme2VBFaKfLHYGN0xhPXLZgDZnq5h70IE8A7UPLBk2qv13PXA
3t5mmN29SPYM5ipvLbk3vRjnzR58zOPVmo/ZfKlmfJKIEtmQzyqVg63YPjNngpZtnqb0xlHY2xNR
eXRvGsjIs0ctWKf9UcYs7ScwCtfzyVqE2Yx98oJLwpjigix4n5hFSz0tVapeJzCQQ15tTeK0VkZ9
r+WkhE4LJ/vJg7Qq+veEzFDp4+N9+TvJe5rErNxlnOLoNM+pjmeLM2c8P5xnbyLenU+YjcZvZgsR
JlaFEivIiwmjGjpFwRjrvGPhqfdqSbrnB0dAgbw50Wu9w03pGPC6znocSmNkFJLDzTNAK0wkFsbu
xp5jiqK6cfPZkYBIMhVYfrIkxLDS5+9IHBdVqbOfn0ThLLXFel8Am9ryUDpymb7qYsQLJhQSs/f7
7Eo+agWIY3aCYF4uduTu19IQ8+wlBR/5zKN1AywbQaGNiYeQHksWwqkQPe9hVnWVvoAv8bMiK11G
fZWPk8krCJJ1Nk40TyNc2r9IS08IHeqeLo6iV6pRtUdUsANuSBfF0wchPSZoGEK8TpPCz9hWK0Tw
9r3SRQAj8ve/EHoDdVtTdRLdSxeNWNJDJYZOXgrA2JGVQLG7dlys1topIhCVDHjsv80GAShgeqVr
q1IYt4+bKEE46e8iQwgrfldN3gOUb7PufTHGsHJJFezwIcYgVwA2/5FBVNmOOUMD8hh5FLC3HOHp
1mmxLbLjJVLEyDJrMCiaPlp4S3GNPCfNpXXAjB7bs/vaavxPcq48K33+0rNXx/o/7GOyqrxwk5Bc
STstP0sIbR/7ybHBRbwHL9brIYdK1zLeX32Brtwhn3ayNzeYdKD/gMnKe5MUUOvwRHYOVP2PNxIs
TmMTQjUAZMQs40+pn3kXOcXF7vul9DDKY8FK0jVQdFTPk7kpaqJW93sZkF0fPoDbenN9o9Binhgm
5TY1EDcm/001qpggxMfxFgbvBUP53+Qiwa5RhdSxe8Dxvx2+Bi5cDc2/nOg9Rgr93OPPi1KMzOvr
btU/rnIyRkwqvnzeqie1rUknDiXWD74c4euM8k9WkEpeGlW4Yq9kKSKs2zddWHgOJcFebwetlMYX
Df45XN16F6FWkyk2UIVUmN2faqe0nW5ENcqExNZLHrABuVeD9UWDsP1MOu6XU/YXbLleNXNEXG12
BUQnb48eG1lGKVeDEsWDu6CVJLAtorxEDo2eJIkhgKdSOLAu6q2D6pVtDrbxMw9bYo7l8XJHr/la
4ZiuCa1f0BE9jsN+eRvOqZ1z+HJGBrnPSF5NJ9jUSzyLLNjBYpYXaTQELzC9yJkhmRiH+BwZCrZG
nS1UYL6f2G5OXWR0xHFaCh6I4aaBZidfWIueEU4Yv9hZKrVEPIMZjkrdeDKF4F6JysHOf9Ol6mo9
m2ukML0SW/2gzIED+UdwPECZ4/lg8EuMzH7aQxjintIV+kI1nnUDn843cFpkcogyYocl5irZPCsW
RYxjjQCKaaBsUaOyTNXbJzWBm+9qJzeMO5AbbiqhMEumlCyo/LBvdneV/wr+oUhYsaDayqv4uAPD
dc/iHiORKocaGdGDkav0xjmoj3Z//0/QxCWQduhnjgHYKjm4RV6O5TXZgqtG19yqC4rpATRq+dhK
JOz3je01CMNQPqF7R/3ywggAOnWgDopaa1aMkh5kWzc7BnQvt3msgUQ53QRvxA/aIbeux+ItwwA+
MUXNdqe6vUIYREjBa1H1vGZNkujFxQOOl77bK1pELP3RAjS/yl3RvzYO6NxkYgt24/iboMLOHruR
qiqnPK0H+SFRqw7ZcWUpvTQAVMByHhjfLq2Rbvlsi6sJu0gwFn/IP3TpMa8b7pxd135VLuOrWHhu
ClakiwpXu/JruLHPh9PvSnr7SuU2qk79XJ5Y81b3zhjEk52zdEYJYB3lzW4DHDeuhy8jpfUfiXXj
ZqU/S9elry3OmtxWmZvgryA+YVAAS7c2l3oxbzD9AVaOnN5QClnOqkJbPnuzWEyauM8oIcqBm/1x
SRz+cNgNO2YAFsiN6BdLq+uW18xyb6FY5RTshGm41OEYWBLwoOG+rMhzaF/YUTbCHYCgYKMLD9tK
XBJLudK8PdQ3W+kfE7ZXAh/lRf9p8/bKvlRYd9BKSq0weKGoDz4uTYu7eR4vZXZ3ux4kDmVanebn
1Gz/b7vdA9wne1pvlemAsErGeVgnOoqBQBZ1QUJ89VEONIa/4Bl6NhhiHDS1krKUqQIU45HiCFvs
8p5EK8reKhACpyIs5lVKQAEMXubsTWf+28SOpu7Y9qa1HeNGjfsXF5rBRBGmpdE1ymQyLV49K1Mr
51lt9QaTsmxn1is7l71PwhAjX53ZSrVOWjKb2ZYSoWDOnpvHLjqhEzmKvnRI0j+Z1Hs4nZNUSIAy
8eMUC4ag5A9baQ2TjyhIdCDTMqSyW7dxpMwDSUW3Q7jqn4JjCXyI9oNJN+QT2kU3Qf/N8s12A1U7
5Yu3OZNX4QGute1MHdNycmgyHLO1nEfzyH5JUbMb3yxdrDd7gDY+lS1X/LH3UiZ4/BaWR/pmSN4O
R7XoAB2gjrtSwFumYMhQwffQziqTbVuFe5sctHEUF1vbAOF0TUs6TUz42KKGEZa5dRgN+Ywi09ZO
6AI9GQQVfOguMBvBJYMqi8V7cvn3P2KlXPqE2Z+JD4LHqjpg1EVspuN3TRNkiPpypSGJY9M8ERUG
DFgnGummi9QhAH64elqMsVhPoyrSe+zwYIAXwps5JM1nq/19BqCp/dvrjKmuGbg6xEAjUNZxNJM8
78Ir1ebGCdbV3qsiGCXLMWFGiMhDwIIArZ74yctEGf51lmqL5gFjsyXgrKnSw3rbRlzUcEHY6eKZ
fxyRDUPjcAlhKqhK97ZtFnLsb95NbJdO4K0PY4L7frogRqmHp9NCNrPuo9OPbpGb98Twn1JBkYgb
DudK/1pWUCsEEYrqzwKWgQskIjwjgt7QBZZKSCcWIL9tdxZrYm0JNIOta5AeqvBoY98lx8nZ7RRa
OP2VEh7UODXdnMBSCKrG+N1EpWN9ryd+RKvXTw3IJ5J1DK20GOQd+Ww4PTgdMhWRakqxtmWQmlu4
oQdyQk43g7BrYG/odcVSXLKkhHSxuLlawUQ/0QsbGguwauhIG9RknlOy/OceC4zwTdRr4mMgyKqJ
TyDKpWU2rV2rHrZT/+gfSkhWw+T1FTdOck0ZnX+VOSj9HTXFEM0TZGep0vZ2sdYwebPUjtAy2g54
Fji/zBhTJPy57ZIZo9BEHiHFRP6v1A/q5NbpJNUxyJlNhu8UI44CMm8o+SPI/u8pDGp66UrhlsM5
V7aQZ+rZDZ4zZ7H+J0SEW/TvbdPVO6Kaqi2XoAS55By9wOWzJ8EpdeA2QLd0DTWHIzbBpucJFUCN
AtSRAJRtMZi1plGge8CGEf//P41nTI11wI9Blz5rV85j0RQ0/DRohjUKuJk1hmzMrUv79gj5/5PU
zm5iX8VhJ0ujEMnnV/Zb7Puf3PP2cw2JDjI1q213VugqrN2tM5QlTHtqZZf1fRIkO1CHPRONkryx
QFCCSgvekDq3TFurClt1XCuI8D4zYu8Fyntif+fg3KQygGHCFmC+T3lhmPKfalp8mWmD7Au29sHE
5h8iySWu/0Cy19z0T3ykr7456EY+E6zXZ0Y24P6nBfPnLlGgR/OJv9qUQQ900X4qjEJHeJUiDX9U
kLmj59kwNwsM45bj/PV3dnFzzhxWBT7oglCu/7OY1FYMNpxWPGFoKeiOXI7q/IgzI8SFiXu2VKMw
beFDuGrv6eQrZgp3unK7aOa3HJ8uMNc74tjH7feZnxJOJ3clWC1WCT+OEuYZ/BUpT2AKeZ935C2f
JuyVsHU5D3Xqe/+A4UfvqCG++9ACZOsT5GLubj306HgKLw5P7V5HBKwasd6VZ3i929inTisnjD9W
OqvIRC+gWOvxERkuFjfU5wlpT0OKrI3MYFtalFrYB5XxOKjIglJka2u/vR4Slb2GBzZHQS6xw+DV
jBijXDkBTGV811J0x+9vbSCEuX7yiwtvHndnBn2VM8jGS5rGTMomHm20HLqwfwGl0IOO1rIExv04
BBNNJ/9S4KB1fVBCApUd+o6yLZ2O+iJvtni1QYKCNr4HJUiVEMnRYBwwTS7zKoamse1EnoOCTLZm
IJtaaA+5l6GmCywKPM52Pq8mdS5TpgUTHZsQ7S6fDxtyjIFKcRb6D1vOmS5PSRNrNyRVYBKn8btG
0rzRs91lgUPCTEXkqHFZpMXHPu7V/oYPDO0XWxbwhw9aRgA4Xa5qS+mQ5zxodIIijmBNnN23OfDX
VIf4qGi9YyZcTykxOL0WCoI/nrCRTs8fBfXoMj5VY93jKgVkGuDIUMlArjeu0MxWPv8k64NxsDV8
nK68YD1qnrgu7TpS5ZfDIhzfBTZygH07oF8PTjAK5LDkgPAKDCaE5zwgWLW4vF5Sbp4iZuqfHtv6
QVc2fF4LHRjAsvwkWywL2s0YgFTmW7Hr+hPP0Ut7/JD7Vh7F/D9EHzCZpXXo7qwAN4W7mjKh5jgq
A7ePHu2ybpV+t9aAT/EFEoknWrslYd1V+OpjYb9cIAgKbbNg/fHt3cGwHDX0ypKvHPm/N0Enoi+m
UQquF1s/zm75WLvecD8J2E0abR5P+/sJFujydWCQaI7IEZSjbRncZpCQL7lwDXuRbMcEcv/SZg6e
ke3lQWqbxQ9Eqlv47PAjg37gegSWbY05hSRB5uwYPf1mpT+QsvO6PiKyf/T0DAQqxPAllIuTL8YS
sP0d/42D6qR7o2ATKfzWDti/4W2I0wo8VDuu7Fu1FqU3/BfM7fEy4JYQYhGCKHYpw5VcceYsK9iU
ZqeOB1+UJ6m29CNw6ZBuHEVgMd0iHFAqmp+v7nd1aUJ6KQ8naczBJ9uAuwFTX+f3dHHRJBqMxtJq
IPIj8JeYSLSF/vrgwIgERJyttH97ePkuBBKynuy3v7QRCk/ydHHfrCexpn8G6J7n6Hg1xNN9z+09
t2lhaFIPk6cNEQ3WXg97QZWOHg/5ViufE9qpgxPzsE9yPmL8zbjrxp7Y4mjPc0GTZdeXSnG4GmOD
FMU96bfZvMm4Pdvtpgm2b+tf7Nc3GP28ovrSXaHfrAbPn5xDF8OSTRaf/4YGUb+p8NEdx1gQ07kN
0i2yP5gJl2Lyt9TrT29P2qpS+NH4dkVHbJCbFnfQhDxOUN+krl1tYgSJTmqY0xwrCT8s7HphiZHu
bIB/uMwzdx/ERraIKnK2sWzYcCCiGcBTIhUJRElb8LXzYTtPDR74k8QG9oacdzMniBtYPBz5QuNO
i0ADplw2JCYN0YEYS9wIaZUWeOm+yc9m2c2hGnSbnLGHUdcRsdU8aUb7+0zO9c0lp01xgswgF1Fk
Ol+65SewmV4Zl9gFN2aojgDCxco6NWMR2pWRUbwH8xsI0VSAa5n45NmgqQNnlbVTkPWg4qxtfuOp
TVktXVomJK5YP7zN1+azx7prP20eOLyRKOqzNAObSBFaDkKKPnu71uVze/gzOGUuTjj8S+IGna/2
sHLHxGeErh1kZXdsPrAnVsRI01fYcPdan/VSV8OWpR2N5RaPFrnA57JqB9raAMhUCuniDICJIYzU
mH1BR3/zdWEheaVVGOYyyMlnnStd2L4F+ab8Rc4Xn8KpFOUeNIAhnYjx1FfKtvBT2L/lZ8s6e1hw
a6nOHr68BRpejgJooC+jLn8Jp1qRHRxipT2an/+bsfC0G9QBb3W1mg079yiaDYYpDy8NnmX5L67A
lSjZwUhAAiG+guudRqtrTmM14EA9MzvuNLWeRZcddt+GDTPL56cWI5+x5kH7pLClO1NXr2zZONj0
80Lm7RqHVJmVtTl9T7k6FBfFm8QSzHoQz0JPARTG3h84fycu9FfHYMRhTLi93tP8KrBrgfNvINr+
P5ofZo9cDg8ot5++Ud9/Dnmz+i2AjaOMwcS8c5mGyhBYvZ73qHhzE11ZqUiU1qz6GrHn2OHY27su
a9TsHpHiSmfkwjjLySbxKM/bWJ20TGe2YM7vU62OBk7MepiEIkEZKcStjHAMQqC4C1c2dkup5Kwv
nIfC5jCiriSmVxYUyVbJzT34MXYpvXUkunYwm5k/0RbOgEbE+mogtzJhCT7cz/x9x9yAz34rVG6J
HCPZh5DKBAdi9R0e6y08tUscAPq5FqTiiLkv8Idpxbk6E+DPScGTJ0IAknHMqgh82rnO9OcJJJzx
BGCG1P5A0yTHE/ZwPsRJcsrgBK9dFwpxSB+4fP8bnhf6gEeaXRowioY5DwcXeTWkxRrG6MXbWQdt
BSVAhVPE8Mzh7VUS/E1MMsaadN+PjyKdCMycciC9cx3HxSbHYC05OZKFy2YtDZmGYnWO5dPwi940
T51k8GWndhtp7e1nxl8AIqGeg3doNyFo4rw+QXxMLDdJ4fgRXFqQ1flBxwEAJHp/R/6malMes8VR
ILwCr8mE7MkyV8yzMnuF/YhMYGiAN0DsvjVkStgHrHn4ShfNX+bOPLLwX1PPj/J404/MvT8Xm3FC
Fq4In2EptHax5zqIptYlJvJJM/AMPPqn69VS4JFjnHlkxEcflIuHBdkqgHmma/+azx1ihnsU7x2U
2Yul5mx86KIaSDWWmGvnhAgROTlyEJBoJsluaTQ2EAJ/sa8KEgvZQJz0YZFPPNHCuKuli/JLfRS6
Z0IeUie1Jlb1qk038KUAV114EXXlotQHCRN1hsEGydJ+aJRYHwmnxdV/Bi5Tz7offdhHgglim+ox
Lw2lcdBXDyT3oxt+icVcgqLd284Rob9Dh/i5DopBSk9tdWuyvgN0k6SwMRSpbwzkPryQviIhjVHB
xUmJl2EAFs0G0nKC5b7GQ/4ASpLqhaQx+SU/cFhl3rcnY/as2AsLYAJ4nqVMZeWi3a17XvpJN34o
F7hva9cZPpftPGr4V8a1vHcaebbHNu4Y/nfgChFkHoJq+90oi7C2fa4pBS+I4SGS4cFdmXpPZskr
mJoaYob56+SxK9Q2OPxf5n64o6XhBm0sDCRWWevDYTgJVenMXpFxIS0NGUP3g4BQmdJNcaspoHl2
/HHBAeO1MCdXdUoTsHVrrM1gqbNcJFBgzd6sxAj87NvR6BjBsP9KFmmyzrYjZfIfYBr+zcoGEj4c
dbvDB46S17ITt74+srICcmdFv2VZ9lA7oIFs5cuN0AEvvcBxnOjeySKEPPxtYZ9V+EXb9y+m4S3p
3FeBqCI1wTNXnSlDvr7S9krJBT9ffFNLIQedz0V+NcOAp/XiogmOKO0AhSYul1zbg0QUTfdfOp6B
SE5DrC02G9Hp+DLpdiujRqcAWefR64hnTy7J1BR69k/6VKIH0kG6C8pxy03/DPKgSGiuAH2uPbJF
ZucSrF2+pvrzDB1Q/wuMUDD3Iq2/oVZcD5HGIMjfwpP6lEko00hhmenFEgPdtXGfJiYHdwN2WbVW
BRYRPwpZSZMxB/NCWpETDzf95MUQbOhO20OmwBBZnV5qKDwUXYnTekypE2sBldz63foGH9jF4MlB
LrvPsyR+9Dmc5386YpBwG583FLU6+25OWW6bTTW/1FuuBWpPbdh4x0m2Chhs9KHm3t/nnP9DmhxF
KSh0oKbtgpbPm7NzOmszbkQTSiOKyGcpPi5+BP5uMLc1kb4fx22GIZTSd4+q7SkV6jjwryZs8hM3
NYuuXONJExReNhUuBWz8PFxXYKprWVR1nA5p+QsXRZpPzYX1O3SDFYv4R9x8BKRQWO0mneNzp4yP
mqflCpq/3CvBH/TOrrripK8fHuJMb6w9mLP/uGo3SqRgEQ/GQ98fBt2Aqc2cHRAraFmrOuCeYx/N
PL8famPR91DAUydZ7zL/A1hZ8OInQDkI8uXQMUSUBQgl0oRCZ7L14jGYCtui4FmVmNe2Boid9PPX
jM3RUUNW4xjgx6u5OP7uW11lrDCGNf/fxWchTWxdATZ502NkeP/wYatHKhh+ygs1m9ntF+VQc9pg
K65D6wKj3oRPxQ21oT6eFj5b8Zug4FcQimmq+D8ZqZxrfM+5JjOzYGtsCNwgOje1SbDoKPOBIRwH
pzBdShLbPn9JpmycXjr6KXtXw7unH9sCTvyb3ZFI2vhGxr6Z/gA2z0ZFuC+gl7dOYVvf93HPJH3s
MrmfanNPRh3F8bF8r8j311Fhyn8WVfuEHwSjJl0S1fdknRwmXyQGOvWsZockg68CTR4wZEKuGzly
UWpYmz03N0xvkiTC+BgtbHvBv4+d54Limxr0NUIiXPIgL7MKXB2yNx9r4RBt+jeEYqh4Bl10yXk6
Mtt86RLsoJ0sSgDt1hTYPylhDdiZvaBjQwUgki90IO6CP8MRUeq6G9bIoLF9Lat7brcF/7ahrgai
rqPD4Dk2bqsJsylCSiMaYEARPdWmCdYLtg3kyFeX3ejIr1uiwirx5yS5zboVyLMnWmZjwD2nsfju
2fbD4pGFalP2AErPqjGYvuY7aTHaiYI09MSXYvQmW6vjGB9vF38IrEKTUgE5rOrUOZmfW1T4JUrO
9Ax9d/Pr3HtcABlZOr02nseqorm6s8h4axhVIVpS4koKB36cEI2f7KtI1zHQUphzXFQ5N0CEq2Xa
QJi7fEbVcYRVbtGNsqYppk3eGWwKCrVggjvx7/Zmfnanu5HDKg3xAlFake4O/JBNzKaM/feQpRRz
7ZLerXA+rDqCThmXosaCimw9BJ51WP13lfif15wul6V/QyyccWfA6Uw4rhfHvQhzuE7w+J6yFUL8
8W5SVy+8xmAHsrkw0bPJO9X7STcS/cHBdvXllzIH2gQnqXc1qHxbbDmSACrA0S7dMxsaIhVKaS1V
M/jrvSgCDRtMzSEFC3uQCxBlon3QYlN7mftbR0+wqLGgbC9hTu6Ld6WbPyruzlzqeFWIyuA9Y2px
j+9G9QYa0MUm0Ld9hSwEoyFzHXRKaJ/f+lbqO/kN/9CMrHGeKPR1EytWthMZXTh63DA0jeIlP5ri
HGiz4TK2LuBkIqtNtFLgWHNFD1icPtPqc1y3VZLoDnm5VT6R/EuQTH+F6w64owcH+s6KfKtCf/1W
VCIVnwFLt2sr2+sVjHUCOG8DeDYkn1kkcChWXP48tFZtRIIREP5v58dQAYUXD4AHll/BEq2gaZU5
n2g+LjrqzgVY/qQA6tx8jiaDe4gMJIAvk0dhZMlE7u80kF/Q1zAyD0wLu2e3nXnTkSTZUb1IWs/0
XAzzhgXuWxJ0RXET9vZ6F+a3df3WC5Wgf3hKhIsIHHBr9Clq5caDx22iw6Pl/+l+tp7npX2azSx6
EIQKSoi9PYQDcPT8qK2krv7bmAG9MENMV1rNNYDAn0LED/31NQLTHbRuA4OWVwqrFhB38X6/v9dz
ekLlbcbisBr6olwckp27MU9LV/8ig0pvo5lGiuQMcvoAoEZ+FI9lModYude+UgeFiNKusCARp0xh
CmSbFshMHcSELRRHErnxOqTafM3CcbWUjxgSPwT9ZIqLdmkmbE5eahHwKwzEE7Uf1PoK7GYkZrsX
SVqPojYAoQKjcok+Lw5S5hy2slq3YK4iFTxzxZlqZACjCzDcbM97sn+2GdjFbkKpF5wbpLYYhT8E
5+FvXpgLyim4Ko+jtaI2bsimLKDwq8Pm1e0CTFP6828bRasnVSbsf6qySKmNkqN97fChPuuExFGw
la99zhthVwQH8oAZvkvMXz9j+2V0va3rslqhj35HnnN3xNPhBLWRRsE4vfMTCctP4NnWhonwDXAW
dMeyWtrQ7QK2fb7VYDdXlCL65FjGZtJ60qeD57/cB9D95IOZYhfwauLyPoA6seZXMio55lTP5CFK
h8FV+w3DQEE2ekX27rbpxeXye41duAfgdncfTgXIp0iQeOqxALuFNpGxfOj7ssSsuUVIlS9sK1ga
wBpaqiqmoFwc1cgIPFKi5dxvce92xKeiFEVp89L6Q7upqiPMr9FOzLzQpcXoSq/GDYI8IaWexNtd
YKV/CiZ76NwRDlG6kqF7EDoFpslxaZWtHYwpycmf4FWGDseBSB7S66wOg7jhe3p4VOt0LMD9yOMY
rK8Kcsb3T7QhSZMf31w9g5oRZGb5ufR6GUII0Ocg0W1r9R8OwmIrbITkYVsdZfZNEqbxCWFGqTVX
0gEXjnllghC6uuYDAmeNOum1d9qe6fk7ysAiCOOyxytu7GW1PPmDdgow8z34jlJDn8IiNx2buQWd
23qTNR1GtGH3hW1CQP1Gh/rAZm7M1q0jnGYufO6e2NlfPPtxBalyaue7KjmPp3JzzV5bEDKC5iSp
Sy1L9TyVNIyjqIHkerkeqZyDiKFeLETMmsxs+v+g3IhVAhtGDsKS1ZGAA7sOocMjDo3w7b1QKJfl
tPUqjuhBbOD1mdFPVuVAQC376NcG3/W46w5m6yzxZfAX5oPea4RP89zKQAVD+qCWuhSxRrBXFGaJ
h7iAEO35ZEmGIuIm/KyCmyWyAM+A+1ETMT0u37S40ymlDgu9HGvmbaRZRNzPGNBgVMID/L8hREzo
qLY4eZ+1r4lFtn8+q2IWK5iMQw0nIkcw6bCJ1+Phbi973OoFvd8GlY3qzrkAvz5m0BESJT+9rYUB
nz6JpWG8rlNwu/LGD5nx7omYXjzCZbQQ7z5acoKymVipEDNiSZ1sFkuY/kdgc3QRHI9c5Qcm3ZSU
4YBe6oofd+XDYMQy0k8V8sMQP61xReArcO41P0c+isy+xNbWW+pNca1BiS/KEHo68HLa1zYsrMn+
jE0ygfBOwSIhWIG9LBZPwG8HlCWNRms2H8deko/83A+cIAnrfKIKu5RIlzzyl2zoyBIfwT2k5uFo
Ek6lwMGnqrpHm1v+zHKM593Vg0GGYcmqKpbu9ugtN+dOEms+CJwm8dwnteHJvZzsJwPp6SiBF4CH
plQH0+6HvhCU12A9tgF0mN9qE9gVVgaW37iqjScPISmGyyBkAz2D8gONEGS+SdSK+vzTR5t9Vfd7
GJme67F3Xee8PPXm1P9mac3vCLf8FWhcwc2RGcvhzzlWyX/EfOs6+IxvxYPb36CTzXn1oSztRZ1E
g570RIi79X4TMyfRoxsrdz1bA4PG8aU4loEUWM/KBIvc6gFujansJOtoQDg3TL8iYNhFu1kvO1FE
RNR3L7e2DCszuLVyNQrpIcVYHze4H1c3M0D2LbKHYzrd77y6gr95IQxx26JJg5JqXWGYYFTjIMKu
6Qbvn3v6DsDXJSlMka2w+aaIiEMLvxQTnB9PSki6Cw6r/pnwfQqK37+oAZy0uDtKc97Jt6Azy3nL
WCFVOt7gJgVr6vwWfIwCPAuhoMxaUgOwN+euE8kt65aZDcUtgi1W/a2GP5cQr0TLwYGsoDfp43eL
1FPJU7fbes7vODI33iJoi2ZlUM9sXA+SZuLt7nWAL+4fjiGkmItdUkNF+/na22KuMrzVOLGC20bN
RTArabroBgdyKI4uZmIcVt88NR7Efiq4VTpILc0Zm3aOdWLHlyifA43IDrNOGj0u2zK/Mx+0U9Ka
zBe0Yrj0tWI9xAUsByq2hysu297hFm7jusAFeVgbCsGcHgXQ7hb9m/C2c1JJ93g8aveQvZsm9Mzw
xg2B8NmInFQVrrJNAUd28bgXad53HOGgfxc00792g4jKBAmivb/HK/71i+r1pYzV25cIr4ynZwO6
5QvP/Wpp4eWoL527RHjNxg0EtlbBtXttAGM0ceE127kVpfrLzyjFd6IVSNsIL6u7KKB8p4j389lS
Sus9mM3xPo4NcqKnvCHTglw7TT3fdOrD9cixcIvv/VDVLTPCLbYuDqtLOCSE7+4rqavi/kWAoyiU
Lnj+/EqyZQOY64LoVYqc13B9uEXQ5JdiheBDi/TyMUmpDrbBBwBE916oobhF1eAiFBm+RqNs+11n
Roxu9G52t6rQU6qXJ47XTpRJ4t4Z+s1NB+2HEiD5ebfZ5/bOlSF5CD1PRsBL7hTMRHKK3VzAZeOI
OTHAPmh11enFMufLJHsniw0J0nmoJ0HfZFlHOUKl4rfYPWycfssqVvYf8hZrty+73Cbk0YkEknAH
PsYXG++fzJRRSr6lb+zyvpomghp8f12lMwVEcDBBU5JgoEC04GhWDq5+L+ykgTyGk/M0wZX3KeOE
nfwYKgPcHMUxwB1Olz44VV02P3TV3oxrQPl7gwnCtZwpZhoQz1uD09hVsxslvlcyhytkRQXCEGVB
BGCzY7Pj9TZDKZv6LwODMAuMFvnVMlXcrd1Y1D3GeRDStqIiWlgJ7svQNukcFfg40V9xekdX04o3
pkmm3fPQsPwO/0zVZRmznsea/fZPUBM8FAZOP+X147CfiKPc7xqurew5II9E1cxk3NpdfP8I74hT
M14NGJr51rmQfa7tUipvlMFm9gxhX7tSQSMWPWLRxKzFTSN28hwQoYfa2rdVo32jo9HXJtAIUA83
YMVmR6bzx/Ya+mzaFwASKhMiR6Qap50QBl5726MXZj3YNYCaXNa3N0rrlpHweNz+hwP0ge1rQe3e
M/zRzgDW4x3JDDJHVEFDnP5niZMWk4SLuXOqOMChW5CKQWlK21XUGwkGE9MPx99jB+MCLBfvYckW
+ir0G27I+yBlj7DSki47vfaHL/CMFEvgPTJHxmuVYo1ANa/HzaT3k7wfLqfWRKVfvegxMLQTPmsv
90Rkx3eAi+y7NxYSYqtgFetTl5bbpU1W/EoSBbfHv0AGrewWta7xEkFP+9QiZ1xw2v0weNcZlNWJ
srScZOcvWiaNYL4I62KBD84FlToUpPdAWkw9aViiL81Tk2UUHV11c37dxrvHvor/JvLEm17wthlH
UhJ6tlB38FAdH/MPCZJL0W6NHl7ipCZSszsr1ynSnFP02pIacfr2lvyu7lASIYG332y0jGfx1KgQ
q8Vz13538GgXh3w5Bdvaft5r+b0fQk+7aRudKE88IdqoeZCFQG4mWMoCT3SsCku1VEznbWr9OekL
6BRm+uyfDhDnr+QZTiAoxj+0Bpey/cEAmZf+saTEP6nc+fOBiKkjJyOncgabBEloYYnJEFLOokBM
FHmtuI0jQVhEwCeh8nSU3ZpqT65zYbORmhAYLZQguyzNIxqvVhyrGwx4Nvp6xRUpBeewQTbDGi7Y
48dSdmaipJtm4TCBMnmRSnbq+Vh+tHOcH5mxQZ1uu5Sk2r5+uJNaKRIF1yhNw5u59xfbiRzuiTAi
FpRTemDawG/b+32GcU4ghJdduL4EV6Ldai+rHB16ueiXmiwyZOtUguOV1623h7mEbz1LDsOwYElb
5uLJjeQLOXTLc3DzKSm10euHuvpulNSqoQNYbOVMQBAuib8oINk3Ff56QV6lTluDTsG3Cuni8e9d
4XFeScixTvK+iTSu8n5l/1CGkArWvvVPNwkfET56+Wku4eA439Dlc7XTNMP33fdADk+NpMdm7Egp
BsYpVvTN9cC/OxXrbExYRogBPWEqryQMwxlQkuikFhPz5ijprPuUz1CRDbdxXcDkfT2d6sPgsvId
0fwoMclZsJtmyaYOnMoR3PVO4NfFNPxoCrM0P9S/CUMNHIuSmzEFlZiBmnSf8tRYlfJIhVEn9t1/
7cikCUJXnesr7JJTp1jfxzYTI3z65cqfmbpk1M3TopCfJV/cAz/+BE/o7+hJsZkoqkPYZvYj0K0C
g5hORGNBPdR6Jizq3vy918+tUzhGR3JDKuDYNQobyhxrDEHnYbqksZIXqJlcAWKnxoYW+fasVG+/
76CUDnlsxIPW1Qbm32YvKbr/W4BwF8htEvabJ0xgp5N7R7mwDfOeXPJtNSgt8d/M/sNo24sXiGfo
Btg24Hnb3z3zDzpNTgynjE6wdkhqFnWskE/RYUtlGd/p6L3T3eIiQprmruLKz1+8nTv5vXxjJa7t
GsJyL3ZS5+FFwwKR8d1egGVCa4FDmWa1tTCPR0i65+yKxu0fuRjQZe7VpqnVu9iEk2Cnowwu0Fg3
641DV4mMUqhQXtg3ZzBJwNaNrNqGH1XfKU0peI3PEa5QB/M/mYVu/ZAdazOb8uNDqxncBmqkJnDp
TFNR1eiDZh0idpCh0i25skxgnyepW49LoVAQZIm4jGG7lQHBcbyXf8VBVFt5STeRi5WZyKOhUccG
ATfdsTwwdXvVKEmYmikkXLhkEke7JafGzW/2CcVRsfZ5WhqzK4TYqJy8iqalbBvEfqaC3T9Kr9PY
VGTbsbs2GT1Sa9RE3BsNS8c4C4AXM+seXMkfTePU4WZOj94m2fln/lSh03/sEK2OgFK+MM2qGkkU
mipSjrNCtbXtlYGOsYizftdJSipgKoY3bhk4N+x7UV3cAujDh4EcWm+Kyy4R9Dyc+sh8/S1aFHKG
CFgJM7FV96GvDFUWdhW6B7dWDGR0XKtersKF5CbzkgEEsSLAp6DaUgHrObEzNKr4cJfXrGKuDpD7
JcJJP+oqH+kn2XyCYe7IXVxhfcBZawbISojBqXoopAtiTn9JVRNPW9SO6RQDgGqg4woVYR/efW+W
tBMqFcI3K/vlaveZgsrOVnL+pRgyZAKwBZbD1cpLa/zdnEHetOM38c3KVio7d0rz7WDyEaO0iboq
kmEuUp8OUnG5U9FdP+ZoBnfrTIAlZcnFpDtPl/PKH9Ex6wZ99TDI+7wvmgUgw0OYpQGS0TJFuH2V
rM1SvyoLkNen6s5ppRg2HW5Pou8AwCDSQmDiRLQApFBDLY9s8zzIBUIG3P81gd4qUahnol/fkr5Q
+CHVProItyKzOZryFK2//n8YZnbb7ztkyUfLPEXBsz+gw++lLzfIVzh6IhWoNpjD+n2VsG4ZhlVI
/lMDXtdMBW7eA/tlQiGVhHTB/fV/CVIxgx5k9XWT65ZvqzIEhEzfsDjiD5B9tBfP68CBkbGP9CuW
QEEeBc09tBSVHTXJYEO9Av6eeH3puWLkGlSF1MaJ9ZhY0UQY7PdC1Opf08qV3QHMmVpqFFnnUmXA
ec4qylSmYDhzNswfh6ly1nYuxTUoflr/t6JmRQLwTeY2wfYuFp4jM0uxyAeHp2i3CzY4daLMc3Fv
JrJrszDpCdey1U8je7pJjCB3cE+ZBMJgt76Mv37vbpc/grRWGVMzD5hytn143ZiABZEy2IuIk1Bm
nPxA3qWEi5INHC3Qx5er5+Ey4kp0Y2ayZc1b3vu6u4wPJTuzMcOJSoRBCXRlF1wu5a6Vy1hxTfQl
SfVSo+QYf3mhiUsb98jYZSKbJFowW6d/wrtjHw3bca+WKMKkpdKvVryMKvZMzNN0ol8bOJAw2qes
cD+F0X4IV24GVREk1NIl93tYddYE7U4rRodWxQHsOYVb1eVTdQtr0r/mit58OnD+hGt1PKvY7dLi
Zd9cIN93w/v19MGitnp93TU+eUuO65W0vXN6FRz+hWyyZvR8qvIE7aQ0CFI7G2hAAU9FJ4X9ui5f
k28Fkpp2PBuHg5c+aRrwchm4puRdn2dfLedMo0zEBwfGC2VRv+iJC5KqD0a6WKQID7iaxSCHDz/W
LK1iZpAzo2LaqbcZ/3QXiMGYTaA1BcLzAvTF6HkMh8iH0isgzHKX+XAaN0uxi4OrptFCCwdPGu0y
yZ63Q5IUz44LzN/r0FJLHhtDMSZHrD4c788qTcDBIM/8e7XpaZ0iAmx6/O++G2kjKYOOElCEcnnX
zD9/aN17mYZlAvCWcFgdF80ccK6te5DumBJ4Bg5oOcI6tD9RDSmRXgue6b6ZClwsqzTD/5UIX29c
blHlSRpl1cegxnEREjlG49sc8bAawutIkuPqgpD5hCFZBLCJHQlCZ8+LFCQuUGBWxc/RUy3Pm09W
714tfEloW2N6ceodsUIioUMO7GyYn7m+6BeLRjqynj29O27qfQk9nqFSGsYB+2jZYB3HXiEJRIwR
NHkQ/M1CF7bQ9cX5W4KzLaHSxmy1yTEIqxh+mOf+sjFiriYvtKr8dul3k89zMjnd1cU1qC7psoKv
mf1mmQCXDjMuVn7zf9QRXOHETiiu/2aRgUyEKwrFXsQuRejDzxaykjo18UgKd8/kiHErFIowJTsM
oQD542EZiXoD4X48Qv1zK+36rRLNWkUkSsfGxyodoVMt4L3XMLLDW2PRF4tG2euggcJl83NUmDWs
UOa4arFhNT+sOSX4qnqIixkVg4UWNnmVzuZYC9nXiGITC4AcJSVKh5HfGWqRoTe+IzFTjaCKSY37
5MGVgRDxuc7fKI9aYFbUS3Dv0p6L8zsTt3HF2JGnK/jHyH7LDS/Uip3vxw5WJPAAZxbtQ6klNCZM
+1p/eJ8kzPkuH/2G1mjBCjKCe01GxUTojyY1OuAPJcjTm33kjv/pHWgIkSthbDU6PSjNzeVRKDmG
NSs+4ny/lm7XJ+d/RvUBzFu514pvY4pk8TQ3ykW6eOZ9NOOpa1qab2MH1FImaHGaiBtaXNycUzuz
THViJ6Aj9ifeZt0HpLYzWKctYw2CKkvfXSFbil5cJMILeghWlaohSvmFg7UWK3WDxW/C39+hjqGW
FUM6cP3oyC1Mx14C10L1cPDpwMw+3Z+X+3cUx8xc/1TphDQItU2xs3ivcvB+FjFbVkaSRQKk7NW1
N8yeLBmTQplyd9oYv4SEwUXs5MQrw5IacUVert9j9h1sggjm6Lq4Rm01qivTvw/x4oNPUMRT2FLA
yzAK8yzvxST6mnfLcNcvd8XC9nBIKvbzqJ+KPTIi/NfsIR4Lhyd2eBYUIh6Zqi5BTT5IpyXokMND
0j50VNckcVSGQ/BRty80KVkx7XebI/kHPc0O2S29nkl7hiqNdGtpPXlSXlfVmPvp/q7/Tn3AWBuE
T1NhsQ//xbfLnyWPMgL5wYC9+UsgCtbltUyo5YH2A9UnAZ4k0NPTfiEmvc+69VqJ6Qc/IBX9159k
G54aQWLwgZmFh5PZdvqiSrtq1fc1ifB68oIpp43cfylPQjSsPK0a/L1UpISLEoq0APwpTYubXnmq
1B8VDelRX8R51M9o3l2Tuz4Zb6ZOcuRHMWrFA2kKwyKASzAS6L3GoUEO4Ep9qemNQJtaEiVEMkvT
dkvMDSKXo94rJuNGhiyo7QNFsAvGe7A6PNuDyftGSSAzxUy4JYe6BNu/cvkikCWdEQJwDYmw38tY
ubJdNT8pkqrtmDn1Ade5nO7fBXGNwcaNzWzaYAeLRIFxgsmIqqIkVkdhZNb9B0ZYbOXY4cUjH80V
lc0+W2tGHhKpQrBLbPPV6Qs9zrg5bdm0kCSwju/9i1glPSD9DzfGiNUBYwzsb/e8v4z6iy7LZN/0
akQ67jcwzQUHY19r9UtFeMxoBVmJAhnJDHitYUSmS4+6ouJHZ0KtfbsqV8VqfwMdS9vi6GJef+fo
a4pYhQoosbHXc55lvjErPy3ahhsuDx9vF/emTs85wvJM3FGIdE/HCPd96L0klxXGd/YpyOW1e9Fv
ZPqmnUZwBj8BnytuDHGdzeDVa6edeHHXa43n1QlRzCq/d9xAsAOoGFRv5ZUuJdwCZlZbGsELf67V
Zl4fyjt2VNiHBVOCHX5gYYGN7io4SoG1+1BQNxzSlhFGqif4Xc0l7EQJyea7GK5/iTUqTlM8bKn8
O/0MzTDKmBq8cwm94NU6Xnpk9fZQrF4O8VPwDAfiopa4P8oYs7gdlzZXIa/ix+MLaO53SS0NRBtI
jP9wXM6dWLqa28DonNHLMw9hvNm2ysA/SI3EN2XtRri631YXC8e7QTJw4fsAy0vF7e+mA137RxH5
i0qAXdMuDftqnW+lZ01Ls2uor+aTJUNBv407KyN4Jym/zZwMk1LSMQTGa63GcYAIiOOcGbSj/u1/
Y6JOhZPs8d24HSnGFK09gNwQig3wbvAliqrcG3aw6MHO5tF3jkw8nO5/v9vimbav8twhpPlLrZop
H/yzKaiWvJtqROAuBpKJCte5jUXWUwtID6x2jZ8fUyi5/v+aM2q/bbgW8CWkI4HU72BA7eRdRSgs
sKZlvlnasC1MHWYeoQXrFd2f7sVmclQ2TrAkOnpW2GxSC9NSQMl+RFAFvVZU4g45vl4rlDaorhMt
4+68z8b6Uh3kskmVtzRvk5lpbI05qVSxPuUOiUISwvNzblvPx4AUCAyKFe1umC/YpvRTdZ7ajPdA
Fnf0Jz+rEWKOSZCB+vWWIExxw3+zdo/VtGFzK8O2dDM6spEia4IqQgmXmj1WQAg6QC7/SwKR7MWT
ZBNDVEHU7qFTzzTQNj3+OlGKKUgIcRN1T4ukHwLDDT996hD6YhAqImuoZ4vFLpjMa1JNnCaCx6nJ
UShYWXvxo/b/MsojBK90583ftDLbb89UGTMfI8yhk4DMBAJU0+FvzkTHbPr8SXYpqARji306igtL
Rq3/TvfR0XP9lQ+8nqftfKp+jNoqdQPBVAtnsM1ewhf/LT24yRscW47yb06IAoyO2JPUlSoSjfxC
MuFQDEP0px7lJe16DhUk/PtK/3LizXKc49u6kObsRQysWwXUhuJI+S7imrrZtM7muC3TBjCmYm3M
/SbauKiWfIqblybDzJzeeNTEXJZG4Aqu6fN/1oecIcAychJINjv6fu93YEZujJUZgtoe6HFKlGqB
l1NlewE/56/sdTK2atAlZYhZIwWKuF1nDy71Db8jbkd5tRkCLY80XVbhWQq3seee9gBnuLVb1Z+Z
B88EW5WF1vtjyn/lmFgIwbWZwAB5I8z4lczQPykKaNCri/orclXAe6ZEAIY9ew9nd6XfTystz38b
C6IH+WwrMZwYRgPNVR4bv9xyx/BP6vXNhz/cdI8ND0wctRMaCt3jPjvR0A3iXqqFfhJ3EHeOXIam
uWhAyRO8GRSo9UMiHbkkIv+lWFC5dQdv9DU33szN/l2bW4QWpNKgjDiJWpVo759rKfnsGq7bd6HO
VFgYlpW22OwyqKeCQAgDGK1Bh5T/MD/cSsIXkfFfkX5hD8JAr+qVTa031GRUGTWiF9GVuHWSVb2l
7ekEZ0CB77HEPbMAb5AxeprcIISAA81rDZ0TfZQzj7PKxY42RHqq0C4BBeyGzCe5BxAGEM8y17ac
no6PZNWsE+MILgvQmxsUDNzBHjLJw/lzV/A2Mvi6EaVss+CIA+tMdZUINwVZ6AKv+6HTeeXGjY11
Ho2ohN22GJhdkp2BVoAn9qDVfFXle2Kl+oghdcFHHSJb1SPY6uXVwrT4eWTyrYIbGJI1NdzE+op8
5MS1/1MJwUYJtGxUG3EbX3hSI9eXsxe/t3+6GOcu+mv9vatYbQAd9RxdEeQugUJbUMET8pn2l4jd
/ljOkh6z16Mv/Vrsu1SNUmkXafKZHMGxA1+QWSg15TcsXwyrIRA2NKAEjYqOYp0sE0c5KmkRCwz8
yP7fpoUg9oWkvcn8T37Yd3cYNRmRMgRc9fXlJha2NwpWWMyOpAGKZjHrdzMqLBY/z9RD2lKeCTPL
08wrD68bQ9hbXOAD4VY+JRejDFQQrTRqQoV2E86a8jDvdCijWXGyyKTo2gFGnAAZZrjVgUBBRLXx
aNZCjWVH9rvp3v1/QfhxOG5kPup5xgJFPWcQZ6P19+irIdb9IDm9xNM/P1gaTwoEo8GiAn+LGhGn
xVgb/GZy3oEo1cObX2xNzuboTpct4WSSMUYNxiDJK41r/Ed8OTx3+8T4j9HKH56dEX/dSVYagJBw
uxq7qDaQbrzrti0fFY2nzDNXtz0E+LYUmr5GQmk5qT4rR0yZsTCy0pTYeurg7oVYwH6vlYmLDs7K
eih+I9XWEEsnKGgrHMSfWGqEzj1GRyMh3bfRBKbcEMJRoM2zqfngIKJ6cNUfnJJI3kwpXW3jbVvC
a5bjbyjFmT9elfHftG+iJvSRlnxZQk10M54C2wya0ROPhcHbhDswB9jwthFfeU0xCJqnWGJM+GqI
FrZQiV5B0u9lt7AFueS3Wmyt+xrOMiK3TfKqJ/6Rh/xZcgqbfDmh13id5Cbd0h2ruZ8UNRnGNXJu
pxNtqQMVOb8R7RUkIXh/7FV7QKDQlHsa021JLh9GjIOrDh1xW03WPlc3Fz5aB9MdUuJT8p3rQgPa
sGQuq2dK7asQUYOL2bzL1IiJTtXWitIDRzb6AXM7X8ZxnHllD+hpBE9+sFDwIdLutqD2N07FxygL
uF20+ALetx6kPk96fo8QHj+MpFmT8CME2xfKEzbtkG2mYnL1pXsWJoj9S1pTi9/SR69kj9tGO1lS
sYpSwok1EiaBj0foBa0ddhQQ9qVSEHVZg9WAvfgElSDxdN1T0ytNnV2LK+NWCWbfZo1PtADiBcmT
eT6hVDD0WMTt++p+ai2i1pHRANfsDjpeAKf+xYsAHOK1KixuFpES00Yv0JJkSf9CPSQqRJPPBb9F
tJW2KIBAVjsyBvTLkDrBgMQmgDJSdxsjkwt2VPgDaU4xys7HDDDFxdxzpv8hhxccumUOp4hAcpAp
PmeQcpbSklec0fLyNNvL5lWtDVHblIyOom/7saese14O6oklONhsX7YFb2oIeEApsAmxhzfNulI8
CYOLr1ylbZlXYqdMOmtv75u+lb8Y6pvsRWC8OrTVeKUZhKOxmZSGVwPA0dsX9TwMz1zVV+GpRb2n
WsoZ/eCO54LjmfKwCzpZTn4mQbyRX0wiMRFr6A2RTxNq1m0Hur8wc/Xkqubit2RK9MMSxbjI+/Jk
yoo+XW8K4Aac3+HreLAn2NTA1YhkAz3yiBwg0SURL2W4Eax3hskoEL3jDZDFqrxbrW4kQFdvYKBZ
HqRaAUg9YDOiuGjwAk/4l89N5Fwlg3LgZxS5zIlEMKmv/LUPj08acUMBTBjaQs0GPM5hg2hOCQMQ
BJYip7ELOz6yhTkjcWGAT80RzlrX2AK6xFOm4iFKSyQ1NuCcMVUD646Xc5bvrDgUnMmldkuhtWcX
usoiZDOnB224hk1Is2mK/CQQrSLXd9wyYaqD5qRget7f5usuKJF51CEYTOsIJxnyZLXqWOcHq1+T
4xZjGelkQojSD1UWpXTqZtQVrqgeSI4m/dQzzyrvGWatwWV9thk1p5OaGDlxdkzq11oj75ePDgzS
AqF2onJQCLvuAN5OARBkb9zadY9U5vpPI9r84RQ88pEY5nF1g504Oyz0p6BdaZPYnzAZmz0cLrjy
ZpArsmWKSGazsT8aH7zXf4kbBemtLt6uZz0FlS1gd2rr4tDZJVmLNmB36KZNS60tQnkxJIssgknH
FXgqDszAnhnUVVoe1U4YgRIwX6yo8L4T1yq8Yv8WvzQKeRF6USnrwuzmru01FJC4MSUwuPdSZye8
vgIx0fbGcWwMO311Za+O0xmkpIZ1lDWbU+AuMo88nG2pLKkRiYUz3CJ7x+/47q2P/VPmomLEOvd4
RHq4POLOhTGlraTdYU6wrgPZhYVHxj7TPqot/RpUCz6B5v2DbxDdcCB3axtwZXIxhVydHO6FnjpT
x39fPUCVLsCuaX9iiWvLagTfHivd+02lUou4oDcoVLJKwXZBVjx67K/F+VwXpe8IxL0wO08TeAJO
x9D3KHeY06yE0UvV7t/8r14Q90MEY6DuK8rREuNmR7pefuccPX6sg3ud9GR3mz+rDUEH2OrwGKSW
zaP9Csc2tr4VlWD02EgcFCNKNog+KqjpfJ5P2TAYyGC/FwukS2gTGwRug/ASNc5aZ4yIL+BpmDRH
eS7TmmLpBwNTn3PBV/ulEs8Djyb/1GDBeEVyNsnR+Dz7H0bBjslgAz8vvlhgNy/wlSiICqnGPzQ5
XDUzScYKqfjN88LdifDG5fLtbuXzViz92UZK4UJjCJqEHauobWa30voWLpagTJyIIcgjcT4mOA/u
hd7dhUmXF1w+agNZKjjAuF6lRJG9G5pIQHASM0BgIDQip3DDI843qCy0dzIH0kbBPitg1H9/jA2d
bnYPriQWrHQRFLr82CG98P+jCqWn/41eVozN5EC72147fpQ30jkL4OT87lBCKOKgbXEBT6QEZj6A
Ig2HHLgFf35HWe4FdYYCIYBTIBYbW9dPBfr0wqkERnq1rQDWv618L3P3L9c8nHTjKc7sobNY+Wk1
HqeJE9/2hpjv1NQ2j0RJP1slvHndo3uTUgJAyJyQ4zBAnrOygtu2uO834nSGHFmrLFqNKuy/PHq3
9+t66uDCXKXUpW6XfVRI2qd0ivjnYzaqDW2wt7MzT6J6V9EE/Gm8qCccZWX4G/SFrO8QX7tvN8lh
IxDMd8tpyq2m3LnGev8UlNaL84+LgxBf3bLQ4RqVH8Ggm9YRx9MtA/m49x1mIQ9JoJtOG+fJ2QqH
aXy2D1IYLDYFTZ/M6ftNgBfjd1sLnre4WQsbUgXokzRf0CX9hVdu7/SghhhxwFIWtfYvuK24876M
y6BV0ZK9KZiw2qVeQtBBuelDJDdiXuKpQQ1RwdrQKS9gAcJNQXKMtVO5fuRJk74vazCaxYZIIfmT
Z21i2ASUaHs9dcwq/ONNMlsvAFSMrhBd6ENPhNwmP++02c78TriaFd4dKW6xzwX3g/MgoIrfPAbo
+0hjLiDwEbY158vqM4R06Zv8Selw8Nqnw24Nx10SC6sBjTAnW8LxIvcZ2qzIlWy4LfmhFJyRp+0d
rB5j77DGdFqeBr4RGQznQcdFCTCiU35aiOvo5HwtXboPqKMp3AxrPJM797GOM7yi5cecSvemtY0K
dpNgk73j0gs2ZlLBEFimAwpAy/Obux5+7cxxkXFzIAHDLu5i0CgNgDqgLPdVt6oyVX410ojv+4jB
cujiB5B8X0a4wDQcX0TgqkHGdBvETNWHrkSlyxcAKSP227FrjpSVPtVuqZmwIUjpDmaaNrWyIg9t
/dfdqkhMKOdh84TdBtEgRuXRW53Xqs0/Hff6Iqhe5PyGFZVfodDUKwgi23OuyQEY4x7zmMtX70he
yO9CTYt8tcEWIOE3YHbE7ODyHUZxT2WNKejNkBUm5v8OVU6umAHT/o7ce+5nBytOiej8HnY2qJWS
4ax04tMa/8gnTYF0FUnUg4s7FahRPtOSsU0+6xzjJs0eoSpPvPS5HjNieuqkP1I7684oxgR2lA/0
P2QbDtb0R6erpKmPTtjTnOkuKc89tfyMA/0iHqnpqIDtf6+EGoKvHMD91W06z5KjN2qOtyh4ZR68
CZbFTjYfVt+9mg/jEFuORFCc7iFE0o4CR8U5WmBCvHja2ESRhXR2XKvDmCktIlQLC3E2VgNIp7qz
HqNsoOFnM6Vn313tfUX7GkSrQVTfTEY9Q1FuzVv5BGeW13Le0mdKlAouCX/i303ix+nXwSfFOGX/
uJybKgi8/aTc0rvaBo5gF2cYAKSusYzllqQ34fC4Slfu7XWz2GgAxmuaKrC5m+7BwnKUNiEWJ0Zg
X8ON6qJUMlT/0kiF051AOlDmxGMfuIzA482YqBIFk0LPv8zvSV0vcgPMzJ+YjxnPVoew30Lo+OQH
Er+9bjoaxowxMChlb2lLdcSVKNgh0tHmXrzYFz34FrUBbczcFuzTmIIQ/gMIdYgeVNLKLgzcBCm3
LF9Tt23rvr11ikGG62uPEmF9p4zgn7mCXwCD8D6DqUyUIp06+f4z832KCMFRJ9BIrkNoZPeeNVz+
xUTuTNu+q1YUVAfkfm3QQw/GxAd+/5P7azLiLqs4qdYhKax/kfEccZXNXTggtwBLKaEdwtwlLPXE
YDZ3nd0gT6nw5nNVipy42/0o6ftJKHzMMgsNA123dSNrK3e9a//KIv7cZpgMjegFFbG9mKHkFmZS
WuqkDs5423gF1xEaW9xMVLg4xIcoqVkZB+sMcowr85nbNNpfBCgtjZBjQiBDiLl1Eenv4G+gmZ/z
/sBrGbkxAzYFAxcDcgGa5hkhKXfNaBgl7KCroJB9JMhZGSwBeKlxoLJAe46iehwUa3m+a2UDjFDL
EHOkRQ4dlI0+CCUul8Ni8GRX7lwGwlOs2fmhqUOXcUgmz1JZe9QgQ428/eGr3juYTDOf/XTFo+lL
QIvQl61AX0xIcbiOKp8htLCIXIuoaPv0jHAwcrjzPmCJ4HGw41BWp8GbC/y0F+XzVz1Gjy3yIjnn
Lx6j4w+9j65TE7EjxMGnOvD9lA9Pfbq31n3iG7FR84tNKtfbH408f//Rijf/6Q5kPD8xBnSHBKqO
WiYZ6vwmNtqB+2ccvVX3NwZJ2BpRTAZO6zMAoPGY26gn4nmYQpnne6uOQKR02572ldDlB+6Jotbf
rt0WioNUJLmMEIab4HQ8VN5Bq3qM6AptIXTRNU5bxqTg6yfneh7HwZUSiUkqjUwre4Xl6T4/2rX9
GfaLpXq//rLfHvo0DsBNwdeemckN8FH+4L71dGtHecBsyDVFOqP6aS02S5Ja9J3RX13KmBDg19Jz
ZPs98RuIi9OuAqo4rGT5cAdIYlPYRUJp/uMJOET02eLf7dApPtC3eUd0w5hflNS4dpZ/GtVE2YBW
rEZl7LGBGnDDpij7GVjHl9mCRIgndnOdjyFwBDadYbiF8PWDv8e3ITfPS8Sjx+K9CtryjuEPzRhE
UfNlMQYVbjrykOc5U544QZmD0yPxGj/z97FH3g2WTe6uNpTLSu/0Bp8+3RLROlN6G7ILMJWlOJyE
Ho4bv3IGS9HEv725lofVQq/YCZY/a3qmOQF3PSzQzga3qGvUu0sncNKiODGwUNGYBegIw/QhF5ix
l8JXeOai9iwYvQqY9eaU/BQVilc4mv0FSf0tiSQ09E61KX2rbBVKzxXVnBZJDeZu1U5uQU8wbH2M
szB8DStyXEEwPW5JQ08IVSUG3BApmgVFa+1MNMjtWO6huanRRDLgdDXExv0zahBBPqQToy31FvjH
26KGpgmJgRfj1wyYApSEzYS4T8zuGI7lPAQFZ9jxWSquA24KSQ75SlT7lAmfSdHyTmXt5V9eV6cM
kvTLRa3HiSh1E9psRxDZs1/dJ12r0A9FS/ZATNNTZdhNCwJ/U39B+rfcVdHzTCEFNiLBEGOepQJo
p2L1mB4VlGpdIBEVjge4d6nesy2gYy0jROCIugHOuDF6dRdplPJ2rxDH0G1ikZysIr6rvbc0ZVHR
+spU53h5NuN4VR5URJ9Ju3peBOPzyjiF/IZEH+rdHqajjsmjKJcoSml+9haJFvWpGylyLDz0lAkh
A5no5F1Du3/kpxjWRkNe2kB8A1YevmctgMJAChQkjsMHDaHucqq0gUQ1HJdFhnIL/g5xfd2ZTGrY
3ouuoDczOXMVKco4FkOTicrnole19xy3dGCRS2qZ74xS6N7BgJrzPxcHx8AiN1EFoLIhKekTh2w/
3Kg+b18RdgIB03zCzT8RC0+O1d5iB1PlC3Q/ZB1GF0N4vN8g8LG33El4CAwPhaKJAfOAto+fXwMB
gHVFaW3xGr3D6776xVQB+OBbMHZHv1eJiY4+ac8Nly7dlrGqQEAQyLJ/eyjRX7z4DQCa8nmAQEUg
NyYb+AR6OClnoV/U1PrjKk4Epuel/V6sCsxARhxJLLxTqJVHIxchmyfGCxQxysTUpc6SfAtzwh7r
R0pitkHOPthnh/SfaWb6+g4wiRApgswkoINvpPcDS+FPntgDaZDwJKIcuK0wP3rmTdX5OUtzm2Zd
Ho0ioUXZ+KPAUBNbFYsAwnsnGSPMlmnsF1zaJ+onuXSlt5YT9tFW+kjCrxJmALlfKMjPzzJugrzL
NYqINDN0ll6GjFakIFx6S/sySDAqWSyvSQChqDUZPsglKF6Ck6Z471z73oZbuIyzcd6V81m61FBy
uRcvEX3cYQB49mtDe6s0jFbajIdV6AkhJwr+c3rMy9Z+kaF3rjeokJsutbPssT5JMk0I7Z3NPGDC
/l6fiWqjkWq1Ou0pafpm7cPP6ClXgAI4oXTtxn+YnTIs0v8DnTc5PWUmwh1bq752XNRKbAAFtOka
0tRY3u1v1/9MkK8EFoHMzfJhHUk3ruclcUF7ZEQcIf+ASGkYDkfqogZeEVzBSUGk0+U43bm253xB
vwQw0V0fsj8B695+fBcx1h4KISLS7wojFzfi+XMnSm6UNq1MVMd9B+DBu77f1XL8HNUX5q3EBwOt
8/fhSLdrZKaa57Oig8tYOB1If6So11SooNqvNodNKhzUqVc2Yd9ZYDYBbT54WmcYLNE4G04UXE6w
R8hrJVTOGiwxJfllEMLbybGQ22Zstc48o0PYPsfuKQWd6Cj0zbNXUzUPzfKiJ0JGMZbyumDxNkWn
AZHUCc4QAttnhrrWASvFBUael1RtmzDBSu85iovX3eu9gTTNnI5+MbxOfMdOyKCpLdedC3A778WB
zY6btnLRY2rX+LHcbKFa6xAw3K9LtsQXDKmmyLlmPIVoeWl8FOnoN0U+L7FZ0caI6ooxZ0L0iJ9v
7NN/wHjxN4U3RBpwJyzvoutkw3iegvGwL4VQacTiNrbdZIJoepSYdFNJCjrb9Dj66ye7L3lj6YEA
38sCgqNssAAKSglqn7ypDXG2jn0kiz5aE0UeoXn1qH+Uf6rr0EjgjIDNWbY6lgVIRxUA4QmN2oAq
WE2ZJgHWTU/b8scBrFH+/XXYUwsjfQzty32Optr/nHueWsQUewHBF/+twYWJEqVx0WOzhc6WRCkb
nk5gjYCxbZoJ66IsPfzYvWEZ7SrQWnQIODlcCbhkd1GPxTmHtu7kV/zmR//RMX6uRBrij7lXCoMr
yulB2rfWQkQLtpS/+wS80m24F+rKnrCjLTw6Xc2kN/NobjvaOmELbj8T+HgCP9NTnHPEyjPcZAJF
QbhJRc9pMFYys2EgaEXvOTV4LiEMYD+R/f7YN6vR46fS9KPb7t5Uj5nmx103uR3MC7fQjcEAA3DA
/wiOeCknI5Bzw1rMmWLicWU+hhW4HbWNfp4swPRRD3wRI+keXvZYY+yX+6VuG7IYQIUgK3yBYW4w
xv2OWp5ZMWpX+g6Up2iTnyXYwV5Q40vu1JBbfl1347xLpp4FW+AGYoS5QqgsdSCC40gcZdYvWjZN
F+ripfKGOda5p7Yo2t12FUSVRAsgG1Ly9kQj+dGS4tek10aFmcXkf1cCbo3CE8MPxSbdc5OEownt
/S+RmPMkKIJhBrXeildM3F0chcRKRpE0lX7gURls3nCYA3HNDFRypxKXEcAhTI67ZqzezNch2Qoi
yeoFdbtMpwuJtV6Vma2V624QeN24RmRqcUUCOO6BmvLczM+sJIW8HtKIRhTjRtnUi31JjKskkOCV
zGlY/e1LDJ9UNxZhxVbQCovhyHg4NuKCG5l97lFxzgzeSHt+/VIiQkFy4JOkGEiPJP2UxYvd+bJJ
NT6DaUKrDRnl3/CQyjL12rLE9AyvMVyBMXg0Ve2c4wG8VPvkaakGYZfLU6fiGdPETCXneHCcXHd2
dPCpWpXMxcGeekF0kQu2EeCjA+vIDKpx7t6j4m+IS1HEOJcDVvfGOVIGa2oI8j+OwqESgLYahVcD
yQZE09Ye44X/lguLeuSf1TNsnnIKqx15mOhMVDlYZi55ZF5gdBO9PjaZcE6I0jBflDCEWY/pTGXX
hQkr1NHycB0LI0gGF3YrGP++Su9BLqbCKSGS8BLVFzm+8G1nNNaYrr0IcV9RgDGCXz6BBXYxhMba
IYh+Kp+Z+Aiuey9LzJdQ9TlvNx/uIU3VU7EQPIFzLbSwK2A58IZ9w7+ToprcYCjWnNT/Y7z06hQr
K4340ymfUsiAYku5tlahmTaRvOYr093pTRhEE7Aj78IoqFULZdnf0jL04odKqOyCxEDN4qDniZVI
pIT0J/ykyQwyAl6G1cO4+HULLAKYoLqJjmOrIfR4rlqxloOFxzfz0pIIeGLIykYPBOKhG7ItMIpH
tJgKRD+K6aJNM1PxoEpWkW941YxgoDUgUFQzE6xbaB+il8twuBGLYKqPEPESoBSIm/mnsSpIAevP
xLhWTSJSdYUE0kCEwpZsroxeNHqefkzp11l+TH3lci3INwvNmBhQcBuclpNTLX7hAZiYzA0GLdiE
2Exw/ANmInJ5yIRFbvGIu1kxbwm2QQn+khcGaB7yU0I5MbmRPiwc5hRXSISzHzzpfQ+65tPuHEJk
QGrQ3/2OONi3OF4tiZg/EHKaCBj7qawvP4uRWOZ1FqEUKwOq6m4rzv9lPG4FmWQFyinor8hyVRoW
jDRQRUtXcFzfDx6J79UkD0t6Hvn9aVX9oeVJkpAsflHvKoc0c0HhmSI9zUZxPz6HY6fzWgzu6f2m
fXrd+6hupwP1m37uF227R5Ie2BLfvoQz8WbGbMo4PMYC0WQgoxxXlgcOmEHoNVRJBrx/cI+HCQX+
mO4LqhPtgkI21K8OxyWu1fR7a/thh4wPvuZIrHj8//pxR0ux3ZchEoiA8ic1xRkzD42abqjDK0Vc
fQJ1rQH6BmWIq7tMijDCGnOWXc+LRQqYfsf917sIPxgJ5uAB5WoEUCIeft8k1CbEFrgrlwnmiYVt
NakPb5l+nqMHAHeRg3X+zeJV92GVn9zMWJwSYmvN6ksXCds0e/PXXRnslt0UsdjFlcSv6xwGjyCW
TiViyFG1bs7hyh2YSXxwsYfXizLIGBNsllmi/AAhb1aeE9IF1cUYR0J8oQ3tUSGznYmOPtEM6VSd
F78piw44bd441gwXAGDMAA1PmyVuA66Mli5MxIsT2KCMKAaJ8I+7AQwZEI0URojSHrNZOUQVhJJ1
8+ddxyMW7mNkjEMoUkwo5W2BMubrmcuQeu/sC4RclQUSNwv/GhtCyfCA4w1ErfUjIn95lIMZgM4j
FAePmSLbuBO7HN87rMFvmLmMvv8Ag0vGgSNKxFZ9ySbyjPRkttupkgSbuVwqwfq4bwV2c0FpX91M
MCGOQjs2ok9wzMm+CU9g7+jZI0JMG2KTuoOlIAdrLTIagoE2Lbz+XuP80Meav7LogpkIUcR/wHWO
OX00OKL6SmLsdDoQSwzfVKqPCm5I/V2m1W9SsNrsTKdbkiUkWP5/4PpmXmDYVR7upxqZ5RPhuLOd
ItF0byztIY7PepJPHzvSje8D3SM/NA5PBFdWLAqWeEKXee70dFhI9zYW7mG5CJTgrz3SLZY7DjtC
NzzPNK+malAUhmeLfdIF8eVx//JWPxviadcKP1NB+cOGpVkBFcjiwGswmdpl7XgnPVV3Na8Ml1eL
757AUORLF+67irPj+dtowHRHKTXF4BschS8nTW+2SDAQdOgos7co/pIJEs+W41h85Q/GclQXwaWq
oDYXXFI9ZsS9i3ZrAIpxxGyn3w1xt+859zI7cKq5yF1Eo2ASIsIo8a9013q4Dj480DCgsTLPfn3j
Ht9r6yXJ9X5bNgtqVcvEFNm0D6JN7Q13yCjxlnv0N+jsG6DM+YkDkOkZucd6rJuS/i1gjHBxLQgk
DYidiBUwKFUaXhvaezTfTV5MfFRGUvC2kruetGSDLfz1ELemXMQC6DPn7fICHGGOjemrfiGUmLcA
NVlArDzn11Yfuy7rUpN109emck2eYUIkMdfpIUGdO+S+AiUMuuTnlQTK7fJ98AZHWBeJJ62awmzd
fXIQ4HqizjMpXqMEIGceS7EaGAtPUaJdJTeujJF9rN9SvlK3Vvuweudn57eohhgSk8Riw6oRqhEY
JzI3+chGBfasU138grsqbm7LVNz9gR7GP1mfVogL/Qg6D9VOmtd+iS5WAyivHVIEvqKokjKEL8sy
UqIu2ucuklMqS7Bf38tdPPcppM2Nmz2LoqRt2IkcmF7PPVH146mPdvPfYiNCAE+vPEGtFKGE0Vmg
8cY/TSF2RRsXgyjXDYfMgUJFxS/e6xD14fNDNE+3tHDVRSEZk5ST1cEtpKg8JRG/OjziGamG7+4N
405yGlGtkopObgTKy1voNghphPr2a9CB6zpBbYkQqQFKpIgWVn7Ho5Zvt9IdXjqD61Bft+zgCCh9
qKpfmLDKF51G0akx+3dNjdgRKCeqOo0yzuBpfyEG45PkOp8VlQ/ICuoiEWlqe+TsbLpbexHk50uy
VtEr9nNwti8zbAfZRaxpBkpUmNSypGhDDEzM+Vs5avydsX2iryOL6IGK6SAPpBVklKkekswgDQru
749HopUYkSEf/YfutYKIfiHmHwXOGkJ5pk42ciCPJpIdVFJ1wFlKzthbZv8D11ZzP5y1cxlxzJzV
Up+zZ+HYp2q2DSoOsx2qenvq70UsdRrAxrWcMSoqpyaCdBzVvKlfNnJpFV2e2SzYLfGC6cXOFv+5
jCbGi4kcgpQDLusdwyVEH7AeJ31ArWPk8C0dO/JLBz3TsjFs6I7nPKE0Dr0YyM9KWoXEnAaFJQ8m
ed0vffp8ClAGDjQWLEZKnsJ6WJn0cXQsqGYbZbNtGSjN0TPNxsEjdnc/GWZQmw0zzYoaaXIlJUd1
67Elbnd9LJyKkiZqULDbfqnc9dUNClBVjfHKP8WxBNpS8W0Ig515hCb32m9qe8BDrvHNHoRT1OxQ
qYZDNCO6TlDl5zrlH1LYLQmz2pWR1D48mBQrJe9xOuzTpCnPRPwMFV6u3ZUGo/AGxsE7GWpUAFsN
heo6iiEPLkSXcGKasqCWL6K83QGSALpkbBVyjSBjM2NEggXP2qjbLUQeMQmcieV1dOXZwe7ey+Jr
bQfCDL78tUplsq3hTNvcnEDp+zJJSnlcnQCJAoC1HpC4CpPriTjBqFvE69zT9Zhcoot6zjNmI3E3
tZSA7GVhFEu3HYET4zR/CGHUlOfwskQshOisYvNqA/YKuw5SUKNYK+Vhs86oUC0O4kEdzLzCMEey
NgFB7enc9Fl6Sp80SxbkKyw11T/nmAtSftxHvkDe1H4AN6HQ2ZkyGu29xBlZyYblIvRv7HmIXDDU
vzs6JeRcG+zuBX0w5Fm3cPqggLd/wfkldR62TWiJNRww3QR7VWpMFYRaYZHQaYJEgDrhxvclc9rG
8Yh+PlTlcXu404jkDCEG6fEa98jew29DOmZAs6uz5HofQsZjw2sESpuxRa8ytf/XhF0znjE8wH1N
A+aEWCXr0QMKSlIw1x0KbjizoNSgNWWnJZ9YPCtK1cvqbBGj8pehJ96ww3QnGGruLTCwF/1UvE0h
sSF+Rsukuxm9fSOezJZT2Uo9w0Sv0zLaoL0hYt3wvGefozyF26LsUgF+IRFegLe9Y7uTeDevqViq
1D1KhNq3kCrOi2A6I26YhllIGdbcDTI0EgDGraZOSFvm2wiESlYfgNWslRD98+gJjbaNPLeQu4yR
lspQSWf5+zVslse8OKj4192DSO93iMHdazIAnykUiubJT/fAzHJO44I5NsiIGruKpli8jOU8o/Ur
XI2gQL7xT6nJn91rBg7iUJt5zRzPdBkAIqy3QKKVU3u3qkffhzlvoFXJpWUsrC5n8ZyASq2RmlW6
DgxtSGYVsfyR7xtlsYyU9mtOZ3DteKB90YoVT3pXfG49dWLcSjmlSy1fBTiQe8ymciogCJoWytZQ
LA0Qpfg5ChXWZLjEg+/oMeSRmoeQ2omzuC/+KBkxnrg6LX+tG7r5sxlm90BgimVRIoHfJQl0Qyc7
A7PkikBVWys/Eb5Lnjl6TM2RFiqM2kleZV39GRSHpYglrC8silNFnUqT3Sg6c8svrzWeprtBF5Bd
cAEIpZ9vM3EBkbJ2HgUE48GQBm6bqhIxPU4BcZXgUsjpuFOdlCYXjN7Cwy74b8j53BHljuLQnY5T
BZR/PnsXISMe9YDsxauuz+jIzM3kBCQSZ5r8FtXXRfskesgeXaYTeC055t9EEs4awD9LAvXqubYu
EeIa+Xv7Eum0IWUoihjI4cRaxOocKlY7ynibSOuqV6ejc9EeThUB9rJQproelgM1S2N0Mg3IN/Qm
NrAtftYlkbB1YCJYKtS5Xjas984szlpS6PielnN+7v8nuy/rn72ULndo3Y2YgNMa9XyuTZiLz+ys
g84ReXNCI2NwROCpqt1wpCvaMLN/e1UqJda4Xg1Y10UbhQIbIjoIdDDCorL1Trx7risAlgd9Y2PE
DToEFy6LmTas1ofRcfqIDWb7FKrCtOpiDq/1yIkixHxD/YPB0gGDnraIFgpUSZfmPvF4GZou2/w8
LVDVnbNXIRJztgP00TaNXbWvSSe2V4iHBgAEXAi46tSgDABcaHZmCV+APnq/tj+WzBvqCMChbDHh
XqVEClvHdhZgVMcN0i1n+WhkGET2WfLSxFIVx+QXYQ2kYrtG7SxtY0kNH/gKxI/trn6F2tMu/qVT
ElANHl5gWwsu17NSm1U57aHfNU2A0DB/7yogLOBJIyxPOdH8H3pjBoXLRjmygsi+MRv9AV3kU6Y8
iW5BrQzm8HLG66WBNTmvKO1lZYmSbcWfrYENIyL0ZsL5hTYIajbpea+12oEK1cxpj+/vcD1O8WQ6
tms4D+kHBZB7hF2+ssfajBhR8LnRDTmlGK8pXRpiddYVibaI06kGl3EquLHa7n/lV6ekhwTFAQWL
PiVEv5LQbKdDBhcx/W0B6AiDdzvVh4Zsqv/+Qd3Fwjnf9LDLRWmTf0BZC3JYFZDnQ89gOKcGGQTF
iGe8i9yvu8QY81EEDav+5eFsu87Az0QhxWtiHgEgATXoXTVarJhTNgQdLB9xlARMiGPT7Gun3HA6
QIcOabfshY7VDlZa3ZuuM8b//Ko9xH8BwFzNSnebEhFxCB8lBSlqMwM6IjbNtvESKzUp8HhpVa0S
RY8Ff8zO2R0FtDGx0bHrAHe+hUztzdvWJY/GlT67bQEGKprJ6qt/ut2NmPZ+xCLxGdT5m4ocYPp9
/bH3ixgsj2GWQKFCOXMVNlrNgNbXMOltnPQygnxgQTd10Ro5r6v4+LE5YHyQUJ8R61Nac5GHmLlq
X46eCkl3ygmAQKoy6Cm6Zw/mJ7h0rWpS12iMDlkBIKOOGIT3rF/odkyvpXWo9Cr2SmEDQqDTmxbR
zibLshirCtyXuTE4J0uYozzk/k9FtcAJzvHnptZLEUkv2H+vGriXG/FVOOCUOdnXtxrXHh1dafFX
HpQkKAv4BerpCzq57qHirHzQAGnjHtCVDCGBh++a+dmXBoPhOvFKFAqzS0czK4Of1EUtAjHGKH7A
nLO0GpmLa8uHhY1eY9gNEemt1Khry4EP9TRxZNNpw3AkzekcawSgEwE0oDc3BzRRmixVb+8PhWBs
9CylCGJqCGZx51yy1CJPO+hyEDkd5ZT9V0+WuMyr+yBOou29zhBEhXaj/9MmPeN9FsANT7cmWG5r
EqZf2/9tntdmzsqNyPBAFpDoXqswDYthCl15XAbmma1Y3Vs/g6LqVtCWdY+f9YhQo05jV0YEfMFx
cZosidVCIiSCWOnKmACm8cZiSifH26Rxxw5/OlvJ9y9xjRpuEkvX7EQKoKP3RKTCx0RCd3pTxgLS
UhEGSDnTE3zwx69yiN/0cLzlPrk9z20o14MCQW5CM8D/z5cawBwQYme3cn+dfxD50sd0sEoqbHVr
NyoFYSsFlQmkXnKdC0yM0z1x383kwX9Ycn6065MciMTQH1nbCc3i7RziaF3ln1i3YkOGkAnrKh1F
AUg/k6LzsGzIwoLGzn3WVLSbMj0aOQJoQf8xaD6G6nIadDhtjlYk6VZ/BOXEU0yHIfU/hMU2B40r
snmDiTnB3sVwv7kdtAarO4PUXKCl2Ljv/N5lOvogpY0TNBe0KG2K/M4oGBTOyFSSPXkHeF8tdYxJ
XJ8Rl4nbVAdCP6BrvR8ZDJZ9+jlJtL80LZlyw2FJMEukI/T3pMMQfQYqax1Fw3bnwkje+FA7qh5I
Xu/EAyJ3DYGTddtigPLRZLCF7TZFbNOWk3OgpJPOn9K3tV0VR/0+jVsxpMWYuG8bWaMnCZ1FnJCr
4F2o+Q9zRBGt5NmLlx+t4omabbwIAbojXCDoZQCvjVZ44KcIduwCAmNZ31NvXpxlfhBHCBBIFECA
LueGDKYm8zTARS3MOSBYDhORZCPIFn0oZA6aswkU2v4hNNgDYoI5FgM8eHCfGFeQZgYjGoKTxWQz
vQc67jjrafTGQ7TQNgedETpyOdmTevHuN8TZedCWI/BHAGGczkivPB+YsB8NCe/hl0gOwILvH+76
3xBMXsN6c/85l7NiWeBPJJ7k9MnLnSDHxazoJTTGXIFlGjF8sihQmKiURcf40e6harla00cu+Lyh
E8os/MSeL46Rg3SynMo5FvwXHxLQkdk8nc3n7h5+9o5etOMaSiXwLyWWJOehM1iqN1eQnK5vRmrv
ib9pL5Xo/QKSHUQoolZ1OSM2ok+5imlpDLpPfijI9lHJkhEtH/l9MWHRgN6Dq3Kz89AZ9R5e2yPc
fvGArz3paSWN7htqaqZLSXlFRFl9lV784ly5x+UGDIu2NRIpzcT40Jf48zN0fc9WE1NA2WHOT4i9
Wynimv9kL3KscmcKnj1gbPU/doy7839ESJ4kYS6FvlZTtu8XQLMkHan9kuPXlWFWR4NbHUd2GopH
ZhQgtKjaJDzdOw6JLB0SMjY6GPvA+WnCQrW7rrz9RFTNFUT1YFIWnAQk5p+sNrlfRjZrlCOXrCZM
zfytX6To3MneShVP3CDrwbI1ELBv0NVqNql9WH0m/nXsb22Wq1dD1ylwTZTZdxliI71AH5PJAYyM
q5W1H2J0ZAthXjMuPAyErFKocCe2WE3aJZGaiwZJsbMBz70a3hwFXJg04L72JTRv7a6In5zQJy5R
amqrKJy0ANoZvoSnIVBKzOau7o+V/tNRmdzezy5OJ6EQozRYWIeE6SHWBUdBQFdm+NoqsCxxpMjc
KX+egIMnwALVcy+6Yc7G9GQM3c4r/bTjTvY5a8jM28l5SW1hAHr79Lv2UrnAXiY23sWc8VlNbUry
9CpV9TakRCpgmeglcC8rBepr5t17fGY5dB1fpa0BdX4Qh3Ji7hxSpDg943n9U3IZHMxTjOQu+k7u
494zX5pIl0bArDqqFWwmshrmka5UtVp9unHiMzAosZS+OfP1KH4hWeNzNkQxsxwwQHCSxlULiQo8
CboGEcbfncd0heJLCm4oRuu0EJnL+fhReKqxNoMkJqt+YfT55S5GosaI2tGmgGqvr0QY4drGuYxD
wOzJwnJKUrC32NCtz8rmkWZA6MVPik4+Hv2EN7cgJwQa7KVHwQGKx9vTe4GVZAJMqnvEH3/I9B43
+IHKfZeAqUvnmky6uXj87ILUt5JWCEd9fGVR2dBhS5GsdRWT+lo9dV3ymBBCjsXoP4BODtQTdtfN
YLMMYhQo5dN67WU/slIBsf91TFrnibzSj0cTci/sE+zAzhPwKEuRnl4j2atCClPs0GLmjRkLsEvG
kXy5wJ8JuozWXLLB/oRUNsJs/bUVd5s+sZ44RtyjfKnsApj8qPxbSeo2ml8oT4xeauCG+l2LGsui
2TJJB55boV5d4IgQtPlKDy0M4haPCyM/wtzK1f1vO/GRAgg1xs332ZN0pk8nsaYL7iyjVdd4w5Fg
VCq3DwPf3u/kLzEhZXLzXTyNGGV6mou95l+mT9pYANsQSfg0Jl42WezKw9h210W24r4+Ghj4hTL8
kIy6t0/aj4NzzXxnA6+vIztQP4/C5UJ0fJNYmFWfHcxX9VfensG2tUWJ3HFm8F7c7nWSDUOgqAXx
90zeY5MoDTqz/meTjBhae4Kmg5T1QsVDkBToMA0h8rWcVS+HplIN1KKhjjjDen0FHSddHs0k2bn3
YRHAleXEo1X+7sCTr5j+l40MpoqxEC+/cdVXhgFBEslB+6M5g+MJNE3f8KQPpq7hiVd5WZXcXrBc
S5bprRHOHFbed8b/vxBRRlmF47LthSYhhaghU7fs6FeZacVtHc1lfrqnGS570/9AJ8emapHYOYe/
IZpBsdJfJqkMukiq/uwd8Bjk3VsWynHWTlnmJuoPnmcY4UHNPOcFRoMJr46zKCWoZ9NpAA32nk1Y
wCNw8GENsiY0tq/Ar/idJs8S+8sOGymfolAFRiZUsMSKoUrcNRPgRm5vjeoVPcJT9XZGQzQZl0zo
DIIistHA3+5Bz3r1T1iXrdk4MjVluDZW7MhAFDP+BkyeU4ynOGKqjKTW8LgbBGRLxWLW16rlUzHn
SAxXIXlK5/L20krcLN1Rldy1bwnkAUqEgDcpwtkxLQ4QSyqwocG2Db98T8R/c0Ps6k7abroCXcTs
MBaYNScVU7krbeCyHDL5ScjoN2PMwFbY+BwJYNR0jDw0bI4jRBglG5XMbT3y+hJJHaDRatuINEKe
wxGw0G6lPqLszkQYf/UOIL+UyC2Z7p1raK3Fufxm9ibwL9a7IGJZQ2aufDmEJ+4TqNpA8fV/M8Hg
OeZKXv5+uxN4WVowQ644R+26TuNhN3MnqBykVe+ybWLSqTEREDQm55iuhzrh7AmNzIwBgPnjkfCo
y9uoOgLDC+3kW0bf6mRzbu7OyYAr5LhRFFojmWjSuhoA7T+8CFuZywxgHCyVF7tgdp3fNwfgPGtR
JSkC0eA3WFWmmFa/OYDWwH3dZiC1+bBATdt0wpWIMtNqUrqgFe/uV1OQDBE5xigvThZsaBqprRIp
WlMqrSIGkn9YGWJgmm5D3osY1ySOxbE+7bDSNNWDRpyBoPNIkwxDUPZPClz15zeE+7JDHgmh85fH
Qg820/dkN6W68gaOWvzsJnAsYMiPXfxUIr03I+z67F01P+qVqCkU5SlTIRTg2VYz6Yr5W4Z9X+p7
LRAgdCuIrZHPPFRsfnUXHK9mRbWKAx66XXTrYcCwWnAbevJ54/35hSc9yFcd4Id491A9NJEH7yvd
vCJTsKglGJD25J/TYDmFUVkPUtc8u6m4uwaWcWaQYka6W9X6WTwVAno3VS+s9Mqo54a+0vZYY+J2
BkZGY/oVeggPuKY3KNtqnGE1uzYUonFDmdARbUC9KBTwFLuJZDDPthY8fOUaWCxsN37vUT8KPIHU
VJ1nP/qnZAEYpoTcFb4WFMHdKuiRrvKo99+pmqmK3fk3Yt3yFPVJ1m14w2CajpkYZfkQTgmwviko
oF0ECtOGS0Yi/TO3eyls2p3JIx9PDVcTktWT2z4DyqXlvn5thuBkmhP5K51i4MacrA0kE5L2xq7X
F9ybibVOc/3ov4Sogr7eutnesOYZtSheKJSCqYTbKJk2wFkCZsmike0bAimkCaavrC8A79vHFms7
4ggfOAxuDT600vqlHHdRH4WpiF9vKolifdQbQ7F3QkwBiJLB3YIb0pVYFZKKCk9DdxTTbpXF1kA5
2UN2V6enugoFORGZwQQ4ik7qLh70J2OMDJkzK0C9o/SYfzh8VyXLeCzWtrZnvJdkDhrpvETKSbKV
cO8Fy9h+o5weLL17r97EbukHJqgq8+uFm2U3oehwIdVkYFVoC6r8xWCQJrnIXCETvk40Raep2Ixq
DIdjYCp2zCvDnM/YreBsnBi8c2JOSlGJPaM6lE4iVG8zxQEYGengSpz5qp1p7PXEYMB0OzE8q1T8
zutg7rWUCrAEv67gspmc+3qM7koGpzKCk/SBkfTYQi6xvstpy0DS6XIBf1R2hczAXQ2bf1HwoB8n
vSTZRuDpvIqTflZn8dydHWzbYbgb6qxmhbetZNPv33kDMQxNz92x41ySDnz+3MlOVrrgwOIcYSXs
hUIhfb43z+knPL3nRufION9vR9oMTh4AOBVwaojdDn7WHlnzO9VLQICsXPWa3GSqA7ebb4yGE9j0
VEXu6J/FECvr4NDoHuHk2+y9jzePy198ZRFpuSHqqYl2yU9Ryc0rmYvxt52HsNpohzseWtk7rKpf
1qjXQEsNiGMHJjqmg5hqcSgndkUGit83046jjDD3wNmXfHVB4J45N0LZfOcDCirc8svVPvIekFNQ
9b0wLdTmv1Pcx0Nl22/Fts0JXmuiOShn4LAWlb2/Oe1O/tj4M3acqMTxKRzLOqouuwBAFV/6Zc0l
Dl7aawstYq4GtN4Xyt/MDke9aeAsz2CQX6aGvixzjly6p9/nftIzDoZ4hoCQAWRm2HuxCMVA5IUH
Dk29tMMLubyXfh6xJFcapMXqymH88zYpibdAtB68NhO54/8dA2+OHlKt1yzbmhl/1LVEKbfmJYF6
WCWZElvlhsC+tahXvPgXETt7vhGP8sZiCepzqucM5QIh9bMYFnI1YWRm2hXhamhTzUC8dCy/8Fl0
3MiYtd+SLjqsMVIVJwkdDYH31XPzz8jPrkvwpjs8aBK7doZZHd9oLVon7vyWwcsaxZBXgdaqPWZ2
+0jwj27h8p6Kb0GJfPGhW/PSmLLDI50eGZgEVl6eHz0QqtZ1T/1L43Vy5JCipk+rxhHxWu4VvJG7
J1yWD1PhY72uMtzkvRudvGd4Wk0K8bugfPrejqgDYn0fVcZ7SR7h/1DBBhCenzD6ABVfSLXQm4Kb
5uWr44V6Tvgq6MT/uLFZAyFgOha4BTi8sWnewMhPYockaWYauH0SFf/mTxf2nPLob0hGK4Y2pZkv
KMHWvy6H1q//W6GTDxcwnKQ0Y47H1YeeYf7H1JkBH/PWbjdVCJae7Vp6A+ch8lYjE1BICn9e72Rv
3NVcSnr9wvu4jcEuxQf8NaMuTyK5A7qDen8IrB+qanI9/UKc90128IsdiHFf34hKwUvPVZMh37TH
UFDj6DCRdTvZydEIWIochyQqKIXPu/H+QBC49qUpqk+f+NPzMp4u5MhLmetflJeaglnK+Rim7HKX
SLh4wP2UKzAXDI1/7npxZZ9wQgg7TMTTfOgvQIcnImS/ChB2gPJcg8u4hriVVuPo0YgJuCk+XSP7
oHJhhCKhTi9QDr0bI4HpX3Lrbyj6jou4BJtId3FEYsX64osfkD/oVi+bHQH9zGu5Yd4zTOj5jovh
N+Z9z/zadrOmhmu67bfCezYk8/b5AtWgGdyMBu1GREYj0XiNHEqaxefPcDoGWUSitxAs1PuMV0d7
iF9e76VA98uQZfxbCrRvWpdk/UhdvCiPoJCpRHJm543GgBJjalzMi/CV0OHAK1g6jruCYZ+ZYqMz
KpbSt0yIfp4YVTHbXhJsv/W6AHxt9xq8WFNj3plhPXMPAnosDRBd7CRO3ZVqK2XgiVSPUwHuLSJl
RR9rWV2Vae+oJbhMDXO5zG6dxbux7FAebmfuoGv9LFJf1MSNN3htOJiDTzh1z4FZZex5XtAxLa7u
n09Q0hxLvUncs97dMwjwwjkDLiV0dFxuQsle2AGbAO/mFUNTBK2SGfkFje8Y+FcyOwajLDi6/v5S
qmZ/vA6//VwUOsy83QNjQYn9kYnwThAQ5jdRnIKBLWQ5lZB0UP7UaSIynLTiLVMERnoLcRo9EgQG
dwQNt6K6eZ7iUwTgd3dV4L4GWqjEfkPXYkBnD09ZdroRI2a738OA6wRp45xxdUWGgJA7pxXWG2DL
BbgPXeTEGrmBBUE9ddzTdmhPA1dlmq4mQW2QM9Nr9GBNnTSxFQ+QxajLZQHdZTI63jOvtzit+1Lg
C8uPtb06tqW4ByENiTKJE+3lQ0Op627v8OHeTUoBGJcfIZiHJ6zO5nmCSD7A5xaJtwy+FlPjOINu
Z+W9wd2Yx2u/OK/UBXaZwdQXa9Ie5ejhrKbLGQPPhc/Ym4IFtCBes8e7BvskqEsuvdy2gyJFkpFk
ZCK/2UF+oTn7P9XfqmqaCiHj2SkJB06oElOUFkXq+VIon+LpNgFdUOY3ISncA0OqWnsBXF4ecGP8
R2kdW46I1UX1as2U8E2f8Uvw33pSLOQmLKc133jFVm5jP8W07g2TQnl7MlJkIxGqknUhc2uu6oly
4sfQL5Aql/5Aa+/TQeXAYXUbY2TvV0Cb4KQa9uDX040Seyi3MlfADoxzdg0RzxvhchSdThqraSEZ
h/yhpeh8W7jw+Wt2Ggi8dkgp0h4vKpz3YtovVm/OolMaZP04uPiYJnJu+tDPjoKzn7fHsxe8ld1a
jYNmxZii/ei8iY32Oxt4lKEWcnmdQX42Sgt6pNDUhgcTsxdTta1njcB4FDHVLbk5Z+GlUtFknpUk
nfkmJaks+EKmzy63AUM7Z6AX7OEP6ogp8/iUY6cLMrHHX5p0QrUuOIdKyUhP1LSSXitcoRdtZfQr
MeJiYUaM+wdupgexlIpV0fDBNI5rkDV5DntLv9f2DUo3Nzj2rFZ0Lgia9zL0fBRgxurmH2kI/q9X
/UmUcYo2CfxYCvQ04TmClUWggotbf4284FVToWkM13YWsgNVgO+KCka5RV1zgMYYBGIiK34L74z2
2rSraTnfWHaQZT/BLY1fj61kk+1aECF2QVXcy5Y/Ap+eDbxFB50TGUvHPrfKpnNNOEF9gCDd/IaP
Yoik3wq0FR6s6qgZdmg+wJi0uQgwPdKlWe7oq6GQ5EQibiW2y7uw17+jrgrd42GyxUGghamPGAGw
PK5+yLkQwvSaREEXsUYujeg84FkFpB78ym1OceaQijVY7rElQ5N8g4XI6mBChrApRfL3HldzKAO9
kBGjK8daI4gvfWY0lEAaSJnM3dqGNOKckXkeXq0NjtkTXMUhWRiWMNeKM+LxTFjoi92eqHEPWCNQ
kQ9qQgSHqfkC2mZYrRDX58U4ErWmOoafCki06KCrs5b04qHjwZXMQryXpYkiF9+jlKfkzg93Vtnc
rPxxQ4IAaJJgiC/oAM/8zEjrGoQDlkuFTBUDKJHGfZ4LKire2oE/ywyEV5TA+CC2zHW85EcdxZPs
q56mzigjCidq0t4bMN9ElfDH4JPhoaX7TdCIJBQx2mfmFBbpNJTFFu9jIpSDH/15C52Pc1Ng/taL
ZDZZc1RA50Xfvy6h8p3m3y5gv8Mct3vYGabISDip8YJrnecJCUjog6gpmLOkzLuTntOqP3kNIvwv
7e/XxlEcndNHrSiiIsoSxoyAh6UucAewIdzRYHeFRcUIem34490eO1nNCDrtWJwU1sGXxOKXsXIa
nFX+TjLh4t6Iya/WkyMyMT2cjtWB8AIf9y0hXJbnIyd4RUyaWn/4/93sVLRAzLW5jj3nwS13Y3jV
D+GWB7VuPQGlmfs1KUL7dEHkWUPvvwI36AWE7psWMc1pv+EYQi1II2lZ96sCgwhVqeDvRE1kBDC2
nbV7li3gxXOxbeH129UX92a2WFPDY1rFqqg5ydri2ApFtjx3O1tvGKZOF/6lDAhGNgWAFu17O5dG
wi4/QZ5cszA0LAydiR+tqW7MpwxKDW6U0U0iAHq6hfwDcJqST07BkIXw77DYHn8Z6F+90WoJ8P/7
/fdCrN5MMAUp+L68slUF72WlxywgPN8W2VhyBfzduvtCopnHevmLNGw2uizdDVwulOxlhKXdECE3
hHFhtXuSGCqWFv2LtsfBN3xSjLNrWkHxbTMPvQ080x97zoi4cL9gH+DskL/gZel586h/wROUaG3m
EOOmZTKmDTL8jw1Yqu9hZ9xX9bTow3IbBSBT0/xWrjRwXRLrXmw+DLBYRnBMN5zeObOm41bcVkyh
+20+0QPND6ALPWKYp0TeUOzKljPbGk8QVZXo4kjdsM6iZy1oNtdRR93t6RgI7FbwnZI+4//ag+kh
FLpTk0wVfSChW+/5GIzH1dFiJb8o6V/W7SWiBQFjjRV0fk2Ctjxana2fk3oSzjP8Bxql4FdsY+um
n3pY2jnFu8yN08s+SNoAoNJW8NlYt64RICuKu3O8TU4d3Ogpf3vsof8rKjg4rT6yPYklXMyRAV2C
9mFfwBt3kAPd9OUrFW4XgspvmndmGAOAgXLSVskG8KFyirgLtY8fwESU5lD1eTNsYowAYHKvt6gr
dBdSUbYxI6cKf4DpKNbMU8CHxyuoyjl6KjGwbkTQikD3fs8QcbD94i+RgsNO1L8FBw3Y/4cSpI1y
3ZTydh4Dw4AQqIO/qmsd5sBc4bOyrFRQ4IjQJoO1txPbbmrz1TEMV0Ciw+bYzSqqezX8AIJnL6ry
FPpwOHCkPjCcqS7W41tYjp7011tqutMAmxc8n37PKqR+hLQPdmsTPf5sl3y8bQHnu/rG4Lt5ByWp
APKb0Eo91z1xrb65f7sLs0m0ORl55AmCXKSgLHSzZoxpTG9CuvBaxTnuEu9Nm6MymBZAEcNWlx7J
J9PCDR7kLhvY8GbktxjirNIxPoMXJC0HkuJoAIYbSoa6mDXXpDCj17B6AwfDWpiDtRHstph2FKbx
06HFErvsjKj58UencLBdb9ixRp0KUs3tHh40Ak9qLqbmCu3nXZ634+GSdLcZmXUHa317QzOYciwd
xTMZI4pwE1J5YdSI7IzkV94f0PnTMq+nGF2v2FuzMQ8AZv6NFTjWglshNZHkFcU8c/cNRHEnbW5m
fivz+rEGjcupHhP6Krvpn6K/NanCQq9xu/kWzrTDoKn5oHEyvv8TvQHe9mGdL5O9yIrVjhPGS3qs
1hEHBTzhcllmI5CUqJRszc5LR340EnubvRAOAZCiASLd39bDoJa3rU0INO2OpKz8vW4sIpAupUYu
AmT4hHlQgFKepgzhUDkPO4RH76LzZZ5/VTxGkBVrFt5s0TdGapbJnr1n1wa6DTOyrK1MedNdlFcu
Qfubh0YXkg7ixthSQtB11Z9UyiPil48THxUJBiL93O4QMLGcbZltRJulVdQy0/8W7w4EU1YwrUKs
5m6U8HEI5w/8ZcYlSHm0vIOpB0K5JCrsP07TyNJ1MMuAgDOfJDhOHMAu/a+MASsmXfrBq1s03TKt
rmgYyx2S6DevrTos7odDaTcEl+ZF9/TYO/UEEJ3MXKpVEa2oaAoXGHXmzevVyR4pYY/VpuCbnYaf
nos84TW0hRl0W81W75pKuflM/GoXgPMYiVkzwQ9PS9RLbD2hwLdM2XpNW9aU39an69QJ80LI6eDv
TuswYJFDFAZyU5UU41FqY1G6sVE2CJHMLhPJNqaNjV1mB9TDSUIhqJdoktm5jh1Q+aEjXDbV5gEV
mDEcc1EMYCl9p1CJS8STvkuAMueKOiHX5U4ScocjrHcs04+cBWp9myVvYcnblNmXD2+QZtCR//2n
FkoYKsSJxA+FVw1fEXOKf+ojHn0CGXNkMh7mcbaGY01RomQAq8he3XsEjH2kgIq30tkcA36eqsFk
g8GhrbHbgXyynuGEryXi+dvqOZdmXns779pxeMpizgBFYu0zTuvJz/Z5bX2MRp6yDSjzQR3D0Gla
ghyxJOzvAWGrOYrQAh1gCW0uQVK+Kp7KkycMxPVPOpjqmBrosyMYVbglwFr1eGe0AwbbIZTysUX6
ZODlw9eaZNWz81y7XgNtOLfvRcZEyqm4FpI8gxPz2dXvyu2PMDkMU3ryaC2G11hEj4JbZZPdTv9M
1mkhzvbeSWvJCfhFQZdDHNHIQrG8S6RP2Y7ktgtlEEUCZ4cznwvXuqjdcBn2T+cwUQiIewGbsc/i
XGHyzl2QgYgdERPZSAatv0hry0oELzdE4on1CM3aw6FfUxBNG/7F/G1fEZku14nZJO85fXZbDIFi
b39I/agtz1icH3tzaqifaCm67cKQPJyqX00751khmmxkuU/rRdX0cLx5bhbuafTICnYwGQ7oSEPe
UY1XDsCsrxd6lwb9qj8YZwkTZ22MPKQMwu/gi+YSrmxDbpPU9Vd2J7OwTPIJEdWAZdfW27tPsMNb
dOdtzX8VcBCtmTjshrjMHHf1lkmX4/uS++uFnKDKpfsbueP50aDkmwThsJ641KsuqT3Ujxh5LIIh
JfyBkuh1T34WB4Qhp0oaxO+2QbdH+ZYDzkkUXv2WRzW+FXRBI6BnCpJcUEpvnE/Cbj/07Prv/JZs
AjcMiInmWfh/epF6e2DFE8oPI+/E4Fr65JmK2SMk+PGjSuj66WKA4/w8aKAZIldRe2yXqs2WcD1m
zBWM+2eohV3T0GWhkbgG3SHRsdpxcSIQTnfQbGZGb4OSXFbjIKS70KbbB28Oqbu0XVMUnuHuHK0h
AJAUx6snh7nU5x/Bui/dqhLCaF82kYCeR1CX2GpDHZun5mRaLeNt0d8BudAlVHGVQYfPj0StAtoi
Y5L0LmNxacRePhBVBhgbO1wcAQRB4S5DUh1GEOzceZ8OphBJ0btIepK+XrPtm4a7eKxB9bwQtYKz
2w34faO23zeijKBQ+A21a4Oi11Dcwj0x6fa5JOUG/rcWphOTXZrTomxMMQwc0i95cQAIGUpz90I4
heNAyeygh8zTkGPZ5a1+AzyqBbzAu1OWnGdqOsHRJR9iErqRDbeUT7Vy6pw1pIMEpVySmu6Oqikr
eRa+mjoeabmgG6zU9CgwISa5CdBQ3Q6mpFHX398TB3dYT1ju/YCkfcVPBWG+yaRPSE8oIuCdYj0f
jHez/uNAVtSkuLaaqCYh/UF8RhCFBiMDq5mGtxfSlTYzmYHw26RJKdvCEtFCLR3b1WtkfgRqcnP7
G4TLZrooNMtqt7GUIjde4iLvP06TayKdzYWTZ2aJAhu2AWEn3qASMAQVNnn3phg1Kpa0v+YXgbL3
tD2a0l6sbyS+XODTe6eZ2bhPJM1M/YEZlOmHbaURWB+nZTmN+qEquQ4B5+dB75v1CVGP5ZPVV9dC
fOtnUIgCr2rlTsvuMbwj8e/lkuwgWDF6QVYZUMihECota7gZRKBMw+8ZzkvDGJtKmHL+4vqlHZ4o
lQlXLfcVLG4St7hey7AO/tOg5eoTo7jQnt16ecWaGwTLIWv/BGjWc1b5Wxxyvjai/MU/LfNlNd8v
U1o6gKUa9Mml3EVrQ3vc3fidSIfY1FtkA8ChzAjRAZO/FJXNK1PFgWOBAeta6b2WIaPnjBliCY9b
E5D1b9WHQxRp47XXC67moWog+ry+vIQqapOyj8fKKIMBB5O3rDLOMv10L/MwgO31uKX5HHOFofSi
+dok1yUWwvH8ar61fsQnOwzCjZjvS8IVWMpux29wGK+/dV/PVvkM3Z/E2FPdZmBwgbu4ixcYRIna
pRhr9IEDzZrJA4R2V/nkk9cugGMSfgAzXGPcsp1OSLKx1HCV/QGnJEVs4fAeZEkbawefDki+ZLa0
ZBYQ86uWhY6YfoHxiTbx8yLXrv5yJ3Bz0JplD0ZEmsc2VR8M34oTd0MKwmVcU9zOXT2uip79QEzM
D0vglyuFOf41PmYCe9S58ZcYAxz8q90HTX6ZuymKplwp/xK5QTzvLI/vqwiyD5sefENK1ALkJXeS
ggG/kSyYhuYpRsTkJOTLEZET11P5sxmFebGk0EwR9QeTyO5UtujZ0NcHpXl6teUMInhL6v4H+pl3
asFCJqYCj+GxQXeYQ/vp9DRz38xSrzPSVVWkuKDMjbhXc18gGO5e4VLL9v9PQBF1Bt6xXEsmkG0x
bBZTBFoo8/VPiW2RlkO9AZHdORbNOrv8hEUaUnOzM67DJABFeNoR7boTvI+72zW8tcP2VF9yWCNK
Otx427KZbjE8aW2naffbEe26pq6peU4aXf/2BvuV0WiQEa3B/NbBMMA+pBmVpe/ZU+lCfbshThRS
wRF+MyvVAmiucI2+8D0BAuQRoQPaWkDnVGKkRfVamNliVqAUop2z7hkJO5wFTfpGN3se4MXVS6Bm
TrIwb2sFYe8m3HfdcyTKXKfEizfOES3+lijJ32yskZNaYzN8dDruNkiS65tvFuSQsdpJJ67liJa1
JDfZqrn6/8v0YVIrE7BrGr3WmqQrT11UhsAKRGLlhGbaf0DBv6rccALkR2hwNREZm0mPYBI5KWnI
o7XhQstPI1Cos7Os5bxCBwyeM8kAFhFb0/MBF1lmVFLoBmk7YoJcKXGsSoF14kvI4TfiOvRRl6R+
dMQWnOA28QRwkIxGpTnQVefqJjJxC+uPbIpojpCFDBL3DHlGnZ9LqddE3IHZBkymVKOM53X5jVVD
My4rioKVmzvOUAuwJdvJ/NFHeYFyl//VYOZJhizZt37UL70wHPxRtQQSlhEfw0CgX9XSoLgZSixW
rD8yT1eyRttKiKeoRNesl+5L3sN1C+3cXO7epO/tQkHCZtTNLKnmwGqba0XFiQQCtQYedUAfkwjh
4aV8zAC/8PHljytiQPIcjGOo54OzhC/5TJsgUz89C1J2sE5M3yycRQUo0/Vic4UgOV6AcUno+Fr7
KHuLwL0m+R3dOR5f97XpAJpWVsbh24UwL6j2l0IOJVHJ+gwJ1sciPBQfOi+PFhDneTLvY8DSKAyp
o+Tx3+6RiLiX2WZuqklAhEbEzejS2qVulf+cEJM+ymlZsq0jSX7DoYafV9togWiYykYg32HZCllQ
aCrY/PFwUUbc1uQ2IyFczq+j+4Lo2vonlMWVSb69SGp/bee836Chkoi15SIBL8JuiRNBm7L6oPqu
gq0N+WQ3AeEdyQBRmqaNSqI6j7bSkDxx87bPC7GjsrbE+AWe9KWP13UjDCTl/l35ZPHgzdH76fjP
5g3sfM/uMm4XCYzXuqLuT3z6v+bYCN3HnEm/3Xn/NnqSX4E0Bika/aVcxut+xcHfUQEbO7GajdeW
8FUBjoR6gckfcStOa6AxeAhvF4GD8zN7gM/+1A99wIAH/zEc/EWjxawe152Z8V3I9Vjh4EB5wWOt
FcTafIFB7IY9CKd8Eg35l/XlzWwpOnWCK1rB6LcZiBNvBiFSrEVaFsf0lC2uXa/LCqYyiUFf7fIe
tP0GEXhySLoSgEWO7bxfM2bR5PwU299PXBADjmK3g6knN+gNEicHq2muICHIn7dITE2sds/vxnd5
yzYHzlELMSinEyRH1+aqIv0LsRR68N8XOeQggpUX9SuBtekhMm/FaQwz/9kJwSMxbpDtiZIj4gZA
BRkIO+K2o8qaQITs5Yl/gQQ/S3Waib+KIHXM1qZB6eFXqFkaPnMaTk+AgApMvoiAmr8PIJOsqhY8
y3nbOxj9rriRDwaewZd/w6nS8mmgCYJ6hPCFxrfIKlIYfsXPWfYkaDclQSaQCcDQWN1yLoqWMjv4
zgjJD2N2jZGGMlIz2I/J6nf8+gUQRokLfMRgBrrtiqlmuRnACMQ4+VnJ/KcVv9zZphpkpxyQYOA0
u53m1WA7IXysHRFMG3ePytaaXS+YsmX9cQKbXO4NIRnmUTJi2GSVd5NF4trruZFs31RPI3qzXlEx
jTqMEEeufni+nOW9Ju6cw5cqgtn1Fzd2rg2d0z6wqX2XNUJSzRHF2BGg/rY879tA9I6qxEZSS6fM
YcwfuWleA0YqR+Nn+EhV0j63oriREZKY6vjf72NaFAtMebL+1CT9Eu742A5BRs4Agq30f2maX6yU
pCjWtfWgQZeONcLltfHt5JSNWiMq60KW3yzsdj0LcXxwZHFzTw7OigAq1Jidof4m0AuKAtTkrPBr
JTSygO8Ml4gyEtDo1ZYlDbFfKmuMf2vwkWVXIRDSe7QcYWnfxCn6sJzZg7daP6ai1bdx4MiJapWr
NGQ0MamptGTNKKEgvcviSRl1YRlEzh+zmD0p5dcfmegT4Hc/acvg7pax8SrYMjjYdYqVAZxAIZcv
5c9iZiKit8RjrMwg/JWLWxpzlRuRqk7g6aLqTl++TbUQL47C+70r2xlAPUCkyhAh0iKwwuvq+JME
1i5mawGNHHO/I1qaoqra7/8oevtA2t3JIZaRNX7cdyui9U8VvWjUxUuOPT/Ia5OKRD0qpnzWNTPf
n7q+J5tiOi39wfijiAkDmwr1wJvUvdIpI10eJozEj/CYFOHASfKsw2FXCnkUJDmyHKSiMujqud1o
51ZV9CCk78rchlmq4B5VIMZCtoy8UsEQgkw/+8x+Icl9RKnzJpsRv5BihxuNivIRXJckE9t22bg7
T2Ne1f7DIXObr26hkc83dn1dvT5yz2eL06Fos1o5wPwP9JYE6Jm9vmrMctw1gf7tMqwhOl05oHsc
hoaatwIHBB0s2u11J6perQSfnuSpQmkmYJ71D+shCuG4QPTqAYerV4y3XffQk6ofFnDWY0KMANez
h1QacmG2b4T+XEo3PWjLE5pe2XKz9boXXr19GJHenpI1PdyiTWOdicTpGHKNxS5FYFzoRfXMuoFP
NVkGcmcBsk1sYIdriAswVMukzEHpfZ+wK56HDf+lc1Irn6kgrEJElTWZWTLmTHQiq6vykaEOUH8D
EcQO5zWs6vOGq3mfZSARegySAUjisyhARP8KpDETMqce5NFMkwxEeTBQlsG4r7kMgbeYrO6NncIs
wr38PTXUEvyYEQUoYGE4Q541+8obyPbQT1Xk6kp8I3Fu+qxB70qjZPr7NASpvEV3O2uSvCT37hcm
EXr0vX+a7FSZiCJUHatij5JwKQWXX89a22G4Dg5GCkHL0/MAKhUrC+pFqlVfsYjI1GJXWRjKEzGR
1ypWTpDAyNp7tbQ7RaKXslpQBXbKOWUuNajwa1CPIAJ8ZkiVUZ5++iGpL66YoIOlI2wxZlBfOEwe
vjcu9tns2aoJmeuySke2uaTTK5GSGJH149GnH2NQfHLe8Bw6NOyYKV7XpiQ3grSEwmxUTXMEe3V7
C1k8BUv9r7AH100dRW9O2GyfUOk68Jnm3flWrux2KGa75uDk/YQKHWHgWVdIXnSM5lsp00IhUeLX
WISdC/FrQ/xnXDmYVnn8UwB4Wz1vVJTJHN13E9J715MmfR2Jw2r3RSwz6hApCeediefin6O4W36K
1UUL3kfvk4Ef7aODLSrq1W3q/ptYD/yBswZ9ksOBz2g7dbiDb0jK9ot93pKz4SZb8vahvRD1ovKV
X5ztvZ5J9jj3e5J6V+JdmJjjsXWi5x7EkDooYABdQJSI4Ub9Hf9k4ILWWsFpTrA+f1u55MreGvmk
p+KAXWUkoO+BSFEULM7NzMhvJ9CGNIqGC3QZQRBkaFPq8il6yOo23L8fOqse0Yv83/qICXZeoviP
V2iuNgt89gGwPwJLKhoPoO4Ut6YloKXcR/XSW3mBLshTAkagY540RzDSIFgORCMjFFhOVYdU+C7v
ps2Whwzss7Plzkq5skD6RP31WrzMKg4NGyZ4A4BxRL4c7qeY0MlTxXrzcwz0FSCUPXPVWCkVWs3S
66Nqb29XdRjZ/JfaBMSm5OpOOIlYQSjMji5SALnpYdyIpV4zcMTqMdipzc0T7qsH13iOYFrodCo0
gbm2kLQuwaqNrEeS8Fkkb5gbCls4XuneyRAlJAcW/mOS60UanXgOjPNDjmwvqMNs9TRZnosxEzUA
RcAJroUGx8xgn+8UnBHXFd6FSZGfi0yMBHGRw0SOvIbMIlprwl3T3zDaVMFE/3uvDv4Dnb2m7HRn
4nG52PITsOcF0O7ZXSEma37dX1ZEckcFYT36/cdR2YQYPquIj2coGmIMEpyW/qnbOcZwKSGCSzDF
MHmywqmqXVsAuiRPaN/IyEYcL6aa48Ekrvxt4AQkHtaWp5RO/7iMf9BURvIqrbjS2K2yoPFYPso8
Lze5DewLFqs/LM9cjcFvL4hwbEAGtIQqH7QyHsyJ5mE/soOn4Ma2rG8Bfe+RMI2MhB8Bn3R2/ajL
2RBt6lD8dKJcAzVQRzlrvS8QenvYetRDAAU8EYt9NskNfmKbENR8wUGs2OUE6tFBnA6u7O/ootbZ
kYK8TQiYKTPXZLLY0b+ubA9OpKXhMLba8s9L22j6F8WNEZmNPqPwZeqszMkHuf/IyiMbiTR3sOHg
UwdA1V6dI92j8VY41sJPPss/9eYotX/QEL233PSR/m2KwzzGXyK0gx1W5VYKH4QxKF4DUgnc3Q9U
KOBV2jWG8xDFGKqu7HOHUPjz/MWj/906fl3BZ7udskIXu8leebjBa9I/JZ8IecNPnIG1i5SRhpZU
5SvxPeAa/XmNTPVnpnjuWeuU0gkE25GpcFzL0bR/8R7tCkPUlKOQgTK2ziuXaBgPsXg50VaDtO8T
igDF9hmj4E+lpxnZLNLh91h0FHmGZYMnBIpcpTKp0CTa380QHyE8YRm0Qffd0zKF27YPy+ribg16
eDG/zn64QQUuCo3OYPakpZwm+qz/LqaHDoWl/HBgd2M1Uwf55wi5O0nZBCIkwwWteIeIIdhaAbA4
QrEnTAxVWQAIcAUPdg276wkBYq1tQynRS4X0qAYDkBHx+q8X0SLJHN7cvbXCPjB6mJxLsyYTRVlE
bsdQg5ykPRl08rBDTcp/60oTY6dk4PaEvH4B2whvq5CMgpShH0K3pECllPKOhPuQhWOowszcR+3q
MGSrepc5oSW7KKibHOzm9D/jfRCffqWt+Sl/mb6nHnqv/zZK5Y6gTOGhDR9espiKfIHkvR0EKtjn
ojCxpE9zVPOuwbbTVlfVAHGJnljDICxR3Qy51a+8g/y2U6ehkaG09Sfk73Kh8IHpQeABNBzoVROH
zq4qwCVQl3L3+l5ft7YPxeyFstTNkADHwC065UW98ngAfl1sC75QHZ7dq961RfEmsjblNmjc8o3p
EphhuzHHMNJxx9ruIhP0vGKBUGC5oholVjBgm5tE2axAAX2xVy3YpcnPQSX8NNAMoJnhSqoxHoD4
5/61kh+ObkepZ6mo1oY+hALd9sD/xh4jLi680pKHCQ9kEDe08zVonK8b1dHZ8zh/65m0fuXGw/I6
i/vmWmqGA123X/bKT8zniZaXuidnmu7oJ71IdUmLhZC4WIfMHsjyNa6/1XTZlCqzyHgtKLflvnXR
CoXFbfG9cclHsMDzaQPMs1PfBw5ZnUTZeAvFztSMyEFs4Zf8Xt0LTFNxM1+KNBJ3zZpBVzqBIHxu
GjL73qQ88y1gQnULxPd1XLtD3sPn0IaYjWzvr3X7aGP2AUFau0xjzT5kx74GIzfD4vqjNHZnRzET
OnEH7HKHnsvl/GGz0BJx2StO/Xv7w0SMt/2Wu5WzatIXhFsk5o8bHmu5JnG0ZCzGzVQY2i8dn61q
yo4Y7OQK6W7LdwSCBtqjGQOSGluOrs3o6ARQ0hbYu7N+bsei9E5C8fbJjh5cPYqFAU5Qo0zwAw96
YPAORD0hGzEVmkemf604O3Lh6/+r4rUiOms+rnVifxOgF/86d0dAa/gCdDCRpb5+bw4xc/QZfP5g
rApwmtubt26DErsDgGZ4k697qo5qXHY0Lmhqvv7H7Q3cywno3LTordFT8puXFjyTVWVXNhrK1UFL
nQxi46ZqsA1HhNT5K/asBU6glxDaKKS9eknyOpKz7fVeADFpwqBbvVs1MINeh+NrOLgzo5+wCgzz
xf6q3fQu9DuHxZGDdKrUbJFeNMGKzcuD2xJ2Y+/J4gc5V4NLGR1voZ7rtASNhHWfmjQyVl7vDgU6
qPCkCfU30JiePrjyPOVM/A1l3phQlkJhmiAYM68TDa8Tyd9WxxAUuWsDYK0vjpOlAFWN+EHmd2az
HYRua94e5zSwzx5lO/KBv1Ukri0+Igk+XeM+KreKlcEkcKBxBvphaPXuLVvV9lC99uTvuFw8kBn8
pofpCBf+uypuWH27csIaq3A456Pv+rbOy+CLnhHQs9uxUUgXmhs8MiG8xjwuLRoI5+wTuPvB372t
67GpzBOhhXeHPzFWIjUKImGy8/DH5ySrTyl+Es23rjAXeyqHf/dxNqe/K7WdkyF0yCSGxzL/BF3x
FeP3o9dbFPqDdp4DQU8b1D6cnOVtDKQpDaAb/6vsjkBd64wwp4nv8w2QBm57wsYIzBwDmlaDa1B9
Tcr1sPUK2zvSLMK788jEgcUNDI237ZI1CvX/JB/b1JbpnqBSTB+Bd8Ou+qNVv5uvmNB+zJO9STrD
JGtdl5+8UBjDF0iQQbmektYos7mtM5D96RrK7RI4EQjRRhOjSyO4GgcvO+izVSN5AmDVhePVn6JJ
MrRop7VvN2dXREa/JBjIzWfKFnmXjsaB/XCNCDV0GV7c9BYth9wJ7KC+zzdAG200FgN5BEhyymue
IZeU/uIVk2uOJqcKLNCNTqh7kJxVUuTUXHons7W/ktC4I64h955YWX1H+5KBfOzjjowj9u1dEjBo
Y1jsEixYL81xt1rAe92fDiA2LHp4rGy+CeE0LhOYB5n69JIEDcToHGCjq85FH8hJZosWQp+X3c/s
0qV+vZxlEXvttaf4+9KF+CCOkkU9i+3YNfZVv8QfIupPc4z8bcM/yGAm76M45FytlTbNq66QtANG
M/ZWhjfjGh1YsYvgkeh8CNUUO/Cr5b1llLODIZLLw8OO7BaHEicSRjIckcbf4JKzFl5FyyFK5NAz
Tn4c284N44e+e2e/DXvfyY2lYixSaRQ4cpySfNomvjwbMgF9kduR1B8nsFn5kH9UitGwRNGmVek/
Ty+KM9ijFYSvxS8/H+vOehlaD7K+9LyTo9Br+d7kSh57fgEAF6kIT/HfJGSKHj0MQgnFa9V2g9iF
8a/J84iigt+8LqGEGOvrU8kTjkLnh3qi+x6xiBf/I5N2NcsONTCw7j88n4dhVPjsVO8PuxIa9Ljz
lP2SUgQl+gzBc8VRsnsv/Sa9T2qCNRNNozL6EF/vdiFAA0cGWvxUmPz800H6yWRa2GmOJWkX0i93
mJYHs3xE+7n/Ss/2zKztTrCi0lc6AGVAClL/A4ibQ+w92NMzOsT6MMDSffG48cqBM4vgDq1N51O/
pRVVJMZv2GViLl2YkoDfrPlum4fdSXz6ddGpLCg+ZO7krIcQmwU7kEGa0dZFTql2Ezh/1qHIi7mI
SZpr1ZHRlc6zZRR3X+MOugT6ImzqMJ1Z5H2gfku6+IRgebnyAWaw9T1zD7sk7zt5GgEDnIaa/ydG
2YpOyD9m5RtDB7CdrII+xP0RVAJxYb72cE57J6rtCQNPTCKU+9cxz7Z40EZ4Zvz7GezkMkaVUmYG
q6EeSkVAiJrxcW08+ym8JHibe3lgJdPAaFFS1g5bwknt+uFAYoL/h1yBrs4hmtr/HxW59QperKSF
6x7YDa7aAHELZaDCsiqf1vGiUqjeMuqX6UlHXXOg11CHorbYLwC7nC08KLhcMJ7dNrHK643wCeVp
jIjaoZYarEVtyCJkhYtbRaYTLZ6Bx1Raalew6SY8RC25b6KTuzI5oMXZnIDPFUn4gauo142nZMfH
t+0MIrwLOpsmDTQkKOVzPi5N16edGJLX3z8lWsekIUaZlrrdBikmU3WeLxHFscvu22WYU34qc+fb
3sS3R6C00OT3J6HQ+ngguYeMyr83Gs1ydd8bqGMsMzGGv/q0hvxutKZwsuPZymTHUqSJjt/WoLfz
k80r7y13wTzOVV1yZPbxhuo2ShQ0mZn1mZx54SSHCctbB+xFqLeP5PrMMc0WGyOssGNB59nrVdY3
SF2oA0AOPzrUlREZw9ETz79an/me+iCQrhnWzipxRGA+zG5hxfHN10uLlkZE06AIkFBy6CE0+Igg
+P9ByrLEZRoAPEw643CDMIne996/t3hStxCQiuGiTnMX5tOXI0ATp/1PErQe5c4k3b8PWMW5yUiz
m/GbuVojSMVJ+mjyKMAW7qM4L7ivrg9rmPFAbecMhNMzVuny9hPPJmaJ5Okv1WJtiZIqFC/ckGFT
VVMw0fGbk/MMWUcYWgkqlzsNEq6Xy6YzaEpeLNlCJLawmITpCQMzEudR4KrF0yg+QT46DeeCN+rd
wUBFEHDuS6kNe/CL+flS/SNvdminx2hRf+/0N9uW7DvBwq2howTZQSsG2+SeyWSxaUSYKM1YEt+F
pMbxJngTH8KUvrPM9pU+kH9+Rx6SL7PWdeA5aZE/90/CgzAQlKwoRwMtMQRLj1k7wozEsJd21Psj
hZ9fZDLEsW6IU9GlYG7mchzhv5obZDZmOfFuvoJKP0HKaRL38gjG2kTvfYOn0EU439uQj+T14ueB
c/3xjRMVcpWMGDgU/sYBUzx393lU/XaKPD7Un6VyLbLqClHZ7crqUhK/J7U6c1sErxFeVyTAiKFI
7kxGD56KpfX9HdQDfCOkzlBrOldsxtJSY1DBJHT+XZQYs0EkbZx6AfAbPI+Se0Rz3dXfTVQoKayY
B63q1dN0UPYlh2J/fUarw1u1lJoz7lIRaIQ1rdMsn6tXIXW3WKQFDV4iSgdpK/SnPKMgbzwyfkEJ
Nf53Ioz3tq12Q5r8WA9l4Chq4gUVz7V4SpkyhVr0Fh8tsWjQp3j/TqQ6tymbTbTzXBYGmSyBK6W/
ANcHSdpCCgk7hJgbnQVlY19hDHVJH6O6bmHbQmnFdXXrveJ2strtwfhOgna5LG6CYMK52e37awhM
A0L7GaOeBb0pUbPSN5sVY6S91KazpkLIg03i0Af0uaDsTorRQWSsGRg7X3X98028nsHrSEnfdCMI
NjCFKx9ovR81e2OI/maO8rbYfnERtxwcR0B2bhXM+fxIk2gIl50sXjXE8lLieh5pSxunuVb62B/h
N+C6r/4uAYAlbmDpR3itnc0OhQuJ3tD83yrt8efe7MNQ65bJ+yrfYmYPdVGsrDxW9wPnLzNhfpzv
FyWNErTAg5swR3Pq9LKOzlLra+y8NZoz5XB7ev/bo6+5aaSaa9oCRkmZuOzUZHg1H/P82T4smG2y
4YQpvipE+Wc9XsavKRd+dqlfXCUb1lfeCUt1WgDz0IPa5CH2o0IHjURclzmhqb8wtEjSczbUvt5G
mqavqnrpu56+XPxC/QpccBDIV2bIWKSCpVVblEG6z3PMS/EVA2u08mcSSHmPBFNwt6PUspRj7NeD
mDh3rgkeiLFDVBGiZ2TOxjW7vY72fbQGc6E/SaxLUoGm6cK5IeV2HpH84i4iE5hCL4RuerQ8P25Q
YQrMmBBNCrhofK68nXdTDuXbiFPfGiVg6OdfiNc7LYedAFztimn0VQhXHvvw7zNCgIPWIWjDnTVu
o8RPvHQMlC415NAPczENvqWgkjSwh3QwdHGWv4nIU0PYkc0wbR2fwN47Bv4eF2zqmUOyPhFk0pUy
9/6WJYOdyySGPJYpmVJGvb8P8h9gAKmrVQD9HRpq1CF0T2BrEeWmuF9naue/nMgt2Xw5kzfSkBFW
sonI88NI1HhqiQ+1M7WWyK3R1ablRCFhbiBm1nH2/o84OxAgzxLnEIh3MyNOiwS09JaP7PC0ziny
WC84BtnxK0rweHNSkDheDyervCyASYzVW6DnLTY9/KUr432Avu/xkVSMHlC2PbbhPvijaJi6k8FA
d8CSY1/0rJZiN7/rLxa2ZmFx4pxmIFW/hll6g6ZG6Tem1JMBS0T2KYHNiCzAIOHpNRfSj2k1y8rJ
BXO3xNhdiN+baNEsmB+S+ELk+/U+2on/BZDOZbdXIGK03sWV0kbccQC3q9TqRhVu8Ll1LqLLEeuE
vfKrfmuza+E6W4GOzwdxdZsbcos+DEnLOUxjB1vL0loDJzyCUQt9Z0cgiLYxWOOYUzrfCPpTjNl2
6BEZlMDJ2HVihllW8OftxFHeYjo427zXwt57o5rrWnz1WL9gdLXF0UFlqYpHaWqugElE3j5YsiOK
+9A9C2+HMIcAPNzS5V5HF/mMQGOWE8yh32kHbb9sV+bWlPbToRTYFQavwZxVx5SYVBQjos1BMJny
4iKxNQWdppABJd53oNJQxf+IjPpxl1Z7kenglgjXstaWW6NoGRrHIeIaYrAXt+8ogNnURAhC9SmY
YrgHYuqyIRVBroy0R2SLJMVU90I+e4fOaJFz1zBv7qvqtnvidaRbx6CRLOaPIJgSqqHJpNszTKmG
KRkupjYgtY3XUXlqwIMNF6PXwpt9JTBO/UOCOLnErFeC2z/pmi2EFH2Fxs+eqT+0oYlaszJoEdjU
cRGlKmmj9am1ulLMmPkAnmej92CugrhRU2C6WOtHSM1hK0va3NiuSnbgZ3uChJDqbU9IpUkR+e9R
gmDPhH0VXAhhdOsyLkvV2scjFKWHeC4ZiSLg47I1CRZdqofABtYy93zvCQRC2+sFoeiAXGuXy5Qv
XLmeK9q56jIeiKcns/R6P/51kizqHL3NLkrbRB4HM+BzSPr7ic0ceWKJDTjkYdFh75ZlSf6qGo7/
oZFeU0tPCSVAeLLYP2qs85bHF6+X8hqBTpvx6DWOf4W1xPrSHKXewxWzzA6AsbroaPe0PAYerFyO
QMnRVr3tsftzEB+BBB/mhwUv2SY+M7LthpVXMsTy2wfGO0kGtSSFNeVb4fJ8QJVXTVuDhoADX+2J
itm737pf23itit3GhP9VTHf6yuWZsP38tTg2KZ4C94WdOyorgKFZuQ+ryQ23X1r7V9jfG82TEEnb
Z2LznmsKDX+lR8JjQtqo4pRIM+A/Zcdbc7edYznyC6JGz5Jodd9wQ12SbyH2Ge2UMVbzr9mV+MsD
RqMx/H8fYhSy8sYNufTS2RiQBjG5rgdpfqlRo8FXPP6Ov98Vv2YgymNzxmX6/+x1+8jo2gUwW+XZ
UCSdJ03SuYrCNT6/vH9rr21pq1llluEWQyMzNKLpJNydFFiY+7TQLB4qGolYbU+TN00JtKW2QEYy
k38PIV8RRKVmAYSCKmOTfy6SJ//I76Yej7J1/BZEoQCyGOqgSrUIXTT27VlhujlTPPxD6cT5H6r8
sVDr07OfHWXEoKoSJA3VaxmNIerHvDs75Rd8sAsBlznXMetbEqO1J5IP5V1xhJcRlFngC4cLxY+G
6AR8kpdXq4Vh1K80MYi8HvbvdmX43U9w/AGyxeFVkrr2a/RJZl7CtTtIXj8FTsfVx46n+zuvDq2O
GxmCIgrT5uvCVzlBn6Lwh0gp/DjZvT3qf0isATKuvQ918a8wggMBeswEsdYkqY4dAxqRSZJiPAH6
wczyjrRhIaER/PJmEsUovQ4ELtBc0/sXNbhMKaUchMlIZxXP7bjno3cDMcWgVsJ3d98a4Uq+I142
GMyC2Y3YodPd2G2nH4nVk2ppb/mU6OQiZBcvao+L+D8ikxUsj5HhtLr+JFz/F9yuGYs23tQ0Dk8N
4CvICChduWiVifgEgAVC6bN0X4uXWjr0c3Kmsm0v3dDRDjnVI8DtR/PApZa5PgvSTaDWB5DESzg3
p9UpDr9zJncffTNAREobFTgfk7YoP4C5UmtQr6XubGo+R8qGX3uWvfrfwCND0H2O0tXcp8W1mspi
LgqhaE3C9Er/qnqXIxbiWmXICfC9CVpFoKsskw1OBnP0p11TJQM0Ofl1xgXb2P9ARbNRNVKueHk5
Zlx9JDVTeJJEXI3KUyiQsWPZ0seEZey+C8bjUgTcP22W+JiIzdVYz9f2ARJwM7M4dT45CaGP2cwN
Mf/GKRlvQbYPpI1AwIFxu6rLXkOgACsPAve2qtOV4TzgknhwQ19Cyp0TREjeV+AKdOgmcn9O9Xkl
fR0xr5QXiIhFs/FJFJasyLChkfbYCYdEC9xAHh7Yfhsc7Y1Rk5ctsk/ORSzeKFex/xwqt2AV4EB3
BgbW5AYw6aSnXYSCEeCTi+OPqIDqxMz9AKHaQDC825Tv1GTvmRCQyuZxT/9JxazfmFTcxUaK4IRs
CXRimkYwYSJR5z8awXkY14Cl4Ceiuc6U3dhpSs3Sfpr9Fb8eLCL92Nqp4rzpHD91I7FFvuI9L2CW
yW+wK5MkkhETqNxTGJVuphAcZ2AA9uQCzVAXSjX1tn9QQ5bBrcDD0z2CaOlUzSTT4zBLtemK1ChK
ty9DUTnWqF9LgAulunAVZGiGYtN7i48P7pv0ssd30iAyhEKJ+TINmc+h0TQ7iMtkyEra8gg1xRid
BZc2NXAfX1lcMgj77B/ZWDKzGKbwn6orbsgmTEiRGAK/eAmXS4ObWVJ+gawgJ6Z1IYu3OEStWEZd
B97BbZmJ/3DrxNiydlwQTyqCNAKmyZUUetXvkpogWcPnc1Wg9FW1hDgHsHJlmCmsYr2uC2/TnQ0U
zm1AzRYcWnSXBQXWXmjV4KSMNLtQnI2Q3yG+A/SsRkwHs2I2chdCHbms27HDEwfAzxBdk+k9MqJD
F5qhw6Tf8iLK6uyF9lTpaprDdhs1fUaS4DcM5J520GjSlkzmcZ+U0B27EauoaaqRRcY0hCo4W2EO
eLWl/SYKXIZC2gE9ho0YN6uY0WF8X/yC9qIeei6to/3bSlyN7hxGLaUA3g4SUBUJiyKTsIPYkk6+
ifi+3TrKhwy0SIEx5OZh7KiBgBUGsYXwuSFQ3zNuk6Rd1MiRm2ESDuXMVAkNvQEjvt+i1iABt8RT
q94Rkrhpl5dk5FWup814w2b40hMfAr1HxL9fRkP7kfcdR+9opx1uXhULU8YZTAWXQnUIAFkXwam8
sicgOnBoNDWmWMNRvEawYld0wnOW7nW22vRFRa8DXARTrTNAvYzwZOZ9sm1aj3y7+NyC9MoNhNcQ
cTP3dnyu9FUlKzHsLJupBvFJuCSdCPUSH6iidpYIIWZGYVI3uBF2RJUisLglpuAZ4F/GjxBU4Y48
/5tuB8YO16vVfnSBCx+x15Q75e3wfMcitswPOa1VIP2RC8OrEuuaytG91boyrV5VvFI740pTo/nq
LxWaNGN0S18YPl41YksghY0mGurzOtqLtbhtQWU8LgQBvXf3RI6e8iBm4UsTMUw+pgQYftmwtG5+
YPUKYZ5d2LSgadRRf8cKjoekbmBWoTc04Lkbr5j0Q1dLy506rcPZTyc+RthbRLbt2SlMso7iWPlo
TpmW3N5/6iSe+Nr6nXc6IMIN7f8JC9dgrTkM2aabc09poM0khsclxkXQHHwcGxJndwaQyV0h+HSB
ltQjXNsygS368VshZo/t2VDbm/jbzZuDofciSeIKAKQCLAcGKHDDIUCnxyUsMDxinFFMcHYphTXj
xw3O+xZ6x4YLtCLr4/TDl6GfqReGcEi1UVvLQuLznbcQ99Z8/bEOxFVodpArY46OFWB2q6G9Xn7Q
s8ZrPxRLAsCjYtvV2NQcl4H+I3uVBAdXsUfZPxGoVp9YzLchYgoQEUab8T4VOgWeUmVcqu6tH1GJ
Q7MnEEJtIUDozrGo/k9UrL6+z7f8K6zb3ZzFYidxks+KxziRy46xfthxJ64QuNcmd5ZE+DbzV7SY
J0GasG++hwJReDrr4iu8Fckv6kFQMO2XOPpwp2P6/LMoh0jjXAOCaXYO+mcfyHKUUgIgofnpxj02
D5jwC95DQmbPtYcLMbrFNpH/u4cTtVoaftAtWOS5zX5PlTW/fLcqheMGYzzSsKC75IlxEnakVaOw
Dco+Fu7sIbkZF6Kk1YtYpNvcaqghTNkaNUqhTva8SbY7Dk4XVpeYzM4gVH2RWFjg6BqrGvuZGU8X
TwYuOstPVY5rlGMSDEbbM6MLSnrR1J/FNkR9zcNWqNLob9aX7It0REotzBwTT4pKVgt7fWDVpJr8
PdGiygONexAiwz1FJ1K6noUI5oFK6ZsFnpjsotR6PwP+SjYZCnCqlTj1g+gubBpxhFRU2v7CKlOr
AdAFieLuYdyk6CQ56PL3TzhAJQar97wnbV7jZcuSarBXs8BOtxeAsaL6p5D89cehwS3u6Rjrm3bN
udP41wMG1iKOf4NjZSiWcovQ1p6t1V8ogH9w2z4PagnBpa0XUuhyusnH5bBd3rOd6nnu8wNKFEyF
ktIlvzZgGIiRuqrFKwWUjPLNKbi9yooXSTlXwIasn28L6TED1jxFqywR8Vta6lkBbgZuQKDeG22/
SgEyDMHmp4lp9lp7rcFUZsHkS7Eix3ozosTWqXZeQcvALvXgMDFsSXgh+Bn5b55Jlu6HRHtSjZZj
dOYivrtaKf6bQ5jbS9jkmG2jmRGYmgrI8vZAWU7nSXx/1VaGHO4Q2NJkO7TPSxKq7U591tKrvEMN
kXBt3t+oCOF0mN9WP9VfSpDCrXBjsKsSOW2fcmwhlShmKd9ndU22xroDO8X8indQ1ZvQ2y4LZCDK
QKwbu3LVzDz64HjWpno1qCHW7MJbWc35ySNzg8+LyPDU0hH/yhymqnCzop/KBpN7cBlgoGFlS9r5
qKk6agHBzNBE13jWMc3ltlMzR7qsgRCgxGqIPbsX2Tycxqu//Sd2OmyJHF3VJ0Kr1fKU7P08fDjp
tbnTd1XHTn++rOkBdOsvYQyMKEK3FokzfzPI4H5BFzOe+rItP4hEHEGGP//GmeWx78UeGFVp2qDa
07tvfATDiZgYmDOQ2Ov32P6uwm1Ze9qih/ZK5Ch5bPRTKTipatISlgXiNnMr1DBl+Y4nxZ90AHLX
Kss+XNaBYVfyUclLAslDMy2SZGVUWTr6eJ1WjKSRuey+E5UMQDVmfnx7VDNyqhmFBJ3XHZ1rrfRr
rQLdlFgGBus803yoTKKJcAq4QCxExvu72ABEyBpLkjt+7+3IU2miXdQ0zD5yBcNkJfL4hbimqIBG
MCEBzou5XNcuxKTM8UUzlvWho78PLdihQq1r+bH2TemRHcwtkwi4Q/h229McJK0g7kEEu9o3MDkk
0D0BYEwjodddlDB+ivRtu3dxvXl2F8LNSnMp0kxKPe2vmqQ6XmBNmALB1cdLDbxgHj+yksLN7H+o
WIrUbaM4WO9dnbl0Jqz3tyj2ztKJ1GRFF/c23EhmKx7Fhepa40kFBF28bxRStoilcOqbwEUvSJ21
zsiA6U1aNPzcasz4ZjGk2rXqttAVjb8576x0Gq/c09X4qlO5NYsNyQuGgSsfDw2Cyzs/a6DN4c/o
hmuaLfhVLQZWdCb9aUND47vG/gKmKY5SuNV0VlrFAVNUXW22VuTzjacge1omw8inXPYrKKERwhEk
HpyIIOm/DJOgdlfdIc9rec7y1Ng+WJQD19LlP+VjlVuZ4wY9GnKF6/4bT6Jk5P30g9QqpoK1t4jD
qaDklsfgH2J29MBisgU0yc6KF3/pvKVus8/8BsLrsG5pXPXRljvEF432ypldxCB/DiZOnNUvXF84
s8E/gpHCo68UnGwnNjAdEpgDrdBHUhMDf/U07bUpy/cRqRrQB6HL76/SQ2SGBSAHcg/FHztlZZ5Y
KCh7+7bFUgKLHl22+oN2XXAq5u/cGXxTVF1LWaZfSEKBkjTM3QskUp52EhOZ1fRZ0xrri7tLc4WU
7bSyRmVCLbzmj5YYuSq8qavT03mzlvnK6h1k3D1s6oKZHdZ3iEx/IQIK3UUXYhgMKCBiP6zF+Z+F
gezcz7SNKMXyyukfR02atqURJJ6kF4n6cya/u2S8rqFxWaYypmXkOGW6+1nW9b6J9z4+sTawJyFb
LUIjXXnItgm3xQ/dmdyw1kqaEnx82VaN5TzYS3owRhxwjtH/f9DyR+jmgNXbcSm9rsFcKvt0zgxi
c1s1vHcxs11hl50h3X5zQljXW2kOGZNUbfmvsDc2P+8te+LIAL545aIr4LvhgfFtgubpBIZyDw6w
bO7QkfVLh96q52kC7DcIjbLNtV6gUVPJJCH17IvKERNPDzsHFb83UY2i/LjcPNss8lu1Nv/ovM2v
jcsI1KcFCYhJaqdorn73g1pJYCyp/V8hqk98GsnHVBed6/QKmovxumIx4kbsu1sP0jmEscCav8Mp
t6KXIXVFbjgOYttJot2PG23RL2SJLRhpcoA7yb1MMSNQPeOavKVvv2KQZZwRfVegpJTBdK+dU5Vg
dFq1KXL3LhwxTYkq83wTZBMsBxw395i0LFdkz998fa82ZQZg3zdutDWfWDsXgD+DZN0tA/lrJfn9
ct4KQUW6X0b1zsQoSS4qFGzCZ9wf/Ad0gBabsTPwHCcsFtVlT8dTEziCsAgl5rjjTsezeQ7NTZ60
K9YGxRat/XFz/QnBpsSBxv1/ApDdgvpDFrFUuma/w34qKWLLwsrsm+MfMgL9YzlcrjaXuE7nHKsM
I4o+/4MlpWrGrpl8WobHixn9ty7GxRsdtBoUb/M15XIXhGaZuaSRdu0zjEbBO+9lnrGCmImPDp5f
GuwlrUl62h2y/lao3ZXO/AXy3JfpqOjXkH6l6pxybzxlyKLuwCUlGCib3bs28XPc5Qnok3QN/Ztc
eBN9kII57VRDvVmwffqdrW1EZHMBtFNYbBQUMu9raAKmD+eV3PKxD4Xl3gb3XICctjLMoybSQbU2
0YXB34vnc99N90hJqDxDS1JaJnUJ4PYUFr/nHOEtQDBPfzy2l9oWOG2MXyoHYsJoArNrkqUiquZC
edLdq4QyNQ+2uU99vEuyZG9JucHpIcZmkgkXnpKRyW37FrtpLoBTB3HX2jZCSA9STUUTX8kG+UCa
rNNH7DAB2GD4hgtPPKyU/ICDAWGaDA48HpO9UjXA63GEC2gI8SuGZPJvSbAOVxi8K6lCfUZMXhon
0nPdtxJAsy9qArPzldQyj4NE3IS3hTq1XfttpnoPMYX1H3Zqq+dkWkJKNNOqcEtlrlhLIma/Z+y1
fX0wQmUbHfSw7Yp07u1fNAUpEOQp12pMETR6oT1ltk+oxQx4F4LAmRmz0L0BZcB/LQXpjlLF0ag3
VPQM2L4Dr1D/WM+5NJ6Uf3K4BtQUEIVcfv5M3DNlJv6+7d8Fbak7Ifzx+sXMzuOZr1gSwF+fj22Z
JrNnixTvCCfJnZbpOZn//O01Fa4DbHMzSAY5qq02X/gonFiT2Q5A7VipmOBm6VfScp0EYpsfFX4G
d2Sysml6lB69w+BynIm2tCBabVhreNbcJ27PFky/JB7WOIN6ysnip45SJ7zOUBYfZ7MYWidGr9um
eZnAbv4Balj2uJj+oL3BbzrklTGPtS4AWhho3eO9NDGIGCMQFfVYFfjHRfG6C/NnLdD5/1Wb/dVQ
2lwfFQKCM2xiGnns5blfIQ9ZKQZVh2bB4jSSSglC/FTLTGamch8tFSJ2KRfIZ86UOIzUZSGfTXW/
QVQdMZTLQU2f0o34JQqxT83MU13egB6+vG77lxKCSamRmZYTjSHO6U222BOWXwBeR0trM2u15Zto
VuTI/f03bRsqV8Ygl2N9sg1+MYSMVSF0GU7zpVZj2/+n5KjnrmNXQMXH2Ob7Gk5uV8L2s3n15dJU
MpLPkzkiflNj7FvUkJODrpwPwsIDD+q+RpZmeEKC3c33ohGXt7tAJ9XlvlzCIx/oFRzfU+Jl6eJW
UZgSFbJo5zFO/qlgwHkFW8SRZeJSMgLb4tzaOctTx9fNGsAdm9B006VVgK9V6D/m3qpb6JcZyGbx
DzO/BQvvDmj+gpysa5FbfxA8OQidjcz39L/s5jQDHyJKg0xZFh9O+CsV2aELxOWmN42WREd1FiSW
4s7JQZNljm7xRUjQtxnGUWdhg3JcR/QUjcE3WXbju3NyKBsbMgPZBpUOHCSoF/rAR5bZaNuDXMsa
OcxKiLqA/yErtnnHcxGRLBSuRPuVikJ/OKnurFllRNj22VvlXeuj+PO+ZU+4/YAE/FdkByK9p6gi
REX4jRQmxLw++p0mtGtflgb0KKVz7+XcjvIGiwjsQoKdgWqy6Dyyt59xytYGGl9ztwzWLPhqUwjy
bPUygJnQVN6rYrK7LZSQZcAfLMkMm4ikL4cwmoQZ/rGsHLGyZ6GAmh/q3S2Y3GNxTz5F3SHPcJl4
GoPIB1Ww0YoBwsziSTM4IOehpR/pTAIodwEKzh7AgJhiTwdW/v0LJ0gMnozKJHL5Yjeyi6L5xluk
BiDpsSej1ow+kS208Nw/4u/FK+GN72V5b38fcLuE4hqI/z2NsT3bzIYtl+FY6JvnHlr3xjvkSXyE
UvsyLzT+/cdSR0ZOrNz1nKAsnrXX7nUnjaEeCkvpbq1aIQfH+F8gTP6w7PdAoEkU5XSqKe6RoLsw
yNY04jc5iCJ6V9FSp3p5bZouJU+5XyJCWdZnOV1MsIWypOLdfmVJvmhS5mk9jmC6PIu29zkzSwwE
5MZZJwjoLJDGDFeBKhHs+f3zt04x4A1iylUOYx6p2mnTsEu339RwIf8caPjooGIWxjw3yFc1gwcS
6HVWSOZm5Q9hswHTzhfFXVf52LQN7nv9z2kVDWEZQ+8q1STp8GGrnLD5QOL0ElNPTV3OnIDSP1Kq
RoSxdTqQFQzdchbFVvSrfauFQ784bjmYU/MYUUuZ4w7E1R0TY7pEikUGS+KhzqKknjb1VKEm4z3R
nSgEEONCYWK0gNJjsZwgjyEVgZXdf1kt06tfrTkNe9VJvPZLjjoBwA2Mfkv6URpBx4PdvoHifizQ
3peoWY9uE+R2TAFLIsL+Ove81cjejXcQrswWwUtwOkP6UDnLz4OQCRtecFoPR4ud9uIUAweQd2bT
87fZrfyedXLarOmU3VfJQXtKYqb0eobvbehVEoImMAeOt0bjI4CpisQzSWIw7r1P07Tig/nG0DDR
mO35hxdBNch+s8pWFxwykTBPk7sYVUoE1pOq9DcrebisrPYJrE8Vei8JCktyhmxgYzSHcrXjTMHI
2YX1Yw/E84L5aQuWN4ndtEMSbLJNNpaa+7YD5mCqdMnDAT/eT8jKxMoSFWKuBq5jkr6bebEb2PV4
8qv36j+Qa9YOZ5tNkfWb5egtmeM6egXG8/1EDlhf0FoVSZVIgjLv0yRamqArTXXeciUdWLl2pHz+
Gou43bHRoAJnX2moEfRqt6OrqJ+9oiUoH2kDBIhCYpuUHdL0tOwWe3AYRBnT0sVfuPR8xgOYqgBM
og1QnDmY7bdONPzmgqgDk77MvlVgXMdGhDGrDcr7vu/mXobgLVTpBZYfUCF7qN2zB7aXWSOdHCm0
oLeXqos7xD1g+eV0QTsh5hMD3njcRwoZHa/6+D/599O7ES3CbArB0eUyxqk6aGlOwpfeobV7bwZO
Vc2ozTypWwmcVBreNoDJzbA7zCF9GlESZuJGNH4shHXQRQ1YJriIPtD0bFzDtk1Qzf4gOxJsPQjT
wkj5Bht6yBKKkuw48USCHFvbzTlR+MpwWjTwp1D/Xg01rIRKjgHnxFUqblGf7Z2cjPFN54BU4Mmj
DwfQV0/iJvuRax+6lFE7Wx36VxpSwN1CCqZono7iEjFxLw73h7m0kdf3Zo9xMVnoUl/A8cwbSStt
//NsKm3Ei63Vz6AySDZydK9QEZp59N2D8KndGskq0IWejauvGzBUxRCIhBVQPNZGZGi7kG2X0iLS
eAIOquz1Ew49VDLUqxi/GZlRevEhJvr6KC+0R3KPAJXOMLKprRkaMAcFVyanGUXLKWa3cyTcobeo
SHudFLyjuBLYQ+ocxUakcUunS2bRqZd7Zvp4gmGUM7bAmL6+gp2ENK7ZEr3+cdVj9NZfwIJJmyJp
i/B5CVODAcjnRuJMzX5dB4Xgj3YXHjgSmk7zU5DOBUl9JyBtnauJnBcJ82kDuCYuLVzPvXmoAxq8
NZgSSv7MVdG/aU2D4y1AE6r/t8A064vqu3O6QQY6wOnmgVIkgLhgK8P9svyitMZQcHG8PCcRUXDx
XJkuSwGDq3e71NcIoQhaWtZM5wbEV00FKe7v+5rNqRyoveKDM2Yncyzm0J8ZV1YOGxyx9QVPGHJC
Lvej6bf2RP5muxW1wnKR1MUVM+UvgDPaY1rXFoPkSEMmzCRIYU22VTqer7MJUNljoABIGTYtS3nl
bu0/yJNGBAAU4juYmpipylSnOswsivuJBC0VxTUqsQ/2Pf+hEvJtjRMz3iwkQELOxYNIqBQTwcsF
+gujWpx9hQpAOsJOwL0RIJNyRZvsZVaVW/3EnrFlphyDVi8bnWg5bcvJ4VUUNl0pf7rNw7wnMjNG
ME2X4RqceM9nN1159U+d/Ub182oGRURZwRx4Wa3/jJfrYVDPguwa/0wjHv2UVcBaPsnoA3PzVBjv
JKtwErWUjb3FqY5TmQzUW0y+Tc1UbwvDcFYEptyDJuAyiAJiovqGpSEe3O4nk+LFr3OvVUokJ6+w
z7MDB4ktryAPyNJSJi6WsvOk/iNIkANntudw6001s4p8m1H6wfhNyqyKs1hOGFY0a0LFF5wix2BC
2v01aCsqGW++fyJgv0F9M3L/4XtFMmiHMBiskjvIzhRelx6gcfWwKoEZgu8mx64LKrBN45hElF18
mOZSaIwRQUTLrtclehyIFsqK0sllH/gYNkeAVQt2K/3T5xj3UvHWGBfyabG1peQV3dI1IboCLgRG
g9Ih0BE27GxXferprheKnuGUClWTzgjmTrqZ0RoD/KDOTtYTk1PjJhh2kKkGr59nq2bO/K/FYrTB
/zQ8BduAxRx2HzRMhiqBdWJqi92MVWqaiGDXvcIISj72JAScHEgUKpkPvNNJ2TbFauCWGajX0J4p
+PGEmj+CNyXYa99qbxUuelMM7Pn1eNh9i4Cjxoa1PGxs2YypvmCjnMJ6JHLF7da2Du5+sg9YxKNx
c+mq307w9yi+5+4l9ber5MKd5u38HBJZhKTZ4kRz0Jxw53X2HCT7QdCTFE744/zXxBPrzDOV8XdR
gGTgNwqkSKdcqVr3YtNeeh5FeaqtqCflXSCNEmVaAj+ufIlMoSGt6X4CSL+Xdn+I+0n/ze9txFBK
DCHSXZS0Lbo0P/t/6wy8PH2I2OvM2gLEQT2GZA7m8QRS/kPaxLXpbTdQrw9VhdaplyV4On2CEqCh
R8pTz3s2BqtchexA+sHfoqMpIKE6/npye+Yek1dODzlO4/9XDkmfoPBzj/8PZ/nf40wxZuAS3FCq
vj5DYuAg+2ZiRadDeMhLp9CQYU6ORyX8KJEHsqpSj9UQWTz+yWuRlbHhGXextsi7s9rujlBakaQq
T8sDZAotY3RKwd7Vs9jAcHLqfE2OUhU3nxsG+r4+yz6Qaz3Q2NwabMrvE4YV3HauVeStl67bECEh
kb7rHI21nLvs8WodwErRzJ+SHVXJpnFTFmbr8q0YsfweFISjNEuhhkMuX2/umfK51KU4vYf/hU7L
YMlvm23/zvXA8GecbRDMus8or31HYY+p1eywQRIqcBv4mndL5QgyZysp3NeluCwexuTTJtVq4Soe
eCiTQuhRsRbIwBsFetOFpkj+p93FG0KrmaBrXZXv/rxIIDXTUme1iByn6ksdeeueFKC+DxXZo99r
3X0aa9foRh8V+MBiOKzTSS1QYor8reBb+6gVXOi0t5P0l29NYaAJ5BcGVckSnRffjZF/1/V5tHto
7LgBEyIP8qOztihxIJ6oVCP3p+0K/uaa/fl5uLQqtkHEQCT6r7wNhAR4IdRzTDni8k19Ub4qCYmU
GzlQ2doYcJTL6uC1GgtZN/7I4oe7XDHKa/xoHfmxHuVrH46UjZrTilrVf9gfxFfXgm1rZ/hVk6VG
aQT0gAZUY9g/A+9O1qiF6715vpCdXnGtdw2atdwPZRhh6/cxWrqkq4wWI4h8AeHfp96/YzHcHN2V
vW/TKsx9R4NjZLJIcHnb/JvvRUVobXT4VedfuesqAW2W7jJIDb0kXinv0pq7GxbHPhnDmiC87OBu
80RU8nW69eGCFWZkySvL7dTT6M80LRqClfz1MOOWd0TdsIzVserzGq/JX3vMO6zCREKf3j+gdVQZ
yikFiMRJHfdBy6f638WGPIY6UU6fPK247h7bq80F1LRMeNPVTce2d9+teAdVlKo0ZZwXbNgAEjYC
PKwwbdHjpF46bl2HBxpCm8bXps73f5afqesrC/NAFU++WsJbH298NGBf3JNJQUG/NSpEB/QRb89Z
76n1EpIlFsnOy5VryQ4LDa1N/SUaxHn4Ncp2gvVAEv0iLJ+geH2CAisLl0iQEwY2dYWOcBj0Czzi
fajjbVoiN91glCq+6FerV8inN4D3Za/vkfWqBcUv/OTYMfn7If+IPFUfFZkfTWPlTwUqol/Id23/
41w+jC5Kc6dbQ8cmO6zQmhOBbeYw8DidFYyVs+RfH5AbMZtB71bDwpv06GByzIyFUMlvwkhmI9JG
dG29zAGVk2/lOF0kY4siydJCFSXaNAA6Jvo7NeccH0JVKTHYoPJwW2Gh7uLC+VC4SJXJzp0iwUms
sQLAiUVfeEGqwFBzdVA+838LP+e4ReXavon+D5vTk+yXRm7hW0OCwrufDm4vTZAKlZLgMVEqZw2D
httSjGhP5gXlvWwX6W1Khsr42URL5jgkse9pqy8K2tVQ0grTkyn5z+9MYY1cQDeI2YFcRA7Nahji
bDLVADhsnP0J+407f2c2e/+GNTEalCdWsJSLwpIEm6lY6ryY2LN1Wvcnmj84ybAf0hhkkRxPa/xA
m9F+ZVtMs7i02F2VkcjC6jlVv4sAeZVkwI+7n60/ynBHIxkKgg27tKJgJC04yvm0KauSbOYUWp38
N0G3tUVWdHVSLYbhj4rnHUZWmxKil8yooVSABpMhAcTVABDVGM3LjsdaSwRg9WaohXtz5dpw0CVX
zHKiLp/4aQ6hGrfucMHRvIn5QSUEh3Rw9dZtnmi8Gt6ziduPQ8AtE2h62tEPKVBAD6G1KLFZzpCR
qAuLxcPeuocZJwq1aybi4UgRYw+FQW4cnYHOG4764NxNVVaCKiZLdeUQG/KnMUbxJwQxnZRFSj8i
JeeQ/SgemjzWOryDUdbj0C1sRfRAS4glcOoQpkKbu8ycQLe+GPrOH0hHfM/ffoGYwtW6m5TwKU+C
9FQhBEZg4XGCDiZMGCPULhqIN1kEDKwVirpyx60QkMzWupzJtKz39e01lZB/9TKMm6ynxPWWTAlS
E4Eo2ZwOPoILd26DvD8rvqt0j4pCfmN+OFRq4SazyE9jSaoOcAVm5Fgf8AqxZJtiPdsFG3XuGeCb
U1Kaqlpdo8slHBY5E0Q300OaezIQyT5xc0wEI/DFXOauOXf28on97q5QAwOz9u7cUkLbSgfuxrQQ
uYRZqeBP9ZmtOaua0V6+e8rJiGRBRJ9yDjLutgOZy4rrfeH2Ybm7u/A/Imx+Dx5yvYn0vpzGblIu
pYP5lxEyGTygPZMSsCBNT8ACmxdjfjrz7TH29InwcIm5yj6coQbjWPrCZ6cg4xsi0XPBrCSlggYy
b0yHB4EmYBX/bUsPrd0QFBb/lnQScb1ZC1wLFArGBDcXZaOnkXtNqXMe0vqGohG5Mg/kTNipHGjB
N6/gDIIDe5CfWAgaZDSckSVi82536yV+M0gEkkdU0SPzMySEooQBmF54LApRDdbIEG5rjMk26MsE
kSPzLzfqGNso5SOm2qJLblKkGysfb8xpZVrDLPeYfndDqn0Sd0YSXso1C28G91BCZOvPDPnkiCU+
y8/SE2Z8GYAj2K4F4p2xyZpAHljX6Iw8q7Z9tyhLbWoaqG2o3QuqBUPp57LTPaP0DpTMaALs4kEj
tjcnFUCVXF/hD95BngJ+d0zT5BubcW+xf0q3vFWwyvXbeoUv2NRfE9oChrtTCR6yyA7BVRlnkIFD
Zjr5ErbczXcKFJT47WQEcU21/auSCg9nGEyOSgH9PnmJO90hXV0F33V6lktsLlwwEg62ZtGl/Eou
vCPRyCTdnSsgfP3CUw2wIKg38WjkmSG3YYi4uWt6DvF/rwX4QClEg7/ricAuPquvXBymJ2q3y9uw
hA+1dhjLmVQwD9VlvxUjeeAD2wRMH8FNdUli7YfMwUIPZbl9zpAjmDSKLbIR8YzCeB7u7HH0KmIX
tZYCoI1QgRDeStAhjGGU+q1Iqx501qHbe4OzjK/Sk5jvAEevLmp8ABrbXoqR7T8gsaP6pQSvxj4p
LAxLfbdcRY5hs7BBQHJHUPa1XBkByvxW1UoZdk/m/eMJQoSgVH9+MYCMnJl3ynNMiJYG4VEcWGgB
aFUwDAO8twi8RCDDYdxtYfORI9mbwBYtYCES1Irh4mbFsPI0j81GDCjG2Vw3MTtvlJva+2AXLVB3
FGEng9cGdh4+OQ98HkpqV7fmh91fLDeLSfVKPNzdqpP1OnAUdDecmz69KFoQJW+fl0xbhYJr52s1
uLJmidH43QCf5xdl35JC+w0fHhgUJ/ZhkyGEp4OYui2oiEaK2L6Q3qCw5lrZD35GHS1t7gq/waqi
pcEHK2Tfp4vWgrXAgjv8nPUbRXdbGc2ZW0swNZox3Q9EKBMFUQlL9fci7jRl/NnPWHSPdFSgJ6eE
oyok5To85253gX8YoE6rzlKnSyhQ4QvGUE7K1J9FuKqdJXODy8eq3oEfvgEjcbq/XIRukKm0hmDf
+C6++m40veF9HNm/bC5Sl+YRXtoegv2ie7GdeuCxZK9GTANaiOGt0SQwOQFT2kwGOlecWoLD65jY
A8zvUYvgIXJZPcsZbBkl5a2sFvsk2ic5Wi+CuXrAPoY3lv0DF9ui1pD98OwXr5QPGpxpChQp2CMp
Lou3N/rTczTdKC+m3wOlnRwKPlwbreMIPbCQx/+YcmMYAx4TkHs2ELXh7y/U2ZsgF6IKuBOOTQR0
TATV+eJ9CRg5k3BprKFRq4nKXX/jiC0UZaLYf4iZ46kNIGmy4DNoJ55UDNqLBoVpL1+TaWT6Rl6y
kqA8ygx+uo/zt7Pz+/qPWnovvcYpsak28uuj2cpmmKVDrTo80pfdKpBr7jNF25KmG1ekTT9Ineyh
bC700RjdKm9LGWnvyxiiYdqRCx2S6gcYQUH5WDwOmBsE1nFCvMqYcuKcWa1E2dDvilY2O+SFBQPK
+kZ5BigWj9FvtuNE7FVaT6q/oqPC3d//m3ZS3o5CcN74c4hQOu7C+B0DGEkyMf0hEzi6im02CQLO
JJD3obykNJ9gRCxErSMEhu1enxp+kG6EaMopVJMs/4ycP4PV6NNACaF95aKO5u9RJzR0m/J7IPgL
mk0ljKQypsgWSbPtW08MCH/4Ag19tfRUOClMQoaF6GqeDUEXKtnCVuqEYwnTAl1y54/CWu1LXXVR
+I66xydcBPZruNK8T7bStzXoT9L4HS5XlsPTDr5VvDPTkj2nNUV+etXwun7rsEmMMFsZjESKgrsc
d6mvihP+gyTXcWFhuPNjgRvlfxeZOQIWJG9r2SD7y9xluHLdcAxPfuux6GToixhhfFvQzhLSNgcI
E94HTY+Q/SJAkCYTZLZXts+DHp5KC/Jz6YHXeUGnQdMqM2gjZm4L3wZTZH7XMiuBbYzqEjyeJasM
QXAF+wZnspsk2zJ003MXadJt3F+UGv2arSwIBfrsPw3dj98D9sU2X+atODidRAftFvi/cP2pFTuV
gA/hK/S9nEWRCc85vq51FIRdJrD7Ry4zZr4Oz5//nHCUVizBCHCfni64xiEMX9NUKdx4AmCP+cBh
25JTDLmWvjBwX1ebJ6hksmKUw0/xkuvspYYHJkAwKVR5MnkGLlZyuv1zG0tAuMgduMfkjt4dAbzm
swuoJGSIaOSmihRiaK61UiJ50bilzJ3JXflIQtp088qbEazPJy3ksZgGShBGitfjh5DWAsMw1o7h
gOjCMNgjqGwZFbO5bejO+Im7J7sZc7DTC2OEQvKFae83pTn0TRhPIPt0wvy+OzQTQen+a0e+kNxH
XC7yTgEhx1AI9DaXfDzweunL4RTQFeCaSsO76JzW8Z9KYCBaDbrzMbST4IAgARIHAZWbfCtdRcao
M0rg4OsphrcMfebMJBkLVZWpdDkFFFm84svE2Q9oPNXkYgW2hosPQgOJ2eBs+I4txd567mcKyTEU
7t/EPz4FVNc7frYMxvnLnUk5yvL6TzY8+WXyhQDVm7x14uh6zHRc67ctIrnrxxdwO2PxMsy6eukF
NTZFPVMfqnO5V1FPKyN6e4LaA9EUuxYW/6sOmS6ZlEx5iKxFH9yfmSNlN0f0EtHxQm1unNLXcsU1
bOMFm+FkyYoMxQiGCHvdrMGGUE6viD5Vv0jENIK5vWzI4tI6NpuYYCvNGeIIlvNQTp1jiRK3DFqY
Tc0eRuGJ75VcBqWcGpcraQ0c5Xl4ib6o8mbdmiT/O40Bh3xOOz7tdHpxw7L/Ee5AKuvpq11uI1IP
8WVziVcX1JlKSEJSM+W34An0XlRM8QjpaVqHik1eBAvaCaXVl5iYVTeB35p+P2qHWW8I2+/XjO7F
nzTEYpF3EIPgzogr7AOQdeOO4P2iRTVfpF1yV+w68zRnZTSFASyb60XjlSJUX1z5EN1F/j9a8FqQ
ip7HIDeKqdKxovGzKz8PuO/3bz7jMk1hbQsKckc23rETDxLS9hx656ok4IfDMODPEYtoP+uRVPpq
zofvcnaiAB2rnPpJqsL5HrJyxlPtJr2r7kNVGd1ogdTva8UIeKucg9NwgJ262gqyNphsWG8Kiqay
n52sC3j341qy6Ki8IR4D95AFL0k6IYeuzukUKU2b5Wxb1bNK3fF7ojNLfoYxVcldYWXCXt0uvUAd
9YzulZRJKjPSHR+Mx/H3mukq9k5VTeMqhWvwQmMXJz7uGZJZx4ildClMIi/8HAgg1iJDyAY2tt8I
0xXEqkI2OTop96lgwJnXgQEXihRcQ3X1e7Rt1dgNjqC2mperNfeMj/zPN0+PeZvoZcP4RAZksBOL
zk3ksasK+lI9aeGjvpFSTJOguIFU3dfeWx6N2597h3fFuKs1//rlxukxp1r32HjJwl5Mq+z/mMt1
D4PVt4OwMYrqqfhIRe+RBz9DL4JUX325F2X+RqeqQX0jeFIn0UEnONmbJDoQp3RgxRe4ywsV8Jlb
T5mhFAhM2NHT3LBxfTWAxmYCtPkIQD6RnIypeWTZEno6dMugtTOMzzqXMdhm1yu8PIf8Kuy30Ls8
h3P2OV9dnQ6UubeIfmj31ccBg2V+7Gld94xkQv8CNsmSKkOLrmSc76XfSxwIzyLTNZ8VKPSjRtPX
CXCuvEjl2EIF16qrvPCrdrzI9bKB6i28shcA5HdzlQskA18kc4SFqnbbyV9AbaQLA+bRHHA8+mz3
RhjH71nxntganUv3qeCHxUMg7l3Q0njp9NHm2y1NX2UPQ1CR2ZWoyTcJcKewWNdXDmbNfzyVM9UI
OC61GhOFZiGSJc6tgn0TQlYKHM10ezKktSPBNqt9B1wpdPjvq4aWeVb6IBw4+oQ0OXeclY8xJWIU
gmtOb81WSZdUpD7h0ic8ZSuIdjcG+Dfo6VfGwFpVi543zDR1idM1gmxv9zDwm2MOxmUiOYigHxKG
EwGG6ut3opp+I9Gpg5DdXd/Ckhon6j9tyLP00LABUdfqE5zgxsO3Qw+2f7UE/BLAHKs9SYWAKt3+
12ax95U8Suud6SFT5zCV5Cmy5i5OWvuvPy978cHFTWH4MEYVOfd2XmLjyq2akBNFXyTP/lTIz6jm
BSP/5IprK7IE0fZcXp+B/89EpW2Tbvr19v7SWvgPo/vS6Qb283EQmQrmzPCM3nwQ41MS/ZGxToD+
lVclsvo+IxqXxWcJRo2s3NixfMkDkUwrWvBHTVR9uwWbrhZCX+18fV+HGjCNxze+3eo8JcmkvovE
yzggcXw5MVZekE7o3x416qD1Kv/9lQ3ucphVM3iI7WiEvw6LTY9WbgPOERoWP0sYXoPquRw2mUES
yHbh1qTtCZajygCYCfe95PQ8srhCyWeTnTn66VaOkbRDGL1LakOwB4Q7vv8kAOhTr3FzMugjjep4
IewYNvLhIVBiKvPSvORZoRxJ72f+YVTP0mapM5ZYd/B5Ot4L96knPMJh3qlDIO2eDhR4JjCQYVAI
u61JXUHqLP3zqivGhvsEcl3Fle6UHwYWk+nDks+ZBGt84te0GYEd8Sbx7cKnGug+nG0Xs/BRaiQi
7wit/9z5D7vKYjfRQAOTlJKSyvF/ITkeL1BMK6l7EmEynHo36Gc0LkDnhd0QAYrswMqoQTttuw/m
DYFpPNGMG+E2FQizaunkjdbOu7Kos2x62K64Gr81iGu+2p+MZv5VdQZ4rxAa8UGVVWL7a377Fn74
dM+Ue/K5vmOqdGLGWDgIfxZ7HFNPpVlNFUJRO2QSIxRd9Tri7M9OLBDKHhdLvr11xkr+AvyftB2G
a9yzP038x9mL0N4vgyzM0ldt7LaO2HsHTXZYCfqQZl9vi3EGAY50Wxr+7FJ9QOQ8han/jrHaQC4B
SEv2po/+/zCpdENCWxLiJ9scm9gDUqA20ure8kChRzDwd4QSxvcR8JBP/d0oH0nhliZy34VYnc8w
BXMzkHNe2A46Ss1Au9SYtKP45JhF/0tk1d0xTW3sL7/THM16v4rsRtwOGL06qW/XDEN/V1rYkq++
oNSMci0RHCxQlG/tx50uyuekumbjvwu2qbZxdpsm9ryl9P8EzEXo0mRWy/9sb5nsK0T6H0DfVU7I
wedluBeifY0D8goBJ/SsheLYBbZA6hQTKSyz6x0DiVgQzDJYxxofeTnmTw/f8VMNUsAVWMUCW/9J
zO8voKOVOMPXMq69eqSnn7vupNfMBtPyzkr7OB6QuRAMrAbyN8FfOP8V7zCCmbHIAGlN0Ay9Mbl4
wM3D78LjmYsYqkpHwpvUnQY1S+iMU5OKB1Xp99sxmdfFHa7nKlEluXDrJHVFgI1wYQ85QL3iasun
EF8eoXJMJKolNc9txxHTJdhpzCEr0LSwJf5uRoPrIxMEQKZsXaqCgHJNIUuDCIpCUKn4f0+Aw7Wh
wRtiuMpNl0d83NW0BuaKOLWy/er7CYi2X942uSap5WPqeQjrBHscme70oOKc+soHXOWN/c/T0yVM
V1AoGlCF+Kh8Ym9pW4RYU10JzGNE512xYAgkHHrp8lCAFkl/Dq5RlB5tC1bdRn0r/JlTfmnAh9m4
MGv+6QyptRmjUZqGLD7oVVdEkI764l7aw1+HiU4TfUO3fAK7bzd/4cwbTjVQ76rrXsTE+Y5r4LD1
cBNElnVVnpGw84BJOTNAunBPnt2Ljt3BWb6jiecgnmVqjPcKkQIBN53nGOWABasuqD8lit01sr27
KcA/fmzf6G1djDICwVgCWgsbGQfHsRWbLm9+7VWv1+CW7yIoe0x6PaF0NOcM50ZwUPZZXnzTPJqs
LmYPWoJ17pFt/mIYCTZt1lFzvZNjy5XPqgbtU3Ib6zxiWWRUlO1YmZVs3zNf6A9BSucly4lccPYT
gzRKOxz9v4V8tgtqO8vZXj/w9GXsQ5ECrSUXbw6/EWQ4T4P9b/+J8RoNLlwAsePS5OlRESTa1qMQ
3OfF8Y0j7BLARA0F3tZL5CMFMMqOKgXxWS8yTeCQZpl1zXSaX2cDuVN461bdObEBkIyFT76U9ebX
my2L8FnSzzU21hi1iLA7bncTc8fcX1/07hNPiUMAFvvDmD2pVtNHLzEFaeQHVKti+EoJRY3QVPoy
PMrV6crETYJ+y70zwoFj41JE6tFwF9Uad0Tc3GLfCfjq0y9hprzSQyp+KH6F1jaFIQddDzw8c+zd
8VgNHqLmUDj7DfEJ1jfdmxyiC9Up6QCfaPzc3go1JPWyVSPz+QORbF7xfPcsbAG/KaProgVaefmr
ZJH+/VHlRCqqyZSeeUWHuiEBOsdSUl50sDTGrfZLbUsHhlNqZ0a2wBow5sOxWzkd0l1Sgq/NCTFS
U7USfGoCZV/TATPPmMxy848m2vu4GwnuXe10vu1bzDplM4l1cuG8SLbC5Bn/oUTopUWwsbGDvSK+
4JjSTnvxT5CSxcWws0Ye3lOAfZPFPXFJ90uY7zVYimpP1wudeJ+XXxA7gfhQFh+dpolLH6BTCrZQ
0EqrGIN8pDsWVPlsRWxADww3e6RRPJ9M9aZuQu+Lv+nGF3S0U9fNSeVGwq8DuA3bNhMMFjAoflaF
+o2OHU7Q7ZUJXhhWAT1Ln9t1ShpucCs9FGiRHh6Q33wVR5Ffv3OhxT21Y/MvIXsl2MiVpg9gHyP3
HSmGxQxva4s/prJZr1YK9P3U0OSHIhh8Ne0T+N1goSH+2+7oA5ROTsE+sSf/bYeVvXxvLpbI/0Oo
rEyDSKoShUxbNj/XVfxZu7j1VoWXPHXhxHBR7hUvIhdAdz6nQzoAmVeEBJ68hcmdOko2QP5J44n+
ufrV6oSzbyFs90F+9FzrF9sQ/k5MytruFJOoB+jwCq3UE9Czxi4gVxl3x3md4gmWfRicxDVRS5fd
dsfP5QmR1dcZMTxr9O1lZmW327lFD397gxqyO2HutWQGWiV+XIR23gNEf23QixFXWwn/o2QhMIpC
aQ8IjLUqAxMcQ/5LRj5vejeqonNi74v3DbLpfbFJHbu/IEUPgSczqfDiUngyzgDguFy/Dd9UoMvG
4IEdyz+QDeJjlbs5MiMxyVe3Mo0syHt2srptEepepN1rzARWbfvpTg2AC8PzJn4Tybv2LKDF/5ga
I5jJkNgwMq+TzLhPaXFBw3SZtZVJTKaC6zRRxvZj5rNkNCqIZt+Ev/GckRgty/N9CgFbr4+5/1nI
e/OHXcqdQOtGUF3OvKfP9M8Ah+5f/baXDh34xkSKBQpGySatTD54l8m5dw9bXarwrWuJ2P+n15HQ
E2EciscE143maytWtDrkP1JlRbEtUpwWzHKuGTrR9YtvUKdmofqRMp9qS0svhcXv1udCECf8Cq/e
XxvTexzXYBu5yZtY3B7ixp/sH94+kOcM3Xlru4O8jLm5MPX1xEQQ6FBvbFwIa6i+kyjoi5O3p4nH
G86xNSHrr3ORXEXF+qUco6NY6jm6RKRjvt0i5beDtjWZWnIiurAfgjhQH4Jz2NChIeuUigp2NY0E
rNQZq349Zg5tFmXBfw/GhTd6g7thrTNGFDKde/8dN/p47FEvAkc2G+rLhm7rqyeViti3fZnS5LaU
DkS/+mBNyNPfGGUwLU58r/SQ4oPmtLadMmkfICT5nfIj66Mpe0hMgfS3OW9CrYtpKf5YqSOZKRnu
RrDt3r8PWvSJjMtRsdRAUFPjuSvlhYepMFW9VNtQS/PCEPj8wY5v3wF7NJEPE/ckbzbyZkg5a1MA
HUDvTgUp1id9ixCcf+cpmCXsKpoo4cSYr4dWfIFrQmS8KJCShnTdzhRKmcHz3MXHjVRKOUtpuLH8
/04Vy+Plq5WGkZzrjP2zqslkHtpXYqtKWF+6aHrypoM7JEZvvFapvwOjk0S7Er3868CpZLxDupqL
Cie3GJp613R/l26RMgn3CFbH/vupE/QfNcYmY3NrJAYaXvTIhmNTcYdnQSSjN6N3HxWlTmvuZOyE
Hisfb43tHV3N1goBpcn12YDrJTj20Z/jxhhv5K556o7GjF4ySkls4CYZCQZTeIojtsd0maAZGDfP
ctrjvgxyG/Jn4lzCn6zP5DtSCU7556xKNOsAo940mL2Sq/34fgsoII5HvPuVBS7OZHkewJX2oquT
fV375qIQtoxXJSJ2WUFsnZYOnELpz1IX8fQsYmYeAtx+2oEDtmubgrR/W4ZnPzvldljYXtmMdSvM
fgO/UWEBB/JhEd7HC+SHIQaAM2rWefoRSJZtKpFmnsbIEyU2XUI3/nyT6KFnbeOogRnUq5FEBnAz
rEIpDDJp6W1AuPzksqbYueAE85TwkyYFtOw7k9YEgyX3DTgTGYs+420P7T+bc65nLd+K3dEaGEgo
UDDM0+2pCE8oaJAh3MbMIwf6vTjBJVgpQ1yvQlpT2Zbpvc2Tp58EdiTMaTwXP9yI99OeWU3r7bmw
EHwpI+SR7OX+OamUutfB2dX0z6hfxzeOpiP8VHrn1ZtLJKIylp6YxiWvzfm+Ks2uKeN7cfGqvpHX
1ApHtzIoUBsmW+fskAttW2eB+RnPcWV9LaOAgjIZVAUObaKGnO3wbtoC1rSBQ5F4oINx0LbX3xqg
WvNhfdAjVy7QoL84lF+bDt2wVYrZJklEXYlrArwYF4bybpBLApKTHdTgQ/UOn4b68hZU34EYpgcJ
Y2pljh310jdUNfNrvRTf8heHpoSwOGOHDK7zqfXqZMpMmx8/JjObcVjoit6H0Sq6eaOTjbJ0mmiR
5Mk4DJXi+n97ox8hxJ3Bhg3M0j2JFT0wfTlKpgwGrjdJkMdJtT4R9VONBGLnGDvNwnyI+qpy4y6z
c3YwvQX90Lx7yQAZre0zZiFzwjiMAYt4suhbtbt813u/V8QS1+YXJrsEhvKEbQMne6TvNqnqJU46
lDg2pB0UOX6DMEHjkxieav+4SbG5lrwI2T1zXk3pnj+bkMkoMCy9JJybDJa8gCc6HiMokvX6ro9/
DFmqeeb2xUcjVQ6TRvPVY3ok1MiCh4AqB2x/NK7Rqqfh87YjBtrEEO8b6EvwA3n8cJZ45ftRExOI
mUd3Bc0/SudyoFs+MeI/6ikhI3IAEuCTjqDyVkPK+/PERUycXMXGvboyDhwVXW1jj5q6UPnZP3wl
F2zna+ujbAFsx+NQdnn5e3uzc2Eqb78NsnjBkFzMWKifMFIcbyuNmGC4DbRxWQ4bfcMgnDSmBk+a
/PcXIlorNXcgcLeGEA3OrNxXYzpw/cN1qQRlxdqPyUmxj5BK3s9W6pIfBIElIuHn7PK5D1QM6crr
IWGQMnUTmRsVneOT2BgBvkF98R+OkWk7oEETJy46FARxu8r3baeEp5/Ld5ZhmiozO7K9dSexAvtV
XyZtV+ieDrLbj9RGUM7aKtG4Q9uMfPNzW7xKvvQgilpNR+hVTYe+bpoRUCK/2Q5Cur6YoLHtYvqc
MRSYI53XYATeJsAo0Cz0cEwBABSAST7ME3+K/wVBM7c3NV+aeJ5PINYUw9eGNpLbZiwDFTEVqzqu
H/kxK5sqBYfKUPT9n8gl0rnekB4nLfvCXU5NSfp1W2h3iqZfooDXla1Ev/e9HMqg/X0dajg0bBaS
IjX47CMHm5luHyE0gTVvKmH+E6lMRCquR2gsUbUcbLQxGWe/HL0SpIzXuSiPMOkF5ePfRUxqkdLY
jfUuxe6vcy+9aDlPQDLY5dhSmY1o1vEZvosrWuwaNvLkmu8VjG+Esd2uJ3EHO5VCHwtZ2sjkEumw
ndO19ewm1ufDdjumHNSLT5eUooaJNz0+V98zMMxV3KQeLH4ozGHH78ZBeTvGVqGwYeav5XxSVUh3
OrlIazVZ2IRvtCIFwvACxTkX4q03sj8V814mBtL7p2RtouenMqmvCOxpUA658WFMF2dwZWNb5u9t
SFzE4CgYZqGVXXqZ9P+3nqyi/XBgXgqsqUCO/cKwofJ2MlUc6jkl3PjnhuCmLtZIyO34tPXisQ5f
aJooeQdMIuYVJaqoBCYfWfZS2Hh4pagycyoI845mF+iPiBnLG6BtteKwvOQ9mi0zXbtH2KUlfegp
EZbyxwYEALSUVshjUxjmBKRQmRx4DIN+EsKRUFthIi2l5oP7ByJUbcr8E/k5EKz/GKTsE2nFzjzQ
jJ946yiNl21tbUYAUse0dBl2PfWmupMoAsDACaDaeNnYL3Mb/HAW2AUTOinvrQ8HrvzIrN9Mc5kk
fkESSXgICUm9+Pkqyse+zVjl5DKBC7dBgJBoD43dt1w9R0MNR3CtF68XqSESfXf9vYOYwTQyfwIf
EsLT7nPAFKyzd/XOEsAvsFwYjSykZEviM1WVGeyp09Yxax0pXIx6H7MRAs5cNXL5RoJat35JaVj3
RcUSiPK0/f6vcd1T/6ZrIOsSNadpt64pJy+klysw54TjM9jd4MYxOC62KNk7+7HIeZ6gZJ0GyCkt
jt9Sy3p0KBNkkgGJlz0ZSX8vgu8Bra6U6JaNUNXSCLK4O2Ea2XHfi2hs8RujQ5D+8yzu1oUpb36M
uRC5NiSFVn0GoH9jXoMWqjFPnQd4b26jvdtWiZQsjzwh31Xkp/E/cW3OgZUqkwrMofGOrChr7S3f
bQHdOC9qpy/M8hbbgkYT+mncTQvvUAiY35yFoXbacQqzl8k77QAaxJXe5oPxUCzsxNJwAsD1ZLEC
uwufiig44xq+ebC0q/N1gcojVurAmcdB17M6ApOSOxiw5L+o4S3PqXFhapDrNCt8o8ZJhxZkvpSv
HlikW4G+Szl52PpVLxkvPHQIfdsEvcZ6GGX492wUh6rXhnoyNL6lryQ62JiWtKaZTsV6iFw/s2eI
m97ffiV6YueWO82eX5daUVVTRaG/y5qIF91J0LWCC51QN6LrLMKGHARBUvSAC8k/F1TWE66NgVCT
u3ho/YPfZcS3Jd7ygJGAgG+1t90XX8uUbIvqQoPdgU5GttAmcyzE9hynSkiKN2GfRefECY01rLR8
eo1smyoKKYrHUHEg7czxvtdgJ/727kpys2oY4Vh6nFT1jS98o2A4aFbcyVeE8hjGosqgadS2D07Q
pEaXnJ/w0DsOOrRLJS1DQb/gDAQmaboxi9sA6rvuaQNjnSeuJMnX6cOLppUuJYGVVrPHH2+27UFg
7QaWOByYIqagL8jYX7C+t9GJDgdpi3t1+0A6Uh3YzsCY7iYIzRr6R7wE45EUnIXxyU4iLRbhHueg
SB2Nbvscvqbo1aUsXp+eZ9tYrFjakH3wBVfYt03IlJpCFTXiVmXumLz3Mgp5GPsYtT6J/6rRvqVU
qzAoRLPy6theCQnzuGlVn3tCjnJkXY/EiuO+aP3tKVhPr7U2w9yEEv5gNZYE6kXIdM/BYGGgqSNG
P7q2mQkh33B+ria24oErEanYQPmXIiQnETPRBlwX8K29ChNUlPOsORq9ZbaZjC174AOgG8DcOV8e
RwNy0BHhO0Od9ChFaE3aib8SE5Nm0tlTt2BQFaiNsAO72y/XRTihzbCfrZz+5BMwtTtoy7p3J1u6
1OSwhu9tuu96kXPjxTDr5cFgevOtTus6FNXHTzgkS7yG/iUme/fwz8Hb9YNmOj+uw0hWOhzJueCU
zEvsGn98lEIpQ0kiCq5jWZQbKaMJTnFPmquugME2e0n9Y9R3skOOlXGUl2eHbfRvF4ZJXb8tjpN8
d8owcjB8xGTsEoMVoC/05RYsElAZtliv38f/6LvLGIqpKX4qUCWGN5HgFtEh2X4UgtyKOzRVbdJQ
I23kW6b0LBjCtgsqBr4+OdP69eOBvhiuPZHpWFr+5RbLlWYXKdIRxah5mmU6eGVgPQWayChT9ZSi
ooTAdqggpZwQwclExWezHXN4+T1FC7TgYc0NdznnjNA4gxBaXX6VkzO7wvo82ualEvutAIqKJHBK
cLBkZ7R/a2f/eDU7zBIq/D5pgPf2bC2ZAsdqlVGb3++pO9pKLhV7GElbpswxTZcpBtgdAoHsM7Qh
jmm6ey7Z4iSn4s7mw2ybLxDFbAke9wonBsipDbmIVIm1Pq3Y27t1yXgVUNs0QMoJmCZhL+eiM/dS
vgBac1inNS6zmfBjoVSjgZmYwIh8d42TdIT71JNi6K8sRl0zoHA1UxB/OPO5o/snbvtu34PUzm1t
5ln4Gm2yaoSZKS3ikRC2EBn+E/3XLcNOz1h1AIYLGKmm6k8Fbzbg+g8B3V/tVztT6xdPPlUmNkk1
1s9RcpV7DAU0W38PFgd5HLLZljwLVQ2vNtAafd7umUMk7TMf0OTjCkOAQMtcTLFJHXx+mWlhdvSh
trQR9EMfnGc6guBsZ8NZyFt250HLtNeu7pA1miXxrLnKsuR6ISkir5f7nXtUuwUlTzKtZ4x2DiPK
fDXwAZ6dV8W1D5pg8iNXtR7qtgIHPvJ/kXYdQZsWgepClSqbs8Zyqw8/PAn0lcZLo8UN5Sg0k25z
9wbz6ew/NckGAE+az42AkfziQwjzlv1cBmVKSr4esnzdQNhmP2ltlELTM3ODXY5DGpkawWpNDdsg
UNSADR4sKcwBRD2aA6pk4F11LzBsnkt2sMhNlmJFgnzJmSGYuybsSv/gR2ZmW297j933pLdbb4Pp
k4qJQFDgyiH07X5cf59sLBYU/D0Eu1rj6V8jDEINRuN1Mx14zGAN9fMaXWnPGLcrmDQ7EopGPMCs
JyMsSmhvlQgQOWXD7Ib1nPJXopgsWNcBVa3rJlpoejiM0rS02nVCAxIRWn49IRvFDpWgpE9mLR/C
oAafvWpDOpaHd6nMgw8w1Ena/+wbFQOR2rXJ+Pq8bkyHZwMF1LAIJa/oZH2eyRe55R76f+nWomFU
e3E3K5PtalBEx1SAfPR1HuLVgVsghKZxS+5lsnkSB7uiNWmJ1An4OnV+hx8JVEhQlv2YxT/bV1CY
k7kS7KIy6CMGkDcuzCV1S8xY3z87A8n5pR24Vh/gnrZwCW0LHTMf3EDAVJdzdH43XzZIPCyjKMA4
G18yqI2egFcab0jRzE2AoB3jS4uTbE+XeBDdh4uK5fclDXSLsmML/aE71k92d5xgOZKNetIBa9CG
bQJrwkvMp+YGkdovWFI+J3ZRhSgqci+hQwIOzGz58t5hhdl2LolT1//G/zYi1jIKYXuKfVYkQG49
zbAOxkpRRJ8GfJHmi+gihj2cwFmQWYAdcfxfRItL5vrciXlSunHXbCypWljyY6Bf/2tmPLSU3CSz
+muXr75Kuotc8uiSKleyUgSBXgAjZnVtejAmS1FLZ4lAKymmklk4/vAffh7NdezDEMPMCo5+0vMq
niJvqEdtONxzedw21H7uGDmRo1iui6UzfKOT4ncvWWe0d96uXVkzTs0/qkU4/GqSjGOKb8rx/Csa
ZvTxkJDBf1cC7klGiqPjmAVMT0/XFBeqXa95jHliIWBG7+QuNNq+lm0HkSXqRm13fQUtoGQVBAp/
MkJohdYeiC3mWX0FgCcHSZLPPibt2H9RdgG1MArq1F3Llz8OIs84/0u1SAdpGc5jVUCnTdrdCBmt
ZuFNRTslmrt4dr/qt6GmxGOPsfniK9mFB0AjnJGTK+SMj68KUur0cZ8+aLLHxl81EeBCAk6Ff/GN
tHB5HNOP5PRKUnsRUYU04sUttm4RGV2RXeWjVqOZENX9RgwdFOfp6bbZIYP/0p4AaP7veW7p9F1u
/DBu4h5Dh8fPbFpyfAyAAyTdzAzNNWsPa2Xys/CegIibVbp6JkCAnt1LNhUmW+rjqdVzES/qcAEp
QMXMV4t6ukUNY5aXM8Vuilr3FAAoqeAODPSOAMdKPS73k6u1eQpxcgonmLc6Cdlxy2TMr3ayysDE
3hlYSarhSZcDO+0TWsuoUM/5U2BuqwHGYCY7yZCoCc/RVpjFHBx0TWzszHRHBba0QryloEl6akcx
5JmS3x4e6+/pHwb8XnMPUVN6dB7bvC785PiAyvmQrTjSOih2OWi6Nlk+ErKr3K9yQ+LtTZXW1LNx
ddUcJFBq0ASYNvX1ikl9WrtlfZ+mgMl/KzQvAiJY6MrkVkxoqf6GwOqBvRRqlCa4p6VLsc3GO+gQ
6bjPdfGrOmypTx20swtSNojyBBZ19stIHLGzDYbciACkBDQrPZ31SoyfFs6qH46tsIyQpXvmq4kd
OglWEJo3ja9kiQEOJSQ4HI55GQwyXd9xFok1svaZqkh8YIW9R/9+abbcexUA2QS5s3hbzMwoR0aI
CidFR0S6c61Ni4IHp/LUH1Wndxz8LXOMbUmFKCZyn0umBqh1qmi2Q/IrUGkVZXRGgJLlH6MILNh7
vGgmsdJpqIG7V9GngCDedqh0Wr3j5GupG8iEqpnwmscBFIzeoLXIkxBwSSM4HxMjBD2KVZoHzNN3
TdmnpzfpCES6eeko70DyZeTF4TrhwvN2Fz5axfWEObNm8mdFlZPb7fq/7xHoCHigxq+mDzDlCIR/
xXcCJexGkt9G6/rzPuiv0sgod2omcAxFZF0I8cDaPDuqxD326oGRdPW5iEB0nwqVycsC+X8SD1i4
yvijQnky3vGcT6NlzZ0/FXbC+w2v0wRpWpKrjHECgFyXHgGnBRlNfxhTpk+B4nvBfCC2eT/gFePK
NeLYW8yBHDjlv1VHkRjd2v+ibTOd6JcmxPaT0mKSSdfoHFR8xt87npM04a5UPGI7+oGM2knAQl+P
HlQQBPG4vu62a+rAUBT48YlsGKig/bHlzmhrO7ytQkukmqjlQiAxyKQzq1N87U2QJvJnLhvSeInv
CiXonK9a4+5lidAS/vuLbNaIpL2p9dVDqips2ZpFzpdrj31VYHW6/612/zF5hmKkGaTHu3ffym5K
QZdJkwBGYqrspNt8TVk8RTOMeiEvgE4jCXV+R3tb1WYRrCnrUB1kK+WIGBJHWCTCppK9vpM5VQBt
8qu+AXcttmMaqC3eF4sVuu7rG2p81oIJALf379Zgdii/Cg/2ruJ1jDGwQTK+AMfnoG6VL8mqEG+v
aUmB43hW/ykoOWp8riqNB5dgs3Op0Sd1LYbDU0FJUkuZsupIfhQ+Lv5thM7+B3WZFiVTxKo0HDqO
XYg0D2q5mcgn8pKZuBwQCkelhAzO+GI3QjkMMUdrSTlee09kigMLyfc6+563I7FmUwMXpXEXRFV+
FKFmO7WNlJeHgETXFtfZ4XO77DORmENyzlHYTLmeMZIqgWyv+qmMUoJhTBVL0jpx+7xCUS+xVArV
oMzF5UQ4GdZewpSVjWfxT1XMiiJEV2BSmTBGMbSAOjhTPuO29uzfQDtuL7YE5kx6bwzCSX3lvNde
1Y4saB+JmLHWtTPoROAHaxBk1dkvHGzT5uAOafvG0oklN7n1wQhjl24jnk5dXqUdvNeEAYp6i2m5
Glw0MMU9SoaEJZkbGjI/u6Jd0TmblbMqgJpQTeKXtbcOrBatVjh3TXFTk2wcaD2oo2LNKiJEsSKL
yyy17qtsn2E4u4zQdxo16drHCCh6ouSE/z5pxpiUogPAWrpazU/CMwo8cSIWVmxtnf01ZpgNvy+1
xdHTA3ADla6LL8p+aWIU3AP22U2QmetxP0SKpo7oTB/2AuRc9neQo0Yo2sZ5I1jlENvE4gdszHF4
icGiY6gAXjjafHSJUekDX5tGbmuNXyshJ+IWUfv4afuNKMPVTseY4t30Au8Q4M0eUCeuLqXp7ggI
u5MeD+ZEbpp88LJs+60cgHk5cwG2lNxMcBTOk5mc0B17w2nxSatAU6oWbNZYzOV1D/011+ynZt9A
Gz37sfgIrCg2zELN+hahb/+R/XnpMRO+EuN2DnVdfm52Fj/8GXaTmNbAMOiddZtNupqHnlhbCpAx
PXHTwK+mY6yJZoAhgXi1KyYg+mqAC/LNV7EjtObPpiQjm0u9qFxTuL9QPNY/Cgd4H44k/d+3KDLY
MeuXuOkE+EbIMNEzYZCKIRG1lQC6kQ4oPtST1o1AULsu3vUA6L3kzILM2D1xAlwlLMqFfHRbE8nT
akLkK5uGG6dI2wLAcON/Pv/x8R2iGFDxG29yJTqKoKjU42qXfsQDL55ZnmaBecF4PrtydGkxo2gN
7jWuqJEUjLKiqJjgQOA3vB641y+exZrrugxgHWwHiPL/ukjRPeAxNTpswjCSM63JBvPjUbcu680/
KdapBRi4gTg7QWmCS4HM766Q4Ka04DUJanwMjcY+9Yg/40qOqDtWBl4YWVWgoG+3nU9UlFcQjIcO
wpPbCqEJTAaqB19nTc73XW5l73WffBien6eqWTlTDeG9h/BemkdbMEgouatVSdu4L+dQPexlUMyr
tkd8L9Ja3eepqrxJi8+rN5f7czfXR1JBLLru7Sepdh7PUKi6H/Jk4eq1XC7a2G3qGn/GqwXzFyU3
voxXO+CAi96YO+IYt/GBglOOybX33DUpClpWJjyzTgTsQ4aiciZaApxFdZE+xCr8QXIO2t7FAz9X
0ox/KJ4IENO/W89Y2VtsU6Q64crDmx7SSguPX3h0nV51oV66iXJIvTTe1w9uPxJRjBfWLGIDbAx/
MRFQxSOS/2BS6R3gCmBbh86hkQ61d+uS9rbYAXAGPD9J69fS1EuIyNog++cJOsHapoDct2Uhtovh
k3oaP4HefYfLAwWq0tM7Kpwvm/8a3SGQKLqPj14mdGbqlHloS0uXfUuvE63iBJDDCxQoLpbQRM1T
bKfCXHJ6rv6/Mkh0esI+S3uHjfvKeGIJy1ThhYEurX1nnmK+DPpwGh5ZwqqWqr/QRCVMt2Z3iBXD
2p04BlfW6gD3pmluFOmGZUresQtfufD7qYyXsJIbckq7KM1VPChHAES//U4/wopAVjRd+pNdVXMK
Nt/2bJGWF+xwn7xJxuyP+9wBxXSGgKU+KnRDjdZpdv/9K831tWxA0YtBSBdo1ahU4xvnrDaMKAf7
JgiBZgCqPM52E2a+nrDSduOzt7gENjv5etfZpYP3ElA1LmJquUZU2obvFH/KyPJB73xwsY4dv3N1
i0zQmy/d8PjuAAYBdoP93D6QszAZUgEPWyaRuPe11jWCXZ6Aw3sqXqsrIZoViDZySslG34dGpWp3
g5MMzu+YQ441Qnd4VDCN+gwSzlBRy4x7AEPmTkHSceXZCeoxXOsya+Q8kCMvf8fjMGi5Fck0lGQi
rtFOaOfe3xS2FxhVY3inYVpYOQgZYN7KWvmkF2i3bQxvkgpGxjvbo/lNo6vc6z3CBafub84QFNpo
V5z7yuPlkAtmKSmgghU6YxYOcqeGDPO5KIaBYCUvT6W7oDP0b43ymER1ptUahOvVqJvrIgrG50at
sQLxPweS6fY8blUfypcCkla3ERFZm4jKDgVVC6p1x3+3rxdOBgte7XsSuMxhB7cTuqaXIaA8gpNU
Pc4eO6Apf0ToJMspWNW3cw73Dj6P9fR52FRPRNWqzkaWZKAwnjuxISGAzT4CiffDy6qGUcv1FuM/
N7R+i/sgCWhwAiHn/pkmya1yaMhhfgeK1fsmmE8efmiaWRPXXeblibr29ytm/KgQeWT1kTLDS5Hz
9TEOhn3LM0dF0eXxNepNK5oDLCt32uQiXEf9yvqajaJ7RzmV8LU4aF0aFbbo14kkyW4XlrBGbpk4
onSbHGThVd9ATl91LFRWsCRjNCdKMWYHVGN2qm4JQkzB2EUaUVZ6jjwq5Bxpe3ZGLmxh8HguIDp1
uMvqfywHPT25xGhSd1QWhnjTojkXLIrRfhYEs969NTSa9X2bZgikGytGi0Q0f34NNw6qB4UP6fQL
5HHAMSJJBUdUETwHCxgkO25j+ReNbGnZOsrUNiqXQmBvDvGSP9sTkmRpIrx5FASATPeTPldtVzRd
UUTlOeUyotOvmD99S4GBIEVpKIDW0Y8SfWwHjXLImsZeKoQLG1qVXr+EdrenvYqQtQkcDClz7V4c
yp2/rnFiBfFOWqdCiMDYQ9pd3p4s5W2BNHGZrx8CV4F5m+dTfrHd8NxEO8/JMRaPwVoPTjZ32wIF
qCOaUDbPxVSXpzxR10+bC3mIvfgumTIp8X/w2t7oNq8wSz/dhlc1HiadYs17jPRSMJWhs7dxV18t
K+2bATLNbVsikg6hMdvzvLLojUMS2la19wl02yluE60kiswuQdnEFuEg66tRBrG9GeRkCyPsMj6d
RgAdh11s/ussrUeWBn4gB7RuN1ezjAv++jMsubqIs7wp4LHqGEjy7+cvZp6HGEUj2fskfuQwD+Ll
HsgTdxpX5J4gGdTkDX5RLO424NQueY5N+WZW9MoDkKpZoEFiyJVJYw275zJuUNwJPT7qrRbnSNCU
t6/PA2m4x9J2yEshxzg82WrsWJGmA8RPVOvwu3t19K6ui9krpy7pSIgtFxjN0VW236rtYg6SYmwD
qfLCo0A3MDXDYogUtyaR+z1Jn0xw5Ejr0cjAWRS5JPY2lUAimNYTPJw09P7sCz1k5Bj3YZKacyEC
WvmXFOsOXsPkKqELo6mQGToMk+x3W9gKsDA5Dfnwuee4ppNAGUFxouqLGMLzdd+Ix/Sjy0/n7N3u
7KDqQF7D4aU2JH95XMRXU8mib47yUR6JYtVzYjXnldcR4K8lf0VTfYbYFV+Hriz4YbNsYtc/TCe8
HAmJ/vzmG+686YZa4X/rBBzMb+KAW1jg2weT8LBfhg03tVyncJznLU3IC1ES4tGTmT28e1lBGvW8
RAFbTwXrcwfzJPHBdQCJmWawNwqhQp5thHoMF+V7EP5CrJgtyJKwd34uS8wgLWkPvzuStBC7ykXd
Iwr3D6RKrLEi1qKVCsaLUyV5O3QyxJp+N6PQVXZLi56wh2pVLOYD3VVB9xOb2Fn8YzoHP1nlXCDr
OrVN5+O+3PCsxKYuRpeMfhybPoHe44NRMWvUEWp0Nw0wQGnLiwZDmT9e54nYdor1arL11dtRFF4i
qxzgWQNOA2FAwcO7q3mEZfgpqtupo1wY7eTlQLFzACjboBR/CfnLekm8JzPnhEkQwlcRr4o4O7g/
2T7Y3xJtCraZHl8eUmmu3pl1pyj/7W888yT/igm8iHdtVNoWd7EkW5R9ozJzrXI5WC7PW+pdir8z
oZtxnhxUcwnkgqoL7iyjF+MhK4jy/tBN0MBV6rZ5CI9Xu2XIZ49yzuLFRBJZEC6pG+a7E5pTK+6V
Pzzd8vUpQHNxUU4P1YgNEIGq5YN6F7pJsLKPReD1ysbRHsGM8RHQQF6EZiBrCnuYcwZUinEmb3O8
YIfytTBfOt7aLYUFmoEX5HY3Lvtxw7h8hp4dhGnPN1xImB2BOx8a3IiGHXqJo3vT/k5zZiwD9glO
EzyQS3ldNGbc4LtulqMz40rc3VnhS6E9M490igm2xbp2LmLXad4Rc8LNxEOLjaPL6OQ4t3m75tjJ
+T9AZfXpCux4+Z2e+VK0G1FY7JkaehpfMLJWjecALoC51GUJ/xgzh88JBuKlWYwqFRB1dlNc7Yp7
JHv2LFLSm8uS7VNdw9wOxqpmABUAhOtH9ygb/BIXIdYLzMck6dY/F9YmdS35NYeYCE/AC7fjkK7c
bHalzep05cmQ85lIuuOVYed9fC2ezJX9PiTY4W3aTNmCH8DGMWUzDbIw9QNmUw3+2QEqSTCxLSII
Wg2TLXt1MNnEO12pouAcSjJCok0GqyeKDiE6ydo3y78B5MB6ZXA0j32lea0YMaI1NfUCKR0hBXDe
xVHgxmZQatxG+qAtVOSbKbX3UPNDaOG5MUbJNOijaazmLVwzrwg39sSK8gHj2dQRquztjqbP8egc
2HVmAnlmGU1N3kgwBqi1K3C/6+Q98zyDYyaSoMnqOsXAZwYFu3bWxa2EYOHWe/xF+2giVUhH2LeP
2x4jl5qe/eGfuHrW7jA7o7r4InSw8Vwnc1lb8eoyazLAAdof87Yd+xG21c+nXjvguX0dMkhYNHxp
yquRdy0lGaAdv92dWHbhZJpHeSamf2wI/xhcvqr9DBOUhKTVwopx/4mtT2mG2Gr6xV0mm3ycjUXL
hX2PZ5/Fx5ktP/OzxNmPdSeO9vJl9Jc6NReF5VdC7E6fFL39nm+rttSoqC+U2hpGK4LygilVG/sl
F91TjdVvrq7cEuUI16FjueXEYO7jdLb4RuRx8G7EpRloCHb+3v80o8cQ5m4dSnpoZvGd0YU1lLzD
YboxyYgpZaDgwRkMvoDaEZZSWyvf68AaAcY0KmS6SRh2z6DvYwl6cESKEaRh6+UcDDANl1jb9fT0
fG7tFauuWPm0SEZMqTXvfmh17LHlupUF8VGzMMK1g78VLZkXhRXLwwxwbJZ97BxqpzILUcvsfeA/
Hhxz7yQLfLM7V6wGFHhtUt85mdC76CqFBPaPttx4klwg8C40WYu3jc8vanbq53VrglQSZNAvJXOO
LiXDBcvcB60LZB+3IFeLPPhXvogLHu0jnP2T/71E+64vbCO2RRv1N051D+ncF2OXW95TyhsBMkui
SEjE1s3KaeJuY97LSxhd+4CYQrhMXqDtnSJAsZaiNXNc1ErZIIcuOvTAWBoOvQebn3Br6x12gIFr
UnwR/7lnisDhD1ySF2oPIZmbxPpTqgPNl/xUTLsqCfHoZwJq7w65JOVSBuN0VAGyg87g5xVDVQZ9
cx3KYJySW9mraksbWKBvgMjvCg64fC4meCrSgafcKxfmXVxGNuUaYN7egZh1IVSJMYDrT1eRPVpb
b8oF8wX5SEZE6XqSGsZASsZt/8gamnZG9X7EUKVn7Fpnt1b+afBRX/hRGWGRMF3xpitfqkedD/OR
gLQZg73Oa/Rfu8UDpyUF1pqZ0l5Sl47EpMkyuCamZSA79epvVVJSvATEwPiVLsUIaWDZmyKgIkRv
8QdOvCNZxctsd6V3e+SsjGVx5o0NMSzvx3SfQetDmQn4ab4mvkpb8xJJRXTqyuA7nWjP4erDHLfO
3s4GqMrxta9CShGHx+Hu89/Lv2lHAYcSDDeujg5SuMltn2EoKZ7RdOqdm3EyTc8f5Q6T9lgXbLvW
ansooDvXtc+ro2qJWMDIWzZfNYIxb/nE8IKhojJpwCFPOQv64doBQMUN2n0ygnzAy34nLid4PZYY
5flqYqGqH1KCs7LpwygFseXLKHbwMPZ5YWXqtPfF292tQkOXtZURxkpngjtC8H+Fn+0TeATb5uWd
0Lgyxu9wOFFI6WM1tKlfmJCOvH2UhqE5pDqmSZ1zyt2tSWXZbGIZJAsSF47jYOkB0AJM4GMh0x2O
MPKFjuiabvV+WzpKQa66TrJ5CUoklxK4KjOTtD5Hk3chM0ipQoc9M6yb5LR3sfXS5Nbp5JxqcOE3
3PCa9iRhE+ktR7gaM/SVm4oyPGdfxRJI8HOB5rHJKpvOQrxwBLX4s+dSAdUs8ssJ3+h6rxjm55Y0
Ly4+lC6WrHQcCvZcI8G+IALH+B7VyNox7G6FlUMxMUlphuYirLhmUHQTgJ4crge8u+6o3u54J1Jx
K2BHBwo/FC/ldGX40xtmFZxE5aZhkAJk6hpurlnU8MWumu7u+VUu/sv/QBEIDWb1tvHbqQYXP1RO
Log0IuQRBvR5JYbBgNBuVyOUADT+jcvOFk5L5cUvW25KXEUsdoEVLvHURMWOy0XeJBA1OntqbQkJ
Hm0vA1Qd+3xdu4ahLEG0NlvGIO0CSGbMhB2w/FbPR/zf9EBVM8UnUDGKlusvtzwdiQJ3ctles+Xg
+NtIypv/6FAXFJkXXMVIQ7yCFpnxTOxZ/ZUVkA9oqNCFJkX2y8KAknQhSjWtGL2XKwkfOkzNltFY
xWeu4UHd9FbNnO02g/BpC3XD/zI+DDCSXh1SriBPE6HBGaYoTP6QC4eYJmx2VdJgfS+57sdArQvj
gvkiXnIcOuqP97TYEKnv6Bc5FHFb2kTU8FdH6h8up4wdowYRbTX6VIcrWbMwNrF9tk1SEBM9jUzn
vcsDUvfA3xCaK2KIsCJVVgFp5JAynVqq8W9wun8refYKJ1MEDmUuFwhAHt6VoX0pYcilMDrzFzd2
mfjUZ8ZpPE/bBHVmOWTope3IdA0i6HXzY79U8/H+wOYkTGgTP9YoxMjjhobKsKZYU3HmLAlS2obz
kPUkR//+0HPZApzngdngbhOB1xtxJZRfQ25XA+20gi+YEvx+5l4GUbQwJBeHBi5h/eGKil8i1T7B
ydSOYiKxJsufoWouMGSNp+tEAVImW8Zg9QvAIGEQxXUzJfXWooWncC4r6ySVlnYzp3eba2+31XAn
9iFx9gEOauLyF3LTwkOVed/UHLqE1X4caH2dSn4UOFtnIIeNjK8jcotWIrjvzSQ385oFtJX18rTv
RczlwaVBJLBXXLsKvxC1lF3WjOwd1LG43znZaztE59Av2zVJ7cFZbJS7QydngnSDdQKePToebJZP
lHwITCTtbcTwlAu1uZ6GohSzXfXm7rM/YghMmSPHfPRKy60ht+vuB5p9/rdmyqjARnzqrgjmeO3e
AJp42IHMq0DMk6Jej6BMevLbbY9PCb6NVQ4GgFyL3C+cSCMta5tnVSAO3BiYANPfSAMdzyybYwmv
bMA3D9pjIqw11VZMVxwGaM+dGRmhOlQVRYOtE701GCbEN+z2ogaGLrdMe/A7LtTuxqD+JYELRA0b
wrer8ePXb5OL8TeJspttDFlIPjxhHk0BO4Lhs1/3b+IC85VnnIrUfWlTsE5jPGc605d7qnzI1omk
Jh0PD0Nsiy2YHKk8A4pGKU6D27G3bZhXTmJO5l5wf7x3iktPIrWKGMFdASfka//tlU3HOTr7KFDa
VU1bIQXVuZE7pAX5zR55m3uhagRdRQ4en4xu5bujP1FIM1HLfQMzJi9UaxEhB9jmAU8F6qtCkAnn
c3RtejT/ECjGhbx8nUgNVSwwrb0y1Shfy+cijEyAhQTymhlh/YhObwwAVHZ7xLFkJfZc8KAm4alv
PPsCkOMdTSttl4xpljG0qpNEQ8ZnNOmUWJ4YZOXFDJ4h6m/MxvZDo6mv9DJKT1q1xXWw0u8L9qoT
75KTwtmiJRIFPA249+wf0+4ApHXmgZSZ9vNDqEnbUCYRt8CZMQmswcb8ollAf1hxatjigVrPw2CE
9O8MetF45DHDy+GkVuMglEgVqp2p9jFVJRZ3ypnlaeSBZzHF6PFekvRVdY+DEKG8gZTZ3blRsb72
OocEhR1Y+ZoHiMZ7SJPGJhNcBrMuoN+SRqRtkfLt1mCBRXKDEQ9sfjsZ04ko2ucaxh8FGQzIXr3G
tzidY7tTb41Xs6VN6Z4GS7V4YetIgFaDR2+Bfzk/VcAMTwZ5Fe7/N/HOz1K+ojDWTGhsI9aojUxw
iRcLsoe3B2Yk4/LF80F4Je/cb0lAGhIePAC87SzmaPreXMeMeM5GhSHi3OI+jVtkH+DF3RAmco4f
ayDNBpHwBjoHAWmZzexMpORlrdNUjZ7lbuIN8fVYdCug1DJ9C57FOOQABoDDCUEN4hyRXhXuFYqR
dMCl2rvw4JbOoUKqLPCzEICpm4HnFpgnQANrU1LP4Nbx90k7KCSlLt7v9cP+ZO1PCyvTE8/gjwSx
NxRibLLS3xPcCX7vQ95G7xq0el/FaV+2Yn+eXj6PVjHqlghWun9BGVoSIy0q6R9m9MN3IcLSC/mb
jLpuwogTFcElgMlQzh13R8AeHoNlQy0kLf2G3XUqdk8MPqRs0UkehwiCBlFwxYhhAbyvrTgCcxyA
s6+r+pZChDFXFbZGQRyOR5T4nqoJgG8BndY8IzciWJSNmUCbugj2LzUxbZUw50OIlB5y9eKFNdGN
T3JNypPIeDW7T2XTUydHt+nt6Uo7UQo5b4vVr85f4Cw8x5/DsCWMpnulk/yciglMgGOTGdpxncdG
8c2Mifdn4LIMoiabvn+VesM3Vlt9Ytg2t3WvINJKSWeFjGBbbsHjxSlxxskg7oKFwtuNlIImNdUp
GDAqyvcvSsEcbizaBcURMlxc7+IzcAvm7uIM16H9bKfME8Ah6aLk6OWxCrE01TFMeDZ/N8DmTatu
r75JzUfkleiofqtjIJp6GSr60NeXv3nsPjVJhyYFEKrSivPWWDYRTx+KiH/QH0cX4wB6W3vaZSEk
KX4DhAQCHOgtqJfaUCfiLf3WH40bZuEZ2Mun+C+v0Bcsl8OloBpPtUhH9n5CB5Zn++3R5gQQMaVm
i/HFBxrxDvK8h/G7fj3JgxlM6uDEPFyhJwt1eQIWWed6EET+I8oEfSb24j2ALOhCj2X8Gl0FC2/U
Lx2wgrAxQvhirb03xCNd3NccZDTghPatMPgpCNZ1lCLP838Gyu6rTb70Fw9ZG8haClodKRFpcSJ0
3sQksaNS2X28a/p+CHGOEKxdZi9U8u8MwhfuiZfpQGDSrwcG9Bw8aU+TX1rKnMAhQ/bDYLnh+e6T
lSD2zRQCz90TODUulZH1Rx9VTDFHjA7Tl6j5bGk7GHm5RwhEA0OT011RTevyPlTOx26qOENBcs8j
HZpqfQD1If1/XJUIt+DBrzfZeBZALMtpNtK09UNBnxziHT2fkY15ml8gjM2QtrUsMdilrVmeHrPO
wMRabCrIfb2KyJvRQvgXuCPe5SkRdcxJeVmY7j7l1rPbbQ1OypEaoSx1E13FqmVflI7kkPzNiSMH
jNdHFBjS030JUErF4TAE4swDRpNpkyx9kJI2evAItXsXDlw+qljVv7A6KZFSPxbNvgzxxm7AjquG
WjFIL0Kv/7KslTjN+9mzP//9kXq668QJY6inqXDOqcoWi+62TMliH0Su9ZMUla9V9fFFqp8oQvgp
UCamaa0+e/h7GHRK5eDlGT849ruUWl7PYVUw5/LStcELQ/B03Y+nBQijDasbpYlGBdsI+zo4/W/h
cygZ4tZkqHayiu9xFaSVDhrGJB+9z9K9ZUIliPcHNbcb4aybjxcixf9In2QrFivWMjWmQKXkSNIP
VgXNzZPE3RH0AISqmEsKmKU1T6qUJQTFBJ1sNnG+pbZOHXugHglpzibIIkHfYyIAWIRqU+2y8xIF
W9nAX2ePMnLD++TeRVBB0jH2xU0W954YAgTFZFllLHubngMS4+jKlmvub78GagC4UnJM27hlcF73
6R2BX3iF760+dkY6AagsD4c1rwC9WcBQ8DN4R7X9lhAI05SpVbhmstH2NCh24wispSa7Cz9XwhA9
8MKN2udWrnZZ/RxKPGTZHzRWFbwv/vTkQ8jSCg7zYqywuzkYLP3L/jvzdumbGIxdAQdjuW+IHzdK
eVJ72WyV1CFHEefbc2734QeAT/evIcy7MFbrJmb4j/qXuQc9s238SDJb5hwbTul7RpglUUsAwv+6
Hd/sB4pPMeOJHl2FerAYiJZ2ZNzVFRQZj5lA7PkIu9l59nKjEoitEUnbFmDMP5L4c4eCgNMY0PiG
olAQZJoHzKJl11NAPU6sPnpcvfHKMlvsWyNbZwkfWz6xChK1pBaH6CI3zEQ7cLzWuVQ52VXIk47y
PCeXHhs5k79+K1F9ZDqhqHyVaEhMBq/Gt72sv/g/OIgofNms74uB00torQ9Rl1l7i+1GevBs2BP9
AdH1w4h5REvOU+2OIQZY7kjTg6JlVytsWt1yM6FvK3KfCjrudUx+JLYlZNAVcYpYMUmpepNT2ikZ
Hqx06GB0voVeYsgrds06GjKdENyh6ax1QliYCS63Dp9GVZUqPHXywQVZh4tj2lFit4jbs7ng97jy
OUMQWyD3UAjm5Fi1dMCQqf6Yu5fqKeAdxuJJUDuTV/7FwA3FJYXK1ZeDlnOK9uSlo0IpuC0Uu/hr
bflrW42JI8XoHndVWfcW6y+AzOdnM71CwW994QkARhMU+qelnpUbGrhYHpaKFOKPiqodZJvH7GAV
Rvgrhd5bxhuLBAT8njCdYNQPVHbmH6RCOOYVyYXFk+cXrUqogxhIUwS7kEZBgDHSb+bqJ/f3oOQj
k/zsfHfPXf3YyBE6AAqqCLdp7sXr42VTi5jX53kkP7xFtJU6QNSgKk43MRE03DIfYH8rsw0nwd60
6px4KbUQzyHkOwdLL7lVAS8wzcvfOqUO5yomOiS2NdMbK38FEYdvZAYRQY+xhY6eHQ5XQytRolk8
iqRzVDTSE67uKdwYCSTldIVye6h07HjwhE9P0Gt4pRD11qa6lcMhhRCl9KYYDsFWv6QrfnLCFZw5
TOHwmAksjbZsebgeYdPRKhY+Dctc5J2CE/xvf40tMI+m65ThkU6jK77AZDMR7bMCiqm3mjiue2DS
3OB//7HEJUO17yQALswuD+l6LpTZBp9bDD6TpWBEdEEAnEOIie/6ZlmQMboRrmyP6wLbLxTYdddJ
4nJU53oH7gCz/Koc60z/vnbg6LFnIDkNayEXlANQbGAxH45NSPjRm95hKpzk0+p1U6rSipc1vxnq
zzlYSAeo42hA9P+ZevtC3BKMoC9tCAey1SAx+v75AAIK0YBJRVdYyBx8j2fkGwxPsF0y9YuR0fz8
ujd6ucmI6dr+5lMuP5qRMnouI4Jxc7ZvJp7NGNPOm3u2OTjedyuH5Rmwa7yqzTSbp7h7MuAm6A5d
+2HJlzA+mAkUOolzQzqDE1KKEYbZp0s7MRS6EI1weoNxPB2z0eJKFhCcNDEGXf+2zenHEhct/RWu
fuRGFG0WHsECWnhvb+V256Kk+bzdal64i3sUx85mt/anT9zg6d2BVOsxN26xcBawuAkbt4uxvi3y
gEtpsE73vTDx8jUyDEKv7EF1q95kuDtx8EERFwFvaKtvxSKKWSsXfhoekK7XJT8pXGc739SlH48u
xjn9rNCzfCoMdaepGqN93vL2BkpNE5bV+qm4fnc2CMh8NawqLe6RC4HwbTOqK24kZtErb2oqVKUQ
I+v5xglAv7l7hTUAuH8IOTOcWzKyLzME9BIIKIkMrp/lGV6RyOGJ0KEflZSYZvqDXb5QcaHBQzd4
6lw+xcR/Fg60TDdJT6+i7RbVNiknlcmhUpVYGmFWCF1oNVeu7e6USGiqZtA5y2+FhuA4RnzA0fej
AqozzDm4w7Ays4W9FhxpUi8LuW3daVXHm/96ryrmueDVvh9FGsJm92sGK8Ki1eXc14O7k+/rEYE/
QGK/DT5SHsw3PQFtmcKIOUjJmq2V7GJfGsw5KtuTHsubSav/SyPXaRoDhOGZ5j+EcIFtMRDOcgye
NyH5yoruFhkgPHgsXbs+KAbIgoyIvbjx9jCd7J4sOCYGD0j3PZ6KmHv/8JCi0Gwaxqzd5SqMLR51
6uhCE+lILaFZJMCag9r/yDXZT3oly3qzfOTundygH7HemE0pM2TEh1qwixpHA2vAeNveiIunKCMy
mPXy185qbNQEHmFjn1Lwh99tDw4noGvCcmPsBpEXFo5F8/STeC8w0zZL/NVHA5IqZJPeGr5sYbUZ
pyzheo/kRoyWy/ZaYpK+ZLSqh3kdHLO08jnTxa/FC9BRxKJvyHHuXBXtEJP6+53Ll7en7G4NkNFE
mJCUci0BAjniNN7F4GFDRWx5fvcyLSfqR9gAQWKw30hkKyDYRyPOcwIa1/VJKAXaNNEtvRgZy4Ny
cpjv3bGgxpUUPFpYvgl2v9Mae0oeBy5DTK1QpUvXqkdI0AM527c006TkxejFJKJ8OEp3Pqh3eNEE
SpIGUXgJ7ztZ4d87E6meA6GHEK5K8csyUGLr+LwmNaEieZmAT/25jqMxgtdzxUeX3DMjIvm+blXq
/DJsWFNGgc1ghbqpXWr5lHFRYgK7XRKWjjav/kfNJbqLezbYb3mgvI5hSe1F2loYGfLbjlkM/8b6
tMWR0DqDcWTgm21UqrwuZwNREtNzn6uclib5Iw2bAOsyoqbdWkY6K9YicoTFmh1ELUBcT2mEHBS5
Lj4Cze2Y9cojMmWrML1seLqD4k7zsULS8r70aYhE1XYcUp/cK76VrG0Za7GH+HEJKXWYJIjXd51z
6d3HRId/PV5/kzUPj97gmTQLv5WIVcT/km1AecpROaPFsoioNZ+h3iqrF4wHXfWkuhKcCqzRMmR3
nKO+4b/Szjnh2qwI6LVEqLThsoTFkGShXlQ4AwbeJcFsMbFtLJrMWUzEJLHQFkeSeAgASccvuiy1
OLP2+ihzEasjqGs1uzwSRFAGH+CEv7CmY0du4pb3QwLgxwkQ29oaP3hxwg+2bGyUfKRjQGAwA2O2
hR6ZXBMIAtvVqO7y9HgtpnwzDN6ep7LWTENS8Jn8Afn6hlTWwY3ujvzcrHgmdUhVzlz1N4sKwA+N
WsC/McwneKryJmnojuYLLRvh1+ewrBPhz+aJnlUKz2J1iyCGH8fK0C9aqaZ50+M1yHIhk8CMyUVa
FsCBxn/WKHQMte09Ijzdln4Dhs/Pjqv0er04dbD+NH06f9yG+WCYAi/BGM/c602cKMYAywJ+cY0r
zgWeamiAtAc5UwlH0p4+Y3EmofwJUJkiLW4UfzpDaWL5bNPJxKaXs7/jljT6/csh27PhF6fm7JP+
PGeii9pcqXb3e0EIqxrnCF91Rawaa9sMzUNdndWW56K9omppC50cgmVxutSuGM8pNSiOp86zQEAT
4V0lM7Xz0b0t0ZmBjsjP6/XOt6oiLsdXJO+JvF8DWXCbNRrxtWP+QtcsHIPExLc+RnMRL8tHQMxs
5BytJa5Xe2RRsW3ipuquXLM7EcCa+wGlR9onekplktvH2Wy8EM1aRENxz7ZNv+JaLIaZWehym52b
LNCFoUb7WrRC7A5uYhr9DLK8hXeMUddLTtU1f/N7BaAsSdj367tA8TEfCzE+X9kC9OFVvQPbuW/n
ASBtVdG+/giCsEfskPoYeUGsBHlUxJCWkyOUo3tzlgews6ZTSMtHUp2qCvM0/apBxmp47OFIDriP
Iy4p2ivmt7kujZs4171HK5wFUN7UOtAGufU9LTiEkODp+LVywoL6B6uSP+bzAqWfSjNkkc0e0yPB
VaQ9not8zC+5RpIhCcc8YTE7RjRwaUbMTNqsdYfJWFV1pWovF10nJeSzMsOvOnF0Dyjd3gGjdL0h
d4+F1hGg1CSnkO9yj3mokWidaLjjq4hpdE70Kc7tKM2uVb2SObshrBJVygLYHFbW41500igyda5X
nXa8xAPhDsmxCsQzHodeROjoawuhmVdTlQiRK4iCDOa7GoP9q8Q52cccoNqU0s29hOGh6JiRApSN
e1sqmM63qnnBxodFLuOf1OVr8zeaRYi1pw/MkRtfILkr1YVtewXeCZVVYwLBPR66kp4SovHcxKzc
FFf62VsfeVysAo7XM4bTTUO/uC/0m20axQTi0FJMwbPbSJjlEwEfY4UH/aO4kC56pJX+H2GGB+E9
S8DP8Qyc1nDsBlp36BICYydFBnYV8emxoEi4iUMcyDHxKAfSyqRXeZ7sLLsMS6YaypVlX2D57/t7
4HNgZqUruk4epi7ac5el6IBV1HhNhX1ustjxoZBFygYJ0//exRMxyyB3cKzypZF2shdopRB/R37e
E8PyugUTacTXz14aSFhP7ECJeGtLn5Ps19ggraNdohw66slTb7ziMB6t0Oo60JN9L4/zvt2mbM2r
AfKSD1n/e3l2X47zQx3GA9nWDddmb57Gi95fQi8J0UPfnxU6e3hTQ9qsUTrx8s8uEHzHVAx2ZTYG
amPVibM2yoLiHuRfgCrhCZkPMTMgXiITVfYU0zi7GdPoY87qqYQrDoTzlAbV9O4vrVL5+ePi4qeF
JFretOnQFh8zgEFyLmKZj2Japjq6chZISYLayveAqlSPNN6i0YbCDO4NREZg2HsAOKUKQy3j9HA+
oilBAOvY/uNQ4fTLZEfoKRCu8hL4D0taqTMDBxsWxO5JR7beyyuW3INvgpZaTqcfB0/Sey526/Bd
HiFiyqHaCScD1asrGLF3Oqv2WPacPRVbRQDPJv+O043kPe1grpst1GiWhz3xCWyaphxiG4hl63yz
jLLalKhxuLN/ggDwkO8PHKNx6uZwkrhQJHG9O1WcMixvH1t8bteYNxQKLSRhHi+2zWL2Tg4qfmsw
w+t0s3AZiZu6yjD8ETEg5cDmq/aqNr6mU+LhnBxgL2eTH8zjT59YmFtTbbDlnc8INt50hyV1vTwk
E+wuD1PCiAzsiLZUtiOBinG5OXucd6FGtl1cDrQYvpiyg6mFb46RK721LO5jiugYO2vFfvQwzAFV
majGGirmGjrGuv48+EVZ29VyEcDgnvaSrLhcD7eLThR9M3KoZ87t94+m4KwEJD3ujcHFEifQkAro
gJx2tiXh+iC1Q4FAjiqiO8J3wPVakuLhkbmi3zQbG0CS5QhQBLf0EOuplxFOy3gWBniYgVYUt3kp
hY290BS77OXcKjWKb9DfzPv1A29aRG55RfKaulKaTPN8tMK0FiCChnMPyP5V+zDLXKY26zS0TQ20
EPhfzQqOk+be4iBLl0DTgMTVV9LiZ5e+Kj9tEyxoiFfG44PXyK6F7IlnPLTXvwQHaxWEfxhmwvR5
cfruaxInCpFRAX4khQaFsTReZCE4jR9f7xMXaLKXezqo1NpER3UXKhe3WdPDtEI4smdVGcK0XIFT
A5MD83cUaHbL3+a/gn2btTzp1Oy/0NXifCkow/kgpUWW/uTehT0dIACvjqZzHKW3G43Qh8VFjwtB
zUqRU9qkl5Rt0I1Tb8WHxUJBquh+GRV92ykFp1ZTf+BR0Mv0knFepH9fggdqG/o8/2ReegbGBmAB
mbawsph3wJPT/DURnaQcePlFVIw79O2m3lmRAwiVGI/eWQ1L+qMF6KS8LRRl/63AbwjK4Qj6p75Y
a3QOTusYOe+sYruLn7G6jjWuGCIU7ZA1s1th92pE/LRp8RnQ6XxYssOiJ/qSKR+CJ6e0AUWK5dsL
aNpZJicmZ9UhfggHh+ftKfeaQXmuc3AdEnPakX5sEh7RrxC7VPUCIuKc4hOlt3jWj5TNIi8LTmbr
Pjw+/UF2A3ORdsIH9RNaj0l8NQuJGvIjhllvARl8CFgOF9U4FW4rb/W/kzgf9Jtq/VuPyPwyl8kr
pUMHwq5fIq815g/3JdTuCzEeKzz8tKFN8oNJXSiK9g3wozuGYdl2ILNikRCn0p9D8SaqvheMS38/
+DtyIlJpdhIdiGFt7xFrKwNwH0UCAnCvBfZseg2aBKuaInX2D2icvMgNlKBqVzMEGE8p1i/f33T2
8ruanD/ouBZo/0B+n7NbF2NDZBzRM964yuDERTZp6gIplBUl47jd4I+7qjIVvwbvJLcoHx1yFLq5
oIofJnoNWCjnVmgX/IQx5bN/hpm6XOTHl1OjY93kyKzTee+sjvRtOQ38TGv2F5jAv8LzVidtck9x
UCmHtqLye5d04rAaB8Pq5oNiHCsaA+uu/ZAVtEkanfNPwtXerNYxwxzmuX7iNO6P7Lxmro2uHExu
MIYwMQJbyx0JmscahsDoLCaIq9RjZ9NdCSz3EjTwEH7O0pE7RotNZyRXZxrprdON8vCHONhH4Ecn
scVafjPmZtQZifYDDmW2uRfrAS5GlNUtk/4i7MngnXFb2NezCYnZGVhLKqmaHkaDZB3/J8mYHHsU
1fie/Wg5mSlXpKopleKJChdjP3H5dDtlHTFx4Nj6UYGxEF8lnR5+k0cz5aDlTxUfnFThbyVqp67x
IZFhscxy7ioV6Tfmj9mA/YtlYYw0jo41sZovE4RlNGGybiRypRRRaFvDNY1LZBctUvu8kx8r6EHo
TdyElpW1Xp6GJnyFfik2+eIcnnPxSVX6OsXa5QdtB3rqfXdWe4ZZzI9aNAz5i966P/OYfKcNB7xl
Uhmon1lDk5iyxq/0JOHT6JRwCWr2VwjwnTPlkJoA9PVcRktkR71ekQdr40YoZZKiWeHyWxO2qktR
NULD7UNFPBGaposuwLfN0qVb+CK0u6sb9XpLugPz4bHPfHVIBuzUTxr+3wH8Zx/RILnkVcOA+JAF
alsXTI/hBc9MNQ5OMpL8hQeLEQ4yK/Zt9LfjnzzSJlbw9lvzHaY75TO0k6IxZaA412GOy84jaDFJ
Ux7ejntmK0WPcCKqX+VJefj5o/gOXPcLHJ9JT/2x0cgtzt0qqbuCMwrq458e17Xgt5iyofCiXnmC
BtbTL+lRPeHKO3Er5FpdGiR8WUBf8MFh12PkNGzif4e6sLgm7C7Jbm1nGIFEa660iab8F0fLPZI1
n0JQsFD0OdIRFHNZMNnk+fcJO3oB26TFigaRTTul8efZ2JxRxokRECy5fFjvBLWyNGYpVRzItqyA
ZjQx4pN3Bcyk9rUX++Dis8JGPWaDyOUEZEeLPsIFHX5IAn18QQhNTqlVhSexmS5yo5GSd4d4wp9z
J7UaXRNn8H4sN9YJJ6cQ9Avb4pEezfp/KGB+uHo8tC3yxM73ErTpLAxjgDUfIcjx5Vk7lFfNccZ5
eFYE7H+EOzm2Lo7prUmsB6lL3elOpBINEpS0HHrC07/JHWcr3p4scS7RiEma7sogUMBs/l8Fwdah
QTtTJ0w4JRW84QgDZk82S9pH145DpiIA8vajvJ8c3tPyQWMaIh7kdXtt0jkDJ/qPG/x6zYFDH/2h
ilUtWyd9kOeg082n2GVTTQuaLlOIf+oVK8FxAtoz25v0H+dXL5LY7malqN5112Ub+aAKWE/RPRdO
EkQhsqSv0lUIienGGxAMx46/AZC7P7O51biY7drajTsRmm11uZz9X4BmYd5WEqwtivq9m4g1q7jT
2JO0gQWpC86UnANMw0ohkNUixNpsSge9scn21Ve6QXLCQGDCgSAu8DkugnYoM7S4FgGNELiQtqXo
lcACVn3a6QrjLqFKAr1HY3Ek9XwV1KQVBuBEFSMnNsNxcdvva8znQslggea18VwAL6/RJ3XpkHen
GjgpsBM04p4+7eXiNz18mnT9d7uyPhXO89kN2hi239ffA18ztwZ2txBSg+edeaWW7ETNumXnfCWv
ZO6JgfzCF5HKB0CIX05enpMiNTFgVVCVhI8pF+nDP/Qhsg+BEBlw2/cOtU07PVEiqXjt0fI30y33
VCkJtIKrvN0rAVr01h7jtLUykM7MFna11JEicmKhIBvWFJXqyYagfmPVea8ZSv8APcjtBgVBDS1k
Aib3EuWUHel4lyfCHrIwsG+NMV2Q8Mc93Ebx9p2wb1Rat1Eu8uITLyd5yizSovUJA1AJl6qVO3pP
je7Jg4ro/1TCFv9CJlxLEsw7FrmJBroIqwM+cI6eWOSPstOqP3ANA354afaHmLk5Rsyzev6Skqf2
Adob8FkdJNV/o4qsSpzRJZIkhj44WMC9rpHRo2oToEJHq8YDa2mKtmAIM02PWc06mmcLHFYiOws7
c8NQI9boseFIcoT8O0RtbVVd5hexRYULBrX/3XTZlryc66TK1F46DiohZMLqonIG5D0kQZ2GHS46
w0oiI1KN7rn7VSLBlJXLXId3ax3HeXN/zQp5hBk2irbQATXxDHlnLqjm+ddF+FDlCyOeHIGDSxYX
dVtP/MotLo0XXP4E3h0xtiV/c5DFFWOaLKweF0I5xkRHBTw45GsH674owM2S2OdwWpFQFcQTN8Fr
olKBH4i/8Ffg4IU5ZlBz9mMVYL+m+F/YbVigLcUp+LWSL8LRPjKy+5DkuAXtsSIdo5Wv3jjOnSh1
tlW8bHipEHsjKapNlOiconVBkAm3mlOi1lfXphRyFiKOpGRN0bVD43a5uNLM6GgBWIE4FJwdUGlU
vvLpWm1hSlD5hNtyfc98g010WI/OPMPP1HZIQLCUQ1oGb6eLPZEhfr8FKQqYcjcTAXDXNr/0MT0k
cz5380PyRhJhUgNERGnS6PkszI3UgQVM0SyC+EXJ2SnCjc8B9ZXfIcqNfUsIOOI4gZOfpAQL4FVw
vOJk64ZgXAxV0jhNXCZovde7ovVEpxmAIuJ6fHiV6vrJ3k/DZrVZSc6wTmly0ZYHXNbLMNrkHyT8
EI3QvuK+7bckHMs4osFZYKFELZUcl8lonPyF+sgRk9wpPX38uFVsWk9K28ooAnORZ4YQugKFyMbK
ELq3xxcHaWor2O2Lw0FpSWl4a59yRo1CyZv8yByjSstRGpObHM5+WfxxVtp5FHooste8OEtwamYI
3Y2mZCCs3ZzQuzddAQxmaBrxJdr4Sx7BzvEbgjuTxug1VBHImGref6YrUUahYHz7krpEocZoLoWK
6DJZI+5fxPmN7VsrpeV3PtRE9nx2Ff6lcOY9FU/A9k+8+X56Lw8cguUlATFnpUEUMpxINmGYe/4J
H0V2oJWIT0woJNUbQeJE35Bd0/nHB9OgWa8d3rRMQHp4IPY3DDfk7Cb0Q7aQJILVyopTdXO43U++
tTCDWk0cQl6v1uGwF/G3VHkTdvzvlox1Vv098Ndpih+xdDmfiCMMevQ3dxCk0UNnzHNcClngGcjJ
R4FiurqP01B73udlT41T9Axrj2gmGDxk8HIMLiwZ7DFsMvrcvvFwfk+84ygLjluKj4w12nWnilV5
mlM7KAUMbty3JDK3N0sb95Qn1xRK8Xdmd3Je4CM+4j6oUMoP21uiHdPlQQcfbv8kgAM2Ee1WGjWH
GBw7+rMLxB9ep3txQniL6LtDWD9FdbGYtf/SMR0vBPCKeX+IFDO5beV/NtlwTZtZ4YDaPbcUHEyE
rbopMcosdL/EUCbtkV1isijzYqPalQkhPij/K+kdEZqkJC4ABEA8BLJBobcvssj9LknTRJPjedGw
srY0J2pC67VMgd8nNbfS9gf4wRUMCDNHBlra3OrJjvoHJOTxcpLWzRtB90vvaleYzNDhsH+ZjrPF
SWH6yLtNCBT6GaoDInFeukNizIYyaW1A0aG7iGswVybCZ8NrO1x8Y0FMKw9+/PJOrxy5B5FokDbn
rubbAxg9F3Ld2SDcf2siA6VrQKnflBkGcShy+kIfBgtZuGmxDDSEb0SsWgPrkB1xD1F3w4TnFiaE
OkyVrI9IWYzCpfWK1p+uuRovTIwpZBX0HNi/uygJMfGlh/TWtxq+5bqzkRqT90hWvpMvdzMlSBA8
SmwYGaaXEPoYN4Mbvfgjv3T+acVTSp5u3Z8fBbi7BiX9KoKubPdkmrYstIxcEiCLw9/KRQABwHeT
6s52Ee+BwQoZn2nJzdQEKj1zdC/VxszaL19JbxnG06ikmBrpbUk/2GdmmB/sPoVv8fqgaipRVH4C
mEgnbxSOYN1K70Lcij44MjjjbI51KowDXsYCmX9nmhjSeyEqdw5Rbyb+CU8BRNAkyAjAPwuC4I+9
QLHngomWRE0xNNhS+s8AfIdNjU2dcvWBdEAbACXf3jF77conFeKA8xDl0iiyXQTG+Z+K6Bl6eB+L
XwIFv0SLwss38RzaaIXJwpSUtVhi//njsSV9BNmUIk4MvGaKp8MCfYYEKNWg0r7wIMDiDFPSVsCU
ZyK1yEIWVKo4cR42CAvJnGECqkimPNOJKpXlnAYmaFQChEPMJbycPtVCfbWW831OG+NhpDiCWCVP
0zaFiCmG9nW/ch/xNYdKzgzjuBnXRXe1tUXbnkH0XE2Z1AzTZFJXtBlwGMhyQwMv3tRSNULnEZwY
3HP9X3/B3+IRQjFo01ipTtik43TqgX+n1oR75cbvVD44Xds+XtGpfiwCuIXZ7W7e1V9SPZGmXRal
rs+MsRHDKPkwbKxBBdL1bSPv82pAZxYAr7N8lNq3fA432mvEDlEVeEdbD+T/M+4Mvo+ELot9/GHh
ihlng0ToTWIM835UfH80MzCXFAgQg1ILS4JBEFdhQoGuSDIp6zyZdt3VrfD8pJXiEHaZ14w/kbNA
mj20CPNYdAItzBp3x/ZhV9oTEYO87Src0TztiaEW2//OhxRTSj7ipICACZeG+uPBG2JRP/VwbM1A
3swC1a95f/iqoFkRWgA1whao/UCvoNTyEnZJlwUKm9kkMK8atjfd3rLT6dI4UXC46jMbIeh+q4jA
56RTtGd1akATQ9DLrTsIV79HwOTNy64EdLtlNnnuFxfk4vQd5RvgV91bTiQxah2RkpY7OnBDI+rz
Q6C5pvWzQgoKgtZ6s3MOP/jHHbHqfzwji7bpJYJjITfo06jkSnjEmQf7Qmy9RkJIqWmohA1HW2SD
32aH1SBaH5Zm7kfcRLFy6wu34OxOH/dd/cEY+3fFBh0umGSxNkL681Y7Cfu2cUp2zqt/BZAd12Fc
LE964BXw06MN1AWGwBvsQ6mQ4pdVK2a+qN4cTE2D+dYLKEG6GaPI88jTKjrBC/MOLHQfFiKyTIOS
B29JLdDfHSlqsz9PmfMyj0pgGEo1ul3UwFtbBYyD2pRE4K49vLt9778dSZYpeKRECJZMh8dItar5
WgmxYWaSq8PB0Jpbq9ZAmqT/bMKH0dKhBhmNVWldjiZkcl3WgIwE1g1HbpbtxI7AqgWw+qjClY6I
WXFaJYU/i4sd1v22Kac8HbtB1Q6mZEXvKwoESe1SEn4a44fZ9Wq1TOMKgxsK39Oakw8i8P7waw1p
2b3nlalLS/Bx69h8pwxVRG9EBz1cv15w+tpXnqT6FI9ECGwEMoN8NP8UNuXS/kaea+qyTqoQH7Zd
bNln0CdQ2AW4O1BKjrnmgIs0gwSgKwGzkNkXApePzpVewmZtPiIhR+0zkh+h8fsE7jb5YTpGVXDx
TgAdSjy1omoUA/6Szd5KW5TcXWWOS9YYUC+FyymmvSJMQZoyjIo8ayRTTKUdy0BJXPnBjpZjvmau
0sMrVe0El8QauaPvLXHOu0uJA9YKI2Ok3irpM2BxLEOItjUlZsn27R1HVMa6R7juqKMW3YQafckt
q/8endjHeyWMfQtH/qNofN3Znd37uLp+PRnSiUS58MOmM6+UhyQO3rXR53JT7cAFzFxPpeWANymL
0NmuznoLu9N/iEsKq+mEkZmzmuZgSjfbkxOe0tmAuMMmTYlrBkw831qYMX0TX2ZCpIqlqiwuxRlx
xYEhiZbQ44hqTzWoe9vYyHP41Gz6NkqBFXw76+n1scT157SxAwk6FPqzjm3lpSwJLIVxUaEnj4UU
gCy+we5clGePx67CugbFIXvDu40DHimROK6SaMMmmaOCGOSbVKjCCjLq9B6b9Rhp8GBn0NoScxvL
xxpZ++8nqQxInTvLUfsC9iDR+iKRHlXgMPKGzebnGUO1ulGejORIZL8a9HC7KN5RCQ5Tf+9Rbp8+
Ul5UfmGLch9cqYtGE4nZ0HUKRAwsVKuEtdA4kaUkDl+fEi556UeswamGNgnIQJdrwglg5H3Ig9bT
6K9T7G5mOOLZHPeu6xF5mlqm0poTfemRyo5TxWcmaYTFYtON+Uisg9FTR6UtmarXfUVLRmDjyzwf
4Bgq2kxc0TCznAHsRNppEldA1tBsAXgE1f1hewqIxfZiPXrYivMmzlfHfWstu8wC3SahNibELUkR
c8pwmYl846wFOBSkqV1FKbvM1kkmZmNezNyMX6GHajXYuOdyq1DBLfRPdmjBrLyjoIiD4/81mgE4
kTA3txeaFx0ZGBpZdfPnfn0lGE5O2GMBRrQ9FvbU+WN/krnlirJIpIcI59nLMPp2oSlrdf30E34M
pvKIA7hJXLrZ/bs+Rm5VYWyvvqAKXlbsBds6983r6Gi8UbahJiVEVbv67POQQ7jPUNq7I7RL7lO4
yWleV8Zm93IamfD5N48OFbTCRsEr3a5PMYQxSQbfKFVl9aEgWASJ/LKa5jUP4bmHEvM7KNEUpYK0
5WTD8ifpUI/IXsBXCRlGKgGzvEWz7SNx9IkFDd2TYNO03+YeRvQ5NyjvbipReZGTd9JuwO+g6cY8
V3SoP9dQkUvP1bb3bPc9j1ke9OLf7+8qkyo8y5GJL5fNPmRcXlwPs2BgJDEFr8mzVKYBEINebc1F
lhzq7lmIsOd4XmV8k5DlN5LJyNMJElUiuWJ4SHqcPK2nz7bu0v0Jocmo1ZfqVBnVHdUlVqKAs6Zi
6TiVMgafBfXBup1Mxy9OGBUXJsl5l6rqjTshpEUBFqkaGYXnfvGJ2jAuQjvAr1jiv4r3I2T/dmGW
FMxXv9Y4FdSssR4wZYFIxnykiGPQBQL1pPOK+hqzad2Qk2m80/ufeYNPN5wUh9l9wnz1whT/wZPv
FxWerpZ7I7prwZo6OaHfK4qJuwk0ur6+dXUwuZt/7w7CgJ6HBWeT7F/7s6f/9b9hhKMjjayCI21j
TJ4AUKRMqo9ldqrVJWhQLefTD34YW4ly5j9IguZ/WTd+9Le4wzwnJ2TwtJojxEEfruqChZY0q9b9
fJlb2Uv22E4JBGmoZnXUYEOl81wjEr/4yv6/MM+rV1P29OGT6scFy4AuDhTg23pKhn+o3UUa/Pij
YcFNBxR+PMSJ2x8L850nRwuGNbW47oU6mEpsPGcNsPcfGFSW/2QodDWT1Ym/yIJkfZFMCJnZAwYp
NfhuWyUPJlrIWSP7o1Ij6V9KTvL319aRuBairJlYe+BJ8K5B/D2ECJnsfrIrawkj/RvNlBWN1bu1
CfKYQK0rDn9I11Co54IPvQy8M0VRW9ejRt3KsgJ9irF2OTSW1xta44UvYdXQ84OF6g7u9aEJ4ID1
XTzA2Q1dK78caJmDy0JkhFIoMM7nNuaF1GZCAc3IUjJdKuNqv8WLfsyhyR33ygErsxeaC2SBhQf4
CXA2sY3cSxLmsCmRxo9gIOCE5Sz0lvR3FNFsdRNd581NBd7aBaMx2kjc+2eIZkcGjsFrWj5CIFCe
LYyaNfOtQU/r8AbtW3sKxZw8LYwwNuT/HsjPTRjpBdKV47WRr/+nj+JKafJnV4d9cDx2YuR5yKwF
6NhsH2JDBmKw+c1eXca79jzb39ByUtOKUVwOMj30zjR0JiiwSzZqzkynwGHqPjPdi/Ht4bmPg9Bg
hXEi9K9fuQlxBYNPmjjX3VyIVyo3OfGxY6zf7Ze9FfLBFsn3gFh7X03sXbj2208pnl8Dup17Xjyo
1nHvXdYDI1dMv6ci5+irv6pWgzAnuxt0LwAfDvlnHxEsw/dWHfYQap7O/NyhEqW90kdWI8IINx8U
xCPLbjBtPivGBL/vhkfn4eilVnSQiOZIAde3mbsIVw1oKNJmI2DjUlxzk6lqivplOf0AVMsibA6A
3JY0nFbegaSgeL0RK45NJRC6XB6OlAfqFSErAnSS7Zxd4SOPEcFPYRjSt9i6pno9DzXS7g2zmu9R
BlA29AG/PFuNbDMdoYKOmjOAxBBglnqGx2fP7A97OLHOFRMzVRFF911vU54dOrV7kgflgyDkXsTk
eUD4ZvTOdqKxhqk1tta5bQypQpiDo6viK7w+8GsZxDMpy1IPDWdF6CGQgTQ5hciV5G51XzJgP9jl
cvL0+JuKq7Ef2WoL5zF6rpUpq1n5SuLA80JTXW79yaDHXxK5E8PMNrX1Gn42rPUfaaUmAl2xZg67
n97fu8zDBVm5g2aSNsAErB56rizNxf7lnPQY20xLnMX8K7Pz1aKZCbvupIfB4oTIHI3TkranuXgy
XtYfitCWzs27JeMmjcBB8raAfSPiqFfsZpugfWMRs1knZYSM+0Of4TlsHZF8AD4unJh5n6sufn52
E4Ao+27yvbsCo0MWAlns/q3VqKBAPa4J5crFmgR9Azz24wLdumFntj3W1RkOUJTSY4oDCqTa39uY
hJvL8KXVL979/DQBW3XUygqFa/tbmRiHzqPMOJ8Nno9qf+fUGrIMIo3sXwFFnw9UOwN7GZbUO6eQ
QVuCt5YCxpnAL6ROeRdHOav3Qz7oTq1bOIM5IReJlEvlsjb56/mhDpBfroVNjO0a9CCfcR5IX5oy
GGA9EABmlDsWLPGnvYiSKfkU58Q3mAqnE2LMkPnwZVAxRijnqLbsW6G42Ul/QXmzUgMoJQa9R59w
cLyde+uT92Bx4mvgk4vXQm2xJe8OBb5yQSX5XQEajUz9eBfHumaJRKeifUfZhMof5Rbz4Whatp3G
9ybtQWQ4xsG/bKEnZ/UW4rIrzJwh7NtwnEwRK0vdl/qRpWoRDJTfvZncy/gtq32rUlZ+ZQxBC8fr
VJgOgvh0jLRgw3wxdsuM+WyrjIOnVd0JM4B41uqJKh0QRV68vGFFf/a0foTFN47EG3rpx6dEToft
eFOtBClAPAznoaky14ovT6+BmiZgUL+0V7df+JjHP0T0k2SEXxIwaNIUo8dxnu+u8o987cb5GiB9
Kf0VuH1cPXLux8aoWeADu3aVUhb5olh8ffMsAGgwVvOWjWLKG7/v+eurEnSfOqHqwjb3u7bJ6MLm
jjMZeoX5JU1cUuhZ1X+JTHUANNK21dJ15koLxLO7hcwZZOBUQ7sVb6zL5/+yy5vV12+J4Dxh/7tq
MsQTYOoupd/FO3DDREHFSXXva9hEa3Od7W72EZmXjXfiuBaWDqUETy5eMCq7xrf/+uE0WITIGDnA
aKA2aaih4WJZyOPrPtBFUwaYfvgcQiZcnTidC2pgLPSqHk/MkGUemxg8FW7+BZDbAQ01IDLFGg2Q
Aamm7MoBGqVx3REx0hyfDQd4C4IewkZhuWbGvH4Aphghqrq7BkHH8Plrzeu5QnmICokTey5tpSbP
1eJqmdGGAxwjKBDjZdIDQmazF9yUhcQJP2dv70pURSBnSXR7gC/NNB25906qDleWWlF9HA+jxH66
covwebSHTPCABrJhwiZVJOuhtZkZpvq+4BzbtWQkR/l73Kkv/FHC8VrgLHdsa9yzr7QwU1CYpoDp
igP0YDaPib5Fzhe5o//lun/Au7TADbRoVPzO1oayIImwEqoIs7BjgmPL6IXljrTw/3uGZjpOaHAC
Z0IYndMnDW0mM2GRvSAz5D3HQh45c7jUD8qGVeBYi1XUcak9UQbGtAMezKEXEBC6fQSzatoJd1PV
bF/adQZlYmg5UOqNSKke9gtcSK2enm2HoruuGGN6KzilGhCeb5htzUNf4gmVpBsCf+VdL2N+9lmt
VMGC4ZEuFEFfA8/ppDdiDb4X3exSrxgAMyNdd1YLT++4RAYJxOHyBvdw7AiTWbadmrBLGTZmH4BG
xBKLh+ixBGT8Az2yyFhfbudXWPfRYs9nEymtQGdaMzb00h4mGFWSvkp1yc8jKY5mnDHX/4BwxvlJ
YjjdYLalS3ba553Pa2nqwDoU57C/yottD7cNNh2zS2MCub5numJDka8a5PAb85Ur8Ie3O3CtHOgr
zXiAoBcvDvP1MNSwGZXRofVeQPX6tI1N7VH+xsKCK139SUOnEC7XVleDf+OQGvSGt7aycot0m6+U
PoTfc1ziFcJ9XcJVLssjsZWTtafTYuRyve4ANOmkxm5ES9Hw1TZ1otqOnIi2fE/jvo33caEd/CTb
t+rxYHhHvdrJf1aBKqZeYdIoMd0zBHEoKRZsgVmC1RGYakutoThzJYDioPHgRkLtBKRJALtIhCG1
22Yd2Ce7uQZrp1Ez9qrXTMGM/sZPRtgzRN6lVzFwr8Rkoa8nmArIYxuQTyV+7U+YOoS4cr2AqAHU
oODjDWY5R/v4ukd+KzW5iHgOZWwIOBTrOP3DAp/UT9tY+v56vN0AOSsHiJpt3gyNA7GjGwX+UjyA
W8//k/2mtftQzRDUWT8NxuUSyGzAGhX6TWGv14Cn9xZss4mbQsHL3KArB7UHZR8nnPXZtrP2MuaR
GFTpMLQ4vC64aWdR/H70oCl5Twoq6Xi5WwXbAHEwzys4ytOPLhuqhwz6+P6aYGW3d1gvL8wBjwUE
A4D7IbUnXPFVcCPOCxcBXVnvHmjgeME/xQe7DD7GXBG+ZHttkqtx4+BJPzT8Bv+Bp43YoYdc/mCs
//Uufht8ojhlnvp1OZ4yqCtK4pCAnLk5mtl1zTe4hiKq/OHmllSpK/1YszaALRD24v9DU7Y2awH5
+KOigx/dCBPGzEYwIRb8I2SrUOmLCnyaW8lrY5kg365b5WovfioxQcAG6jiH8FFnp/Pl9ITBbjF5
1UVNs4Hl/VIxaozPG+1ApNhwkMOb5cMQqOFlLCpq+CmKVbwnIQtudTJGjtSmxG9esEAht8to68rg
4XxZtSRjaFbVN7TQszsU59rS66Xyj6AWGKiGYVuIyeNYfsQfuPIRjhPy8vdQewAqKBCZTFnwOdF0
XN7Y5BtZPbxRvOzHaLR1kZQn3wfVrwE6L2NGKOpKrJTRRs/yYscmqO42iACVnafXFq86d9SpD8gT
X8/zWDYjYSu5q7ptlLAffyZPkeXRW+VPBswdG1RDe7mzaHMzBTxZblGRw7nElXkVnSn/CeRxCelh
QIVxIPqfjd/UBw8w2Ir2y502NaXtc8N8s3ziTlGE5uvnsvBsyspj/UytQHCT7bIHr7JbTvX4r487
duSJPka5QW3l4tZxYAWgvxKUrEBHA68yvNOMNVD/19dbqwABbBHbUvTCmVDQDfb0shq0+shYU9NQ
n11f2fHNgcbcxtBML6iaZ79cUSPZ7jIZSW/usX2WrV9gt9XyKBbmioO7FUdpgDtEi69Y2ff2Vk7D
SkZU4YyH7qQL8S5CsTIOFRKvz9SqxUHzhV6FXQTUnUEN633j4vU4eYDleFtZlC6gBWYH/M8jnTjp
rzzROB8D+D1SC78f3S9FPOis2xh4P1kWADkLzzng2CKFU65CMbkq740wCfk50S/q/ri/M9963IjG
y1AuiL67KMgPfDYXCptK2C7himQBGrgJ5eiLyERRdWXY76rggvMRDmDzqS2z7oN8uuNI2snFPR36
BMMxTFpQILNtX0o7zFTNelpv6o5Pfm3gxUNlGbWNgufejMGTkb5mD338Bb34rOIgR26EfJE9mlpc
XmGUpoitXJ3EjmBpU52/JhpirlAMFbHC3Q1b90JJDh8Ptb8bp9WJV85edc5ZAFrqaq4HywC3zBST
xh89ZBGfzFTzhLpjMwIB57C54exGeumNFaXxD1hkRQzjUfSSiwYv8CiEfAdm6+d02sX6aj+m6vAG
jQtTLPtlHGxkAEM2p6UPdsYdAeYVtQdYTqo8SPW9ITqVOlzi2GDRsaMXHcaWZWErs78OnWS3AaCd
xZvu03PXTXTWCjDEmloz38fpAcv1JwCpFJ7kQLZU+JetnbG/p64NKaflDqkAvtiBoB7v5uSCDcDB
63yhrk/ilUg6NIZFMMb+Hm5pi9Uqitfi82RGDUCO6qvRU1bBFH8sR1qpHgdu4WY6CNTBRP9p6yEU
Er9X2Xfqcynw7egbwYvVnglnZuKeZdTIpn25U3T7ysaqwM/IPTjk0MKrJoE4JWyIVQWzocR30U9d
OpTp9BtP/SgfFQXh9EMFGPLuqiUFiUcCr/KhQy2exUap2i7E3Jw9OA83mQGJ8mDe9U7QMOVo0GEu
MaS2/ABUTEHGnElF7VoufCnBLE//reKl/0m3D1Z9c162AEd78piZdprkKicJTY5qoeYXmW6YlE+r
Im2Klo/K+45G+zhsWX4xgd7ziNjFxkR1D5qm5Vx0sAvAIQNjp+w0dgMKz1hkyC1w641n1AUz1Iaw
yVjSsagElhykNvdIr6o5U5cm0wPzjMnzAZV/Murw9Yrn3BPz6A0xlD4Zi7YiDM9H2ZmcU4GY0DAi
5pgDqETG7RSOzuzzLlqmfD6sR9MK3fuX0dgfLXXqepWTYOk+H5SgEqaPFm59Tspv8Mxwc30Spe7f
MKV/JtDkrccfpiSFEzBdF0MOAgRyTHd3Hq/F0/AFe6NCKJxVI1OSJ5eMN1P+emWCAslEKJOEQ9Ed
Nom/CyEFIyv+9gwbHPglWerX7C3SZyfrbpUXx0xNVyH8yZAsG6mcMPFzj7DfQe8Gd0gkZM6t4pNo
+YmVe5tSNZgldCBP/YR3jT+b/eLxlCTJkxjBbgxNG+yg1/N32SkpVYgsc+3dACHWS5/j99zZQuLG
gz/GS9oYsg/xkaXrziVNlirZWl3IHsPt2y1NI8tL7ckBuFUyKoZF25AzZwCMkt9xnPkaV82iKCDB
FKxfFFIfNmMkHDimKjANGlnN6vKcQYUd/k8VynCIMYkBF/dJZjd3rxGGSIawYfyVwOdfIz5O3+rF
VFW6Vsn6WJRvGlAduAhdvZP6UAWaVJNICI+NoYZCAlh4gP7ZpFGZXQ8qalBJU1aw7X7WpXA0TpJ1
h78q6PtS8w4HHwJBvPfooAXKc5yU44ubiBtifTXDEpgq1K6+1sbZz7lY5dWxRYDOAyoMRRFBq+r6
fN5CclNyUJZLrzsk4BKr/5aWdOxTGvcmzaTfNg/fktzXpZVFHGWNzbHfyxT24O/xAwUsE30i/8H3
FIejoV0NGWVvF5Coi3MzzvrAJ5QJ70HuPk8u4LW6T44/XP5p9DEprsqg2mwkO45Yq55gd3X0QMbn
p4ilktetFSq5Chb951S78rp8+kWtEfiBF/HFrWbD202gxY5/SDWZvWtVnTVQUY+2ftwfNZcwgkr8
AvdwHPCXbrmoUF3fkWBze7k6Dj7GuysyWP0/DE2+rJM6jyfgB3SF+bpmgRJRXPvHakAEhf35wcEu
idNMVPR1mMOPoCR4EEm1oRGhfTLv6P8VNb6beZ8IdRXVY7F9UF0IrDco5fn/SCKeYnvi5vsmv6KC
AqJ91wILdXxsMOADvUgBXuaWoCWLEMePzdonzzXlvvOzVmrQN0FwavVY8rryRs0sq/tnB1XnKUfp
bRVzEpsL0KaOQ7r4WrEqYJYsNZTw6a2ktqueaS9J3MLsUDBjrtexzJzrdqt8VBkNyXrFz28CHF0M
1O0O6us3+Shy2q8LlRf2XBYxRXc+ej4Rx2AU33u15DMM8w4i+AD//HxWH7uh2l1XsqzvxJvFQSFl
GEzHkMmBK0JR5rFRy+rjtwPzFXBgfqMZr5pZvQeiTGDGsLXxYPIuLrNC07MvbneY5S6eKUM/bx9f
22VcJ1OKKQ67OPBnGi3CJ/7yQXoJWtUeoKeY78fXHJXuDM16gQmeyXLiH4J67WgahJlRC7I3+V+f
1eScs12ht2YwC2L4xeZDlYiZ9nzxRIbAKk2bAWF2BrWkSqX0pHAv3nCDN1XydPfYEtqLGtlL1A0y
LaAIxEnyl36wAta7x8FpT3RtV6mA4KqZ5/daW4Frmzmzc+CVSoT4GkEyNq6SgVTPtLkuoeA/gIdl
48BxM1BDAz99OGDx0RKE30MD3qbeKqyEfBavs3rR3Gr3lmtUm+7odBNGiTbxT3Nj0mXiDibPs3gJ
ZJKGwdzSZUYRPVo47TQL23r8i1aUaL0KiUNVsa3OgC/7huMfgC3mWVhtrln6SXYXSCWJFhdkxAm+
W4vKfx8v58+Kre0jEQpxF8cL2ocaYQ9nT6yThQzXbYZUlXXYQZGogGo9hN6XzTEWOnmUGTKx1cju
5ODXTQknX+L70DFtRkb0OUmlkqM1zroLKMZfmKLK5RkHxwP+8uIOCXPRQ4hWC4UeXj+FSrjMACWk
KvpoK26tmCMQ6ARdGy54jtpSnP00Un4xx/z44ra2zTMQIoqsLLG/BVD7rAJ5F1Oav5Yuk7xRcKta
pb9aS7YsAZZACwGnV/dyDUV/YGretWtbJEdAAgw7pzaMwCqumbkYNtEJYssdeMt1vuhhM2NyQxfd
ic8tHNsEeeaeBVxGp20FKXH1UZnshOSmAL5DqfpYo38h/3gQIh7ABOyeCfapciTwNgghGSEVs8Nm
JFoHPnDO0r9QhYk+UXu5NYq9NddlhLAvYuN38O6f8cATemex0UOriCnzowr8/i9/mlnow7pkVZDx
jgK/2wk9OocjS08PFUyDPdw2kQxj4PeAseKX4klWmUUCdPZQTtIHcxVTnZOPlvF2pDZUAuUxf44e
uWHJL2vPzWLlruvPBXWXkHQKOiXQhJd1FXJDJZlg2HlfANe+nVq/iVXvAUkvtW7fKJrKIbrO+Vmg
ZOP0ufyU82kTHCeI6wI5FYXWtvuIExMfTVlWFD8UtR+eH94B0zQVfvigi2y00QfF6JTvrkuDYHGS
833Hc4Ul1UkmSzm2McY3GxnFhWj7mCGV2En+UBwxMIJOuuaGmYaSNgKNKo1KDtBpfaw2u0moxhS2
4GWWJmFGPLeTayevEbwPPSMnQ6mUyAmzxB9gXu5RqjlzsfyQIJrm5WZCwRzud4f6t1EtJy8INEPC
/tRoeGBJFKcdyoJAknUEs2DeC4/ImvgSddRvmBhnKMTMbDLJEBbBF4UDU/D6TEcapJMh0r87k3Q5
4GizUC3/ku9TBYMpq6eX4wnZvj1babHL2URW900YKUPk8cpcbZo8iMc/XkubT8GUMbJrnRszovd+
CdRgoX2/3x+EObK64BJ6LGclIQ/Y3OjVB5b3d4PejhEeYSuTZjZCk+yIkMLd5u+t8lNNBavWXAFg
Xo67LjrbihtOGUSqdvv8nJ7yUhBrz0rC6KBCWBWaSDaqsmbmRSkHwN+X5sYlHilO8ocJn3rXaV2N
/dSVVm5KCfzBN/+iT3j0csLwhgLX0CyTm0WghwHY2M8kgNBfqJd6IL61xfxpTdY1ijxR4wt4vNC6
xJSe+r8RRvPTQNLoCyskDobWv4nRCkT0cwCB0HuVL2BtDG0uYoCDbe96bN7vjG6tSDpVmioXBW11
EfEh6+OolSDMIg7dRIjaQvRiXmciL+IgUnHL6eQpA+DIA+av0q1KIsJDdRID0P/W9Ku2S0v17+EJ
wzE0FIdLsLOcPg/MeX1wjeKMOwu7b1RtYLXK6jiMB/3JXW+1ZpSceZdAuzjq8vfbjPHqM4+y9y0b
nYbDoyXiUN2etYwM7jRdYPVr807OuW1P1sPVEHqTU9/t1+zCjkxpJzc7BeQDXuah3qjBRW2TCBEa
sycgYJqgUV+r6jo2+6fZxn5Hf3MNRyBykTZL1ReJ4d69w2ZQjBlGM0eooXMwDxqEjiRZA4NS4O5I
Li1ytfB0SUv4qKaYg4BIuXYNNYqupSjWjDLcCcSNJDJB09h0l9ELoLVNOkev8/gzZ/Yw/mky6B0y
kYfUcwtMfbjJ7MeScS+mhg/9DmVHnz7ZDLE7PGaiziLTJ8gPhhNeI4RthldbGJP/sui61E3KBOXP
tXlbVn4jS+qnSV/nud5L3OsSKirYtH6llejykmsOFXXOUC3Ja02gHyKkjXUMSoIYq+0o222TEydW
ET0uy0atwKdAs3AMmXnOZ0GWNpR2XmXsz8SSvMvz3j0A5lVPXjDVku+qQNyS+neK+C4PyvcCiPxK
RZv6cY4rBDNUkoAXh/m8Q2kzRrmOfLt8NzjJPzSra9ULj4p/WeDAdYQDWGUfdvEkxplGAj60dsCe
8t+1I/s+FdrQ0h5UNxGplUm956yv0QtRy8DYFVkkK9ugRDdaaad8+DBhuMuRT9TMWKqPG9KcNy/7
PdENXNHukqDjmCJJI/ssb2/SlzhMGLS2hjBpCD0F8zap8l0IupNITltHwNuQiSJ8FrWnR8TNmfF0
CJygZ5Lq6Eh8QbMZrs+D/pWxUJvUTb3J7oTu6bahHBxXOkjNQ80mDidjsmcBnWjPfs+2x6MPJEvD
wC0HLKDaAEATt5vHf/9/b1XXvW2+ELlpYheM1PSPsVXhLzAqnXJb7IdtB0VftC/BfSRLfai38+JX
Q7wRTHj3k+6B8g6CTtammFCKI5u8hULpZTUBKNiOYvLkSeld9bzZiEEp5cmwnfaW0TN9sFjV1F41
2FccPdNouPGYaBed+YFwNekW0+485uJl8k3yfojNO8yaBD4J15wyexmAlHptgCR9n8/Z0J5j6Vq/
VTY9wjUL9Nb/XYYAx5n/YRWjyXEac6mFEsvxoaOSOyOgJZtlxG/7f2kZKtraghcRsoZj9OsC85Sc
UtLtYegkPanDN2UYfddzXBbmaWhayuZ21E/vpCdi9IzSte59hzca5rseJfDOcIffKu8XpN8mcWHQ
cGVC5K30Ua1QLoKFc8vZbpp0+IGt1mbQELs9QCUzm3fIuXZyO7m/1sHYYF/8si5wYu+qKf0NOuOK
zjE4Ip+CeFTxdB0qL87t71VlFGn8/2GF5shZ1y86poT8SHBcSTi958rF03E7aF5xsV3W4I9s8cSG
Xj3CU5WNyFc8rY3j+e63lA6cGIdfzFkmrQXuOYDJYzJogwuSjtimh7pxTnIJLTzwQQL3GiLvBCBa
QrOX9YcIMsjC0QQAlB/G2jQebtdgfOO2Mba/3hyNZhM78IeY6krTMFZ0rGXNtZqHC0Eo56RFW0bx
heOu2ICUslcNGubgLTYzLyZP5AEGgwi4edMZHWIwzrRvZarHlLOg24k9vz0gjvHkAll4A0QW53oj
Jg0zB9LHGHV4npYurHAd12Sb2XxGOPrCLxOfG1o6o7zMFA5s/MgBY9ZdDpFdop0mHxAuZwkmTQ76
Z2AOsbj/n+ZCf9wl6/aYEztPbLI5joq0SdO/0LMswTJyIQlELY3oBUewigFrTO/vElT/m9czlW2e
6WdvbwIYEygGLSsr//auIxzGvzmJd9rORaeWBhtrbRgA9kHGEUgjQFxQ3cZD94j8JWD5b+hJKZnj
4RVEPLEaA+lAl4uLZHRMU5MtrLgkPliRVODjGVpy0xTNBU5oJkJLwJAoU78Pp35bc4vf5Z92khNB
WIHczP+rGPH8il5QjmiYN+/JyBsP2DAr8fIHkPzJsF68TfSoEe1BrFOu2kni9Xffyvp3tEyW24Zk
Yz5cq1rDuXipXBZRjZW/G5GmhKutEbbBrd1EIjO7XcfrTcxeXculTmX4VRZsqF3IXGDlsHSb4xdN
SvyATQCb9YvuxrJt1apuLbCiYKx52fKpXbxZtRXojvaqeRxMBESP5ao5Xa7Bx7GZLL5K/6DF2C+8
u4dmvUCct5Ckt6C3hO0Ote8p414aM3iFWD0JCKNdWCi31tv2H2MXBi3avgFPDlKa1BCtRLqonDh+
u6d/q+VUx1DyVDRIMK2Dyww9C217x1PeBgIu9dpZNkXwxDUPt9QP/ozTU2RuNpyjjGLzIyb96kk+
ev5uoZwfhg2nxNlLhGH8goS2XY+wr1tzskBq8Qry30hiotQusR+UQmj5TU1JOt3AQz+Gs8I+51Rd
u8yLm3k3hxOqVQoDh3Z5DzgOCWLM7vr/1hCwpBk/sToxxKaYdjPQRptjRpThEsSQBGMbFWu2oWM+
mKBqgRZPPqN3bcqiHEUqnI5Gw/KohhxP3J4/RhlmAFB+qnpNtdw3YWDv8FoM4vQNdXJYUp6KWvdz
F52XCsU27gIbF5N/39R68quXol0xwXiBtSrhGH/JX/MSMC9ThTZeCYebR4ibVI8mY1CHdPfgznD/
D9Wl9yJtDvszsqFjfwZQcEF59jyIqGbiR3HGpEfTcM/6QC7AVoZ/rXC7CJnUodxjOlKy03BBD30Q
n0zspxLkZDzgNxPE6K2rM+/NboIXWkYhtV1d3cXq082u9vmMqQiatEKg/2B3dOKsWrRvZreTWpbl
USXsoRmlIRPNpcaedKxbgBCOtDwW9S6nr9RfilRHmhtNvDmED5GH75W53+8y4EHnfQlY3SeAYQMU
yunkPy42SZvL36zfqIjie7+ljkp+rZrx8ljshnLIfMJZ+dC3801ut3lCRsI11y/OwlcdksBApQ/N
d4YmFn9X0h6ncte+fk101GzWGyM+n4sbsR6ZT8VGr6JdZh3bEswXw+aiKaY8N5ou/37R9xPyMUUU
2S/o8DxsBt3kUcWzHmMmbtJaIuG7KBc9bEd6gEf+F21hSQxUpCuqH+VM6yZYfnfDZhtCfDM91azK
Wrj+P6QMNDOnMx1gykqedjzo2S9mlXSXnluqmcRkpy99dIPvMGG7KvnWjCQgKEdZyffUbiisiiea
bo6u2M5zYfkta8OyAoM/jqEaAN5i/Ud03dnTo0QkqUfX8jJn4Pe5ETH2UKV4o1mNYNaIG+dnrF/8
euJUCBSYEebtTte4inoOgGBjrqEaB5jGVlRGi2prgsW5C+pfzV1/yDQ8Z09nciJLm2Q3Hsr1Onlw
2AETb3cZokzCJiT5q4gDVQasG9gqFaBu9ay8yF3nlYiPwlIv1tUGUHp/GqDTJToImIOljk9jkM2u
yuvY34GHL/TG72GMl1QKpsKiV161fNwJ9S8kvzWVR8swnuu6z8T2D5MjLSXGQQufOxccKg4H8K3A
JzE8ucMRKHAR3UO49MybqMroeP92RY9cqI/kCQfQZBDQqSt1jz96iBJb1amBwajsUhT1Ml6cO79V
vU7iF11Z4/kW2usRczYeFQ22nVcy0APbO6lHe3MqxKYUBuApEaEBzTBc2htSjBaoGRuAWB+GCB3X
ZKYXKhJsrOMlsUU52qRIdh06r0H97kpfgoeP/gsyjOp9wxIA0JSnN0te4NvEI2TCeeK8ESVxjN9C
VFG6vI0I3wajHkXviCa76wdbgDhyiSi8LaqSVbgQmXF0EOI6HlvR3DT29Tm8HpCJ2a8qH5Ki2v8+
7fcYuI9dYH1OQvmp9Bijk0vvxKwUwz/GNY+E6GyYjm5wIBERuqAOHZCGuKCIFoNpUK07lK14SoCe
mrvo50ielEtIrtUHJc3BG3k41A/W7/DIhXSQrEmCaOyxUnT6BDUA0Gy7uZUUUg2LIsBe6Mugoswc
XtSNHSEju1y2jpziqCAwiGWsmXmAht4ZfDndkXNexvxLwTyIYmVmL9RS3aC57e3iOGqqj2NoyAsF
HT7vn1kFRmTGW+QFluTpn53AQwGHswR8+vGeryBp+pczVYExKtwxZYsaegBPj1EgCBbFIZVt0VRR
TCFvECUFBZzEG3I4qUb7gqc+tOcuknGJ1iR1tnf8uwDrye3zGXAVxvzc49NrMDlemdE5U/VsQokZ
WnzHu9fIBRH6B91Z8uEWonIPp7K31Trleb9N2iQaSld2iBRX3iDMj5HOtGNpVB5CeE0Why7GZan8
GPui8s3KqLSjO3+W5R//4sJFZFiGH+ud8cDw9C1pWJlfGqNATPaDZFeI0cZCuAyXG3+3doPu2b5R
JkjHs/NRXU6o4RzdIh1cBtWAdFN2DHPj7U5GR6mmCXzyiKk3P6p7ZTi6OMsMfNJCcxLYJmjdiTKy
8h967XT6sFtBBrMAjjgP2rg2RxHFn7xj1Jc13pPmNflL8NYK1s1rvwyDJPAtK81dPArMsHXZGi3w
qFfGg8DQC8+1wY3meFEjneGMmtGBT5ZgfXcSBo29dayOxANE2KqKlpnv+DhUYgqCEQ969ib1aoHA
HfHLPnmpqWS7xryh413FGvaS4YEozz4GhLFShDhWd9uqx75+/ZfW14Aoo3bQVwDM0HXac8yKBXHK
hxlvYF5h3OLmqdBLmYrbFL+C8tkVYSv5tpM/JhntXOMdKrQ6TYkSqyR80GSXIZqqWyufOEPe99Yf
7MSm+l7scIfILEWgX6inu44l+TOODBh4LBjG2SDqa/7dTwj+mlk3AYTGcwzrBNPZOZro3XXcjHYn
RhrgbM/le+8kwNmO7yD2X8Netn3CW1h1MORICUaowJzS5zdiSrUPRbWsxo3LiqaOE0gqAX8g9TW8
dxypLxSg7ZF3bRar9nnQlWFwW8L4FGuW4u4Jbb73KxgD1pQThsTEmP0pj5N0gBuOA9GQSrnkg9A5
OuTq4KjrpktGps5qeFdB5HK82EqaqyyCgvzfSQNeQerbGreZDJK4huJ3GMssTEh762oARuNKoNFO
Dy+Wmuk7+l+416dbAd1B7Gs2NXKhRQ/TZLpI64lFRNowbryde8mfTXlc3NNyi7hxixcFYcJ6nlLp
sn9fiQaBGlo5ZpAhaWJs3EopzLWgoB3Uam5Uw4zl7fQZcs1CQ/Z9bZr5JrQxmPQAaVrYG+KlyAFs
Fl5mEXajFIEaYdMGEXbJSiMLvcd2lTYcXrPmdMU5t3D+Ssf+3QXI0nOvCrP017WBhm/idyTzteCR
BhpWNO5fmdCI4+yZN84zVj2isMKK0nSHkTceCSqwRoVkKKAxFLT+2Hc0VBeE2M9AcqdYoj+97fX1
Fsga7GY81cuJWUCGYqpDzuvl0/T27SVzoGapDI9ERJsONTKbZ2z9ucCKTUBTVT5crwfezPpUTwXi
0o4uZPZ3eU82IoIcjA98tLOXxLtim3CN1eXi4ORO3nRaE5k/rxjT6LDjhf4Yb/lBjoo9W6iv0JDj
YWmxG4QM5SQBf1wCZObquILxdZoulLLFvUqjbgvVtx31sNy2J7YR5jfQmjB453Se1DlHPr9p5nyZ
sdr98hyjttgbGiO9+6lGpVsCjldbl+r2Zduv/r7LvWYvP2u3VkLyYyixYAeyD0jGA40WPv10SUhU
CLIyTu5C2B5k1bGxlQXvvU8a1gyZrPFHdrubQbkECRbCspRiNiyXJrk6EN4ZagCfIB+YSxH7gt6s
+K858qFOVv4ZLgGfFgWKVxHOCFmOYBBripyoDnAYOGW4sKQdMiTxDvWLznu4FOb/IZv+h0uQ3hmS
Bq7juJiOeihf0VL/lPY/fw38LktLA2ZYe5YVHIwxFXUlCV2w9PIu3BU7qsMxKUJdw0UeeXQlPsuU
tDN4pFWoSzNYgm+1hP2+DOwOUlrkWxYAzDw399i4NfpYBH8GG30nPSwZ8z2bzs6FqicJ6p+1Pc0w
2JCAodWD0M4hc8E1ufTIXgslRY8GXaM0oVFyYR+5+DGw9sFFoCvaI/Yyay+UtnBtYkrkneDnYi8Q
huXYuo17xiNtvyVAXsyxVrHxYdm6mhnP0YzM2Uod0UlcQUPTn54WoKYOl7+r753FdvvYfZjOn397
mcetsV+WQVzHu8+4PH0nv45WCg/Zg2WCLMcyFCgCqVSpQpKmzdNqCcAK9puyXwp2vpE+kjjux1lq
VLncGHoxoKKg6/rA5vwZeuwVzO93wzoEjoxwS6dBfIvp/xRhodTdDrSLMdSqHFqu1aYFsoGFAfNd
aDq71rp34xse7G/XJUKsZdewTIX2oY0IznWYzUoxoHzcGPDvc9cvlTAwRl8caaa+IBBqeGhDg5EE
zgg6CUPJcfr3fp4Vomc9GG2DWN/mkZHHeivMB/nS0KvvvamBub2W7CmJQyhlTYXS0Xfpo6b5OsAL
uoqDBwhJs2AvPtVXqZtuGmXHnZ9PCI8B7vrVudV24/ZqgsvLQUCO+Xo2rPZfMfTD6XOmh+E2z2Oa
QzHx5hf5p0+U4AzIrS45ozgjDMaKULGFuo0jUHKuexTWB1QyLJfIeYmAdOMvWTgvS0Dck284Z4Yc
39HkHitDfUtdqpDT8SKsO0d6HDm4nS69mG77lERIJiVZPdae6YbDxNkrtnHTCDycUANpBIpaRcnP
inQYpc5fjLyolpFdtv4H6fFYavw43N5Zdl0or2eZwskU7+/7+xxXgNVVYEJI2ssGV7oGfbV8Wcib
0Lzj27r68SDDF5bo//UXVtTy5HVAs4+nNJJFttFnJIHzv1IG31UeWovsi1b42FqjlxeWX3Za9kIZ
kGYwGzuGI35kSPPcLSmEoSlhvp06e6haVo4LoQyxrH5bJgD9rMMWeD/5UGsMQuBJkvELzFj4xk3a
NvKIZ6vhhqCWZpar+/rkswwJLESE4xYt5gaYWCTfJutAfYp2g/uM0oqlEAhYRB6Gur9cRIf9Pcb2
lr2F1V4GUv2PH+7w4CAKth0omKbXgkst90wbYds2ro+Y+RAgTwuylE7HF1A1qPtqZyzjk3/SNAec
5XntTRq3/H6o9O8xy8uUMPDXpgYMglk0VsKbcnnBjaXrph6xBzPGHz7EPsk/pCVbatzH7jB5UCrX
dXqrZAfbXUkHAtj2KcpF8VKvXgzFVqEAfZoR97JA2Nb2Bg3mAMtpJcTh0bZVssF9YXHrCDlcv+s5
n0APgEciISP9fDyUQsmVsDj2lnINpNBKN6CKerCUERxZO7g9cnxLvn37/2IiZLrE8Hmfd6oq0hdV
fNzLb5sijgI9Tkur9ifubQI+BeCja7V9u429B5dOXellkURpjrDUWqBbD5SxBXQzuoqWecwAJbdC
O4BMFbBZKMt3KYQA3uAahaX4vfk36EJ9aax8NPtT4fh3WsEpjOE/x+dXgHhKWZCUhdaJtswsaVXj
6pFZAyo0ZWlb9JE+1debnsH7lBafG4C01v0aL6d97+eyFPiqWvlPGrNAnHyVujU+oEjZ76MhBgWO
l9fzfIs2PLKez4RhlKRpdfEf1Nl9a7XjS8TSrxbN6+GFglpOwgK8Bx6th8Vtbr/eygev1JPAzYo1
t/c24bIorolCrEvjQU0EZOeRX9puixUVN/78i6CLKNLMvyA0NlrXt784SRga0SH4ATbC9XaiMf/Q
yyWd0xGLpnzM9H3pZWgfdW84DRYBKdyaFHb4p9LKdi2rIgJUiPd+GEm1gP/Q4deha/4QXHZpCVBd
Fl6eMNsinsGKp0MRRr9FdiDXD4kOU9yLWPXQT583dxARASFV8rNFLztqgc5qxtJF3csFNYikTXJN
I1L1y1GiFrBL49rgiN9/rrXeqJmMKW5ccoRmIfIIMOzFCR81PYmwGrnIIef57t6eDKGa2zfI6g4b
E+PpsQIPCHQIn4SDKJ4ek6IVZGUYYSojvKUjYA3T2rYle5TSuTSKSvR57Y2XR/EQ+l0+cJpntPUI
cigbw9plbUFCQQJEvm5cU0apE41Vx7+9D3+kSBy6Pn+n4fFKQB96y/icxzIWnUF75yb3Lk/NU68I
S/PNs+GAjnh4eOIJ16ZgJDS7Xp/v6GnOiO3+AFtEcDEWfOw/KBDI1ZYufkI7NVUwSLPnAzhtzI/U
GkgXbleVp3hykwqa6HMXA5Deh+RWwWMq6H2oYGnbgWIyae1tYAd7acJPjIiX9zbTMNh+jP1pZSCU
OUo4QeuTS0AjFwcFKSse+KB03lYBOTRh0l+84cgqamAwCOhktR2KKTh5k5fxwtgTtXuTXgycDY/d
qAKcqMXHVhgSShMzjyvEYJUmzqD1V8OLMjOWfFUsbc8gpp5s6FR29EpyXnasuqySP5G1fCm1rcHb
ziK4v2PWnq1X+g0fTAdMyXLtFKLxaKx6HpL2W6jXz6qbpjWAV8de07oBPbExXlShNR8RdOkvtKfS
InLxMXETXwtw8PD3EDzAPbKUzBdFc6/FGUqW8+tLMjv9nPPoiBk6O9ApZJtj1dF5L/JlgzlUMmaY
15Zs57hYFyhJLhuoQ/jfas7EJTtFcsCZmbvJxh/xC8vmmvvyS38bYI6v82AJcSL7OpRlAWkrjqjq
vizgxb5OOsSX/nucMV/KjHYbsZh3E573s8RGcuPBkm1JszeET2o0r6ld1SV9Im+2W1sdo+gSGUoM
qo73854vxYyCXhfGvSywXwaa1TNkr7pmLsFa5/2MZle//egp3sjFjnbDdX+FzKEcr8AcVXKy/er9
mFyA26VpeOBzKQWyc+YfuMzMrasUWKL10e8JRsHFu5eMZ6gbONN3ajbEOCAfNwfs2TP/5dt12tJD
XFHfmORmwBr4BpGnbdyahJxfU2FoW318WC+n0RBdK6sA3rgOobVI6ta9XSGIYpWosr2D1e7NuPoL
pzzTevxbCVIrjyifDJxeknCyqOW0FsvD8XD3S8H4xUV7HhTIIw8kxr+0YJIC6HzFWEEh9FbfQbIZ
tjDPkhLd92vigUF3B21rX+6wIMmWZoZNie3TguDjgMdY2Awx9LSt0tTuNyO6kvmM9G1L2R6QtcxA
TEtVeEhw4BTFUswklnDq9Z3UmbaP7u3zx553VSHfiFyyeCFIaXq+rduzBd35webu1E3GG/jKzgZ9
HPReH749an475dRYduMf12Z6C8DGTvnHBMQe3hbydysE9S31nLIui7whvHclBlzkc+6BQ4vnIGnw
uRLSd9bPYT++b+afUlSSNtPXU622iSJZh4IsVWlDJ5bZ7yKXPc6vkENo0GSulZc5XN06DH8YF+hU
7VQ+pdSAU0PrQ585M/o8LzaBd23csIUimJj7QPAoNqP2AMX7bWPZFMjqOmsq8Y6K1dJqG1tXLF22
YwkqUOOcqes3jyiwMibmlNtnI3C6/km5D3qYw7BQ2j2js85pe8txlO35/T0jxguED2bQnfaovv+R
sGZY0z5dyo5p4KcslHiSuqTeXcaQpR4DqnaB2lI7slXM8uyrrz1aDB8IXEiyiHxn2RgcdE3yK5bo
mDu+ePnqwy5ouaLjywaHCLQqRLHPlfes250VPOGsAS1AiBEyNHbXNYqZUPvnPjwHbzfb84+D5/eR
BLs+YZAWoz0udFB9CwCcHmdnlVwr2L1hEK/XsiRXoYpzYyO8d0tHVx7y2AbFsUZFk3xIK8ek0hM5
SjKnGuhvRox84jAYDCuszhicYPawraITl8XbwxSjmMxOvnZZgpCkWwe14Z94eoBNxl4xj0X5iYIA
diZ8KU4TZ30yWZ5euxup3pkuSTPS+J4sqggag0uIAbwFUubjyINpHQ14tiFu0S1sP294SdMLkESV
IOY2IyV6y5t4UBpomLvTtTxh1Zm8NGYG9yjkp3aMVI5NR6LVEtSixbA4VNhxDBMyqnQvyPnQ8Rrg
N2dIXzZKlOLnc3QGksNWD90/xg58Um6DgMbqT+ZzLy2Tmlxx7RP3o/O4hMS8+BNsdnHFG3gYbXd/
/fYuYC+TS4NfP08QMT/9K0loRH1nX9cghUpEjYsMA7lynweP4eGL2pjAF45TOWzMuUdyoGEotavu
QLfTPsCkTe9v9mcON5q0M03OY4a3i4InewG8P73Wtsi5F76yow+BGYpbaR/AkeIVumPy0Y8IG9tK
8VWz+Fxs0h436wmOlV6lVA0oaYxuWyJmlSpyGK02zhUL7wbkvsZN+vR1nlVgPTOnomGUFkgFewaT
+o/rgfBz0cOlyvoqAItWTFFqpB8++Wf+p9yMcaZoMQjRdLR+208x+gjkufrgwubjxF+VlsB5AyCx
sPWig6f6D1tlMctO2h48woITZyfaV1veBZRFSpKVY37CPliQHOYmk/NZJ1ElizHgrX5D73cbG+jc
vao8nwna9B7PbCacWe1+Btrq+xKXoqFrZvxWMqQbMlc5VsV/DC0K+kzcdt0D5LstB/95x9pFjqbA
s7qHdA8aHDhfukLHLKlLgzMd03EBZeDQYLsR+N0wW8iFnDyhT2f8JVJuB+3N7ZR78YaIHAm1L0UY
PXuMFV5QB1+BS+JHfBOQeKdJyeeXiO91UjwFjZIjELJ8Vus2+nCHVb2pI9JNNihG2QiNFkeoiFVT
825WIP715TrxwsyhkSgW2RsM0nYtWBptoUvmFMyRHdBWeBeKHnVoQsMxpxR7nscmKwaZvu7MhjBV
CO343nbRsfa83e6/8YEB16arS8iMXOm/ka/nLztO7WH7TlK8oq0zzMN1hf6ZFXijYX95lb38bqiG
7NYNhywv9mAN+2ds/WpaVDGE3MP+q2GYlAAMXoqFlkJAAf62ujDyydFv1/zlGxYS1aIxcEskUmLP
o8HcywCyqXs6x1rWYFPYG/UsKtHBcOOSp3GEGR3qcribN3ICL8oPwNuHG0MCGVZXD68IsdljP/C1
4Av9vqbHmYoJONCOLwNdsAxnGzmmVJAfYoWyvqTMW+UQf2rzuxzLpPY7CITe9n4POGOF8F6Y+6UJ
GROLttfntwk9KpyyMAPpe5VINXMafO2zgUo4wQCMMuOgvjQqUXvDvKXUGoVwv6znQ5swaIsugTNr
3XIBrxVhe9/mZj0QRDtrb/1bcbCgl4hRdVXQgZ2OKhzrjDBy9/iU0Nbo2JGhQTuYnPVn9z6RUa2P
YsYjyTi3mJoHzXANNZm+QYLedqpApXopYzJHrwU+ZjeGfyUwcohsSX/dwYs6l+oLTlOKZ1ymjvzp
LZsETD2JmV60pFVXFWqYcugWXHBJJrCHkLd4MBsY8oxxPnGI/YPD2JPoo6ieEMsrhQi1+u9Z+jHJ
z2KaqPYykhUHBuDVLn0MY9ioyhJlr7fbNdRmGAHg3EYQkmF4ROrCXRvRUxy2eUl7SoAI3WtP/ntB
OrSfdnuG3+5IArqkVOkMsu1ItTs3lUtK0GGZwLmqIJQ7uvqHeiO3ajRjEnjHQ1dNKz6u1TGlpVZA
lL1MgBz/FpWjCCVZJwBzoKKjo6rDxnWXwkajRpfI8g611DR7XY5kALnAC6eFQ9yPyPaHNt+tQsPc
U8DSZISuGp9XbsNuhd1qMVaIQXVDnWsTaDHAO0Phej2Kp+EkHN0ecMsf7TppNwNn5P5mLTuttm7T
VNtxFHrkOSyVRzQlXt7aSv9TG6sHMSjHIDER58Emz+kLcWwZalJhhOmgvgnd57syMx6Am9Z5vbMs
w4WG4TNNd1wL3g+N5niu8mkfWsC1eUkqXvzBqEqZQnvsMMyDXFK+EmcERIlFAW2k7bcn8GVsbk1F
fPpqt4GFqYGCWgkHKI4YZMO64f08aF3L963YrK+Fhp+qriY3ltsdqUlltLgz/2oKOt52RtJdLUid
hMJ/buTXQUwt/4HAAv33Lc/ldz3KOlherG9ocpd5e8Xvs21TpDupBmFCAyXal/QmFN/WqWgGZD0P
uqqmmwZVPGxMs+8tzgVueLdZywxVaz03sMei4+IrLtPoH+vBAAZrHRsJMpx03H81fyzC3ZblYUEI
yGyZev/JFIJ6LIU55MLA9N1rsBZK4araU/PB+wWaFlgYBWG8Fmy1YSZzBcgrrZ3/5gCidBazitCB
nbF6FzWzn3fa/L0cwHDXGGlbUEiWz4T564m/7eFggq+D22ZcPyYpClaWnLh/L9ovEtMkCMWuB84a
NZ7Spj99qM4bnD3cCzKbl/XOxv7KAaHbEh8KmuRyV3CukZiYO8zOkJy4iwG3pou1zI8zL/+xpLNu
LyId90oGjZoGSExNeJGn2E5mL0XsFj4U/DBmupYaVFg8FoNBCOie8qAgVYbxzWxWoyiaVjySvI8S
LNUjxRvnYE+Hl/+gXfKe6ogSCREpLwsI6VWrd/kmkbjeUUYzaQUM3Yo+2qiX8bzMSySAu1egNrK4
iTTpd8jq324A+1f9xtZAP01NV2Hljv51yg0V55lMRWn+FSjCSbEX1W6eXyyqLOnBoIveKSnyUSbC
vksSWoKzHXYPdQVJmb5yYfzXJTXU8BZykuzabvzKXWl6LWHWrgU/9xdSkKMsLrERciz1rLPnBGIQ
kHP9GNxu5Ji+9AP4HxITWcgAOuEPM0Lq3aRschj2sTVPaYuMc/EZEpN/Q7ktC7bGQy5qgw2pRs0f
LQh5kUX0u957gkoXmLDwovTgbX9bAY/Ikqzpd++BqfaEkg2A2z7xMt5iGrRH8Ril9ZTfhqjxv9fc
Rr9hnN/xNeZ/t6PmArRkvrWuvJKaEomZ8tR3aa5hd/jTLiC8axvDJ3NVCy4a3G/YAaCpWijhtXHM
vlwwe2zBpmP76NSTI6keRfSa9DtF5b/Smmpow5FsbPAOWFWuQI3k5A6D3GoDPwQ+dak3rDzjw1Z+
2z5OISrH21rg6uL0mrTK69oTuzicmHoPOMN4RRLN1VtCkigbqURWaYsn1WIvvcm0r+nTlnMJqUlL
/R5rvXqwJO6zmvf9KpN2v9EpRvJo8PRyUe+1i6D3JNu6hvXQAeq3bb+aj+rYN6X2bvO4m8Zy7ePL
rjWRxgSF8ldzoqqmuDuzfd0HNtlJIS4PkN5+QlcEzC4lP17PdB9VcI4RIAGXMPWtH7L3G9i8qL9n
lApgl1Y+gzL2OoQZljVTc3wG6yqKAc2sO8VFoU7LasYYI+1wQBdubFomSwhzYOOI9gZ5BDNNUDEI
alf5rpiISdBteEy6jOIaLW4H4G4rMqwaWgXetAuSNaupkWmqgnrAH+4LInAepTsWfCfdImmHKUU6
zScE/tYJ9SIasWIvVXbvYh57fcPCdjtaXo3GNKq0R/42wSWMlAk5BQM7t66rWZmJzsSsBhoYZJoQ
x5n+ZSUvCIokNMUlbRLXlK6eDVzPcu5TD/W4ufsQrM2NMAJcOvSTfBrBaUKSUsJfc9aBhSOI8K4j
vDjv5zDlBVggwaOoGHye4S/gWkAmR/CY0nOUWoWAOBWK/rtSneW6Wes6hugnfQKE6rqhvFb0WZJh
g2XU2oVCkjkjhA0IyirR81MAyv4m3XzMEdda+uU9mMkwfmCMeg6y4zD9HIs2vnJetSbv7+vAddFI
DQrlX4yA2G2AJr3/zD9hVdxuDYpqtlK/AC6FF8Q0ry4pXUpCBpqYUnEsv+Z3Uw0wJNVmboJAdFx9
rTzHIm6GKy6MwW3/JK04+ZCwy+aAeJ1SxorQHpXejxxvJk3i6P6RaphYU+5dHWTef50pCMcuS6b6
g9IL0IkuDnYfMfJ7nchW12XoD9h+8lgsExb0WGDPldSlqfBQ3jCqbc3EJ8+qyTZp2DT3IDdvqLf/
ClZ4dHqq/+Z2HGQ7CcpsEgRtZtILi5baESe0DzYdsX1XrTuLS90fGovUjGzJAJX54Pt0MD3oKdiz
kufad1BUGoXlyTMp8WsbRPDeLvuhflxLvoSU8I/bFmvJpea7P0lYFBPYr6bWu25ZzWff2QCwTynn
LLw+DT82yooHUmrCVh41/fOcdUqMKou6LvVKrEpGUbD7twrOMrsDqldqcEaQ24WS/MGDNOwusdIs
uaMKkc8DIaX7Fo/uFRxQctIUweOztcDqXWrdRdOVdLhSlGgAPR4gzICUX/KCE5YwJeJQrAUUdnQq
wQDJxzQ9IAxePhZugWOyPhTIuFjkY3ZOsVNljSvHggpVZEQ9FR4+z4Fp+oKseOsQ3F7Yj0w8V5jB
k4h1e3Hb7U7E8FuuIJpgYX2SiTpmtLplxJXLL/jTbcvGhISacjXaNx6q1PSzPvJ2rqYl9Ni5kukx
a8/y+OOwDRc0kgS4dSQKSEac6hCPQE1yjQ8mFf59v5NtW5aI0XXYJF4NiSDbCnTUd6UgLzuDD51z
ol2XXgdJun1ePp4mKf6vfjHyk+QGMzugFV87h0gZwvKO6YyhKokqSmXX/kh2tZaZF+EhLPJ+BG1E
msZkFEeuiit5U7WFGG2b22KskwsgQ0O7mVi/6ymuXpc3JOGIHrK2dJlsPi76GYYON7lfqga3uclB
LhnfXs6a5LC8RZoYnWFhOeEueJsepaf+SjjkZg9OZc7dH3DTIst8qMlmW8VyOgfBhbZL9cYtEK/+
VbOYXzQayOIGkd5j5aVTH99CSKoE6xCh3DzIKPhtBeRBmI/MD4sRPhdjA9CGPANpiYwjPeRYLehL
0JNrIcYUY24Ruj08g8qmfP1lKABKiMP0f7NVW7cPTAt7fLyIyL/6RLNxoWIXiWStoC+FGkP/ZDxU
lHVf9E/gKOG5lMDOnTkpVox7I0S0kXK2k+qsPIq82rx+SVYjbh+yUQ+jREHKdoq8OFL21Gvy+xMF
ayNJJXEfCOmwLFDGljULRzznT8YaqdQAm5UShswK+VANkf3+U7UKpFfgLCfcytJRAlB1hzqT6lZo
YsGiJE9mSpXad7OoHnJQUgFIvuAtRM/NRzRTl9xdi64mAzpgMLIHQJYdTYZlK9Dr8WJkyjYCc+3d
SENKUPHH09/3kjbKgj7yFxQfb/s3d999EPJD0FlYZTS7trCPbdUhbwPXZgpq3jmCJT++JOvvjHhv
1ix+5LZ4Po9XsIW8N+KmP3+zz4TlCSWXpeII9cbAEM4km/whXZet0aYquad80ajyqgz+YZiUbZLG
KnTixGFkATJnavdnGn7zmDxRXspcoiHEZSuBAcIKbEcv6LdAFJ4TdjlkFpUyjtfuiVMoTeR44rwU
T3TQdAsV/FCMnjiCl1aCLUVywWzjv2cbZXFvNCiLxwxl8kuxabaGeqMI0A/qBmNyn5/MJt4z8zBp
te+fu9JTfm/I0BDpRA6lSvVHGnuoXnJXlpFnXQYKnpBPC/Ea5IkQzaZct9OSRnRtVMFAZY2OBkwo
pCJiOL6R3Ub+wPfluePkdwVa/XxR9we34rPqjOwz3G/wq0ktJxfRsx3QvQCIURKG29e8B5/arenI
p61lgJSwa8ayDEfFYkP9K4D2jmj9Vft4pcHxjjpdfsmMVkDwMHwnE9HMOjX3XqOIjj5GiSNGpfZi
Uaj+6rJqGrw3IInZheYl8T8boVFgSbdmMCt2Jf4kxBhPFgHlX0DwwCz+6l8kfSS7JSCvHOEv8hK9
NDkpBbSYZuL104VG0LtBCtXJrgR/kAqkQ4GAwqyBBqHesjm/eiBFpD/MKGbeYs25/FOQ2/0Mfj+Z
nqedpW73ehmx58XJsk7kWkN7xBBsNCdPZ2vLKJcUnGHnmjzkSpbzgb5SD+TTS6d2s+GMHgjRdubi
OmjOPRwTHN2FB0NmSDrFXgQLVKJmF29SXT6tHkK6Io2/+AKd6/bCzZA5R++CTO/L/EATK0NktlVJ
16eGXrQ5xB++3KsD44GogItgH0+oAwKY6c7Qyx+fYvqJgKBjNWP/PMRjfLokXnpf46xqnYDe0MyN
7xiWO8u9LYKX/Z2kUfn9alR+eA8kviMj0KWRg0hCES7kkDISuScr6eGm799r/9Emm6mgAXUaiXDw
hOh4DhelGoRRTd5AhjAumDT78MJbm5MCbrUNDcl+NsLoIrxNMHUvpOh0pvIFC7NEAi6DElLu5xLc
2XbqXfVZJV1t5+pbmHpLD95k+HgDsLGfUdkekqAcajv7QA8BT7oiIaj1Pdwoe/Xp3z4+2jUkDPnb
UYtEoJ1tHKEQX8qh5EedVtB1Do4mkJKVISQ8B1DZ62SQXJq+djtKteWsVUw2TvHsKlZp4vL/r+hf
pIwOi8SSxX4LYe0UGrupq4c+XjNaxz8dOmbCcAmf+WrICyEoAzNrQ9f3rAZqiJOUrMdO14Tz41Ei
iwjEzE4Za6cA/XywwbDCGInRi8EgPfSh0Ya1WKo8eoyKO50dnQIFXfOAl3I6gB9rhYoyAg0KAwZA
UL4aI4o2vpLSdO5kspWKVAT1DpQY+725K3c+w9253ny+vwGe1/H4odbjj2oAlND5IpK5FZO7A+z0
U+/aGtH1QSAumOvY8TP+XcZcemdZBsozLcshlcwtOrWtnUszc/IK0CGnY6KwdnVQzamiVgI5u3BX
92xVRjTcYw+bp6rz2NKRnDHoUfgFMYCFyw0pdpNI/7waQnXsmvrWRVrQjQrO9c5tA0O5OYPsQqf5
TxD43QV1cX0efvJo4maOISh8gSgTQRrDWGTfmjnpcMZqVsukgqIXyG+3TGDUSVwNIftR4boxZ49F
jWwl9OGzzeX8MxgL4Sg8FpFnrt58kr8AEW5zBVOU+1mkwM5SUDEH74t+Ub5Wv9eL8dUwrgbECgrR
ftxSSZ9EaE1iapA8OEvctV1oMfl7aIlyPorHW91jBvjd7kCFIShnJ70WK+f+fW8i/ryLIPEQ2Jxv
GR2bg+Of2Ri1V29K+zVv/yHwgX8xq2nRRKKi55MPnda27v1TFm+vnfRgyQexk/i9vMklf9128fYV
fh2l5l2euS5rrooWqqj1qC0fLFSfXn5xDjCN3W0BAtrLnB1AYg+jTjb1jrNaHYgDsCsh2rZ2QiZK
7csS4YAJUg+k9r1c2RMgEXApKYRL5cZdevkoAGaxlHfYXIQAedij398DYTE69kAsV6q1XEPOwVZ+
5I/ijRYbr2mdYK1+G2/6OtcjZCCjzHWdE9FiGVJtlbpEKd5PBlnTVenKJWPxZqIwOV+9uIdRBw12
n6NLBb9+2Wxon9DY6sYL+2lqQk0qlrklXf6MjPYoUpWt5jHw6naKV7WFNkdXLdrWVygwpSuuasJb
9oIFtUSjzQwqdYZ2r4/0p9WLm/FUNHBejI+mDCa7QwKjUvzTZr/7uhLVaLuOPQUJNY8turK7vNs8
UZ5C6lnDQGmrxygxbz5XmLaaDMtl1rsx+cMTEKkOowkqhlDQIbI7BYS955fBURAQQ4N0Z+0lM1Kj
+jy905DtWVuGX75G7/b8i8pU0EBpmS2owoGmgPJmDjioOO1JWL4/+z7+liHKoDtna99pDnc4SaBx
1r6qFgDFUea3QU7Rw3iADoeZonuANemehv2Xyt2rpogB8d+YmsfD4LNDD3KsYgIKZ1408e/+hpGV
JvHDnC0LXg35dFdEERP8Kzws1HMuyrQCqCdg31KGLfcjQyjO4PfKY27Opyh+LE4efSiABuQdYPQn
GzEQndUq1DPlu14o2mcGvKWetYHJnJDZpgVjHErgBq3upJ1XGLsn5+cKIkSV1T6ZZ7MGTTVydBa1
7wNiEYg+pA+18XYo7WWBIn5T4qFBPGArP+XS2yx3isZbAAxZYWVpkggxAoLqdxiCItvaXFpqdExD
iMlLHZAQ3eEvSOMrtnKfy2+fevD2R7X2QDDN8c/ndmXWgdXDtfsWyV2brSbMQJYjJRX7DoALrElF
AhLDs2tDPaa5J1WoiQyPlk7nHlOe01QsdGFTGeAegqAtvlSSUZk4pDOdR4orb4JYvuhRHT7krjOx
9Ebrp0iZR88WrzuQ56KHQSTEBjolPiN9Q829S+qOhlNWxi1ODsH58PFzhzs8FhktBtDlGr75BLAF
5ArSXlrFHEkPJrbc9FduTDUNzB/68CqVXaXeh53Qf8tRqF/S0UHcXjcI7pxbDc/eoHLsMyC6SWah
PusuSyn2cD2jVSK2tFv6G8gi/UfCt7N2fXO9MaWrWu6BFWzSfpQ+eSbUVQUCNQ4qOjkX5rVuQGyP
ndeIQtjr1l/LhHUrTZMbXnUe2j0W+bxoZI3HN6cFpCkkEoVjYQuSs0e4StSWUlj7pMo6PCF6lKAU
d4gGNt4aaQIlqCD537k7okqgGP+1iLMgrpO/gMu+2lcJnIpj9BbFYlm+M0iCU+7rgXhk2xuu+ov0
yrQqnYN2AVNbAEScKIKaWc87ayONFIxg2UJ6jp1io024dBvUYnBV6O6NoQNK8lMsrB44zifk0G3c
2MgsxVfHsCziVP/yKSLwBOXGuk5PAyRbnL7nasc5IY9sR/6tDEbfX5QLFGu8sJXU9R7ZQUXtwUFQ
f7doTOQYSA33A93OkGjVNnbcrbzvjTyPzULbuER0cMSPDNbm5jYnWKrhyVi/8C39FHttWsIEFv+K
uASGHMo9R3qD3611YLKSj0Oqqhdw8DMMNM/FT+wrBi0yfqTjjI8LCDoYUZCOuPPVyi1HvPrvgZEI
0AM7C6y/4I2JHYNrnAWUnsAfWSSXAXtaEI9KektE7qoL4OqXFm7bu1wLDWD54/+ZITnMkXKUXMU4
xum3fYOQuzqC7YoUrc3w0mRLuHNzVEfFMU7ymhJBURYpBSXEmMBcK/HV6KOFfSheRYwXb0p1Ouyw
GBB0SmLmeRfaMlyhD6l5XT5uqXVtkxIx/zzHADiFLoLGT91YsohJYPFgP/UDPdxeoWkdVihdfH3Q
J5gUgRL5sV9ZMqB8EuGBUzfNX0YHyRjZxdMLp9WJZuyLanoPYiKoeHFWKVxwx8HHIvF/PqBsQw4y
zOCUA7OmVAz/QSwnU2KhOZVGa+cNE+rnZ0k9UldOddn1yFfaESsxJ+iCJ6n0+wFhgQikrBdt8wwa
y3Aa842p/6pZ7RyuH6R9Cv1qxEZkbtBQUHUXcXICMWi3nBNFVq8bki8MOsjki6S1UA06c6Xzff7C
c/DmkeDtZIwoOoj3az0qvBwymbv9tpuvYOg/DItmELRP27R54Nx4xLw7/ZDX/VrIeZpz0hEB9hgR
h4fApFV6Xkde8BnnNC0R6L4hhaSPCc7vNRS78+rcOfkaU9wtDNGSCx4bC7hsTnpQL04CGtxFGu24
hAik6OIpYX8XIrz6AOkeWo7PoM5S50QlLFXzWd9g0PVTX5SX6b8leRYyrr2Go97TIkOMtssyFt2E
qJ/HSYJ7N5STKAwMe1iqmbGU54ZHx66xjt/p5+kwSKs760F6fbtk2G3VsyvDQYMT41ks9cYDvHon
bMTPohZTqLkkcgqxIYFklvbehIVstbk32duiZs+XRl9fyK0B7fivFz9ssyDkvux/V4QVWNGnwDU3
AcjqWtq7R9ycTOvNcgW+gjWv49QAcocp6DsmTNGSYT2sa/wxqX+s2demKT3ao2NYOtBNzbGCclJb
l1PSNdTGshDOpnQkD1gSBO/68Nza7xHzx2V+pAu/ZUxtQiwIZDUIDBBvGGpgsAd+BCZzKnG4prsU
LLZrbjL3xAse2HeJW3A4rk50hQbxk9ZWrGbH3gfFobJ3Vb+gr0ln9hL+FAhW41d4x8N7cbzuVbmF
O81GmP4GPNOe5VamwsWh3DIctTjtJS4Au5mszKQ1jTPsy6wxaNbZylBNziofO9PERk1u4WuTtyYL
Ody8KYiq11bHEZZm6JL4UBxejCgmm5/6ZBEsl62eN6ktj4hYuA8QoKcsW3n+zjxmPLCZFyHb8spV
9fbh5dh46zt+6qam2bolUNHOPRBx97nWwiDnl9kG8T8cmzUH3IyZpButF8rDSJ+GpVAuY3UE5W6+
pI8QP91m/VSOAte4wZyglYSQL86cCaRn2zqOq/56bjqgWNu1GSILk3A/f4ak1jIBxf/EEF3aNz85
Q7z8PLK/5mwrNMN9cuk/55e11aEQ5ViYnG5gSCBTo0SOChLM973AshYFxVWAoRkprM8ELWO4/07J
oAwEDDUOv5cZ8+xNhf9NpiWyXMiRHxY+9mr1Qm4F/hqzHNJR3tkcYP0gV3yyidAdT+dLeCDDHtck
lZnGknK+/6g3BvDFjAs+secDbGrV4OqBwwdc+EXrMyhUeS0W+gelsK8u9wHrby1LUTpOWg5jU0by
/WGhRnLZIF2K4BQuDubvkVHOJstd9FjhA1HFzZoD7AZz6CtCsRHg4/Rz3e5C+lZ9uap/7tAQwRQ5
MP+xNvIorp0Zrd3tNd8rAEIvYvCf4Ztldlu+LqjrJPxVjASxcIXH86ftXfskLBRW/X5xgMPbPeG5
GAS3rHU1rxOWGYqp1piSaTtEUGckgLxLfrMAE3STK2NtPoS55xLrv7SO75DLNISZMkFbanF1Bl61
ZqO4/DUb7nspcxbNhS1ikbpxXA1GBrJkAjHfDVilMgjyiVTaqojBXiBVPRIKvtUiPDbD8iZSK7Ey
4sbaS1IBxaT/EQ38+1vCd17B0iopd7YckqNTwD8aqT4rJ5baFgUy5XA4nu7YCS1uqOgjkYsCcugG
5sylYEWjykGRaCH5888oLAakiY2oP62Dfz49/A5BeEQYeQYEMuPX2+IAPLN9RntnGbSBkfWtkGXf
zeVZ16CbkWBiWBf+CZWjZTQ4mWSc6pHxUPb06mvgyOFHQxykqMrI2oyQK2BGSHZ3yH7uZ3WUqjbV
gnDYPw1LmvMhygcI/PZ1kQ+RXsrj8DY9Iwj392Lyq6FnUQR8f8qTkvN+eCQm2wth8nteVR90fp9o
LLgBhITmksQCJpfGfQ7cy7S7XQyf23p7PSwxzOoV+XC1HDtXPw6mOnnfE8Iqf04qcJSZ+fK01jeF
MjTW4VXj0YjRQ/11AS6FxnUcoZLmILKzX3LWUqXQVH3evHlUiNrQ7Tk/FhTpe/r4jf4fLNns1ds+
iRDG90kqXIxM9w7/x8SR/Wph0TWWjyEEEqP2uVw9MvU8ehqktPmQPA1DUqMK/jbgJ0RK6extRGIh
3zQbstrjOTfB3JP/fxRXGiHsWWm6MO+ap5mkG+syv8GxMNN+IYz7UmGGfPDIipNCiF8s0FGR2X9p
pnL8axlgDTFKLoJvQFQktecU8bvLq9Zm8WgWyjM4YbzoR0czYDnnJLEzwvxU6fOYBoHloS0P3n6L
A8xTRCKBgOTC54DYkWQcnXiseN+ZsKM1PaJsQQfsZKrBOvkpH+uvSoXUqfsXA+b2I3FYRNpYuHKb
Em2vWEEGKpSWgc6wE4JqyWyMXc/lREA2x6mdLn/8UPNbd2/5KSbX1Fs9+gOAovjRmzj1X3oohz3h
9wm6/OzDnmM0OfjHcIBr11c/ubOvv17chZlR+5I8aMCU+uCQefNp8XHEbdW8WIRzYCsC5uz6Dtai
hlxAxHmoyndbUxC9a3U1ubsBv6i9ql7Cov+abquQvqH5CtVpH5hB1RRLaIr/ocmxL+qFP75kJo43
rKuf7CvCAPaH7dPxDnruSnlh5QZ6fOEEYNh8B84/5i++ECSs2Va6i5VbfXCJYZAKHKeq7G6yjdyd
Np3nQyizowbHn/3KcOca3kEe8PJg8oBi/GQRD674fVynlDGQ/5jur7pYpO05XmnUOR7kaeNSN5Jf
f2sl2isBgP6cMvIkeo6W2bsRYZv8rdh8cPn7QvRTo1zisU6HTr/c95FWij/QRQRIdz611IfEhgIE
SqnxvO0CD/53uF1gn5wlE8stPig4Q6oqLjXmYVmtP9Gc01S/XxAvjQNI7i9YehaRQ6jMBs7NK34p
Bx96opm9lHHUXTNQ5aBpyEaDsgs9rpFyYv88lTYnll/9RPM6GrkaDAsMolP5gullF6jOUX6xoV1R
tkdIIGmFC5i6NIcKYF3TMAeowTgpQGOY45XCSPI7rzKhyRCb+jlTVXcuq/7xD1wEuSZEUK8zwixs
TsoX75f+OH5M31vkevNX+5QITN9FlylMAGNf7ah36FJEgFZVHAnPChvmeEBkrKJpLmXcG5EWVXyd
fZrz8E6wwrs8h/bNb9Wfrhq6gHpjeuFk2bOHNOV+2LLVN9tdqILXEE7QZ9DuAUQGAFobtHMan/Jv
pM20LrnNvWDt47ZO9WSjbQNRkmjktCK765ErgCE39p1Ss6X8e71rILZqlMr9RaYCdukd86q9UJYI
cRVxLRJ4ID1FgSKBbCG02/7EW57xcBhd3e3ezFbY7983XLxcPE5Od6e2w2kFxYc54CgYHIgZB5nx
I0b7UIWaY16cPPlzEspNTVFNp90WzHjjWuufwFf31ZGjaSaLRa2beXsQM3lLJleJKVUWvGALnBM7
SxVrAyCGeSKB2JL/58f1yOzpZt1yrZTZGlfBKM6axhlwoaiBsTVYfODNE+CrtYQo6UclPSE7Gd44
sRK/HXeVVG+yavETYtqpR7M7i08ZpUYn5Egh3bNhhyfSKCM7dSzXJ7CP8g8Kh7HTMTVhnmCSAWkW
bYa4sVJztsvLrGos+n2HJkmDq4lHPMPeoVZKpccR/BOAY/YYjT/6JiDFNReFHms8aGTjJECTDJHG
1bqDnekLPiWKY+k2+rY6rqyB+fzYhCo0q7Z8wVje9nRY744Jr7Vkx6n8Gjmoe+YvhW5BYNslxy7f
9cYeK6hvSPaKRtz2C4N9H7kFOEY8kgK85aZbF8SgKUShw2mixPPPAs8Z9egMBFRdZeSyBEb/FFi5
g8BD1fZRvcVG/YK7syoFdNpFSPNC7S6KTrozM1jia2DPPAoPE4NPcOegkLbNLUWBgDX3UVKUeRRJ
2FAq9RvZvQeiYoKBhkWWLrOIY+lXSkscOCeaUcASeEWpVIwyvxyFAXkIEX6oiDk/Y6a2/LXIlwH3
5wVS4GuQiOlQ9bAMtlpGAaA9fqVwpwRJN4NKLpt59/TAUDV+JWdnN2VJnjQ/J6rDdP1L78+FSApZ
Ki7Ig7/LEzjisoN4rFb7RzvRin1iGHj8+5s6C/LTuU25nuKTZBizcD7wc1CTH8M6/b6diFqC+2yy
TOquGMyXOHOCjR8ogTrXG1h0MRHbZNIzwF1DYmk7sdGmkqQhk/butm778mhiHn9HML1RjU2olQGk
Hw46FWA18m+xKLJRR3mjHmzuTZZftHuW0URaOh5mIRLSDQmJoC1H3P8VYqt3Yv+vIU9qx3zSbEwx
xjl6m2m0+tgBwMCMPwdT9jFq+Zhq3J+xqwCqV6eNxelLZt0t8s+uPNPiFXT+AqzQc89a5aIUxLpq
g/hPS/5bUy4HK+Q3zyG+Kk/mhTsnlnrSsS7qN1sj6r/pXQPui59iLviI7/x3WhvObRvUF7CF3oni
Dl2wOu+LGvylHujnD4azB2hYrr3wvvGZJvkh6OlxHWySZF//JuSIcjJS8Q0z4BCb6FrYsIZD+NoU
9Ko+Lei4vM25efYEhkMI2jyYqT2kd7q38KLXEHCEWvP2NxuRQ1pgGmGAD1ODIRYNcV0Ptt4tXGKE
r6JH3BDUl8xlK0oGmfiDDC+ktC7hhMbiZu0iMb3IMFK2QqsUcIi3mQDzRh6nMMzGxQwmRZqe3mhX
HP4dqOyla+dSBaaFd91gasiGSnOH7adL98hLBzXf9WH1hdEXqlG69ySqs5rYYD93PxA+9g9fR6KY
zhu6o0ePa2H0nC6BvzgHtJ+HotsO0JSj0k0OEVR2bbV1vZB1ha4z3grbhOCg6iCb660z4eHe3sZS
mBK3qULOfaynSOqsQ4gUAziG2yor99ihcS6hBZFuAeOUs8d+2MyveU+p9ZyBANT4T4FkdDMpI5xC
94qg1mdElYF3wTILnn+M3wxezF/34lCGtNtlEb8U3BNtPkB/hBnLDnQpBULgbitMdgu434sKGx+y
UOqtL6g9qAjuLHqgYrJ53ytR++EUuhdjTGS3s928yjwsa600x3WhdVcuEnpnzzgrCmUXvJIjuScp
PM3S3ArhjFwatonytkTnbrr5UUC3YJLwM49/m2F6JUhzGLYcet2RD7qFk/OyY3YRj3dBVtybCR1m
qStE2/AlcYNIUdFmzsEtOF2B0TOJpfCDH/7ErBTCmKsc7f1+Da7xl2p+np2Ex/43WCTTeGicrNcU
L+UvY0YNngp5gWbFBySD28Mnh4wlLvZYJtEfj4CTY6CCKZF7xZpTIUByFoeEYZHrRZMjQjoozKt2
LmZGdMBHz0VIamgVrNuvJXqDE6gj/ZmdXPPyncbCJfO/M16A82IuJsrdkiI8AMO8NJlzC694VGON
ujFOPq1PGWNvfQjjryr7Fj+Lq96fcAky4QMyeeeEZf8+4PQxX0tsjhbqkeCtsFNcMakaS0EbZPv8
MbM9h7jY/q4MCI4aqN1kwQ/jylKubzTsLkGrJQ7PSr+ICphO21rwZG4FCTp5jJgpBGzRgpFCpfRx
4EHGwXzE0XNmkh9T0Fc9WWZnU7US0GB1FAy3ywz1UZlDVQOkEV7QXv5aN2lAvfk98G1FQBf/XnxX
izKme8qytVvnvChMo0KrFwpunx/fm0ymJmN6lKU9v5jvictHmjfZhY+wMRQYrBa7P3dF/LtJQDuH
x4YGH/3mBRdNOWcmHBMReu4kPGklgbf2gnp8EFhSZdRw4UJF41fS60TPiNdI3vLu9tWGahKg+imR
H+mykQ3L5o0oZ+CJS/EWOJq7g/tY4eZQfxoRSfhIsn1vvKBE+OLilCLO4nN0Boi5uIy0/cDSS2+m
mCx9ngyOIh76KTigdjOplyT4Bp78dDRz7wsFdaT991g/XdCNX6ubj1CGAmReTpdkEkIZWb/q/ucf
98OV74KrfCCL3faQ/DCz2lC7Sxoc+FgiTdOvuB1R5II6SK/9iiCvozs9bgF1utocX9D72l7khuQc
FqeB/z112iLnrkWBUbkOxY9SbUbJP2GD/K/DyCxWGaTgztlx7gSSzUAR6GQItjBnD1mZBsBiQamM
x54Vi9xZ6gXQHyvj41yBM+5Jlujif5PUWDy2FKPgj85AuNpYxPlKne0S/YOmy2AtcHwkUoLApp6d
5xAcw0kFeTmNHREIG6z7n7COEKGMtJ2CFmaRo8v6BVWJvM4MsM323l8ai0qP5eomkd29mptSw6vb
15DhZf0H2lZLLkvs5NjtOLxKLtvw5q1F/2RYZWcWBrH3d3aVPzqtodz++5hLl7Kr4UjqDCCRnjxY
aACiCY9f0i1Id7B/tIzsnhyeQ6YfbakK2jRcOkn5j5J0eM6n4X0/ZE3EpWn4HU8/kBrN8Bn18oiJ
B4upIWj0uxHpLYb29t/OPbyw+HRS9U43b+bFY2kVe/X/8r6VNUOTTnYBR2L3Y8bx4LELtOLkUPkR
Gi+lPN3zGQfcJbNr5LbtDU2I/UAJB4rDDt+O5Z4+nl6juVUaLJzU7KEBeYnxydE1o3klEFBcyRtf
h7RJd1XwNjSqEP4mQ6VrWi2WsXUv+hNVOdI4PciDe2frc58W80/6H2frzjDQswB0+A+7CG1vxMw8
auJCld0wn4JMVP5oeoFPZCVhLaOn7/dZuFrJr3kIFD7pQOkVMw2qCHOnW0xnEFrCuNFLgCos9d3u
9R2YTAJ90BehYnDh3ttUR1zjiOlROUaDT5AX7HmJpE70VZeoLZjuU8E//bRFWlavtXBdabC7Cyba
WDosbphHCY/Z3NbAZxTpIVr5OLfAWGhpLGF36kdxbu5VuIu9S8UPnR9xSDGAXOWVI7oKxDIRg8e8
t4UHD5jJSud4ZbbdtrOEq8+TPXVFUpPxCGw+r4xWe0Sm35DFny5F4qb+jw2b5duFKxHzn0Y+MwI/
XrNCydFyoGkzMEFWXKPPRwUx/PSemuT0b+Xl60p2F2aVEaP4AIYnAvK6HcBLD6mpFMjUCI3t7QcU
tK9kLzidllusrBt25qGKw185gAISrsSj/nTy0NjeoUyUYl1bu1S5rfQiPfx+fGa2DF/6MLWQrjy0
t2n0R9BhZFb2lN+h3fwpyccnT0pOr+1BaQDibYefv0wRihCwsreASk/IdO96yQk/UqiupXv33rdd
hq0zPaJl1wiRJ/fyJ+5bpauM2BDCs+4I9HZJinv2hmWrm3essc5BalgSzoKYrWr0E3yd/nUf9YQL
tECi3LW31Htis2tjb5hncie1VX2hNjdSi50lMTU5MxkkAqFLHkZTiJiuBvTvbMqr6C2v9ywMS/hQ
ufTtsRgZJzdmCGW1wQPcTJ7Bdc+AJA/i0JHiDzzMzUKclS86FyAqYBYB/cAtfa7JpTGpRqlbGxhT
xP/Yl0Gqi++2bTjBsSSkRrqI3DaSHDXuMc7fcrsWByYcfoaL7cLekNs1ZHaQpBDS8hDFZvokQ3pz
G1tshai8pkobfsKpF387/8Q6G+mFKBFSQHjHlAyc+tjXiB8tBvSffWvCJJBEArxhlex347dNE03J
c0V6QMlOrezf0g5jg0kVhxJ0Cx4FqQBPHSYiV01wFC0TQhGUzs0iPeyLK3JUcKdDUiY1OjpXba97
iYDDsweejsUpQCKQ6EEwwOFu6Lw3D0GCUY4J/EgPFkJslg7rZCc6kKY5I6GrGgFJHUgjsFyIsdHg
ygpc/8kFp+m3q5pTTpB7JmxVsrfceupij20Yc+3qB8Kg6viFpqtWi6zp4anvpBBC/zLwAy3zqnzS
Fk7KK2cGSDhofnZl3AqIFZz0CmtONiCykpDTwpW1ppOJqQEqnbXnDGDLm6ZRVd7FAeJ32EP03fgF
bvljRDahGZJ/QvFtMyxP2R74DhWS2q/qhmi/22EsuRjtIm84tkM0mNJWMbgqKSMoSuop1RRTIK7S
3OTFZ56ZArAiKBiAMT2G1aFMVfjYRuY2ixYg99wKsfaOrychbo3M5C+69qiZZ+0gxdy+R+PzJpWy
7mDCe+I8k1OQeZRvCkg+DmEhbVCf3mT64Zuy4Ksgd46x8CFzewhu9WwglFKQ0Sy3p7EDfZ4jcE0i
vX84yiC1g1wptjWWqR/HK/+DrOvjOFL/19PGFcg15iy2sBFowEanwPu7zjPkLm7JDour56aKTW2q
tnCYPsOfEaXvlEYTe5MfodWDyEU7QfcZJfBiVNtBBvbMj5lDNfk+H6MLPdAzdp413YKxIK9z1SlD
C3N/ZRhzp2+xrSePeKHzG9b22FPhhT20qP6L6QBQ1lb7Lu3G9mgRLsZmr7kKnRoWrKfi1TrYDJZl
cwOPHbtNeuFnKJiQ1lsBvckCYhRzbpBtMvRCe422tms4bVaOLFXz+9jhwS30k8EhTw3shctiz1u3
pvC4ZLwzbR1dJUwl/UwpG9fNaiqb8Mxa6MAUmpDSdjlMtiut3pgISeQlxv+dX63HjMzd6CtWOlFu
3EqMU2eZofgpx7G2x0i8jsIAyqSOPGaZHopz3rbzTSHQ1s0Q7HR8oMKQlVRxHa3hCn305ZLHPJrW
Rzrc8/7Kt224oVKrH60mKJXHkRxI+OwFRvmkpnLtfqe+TKXIkKsllvFOwdj/SG4l1N6JEmChL0//
fGig/HDD2yjuTHcbffGYZEB9seNcXYhZb5A9v9X8utNb7+7ypIqE/7hOELd2yYZrN3IwvBtPDC5K
Qo+XHxed28S6U3QEwEfMjrNLxEmHNhYMM1OpotxRFtMBk+eXXx0zDS0M2wec6XH+HH0siJ8uVa2v
Ylr7+6I97iEBd5Ocn7DnELFSG3ve8yz6eA3ZOr7mq4WJZy5IaemUFHVCE0PcR+FLgNcXyI+QnUrZ
UypFyYaK8DD8CzdivSFYdjsM7PiZWWU9Oxi0hP4Oe+4xvic17NTCpA3TraCe9cQNHLsoUq43lRjx
rG0852ug3yg/BbNlO8VWiNtu1+awksslOlxxWu8FQWermxqavFlcZnAhfnZC/vqkXgg1QJNtZ16U
s6A8CfLemEJeKalnXEnRruXTdp4qhHjdCZlEt7jXejuaTJkwBz8hgiF3kykx8AwA61PiElw2w9Sb
9uzzGRTpPBISi9ku0vpdX93zfpO0Biz2TRUbeq6s/vPL8gqIX+Y/Bf16ClHG1iLTV+9ddHpQeXjy
GhtBtmVkTDzSXi3b6VgEYOGYqr1HIfpSQC+v6JNGWnMZatn27x02U2AAU6TkbGFqYGIbBmXmLJEJ
fF5w9tOFmuub5NwSigF+O4VBGntqFnTflaityFBRQTqAHqR4eXF0fHrt/ZbKRxEGXN8xFcP1HeH2
KwMl1c2GtPH0mtdBKn1CWfLJDIuj5qOIv6Ej/Xyy8sOqKZVp5HirvBxR7ZsDj5FwBHITl9IsaM1E
rnuMtsAT5domNTTVWRvsf8buZ8tKpqJO4zuVNtcH0bBZa+8M97cPEN17RGLj9cwOG5SWrbSnhCpl
hK28rmICojMUC+9IG1EbR3NG6LAFXvitVsqM6OpCCDgrGy7ZeavU+g1Mk3y06P0Ywh+BYMouqye3
by/R+N0g7+46oNzMIIOfgV0MmneExt9kUABJFoezZqnf9k9MeW0F897scmRUHztJOyyD3NgowIP6
9WhJwn7ZvdmpMl0eljko2DHsa/kSMTBaUDqZsK4FQAVA0oxHfFtjMJYh4sc2D78Uvu1Yy3cGdXpD
jvhzCS8IZeuQnilCw04SASrEi3SLx6iz9YQrAdFqA0AmrRzG1/pWnBt5O5DpXXXG74UMPQ5plVR/
rm0fPC8fum8yJymLNJdwtLKgM3467gUuw1lgYFsNMRqVA1TOs+P7OB6DKYyQdygPf/FyYBZ8RzmT
Z4KPc/d3YYiOxB6fErXu0aLFqTdAILIccF315ogl3LEbR22D+rBTaBYvkXUAC8yO4Go/IpA5MFad
T2stZMsuQTv42M3E2YIy1ojm15xGKAXMyMWvPnbpg/+Nnu2wC8wU4d7sRrAgOhj1vHVIAQikPufN
rv4FUvWL13nEDTb0hW8Qy5Y89wrH/MTlSvSmks4Lcy4XNy7lp7bOL0doVAVQEHnp3w2ZLU2btET0
IQgj+nfInbphk6xBLi9C0Pl8gGlob+wvtIlEpwwBgieBHsPwnYlShrw6IQIGORg9uc0Lx++61bb/
8gWWpKUk9y/vTFlk8DUrzYoAlLqGrqrQc1/aqv91J3eF3Ji/9u8F2RfrxTosdzGSTrdcmRuBsIjC
Op/fUxxdwTl6lXwOVV2QoJQM/9x5hP1OD/Nge+JblLpqo/tYnScurvl/FvhdjF/v927opgbibau1
uQuIB1dJ3CiBG2S7PXU6/InJHZDHadcikQaZUL2mtakdIVVMrIDDPyn8KVkmQrpreGrU0IJeW5nX
S0XPKpas07FV9pFdjWDlopBolLmWRqERDzcfIJWi5r/1Rx7QNlIAtwbggV41x0pysiYntUMxJmbN
0DGicH6skdbbrSa2Ge5JIkWe8pZdWwf5BSpaf7OImXSl8DMVaJFxS3wlh/uS0NpN5bIVOLV7BJv8
NYqapIhWqAvBN/gmCEzRTi/QvsjMc6LCQl6gkAQ0QjR6oZ8Q9IcO6PCQWpqL6oMIb6CpHY54sYP+
eBuk4iYy/LC8VQOR5jg9+OtvC0W2qj2N47sxXHckfZXDfUr+rr1r+qZYYk3hPYgjtF6Jtoy0Odf0
MpVZSn8Lpd1+ZMiZO60PDfEFLZAoXaI4ImipKjcYMHm4/PotM9jsNffIrOmPdDL+mFvVAch47ez2
F18qtx9HfVGzz7b8Hvk+SoKnWqSzu7DKBJ/JGPnfZ0s6y9JzE0kfypv/cmqRx/iQHk+uQig5vgMT
Dk837vsNCghGPKDzBUNwV0Et4wPz5tx7dQJRKeRWOj5+HELaGb5QS0JK1TaiIKjFC6cfiKatz8H/
Crsy9niaiLQPDFfXfLvfuQsj8EB8i+dwOngkvQqkGzoZ1s0XsRiZrci8IPRd2pqvDXtr7nm1atpQ
P3YQy26bCFp+DYlOSYwf1ip5ZETxPegPNkxRiG8bXJtE+UpHMO5O+8YIRpi/wRrkyy4ua+BX+g5J
DWNl84dKFXmbepLsMdzEcS0sOJ0saX9ahC6tF9NPSidbHB0N3x6v8U6zPlleV9pqL+7TFkDtx3DV
CM63jQv9UKcCms4vE0QTqKGyj8yMwbqNR8YA8LRTsmYzjQH4qnSXkjdxW7/UM6MmIjH/jiYIqGF4
CRbh9KqiodChW97SuT9q36byXh9QdyGocM70lgpcTWs1Uja5P5pzJeEu5dk1LdFEAd2QpSzrgX/u
suz3gSZCC/ZIz1Nz2DgS0ZaX8bD/3av+4f/6GJ2ochUC78OpjsnpBil+zoo/5T2ovvZfU3/uCJcS
PG3SrPboYUyTBHlvqJ7TDIRdPdtCzDqzUCTSUdok/lgiT86bnIb30fRuaCvYkVNrOXo0I/RYp9f+
hOWMXhbUiRHBYcyLcjzwBa/b9E9F5FqZM99yhUgjChstlmUQWAC+II1e6EAGMNVSiBJl23txINmH
sLsLtkGmdTwhdNdKYUgi/Xs8Z62nBL7XEt8Zc+RLkZTyZ/qWQTNP4mm0n/g8XMGVQXNyBh0vqhRQ
thY8X3zc3JRUNUReS9G1FlaXQc4Zzn64r1JhmSxYAhB4re5IDGIG/5z0B9xJQUEEtuDfElZ3GaKf
nH4y6JqgUn/0xWr6fZndiSGs28aY0wVygge+W67BaqzcODNHJURvdg4SAGvc9a+6ZDZJTJoH00DO
TWg0XBvmOrISfcQHG4NOzkIHLryv1LMZu4s16UE1URA3ynLJB3DVG8fjZDnMY8vsSw5yuT68a3Uc
DFKTHtq3lZfEN1IrBhnjF2XdI/SfnJzFPdHHCdCVJaAO5+A6SDl0Lm+j05G+gHheK3/sc3hgHQYZ
SACQ4quZAJ4jIqyhXW1/pHTR0C4c3zUV8/t8/2zMQ/Zv7R+WG/T6bsWe7Ng0o85C2x5YL7cRdMkm
ZLk8uCYOFd+Ueq+g/iFucAvCEesS73DXWNuCMKQMULB1+psNK0g0MDnGTHxbRUFPglWZt9DASTRD
1X2rqJc6Tw/1aPkLR9zWlMhqdt2SKduMByRwvcnmKOEx0P7PPJNoBl3LMU4y9oN02gGpOAj7Oc7J
r5LU98FUmHDutQ8FJ0sldgCRIAh/knJdGdgzslZc0G3L7ILfF4J4F5DAvc7GJ2Nfe86xtcFJ9tfh
KIsN3Faveymg/5D4pNckCe8MoVFBKFPfY1cNLbkO4TShEjzR6fveTIMHrMk+ib1X8hsI7T1rj2ee
dAcia2eB6oC+Wf0OHz8zoFTYiW3TDOsWI8xIMdVUhuKDFze2MpWcoRUionOcQvPhUkf3RHVRvqal
z2quCnRBuws6S3odBITgcSD8X3l04GAASQgsHP8a6bXCdEXYNWlefsm67mXqeyLHMhB+W+jarFqb
whvqZ6eVTiUtjNeFi0DxFFJW6TBn+EIw76bEURD7lSB2x5iqI4XKFtlJK7n7U12OUuuib7DKBYDI
oztwms2vxz7uKY46ZlraJuZj6XA/tO4JdHPqucy2yD9sHPHlspUGYWgS3qEeBX/XvCLyKsZgoc+w
E+dbqS3BiFPY2m02LdSLOvsajxtaJPcYtT4IW9ZUb7I5jC6pNokMEHB/bcaes3lCrZqChJZNlBhi
7kQJ3ptOB4TYWVJbgswxYQ/6nY/TL7R6N2kw9Xy2pLNrbkI4CymoKET//c7nlcz6bxm9TN9qxxs0
m8vaJsL2OnROvBiWEGZlghYGiQAj3Ys1MhP4Q4CbD7Cy7rODstgOAs/YSRQMoROAf5EZkTkqmSdE
Tq+aHG1N0QQbVenGOn2tW9rZh0op1CvKghSvoEhidgsCPGYYyYbNU8994sAGjcmLAxeYuFjOuFF8
FaZGUskhpMh330mEYvArt7ad+4ujr2yDh/yxRxTz/3ghtB/daJGh0eIsWejCtqh0so9zxSmhyy5h
HEDuhNAZ3uO2TEonrlwzjzMVI3OMoIKLG0ww8toeBTih0+x7FyOl0QfuO2KWRRjE/+pNf8z5IFXr
P6ZSr9BaT3H8pg2fbLgSr4JJDZ0DK+3gqywC+xIRLaO90DHFmOpN5QSWBexqi1Z79bHRChKrrY6h
ydWABlTh5ABs9zXmga9Wj75YVhIy2WZlE7qhMkoj0oy5F7Hz6XhrYf02awR5HJCe1+eKnB5Ra2V7
CAgSIy95OtR/b2A8c+WKHi1F6qT6F/SisNAdpjq9OTfE0gRJHHpcrlAv+iwuWMQBYd+iLeBEO/PV
LnWJ0UYKSOJTVNkngmXiG4Xuu6FovpqENi3v9NeYgUHmm2I/qnptsRZTmHCXZJDi6LUTtJU1sD01
ZUtoQyYnAHXiWG4I34lKt1bxij6xRC5sU9Mh2gv2wuBZRXWJaGrCYChPaIO0qQ9paLm7tyfv+/RU
WKtJD+ZXvACVTrP6Z0nC0lfDSLfTFIzaeFOyIpPbbM3qEuodLgKdTfYFtyK5bDfm4MKjvAgNw3s7
iOe56XFu9+tW0lg6mYn51a1WS4ggvYzfUyHdf5vicMB/v8QlRVn1gBaUEufOvVbnUWV/dWST3b7t
Jc7SnfH+3BxzrSafvp3taRBsZsbyvejevpUqbenw9f7vfI7H8PbVcIIKyNR80Jk/OKD7IvClVl76
3iCcVAcw1PdD59L3pjra23XbyqyMYs9lE0bSlfw2y9RMhk2s0tztosJXnY9q1xeY165yujEtgovw
BPtBKqv+tLe5eLpl4YasCtIv2lHW0Ex/JSNWYz0iPHJrjwaDqYC27/sIor6+yo2qXYKvO2IL4Y7v
2RVPDf9u66mcjH+iGBDol6IWf2JTwVD1c0+kHl2/ZfNz4ZQ1EjjsqLplAFrRXJ9Z6JyFKpIo+MT4
aJQ+mL7Cj6MfzBHNWuWyyFWF3WDErdn4eEqybUtXuicKMRcuEcISgfbgAfvkRBfrv/ac4pxkc/t8
/LG/I3qLDMVGSE1eibFqB2Y+3veESNO4UiotTpJi5zRDdDyEvtfd86iCH8CmqpQxTHIENfZO9pC9
2Cg7eWUiNM4Qyv1aBXY45amn3EorQFElEIocprzDdeZGyF9NtheudPwJ+JbYhgMPRSp5EXWS7Z0X
SHrGLIuciILUbqBaj8D78eATBD4enZBS4t8/AemPfA7SPBSgw0dS1c9wb+UAT5tZwHxiP8cpdJIi
GqED/MRp+jEJcBRqx0k6MRLKVN9eDSQZU/TJPmJkhaBPjbpXuyict+Lk4EVV+8hnn8jPC0S4XXvH
4AsMy9vSJ7gbIWpfCYsMzbX0/ABYuHecQ3BtbyEX+5cx95U1Dn0A9r/l12xtuQ3q7V/hf7CbW0io
ZgRG74y2/b8o6IvVWw4EY9Uvaki5q9XDr2hrPmIhFf2oGpoAiMKWWlJiSuJZXt1Dvd9x72PK/qcF
+7foRJr22SKmDSWeIpx9B6MrPg5cFy5Pj7RvDJW7psYxXrqzm+4IOPII0ZtOs6NKHSAJiKJ3I+V6
sx8gEUIZoOzEbPl/Pq9VmksBN+Q7n5T7Mp9fDmzaS8YEpaJIcI+4k9jakI98tWztWwPXKARMi1MC
oreKDeRAzi7++80rewyee18isIo8LFkf4f5sHQ/vPW7E/TGTWAUHPepINEE+tjDo98wkbyeduWbh
JiAviPbcNul7z1Y8EDDEO+KRUD5MDp/sRuj2RGA6hORGGk0yf6qmm/fxsEg5EhVImOkKy7nEgtLj
eLkXoVsKXPE1zJE1BolG0q5J+utoMz/mllAkuPD9yYX6n42ShDIKKLtudc0Wk0yLEZFinZon19q+
On8oW7sQjCuJDCp2BXYtuWPWhgVtPhB2STbj4A6p1Zom4MhIJ5SA64Uop5mfUUrhGBzXFOEXsylu
kFfJiow0FXDxwFanVN9Ty/uA3ugsoSZbz4Dz4kStxCANmG/oitiz6YE2kZicUFdRi0weXhnRoada
C+5WwMoXTdXF+D5lBZpiKMpId1MynGxBEVO03u+kTRAAxa8Khn+EKzdSORmilreSfajrhyIadNr3
U3SOGA4+vARKMBrIb71kGOGUvIGQrECarhW2we+QMnshDrbL/Ywf9Ha0YFL7lKyzAXtxEIAc9LE3
CqpX0mxMlJQ2iBShUu0Xlm0Srd9a/TcQP8H80e99v8bSMFP3Zr8eqN4o9OYUgZWK7jrjZhbhi/ys
KUM+6URwBWZIzBb+a8YO/Tcl9jb0RBVzHZGMqnI9cfNYUAiPDIXav4b0ZHPDYVUOBthlEcPyM4G4
ebnLtmm2zxyg34Fo6zsrkTR6ykBw4/75Ds3ZWTOZMRiGDYc8LoMrxfvQIXZjAaywfKJWrWMDqCC3
aHVUmKitc17qCC/KZXDXmiPD+tqqy4rpKm6t8Yo8qiA6jhYmkvNw9rO9+Mj+TSIzAMU2kBQj1ntk
x8ZPQYWkstzhJbYl5zLXES8B1F3xjOEGvu0Yc0RWsqtuY2fZM7xgwQQybscjJpGUp7ESkZYWb8CE
rVgZgO/5cVmsJLF8pwYbMcCQsvr9tYoFWkx1cdlWbvSyFzZ8ivsgwQCy9YCwLCswwGl71Jh/pBtM
4TWqiyz6nC4rJvPr+TCdGGNPUxjfgYiViJvREvMBKiSlUfDqlAnPvc4vLxsAXKQRwUHceBfeWw5D
Pa7pg4Fk2yeuoCWv5RD28qQplbcH2ysxfttxzyJmrep8ct+g3eSv0TxpHxz3bYnJo+/SrqgOa+4X
0xl7tWXaj58+aQ8+S6IwyUpG8HwJHzibq6nWTpdTU997lKt6VMX3mJG7dfYRBFWN9FYC4pYs7c+/
nCAligWU/FBfD846sCdPt+go6CY2i1VL6L1QpomY0HjGyftRaec2xGH+EstE7WnzXRWTblDeTqR9
iEzZ9B9Mjqszku7rgGIwcHjfz8ydIwRH5OlOsxQxJgj8FcJMPZtLLtEC2dMO+MnPAFpFW41A0Wvu
tBfhxp1na/bK0EgVRCYvSvyk9r6TXRhqnp4J3VA7BOKaFtU28HEOEIRbfh8cMWnZ1jugehys81xI
eHOy8U7YrS6xUlRRGXwe6f8dmUXcRe7zyD2LQIji+PNu+2Ua6hgBLMdBthj9WJPIu+Atg8PcN8kU
91kNr2W9DPdebHvWNo3+b5l2SR0Q37aqOled0L4DUM8ZzHj5QoHjhrycilvCZSkZRW3wXzh+wgpk
XY6PhKSL4TgYbQqAtBGgzPR3bNj6Ywe/bu9zuFk7HqZZul6uPYl7jHTU1F+af3n9SAsIWsW5Feco
UJTuxgz0fvSoGtlai2oLtac+H0FpzoVA2UvoFdhUsbNZaIkwExnCAQSbrbQwpTmoWFHsXVcOZk7g
4y/xdGUk4W21dTyHWjhzwap0+fAlz46Ii9GZ/Aq3fgos+8C3CUyqQ8o3H93PdMEmPC+2Xz+1wNsi
Q70QHANtyLX/EWR8jfdIl+qQ8C+6Gp9hJhMvsunQyGkxgomSIWiZ1KTxP75QwCwlh5hH5ijpTYyL
Lnp1teTzQevd2TSppJNfdNsGhGYdZN/lad7bCAeR+pRITN7NBpDkceekAAxLvsD+pXIdbCoLeGCZ
zVMZfzZqAYPSNt5NkH/K5EqQp00SB077IU3T9cVA5acKSI/f4D70ppJiV6sWTTHfjd1m8fP4ZrOe
O9yhbAnu5ELx0Vd/aTxSQU4n8mavurUMiM3N8JoigN2MyTpmyVXgdVFGaOBiRdg12qk8CiX7BqvH
/MnFbnqHmg2l8ve5VwbYzOQ2Mme4ZaeBKt+/dLS2G3JNkWX++aLJXI/MS2wkO4UijLvWuqMT4ju3
HTD0LsrYeT/MYNoBB6rGUvIzop1//wuFnZ4uo4wR4DwCmKEVIzUBqdbDw4uD/meLZQ2Yg4Knc74i
W14qlzqjzzuz69e7ZvQq9kYuNYyHCplQjeKcU+ORWCiZgDGNF1PRRlMWJxAPMAc0Xhz00bU7Sec/
7JKv+ML4m6YV1uVgXhymxY4JH+ahyFZ3A9x8LJpZ25m4eu73EN463XJhyW2EglwM4zVNirFFfiPX
sPXPqLlpIedzycLPR73JkxWJnSB3RcQ/5RqFc9rGVCL6eFnvmiSKMRTr6j1Xrk9AmX2575Ellt1S
9HHe1mD/Q7ZGIDM6quhAmG9t55c/MxLV2CyV/ijTx2/vb4P6gUOYR1Zc3vXqx78nihUK+7/xkyHh
WssniBl4bcqrwalB0OrDK2NNefx+NLd9mT1x/B3z7PwNaw/At9COGI1yYJan9P4Ook7MPdz0PcNV
1GEw1ra1TLFl5D5fBfWYSnezLmNvUz5oNns5yxJUBGrmYKXBq3WZckE3krOOCWyOB0V3stQM4cFf
yuJiqqTFM7IFF7DfYIld1d802q+0CNmeUCLDawDs6K55lJgD/LLVY0J9cFabw/AlbfBdNYaC+Sq3
2hBs/T9OXUMYbuxuX2zq1Spf9CmX65gksklqW9R6WY7ikg9CtcHoYe4n3AZeB1INkGQwU965BqyN
XABWXSr/QxFFbYxkRp7b+8Nn0OaXnEvyzXiCgroOVNzNjsNP6keISF1DQPWcRr7cRGDqdnoSrGdY
+23lK031k8BKWYNNrZOb6sk+Pm2RBDG9TR1ZqPSsDnxirrjAUmFZOwk/ELf/TRvsMfD7/JbR8prp
S1g0QBqTjxUUnV9ouBvNLDHkkI/3QWSzY4ABPwL7EppakGTeFQw8l+79o5WL04QMTk8xJwhtdEvX
ExIo7z/EfRntQd73B/VfpLPGHh6vqAVtAY3qRbwzM2/bpbDsPiVR8q+C8q2IVEhfBWEsea/q0X4B
4CfST31jqpSsQEffVVV3e8L4aYR7TvIUqLgvrJJ3KSpK7w7vmw4dlqBte/zOQKOQ8eVNlvynZLS8
2+zajx8YOntRferWLAf3zrcoi0Fq2lbMjLO57uGv32bTEp3GFoR8Pa5Hzu+k+igHVF27xLTqE4pN
REVdHPTQzwOmDm1jWBXUjVNR6AvtIMwIEuG++vavpmx22d16LXhPQykTM4F4s2jxCi0U9SyU+F5R
BAYjQA2U1uwA1qhbqMUmVqM3WX4O5jc0W9EytJOeE0gzJ96IDozRofjBUDgmGWl26DrTZL+txXU3
+KXWEYGksywGMWAcd9XhKLvohjPWUXXjtNIQKL3A8ZoqA9CbKviAmtDXzzu+RRlso8SeJBdHFONc
LaonF57m+qs+35CgplSrkz32tGcdmBu+FswRv+AnuxennCkTT7asFN7ntnYUb64uxZNzMviJfAt5
eoHQzHTAPrSjRHiFz0IpJFpw5w0B6hCGOiQ/6wnohE4/kwUoWJm5+SLLRWYboCoZVxmnrtyzqncF
LHrQuoCi56gkha/MFnFO5Ul9lihFbk7bgAsAZOMUPeqWWh9xrB0dCYa4TbvPmTrcfvWJ1XcgP791
voPVaGSMisObQSO+Q9dgim/gnSXwZAKV7/Ymg/XGx82SWFutx7KsKFIpPsUGDWfTBaGqjtPQ2ZA8
kQL38fw06hYvPCCU4Yn/1YOSjUybFK9UauyWJfAQITjmG7yrBZowIVPUEOxo8/l7BV9RUcdi32Xs
pKQJoMYQ3y+rfq1hQFdFPU0IQONYcpX05/Qg5uRERtCAbebYECaY3siF4FmIyZMd0hgh570Sx6DP
9Gect3ky8MVc5KaRD2NXyJ5E/knS2XNcncnf8RxiyQgJ8b6+aULUBEQpJqN/ZsCpSd1R+tuabuUT
60Sgt22rE3B+l3mJA/yxHNajTdct8VwPmLYLx2vwfbKFrZW5GJMqw6ISl29dq6k7fmwsWtUyLaDQ
CfC7R69tdbdZ5fGpM3Ez1uBO4aadenLCaVa4vda1krL11v5mlDwDZEDinxPyTaT0EdJTmNmDgUiN
PeuRaSTLYh7c3u8SV+oabFVGtk45S413uYsYSrLOd6YtEeqRA3x7YdfJhqVFHGkOc9FGp9r7Uvqr
ZmNIscw5TmCzE8Ih3bu0a/6h3/Cn8LBXqcA9xYzdoK8Sz3kLuVbSzsjva7M7gwo/W8EwZoPodJxO
Yy3Ho9YdM2t5V0p6EuGSGQ0YfuN/191SnrfObk4wR4IuHMLl2GgQ9oRxKY+ueaXe897zBf5IUZ0A
5TzBoTnSsFL4nYssoxeah6+j8AvBgOxDI2MCbUA2WE3rV/E++8efc4AyrLfGGcLF2MlMwutmulxx
/zdMpcDvQ5QZeiVBGUvMuUYYFbmbWu2ikRTugceqMhFU8pJ5/JQo8rrH3fRVRiZNagBf9DdJtBus
N0kofw5z4ORyUmlLGyF6lGdvGjqevjgghu3/wQasMi06VFMk+ZezK7VSLH3ZbLJOu7g9jPYoy3hx
l3U0PgQiSxu6wm0msrmycFfEZpkREQKukau+Bm6dL7iF3DgTkrdFCPGRpoom8mFItsLstFCnvxr0
plqF3f2Q5LZOZlTxL55MiD3sJskmNoJt60LSge4nQUBaB6bvm7L4A0xw9taP8ajhBEjbyorE3IBP
UifRs7p8qOzNTKYcYraNfwpxs7On5VBJwAL01v1IBL69S+S4flhNJaIGeXr5+tgRdzw0rnkB4v98
EHXcJrbq1DVnanmNp7CDB0rdAkSv6rgwrcjxhpHkHuf1MI4XLFIjA7qw3NrxkFRen/eJne7sfrIn
LLnOvmEYv6vt5chrTtqR9PL9h/XRfHsBrsjuxFLGT80Jx+vVzx9PIsDq5NGQd9NfqsGtPwXSzJEn
EezB1+Ko8YTa7t9kdiAN6vAoAydx0F6RmdPdKysDNiTaiyzW7nFBUsw7sK7FEn6RCQRmOpUe1lk/
p2xGhRIIO1QCBYShueF3yD8Wg1djub2No48byCbvM64/z3l1iWH+dFmxxOi+LmS23U6S26kTLYQB
dTSvS5F2d0SZT/Gk8gYpUQbAG+PP2DWB8NY0a6ND8aK/Hl65bCnWG0kg2V3AtdBi+Xzf2AazuY4F
3szfzjQIsX2i9DjFfR4TTAV28s7wEFkPEF2Egq9UIDqAY5yvmWk2xoZ9CD2efj4Z8Y0RY2OKLkgI
EZz4nkSwX4xuCBNkNg8fJ1xQEwIAJf1RC1OxwJkjFdTZfJ0cOggBmXnp8ynZmcxmRq58dHE4Qr3b
VVoellgNCf7G7qsnZPcKeTSaIylbiaBMc8mm6IsRvrb+LURzDIxZeqLo8yLPaWFos8OlR2rRV1s3
+F6DvssBNLM5RLGW/dzbXYlFGi/nCxmagzs21ezuhpEOkVc7Nykv33CmHaNzazpVUaeBgG/+HE7e
lRlYB4ned1H1topNZ0SpDpInZfrRDx1r/j3d0PIls5g2UQM1LvE9ZDWbrLvLpXBy9WXemLX75rHU
zLnnTD7uyxiFunljAfJ8lZaseCVNS/4aD109cwapuJbDTLztQMaZWnWyPjA7hA5RQzNCAn0FRUGR
5xC/lG8LHVj6z+XS08+LHTo5BT6xJfcTdQPglgxPSN4lyBTuJ242PQpiRoaj3OmedygtltJN+H3F
yCDf9i0/avIj/pqs7r7X8hC7VA0ZZ2vObl4hv6cPXDkLv8nx3usVp3VfuTbjom/VHAE5sx/ebXqF
I4rK8rW3HSXaAM2ciI0Q1Jy3JC2iag5K1nvNNczsPZRos3hMAQYElRA5izeGZGflruX31XXdhT5l
83pMlQkBvj65H5Aq1Aaj/x/0WhgcCSh4w7tl7Qmkw6n3wQZ2kAy1YHKRQdUZf4PNPl4eeRzQaXyl
mIQtQ3gdqlZ7EPg0GnG0T9LGKSNnU34gST2eyuNUiQngKmAxax22H9JdeUCqlc9IMdBWUdus3X0+
kJ9aRrDCsSCs/Qg9oMvyJVOIC3uEuuHHwzNR/FLJV6ygmUcJCn6idyav0ff512ySy18rzKDk5RHO
gskHV+EOmkXqvl4KYo3hHDkSK+mBd0Nm702wUPqfay/KTgdI8bmYGcnoHXlnMklJq2/XIxvWsWAw
964ybdhU8vNycOdVCf+KpG3NUMsnGZVcfatOKkgDbFxEf0icYQxumSbvnmtbB6d7FNtPXNzsTYyA
3YnnlOgAZYYNnN35yWq6GurGfbfU2XPjbPXhhnLOi223lGrJdUzGo2ycnGFt0rKujgYfSOiv8PVY
tloylK3RwwjA9lsR6jvQ6PCoq6VktwgZtGYipX/Jk1WFzGJKA7GJexwDn+aK/jNqxdoj27ZUCoEB
dKKewd1dh93wf3ubBnJf2rqBZ6cAk1Y/GYgLLI9ZI0mmqVEtaMzNP5Qwtayl+2v4E3pZf2pbjLfD
rHppCwaMbxaGk7dRxjViGvw1+s3m9UCDOZ4GV3aBPcXQ6VF07aMEGcY++sKTPLZZ4zCuUQHbzI3A
7GhqiLx5IkKNPcetOGOLYT1iVnaQqhTZgFFugP8rgiczYdwztVIOmQH3IVgI2ryCe3P4P2htcXNl
VOipzIbkCksbzVkjnG9DeIkWM+NQSpXsfljdqhkhw6XUiAwuuGk2zk4XdQAfgmf7g88yY/gnp0iE
zDV+rMznF1wwRT0eGzDl0RbNRH5pk6gpnNn/hN6iu/SnkAFoBrg9OraUz9sm1Sb8Hkx0BhhAsOgy
eyRoNfCHkdDgiDnFFRBfFDMNg05GE8ZyvNLJlkUCs92FJhqLqIKaIGNKH3M8qRwnTecM8nix6OCK
5zjTs8usk9+9RsBCCCIPbrSKQxOeH8N4vj8gFfZs5kqvL1nGfUy4C5cjp1xv+UnR3N4XKUxCFpls
EhzOirxDyv0kKp2UzW69BfsOa3CQtLjc9P7L5TU/57LeljV0Vg8THAow1V/pitlamPgsAuP+CVro
P6lGgPnPQ8kzJJvxN8R0DmymUwxPIQkx6ioFmJ8fTnuHTIRm/M3fdFwtl1ESMD7VzKWSlzIURGti
eVgJGNAxaCJmpFCXFCI+cVQNZXvVsT9I4C8z6mJXFUj6DI0i4e44NiiqAEMXG5Q0twYG+12Q6i1w
9DQlqlyaZNdUCZSzJPNY2+8vp2AJYwOJWqV8oChVE2TZAus2CMlnqWyBr8ajbshKX/V3nufXOmJY
wAcQNFFWCNlqTeVjhmaRnrrV7EYhX7NL0uLMegeq0s3aA+ftWEZKj4k1iooP52sZuajpiH91U0h/
oRC4zMf6qx6650xERubz9d7wGqz7mYDbXg0uLaQACnJldDAbn6IWXvhsOfPpNq7xtFh5l6GlI8jL
IRxl4O3OLSWpxXICW8Irv29HBY04YWuaHjblVRnCC0FlvfBgFo1MzVQ63fcpp37M55TQ238eCYpN
e6cP14wmwdqGxHXeM3NHhQPhIHXLhpBdvQg6MfN2pf3X/EGBN6gvPE1+cC4Jtt1Q8Ra1pfeYB+Y7
daHUyDPHVWtocpFeNducaDVmC3u8JNDyld/YjcAJyhf9lIAfVEAFGhX56eWTbX8LS48a9iNjmczN
qyZ8UMXVc1BLIMY2SZvpR2h9XGdawj5fJ2Lee5iTqQa2BzRF+ngFcUSjbePLKF5LrW4kP7CmjqRf
dsX0bgAYcwTdw2paefWi/ZOL2QMUkJ683HrGgaEscH1tBNdHDx5MCUEyKZboHMdD3hD+6X8GKi2k
2ZHdn5ov0hPbzLtVziCxoAN2sRpWTmMTfGyyvbXgfhRLs2ETw1wbpPwqRoYvYVlfVg8th8VNQFE6
2NAAX9b7iq6W/Zg1vTu8kVpQE1UuqDcuaOnatn8eLaJgyQSwJB0BjkjBPd5xTf9fm7y2mcDym8UK
BAsDJUeiQ27K5uuij0MxlVQGR3pSYLHpCm3XLE2Gi/oajkjWUWlWsFDH7XvLCrUgDF5EcJ34dFg+
IRwHAxXChbAqsg5SRlVyJTNwWT/y/JYVcXMcBSR9OQOFkPgguuough1tK/717Jn9ZtO+CwATFz3c
ElXIuqlM1INnoChSnk+f6lX0FBfuHQPZSw/wDjJb3Wa1T07K9Zdngx0GRWw+XB/0VbR7tHRDabbD
W1syDI6+vdbp4SgRTu0iTaEoV1sgMR4JBRCjhHR6ChEK85igD7THxiA/Cj25x2xqpchva1pTAUAl
zHnBwK3Pvm+mj24vJMAxD4XEGrGHbLEURQCk8SHImFEutrVa3aongI+FEABO6Q7EtUKFwNEN3Jtx
+pYw6JckMBbFP1fe/jqhZpCsSmJWGr0wsfvw7GzmvubZ72ftqsqWAZ3rIhSUo5TgtWNs8KV+ZO/N
TpiGdd24hHxuDL0zcmqxnw4CLiAueYpPe559+pgTNY3B3frVO8oyMZSelwRu7OtmhDQgfFnLNNHU
D+7a0lw+TTEJsbxEbDzRexdmbSfemEmVhMKZAh16JvXad8dfTIBV1BqbV1EjPx8N9NGOTETskNw/
hTZfHr//Iq0LiYrZORQmp+dNuQT+0OSReyE1lxHY9Fog0L6xZYjo9KV+Y1Au/cCJf/xLJa592fc2
qGyxYRrSdVyqO8jYqcFZl8LRDI4y0DMhOPj1et6AhyxOUhqd2ACTdX+OGa64YpZCsjhEBHvgYIBy
6jjQDXb/NWF5bVprVbRdKATNrXeRHyB5sKK3a5tW9uvsHrBireiN1VAUiR0GP08k5YfW+hLVoCvK
w4fLdmNlxRYWNGvYHYQHEaUAJ+DZ5UCP7D2c4xwSsmYU5zzOJ7plFmChksgH2J+7BJvXO94DIDkv
xA2Q/aEf5Hxlh9XaGn6F1tdS2Q2FzCqXrXKt/pjATG76ELNZ4MfVmJyXUUs43/Qflr+PXVZL5UwM
XDVkDfLC/ha7xXqLR8T2GVmBLFthalUtmyMHN5NJSbcWqeQMHccVQ+L9yLZZDAfDvzJa8RnmtPfr
JxJnS/IT7ZkKGtScMm9qLCnNZQKpOsCyHo5HeZt7D064/9iKzjRhM44ygEzKW9XAiNIqlmJiI/0F
oDRs7xifrWlW/lDNdPLObumfXPT9NCY2TwwZr9pusEjD1gI8Ad/oYeyVPgXjF2kANoolQKTl/iAY
toB+KM+z1x3AgC+WtH8fyxcg+G9lkJ+S7qkkY3j8OWaEpQhGyWuGFgy/H2QcaG7nO8iY5gVImAQ2
54jZSAa6EH66NocgAGsy+0OQ37Y6kvMsur2ceubLWA6TXpK3nNWJlFFLtgYwjVPu7xm7va6oYMPT
Vb9GA3e0AWhMcmxZ8/Q6+2wrjvbB3qI08To+ptX3m9WbsTIh1LC/2D66S51tlL0QHhpU8XEVCrKR
bQjO/KxoiDbVvUQODQuxcvPCrjMQNTRV6PYxAhXaaKXYeQUteLVYIfHW7JF9ty7dUhWvFw7gEoid
/nzJhW/9SnLgU5lpWI9XOChDAOxiSpNkpeXKK+NKihwllpKtDni3I+kTz9MNGnlQiEgVWVYYgg+6
qU9WZ9s9PzFy1kgo7aMijFYBA6UoczKO6pCS3B8H3+0FgEvzXBcAVrbkBlYKhshiKXetAUC+Z/Yw
xdjZy2K9HXqJ+wRuaLAQLWaXmPBF89re/P1HFGoM1MIqFgiaGbMDhUk7WBv0tHYgjIvCCcklW/7H
SdBKSciKABdGfcgk9aExIVS/IGMCY7d5whBAw+w005ABeR5XVUkTpwlbghnkkBXoQhKSDfNsavmB
jzz6u+B7jO0TYj6urzWCjDCiyglnzvtU/PlgKm2aeHtgvZ6mqd7gZxdFBT09vYqPTSXb3xWiAr1X
IjBdmgzNknwM+0T9q6dwAp1x3mzv/7IJrcPsdvYPfD88o5QpuJztLSnRxttRk23kVl31LY+Mqlz3
GqlHgktDn9GppggJgshoeJ1+o/6i3fj6w6fNtp95TMmsmA/qTUHroLT77dXgjUGeyxV0iFYMOkH4
Z9dRyAyK4DV6PbCfVMPTjWIwdAKOSwmh2WRyPyyL9ZhqCSjr/yAAv4ZOmMfNM8SF5EG93KH4H6Y6
PQliqCVl9pcZhJs37frWUbNqXDtmpbSwtX6iYR1wglqnw1Nx3M40hdmcPWYhhkNjLaiSj+JIIQE7
9dNOVzsU5njkqgGHqZMuqhNmvbcfGn/vEOW+lMmPO5tm4xFhWluZtlG0orJtUYin10GtIxOod9L+
dyo69j2dFPuApPUXc9CG0uddPlQsg9miz9m5SXvUkRTqqLGkvt+3SV1jYOz3AZsyGZt01vWpWCFy
sMo6I/n5r3Nlw7qtrd+HTGTBhaqeA4LE0KZXYZA7z6sYzxEiI8t44IG8n1kKpCE6pR1r5ndtDgvS
2npi1PUGvt1xBznqe6gPT+waJi4+pFqZC3TkhnRs3A7+c4f8GTPRzdiqJsNXkpVntn/cPp7wGWvU
eOLi3ZcHul21PKLNOF79rnKEnTfdbxhAhDI7L/pkyROD6CcVDiXyp1n6qPJTVTtQ7k8ugi4hHAHo
MzLDQbOT9j8i2aNdG6vV05zr7HyjROtFn0a64W2bvW6RxWv3R9Nb8EwZ+V+nrENWq9AmW6T67tSn
LcAG7ZPCs0keZMQ6VEYU0hpTTs2QI3wo+GrjdalDSC3oxkgD1lmjb0aFWS1PAA8vUO+75se44erm
RNh3HX1cpkaWdWosmEjrjKAzs4vLm8nfSHh6xgajNBlA60uzxe7Fz0PVxm5Z7fLecgg4oaq9/SMW
uPQn2Xr2eA5nkvYKx4i3+UMdDoh90VSOpL8RZy3C7G5jAbklKY/8UE4eB0oz2UtWKQ5cV+TDAknn
48djptG5cD69hH6OVADvZ3xonsJJWXi7MsovRfZhipqHB0flDobYHLSDXq1rZtyyyAk6iaUaj4Et
JrzLxsY31egWPA08Y4oyFkGXTh8o7q+tdwtccf2xIa2KbMjvnfBcxyL36YghFTSpX8iwf5agiVit
MWnAQsa8WH+5ePjlAp5HDoydQBYhNTolA7X/cM5pZlzseO00Kda9BeCbNnwnymbSqaYGmoxHGlhs
Qid4UWHYggtGRjPN/HP2eeqtszkh5Q5zG0+5A7v/LneKK0hJojP0KOJVr6ixdj0PGydoo8iLGo2E
lsVLywGTS2VV3zp64i+D4f6sMYGx/O5mrMuXmNm47069msTbWdRZl37nEVi/58pz8N7K6I4dh+Se
yhrif6CEMT9ykRMY/gxHzVHWiltmNbRZDJrct/FudzxQqVbdG2duXTAC/TSn3r0nFlKef/A6zAnv
BfTyHBAscXvQEownLb+moGqN53KnuZup9zrWGPtWDQhVv10JLQk2frYh2+z8EyqLA3/3Q0xi5V2v
L0jaIGqY1q+MbQ/w79Llu3n5fyk/XuYyCoJGEAI08DHSt/hI4lg2Osle4mnzAnXYwHorlLzT4v+L
ZSFNnDewKszB6nv4XOCFEO/AxmD/1cKOV3yJmYVYvvNG5V05LLUwvKpvJXbNee+ejn2IcZw/hIhQ
8E/pe3g2zt2IX5f9fpA0zYwRlnbHDbKECjV6bZWcQIfK5XljljLYlS1t2JHpXhgtG1wczADfP0JY
vg6IaRUIzcxij02eYVpL/ORNS/b1bQKMx/Gt/0tg4XqHcoaY58jemAeYXDQf1cnfaQ/EF+KFW1rB
spjyi5EGkD/t6wdCoEK1ZwMxS+sm1ia6IuyZQEeygl8rO/v0gj0xsHnBNBz2pXWU3ChlYYqcpSzU
fdUmX0YeMtxCFchfVk72ctIu10VeKNXxgp9bHy1C1zG5EDDiGZlZX0FuleSE06BTFTe4usCUt7XW
yBUeeONeNAtUnUmhIz3tSMIMTsX0Naub7Gs8fXRcLTa9SFriq1PBRjOPgiK4hDs9HR6Fb+BAZqrf
qT1T6sTIKlKwhAqYc/BMz5nWKBxoFi5HxRCntz6rM42ZA/qqbHthUTtNFssd2ROoM3JGQ4EZiQIi
xIEPmWvofQznBO2rSX2jYVMlZVZ0EViK1jEc/s1vgVt8fKrcd9H2jWg1OIdm3IvKp/QWwP035BF9
5NukI+3zh57qlCU+itJnM1yHxMXtRcdUUM9aja84UOTtocyoD2TVEGK7lRI00lgWtJp5OvVhu15o
ECE3tvZQX7ameDmQLvgNLpRiCFnDOdcMAGG6Jklx55MFjQ9s1fOz91GA39zT3WoH9sZKFO19klkt
VHY7qLTiLuHETU0TGd7CjkuRiOUVFQjBT7iX6vn5UKvt5yahTv/BCuXOvQ4gUtAmEr708Txyi0zo
MO/8mUx+5dPu7YaIlw8HuYIjTzIaoQRq+9SIMMGpizDT/5F7ndjUBzzT5nmrj1wTAXED5hQGsOfs
X6ASwhcage+ldG8L/hO+Cy/W7pZ4nn/+l9i29Oi33g2G8g2XOSk/yosMdyLgvwSouCQTyu6g/os7
zD0DDcfowzdfhT2Dt4SFy7LSx84HnT5zHpib0tOgAzWEPoSBdWNPlqUdtMrbPgCv1VV8tQSratWc
jsdpEJQbBU+rOmaGLbmMCcM4xiMgeFTrqiK7LSsgYJpJkRnT1DdU11iMslJ8Nmn/LA3OmZc1UXrR
h8RlwHYOOpAtucUy/FXI2uDPvlgUtwGz+imhqRVn9ZRAqmZWfsJwG0oWU3g/49QzRjoy805uAjNv
CsttL3Y/ksLomiJlGToXO+7+bli1rzOZstKEiK+VrtaFJvEPdj+fGCAsUQdtVoQawad2EHBiSwY5
C4PnXmnQ54/C1ZGPqTvmKknw/X0hKoQwpoWvkwUmgrdrKtTfAWVLg3Z/SJ0/W+904Go+VYrOfIeC
FIwPW5K8/KUDOkXJGCXPfpvBIfkGZLH/sEc3QTkk/qEvGhrbVUlJN5I47/68BLYHnFsjpEq7Hgjz
Uxkj5A72INqIZcrNogb6AB06OFoB1Sja+Y8A6ZpPfrYweuoMRoQRmGbJzUCjhmayEdpmR78ZH+cJ
ubES3aShbz43DaiX/giO+n1rLNu5iHUDLNZOsX7/quixCK8pb/7rGT8RdXfkDtDMIhZXlMFcuhk+
pm0+muGka/4wJghhaqttV3mozLQ/QBiGhCOP8Uwng8OCAzjLS5C7vUx6TlLUWmNbnDnB4Bmt2boA
bPy4tgHGF5zTFT60oWrtm39ENkdZBWBBtgDa54NpaRRU1VERmWSVG7v53+ddR5HSf4X/CuBdHWej
BiWdP+E5skaCFVR2oyjaND2OxWqejcoyPXpGChugFmBJ9TWoVmM2/wlTIr//InImiygbkjrCXvq6
CFS/RxK3J4oQb25OoX65GCNxg9e5/ZCUv0NzIQwzDinTIaz/ZzKW6Jb2ss96A4qgq2AZyacfiY6J
pv/pgj1jPjXipI2yFYIJvwu9n3cv0mJsxyivWwwjIWOdGsZRURv6TWVbTCcnzGo/x6Nnvi316eAd
St8aG+pGuZ14R3x00lw/VZUUadbObz/tusu/a1/QchqNYaIdCWaEi+77xIEHMTUvnewSyIWLRE5G
lsmKoY/F7AJaJ5CF0Ahhh/VZ1rykYubV57r2JWrJKfe9VbRg+LVyUNhKvZ5VVqS9MC/BuTxDDGo6
AgcOIvuCcqVpFmZykc494RjnXBiJuzogQ1dmUWyCOzgIpo4kxtDrsPtSKrcnOA0tf0axFcQx/oIW
9XDnbOam2mP5vvAEBohfftlcs48sTQUFdAxotRh7c6pCQUyi/j5hNsivTwlQgFmizL7iWmBpA2F2
PSFNElTg+tDk60TariWEUYtSye/3oAHod+58zxJhmZ+XKeTbxR9lFS8PdWBigue2nME1Y6z9uyR6
NHidJPQqLVH/rUUXngycKQ+1bcpRearu04ohPIhQCrRpadDhQV7Ktpj4ucpAU5kWVOdgKY2grbwS
DzTsLGDFPxZ4h0KixeAWEwuubMYAMoHB79zv9Ghw1yYoD0W5AijGmfacP250isyyuOm4wrAqNeHd
CHDhdsaC3HfOvL31mjGUZ4iWu3ZJNBbeTTAtxrdPFZUgHyliqIGjmbB9ckZC5Ycbo2Kt1VnNuhGH
60KWgSF8CpBvMFYabK7qXqaEM0z+R2KddKtXzOc+G8fIap4BGfMjzdGSy+652xNL7n+XPxAV3hGM
qOPc/kmHA2UunD8T9uc1HhSOsQN2InN0aF7AUaKgliDYSIqbjj+Yv/pKoK7vDToJzPscIyk+TpKM
/aj46VPWyPjZ5gHcf2K/7W7VtknFUQcCYWZ3nciy49HHB0YDbsUuru6UMrlK9UrufNVKXvU3siSr
sZCFviFMoQilaUzgFpdrlOn4AX8tm3oNlRAen9OpRYyKmQZJ2Jd+4ZuGj14DuvP96XS7xroy8kzy
9bs8TJb0ewoGPDWJj9HlBcjR8riQSuc+ldk4bNJdxzTJU2hWn3u0FM2OEZXuKxh19zm+sg/Gsy/I
12dUlSr80zNIw7dp5RDnl30msi5XFkFxjXgywKC3CAZ3hJhq5N+hBsh4wf9j7yIOOZBvqPhsb+9X
TYpfogK5YADFQ371i9yDF3JgSIpMnnR6NiAmBMBSBjFxPZCxd3VkQrxhmGbSZLQ350hCbAGpkkUW
ugMckCDgVxV6BeQmGuoAnPdzrOwI8K13nJGsXHHeJJulOdOambrAd6jIO6N3ZQXXT6fwbA3LPHnQ
CUDXAyiv/Njf2Rx0Asw5c+OfFgM7m10Pn7OzUBZ2MYk8n3rf+KynJvcEkoMM3CN6zEDjRgCYudJz
X61GALnLlOeXwouAqYx1xHvqsYut5vjIt7GAGh/Qwve4tzPIOpd7eCPsggx8PAVS3cto5THjsS1/
rUppEM9ScYd9gDUXXSfBKi76J0G3KU562dCvUfMZJY8+23ZnqFYPbeDXIuVnxyN1hbAd2HHWWpRG
LnfJnayiTePvoZBBqEC9r0BTccB4sbuv2dbXjYGIhruhgKSrUCssTiNmcWqxBOJWC62yMZwfOkHt
D9aZSuZ8iOzUYrcItKd3tms/3oLFBVeK+PU41uymYhsqGkrj2QKFpoiVFvADmLMr5Kus6sq3s2Ad
CC7+o5o0V2Hl0wC+T2Eka+M9KJjlkYGLTIgbvyAAGHEbu5CED/uoGXwuBQQA2yaaRrPvZOZKyqJW
w4VLCZAbdbTYJMttqzKwHUrc1SDCuN0zmujwUHIDGdI0U0WE1E+UMqOOHEW3f6OK9BZqK8zkLIIU
xbWUe+uW+7WidKbjKo3HTeO53xWTRvTcrj337AMaxuvLo3NUnYZieFpF/DB30mtCEApuqay8c81P
4KOA0CTic2GaGVatgIkwUfjzqnMJH7dUkDhHKFXpC6QhiYd+yXUdnPbXmzjRrt9hS9hF/pr8DC8A
BIUBXS/EWHURrt78A/+WXvcY8yXzAGB4qwvoMok6fKLqzsqq3KZNiQUvcjIFH7Jb3690qfjoQmxE
hB3WMKOd/pTSNEuI/2SUYxpLsyWbIyQ/NxXEn2ra2rTv70/o+/RkqLS6gjB2+PietqFCBQ28Iy/E
y5x96u9BaEK4vhoYVuXkY4xQ5zdvneycCJRfSwIGcFBTDFo6ANiCK0Lm8MLfAaLYOWcG3rGBs2b0
x+e6iWbETgrbzH8F9wCDTueUxL2RsY5Rd6yI7oLgXnV/+o2fgHshKwMDKvG1CWyNZ+VnNdlzNuEz
ArdydlzLvttXlazQz1ONwK3hOMil3KIYO9fRMn+vDUM/LhXKKWrBGiGep0Td3n1r/o1vtGB+FARh
MIyRGLJtrdvrORgAyWJIV1c7SyXXF0RXxB9VdFztCBOZwiPEnkWFAiolaYnr5ahpgbErYioft9/Y
gd3/j6FSNNawMG7wSc5M7o/5Ocn/C1miQD61VPfEFp+OQknSuokoxXqGMUu2StoWAbkcOpZoZy1A
1aHq+xZskDAttGb49Zb0KrYz0SgZJzYTK5vcdwpojOiMwF8xR6kmGgGXm01PvvdjGoZPfES4nPoA
zqhVeM6VBbEJd265AY9RToq1T3kxW5KY2dycodCSIAf3dQSr31pTFYC49PooV8xI4oARnt4/S7Cz
IRQ+OhLfS3FUXyd0EUqhD4XfRZkn3igxLuPTYhUM9Azei4h6fSCLvoBXfP3BkAHbVnmGuXwBSFoa
6e8+509WS6ZRU5U9BCDqx0dTYwJNQ3sngXPVZ7MoENetb//eVt+T2IycumbyvS9aHLBGJfl4cSMp
zi1Y14xmb97/1q9OKPLLzA6eKxooJvkB0z9X5kiJJezslz0tSEQsfaXJKnWoext99jLz0MjuQC6k
T0DZE56ypuxkcAqW1B3EOoc5dpv8Ov0kKsxDV191ZfrIQcuNQ7uPvEouZoSxGnP7c2SJDsBLVW8o
sIofpsSOlbZd4449rjYEX9ogzJRHf2pvIyMzYaEu9N3f17UG5lFR2eJNQYww1OArLC6qSqNr2cSo
QP82hqu7iEySph2pkKcMRvrHxEIuDjkg8Ohh62j5/egilIyV/qkhATp0WOddbbE+puaNQNU2LzGK
q0cORHrbvWd94tXtQLp7CleLNvuOGadniHAYTfYAnvWRexpm6p50W3Qb+B31h6iPfGb2/aId2a/U
k6sA8WcQFuZH8wedta1o4BbTF2vbWTHfIx6q5elTBc0BZ5TKTZ4hbOFbjBOmkj4hSTBUPQ3XADxb
IirQWt7jlgfIQvOZqc6t9ZRaiKR7X0Gg54nlGZND7ut5IWTN1otVznJky0vDePL6rsF0yy5X9ycv
BvkdAi8I1o5WnJoAEcv1OV+SEQn4VsElrUyg9fU61HgUgsFykOjvDLjxf6w3MyPyV/PFWD4RMcmo
MhhHHWLtE8fKgyf8bnWW5I6sJp7GTu9RPj4/wPNfAR+iQoOXyvvnR6uYG/O+8h7AxiwsKKKjDdnk
K/IQ3B4YBh+Usve9qBAr4gXlQlI6n9pWV40KDMKklZyOXNjRQlRXgnWAno2j8KptAEmk0Uo1eb0O
TGbl33t/3ZvvWCmIAmzlzBqeSgHoPbKFGZx7tB+0XCI52PSWpu3pBGvXwNB4CAj2/vGiLVZ2tjvP
nbXjfbsJR4BBzDjKIJIkJYvIuWZ11o/yv3qxx4KWJR4KgSaVtYOPRshPTWK0NTVtISPEVOWLYc0J
vT4BHm22v0Lu0K1LrE+4WsaK2yRP5Ath8ehlFhVx3Ny3WkRsVFNZnil2Ot8uVI5ktBxArjj/lbg3
1CeUuAAS2sllwda1WddvTvWYI2L1R4F7vteCQxQn2vynKqeIMQVlN4HC4SS3WJr4aXKOW/HJw4Jn
A1QYmSktFlpZI6GIhfslbVZot2c5/RnY5OyTKZFZ6h/HbR6iFV+i9/f01O7lJges4OtqS6tuUeDH
vgWx0JK/DdjeFNrUGIyn5+fPOiaC3ibbGLAAFfgnD8eT5RMb1Db/Kgbx5NdB6RBP4n1o/aTQJREz
J/sT+JTZAl0UWPYgeQOtpHNqha8k4uSz8TisFcq5FCPvuDi2R8TAQkqfn5i9sx7G/m6sZ6LrZssm
UuQyOm8AoCjd90ztyxxq1xXsB78QZJP2V9v70zueU2PKRS6i6ewtJ9e18WWTJFYDXviXpv9j0z6r
c4Yv3pUtpV6ESIzd4fsQ2avLL70SrJpZp7H2U+I2BAFcjFEAaBjAkPd1Y+5kgiwQznATVMfBFKzt
SzOcPQqG5aUbplVP2d5Sgy2tGCs46EfTDI39WVOG73P3uqD17wwNbILIPuudKyzbJ7xXsdE4qtuK
+udf/Fn4OQVFP5Ku57sdTTmq+KToljQFA1JY4ZB6df5sB+vsZfHdSTXgmunrDtn7OWvgZUl6xALb
MvGEpmgDAvC2e5i5LrVLMmSG96Qvfv9s6v5OjiRqrIy8UtTej3mAjIX2EsaDpJwlOx+L+ACSnt9q
8ac8lGkbYJiN8qxe0YCV2qWu+r9ykGJMKXIvrRau23AAzrq/1fB7TtiR2wOFxki0nBA4mRAvh6Th
KqrKsRWyzYil1OnogNLZpGGWMhcKfqrfool80OjMU8B1Ojp3T4tLk8L31Q4gc8hvhXsB3yJA0Sn/
1G2YqYEZUrEL0vqLLFBxABJRS1BIXr2xBkoyMKlmLpyw14RYrqvkYNsAiuBg1rfqeSZQ0OK/U7Er
4zRvl/7dczXU58rG9+ff1YAVHauNUZLjHDG++jh4EZi/72KGYBPGvDepa3pyFKzr1oJyUwE1Gjea
YjECfMTkV1j7heL8m06l7grCE6dg1hh1AsV1VJByoXnKswofc4FvhMCDTqW0q7bbNQ/818zNl/+w
WXOuJG3jbF85jiiLwyIwN4KkmP5nqfPZDui0jBhaoeZBcgAVP92j/gCERkW03zFRnn2V8X2rK+87
KsrvskC49fJfHZAsFsss251+rPxDgliUAmQLu0AOvZd+x3WxBiPZgTFJR3VcK9AX4ZgPd9/3qugE
1TXvkbwwdLTYr8ahcZ1wExEhS5XSdgRKXzxVdFgJICWT7zKH957eVl5Hvbqz8HqMGi8uxCB3pQgX
rVfCEe60uPpUCreglPMoKs4DoEssRuvL9XIy1w1giodBMXj9/SAkxczoqivaz5fbpEni4nAlXj3b
61ny+li97p7FHXdHrVktyuE1uCVlAKoL4iB4Bt9QX2oKKPkGkA+PCRM4dLgsJn/C3Y4n3tsppxi0
fbGT8LavuMhoMVWkrujSfsOPDuE2XGn6TSumz6rFwssyDHiGgcZ/notP/HsqTH5wfhQVIW7Us01S
kaZli4Qjjy/yI92CYdPMnDjM+MnNZ2hwfQteS233kFpePEVxz/DEOhNFHoAz91vgUmyqapmwzekz
lfHnWdLdGbTT3AOg8z8T5twPWovTLQuOZQhryIsE83EIdxzLbdnoekX9J3Xe0k6uKkSMyBQ6X77f
0qWfxjSH8d9uwG87rCJKn32fWVvto4wxYBgC+Td4A+oivFDwZZpd1tewvG5PRTtFBEUGRL5aLs5T
XRy85JUvMheziebqnngoHLmOkLm+RqV6QhomD6g1JTwOSL+7kz0ONLawBQQ0uC0qB2r57pkuTmbf
Ys1lrdijZHYazNhSpkwcm9WSpjl45u5o40zHPiixuy9COoYuGMPXCMNHeykwVkoznBpmFhTWLW8S
T/Nw2+N/KdBNW0LPzLyxvJz3/JazclwGvruCtjmQBA2XzFYIx2wumwB8YdkyRXMyvmUKbFFGauox
iaDad6CYdpEJ14R+87aQtdJ4sNpPjMhTVQg8RW9l8TJf3/j1CCa5ESn+X0TFkiVoY/ziLh2qBD/C
IY/PQzmcz+shoVpiT4L+93kQkcI/uZxGGHRKCc83mEPqxKe8fwFOY53liEh2/WojyuHys3nF5Bhn
gXnNfAsFhgIRyVwR/e0VfEezFnpo+2tl0Hv6hOI/2oeSaX9nsdyW5slXO0HCWOgkptw7flFYc6QK
AYShe/0uSKjtAUeJ9jOLdWak1RkY9nUU0m8MbD37TviLe/6cHLvGgQRLZBW9TCPFK0vEDwUg+hM7
bE+9DYSIBGkzyp2jIVR7lXpvc59W7ixSA9Blrk2vzcR2EF2oSwA3GcDdix9TDLQJZtfNCTDtEJ9f
gQbS/xs/In2VzytzsIgxTMvfXR9g94GMPPrDOEYchpZ2fdO1l2sw3X3GNvQrF7mkhqDGebk6ZgCO
oHz+IzXMY3WJ9qstnuAZ7upaosOYn0+bGLgyCl1nKVi5nbBOm9arzGtUYmXuGLwK5mIbiOOs1aCh
4yL3bGL15g/qE7Hasl3OjqWiqGzPlXn8b48q+Ea5rw+BJOPMjLMMsLlQWbcSXn8S+6uhRnV9cepH
957iYgkEg9ikg8U6ZjvkUKIJ9UvxeFjzttbMT++rxrVVpwmUd2QMKeEfpHCP2BaRTVg6plpbVzwx
LtownAZWHNknBWFkl0Fzyh+27fQmuKkp57cTe0Tt/2i8Rec9JnRo+mI5AFQC0qQmJVnDL5GBkvJR
hKIdQcnT6pGCwniF9KcYIF81Yiw4bk9e58jvjdAJDweW3C0N86ZjfFEhaMOXdC2wzqyAg+G9yKAr
6rX5iGYa56yBWaYRhf1f4PcCs6w82QLFT87BORhBSqDkA5qU51NfH8fX786nJtKphjatQ9RvHhcB
6ZcNaGu/D9BZl49dQrsOpKLonlKO4IO490RJAHVvEFnUrqdM1WGqRT2FSt6BKlEzKmoGVmb72CJI
BlNocfKAL52+QsuMk5+rmG68ECtTY7SC/wDzHkHCiSgkmIXaWGx9hbQOzKirOFZAKGifHk5sM81s
kzEMqa6yqhH+BmXeoxOG+Jn/aoLayXcu2/+GY5m5NBmiHb5IbmO9kVa/H4xbP394Xl583xv+IlRV
brUWJfDIEfdEN/PQaJ1g5qcRYVePCP+FB6AaKU8vg+hPqkzjlwgy0nM9Y9cOhUu5uNnNEM+I23UW
nfyYJWIW0q+7fJaoA9Ukk/a9Bo9DZCaS683gCrZhGI41U6GaJn+npp5n43Q6f5vbu7Ox2ymLBXRa
gtJXEeqB0cGuZog35Nu44KYsmBPI5Vpjoyk4mgR3TnQMlnsuwjEvlOxKn6rpygt2Dzs52cCaGhTM
QWQ3EzeI3G61dxWsHwbtqW7jnxA8TAeOLETx3jAOxTUmiShbLAEFOEUz5fSSSRjJIXh9chPYdE+s
57AsBUYu48id8EaYoPQi0QtQI2xW5Av9TlbXMKSGbDGhuN8dOjJudCMUCxv6eHCLGINHNEHkY/pb
n4RG8fkF0LKTPuv/sKCGJvjQ+TW4+U/14FErbUQU2CeR4BKuph86fEdkVgLVwvJy9fEL9BuCbENt
1cRrwkFE0pL/1FNK/jHWHeNNWavSj9H4gBbNkVPyneuGKu+TYNZXRVbotnsMifY7ShulEzIreQ/Y
3fDJJakHzhFdZLcxAvoaBvhFzv2Rtja7pgAq8KnUlflFrE+tQXQwiG+uNREyU0fIaZXu194iuyXj
ZXknCtvCIgwe4wV+qbQ990WSb+JSA3lr23wCsO+WXzCfMrFyqRvPTekW8eXCX9WR18BJSl87D2gg
va2Nx2YtFo58iQO7hAqw8nnQIfE5gExpcYKMGSAir8PVg3RhsZRU1HxQo3xYgvsozijK/whLFPYs
PEZoP0bwGmNVcDgKGJq6wJ0QQ5zlV/Mm1JB9kqrS9HvXg1Bg4dD1dWr6K6+ph98GhaLfJE5KAD2K
N9LP2nW1IeUhxIP7DOEMMsyhXnuNld5l0NKWeFzWyql0YxXiBtrg15K5KfzbBrZNmR+M8H4LJTUu
cM/pOihIkmJTteFdhhdiWjv//tnaaQBSuOs5x0AG4ttHVBr7nIb0Mu4rsXmllT6lkE22IXEv/PDO
/yvmBh/iIrE02FqDwdNEycdXQXEZ+QM81FuOcc5DLQ4GhEEgvCCsYPpYbln0FZuEK1U1tvF7AliZ
soK5Mud5Do96SJCTTdldEpNk/L+yS7btJis2aBwv7BpWqjINHBvxHJ4O+VMou02ILOI9LOKmOUMV
MdqD87jwg6zVy0bMLZl4czALM8NoGQ5V3ITGM4px4+Up07B4HNAq1/g2kkX4BUo7PtVMlecqlu7w
cARBpEfsY6gvrp/Nxb5i6aVy0tYox5szCAt0s0heOczt0tuwelnKDRzwLJcmYPzAWo4c7yv1gQNa
JH+pEJsIZQxt1kNQpfnqpS4J+4qWEOXFHgMxmM+z3fa1IY2jK5K31OCFoONs8/ToqgiNpQk3rlTb
BMZmv3TqVRi43u94yhazUaiI1mA+nAxT0yHGl1QgMzylznT73U0Sx9BmmRJD9jHpI8fv7nJlg0y4
0FeAXs6Hrs4QWqAxIilGnlj8Hjnm2MGE+SaI0LyS3JvbtAecLcOtPx1Qo3qboswodOLhemp4rZT8
ARNJSUbudMZAdmwjLMTwQiCnSpwQyPCahRW5F8/orMVOkniDojRrq8Lm1bsnw7I2/QS5mdpH1ZL7
Gm0ltlJN5TtA7ZC4tgr1uBmv8PR/56yaP7Xahqa52lxlWhpwGVunRac8OiMxO8x3MhLfTpLb0Cxw
K/ORCxeffI2uYNcs9pMApCkU84/C/NaemUD7ucNGGj97Kd0AVDnUf8246YUjKHmiLIZlwurWMP5G
MNKdYBtDxzDVdtvtIgjtBbLrcf1+91Y1jw4qga+xKBKaq/bNJ9/ru2kMTwS57Rrm6ESk9+VmKEpH
ggyYJq3h6aiMxZW3lrPA8yem2NzaD6d+mH316djGz/ouFaVb4KKxHGGk6JIpXoX3Xf1aFLoQJjni
rurg9l83a2+iTj3DxiG9pLcQmIUFSwpJMF6rVD0r2kl+TObQjtrrY+KEAacffKTJkX8MlKMr8z7p
sbTnVfmHn0wYoNZTAdVGVphP42HAAWj8TkZzCPJ7JNjn4GY0dCvVgV4NiG3BMGhKjhLVllEFUET9
eQb6DY4rsaL7RZirif8zBYupQFGEuZPbQN6dz2WPvMpXLKGm9t3Xh001Hv05hZGfGvuXQcJTPPRN
UHED1ED0ne74KLXUbeswgVukjuH93ZSKNvcw0u5Smsf1lywEsHjObtsNor8TyprTHPXzz5L2HwZA
k5PQ1VyO/vavDDabd70uy2kD9+FZ/DgUQR+kF9fSprB6fQYfUWWC14dyINEHeEWYvd41q5uXvVGf
uWgcpZwL+y3tLscnzJSqQbCGtXGnDte7qZVNphOYqzyf01v8UpZuldELbgKNh7Lw7uuir+BleCxp
63YkcynBlAV+a9WwNAMwBDdPzINceGYMxP+hxuYk7efWFTSsVx4hCz4WmoQxjIkSo2XLiR90pX9f
M4HS887lDkuhk+/qaod1d1bAYPsb2x18wfM3XMhSFVdilAitKaAxek8tidkHqNmeRJxnuYRzil09
m17CIwq4VQgsd32y5ENCwWieSTRipk0RcehBnn7/9ybJUD8jvFOkU8TN6tDzeHaVmopb0vJU/3y6
/R4l2v3zM8BAm8q4JSxAs0Q3Fb2jSAJL9rDKrdi3q1h08k9R5DFbFnw1bI3kTVVuOXPZWMvvqPn+
vqMgj8L13aVRI9qboB+nnrCbkvJ3EyFSToWh4WyX+ybu/SDCtNxa1tEiQNng+aIRa1jKHexOnSUw
qmwuBrU9HTmnYjwK71rbX+48pKeFwLnfvPCz67HmzUwCMrErMj2Gi4vxfQiJ/wNhVWCdVd+fZ+XJ
Wbk19O/iAJHK5OuMwvpQUCVuYnd3bgEA0ZQ0pggfIzGjevnlgUKJOew45w0BsS4o+NjdTcN8Qm9n
CyEGUo68HzpImcPaZtVcQSbcrOEpOTubRAE4DUv2BIW1fuhIfS6LVQr6M7DkXqzSnIwzRFLDBjYU
8uS7ebLj90VSPMBYlwYb9IsSBeyTyg6EtGFeBEYPBrFa2hWPDzcysd0oyQnsWj1vmnVjTyBqer+f
hlwMVHTIGr7mPim3LQ02sMe818dgEO9P/SR5DPV7GJ8OuDZTUpotWSTK6b9I4LJXo1u0FGoH5oAq
MnX5i2H3GPdSetccQVcBvnTQ1cg2aRmOfUXOc5Ie8iuVnogx9mf2+NXeUq/YN0jcaVmA82qXllqH
8gamilBJOE1wgQqa0t/JddcojuVfXO2LdEk0btSoXpd8fosxunU1lula7+DTtoplD2VHfiBDLoR3
q2oDuTBWTU8AjxFnQON3DMMj9V7TlYEFH2WwKB8HVkFw/Lgl4FA6yFkwaC2dLN1cR4oXKunf8l3L
DwiUraxuVsaKds+AaYwHmt9CZw6iCN3iA5pJEOJzx4rPGx/DJ1OiZzpTXoaqHISrpR3TbcspIgpj
ntx9JnonxfjiqyIZdNblKdXR5XDnBwD+cH0OfNKRMiuNr79Dj9AtIoO4MIBMct5d+NtNYQyohyG+
y+OaFHxdjpgkF+elkkTlbcqDXk80m7zVVjyFBjehurvjZUnkcNhn0n6JU7n3VzHyI3/mDGlCa5IK
7z3z78niIrdJ8Sps3tDng+peAkyuPjkNFRDDam0Rx4U41QkNlJruM8CQBi7NHHPcKMI1oas7nDkC
BM9ZiuixdcVIsuuDFNYsU0UuKpZ0QkGn7nVsRMIhcahKQJ/AqjrDH5DvIXTXR++8nAuhvrqOXvHx
yG2x6RwHfucjl88AaUBS/R05d/9dyNkKGSSaOQe7c8YRR7LijndUlgeyrCnpE6jLKTcg8hl+Zd8Q
9VpdcHhXIjegP/uAAkGq9+nm+nCcQ5I3zWD1Ip4QhJQMdVaqefNKQNRfrlrIAvJRP5b2WnLpdNAc
mxBFb+adwTcYNFG/7qEo7JDV5YsI9Q9qFneC6/uPGXWbOAzMJ1134ApIcSgXA+mPGuUx+Y/L2ulE
6Q/BY5/iE4HAREp0l8pNKy/01wTN23evW98zOsiOjNvfUj/2Zu7OUi/v16YweN8sIUtea5s7hxCI
UvbcLN14t1amloADzxgVR0lRaQ99kf3Nm2pnRiJkMv3dRbEUbw+c5L7rRYgSOtYVHI6h5v+1kr1l
oKAJSvFzKDUoQZ5m6qCa4zqnIlYA3eFQonWQX5jsnf2Wud9ctavIL9OICqwx3gHnCXXwPwvfKP3L
gEOnYCWgVic84JsJ0yE/+3Wjd7O364d6pqjLn9CZfS8SPLjsQsHVf+4h26rvmFLisy/JaEgwx1UN
OJ6mLCN+QDGS0iAzmc1lBEffSlFCqdZ65XcTDPjS1318culC7P5uZE6QQXo/hv0HrfV9fZ1gojNB
PsFtrQi0IfeLglqbJumpAS710wt8OLWA0/v1wt9xw1UNmOU/IKUSV+COenS+3t3M1dPvdmnC0A/L
ZOtA6zkk4vzvdovlqFqfDesjTR9GyYM5AN+fULfF83wSqbVqHW82N3pkqOx8G05060Bmid0uhWmM
lFpPkUtVG7mqcEtYYHztRcv/xP7V5eMtjVyQ8sg1R7EHw1MsYMr8mv7lPyqihxug90QPf5hV8wIE
fSXIuZv9YoAUJlQ62LAjK8KduP3e8lkEt6efp1ec5u2bgaX/uUlW8D+artWJOpZjg48pRV+qQFa1
Gom6tb1Hvhpf3fxpnlCYYxoc47z+RTcAAxEhnnvUqYJuiymm3boLWU/Bw3LUHxXTj1GWBXRs7FAw
i3YfT8qKQ6y7w4DhZLskP+f423EuI2KIoFauvA78qEt5i5WOLbPSEeAiK7ydZZ2PZB/RfKk4ZyaM
xPH8892ZwF99PCyxFswz0hDk8krf12RYkDjwvpuyyrXkxVuYYtABTYhndfqa3h+ly+CejNZJpqZL
qCBNxYOSnxPoyNZCvoQGOBsbGVrR/ciNlTVCDmrdx4yDcSnVXaU6y9D3MNuK/dA4dw+yTh7on3yE
Nn627IM7x4VcPlwWuhmZWBUrTOtRifUP6HP0N+ARtnbro1yEz85Dpdg/RSZZyiwaS2hoDvNm3F6t
/+6KPqN7yBR1mh7HBAhSLVAjxJ8Wn3l1OdYrqaJWHO+mhSViKREteFJ7yxgLICfujTKSBcjsEvYq
RbVsJn2uR72imcheVYBaHbZse2ydqM5kcSZwFKHVyQWuQI6fl+G6AesxGlkCZHxI/SFc4Gy0dUyt
u1mDQNH4LuG6oojPDkix2NJpauAR0O4kJEgGHt/6srQZ50U9jWHFEH5oFVqjWwUExeR9shey62A5
9ApDr2NMd7YdTZWtKSd7qsjVsmkK8mx+F5nyui2xHzmr6Qpj6A8/tOmo92cu8/Wu7yJW7MiEaiVZ
Ywki8EAb9b9+mo93rAO0ThMT6oyix6btkxjMlf51pDw5TcP0Pvax+6fuYawvPA3Q+N1mXlmZYXjH
6BM62WZVw1f/c7u9sJPNz/Oe3pAaCfGvbIkQSjIab8zT0nwKlHJzzNiQn/Unso2keWMyRsFIqDBb
lExQIVJDeWvZZVl4FOJAR7TONgqp9r4DXUi3ZbtkkRHcUOnSr2PW7ekpyezEjTztu0swDSDN+s0y
bOYwOy/q/ud3m9FAJj5CLeD2vOnn8CnFV19jBUTNJ1zHfoK3bG4qOoh2UepvtXcN6ZOOhjeyEukt
9jnprTHCskWdLB28vAq205rmmGo+D+MLwTMQniuBkMQanG6OzX7v2/5sucw00yWxmVJTv/26+lQp
/xqkheDT8Phcwy1xWKu6PNNwI2+iz5gdHkQUvbTWmqOG8JvrFcSKw6FuevC7oXxwgwHxnMjk7ovR
dQmSwTdAzIrGUxvAIqF0dc+dJ8nv8b0ocmDLklnu19sZRUJgIDSf83+gaWnHe4vDgmRw4Eo6s1dC
aIZb4Vn4wvjj18I36veYfkiZN9LX086HLmv+GKPbQnATvHdPia3l82OFvRYJoijy5QkjRqm6bdtd
guKs3suYM9gL+HmwIAWRSdj5YxRtNU0GHszBPHbv9RpYiL9Lnu3q/0ND2Rs1R9xj/t4h6xTG9RjI
TccWTp2/qnziqCLd7YNDgTlC+brkVAkz22qnTfhw7vFzVxM0JApbyG0RADZsiHRmj0+V1wCicF3t
vk9pv5jzVidUDl3aIKZYB5urgEvPiorEKmhOJsDFayNnhiIJKA3C21oBlcSiIjbjTCsvZlbX8AQ9
HTxWM12AtvYolDP1NFtBhsNkx/BXLhxl8IFoXn9PGnicF+FDEms1zzIuoY0Ejvy+2Ns4xTGkv7kV
wnwViPzd+MC1r7szXA9cgcsEH9FMiPAct7ktbgVDGpow5ULw/6imIzSOMzXKsJ3+11UbdLIaQQjm
xt+W6A8brWJr6yfmmCSEZWx7xpctNT7qOWZV4JLqaZmeL5gpTux9Wa9Nm41LMQWTyC2NApa2Dt5h
UzpRp3dpPX676ftLjhuGFtomZvf98F5CQ1K93wNh15ucyVHfV1J0vnJyy+TjmCIokdnsDLSJPmaV
fpyjVr/IywWRolGOYJlcMy34MvD7LYRY1K1oNG17CGssk3g85/rVo4jHy00yOA9EVrDQDr4MYmiU
pQxHYnKZhW313jP6rw6zbkFo3fgwPXZcCCBroRL4UBTDLKj6jwbeVx+NmaNXnehjfdQ6ebmcX34w
Tr8r908nS/7AXyzDtvmKYZ078NVzM0N2Lma4pyvB0fOlOuC1cAtKnv8Ey36kGVbNJP568QyXcZ3v
bKi4/sbr8IRt/805fnMPIDFa4v5DLoSOlFg9ekjma+Fqi8su8P5Vq5FfZ3iIcBlWmnE8feIMjP7L
rv41M2g5zeOBhTEZ7Ztuw9mbmY+zEyCZ7uAa+NWYMRqEYNWOomYr1IaLvunsaw/Fi4uch8NGLa+q
/PKdID2qD+0aDxGmsV/GWyduFiYlVfLgas0+7kR8Tqh8hWxwAGd1BAXsjsUkFMDWQadq7ko/Q1pP
jRZRHgHwz/aiXQqj4LwNeNH4Kc/exYN4a+5c1Wup9NqZ9OwxFKIgxkfYZ9tkyruV1hjZ20pvZXjW
QvOjYwkrB+Zq6vQx0ZMunn6QJtj2uOb80h7qWz5ZgiO5mB5vu/eQpWg8FXijKDIdVhiFJ265xa1x
LG7AvsB3mSKJjA3eI3+UhEutoIxyAw0X9SYhtvnit1sau84ZKWo9AzMLfT1Su1aoiFzPRPCAjIj+
HRhO3XwulVCjRmdOyAkuJSAYiZLYuS2aGrjELVlEfynOFrcIsCxbQqgKoaGGTFYfX0zoHImppLmv
xPyKx7v7LeF/iM6dkz/GNu3fjGzVcHA27Spp0rDJjzU+hJeIaux6zrhS8AC+LjkATEnKBf6oJYD0
pyPAWd1tP2eJIPWLc3hvRGmovakxg3XcNcyZeM/dEUdaJVT4E2hC5ABRhtwfc+6ZF1jOrva0RXB3
Lm/cD3U+mbrIesbWN3oFQH+Du02qrEcgQLHlp1DqyUTLyOwqMcgunEzZqdH6tU7xGa/DAw2hIP+7
MArIE17Js7drzweDaoAj6ppOR0QoFgF+nnpx+oZsjZGeULnj4i6hWxppqhUPyQ6cAg4x63tVRmXJ
VgDLb/MBvGgSjgGQAA0O3h4QTjIUcjGc3bDth6WO0fA8bc7bDKpoIxsKG02Nobh2RnNEGJmKGMjx
0PflIpVj6IOsUMd/Q2vKMay1UA4drsAZ8cUO52obyUlThoR5iies9QaPobko3XcP+DzEho0gTiZ9
rZjMUjnOfdCYM9hUSqX/dAuM2k41PsCvUqflL0J19GK7cHvndqmJFEnVLmNyB36s6p/MMQ5Jkpdg
Y0KM+jUIQMvz+O/K5PWS8PeGZsCXKT5dfXflcUQgN5jVOrgo1gENfkKB/TJXcL81xGr1ZFRAiR50
+2rQklZgY8NKZ4P97BJ55fG32W2m7DsfbDAXfs4gQfm9xBo07Rkmz9TDnvQ11QniRCSM0jK6Wc+B
FoXvJrckU9JWwcotu3524fAp7Unf5Lo+TdqtKcsh+nwmaRiNbjTD0S+pFjaaLrJLWARkqlYDIzB5
P59dBcezTi2yEWG2dbtUeHvXyijf3+WJQdw/7Fju/1VZCnoI3OyToPa+NfHHBm/ozkEjPYgCFgNs
zRgLJxns7k++7vyAWG/TY5sOsnvwmdTQOtvQgATgPjBffG8s3A1Ngk5nBr4CRgg9sX/W0vbeyRx5
oRCzgw9R6dJV0YiMpWwEMq2ze0Cq4VD4BWjTLfbBsMFKtfYiiN9VlQdeVT+0i/ciWxtA8mPkQGrB
l86hjQX1XB/d88AQvTu2tDGSyFjd0GDNThq383PD+mmB4W0D8SOwicLHhiKOP0ZyDaF+ikaMyHoK
HDBAYPESLf2Fi0u9jLMN75tjoB2tDU+pt+PmMpEweuwU89r1l2sWK7w/IHU5EUDsrkTPF/f0dFbG
iKGoMFsTyrLE70WsccVrzkzEufZIjLqjJooKf0DqESQqBf6PU0+6OaZrR2G6dy3PSVAAGb6zIO8V
ChaSwqQnHwxMVvhw34AnqTl4QS+C7162KBzYfNKGPQ8CWPownc6CAloblo/wGiQM0PYiLK+2jCJy
0FT1chG4h+jG7rbXgKoEyC9Tphi3UK0TeUlTQg14ua7oKSLqP8rxh4XqW+eBT+xT2kSfoqFktpSF
d2goA+223Qu9/RJdZMEToAzchUTTsI1k02CBxYGqtinhd3D8HXArtg5hvoPCqD3GflEQnmZ3cjIe
aj5ytoljWoXqxp16nNUkpNnon2a9bJiukr0mIOvMKIRSMStcs5W0smP8wIu2ZMXnucDedamogb0C
3xpOKn9ndeCDYbA5kjNN4+F68OG/k0Il1pUH5b2eRD+WBuV60fx0uGPydca8N+Zz57VOLEhYcstQ
827VGq9Xvk7BRopIk8C1YjUOvj6RUGI+4TwIXT5t4y4Bztup4roH5QnPyxmlvoNq8jkSv6K0uf7w
/YL9LYSH6Wcx/NlEOzMwe0pjD03aJNqv7+B8EfkYQbqXhm8VaBvOHh4eKgQmXkaoLDy9YXZ2t0u5
OBkVQVy8vFFlv8kpBV0De4Yt2Ika2lCsLkTbRCjh5N2iyeNy1Cvm8yVh745T5Hqc7uExlkU+01jQ
k3UXtmgyzRYFaRvux6umqUWnqHJQCdKUIvfOkcfnTql77xqhFpLXHbvEWgGA3PibXLB0N1+/VMTg
Ur3xUTSiQPQSgXneXQHwIMfZUi4l7iMxZnvnBtTmn6u0iuUmJ4Eu2wUo3c6LZgWNN15za0Qmxpgj
WvO1c8WJgLUcdrwVmemE42rgC/xa7dfVCcPlWhdBCXkt9MfqWJDhk6Hq0ogo9T+6vKJSr4RM0nPi
LPwxgIIUTTXeCh73eWSQdzyOumMaKJ9ymDyVrgUFZkeIyUGij10FqLoDSQmlmWzsy7YIH9Va2IE0
6jf2HVP3tZKEsQkgpiqKWAIA6jRIvz3unnQBKQGAo0M1SAID8MBV6rI7pONByQPBA0O4Fgj1nvhl
IW6l2UTtZ5nbgYlhpwSmT9HjaQDedM9GgyphqHXbX3ArW/aYAMBxjivlN3P79TmYHGkB2AyizmrD
8tlIY9Bh3obKHNYqEnRHeqMi/aFaITWYE1ivDWq7MfkOKJ4Rqb4CLfHdTbM/ItUFhHvOHEINrfjF
dXJYS2ckvFdfNhU+WsPpJUesEz7wb5vZNZha7rHwalF0pD/IctXoz/aebpC/Rx+siAypMKhFH3xo
+zxwo9PfEXMtCzWQ9bM0dN7Mpt8E8qP53bxFV+FIzjn7XHl+7Kc6cw7EriHBdIjif9btDnxEsX5h
jiYjZKvpFkl3lX7sDp0dtr6aNDm1YACoP9Y3z/NYc0hNrj6kcovL/aeneiuSrPuO63fQMG368PMk
eJMKEqGM7tmYlgz/m2xwSBSjpFETM4EBW0jyzf24cCuR8bu1WTC0ZUudK2onIv8vuMSPhUPrdJz5
mYvImvWzOs2SpdfqAHmV3rH2RBbSNHpQv6+vJ0teAKxMR1iFSaiIgeD5i70R3gArEt6KPXclRXAt
vBOb1M1LcKT/nBudCZBqZe1yLwbT8MVtWKr16CnG+SwjWKmxslT9xVFuMh+ch8d5hcu6WRCtFHwt
I2nNidnXNXEDxF50IfVg2tTSqm7Ki19m4G5Altfe3W00eSgJyDQtWwzlfBn7hakjH/i5zH30IQAl
utB+rDWxwgSaP67CgYc5ckZ0DC9/2L3Sd+LwLh73aSNca0SpX96fj0IXO4tjAoVdS38WKkSF1K0E
Zicxp1/m7QtfwvhSoG77Z58jSRh46Ci6KH1pI2HadoO67TaOMxFz41hyRm/3e75aI/lXuOfeabu+
9VLfbedxUEQnarSng7XhJuJvxz59U/dz5vyEP4kL+iu2BSmx8LnPaI5mPzxY9RB9VLHmSQrYGVBR
h3c8gEhVQ31FiGAo4mt3Pvah3IdaNwuvigS/VQgBmWjBuGAiyIuPtbDBBfVP56RIEH+c6aSgvrG6
GCZLWCvjbIbWvvIXFiR4mR0Zoc8zHYSOmTn3BAdm6ZuFZNaorD8vISrSrKhXzWIT/zodLyCddBID
a7eWAJpNy8bGpLP2aQ7h9rZ3tBdEzTQPVNAQaXEnohDyhUpDaAZotDcCI72CcSMOLvGhWYM0XMg6
Yrxr/olIPTQELcl5vZkFPqPsq8LMaPffKnicd6xPJRPtj854kmuNcit0Plwfs7pjhwFDQr+MEvCt
cWucLdTNoaq1J0lYa8oYOiWD+Feyezfge+4ayWsVWpN/uYjKgzF1biXjZaP/AmpIRvs4UgIjgA25
bO79qANK4FGzc+tiOFiwTkgiwOPkIZqYyfVxG22AMAHmM7GOB22hS1l1CdQ7IgbyJuKJ54VCD+CE
5qxIV1Lj0F5eFR8MwH5rtvr3zCRtH7DHrb0UH4oEKSCid1jLlg/spGmiKFwQwVinuOhTpDeBcpvC
zB/S0U0w+KSAeEqI6aoh0jC8g/v7PQq/o7fdnLnF6mlsASvKTgBSEgnJ1WIqb4sqa/G9YoBPRQGU
F4j9LC/1HpXFd2ebQ4YKImF1SsmHlId9fTk9w0L+eJeWC9QIuq9NbdARbUNddkyUg3359izPntun
Y5IRKkCHYVsYQynpwwlNW7J/10r7B0BhBUg0kuLbSk3DalI+cJKTcq50w/B2rL1VRFGrbZP9rjhX
e0HLd8q8AYOn5OkrFNR44fhxG00vIQD5ypIor1vyR+/FyXCVl2NW5rY5HPbARr5X7cfaXiryRQJa
b+BboMEAXjHt7dI79jcLahfkPI/KkKfhMab+3PWO21umQzxXesWMWduK+HP9bsNO43/vKxoNDMM8
TJy84ThER2Q7Cad87D2mZ+GSnoCfDX3jUPLxBEOVTTf4XOQr9AVq8JNvigjAtexqUU1T3beIkA5K
50+eOUHcE/E9C4WZ56g58DtOeP91U37E6i4ons3t3agCyXDjd32uKCXN7rmJ3NuF6vysJ0MP72ZK
kjW9IEeAZFUnEIWrMi6fB9E/VgqmpxU9kKS1YD90fF1VOqvs8OL9cLmyd6xYa8ifxSg1PhRrdm/L
V4EVh1ev4/7StRhHX0AYBNH9rP0GO/HjmIgJrflt1uahm3BNgEe1JDs9c5fvc1CAR99920nP8IaW
f5NBW4p381FXbYz1LtPMsUi59Yaf/eE4krGuarsMfyafy0UPLFM6q4L7XtfU2DFf4IZzCNU1cn7c
Qwk6amF3SIPIHnQyzz/oBvLOInrkEcr2KFJRhMp95lyLyu3qNxVgVGOgdwsuev3WVmmGqMPzVqrM
lmFBnhuz3c+kkbcxIxGrF9fT2AWvWPk/7hxbykxUTaQU7bXLDpXpuOjH1D5gMOmydND2qCe98ltk
YnLwYUALU/w+5CZ6uWTRWFeEH4eARoLhgnYRXYM9hf/9mMaHZqx+EN6ARCkcDd2HDDnXGi8DuQ4d
RtR2XPmDGmDk1tZpqWztSSP3JTKjOWwLo6f09Bo2l5hpbywh4gzFjf//WrSdS68DAJKq5nzYDYN3
tIco/2grKnH3ptDRJ15uPpOSGGvZ6UWtwGGEVo3XwdKl7+Ir76wraGqNPkE6UTR97Rb6Y1y7JtQI
QzNhO/ASvhlifgnvhaVkMH4Bq0erlDKEbiKukla5adsLU8aL+/jFs1lVTlOWPAULLW1eQTvUNa3d
lCk4EKuIAMpA0MNXnqGQiMXK9UUAhifSbu5Qi7vrcDlzfJn3DUaLIoTRKopf/KCoiKzzQsCIS6xG
ieOv7qEeC/kOGXk360orz5SdN5TV+tPfSDpvsMaYU+9QjfjNZGF8eh6n1Wn1wx0D118EpwR1gt8z
EqWOzLp4YIGUM2ne86OY+IZBdefYLQ0JfbfSyqHEsKrHFhJ6lu4Zmul57j4fLYosrf71vaQFn35p
2c9qE7g6OicUGj8oZPSgwUydrkYG5XMakIC3xEqFH07B4Kg1+2KAEPWEofTNUqay4SE7Izwvmk6j
VE+THQMxQDWkBsX5E7P+6ctGGA3DbbGqhnVq/ijnx12os0tDnxdjDXINQ06FDhGbw9wfX1keaQ3k
d3QixYdXH4vzY8Fyjtu7wKZUV8lW/fA4izg//9kIXgPkxVriZPnf9Q1zKzVw2RT5x1TERCuXg4dQ
323wyb3UWsVyIgf6KPdLCO6vg01400RcryzH6R4bQH4aMyLQMzZYxGkJh1yDOK4g6265MYnMByag
buOdWesr3gMqe/+Qw5Lcy9Ce8vea9XwOJxC5VpphE40+HjNuuYz8z+HvMqtQ3DgwcdaS2GBc6EHt
9RMq9N9L4Dd68W2Kn0dUR1Gt+wFC6r1tX2J0IZzXULkIzw7GT4bFeDZJ6J3oD+a51dhCc8oVegXh
0kp7fAud9IzYIe1IOJWeIm0TfwTk7DMWauE4Fn75njHnkd7cDB5CA3QPMNI3h9RKF9TTtYlPIQcF
5yDxTc4htx2hgneKzALZ7ameMYraIQIcMSi6cZY4Brebl467sm5JcqyWSNlcidnreH3gcG/F/vYy
KXbI0y6gCDuE3H944bj6gwLuggmxvc7vnADw2Pm97KseRJQ+4w0KFs3Q9csiF961rFz0dKfaj/GI
0ckRt76HGnfDROpKNcAvktYmfE9hYvcdJH/k8dxoTk47u50e4tnlTD7yeQbnyKf9hO9fH7dK6eOd
1McfYCtNLuxINqyJnN2o6HRzh85ccbXJllo7XpSN+Lkuebp7DdAkGLSDgbDBFW9nwkeK2x7nwYQz
GQz19AE76bjIubp8Hiz9dLrMsbirxQv9xHmu4nMFQ6uMz1pzW/HZcnx9eOG65t2wZa6icrTVBa8s
eLAnVnocgrTfPqe9Dm/0hFIHgym5tazNNpqJj4SaHsG144AoEyycm7iwuM4L7jmxdO1zBctvgpq2
G5NlaKUyHOGPs+WDOljyKfjf9xWGhdZNUt6I0v42im2CoxFqemzpvx9ZMGa3LG3Vgd0fJxhbjxVC
mxP1+wPTpl6AJEj6nBjpxgXgQyP9+ZFYlYmRSO+gpu0rNvlhi4QVdTbjvp60hyQD9bsAAEOXXZtx
PCykwn12vuO4qaTd1qI0T7USuXJ+MXqaF9BYcublWrs0CL1sA8GvH2sS3xNU2CEMu9b7YewtPAmE
gIzydrpDqRVf+7W/wTnlZu7kFrQpjYzeDoEm3L67ZDVLDCPHZYBIFZ+oEKIa7Hkqs6Sz+TvFW+M8
OPxwvRuOkKuwi9SpzNCpxc7/Pr8jA6/vc6eKXe++rzjF9IBNJIio9AWwVQ2nJ46MLSXXnQ2JCDXs
hPbGg9GeQtMqFO49QJ6B/Hope6t6MtZj0SrZxkXig5JgPkt1o3Wkw3XgDILJeYg16YLJ/9tJ4qvo
HmD5qXd4GEdrO2NXmTRP6lP9+aJvE8Nx9VQtzPMvosOEnPcRJ2w0q/XJZ9wgiN8G87tDNcpNRODG
SHtmfGmNnZkhibv3F2h6mN98fJT17BCMj7+AR91spWuVArR6cbEyhl3/rdn/hSTWATIUO7WVngPk
7EVyKDJPu0r78jXEt1AYZyrq3/wyYrWXS2yJqh4Jtolu+2MirXbc399nsBnbG/eVrYL/tMTRUOrU
YKb4sH2MSycSgIorhI/5s/16drujaTKcZVwJWVh8zlmqi5MP9r73GFlUwbzTG0ESpUMFRhYKgWiY
FIsU5hiSgt4mf70bdEJdddIZqIy3TJoYN4E1lIfzroh0EWnOtQ0Ab09nbpco2r1oLEaRkzPbWyMK
apMyMeT59xUeXCUQQTyahxZDFpqZgGRVjo/FOar+mJFHW8MVCrUfQTWOEIpebkGkCXoR4IIHMqIl
v7hXf0WdvY3cTan7BUq/DGd7XaPW67Avn5uf1fqBUKD2AXhcWZ+z4Kv870vsDjTDRglw46IWgOb8
h3Ey6+5onViurWYKWBsAUq/Ose6JijpPRy2PsxYyQ/yHl4jGmlU6C7e2EAEQZswaZQE+1aZVTDPf
Uo46znVUXfajLuoHUWVga3EcrcAwcGFzF7xpMXl9McN2aWGuj2m8wfugGhWz3BLnoHjEJkk5nuno
do9/PybQ0enepWLkfo+twpcUvq1kNEnn3srEUvBMDdVlL1MveS3wYrFWyWcE3Ks8PHG6dunAVnmi
ZFnXnmTc8bkAyritwE9pUAwpjFmDFT4jiWYsdLzANYeM5zlJzqOkEmnaio0wHUsgjUEOzYJoQXmR
E+PEXfWQ7dNNb6ZhQL6IquGMGdA2Xufq5w2h323fNFqPcBXJYjmrS54ifOoLWEr3E3up+YSUqH7Q
KJHGrQJFVlt+zk9/ApiLlyvuZ9YDSjq0USm5oEOfrjTOeREY62drc0jtXvVcIeEhPsoFzhn/xFf1
r7jPHGz1P4VTHvSs5DEqzhtC5PjFSzHymxumdaFEB92oFWZ0z4YJyNpFnrBS//58p5HZs8xsLWlr
6ceqCO56hTHYZVGmKGAOrJ49UyElKr3asv52dzYPi5/IQZfd69kKzz6HTy7box5695EfP89GQgSi
ksDZ59sHHAI8SUL4gDnDHuwuA96i+BzxBIlRMmwNIYXmRWLFzwJiRdh4z3Olv8qmxluCl6tt81pQ
8GbYVvEp2q77qPQB8jzGBpLAUz6hbHQLUO73I7C2qQoXQzV9z13IhZtY+rbHuc/7cMVWfT/WaMRk
KJphpPBkdVsT+bZtNpeLTliiNVyXxckwuD5vZ5EfN0z2sQ4f4sotbgCQ31yID3A/rdsRVFIdUJNV
Aa0GWgvM60PK6xqcXX/7Ero4U7CsRJNbuxoBfMWhM0KpJoKZfsIWls5rajr5v2LijwHKUq3kSjHm
+yR7DtPpEVtSCtQhZmPtq84zPx/6+S7adtiDh4eP8cjbR6B4aX/kv//BOLA+M2OfHkhvspxnfYVh
9bgDpe2O5pmMuxfv4KY6ZYMujX+/WlCe5+BA9pnXB0Y1iXz2nblLxQiKFK0TiOHeW4vGC5GLls3+
4hPuVSzTBM8tfLF8ni+UsQpygTlHF9RpEvRVPHVR671uQ+8boj7C8jICPvpn8IK3TiwRTAwW9lUY
mYBUsgLovSjPsHfuMsxQvC5s80itmMDJszBpyFNREsvDNTdVdeI5psU7oqcExkxA12K1IItp51pm
5qG5i9TbLalcxP61NGQvHk2bDIu4xD46rQBRFTmu5Iw+VOlLQ2Tu7URw+HpQVl5K5FkFFAAB8lzc
aKFFjnVDE7Xjcth8G0x4N3rvVgmet4L6lOKFkjR+tovEC6SAsYv+qa0boiKruXzZcDlW+1juzmwG
/QQy7cTJBushMCH6OxMrf65/H+sk34rgPZQ7DKiFOMHUmi40b5kJhRsYFS45PpEre0pZSG6q2P60
yVX0C/xeVSmhnrbxAkDB6FO+KHcmlViA+4/d2ck1kh8x+Nlg83Wpf69/xRXXCY/TvAFCDmEc77Ik
YjVKJSE1HPDh8mz/TbTBCcOp/atDTizpwin/wv2gaMV3WP9UhU5S/CrXr0bX92flfBO706fuXaIf
Y5bhYSGrS2atD2me3uFnqHcWUkHm1MTbRbqo9eMQOFZXB15mHOhjFReW0UndK4itK10zSsNlYVns
/UiDNVlQEqQqnvSMnmUqwa1f7AcEoXeHoRSbsIBAwrYtnCUKujANK37TzHV8DGI8dgG2rYrR8GOy
9U8hVlc7Hpsvs61eh7p/9YiK2fLbng2QOUAT2lSg1UAqufFjkdCZohVEM6JXIlMOtwveD+2WgnMm
Wlv9jrjTf5YKTa63Prf7Kxy5aDpNVAke4rUxqSxoTmK3d08x+zoCnXkxMv2oc3J8MQeaIotTwZkF
GX9lR6p3mFXN+s2FrBJgD79usCUuFZOqZUSyrY9AfKuZBT3nBgbu+Jans/f2aWu81LCElvA0Lfqk
YnXfIKuzprOyd5KmxIuHDsCRwr6/VGhTx5JXooqWLUb0QDdZEvf6JrwCneKQh3XEHhZqfnUJnNi7
tNkDnhYqA87UcJHJF9hij7AXQ6/9JywmM28Y88AOevXsddZ7epiqLDyEUOHxlRBJAxNL/m+2Hp2F
In2rAayBvGanO+Fp9xobsyiP8O27rEx2RD+3xdDedDuYBxrP2I7w237gKhuf0/f237/9GAy97GRH
qLRKklcMPZOwsYb9Cq7OHI13KL1H6iGiZYWxGpwh9DOJdbotSYmINqDXTZ3zvMw+vCFXV3kMniO4
D+RuwjdDgzKZlb3Qs0+WBlLWTraNNqL5W37N0Z5WeZo/42uA9y5fwMUOWit3Y2X/NbVRc9gg66KI
lhX9KcaIkvAe0hd85cZI8Os2YVKGWcAeOMYGzv5quFMjCosNlXkfFM6ekewHmyhjRFXqtwCQeJif
QgFjS7dTDmMGOia8NUlnJj8tbDOH6kMameXEm/6EDd0HVR9NubokoV6ZzYqrXJdI6Sx5C5rDuL3h
rKbrF2UkZvARkAr5prDdmMDUfccDSVL3W/quf0OH3mv1y5Ro4Ah+7ZXntqoqCqpDdqFt1EQbTKse
TDPAQg7QwonHUGRF36rRzTYGJ8zU7uiSVBPOJ9iJ0EFtOe7bhVRYEdy1+0fEXp4ZKLaibvCPJEFc
bFLYFbSZLgMiKbNjfsU8XSa3Pf7Y7+NOeuPDAnPr2oZlFT/KukXvesOAS+r/HrqzH9PvvDuZBzJp
3i2gkUBSxvK0eTc1jp6KhvVe91KO/j1pBJmE9/w6PRoVifJl+mjVfVaCKxwqYSXdKa3/WY8NRydu
gNCTwvlyp9BjRZO4amfwVoNAXQAmzRPC2uvVcuF73j4QMjVxgZA9nvKxEB1CJ598vKRgSo6hg8l1
uBDyfFZM2iN2UAA4Sj0VtYMK4hhbQMNLzV3x1p7XXzOCKZZJYfHC6TUU3Oel/KWX4grWcICAWuzB
9tGqbbIwdCLv2CuLGFT6kg0EcRiSfwPIjfOFA861kny7JyhL+rENp+XqX8X8eUdL8PvxkUzZ3+5b
OBy693xGo1c9KfaVK2pelkMj7oWec4KSm/rmW0gIs6pysC/trMaW6pv/Z/ENuiaiXPxhqHaTsXXa
679tyrVTW/KJhSNrUDKZ3F895K5h7qlRQk1a3i1froDm+p1T05ulMF8YlhUY8jpPLQF3JWd8fPez
XQW99uEtJDqMAGDeQxpYRzRbo4KYnhVPfo082fIgHi22+mQMS9GxQ01K6aBwj9Aspk1loFe9bCH8
Dt0+mTAVwjHj1KzhdccNfz5OIgUQg2WBCrGeNYhlTnixUuAiS43AVvRbrVUmCf5JiyPkIH5DMj9+
f/t/YtPI1wvxC+HB+SH8/48iIt2XHVYE0FVdv2mWzJYbwXJiwA+Tv+olWZvT4N8DXKhEj0xYjOqy
VF02093XztdEz06WF8XY6wl3PKs08QjDC/b7gVh7jt2k+S5QflKridyUlsryaAcZq4NLracDIyy3
LMXUZI7WY945ozPBQ9X2dbSYvoVNcjke6tF0V9ySG0CmBIbh32Y2qUyNdBCummmu9EorYLIQVlTE
0NUwn2VKqA5k/T+oQ/J7nHuzx9DyNmKjmUjySuJVTfwtKoDQE8+krZHgi9r1n4v9wGE+PD8F9oiq
teJ9aituHzVso3BH3LzWeIaoWrZHz9WnoZsvJHitoMDnGiamfsmzFyhb9mPkg2C1UKPDjFY/vUUk
+bMF5rQIpNdQOC0ZsJIv5BdL03YbbjfMZ1zX74e/hudG/WPvqbzfMm4kp9WGaUAgwaN8JQU5hkrA
SVYi3dgxd8jGGt8fIhHcxdMlFakgHmak3pMm3x9qLv4RRYCulqEyE+C/Blmee3GL03P0RAPvvext
Rd45BzRPDZdEkVuBanjRFxOl6ysMVALRsjQWtXBMQ0xTiZxIc0ahccjHM8R5se4AiPccvH12T5fy
WttBKJlQy9ahJngUMfgDwySbYejX97etBnSLB23kXzLGJlf4yiUUEo9VYwEfjCgUfovp2XYXJ8ph
8+/8YorNIWDHdl4OgeKj/4gvqKPeKnjpeZdMVxOcppdwhxNoTHrOUjtulGf12Gfo1ItJ698CBaFQ
mK+bD0R9HX4zsviGipasFExk6s3EoTmA4eJwUKAfD9W4RXzXpxEW7+3e/Qm5pqWp5qTX30MhSey7
blWLDPVRMx4cCmN2aM1QDeIR5uRh8JNwbnhRl5WvpXL9B1qfERQTEgh/uaGl3QM1YaeZtkDPaeot
BU0oyACUff0tMEt77bBtG1XXj3MSjGYFilR5xpJjUfP7VkGEKHzUDPMPR3HqEnlC3A2uqL+WrHJQ
b88iy8lRRCpFoBagV7NFbx0PHsd4Bc67ejlxenxd+L8f6ofF3EZ/hbRgyCf0PaLgm8r19uorq137
zpVKOW/S2fi0cUiB1NNWYqtE5AD84TB7L877mCFNKWHn2nvdFTcNiri2U7WfmP09Whs7M9UyWEYf
8rYbkUGboxU34OQInidUts0iiMJOqONGsNbKEt9eS00/V2t5+gS4JNz1tVYa5CAU7mLmE0MSd6Ay
rmmp+lPSxt+N27wxk20cYMEmrjDpsmKXD4OyY8+mTXtD8wkjD4ttlT9amrJx950oWnXPLPOar00o
0rI6EUJYCr18OfgEBDMrcYGHyvrwc55uCghOCbSlaVBUwxiNrdgfFoDM4uYYIE678b3oJy8TZwnj
I+DeH6leTs1sIeca9PXv2iAlGDNuMnfzAziGRp1QKcmgFbDDGfrISi1KU9G9e6vl5c/mlRgwaPWC
yLqGC+wzgJxxDXBzNT/teicEqzmr1DmsDRSZ3THg6iE+yQwGtYBDy1DXROg+UW8+6nxRbAlL9Pdy
jjN4H5YD1JOLRBEL7NM1iCzDZ25kj5De7IH5YKLRBr5EVlH/GvYXPX95MmVvtn8YQsogtAbjf8SV
k5rTZR3guV2BYubr1lBNS8++rwmGWvlj/7yIdDVtMnqDzgDS4N883sW658b5LVI9a3uJg0FKQKB4
j+Lel7oBZXbwV/mkS0tD5lUpdQM29ywJ/nyc3tyDmj6GFIpNwIgY0sY18k4CICv+mqM6a3mlSNcw
mZdFR7ioP+hSn6EvpkPNZbxIitJBXyiTe24Rl4a9DT/XkWel57LhdeoL4W9IBANCObwybsJeMtI1
daa7Erw/J3azPlhDXYBeQgiXVIzodjokY9OJsqoWQbhvLyRJGCpSgifvHIQci1RrJ/cxbaGO/dds
KNBCm+mzHhuHNnZvzx1DH7iB8WE6xZJ3EpQWaQDGKpX/5nJKQD4pPasQkSEAjBBq9Ntb01c2lYEo
3eyZjnIOdlNjG2oX7BjzzE8zY2lya2k1vHX+2pIep504teMtReCisWSkwC769Sm0XXpgfiKjZe71
GQrgf4NK4csUhw9qKntvRuBIly7ELKiHfR+3Hv+/o91JqRisvlD9fJ0bKZtFerZik1E6qkKTYO0o
ZT8YYcYEnI7l173BFo0sm4DNxqEvCBwdms1G+n4urJDOrna5Jn5lMF3jyAJBgkDpSon7YzFjM7xy
Us/9xXiY0JX+jn0d95HfCqB8VrZ44btBCy4F900up7Lz6lKbhEwMI7X/K+JU5hp6TX49JX1wqvem
9N4KXQjwK1AvUSIUrvzL4YYZUEKxPXLhKDin0s/VvBt4tBoxzG//yv7NlgHM887Z9FzFJOP86//P
iro++bt1c8TMgnPlpy1gC5xI2AGmAaY4cx9NrB08M3ufrloCv/Ftn/Dl/eXxdkzHtGRqc0B0sUZA
e5ykOI0/iNNQpbu1Lk00gEi1E+gTL4ohitaOF3a3hHR4N54ucrPoVjzD6i+gAeNNfb5RTD7TB2dP
7zGDjv62F821nTt5Y4rwMATokF5M5ia3N8ePZ2B/EFlrTc5vl8IRwqY7JQpLstzqflVbjT1Hvrk4
QsGKNIrdRatlwtUE8/QIYXz9vH8urXDzQBlwllbv0JfAxVniDqCAxca/tezP0CPcJT4yU6xGvRiP
rKK8yUiSyFY3iAnqZP+SMR4+hb+TFl8DU7MRNuB3aWwqRd17CVHu6h/78VBYkX+WOOQwIhOsr9+J
mYJZY+R0Ct0shB0kfRBhtwMPSzKAf2Kn7JHMk5bpBeSRJDVKxl+/GxI64ZEAI3GuARDBF95rJced
KvlWqI73q9PzGOzltZVA3KVUJTPXQHtuxXUb75kiUHT0AyOZPXP06TNq/n+DKlBd9LQsnbrihZsE
27QXHn9UsR0bQAHwiBtCzm9J3nfsaNHATijRqHTkDEps6vEJ2dUg7nY9+tbyObJc9SSPk3GJjwqX
AkwAPmSPmmeZhfVzjH2QWXDpBKMWvQ8X/LKdUJ7cfdffRNXUlb16FLpLOd+A7fF3n1am/xWkkWih
grvT/EVOOZQu3LSf9wMd5fioQh8v+nbDdGaC8+bbbHUsD/ZevO6D7x3hAz+qvZ0XNg/s+Yqs5445
IIuNMESua/i8GAEj+9vXq/fyt51G1luW2QBop0SLAp1qLAF6RNSRhdUp2ITVTnKBqESABxel8Uny
UGmC4/sknaSV3HOb+9gnLU7MLmB2hxeneXmksoWj7G0uYDiaVcRzq9xspNpGnd72ktvdTbEESZg4
j52FAmRhrTBoIXlHw8j9rePh9Qr2bAiKjAb028mRCKaGoSEzWxwY7vPfkWrkRNPT8uYYWexUAsLx
p0nSW1tGphVxG3nkxEnAbj/+m7J12QU+jw0Y4xoHGXCmcI8UU+796Y/nI4QYndHQyyfW8Tj9iZ5l
9CyLTk25J6WVL0iicZUdN+dtu7fzVX038pOFrA+hxMAUS1mTdjnkxzpaw4a5SwXOmb6XiRKarwnC
m0NXQ8FVF5TsJ64FDr9RUp2c28ubHO1O847HGD3Dtc06Aq9Wes/YqGq6UgFZkNM5/3RTGagVnzb5
f2i10DgO9UzEqfb14HhBANslBIZiVztFyTSa5N2I9VOo5hvd9qtRx+9PDy7Vzb1m/zdNHOm1prJD
xbIoUjH+3+pE9lFzXele2DN32nGjz8b0x7m4vl0f2DdFVxe/4RBOfsWOC6m9nCKCjCc7ni03kEGi
hUPemNHCvO8dbOKLuJRjzexfNpnO3on8Co+LJNKFMQJI3ES5tEzMoWShWBMNd6rsXMiqmM1uGE+c
Oal+P78pabWDTa4vRPj6HdNkZ52PW/WNLeUKx7ayp8o6B3lBDdtLlgB6k0163hc9/xCGtppK32wX
0L9KBfy/jNfVqwXEl1Bw2ELQ/S5xNkhVOepMtletrJs0l9kYZNEQD4BHdF9Xh9dL5L4bfSaem0me
j8DNcYes1mTbMYVUimSK07ZuHvLUUybbjUThhXc/ZhaWKCgz1kFb40Anb6gmRmAObXXu3Dp9xCcR
I4J29pjX3SbnSeEk/Gi3lCCrZtLAne2Kuox+ZrRNktMSmKU8pCE9xHOgi82moidSqqA3JUiflcJd
Cy3oJ/uwPO+Ovx4WgfkISQju05Xuc+oJg66MAEQyvRXH4WQlWsruAFkJHQ/r0dtUtYczxmsnsgdq
59opF/QnG5MBi3XvHWRjPfnSZMacau6drlrrac5FGg29pC5QAc7kpEJcCPbcPzcXU0wf6bIb8UKy
uoCDOfSU3tYtA/QvJskZs2prFfF9y7uZ+DFKsHDEYicY30T5EkmOFq95j2SJlMEDI7erZpcI4cfi
GksIC+bAj7VqrVzdw4EcI4rvkAuYlJjXXAT/rVepC7Kodcn7+9EDVsg0h0u05jeXEmxz7D3rNmR9
I1Vtx696VIyt8rHM0hIMAXFZ+42N9dIdLd/OzESbQ+0Y1V37AcgeDs6e+HgUUgca37slHV/xVVIG
IZ/Yq9v/TFd/Xq6XN72r4TObkXRsI7V0wc/t8jBYNT5e8B5hxQQIqMkomXQh0N/lH6B1LITknagp
2XsbQHJkR5YjCeiKDANebK+VQ+yttCRkbCBHA743/k6XALOt1BIBzZ3CTGo0Ey8hfm6M23YeWmmH
HJOvOKijIchUlqhouBxQ9WhPzh5HchSI0BvDb/oVqpZbFMG3i4Ka13l/4uJH9EkqUwEbWMYtyfx2
iqyOR9iSpFJsykWEb4rOJw/Dn5m1h7S1Ehrvhe+dH1QeNo0pp4dxF/zKfV6LiZifKoBCB97Sj49D
iWY/P6FWAekdNRtpF4ay8KTyNSpOH10XOKteAE6qLCKshAMCkaBBxuoWfV+crcen604Y6TkBYkkq
SD2tX5FKo72K+AYPAWv0HEQ/w8WQohn0mtIElA+WWfm2Rr5DKwREOpqec92QrNx2F513YB/HlxIp
5I5JnfMMed0z7BVbzVOA4GQMn7cYa3GvSBkPOTz6xO2W3PQlEfVRFqNxFv52IcEeTeL4MTygQHLy
9Es1N4LJBUXa8TDxFX8Y7jLFApkFklJyIHQ8s7sETFJm1w8PdXi/D/AcEW9qkKYrqG7Bq08DxoyW
20nlpl8DznGUkKdzQvvE9hL5AoFH9BWHlxWERp6Uk6ZNgM+wZptIInsBKtxcNq6q4U7gg3hbAd3G
JPdhQ9cJZpMd4akeKkEgAflwjRZp2JMnWD5KtAL1foh7uk4iw7F1jmYGSxYcZbYAVNamwA3RzZc0
SZTBh8b42/PW4OCCo3NImmYbSF7b6FzXlrxKWFZAf7D/7QUMf2e53iz/pSRBzf+1ALGeSgNkRkIj
63cvilvAM4PthKXmf6MsSqqDs+ExfmFVYqerd7cnUwiHyc1GaR7JBb8nlhU7Jl1iHRaOSzjzbrni
wEL/gf6oO9D4nV1i2uLAPDNI8v8m4oOS5VcmR6itSaK4RiAmXq2pjCY1hnNhkebTSzDpW3qmeQgW
BjFn91RbQG3qI4nAIE3mHITZKguCEthnNtf6N+9V4CijBRbb8WZQ7C2W8vt/NHxQICUjDmFxSeFT
m5RdlYB3GYM5dL8tu9MnHkaxgZdV+SDpMlpiQSogr4gTcRKBxx0lMBDBwKODNt50VtQn3cTt7pCQ
IFOfpdyPWplD+gI9lJBv6cTPVxRh6JgV7l+BysH8blXlqMUZ33dc1FDat6BHSijS3xwPiVpAQQzE
2gUa3bz4Sj3+hWtNC4FtsadRfhJ5ak69tHIPUKeAnf73K4l0JA9LwFPepL0IWvcZ3e/5i0huXJfp
l5gks2nD0fJQ9Z79yWyCKPuihUXEm0/M8A0+T/FGxLl1ZOK/nZt3QE3dCt50kqxW2ZKiSLoqc/3W
gPJvyF0CUAwF8FwjXJzUOhZ7npbvH80+NaGdOext2PiNXtAGUQCwGybfkCPB3k+oBu8g+mLTYmQe
YAf/xBRSxQJ5jOnFRD6z4vcojN8rzbexnPY47qstCN1KemOWcWtVLSz/EyHhWAKnuREO9YXqP4LN
Huz88CgpP9ZPOMwdOJ4BSDYk9OIzGWytRpkrujRIRBs6ZKamQzanc0DGVvV3zHV8R9TLZD9WZcqt
HdI2ELSAXghVHDouDAnmUk+VyXV+8qmMsJFl2/8Eu/ScpayekEyZLh0w5toFH89QnGVenUT847yF
ZNKmtmFMQuR56joHQsOHxXnb0wruFfqG6IbeY5yBigJIBbdzGMJYEGNIXVLXQBwpJT5/zbVQrly1
/OyJFZvwDNDJVk7PROKiZecmk/3jtw5ipIPB+J0e0/IcPJ+ruu9W1r5OfTDsYI+8aBFqZUrCww4b
I7FnDC1+3sgBXqqDUEvkIOIyGGS6Q/PU5t9VGGOHYtC4A03JuvZGY4FcaXSz8+pFSy/iDyY6dR/P
gGFZGl1d+Kg38nIsXh5wa2zXx7iMpFFeCj6nDuCCfi4ZEJBas+MuhqlaP8GaBI2IlJNvGZrS6lDu
uH/OivvPway0ZZ5iDyLUVaToX7/ye8FcgUITYmx4LpKCo8dJEk5D2a6blDEX5tfZBV5OwGcH2hMW
VtnQdiahF+h8mGvuSmqxjlspsn+7Hxx7QltSNSQzdy4o3MZMd+LQMg7Oyg4jgH8/d/7V1i/qAMj1
jpiOWpnxOnpeYFxkKjIewtEMJxeSRfelfLPBJzPWvNo7me8G5UOjynJ9NXhu0UfYbO5soyDYGdgM
1kH2i7TDP4OSkBNF2/cKk7ElYSBB0jybTza5VD0K8ARGwtdbcp4Lt7gM2f+0jA0qzO2TksmRcSzP
NadIrK7bgpOCnWNGAT3DxqfKHlsR06082NpfwdRSzdAoCZfmaakVrhnZfcb6RZCHyyApwjBHmcvn
uUHkgbZBHYypuco0tVFgCv1IongtjJPnpee/j/eJzVLDLp2MxxYrkLiile/x39kYpzPi4yFAdrBJ
pZm6h1Ro1mDeWXloMm+9sQkQIgqATntYONzmzsQEqW7J4lZzD9997m2mz8+Fyrbp3pp3vTNIjSEY
plrLSPfxdmdK3VwJFB7c1cbKy90sp5lW8h67fwSSA9jGfh2PeKUHSEobRwtcheg044FcjWrMpTl2
bguOk37GnjsW23dmYFZJVlUlJwXgX0pKEtd5UrRcldr+i0aJ5bWw2fXTOeNocEdJtxz6p5l79ILj
DGmHil6sf7wJ+KOzb4NIm0rUEDRK2YxnUJ/gzTd9LpUpBxfWyol7jrfmp52ogbcajFseo+8RDkM3
17GWgFWS3j0TmvNqbrZwanN6xkMwEO/Ke40WTS5+ebpxZ/vhpr+i/yExUdiNf/KkeGuJery6TuvU
4DZ9fpF+Q72NLFJmrg9n8ZRkqzBYqbpWN0Aa9TduQ6krVnRDg3syeMdjCEWbLjV6eXEQ8GCLW520
PNxQ9E9L9lAGtebwA+/9qHoO3NduMwW73FphBMY7INjyiItGdODPN6p7Gz02vp9/UaObloNlmPFa
Ck8C2GXI2i8+HcOFSHc9A6j8LRhbXxOhB5f7kcj2jvrxjgEVFsXn9OId+NKyK4uz5NdQNBfpQ/BD
ZYpdvh+0yiy4wwXbuGaL690zUQPd8/wmdWHzLbCD9zTT/YOgkIKFaTwA8KAhtYClQqllNPNjeRiD
IzpNZa/HlLplz3OqNMOo2bXliWnNWapDgF/16sikTIy2X9iWgfk0sqW3sZDfQGeUqMwVXdhTcdgQ
kQQwrs7n+ea5bP3eEFW5cHHoC0/k0A1u/8SJiCJQZ2RQiJqHZQtYnYgVtp5SWwDj47p3seIKwwXE
iwaHNjXDOR0ec+W4iSr07qzYY2VuOEZY/h05+czMgs0XCVBQ2jotzpCa/4yCtSFTIynfkGATC6Z5
swQ0bir33wZE8jBbSSpjUcPj0adv1oo8tvb2c0+kq7ExebeMdZpuU3FYHHWIUGmM9a75Jd+5mgz4
qyIPyrC9lkTm2Zj/UtOUxXS1HYk16acPLko4PGB2qT8s0BWLj5pc8oPjgrxJH5FCsvAYM29YrmIp
eWQaydGJVCi/EEXQZaGVp8HzH2HAPPzOdYO860PXK9NuaEFUDH71woK67BaxoPr0mOfAh0P/iyJp
J2Nth/7ULWbnue0eEQN+/NyGI8WbmvDuvdmJKcGxLk/EqGQHiTSi5MKv4v/9O2ztms/tBiCnpRHE
ux/z1DMhEDGFzJnR1qmvHw0YjpvHxioari79doyR4dQRBCn0HcDpgm0qsapJhYdhKMAOQjR+EP/Z
URdjNBfQKwQaaEeThX4XWvhO7ExYfLiQpqEh1eH7s2ssTu2kRtzsoWpyeWJgrAedqOecpQDAMBLy
OPJuUemh0jFzrKtHzuw5guSVXFMrlDeTjSk2RFFbZNiz6xJBp4oAKAvLnyLEWTz4p/Lk8m6oJlMa
SclcnydMT2XD4osBrlMCsLpDvzMGUXtATdFSGNLIkUJDAl6FKmi97J82eW9znN1aLvnj1OXwd0BP
huZ4k/76N1vGEXajufyGrGtcJxHvNcrne9E1tJM7TncBG840eWjraasMDiX+IAlzfOipnwcWL8Ab
np6fjmu5XbbDjyH16yzPISB+CQi3HCs7PYvYcptupK8vo3HaAoZrYrZ8EYmu/1u6JNldScGKUp2N
6E5fGw6whm5+QGw4X8MBYL6tREuebrCd5776OJxxV5eb3Kx23hiAwBZsQW7pXVZzicWY4Moz2WEF
GIMmR7ge922CATBwGmgl8sPJk/dScShucUXIuWt4BLLCYnYPNfzxJV/P/ubuhQOVXxJiG5SG4QUA
oLBQa3ZY2yE+Uu2t0h279Ze3htobJR0hg7wDVLnue0gLbC2U1YCuuDxf+TGnjMLiwv3L1aql7zgA
eRlutGn7xktXBl367YsAnUEZm0iwNHpdDzpxNKCTeC2dH2EYjxUFjGwvj7iMsbtxBNiuie0o33+b
7xk3BONbs0XZo7SHJRMT7Ya8JS1lidJ5bO3KFhcRw7Pv2iZ30Dl34pMIFzFHfRvdkcTyhlPm2EIb
m4WrB8Ep/7+ysCKt59OVDjDW+kdk9ICW1ZQ4jF2+4g87SuuoECSeEbgGY1FzaTHfKVl9Y62PJmeD
KY0p91lusg+WQpE7m6INcChG3J3ZtAqA1fx6h+2iQEwJbgUBTsY/AJFKuEhVjdhfOL6IcS9ci3V2
SijzpUilIGwdrQMNA9nBLfPEl9Do63T2gUyX/aAT9K7dJYqjQy6GI3D/T5NiPcUohpLGCcLFlx+A
fPCCaQ/OWEjQpI0zPZplmrUqCIuj5KDof7tJRwJY1BgzqUe9x8ZlLOR9CoG6WquaFyRhUq2EZVRn
2/cODSFOAzZ3ucdDDv4UJ/azPsGKPSIfET8IDpLjjcUpghEs754LMMXhd34D9t+wg0kxP0E5NeUk
c4iQmT6WhZxxBZFSA6MfxAyjr6AWb3AoQEIIGf1M5MGYFdSvBr31rs/O+uqcKOmCkEh7iF++nPyS
LyfL2CKsH7b8CyOlxAnVCzVLMUZr1GSx9KLwl/IPyeXNf1OeQ1W2Vh2aEyrJ5C9kYjWxN+5cWD62
ao+p4wI/31TC+DWo9feLzQp/tqqJtE2Xfwgw4HwEwK7diA2BItNivGJCYelL4k7ggm3sFpZpA9hY
Jqg4uKx+f+dp7snxm+c+NlVrQ+rDzdWh7xnC8VUnJZG12VlBzDiftpTv+GE7E8Y1cFP+zcXHyle0
cKp6sAK2TYFVYoSqlZMAJf6gbAdVuTvgR3cH+VB8v+Z6a3/HvtcobRlt70jc37j2ghc+hWPmXvja
ncRPz3lYS5Erx3sZoIWgKv+er+GqCU43vlrrcwj2X1TNg2kjaPScsZsBmEKVRcfg/qgu5z3r2i6V
FriI4d09duFout4NPmbw15cGuaJCu3v6M1TqNNhe36J0563ImXaj/fDfprb6cYMzTI17/CcuGhC5
CfwrHkZHdhoKqgXYMDnlPskZQrxQXNp3UoWOimunF4YFHPR9svsK+KK+l+xE+IMJV9PxpQa1zPMF
t0dNtkd8Cg4VXTLEnrQQVo74ge/ItmH4DU5aHVZ+PXJkTbs2IVtP3HKg5U0KYd3p0LkxtdLP0I/w
hCkiu3EoPj81WVr/6OgDT5Odi96ImZGkWvJQn6qgkoADB1ZIWlFDxS88Wd/TnEmck3/0d5/AQAUG
TDCohiMzyq8iFPk5Svtyt4oMHteW/4y6WRRDlBCxpOFrhU3hJxtvIf53MQ2GoGehT/umnbUk3x/+
o3G3ConsKgbCQgG7a5D9CyU78fBT/bUidhZHHWGHXFGd0iwhPVfAqRVut6Qt9BwU1vzSYDw215qd
BL08LavTOIEk2F/M9ZHaktsuCEzkS2NlDJ8FIDTp+1h2EA1bpPuC1uhGvJZydghNF/lvku0mCNo8
GEEDTtIeCju0vA1V2A779JwK58eF0tGS/PrPrVwnUcLtKcqoDRhqkwCUlEj62XHDJPNIBJDuU2TL
00VmezOnW6H1IPuxS030L6GD93RRCCbWfkQLtDfmMl/IFJmXfRTd60sufXcAnyhhwFkMB5y9mQac
QhsyI80Vd24CD0G4EMdGcKc54OotzuABSnhXi7GEny7KQhZAFmpIrgKvdLOM+o03kHa1DFrAKQ/9
srW821imtzaehD3MX3opqtqvcOuK+NpGJ8pLm52zx/32KUDiFYC1rEOif7fnvdQguPCCPM8jrWPU
Z06HNEcjvznnohhS1YA6EJKrPxRr0DEhsGnNNWRi2DFsuXwHLSbv+2GVInLieKAeUAznPN6CAUDc
Hlznykk4BERn8HH3YN8pvnDhLWUZJQWEAfB6bEpX05WZw7o+flvHDAkuSc/UifjIv8sYM/zO2Z+d
Ldypw/1rF1XUINmqVF9B0QBGmgzYzWlt2JUjleVjsNRlgSZE/rMZ0gq/570hUA4VI7KF5yBhhTuV
Sr/QCyNDtQBGN60Sm4RaiKpp+1SJ4xKtmhu1PDXAJYw907E3+TlFUUnctQlYfadsfH4CiPlfuzJE
GF5cbl+qXcs8hGY2qYsozlrs/CbLZB8ZYM2edNn7S4C3W1wJxMHrwL0AV9MRx0Q/pG3KGECOcHMW
OENZqmg58IZCaVO+zrjYp6UGxkWFwp+6hUHL852Rw7HGJ641w5sNChBSCy+fG/BqlTh37QHLAqzW
nkC0cMpizuwe10qGDdqJHJHqxqxGc8DJ9JUBS+kX05OsgIyxNSpIYKVge0eLJXpR8xOqVUsumkrz
l7iqyK1MxfN+Bj6tJW3B5qwXNNTLeuLZmi2oqrI9aXgwUJE42Fqea/pLS4p+HhHq9/VXBreDAT+M
PMb/cRn51GYO1wP+7/oUz+1IRMwe3M4axjuQLsBYMAMhjMYuQYTnnd8eNb8BzoL+WbIzhpl/kMGg
Bot2sMjknGgvOcudZt+/PlY5tyvdjCorLDqqSv8ctuIdyiw/DBdJced+EHUdmRDc4prChT2yTy0L
yChFp5/SaOYz4J43o7FxbEJ27/8jAntG84uGKhajywqik5j6xDpIj/DuRBudbue+D6bQKiRBzPty
wEzjDnBgvFWITV1LwaHhg1NHoaW9bP6hPuQSep7xiizIdhDaMMZqMtnz89W2oCXt3lD7M3EnyTir
6XNvHS2LcxtclfpiOrFcgODjJM1kCm8W8uHtw02C0vi8nrP61ebiaJysPIf/Xu3Yz3uaeskpqgWF
kvJf2YIVVP8N6Tuuicxrynn5XIxvK+hA6WkvDq5Naxy7UMPvthmkUnQkDnYH5X3F1F8CAQfVrSrP
wmVC2kZJr5VOgZvvampczlGhNN9stcUKcUkOWs+bfevWSx2NLdI30EnbeYkQd6IN/CZ1WvW49HHq
k+GuRF+8mRKiMRaix7BungY9x0pFctb4sfAijhmWdNQTAjrQNZYm/pN/gw4j7X81aieEGA/DeGIG
V6CsAt1N5PsszYEa3V8T3it08RIQYXlKuH6y2kyOibbUpvcmCgEYtqOXXbumMEZp4eOBbaVjxycq
Kcu+7aKxFWhIELRC/K1kW0x2l6Ojxyn+RZyx0oMa6aT/HAhXT1s8m87R26iwy9U5TvTLKrlH1gnW
NjE+drxBMk7lUMhc4DOawVWLNmfQpWTk1Hr4MpQ5fC2ft+AD54yc9J3MRwPoYNCG2HonlXvpSD7W
3q6T3DC1mYvE1Da+ECwU7ZWiGTyK9J5p1fwrbqmIcRERiE0YGLWy2AiUN3LEXUmT/HX1jcQFeMwR
GsOGyEbmzQzmz7dsrP9pJ/S0CxWPT9VF2rQO6DZDfEk/oRpKP8LZNOE6QoyDLT+q5XKWKHY3sDkQ
E2YuOfTLxdGD0RDwCVJu8sdL/9W8Eds6xikP/VeUoH6LSM2I2pt+LOE5x39b9ezOEu6fXucS33AN
3w2L7O4VGrAKX30ZfTTS4KmzjGtm588p0bzFlYEBiqMAHDkIs/xOXgjCK76PVpYk28SddTBb7JRa
jqbd3n4LhSp/O4QMvE78nnZkS7VPrLVcR57DvZ61T9gCz14JJ5ug7IcY8E4G0JvF96eNnJkLsN5Q
YnyzcUctr6ZIeQV4ovidyfipQwnKa7j4CDyJhYdlUEUAkTXL8wMZtSCnvh+IzLfBKJb83jAkWJuD
SKdRcJSkebF3RdRb5rVYInVR8cuFXOIUGyfSgzQB+kISAu10Bt1zJCtbbyH1S/W9WxsnW8dghZBk
IhoyxNdlLmgFsj9c8BmonmjmWDEURI3bxV4SDTa3eH6xbimJkYxrc5ivaoYWTVxW1/c9uTNdjpeN
UseCN46ZkRVMrXLdj2Q8r4kUKhUKY7XQUt9kYvhbozFKbgHUJP7YHR5hlQBulyN1WoXw+sCFvvVx
J189eY5C81TN5N9LpBgbcXgQ5okAsFIIMSMmvqhAneTAswNzmIkkgyvlcUsa/skemnyzyYBxmDVH
OLLzIRENy4iqnNHroG5mU3NwDbFzi4k1vt0IPBLuJJ2XVU8iedS1Vp/m5H02MEFYLdqj26KP/mtS
Nq3GEsw8umxZU+7o3kvatT/3tnm2r7eDv0mHYui0gj0V32Lo/0yEU1NEIMcThkiRLoJ/MWAAEAT/
KTgOb1IkkG1duWiEXwkTKyxdIv43lOKQ2191MiNYgkZlZHEz+gOaVJZkJ8DFWcQxIuhHcGd2cAoF
TKNUHYYNfZY2xECGhFmwSnr9YK+rn15EGs6DgPRKA659aHelnJ4Rbkt3oweMot3VpBUM15wkeZr0
9VcjhTWIQxkfBlUa1UeqNYwBWy4BFicXvo7dWcBy0BKJ0w0tGT6iUJ+3R/R9kqC3pw11MZSELQl5
xC0vMJozGtq4fbQCACof91ZgFzE4PPp6Qhs86AqqWgnSMoLQN+8wZSA4Nvcx1brgJ8FvTOVLh5Fo
pSnltN0WeWSZAlDCWm1q5e3reedJVRW91aGoerGXh5BNAX0ygXa2XF5qz27q8A0AqJXnQ/j+sd/4
5xcdXJIf5Wyun51I/LdFUv9HXz6b1VPBqWeZoG0UuD2qUppQld+M8MNetIdqPHAAmWDKQt4Q2PwT
PxSp3PqFNXOka0bbqIfIwjZSRMzkTggHiHOPrAFZGfEWA7tZX7YEOQ3BgW1WqOd64YTppeWHqZF7
7Xr8bf4qMwPnDKaxgX45hmgqjxVLtK5HROzczpLln3/RFB+36Yr9PMwQ/B63q+27o9nFhZJL9bMu
zI2UyMa7p6OtricBMUck7lVgQb9+gX7kizpr1sFATo5nMUJ7FlmnCCAtzD+Jx+3fR3TOhvA/iutg
IbtUqqYZS4yzcqGOFpQwk3YGaahmpCLTGFZmTZ0GvzdKp1pDJlK5kfrqedkX11ZGNCi6EeZZcGLP
A5GFBLMCwZUL9sIhIsE32Zww1+8imKXj5rrFZMd5mTTC9kejHI+36uTXlmUyedzx/8Te8MGdWahx
OxrmvoKyLRKmMK+Z6il3+mxNeQfrHvIoS57OuxwwlnuByNdbJT3sOurVFyoHDsdJHhyFxVvzttiC
p9/3LsbptJPWUWjgwpM6XMnJznT8pAXTb/SL8/EzoK7OHH3kY3lwXiOhlmbns6haE/rl0amCoCRD
0RQvvS+t2M5qRqbZqoji9qxl6f2wP/ZzhrsxVpHaPjhAHdrSTwJ77iZD0Tz2G3NAvzKHGsleqXEZ
Xz3ltvjWo/Ic3c5E3VAiNULQrtiN2YBbdrnrSDMh6jK71Bd3gDwtdKOe5pg3JJflx/4ZXSqf/MCG
fYWsA9+HaMy9a96zVIxNCm9y17xvHRDEa3VOG2xjUxQ6OcnDbfRmPFbDGtm0bXJGzfL/rhcFa0k3
faIVWLVZRBESgKtlKRCG1Tq9Qb60ka7Feh8hyEuakQYKvu9ueOVNvCu2qbnVe9Ra8+v0PzeRDEU0
hB/rFnphhBuK+bCKp+DSu7tj9XkLv7Z4rX0xxzFqFHm6czDX3ZYb7EpPY4ryZHLEY6m2xGkHoH7W
ejDDZcZNdJ4jZg+AyFjZd0xeAu0vWK6XcNsEp1isaJxsprelnGHakd/pp95XtB9ZMkALecVr3qwl
U1Rcis3JiRJOM0/lipYBedZLq7OZMIcp8gTpZPwvQOaoUXEv7s58MYjJvEUVkAWZMHSOCQtpmNYW
t+5AzrCU03EBKvDYSsBHrI+Zz/9Xa2hixfX/3olkTlu/nkh8Ll4BSk/47voBE2acomc4ff1FWHuZ
ZWpEp4cNRUtFV/YjG7aMG5zs4TU9EH0tUz3RFy1W3DtpNnAHn9HmpgctgQp9ypOaPSCvSfyzn/d8
bLcfT+RgSjU/Icmp/qqYnVTmh9+fu1LiJfuLdAAVtgsMMNqjURtIfB8WSk/57dYTzJridyCCsKBN
NXjE7GC8rcHSI6cfDiLzfZDae/vjuvNAzJCzbrf2FQTDzcYCZCTVuBkXlz09DjwokmA+Z5Yjl5Fs
1TQqyFbq6DpyhwT4jJWe26Y/dlJmXD5isqQMTXDrTkRsrKy/8qYNeo4fp/dyOdmjGvCxkV5uXYaN
k0Dy0Rn9PgimK7MWFH3BWiZdl4XSnX3jgHFU6o4RXX0LwxSMCRhUh9AJSJH3TKaANavYKwKdUTvP
Dq/m72VPlh10yKFZjH/EKvG+Mud+fsgbPt+O6AtRfe3myuhPUhGHxXE8dozQ/cA9WXhnK028jzJO
w4fzQgBlwN+5VNy6QPnRiIDhhDDuB6ejm2ycpnZ52GePYzIGjZjx3ZPIgspTXZk8uWm1PLdddfPm
XHXxUei17yr80pGbJT+ArrAgouGcDV+QU87ndl03NmAZS8WIDqCmTzhfK3XkcoU6j//cvdCYajLZ
2EZbeSRv9MHUYhXhcGJ0gibxRi9Y0ILoUOm5tRSmDXpNca/sW54pZMaS1IxIdgAAE2TzsICo73Bo
Co09Njt04EII57vUXzJDC9ZRyHfX9qszJQi3nPR51s7DSXUOMH2s8tNPvT237EwpFMwUs1Z9zsq/
a9B4OAec3Px4u6bluheDzL5ks67sG4vck9Xwg550HeyQgY2PabaIqQ8krEIZmwkspzLFNsblHSVD
k0O/X+6u5QgTdwTej6LjLWh9BMLfrzkK5W0vh2BMafdlJeVQxVmrbGYYeI+uA0hU9Z5kZn5+QUp7
45CWFmVXONS7M4yXzyT/J1Ir97Zwi9hsiI3r/h3JUiXDk8V+8SqMZbO2sDVEHQ8ni2lKD91/eY8k
3VlnC8wvNeSuqUpJ9k2VrqD7vHuEuiHwVjaH4XeCfUN98NDdTpviLlYLpWHk8/2Nj/lBnLiCK8O7
LmHe+X7iG3SLwAcNgVsSV8z+k+moZ/Wy679hWzDCzpwdGlExxJOPaJX6m7VbKzOJ+jCka5TuZj33
SWenRg/mog5UZ2RldMmmxOFZGbkpZfFettdd3JcLfVToc+FsQA+qiehe2Y3n0wIUzsldyyLS3Uvn
T3EABNGWjOiJqLGjjSmy6d0Yyxwxykdhv6knFKukRUwvJzcYQvue8/MYRJ53MXaL/gz78u2w3wTi
HQtfczgf79ZEottCCCynQvrv8J98ZrZXWlIUEDCoCjhWZ3tpSM9lY0PKq6I7R6pEfFxkGQb3cS6x
seArEyNQtc2WcArNpnz8U2WLlhbYRL2P94khgm7Qr2+jQ2/kaAEblVusGoS9bw+MxkDCmUzDn65p
AxO/NFrCEfxl7YJo0GFJhZXGkO8KlG9Zcefoxpu38tB5qq4oKj0c+tjlxnabXivV+DIaXKHMJ1lh
Ss/jmW1GCQGA2cHcTJSSD6O0FcIrkvEV4XQ7+iHcOb0Nasw0wB1w9bawMPmfcAGxh77RiWPCtktS
HODyYOdhdKsdQrPlcVBbQJXWXwngmJgHJNE5F3591e/N97qiERVCAyzHdGE+BF/JaipGBQzmnxlA
PsUW4sHmVIrQbCZUilkQwjgc0m83/z4PEhSLONqrS3iMdwvYqT+4/5uztU+A2Jf8J8Q246XVBD/i
SrjV37IrKrJ6T1Sl2FGpGwgIy68kzluv8cI0rExEYPm7Sjm1cPdb3UclkqUnx07o+cUsu5X4Up8m
T/zwdRcSj3+Dx7L7ML/Sq9vZ1gzadzAev+bBK7U2uQjm8VyWJ3eRLUM2RrCx5ZJY2cLnFMGxzFFa
xLX9RAu2yei2V3/Vu4zBBAsz7t6EMWe0H0kOJEoxueoBT+rleeonqGe2aeTBHKR7pFbqnhva3jvb
R26LqWNBehRnG4bYh2kAqdaT353NUz1o5dsXAWZyDc13VFQj+Qcw3DwJjZPuJtXIMM6LTSyQBRot
Uv0l2OHqSdUHRTI0jFbvNjb8Hy0RhBNXtINbjNbDY2SzJQijzGunlQ7DE2C4EwjwPzgRvne+2gXn
mr4w+8VAbs1dnfvUMBV6p02DpxWXqHOq18UMDjzKXxiy5SFG42nh2fBIoJ0De7A2IzFG7uu6lJiw
s8888xp3Jj91Se7dvISYVdRgxwAWxx6iq4YvZgbMeMcFgYAwqqhJ+0adChvEQTr02G9rHXvuTp0C
w4IMkddFV9f6Zc+uKDueQOTcBWfPRgZ+tmxi/xpRDTC/IjtC9RkCxJhai0k8g8aFy/itMPIXFjrS
6YhRWcw9EjxoF0NHAft2fJRNni9bbz+KglDu0ruzt67JXejk6uWwFxG5TCxltMNjnbYd+LVh7EzY
hmJnq+ZO5OJKwrZz4kMqup6c1auCpMR5//BeNXTs0nvcNbUMsecLbsRw1QvKwhGgu6EDVAGzk95F
MqHdzESLHGVBmV6/HGXYUcbq2ioEhWrZJbY0syJdWJCFgCfnW4s7/FBH35JksMb3eOON6YyVrQFa
zJ8P/9+gHocm2sR95fsthoPcVmR6+7OzCpTeF/CqmGbuL0XGZiPcKly3tdrRhmBwh/ZAbhRSbE7g
srQDMD5dz0kcCg54bgcy42xM004vQhxVfHWkTrARXNNlQAhNJ9ww3c5PC8a2c76G1B8VowHIoo5R
OxryD11Uh2neEEpMvUpiuP0ydtsYv4PfS6I0idxQ25GgLY0L9PbvdjSCtyKVzHfHZ7bRIy8Zar1V
nOv6Hz2wKuJcl4/O2ZoTqZC8UFokBS2FaBEmVGXW3QXrgCEGCHWypS1E6zflIPd5n8KoidlAsxH3
37ZCUwidvpJG/1V4pTtZ3oxFTcpdK8z4k6ZZ0l9wL+BREtmlnK17LR6dFwMo6LSi+uIEYDoYINJb
LeociHeyKOTwOlbi8Ug4jySMddWSJn2jrX30a+7KX94FNk2PnLxiTFDmd9U34I2EeqF3KHXvuEU+
gfPDAL67Wq3EJAcE0pgDbwbgnGaMuCrPfs8sR4iomyEdDIdVgm32FzaHa7xxhSPbhFhP+V3ixNZ6
v1MB+MYhUt/omW1DyCWIKIcL4jY+dkXs0fEdlDx4dgOXDKW7tf1rVp9/Jr1uYo0gEw4des8IKrKN
hUylw/HSWDKxMKLo0FVcMKJVqhldjokAanFBKIFnwNhfkHtxW7rvuRITMsnTFjao6Sta4Dy2J/iN
/XDBR/ausSsjXRgKH5PQG68U8ICSrVjhxjS7Vfxq3nNpowZ7Lc3dCPRAkW+AzLzP9P3licy64zmo
/kCLKdn0y8YPjw2ZkzSglwBWgJji3WiB8tfszOZejjAaQXLx+4oKqnOkz8hMz6UFB3ZjumOz5QbQ
lcd3ibrUz63OEKrNnuz3dATpsiEBkOneqAW6ZmOEuciDzV23IQRN24V1ifvX3+X05dvtUy04Qpby
DodX5UeZrTo+tlpm/KMR4E7xp+OuYHZnjuF8Hbaaa7xeuQpix7DtA5U6ihtmWpLYF7frNI+Xns+V
xwpeX9huG92Qhm3Lt9kN6PzNF1O5Wi1C9D/3vloWpT/hQtHzk3ZkJJXVmA5ZysM/MldapK0VvZKO
jVqs8qaLoPlIfH/dhfHnyu0uNSPvg1qDCrM+qqJgXVWTyIEv4MDOFe2xoHBNUApVfcgPIblesl6r
aQpRha6+rX7brJZkGGRC3rFRn6oZNvqufAoIaRoZXmI9bkohycEIae6UGQhihwn9W1B1wmtpQmPl
7UGkxLhmMv2znXtAoltQZjCaAzYKO0rX8pF/9VW8MvSvt88oMdE6wRaj59RaOPeVHwpoApLYFHPZ
nA7/lvg9J/IixycgE53JL/tLMmlYJTn8URh5uS5YGkoduIQSKlC+WXreZiDNNpZlxZNI79FhOdsg
SFn9gFB0acKn8hV2Ik1pWF/YmqzbXz7S4xxY2uey8AY/wO0VYIU55iTLvsQvnCDjVMM0j6wKs0Gs
FjkLqmxtvoqCJiJoMV53dnQeaVfNLEbrEUkOpDAXshMb2Vgx5gV//W2LHDbHVnID6ITc8duIrmHw
EAbDdXGamoc0/QKf+lPIQLc60yyRKWgqC1nCzZ45wh35GrWWf7J0VD16fR19Z3PmhfHuhGwZq1qh
WV62D8UHNLD5LwDYGrjuzKXZyt/CPa616zvDHuoyWHfijXmoeLLqU64eTA38NKt/+iWLeelzMYuh
pdm5g0vzPIH2QnherN1JgO8PQez2swWkv3AJHoFBBmOvU1/zHFtuOUx5IeBdW7myjKAHWpHNKUiE
KWqWkucJ4yivS4H2khLlhHzmnL+oL7tZDUK9C61H12DyCLxr0KmMsrkWOxyG8Y9hzL9/kljv4oWw
gQD4LR9IuCUO8IxL/OyQOVV3IkKQO2HJs67dT7WVi+Dtnud0eFd+tisMsygTrduk5AtWKLL1EtKm
CYW6JPz7hDVUWrg54DdgCOh9GeW68Ld1IFsxwbu9oS1K/6IXluLt6paZN95wUq3paL5ExXoFj624
50QiR+EsxxmvwCH/fS8IGWVRh7WtHYgiibgbOHe2EvP5jqGYKgYvVWeZY803s6AXnuARypNKCuK8
+81dbVkjPK6YtHnqshHzwVcgGT3247drIDSBnKCeZdkjKLBtD5VabJ4Ag9cU+ReFI2CubrRYH7+2
auRJzkDsb4Bwyz36lA9UYpOAkYrdDz3OlJrJUpDCX8ZUW9KENYlYyBvGSVkhG1fbGwCMEum0n9gB
OUdAA7h9RvX9Ys0rr1bKk/VQ+qbxG/ULeLGCWXIlmor9IoyFaFA4O3rrXPrBq55n96IVD7S2ZV4f
UDYri+NwvNBJzRhcHEKur4WkeFcicWzF+hMOe+mcZWK+DzKWsM9gK86uQ9DT9Uk3TPyPKUfFbijR
qI726zbKGOttCA1/osBMz2xd3KaMMXPiQlkJs+QCLxGR6kOXFGJZkJDDDg9mNQK0Zxa4pY+k4/Df
rxNhqJl8yYkFZouOHHoIuzIik1Dj/Q7QRGOuhAmXA7INM5IPyVhWflFAbsgxtSiiT78xosFsdibg
rBRsTTlKvNJ7AQ/bnZvUZPlPeNGjq0+wE6qAzGFBkq5a3Uy80GiCnRbtCXFBkoYngDUa6jaqVh3I
SPyqiH9fjX9IKjztygsr6bPeXakZoRMn6mYe40pLeUqtbwQhtKkYRcplsR9mtr91wlS8wQEhJK+9
DgUZ+jpDMLyhdU8u2CEAu1bLyJK0j9ljWCIuUrKWJM17KxyXCU3Yp6xPhNNUb02Wf+Q7ZaxktJgq
h+QS7AeyZBNLGuKPOb8CLpCnOHlMNmVqUcRcYVIA2JK8+Xzvsn7QxzqD/1JpNM1p8kLggsr1a+zv
OCWy+4R4YKLSRIt63xb27ZxFj+YCFA7DmwCBXXS4LxC+j1wUY43mHHzvp3gZgfoC65EAiviuGFe0
4bFOvibmhQmvsPrsCJIxZUSJyrA2FqFjLPkuy+4ImYnScNZMUpnvfHAHR9g06QmhZPwKElwQYB93
sHZFgeken/ETnCl9nVHPcLTAypIeTTzQck8tiL7zj1QLY2HJsG21g/+VWnUh0rNVKcvHMSIYbI/O
B6pftst6KkXR9u50/4Pn8jMgMiZhA7ws4O5k777xKWssJ2W6YjbcEl8gjjvYsQd72NEBHY9Mh3I4
SOKFgX8pDkJaReM2Z6UzPjuqK+lOhLVul+lwZ4zdgM9kRw7+aWMyK/HY5qIkgA7ydKtP0598iyxi
rzD1L4YaN8A2vx5LtulDF6Eg6C1+0VmacBEMdj4lNeCYjY5molctGyZUlhlM5MpKnsyJZsSHNkG9
XzsyxdC5hlzPkJzc3pNBIBwsVV90S2VDX7srvsB9i+xj1jTkqiI4iaA6P4/APUfA3gp/jkXETgQi
7rLEaCFYRsjJwVWWQAmQZ+QCJYcyrqcduR1OmF4iFAgv3bmfv3/jdlUTQX5e6xcJ5CMI2p80F0mR
gFACITASQ6hMIGYLKQKaiFXKYewlaJVZv3Z/PlTv+i/BBJ8HDHKu+RE5hPjD+AqL21KOV06rjQeX
iVMQX3afjvttUrW6IzhZY3NkcfTlzHlHKZozB4ChIHow3tjOvS7/qQndtKNdPVzCYznmpO9eyO2R
iDM2eLRlkUvqr42E3wzMzJRcVjNKLfO5ZJaFhMP2oXlvZj3m7iCsJGJZXYKIclAroZkFmZ2uGWW5
WqFJF5whkTfsPNMAjmQUyZgZ09/UK+HGyPa36xU7e4ZxETD5scdqptC+nmc1hUE/mBLERN0+Dhgg
a1MJWgIuTyPrvKonqwT0GXPhNM4m3DzlXirLIUx4R/4O8/Ug8y6rPlOHQiX7DceJNMC2f4Op8JuD
DjIsyNJ9ZsmOhoJG1tpWQA0rguna52v9i7gShuh5BDIzAC+udVoxYIM0+0m3TnXnJeSuz1pnKRB1
6yrA//+zG0j0hObW6EuYnTnPzJc6IrAuothBVmky6OX7OdWFgYFxHVicrt0dMR9Xx8LBzvhvZh6b
vAtm/cg2w3Xi9MpCwo1fETOX0M4GR6iRFhCk3iDwg0KSIS1FFpNY809EGdmpKE0ly5Mek6jdQFZI
C/KSUimG2uGD+rlgItbMyYRANRX7lmMBUkVn1+0D3KTNDwbgTIm/WFogSKd0xxRFleVLwGsV3E9s
9W8LPSzcSN1aEiFdkyRKqngal4cGf7v69k1VpRtk9vhsi9gd7O99kl7hXP7DBe4zZfXNbYjXGlx9
ie2otxLqcnAPY8HRqn4QfL9alZ6KlMkVup3EPRngYeIyfqMW9JOVh0VCK1K30JDFdCUkVzRTxpYp
O3kW4TTBQ8YNPRwsPqZQUeSRo9CK0fSuAKapV9GapUa4fS6vQ7KYiCVPELoiDwe8WBLs0eiNi502
UUytrbPY142nnvdHinDQKbjIGRsmfjyiVFQGxMnUbEEFeh+ZkKBsT0i3shrs49spd5bOyKrbOVLj
ISaFNa7XIEojFIRrgDG87pIx5u8I4rFj2j1f+js/7Ue3cl97A4TbX6JafwbrZCgYrQt0fUjh1Qls
98CUW49q7PZa0qonwE+Txx+g25nSqXoe7Wphh82Lv8QVlEy6JUspCFXSkB82GC4i0y6mIea3NupA
Yx7lIQSuBJlthdXp7ZbW+hYztM/T/OIH4sGtw9RsbwgACzMbsWUwUYi/L16d5hfSfXmJ1ASdYNOw
yRoJGl5q0pNqjsDsIHwl2kdUCAp2U8b9xXisX13c+KLD2DIexuTv+Cu34YNekEcyCNqXLYum5dYj
wNqIA//dG74xh2F9Mw97xPIeKSicRdsJIYCgrr1EyB9ERhOa48kdFRCxq8suMFYiC/bw1fGfsjU3
Mi2Qo5WgF5NWnUdxiMCd2GzVTW91bcWjx8Qn54Q51dXOZSWMR3DZY/DLJOCczw/6SMFolyk/+zw6
ufVEgeqpDFSEE2HcgSz4nEvB/F2Lp57AWM2uUOD7Hgc5YhPrFV/hztUQcCWaFBtoO3oBh456vX+3
51vXppgMiLH2iJc8YIrm30vwMriL6VZ9qWpjsOt3wq5zkatjaudDya0QFdTE2VHpBXPwKkmRTI/W
TftdE/PDnE5esJLPztoQp7AVaon8BqOWLlONbnuT4oPKMzcacPY9O5SXcXl9QiQmLOT/eQ5OZGd5
qBO9YSdueXNUWFkHndixY2r6V1/gRGE2PIZbLOwfimYBaWa2N3ZWfBWuuesIQg+/pxBxAT8RO4UD
EFeyUDPew2kADowT3IdjR32C5sy9fs1Jzv/I9Jd6CgD9k/cOpk3qOuFJJjGKDSLu0523inhLjV/D
/6IiKft2/aRgv7mBjfRbaNKrfx1bJifc0JFJNqBMTaVCBBHySXWuv8OTYq01ncWsyOSRV70vMDSh
hfZUNqz8UC32iQCIeeWZftjRJmJOWaeCqkGtqlW6nW3vSwIhLPrxhya3s4PrNT4Ouvnl3Q4PoQOq
UoEWMlp1Fw/jEmPU7nz8LdRWmgbu8S7OgW+2hrYydVHYUD93fU+YtoQzO4zhGqKxixI96vnucG4s
VxLfxPWGgdsDREoPYaebkTROtc1aM6iJGf1gOvOUlxJR938AVim+p2lfzNJy7AYZ2ursuNco8b43
65hExnjAlId64zYfX1vaQJZW6PCZwtuFDE6A2KZPPLTRie+0vSvIEyDywAYT4yc9YDcaSmk6j7qI
UHrsWLnXOp4UdapgAd8F1kxNVBVgKb0rXmz0s+qeZ+aVFo8ANMCtHygqlk3DcY6+PDPqHfep2eeC
IDUSPzi+yKTxXfe7xFZ9sNol2mMWKFq9RkTvr3+8on+FpgiTsJMqcfVKHt9kZeROUzZutbE8CxHP
GZNC4UZLuse8Ju6ONNq672Q0yczCMOXddOj00aBgLW/F+hA5bmOhDGOkABgm7QOF+YqYiRLpvm3U
wdDnVDGMxM/c7uUBgczR6fcvQTSaNz6LU1BxqT3MfwBGnjZerhtdBa7toTToUqgQu9OFXFIuKKlJ
WKBfEuc9Dt3uKKmhx/wtMwFhXg1diiFjLkhsYxz91kP+V/m29KZNHq7MfTdNyTeEBvr19kFA5Feg
RegOKW9MquzbBUqoSBbcx0Z2DY0AsdO5UU/YXBSxIei1p7sMkUpEty5kTNwO5vtvydVysQLe72Vc
z6PtB+CYJ/FKyrdK/KQqA12eCEMq6iMUeBDSvjCZLRYSFm7GsefztIu9Bq0qNO4MiaB0DcPPZw/N
w35X5sQayHQ7skPVMgPfQgAyerSHxtxJhLmn+28n8+85lbiEyqKtXgO4yDGaV5+QyYquqILeRnBk
hrL4qLqhI8N7xPJdsiPZKMW5IaABHYHGHz6JG5jcJkTkA2dA8MCfKUq3cwGj04F8X9hOVMXo+pwJ
7yjQPULqIgfuznJ2EFGQ9msnkF6GHbZIqbksZCoEhSTIofkKuht5CicYKLR+qzy/WPlr0LXQ1LWN
jwBEvlIaBzli6Re7oP9ZaXcEYOoaEGX4tcBnSn/15RfS/+vY0kMwret/I5bSf8P5ODVQ0wdEZrWa
ZQ4ap/oCNm5GOVGo/l8k7/z5QIPO54PLvsms1UNBkDq3ptMT8ZhaAlCa28ss/LcWm9go+BeYxhp4
wgdXFYobLKqmhmqC98IFBNqrKpMgV1PvbfQLyonWpymEhpKtJ06PcyLfqOMTTJ8g71siwrG7/e0X
QHPsCuSxgdycnzzr/iy+9/8bNhgk2h+g91n0rEUZRdZ8C55UijRuBvoTmBCS1yefD6+TyFps34nZ
NTFaJxSD3qwWSzb6r5g9ipEGqxVgyQVN5Lbw8gjnXLZyVOAceoCihh96HVe9RdePD+PUPqp19Pv8
75Yfj94v1UllqxS4kAAwqkhwqzSS6zszCHf8Je1XiFOjrRTVA0j5swqXrY9zjP/zzOkQgbbk04Jl
OMf3v+1G9ZYs6egvU6HbswewTYhKzfJvbbhG/ky+XyA3YmC6dSOx1PyUM3ZvEawzFA+MZxPF39DD
i13oU11YG/mSdR/iNpFdPtHup0PYGbgbCpELurDJV0UNlc1JuIy7HSvmodlDrjQpQCWJirdMPO3i
Cv456T5s1afH7X1iaYg3wEE+gj0Rcp5nYfkDpvVEO60ZeVBuvczbipNop5aNoUie1jFa2gb36z3Z
x1Cg+e3ppVY2ihEeHDHMLubAE1a73bS6/9FcGQ4hvXjjBTA/dvkDW7fsdY7+Gcf87uL52o0Kc/yp
PazJ8I0ETUE9+AXimQcXj99kcXKzgiH33YT1RB+rl58SnLOaPn142ikOu/sqMl9u1dqm6tJluQkg
yvw1mre2SDY6CQ1TL3cYWctyosMoW9++HkG8MVFeWnD10LHGoBhYoYyoH+nKPV0oh36wgdYSh+A1
yJCvuLfcsp3bfj7uYX+vEqoXfADw4p8JRVV/T0ocsXenjzlAh58O41o65ByMX7gN20ahyzY0sxcJ
64bNMjaEONEgxvI6BTlbNtTyT9e31Lxvt5pISMf5Sb48wxatDJ20brkTc42h9cMgUPRwfkJEQO+q
orZUMbDQTZvqOI9m2XTtxDdJd+Yg11W5USesiFS3UUYOZINy1kaIUXZT2uXC9pTPhYnN4L+dKtCf
kNzR+fQhOFfnnldS/+iXGzuDeu5VKdshslV+vpnRwHLs+3/4Ug5a6MtyVoDBGF6cxBwdYa/ouBem
Hop5h0vXQHv12KPgrOJUnIPsu1njkC4nhJZFIhWYdTCKuTcHAA9hmIOJHiH0QlaCX/VYmD3tQhRt
gydX+qhWxsppbYIFXSn/oV0mTU7+FzhrCMs6F+AIYnoe0lBHLV1V6RE309zCd6A6Vp/LPDpu9r+v
m95A4pdwTs1LRA0rC1x85WI3NYM9wOhr4QkjsDXp7XeSxKSgsXLU+WEa6CSu5GBaqWJDP60Euyhs
vhqx7txcGev4XF7PxnXmJnjStsTo1jZpip/jq5nGOhLWaM2C8goXdfj9EzdiP6STR/s9xFxYXGky
D38S5b1wuj1qtu/oHMnwGJK+H0Z8XmtVb0vsno3HmHht1urUgdr20jUuXGJjx8Z9CmKpyYStpVfy
DoSpt7LOmoRohSrMII2jFMOHesMctXw0K+UzixN2upMNupTiWOcrWGiiCmoePGVtiRPDEU9Cgxm2
532ysmcIdiRpqQvrOXqmF2o7AEgOtG0mnqfXLHO/UTYKff/xMtQDOh/lKu6Coe1pbLBUIad8EY6S
hBLI5d3hGb73mc3pcoqaS6QAcoPwJyNpxRNHpFTnI6mwZSyAaq819qprXAguzaPSEKm1IcxyGwPp
xRw5eLqu8Rt+iwHohq4ZAUx6wF4khyzNWVN9gPdtPynsJ2dLLu9SUR0qtcIzcqt1yRXB5BFLFWU4
qZ78ZJs7G+vdjtxXJG5I0Af84B32/IY1d3Fg+epmUZp+n9WsYmj+GjSOFoh/ul65W6z/MdpUyIth
rvidNxCrGen6Tmub8RKBmt7E2NOZ/m+5rqxNJSa9+2PETRIo0pGvEt/8voVh6zyfycPVdx8y9pYe
BmhVAiUi8jhmBXjeUnsvCw/acTJ9ys/ZYdVR29Tb/2uYa8oJAOzLVQlaB4179rb9yy8lhW0uHJ3E
RnAW08OJtVX9CzPlXPWGpDdb4K8Nai3wVhQPRpSQXLKQLhFjaMSpke2OITf5b8liaLy8POERCj6D
IyaSreb441aCMWIPCOCZEhb3cDticw6/c0C2NFdbyRujyiIOpdgORZWxBeo3KuvoqAyPgByavCPt
HSUHffWO4JEZGqARvGlZ8gXvWeMYGNJ7YjCF4Hie7J0fKbZikBSaGh6tG1AoQ4z/gvKnIkijpYYE
DE6/uxzDwf8HunRMArk6gG76tL2Okt+B19XZQbYrh5jFDSoopGskuVductKTaMGfXYEVYusA5cyG
4M78qaPCjksXC/V/6p6tMNHqZ+kXfA49rLxdfE0VKcKz+mRrBimggYr407pXLT8acO5Ron047FGJ
EifQaIu5M4qZQ9rIH0xpbVk34UR6NQtFyYxsChXae+qFYY4dElOcwtW8hOSGubWP9ibmVgXznyzg
gAuWs1Q+9jk+hGX46Ze3Lggy9jFBjzD8kILlgAeW1XiO8e7uugKYe4AtJ1PYX9N/j6tphd99q4E5
iB3g/8xXFZO5Cyi0s2EKG2+NRLvUcBd0UC4S41i0wt7dnqoPi7Ia7ldIZsd4oeYMu7QC/s/wR99D
Khy/pHx7qyW4dvVItGolRNTZg2OXkKNlZwWepokTkF1VFHPy5Fq0sygpl+0GpFAf3Nyc+R+GDRn9
Q+5UaWDdTm1pnVGBVmSjzKp2VpniGIJvar14rkd1m2E6dxxGKrbXNthZ4Q+MT9RbMNhGvf4g+zlh
bWht1zgKsTHrug4CrGVC4COmCF1VVDUYihinRtJwsVY9hZsE9sODBf07190QmW788xRQfZwzRo08
64tOd+jHQVe4BgjEPydnWHGWfCNt65QMK1Ns16Bm+k8GbAB7XjzjrbsA6cda7SKuFrgw6nn7wCfC
3hISMg0pHpHxcY11yXJMMm+rtL7wXWXfKg0xTyhlFkdCPAXXgfKpEr+Yl14NM77BxoidYmV2yOLI
EJ3mph9nBJf0T6JWxBmlMsIT56dIyd86wFbV4tOMChSns8LYlfRgiW+d2hOP/g20prOhxg+e8bIE
Cd/rMvL8DFI4dt/ZcsBqM1xriJUxdvjc6y9MRXYDF/jzU43yEO8yusdar5OH4o2Yk9oJeLW8YeTg
CLzf0usXcINy5hGBYaWjkYKUDYoX9aUwbdfAR22txccIrXYEKeiWl4TKZBKeAW8lRapILCa24jtb
lQZTIgEHeFXZG30VUcSjQSZzxV/nIbJ/IfsnLOfzmWeYab+kjJdX7VMcEhLjejKsEYUtPPUxaDkW
TZAHBUWCcMSwpsc5FtoWGOZ/SsHpoRZbyVh28BAZ/cBiR4tyuw91bEAtHT7QdUuZGhjIfMVxra8R
r6K3GNk39unPgimc9zGsvz58Y1McJ82LrGcPoslRgHLQdAZtGw18QquuUeWwN51gYKOm7OdX7xuH
8i6BbEcDcU7j5+rX8T7gK4ptBLqUWTUamyMiO6QVrWMPr2AGgmnePs45Rab4Yxfjtq9KiT9qqMBc
0viw4Higmc8a4FzhOKrKWf36W0FIC8s8sMcQj6PMqUt6CO2346Ev8F3m1CnYQMY7afOanK8Us7hq
1bUmTIFxnmd3yGIY7hyoB8Cv4jP0J7uSRUUNKbb88U8VFbLKIa8L8PFFctAtkFyGnXm3nVtMdJbF
lURDHbwPcGSWl3folehwemg/JRWXgZPXI0zoQOKFlORWbKHdUlgs5etb0M6OYFJaLA/goWrFf9Z8
DRl8fEGDEpTWjQVt4ogLqHDikaUGbtMxrRgsNc1DCUGASPYdruJfrZQX7kKWBdNVQZ557tP/x4om
MRhHpaVEvgJnvMamw1LZIVxQECyWh4oGcd9nuMP4lxPCvDM3c+f3KGl9rIC5ZDTg1nhdjHivx8cT
XqcQA7EI9ZJEZcMpTDmB1t40bA6Cn9bTqbeKLx3vkUn70FjlvvI9Y6GjLZHoM4JWpNNAFHHiB/nO
vDAU3vvpkpmys1oO79nVYTeGgvyHEBJeeYBJNAPG7KDAEEjcTi+fSw1+YfkukT4DOljCyLGhmt2z
JGGiO5BLLJkO0oXGk9bZRac44NTcXwFyFwe352xxY2CU7Un6zTrDt8oejZ2Wxco1DbFWKzBbUylO
ade03AM4XTwcThNuBwMjexi0A9/mAaQ494uNZV3tCcePzVSJiNx7ke7iQK6IAIIkiNm6ip6WjgDd
X6PemjOZ89rtIh3uFxrRPD+sb7xax83OIF1dz8zSEl2CaZuzUz6GAgY2xiI9N2Q/nk7Sr4+Rz5xz
qK36AfMSMCMB9RuYm0sik+hq+69E8d1QKJY0OrRvy36Xabnps/S2z0W/Q9oQQxakwu9LyWEhLsM2
b5tNRao2U63EixCPd33DVRXYPBXxTWGSCtNYxWUE5Az7Eoc37nBOb+XL1Ba9Uiafg7T/4nJXMbNu
GzC0ev8T6cztb9ErYATziI/m6imoCCaBLxzhQT5J81kYfNlLZfOGEaWpEZ5Yz608PXO4xoD2eXsJ
ETX+1SmPF6d7YpEkLpqqQf7iTASBluxkEy3JrClc2IUdG639TIU6MOnMAb85Dd32m2XbuvgxGUHD
duGv76B5aR7OV+vYgSMEI2sAMRcwL6woGMwXVpP9QkStSGJMR+ADNmAnM11lPMMTXG7qKUlE1h90
m6FJoNA11F8F6XLOaMQNMNt2KSdpbv7WHptp4lVWeMfkwDJOJ0S9FT86YF/0ykUn1kujo0Xn3u7C
+0jDA7e/TpS6Ols7C22JzuWaqhtuZpNAMxjLguKpi0CDKt1Y2UDBxcUDaso0o4fbeNiL0+gpF2HB
6N141Qv/BSUPzq7fBIGpG8/eTluboJhjHL15rGBNnEcWDx9dQvBalcM4GLSL9TYj+5WjaJJMkvBu
g9Q87hoSl5jbP8g0tSWiJLSfDl2f3KvoL9e43eY0UMpVLyF+ZP7MhoOOYg6p3yHOWRW04eI5ohoz
Ba6vW9k9TrtZbjGlaqQmRq/V22PbuMJtD6zMLEQvuHUOhCPAQs0FshC3UErxAgwqtlrPMpBdDbTr
IxeXEjWVXHeH5FfES0x6PIXijRMX7hPbaO3o3XkdNnz2wj6mVRjEj2pVF1/qEBbeaXJ0MXL1k/3R
a67B9FqBAwNRnf+XPvps7q69vbwp5usF5tHHWE2aGKvd25acjaegafcBgp5jzqnkolkQopEcuC5A
aG9wDpABWztOSTVI21tD8jB+gpaMECzVga/dBLVe6IrUc+SxfiJvtKTGGdgPhbN+YX8lmnbW7pSP
63lr8Eah1zeeuxcXgDtKKcRIVTu43ItDpc7BRNEaNRBYuXJwWvD9VLH+4V0KZh1k5CsN+yt4EKTL
nSJ83FgZjPnHvC+a+iBT5cPFW/bXic6V3793zEEBqO3NWKs+nGyfLSgim06d4JZkqllSj4tRcR+k
uLUXj0aGv88b3tfuRqqWB4ndWqvgOlhdlPFC9CWQMPK6sficDb4k2cTbR7BeYq9beWMmRpx5VZNb
a82TQR8/ZKvDPSZ2j2Z0+HTa68Erwbocg/M7MzkDCJCV2RW8sSDX4ZP1zL/WBP7Nk2vCbaQZIMsq
DINc2Ft1dkYor8JJRR39MDJIuJohjxYsayeo3I1eTgNnGpPVD2wpe5p30zGVJn7bwtvUjHbhk4Di
ymvgjhBt6H5YZIunESHvJSfaOQZuc9ZFH7nPiQ9kTUbMoGQwFIF/zfVIPSaFYadNjSByhyJZcOw8
ZrLhd/Fr3iEcdYL4br5qEsZXwxvWvfhvD2oQ8iaklLCPSBaQxR51h5gxL2rjG2tulWOujT9FvijZ
5lmVL6qFg/H9CtmoikNvrtYmxhzHIb4I8Ph2roUQicKP9csgNbYdTXpl1aBzo2yjCQAnyTnd6G8a
fnTLrSQByYcOHGTHAaFK/1gJezzHSXzagsPbe5qNm7/fMHdgqxBh5uth8i7zmvNZtI/q4uoLNbuN
thSCvaFr67uLawOIJe0Zm17dG0yf+3CqOh0JMYsRu258dBkdtISBJ4NABJX+rrILmzS7Bf1W/nuI
OXVMeKmxIwCMvxpIMXVUI/Ucyhz+E2GCMkQIDEK0RC3mFS7HlV0SmzcHAxJYBWgnv84JEfFh/WQt
IGaaO7zJ+c19v4fV0RjZrdji62fpCUEeU+NpyRxGz8Mxb6eWnZgmMIF/Oq1y0ILqbhZVZAcmMpXA
CPSD1evi7oq2S375d9gIkUVuMu+/7TczK8HuozDIwSR7qlHSWhmH5JZW4zanVWYBRO82eoDzcCx4
jOZGuT7TitTXqDpuSx6yviUaVj9sxgfH26uqvKq6iH/Pvvkla1fQ+9c+bCLSqsSSzSUNvkRSCXQL
H3wEMXCasHbKCORviEfDePb5T5KTE3znL17binLTu/fh6fVgJEbmp3ewcG/UO1SA9u4jKYKsCNji
C02lEZlxCrKtSRGFT/e90RFnut5D2z+GMB41DghUCH2RvHmP06PxnGLI55/qCnJgLTPTB7w9PCuj
Nw37wdsvuazzpd48PumXEP0S6T7CuUJPZKmz3QxjQt02SVIZpIYtqjK40+JOOGHBZ5DEi0idWU1g
ZyDk6Zt8ACURwz1u9q6DNpl+PqY4WCv7wPCTgt+0A6ZZZXosqUKRpPIq0hwHIKij9jZus/Vm/Z0t
zOo16B35TPvg1bmgsVVCKlMCRNdoitdxFy0pH6GdlNSX0yxhr03CQ/YvwIA3eo63pZfPp5QbxPN0
UiwDipywr1NMNA5BByyECf3fbuaPsFuB98M5rMExzrI9PZtev2z8+7CIW+URsvWBrSAbxjNSyQM+
6B47Zo+uqEzmzhmakFTYV671fJVCDxrXi/2M9BhXhAlGOrbJPo11Cln5acpk+XqbvkwtJIbhJumw
OkdKeTob7tUHX1gV2ap/g48EUtKd6AiZFGtzRhiC6PKRubh19Bh5ecAFTXzZxONF2o6aobv43bzU
oyw09vwrm19LhrNbYmahOl2uj6ziA/snT1W72emYX0vK5A4f7FWmAtSHoKpyB03H+b0Jc5iwD1cA
hHdUUd9cqR/EhrVnIF6kq4rmNr7C9z3+42UoQw8ImM8pN0AFRz84dOvLdQ6WbLs84KSLmtT7CPQP
hNhnUY1WTuBPYD/O8hcWqYQYiiuxoGu61OXI8/4rjwswepDGlisddGSAIYuIzFfZ1e59P6g73hwm
GZTQ5iU2De/TVt/pLtC8bRBRPkNxPlakccGY4Cuc4YrDiuuP01LaZjhIrEX9T1RPTjnr01s7qDIC
+30oEZYGPXB6+nKBD0m5PuFWR43uBL5/4hu66j76mM5CvJ+co0SFL0oYE/KxHGovfjxxfd9aBwUY
p1BJ58waSoYieBLW1AnpaoxGG87HIdlv1Ue+0wsYfkOWb02MPdRphw+NW8FAHX96zWYn/V9Pk0Fq
crDu7GRTRWtC4ojJcQSURySNxVu2SZU6QUNLAT62op6h+Zcs2PsNPUYBiXlZopmfjeNNnkFTNMTk
FNtfyXVFTnENgVpf6Um8e3dh1huR25XN4e/GlUl8+oaVpsO4Mv5BC282aMEiedA0AZX7IrfLrr2U
9NtYveB3i/qE342M2j/nicyoU2d2io/LmtKA74K5jKUiFSMRNTdYgHpGYe68jrAdT8UNt4XVTV6D
UJt1sm+3SXcMhDJPEdXBKL3skOYmFcXMpIAZJlanJdRR6GcEa03CAD54tWj3D0rNbtN9S52wi9fM
FmdVO3KLBGuKemO8UkBWaShKqZuaLt0PWamBSij7KekBpbU2AZPGbSIXiI+z0DfepeOWX+opIYBd
m3d4UYeSkoulHuwpXlB3sdoOAPRawGaS+hEWayQGGhrB862u05c99755hqvlLQMTbU65LSbOTGv7
3H0xGmxZKu0xDBZoPcAZt4ctekvhpmy6eP+Jgct05+Mx3S+RyMwWVFXGhl8c4oY1sjbKFA6kNDGG
t+dJqmgRZmcv6ZKsQZ1tl1O2CMtPoaATg1Cie+YENcqyFi4Sk/dVtW/FeMBOABe4l1j9WbPD3oOV
hQA8LEoZRA6GOi+k3vFYgZ+kt8mvM3B5Y51UGJ1bbNBP/puuQcwMjubgwKbnJR9x2PntnlT7hp6P
5ba3wYvYpABrXRmzcOjU+gcMVHG0kZ3mb+2tbVIcn4gQsO2mIVLa/1Thd/dENzLcVDlK2M36sgS8
/Ewuo0wxXTqh+0/C316tFhA1Wt3btFbmiC5RWj3/Vl6Eawc8Ka74QmTx3dNw9yl/0DiGCvygZj0X
gw8wsM4U8JSYbUDb7ncLmKgjzgDLafIENZoS+5FNamqcB1IvINOrmk66MtEK8EjCH0cemxAxteaa
8+JvDhm1o05YgFxxqswXN7yr2xs1PpEbFCyt8tTjUqv0m4ks7z3RKsib9+J1hD69FSsds9j4gDBu
+PokJPVT7ezn98tb4JMbFSV8EPwn/eOwVZZznNCeWMt5RH5x86No7E1xuQnKcPjhOG71I50n7ofc
W6SaXpQbCbqjtWZU+7OnPp9S2QUfidhlpLWaXL4ie1LrPr5LBPoIpdTroL64FmQ9xaBiETWoJylm
fyaGW1Oh7ANV4GbL0o/ldirHmcH+lA6mjGQ9AzjXFFXYdKtYESeXwoVf+3z/omT3+tAMMgxcfx+j
COSbZx0c3yG2zg+xplZAhirvt7iO9TctbWseMt+MT5ghF2KIc6BGS3Ldy9qt0h/vJiIM7wg3SM+N
yjH3YOLC61Dk44Ka2sIgryo/ICQjaYLn+25H3kHZMPNZ3TkbuSj8v/uE28n8kTrJe6WOIjgMjmxj
kW8wDvkfozRv89d5J2VKiwBY7hPMMhAMTVIE4wZe7f2jCiIbAPtFbxOga2vZi7QjeHBEWSdLrEq2
rSnYYBUr2Q24N5xM7Cd9LUJmMKS0K3Iw+zx5fFYs/n/y3N7si50KvQVayqTRm7Dw5Y1zRQA9ymtV
x/9mF5UNRS9XTF5WVzaAAbQDRSNm/wopMdvVIJsC1/V4h3hIa61VlsrG756R/peziVyugk08eHFp
BimSltEYfWMX/HeXr2n5LK1Vrkomp2jP2kpYdS2Ba10NgmSawX1wKByz+BqOsFHwKvOy4rBWgJvK
wtwLJCUO+rKSWu+cOf+UAlfBHrmezBKoiu6FaaAgktuTrns3uwdzZ2Pe0TAzApVovEeG6VQy9yX5
UTQAmSF8v4QvXr1bERSq7vb+w6YFiJOimVv6BWzO9k+WFeIPvs6a99B8uKAtD3XfBUt5trCyW3yO
+vrQW0XRmT6wpLytsEM61BN7w5sB3M5Q7UheknaRSEVVo2Ofzp8w0LL6/y0c89+m9m2JGowzPwv6
ApNK+hypbC7cMDr907dkeK3zhY7PiAtOdU8ZQY2LHMa8GBpFWAUnuxpz5ocIkx4cS2T9qHbwLc+a
241u0et6bkhu1US7CpdcLBxc108ESQWWCXBi+fopTLeMsK/skjVYFR0IJsJ5HavwCXmfL2GYmCKb
wKjhMPIuF/M7TFAneQDTcZhTaLmiGIdP9ZvUvhsBsRNbe0bz4fyuYOD9qbwmmVc5cbk4NMxFwaks
2cHnKczDhVjXd2zur351GVdRPrl1TxmroykXTVmq+WhmzPZnB7kA5MipFZhf8+yUKSL8XhdrdXBi
RWx9ujKcfuKYOMfoK5JL2dmaGFyCFWvJ2ed66UPRWRwLnDngx5uNLwhPdYSz/tkz1VHkeXEwAJMw
gaHsuq552Nofl7UPcqjVeGSUMMKb8/rOUFWG+TFdVPxktmJCSRKTv7/J7pbGMqxJ92JzHwf4EIne
Z21XVL2w1t7rvcGleSm2ilB94jVx6vl8JDFIDy5poB1lfs2pnbktu1YecbYD1MsQh0zlTtIXqKpm
5/oO36xXgSnl3HHVTj6by6BQKAVky5NCxiBCwzeVV9hbvRndhl4H2SUwnjE/h6U23eq/jGhd7YrW
bFSCPa5T3YKQb0SgmOjhA4XgEI4Gjo8MppN1OXc2xebR5/kzr4bYmb3Qpsve/AOQayS3IDKJkGop
DocSCsJuXbsVyScyo48G6Z64gI+dizRpJEjLoAyVLhyx9zzT3vJ3wlX2+oqJS6BIy23xlUIBz0OY
/jgEVMZH/+S7t1Pq7cVClL9bm8/qMb2fgbhQhJUgOYLixnDeZwnryTeP4j+yHMz6NWm9hG93FYou
haJPEnLlsZbogcmV6p24t0pDJpBBxIGKhpLA1NMrJJJZrjvJ48KAdhI3+lhFkRJWwSznTpBPgtlj
vNxr8qpxTO41NNIil8kkNds9zvrP2v5c07TTGi0S+c3rsvrekUnBYll4zvCkebNJnWkHuNEP3ctD
CZzNocbl3YZ2FxofcnooqNWb3vp0R7Q1MvPuHQNDCVKSUIy+M2BCylH+RTbFzmNh2S5vVTlAGF/j
3shqVMGzF4ADez50hSR95l2W4xCB4jyhBA8i8lD35MgCnyWT+qiS8yg0weIOoUhbYSOi+Gq8eYJk
2at2mdsMP3lG9telUYE2h9jOVmgCNo+VGr0y77KBzLrbRW52K8RBvFYNb6qpnxWRku47+uRB2UyX
Yiv4/nHFjZQBnBMz/wAujo5yDleMOY7VXIBG6mRVQUQPRq0QsXXIMvLpElcRhSt5zdmuTzxMOQQQ
y1uKSYNNoCxDy47Nm27lOZ6MOpeRlsbeo8+vaBdQVZAFbAv42KDzjVj2uhxdXih9ZvpLjp+Oy+2P
xTKK0ePAHKd0CH6svO5lx3dWu8zfuv9sCY14yHAhjksUzNYX0QpDQtkZq5nLo7kh+nh8qoXDuWqi
AuSH/oZMEBUi94sNbbcK9UFfDytwIFoJFklt3DJ4LtWnEAWxsxOW4OTdLl/Wy7pkwYsVZCBBuZ76
/z0T1mbRPxBi7LIO2/1AhX2/rWKodVD+gL26awWxU1JpuU0iud9V4oUmMfT4gjqbwsK5dn5tVUJW
pwxyBHYVGqym7QB0ybjC5YKfLvDqWVz1DUGiJkM5t3/VLjUd6w6aCODjloL7vIeervZ43hopcdwr
Xab2uII6YTFWA1kUYZ3F0QigxW5DEjHJIzBtwNtidq+TMvvSCgjk52B74Tg6EhvRWeWGpGKoGxkY
QhUnS2GIwIfqw/qE35maKqcDypo35CMfq+qururi8ChfxDMinAKJe3f+reSkKUqBpVh0O4rESInG
W5ABCcvuh0yOD28pj9YOwUqwNy3nuuYTDaAEFHVCdR19j+N0NqPymeJfK7wC978fTBsAAZsyDJSB
DZuMPSO7a2WZ+s49JOnUwTXRqQcUOSQGtGJZaX46s1hUQU0ZYZMR6BrvJEdg0CGzQkd4QyhmEP2x
t9rrZTqY/TXVa0QDGYz1vhlmGnOHV9GMiB53ZwScprlx6G5pdQlf75ibnPlB7iPJfj+GucJ9KZL8
zLIpl1OKCS1uHX1sCaTMPztyuUmFjlmV5fFEL9RqvwrVmbH41/6ho5HIoSYcP3tWuI0SHytItdfN
+GBmsBTo03KFSQ7d7vFQXTqsgVszdxXlvSwyVJdTXM3uOR0U2Geu8oni7pqcCdg05zygH0uTBtEu
YvabndZJQVdLqMEHIPYUUM9armx4VgvTDlM/46Lh2aH+gKHDIG6UtkYw/X3/64fumvuuwIQgfQnk
NtXrVwcitAobgwGjLDT5P+QVV7LMqZ/BPRPAtTCZ601vSsrzA6vX7YxlsnJlvVEo0K4cg9B5BTp6
G08hhtR7OcVerAEVGrTml8/snnf4HtXTuten+ty80GBHxToVhOTfSyFduBiyMXK8m3eyQi5X2/ev
dvNOWp45zcRoPKDobSASExE94a+src6IMNCtZFgBkK6Pb01rloa55u/hlzLI+6B5ru82UuE7q+li
emLZojvlmJ2jzmDmcLO+Y9B8vXWvWPO0qPgWLm2j1DW59J1f9Tn3HoMXhpgpJp/IJa7eKwKGbCL/
4JDqJ5vcc5teZ5+GMO1Ur89AG9nCI3lKJcZoWMqamU4xINkAsuovIxee0qvfp9mRsn5d5BJv+6EB
A04VicRbZB26FvTCrOzm1u8FXLCH2OBz5en9LdKPAkhze545kN9WFydg4dhvpMF6VlRiORq6TEBl
5Vi3PC41Stc3vM7GzFUGX57MGQmcp/oVXFUJhdJMt9SJTVRmdp5JBpLnpl8Xi/L6B9XlfEQQP7g3
fMjn5VBpHnUnS7Z7w37pzaIN2DZORIBl/rg71l/24F5XO+oWrmPkPdH10s9cEZO+sTieO6DlpyAj
sDLoW+Hm+p5j/Rgvx7eVwhrRzBeew5LUyYxmnNHaPllinBBKjxP/cfEz4l1WMKJde8RD1TD4YCbE
HJ2majOnI6Stp53qItK8Rdiru8IWatAvUX53UfmRL2ZvzWcjoUfLkIrwltLX73svM/MVeCCUGhcO
kxH3SXn5rDvzLMdTvVMOMrrogkH5C2wRv4hF9IPjHwrVbewt/TIjRcLQhxHF9jJmVHl73ZLbyi1n
7kxlmMCX39ABIkT3fHhePdGNvdMc4tZsKVIaPMZbHfzKJCyWD6+nXA9mPzD3aeHq1uQjkinzmriR
NT40obj/4zf4jfii7Pba9pTFtE6a4m37K0E9+wqoSkUu0xUwDsGILIlptK1QI0Te/zxwGkwaKh+K
6BCdTNRFtQJCGtcC1m7vJ8ArlBfFJGCvpPoGIcPC6ttqHUZKPH+8fub2MXTn0R05tVRbYYhL+WbH
YEd7tOVBbVEHVnWT8k0A0zEtg5Xz/ErwmfZAsYijxolL2M1Gh+HZLKV7NC72EmfAGegqc6+XBZvq
il0dDdPAFsKnG5lPGEtUD/7LtugUCcsjWqum+o4HBnta6svp5oKqTiyccmSh1PlU2FwNgiVGzVeR
2VeJ5ok8RJtY6GmlLNAPXYjSiNaBXEVgL81D2VYBaC13+QC07g6/WvkC9P6i6Dg0/ZzWOPkru0iS
mcaAN/iM573wPwHWWnksIclFFyVGFscuQbGdMQDfxb2WTngIkofsqQLqnZcZAn25USAbkzQoDSP7
MaPH2YO+dP57loN1su9fNP0uPm/izzkoa7vsbWiuFvnWtRQhowaZVmuB8FO9leeGBMlkLbC80P7J
KSU4OyVgL1yGxR0e8iepd2wFBLXXQygY71nnqDjueF/b8OhQqoWKE7sqRw9CIq3nLv0Sh60hmbO1
Pj/GECcH+DIxW95cLattWaiby1VjEzu7Lc3A1AvXg+p4iyNR8LUnm8qB2MFs4LxbqCj11GhUX/yU
u7YR7s3RbdXHENAy8LjQ4azBuDFdFR2rZeQJ07l8DnpZeqN1Dcmu2ONmyScsOkGs7upiyr7ZTapG
8/pKNjuy8C8RnqubbfpM1h+qN7r2g6bvud8Kt439I2O/vyKbRBORHaza04tcfyrLfgZwa++s0RfV
m0mF7MQqkb8q/K3coaGRPOJF0QRmQqZj7FcLYeO4doFqqa5qIwT0mKLeViHRCU54c/RAlm+Bfj2I
iVv9yWwmlKTPtIj9whSyMMIM1kY8Mj6p5f9yTiAhZPRz5zhAS6+WnYAMMd/PbRHmwI5NE73FaH+2
KMLHdqvWN1PTbKd07+gNxifRLDmcOb+hOWN9n4TzwVTMoFYr3p6OE7qYtUG4oa2J4GoZvd1BHRy3
LnnIoqSHQcnW2tDgfhODqOypQuRDWfKfrgGGVKM96YTkb2a43TRxSMb0qzAshk1xATe0hH6TgAnc
/xZvT9YhKMKbX9v7dUEMXyIZiE6KqEPjODSX+VjLu0z5INqo2gzeC5n/o3YOM1alPmYyBv+NPm0M
O10aB/TeccZwwLy011rgymfal2WU1Vk9LT71vGOLp2kx3OCZRJ3+a4Bo7ke0nQZWEzu20jphVOz8
2fqJEmoEAXn6m7xFQtoY61X8n0BpxJ/wIrLbZGz8kiVKXRWc5YnIt/jqKH91AbvNcnVte44rPYmL
sdckzSAPWmieyfvpy0FnbZl6ZTonMYCOrsbmbEJRHsYmTFdDPNtHeoCXFvIfGUlwoKZW8OCAQFnf
kLMLTHtbXa39wK5/Sg6frx5o1KZc2txWlc2Fp/tblvvqDKUbNMHBgVBAYY5xERZ1hfXVHuPavKLQ
jCGRs/JSELdFkizSpIXzdIumPG895VLm4nOPJ8uwFxdDxEIXINZZb6HRuQVbx1y1ye5Prw7hohwJ
5/dhQv0+vWu46wC9HEx0fMvo+41Tez4BP6lqHDfnmVolxajYL85pl86xQ8Z0u3imlKvsDvznAYTM
0UroKPZKGtvt9lVFB/GXQ0+C9W8mrQGPzEHmp2cE39KGUimRehkcFzX34D8HTO86Mwz4GHAJnQgd
vGupVxFnU0Wh1lAlZjLEc9FMV2JymMXhIsumDIozATxraFORX+tMYPFo8i0YEJyBTwJhqN9XnBeN
yrIWrcaR3fZqiOqeAqwJTbsIxpCnlWZKKPn6uy589c5RbFtNjfp+JB9fT7pvYndFnNE50DIhri5X
hZFxecL/LFkiDBdd7Tr+QC0MZUSe4n2VyUOa5oTFlTLKyYeDqS9J2Dui2ppZzlxwEkKUvBavtIbI
vDxRJ3Un5r/Ab5PTxm1aY8C62JAGrg1sulZENz4BTLim8OlIIEHQa+9Q22YD1aLPEx78ZahiGngs
veVGHbVn23D1HH89oy7pFWn1yixFu6DHNY4IqUxKHgIvUORmu54l536/1iHNsiXaBhfGPemIVVhR
w6+NJOH7VNy4S//56hppPatp2XyuMxQZ+qFGhlT/vjuOq0KEUNO8BhxjqUFQyBUlHqTnt8g10dD2
1Wou1QZb6fF/3nAVk0k7dGyJ51DImUyuVG6SpPK7wjnhHL4BdzmX73XdXFpmXRKRiHdOZ+pM8WwD
DxK9s8ANjAugUE6uIV8L5yjcKlZu8UJdHNJD8xluMv2+FfRLYkPhKUGkRLRyhguEcPoL0nVBatVL
gWqwFu2PAtG7lsIooYjhRS9gpz/wBxMd+eRghlvwEA8l5wmXqLiLCMl+hw9YrGW+ZtIDZBAIpMz8
0BF7nOEREv+Yi5mRkGC0SjyKZKaVLsjZJ8+CmTtnfmhb1p8gzk/g9f7+QS3eoqHKsc8ekB+SgVPW
ONYz1k070G3x3xVOPrP55CouqxwJQrCZL4F6goxUQyW1OFoJToj+50ZVEgsNlftDzeDzy+frha+d
14Q3Wn3wEe7VSsYQ8eu8Lgq3r0h56zVDij6meMoa4wr9pe0HNpvKhwJ4bI+iGstmdXCjHPdGxCr3
4SjUoUC/8/NzR+M0vos1dvywfKY7Y1KnIfMpwzZ2AW+DxSb3CGV8CMhqiwzdk0nGuyEDrBLu/LdG
/pMJPd+oku/KB3UyCI6zbkmcQLad6mw/Yd9RmzUrjv9/Pxdyc7BxU8m77itsDiDnshLjQLWA/Il6
k1Q2S/Ru/C/FJJ52Jqotswd7/W+aG4thO6yFJUtMMGOwcNjIthyC0EP0Qt2kRwu5nn1+PBEX9fgy
gnvXKwvytw1KxyDIIT5AScmGDtdxPEC1fPARWsCjyz5MQ7DFNVnSg5wMS6Wt/5ejTZqjlglOV6ZQ
FcFOYlgfu0UwGevQSh+uc6cMHcehKIEXp3QkEjybYUqMh6vP1mgFxXA3hf/NKOWS0wMi9rSNrOS0
9WWYuZ1KgDKaJ11s/9LnZzYNs316KL/gasJZRyVf2DnXvT//VLxXzxDNYT2NdMULQJ4bAqvBqFjt
qJKZONTobDR/b4y7XDntlqBnpt+CT+6nq5BGMsS70MGqUBiX+f3slKe5sTwJrJC/csiCB/5CbUTo
Hh1UVHhLdMwbZyETT8/Wdm2H/9OcCpDZQuai6RPt3jtw7DYkNdjUrtsfbETJbDAU0clDlspcoNTE
888du5+tRiWzis73ItwWqvBAxotCivU1JQqxUtMSXlPlLhQ/KwYSzm/n9B0E03eXx9ztIl4Ms+42
q7ItzWSc7QqhVcSY+BWpWD6gh4bFi9KbyoP205QSZPQtYqiRMwiDVOlwkvb0670WlkWxnRXlAMTI
hMKYvgq+KPPMOJips2iLsPZj9D4kbE0T6uIK/OhXSB4sVyUJxigTMF+a0AwFZveQZB8K0HnMbcHh
z916C7BoeQa4gCJUI20FNtCpA/3W/twVP6GhN+hVu8jXhCOZOLbfXOdLT3x/U32Hr9rqI2bXWN1Z
fMXZjl60z0MolrCrJ8b3xj5HcoNRLdXnLimxEXrc3yVXII5Vir4fSiKtOsrU6w07mXdhWXLr16NL
EfWSBxon/hgCMmvmto61rXEwZEarkb8tEeUoE7FjUQ4MAIyeU50QYaEHYiLFVHcdTJ99/lkyCPVt
qsk8K+kz0vBab00TBwJvjaZDUjRM05OAl7pLXLUCzCFUBEQxiHbPWMCUI1wcy3Q1XHfPqYQuM5HZ
s7WnksQbyreIgRkoLobNqb5AQ05w0AObI3fFnU3n3OW1J3duHA9Jpfl+6wiwKxb/kt6WymQ+9rjd
zHOKl0z7zGlYYpE59WmHxdUyKUM7iMc6avdXGAVC7+ccH6LwfwX0coXbQvH84ARLY53kynBRnjyL
rd9quEV6Az6TAn0FjjloHCx8A17lyeAiOWsAuNIJAChV5v2gxRN6RM4dxkcZFCkjLlberDSXQF/j
uh64UTPSL/iRr4Ti87kDSo89QAas1fzD9UtihC4edHk1b0BoVozkx61mDJNeFbHmuVnwnRFEYSfF
oW+xSXOn89ldSsElGC/wgWjjPbW2EBVvAmDsjEHOM0TD+zXl1ihLEvz/S3Qvs+f7lOhTo1NdlOnN
anTWrmKCoA6iMp7+hgKJjzy7lOkDEMx2y0SKc1tshHiDfQXIq20++7QwNJv4+uPjbYr7cXX7G+UU
Tz10tiQRbjrcgw1b66iZKBYJsa3wAHX5lNQnjZ02LxFLEmb3vmEF6vRFnDQPJrVDdkPq2TC7TH8r
F7Tr86WeytJaShD2eO8XwbZF9jPSdTN7LosD3SLMfme0nq84bD9BDFYmWVoDe8cuSDaO2iF1D0dS
TOQ9dsER6plytpcXXNH2dnnkGt4Ysdgsw3vvyHQ+x1px21x6KtDKGAXPqmvyZnn3BOtda6FRDKpy
g1ot033IHlN3L85o9KmeF0j2/QlW1gMzO2fljDjlefnDhyq8MUl+HEhrBNkrZpu1JHEGAX8dnfph
yhnm870xFSSA5twukhlNatsyPJu6T7eXj/XBlc2NhbmLggc8cN+UC06nPro0x/RNlQ6+6CBDUcYk
gNi8ZzvAp13YCa4eXLRBJHA8ZZah1E06xy8+aXjce6NaEVFij3AqA7HN0YIfrWRvVCR0vVtirohx
wGyvuZjXeL/35HQQwLSQsF31Mp9Raeouxr4lZQxkSxxLfDynrQNFf6JvZe6KjwSubxreKX7aq8c5
oFDSF4txQyadnHTzKlBOuP3J1nIoepfRapoabjJT30wZcMU2KOD9aLdoD67sd9VqLqh9WeucqGFd
xpUxCtjXTKCn2bblclvqJjxweRW+vZUmVbPfZxFXE+6Yp4u/CuCxGMEGdm0ayFHmP9hYB/wZ83E5
3yQhtf8dBYA+wkQEWEn7Ijb+m0fmNcdqb/2mBEI2afRrTI5LS2lSKqtO/qjPAlJMq1Ul5y2jfF2X
DwMW80HiFoWuwM8vdXUf7j6TV0a9OCdRNTiHCjb0mcy4cnsdyPfI1FaBk5XxQu43OQi92/hsrzRW
SEhgtohmLj+6AGxEKgZB0sA3+KtT4alkzev2AHNiktT2Dh3K/6qziTQFKK6bpYxz896+mPlZpqn6
4aoEkJu7WgmcVEmeRnJ2Z0RbcDXtc9pb9SzReAfGdZLH3ISbfw4VozgCApHj12c/1P/2JOiHt9Ol
yo6bPYaLGYdzcv4c70cleCJNsXG9fKINKDwImZuri4JfjTpDjOaqOYMCMTOI58gQaE5XgIV/bJkQ
5AoOiLIuLg8SWtX9qyzwPWhIK65JFAKxAw6zqd3QT0ZY1N3Gt4Ol9a0C6+Iu4ene0ZIe/UrTTUvz
LAfcFmyMvudDJK8ebQwj9LcawKWcUaeH3UdDQBhVQnNWt6OdTaJUSpeDSNeYPD2OtYX3s/A05bO5
o+ObqsEQvItcDT1oIMViaexeMbArgwLJgfG3NNYjKxmnisYlHiiMGoND0n5jr1o35gTB2TL+7mqy
pifUTF4gr+T6/utPMaDCv4JPvWpaOncoTqhCkorOtMPyJVuaPvffBIFU6cyg9yKsq+gtSt+lELTN
9v3J+pWurjr63RxnENS4AjHWDQIm2DHaN600LyY7G2grGuknYC/7dmvWMLdXpZxok29NLvgxDu+q
FW8pCzuKndASb11PPd6ByhY/vJ55M0lIMv2hlgYrWQe/Nsq0aTT+DHvcHtmaUOCBkwLDBu09yTYe
j5y4HjmAe9ATcvwkTDPYgzlNK0j18O1Bh3jkjSjOyG2ysOgHGOnBx5+A1X9rbsckhbQ2VcjgbBkg
LrknVlVuTYkavi77OSTrKVd4uS1KhjmphwIPbeoaXKb2TbeahFVBZ8zFaAXSKlsqynfRsXlvWVD/
/uFARQbDFwvtc5Jy5LaJ7RAnUAhZpCkgd3jSViUEfKJAMx8kJxLyOVdrEy/M9lmlVhUJAAjhJ8EU
G145nvVa5iDER92OCs4MITfbZjIXQfoq5UtXEGy4zafWh6ykHk+3rghvYoHootl0Af0gz0k61Kjk
X1yOL5N4LXNVifse2aXzXmi8HWiJko8tph+CFkedAlhrfaqBjfEAvBkhnTHZIjD4OM4K5AVbncnM
shMSs64gkUMju1vGvBsSOjoc4BZBZg8iF/3XDWp2dM4k/bzv3GP4LAXthiLCqRvHZMxN8cbE4wdv
E1ETgvE0AU437vrqyr07atKwUKBh6YcWK+/3WXy1hv9qpK0w6Q+r3YuuOJ93kU8yBOnwpdGZra6x
+3R844lQVLv2bjeCIiXHBG31KS0UnJvImHv3EkDTNligO1sqnvPnlaiglpk2B95JzTOw45NMVrXS
cGywlGxnDrI8WTONYBgYxVQUD1bxloR3RyEEMh1ctIwNhIteXBolFjWpGrNCs3m9CyeMAYocqlkU
gdeEcWVyObWhvMLLBqgYvq+IPQLk+Vg1lvDRjfWtJNAqCEqjVRSEgw8vPlJRbMIzh4zqt9HMuL+W
o/5XXhTcfMne5rimPm7O+KWx1GzCeS6cxpNhjminfDIQ9W2L8RnZ/StnP8xZR7pIgli2gSRM3SeX
mk5WgVxL+THG8W2QbXtha+auTga0MOupcPpuyeqez30muwwtmpxfOEtu3+V/TaWHl+NtYRfigEX+
uAHe7CMPBqVIpklwaHoDD86cag3errpDweUVIz1WI70KQ/dUHh51Fi4wKAiJbZUdeQslHZve9+xW
RjRlHDSshmPOCc7M/l3mNCZ4Z3GyUIY/D5eZNN/v2mluv67pDIgoY+QNW/5RDLumXzJu7IotBVEV
zayiWq12h314hvTfCcR2Y6083VZnNa9fUtVdxxUk+zphCwjPSiE4n0Uz/yDnywODKTU90CTLen2f
9e6qtHH6HO9oV2TciFEWnBRTo1OFYrbQ8nr6e+EtCRtQrDfoucvHeJdIm30dj6xsEadIsIfQm22V
4nbcwmaQ/o1Y2dd3w8WEP1EUKO9MftibW6Y9XDg570gD3Yq+OzwzLma9uz3dz0pQlnaTutKj2kY5
bVzvxnk4+qoOwsbuymLW5stE3oZSf/cCOgNb0e2Qj4Uxk/J8uo8XZkLK1fTnNn3tVSwVyjqA6eBp
WUdOMeAiDYhr/cO3g4Qnvp4cDfVmE9P/R3mCzX1cxxG7pcZcWH8mrYGAtJ6X+fkxtcwYaDKVHmGZ
VaMIRCy5IaeXDpySCmDIOwXVXk+C9Kzfj5mO7e5A859u5wltPXvrnLg6CdZvmuqXxq9opDJuxyvb
4fWvDhi46GBLfj1BRMWIjOdsXqJmA6fKXDk5zvZsSYeszSotJEVb5M27RqOeBymiWvayoY0M297z
RqCaEaHl8nl71l0+A9iO7ZZZq6Xy9rwv/YfMELx7uifNzCViVaURVm/LFhKpxxWR2v40WAdKY5oN
/KI1rjHpxbpzR1VesJIViQOtyh/AQsk2Jn6RHIztfEn0ZgDN18rHrbrADGv5ARvzOm/akf/kRfnq
NzM0hJf83A9ZIm+iIGH65i1Ek4eM5679u0zr/rTd82NLgbUKr0fmVCfsbzh3UOWpoYEkgOGvXzyB
pvM7ave0l+d+7OgJ/GeKLW3Vta/RADR/AJK8gz700koaEzf56P0KuOCUUZA7cpDtyqcvqH6np3iw
LN0pGRLdzz2K4QPmgvMEWer9Z9wzVa7ZNnty/gFAbGkdJUuayes9EaRo+pFHaR0u7pzAO4kbMbvI
FRkccLsO6spxUz4X0oCpNFZ2kwH5hS3iu04Nbg3up0t19+DxjBCtNns7M2h+ukVpjHfMf6yWmem5
N8HtCFtzQKmt3dhA6WNATFXYWzTCbh7x0a7ejk7c8BLhb8Iji6LhDjggbcSDHJ4z1Sg5FtT3dxNB
Binm/QJISL4K9isrOwkcNrBzGsGb93pyFHmWz46MRjRcyTBuT7I+Py3DvtzuigtAjZHfZ4OHHbb9
ISSK7UQ0F0uJpWO5Jyk/MG7UdJHqHbfoL1BBjfZNBZMKdc5/IzyfgYnoenemTIqxTSQcUN//fPkx
TvNEUK4CpfB9JuxvREhZhqseRcP86OvbjzIbTyFt3wd5KqegimTnS65VLZjH09MhBapJ+totn0pJ
vTYoi5lf9QbnYyMPNzNa3PpY44V4cxtVIwnPXc9VGGZi6FbkHT7gJPWDR31t1gVlMDg/BItdqdVr
YMKDj177NLzFV2rUvXrwpEgp0cDKxkAEnT8ONZBbfKwR2lTUZn5+J9rmGgBqzMKAYV120a8Gtn6w
rjdHqhpW/UE4PjiqhBKQC5khMprdTyKuSOIK5TLRerRj42YnC8CzI5iE3wNCv2paKVBEtyLagS1f
z8XPrHWtnMKYh4avxhEis5xkFXV2uEUdv99eQmAajJO8Ple8ylCYyIPxgeGrjBLydOlQo2Vy2tNb
ZicPlxzUAR7tv77gsfRbiD3BPnDW0FwUV3ROOrs49/LB8Xk/Y8lgNRBytjh/hvXE0YPznVOI3f7m
8xNonfQvgfZgksRE8Xiqx1I1ojGepdHICbPeDPVzONNLdvNKCYIOur9V4r2F6sjZVhmjSk4KMere
LSqKxbBqMel51HrjXp12D8qZb9Qm6TEgAJcqbJ9SJa4y4Om4g5pfaKudIhitx7r2b88YLcKQ4SKj
LxOsvo0fvCGVfy5gMVjgmGDbCMzwqg/t3xG/+qr8jxGtwW49RLNbeHsZ/8ZNvsv6wwVQek1Ix/pV
Gs3dXYbOaGq0x4ZxoeCNRjUeBvmZdpua+4pL9GpiCMy+sbeCCnaIROcXYEooMTg9jacxEGZFO1WB
0M+OLMHZOFh9ObH/vGfwy5r4g9wVOXnFj9j1H2ff8ytY+zQRK7LKGbCnEMt5P7J+Q9/0iXaoVJhG
eIi9x8xawrTRpdFBFPbQA9dm//lSrsQPd8asnKAPUOsM0ghSBBePoh1DebNEtBtHQyDW18O3cR8a
U2O5AfKq6NxKP4Klsg7Zq3rst4MdecX181wb9VMSp/I+FP9TLQv31doWdWHAOxLvmB6ufW14Vb50
arsnyyV1XNf8vpQKugAr2wjDKPV/fdAJ5SpygCcdBkyzU+FjfSie6qAwFvuJ6VhvHiVa61KPwzUU
VX+nK0ViHkSO82mmErCcBsfwAL9AodKeGnvorptLxjRGacc26ITtf68wHSQF6Xoe9DzA5lER5JbB
C6iWFDvb56qt9dvyxD0oUskQbdlI1mwNZCkaDn1jlUvL4dU3LeRJ7R/ygiYxcyyG0KLp6raxlM19
peJmwF2Yv+pEFObk3QLRQw56cpNIM6gsiWx4sncpOY34pO4FfyCUfsrX+qg6Av4liiLmUGpPS+0q
zUQznobtTWh7rdwoc4/g+6VFMazGlBhL0tIROrlwlvOor9GZoge4qvQJZJrpm6oXU9ReUKr62GMC
kFcsvZPhQsR6T5H9eFTcKlwIicLdgg7n0pGcYw+CdtnETak/XEbZtsn776qoCoQ+ujZcXR3rRf7U
B3v0mKJC2nfQRtWnF/jloIEAKFqFSnc6rOs26ErtvNn7nNDSTs5SqzTxs03T/AAkjfPZOV0FDX9i
JEac5/4EfE1s0SK6aM0yqDhhSPTNnCpaDz9X5iUygCsJOoTKQyqrHzs1dJNTkqs5DJLOrnoqSy+H
zeyWdoyusS/XBtCSSx55WtOsSBMwG7CWm09/LRcm9UMZIrbP3vzws+Rvy/245B8YVuPxSePYDJlS
G6JKC0m5tfIqkit/6fpBAqGQgC48QTwpbBzYoBotgzvcKCQhh4JZu+JtZyvwe5nRMypWTBa0l1e4
3cQEBxHHh8XAjj9JzCvMbsK7qVsUNwUinrcsL6YIMZSLUObLqA89FI4wZDw/Lh8GxbvT4kKmH3pU
cxlgKdSnd8Z0Pcbz02hgnZtverdEpwqH17pUy7yTdPhf1GbeHhoqnVPiieO+lcymYfY49Sxg4gSJ
o6rk75Q4c2t/fKx4DPDrz22TGYQRDN0GlCWNOAf5HIdi2mqlnUmvlEAIsNrs/bXS47FL+fOOZpZU
QNblrqNTUNHhzxIMRg/4ynx5OvivtzcPdpZoP6ooVBKO2S0svazB2sBcFvAjvTOWWTwFHJ5I9IeC
6OzCSqCzpsSnQDvV7bf3kgEnggSaSNFPdIG/2tZCrm5F3t81eLi8GvloIH5YGvwGxlrVw6OuRNxv
0S0EUQR2fACNlI8LrHLsBLxye/PWFZtR/UD2MhS+9LGB0oQWwu1Ka4qUsWfnw2UVyE7n0NCiZ5xR
YJsRmT8yrEfSoUfejUgx7AI2Z1w8IWj8ViPIQY/slLKRsoYGWVx2/iYwSqiFOcjwQtAmPXovZNQV
q4Cf9aLXBfjblYSCvGjbhvZmDxxER6XqRyNuCsGHyqyPiagLX2wCMlJt9s96A/cdXgatxokdMTUH
E3X8MNAUiYwjyg/a213F/RJ1v+TD1tYLJmLvrtIMziAE+sJUW40mbTD93b4PeUma8X7tDZdXf+5q
d/v8nhAT/CY+D82aUz0WIWyuAX4RA7gmUf7t4n5ukyrS0pLttYvLeP7ewalvkpoxwnl8Vf/jjK7y
nXeeZSw4hBzsiwotCPHuLUz0qjJ6H3KzOwiMzDv2TVxCg1KRHDsZhNCafnpMTkS1XbL2eFamh7P7
OpwA0GyW/Xi5uaPBhVvjHLlDCdme5n6Bna2zswDdwWDwNg0LLScYe9T45EDzxCpO8xmbD9PDErPP
eOrd2ZMEkU/oUnMGpCp+OvX2T4vrxGWMTfbN33XEeDjQ9CnY6jujwcs9XinuLqHEbCohy+w3nJgr
r4gL8RouJpvf4huGpgRCJe9YNTRzr9Ehc70Ta99CN0vRhHKZwh3Cs8wELOWnO90n+Q9X0sVmMTzP
NsSuN8ECrEb1/ZXERol9axU4HeH+SslNIF1S/UVlhJWzo0nsqMPWLbNbEeuOWYpCsiy16eFtm1QH
pTfRRdzNzRnIB8uw9WJ9jwejrrvOr9rXzNUZOWyHF399EgboGLMD+myIkR2Y5eKM2MpAiiAPXRla
JIHTKd3ffVPjVQkVxFhgGsuenoqav8z/9hYWI/I33TnfIjUaa8wbPDZsxN1kJR6vhKIPjM1rjvqX
TpobaUx5nOXdKiqgckP7X5PhgyMkLxvjj0MeM01eJZM0ZmUXNKiZz9cZ+ib7CO/xYmDjqNytAzzN
Xj71rfcB3JsUfvJoPP6uKR52In/9T07aHe4S2LXjxVvsBAIu0TWjNH2IP/Ikql719VXvce0tSP7h
QmeiO4af1th+C8eg6ujqA+lFNOMDj/NulH3fdYAvtR2ifQlgEryvpPWHFaHq9cnjX/dFZSc0SMvN
w+L0DSfYfV95sRWNq3WUvBn3s35CVJfJK+5bfZ7gm/0fEk2PJgB89Nu5Jx+IeP0zNzmglJK6TZAS
+3QX6NPAlnQIR0oE0ZJG56WAeU7bS9dn78Owt543imEoEi1dxtEqWQxJfod1PzGWPrPDiVMVwrh7
cDiaYMtHVP4shKhk7cy4TiIFkDTsOQM4lyvEfyU6ZcA6oSoFgtQDLzM9I3OTvD3trggbpjZDBwyv
6j3Oc6afFNkSymHy2q2Ahaq3XHTcICRWGG/BDTT/w/bXHVZGWvY4nJSz2J6gos6jJPM4uSABcBlb
zycRWp5UBGEWW+qhnLUXQDNJ8HibM88El0z+PCy+nCkCM1cXwCq5IDZVo9AXP1g/zqypVrF67HJd
FuLLfEZl1ACJe44UMI+fXSZjKgoRxDaXtjI034GNuDchn7SKejRC508PlB8pDrbDhb00iFNz65y/
A1nm6Kg0cVevpGCP01TeaxQzF5Pnp7O9UQq6hYUi2mHeoePBT/5dJONDOIvvxezJ3gPneA1MSeeo
m3ryGRSepm2qTTQLOngL3op3mekrof/qywlZYU7H0u6QjSeuHeSPueXpEwvuskKz+HnDsGzHSPmu
C6PPMWLlrK3KFcZzUZtIEnIkdQB4Q4YwCys24lM3eZ08hB3r5Qj/g39ieXKqDmwJ/daX/SSmRYJY
JQdC8DemdyXQO3uGENtWGGh/F6NI2kzAAG+Wz/VuBkJRPJXfDVs9kg0dh3/DpaiqDED5WTB/Ong9
iAVXaa3m56L9Hm3YDl5b1SdNbcdj9aiSnJZA/UrJupe+JT8SFs2aZvF/q5uzKKpIgbGhJqQQs++3
WOf4Bf/s6KnWgWnl2YSquu529yWoEihv8KQoLt1MaKhAwuH8LnEakIHTJLc6BPCufA46JC0pkX46
96A9TcOK9d2IbOwTMJRow+OdRVDZb05EM8wYqubYX4h4C43Xar0Liwbn1qqoGPdO16VHCNiM2aV8
Sra7yfStkLKHV8Dd/LIwDJboamh+Rgl/QvdClbnaWT3MMCINZMSJTFgo9+6IUWCGMlJ1WCCs2y/M
YhA5AFLUzYSrNxcEpntjU25MS3vc3QzqfCCoa8AjKMT7gsGTq1u/TsFEFMNsZmeSUN7PmUlLjbz6
WwGfQLZBk8sZS+mv0CxZ3L1ifcsyvn1+luQplrg2wvyxo3TwM20b1VBQs/JXg5ZoUT/0jPOb6D5L
/VqUMsZ2+AXk1JZOG4oWicr0pECCKIUoEI4lN6QD/fMNlpC4csLHxuHcC2a+lfCs7kHE3ZJy3pVL
pqaDsaLdckH+GD/Q/ulRe8tExCWgbj9towHmxhJQWAg7KS6JWS2zLjGXKAqF/SfEmY3wju6mBHDk
Se3C+gisD6UrdLaPX5YpvkC0Lf3XOvXUBjsJCLAw9GkTAASinFywErCN9DKfplH8pa544oR+7/lp
e19PF+jhmc7mHYHiIjIl1nzAWcVauUBZW2OsQci8xkYMITMsMkt/8Awn0a00xcTe+orjv/kJSPJv
sp5nuT5G5hYs/K8jMZj6kyYsRJD/cXNcN/814tyz+SSoJZWb3IZmHlVWpwKgcMQBnHgGHYLU1NbB
Rvn/P8xG8jtKN0Bb+poAFc1iEn2CWaO2FhXgceE4euECPF+kh2XG5J+0rf9EleBiHMYJtKk4dWaM
0QZ9dCMAugBdhez88/NKOlL53pMJRKKz19b3c3WU/GvzIZy1Ij/ur//mDMpSokSK7mD3l0ubek/R
mTTFuKoB8FxLC2JQLH8p+cBlfkr12AdY9p2XsuwpEm8EKs8dJL2cqb9bCCZvSKVGfroV59gg7eT7
PgAlMH31sWySeHa/kz1ryJLwhwl3/150aycVtqpxiU8kymf6/k9cf6aNuNSrCXhVUox88kY5XyUV
kZwVm2lpIDgoyM4d6Q96yF7uIxueu18smDLUO+BYyEVDN7WsK8MHId/N8rLIEn5W022IfVu9q1d+
sijQvVMQqSCOD8XlyNgZCq27DGxY1lWe+zhsWfuflYPJTzj6L6lbosvDt2sercB2b5GWofoiA+ac
H1YSpt42krpvSIAWaI+HrCYgKVOSbANF3x/UyJLGSHF14sk7oblu50fODtCexFjAGRX+ii/xeyUH
jMUGg+F+XWowvJMxBKYWPH4LZjO/huJ8dcbdLY7yeBbsMdznle792vu4GQ+Yb1vmbKNwng4PKmpN
5tNnGM3cnyHpcXPPV7M4t1Rb5fAgyjz/Fx1+UAb/xQNk833do/Yih8cl2AAnMiu+9Xerg6WJPZIp
bnTGGfqcAkx41HjrwGqi93cL1MwpnWuFV3lTwA7drk1RFiootjD2Ehorn34GC2R7radl7CkeeTJP
0n4I3NPVoSTX9o5AyevbrrRN7x1ryUSbjmKvuzlJMsDQtnHR8ykkbutOeHSP68wCugTvCuTzpC+D
QcWVYvDXPb5NXuCQpKgDT5Z1iZosFe6zIFTz+Cy4zksJMveId6PVGwTple8mQeKPChKYx0ORWgQe
Eoscjqs3nvTJlmB0Tn9YwFZkMgJASTIN5+BrJsWX3whSG3px96wVsM2hZNWFCwKWkJty6cgF+EGn
aN8j7V1F40AG4mZ66zaFG53pCUGz5oiaFIJ1frmjpvlJ0JPZ3nRrmBETIHmf0dHekFZqIESDU4Oh
USIGy6x+CerNw4jK4LhwfMzMiwUzQC1hjnHxYCwjfpVGhh10RJVLYU5tORL8XFDAdIg574PysIin
MSRHTBfUBK1c6j2B6ApHqqEKrSwfx3hUtzP6mxreco/yHdU2s05GjbjRoCp+CnQ4IjDA+TfDPsiP
9xmhKUp4oSOFR/JVRKWc31A425BrVf87bw6puPpkVPXQhVajFuFiABNR437hOY0s44YSF+7YzUQM
KApx7/0gTBYyQy6EIffXPc/FPn9sPabEaywxpJX11FuHkLNHs+KxWPkAMm4U0pSGfSPHcMJQMsAb
3VkHTM8Zw06NlTcFIXUJuFtqogF5FYN1Ev3B1+PHM+epR+V0zZJaM/Wez2UdGv6YPgE2QzgrNl1V
DvMgeb12ZPU7GYnPHHF70cMANMpgmp42sZqHcEBgqsLShoyjDGB92h7ZcQyiFb+45Egap0ucYCdP
pJ/ohuDkc5rusSV51G6qtsIG7pRuVROs2dl+FK1kvBV83TwUwMsb+yzicLg9kw+pyCDFLTQXwaTA
6D9E3KaL8HtUQg/rsXkDcPtrSKf+JNhDtHQtKjGZwGnWkXAIL45zFkUgt+qdSEmoCxw6OxDakmqI
ZBWAE7K5RM+FTxZCZXGm99oaPvWgxVYtzDiHEJtLho2KpNNw561pJpTz1DdwdbMcS/6ozPhsvKOZ
yKLnnzVPna2CEFY5TOMYVPg1/lBJAOVizEfU6L97+3B7wBHkWe5ctPZzaLvHH+aKGGJ2wJU6rDK1
xa5/AwDTTj43CL8nOHsrw5AlUn4hg4qD1YP7m9dzNAETjbZlXHOrIn6naQX0LvOG1Z1r23cwO7ff
a0FEV8qq1Ro4gSGpJyaOYllsXmAkRwunBo6doGnA1eW4lZNPrWneWVHkfsdHJ4sRyooyOVi8bntV
FsVsi9bdBvMkeZdYtoYIoT0ndr9wPDvLmb/qE+n6geIskMMb3LOUeQdhhL1M2rWh9jVb0OXV1fXK
jjw1LTfUnwOr18w5dWe7cKErWe9oJ7/SPl3tNMfU7unFz2+4Ng9y+LxyhABJXj3V5+lEXBOjWq52
VGoHmI1A3xqaEQvp+JEahmnd+wFXidDUwOliBoxSz8owvO+Aqke0ezfcsQitEafFMFHnWWfYjtRR
s/lg6eJAy++U/0iqlvTa7b+MUwdyePan9354bVhHfGQ5IObvsNxWMZnhV0hP1BB03y1G4Cb2y17I
fDPTyt/SLzKJI4B6JOkOmXwMh7KGurj/Afp28tQLeRCGMqhXyB4LfT/kRoCmo3ycfX8IDeKw+lFC
6RxPBX1b9OwCHC/rL0cpoAfcy2Cla9p04lvvBTg2xguwbxnhkA8dANYrGMo8NKrKu3H0puAnVG7W
LIi5GKNHetMLEOjSUeba6G25dj0v6albNY8UJL6NLb52RladymzntVhM5NuCc0DEDul2hDxTfd7i
eR6O1hw5kpU86gcfT6eS4RI/tZGWtLnGEsofeOrPdWC58bDUxlyoG8si2cHjIKhHn8gT7siaqgRZ
fzubUGh6UOtJt1/DCtH+1sbCaYZ88TInXMQ9N8bNfvxpL30J7jwOD0BmXQ9TW2TNrPhTTq/eQFaj
nFIzfELDsjKt1PhBldgTBekO+nEulwK/WYWwo9GutEpNsLQev5yJjOVFnuSJSlT9L+0gxbZYBFs6
uJgpcbodtXe5+gHumtx+TCBHACc1cSedRl1BNLYq8K+1Q1PDgvgbijTAB9BcX7W6UA61afvhVbzT
T6rPRr5Qxb8Bg/ri9goc7bwNYiusD+L0c1LErQSFvGekBfefFfIRi2dZSvTquHEVtom2we2yPKgW
vWNgE1zB2Gzv/68G1Ww3LvOpQEBphaFisYT9LP/y29EtdjhhTbfHyZeiMEuDz9OCxTA/5wAXAfDD
uta3RSZ1t+RAEcG7UWpECvlYgIPw313+JTMfeb8HEPjDo9nd8dBlgi9yuS6oiuhEN5vE169o82Ke
cBOO4ACV4tIvznUnEo+HXUlG8Zb+NNtd+0rpuj0aoqcnVVg0LRnlPDst6yoOExXuePox0PHmneWG
mkKoVLNLWoTKzHzLqsOFUhpulkg4QU6xT2rLJw10a2TCdR3lyFoS46J20phkNhFuZiMdZUfrqU8f
AA9Qw79C6Qyr62ITVqPn4I8bNZt8OYdLlwgiiTdbQA1n8fkyhMBle8xzP6vH2dFip6lrAy/l5C7x
Ph5ZZDaLc7K0l13Mxc0HN+mGHbXFCzE99o9mN2xicgqThUJH8EkAXL3yMIvJELvBmRplJXDoqoel
1Rnmk9SKaFDy6sqPqREHT+pDLPqxgR30GpHKgPQhdmuH13LcVy8OC5649gts5BEexMB3LGgDsxKs
U7x6MT3GoaNL9wwb+2wRh+CO59xxNAoj3/HREmamsQJJuJ2FW2rQBRjJ2QYkkfDBVJHCeulbSjoi
LZeDKTbNY10ZVirL8+YZQ+aVQNHuG4tMcBtT3zPQwG/jNPa1L5vzMwPBhW2t/yuJHVdV+HBsKw/w
Blc3qGizhCGpdN/4CTEz1HP4vrscsm/4jrz/BOKCfvvCI/kByxK97OZjnsldWgY6PzbSCIpdS6vX
KsgZYQrgQnqTVqsXTVX6duL0AsqfWAxm8Fksmf/J5dieMYHEiSJx5HYqU4QRR9J6buvMugAvDgs8
zJnoomffPxcbAYcZNuHxMDbKMsU+y/9WBNli1Wb62CZzciP0pTfKvpHt5gpm36fPtJUUWQaEHpMR
u8EXmqEu5VMiotRRZw5hK1a5ghEY9oqDFNRj2yYgxjhXfgkUf8KM6nLp6XC1jatwXLpdoEW153x+
l5PqKnzxbDcBC0B7IXaRtx4GjoSspyofbeA9HI0BQVmA6tH7xAdBbpcfmvhHSu5V6Ex4gpWcLwQx
7TeU+luE4vD85+q5koE4YPFgqSwtFZLDavNLJXaFal7tW6mbVYOHAxPqZobrBUOB+s9Ot0ckKJIN
Rq9HcINUZwx995rF4Wou5isnQ/2hu05Eld1u3aQGZYCD/Mw7loZ4/eb/kD6f1oqv22zFK9Ox5eTp
YMyl5Jfi8+noUI2ixjr3nwr30kU2pPSIASeEV0xZPMQaaaavHDLDFiGVFsm/BxUg8WnmdCTr4nM1
Aah0jbxMjp8ORZk5hHLerkAMf4KLogJE1hdA5F9D/UHjK73BkkkMb5bhx/9/mc6rv6m3VmAJ5/+U
EzyQ2e2hXQtZxW0DUnpfJJOGHfKNvPG9nRYaBOg6AG9vn+Cma+Wdm7+JIlvA28zci4jeb8vLqDe9
i1+d11KFTHXmzLHnTr3xskvccno8ROI0k5yVZB0YuUi4tUC0eWZ+Ribu+6AL6t6aB/jYhKnViGCg
J0QinbSdoUZxZCcW2LVsUmeiRApuVE8WFE2NVb7znyiDbfrczVSJwPz/hMaAUnKmokuPCqjNrxUc
iwB3YuFohOfJ2qdPlxA/b5g38o84I2t/1VnKVEuWp+SzO4SsLItPDx4DCyBNwvj8R1HrR5D6BJft
x/H4AFZKlEmBIUuQH2AWbRVPGswFlOSa5awq/MvSvLdsWmt1/h59oRqDWG4aYPtfCCy9hSpoBxSO
S+XJogAUtEwm9NJhta9zD9YE4NFL3GuhZqD5bLH4n2gDssaTE5WMxAe8uz27iIcC9yLAHBjulETo
aGMRAbKJ9t2MEdu9PdgI5PY680u+hbzHutHQu/fb2Xq2r0ZX/6Yw1AO318JTACVDE1tgu9Q3RpGP
K23t3l+4b1tSqwu51C6T6BIeX492ixj7CG73MXPvqnmn7mevXA13xlU/ckSGrvWPqqbY9y+xZ2Wn
zhSDw6bgzDYthTo2T1nvQ5EkZK5KP4uqVuIqLKPQs2Gs4ESRXZVEMOo5MGuDbU5bPKeDqmgYBHnT
8t/+pO20B3KCLb5FVs4/aEQUSvklamPTSeUuT9axPcNlwWy0iCKPlirEuV7qUNsVzJhGmexSlQNy
ao/Eg7wcVvnpZh+YXjYDMYh4si4i6Ci9kRdqYKkFqI9P/za2v6xYeWZy8i9kPn20aV0oDbIjONCC
zSNNYRfPrcqSPj/TGIczJv/aiNrLd/qtKoLUb9xeSzHaJrGCxqfzH6ZbNh1MMISUyhaheYP/wNcF
6jG2EiFiJbXTVHBsbnx7EHMXRyrskq+OgsoUVqiiLj9WTnMQuY6lVIy15axeL3ZPxW5qfG7odYAS
wcf9SsKyexVao6Ud57kgF9admEjp7S604EFfxLzPZwn31sCx2Vaul7yzzY5YiPEx4148luCZI3GS
EX8IyqQTgUa4AYP1bmtRxoTDikTpuoAM7NkhEFkP5JFyPPmGsRTPOGxdsXJSQdcrwGb3tHy2afEB
KJBJFmmxNVQf7+65C1chqxhT0Zq+RZiuQkXqQ4KOS96nmtXwqd9zQj6CxcZfWRHIV/R7HjRZjrb/
E1gDXEyhxzzWsozYjTxNj+HNcPzNSqJO4J/WF6hhTQ6VFKhjqXxK5IOSL9nVc3CjCdItdSFFU1vO
CBMkU6P2J4wjwfEaH6RGlp0WIs07hYvFhZpN6GnuH+9pzdaOuJsXnUTFZJUyCcHvMtYXxtdp8bOK
w0Et4fU+Fivq0LjHPwBOMrtZF79C6SQeZZus8XqZ7OUpjh/fhtbV8i082bKKM293glrFjV3nIOQs
nu/77/XneH2pvrU1h314Pr44dDyPRVG4/pn2CVq+00jILkSZc7AIk5DVNTnGvPJSoJPE3Pl0aHEg
/1oyRfYlPMuA2iQDtji/NmqF7wheTZ74bOHYKqjThP4Cu7ND0sEz1aivHc5WoI9amnKVp8mGla3p
Y0knRvhTazDOK2o6WTrhndZ9zMe9+ODejX3no0vsw0Mn9BuSX4O2LvGZxpOY7ujT0lwq5NztUn2g
DE3Ra0ZHlEjm0txM1xH2DUTm8gR4kX1e5R1mnmd4iPz0KEXEIHlViiBQGdvjHhRBYkC696+ycfed
B469Vszo7Civv9Akj4TynLo1w6Pf6MAOo8+3V9+5w9xgOYn/L2Hq2riODTPigAuPV7PMe6kKG/6K
KweDwTIUJNmdy86ncqCIT/qmvJNMYSpM5eDRdl/mxYAbZVaB90eT+MxmSTukAppFy6r1V32dm6my
QI+S6+MyGajQpkytFcGcmOvGZbLsDbpv+PMBqrnmRiWa9MLOXfuOZZjDt8vVkkXObMczb06039UU
4SBn0NeKlTaTbsNy6ulEWuyGbLHSUO12vZjTuzVVCHHkUGPS3jKiHa1f6rjJzboMQEehKhSoouot
aL4NoLUt1DZISr7oeG2INe1/AGgXc5l0suhaCb8It/+FVl+iXs8pihbr3M3ER7w6Gjq1Z+F8+Qkg
+3pIpjSvV8P9utTizxZJgJsvBl9+PTnkYQP7rqNQ45MntOnwb7cmLrs+r1Y8KnyOAZ6f1LYNVt//
N2Y9+nuDVW4ef3HHHvJqJHvOj9HHhMIMpPYmb9mhwQpAptyChh8Nkv8moqzEbHonWRJFIN1ZilOm
V+UvJJaPAf4fihrVsuhRTLXn/rOIj4AYoBP7kufNg0bqOP+aqmhR+5pPiOQBOTmthsip7hlUKBJh
pZ3lfCh2B8ljdQ7Rf8vYcgLKxQKfEQYJp2BccwqJRhsTfxP8ffDlKeY17uh3w9OYR9LhyQOJFcM0
Oq7S0GAchq/RRF0XAGNyA2jDyoBzBjYRHnGyWWZl/NNateKpMyj6HDOpl5smUOPUC2YrMIpAbR6Y
H8uu/4Y3bpK41I53L0XRvj/tmBYSU9puOYhbbTqgPrdTfUYE58MDV9uM1MNMFT0qmJphrPPYI+Oh
KT9blYAgpsGL+DD86r54YIym38Q4FBPGzsD90r8PBA+tX5OwHtCWPE5w/Obc4YVYNktt8XD45mlO
MXGdIwh1c1p0U2/XCZnvhlwD9jLhN7BnAsJ/1UR+OtvZnVjlykUftNohqJbsuf0/yB6DgjLq0r0z
0ORW9ii1sRdwgmWgeLXMNd5tTHNHmW0qQkfwnN/yAa0yOHPSusDU3l/VFJpaeeR5Lgk07Pxxk14G
fBuoNmJscP+tq5uiTYm6jVsYcYbBO++rUwghI191rzMLbd2y0rUM1ndZ3u/km7zbmTD+1CZNnEip
Z8sp9BaJziKEhhXRr9QBu2/ZxnLv7nMPQZAhxxZNN0huKDIZTd0aI0AlxYo+11dWYOIjWVGOjcho
vNEaxDy5K0rZjPA8lbIxIANuobE9VLuvpmYi5mvQy7IHNAhXFFVIeybP9Emj11a3CfvvgpoPm15b
ehfexVRYp3hHmoNQuB+z6dF4B1V6IGqk0QlXlfBNLzK7nM4dYQaFNjxbRKd5VeG9Z1INBBJqfk/G
vTPgD/5dVy0VK6x112L56ZvIiTQlGil7IU4iEWGtKa4XvaJ1MyRBdzPujml4oTZOf9R6HL/qF+UE
luC4rb2a0Ig5H7U6G+VHy1aaNYZDwu6inSmkm7dzFhtltX4dXU35zr00NZqUVP/xLg2DcxebbkE2
wxusvPSdFz7YeQz67geY2UFDltfMfTUPPcYuUEq9Bz+JGKXRgRcYu5FyCgNZYlvDwgHyTyXafu3K
f7vza+6FK2k+02GLvahjUYeLI3BzjdDgi/ctrr4Hogn9vAPlspNurQbuHxwRPu46XsNXrAJpDMom
BEhIYVd0V/NlTU5PBHoRn1x2hVCWePb67qUVroOnR7kJlTgqdutxb4lyy8blOwyp0EamShNtUJ0H
iC59MSQLym1U6uruebI1aJqR+a1AjM3zKcHq/kGfgU35GHovZmel1Wvi6EGCL/pQ5oqmz+lJ3D6i
9Tm1LiE27RVjqwjZy3US3MP1ScIPI3v9XUhCpfIm2q8cm1zedmu/WvBAF4RNUDvZhzeCKUFtHisa
BpaTpryUIEvskBPSYjBiX/8SgS5OK640lshScvRMloDAg8fK4iLBeCJHhwR/Bf1e/9QBnPcKKa0d
DjqyI4gjqRgmDgk9tdNybkzwGGL90yial8fCN0yVdOLSPeqHhUZh9/1wR+vL+FOEBlpObf1VJeDP
IsyxnRxM8DQXXOpQwGuSR01gH3Nx2QoY6w6P1vrm7rACaff/vu9o7CF6LZSA9LugONL5MiUshsEr
OF3Cy8KXY4FIOaAewq7reLosC1AzZj+/SfJeQpJYbscL7k8hk0GtxfG8CFJAAd7I0XHL99zEU5dy
Vs5k+3pfshb62nNtLqOm9xfWQNlPTOKmdflQxdANbZ07Lx2qqATqwSiek8rQEjdpuSltZyeSTcMN
kKyQdmM40pARgmzAJ+/4qtnk31T/Fq9kBdFdGH2oSspQvF7I6JiA3Xrd7l2JtiyPpalBr4A541fM
hYC8oB3p8848Mn8Ur2zAwUokr1Lw1ZK+nOUNM1ZTVmrim2quccP6kS/33bn0Ha9sN4QoyW59bdWt
lJ6ZotTY+BZlrxV4UlEwQmMKTEbPPsyplr5ZLCPc2bgJ4lUNsN+FypOa0j/7G7NuIEOZ7k43V7SD
DqsDpkEIf6ShTpou6IZNS6Occ0s1VouV00qUR0dbyzgzSLVxh6aQ6Qi+GZnEG7eh9guaU/RYFrVD
/w7E7rfKPIyEigBlpmlXTR7VxXdfr27ByzZo7Z2nLo+itAHGcn/MzUVU/n4B+mp1/a1uY2bla0vu
tO8u7ZM5JFaeEpmaco+jRzEipvAfmf/6t5J1KPSqJOC5b3KnWZn9dVP0sQBqZwnac4ov98N726LK
XBXV3oy0liuriIF0yEqt286JhasK/VVwoSp629txiwF6wR3YZQc4bm+MM/hVLSYvEWT/dlyTjKHD
sgHtlnZEwdVlq8KU9H6v919FtfaUg0uynm64IPPU1X1kOLEYC4qMEWq9iWqM+/LZ/DIEC9pYFDlG
GgFOioz71ODkn2UNaYtkgtn8K+/xW2EvuOc1eqhA7PyoXOwwCImTNg/rOJzU8SlSzIUfPmrB0vTU
0MJASyPwXUetyXdnJ+RIMXsUD2IM00BMLTDIZKBnHWnR0WW5dMt0LYRJNKzJs3S59XhlbrHTtFi8
7aBOopjQtPCXrAlg7FE5ftWi1Kihj2EXMM+LKOgbculJhr69Ui+b8oS4M3n/fM7r+cCRaVndpFqi
NXs4/UDGQV40Y9tucJfIXPDxp7suowS/v5k6szhMqAKEAK1sT8BX2z2Rqafb4CdoOSUt66xImiJg
v2GxLN0h8Sx6hwumnhifNMh16q7AXo98TxANF9r1fgU5kQjyy0mvSLrFpxQqzqECxKiXAET+eu+4
IKxrlXY58qTJelaNYnSUkn2MGlz332DknfKA3hx2wW583WT2U3h4db1kgWiDr6UIQFw4EO7aO6rX
ld1AwsNaOxa5jEknkmTHpGQCldmJ5nICy8n1zhV8478hffHw0aYKfubhkmeOLKEWq4l/UWtGLEvg
2cdMeNNGYoLDBvSNVXJRHnzzHkBl3/K1SBvwvGZpSWWrHDwdcSku7B9vbD34efDz39KqVI2wbnHJ
B5ycBTsJdVozbA4NQXiHfkBxjFzFaiE16wgFMvZqYF9WJbfEpuTfmH9UaHZTFPj5HICka8zzqvoQ
47rh/7V87tBm6mukjNCifeSH0gzzM2vhtHqn0Vr7ijIFogdhLbfbB+7BiRjS2trLt2zy1Q7bqEns
GI06FANGWrsjtiqRTstNeppgo+xFnw6hYjaOcoT762Qv4W1xFgOvbmZR3RbSzDLwPdT8okGDKk1f
TjEUMD4z0utgYG8hB0snPYTC5JXG+AC3nEtAJLD9ue1nslxYAIrCthk3sxMGdyv5/AFtz2nmUXUz
Z4Rc5Y/wYz4QXLWZCC9geLuvJilo99Mjfs1rlcen3kyUco+Wfqy6Z1zLas6CeOepKSFetAxdKwXw
NVnBeEz3/iyiOF4MJovpzl9EIfrWfcNMCg/KTOGNlGfBC0Hx9AlLuHmEwrKc/9/Dygiycj9F8Ull
kmTZYQ1fIYdYMslqW9vJJ69LZp2yRuMnsoHJam5gvIlevpD04S3Ps1tm/tEngn4+HsPaFjGGDt2r
XCQOMjCVkjw/SFegUmQ7pUtx8KRXtIyy9DAxzllxYfoI1jbsGfP9Y9jly8arruYCEBQK/rheATj1
TOUBQiioTT6H9NrBBDyYu1CHvxmgS7qKykiEdescbdcGM6EAolDgtPwS9JuRk3n8XZs0c7pjbLqt
ZydMIlbaEi3JJKGMJuqIJYkZbFm06yNcLrQ72WRJoKLQfpiZuSfl7scDTKCMTfIuZ+qiFt3cXxyt
lM1Sr0WrsV1soHCs/PHVRCJ5g7yKQNh4IiyvMDjyRjtkJ0Aot8R1OmIM9+ds77XOHumy8lkQkfDU
4NEiSIgNqyQtECTBEsgPlhihKUuV7xlNtInhwlPltJ1u/dTLCj6qmi48P43/rF+wQAifJQxzrldx
nXGcgg9zgluHJ/OS8jU9RaT6HuCdvvMe8nnO0dGJe0EIPWoRi8GawcGT43TWnXedHmTuyLyN4OIM
uGlam+q/dDSz+sHC36qeCfoJAjdedEOnpQv6/95qadPwLmXH0Cy4b+LYywl+F910Qf5xRN01vq/c
0gdkEliVCqQjdrkyDKxCjnd7rEYkZKbEF7ht7FD2xPiJ8yALskR0orMqHu+NIZV6iQm9AISq3bsu
dhkryPftqENp1glOshfhC0irH0LgegrZhhJXvJX7t8mmO/MWmfSZesmCUPxxSop6m1Jvj4kdd6Bs
t7SIE/ZMKmeiQ3aQhAP8MrgxqpY5cvs2FoIb9z0Tldc+EMkjFwaUYhYk+dNRgrwQFh4hxirZGkaO
b8sXU7XSZT/x64uiHO8I4SN5fVC2se5rvlXAAr68sJKAxGUoR1eFVZHOH97rDTOFWgQuM+crnn3/
EaJfFeiTHqcphEJ8v3cf9wJtJl5SvnnAlVQ2VgCG5gefzsRBlnYESyYJFf5lIc1CkkD+bwetR2EI
jAg7evVmojuou8tG7eAbUYk3I5V5j7ZB30ZnU3wGBm//O2xY9MorPjzTIEIzkf4ef5jIkckHIwvD
lpVNcqq5W5V7O/jgiR/ospOrEEItcLPsgWOlPTO3OEhsSZSgO0bFv69nNdJEeAgY0vpxIrOX3hIm
vFi28tO1YieQ5rmFIeCt3YzbsnBHASdBk28i6Y+39mwYz83Sm+FhP7EZH2BIc/AlwoKByoUrdNXG
R8wAP3OJgk5LFSB/WQesTRTp9f2qnAsLNcROgRsrOf8i2fACSTRb9BPp5DTSxpwdEnTzZQ2IcWO0
3mzVUyneoND2a0Wpy2QtPMr7R8erVNFJy7an/G6X3QDHeZRYcfVwK7zo0U1CDiJtzK7oJL/wLlqU
Sgyb280UMv4HnYrJgZlpZKtvvkYlU81DihEw/JeX6upxRr5bNpWUSOo65V9Tl62qrT3P4wUtBKOw
0/ajIAPfsdnetoRYWpKFH46eb2JlNJNCBPX6FJlQbUGQroxQISr+L2eGkM46fXsYM3YY/fPcGV5W
3Q2Z6k2kw9+33mt3eu5TN1Cvc3m8RKsHbgNcGlHElzD2SH/tbi/GFo5HzQTKG/3xnvoMmGO9Rmf2
ZcrLe+kadZfAqjgn3blzoxqyWc6lOvwvZvVZpBiTzpX1MzCy2JDg7Qh5VQyCccv+L5eXdCakOjfn
DDofuPAy8bqsGkhxUSU800pF5O549MUmgubdStNWy46+9NBpUNCt5LNZJeeY0vosCAus1fjn/KjG
ppmNE+5+2lyoU3Sicih0cVya4zy9NUD16NcuH9NSkPt+CVf2H/1nMmUmZKFrm7R1gp3ccxYjiQvI
y65x0EhtR3gsv0P69QHTJt1E+BbESwBr5wr7xq1RTOr/Gcgw1Q+zraav8qnGMOUDIK+2m1y5XJ4w
RLr1e30/WbZ9J/6tFbM/lNcRsmMBNHtOKgQs6OrpVM7sDLi1PI5eXIxBS/W6EaN26tQoe7GE7iyW
NMIbvjJ5ko3ZzxRNNl/Tf/Mxds5PK/L2PgzSTN0zbkQVITkwOw7iCEd+YohNFpA927x0yGC7qLju
r+dvD8BLznRFX/x3bRkZvLIvY9MO6N9T8LUNnc8fuybjGPzY0b5NmVAHpfoQmgqMItZ6buNlnflD
jCvFlRzG9S0uEIgls9DhHoQ6ommX6p6eyGsTyjJmUzu0/mIII7wxN4ZM/ha5bkkV+wIjfeKzUV+s
+3G111ZoeMMh5fWRrdm3AO8F9tTGj0XzlMUMmY9zr83/SAM0Ia2/q2rIbH0NWOwAPrczkURMllIB
mbqbhVe7WgSujw/8KHbQVdFTD/WagUTdE7swD5fXGIRunSQCuOj04JjEd/oUCsTHRhUXudyALn99
Ghw2J9OIPY2YMwn0588jc2hiQoiCCiZmBmUh/EXEsjaqZ0aiPt5tCO3T8CH1mVqKd+Ebodl2aKF/
C9TKeHMfd00LolNTdklnUG8mKQ0XCMJhJGXcxuQq1/dUeJrZo+R9sS6ES+3ZKiKde/aHmVclnX87
V5DwvFQMl2krTL4+RfKKAhmakyc0hBBO9+08I/DASZI2HirOY5BPFpt4EAe3qDl2L3mfPgi/wWvx
3UYlQY5edLvJR8bJdMbpjOY8OdVu8oa2h4ArGE1mmU/pA+H33Jfr/76aZGoU37VitkVpTB7wxP08
m2uRprNvKxFJ7OCbE651GWwOu/nUBb7tZQNKxaScMGVIqFTU0LT2dWlgarbL5pebtyNeKA3/ieZP
m+FhrN5CqSrZoppsERkRAFRRUccJUglyQjfoIb5J3zWrKHgepcus+j2U0u7UJht6GrBbtEX5kndi
qXCszOUrT3HXEeonFK9WWp9VwdFduLslAXbB1dOE0NEvkvmvhtRR9ixNd3AyNpTdRHM17c4Of3Lw
fcn0+l2G/uBXEejMjNqEBMI2AjbUyfBEGfdvKweRG/aNfADdiGGGJdD29i08A2xx/gZroMPDKWfR
p2jp9FhURqfix5ZEuTXGC2uW0x8YHIsvBie1wHCYSoOuPoMDihlMh9t3LhaVV2aJCKjfCQWnIhrR
qtPnZmDSTdQoSoeHFdH8rG4GkqSbQ0brywb+5dnkBPvcbhi4dHBNRBPOimNiWERinqL8EzZlYq2f
mlmiU0GzeYLdGGj3jVW+MI7s5jkX2TpT4iluHuoPnTZ4k+z6GDoRnywIaC/7oL1GsXz54hg8vUg0
JjFkYSMGjecwTufUtYTtQ1AFIVdaSDiNCeyJEi1lQtNMnYRB9rf46WQapl4ndyv6mbsDU6Rl1rig
VYnLDQoAN6omddj/gJ+57pr7quy/asWlZ86EFlP/AjExSp6aOeoQEJ2t4ZVYy9Ol8eyEGXrPfpFL
KLtoZxTE3YqJxko+upDlLifWxX4pUlC+B5nAIqXIkInKJXBDgv8bUdc8JjiOZrRh0DiI1Vjp4oD8
GZiqxDFulS4f+7YRhx2sX/APtl7c3oZ8pCz5UD5CPOhqR56Co5o6hu5Gi9QaeIYTUxG+VPuCIq2t
Bk/pOTRuffymB10ro9D44A4BZya2SyQzrGMd7KY93XlLRLms/OR4NtsWrjE881V85rMlJEop8UAz
vsJS8H76dFbx/cVVTUZXCp6T449FwRi4oJbBayJgo64oQd2HsAq4bVzjB4M1UU6GB2SFbdTCkJz4
LEpAnh90IXjT3twYBTdXBoCxzailHV7YpUht7kc6TSVJDslRaN78kCm6ZUAyRv5ysrmIl+qoUqm/
HZh/pth9S4VnKVnR2vt4UnCJLQ6rhYOQ5tXRomFaPmf6XnNFwEWmykI6QIHWlCztouaFVXcU50c/
9yqTrUpT3ecrTNR82z5cYCxNWjmuMFxBueQz4O9EZvNS3DPmI7KxOvR5IKt/qOLVL3NVrRKJIIKV
rB73MJ00qJJwGXbgeQMfygdqGX/JWrjTIwLDG2XkPkGaZsbF8FEZ3fPmWkdP/6DXyU6JRDhXkL1n
eLyqMarPIbOuo05OGks+lERKlnvoeBQL8pWA5c+mYY2c+iXNfupIpQ3bk8LrZbHM/8OrR8Dduzln
r5zpgze+KopjSrcy7EA1tmlzKOEkoevkkVXIg+Eil/gAd3O65UzbBW1nFZE5TWnbxHP9T6yj+6ij
xY9wkEWVwBk4mSs5uhmVP2VC/i9nzZVzUv4d8FWCQpQY4I6DIyvHg8uzYOCL/rlptWHSXLRAbE0c
s6XYEBIFzERK3AJpKhPb/MEN08I5AvAa5pi9KRktJJyFhscEqQBpXAwJU2sX1GANmagNQTZfAaDb
/Ek1T0RMUdn9KY9GR5bo1cFE/XCZEEw7huHyDEMJgCi26mBKzhc+dU6ZiSe0ALr3J8z44nuTAGWe
A0HaqxEqa/zHmY39qgl8RPImVRnV0xy+aWOGwOOHaMc/b5FUUxI0O+6TBxr8x1AAfnPuhFC+nncO
rCBerHLo2scvI8sA6Z16TlEPNVvRWX3TSBNKm6/6Z4uENHqUMYsa4RPyPcgL9jnlJA6U/2BeZ28G
xxJv+xflKR+xpOB8q9WoaYgecbPr/BJHq7GeepaHwB/EV7g1HEM1oFmH9dyBLLaCAe+fj2ifirTa
bgeeZ7QqO/PsR3tcgsKsUTjzLtWIgAy1zg7QxYKiEee/tz7bUQmkjZPgbFnHJ7RiUZL6vOWi0+DL
nj0yQ0YHFmOqEA92Qx0RXHBa7OtVbGt3MI2+OxITL61tXOvRccXCppz2kUAu8gDGr0jNsYvO7ZaK
KfpjmZfZJcISvtaYKnBqHXxoOkqbmLNBE+5n0MQA0sb5+t/DGHmE1uWUTU/dUzja4x0Z/cSuPV5X
R8AmHdgFG0Tmd10MSSOpbRmnzOLEBSLnwS3oFTUS8ucwyb+BxrePzOrAVxAg5O99q52LTXzX+T6r
haUDsgJcRye6yq2j5LQ0YzofvPX3LMaQj7hFc4V//LuPdRcxrfFYnCVh9OmKqYT/fUlByI1kj3OW
0x9umPl4a/LC+YAum8njTzYmc32IgitO+t4f6a5XA/5MKRVy2fWoUy57C+qRq60iWrWGjaZS5eF4
IXfhKfbsc0/ChskTXUj9P+OhTUNOr1+WfdErUU4l4diQVfhpvoqbInOi7w7Gfi4fUtFg1JuQpgx5
zkJk4LpSeuKTg/wGxqiRa3YpO+K7wPoj+oNzXngBpFhC1blHWVdJdKScF1hGLFP9oxh/9RSAs/d/
bOsVAMtrXKMJymvJqSliIsjroriopKVuidRzh7fmuhhYi5AEzjJuKEEgZBwq7dwWA/oNSlDCExYg
ALVKwNxiIpddK538tnuhPjwtgD4ECX8nVitnozTJyJ1JA15omdZJ/urmrdmymVf4JbVcrj5EwQal
0K68o0Zg8RRJQffFWSuTZtZFD8Wh8kW0BesGV8PGsXrCcK81ZbE1JW9xW58fZ8P5v79Z1wBzlbgY
l7N8zhZRXqqav5jDSbUcI8xqgBRS79f2QJ7wrBMs5SWDTxJDVkcYaQAevxpMP46DadKQg3yjPOUn
V47Kc6eaTWAD6NPG+oZkpRjw22I0Ppu5BsvPvQUohhtIucIWHNxASi/LUmMuhkPVDLce5eeggRnh
jfJUAv4xXdnPHY0dfHqpxdvk6pviuX1GCDusa+Rc0IkwBOfoon5gSjP5WRm4BiHMep0JnVtrr+jF
TDR5QmfKjzaQuFbxFLCWsNykjy2+yhBviw0hJnoSw2jeEqtn2D6sbcIXMeLm2sCSzfj9x4agKpW5
pERjT1FJomfWzrsf+6Jkin/i2ddcXdnIjC9cSV+cPQZ8FnzGYWMlMRvvkwCghQdMNXuxl3hWLEnM
pvPukwLMOQdWyYdcALkXUndv/tFHCxgYZz+Hb+0PbD/UnbZWyIMHSYMTnV2B899Yo/JMR2jVfijV
SjK0nPUyxtb68q1Y7NRx+EOdpJEQFpBMOrO9Qam2pZAJ/o4qxQ143FA+QtY96d6eksNM8uqQouEt
6MHJQM2+2fYsewh8BWs7kIim5B4lvL79fFYYSW2hD8uxvE0JCl+mYBTNkButUYqkIoiaFpO8jewQ
1H36PKvV1wbAY9XzdtKthr8CTgeZP2nM/hLaMw7HyV5lxx30KFqiBPb6/beAq2G7p2gocqXRXjOK
c5q2NtniFyczAgwwl1CLQwThHSmISA/LDySviABhdd2KSRxnVLYImwTxa7n8SUB8mku32N3bCbNv
orNho1oA/MpdzItMvfNQHn3OUacPmchFfKrhjSC+kEsbwM2WIosShl4mUx7xT1Hyks/4QXUwWx1n
H6HWXN1oi/JpqjP9PJs4X3sIyxFUSw8eI7K9e1OKsQQE0Rpr2iZ8JtGG/CRFW1UTR99vnyk4go7n
nkkp4l4RwAI2vYBPF/kzSLpt5kg9ylGpzLY2V6AW8vWy3O3EoLxOmhwuCt+nXaU+JxMpIXwKZ3Wt
N80C0DnGBonvIXaqQRuZqK4c/ZJPlUyOvTQV+ndMg85Dq+musDioeycRv2WR1VHnr7FA/O00/4VY
dIuQu10Guee8yIYmteeKLDs8HeOGD5A5hYkwgbBc/mwdSAtlNmlZC+cghH+v0VI58nbJLq+DYCnQ
znZn5QV7d8tH+e0d7VdxUrUvET6BjORbO7lX89lYdQs+2uJ8M4iNNS2/25aTpfva8AO8BO1luHzX
HNWdDUv6U9cY/F4YLPb0m/p0Wkchk5e+F1BFaOoGvwmpaIiip186AygEIO0M/EFHgOzbEXyIuvDi
AndvzLmeZdJMAAfnuV4jBQuYfG55sLlrW+TXWKmJ3AYscyY2hTqea6QPfR0nYIkCEz/vzXgLMMfF
8fj+ujKr7Zwr1fTXtEJ+8sElE9F8iO4bdpMR9rKVKJ/9NYLF+bIKC4zEpZ1bGBRj3Q/znh1vgIBg
CkPNahTFx2TrKBUtBfWZwteZrIFimtLYwHxStX1bCE/nA2KkYau5K5sGQ6nHtQH85gBCQ8EBUagS
OE1K1IwsS49BaGTjDb6DWwbSA3ISNOy9Sj5Us3Ltbz5YwZGlFD0y0x+4p0+sflw/cO4f+04QJgw/
FAocMJ0jWv7Ai1HMqp3ouIBxgcPWZGXdH48uXXdcscseXYMJUI63Y+uvjWm5fOQeoCV5fP2xAyx2
WWLZJ/9Nwk+Eoq8TGc23bfO+ZnaOoxGlB9BBXu4UOw5xX0nPpaTxeT/nc73EFuJvIaTCvMpQKGxK
4gv7RKUFepIc/+FN56ZLQTfaDTHGSkmUyjx3wD0YoYIQe3rswtMoA5U9nNTEB9d5X6wM3VhiwZTM
PvMieHMaY0xm/mUUTgUd4ImgfLaNOW6UWQp49MwtNVCFuTF7+yoZFUdn6AXMejMkhfGoP/e4yS8L
fFuZXFo04jSTAaWXaHv3TKVZ712m4WnKUmI2OjB6jEu0f5ce9x86FXVwhapg9DtT/JJSBbWk1Iw0
UyycK524wL6Euh8olqLLRPk18VpkYobpWww3wD1Jnje11pcoZqdoTZP1l0j9N6sNTlXY2GZahxJs
OONjaxl5oK/oXuv+0B9MytDryO3oLid4XDBGNehHwusfxDo8UXvAnOhyuQp0rHQV0CEKHbh31u3l
Xjo+baaxlsVWH1gbaBC0wRM0R0zr+h9gT2VzxrkGAXhGUjbtInoTX5ES4NxgxjVmSfL6Co9Rm5On
FWMC3eXfbr1fOedgnbwngHdaSs5HoAoKvnReff0DzYnksCPyAWRGjdfDvdy46yuoyjbcnZzrt2ZL
wUwoZLCIEAigVt+aTDJM+ICtPTeMf1BtcdJpbGkFksNreriPZK73KvcTYvtWO+IGOPs6nldI1HDb
ys3O/+hDJ3SItrzu5zcx0lZBBsBPkrU5cewZOlazJOWLY4DRoGd5czAFcfa93oSQyod5ehzz3t+e
4cBXbwyZ4yADAlqAPjbpFo+ar+Fm7tmUoUUr5qMaQ6DO846B6ByVaMtyZZJ7KyJkuN89ZIv9Bw2e
TP1uIPDeBlVEBzwOD+18TmsU2dN6ZRCff4bvWSLcydsPVrREbDbn73LDZm0ODVKKJYJ/pT+sO1n1
DvZhElQJUvQQ2v9J+QNaG68evACZa6gojq2jdrET3hcKCBGyiOF8qHrcW2gd3W176Bkv3FI8CzO1
ZI86v7UfbNckAqScJVhNhUwoHWRj/LU3FFMYsIK5CXsz3ZBTBurSiMnm1dAC+Y6rdA4rbY3IHIcq
/r9DXl+5FzxC6r2XQGsVbju2gpCNr9Xj+KMafOeJsnZKagRGi9cmEUfUJfVBJxuYDyB4y05IFbzj
06SxlNGUewnLIG8u4QczaJB3VIghy6wVGnX47h9UGg/REI+DOWZWx3Z99gXnD7uG3loPKeDViuoU
SBc3xeC7Pa7tRdLU+EuUTG88x/Q+qXXDErxO+c2EI1n/cWwJvz45hCzoo2kfINNLsl63ANFBgDvv
8z3vAgjsmfK20Izc7UEPg1rphsbNrdV4EaM1qcjjRGEafEIfnpW9IiwLF7yP8/rosEw+D6HMnc5C
jpEX9rkDa81KKGxxVW0fqjD3i6kRCD01e8Qol9iQ658+ZsAg6pRk/JfJwsX3WQC1X2KELnrTCDMF
fTB5Ad0VUJrA/KWks/tLIevaKZvc7BDWg9GZygv0JhKxyjS0Op4rwpsbdcwayoz58rsMZ3j6SOAx
57K4AzR2eKY86Sm1x46Zby9LlpsEOV6T6bIb4l4/OglHDJfqFm5JGFwKsjWugMKDM0TiHFr+8qHq
NNd8bqPPZ3ddECqPpAhSZ7+OfqYJ3ut+vAACrVlVDYPPd3HDCDlgA+yOEMw6rtVFt4MveocXfJDr
uMrBeKD5JJbJK2BzW9ICprErbb+fh6evWpWj21lYqejmcSyDDz+EUhLQHZpFGEwHjW+rddlYaWZb
8DCsWXAsty+obpD/UX9wpCwcBH0vNaFZaerI4ci/IaGJ753f2NWiXIlFNQC/k0s7+4v3rg9VxeH0
lneUg1lSbcs90Gv9QHGSDH7rcayCr/02Cb+sTK/zIlAC6nW96fVkWD3rEyYg2tVPktN/YHzgGkr0
/ZxsjpL4Q13QdUQAVoquGTE9FobgwvFcXEoUR6r9HLbC2m+DA9WOJYoTOc9Ic7MvsaaGU6Vib0zr
G7BzeXcvXweonnJv0KVjeQujiw5Qu/nAdnXlipcQ50G7Y8Kvz1YUnzdgOUtJpkRr61ydUVcnXNwm
+gIIW5tdX7TiLbE/YBe9iOSjr4DmPSIaIPO+DvNIYEUZ1GCNS0xL5vWsXVuBrx9DYD9w20WFtDWJ
vhGviJuZ44X1cN5nSNMkxnBrDputi3nsQkY+3qJ5+L1ETrkiw5Bsts0bgGhwTh8jk893dNShaejL
b2mtyJS57k9iH1BZlDYIUT66x3duy4Yh0em1bSt4fAS1cNtej0ngGJrcJm2Y+5lHgKiVK0IZDrHL
QGn/M3XhJrESX87tM7Ul9qT+hEV2HdaSErBbve0YnIKj8Q3VHxbooFbrsDS8LE+VcQK1UFzX6mEG
IauW9x4cNv3XaSITQcKxRoXZnc79u+W2e8PPv6OPJhFITO7iG9BX6Eg5OYXMhcdWMaYe/NCGodpa
z/9/u+ki5O+DmZ/hErQMFZvUDpDxo5ZqN8Ei69Vdzyi+xcSVjlsRXL3CLilepft5a2IYhNaVArHC
TEjrtrhZPSEiLGJE/ma+OMdnRrTFiJT2QPZeBBNew1GVNXKLmhZGNTeR9X8gF44tqOC3xiqBCsd9
cIeaGVK9qucx+PvsknWhhzAmR/9N/4foLuARLeQGL0RPbG5c61BZg2qE5lTljF5rqdwRq31Xa+PV
SFvHiZPPmFx7GA9M7rKoZcTKhTJheThv++iNnRUwIo8BDA8a2S3cmIKiGhVotKMrZ7baM3L28BKx
aNnf1WYKnKhC87QCMvJ59hJ+gSeDC2aYzKi/ne6EZ5t78uSjjFIhvDfiqro/PpGrGxiTZWXDsuU3
XrF3Rmh/Dq7OlHkG9J+0bU0FVN3tE0MmBnHEqPhhYbaY59W49LdQK39iqRAvkoBLPAJ8+0C4CZmd
MXKFuU+BMKMAVe8Yiw49AhrrDC1PkWro1Ex0Q6I1FsusHL33ZW1Cy+XVLrmQSytw+FnAUjowM43L
Yu6LPXwVQKKwiHSrib+FmLzIp37LoOr/YP9N4UdZzAYWJueEBD6iBMLl2zOMQbLQfdA8BZve3uOi
r4SY2ODOI1qWxdgu3Qfpb0Gv4SpWo5YfHOfSB2GxjtvoLslUXTfzl+OGmMwGRGr/zNhVyHxVwOpr
tsK4s8+jPAeVHGOtm0lrwSRduQiZ/52d5VeD/FCAMgEtKwV58DNMxe+4HTDLeqDqmVsUyDaCnKeM
IIphntdPsiQB0YovuDZ13zjq0i+AVwHo0LVC3jOr/Ce6jU8SXjIVQf/1uMy+NzqWIpda1J/0DWms
9FXvHxIZ8SpdvCq5u7pafmTHydUT1pjd8BHjL0ipuO1EyZ1pGLI9Rsj0nVxvdtN40ZWlobyNjOng
ZWU8HaDosvCfO1z9pcHsoPmR0Dk7DWB3NBXj7f2DZFxNzQZqt/52SB5QR3IeqMTHNvqgOJeldKWk
tviQFffGE+NkaEIsaM0BObjE+GSuXV7xo/bjOSCgGfxyCwvUeNkXr1F5cYVWjYe5xqko31qHC8PU
64IUO7aHRTAHPCNJgYvSKW7U4GsPvgkwOwbnMUlARDS89rjlmYv2+MejfX9GFbFjla1hgGDq84zB
fuyg4dFGvIXzQzrxvFGlgFyjfHMMK/CHeVvhQ0S/yCUUacGd1IPr4IpzkCcwhQR3xDFtDW3FJTTj
gmnD/A/X6pciKzXfjnJKhJB1Am5DpvrvvACcZ9GGYylSK99CHXUbbEwLo3KOq/VytiCaqOKxjmmZ
p4hIkcVnqkWERjl2Oei5D/Cwsh3MHtcXckvxcpHA448rDPeD+j28tRGy134Z9ezIcW2LYqsrw7A1
x9zxiSXCPgs5qcf+9BRm2vXSdni+MUiqzRWlaTtIk98bNlo7bBmgVfueNQoLkHjEd8+ZH7FAbf+6
Gnu8URxRiyQqvos/Vu+BlWIxXzmjN6YGCssunRfrtPIC3o8bO2MWZIfrfWLVRRWy3w7tCvcG6+3V
MvSFabxD4av31+7KgD8sbr0JkgjFRHRQVIkeVFrOEh55vzgbVeOnGzFLfIxbEGf8ujZ5ihpNV5Kj
aXBJUs04W/KtJqdENqvcFuucVO4IG8WlAomkGHlmk7QXnfXzClEX69MkC7XjThy6UH9bANT+ZbTK
W/llVy/YwLTaYeXbq0O18cynUUtY7mADIc9g86xz9FOuBTFVaUcYpM1kFxAojy7YD0aC3WTGxerJ
qTpyQa1L/eVANpKazhdXZ9z6UUojySu/iYfTUV6sk3XJbX/pUFCbYR8uFTmwgpnUk2w8bJSU/I+W
DPO9c/pmt6ejSPSnghgtjo05A9c/W+VQ73aeZge02DFSykxPUsnn4TL9DquagN6SRLooh6cJ9j54
FsalLIxHRdEfL2IX1P2LUoY70X3Y2a6V9LLilMDZJL8/mkuE6bJ1X+bKaz3RIMGuUDBKoVyysvsC
vx+0VaP2b0xYM0J3ndXjrMmIsaQ0iaSODuQu4nQn7yUqc3nD23IkAWtVNijGhqt6sjlvOq9Kkc10
5RWsYncCk3oFlF8W/YrVzu9GBBbU65UyaaiwDk69sHs1LelW8iBQKh7UHERJlcOYM7XkZkpInKot
/VYv480pWRihD7Cv169HwxJOqeGH33fK0A8khFTM3sEUiktpPa9JoJ7EzF8icLQ3g/gTw/8QGM1Z
YC4ON9HAnZVQJR6CVJ9lmFMocKixxlA7McKAF4DAGdsFls8aNG/Vwg33VJzvo0o3txxO2L9YoSc3
ajrSz/lvHRRa5h9t/qW3T44jNHzoqGm7sjwpojfUFFE9FJXIQ/Np8tWYk0fqYnYB4Ec1BCns0/Ta
lxUuJR1HNSsXfSRYnDnOY59IMmSJdtCLvOrWekDP/MNlt3YO5W0wjgM3CFqIOaHPfulSXzrqRwMu
GCrrvy3UgoqbDemWxG+fkr0PlDSAkrd+Gpua2n47rnEsSzbgSkCCJ250uEO0vZHNXaXulk9u8Z0B
Lh3FkP9eWCaU2WZ/RQsh7YSCmcfeDuCokLDET+2c+YsZ+jIvVnvQ8525hn/Ncp4LEJJYSUhbAmyi
AdPDkHZpNdjYoTWMv9WMPuJjmAhyXciSi7nrrIrcLzrDZ9hdipF088agT8yoOevJIwl/n3sfOWZX
wnbDYF44blRFHaF3t1GJ+iBgLVaNkCoTNm/cz/vdJIL8A/uM2gzIFJMz+u8wy8EMTK4JZTgqEERM
5Ja6id8pdOCJ1Nmgnt+Iki3ul+IY15/oPnrRKYJ7XE0M1k74U6UARANP/Ijd1oF+7snZpQiTqnWb
nr4FJ59EOgE/RP1gWyjoQFgNUzPT5yBqelfrE9IAh4YLW/PMtuVdE/2FZjeeVhuGfT9sybypFPYf
CcfOgiuvpkF9dDBba/3mqj3sGh3PEL0Cg+XhVIXZFtHpCSRx+5QhtKLgluYA96maFw5/0lzmXxhd
3ofMWCgM5llz70glC/V2QVi9ScS+xnwjEAg6AETpdeYC0vX81BMHNNxq3vj135xIhzxXxbSpOWRE
JlNdm30yQM1qJWSlLuy8QsQqnJPFrAMX6R2aRJ7I+PI0oUkIuzlxuwdiP2ZCLxwjN3zJ4VYf9Gzm
5UG70sJt8FX1B5/K3yzJv4q2XDIf8ek5U9bsgipiZbRyuUWh7n5BDZSuo8yf1OoRXd2kePXb2dYW
74Sp9AoQq35F4Sa9ksKPHfXxhrz754CMw0cz5o1zpLS7/AjYTBi+gVDEq4Wj5xDGTxxATs7H8W2G
EMXJp5rSISqSG+fL+A6zqC0EJaNBN57V+yG8wY4d/v7FFhnE4a27hw5QmxNwsA9x1Ye/UVNKRavH
4ndYO+npq/s9Zsy8a6Xnz8fbPX34nIpys39cQxk+LVk2iqG9SVnnr2zsS9y9rn0BWauZ9LwplyF5
tWRLnCG+ykj49CfuEDu6IxxJ7+u8S3Q1wO5QzqkdX8ytA70WF85uUqXTZZwJXvun/XAfc8OcJnVo
EzFuBTZb7RLt0YkuHBH0pIZltPWY51h4jDbkl2Alh3a2Lcn4+3MD4+kmgtgCyHo6yX12bZHe2Myl
KzpJZYohTIVhcuzUuDXQ24WhC1J6R+22nrR9sMM+3rASTtM/B85oPylm1wQ0sOwoUfsabJE4q4Yv
tYREaHYglptmAUc1i2Z6Y5Uj9CQxWqoSSgw7hCt6zAbQk7fNUtxfaIiWzVwWkugW06+ZeACTv0+5
k4X5rhZO5G9khNcjZFgJKggO8f/JcDFmH1GuRM2WQKitZ+KC7FJqbixYpN7EZbdJ/A3/0b+Z6H3x
5bl2n8ifVrXmk++jtApcvc5O5zMXeNhhLXCfXJ2Zy6RYsUYcV+CNqUDV2VLLmG0+bhLYuNT+dUs1
BeDpJhMOb8Rbyeq6TSrinmpnJujv+q+QWH6wzA/q0XZWAEbPtwcUogv+/ad7/LN0RAVyiRshW/Uu
XfNhVoR+48kzU1uk4sLFyuOtpKv5L20FjFtEdCJAaNQEigy94/2jqH9PHe8JQPCP0kSPblsc5Akx
SdTyFkLYg7/2aH6QKl4cIP33Z836K+OO2MN0d6bZ4MsVes+T54jNgkNjqKI3tRgyLgOq8hSD8pcw
uxV95cal4f806qbPtLZWapvGpmUm7MPCZRMVO3k87OKHmd6s1zWF+6UteOJyVZLVbp1NHtmANrrR
1jZtbS6biv1/15UVCtAOi7dnZBCahY2SeoYxPBEfEeCYvIBuxxV2mey+8/c8iTIIVZbzeAZgrPsz
Y4zxakPWJFnA4JZW0UVlwxvNtu0IOejz//wuH0i6CfZTKbAi07czdf07Q8uIo2jDKENaqeRpG0ts
2HVk18V+H0a3VTN2Jj80+dR2QKz33pl8Pm/YstjVx+1Pl7TCodf+qoqLhm765tgUj5Te0zr/iuQU
0OKGEqaswEwKo5c1ihmEcgkiiyg/6/SV0PWuKpIrfyM5WtYcmFz1T4XRNd/dOzr+oJxu9HB/wFpE
269ELIrTfmX5+mNQ13+Mt/p1gmzlzFEM4woyzl14psfJ8tFNQzPB0kF34nxhZjsHzPXljdYFKqeL
ku0U51uVhaQ234ntiAKqPSJp9Ly82/TcTJ3V0FjFfp2nee6a059QBOhWUkKby08C/35oEYwryN+a
JDVmMtShA6tYNPSveQzb9RxYgJruX3do9eVlCHsGdGjZzhoFWUfEqssXg8ag0ir8LtU6yC5sUfyG
BeEzxYkHsWKnPuePYUzEC0kI0uCo3l5w5hrvG2J7aFhY5Wd01jKQrZNtclr8ze8RLYJF5sBK+lQa
RiNfqnu+CaPMAZkI5R4BhhM/W5tOabTmtX6c5F3J0YzV3K2ijYPyt6lP+keQzg+BNIlEMLj8+PEp
iV0qe1lME1jj3jjZmqMby69gEKIXBT0D7fWXPZgshD6uQ/E86CDX72CWj62ahlUkxbi2f4jEO6vJ
ZcRkcSU88Vis7sgadr7eVA39KFl9/kRRFiN9BEOFc6DP3vzoUTR24mJKZn0RaUghhtNhrPJ0a28g
pvLrpFPhu3t0g1cZiG5QndPEzLzueP/ACnw8EDA1jfFQskmYSjmTEJ8xfa6zri4j/arD/uz3C5bl
yKVgbGhcaUYIWRilIKGlmOj9HCCI8wP049LPvfgIHmdd00FdqkJ6lvdOMuLeNMhQ952pML0bZTrJ
6zzAlr+SE32RSJj9lnxjyk0pM/PlLyVUpEXIQEmFu2mpMiqEvLuQ92YNdhjl4r40qjE1loohrNhk
jGLH3KgnVbWSMKZqxvikxCSPEFI8n2g2m7kcDD8WRRKyuDLDU9FeWBp3v4kB/J0yrEvfeycILqKt
G1xvffUP45vNQAiciv97A69t4TUGcHHedKt69T4yvRTUeJafmN2iGJk21XLk2BGbtSvIcb1ySrEQ
xVgU2KCeF9shUxSOiJMoowwMfjaji147TY/Ztj+k4akSfSYHSn+57AKAT3/Ge6Aq609GLjtFjiun
UUsILJ1VCBEq6pSVOEjv9BKpZAPc6cgjWLMqwp5y/iu4L/jUZ0HUY8FCRyO/fxEPIExuXi2NuOjv
7vxeSIsci8QyRnAB+pd3+h1EwSkwqZbVI/cG9ZCiVv/ormdCNr6OPrHxC9VRo+8xlp2h4wKvpgZC
EfV7MAah2c+HldQ0TfMgW8Pya+NpffRMDfYUKelxE0f/Xo2hKU0+lSAlje7Q413oIzc++hYN7zx2
IzqNrxJ3zkNFPKRIqHMzVc42FchXwOym/sWif2hMErn1cMjSbzMXUZErdnlYAFcP32sLIM4Sai/9
NDzcFNSijOxOGOnWwK/V8nhWDnGkCnikjfV30Yqha1U4e2PM+kQjIjSrBvmcQ0rqTXNcDqeOKC4B
G6pzgL3zGa8DsMS3vG9g4YSp6eZFHt3Qad9Ojh5//LTZschoIxaKDuFsG439YC4106vYfG7u2tuC
zQoCBNmntcDwqX9Mmw+LHbSWznHfj15hRlOQPojeAE1mrOVzsN3LebY65/gP+Ajcsw72kgI8EoDv
WYBaQZ4/78lGISoOynDWGzig5s2AHQeXjWMUDXweSN1rRG9Z4rVQxfPksWtz3Sh4lJ3xx12vg3aE
Hf75LhHmaKZVf5kVUqxDs7e4H2jLkGK0IimsuI5CVQbsch7LlLh3VkHWDF7+cl3cncRq0Ovc2nWY
52ey4+79feMSQMTDcM5dVIYqW6DzLQfN1zMrufbevRkPYZALlroPDNz1XnpVOyPNRjTyiBEkxQea
klOUK6fB4G/e/7YhmkwuU0pPYzPOwbrpC6wxlTuJOjmD1abL4Bjyvf09uGbCbf9IYb8rzewYPykb
MkCsmAHghlsG89a+X5ROEpdtYmGFHaYzXfLnijIxFpxjGZbY3Xfk1+2kpaYkBL4Vsv0imWjEvtPW
g1T5cweCNCy3JLkIbyXu3D+fNApvDVoSAObsL0wkfbGYWevhZVzjrqDlrJLH5o19BXrAii3c+uO4
/SP0krESDjII/PjqToLe8rdcuWFHfhQL0ApnuOC77NEFH8OKK4M94X9KhS3CaFxy4UVcJxpJ2Lg9
dcsXVwpOk984uc7ieExb59pEnnnjbHXfZe7ke0fHcCdEqt8WbRndaYCYyRPqH6NMVBRZ23c/Us3N
aVZobQON1Qx11VviyR3+AMPlYMKgbv8au0D52c753pKMptP+pXl/p+t0/e8hD+hWf3UpZXY3enjK
1qEsMP0n/oy5lxK04Pdc73teCuOoXhVkBhzlrRBKj3KlmQ6L4QKbXbjf1B0en9U6ZYi3NbQAtAVN
Eg4In+qn5NcxepWL8wzgDuvt8b3s8mgeI0OXZxknR6+yUheWORe0APSX8nIWNcyuKY0hGuhIFwHf
IwKa9oDn9HZ0Ul5K7r0/n08kwUfZS1HIR7Z5rj1QsPYwUf7sIKoHgfY9WQfytFvOZgT2HUDYdj8o
bxDP1EssbVtWFD6yDMZ6EjW+I7b01Kroe66amkfR8IrGTESYLnOS7ta87/Aa94vL32LYoQvYIHRB
fs/7LNNgAwlcv7mODppW2z9lpP/8wQFwXfeJVDoudEsXegcns8RVPTBHNCFo74TkR43PNaw5RGGy
34weisjO/QIaBhxaPCj7qI6qHGpy9h0aLWIzy9LeM9KESx5aIf7TvJSFGUcF7yWbne+MERiA2iUL
/V1W1X0x717b37aC0+TuV/ggwrxHhsWM3zr9W0nW+Yqj3m/iGfQNYfTLvUzG2zBj9y/di9buVPDW
XE2x6j3D7QTrN+TwvVSx9wkAk29IWnmKpHKnKzxhBWC81Zwi6O+r16BjYgOFrsUo18aXeHevRqX7
3qymZly2M9eHEykRZ/05OqbmulnoG7akRYsfZmWyusyb3MXuSmfjg5KOAnLa+JsmYhvkNCr1fFbK
+G8N0CkAgS8pqb2XC8/K5kgd8RRS85gy3rqkTJBC6PATHgy6hSdKVtHEJqVWWYE1XEa/Bfl2bjth
Nx+tbf3m1WXaVqldFUvD91pFbIfWrQINe9HUTLNGB5nl9EgBm4D8Ae7n+aelq9viOAxz6dw2Wh3J
tlHOHue5K4SjHUwKoPy8m2lPQIqadNw33pD3wnM4fCslss/bFpJoS+W89isHZ7w6gMrBf6raYZIu
NUiBgnddgAc7NnrlHk5snFmHoH7eNqILxUvKTstxSo0T+EWu2fKa2uxon/rRVusvQPV6bU+GFZbe
BuOHAWezgBSzmv2BCunPRVSyKp7VsQkab4ytQadPY4be8OdyW8x+tAft0MYnbkbzmdHvgQahiXwC
SrRQY3WvVfXgOOI8+jaJLX/3QmWEhBcZtgRuCbWq+r8Drwj7eyTOKQpGD1q3F67anT6XGNSwx6SS
6hFFy6aHhFdbRJt5SWgbRncotbdrfx+BTdaXJ7HWT5Pc6o/Tvc4fidovzv0gSZDJSMy+mywyvQrX
+txAN/bqZkiRNEiIiQmUFaHVQZOMkWTzs9SDzCITHcG5NWaI31AS3ZHNZV8BBQXt+KVld4hCKoWi
Wsi7cmpW++/dLTVRyImcceV+D6065IRTuIDmLh0zvq/Cj/HfTuAbpol38D0nkvdyXwMiezdTPO7g
w+Dv+4vLEvMTaYZ3XM/kj928LHSSAbMS8sZykVYzHA3iW1KXsXV+WS5uC93gHiuHNigSi6biSKey
h7flqCX4doxVXO5dOc1DoSjqfogRUakbDEWqgwOPwzySmqt8K135jdBiBM0m7L6g2Gjs5McbaGnS
J2qJVFzLQMAPoTXGNqA416ax2UTitUNIcDbwQe8Mqz1XiTyN1GjR9kAcMUZtnJrjP0gDWsiJ105B
JGpGYUVAXRYUkO4b4lLyJZhhYqrRmpRxDZtyrhx1BiX4oiOq4b8jP0MKK+/Zxno9hhgcypAqKHpY
Krf9+0aIph9dd9D2j+7oCwsVYCq4E9pk6MwHruYFMjxgKxFR9KxtVrp1+ikXdsCxTx0L7eQIxdab
MeXrIIqHxgLdRJnXwOmIDLKQC5JSsDl80ucngrqjs23+nWfXl94AtDMCAwyG+mAuk6QZRMxXEbjF
+lnFjrZhvUndAbBT06pjrxB8+4IZ7iGZRkuf0c+JurkHr41CXLRN7MT2mJsKO10at3ZFH2vEnOpP
PMjsDdiDDe9FRv3i86iQ9NSwiz1Ob0jIgXBQ/82TH2maKTa9lleCJNeiAmV4xngRbOKtD6b2LzHI
0HJec4tS8Yey5DAnUYxcw31i2h3OgptRgMm1saQVXeJSqx6GHEO471+ZSZbwO3yYrRfmDDddDx3H
6dIPEsBoBHtF4Sn/i13x1NblivbInXDWOCfS4QtGm/b+PPSjtnucDzps+VmAnnM0cKbXGUjGcppM
LeNc5tJvmIgepKbDCIWuLJKxNwdwQhdxJoJBXED6cRygqydCJ+pklsy/kFh0hEsky4gakYGPF3pG
AzyIQ6gVhPTYNa/hskNofY6A6GubWR7qHfF19IR2UgUsZ4Hsj+hOi2pCLHCHs90q+yIyzhD4i3jA
/d7qSajGEUKSESyh80TciFiIZVIYnn7Xyg02HGLBk213giWlF7FzatnZwr984vHtX8RTwLcdSRTd
g29cWty6Hrk4If0Fyd8Zilou/Izug2MUDHz0AQ126DoP3v3TExucxs7lkzuro0VfzgBCWM2WZETz
XA97SsiyJnHbJ/dI4Zl9p5GlZkvgzd4K10N74mF8kM4+zIDdOIT8V4U7UTYtrjiz9n3/hAT8jKUd
T2jaF0Mmik20h5Cj4XGKZfReN53+eHAs3e2nLTA6pkt+JF581yVxmlQvk5PkP4A+uQVVFSC9xG7V
Q5qUfgkPMqq9ghCpiWlD4zF/sYSANFGJP52m4msezsZPMzWGZOUUhBPWQUAxWhJ1kOzuoRgZXeEj
fYPYOBaYOXm6kciqr3RDXBbsQz3JRWVnofabbYsYrY+Q1sn8m4D0oGwEQtk3RKMnk8fzIriwU3XY
FlhL4E4gx8/5IeOb+7Wt+IxTixrvewNW2keazYYWrnc+qwOcPcTP1h/CjalJKKLLDlgM9bd6hW87
TlwYzFmGeUG98VTImLjzkxchDqFJwB6KLYzF33PL9AzgiKLwNgnJe+rAhW7B0e5pdAf5dnTKD3F3
G4dIL0L+sUBYH/TrBj3YA42TM1gNOTfAr/n8xFgWIsss0WDXyuIu2hdbSE1pdcqdvZbb3BdKKgOg
9vHCq7PCqUBi1YcDHb6mWI79JNTMgF/f4YyS5QdJ4Gy8Xblvr1/0inQns5OsmEwEPhElH0WejCtm
kPRTwX4NqIT6nQ2vEak8fUGqmom60+4O8BQE0iTwwVc9/6D+lrpnQLQ2sTOK+5CSR3zct876JAm1
MNrbnXsvLPwKmXY6VIhhGKWSOyMFaJKzJfev4BouX5tGwkuEjTyY8qQSUU9wYmmuwvFvWICaTek7
75scGWk0NNXH2b7tbU/jgP188pQvbuVIi2wThhXV+UBcDeN/76Xo9KfBuEArUIwMsbyQSNNkUnK/
jgzS+8pRV03JOCUnFu0mj9b5Y8apDoVSKB7oLiAoWKx7yOX2BeVJgZHUzmEF5VlMjoR98mdq1S4u
bSbjcpHQHxHHjwDmyXzLk+Y8LsDq8QrwrcBDKeHiYXx6nJTiwC4wIolymUorYVtevFP3Ru7p1UGS
x5o+LdNuKQr0E4oADWBp5OGGE2y10jbZwpNkzz1QQxlcy74E1XzDvVadggWRXQioijE4Yg2JolrK
9wAY+X1KKnRAIlVMcVI4xE4eVQwyx3gfbAzqsBmU5P0+slan4r602j+zxTH72fB7U2HBAhvAA6oM
h3IN/nBVHT35VgyaYsQyP1rwBZurVgOM4KO4A+cYc/beUDcPM/VjoF0On4rfIBGnJNQKgonSboC0
sKxK3rHBVdp7sdHgNr87Gncgo/LUS/k9v8Lwg1dfomjotGfakCI8GbUaydkTB41pFd8FdxGl/yfL
6BFH7oce9wU0qpMgGOqCGbxn/QDPphQDGFEqrQFT8N9S4r3iV3psgg/qKHPaluIPD8623nMuMx8X
aopHTIhnSmFtlvkym3eMiNkF7phkPTG0QKCoXhLVtHWQQ+odUVKSNzVtaiJPGOFBpCeKfk9RYPYD
Ck24pVrPzVcQuf7GTGulnWlLtDljz8jZSToYvqn0T5aXbziXb4Pz1x57fVBVWMUUM+LcIGmZ58Uf
3nYIEB5OH88S8UAQNHw0qXdMVK86uy/jlU24Fcm9RDsg3aAEruApzZffju4r8yN/fNG0a4uZZPn/
Qwxg7ICuYLVkbQFSQHpgt2A6gOz4mSSjP/SthZc5HHf+uXYXzV4eqIjXKuKr6//LlVZb3M8jcFZW
kahZvkbU2JoH124kKLcj/cUM9S3Kukn19X49W3jqXzUIFz3H30LFcQY76/0bxktOkpOjq2aeUULf
+1TpDR8RpyikhKEwb/MEJVsFpOypNenDNU+6Xx9+c2e4dmBLXRls0IjiM5tomlqW4z4ij0TeENNm
H/UvvIvYwwDP6IJC328VM4hxs6XDMG+wCUcE7IrbO6GekBKx2l1B1gomuea8HN8CgHawy9LDcdU/
8m01rOxUDE9agtWwmN0Ze4GgV8KPsD7CGwIdUAx0kry9ngBleyrpWVZA63fO5AVCsNh95Fuks+bq
MynPiK5Z4X1UACoMPO55fBDVXt8wPuK0RC40kaW1OLHQthNy1GN9TM7Yey09YLvWBtx7dpurnnzH
wAFllTBCigDs33YIFXFhVuAjA/zlfSdzheDow+zgfuFjeViL/g6fTUwKW9tHZrafXwpdTO4w2Yov
IOip5CRoCxZyF9dMI2q/ONdyX5rd5bvh/g+dz5UZ9MbU1Wh65gKbTTRN40jW1AQ258cdN/mXx+sh
K2KFSQOGPgIMjGhPeXFpywiWLMVKo8/yltlKjpX+ptAMzje2zvJnRO0GgS8ELrj2TpYjZ1ytokGR
mDeEkWjcS1RbTQReunDBckuLIVxn+Rre2/IFYXq88e4V8Ieb9u3yReA5ADNwmKkABSDlVxQsaE8S
9bWrvKz6ELHDQcr15JzcQWdSvzhRAf9RFsEl6QcUDwjh4T/sdJaRgb5Tqxsw2x5GcBYJ3yUzmhKm
Wdcv5LVkxy9DvIFirmcGTfKp32uLZKPzGWjIdCVcF6c1uN49OOnulcF1Mj/rTLSfEyIU7vdW+spw
+GRlw8bq63wXyofVJDN4/9Kz7kTMVqYxktNQighWCSPoHgj4QcX1ts5Xsk6KHcjywinw+02CFwBE
dOXZLuEFi2ylOtCxbt34GTCgmtF0KEiVQCkog+YFrAlNzs86T8hV88Iitj1MK5R6NCde74IKtbDf
KOrtcxkCfZBLCU9CluQtUZdZHQVdWZxnZla0XhDzrCEYrtVBCvz8d7evQX1+eMXXOeFE3WFF4e5l
9HjhI5S/UFuvoafiCax4MuqBTfJlU1BF7wD4v9daxxwPU8PEJSDxFIzHAWxuq9oRYb55LeZVYQ/z
GvSSFOSZcah9B6LxtvoSqPaNR4eEVreveFa7kdFCaprVR91plKYNBWjPL6AoLPSUBuZJa2g052jC
3pHtMET3qR9paUuE5qPA/qZZUzwoez9z0jpc+Oan4zlEU96K5nRLW22USHUN/obhYNG0yGf8R2Ek
kTkkbzc3QhwWL6OzKc81tMruq2KZeN705hFXFZuIm8wMFrBTtBaL52pAAHg7n9oP+hZKkLF1ioWk
ZT5Wb7DB50syqZMJOoObg4sR7cKRxYcd5RvNxk9DTNHgLV/hAAmbCCIMBXRodujc83CJC9vD4qbJ
fup/hBj8nF+lJG7EVUnRkbwsST6RrkWtj3107NQRJcTaXbfYN7XAwjpVjWl9s0E86aXCSq829WEp
OF4Snn6BCFdMDpuk/yOJieVlXlIAvtv8l+pyeFoBRa2lTh2/f08hmt+/fj7SXb2s1WMiCYEvig6e
8swNhNgy4/1IKaCJmSvQ0dNNA2YL8yGXnWj+tC7pvV9qDo0yucJPmVAI9mc2oUTmxlTSZPUjySi0
/SE2TIuv6tkjj7V3i0NeA/vWjKchFUW140x9EWhHy6FNZ8P9HAgTmiBYF4rTcbZry1jGfdF2mgh5
OpDCnOHtIC6hlrGTkxndu5gc/2Aclup8zzx7k8jypp23XK//d/W3evM8Vw78A1us9IjNYI34R4kA
6R0CEGys9hqRBFPIevMGL1r+0oK6644y5k/RT9NTaeOXQPVQLkbFTY8qxzYYtTSgPwcCbXn+eXF2
ttMataBkmpmLaIdkebP67HplbQMF9F8pb2UEcqMGYwHu29NsOmQq8ZwmEIiWBWGgYiZnQWfIGVqS
dFVOJjKrwMB6qPG815Q+wFbgWghb+6jLeWknk7amapbfAT/rdbXJrB9MkDtZ+Qpjf4LieJTvk+XW
B6Fv5DJzdh1Y/h1frKNvUBRVFxPNkpAvBgyBSM6ciIMPY3ny8Q0PkuXqK+dbkYzKfvGaJo9EEHAW
Tpwg2DSX7cxrMSQb2RZc8kBQOOBCJ7JlLf/7QYZ10M3nf9ijM9ASriKoSsFalh3mo8gYAhYO/4Nw
4W29XG98bXG6wuEKJVzhl1PlFcly6V4vTFUEihhc3cwfqxHLb+txReaoM3qeJ+5R8okk+Tpdu3My
w5Oev5oItbE5GOu19L0abcX8oZfmJ4n1xR2QeBoAnjbg++6o4nJhyFedVEFKjpGB9InTidGbSVRe
5LTAxx5L0q0rd/Ke6/dAqrHGfryYteTycphKfFEcJto/9Ron35zVg0mIf/0k9LT09wQOV4lO3K/G
BzEvQFeu1jjI2LT96PnZ9Nupf/Ek4aDc0WXQaeKh7xyI/GuG3dfFv9JqT5bZBgTWboo07zGcMAmD
9PLDjS0kjPWPAfnywoRy63nMoyVY28X7RMrMK5VCNJJAg/Jr+/IpQo9N5FVE3pG9Hq+TSdNPzYuu
5EpzROI9Lz3CUggdUAJojYkp5dpBScWC53wtre+/ivjxGWdVvZcJh+0HTEHiXhHhLp4n+WcAXdix
5yDpvqpRQxNIY7f939gfARdWGLzn7pyHk4It4PG1VnN28sd858cgGmd46uZr9pcIT0T/PzRw8vyV
cTiVX6OLuojMPyfQ6otXgjKsQQvDseuFB/kW3A3Bhmns36PPNpkOsBkAom8P/m3DaZoRFJIoMeBB
yFU0tXD4hh+6IPs7i49uC/W93ADQZmr7oCakVrxZWvEe0E2Jp0fgKaRy2LXGRf+qrgSMcdTvH8Jm
AO3MOG34yvEzSrPYT53zAZZoDiNb11MDUUe5sE3cCQbMqWG3MafA72ti5vTTkSss9BALjzmLGDcw
oakky1i3TC03nAtcpES6VALJQoM4raB5WF/4tACX3jiPLUTdHgylIbV1O9zvmkaKJowh2f6mFL61
9ZEC0wuMpGXgwfqQXLws16dVY5/c8k8ffdn3rrFWUF/aMOm6KciWfnfqQ1VBaeS6hAc7M+TlY7fL
SNCPmZZz664dwUhFiRrPLRlcuIiwPGFoPc3wdrvBwQQJ95yoVDNQvhF11Ay5IN7LdJuknDp7cxin
IZud3xeY3r+xqaSEk/eQ5KX6WiHiDlH7VFxRfcvnm1QHN17wLNJz4gYU83TCT7L9IPNaw6TKC2C8
OcZYPGJhcFtBLdUH2QA6jV29A+wXqHJv6IPEoI+8qqIRHUETINA9wA5sxhosg3Y/bRt2EqT4xESf
UJeTOSEOtlbfgYO+FuSteCZs67foyuSdwi+ZZgLUELe8VxeGw398CB9/p22068tuAP6U5o3iyPcp
t9SS2BkksuTbdozZ8XrIf3gN/dIy/pdiRIe7zoDoSyA3KSWYVGP+3u+NgCVzhbdRb4KRWySPck1W
RYiq+4ChwjMVpu5JXugPge095b9zPCXnIxbOX8x0kaWj9WnP4MDiEUe5r42XfOuX/PLjk5VwZlzs
cxzpKwROC9udXCQdfk/NTkGGm/cc6x4Ul+ciimHj2uuLSTByWCZyAvN9t8V/4jLpWQ+MSAJ44/P0
OjmC/i0QBuE3bbzyu13sgw/CqZV5GbOYMDzMp0OwdUSoGFh87KzUGB3ROYbF8Xd8ivJ7XJNug1lY
G57lNMDPGzg6qVl3T76wGOatuygKNKhgNaddLMo6BT0yQc+rwo+iLY5YyKMu7AzfbM87Qq69uT1v
qOAcgC4QUykWQVeJKUhbX5I/sD0a7N7GLYDwcWY8vaegpEOFi2FG7VAPBI2Gxi0hiC7jClY5g+XV
+n47ttDWIYSsslNnZRie9DVogUPKcbAJ/+5ME9Qr2BkBiTpoChSumSouyFUs5Rkdwmn1AJlOVy42
9Mx1XEViccsSZtKFIQezx9imSGnLwOFpicqp4ZWhK8bUNgmdZ7FQUpXymA5msPaTtkGwtT+WxpAO
Yryplmoi6uEz5YhU4fGGitIaNDoQ9qT/5ITfniPPs3pNvhU7sNQTvkvvTVNfV/SlfOmRXBMK7+lu
Hs+wQ5F7g3yRLPBDi3gAC/Aq1F0DrW5j8y3h58YlMHb/ej6ogswE87JU32x4hCzcu9AyWZ3KIptD
9zn3YIcS+xyuzJv94jd/tZebl/fgiE0wtcjknSBNm61UDbYJJy9w7VuTcy897zK/rvhXlL2j/tEk
QOJGpv4KFQwnbU93HHHDSv2kBmrzA8rb+BXzS80rLbiWOpkaiUgharDMsjeprWkerpcq9ozSR/6d
y7+9BRV5gRo7QxmEaX5dfiYo8Gx1nGE87HYkOpnSk5UJw8wU8qwkZaGRvdLqT9dk3W/HTqDc3uVM
y3xUNANzc0Lzu6qllHgQw/pFEq4HuW9K4/DiebTe98Ld/h4+g4PmOMRfJzuHxNw5pWIgHtuF0UxO
SRXSMm4qEDMGivwKqbPu9FFn0Qc2ICp2VOOU7m4NRHwpifdZ6vi7e5wSM+65xoPCnzVP1e8c62X4
bT4EsZc7xwFLV7hXYSux4Q+qymGF5g0zIbjE3alHTg+xyGEAr1KDtCRV5k8exmBwivmcwofbyaWK
wt9kLFEF9QxKF6yY7CqoDmmmMvv+CXc2wbQHzEySae7kkkgurcV2YUmkLzUPNgQETvU6dlfIotmh
2/PeoPF1fp8pu5tCxdcmm0Wfe7L0kjlsBHqLkC2Gl32S/Z+z0hqqZoaJ5sDnoUA9WUUIL0igt17j
Z8pslI6DOapIcybQsFQYRJi92iatrf6yhnL5s2pBbQIZSXiw1e6b8FQUAtWIa+yApZXyySyehBCv
onGBogfO/YmQnMppOQRjbD6CP5RIwL3xGL891lXQItEmCtGIKx3nVKF9VHR2WFafIDl785LD1UQ7
huXJZBO8uVe42K9u96N4PE9N2So6cT2NPjfx2aX/k6r7Es1YLdr3YrK9dWoAzFPt5BeCbzMeLZGx
6pY3yzLHzzXybzGxiozoumplwJTHAikwX/xP923CvHX3gLdQMDuBfFV5tSrMNs6J/CyPYgsCmqEO
+z/FFNsgIojsk6ax/V65EpBhiSi3qQ+xK/CyAObUTsjaIS9VnfOvuNI9kp35ktvLKEeSOnnWD0Jm
W7R5zqb8LJ+ZXAt1zQDnQrKwZ1tiyiDUtsXr+xGl9fQwbaNaEBpO6rawTqMr/s+vL7LVzH+2PTGL
931KJC/CcYbDr7ZL4rlSTMCHWQpga1hwBSs+1EndmSa5gQGeQQttOb3+CfHAJd+45wkVIBI356bc
JmKkZNlws9vlgztFBQnP8p1D/A09/JW+LJpqFHb2AFeQXMNQ9JBTK1zBly70+meJZlstlAn8SFJp
WSBz8i7Kmi+ImxxShtX5XgubGd/kqLgMwK4C/XQtqhUM1E4ehlBYrwViq9KUzvqnfl8iSLV5yT9p
I4cqmp75qYNKZABFtT0eq3ej5HNiPBeLVY49byn8EvoWJRCwNIFQtTDq2WkyeWZGBbaLBUVuGsAf
0yCP9N5dq6v3DCV4AvaayLN3i/4Eme7BKpIuowZ/Tr48O/49uCoYtgX5uUDNVeP14fb8CcFHUIDs
Od30SthqUvBLLfhp03jfaQAHzx2fRAY3/8B2bilRgr4SByqQXB2OVrsulVjy1QPoW3NQd4c5EVzv
MLO6P5VKx6yDXre9rNnlQ4Bpdt4XqjF6r4ecipVB+gcQMt8h8uDD4kUrIAbPnxKXcNELFbdP32G2
SbNvqUv5xuuqE/bySw9qcTSS2ix6TyZi8cOb4Nlz5lsG0sIGd3ujhHhQh+AmkJ8kugaBqdvnufPd
w4UMwAxmJGllD44S+iEF4FZIQ3EYSPuPJpeEr8ByMm/oMk16ltRxZrHDYrABWRzrfvpARWSi9evz
GuyuldAzP9caokMRgPYj2DLuVuZYv5TNP3IxU1s6oBqzT6Akpbtn/G8m12T+WjPchijX8nPUpW12
vbQufJiuXnMcO+0vmz9w3MF5H1QQOT50ZYpaQz/oSZszn1Stmo12dgMEr0xHR93d6DwnV5VZ9p59
30VPXALzMIbGQPv45frb9zf4r4XG9iJTJw7/DDQh2wDgssHrPg2Y0JrMtt21mE2A8Ov5cuhHmuF+
bnEKQ8PZ60QpV0CGCZrijNG58ZFQJVbx2cD0DVgbsDmi5sG617byeeFgV4niOEGGH/84bxHkqfZV
XJFBDMMWPCA2NdRoikZtQYtIUqgixB9fWW+pOT5vR/ulpSZjqyplX0+rffTQyMMHo4OLDoP/UH4l
vvSHlidRErqYnd895q5a2PeWoMqn+dunWEg+iZOo3AwabrATf03ZReX/Zs3+xjqljrkTtmAZ9aQ1
FLgdcKUnEs/tBr5X92QE8qCPtKgzFMQPiG369gyUJrOV+u36PMaREPEBgQjA2DQw97KJdl/2/uiD
7GnV0tdlW0DWIMTtaz8f+onRWUyV3aFzwtzpbQ2AFvLA4737I/+oetxJSe6RmRlKy0YBB7Zb6Sxv
fqyFDrLLxso6PqvRJnGMBJ6JUuz/jp8PMTKKJs13zvJ+Rrta/je5sLAv7/x47ocELPXtl8xqsFtP
7hchjhamRhZYDmYiAxmKmyiy670k61ZiuFheB2OYHQVUUNbDs7NIUKC4bgBxpumPRcQc5hnhJEk7
HhWbckP3Dx8FnGYGGl/uzT2yGl4/VBD+vffa4tBE/SXlhefft6UT2kq9L50WcvDLtxhRToijW4+P
E6cd9dgVUn0qJnB2JeEw0vjOVmyO1HKw/ndOMocdWAEspw9I/C+BUytyz39AnQdXGxnSwR/UuXIf
xiwL++nVWmD08UTfnShy0gQij3AyLxhI8TbBFXg/x5D7eqpc9+UB+IDW2twcKFo+I7/Maayk+Jcx
6IC+D33N+k3whUHX87+RwPESVh3hJs6bV9iIGkrdQ0cYWUUcLW6q5ChGjFvKVcU7gXQg2IuVwzw0
vLrUb7J1E5PZCCK3mmChWWs0KCfxV5VSGFVlfwu6gz7PuBCId1ocwGcsL9pwPWSh7Tfh0BjXyhIC
XLg3ba9Ul13uHtdm/zd1utGKfqX68BbE3YppcaQ+D6cNrAyPIpMFZAIKnP39qZfkLzNRZI3yZDU7
51GJPVyJjsZiuCr7iXOfc/0oEtelr20jcQc+GxPT8Y9dwCR5MlmIeXVpiHiDZG/+UbixbKJuZ2DU
/SgN5yasUHSqZ6yRziaKVWc84UlrgV+oz22cNn4zEFiT1kNRz++8hGxB+Pq8QEZHvp3LZzDh/EQ/
HN8Wg+wpVgvmbzI5M7kEXkfwJ0lr6cK2HtqHKbj1zRkWVttaLf0wM2OPn3nytB+G6ozSZri8KmZ3
YR+YQOLnlPW+p2xh2mh6msJsuVTHjWBvZYLOXPIUUmaXVIYWzn0HZvbXp1V8nENmjPAmsW2xdARr
K8EvSHE+C5NZxBVO9VdxIDkgrVa4yc6IOn79DXS0pOKXY0nddWTMCwrzgv3TjM/E5glWSyxuhzRA
kuMy8Bs8J0GxZTY+SyKHI66OZImHCQxl9Mg7kjY3HwDyJgaNjB9AK7EQ57TpE68Ak9J9YZ0Xbbbb
K1P5/GcavQUNnWxvSgZHD1kIsVg149lFFtJ6qi1drUoluEjrLrmzF8VrCFaKyclE3AmHyvzLNZwH
O8BVc0ZyUlGi3e1tiPOj99cm47PmJC6fhNwEMTxKd0Ufonsq3lCHh+ZC3X/csghtVB5YW1TzUGj6
Geui9pF3JJzx1V6N0v0swgos93kOlwhTobifF8yIuy6UqRuX/E27QD07mO2xsvgtIN7waJ2aFfxo
wl3pfOU8Te18RtlIUAP2R09cdKGxdTkvqIvJV7PhU0c2/1/El+O0kaBrCm94bxZWdYSS4LYtU3k3
Zk2NIy9JqtJ1K/4P7twDvpxCl0xYL7Yn++xya98aKqqrSmy/PGMUR5gfA8oioJgIw0p6zywOSoxD
GO59QTU4ZCI7U5nfoTWLWCW+5riYHwSEF2OWpFXnSsAfzfcgU0MHNngRGOr5QBpOA6gA87Gt5mwl
/lqZA+MzuvtGEGcnsfhm7RyCe3Zp2VD+7sjfR4VM9+NewRPTLL0GXco+xlzk8nFLSLQlDWwcfB3I
DBwVyijtCy2jaP6ad17MVQ74DTw+duBB4+JOSQnegwYihZV/WQxJt52ep++VYlFsVUZKeNUsCbFi
G/UALXHJ0nLluH8oi2EwGz9DWA7rGBf9i60dQVexjnvLhrQ+zZm012SATXfqgzaX0dKLQAYlt8La
x5ID9XAsqvdOF7Qv2GQxJwyVEIqHpqkrucKFyy8iTWnxMLxB7stGXU8t002U4TNI+5Wk5GAPd4Vw
FgO+aBGXsPLZTgyDiTo4IP5DslQjs07X6Xy82x+qTeH/TNO0PGgb1Y94LI8xJ3K4bCsTxnT5dQCJ
oG0zeyfWR9lZPXE/HIyEM81GedM9DXY6wzSS+yFQ/gZ+ZtpNd60zqHHvO1wjhxhW0reAhvfUAF8P
QFX7O1GQMYmhG/2cxgraxMdx6wYLRU+TzsRxWzUyoDlhrCtka5Kq8UzjwPg64XCnnB+88E1//j1Q
LhvdQVAoMpFhT+sTY47y3QI5wJQHg4bSQW0Wd2eDp5qS4YPC3DsPTOJHEsghh5KPQ8eKxViPfLLs
CJ6fJBid5UbYnCwWIuGgt+JnkVC78E2yRJh7oW5+h081B3VlBOHnh4tTJ3Rm66UTPqYmqJkEOSoU
DaIT4VT33SPiy6Lqw4IAKO9ehBGEMPnKA/8y/s3XCOsYDDp3s729S7qddeeTD0nMiGGF5hBuXK9p
NJaD/dUaffOnFwbCMEwQvBuUE0HpXFGR7KkQW4q+wOZ7jpqoTO7BDwCM3zGu3p8Hd+7hhuSM4oCq
BBDXWMlHZaGZwARpats3IYlrjSyhu/WXjsBbyzmqSNduRKrBRq28VyOviNgFf6TW1ygYhJWY7N5L
ijGNqFnstcppyWODnfcS1UR/Gr/E1mOXcaE/InolTigXtyuPMJHSN2HkBheLo1AbxZ+YN/WYU1bF
zdv023XE4Yzr+SSUtaEDnVxD09Roi/CXTBBAafgwsaIgC8H95KudIGF0DEYz5gwS5BYTdRyrZq1/
xFwv6fDnt94c78uc1gvvOtMA6Kx9e5X2cvMRcN2GV1hEKuqaQB7vapsXolfuurlRrvG7UgI8pGuY
PxbO2AKvt5sNaFufAetQSaLvRwK3MfcJTimi/1jO3jcodcdCUZsPfWmhUgu1+j0hrwtKiNCuUjLY
lhnZTeT1Gt7Z2sv30tU80AG/S62vOf5RDwc/WjQ33qF9/LwUaq0wMWsaxYaUM/ui/AmdMVi0NZLW
XCcu1HGLPcSlwE2FyJLws8l+2Q7+oSXlq/E9mNcG9zL/FDtACtwqOdELqVPB4ZgQjhYU6aD+UEnD
4vZiaKvFat56xVYB81HKMCMrmQL2PhOb/uXaEkP8RPyaJ4KDALhhH3Ts07lri+ZaSNKb3vXKXBOj
RTxCG65j9OYG3mli1RmS/U7sxIvy1iNkxBeM9UwibcEB8Umfr1ym0NVjzVNFVsBOJJ+o3nGkZXbi
rFh8nS0GG26/fA6yiK/UHxL6BlMpjYjII1GHw5mc2c/0JX1BI2mUg6+pCiVuLcz9QJnyfOncwlYX
j5Xm6lmd6Yt7eS0Jf4n2nPCW/LPXsRu0rzUvMj2czAyjCtTKNgkQmkmydVlFO5P2EtITISynViiI
NbtAdccts1Voc9fHLds6wkWc9M7nvtlv04zmome/1S2bppjYAzzCSD34AI3yWO6547Y6Qf+UnW+u
yaNe8/ffLmFuhFvDI8BYLx07zwFSZo7C5cYhlMS81keo6IwpQnBN9ybKZQ17o7YeFo2BWsiu2+CA
+XkjuIiDTmC4latUCLEAUTZriQvnqgnQgxAppJG/sd6Pyo606xcgjsycCUfefIonPzdKYUboHk/u
pS99YzfiDlTLjk66VkzMH1iU+A6jfXHe0mvxeK6Z1yZ1Nw88kNQp7CcSqXoXYVU15KC7aGvU/6r/
apVpfRQJDKoIujQkh+N8VBBiBp+EPsORjtUHvOmAfHOd2Hvqye0jUbCJTh3g2WslKHgzIPzgGdJ7
KcMYbdCB2+s2ddXPTq8+JLwryjN6NJ4btDlC0nCzBCRZ38xMIyDi+dNLGZWgJ7IGH4OrJDNRbCy4
yh+jTSTveUez2cQxt/usWDt9njsk0jPGNdYHvYMmDXkQ8DERKEPSKxZv3goWKWUfdy4VaTf2eDdC
DpTbnioGHypx2ppXipZVFTx59MFZBgrk0GPperl25SQY47aHlaMWvurGMnOcMifrKvfTwNbnWhcI
EA8GwLpxz3DnuK/RBVBXzHagJHIM9xXyVmVuLemZ1PKvutItnDgkLSD2/83tgxgk94xvrm0PT4/h
wLXplvpOgh8wuRhBtxIePaDRM3ktVG01zHTw4SmDMsHr1uq/TIvpamt8h/ERj/gUm9PPGOTaqnBT
uufsTiVpcKfPOksxzE1M6Brsp9qCyjHvN7eMsWwhbPFCCD5FuCqBE70w7iOGiFmiKmOVc+vlHB/e
t+CGZ4JV2Z6nJTzhb0ez0J0SMMd7SXa0SjieUmOULo8+GFdjATiAuyRAlUb3BkjibY8VkWiTPXjc
44xn3/lb1czFQUfUEJu1U1AtimU31BdCSc3Xp/7Pb0aaJ2YHxkYT6x1MqjpnZH3Fqmgf01TXiAaM
K0KOxsfG+ojl+Vuwecafyw9LQzyXeld6jNM4YluQrvxkFL5ny0XjJB7Z21kCxV1gOhMJ04pjckcA
yzm0EehYh7KIwdalesj4/DBaT6dQDaS5nw5CXlOioWkSL80mi8GWlOjPEO0zA3ltSxoI79VJx7Rg
VnpP+KnQWpE0vYQmqAXz+OiOnn0rDbOSxF958dhv2LAbbnGHRYJLYo3hIssmpHKVBKQQrN6HqIIb
wU6p4I+clXBh38/99+MQQdED77IreMFeHvFlJcX0igTOs1465ZFJvFrzCABMC+iBGVcKNCH77iL+
zH9/jLf07E/Lgd1FUPr12ZztmfwwW+MHySyiW4b3qO5qy8GEdqY3VJJMMHGcBL4V9wlUodZnOt5r
pYT79U1DeI2ZpRHXOdpPOr81wmo7TQbwOkpjIFVzyZFaY6jJ+8dSe9cOg1D+9bbVX+ZGtM+0BqjG
3126z+3TYNwIMJGPIYw4S8SD66/AUHA+AkDWkd94dfPk8YF8M81fLdyHNNZoBvJC1nFCEUsdY+FE
x5sGYCclrRMRUL8xILPpRI4x9RmGPMAdZEqcPqzISvwDGX3Kk7uFWDLcYwaarVlPKt/+4XuZvYt5
Ge/8HjvwrgptWwI1+0guNQGmacPC/iXBV6cRkjUHX5SKsRO2aQzNczVyV8F9x/iUYzdtD9gq6rvb
GK/ptvvruIzklm/Cd2B0F4hdHAGMga+C+cBmUHZeVYu4CME2hEOqooDHb6hbGcdilhUEg69fUxRS
FthoH1JEoSXGSrfsIh+HSXmujAJSJ2yndft1sDXBgaQ0OxZGWyGyK2sONt2eOJ/gmu9Ozb/16Uwh
R4Geh7y5n+/FcEF3tQOio2zgU/gX+3vgOM4xB1VTuTTCgiQf+JwGOJpZFTMq3lzZTvytUdU8kZTM
i83TKo4NafUX2Aak6rXS4FvMnex/546BYQCcmj7O/lQPGtiv4dXHnbHMi3rhBRMrIJLwqxNsdiMQ
QkVmoX19R0rnDci1YC7vez36SfTOGHriHHmPVt9Dm8bj5Xw+j3pMBTu7RJp0vbtXktrcNPcWDvAO
onq5fJd4z32Tz+ds2Wu1lYDlGdXSrgVkXXFUiprDD8bKSiIekVFeoUy/hPlxqmzFH8uy0Ea15KLb
lYx6eAbgmWydEKPulge8AfmzHx+rKl6HzC9Tp/4qAeWVZp309EW9GRPs303OJKQFx0oHejtt7NBs
RHeKjoKLC8emleKanEFst5Ib59q5ZtL2HfTweSwmkZmzo75NbY/2XAfzMzZzsJTpfyTEgZZfXZiA
QoUjSI1TMYCpVf3ueilkWq57NOYeCzkvSWhoznPLAWSSGYNN6b1Kwq19FBXBJbh1TG3Ddz/ktkKj
qlduDJTZUIQcDyxz/M7fGvOVimBDikMxWyjmv3YGFxh71Llo9/wODLMq+1w1oeY+sZRtiHBdrehp
nYng9rIKN3IFtVXRzeLY8Oh3yUaiwhcCUAdIUJKIb+N6xb2Kjw0T9TcpRH+6HOSEN0NgKs77qexS
7gogzqdh8IlAJK8u6rHbUDRK/NmhRg50a8vuaHCP948Nrq0VVRdQ+Me4egegjCagjuANhgbsvf3m
zFx3NM2eG0V4tKENYsIlob/yXWE4h7inlEiKa0HIcn0qPf09CtlLl9MUeFwTxyx07tjAxysaaBrH
ddT7+BeQKeM8ywf+8l+W3Mm/qy1dQ2rGVgtkgh+k6pdVvi43WddZlm5FCPpTKwrjcAdOUATnsZ2q
rFM1uVdJ0DMnm1okvfi0CLP5k7MYPckYnrhe81G9qpUISK5Bnk4QZKMdJAFRFS2ZEjFoJBk6Vfa/
sFqG846oEWjbPhOLP6LoWO6UZwMulsPr6FeH1XbAMYSkK0HRpxC7cdouVeiwM0BWLKYStRPHgXJ6
Y9/M0ov1b8W3zpIZHJ18TREJ2vKpMY0zZ0YGs5pxvdHeRbV4khQQFCO+esBh7UdzajeYWJfW0zYP
7HWCXDqUeDpl6c5rcWcfduEuSjMKc0cEPixt4IQ+MoTbmuN9Tqt/sEMzKzmOB8tZThzTikCkmkaO
hBNYhwWd2zqm6aMuwVLDl/2ymy4PPQlkrUIvi8Tml5gsp3VAW1V178fAX7Lv7FeBzE8Dfz4F7UWS
+pCTtIaq1I6ebtko5HW1p+bt8aMJ7Br9rwi5nX4XoMNREEJH2IrzDiwzOd3nL4i8eZuVyZilQ2iH
J9cDwvjmrScJHgLNQTdCFQaIg9vYiJghcQx/3WjyTOqDxahz3GAMhVazWT82H99QbFyn7Au0bswp
nI7SasqOtUIuYfI4VAonfpBhAKs26JL1Pvx6EChi75ME31QJ0fPHJRYp300FDs4aCEBNFOgB8dGK
foPwptrwpj/kkNZ1Bm/fNB//Bom3KmemrbAkNhTvrW4yB9RDldaeWe3GM09R5l6GrqymegVlTQ11
JizTsjc2zlCCbJaLPDX8ivOyvIQbQLyvnHRk9kL2W4k4IUGvqKhL3a2IBcwKIxKt1EM7kmx4M+QS
Zv494likn2F9pB0FCsFQcPu9hjvJdAr+UqYmIdLUaUQZ3ALbP87sPXBFHqVVzMEn0UDSmajBSEMa
qa+6Ahg936xpRQ7lQYM5PHMxA9kPlzz0FT96uI3RD9FI65lB7pZyVtn8bmQ0oK28X4vqtiCtSD43
Xx1EHFziNbcJCSdW2/5meyrZawahlPrRKoQd3712Dms6OziFtZuPlP1VOpAJ+P+aI3aDl2exB9rW
B7W93IYd0gJY1nbHmz/kHY0HxoMc2ByWPIIWmXb2nuiDwcBV0oBoU0xFnGdqKkz7kzBBroG9ckmo
d/5qxlXilqERuMaE+ZanpSo432CGcJycNuFLmBNPSpR0qkcDrNbBvefwkTUj+9m0l+nNSoz3tYKL
Bnd2BpfCLiOLQouiTnKvwLNecPubvQSmtqvRUCXPCtBKTB7PaNiJ45hIelOPLBTEjcUq+5Jprf0o
myzzpJavArNIiyM66MqXKRr4SJS69oD/CUi9fw/KEBdJImsdmwVi3Y3r25vL+C48ZoI0IOtQEg/6
hxBE+gPlZeptqeqiEjGY6r2TY4Q69w34tf/SwP1F0B/jdKoK4l4xx2whRUzM2FqDqB7kXwMTUFN5
KaYN2jJ7lnRAXdTtD9E6C3/B4zKJKEgATDlcpJwSW73UeR+mrpkVzjUq1zcGJIBSnFyeHZcZnqei
+lKKsAE1QTLyO9+sSAJFW1KKTcnXF16dIiEvHCNm31DfxgpPhD8Mdd8wzSJo8ZqxniPre+o7MVt7
ynOXCKdGW54jwE64seG7VWC8adntDwPDGY4jXASjsDeVyvg030/73J7khezT2L/7ehSZpmXZMwTp
b+A//9EWneSC82lvxMpddda+MjqC1eL6dg6noLVVdSy6KiPIMm8138DxYH0F/SrqDuF8t2JvQsz0
p4+zXH+9zJGfGHhv6ZNC8Sb7tVVCClYExy38aDnMdGrgUedfmJinziSuZW1z9Q4M4sNm3QuIl/el
ARPfcS3nL1WCfEXl1mIrxV/EpRQzRqPPy8WUgucD068zOY7rDFU2PkHxHv9uAOTYtx29HBALU5JB
uydDSoQC0NsoRWsLY/ohUTcOY6iScOynUDpzawIGBMu55O2gCbloyxyh/unkfrWOgBAUufwCbw4T
0nFY5Br6HPXgQW+kU1fpqg4x8uOD3LcFzoCAHz9RmGbgDYmT4aGSt55+xBTo3LmArcg2CJLdmEEC
XsFDV3uVVvFTfuOkgwhuoXWjY6z+MnW1+vtIWLhZSQX7goP0L5VoGu+n5DGGiicSUYTVDq4j13sk
ko2iYPBdf22UKtY/Yf9LeTNy1/0KYOztLe/k3J8wj37u8gC/+JhwGZZ+1S+RQHmhHlKj75NNA5+g
qqC/4RGv9QCmKHOYIrrsuV7Rj2WjL9/qdq1aO/4Otc49+y8mWoNdnVrxjfsBedZq7PDIi3svaSQg
aEWaunvpkVwN0JprJdKhDcdPIy52AyzC243lk2zQxHGwcpjcQPFoEn/pSDuaYnfkVKgkA72lnBkl
C8zlD+QhnygybrqJ6aR2YfvJkC57M0+zJWX0BlSuq9FgQWphTIGBl+hPq0JX/j7hgTOcujI4nh+t
NJHPkYLqyYqYbVROOiRlXo4TuK+9AKxZV2Gn06ONHRsZUEtcbQCNEAmRBk6JDzn23RDzQkNb2Cuo
lEE7gvYFbElwH7FeprSKs2Ie50JGC5plzHHhO9BVYtj6iZS7IBDwnTOw9mxun7/tA15fytv0pOS2
App0Z02rlTvyYMroa4WKBfUJcqz0fbjwk34M2nbpZGEqW7t3vzDdv1yBSxkRgEaBO9UyXN4/oBOD
KC00zzBvJTzBeZZt+WGHTNdU9afOiUluWuToEDqIDGL6qIcYkdciyA5Vv9A7cuzunkkeDsKYaFkk
L9h8AzUN+uJUX0rTrhA/lNX4SudK+l8UETN4OEOZcy7oecTBwMxSsfAHLtwgb4TY47g/wOzcNPzU
XOfA8sgNWU9+tTsjo2Dfe/AmXJBe4DtcnvpZrAJNgj++nX3D+L6khJuuUDlOhkhEsa4vtixTJ2lV
/xkH1vFuYXw6byRv9wfcJ02NboEyQsQv2bzJG4sIboXW3FJMyIWD9jr/y3fLF6OX6uWLJYrMlQep
zyGNTNBXrT2/9K0RDZUmhCszyMjsCz+BoH5e8/Kt8VR3Wtbb7buaZgz09antIw0hUxwJ+VBBMz86
9ypsKYWsK5n+o8y/OUvxlsKuE9vxSX2I4BG1IzjuMgW3Wvzgx4+vSleu1roxHkmIAkfmTpUF3Kng
lpZDHlJ7bina+/9FrXoFZUV9HJ/nPyZDiK9FDy999Mlv0iynMeY9lT7saqsCpewXt67wLd8rb3k9
sYSHkIA2Fn/AbLsb1D5hkpStZG6XCWabxtGQG/bvs1buaMGPiNcsMdIk8SFU1n8k2PIXB1z2rham
yppb4OnOt6dV1Ss1VO+FEckgYMJvbp4unJLHM1p5SMY312ya/1Bh+23O4xnHApu8Bmy7SCTlAccz
lT/Hmn8xgTTNTkyzUNJj91gQ0kctaijxyMg5Gua+JTdrxAbeKaaFr61t8eUUx4pDA3WpX8GEXZ9i
tqWE/llgaT0TcdCljB37Rz9yb1oJMAIuStUXApdQ/bvEJBaAPKp36e9YvT9Lb0DtDXVLulveAlEt
Opfa9pnZX+j5jjIagVW78EinGwHsU3dO6qJKCvlWOhCu1+HEu8NMiBUIzyicxmX2AXqxkBYxnGRz
sMkrzIi+aTwdbqGYsTHU7ihUkkU/HRXy3SqVPgKvEVQuS3b3GW+oLPUIx7RdOa/gu1ldYkVYqVXR
0gUTQsq1qJpWEj6e0RJ+oT/UjZGx2qSSxWBpt4LqUiIHlejbxYfXLAa1tysyRZdmyyhNMt4MYIb9
BkGJogyvyj+NMbwaBiaiVuQqqCDFms4wtQsimp4IB/hM0MMFlRzm7WTzDHrKrk5wNB02HvHI0f0T
2SRxfoVYMvcmSEUqTqM2E7gCYg8W2Pe25lCa/3rZ6dAesDgLQTHFOvqjINI0+vuXRGdsnkO5HLc5
sYtycpC9ppzELlXrxa4yh94Ro+b9/H79HaRKq8KKHZvtu9J6aGQtBsO8tMCJoTuVUT+SQr1kBzev
BKLC3uo/bADkQ9y048Xe/p63JqLp+yvBoXp3T7xWUHPTKRBaKREeKvh8LE8rPkUYH/A8yAiva/zJ
9I/Nnb0QXfA7TGRSx9xskZodrhWRzJhjVKOlb99hXMpp9bX7vTcFz1Mlh5ZLBNbn3DuL7DPvGEFr
8wb8t4XciqSZ2wBF+foCbRhSlX4/gkzz5hKJyau8+lkKSWe4KZmjI0fLQLM1dsLMHOiJ6jkIWfKM
KwrgbcrhC/w+s27igXCeXDlYZiNqFMaVwP/DsIzRT2S8YMG82gGikgNzJRhBaf/96E6V+UGV2f4e
pSUbM0PQVhhD+SjjTci7E5f2NPfX/dU2f4A09e9xytTi+YLIfnlsvb8Z4gP3GyCLJG0UA92JAS+A
+SsihzZLd46HvkTiyIAa6JjDhaDY6CJDX9YPVS08wmZ68b4mkEZUkCz7RKzlnHCL2UBI5/xdNt8p
6nkAF7ArY0ysUP6V6NH2sxmFVyg87nWjgif4sAs4yOFAxyLcqZuVhcEp19/ae/Udh7DF3QqlbCqx
IBzWc9ZJUixVc8imYF+PsUz5aZXZWY5GjMwefz9lemOSygp+9Zn9YvlpzEbSPTNjQQlsDYZO+cNT
lZA+E5s5WBC7TtdpgrAwlOjyi+SeQ5oUT8CseA0nBZFfElrGQ5nTemkvjSzxBYUIFonqTIpWazhb
TtNjjfck0R1wRY+lAItF4W4dtsKW+1ySHVNS76/Xfqx43YB7HArugIvvvVF4dcEzKo7j3uEZsFn+
R/QubRQnGrymmHYpOccxOVSTiCYTQWovMmcygZn1kXj939K9S2Rs/HLnSNn4bS5m57e+LDyp2QBN
Xur+PjYWidD74h+iSvVW6cWXoKvCYzbQUUD6Z9Swsi6z4xtPI1xXdCWeit8s/eqN0qpncjeXseZN
U86Bt0XV58vBdWfLqpFowNV3T0+470PZtUkYn4khxz4c/uW58YzvNz5I2t4vOoah2yaSdVHZ8YyV
JMWi14J2QiXHqpjFEHi0DpvTR6WAZqfgWu48rCfz+2lGYdPHv62MejIuF1/06F0OKY1UIYu4SR9s
5qvOQtiuqnPjn8twxXq96oke9yVmxmRvsxYPfJi8uZvhguJ2zN0P997WgVRh0nXkLXRrTU9QV0cG
DI54eyZmAk5cgEb/47+ayVC4jRgA6CvcyRDfuf2wQHLPehitfpMUOC5WRM6yHMq6DMlLD75p/YQl
bhNaDKOGzzjKyZQx+RhNTHvwKfYYhDgP+ZQbfPN4w697hFWogK+0XPLTbe52IppSJBEoYCxm3bq3
unK9a3S8CbwSVEqeMCOCkH5tR389ykz6Apl9PuvnY2TBPmXp4owWAATdJ/okrabO61vK5/3m310v
5BEu3tPBqiaGusVP1LMXBmUHhv8inBBQ8+z2qOyNhNMDbdK37TepQl4XSXb0+D8gGmTKauhB8luh
QToRELE1z56hOhSCjss5Y786sNHSuH8m/P9xufUPzK4WnzXPHjeHl1X5NKggDvVAOca971hEEjaa
R5ZNeneIMqQAwNsdlpl6MIfEISTl5gmDK2puqH4mVoYm63TCUPtyA74UAb+vus8cVgXp1pxKBvYV
3a+eLoQoMb3Zu/7a/n0I5LZy764W8xNL2SJFGIzk36O+uWZyOUgIT5PPjSSXZEyzgvy3lOAXwZ3V
lIXp7XBgtrRD/jR6md1tuRMfXtApTyiCVcDIOiQTHtJXYLAmn/ZUuzjAdcHvNO4omsmSWVl+I2cu
6Tk1TmK+fu6MHA2mxKJKnA7MWhhaX/LLQQgG3PQEyJ4uKonlMMOgRkN1M6D8uG+etD737uEmxYNu
b96iv17JoNGW52bVWsxNjNeaEofkNN9wP6HYl21eBbSSkiMvHirPm+MPQINKHgxMQi+3fnhM8gvZ
mnC75Jhi4xy7uj4rktHdBHeX6wBVQkk3FQkHybJP7ic2ePVDrpaRjhO6gTr0CaGMK/wwkMvUNzhU
2lxzERMcULJGN8T/hETW5HJKSd3XWJNItteBJOf7Buf4rIneYxehnYWdusZgsegBgltAzaGsMyBT
vO9VRZWNnwIzrTjzeimY8FQifsbpgYzbWEZl61EPms3fMo9MJPXC7LinrjykyVSYqIQ6Gzfk3i7Y
9zGTaz0L8DlrGcb6L858FZet0ZspFX20gqqIEii/8/2Ow2kUDge09XRxGGv9DzwfQpvVk3aJHOfX
BphwuHIJ6U8gcwiL1z1MPPxQOqrcTeI5dD2R9c2s8F8b8cxQe1dDa3Rj4p1JlpTBxG3aJLbUVdVF
ADfbpBxhrYtoXI2iVywYxDvhMDjpzbH7+zDNqlAlnnZDeFHvGtowW/ZVXEl5YA11LnC8DNc8uiPy
yWL5dRfiCMlJYP1yzPBxEPu01URIvV/dlkqoYXcVcRQYJPtr+YQ9jYFr2dpWikFkpcbs8vv6HNAa
/rZGlCm5EQCVP7/CswyaCNR+Zmelr5k9Q4TErFMrpwDD2Etaxfry+afA7+eNJgTIyRsHji6egp7N
RXvRHasPLhQXDT82mj3C1zpnJxcoaiNa1QchEhjKsUEtS9fevfSLHRoJQenZLbHvohGMYS8rXqy2
d6hxTdDUBU/FAzf42xUHOnJdA9+fZ3SF5yuZqpbiMzN3lJgeG93THV4/YhWdGt7XQOMyg7GS63+2
u/cC2zKvjXkONqzdQXBliuyfnp4OJCA6A1tFgryde8cudibwDKdRzCsiPeU8QO6SGior7MgO5wB4
88jWjE2SW0+866Rn3NiC/UzhKwNUViT1uYqN7EZQ+BL6Pw1iqjftDzWV6//rJBoYnn+oIk8oItqH
D2nJoGWmh3mTjRneZ8ybWdDxUGvMhgwbD8PzCr9FMl99/TaZQ014XJTTgbcXOrtJIyIfLRKP/RzM
UmwNM69iiTvWnX2NAy6/BUwfuvRM35wiMg+KfM0FOgqHL+dwepz2Ht0PE43iHh4WTAxuJasQqeex
N7sQL7NQ6RDPLGs0dqGyA4nrdO68wcV9RahURApOK1qPQ3Z2x91CtCuQ9NsL5VTmc8oXOQ43YTw3
anAUrDQ91/WMFy9pyqc23lyeE3UxRRPTawp5uPkw0Mw8dX07Zjj26f9HUArNDDmuTBAOiNS/L1uP
o5XW7BoZmghNebocRrqUC12m5r97ufWpYXdFSiJozsb0IKD1WHjyZz4VMNEMIz440FKdXGrx3cmH
iYJcceQGNj+kyZidCA0sbIWpWuvd2k56eKGd/SSl0hlGdcRsmVSxtlHXns94EJyJiuk+30n5L4j6
XKE/oKQ9XPnLTinIqldndFsLc3z0iMnNmfjLk+tSE2FntlMLWFCYCKcOtdkqPfnw/KkRaOZUVSpy
HgtUoAD59vSro2Y7BjAVWEC9ZI4ixCdzkOu/bVJwWXpZiTrY9z/bND7z14ixUaIq1blY72qQfZtb
azqVoLZPWwsdNwlsKdjNfUdCIaZ8FWEjIF0dtB+oz2cWyQaOApfGRapKw38TxFKpyl7UGm/ObE0N
23+W9u0VfH66PtLweQjRXzNxeuV0ByX3L24eboTIUg3SM/U11F9KgvLnTUmeyQZ9TIn58UStEWuK
ddqoADDsvg/heE5XXv6QCL4TmZtdT/wF8EXSQ4ZhyM9UN8y2h1WqGCWYWabaqI+HGYLsyEkjdacn
OGRcc8Q+MJxMHnt1wVkCny/Q66goHwRjunpBcWRY73YeyRr8xic27fR65vvtC3TAxSDUBnOABT1p
cGOTUr9AY015us/RXnukvG9MuZKOZdUhh/AvM4+PecaBsy6sH6WqkCI2iYmTe6B6zEZUZ4nEG7uG
Y+Lx2BojRkc7sRe88M6W3DzhWcWGDSVbuy5z6xUgFVIH2u564YiQCM0DMbQuvAmRyrljlv5qYnQk
qWKVhbvralKhbrhrxQq4lKc0ElZbROpOLTXIw+BC3HpuoFnEF6+cEW/3+/6PGXzvmziZiOFSihQr
ouIP2dkUGBHOsSkHaa2tJYOVNMyC9rYKoXNB/7oNX4IpN/ArkpMzZG62Md4yMfyH02RuTBtwXwYq
zdJbkgJHgL+OeUMy7JiXZw/kDRKSu9MEDKvWCPok15XJ2qMh3yJWuaOD1ZQK7ROkm4fZsSZ84Gbt
2izI7FpKuNUzjtz4bE5Bsdw1gsYHUvQiovyGyVNhJJMFyyDfZ7UNRd/AQo1GNUdjL9LQ2P3gIdqL
LEfoTAW1v7JhOdQsyNWtLZT9CTcvG703od++G09ixXOKpHYCCIIBgVf3sbKc8uIWFYmG89M2ob6z
zakChKBGOwf6nTbnPgt1VBIY7NpFt+wTJCXxtJ7IGdPQSUN/+6PToHyggEzG1f+fMWPLk4W5gFKd
Cb40wA5Qz0zzYC52oNfllzKTSbz4KUnGOIfpEWUWhNl95e0/GlaWYJTVvy3ODLtQiMUl04ZefpRS
iTTDhC7ofFMpYT2wuF0DPhrgfcoWOAmEz+uJWs6NCcBwGVd9/dhtEFLqSMgd6fR9VX4a/NwmD8dv
NZ2wVm7MR3K07rXXTSiHeS2vaO4oIJQbuU44VxPzNVkjkECwRB33h9EB4iaa1D8ZccZZWmX4sTkP
dRt7W4GbsDHER3D6Ru8a0jdbPX7k/ohOMFME/wkdg2qOy6KzZoQHjeAILczufeEgQcjld0Im1v0l
Eodq22cdhk194IGKNgIoquVRZchjvGs4zBH6btkLLdG8DYbrVIfToh/JJ0eS6Gotdqo5yXip1XWC
iF3LdskjcJ/EY3bgSW9dK9LjtUiia7TYgkJdlBfGHBg5LoUP8I8gpJqGBR5JIAfYmi5k6E/fu1Xk
Vglx4Yoy/pia10ZNgx9tycMJNdEUf+EdcOvtQmAXQzTQkomGhI7dTDbtPQ3h2yAfDisjy3d0700A
bEojZMYEBUD2X0EVFSzT7UqOgRByu1ti/uZFQh00eQBZCeXJ+EEMbW2ujbFvanIY59vcu30/fkHF
/FBsTchAgh7vMdYvAYAObZfzuarT5kT9mHcT5OVHeRCXp6yUBt4MkiNPyvq2tIxW539mJp1miTJx
kLY1h+wQnYFZNsze3WBlCm2qaZLKtUe9mMO1HYAnTBHMkWcF481lHUaSrLazxqFkKt2otU9bzA1l
iJnSuc4DxeS/EMmO8fEPCY6VXpipF9tVpAPIRNVDshyeir+vil9GTFhwoR373bU6xoJF1hhVEEKq
trcKBHj8rJB+2dCxVhah0IZq3e/YjNTlxtAgg271sOJf4qsjQq4zIkAusvo7MTCUKsXoADkeQVVi
vt1zVCsgs+cI4o3oTEFydVdbG3zjaCQNJZjDwUeDUBWs9EhEHSqcayNOzdJ+7plg9SQStQuwRgDy
xnjZCA7HS6ooGDZ68MPrt7W9kWC4bVQ4OVL4v5PrQU+xlewT4DqA1cKc/aCmHRXrQjpd9USHRf4T
/tF7v/bItoypJp2vZhrwwpbhjwXIh0tk6ILLvzH0Jd+rtugY91BvWRWEAWPhtnBSUWOsAOCd6tEe
fPyqmhXJ7BBDqEAXAz/9TRyoUljklGMs9Q/dFNS1UExquZu6RDD3dC1An7YK1O88zdPnFcKuwlMa
w5itGnzDZdGywPByCki41Q9c5Kj8VDUYL2fFq5SqeZMGe07ID21KbEMW0SxTancMh3YhevfdoO/m
89FoDLISKaYk1IZG7cs/IU5PiKaXtVGn4JMYJt+FK6pxGbBbQJHXwUIDf9vbIw6Li5+LnNgaPX+R
ilCntR6KdnWgpT47MbtMQv155dXfz6abXzzGnz4wXFYSBDkBEgL8AsOuI8a7VF9jKN04N41chPmB
C0ZK8Mw91SdiSNk1kKgM7x/1YzvpuONFwXHjHxe2PNvISUKz+NXTH6vNPyeJg7d4SSsmi/VW68DT
1f2gVzDbZkNUytfyRcTkpCvbnrxLe6l88TZBDYz67zhayJDWIfcZOAsOPJ34U57lVauxt56592ne
whUEFEr3vFZUfk2psL0cIihDB+nEmnAhY3/tFMXxWuDZJzzJUOWJ9XgZtfASDqz3l3nMf1pin7OJ
5u+Q2IXTHMs5IPEzduaXMSceUBzAlMRHBm/JK7qdr90cGFgPSO3dLeQzx6domkMSclJSRZCzB7SD
Ldg8pGOFHL7fCFfeccxT5xNWAx1OKZ/kC8BGFyotNUcFfFUGVGb5spCpiDkniIntCBHDHkMCMxZ5
S+oPGe5H+IG9FIo7pubJWjHm389isYstHNgzenGMV4wUDRmDlL/048BofO/1E+x+zuq9hwipSWqr
bXnaVHXl3T9wZIfr7E+mAgT+QqRKjuuTOrO/KaFDntyetLsVpBqv6Ci4lK8TybtLoHgKBiAr15Sg
POVgSJBTIF0FzqGIte9IqyyVScCDDMUUKA/+PrCucS31XjkkMXYR9DQCJRKBp2OKrSbvhLGZRDZk
zQTnRJtLa3m0jaldZgnSC5NEo+yXGZCyFfzePGI6uxGdTvEndSurnat4tP5Gz3QRq39sn8R/iPp7
KNDBoRSyVXAJFrbmSMoCwZJUPAqs28oVCGk0JY0PRKkKS2tBlChFXKI5i8nbJTf7DjqVL5ilogYA
lEiEk7QIODDW6+mx/ebOneHCx9M5HegAw1/KFKv0/RE72shUruW29M3UbpLF2Yi1n8X+9Zy+vYLr
Fpi26JIBFirOVXOgq2b1Jrgk27W0GNRw5KwdnVlgZJfAy1NyTbPz57of+61UahOENezHpUT8ask2
HDjGgGAmQc3q7oKRrGkAnfEZc6l+ZFnh4yb5295SROCcJzo98xYhPYMuoM4GQXxi8Ld7i2oM7tM4
JxqFfAJSOT9BM9oE3lniOApxP+kdB4l7MRkYIZFJE5CnBSouBgIVBbSXppg/ioeyFU2JhGyzj3IV
OSKylaeji/UieSkPnbVx3MgDlrNNta1f7upFgBNSipm2IWirW2tam6RRN6AqE3i/VkoQVCx1ADvl
sdOO0ZtCFwJbObRV6mAs5fe6cMBhKiNkY9nGOmzQayb7j0ApEGVWrj/Q9dh2/m+alujVCHNgHHE6
7Om3ReDH+Ae0BqpGQxBh0RM3y7bNU3RHf8aMYFeHVugiG/i7MV1wEzd50mkQFFUCUmx5OyFf3Wi/
EU8zaiuO2aDyI1aTROOoK3Dkw6lTNzqOHswCOfL20ZjIk7Q+AysdMqoC2f2/jQVA/GwCBQE4KLov
MxrDa0mZdFXECJPVo4rT+UkhOp2Kx/TFvlx1GlXrobdLe+Rl0zx9X6szbICMKUWZXTVRLfS/nTQ6
62sJJSuANB5Cd8/cP+U1gWy/aY0Lbd8DLUryE3eHy5J31b+Ko/0YN2u1/mtRK0r+SgLiYsdosNRS
k1S29ks3/iNqcudeaCrifh/hOv7PSBSo07hvXRgRIPg0m8LIsu3I5YOjmzPjE99B2O2gc5q9dVle
e+e6nT8Cl93QaYF9244Zy7FrYc89Rkr04fV+7ozPwcsXQv5/it0h9eGjUQJjWcPQNQT/+EbmCD+Y
0+of2lsGeVYWNFJxPdA0+cy5GvgZC5kag+n88q6xt54mUyrk70f9lLGVvcrv4GC48pqK1uwF27mP
1zflMjQd9rQ5E4nVLD08R7xEbgMunjuzvTk5QY2eaXT3rTj1A/ko77PraXNNyRa3Smq3avjAvEII
6HLYeWnV3Y3bDN7y2LsGKKHK11uH40RH3x9rbkHtp3+2w4c5hZ627JdNTsvmy4jx80+kFx71Fs7q
PMcfAjwitgLO3i0yIiLLNLw4nnjyN0TP3unvd7FZ0L0UenYgEKdA5diqbx9niS73J3z3hvTSlrVl
dV/GybgHyk8VWZattRGE2WmNkeM39wGbmSTiZzU+AQWr0AaEQIiyg135TxFOU25xi3tqziIQ3O5J
OAY9/a2++4hdhJ+bzXnQThPa4eeXWZKN3I7bXnWjj/D5wqMfNfM6BSx+ABhrHqgYJ+Cb0o28mItK
+KbcIhXFpb2Hvnb7vJc0yMNkviTzTHWw3nXWWKsMj4NXs36hb7VVJTM48sHh7sy23m2X76oOfbXd
iiB8XGa8J5jOtJ7249a31sHaOyb+SNipIK9Cz7xy7bUDFmIP5H8/ooM1V8p/WknrRu98dbPOhh1a
eLzv3U1DN8cEpmby+MK/op2nPX5CqXUp6L/T5nuHVby/KQk2ElhrBjVJB/Hezpytq9pJDavZvIcL
5vhzUGyqZDUJDFKL9BJVaVVdLqCnex74HYqaju40GF4jK5hCAXL1JTFcVysy53ufJ1/96SCuJN6V
8OjR330sa5dOpyBjaVgdFD9u4NY3p1a0nY7L2jSY29yFeY81qGYbyn8juPaXYEeiRxEAhhL/Rlhp
DsponmEHjQOqQ+Tg196ubyAhk5Z+Lq+Lj1AF1WHBQpnAk0gY5esVLVPN1tDBOub5C8mocHV3W4fm
zPDAWXyH5bvPosVipV87Y3leHTxuXXqq55fuN2LXx3b7nvdPu9XCG+/yOixwyIx8qBgkAklJljKe
9NTDKAVIKC6iE4bE3F/KTytDtv9wUglOUpTHWnLDSFYYbCeMgBTpHqyYgk1mH81PNFBpAvVtnghZ
o7arbd9IrCHGfhNCPLqRFl7jL004FHlE/HVC5zTZzcFKG74tNcEKypszomMIfnZDtnIHtzMW2mkP
CQ61Cm0R9HI4UR4i10iJZnMcnCzFUZJUHN64IBabyn+TJLT5FrcrVt3H/95Hh5tlQqFtBX53lyVM
7Xnq/kgH8hFfQ5POQPP4oW5GheDRdKcenF9P+e32jnGrRAqqEsw+0JK7Wqufm7dx8oNG43lOAuvL
gA13hYXvQz60rJcu74dMR/WoHjijdhjNRQ7h7JjocUSG1nwrvm0xWTvtzdT/IDzCqR13DoemZib+
4pDGwX26+uS/gWaYcN2Heo+bdWy9NFURwqSUTGuS4xtBUmxa0dbr6iKsc2iwN/QTIYomZk9kcJ0k
kauw4dQvcHx+iYrwblSn1cIeNhS+MHxPqn9fZNddCgdKhusRwnNZNKhL09Z3dUmLL+rUJECU4Ct8
I+R7j2JWhtKRRb4eJjXrSOGeAhFR0pjYwhwnrxu7zRzpqQPvNrMURhHjX+MvuZvoGleuL+jZ8YJP
dy5BaGGr5rEksKEbpmaT2N64x7cclOlz7JRxxrsAGedQLtwxCq/us+Wgg51qgRljymHQGvXA53W8
zAEv6RsXxRciI/NnZMXdlpb4TuupiHTixn2HVVwx7vpGBBejwIswh/GpSAdUQdj6HQxySWq/RXQN
0HOLfscn+udTOrFWS/MjsWMgAUbomrMsQh6eTYW/VM3/h4MjmrNPKNV0i2GQX/LmegwqYBXrVdbq
XIqrWScbn94wH669+UCBi4EJc8ew27C+EuVRMm3EclBJwr55GoS5A3Hsq/KFWwo++wGxVjshTuhK
MbhOvgnwqWUTCu7zqAYlvePLn9uU3juTdJrriy2owiE47eU2sZB7IVpB3s3k82iaNUlcYmEZcv9i
ohbnPIAxEI/bS9sau8/1Vixgag2qBoOi267ocnyiNvCQQ4+MlhNXCmfKsLTKK6dUVsQREQlmOsL3
czWvQ57yTA+nEZz6OIIPpqZyxsVB/XsYmZtEX7Ojn+XRk7If2Db2WBYB3N+FdcEanZZdrYaNaGRT
r3vdlxC4iQz4v2IAcb418k2+vZkM3f9LSDfk+G8pMnqxx1+alGgRnJrp/o2NHHhNXXBkwzep7PhK
xdGvNVMdsnefDMIADXk7LTugsk6anuF5YLp7WmKswR2+lohJuMSIhtagyDnFfxv27KXW57mGRj2l
CfPyUZrI12JpzX3vTdcR+JuNjRSkjT6q6IBnfRV1DgMv5ARh0MQlRv3PNWRuMNnRD2oxF/FsA1Zo
aG57Ju44YbGhFDTAeIViLptrI+Z6tEIjV9orPjDTPfnNajexKhRNSW1bFQuiEZt8t581mN9vZK1J
UYnRE7vyMmm/1SRbcPtfThIVPLEV0eRHpvKNqrImpeHf+zoDosHoFLYJKztqEXniZcNF7ip5c36Y
Btjo9EzfMmLMqHkMJ63voODJ44H4+Z4+PzmjwY0WpQ9kQ6Q1SESsf/vH7JkQWz0/0sqjdODyV22N
mNBpSPuRM8YkNg1z3FximCK+N8+RQbbY3jH3g7X8l+KqdEyE0XzhokT3Ev4lTf15bmxWjTKtwfEv
CW9/i3h3IAF5eFcs5jrt/3eY+0Jps4Z6/2Zv6rzV0PH+Rmmc6WOzQtHeh8otAlWqRQoEe5dkY7Nq
umOPWYSG3bTXOfQ6pOIRllyP8p5HIR8eEj3eV3ovGFJTyeeLh49x97tFjzfRwvv6Qbk99nHVdWou
ApvYIiL7fGQBS6mWYSlqrYQWyvL+NppqcAr993QS8rrjSplN58/oSj6Jr4+qeQjGXSnSsZgumK13
ugIiXjcIUePWf0Po6mp/DuRZoOg6y6PxmbeS/5fNYbfKsZqr6B22cGJXjVZU6wAJzaDjzByN4zq4
vAuYopjUhMjXIpIgXsl0HUu3iI0bN+x9/MunOyElfZ5ZMkA1r51hgX5O+fwpE6bGJAUylqIglB1D
4MyxIvIJWtQ8ob7FEjh+W5+nx+0/i/UbFGOhuqmE+DdV1/T13cnlwPOVLOX8cM7Gxw3MXl1YOKSV
y7rTPFjQ7kX0TExWlw1M4Hb5HmxBP33TxgAQDINBAF0nvNtpSp9OstwvDaZlaERxj2m8H1e1IyzQ
HtdHQunJ0smHVCClJfEgcoIPVi5yiUfSMNiETsDm8H0Xs8YaGFlQ5L3pFIZWfX0RYGHnWX47vaJ8
chNgVNRHagBS4zmGo03lIZ94HMyxhDiajlIbwKxnE32I4pzvhjm4XXIJBV9xK2fj6E5lv1lWumzA
UI/WH5/lLIvgwy2K7hLBtvmrf+qWEIE6/e0aXhWbDNJPD3axA2b/mTJK6DvQxHp9vbAtytQgMGxm
WIWxEb+IjrcvVgJjMv6UCYV64cT/bfKSqKWxgBse6Qdr3qz+x1XAxl7Rfjck0IzewzUYlqNL51YF
Qh0oiJjPS7deFqWNHAcAzShGNljUZkJCctiMHF++48kK377Gi15ANp3OeptDI/xLHKhX5ycLeixI
IweR+PwgxjjgnYBHHlH+U9G1Tj3S5vBpp4chDp6nVPcZfzBjN+a2ev8BYuzh9x3wtrHEXvaf39MQ
JHiaUKZQ+18pomIxabPn6nlv9n37JtjW4gRd9d0t4V+Z1H+sj2tvu8k2p2yOcZFeShCjpHKDJL8d
g4KjdIofJyRAhB/lfRXTyVzPbpP+0oAU+hK2LGB+shSwV/46Zf4K95u2JM6BIyOeKuWS1H2KXegh
XZ3slB9p1sVvozegLVJQqFNEH8WYXlkZffGjd5Qj674gGcYFpU9fDQao2qPUtw9wCJO1Iha3SiAJ
IJlPdwXowgWfx7EZ0ytHdvjxigRCEono4ktrompEQhTiNwAjEjO5Qi6AwiovxkGcHQr9TafblX0I
YwbTkyqVAUwcHwlPxW/OuR4Mng29FSxQg0wOsu/8ThJBAY4psCfbo90xop5j4ciLMtqa8uUk+hZR
yDVOFQQ+EzT1/oZICfwPwxXuYDwUU8W/lYmMC+ds/16qo6pSJe/5ircP9WwzjxbUTGUw9btxr/Sm
8iv/r37luy/+yItzTyGvETwfREAVfS1R4FwjMYxatJB8QfB756B14XQ85bKWe9Rdg5rOEsb9tdQV
7IVEFAB7HU6YWZQg1Ryk/OGb5CUSKfM+Fr/+R9YlesTexeOd/WVuqnQJ3pwPl3FeEjRfTWkjOjiF
diQtm0pydOBUFQ+MRFaGBrZozOt4Lwa/KSVRE6/GpmsMR+Fg8C0wuyvX4OYyS/aEn90WSnyDeZTP
19sDgN/86KERwejneLbeIAI3QtuxPFFjgxnppiKC391GxV9P/C5Qjz042SnSVea9uhOyCT0D48Vz
0HtHm47WpCNVzDwwOSEzU1RC0BIrgjmHCzshZIxjnnCqiOCAiuGUu5BjfQScceWRGmuOWsgliK+O
Sf75B1v43+elepPxyMJDGQDISMZ4zrKMKxK+8YHnsijn6oH7FnKKjo7XMf4pRv9tmS06YlUoedN0
8o1WEobYlZrqZGfdeSMwWQ9n+zu6CFw6SQ8G0kfvqVHmOHiX+ngB7y3aKY1AsCVNnkQHWH/L8zbn
c1wYVkeaKtYsrkxcZwwgjjvWogkiZ2Q9N+0Zk2RHvKvMjrDpe8oI3//kT1WYeFI9F2VwK5X5Cw4P
e+cCsQYiCD376ja8blIqqRHW327AAcUphBEd0TT8e3Rq2A4doWKsE8zF6xA4af7Hk8Fd/jTK19iP
SZm+KtuBC2aUl1Kxyd1PQfHbSjXc7AAZHbXQxV+KiMhpwXCngyesM8iG8SaJ3oIHyO2jm1uIGCRo
thA2tnu4tRpscV9/onl4+fqxvyId8pkzal0OyptiTDcxQF5eCVtW/1teu433Qdt/Zrm2EylhL8Z6
6UF49au6t+G+wdGXY8lQjKGHMoD5/A/X+zJfsMuSdy9Ew4HuQzCmBnSvEC+o1UYCRi8/9svMBYKE
6gF0C61x414+RTJ7e8ZNOJwG2gd+UWESnTpp7TZcJwisIr/Q3TzIRCzQprGJaBjIF83W5dMgRjRv
FUfDjfBhZgFDic6W6vIKBwabA46HIDWX+BS0EtQ8K35+HmQ7d4j5JiV9sjgjtBZK3wVUZXxXqvd1
jDkcb2+A0il8Rc2ojs/6YP7bHhHNLTxLUz0ilL0/B29IAAkHeJJ03YJP1zhcIukdHCtiUCwyOAqr
Mx7ENJPrGyx5tWvsQJgjZ3rJ2ZCexSbtoVdfZlQdAiuVY7FWdHtrz2khHA1KuvsbbNDt32kMEfTc
ArttKfjDhEGrceFPeELuX2DycFgM93o+hIWcvHIhKkne8nsrrW5Mf4sEJocLG68mhOZlGv7uKQ3K
KBp4VjIY2NjIK5vFS3hINSUafG5xx12eTLlDyX1U3Icp2avpoSWZfhiwsPYGSzKmuzj5l/MZWVLo
aDjqsovMHks6voRfSbeRkqZmaNOqghbomPks9WksXm1X4MG55N9vQAwIgab4AHbU5al6p7OM6z3o
NyabHtHeW9/k6pqEKU5lSsPdx7QCnlE7NXdcrHv5YEqhBqaUzI6otCuiq867QMbJ7ZziR/bTESrp
NkTem9Z3YPNxZnePYaSab23ZX+Gh7dxqTRUEjR0RBko7aKCBKjKwfT/yI1BycQZ190gwvPSn3tjr
yyKyKCS7cyIc3V4UO+oGNfd1lGN10a79Yvo8Hg4PTXoGX+0z+Y3eUykIv5aPUXN7pDYdXVGvcQzH
0xeA8jJQq8r1P71o0KAZHkyaFRuTundxRtEe8ZHLk5wJxLICwCtjm4m0q6QS9YUgPLDjfVubUHJo
RFio8mlG7sT7QNWZK6/UyefWFIwckTslbQQCW21hy12xPjiYvCZfYUWP2hvPWa0KnEbGqQasT1/w
PGpOe5kTcBMwRsU86IJeuYeVd1Hx9rr6OSy5KjhYRmDxGHvYpyGfCW9caKQ741J16foF+RgbvxeD
a0O2xodGE3udw84oXcf44K6rtGUMa/+815aHFdV0nor6sC1d2TLmJqW5GqUXrMfWHp9Pj3GmxZQN
hIloFQ3iGYlLK7/CkLzsm2nGS5xDjUDl2eA7qJlsuo3R5tATyPPe0XHsp0LK5MMLYoOzk44eWiGQ
UkTVp7jBtsDLtmFswFfBXRIqEldnob6GMTrx1scRYwNTes1ttghaKQjolRY6219l1sTVre5/ryBu
oTicI+O1p23caF2X+JrV+fIiPXlmqzh2PT42AM4Y4pVu2gSIuJXfm8pq640u6nWFULUJ3h2j3AEk
OWrZlLm52u7tw36F7EQBEQOwFx7ovfsvMHRSa+SPk4WjUX5nKhFH7AlFeQDvoksdX0CaukzROBNF
ZR+4S5W7AR6AS+Y5MXvC8qxtFQhhndTBGIElleZtujsEDUh5gp0jHUlmRv4AxHJ7+yfj5R6pp8vS
i2STQ3Fmp7N4+MV3WLCwkHvsTzDQE13QC+2Z5bbPPMvCaKLwbMyZaMYawp39ZFFos0M0zrDjB0Ll
A+F1am4gOpr9FyhKGJqrImr88c+r80bTmilbpZyCaLKwiZXMAyswLtgfD8Y415fMT2bfC5czsxfI
O17TLLtVIK3pP50FFs37P5Y70w+fhrTDtn/pJbo7Hb2EMT3MgTcSHkGeOtpJiegd4RgDszOfg2rl
yNX8rNphnwWJyNLL8TtqceNu6r8KgNAL0oPU9GD4M4PTi2uVti2C3oYCeh3snSfcBkKhq1GUkyj8
uIm1EQc4qmuN13DLF1kyrVaH5z4HjpqdhOKAT3KTz/Azw5cF1m5tbzZSaVcJ7moj0zSGhFjsMRYb
lYty+3aW+Z0tNtr7k9vws3IB9WfHoCaP5nBLfFObz5w7Nog9S0Dk/Atey6XILGjX/IBgA+q9m/p5
VVlHaoXh72zrzMT6aNALAwQW6iqbM64ofxv2rByxI3QJ960nSNrjwFoZoDZ6k7pdgi/boS6Le3jl
UODGhRVYGoSyrHUlZ3Xrfzn8DnBb5lm3jxv9FwOOygKeKoLOghKb+wOW+J4hBV3FXrxW+JJ5wleq
ytDF4l5Vddu5KczIlWzt5Zut7etYLE2O+rfILqR548AEcYrhix8sOu1QVPAPrBByXeC0EWHhY976
MC3Jcc0XOr78CRl14Fm8wrrZNClXlHFS9qS4rrAVRXPYqQ/vEWv0R36t8tFFprRKugDysTNFo56U
JzF5SKaGHr9knUnhm/C3zxcb4n7TFkNuP48bgbT5chTU2OlfBGxGc85l4t0Xg5f1JyYBSMzkQnGA
IQh2Yl9wigi9TdNUpNHVK6u0hl5yZ49DsTfs8uHIzGOTfT18rYCSx70hp3T9Q7+xb8KSuPZHw17Y
MfHL8Pg3EsWrgnQCHYV/y4cDRlAz1DDS/91N0GCMu7cKr0ahDI4RBuXYU0qyTFWpdQhUiu2a+bME
Nhr9JGZ/x0k2802K5eT6S2SAneiCfNQK+i/vHEdJrZkSL61Ct308fi4oFsHampgNP3FuT91pk/zl
vAaUceGUl6dgOraSfv1EgLr+UbqU9K4KMTGwqNOIu3QU4zVamdnLlTZ0i3kZn14ABjE01yHKQslr
rWmc9974XCNTDOlGaRvhBPHODN82tpalm3CdX3H74thxlunbsgounnVXRmhVdn95oohxEIf3ufs8
4SMM6X1GFciHc3J1kuh66q9VWGnD9NsLm9+685s6U072H0n3gc4ju/mfre+V1OHZLhXSJ5Yfw/Xe
XkAdjDtRMKNWyQ9C4PC2oDNThQzqBRcLC65Hv1sP+Q+DAadxX9V2ERTVMllz1WTaWWiYUIASia4g
mLnefmYp2izWhfcSVuR8YUxvqa6VMLgamNTQiyJw08EOl9Pn8x3a/zpH+je/XkqBI37tra3Q8xy5
fgcF/NJXSNsmFdPJW8RY7RGj+QuQZFK3bWlWFIvcyQGZa2kojwbaPayefbjGVeZMdcm0Xq4bwVr0
7Z+Lkyl/DjamMNF12a940ZeiPp04yLIXAtj8O5bHA24PoJdMLwXNdclX8YqvaE3jc+9FidMbhwEn
354NpVkNrmOzGVYD02gigTaTPYbrN2BnrbbBMr0ek5tu2qNgrRWKx5yysiTUtoOI057LXFAH9/XB
MZ17kyHsIaQKSIv/2tKxyS9hY1a9VEsXcNWJDXbanQOrUSKM8JwFxJhzdYgYkdUDSWO9R2pfzIRI
mcMT9KWWqhvrH7Ha4kdnrQbhoK1Q/pSNZgICuHJn0h8HUJXc9JZWDgmxKiz0hPGWxu/FEMfr7elt
VGbV8T1r/a9OW8tU2rOZp/1QRJOq+iNPT+D2l6o2ycFFwqIMj4R2Ug3Xe55gkirRcfRrZp5zhob6
V4g8dlyMUzjRUks/vVE7Iymo4KLSSi8N7Oln8TV6BwjCMsCxCZ0QiMlXVi48iaH80mwjaGtqKXzn
rIvLl3anLubcGVM30zaXoMfFp80Ii/LaXEu2CoXuxC0zwMCR+aVcgmu3T0MPmV3EF44OOzd7nhfy
aFkgk3BemZIWurK5WpuNrMrxE58jNnkkKxYxvgGcObIZo8UbFz8Dbk6WquZ/rtFo8laUVAl2LneK
srti9BaVy2qxtJvlspQ/0NYArRhj7LwGN0dewvBLA0jebXtUlU84LwT0jMR97YoEO2kjT+nmY8mh
5CkbjoAo4kjS5WyoKfcJE1gP6rYgNUmEv9t7JOQu03alR09TzbToToVKxNgQl2D31zn4HqMWO9yA
oPvl13agTo6w+GFdYNjiQSNirdkAJTOP/nBJzubr0teTb8VEvQ7g8yFOUs5hIqvQuGXx0w4uVqL7
BIsneBG3/il5k5hJMy1dRmcHrcfJeryNYUOg9YcqsAYlfSJvqWGFJTzrpkD8LJRLGfKm3ZYoMyl+
FXcXiiG9XE9AmRDGsVq1iyz/e7lbXJ1uJPyRpSNRWw1ZTlUQ7zQKRL5Gx1UznCSocZwfFtajNB+Z
qMdGamJxN1QRZNkKoDua0ZcbA5QJPliV3Oa8fe9XIgi7x7KIrVCvV8h9wxTYIVbNcYdTL09RtNm9
mal3nunU9HKKtzSaLKHz4qHeea7unEkjq70fAGkjbeRokalrWwKAbLQHYzjeQAXcF0VZo3Rl50L1
g3AfJFWKsu3VuBNDDw6o6ou/LTFr5NXKPYu10DzZDwWu4nI0DUedn/b0FyMlRXxqseZeMAA8sClV
YOrg4OuhfBb5LkoONHLQMlXYce5H0ybQr2uCFQ/4T6wQbzt/YiJ4VEDkc8w38OAfL8y42nvpPDVG
rvPaj6ezrVWroiuuKvLvphsY9lFgPWJTt9/dL5nm3L25Exxt3foOJDLYGBWIwxs9Od0gaCrsWodG
Ozp+SXq9ltoTYnFezB6JMi6Zqy9aMpU4oIXwGF04aJ7myqaDv+rd0OMsz+xFNObYNFnQEOZhAo+i
Ym0NXoeR8+IuK1APqCIc+g6/z2mv0ggPquIMaa4OdREpSdu5/Uewlv/lGt3kWEhf3JuspI3wzb1J
3jKKLBZAN3xTQitfdEzRVHX/Sd0+m6YtbrrFF4phe6RcZOqlB3RGve/XmYv/QW2tmiDrrutT+xHl
wOquKN79Us7s80EjshL0BYzzWuFqXN1wIJ3K4qtf3Bg/a5va7OkyoA4gPY7wOn+E+GGEYEI/0I8M
YcEfgZf+DWf+mw3mcKaXgB+75e4IN/qhMeiRsjNCqyFd4u2aUxvJ3VBtmtsq76Zr8Df5sCJn7gMS
xnVB2Rq9zCDguORW3YXk/gEP1H1MUgbaD8yTYlWUbvmvl9ShDemZ/xuaegCeyVcfNt1OYRP02DNK
1ME975HraGv8GTzuK7L9ip+333/uMZ7leZ7aOoYmbfgUCWgLEJJXaFYZw+Rr/rRXjIe8C5myUK5o
DN0vRSpUAhk83eZR9Gp+hL32aRPawD+KmwtkF8nm7OBrgaIwUWNIGq2MuyQOzq3YMGKCopMhTWL1
XostKpVLqRUkAfQnZ8QvgG4zQHXCYT7fEVYncTXnzkG+Z7kG5V+Vjo1PgQzeRQujEaLIBgIrL2sQ
RJwHBuRKjQ89Uwf523ARroPlqiu5aBdne9QlFZkMNO/2Pb1crC1NGgeV4L2kuvcEjv8pFYkg5ax0
H/OxFQjNGk2IzHuWeEWlaMHvoAJcvVZ8vvLkLoRRezWKPML9OrRaM1Tv6wBfepfUn36/jcAOLlmH
lnnUiSM8CUN5mWdiXmfU9NpmWiSqDrGGWS2HivuDN3TAN98UZPsMfjilx8NWvc0HhFAOMFqL8Zsu
5G/58FiP72IgmHSmfpfE6aMxR5OGJK401e/XLT24C2Mvh9cNogZxjTBJsow/ozZwHtAshf0fP22J
bW5wTEFjiYI1zu8C0cCPEcrsKKVoZoLOGoMR8EWCIQw0fLouIM9xoqtWvwg+JFd+bTUUN4OJrLnj
ye2ZDYDQIyz2P6oKD5q7ZniFTR+encHTd/33VfGhkeFWPpMC3LE7WbLCRpK+aElcApzaJMUTwL3I
I5paj+GiBQFR5SRH6I2SpD5e5rQD09zppBJmhBxEiN/LdIyNU/j8wXjLjN+ZMde/UP0Qq6B1C2bb
uAHQKLVgXoLSxsT9WF3Mxyeq4ZBfQ1dUI2VtShBCh2AiPVlNgBw3GC5V5buPkaR6E6ubnXk/SOYA
00iRaMfUpqpI04S4Em6+Ke8CVNYG2968FudSAvglgw8z4NpJh4bCxmdG9tjDj+Tkci64ab+x1wrZ
eix1DBnVSGgludjXitDyPbN5GSJeVE0V2BOW4Wc2oH98nMBZfhmUVBjQRmF5FPMKhLLbkwwg1oWd
ZVd0mawlO1h4XP3XjGD/dcUUIc+ucOW9vj6ItB3DECnLHIeUueZ3Bov2qhp/u9LcvmtU7wDaDEXR
4eppGHTLcCJZJhrweIfGn0BJU8g6cplWKdX4xNvtAU8EfC+gm3UBWfF31oQsFBQM6AA/IH4Tx0nC
79BPYnq6Wx2wgOmgt0SE9rlIHEFWrsxPUmgKPXlO8SqLWQ0GlhC8GcXG2rZ9MGnOehytVAxhc3eU
KjrdD39R5KGknvDxwaYNDsW8l1+ozm2PoCwN9mYX4pDxgFosZ1dbGNyNWAxZufTPFa+F7y9yDz3b
qskQYF0s62iWjRaDLQ0S1w9rqjljt9CGwCq+VUWs7mTIF5ZXW3UCyIq/NdGe4w0R0NYiawAemUUx
3/VodcgbHpmqQbSzq72e6gAgG0lnDZy7g3vic4ai+0vWNti6q0k0Ghzd5EMZwqpjHmq9mt3/S17W
mN9G4GMhcqC7UnNxOFJom6IYGYfZkIIp/ouRTFy0oQALXgRt41tJhytZvvsPpc9HCBW3OmngOONI
Lqdcw3wP6ViRztYEjkNM2+GXmv0YMUG3Pyv7RDfA1uPWdPAa3aVHZChNLZbmaZB4YX2UvWc/qlSJ
AGABe2gMYuHGeeF5TFfOGisX75cJmmHmRKTz3aBNEqTn9j+Lh9LPPUaPlpHMJCQc+nq/X/FtEpPK
/0cwk2XB/919MYHOju108MGRHfwETVw4NMCC8l7ecXbCxYU4me2+AEtCrhL+RFX7Q0oJW4Lto+V7
1UGWkGwnk5H44Vr3RgketYuGl1iBm5B6jh1XrPrvi42jiTrltA7TX3qH8/KcX0tW8/YMeRF0E0+h
S/R2bc/iH2RRBZkPWRLQSvzKtN7ZgLnAx8HD75xbTjjaCmikcO6zGnZq5SltXHMVnHEM+ZnZCuXN
mRruvl1YgIiRFlA3zkWUlf5Pa0QwbYQmKqT1m8Lp9EyfKp23V1BQlZYHGF3vsWRKOs0b+H0cz52H
Iig4OzMiMXDaoLEzWSnOG6o1D3OD1ZDPiRbM1Kt2Kc90T8C83lbHD73wCFSbQFAdcfWaXNcblGcf
69fU+qcCbWwD0ReksMvXn0CSihDtnqb0LwzUQy4OvaNnlIlaz1yTrhlXsfk1WGf0sHrCMMxkdw1I
SXxd+IL5Wh5hN9fABgCCV8bRGLRCuuVFmcQ4q2X1elNwfjm5g8zkb4vOh5HGnppzE+3W5g83fm6P
/IQcIwo2VFvCho4fjUi/W7lgNCf2SIiqTh4/A38LS7vp1xYp5YPbt3K2e9ZfwBm7wtI2UvzYAI1O
MiK8aOxddhNLgOLrQ+pGZgBx0dTjtukZXv/EjrfHZd/qN7wn+uvs170n7Z1dMpaZmJIw0HhiXQZw
uBmvXu08hDqalMhHDp4dYzcl9Uqg3z9/T0/iA1CHDFUbcZ9O+8qU/sJgKt3XgmjhcJ9lVWPpYj/l
0VlzoITVrxZdOpNheyRCgLEnsfvsmdbWVL/z4R8NUgIkJJ+T5ujfKEf65VgipNKqs/r3q4tRVYMd
TPpezEcGrUWO+tKWXre08GUQq0b24IHp4vlUaU5djUsip8Kaol/F+wBQ7O2cJWjiQTA8NVbKZPBf
AtvUxztwMmpzk1Rhn5G9NpGL8Cs2ETlRLmx4bsbfcy08Y9M4D7FDYRSM9dl3Cg8QkSBAzc5Sb+oz
HHV11nJKv0jsHfCfIJrN/+qf4CjqSACjXmLaYjToE1t4tCVYbdYda/aPes6bPbQU1aGdCYb5L/d+
3G6pxYzV9HaSYjOiOt5L09646dtrmEXzXxu+kNyJ/D4eS2cGNnjzjOUEV5aL2T8wYa5EtF8YkM7k
M4Xy+6hE2YN1qBmnzjDXJ13PXR1/MpZKlYmXma+3/hjw8Yf0RUcY5qaowhpr0M8Ui0aqi0h2TrLl
enq7md/DPAwTqkKyWA7QmcNI/+tcRn9W2xUL6aUR9/5UkZHgKfqdrRRjCErj6xRP93T+9xuM4QgY
flfJhtGPXs2ZOEOrJSyDNBoY9HXDSnwGZJtFrLuqXRaN70yTbefNHrpGNsGVTbsCaQ8lBOVXz3kM
i/RCGpKxDMyucrDcYkrwDq+QinmN97KJkgNi5Om0hwgLirKCecJWr4FAWfHPCLQ5UL+gYnlw2PWe
3jNZP+3oB5v1NcHssJQapwq3zOPBo2mkTiwguTC3iB0woOh/iWUqPs15uBa33JSKz0zk7P6RIXM5
OTNv1y9YYP3WCGXdNWgIgEn+U9B+dSwBI+GsoxxgqgzSouO+zaaNxQ+NKMoBMm2h1ZBWENOspzLV
DXbCxjX5JshtgtCIbBOVVb4yNvOlOQecsBc0Lc06ebroWDdgMyRjZkXqR/MeB9j5/L+llOW8VeyK
TmZ5eAvrmp3DDenK0tIiqFgnIqnwMwA4/WlbKrTv/93YQp3c3UbM2Qnt9l+rWpR1X2cA98H4e42a
sUxoU+XfmQiw+QW8YN/kFxjaQwCVRAK2gHMafkLpm8DyFr84gYUGIqcePZ2nB2s/DXZi1kAuTpOn
6bUgBg6KZf0iHuI3rr0BuxNWv/1f6t9XEX28laK+yKF4zyWGigwW3AdDlDHpi92nzkf/4jKUYY57
78GdLW6Teks6gPlO0B8aV/Z+55OZqBuvzgk1pf99QFjekGDmr4UGIEWZu/VzOLaU6sjKqIVgjD5/
QJKSKxsebLwZdjQJTH3VanBWjMF/VG3rPusHFrJZFHTONWoJ7TAr/eZOuXBcqh5S9C9/biny0woU
gCNrt9e56NDXl6menU/KVAqVzYvDv0uP4Kar/wEKGtELHWjvUD0VP2vxfzmvc2sNTfnxOmARyam6
jdmTBmHKpJLXW8QPXDqs6dOX5+HopApXxS8TQWlWLbd+z8VOeIAn3xCS7Hod7kzljkm26p48o3c6
3n1S5T5DlpCJ03DpHfaSB7HUIgplILg9FQtisODfFtlGdp9WJ/VvwfUrapxwA0zBulQ6WYYPv9tX
C7uTdXeAMKLKswOzCyYMC2dx1uhndwlSm7WVNA9+09MqPSigxvs+ZLTqL134XGhi+tq7VlyHW6Sg
/OMZwaXPeRPGvSNcln9kHMSdPIxMt8u9P9H1ILF/CFYtH8sHgMEbUswTjUwM1246nCMmXzecusWC
HlX8Eo70bzuRM1MxYsRWlNI44SyiEhCsyIRuiM2JPG/QJ6iSXXP940ffsuDjwmeyLtU69yqdylIM
2NYTMwizeWlCPzmcoKood4dLRiGn4GssOyNfaRJyUbmUe5ikxf3IfMoykC8SXowf1/nmXsJeyE0h
iVxdNK1yycpb0/IGsR2oIFkeM5THpEZg5hR7fuRNly28XzprDlX4QmmW2x1Jn4uEMi6Mu4HEshB/
HUdb+luGp/Rh9SMtVpxdysbf8oGbYaw2mk/oRL3LWGcgRmAAJw0Y5IpzlNZcZLCY/8elsMDmJ9C9
kREB5Ed0EeWhdQ5MEkxNFU5SpVC2fN1y7z+9+QgLOhBY8ww8yQXDS4b+Iw+TKh0gHH1sLG6n1ZtG
bP8qq4CIicfxfLaffqK0B6RAJCsBknB7ljhYG/KFwxadWZoqcCNaCBsDYM0DyA1szj4ImJN2rVLg
6E9hhjUVTTg/DZOmOFoZvwncLMry3oym43Q7PexzY8BrQAB0BYEjlidmCxGaYoxfKFSZDk03VEpW
C9hZesNuo/tZ2vV5nzXMLMMeHyrDyJ4JpEfNq5k6EWhkDi8r/+7kil+NNgtOrltYGE6vxKfZ6AH+
HiT4S/Qyj2Fq5IGg07ouV6ThHpO11bmoRsdzms3NFsTduQ5yQG3/f//cdmpW+m1itpUX6OPcDk2d
J68ZWRteWQL1S5eCdwyhw7uT09RF+Vi/7Fi1taf9L2u6X+qBP81EBv1HcCTc7v0TvfrSxJ/THgbE
nWEM+/EqwhWp3t1B5Swr8qBgbp8f3tsWUt1FvN6ISVk1zAvqFI2c4OJHuLCShSlidQxWKzG2bMKJ
9R8VntJ7kVu7egY8rVQnWwhcrwIqXueRxUJPFHPKWRg+hjOoFpP4mEvt1awuz04724L3+eNi2qiI
7JTBnDMxiFnkhY1fE9y3+XvlAdoJXG3mj78Q8w4XzB6CErEJq+nLOMDIEbG0CN/cKc0WBmv59GNx
FixGnwsVANtcM0hbIay/KseGOC6KHDe9evWR4aWtby+QGGQDpXzyhNAHqtv14iRSZlu5dz+9/6Ou
rfxVI1Qwa9MMvSaZ6j7SabVoDC8ZUOkQAxCyS7uApmFxRgLPS3xhG3JFJEmX+h8iM31GcNSatLP0
sOQ5qX0NUHfm63DFedLq4YNoa7FpRXs0ziNiJGh2BOmI+/taHe3TA/rngJAtygegN6Ord5A3iYnw
PT0efT2iwyLTjprxgTn3JQFyKLN9SqWHDvNWfNg5+SCu6bW4GpQUZfGnChDH4AVa5iuxQIfvI39G
bfHcV2lJwoIJB+G+MFs+ML8ZFio7D8mA/9GITqALaF21d5gKr5gJ7qvbMuZSWzDA0+NkNEeeU1m5
hnB0u5vfdg13/FnNdeMQR2t3Bsn+vRwuC0TjikvyHhdPiR/FhDsHxnVdzDTWi8rUNuERyJGOo3g6
T/HRX1UQF7kd0zXY4kPRxKwHOX1Yu5Q/bzxvV4ZKcSjdVNXtg8jj/EPUtCt+8D/CzVhl9IJTRugS
ACsHpuXR6p5lkMjl9vp86/w33uV7/Jspp9YLkuPtwoTIi0pV2w4BE3yTi3G6olrTSFnUWMro4ENW
3FWXaIe+Hk4tC8ktN7RTodAmMDBrQjgTyAGJV36gK433meEa15pExYXN6XHOOv8ewFO5eOkn+5TN
UQPN1pt2wwwawi2FEQqFgjetrO5H+pcfiv8ipUdDl7R9jReRqzFjgGHSOE12Z2TAoOfN4Ki7iX+1
HcpmRW5s+XuJNa47w5Uv3HCLpoBsjKcEA4VVHzd9KCM5oGr6wHTM7m/fW0deen/lnmirGb85hvg7
ANEw8YXxNYmiQbed1WSOcr1jII7Q4gKOEC4jD9ZbDncCvOwAgm6IiPasmHJgaURPZxTF3HDmnMH/
CLXDaM3gs6/7bl7IgJRqsjN/1B7ow3XUWSLr60w7sewuO73viWVYKXWViquv35/5y+s5Q0BPfQgq
5vbcOiSU/4hc3FwnWYQRQiJi4JuFsQEQNE8mC7IAFBkmQxBKsZ1ETk/UNfTodelm8t0xWO+Vjz/f
y5Mr3Co6AJ1M5fO+CHXcLLSR6VU9ljD8JphpoeDV9VG4VEqiALMS4cqq85DfeKVvuTeKDadit3r+
WJXoanWbSJe2IyVHYZw/M4e4fvbQ07GZrZ9ppWceDTN5rcrZA9Og3K0IkhW2JBGuPWjn8YdsRdcZ
ESICSgAPXWO0YKFKL2udztINMeHJ5pZyGHp8Povxhjy29xmW02DcEZ4SR1BwcKiUTSSGzed2QjZ2
u9VgFsl9CO4z0Fl5MFlBmrFzsN18gCaaDntPQZpuU7MWsldmP3Z/cYd8VmwN2oprlDJPHvQqiBu9
ppeVKjyCjPDwrn5B/m7jCjaeSCAJiEdYwtPc6lXC1Dq1Ix8QOJ8tJwFyi9w3UCyH4OgUMg1qfzQg
rzbG1RyRVn14zjW6lRatj79LSqfXPW2ft+TksT7Qa0KteZr0hokEMj8bCJbzJM06UCUwlkIfdXn3
I3S1tRBdy4p1I8PPHvFVEzyRqex01TN1y00y3RU3kocJSiuVe6AN2PcegbNcuDFJZ8VPB85BGRHF
9+DCr6Q1O3s1RuaJFtFrYF+0pgVRzJx3+waig5mNpIx+3tvnB2yDrAWOnWVsyHDLwezVgcTNDoAQ
AzzkB0yLoH8POV0g1lVqBdJ3plLd1K08cL0de1Bkuk+Pm10otnDMvZftQfRS82k8gK7scSHqz067
pIFlt2PDS47bVzl4aTV0jKstXhsWutPg50kod7Qh1M67Sfm2qJd7Q+Wa5gDNNIbozKIRuCeZql+0
2lBZttF+b1JwShcHoTuKBtOKcBtjF4QGgypGGDyhVSM0NIWd5GU0WZHEX7SQAA/A1zN4InXxAvR8
Fvq1O8FW327WwDzmOJe/VnxG9/Azq2yeFPV+XYTjoZv/Fz2kCh7yjy6/abA3a4U8Dt7lPmXV4eWn
AUGyMQKhr+en3upBaE8hBKLAzSyByIFPtk3xx473A+34ElC6Tgkc2NUxQ6qqy0S2H98FIQWzjdyA
mr6GI/bVxyHC9AykX2ZPk6OIUytbe58a5wVCr6KYQAcucOvd91iurmlFAQQM7m7pLau+0phmjQbM
8tOOdsvW9Au1hBNwohhlxdC1UYPbIOIaYNrTiEUEp7rrwN8eMhJRgKiD0/j75tPWMJ91ULfd0lBj
mYSMWilm7KYtEMqFuezEp/KRSSqLjJuS8CZiQmbdoqbWbNUnb+G7abnGLom9u1707pbesx1bMys2
B8URBbqFmCJ1bMWlwAsY2wn5mLVrETMzz17K/2P8cdtU1lwhVdiNbeN1DpG6g+IsElm0eqmEan4R
Rzj6BtzDxKupO//KdvndSx1X9NWZIKdNXl37dTC55qwC8rsxKeg7htKIwu6Gw8WbhstkElPxzz2G
novSEspzuzYtz+Mx2u+zBUR6MkYFcekAo0sRqQdvQqq7Q7YzBJODppAOnbwkMPhkcFHJm+/5kU80
jcDJyww6+9t6IKRRHaHWEE8KO0PK956YT+/z0XWMhUWJXG/plNPkzk4Ng5WLOPUbwslAOuhxQkgw
bRzjOE6XfTdVDio3txUmUBPHhzU7F61K/BXfzvKgYIW5V/kNWA0L4RPwnd0UEOkU9Q2NFpOtFoSJ
Mm4Nm+CK5a72Yw4CwA2Scu+W5ydR5w2uVIf1IYH/zkkAPCkLz/OWUBMWorCLcxG1wk6YhRVy0xzB
cDEYuYwL/ZmVoytThb6OVHo0jPWq/4UxMSvSGr1K53v6U4Qi7Zq3/xAMV8LQvRN03b6yVDvEGQag
brvn63FE6mBMr4x/mmOHzrARO5BZNQky4WtjfyCHrfXYJPVTKpqwNQco9x97Zq2OQRhnAN13fPX/
oVhn/LgUOabWIfKhPpN/vn9ITAA6fq3kd7dTE9x5l9s0pY2vWdQG8W/l0d3dkOJfDoCGHJxcHVog
/E/V4XzUH0tDsTBwm7GSdwj+j1J9i82OY19wzRnmQYUt2GZQ7ydOm13QEuclNA7NGj8Qah/i30rT
l3313bVSXq+mvj4pL4x7g+2WszMq7boFO/yn1wHvVVQL2HLnZcdLOoBO1pS97W3pertnKjl7Sh1/
2ApDl0oPzC2W+jkLtyGsdh99fEKsJUQC88ZhoiL6bPoHXqU71UlglzWf8/VWzleytWPjZiWnM5be
fld7JVyhwKx5Znm5mFhTowN3NG6vZmmhb3r6QM36VRMueRStjRCfqPfwA57/YN39eKsy0Fux6Rw2
eUsYuewmoKA0UMbo+Y3L6IBDGKYZw3KFksEH5K9YpXF+HFoMHHamqSI7uvjO5Qb7aIprNX0AdFT5
1IsZ7Fma/8lahH+ncf4T07vj3RMmJdWQy0V2DQyV9GpEPRd/RbvQawm/5vgPXiljHfgTykjbIgJj
ExJrU7v1epwF6vpRP9Fv4OOO52/RkD3jzIUx543+UFp7/Mygce43nMKVuY7YePmpDGh85Up71cJB
uJJOqabbuGqlVIc0YPi9cSQYaMZaBGymxG3vCSQvUxehqRDTGtGesTGt7/sZ+q8wbX2SZr7Ng+Q5
d4Dtzzk14y4pg79gKXguxhfb2Pgp48LybxdcJc1adOcWrm0G47/yxiAIjb0eXfTGbPYqMk3svECT
guyh5fI5azTp1X6IpqmLivKUSJu20KqDeI4wF+gJeCBdEt7CBWHCVURuQFCGuHUycQWIweCjvw64
/oEHIABdCAdQwL4d7NNZke9L7y8kjc9HyevfJidghOvASOyoNckGr2RR8XExaT0hyAcHARQSOdeZ
TvneGLBRSlDeGOKNAv4JZ2TOrPmsPYfhOP1n6PatQbj0+EUEWg4DjAmq8yIZz8sP3FPdh69s5C+U
+oeOR41xbw3oCnZY97zQe2OiBzuiosC+fAKQZHKnBDkUcNFuAV0dDTMZFzRXCUdi92ICd1hSMnhb
xoBKkShRMikbzvWh+y6iZ+ULTCLU2ZyZZwGZJy3VSjDHocuRIWUYk5KtS3x+4DH/lra0cE1Oom3L
qpBbmx8MgOpK09OzvZVsnVUTD7EKmvq9WWBjCVJWskZDng6nGZzzrAAxCJo6iJFwuK1reOc1pbzl
vn4u2GKaNoEmfS1jjt3MYmQEvBVGCuCu7Q+XKXf1nMBWKGoBK5WlEyjhRsBg2mZq7OWfcetDKnfc
PTI5hqRtTBU6sbqo/aP3jXa9gh1of5DMBKCwThGolBavxSMzfbJW2clHNiF3PCXNbegBmWivsYPz
AYOFvpYn1DwCFQzlZT0hyFZ+JqRfWYdGEnrdgk3n8dc4+/wyRUBoCn0KmVYlUfSSv25l+rJqpyht
pfRmom1rcWQLudSyBHFsF4bAsQLWzXXxGO1T74xHvLg9qNPfY97fHMTDiyqlX1gIdWiSPh4aMMoQ
Ok3+/5fUQMZy93VRmH2toYVgRg3W+cIE9nIGysGUQfAjc2ux7nUIC0d/qAh09LGcvpuQQpKV5xwG
KYYdB9l8qK+7FvSdaLqantt7cqtqDYDKcvJDcxQtIDKkAK6laojFqKkuxmI+8ewzTnMVrlkK7i0q
+mJnuSRyrl8XnQkIIheq5Ob9vvbpy2rwD8tLpka6dTEQfUJLEJ3B1wekr2vPIscDiysPDyS4OXNA
8aPH3dvOrKXzSF52AkT5BFIcye/RYjZc0EX7FFVinnD/mC97jP7BQfLrtXY9zWNSROPInMVTZUYE
eXYFQCYsv1zBh0aTuqZM2ueWyE1Z+lD9TqRcnWz22XWEdJJdIWjICN6qRQDCjUxAEmH8REccfzEy
C+iG/IulI6Pc8fQecMFmp0Rbx1fxyjT978tQsWmeh1d1NLrPVBNWgBqCmF/9vDb1753hcIml/qGs
vtKeFPpLWlAgcY5twMpScXc3EGV47rd4g7hLkYZ9nHPIQle3j4FQWcq7Ar0MBWbi5MFBUKgmUQiE
p3h3rEeFWorfqqsRElQY9xYr1oovnFqe+t3QG46WbyCRcEjPxIXDitVVZaYfIF8ZuxAiCNgsvW/n
XjqFiiaFYbgQ7RiWUomh16rmyJ6oGnKuEX9V638K6JiJrRmkv2n9TzoFvIgdVqcAXmeqtDzC7dD9
GtWWk1obw7wqc+L5fwkpqNy8rkySzO66NyuqFsIDqWpr+yz+OUDzQvjvuE9/pbVhizyjYTUQUips
OKyWVOOYkQwZanwBBVSSeMAjycgnKZ+nPIVcIvWcXEhpaDWLnUhBgPKIwgTIfwmRxyXE7Zhx48aR
cO632rry7aiBWkLrF7COgc5G6Ou02eWu7LI2Q1n116FToaQtmq02SpWt1wHTITBAuh/xR2GbS516
kJrf5WhJ8H3ln0RxdLBlGV4qZ/JpF3Jc4PVaHw5pQniIWffaZ6DToNpwAmyd8tMhh/YAd3AQ5Aa2
yoUPsyBPpFitlZ6i+tUxJYcxBRm/x7pyPW99qTZKYMDfJ5bXuMA1fK1TnVodoL+5WsH4f6iCuXTn
LVa+VAcfxZyfyQE0EsQYs9IAgjmQ7744ouTYjpIJc9eD4nr6Pkc/ES0244IsnE8cQ1kviKU+AynO
B8L2h8/jnLbFI+DbmVdEF7RdxaF1LqazBeR/RuXVkg9M/mLIlyB2qMS18DQZPdUshPwU7Ob9R856
FuyXnNIA2zlCrlj6ROi0H0KoaVmRmSF189I2972d1MglByGA66AZvqn9ZIYXGq47URxWbw8d6f4+
JXsZb8jVgyqC6z9qQd1asFXCfiOFh+hRAjmkuXmxj/4BC1HDVKnIanPfVUZlakCOAppz9JnXHQbN
lSmVl9WyegMiHY3QClLNroUFZ6M7cB7isW1zXeS4FnM8f/Qt65BmhwSLs5o5M2c8miLqvNEf3KQn
YpSvozIYCA8Znz1wB08/jqiSA9KtAWFype8XaNYOiJ0qyknZ84avW1F4ZyYy5vlJG/p/J3jRjaSv
t3ZeVoUEnjGG22Rcvvdahpt/7zHN9Mo6JaMJqoTWnpzWwIi47CITynPiOEliTfl3l55mUqkpvqDe
oYqDkgCW2Ks5V4+G5Uzrr+AdknWU6wmFjXATFYsP8D0eEtNwehysE0YHc0MnEbgzzgbpYl4cCWOC
xFlOuSZXsVOle5Hf7sc40ETd1oD1I9jfP+GVonizWskPNRm8qH5GcDfzogYOOkhyZXfUrSKX+g3c
66VMYy5vTqxxYHFja8e74mA8rqZ2eyXiqFwyl7Iypz6g/ETFGYhqJAg01mPygDzROrsjL6a6s/T5
1R3YoqIWvhhuyfX71O3kSCOYDzrKwpT73q0ob9iKJzthsWR2Wld3SxvD3a2nBDG67vGVndiySgo9
JlzvwcrHk3qxjVXkQFaIllssSoXF5tCgbvKX+hufvNV2K+bLRlcg4pCpejAM0mkOpEPSfKj5dML4
U2zLO+GKwzH9w6HrR/Limf0lKJ/IbInYU4lrSb/Jj3tFRSpOjoaAryGKhYA3auijxy6crcGdOWcs
THoogOJ8+XHnjg4QFwr6O7tIzq2EE+qCD3VhCywcwUfcAhw83PCPXTP4jVsLnkyIIfl9pSX9ZvxF
9LacExTbBqYU98NDkMhJEi7SlAtSljqiiUhExGGe/N4/ZqMRR5Zjlg0adkcpW1HugfWlsnhaWqv5
KHyUpP6JdN1myi+2XTtiAihK+visQ95tA6y4ZMnDYv/CKJAoAsbiOr1I6sSnbtC+ij4e91xS5u5w
0j2uvI4Ch4MwWONViWHFQ1QLCMLPStT/yCx/14nP/RdTMIiPiAV7swxRxq0LOoZJNw6ZdiSnmZ+U
fkUJWBi9pMv/1YO23dUqU2V22jrUEAmgGq2r8eUyAHYjtAQBhs9WkQANG4p9XQp/EHctTcm3Dnxa
xuBIiiyS2+ZUmLVVnc9AOFcKGbZuV8HlHYJdhMO+JM+eaZi3RJtzsyq+I/R579ylzDkqt3BH2wOg
PiJM9DQxF6F7s/UDqNAKsQzi8GTrxAf19kid5PcPYtn3m0AJY4+tFHRSA9T5wOMiVC/YgKTRuKro
6a1ZeVvFFswHRL81qpC5bnQ2TwfkT9rkhBaouhZte21QaJCYbcarwnVDDABgBkPF2wscD7NQv1rH
iCxmzDGImn0ZLdWXtCms2xgiqzBslzDj+yCyBOcSijtA/UhP26GWkGc5AqsrogcOjJKWrPis15s4
rB16Z1QC8XgJjjJacwA3JM9l+JvO5WOODnybaH1Tlp+/F9y8qniAlPOOqF2I82j7rddq8pVmzcZO
aOUYp02Orn4rLjLW8skbwzgdpTk3K9N8BV2OQmbEz5ny84rgrL+CNvFNNR5ZYjXVwMAHd1IrQigZ
Af5qRvPIBvrpDloj+olDBms7aFfQjToyBcsnGvPPZ3qA+zOjEoBmTzNHu+YV8Ov2duBos0hO3Dfo
NVaD4X7bo1wWEIgIRVp857g5Sype2OmCYcDuaY3vdttJmAS1Z6EBnDNFGAK//sLWzEE+dj4NcTkc
A17eJNltw/axjDlSbEBXHqtke4obgA+iB4Sn+saDGyY5t8YndZYFKA558d2q6X9NmOrCo1G6iL1A
wb43HublC6kZ/+xJj+7BPddh6jOtEHtU20mRy8ALN7AJRW0Bv28SjRrrZJ+G89awYMKYGc9TyERS
xM+roDPa0LMEU5DT5qsaAwVBimkVaaT40WiY6m36r9Qd/hTE9IbaF9aejXy7nUU18R1OOikPZzPF
DTwGt2PFTemRSDOFvzdluWL3BBOFicABI11HIf06x3UJH4gApZhb9ATmSSxCbvkwexkNan6B+Ypu
hRtvKy1/P+zNK+T279XG4BtC7s4VlFkpkhzdscdnOQ4yZ2hywUg9VAbSxX/HG/9Yjag8E6vm5GUb
pqZpSIFiHALeLxI4rapCzfhjFVT+TdhHc87jhqjkvivI9sBbRlA9V5dJvQ/r18xyomlJxbotHl6Y
O5NytJKOgbz+huc6ymf5DWEQlPauwre/2w+KvQOSf3/FQsYkLlCwBKBAtBpK4uoA/MUji3c75DQ3
SfHCF8qF2FlvTjc1EC/Xg4e2cfc+tbWfiqnXMWgCMeOvtefPyQiFkMmk+YeJgKLI4uCzLap3uDbI
ti3PKOXNtC6wpfbhoo6ihZ1twmi4RkZF0JeNMYsMgcurkdaIc6ec2BZxoVX8xhQurVaF77fEnJFd
Jvl4b7qZpQXoirMJpRv/DUE9rST6DwSJiG0I7c0SyQea16ZZxiUnTYVr3IZ2oSfFCOsHTjR9hRId
ATWkBxEYLFOA7M3i3se6SgpLmEdkd3llMgxHlGBWW0fcXzL4C4i24HHdCKoNd0HqkSY7Et4PFicw
JkqWMIvz9g0ikp8WDq+Es1MUPLsEyEzbVK4IhJvbJcpC0p9FeLnpgr3b2QmYIKhZO9uOXyKlLGCE
iERa1Nx6ORdBOLwvV5Hoknu3ldgLxkF/9uZouiTrV+bWgfbRGeY7bHi9L9afafet6yYAm/DGERzC
9BnZ8NUfseTHk7jCygJjPR7boDAXfmUbcVAFUv5Z/9vy28Oq4hTQTXBcLaLxQqJAH9+hYBcAEZr1
gPhO6HiUQ4+kCAyK+0/KdL6tEOjMD75eOet5UG3edN3bFkx7rHJBH93ka5mQWjJyqGdkLmZZ1Zyc
0OpZlxyLYFMho4pv8O6AOzGBhD1B4KrST8Xpg/lsN58wkz3JUX9g0th057jcnAS2BGZGBnkzhl8Y
ZkXZmgT6fbD1zMkG7qWNmGKdOMF9xKg/kgDUziebM2+0tIWrBmtxxCu2AwSey3i8ip2GDjV7WhiA
fXbdn/5p+4zinmCsLcqw3cp3XR2dkTr3JbXOuZjwd9XiJGaC2k0xx3tFLQhq76BfUc6f3jLavYJJ
OYfC0QOGhHL5U2Rjsauwv96yIhI2U/89qxKza+XDc8vR8/0RbaN1noRr+007wV0Ea+xwPj5TivFp
3Gu6mq3nADSfm2LRtTlUvZSxPxHeDQHpCnIOb5/slILj3Ob8gpeA3gLsFPCodjkfPGCQRc7wGgJR
wbMDR8tiG2gvqIt7faOpW1xKbZnBSrYsK3QyECmzdzskrKb+596lJbUzz9cv68H04Zsr6SvJI+nC
+JpznxWQfPTh3O6raFeqY2YqXJvQOU6m9/UeJQURltjc6kPjAFDqXYa5tzJnNZoxOtMxM2IBuW+o
TXQy8jqnwSjjRv4DGk5IoFEJW+UXmTbJfeedseIgaQDb3iEkMQwsb4crdk2mHN6R65nA+EEFoJWh
7G2mbDYhDBQkDsipYf6ohmzoLUbcP6OyfuIqeYp5Pl55IKgoKcRzr+OAL9yv2LC4NvMs4HZu15LK
FDBcpIZYQAX0k1UepmP/dFFgau9lzNw3HfyiAjoEkEaKN+S4avYErYqDK3jsGofxwo3A7S3O4py7
G1wNUvjoNswARFlwV+uyD5EmW05jHCQw2xyF+scv/EFGoEJlnkzhWsOyPAHm+3VFrukj5OsLboyV
Iq09MjWdHxoetlkQ5+3IKAmD6f1XDP2OswFZWNb4KMVI8nnPP8aIfRFDVrX727LdbWnDwtk74qg1
+s6qIU8Afmq/3Ota8dVguYWx//LBGJ1iFNHcIhidRV0eAicfyIYQ0YTD+sqRg5/j+HQs1Lubvyxa
R9WPRxlVKbLUvI0pG1fncViyIN1r19L89SDPNUcXmGH3Mt6gJb1TzPpxyJG0JovqE93LZ3Wox04M
VMj0m1fJvAkioJubgSzmNcOtZz08FQmI+7P6pmmYAyylUnulgC7hF+hFM3T2OF2Ttx9CeAbpUKbM
JtKCCRcw6KXzePofxmAD/DX64j5mMJGK5OHHogWSRqQ72c01vvl+J2Skp47K41t+J57KVw9spPsJ
xGAmFZWajLPOU8dy/BHgiyXQDhzJzcsuNcEYQF0Njg2X/8tWuVkfORK8wcnQosk10uEcC6Ic6/W5
OXf611T5llbMy7mAPtlyIsDgq8kN7RGbT56BskcBMxvBSAKdp68maSghuOnmCSBJkU5o0St9Rk0N
lANOIJwdAjbcwFLZVW0esy4PhKIzeyuIhlI0Wdkmu/rn51QyFW8KjnPQimvzcwpg6VH7p2fVjvx5
YDn2d/KDKoG2rq8EnlojnAGqga0IF3rygXkwpcTtxI3vPPclqyXBEI2Xp+cDoV0cZtvDj3J4S49d
Q9JDGRz2WuamtcNkwzhSPg4sDlFQNHZgOLkP5rmkOyWeLk/Xe2srBRNMmvAFi6oYfpoDLnKaYoGi
YmlQbjZpb/WpNZ5IJ3vyCpOB5kPIPXAMM1un+cO7FVP8lKSX44jFqOi+gXliyUF7JrtW+jA7XtAC
G8YntTYiiWMXntNus1t73UNCH+QDf7s2EBRIyFI8jmmn9RQPiEl6/5VJavCnzwlmVxJYzpXmpUu+
GHJxAN67txa3vrC5048lBoLiMKkSpek6FZq+XMQ+7CX61oDWicYoNGO8AetN5s3CI52D6yctGOYH
ufLyIzvY55ZMpOpE0so5JYItIpxKt5SYkhjdxkdepD9Lh7K6azM6tc3wov5aH4DS+j2sngI4v2lj
iUrLcOCQOHEWJ44kPlIyAGP967/Z6o2TF/GhBImc38/X2oP1ZaimWbcpI9T1hvUKEVAb0KbI+nA5
96TEy8aZm3VeCJwPdEL2TQt9j0picQj0AfqpHOi3gvKJ4j0OctT30968SUv+EIHCEGATtSzKM1P4
yKjwGL3y6bLosz184lYoRS9UcEvwCPOmBqk9kZfDJQV3D3637Ztb7gil3HQXBCp9dJ0UCMZV4rEw
Jssl4mf6Fv/9WZ91r3PQAJwB5eHHl6qOUIKWNLuHcOn44yXDcCZD5/KnGfYZe7ZCux5GWsp4tTQM
ejfMmf8Z/JMB8+rXH87ptFt70Ej3+KaxMYmhTMOqk3UMxzrYYVBPC/LpmPvdY9KrK+KENLPyZuof
5JM4tEhIFw5UwE2EOmSRKdXSUODsU67AgzGx588Z54WaZjGCqRZCpksLoqdPYhKbQtDBvxIOk5iR
Ilss9SSZB3q6FnKWki5Q0iwyCa/Tyhm6lJex29gYz0ViqnN3+ZQp3McS5IuaUeZP60T6YLyAorN+
scoFB73bkm9f8odBhyG2x/UvmtBsys9xzOFKmYph28B9cR37w43TKC6suxapbMyoWFGAqn99ENGT
WgT7xSxoyZQCA8qa1VWsMAvLQqef/+nputtFsuM4Ba0Qu8FmegQyMsKefysMHOBCwBUQkcU9lcWF
2dtHLx/IaOCbAjsXnCBfn9OlRCVXsEXd6lAl3BTYUUjaC8IaHfvgB1cVPfW0Pngl/Trc9RH/BoE0
vkHpJHuYwVF3MN64RvKQ9Q9wnTlt4LJUlDGIm5mCB6hsqV4rHjhoXf+qo9FkPt93KGPoxrlrpyag
m1P5JdU1p8f9kCoJUjo0TcQLMAejOg4YvM41WGwhKnie00VE9M/JKH0JwGO/5mobRpt4wlwpspIp
8JwTjTc9cQGYdAsh/+/1h5aGGyo9Qo1JoWLkYpxXos8VORjKKzBAi9LmjRjE9THamMujavqym+5t
BNeL+JwrbESvZ+Wv5Ga+wdPl+GudSr0n3REa+Y16IMpz94UG59+67xceJDr+0Ht6qEDM3MyJQdx1
ZYFxrGtaceMtXLsYyOrGJbpsI+vMqnH8U7PFkKgdlnS7i40zTSpbrtzpzokqUSqNLlWwNyaqZSrV
0GBMvlHtbYJqUi8iG9zMsE62CSNdDmTd6AN/kucmZMIFEjBVjD9s8TuJY3GWS5GftJuTcbyViF5W
vB/goF3hbYhfajMLD5pRRbj+JmSjBEcAC0BoxFY4Th968atK49iGoAE26UP9OqxMgF5yeVjDApPh
x4kU+h2vVsP4lyF0/lcwqrT9itXQbPaxCUcnXuWs6+M7+Tq9YndVJxEM7Y+8j533D3QAIdGufqyP
8D0XnGQoPzR3F/h3ph92Z9XJJpq7JB5B9gqDpTqmTMx1839+ojA6rviiC23iL7zPn5FSy0U7soGn
cQ/l61NkxNA9uEaRmsBBOVKqB2YJe/VfeCx5DeoyhOniL9SNFcpbQLjijX4zsRQ26Q3k+VkT4nQt
uVVdam9HH1AVmYbKvFWL84hZ4DRz58r5e0kxHtG3yUZnJNrJ6HRKkhP6sozEMNgqvwqLK5+P0EMS
iQn0cCekAANe/5rTpsnY65S2/JgHSY2JE2wQ5nAS6S93u74IX3MZORJhdJz2Tcn/JjtGykfutNOx
TlF/AfbaI4LqqLug9qTGi2audgWTWR9XSOnwiuBoC9NtD/3Q1NmrRzu7gswbWY7H0uIwJgyIXXIU
IPeFmSovnLffJR3IlJ9PDuuz0mpi75JNv3P/T+Q5PIPWn/nF1HG8aI2mbmN9lwNaJ6Ct4dHBDAyR
9o9FyY/Ovvipc1l3OOZj4mHgkLz1IOqQnb5yXP2ltkbUQDsayHX27rnJh3uGgg39KOX9Zz3810+E
wATq+9qhwm5WwPc9z6f3uBXAKXqUx0H93FbGAykmnFstW6YilN6aYZYTx6mjOUiPuoz/aCJH5j8I
EZa3s6mxbckLHnTcxU+UPWE65M6gG/KZHnrBFGlEtsJbiKTDapwASwdDlTLlDAA07TdkGcPCegsl
CvZpJF/ZhiQSRtunxgtkvknLzJXrh+TSuPylll7ESLzyJApGAWxd9r+St6Vx0wpXrROnSnhCtES8
KDwxK52z8EeCp8MFAduyDtOtqZJ7TgK92gJX9VX65k94/WRD8mgbuLXV31eTfGogQKuz/qsiAEFE
WA/XWufnOQBSoEkNav69/OdksyXvfsbIjqF+zQql85EMihUzoe1IW0JABki03Mgrgrcu1x1RuMcJ
IDjuuclwhqxdYF+1vl430b05p2sFAHD5WVLq/QqliMp9VL7JqUiuEQrI8osuxk6ei9NMqTtmiBlv
pTtdp6xMtBmAUTgHEQUbG/UvteEm4vAOSC8I4QD9WJdCoyA/Z0mZjiMS46RtrUgyhZ5BhewgMR6L
sBCDeY6UEiZ/ajOlDwoxS2jfQHH1BbirbLU4P//hQcWie9IwJL7FOTHhwDPX/sAAoIHrYHt9bNn6
r1motelQlx2moAiaBy4kuNd2GDFsKCu4R+RBFpPQVvHovnc85EBuFISsyqjLXIOuzwY+448LhCPi
/f/CN75TVO7/pNK00wwVNFxA6aial+H+8p9zLQJDDhRlcDt2c3oAoI3YMhHF3Ubj/kizo9pNoBW6
XoaQO1zxTMVKbCFJ25WQNkvKgECoDpOHyDEaqGzZPDWybENiWjobE7rjXwf9HMC6pWXzYu9txNlt
jhkLnGlgBU5vQLU5OPe4M43njj80iUF+0l6mImD2LSZ0duRajphZ883WjRuJL4LNgstwHWMbj8fD
mk++FqyoeO6E/CdcsRitWW3131rDrOHdfo5PzPWZw5zgdhvKdg7p6XMj9NbTUJvdhqC22UQktbKi
BfmQDXdqOcS4cB6I/TYceTXREzdyKlRPi9uG0aDXFJeq2Ja594YF7xj4KlHd/jUquAMXmWbC57EO
DDiOsBAaGHss/IDqGJZWWHhuCvE3VhIwS3Kf4IbxDCnMAmahfWChkdwut7yQEOOrCGYuyDIPo3Ke
yZECHlbSWWlyoqa2gSGunPvLx2G7ADCGsi0W8JtBWY8zKx78H0kGgEnspTcS1zaAUItlpdygqvh9
6/+KbrMEnZgd3rEyCzfT9IB0o6hM5qwFhUbefMbwkA3kOyJY2XG3YSn4IW6FUY8CsfhL3pvXT/cg
mxn3eWEx0sQporPKvNcBWwMTrzjm2PaQonVWeqF8I/WfQBWVO53HoctFKsgHiPZ/dCsfVNnl+tU/
E6KynWBAhBf0zokKALutad+uaaBklTc7rkbvSRtAzu9T36FCavb0fYdx/6N2AX3gYc0UcNtsbkwL
BJ3i6VWcsbwqnV03Z9j9QCDdiYOvbYpLdQYIPTWo1n4IbkIPf2QEYz3QohPC1dL/1W2EjzlVZtUv
Z0SOWxCWlEv71G7hJDpbfXAGFNHM89ZuySWCqodYgJaWlxx37MLZlF/nNjJ62ph4lZMCdrP4bTIk
M6STxoPiIS9rlDKXMJXKp7DB/kNfxOFDsqxXAe8XuPnCsColwUY1NWyVsvHpREuZm8PPeR7/NOqd
FbAlRGId/yM7HBx7D3Bg3E2yeLvdQDXGXkawjNv7Plw03urZfls0wR6e9GZlNr3OQxfrUGi89Rae
4L3TbVYIfc+dSWZLe55KWeowsrm7mwu1x0LLSK7NiwnzJfTf4SW+oMjialE1DaXF+gGhO7bQUAQ0
/h2+k2axyUGtUTXgvKQcNg0zGOO+a4bDfzubUt7mu0knFk65a6SAYeODE4Yt2lYZHgjEXnbQaehS
7BzFbUqIk+hWS5k2W5o/TxV6KDnUCNh10obLeKEkm8iJiy4sbicFs7CvfkmKUpMkjeDNFBTkGUMK
fRdLki44uT7PMTUZiQKxjylmHQ9RrSt9Wnqwt6QYSjcjkZ2xpawjz9+e9wPqQ06By6in8JA+IrsC
GsB23SJg0HFIu57p8+7Cuk3yVZbVsmn72mqRqjwrZr1pWgb+Kw+SRbWtlHvdLnADshLNBl+0cO7i
5LU9sq5fodmdlc1EgoM5kc5LF3d6umwuRguDXEvJZgOg360X4ftcoMX4qf35VQ5HD91Tpxj5GdYH
1cBGqhCrn3vrx+eoTFhU3EAVbx2VlY38p8PlT4f4r4sJ4kJg8ZDZlPxbefDndFTLfeLlRGLCW0+l
a2rER/b4GT+8aSxPmeJoiRwWV0iThHbeV91Jb6oX3JHzDqFMgKn+cLuXFclSwcnNCwolSvMQwhHR
xPeTET3nO9uUlfoTHgZKr6ArcCG1tHxqfB1RDDiBsFIKipnJ/sWVcutKXgiMecJTwdxmPFA4+GSg
+DUlHVk9LfpjsuFSQiX2M/SmTlcWJuluq435nYRDcePGwZwyTpz97JwP/wsemgjJeWxC2RxUQihs
L19hqDOsPQd14QzfNzdXleDPLs5yx0Kn6woWOuFF5cgMjc0B/QxXdMewy45eIZ26h2s4uiksFFYa
DAJpMC5oBFAwKVJJxfrSmxA8bPy+5M+5rX/p6k5QOHO/IRJSMKMiHlMdvR9NggGXZccKoyMXrRy0
6kvAFHTbZl2MOSCX6+aeXrxG8XnWPvVrFatp7HhZmOhfo5iD2mkONm1uxVfFzwyAIp1N8Hgf4ytX
tGnfQNqQW1SrdEp3KTgU9oeDTOuY/qjh6CpXmu/uL6FMC3NQGxbQgo/IX22vNg2L3SSAlpv/YrjL
saCBuUV2P+9ZJi0Rq7PIMlqjBaTtDL6yZApBgMnpqrhXQpxyL0MQOO/vopbmYVk7qgabgqcMJZm5
SljI2qrFG9ZHz9NMHcQmyFE6g9b49hkr4rC9NYaBYfQgQCvrACP8DBj/1L1IbIpoOztxDQsYg2ar
FzqYj3HQW2AUE6AzV25Ttbv6BNjs4ZJGMTb5lQp/mMYvoNI2fXLd8WnnDsMIM3voF4mUouiydI27
2rWyRvjTdJe2rgm6s+VYI057riUguLPJ9Afho/SZXLqoalg8hjyHgUbDCpSQkDXtXivV2J4P9wV4
zZGg1S10uj7jdL9F2KalhZTTdcbV4rNA1SsBjan26G+IDL3p7AXNbU9vpt6EartX4ZnspHWsnN6P
yMnprofzBuvfnrEjZBpD4y9ybv6PK0gs5O8nxLzdkLubhhxsPId2f8s+VxHBKCRKxCoFcC2T8e8h
qmcEI8/yeKp2Bll+Uy21qxOHIMi8KvpizEqORKOalg7yMor5osimGHSQi4CRgudWqGpIGRNLEdzx
YyrIf6LtzeuL1GjhZytdTClwaC6q3Js9vfwMwzMB5uxSw0kiEnrYd5eeh5my6tSLVJBo23u5peGN
kiZRUpEHNHE75rkuALGYGly0mkyoDIJF6yx5SCcgCROLfBqz/9Q+eoMeUNUmKSOEqmHfP9LDem5D
+a7gETcVtTMhNNdgWM8xsVfm0Jk9DqE5GGLFgEZGCY9D1QQW9C362vSoDL5h3V1+taWc0zd2QZJD
ZShc96RwfTKhMHkMOugyRdgpYw/51XwuOm0oJLIHx0mAVEdZGcjcefLfn49DdKGHOowjW9dHZCBm
tnkTXJgqGoNvBdB0g1Sxh6Ef/pc9scQfwo7+FfUq3V4U0zwDkXmYEllTyL77W7b33k1FNIdHllvs
gumfI3Ci1+JRCqr2c/aa18OPiTJ/Cakc7Dck03of7yEp0YBPGmbl7SLxZK94K8rOFdVRm8rO3Wgk
+iN0Y47Y7NbCh6FZzE/Iea6JfoIedm5dcGznwSO1GDLkO8aYOW5SNt4Oo6H4ThIRbqds36M5F7ge
J3LIDCPf5rolIXIoD4FCNIragDofRKcgZmlSZy05Q8N9MfL8OEEIYi2bKcivnqrE4pfGXsTNHUMw
aFI35jGrChzRQsQ0uqxYPhR/Y9R21BkjPyzOmWVEfWRgEJCfXzz746kBEvm/VO1VGBQZt3KFq1Uc
jeGJESezqpjCBBMD+lXkELGM5qRe7/AQ1Y5TaPN0WwmuVUJiFylclLBvH+54rftqqlvHrNWQmBaf
qMbIHe7zqlTPU+zVEviemmbcVG3jkep6ansrgP7+VJFVqOukJUT/sbCIzvnMses0ETMCEcqpIJrs
dceQU0BDhJpEZTv68f3hkta+i8Ss8KdQo+/ktnyhRjyAcWac4APwr2fA/bdXPZ4ibWBEBWzrm7AL
lMPGOywCJ+gG4zQ7u4c3CoMt78oOtQWKlF8jRlBgsVpzRWVLnyG3r7MNOtx6b8RPU+cR1wKSrDPd
H8C3ZK4TosYlKGbjungyT/nqJyT75fsPsfnd8limlsXSPjpAQHf9DeccNiwLarw31JCZWyEdiC/K
6B3MQk9ib5wHJ8gZg8/DnjTaw8ssS4F394XIn/FePo/g8tzGl7WB4MOr9M/ABDfyEWiHbHlcmkO0
33zG9eY1NOl4TojuQK2xpeNxSzHvG5z9Gql+VRV4ISl+LSFlYLktIA3etjL0/lVZbI+7y9VmJ50H
k1F4+0tKYHIWtcpo2MZcG/emRibi7UHi6v5TMf3vO7Eo3qtrDRtvuMyIPsHrNX5g6APR1pKh8vpF
zTENoRxhcJeIrWFATOEgjJSCRvNZzBJ2BZ0Zdg3itBWgCQGUhnNjKwyrubsiaoQdVLxH2L7CJU2l
7VQYBeWJJ+P8mRWd88lEUnF6U6csw3djW4uT5ZeuSziIlnw/tJWHuho1lSz6D3iKaR7Oyr3wXTEJ
VHZmPir54+QZfbcRyXYbz8MKEZ3HyFzT7Qd7D4r7LuQw4oI+H5ecsxUQWWhaSWPLniTnVvKvIF/J
hhbg06rhe03TQa8dF4wL1iApObyjqgZf9reHahhu9MucLfIcCx/nSa2cKbatAJ9FFibkgWrT4d81
EaiCcS5+kHGZQVu383/I1rU4FhcIEnbb0zzJXKHt2iKuITeS9xk1kX/2CNjbqadXg/3kKywktN1w
yrJ8oS9w+HpOldw5yugtmfw16Oqzgrv9SIsRdn3bxxUdxL6URtmF4XO1mj/S/cf54bP7hGkNpcXB
gm3ZqLkcyZGEFZgBbRiGy/rFN3hbJAGRnKI3o8dKP/03XHnKS/7Xex+SpHUpqJy4zBcHe2gNsXo2
uM/uFxRgSt6Rrgs15SRU/1LdTNtHCduAQlkQgY9ELHKszDoiGPGvpuilCo7QvggVASte0Jv5PbJ1
hkTFug2d+hnegU/OL74dKgsE6H2x+MVMk1LD7iKpwHVN1rvvqY+J+lsOvqgwV7IB+h4nZQ+6drG+
qXBI35xKlb75HALSrppMxfnvLK4oHvQ1Q+GVZk5jqVK84yraQ10Bhk6CfZJlGOI/0yrmc6Ag51bM
EZXU8/MtYTZkdW4LQarVAbUJ5Za38PMqtnCFALG1BbWkTD7wnoCtblEgj/WRT2HQeZK5qyIEJO4s
2la3H1IboMvECRpQbbiQiklZ1OQBdiZ6DWVBbfQ94KX4+Ggh+whLN6h5NtbHboddTve8emS5dbrp
1oGDA5/Lrhnnyxi6RnLB1ZW9/f8XMcG3ZqZhzK/pp2pSGi2frKZWKsSemwOX+1q1n8uoPDUc4NUG
gW4PLgKWNgUiwwT/okrnvz9RfGxzhUqxGnjQb4SjcMQkBLyaK56X+lCNDw/ge3DuFjaynSTS4lx/
W9WK0IQVgl+/PpfWYSQ5U/fzHdC3ehn+NdZakPlGVilfo2foZsg9GbkqnhHel6t5NXnpaXOviicx
YqMQJwOO6Kakismx9gP3z4iADfb7mUGp7vrVYVS7H2Y+UDe7TMBmHV7byt5JI03gZVpJK3c44HBU
eH+6rk4G1jR8PnuFJCnOjvjyj1+KQKWMWU734hWe4rNRFnBNJjLVvpmUVlINzZUzyqwUOSn+9ZiN
JCDEDDtyXkbrcIsOwJB/R6G13MomuVJ7idsmYpiStt1yb0wB9Ea7tcXh1sSzmnknlmwjM47jnS5f
73vv2kFXMIvFT/jfY4qifuDDxjMYirnw4iEoVFCA/cYajGADtY69aPEh3iJ+/VI5/d3lAlAv27rZ
5WyaEVB1yd8xQUXpK5H/gFwGV9BWYBtxT3RVxwzQjIdUMbFLrIiCoYimKMRdIw+sZNSbh3ikLvtB
zKyWRgqhnNF33BMDQG97nm+b+ukFtA+Zoh9Hkl1Bx3Btx0+OiQ/+VJsRxLvsO1j77g833PqTkj0F
oVxpz6GTe2lGHgjUEZPeZjAoBpw/LzkPvUaBptnlZbzrncSuntktFXwV0H7gyeny3BQC1/7i8HMa
QaLNPQNSoJBb4fE18lkGURUQW64FYgPFZs3HeKOTmC15Yi+nDaTzb8zcDCvaJMT+nREJsKUI4uvP
gltCkvBWXklgOALbIbFSNW7raEDQIwYYkWfvPxnOvMT9jSBx4BZbwf7gVLRF4MTLZmpb9WVHN9sy
fNJX3vvwgDgD+yttw7axcKlANRcb5Ut0ruknrwXyhbi11DMaI9/vbhVou5bEdbvCs01aiyJrhf9O
x3nfZypQX3GUd7dEKWh8I8NB4r8sS2Ftn8AyPd1YDkEPNNWY/yLb6ClvVp3ofXPOUwtHFdKi9vyA
3U0M5651bkLdmNB/OEKMSrZZLluyoakH4V/M56binQSgATO9BFk9TW3OKnU9Ba3kq/DwE1NKTGKp
QlpKlM2F/j68xrzQmjOtp0fnpaKHpDOheKNPn6jokLk0RTU2Fqnuw7EHSV4kLJnm7tEKQAcmV/zC
9G8JcGbnqTRoFkzi92UF78GmzdrwKxtEBLkjAGvOaxZuivATYMLWT136iXgqI595OkkxwbyfGTYz
P8Wpc5yWA3c8XZTxDBguYt2Iv4dLwfCmLoFEKoGY1TFFHJp6MhDVTLMxHmlN/dhEfM2uSw9KtwT5
W3wk3EpMzN4ib8zuJ+gSuBnaXKaTdxXTYi5KkqhQ0Kheuoun7If6eNIOYGO2MAuHFyqrsRTl8kOD
Cpg1/ybIHsOUFY9B6PnFwpH/H6u9J1+Ew8X3K+ks3vOe26jZVic1caotJhqNNv6DbMrn7FzRXMuz
Rf3rk0i31+2sOmErUjoWzuDPocPyj8utI8U/FhaGHg9u/KwFEOVDVLHN+/7S5j9XuLS4k+jdk75m
1PAE1B45d3aA3/fEZ+bjnvNNmDELh3Kv1VImOVEl8+g1mU2lkBK7sMWA/pnhqvr3PxjxtNqpOnWH
LAf7nBKFaVE/xJMrhyUSUmnAtsBMrQv+pykWlqY2BZLO5VU2WzDp3K0u9Lp849UNhsKPRTfE+geq
YFebfxNZCrQC5g6W3yOSuEjf9Oy+VU0kjpi6OP9PMe22SzTLimLA2IUSMVl+XEGuHQKzzTmI1KcH
E3GKhxv7t+Uh36Bxm04lFg5+pX+QfAaDIz3/2VCeEFVwiE7xdDTNJQJP5h0nY/cSE1ppP6WXADyN
uBRjENNqvuftTpFGgfAD+tygNQEX0QU2BTFGR3Fn0LHvEskoiWX1N2MXtsl9gUZATu+iXlsdWpgy
3fvoJXA9068DpO3k2ySmrpiy6Zpzz+0k/e6N6JXeTB1a1LX6kuFQ/lzKfDRJDTRl0E0vnHEEUQaT
vGyxAsQ5mrX3gNGxA62Lm3xU4RwE6Sblqk57e9QG5yUt7/qKGTUPjN3AfzZyZ94GPsAKHtSsuXyD
FeB7hR3y2vWFYY2q8VjbyuoVDMQYhpybg9R6tzLvTKucWmHV0jOF+6OfaXv8l9ccwUwH+4VRtP6d
u5NkYeQa9DH7fNgEqvJnGL8yeb90xAwQm00FKVpOUZ49aScmKJC9po4myx2HjHThq5sH6H+Km1O7
5FLBL4hES+tjLfYAMPyKAg1NsHkkshUuMLZH2iVjeox7jv8quZo4Hv001AFDBFmJ9jLQiZQcWvYs
bog3/wKxa6knc14bmXOr9vgKU79TZSBTy386SNx/J/YG01xI2MI2Ymh1Muxi/hZebCV7n+KTH2Zy
lUw/p7QXRhrgdVzBuadCsetuhcpe5eSb3QDSvZ1+b5iwHOGQrVAqdzQ87gYJbMkKBsRtM+NNkIYY
Mo9mSujZA9wHxO0kfbkVTqe/VyixFf703FfV1+LdW+UCcuOdZTnCUkjScAGWLZRLW+/wsp+ycrO3
nIAEYjgC0h6p7wKCKTMQSL5HANDP/Oye8cFjUP+AiMcjN6a591sGiqDMo/NDu8zzBLO1BKH7AWlB
qdG8XJKma8lD3RBLXevh58YUy+mw7cjBUbZIK/p06r4buq/8lyRCt/DJPNcSK40QXI+Jc4+VZD2T
FNDlQ9iZaZ17YvYNPRsI+hJn1jElpt3Y8O+py9q263yQu6yMStDJ8u2Pkn6udhDGCGm4dU3rTe4/
Qnp3eQktiPa6IBSsI1Xzlwlto/sCUyASd0mP+FoDskd7Xo2rCteNRakrlSHfkigV9m3EXKZDzCah
o7L6gbSWLyB56MewJMq8wbRAvBOW8bchQnFVzw5rjW0OJXfvUWGaiYwOGNVgU8L1r9vaYchIYPiz
ZOvQSGGRL6RiKuXsSxJWq6vWlG9zfMoPDlEZNd7hCL/0P8ellNYuROwvRdgEN954IgAWySxwMbbU
EMsHSS5eImdO1EScOikPfS9Vx+Q9qVFVSoiYig1zb4NPvCwD3yP8TxlBg28u/dVwIaLRuLy2YZyA
c8gfrUHDm3pBha9Uw+2xykbMvQAbjv0PQ/d7n5bG2fwEzLMBVzGCwhP+Pcxgr8GIpAb8S7Pccohj
jlISbrUPWmsHL5MGf6Gs0+CpVgQ6+7npyVoF5a5WpCqBrt3/1GmF1/XhY2Bop/EX/43AsnGjGZ1Q
iLocebbv7hLj02fq4MqsUR3p5KUlnMROisRCU/kAYyR2P5JGkyJETDsmTmNpPvLlS4nwx+1/J5Cy
TdI7mJ8P4L3KYZB1ZabnEEtE+bk6xcpsoLnrexgtWicGZgzdTDE2pT8ps51NM7KYaVgczsr+2aAB
7jjlryhqst9StJebzKSO2kIxYqupWJRNsFb/Fed3k346YtYMj+dZQvTA5rjN4GwG8//m7SuyyPNq
A3S7KtVCnHp/DObgelkSUemUGfTtBZSxXpVNbwanPZBvbBwmV+zOA90LFhYJnXoGHDbx0VV1QuXG
iQ2kFpORGC3ArZDdRAad83usilP2CI7Lr4blyex6cCWetKi+PLPh3uzGFV30sNIHNuJkA1FsXcbq
5sOQBXS2VO+SRAJfqq6pGliwFHEimzZCTCvjNUomy68ezYniLhcGo+9CiFTPhuJRMPE1/cJHELEA
lhF2tAeYjCgEsqb+p3wo1f53HRbU+H59s6qmdLVrYW9tBgJBbvobHfF+Epn5AmxdIn0koHVUVXOp
BAafxk2pgDSeCTVVCgU85nopN2ZmepLvlqDbPjqMIvXqShXZ+0p94eVMmq5zY+xftTHvjXKkF1B3
nPRQIqD58TH4GZGX9w93X9h6behuu6e/Y2mGSuAduoWeMRtXlBXq6IOIxJtXbXWOoESJ1urbS64s
yGIi1F3zfS3FaSfYST1ygOVt0O8uSJ/q/egNQvXR/ycoBIheB2C91/8wax+JvzSNz9Y1PzZfBHop
HgrTxDyPdGSIptRHcDOri6GEqt9+906x0Xn8BjMiXu4J55Jyd/ENWPofhYqIAgeZ6Yae3Vc9qJgB
sDGj91WyJiUekWBRzTY8Zu8UDe0bSJRWa3MckQow2oBNQRUtpxZaN/oK2PURhF2miYoq7U8TYQiY
wLklyLhft9kb/ez3YtT/+epvmY03Yq+4lLG7ov27aS7EdKcLHyTKWoiQosVNCe/KUzCck9uB60Yj
Tph7igC5c4BFk0Uc1hT562vw1e4GVPVZcJTc8U/Y+wRmytqz+6M+lyL465UtXbkl1Blxuxwkds1f
obBC52ptpM3Pd3nMHIywo3neqkFmkLH7+D/jbhK7lL5QQImj7Ok27rsYFn0RrLlhIT7CU3547/BS
JEoLtWtfMZ5xve3E2pZV4Rw3csOzIWXznmukE47i/j/HFUPxa2SO4t1oobpKTyBzBBUBlje90JIB
0uMDPExPMiIx+TfN4D1js+/1n490RzmCLOVZ0Q2R13atdF0NzHPsaJmX4gDn9eu98tuQm7HUbrx7
qO9/paOp29LVGEYCT3LQA0gg8isuFTVEq7xrZYX7vSLc6vndBcYcLoufPCM7QSxqST7lw6a72DmM
XTFSKsALaGZmIqGui/tNDaGw93UxD2QGpfEMweIa8Esl6W3sIRgsSfBF891wBBzctkA1tyXayGZb
W5S4YyzBCZvsPmnDknUEx6W9Igp7/hsy21deqqsJ6E2T5i+C6qh42x4jlqno47M2gDVXxjSMFWkG
PgX+GpwcUfnjiV47uzwZXh0D21V3973WF3DKO1FO40iU0NlwpJywr/kQEB2GEF+6TZousy9ggvsB
GweTU5E+hU8ZJu56Hd8tdu0i+PVkoUTzbLXFjc8nwW3hwLJ7Q+ktg04S6prHtABZFe/MQqIhOJHR
4IPo7TBhSEOGqHEOSnmneC60VlpQq6T/aWlh4Wo5tD68UzAs9fPSyZK+P/eYKAxenu4fLBuPXO7n
r32S360EOirC5kFrAPoQNmWjiyUBehLNxT7VrCAcLB3YkC03S6zHF6x3qhK2sTzU9WfaH7XHcMIa
RXCGfyx9gHGhFZommat+CfGoXceGHTsuneiVJgwOqAagbzL727wE6yrUXoG2f6Q14pqJSNq/lA5t
umguLbiTO1wEcVcdiQLTcNEQmPJuJ71TzRBmOzFFYq0DS5IQtCr/nGs4JSQqVIYAGrECCL6N9ZaG
2VbzsogJNWfIlxc5nxWZwoKg1qw8D/58WuevTbmDm+U62H6sSJqtBX1s5TenXVYY+H1NwT+x9fjG
vIDZbuzcB3ervwN3QZE5lvrx2XtIqT6N2T9yRl7fFpEATODvcbR9cG/zdy2VssWRKkVF6Fjkr6Ft
TT7sBO5Tt1ElLfFLOxe7pSJ5TGF5LQNqMjZUzY4eCbeOvzaA9w9M55+sUrrrBjD3F+DBfMbkaibS
s9ane01O0IZzHnRJLYZdLVeNqFOa6nWlJooy1K6dqgAvqVM3F1UZ+kA4ei40VHkoKS4bdrapB1F3
pKZ5sr/TKunrzjHBy+wBs82F2DDOQLNSsAEVDiq+rPPWLElEi2/baTiPi2tBEr1d+mEkdBED2nMZ
1Dg10JAWvMsarc9IoQUf+XJ4X/zvcWp2owZTnRBplPQ6VCqB8YQP5FQhh2leOlpllgBG0nktr7V+
eAPigXIHGigH/ZKsgRH76plX9u+wos7lgNlfTE10TuYP/jfWDTPfjwYixuNm3VtnGM567ZjJHUd+
KXJnpGh2B29k+BsQunz3s/ayoPYUPX0tcF408PTrpKrGna0kd7PNyEJvGUk96RhDjHpt1ecZsdsy
y5FVKGBLBWvNJVSEy0ci92k03gt7NLN+h2FBuVDqiUDs2yAr/3KVVC5Wqi5sTNfW8Z3tCfwy+PK0
8tniHMXkmbj7HXxUAGznBcqBBve5BNyMrBTc2DJteMK9pGyqMEOSIh1wdSypks63duQ6xj6hC6RD
8arws2klG21IG5BIK8u9Sqgt2fvkcp7MZALr6j5u450OBa6ZrNYeKot1iZ2RMz1QEKJJ4CELWTVZ
hGRFUKtNnsYnGqyZpv1IK3Dpz239XHq+Hx3Ekm37wRa3cNyF/BHy78n9uUqsIorKI6PWGFG6pors
UMqwWTc5iID2GvYBm283P/Tl7txvz8swaampF2yHNx0dmudyLN/olcJ2L8u6CaboEFLHDuiaE7J2
fsOQoRvSnG7ofwTOFHyp6aRwYTAiMrHxbZ9rQL5oWWEH5sJPdRQlilG2fHfdLztfCDIGbx3Si3M4
ybG6gkAEKuWx8Ahu0+1JVl7cctYMP88Fc49MtssyZzCuHTU6YrvoJEonKA71EoP3xiK1WMwlY5Et
Kx5CJck2qm00StLqWPJig6iEI9OT4gGxxPi1ydbfNTm/Y9ey52L0HOItx60JAT3r/MKlANe5zIpD
nppjPOk/GyPFN9/6PImNty2SGwyb1Azxa99LGUpLqytDspFRlXJnKuyXaa4leT8loqOYmese7PBC
rgde7sYL1K/hm6lL4N5ZU+0kipb7VAj9/pPT+EX3+FwhxvQxssvfhaUu1izweyqnr40MpVNisJou
LISy+qk6Gv8PvnDu965ndeBxd1j7U25AIxmXEfobDll9UDnXs+hGYSbKw7V6g1ey6pS3orHhb1t5
xy6IA2RKk4FLUFS6pV5l0VaR4vLjU3lUq3WRXArW9ga2pr0g2XryJ82a8ub3Ngz2P3aLlXsGOUuV
0ZC1dsgPQ5kPh9RQqGztAYFDkk7xv3+x5XZV4mwmT6jFv0/6ULrxCEMOs1LfE9Aa6/RzVkSZFrVA
rqYAPMXEoBvm1su8ejqODOWbgFyjy655ajKWSGuWWer+sUCgG+27HjtlYLqyYPPfQH1E06GYkVJc
G8/qrS99RDSwQGm9OlEyfTYRPdXqh/2LWN/HmkAtfsrk7KGTw/Gc2F0ubd3RdNueXZ14XdERudVe
87jkidRMevXm9ng9fLrMSr8dCRH4PPVf785oy49E1I5MQnAEr8xdHx+5n+ufOcmyITXglfSyqXb8
0CHENnNtqe+a7PNoDCxfvo144u/s2neWNixYeu1IAEvAexnXPnw0Tb+yvNLH1PIvDgtwpgmR2Yx2
eXRgqakdfSSKoEQ3N8PeHUxtXXSVnbpYco8KEMm3zfg8wlTISzIRgMiciBltH9Tlj+pUfUqM4EW1
cfnt4J6QG+UHduomZZIoEdvDatU/a8S2US7EPNqXwUJfjjaxWm4uhL5/IDtW45l2J4msaCTwVcXF
aBHcZ+SAweFjKeBooVeBOrKR4UvFYZzhj6GVYKgshzWs6HL1lABMYywK3EXupfMlQ+weW2OmBHwR
INjvviP57eBjfgc+fXim6i2mJ0T0lMU9pqeiOPur0b/PsIq+Empo3wXbop3QXjN/fhesDKsfDmxB
fsmW5h4XgKn5Vem9Tptc3GU9Okt0xSoyX2dy2luIwuafcB7j9iTJ3R4+Z2sT7B841yD+Zb29o2vg
c+FGdlXpEfVK8wcuBdVqCkjPdjAVraqlWYwF9LqEyVotAQa/43n4IuNX+V9q7EO5DLZdTChtw+V0
XbPHoxJOjVnQr1Byw+w2oY+XqgQlVOSp3d8xeqDcUsVQhcsd9oGbPg2U3a5NUbRnNEzWwU2dwoiE
AORjevvf4ucxoMxcuZZoiP+KQbujVbFJogPEJjFXhyrEF2k8XPrEthPyy+l9Pbagw5nJoozWzm2+
+LMfVNj23yvE9bf+LXvwTOc1oB12EwFRVCImJdC4Rt8YKXa9wUi4OCSf8aRx/Aq77m7rDzuEam/o
RWLTF148nQ590E63GV9d3Lt8WnD3SinvQtW7rykYzfuoHG7gIQpA+wtXY55z4cIoLz6V0q62ySGq
jHmT7uyBm3uuYI14N5A8E7f0o1DFs7b8IS2LygEVBVFds5acUDhpCn0sWJ8EXt8o7iRr3VNm7dZd
EITWDazLcX74RATnx2Q5+s9MCDXKwlZufiX8cZteX4zVVuBVdLV01B7AmRaGYPAjVyw4GUQ/72MD
4qVV5RmYZlHT7cn42qrF2QBFDlOpn0g0q2ngXPKush7Am0Jf9PvIx9KfZHUED+lkO8qUr/H/A30c
jMHyqMwh9OrQ8WLh2N1Jyq4P/TBX18T7uxctG0jo8SzD7nBJeaGweMNawznMRkgNE1x1n8asI9mc
aHpkC09o9i6bhm7/soNp50HOVm/ZreeNjvEQIiPf6dQUC94gEG5hgAQ9dvPk62uSxODfmF+rWJht
BmibyGZm5kLXQPfskfEeHQaZ8aeANLrrdfAeYX7TBg852Ke8WQ13r9/N+SMikFlqpQ6D5hzdpNVn
dAwHk5OD9mGEKXL1gNe2MF2asChAwu6lrma18xdZhPzPjZcKY96ngJwJPy+G5fp1WQR0MyFWkUoe
djWXZeGJbx7LcxwzscBQV7a+BYm56jGRe5Zf02qLkwMw5e6GsGcCnQwpCoyJIRSLRoaD4wP1xuOR
s0aNDw0Pw9C2FTtd+77QRAnYDw8YWHd1TW5xQng8y9T0p7zGWmCR+Wc4fAVLaVE9ImipaACb36Gz
ta12ft6LiTsaOT1OgD4Ylyi1sL4HKezSnWRS3ei82k1y3seccVgoGHQhc1TaydwDyoN4KohVFxCh
zwFJdDRwjehpCVxeBJeLkz1fp7EkvlbylOy8BehQAjATRQkKeFin+4Q+lAs0ADw1vS5oAC+WPfhF
n15BEgVAkv6YmEHuoQiZQMqaOJO5+i3o0fMKCNRNLLFkULPOeFScUh27glbBGdjMGXs4Az1qjs5Y
Y7MfyiM7+G1+GG9bzVq0s4OHtPlMrcW73XL3EQfvl8lw57JTRCHTBI0YAazc8DIgVy/R1mHv1rMi
abD8cywfqE//IClknkQjIwZ/3uT5HY5fZ109cVgC6kW1W41zVpM4mS3U2CUMXI6hDqQeCdxMYeyn
q9rNwSdcTDk+q2r57kD9nrZ2Qv1SMUrOEWG5Ha4ahpVopHCf39obXOWQMk8yV2rhkNTF6/oNliMv
SFkweyRW8UiDLxVDyxzWK3bDbW+CGmfjGOAjdhP7kKfpSTH+yxFFiu1StcGKQ0ietDKLlirkZAw3
Z2IUzlN327QfGk8vOZc9efIZEy3btRxGZCbD+emWcXKL8flkO3HopYnRUD9MOj1FUqMpgCG9yBN3
LYa+A1JL3r1vjwOyZKCAgTByCmW03XPiyWbsuk6HaZJ0C1FOseUy3hyL4AQ3SxdP8yHN1Y0A0D9z
h+LHk9YnM9fKI15HZ4Os1nHxRHm2v76+v60Jo1sU5Dz3nakrnQGbipiVLr0s9KWr0/a/vxoNbcAt
qx968GLZ1scMD90a03lOMUyEJa2od/S+JqY+7e/aEDmJE0VJIOqD+K7Kx0VyGPazhIbXtB7gkeKh
wB+8/PVP0oersRRl4xEj/nQz6pLjislNiPnGLr1Qn3O0G7u8y/ADCELUXDyBIA/YU8Hv1sG0YfFe
z8nUKbPmbw6weKrVBycpyQ8VS+5cQzsKC3hkfMJt0L1ScNXvKJeVTgXJFsXkP9rBCFt5EZbJAABa
T59yd7ibUJur09ryZecUjQQ2NwNrssdj1o2cpymiiYs9if4lg/JtYBeW+TvZjx75aQWINnenhKsk
4+94w7RFHFETXfrsDqTsd3FhLYycNCeVaO9qTEkzWCF9DBAYFJPBz6mu9TlNqQbAXiJQD7/V17tp
1n4V9aE9KNm9bjML3z7Ud/yGsgfe8ilZrZT4L95y9lISbE6YD/HqISEiL7yUMSDP0rXw1T2ww0An
skXhEwyIRcUQsEz7h3I1kHjJzlPdJb+DJsig/fGt2vTygZHtyOjaB3Ml7RSce0A9jpY7urnMVGJa
/Z+F9cKyosRsV/Z7UWww4aZ1/gQNQBdCRDnn9Am/3idhm2OLmCDaQc01ER8P7IpolWw2U9HjucQe
xSf3xlNaT/WyTIodCAN5dHlQ6mWnCx9+9OIq3Nsecq4LkRtNkD6yNYouDKI9UXzyyDVgpCqkbadn
0tmRZ5Jp7+ndYonBDq9h4eDWsOMQnv6oRCxAkBZhk5lsuNNG5OcCtl/tkZWFvKvqOzjnwWqnN/Wb
T7bOhNqbj5WLZcMedtdGb+A3U9WNOkMroNXO8wPfTtdB2I56Wz8aEgsEpcBqlo0Ej7/oRW1RjoE0
YI2phBr5PuifPLlsZJL0bfxgelJMCVejvAGvCSx/cKsk3Acq3dxLFJQcVihYCl0MryIZE+bxK1wE
tZrneQ2TtTR6AqB261xAsG++FNtyh33vshZ7790kMHKhch3s0+T2/dgv2512P7SlGRDgFoYUgGF/
w/Df3QfNTnsjeCKbVFa7rFTTEcmRjgGiyUvEFi6/sGEJeE3PrF5YMnbpHrLnIwExWZQaRgN4+QG0
LmttnF/AjBuqbZXGZ2bpePg6pgL3KwvgKGa1QN5oK8xV833ScwUYpkLjG/cYMq967mApjFmpAii+
CAZJtsSSc1ILu8gY0+YNu+BYOklO3c3KX50nv5vNaAA7hYXDFrLL7KVhiFispb8qIn4RG6wcr5Xe
EGh6sCxlqrCEJSs1m54qXGxvqFeCNciaqtnTbfhJLAuO4yhchj2v7c/HHPeFluJfvyLdu5n1yIT8
TVW/uGh7UwxJb0IuTwkW+Ml+hHTJCKu1s2Pw407JEzexLBd0se8rrpdMYawMK0Hzsr735iciFcEi
vyT2hYmUXMpPUMr5WrsTcY12S1DboxEoBIjIjWtL0JM9GrgPca/PA/+JWpgZ3XF/kgsXLIP+WHCF
ciQJjpHhmVRd52LhvmmlCCODoDxlez24iWnboLHoIxrkUewvrV+OlWuyS1TkUIGc84wYw7ifmXPB
8s5mJWg5IhRBg5IB552EnpLGf1eysDfSw9T/+7phhfweWmfP9/1F37cf+fP5lUfJduFoXeP2vKxg
z7Mi3q9JjFCQZlbNjZjx5Vdpi0WKFDVC/tALjoHjACzrsDbHxg5np/2oxxc0C7Qz4PRGLifPHmks
Pj4/XjCm/mlz+W8oZEk47KRCBEvyXB899ayYm736Uj/7rX8Q429nwzvZwj/iXVGFi+jXIk5myqLA
ZtDlPX3KQ24CPxIZbtAabtv7Z8U1QbgLsNSfHH5CR1HXd8Hl4L5dYVrbFB3g6PZV+cYtSHNDszTA
MbA892OOOda7aPv8Noahn3cep9kWjvCC8zWHlQORpDkPpdyCG3OSfnLNv+D9bkYS0v5GQrsgNwi1
IrNSWMqKOWDOtXlWQhxMtaeSo6LEmvFNebjUj2PpdGf8Ox70LqKxOAV29pKFMw/y/gQk6FqGowml
czUBo3bvB18nRQHv257lBQzfa6/BhzLkge3QCIXJaifX/TOfyTNjdVlu1Q6Vc/cLxObTVluCtyEd
+GoBQa/XtTdSh4j4214Bz7NFAIA2Ibm56tAQI0KED/7mzM1a6oE7EN/xg/CFFT+jMTPzzUenXxDZ
TkbTeR0RQI+IfI4oGJxkIBiMm57/il0rJWoo2/qNazGkGRE4g3Cm+zpAECn8Hi3bkgUgXp4sb19J
qnn0fmck1YwV/XORdRQERE0Rn9TBATFoa0FXFkSMhXYHYiTKCQJfyhcGJdaXaLMB7uypo+A5NX7I
cGLsCFjs/zwb2cB7h+luKtTAK23rmfJ+qukqh1XhMHxoH6d7UnWp+axTyE8UoTZpf3OADRblICIp
m7HXHQXvXWaDENiJ7iww9HnTgJjDRys1Kh09Bh9L7IauEQ35KeCgQLeao7NImgdPlhzV9HHj+kVq
P7x69226weJHt6oYrdBRndbFOTDORG/s/EGPfcI3D8Ze2t6RV7nAs0L63iGW2WQ4lID+iva7va8Q
P37A00ivXCe5iA24fNBVRjAZVNm0Wcq+I7NwjCDOmtkkj6fvJs9cO67hPGol72cJWk5oHaHQvb3w
C1hpdY3Y3XSk8ltDB5/N3AKz1OFFXRsmBG7gUMQbW3QCiGVaWydas79xOjLKKk4/eqJIrAifzoXk
GVDdfN29xhJkSTzOTdQT+8mzqSfdC8I6Zg4XXI20vlU7SMHQlmWFphNjlipwuXd97icdtvR3BIQy
vjo2Q1xkYrQrgDrPw8Na3A9GO7UQTh9xBVR9d0hwAJUvlPiEZQN7eJlqN23TTWIMyRMGCJr1sB1e
XyeZ93RKvmsgdcTUqM2rF0SCzqXqe+6ZGqzZvcU+Vcr8b3BEXg/LaKpaWcSWWUrCM7VCnLrOEC3z
j4EDQhzLR7lv/Jjkt4bPR79OFuKfOUZ/3RHadO1zuD9s4UMqZjpDRS7xYME9O+/qGuRwYXsS/ML4
0ukUQ/9sRNyj77jpyUJjYGCbplYl4nYz3V2lgrMZdXb8yVwnYbbgoJnlgd2oqEsuJ625QT4bwL1J
caDzz3G5YBozGnDxqodEHrJ499sJm4Ol3RiIlBKAf7hTb7Z8jWkH9OF5k2C6ut3+K/HuCoZ0EqYZ
4iLOdHhIG6/Rm+lC9wx+bZAsTmLcXaPew/dQzAslA1dCJKzd1VfHzF1HKmKVpEz/JCXrH2PKCBkW
MwYZiPqqCNQ7F/LiLYNDFxG9y+euekmKb8bwUJKLYsoNS+4QBBxOib9rIHEaRHg+QRejTYxuLKbh
8P/mfdzM42c4YYUIny6thHYi0MWjN/iEnERm7G1MlN0eTV2EdosRMLLAqWEhclp8uUgoiDhCM073
wTL28b268PTkaaTqCH7VdXvOpePC/INmWDO8csMqqvyVjrP8YarA5Fa++QDjBY5JcojflLKonOXw
LaHfxpRL9194x4HYg3j6oNKjQ0U8sDzO3w2jS/ycEJCKh8JaDKymVVKYG6lHAECHoWH1U8IwIHjq
mJw+IcJ39ORzaQM8ruAwvX1xgZCZ+qkKF9QAH/0upZdHzrkW1qncC/rQFc5Yoznm+Gs+lHHTVSPr
fO3MVwdiKjRhCrSbSc2nWNX1E935JrMoSpRPjs3lhCDkGi1sNDqSxggZuvz6qzLp/879MlVeCIas
LC09Dfb4rSq5C2Oi3b1zeYvcq+ej59xQPtVZVoo7ovqCkGGLsL8QAa3iY9X9Ity/PR4Exu+x0fMv
5zQAK48DaDA3kYUuCjtGynXa83ZT+tFUpVMM/a34Mg9txTbGbfACPxVqZmOZ0Q56bTQR8TxwJBaN
Vj+NoxRcwrhfeWqnvCywsV8f4XZjaa+GPdtNZ9XLPS+90NKQunn7q5jZnkVrPb6TgXLUcUdbqLHr
ENtTnqnGEBaxpbLMoiAodPDT2ExfDWUbQVUm/NbiHW7J32E4yvLCzNT5ZNlz+pBPyIE9QnJnzMm/
WAJDYlXI8sXlu0qXCsxZxiXZYNzclAEJidPgrOeypDZ11RGNP6We57nHcZLeQBCwShLsWQl3hoaP
MgfI8ECFCifyoWZ/lqP13x8KLTHmpEgWuJaM9hHRdSXvrbnom4ZVxWZqlMYF+bw8xmWuW58u39Dd
eyoaAaQB86WCtCCR8pXYXkBJTkyRBB2lpM+hDpIis/VgIuink9PaunM4/uKtvw5c9igkvnA6RTcc
Wc4o7CikKwV2lj8C9O6j50Lh7Oj+4GQed9WjMXG3U6afI+Uh3g7oQ1ONq2a4aQXSYIrvcRHT9zpL
h1KmPemL0aBVfuFbM0Asvcx220A+riScNkjA0PeUY9X+krg9nv1Ns/0MJrYoXTldXByjtDjhvj/2
6gFH8POZ4Pf2D6TsrpqROolqj1C5av5wtF0FBWDyoD7oq9ucyREA/3HTCHNpAUFm8Gqi3jxjgApH
KErTk+J054kPAA8dDcTE6t36RWRQoqOYgmYQ7AOD83fDgM+FXq5Jknuns1TghH2yifBNfS1bStaz
CYqySR7a3LlizewZeEc/u61pJyxoAHefDw5/iFevfWkbhMU/jVgpy84jNZtXpQJS3s/bWnadYdNb
sqm/HNjfWBEGkZf0pO5cz+WjkkO80q+dHOEebSGh/HLVzHVmqTkZCP0Pz9GchjXxjueN5IuVeI1c
9NhUnhhOHejatnu1rw2WP1O+tiprLRr/zGgogPwD42nf4CGF/XCHYhb+ltXyH+gjTyOUFI2Z+/gu
bsmVSqr4WRWwO/Cu+jbB69+J3WGXsuheAijaucGpKNmw63KrcuLBlNmXJwlZkTqM3mfq1uRrHZ0l
Xn62w37apfghWgLAtR7xNdtJmBg9+0f5dUm1VUmxg1QHeCXAHu/4bPoJVb3luQmUD2VZB6XP//lV
LcInrMSgpfAU2HYBRDviRmxBYSH77q6UqbxbesUFWcUeSfi66JXINsg9af/JoK3r+y+5vaiMwuW3
tHOlzeROu1SODdAZtcFdmWzR5FUjr24Npg16i+4WrK92GxOi9T31uYjrOgIF9zHM5DX636No66xb
VoADuBx4XmT5ZnOU6cokgtHmWLhkoPJuNfE7bxmuHm0eZ31YOavxcuRZmKqrDEIwtyrkZZqREsMG
npzNCFxwz+pKvhnP6P5yHBLK5fHeM+zPzF6KavfkXjGA0qF3VRGhRp9Rd4JRePZJ8/M21RvjtNcq
baszXNlICWYU2nXoKQCAEQDuba1oqZaGdJ8aVIXnxRyOGdDv/C9OSsukdv5LC1HLj+41C1wCKE4g
8LCOAYuwnQJC25qr61LXGJIYfhBFuEq7uFPlkbJNrYnp4SX9MOfsoocq+QfJUsB9vppIzO4Iknio
C8A8JL7kPU4WYBwHGi6a/CgGaXNE/O0LQ17lj6BIfd5a27C6mbFkrprqcXJ/V1sesCW0LBjmhpFD
47XWZNAbhrmNqy244p663Sv1eBDdoOp7Vm0rmRBaeI+tTVeqhI7n8yvWEOhkBn+IjK3C5crHlsnv
7Rsu3tt3z/0+dh/cOET3jVX6ZZi6NuKY4Ih8bLwXmvamtkd6h1K42hDiT1V89aYoi4SSTMydomjg
q5yFSIt7NsKCSs9424YDsLtExod56/4UR40/Udpu4zZT67A3kmI01vcTE+P7lnGE2vyZAG6jeU4n
K7RBYr3PVtxFN4mIA2gNQr+RMUqm814jiBHD11xGxhcI0AdlbwG3vogYXEk/QPs979YgQmnPVAqm
Amegg/3PM9/qJMascL9N5VzrEukaaQeJoDvCBA0VGdpU/T8BWHKgbc5nw9Hn/WZZ58jkhI1zI38v
dU94n/4nOS/4FYLj7hFwWEGkKzKweyOIi7d8uiCFmRYKIWFAg2qOxyKxuJNfeZR2M3x6O5wTxd1O
RN4443gM3uNwdmy8iXcQNarlXtCrWOf+0hvOmAVYzCfrgfOXTF1O3fOIulC05ZIRhEG54qWGp8Ei
bECvsjXr1+KvkdqYaZP0wEOwLh0TDnFB1ermr4bsNB0pWLBCaePVckmFEZl16p0l3VCa/K2GnjIz
XWDrJ9WvD7J0PnOp/kunJhUViXTowb1hd81+yn/D3F+IG1trDGxYQ0k2B/nrD+Y5GkAN2swSZkBn
U645tfyBkauj14OOHVfidhRxI6rcjeVKzGwfhi0ZBikefAMzhukUfbbXfphPUTYaLOW2bvaygGhb
ZdCq5fx2ji9wnTP6rBtbNX/3RW7WHkqOB09L2fSG6rGmy7DTi1AxAkJ/HG03FBYwAAj+3Pmesjgc
PYOymHetUuGDF865ZxWelzSRlGVAKL04lBVpqu0voq/zhczSYab3fxGxor4uiCLRe1k7Iwj8teGO
yKUiV1pCBeFfaawD0lFajwB71lqIGgJ02Hwff8fRpRWAWU8oAd1babKe8iDB2GYM+Tl0058fLLP1
4kNzEeWhGmyLVbtDU8fH71Pv417R47BqW+gzGSEjFDMuFMpGfkksZ7IWrLbrjvvXmYk/nD6KS/bQ
48qqwF7O8hwO1crMDNPVKKgD4S0yXzJmN0bj8qa/zAd8lMfgZ5cpnPXfG2+lZezDH+PPV/Ajc6a9
N6pqkz1dZ57dsL6ShDUEm0KH5KC9CCdKRy2NxF+05yRwiBP5nz4tQEAzNMqsPr1qZ28d8vdINPOC
eqXucsNAy8s2i/gUs1gVjz+vuyZYZ6AIAvTJ9Nh3AJK15TNwHqZYn34zicC87nabi+v66Vfi7h/y
VxVR0PTmD0QYRFe+I51aJzzTBeE5YPgIAhKZ34GBYt0NRwkcQJablsTs7nZmn44gazg267di4S09
NVsLsR2QxSfp/L2qLcgRHPEwI4nTrqDxAZXqfhuvukn8Vz52iE2ROPRhYkmXmf0A0N2sXIj7Xzlp
HVHoPzYq03cL0H06cMqYdJz+prgxg76cI1CltiQespP74Ru7ZRWycSlyzgkZuGRFYbOgNjI36PlS
+Khyoeu6eLhB+ff81poxVU45Eahj1TYeba7n2kmjMAEEXERIBzd5Tg1C2g3JHzcHnBEfCrq2eqHX
kryd1YrGFfcCKtsttHUzxK8vlRl5rzAprC8ladEN+aNX4fraRc9JQ3yKPiLz8KBp6aTKJNz9mouQ
NTzAkh0OFvI7i6kkpH11wUD7Y+fu+Rb9eTRdQg1aV9h6/J7F1xo7kVk9aQigN0ANCbCG0ufynJ6z
+OlRzNaVDh1vhmZ/4+dxGaryoI6USmPNmDDcix50Btmt70AbsO9HdFaRNfDFS7YcdNUZ5LJ/Kc2m
uT2fwLbwlzrkDEBVSenjKJVqf1PZLqZuYmMOe0Dj0cF/cRMEjN63z3pzHWZFV0jywlpAE3bRJzjV
zqM8Aec+VvzR1vojQgPWnfdY3Zjf7YXuGwSbzFj2RWoA5wl0bSLdon6v6u/wQBZHmImcD0CoYlr5
o4hij99/LNZ0T9R0h074aUEvAZ3lj//aZCj0zac2KCxvQQQwZNHOI7FWPkk4B3nmlJtMM+1qLlva
8Xk/B+/8xeLkdLrvdzNEhbWATSHFF9SjoqoaFO5kqGYpY3qUhEYGGFgBeiyx8QfZW4xTeZvHzLXu
wbKgafkKXmgf2ugdn6qHfezMin7fS5IJX83e6kdhAXrSO+/RyPq6wFXaSqV6BLCFha++j9ksCT7c
Zn8LaFK1FLju/3bHam5UCqJYjjBdXdqwJnM6FD719jNwo+y0lpbcEYhPv+y9bJTjcxlNA2mCCJFq
SKk5jULdNGpgjaWpXhgqo+4jl4AgsqpJT6MCO9pjSDh88ABQNU+uXxwXHA/2wcSsjWlBGg1YTyXN
aByUZSbtF4wjok4CLIGRlFkdZqOD3yEMt1ZHEm2Z3ca6iyp8g0vrDAHTomyj7DIgCbM3B1/6BJJ1
m80niVF0SaxiNLEx1ey41ppS2P5vQJIJCL+GPgDt0H8b3S60n2KQWyTAMra1GSNO3kiZ1lT15RMh
rrgoR8CTg/tKgQWgZIyrjUDIF3IgVgBM1CJSlpWRIdRn6hr7d+C4POd5bJcN8LqhikQ+tO3XGQQS
M9AIJ/blqpEclUXNoJ3OudgKi87nqjAnpUgHEz4E78fttMGzSHy+PXIR6XB59VW6wMkL/j4yHv5J
MYmBqsNjbJHWojWTX5SHILyEGYAgPu2zECdw6uY/cpXOP6HEyUMVdLKF5TMzGX1y7PCK85YZZXZu
cSkUr5kV2oSCt0DCGrRNwVn+btPL3IrRBNatwH8bQLmD7o+aHKJeBcB0ZI6kxtvcDxXJ+hR89Jy4
4w35anqjAcpiUn5CfnMH66XbcIA9oAUPdvpfUNmbt0u+ejxyBkelaGcn5IbyB6r+8SQUleJnrQgz
bsHWJhCy5fE+3+PNJb6p5JePZfjWdKy+yIErf+60rMkW9JFEcgVMkh7U1G1ioiFBJDgjLpuSDWfN
r4aXAkhGDPAMRubvVRb4KJ+jsgAtQ8izsDDqvkYTwSdc0Afd6Y3HpLhkI5d4b3M2yqvepXc8QPK/
lzg9tIOvqh9oau0uh87WKr0Of8ZM3q6I6cj56HKh1m0vnGQ2ivGaCLBYNTkmbW1tm4kc/IpAxc1V
NNmUwywJByQUjTyaMuM7qEKgik9XQ/j4cHzwe7wLpp7YG0jT5PSbiJ1Kv1oRuPFB8glqKwLzlwfS
StYOiUYA/qiMQwRPqSlPzYskSxgBecAdZSnFCYbXGu+0jfoXuhPOZkXqHeeWtsYCspWKXwvkTdBy
iSvnUWhZ9dwueS9HM9+o6ByF3u/kwuGt8QVZD1aCD+Ys78EQiMWgLrGibQJIOJup/XFyQHClicxI
VSPWP1uOuLPnprNqN8eClSWpjUtGZgEG7W1Z0LVMp6pvjwurYjjNftlhv2DdDxvKVPuA3ll1fuFv
ATC8s+T4rh2IbMj6OWPmZl4Ql8qsuINGyJRhI7dklH+cgKcHYmcifVGuQK3fxEAPEHxMTY9uT5pt
2nONlDUaDxRT3O6SIJeO/G8lPdxs492v7wxf0ALSBtEJe3Y5Iv5NNxDcfmVwoE+bg+UfXz5W+YFA
azSxndKeg0OamRhkJM5EWP7IM85dhy2Hq8vd2cUsLk5HcS+SbMEHqjq8VFDXoCo2jMX0g5fUOtcO
3B60gsFcEDpSkokah6c7QiHXGhISydjuJeuvOPsdmGITeTNc0FuTBO540b5XtT2OXoDPyzDGhwjv
63w/sM6QlQvNDo/PkXhqHEsEO+WL/aqkAZsoMSBbKRG71qqlvraUamqt9DVH/2bELXyRICIvWznY
s4cqGTgmwOtbsyAXRc6TVkMK4fvH6p3wDyU7tKNJNhdX3CpvMj8RZTyiioewYLWug2wS2DNw+vrY
cVbpM5C/cmF25n5/IbaeYiQ+adplRrMXVCkt9/pK5FOB+6yhNUDFtXpudT4yAkRBkoifJ61kuEGE
8/Fiwb+75Wg8aed/EjDRi3j7eUGAkba1RMhNHw6c/d1BOz2+TqP3sNctt3XdlOMYZAuyREIDelGB
5+n6kOdNLgqE/dPR8y58J4TTN++0/iuwQg2t3lIUu+LY875bt9i75zwnKp6Elqmv/8s8v9KZEYYa
RR0s9BNIBCn2PkGCzpKXhIZCclnf7M41SC7PeHIKzezUqhippApi0a8ZpC6JxXh6/w2WlODMKoi1
ntXzEuQUSsJ09wv26tvfScGZFDMmb5InhRjl61L+aDxNcWdJik8rO1IutvWz/7Qjxe2bMaVlg1q6
1D6C2gMz58upLm1BEz0DN8469xYJ6UvJ0qzT7a3eTihcnugpPr6/lriSppmTdeh6ZU0C4O630bSC
zy6nhByQPxkJPpRHUUzmZSHee8hPbpcswMqb5VaX4v5t1VZc+vidqTThk4lTa6PEJ1Dnj3f8p4dp
XhoHFuaPjI2T1qk7ieK+f5xHRligspIA1Gz1gTGX7oxpdQgfv/2adk2GCEMrn8ixHcTY2rAShBMJ
ipbkIwDYZZXyz1IHFhsMMUSIJgzP0z3giVBzoWVBswujO3IC6F+qvbh2z4fqXTYAOqmM4mqlKB6j
CgUPxrZd35aMyXz98EQocxBKB1OZrcTdQEce2GELyCBrLslKfShYKuvfRqt+S3srBKfhuOOAo6IZ
fp3VfInvJFzBiFXiAF4YRH43lPBh6NSgt1+cpdfvjphalqiBK1+ipJSR5p/UnyTa4xJ9a/Eh+IER
f1nJEANZ59OomJK9d2rHuZA39N6hxIieOXTN/qOLDtj0j2LB4DgJxdBasroDW5RAIt7y8u1h3fOT
bmNTTci/58gyHroslSU6kChwQl3c5OMXzLsTcbwL7K9DSU9ipin/6cbozhGz2URDaMZgyTpi5m46
d2Gppfp14uVfYlp6pjaJSjXYB2qicx3ppjO1Iof8PG15YxDUe3bO3dIQZmawLS4uMB6ltuLSM5/y
2sxgPOJDbPurFiRikPOEMljbSs8x10HEAUaDUgzhQYFpCgooiCQUzZ0e/QfVXFdeJWNz8PFE6xMj
zyeH2tn8JsRfuPg/OTIEKlXuejIC3Bj89ry6bE7Ez/4JA3Xq9rZWZyybuWwjdl85mlNbZEb7FPyD
QvSRhdjXL0zk3YujVXmJP8P8Tr9fvUPQY3PB0LnxjXdKOnPGDlOz2W2hJ7WO8VdyuCx/A7quL7ys
OwBOcShlkClTghHteFqTwXF7cZj4j2PVkWQ7lcsLexvRfPneo8EQFv9zkVJ9lR+DXaSuqACmypER
3M5OFdzguwfukWQLECIGhzj1gu/u1BkCUhN7lxzeuqLxpNV83cX8s6ZFyv9zzPGbfuqu3HniBDp+
33v+VgSFyqMJRl9E02AF4YT+Dj/hhMIsxfavA/ae3/8grCU1yOf3GHSuZXprbwiK2tEZ1Rg86vn4
00d/OWb2RAhpCu8ay4OKVO+Gkg0VExGe5aUD6J0Vfz63+CMkTEZNEmQpNKFI9ljRu8yeAujXq8eZ
4PhjOU/virCUXCbA+Yh/FkimR4Rb+9DR76zpK5R9eLDcZ3OngQQ1rBZg4yqZXO59IiR9Q02Rvf4W
kF3cwCQerbgWGSRkL5WMFfvAZ+dD9+UNsb5wY0KbKgIwELUSpDRJyohU63MAQFK9B+cfM0lfqJcx
ylxcTZQFOLEMlQJn8OqAx1SiR6hlxwviY7+brrXNAIaVf5zqQ5wMZjrXOdkj1Gf5UN/zJbted2my
HiHpQJEpz/aBfyTU7eIE0zz5xypmpJBQHRJiub+SOWeVCX0ui3MZeszhIsp/Utv1ENoFVIWP9J/A
4AfI+5SSMB/UG30jQ8nQH1OGb0B80DCYSnMRD5bmA8X193A8aF5hpD8uUUXxr5dfyaW15nHqsZyR
QjeUgIEna7FWgJhozuUseeg2FGQijEbbOafJDeWB71YRX7kpxAhrKY6EAt562u0lFqCVDKn+mig9
r4KjQcXhTF6G2iukUdKesAnLbdtrB8Y3XaC18Tp3F0BH2+VjN6QcE0MDtq8IMZn03YbttQreRVkj
5g0WMCNN/iGOYzMF7LL7Pi4ZkcB64O4diSWGgZ6Hbd5uRp8eyl56DcNvjhp/M1jvAOpF0SRuEWGf
JMkFQtWMw93DUGgrenKwKR48oRbGWDfw85gf+LJpwDFxKZp/kuVmzgAZ5sFWkxmZL2abktR3LVPv
M9DoReAkT/s8E8aXt2XGubUyTSuBvv6v07CWdJ8togTcJ0AW+x5x9VoYBoEy9ao4MQ9EeMqtyJUs
tGWUIEnl1hrHOScU4fHL0nsYtYyOpMGVqQMa+psI268MywofUL205PEOt7vX3naFY2I+77DpOpQ+
PuRLGN7CXzUdQt6TYSP8sfyYzQIvK6LkO5cR0rABOKPObwcRkDMfLxaguebe7Xs2irYSs0ImzxZs
pbEg7PzHS3hZ4YR7DWSo2tIxubIO1JmEF/dKaJSzuWwqLGw2WIsQikTAgwyzco5Eu5V5JK+2XjN+
P9cOFsWB0jr8TQADm75bJN3WXEz4TAQ7ZoTmxFt667wgau0nGzYO/xjgGtKMDAu9Li+7ia5ACY6k
KKesVZFkEkdkaGV9pV/9DNTqeP9npbAZsFad52ZuohfRFUlehMscgvxPbopbHJwcd+QkbC8mJdY5
YZf8IwZaaTR3miNePzbp1avVFUXq+E16DoPabSK/4p1Wo1gRSin+m8cpN425rCGp5s+Z7Decacu4
MyqIueXKvtxxldOEQP1uySTvAssn8Pbb6gzX3RURzoZtoUegIhJD850UA/Ewyqg8A7FVTKfLtXTW
00cw6ITZKAPkK4ni1oOvLWQsPMS83qTQf6TjlNKGSI8WRs2hlGe9UNgBaN98gx9bds78bWDGpOKO
fDTQx7UbDeLpewdc5qvXC7f4UQy7dAhGYRKpKm7JsWxwlfcTBDvAgpnbWjdSrjPm425vQhAsNWJe
HnDfcmoNqxC2zvBJ8AxaTdcFonkEtlKF20bPHr0ADj/XHowtE7dkWyxdAz/WNdpIOKqYui3ZwnIh
rZSNQ2o8UhsgmT9Y6uOhEhmk3nr7lltZN+rp6wr2Sidq5FtLS4Q1UqrcNfHTsPkgXprYpMftzJfV
IIg36k21YX/sG8yBQUpBJzP3g3Fd0JE7uR2qg257CExH2A81cXM/YVqRXL18LXg07Upa22nQ/0xY
vMVQ4Y6DBMC1i+M6fNH3yYHC9xH+4gaSXeIKsYAuDlYkHuN5JqEvhm1sBI6yMT8m9fbkvPwxxrby
Ai4jGPNSMRcRwcMC10xAQFppDCRcqp7lp/NnBLC7Zyq1byC6YCUAiXU846deuMJz9Slo3vJgUrVU
UPXUaj4unkvKciGi8easpo7Ugh1Na5PHGVcCziFTxEP9XKagGEqPXFQjpewh9C7G9o8L3lWwgHWU
R/pej7z74yX2XxrMOP83vaIqzCKQYlIFjKECL2OvbRSaSAvD3/1XHNlSYwL24tGHTNRf8YYA+qHn
FKYafmZlotQWonfjgxST9qR2qW3a9oJmeLXtGjUw8FmXCZQXR9BcQGsT6FL5KUEUw55/rbNzFjxm
n5ckIpw1Ie5tr92l6PPIK9wH7LlHliDA3kbLc8Sxncz/iWTduF//EFW+WYaTtKNY7ftchyvnhJpZ
CojjzMdh5BhLM0eLR15qN+sDu22EZy1+HFVNapDR9zR8vcN2kZ2mDlt9CPx6rKybclDH4CBILAd5
0yT70Tyiam6xyFQzT0cTrYnz2Q7AAFNU1qUB7m+4aq3gjz0jDvfsMFHwZUJkAgmFLSKB2/UA+n0Q
o6bdcr8aVs6Hnp2JkX9+vcpAfRfYbHu4zAgti/zPwFmoo+I+bI0MuYtWwX/TlNmeLZWeKy4bOusJ
VlCkkg5sAdiGOasYNqrb9hx9T0rjdz553iZ6VrZgr11VOb2q0j5MjcrXniIYGpdiTdoIKIANLMNn
fAj6P4lg+rIdVobOVtuCufKUfjLJIoRQZiwLaHXjClTaUi+dLz1r3EFzPJC9BAW3cZV4qMIHI1Id
SBw0/3/ojyKL3CrU/PbMQmS/5iFjHjkknT2lxASMt6afhl0beoQhnQuD37Dukk4d2U8WlKx7TTJN
hTEFyxNoNQXPNSgkIGhyeJYJ4CT31BdlAEYHJK1FgiVkNOm/yX1QSGLtEZD3wOL9SedkPkB7diDn
R/YE1mX58jNKleVpARAVvt40HHKD9DIL/ywYu2gatOTklr7i5KJd49MKRa5sZHEaSFPkzRNp1bLJ
nWmIAKPz9icbfDYGIlxr0ssR/wtef//9zRW80eOFQLSN6h+pNVQPeChlI1WJHlzxvvKdgpjdXoTL
esaSCbGIr3QgMiV2d1Ooz9xbfh3AGIBBuQOIlF+0X0lhcfvyeMK7Lt+ogff7GQ3CTyUnhkoKhZwR
jrwjEMOdpdRfek3iecyfn2kQvKwwaqMMa8XuRTl7zXn4C2rU/3PgPXo7HpPp307RuQv4H2BjgfxC
5nPeLs/qJfCcu56U9Vak0sbEnBqJEkkVjiGFGNcMYxzYS2Ka/zSEsw1rVPG0EKrobcB3jBHUmZgd
csjgguHeDmuMPeBmvucPoXWz7buhC7/CUQ0R2R0eRroNy3gRm0Kt68364T3tbGrtRgAGiy2qt8cD
Mxi+BmL0UwHuzpCcG6YMzjzoLcg2wTKvtvA1OtfPSQJMbIWlIxrmkFIPKKb6EIUpZ9JKLYB4lcoZ
IpFBMBDsXH57kSip9euggrx3CCpNB7GMZIz0n91Kw4iTXSYpmqoz+TXhqocvyXLU5RmBGJwJcRDN
28f/ROw2fdYP5kEbLcwP7ffTrH9eByL0o+a1kb4iLixbPQ0M4hNz/l4MFHiC++IFPC1fpgOoHznO
kySfdmVOCd2TznL0B2mLFLA9fY2LzV61E5wIUMnax3wOMFpIJUPp0H9pT4rXIonSJHJrbp4fjF7Y
n/WKc8ZOW4cUcAl/KA28I9MNGShmtpTIDBdxoy8gHmAMp5BNeEjX+1V94bJyLmzqkj3mm3tglopZ
N9uRGlrgKG+h1bkuAHyoqrY2SVR1tEnU0nrTctPbzWY752AaID4ic7JShDcXy7m83d1BBREZwnCH
6kkThk8/TjH/51ZkeNBesaaZj4B0kO56TTqWgZRt5lxhacMwJcWr/O4kqGgwcUYB+/5ljZKrNF7y
c2Ia8V1tH2pmrCvLjqRenNftlUuBsJZovqwWF+o/bwGJXX+9kS0Md4jivC6wtLKLnTxM5szZM94V
1KUakjxo7dhRhDb7rsPNmgvhzmqF5oIgVFUw3z5NNqkkzgz5IugiHNh/UtgMsFEkWXU2s3gwVJaM
b3oBlKcxRYLoKliPo1lB63enN+tp5lfTS6mseq5mVwl1maLGTff5VjJXXVoaAtGhd/8K4xRQtd7Y
bUOeKp4HbAv4EqsgDMYvA7DAEIDq4KKgN/5TxfGErBoH4XbNntGnXb6okmHoCqfoRY5le15oqBFG
PmpEozeWtkqO81Tj61dtDuCXXJ8jy1zTj+7yZRI6xFe33XF7bEU1qzJA+6A658IBBSDG1nyFKRYt
zep34ZBnYISQkGcO+Rxe/Q9JUssMbo/tO1b2dq3cvPh1PTgOEK00bcc6ZybUNgRa5QFnpnP/IKXU
f4VpzBuNVgLUHJqYnfCMi3fvZsrONpcm7tjhw8nqG8ytYpMAW55WHo44hFe2ZedIFmvSERy7VXmq
RchYruZ/fUc8fopyGHpCQ9azBhrQMnH3G9HiglfQh1d8kutXwqS5nExFmiz+9fP+0mbD1lOsanBf
xQi0OdTGDFFt8jGWVzw04c/u4V9OPY5xkp642ZM886BMlTPR3lB0YdqpzT8F0owZo5qD4hDKKc3d
x2CMHPpbUzzFXpMowT9DmBORA4/GYm+73f2dJlS0tMZDFTi0XCLLfj85MBulAXECEu0sEK3Tt9CI
WU0g+lIRLxpiawO/EHww5oq9aym2wVJL1hEX7H5mTexWNi3QltHh0sns1l46XNVJjPgmO4vIZ2yx
11R9CL8IulHxd4CA73RLrLoL5vjIKR5BDBEoUA0uUR7GDSWbM/T37hINlklcVt9rP8H3JfjL2mnr
YnJYXrt7iez6hXEII/h6xW7w//Ez1J8JW6DdrQYBq5CFiTe1EOAjlyT6+Il87eGKWLIpNx9gO8Qv
Wr/UGyq+er14bjmyV9nNRgSgUDmw6+zEKfVyEC7c8Q2LnGjT0zysKxLXK6TByr5Xt3/Fz0N/gV0M
tqEqkt3E7N5AumaDiGBx8t2tQqf68x2geHSoMTrUkrc4f11iv6MjePLqWmSQzKGIvA/RH5jyCt0F
nouE59BWhJKsOsbs1efVu7cmrb7oxmHyRjYl/PvWiH1+NJVTdZq86f0REseTEJhdt6xj4uJhmSdH
eptPmiinLJ4yM5awMqPHZW4NZDnQ660gt+R/slEHJFEqbnYxShoMKxeTTNbYXgFUXWi6T59Y3Fqo
F4eb1eQ8PtIWXKIKA4Av2KsA+jDjj/oA4iWPX2cDvAJyyC1KKEBtJOllRVDFXqoIawOMaWBCfALU
Feb2EN7v4PmrL62oEcep/C4p2ezKSaJ55aRqs641HW8LQgDr+7Qambf0Wn8ywygBBYOpxTRyl4x/
YS/EI+d77jw5E17/m1JmtHy5Ti+kTRKljyk+gnhX/yBEvREFuSZr0OWcXjjSjTqfcq1EdDf7Oy3b
mWJIIPEhcnrKxCR8ZyCOh/oaOfKgrVUILAXPD9fKKm/m0bfxP/ObcJVhXVVhrYKCgoRB9QDU/RI7
7hHcxcIggiABOPFS+PknVYAE84yVD1BCBpAmLdvBbhGlXXB8ZCOj+k1Dz9OYWEKpBRYcx2zq3RDr
/2RKkm4Dag10C8fT+GJ7lgw3/BMFrp2qEahrSCH3kn6g+UH9bnxy2sz563OzmiTm5uaSzpjNUNwE
MXjRFmLVioUXFA230WlxFSkfniKyVqLB5ZCUAMmfedk0UplX+hantdg4+OTWBbG8UgD1p0rwrEs5
wPZTZMRAEnG59dLJlpW+Of6ZfdQjHjr/lC6kZZhoLdcrN5u2LCLPzXMZoM9YoRKyuwOIVEoewt1i
ghCsnVzU00Gw0eUCV24VcsABkBtalQCGDUqBrnWvYgtlv89Lv0ato0AgoIm1g2VE9aArgcmvm8TJ
pqKzQkCsS0M3CFvcZx8QqboQs/iqYECOX3813qLOqTRqOqFwYJqrw0so0jMZsF0Z4qTO9yP/bQBQ
71yhbhjxdIlAiNU5wbVcr9sPg59O/oGD1F6vbibwf5lRQjte6u9T5oK8cUjkh+hqmICI/lytGDay
uSNp+H48O+CVxDBCl8A0djL7vZeg/VgnfyROX4380L9z05RP3YIwKe+615SacofCVPJ9f9xFaSM1
WIkUheOVsXm9K3UxiolJrbAGuV++Iy67x6pySOXiftSeawavTyigIrZJMTVXErQnws3Tvo+lz4wc
QGIdm1WxAZUjNxjSQmVEDwjIiItm32ZfCMcSI0UKAKA4B9IIysuT1zWjxdKWSzfZs6pym5rWt4xt
XSM0/DaTuNo57pCLPQzMHia1swJeBJ5rVIcE61SPFwQLDSI2uF5unYL29DotdqAxhssYB8EKRpcg
6ffFrrBjW1UmvfuMnyHbBJ+GRG/6MZCCdDcNUzQf+PTBvzYdFMUskKVQtL23g53Z/FLFr1G+nSpe
GVfRjC/f0QPfzOtKE8b+MwydEaO3GQiJy0+5LJjN2GIMMKT09H76CvZ8lPi7/7JqzyDtWnlRu6iE
4016K498A960GNtsQwXLS+lw3gCZqxbABrUVlUOWi3VUROMwhN6BAHeqXMkJ+r70pE7UBxgTZjZT
P3LWOIBmqzFDUqr1xpRI4lXHcc67Y9oJkU+eE9LXhtpWJ68Zk/kLV8yW5p0UT+UcYZRM5AwbV/yI
+VyOYhidBGnoW4tXQW6cB2IhM5jNMN8ulMZW8fGo0dtq1CbionVjRlvgbQ/2LsLFTIf/dWfuRwVJ
gidiq/A5qQaNLdn00pq1zZ7HfJhsz63NbzjOVpceAobASi6jF+dr6WmQDp8z4JYqFJkWt3rD0fo4
d5hxt/fxswe3+bh7pkXPmS5uDi67Mq/t1eSXrccsut4UauOIfnMkJxfmbabnrpvAhIvHdFRtoy8k
MLGFAOM5jFSN9kEylaYzOZOchD4Or5xkTq1JdQ8jpqnApmUC0TEvRS88LdZmJwEgbVtRF0Mayul9
Q/GW2rypdh3lTlcQd7hSejFVIC6Yu/lw8W3apwJRWZ3px0KqZHIvDHWe1urbGdbM9jNpalaBSeO2
31xWSQoCFSnUk6LjtNCPk+4ZZQWlS4zSKq6JOLtH4cUwvO0+OC/HM9dtauKSAUwjzrj3P3lBYJgY
1onMX/J91MmlmPB+go8uisLMKuI41UGq1LQ3Sgk1VnhZm1CJvSNXRnKuhH1/X/qWtmXCGUZKOJ/4
D7uFB4Cn66OwUKqBIgQrS1AqCI4VvJjDHszKncDaZKACPHjuCPIN18nsPNK4d5+3NG5RhUSJ4sp4
LQlwPqwK2IG+OpZuBqDLqiJHzkUK0bl51cU5NfxMuN9jOEXUMj0lXpGKPz8tBon+w3EhjkuBYrND
NAiU3zqi+V2a6IMBlNWZQ/7KovqB1Hf/Ef4GHZeLuY9JZCwrlmSVLDpXDtYGe5pwlHrVXrS9PCM7
g1fyV9i0bS95TT6GjvWFhO8TveMrM+Zweb8lt2kckgulvQie6KuC6ggbQLoMY57lFJYV3brNsVSu
e4YvMtK3+PcCXB4RZfrrEWCFs8/iouvdM66wwBsz/X53vwDq2h5MZiyC4+L1agyhLV5u+f6kc70Z
jEhvgqIEdaPbGEd93HQekP8J4WCzmvjty4VQvmwF6mmk2f0I6yzb6Xce9cqk2jY+hXJeWl6h0MqB
UhUtoFX9p2jolhXRLQCijinZNqYAvxlqYz5mH47Mg52yzTRKGm+HFMmGQq4pRTXm7Rfa8yQkE5QW
HWA8jnJqB7AaT0ezuVl6/OxpQoN5E7UaUWrEfy1U4p6f6eXhnbXaR77zHjddOby+BQv5795BJUoC
cUuDYUOe2AcJ4c03xmFQMiKBzvGYsRIu0q8yG/SEYAEUmijIclm48dLa4FIHuUVpqi1spXi0cQ2t
o9/wi2dRUsyEn9fewEFJEoeRsSmuQuyXJHUiXYUQrV9y/8IeKwkfw05PMYn43WPIKESi+tN3PLXb
0Bcl8CoKM+GLNWwmayroNJXSJBOdZEyrqfYoUpZ6XPQ/meql3n9M+UwV414jXJbBuvV0jUF7yjDh
YDh2azKq3gcCBd8/P+ihpay2XncNaOVoxT68KYlbNc3BGbdx0Suvlucz0metBea4k5dpO1ROy3lH
LjIZti6VC3QXfcwv9SZGYGNkyZmmDGFCp6AJc6czJ4iwwdKnjxHIH992hYjxSyVHX1UkdQ+4mi2s
FzLwGxinS73Ks8yhu8FAWpFhd3EdbkL0yy8g5YLff9VO4zNSEbEO8bx1WF3kyLfWYqaoFDtYKzo5
9/s6GU8MVKtEniHiwD8hKyXCaU5N8aYm13IxZ/3WqRka6wm5iHanP3HAzQgTwO2GHfHGSIwAXTKA
7m6wIaATdXDRpzq8PU6Xs2Qvw/whqPO5W3O8B4wq0s8J0RBib7orjPoEMbdr5lYN/WPYQeEP5vhZ
bX8aDu9qtrgxUvcjArGGRi5ijYxtefL0JUXxVMjrugX3XmzXOmkPdloQveVfbimFo0uMj9Bw1c4X
V44LHxqakCPdEPFyTpRAIkL+PdhX3YW/AjFq/YCO3rGXv7BTfJ/vGfESCPWRwuZEmVYz4KthvSg4
Uuwh0PpTh1CIz7D3EzaP2t51zoWOh+rhXeVOqNu9GrCdfOhjg/RTT7FxnYtBRCRHLV5EYDCdyB9O
HUjukmJb5VIfSzb2NTtvdLmzUHokO7JSneZqEqFPycBMrZ5iLn5omcrUad3L2gt9PqnYkAmAUzM0
rLsP+1bsUSzvBpvFhN55ulkLF1ZNZeaFcOdJVVXJO1RLffwvXwmQvRDyCqRUfcx5ppXc99o1dqS5
BLwpZXbS3poo0nUaRrlxy1dmMNhSD3g97I/buROQ4CEyw5ljN+LaN1LFqQffGKDFt44JvxmCaqDe
qX02yK/Dr5xBfyttOU7Yp2oBA0BGLi/S71I537Wc4uJePIarKcUcD/lxE86rYbInO7ST1rZX2Y9t
UPvDqQvVf4mQ63ljOXU4U3iub3JqsnIDhJrNMgims14Yr4jbg0KoFKya43GHvdPPfhPdsFc2dFke
lzGxx5tE/u7wXpaw5HcKvySUHA6vGPyvrlXFX9LWqdl+InwZAN5G8TMDyuv8y67z6HxAxv7Qbk8o
WBY6IRG7zBN+m855ZP8RJzhl/JuMJZuwd/h4bTmOTMf4WQ3KnYXpYVzHqNxTRlcVnk0doRcfkwZ4
/p0ty6MWdRVi9W01+GKHFApN8IQyd3wol5hOz/XD/nqZyVg11AJVw/rpekMYByCACbDww/Nu7FP6
ul796LN5XszoSkI0d7huy1ejOVVmHDxacq3ZEzuh44CeTqpXdGHdMVm5P2AcF7Mr1/hKXE61K9oe
uuzpczXR884QCfuS7NvN4Dsp82+egGe+/MsGFEnc8Na2H+vM7r4U9j15jQRDy1aWYh60TOe9gh2O
lB8NWQLtz6/t3gju4DYohGNf9jrNct4hen+LrDyyNWmtBsyoW2ozT/WaPQhNwJ6MQOTLCyzzd8HD
LrE6FmXgDvrwclfkFXastd8JhftlDhysqgTg/yBrezuxd59JF/kv8WMtyTaWoapQAJxvaYxHtEOQ
CqgU+af98nCNrVpTGAtj4FJOeBV8Zv1HmTdcGKlhirsivO46Rs1MSjtL40Sj9f/wzYjfDeXhr0MF
YhYbo6UnU0I5z8snoCsUq6i0OWz5lEA5AWnZpM7EAub9lKFv8903XivXJso1jKhVrdwjGUQBJ2j/
cXYz7HCLUeNKcz1SLqMKLB2lcVLXtmgMzsCxf0cWWkVL1AvzNQHmmlyqqqVs3sTja2rSykWTOm9z
3fdc1O5a/c/NRck9WGX+Q414qQCh3qffBxbr9qTEuDrSr0yXcR5Y13fkRBSddar0NGuFQcG9VHwR
p4U+WHAnhaSn5C+X7F9483mH/wbCFRUu/O/NWIBFo25zjiU6QivfIEYp8oi5zQa5F5OrPRpg1vo5
lAAYjoBhvaZxXvYo/zn0BWsuqI36XcszZYcUNsrm6HWB/S7JsTt7suW9Ujs/TzlyZDde8mZQRLMk
gNSGykiJmpxXwskBiyqv97LDw1+jjn2kwTE3DAl/ijE2Vvrs9AffE+wwrXj09EPd4e2aVjgNB955
zGvN2GF8FQX3HJgmEkcW3szztop9rWA90wgkbCtscrafGI2op7qPMpZDdIch7efiXVtxQ+c7fKDV
aEZzzNFbVDWFRi9+DcqybWKhJVc0QlHbFQGqYEtmEgu8GDQisa4LfJ0rBT6soXa8YD6mYRLe59lX
Px3vb/Y+TsYnZSaLk71uXB32gwdVCrHxw8AplekWZeMe3f8GOTnxG7KUS2P3hSdkzNxGZw41dYaS
Tf6k3NobjP/NUterApxDi4KOjjSvsAlbyMxqGvyMC04QUbuIeeoAoIrbd9X/plWvGwQ/+dAx1HCZ
/XAgrsm4EJ/mVTSuF1pI6Ts11W0G7BfZobwXLeiBfV7XifpfJISw/yCR0Kns8FNmpcCIfbKjQHnp
+wzaBQacG8XAHk7rT9i0TqFiVsJtvfmXWCd1Qtu0FP2bvijXOJppC/8qonFUja+CkAzV8kNL5UNO
c9iKp+qwxD/X/Dp7NmhssEqJHo4Zl+xI99lr8B/XFliqTghcceJOZek76rIrf74++Zf3msW8eBPs
IHdxU/8X1NQjSbQcE4E8PhbahlAABRSyPBxLEl6wDij/Tg2QETIuQqzr6H/Vhj9bCgqnCw5jWKEB
eo46/dRHIExzC1XLWQ2oFo+VJDqHfoLY6pgGjTiGruk1iIFsRIXDQAVV1c/mfsvX6szBdaNgQ5pY
WPBGVMCXVNtuF/Bk1pbZJAeJx4CW3wAM9Ogec43ZJHKdDJ+g9XeA1qEHDk50vgrDlhE7nQVVnpom
/Tkb39969NqowxoGjVrKYUvB2E/BCixpoM97gmHMNw0giSU1Nd3hjyAurVcFXcne7TBqQ58DCr4q
zPi2wkg1Z6JDWRfVl29h4N+sJ0uYsCM42vQulmdKkvOzsOyQEjegF/KVOiejv7sYed/+g0WKrEzj
M/XCxXpd8en8LWOuokL4vbL4kSanQ2dFJZmTWxUZDEnlRYNoT3mPOv5V9+pIRHjxC0HhFGWmVR5A
TW0t2HaYD3xMzj3zUEB4klZGJPDyp0KvQ8jbxyZTgSTHkSXKrRn6F1HhEETT15jRKfYoW3dXhr3O
+dTldNoIVAc8RdRCt2IqY8SKjIjsNhj4CLZaKIYVwAqN2QaICB3sV43XZpdrLCVVXAv0vzIYhliA
nVD61QbvCrYqZGNTN3YcrIgDsnvQLJ3OwEguHcWBj+1yoGjs3bNtEfrEtMp7RwEf5AV5L3xiqf8u
D6t/Miw3FdW23pcrApGlv5IfStT0QOm88LKH5afJ0NJU55F354ftZl1AfJOj341dSM0MY6xFytr+
1+aN1TtNur+B9ccyNZZxQc9/kEL3U7oBeEwnuELVpPYobJQ0DjXwpx/WCI4zdulxZn9YTXCkEcKR
UWqplNSTkoK/poWKxYa2fpOLYYV3h8h1eFcjbqcCYSIDOU6bTPwQS0PnVURSLpBPwWhHYi44+A11
FP/HQhYi+1Vi9RpsM8B9RLRh3A1twIo4F1cFkZA+5ZSlxEO6gufrnGT8m2eZ1r5Y2iXiyNauydS+
/DkGLQtyT0KSTIc61+8YaxfNI065GwdHXB066yE3TSNOn5j7e2cOcy3JpkiwJYDcdOrZDHBgCaVC
mL6gAuvD27Rxa4RjBwWfQG2PaZO7bbfWGudd2sA/c2qLETSOb2YfHdE3F4Fz4Y0LC4oqwgLJxoyv
CF8IGnenn47A4MSDmL5WfjkoAJKb0qho0Bhr5g7m4GUUQ3Fo1FYr0JpLwIe5hkTUB+GfzVD9yeUB
49HV4Zaps6z9zMhRW5SzdAWON+vDxXoNgu9owDQQMFEKbndabaHTIS0kXm1dUeZL/k+vpMRpFhYu
bvQbKKjiBoEy3sPkkCe9sgNtzhKiNPdaN86ja0sdAfmsFK1K3MH6KNZQOF4sRsQ9yeTsYG5vUswi
xIPlBeLemOSK+enc7PBHlYcp13l1BB30oUTSuosTLXB+f9o9D7cHgsQ8pjazHEi15Ztj5Tp8OujA
7pMp70dY06+ujiN8h+2vzhdbHybGDLH2yFl8YORcqUzKGfOvyh6O6fR63LoA97FY76q+OGDCEPos
E8vEtIcwgFQuXo/ouo6cJWGfeLZ3uv+ZvAjyqNimkENaTwDcwqKCMg2GpfPRhebPGNghrKgaWBfC
Jq7t2p7tlr9aqICh0Ne9vKGbXOfUjV61evEG5l3AFC1S61bhSEolFo54hLJGMAIJoOR0miZxwf23
Uq6vLLkrZqXsC0vgMlt4yZxK29sQtd6SEcUTOR2a+elI/gN1OaHpbr/y1i5BUYS0xMHXtVYhI7cm
guUeMuHmVoHhMCkjnSrT4Me0PnXM48SzzuyVwlyZamxQmwhFMEFlezCy7qMm9pk0nWLsMSzsSqaq
ySubMfyvetuS7aFrY6PJOixI1T/OII+d5iEqyJgHsJOogCs+SSEJGcMGElNKPMByd0rswIdBRjAv
zuaBqTvv1/zaCqPmSWm8i8J7gwHZ7xXaLsND7pmBSL4XEzHk/xC8OG05Nuj5Xyj8uAt15KnQNk1f
1EGIP0lby6hT/OOQRobC6uS4JHShxy0VDRMwcAYLlYqBvcGQKbTJAqlbm+mC/4nhPCotPLB0N4nE
UHQ1bajye8ZYFimU+Zyir5EMVdsGkFucuAcGIvTckstPh8mH9LNKl/kEp3SPETEeSpDiGRt9Efix
RL5ba8yIyAoyoLd9b567pUGcIysHFQNoz9DyJnKtt+BtCd2UKgAap7NPBMLJACGDMKlcxybyNTfi
liU70Ow76Q7oWccmxu/OWuDPQd12w/TLxA304z5+zNn/K7j7WZChJRJ5phvmIim4+uZKujZOEmfr
Ld31JhP48jHxI3rE0GuBjYufsXQWbvl9gXWZHkXTbcqbl4cVSSniCJ2k8R62v+s/QF8V/qE9iTaz
tNi9MBpiBwNcW1EVb6oaZXtLTTSH2eEgcb5h960Cx9/k/plrov9LqBVCmupHkBZCKp18uXLxvMFO
Oa+bKrlZgrkxRCwEN9GDonY/BHU82OG8EbJBZGzBsR8SpwV7EghsZ32RTCA1ouSjzLOgNUNqkhAc
/FHBICQoMFXjlbG8lbCY7Y5BWATxvLkkG6k/TuHedV9lF6BJIeSDuySdXnwvzOf8ONsYCXZxuiH3
Hy5uxWU9B1d07dhSISiEhii/I/v/RTLqasxl3Yk00p1ZYt3r7UiYm4DGy+fRdxvnr7n89y38JlIG
cnAg1dyWo7lWZ8vGewjk5uvcchZAsrnenrODPz1BdMa9CHw5dKFjehsvMuYXlZNjlSIKMhFzvLxs
XEfMmtVZFhOExe5JpD2VXqR3xQyn6PHaE3P9o2xg9X/hbPpRJDZJ4V9LZYz63WrsrcfobZsRgbV/
BTobbUN+hOpMXOVzVaKB2XGLbY4RXfFQi7YH5upYd6+nDRxY2VT0a0xGErRPq31V5HuqtoKuxQEH
lkT6Q+P2Pnb8Z535T1Itb1xQexu2ZoOa3pS0yE29r7xwRexrYMsKUv28FJYJjCFNNCOb7dMSXqFc
Xhw8ZAsjYiUhtJYBRO1QKap1cUyid7ttNo5T1PUMoWlg+2FXsUIshdJwM5f/CrxCKTurLlhbvb+k
CIMGm2988Jbz+Ampco0noeeBozKvj8EK1a2IefijWWtNpnEf8jb5wixSySl62W0gSh/4+lgVXN/8
Dnoz+bPT5R2waGXl7E9p/Tcjs+E3hFSZJ+81ioRNPYuqO4r7yvzvvO3Ei4uH8Jre3CSCdiVknchJ
YnQXAmsApF9snXiRIeeDkzKkUxE9PPahP9+6ksA26+/Rr/D0Xf4j1LYvSPaPjgx7O+sqYY15LrBa
GINpmx7FsuvI0zPjx95toGEyYLyyYjWcBpLrJmc1qU6N8hMjy3PXQ9TrmAFkcBHSoLBp5mA8K1qC
ty5A1yz6QLyQJ4KoHXxZDQSD2x1A+MILXF27wOmoP4h7VNcH5lYKh8nLZFGpVsU8Ag5s9hMyGeFd
U3cc12RJr58EfEEPOlKCVN1w4cd3Izz6uqAvCt02SF4deWbcE5OjF1aor3UIqqLm+GlR96IlQoHZ
eoPExITAd66eum97J9r71Gx2pjWXJu/28GEDwEBQGkKvnvm7z5ZACkPVIlVWDa5hEYxKiu+mfl2l
43gl9hd5RlABQSowzSNMY3c2gkEitLbsAEz/sEtZt+VAfMkmLxVL7dAvDSl77E6iKoxv5TlM2CdT
wpSZbOzIKbi3Oa25kyKWo3cM2bqRWw6y1azQXYaDQdZ5xxshNtaBrGenyCQo27/CbU7Sp85WmUUx
bBgOyFaZetYBqNxV0m7t4vcmA2Xlc+1w104jETLIWToXDCd4mBZiry6otWXCJMwYJHgFDfdV7duw
0k0fxkqDOLdQLs+C8Hwy1t52pQCvQnkZiKnZ4W6tJ55QgXoPlaLNpb1lSAAxBrm700WsX8QoPkjz
HWgtG77xVL7odCAL2g5XYVu9PAp0odyMnu2Ipm0Fi0Z7RCa5RDi7Ro/p40KE7KCKWk64cpxspEVG
2kCckhKGyY2ng18n6jGUnixaLOCCk5zkMuzSc+UXEKRQJw71kQ/HAAzluPumJgznKDoZt2jXCvWc
STrPvrotxlnU1b3hMoPf5a7UGwS+Jsd0jmVO4d32BpYlmIPBV2FgwnvwNGI+zxstEFGO79zf+IsA
pBt5OItn11kr2plXL2evGvGkAT3BTyRXVFTElo86h0Qy1p25Zk4mKaPnOOhlM0RxzTj1QtHgQuGT
KPVzBGEbTzc0T2b1Q7YC7KwCiOSM9vNPSI8w40IaSZ8z9VDIrT76BB72ny5rIw2OJ0y5KqEu9zsj
4DLyZWNiHiOImQTEwE2XnxIm25tQMjGlzltJIcw09yBk0MZDpjBCfiCiAFscmonqW0BbgMle5yW0
Z4sRjPUL10bRSMbBTiURkXJZ2iFm/n8VnOJdZdyr3bj6GbOCy4wnm9wVLAYM2x+3pHmMUcosby4P
LQDB40fa3V8Co3G4NVKiwPDgAgJMkWpwVHjfPQtk460u6XdxkcrZeiVauTdVqj4YS3u/K38eyfvW
L3+aq9gJPIDpIaDBmbz0bZWPozxz/PKW4uGgK2JagGYhFlHh271qmkPg7stoQzijdEZbLqRLq5Mr
m4jpEbf49wk4BB5vEW0UVtUMFWG8dVOGFGn8YVPLjm4Iy6OXymzzaEji2C4Vu4T88+EgsM3/BE4T
YZbpI3Xi4/dbHY7IEdaUdv7mRY/e3stKGrWmeWrUg3DgZlGomUvtoJggObj2h69QD1HT2PQFsy58
MoZ9VyJBsdGeds2hiC5UM3H4mKJyR6SMdm+RVZpq0/RdqK6BX7IxVWdt9ZROSw/UQ4i+Rj3NbKX2
pQERNux3ttcBzd+v7ivQjboHoq2nh8YUmtzi+uIXzR+k6US8/VfOV4OQnCXCQQ84l1aXwTMSZE/l
U9KZNTF/WXKQr0tSgeD+DMmAvcXhHTHl0klWRO6zS+/iXyw+vSDpiJRXRVOEO5gcWBVtmaye9p42
Lc7Ukr/nUT+KExXfscrouLMtDF4GgScfhpLkSJnGvtxcNt69tks+hYPFa960zCNVkkfd5lhDVNW6
cWPUyONQIHG8tT8EcqntsTVE/+/6Xn1OSC1jGMQQERry1zs0KJh1ePPzu0hqhg1vp6t7AWuGueGz
TGXFUqUPXHfpiV6U8Qw1l6h4BzTQdLOlbhnA4Aj7CQG2spn0Q5WVJAirOGeNhC1FTSqZzCU8I0bq
7KBbVXHXMCw6Eenyj7Q7pwwhaYyo7JI2Yg67YLMUelwO4L5jlW9lPJyUH7215UoQLAsPL/BU66mQ
S3f6ngmv4qkx+nnBu/QrFLrtLaVqhgs4kox7fUCGYO4FrOV1kUuvNPf2BIx+6wQ2/+Km153Rjtxl
Kv5wmoTEK6Pwsk47Rrm2ijJY4xDbPF0/ThGaBy4mGH4tvtHGLv3SYesvWpDM7ZNi/Jq354Uk/kD3
zfyydWEh/sC1Zoa6mnMlMfT6JE/0Z7uX8JXRt1oEURKZh4jTe01tZa/6o8FX7XyZytpF1dupVdfP
b9JNaePHoYNJ6R3xfll3ffSem8grL+CTvKvnEq5q+ezLUNmwXQs4jbZBsd6k9rk9GxvlfRtdND+I
WfNY5dAo9PJdDSk5RC2XD1dWKa0DBC3oHdGZ2sudG3/w36YobTfMbVZQW7pkWg5KyYWOaP+WD/2D
hHyL69p5cvD9ErpiIUMajSHBBBRam/Lfq7T4bMBn/o0EAmlh//2PMZkCRmCFrWZ7OjJNhpS3Y1Le
gNCepuHyLydAQECESSx39VTHi41WC/iaJqOZ2JAPD0CFnXFaXwf/Z10TwSDYV6sJ0UOn6rYeCFXi
w0s3ZTx2Gusu6hehFI+W18DeHdXXEYAjI4wP2v0m6kq6zeNziBDvwoHrq/q9WY7z9WnHthXVC8zb
KMfR1w0kldvO8VRkHEHGRK6IYUxfnk7SalHV/iHcEgsFFmTm0kD0Pzq3rZQ6lYdhXEPbHuJeWFWw
80maLfyjFyGlDp3pq+Q6jTWuNyCglwjmtHeHLq1RIi13wYWUdXdCJWlkhUUkZiipoiKJE9vIZHcj
KSBOv03pTkHbDoAvgMYQKi2d83V0WIK9hN7ADHWAyhLMF/ruMiieuUliSGTjBXmiVJ75h9Ab99IJ
ZJpWfR+Z0fSgDz52Eyu+6+pmkvcIO7kguoPdRduqByqYu0GL7l78fetK0fpVq5MwK+hvUHXCA1bZ
4/C4Qhz2lXEoN6a44SM+6w5oHeZGK1OPj0CcFca67HPFMw3MVXvS60BvgfwO8FSsD9FMqqfSVkmX
IKTDFIc2aMzGeyInVAfwav3Q+VIBSmIQheiGUmXiQZypReylFtq3wzUI8aMrwU8O/dX8j3RgYmHr
SdJRJgxoYxktnx/Yb7ppCELpqUFapvAqEhun/YttjddKaPfFeveA1WUL3DPHIUmNR0eBLhVFq9HX
kQ2DWH4UBsQIe9Ks+dJFaGecLS7zfckt6t7h0yNgkrUHGedHM0hwRaeQSGfcEjS67eRpAJ0iDMOT
H4E6XEhtfN/qK8AgEBxYDEnAntRHGPTVb/sR4Y6Q2D3czONrxxbQ2/fWlDMxKg34zE+AmyX8NyRj
nU2XwsQvTU6xuq/KUY6zu63+xpcNjooUdpRzqg179gi7IVBGKPd92m7Z9h/pMUO1NT6e+r113g20
WehXG0OoKtS+P2EhYURVnzCUqXFm7HvKmCm7SICj6GMbOtEw/kEHWVmXPdoNxscD28K/tF2HXm0N
y/c7fCIIvbCYiU/WjJ0zAyS4POVDWevpSNtLAxhW+p2yJkyh1sUmS6Ld05u4m5bd0rvXqDPx3eDt
T3DVjKz9K1iRGKP2bwvDPYFagUFXHR6JpPhbKH7mVtwz5jRotgZK2nF1w6RZFvnDfcLeMjC/xysS
RpHkkN2/AxtD7apVPeviDvgd8jl+MXL+zm8kAVlUlgK2FuAFGOu73gImJZYTMGTBzr1vcy5ROzro
RJcLUsEl+MVJ3dExhfTVkQbYclB9lJO1uV01vG34vJXDUIG43K96YH3mwbI9i4u/67lCXP+4iwJR
wK6yEzOt3i5Sc6upMq+78zWVvbbqqScFhwohJjwBp0Ju2Eidi+IGCqG3KHEHWPaQqeJrZxsTBtoc
j+meRzs5uOM6Z3effHzyYCcFVlCsWOAhrMjAE61YdgSt+3PuOyQLeKE68hOyVG5dpwppnm3nyzZU
o7db8K6Nk4YcoUU8GrnuMRplTXcEw0eq9rpcvI6T3v4tgAiReuers7Bb0jyFQRJ5YmFfX171cPyB
e2KSmVNCTX/+nTQrBa5OcTLf/L8JQDsVr2P7m2I+ESovldhYjn/InubO3RLeGCb3us5TZsQ/hpFq
18Gb/IlPsg/i7yQsMPOhjuVxgwB16TflvZ7mS1EyFfUgABRB7qH+uj9usCWTGUQUfa8dYZtho6oK
jV7EsgFface53gTKjSc6s+Gp10+XuIMscEwiy9Qbbif9IjUjPEdRpt87B18Z+k4TgRsa6lFhTiZt
r3WLtJnQr7s+3BHp+BRINRIilGbL5oqByWJMMmTjKM5Hj8veE1C0OYUhdyufkdMMEhrlG5dHEKAf
pMKSLqhOUVW/r0cI38coQjwFnr0Q49HnfAPkiA4rjRs0SBMPKBLimVZ2QEJ+T0kFt4hhfQIMFV7V
9fOWHiZrYzdL9kY9arZK8Y7XxWyNmbE1ZI/cGz51zGVn3IFMF39dU7te+gIqL5DAm33cAwdzoLvR
42+6+/3TbdwiTkTbboePIjDnVDhMenTUsjWOoMMOcGnRusfnXmqnkSDQ0SxKUDuBr0C3H3jufkPW
88eBno8YeKIcE0K2mkhWVQB3xFE2Kea0s8VbEeXw219LcBc1rbCcVqULVHwyFqRalY9EK4fqExYo
W5qQ35VNJYcamwX5wwZJBl7DFAfUkqpaetNNKoW4LWBlIQ2uEhOWBSwq+IwYyVOfYRtP5Zdx33mR
PSTBQ7mqWd2YhG10ZM49GwUTSuvDgV2l9qm/lxjjnG/CVK5qjGzmJ/+xqW8yqV30YmyLDNi2v0Tj
vBeB1hzByHe9zckz5NEICjJjR8CcAGhBqyGYEMWV4tsYjiM/6N5hOuBbTQMMbT2I9dYFc1b/aofl
tIF52pTaT6gI1sHwZTpxaNtup+5W3LxFFSeE/BNaSWke9PsVVdFp8LkshA8QqWpSQxn3KbdMxsA3
FU0GZrb6zdZI9z9Gg4+CdM19jNYNpiKp2FW8bKnV6DSGmeBdp1BXhIMP7JIkW3zKHkNdQKHz9/uh
7J8GiSlloJBknIAKCMEepoFW2ekBdAvHs1ql2JrzylxsW/Q+0SzbhX/jDaVTKPlwQB9pIL4d0Th3
zWVZc2V/l5HryiVHRnFquiMv/l3yR7wNi1mvsGiF3NI2hsJZd1m7qaMtk9fcJUDyj+mLu8iLlRMb
tipKxE4CCg/1vZ0Jgrh2yxR010MF/cWG5LKgwp1vmDybWv05qvWe90/wACXlXgusAX33hstwCuVt
+M0Cg0n7wE1723V0FqPBddSyJCuTHlN38YMYL2gY9xGgAbJkHnf+S6uUHWeVznIkSc7CFaYaZmch
Qf8glUOxfDf98gLDe1+CdqJbokEJbnUxBBY8vRSECtANyf8AjQHv24jyf1YFYQw6OzifHpAn6dB5
u+EdoQIRinnz6z51wjaKkm02q1pLoZzbcNE9bEJX7x4+wVmyan5MGscMW/yNwoR2LlQArj0lvHJo
A4F/E+mj+KIQgmVrhUtrbzspvW+kr1GDnfMHV5qZr8Yu/3ZAUNo55+EP90AUaS/vt7c+2xBimWR9
0Rhm5UJxOGye6a6uHaa1+Uv0AdcRmHZwzA4vJ0j+tgOE86SqjF708sfivQcEnG4qJz/YaQpQDenW
QDnZ0puLILOrObVqZTKnu3frUmHKa0+1FBXTDQCZG92O48nNXc9loCAdqBkrM2e5ArDv5rVpjDPl
dSFdAa/ZcmvUfg7qEnfrlPnCSrBexrtI8OM996ZDbOb+i/pv3don8x0/FX1a7+ta0pjntWD2hJYp
ClhMkSsHgP6pFJC3G8tBV5OCv39Gp27vUkfyODDlwnLBABZyPGKdYuMuWkcmNMlZNKgG8Aiw5EdC
jd2Y3de9DxKtnQ3PCp4BaD/q294/LNrT3GYG2Dwz9DCFQIx/gACgTrcgM/IF6YH29ZvP4knGQaak
qQOWdJwB0E00SxMN4NUPkvq1i8HsIKrbvaIf1Q/Zs3u0SX71sQLf7Aej0g+WTv4/gXZ4qLkKj1Ym
UkfHdkLmi1Z4ghjAEj7oY6/7FMqA0LOxFbBaYdVRmoSWlOrPolqwp3e20CSWoYap+TudH/EgW9rr
f7VUmYcb4qOtZDHjiDX1b2KNE644xfWkEibBHutk0FVrCd2IbM5WD14GbqU+6rSx43YZNzsegN7Y
Chyb0qf4cA4mlaGonu3hOUF9Bm2bXK4lZylrMMPs4ULlz+rXuDLDIEU6qMI2IprjX8I157ySAoP2
ZkS6yO2IAqnCC0qmV8UJ57C8Amsx7U55XTesSR2SdBJb6N8OQVQ5/IuDJFAneYzCw72MTXEQCWhT
WQFIUR1sLgxPnR0FJQJK5ccVtjYErEPXrP8q58c7xMd0ql6p95yJt464xEbj9BTc5Nu5CYzmyWnX
SugjNsfJtCOUAVkUXn42FGt0i2DoYRxf4ZcTd9RwCn7zJB3s8I8TSDxerjZ8/hslL80OyuuLCgTe
X0j93AIIh3Gl6DwL8kPlooxkVd5Ch2M5JfRvtuLYxojYGbUTaxtaui4/laPx3+n/1HPab1FOqa3V
iuCWgXVhEtRaEcDiaIBNmyEi7bRJErQ9zq+sbG8PVgtHq+OsMv0mkUFqhNps0bOLG3l9jt+WBPAS
TaJkra7jNOjT1rB+nHEbuf1DstpeczlIOBUx6cTJT2QY3nedyRmYxiLEl6ZXxFUX0mmVx2ru0G2l
QPBC75+e4SiIHDlYpQ24w/NwRnl+Oj8y8Bx/G2fQzEaoq5+G9dsqmOimbmPdm8yx0TgfTZlgUGR7
zdCtXcugscZ6BrY7uNP6F9ksP+HerbkuQsWgcAzlU65vOTxkFfH3rWFyR6z7zckodlyefAl3lyvW
W2cheZAMkApVZv+Apo+0jTwZx0r0HYXtqrEijaiPNz7dgbzC5Qc0zNpz3UImxic2wPW5w+7duFvW
5HoArmEhabLv5bwupox0iZTNmQbz9KqljVE8S3MTt4db5sk76zkrS8StpDDIdY5QMp8f/BJvn7u1
WKh/uIGnbbM/nKZizpXREjmWBW5FlXXF8l2ZSFOiw3iw4/vCgKIeEbsW1lJjS4dbPDuUoWuQTSTG
wypk04Lp25GcI9JSHlPcagicjXuxJkVZKzJymqqn9WTLInialHLcXWGo2H0KjwnzGPz2MIYZcSqf
XurEWqLSL4afqgkyMYswZdZbiArW9G4/X6AMnOcQZeIGVoiTKz3zfoyTMEAU6HNelKIBSz30XvHM
iZzxgUDrpOCfJZjn4BQxuIKzOKdIB3ReWRBLyhRxCvL75n2MwJSvkg0TTv/3MJNa9cSaUpbJw/fm
4yeMyIfolkBDVWQZOY4yw6skAetlD9jZWjnBY471fmYqrrSzCTuHZuNKIEUUYhHtHWFAl3TI0LRh
DR9YWWfOu/mkQIU9yXxIK4z1aS8VRcDT9mLVN9KTpbM/0yqKGvlKY17BlK56SX+fxACVmTY/LyEF
ZMIh3THvO0S5JfQNDEzj4xtNDuvnpFMgbVz34F8EIAyK6/axCdD4sSS1whSfSH09nXm1vZtMGwtW
yMMHEHt5TH3cD5kPy/r9HcT4/NP67Zu4yesZprBxS9Y8wRibg7qWiuB+pzhWRYbT1/ubRGMDc8A8
Ii5zB6Sa4ueL81LuS1KRvwd7ENPyC0oklUCZEmVRJz4lsZRbrgM65e0TGBfgdabMom3y6bZxETgt
fFHM2ZTmy2Dz7oTg+GKyZgP1MhhGuTxvQ3J+WpBngAuc6L1BNXidR5dC3TbRSK0JxKg0HdlNf3t2
xA+GSrSOMnKs7UEodMYvY1/mHU5+dH5EYn4AmExcM/Bzu2gg8bqkpHLKP67SwzvH03vF9DIVtJrG
jUxuWzS5U69Jyv9G3Kb7KtkPc9APRRWe4KQ8KVg5eJC3hSSnFbW+SIuYhtaXw6q7YRVbMgRU3Fl+
50SPxULpuegI6NmGtpg6WHU5J4H8iYdyiOoXCb9hQFD0c+AloReuCSkDrdc8XFxNyvp7GINLmO8P
+9WeL9kcCT7lpgn2WElGDGMoPW60lN9kqPit5phLePk46nh2zkQv8iKhUGGWtumdQkx9D3U4gl9o
gPo+tukCeY+anpVIACSxpMYR+S6dEpUVSgkyChjuDy3Y39v51W+tZZCt/wXrQtJHvgRaywhCUnZd
sDerop7S0PSQvw91I5GgDnyI7sjcH9BiV0oxYeeLPgrl9saC8Sk9r6qMiF50oWXbpmwE3wlm1zx4
8SH3Aix1aiTBguJ73rZqpEj5q7eHhSMUP0c+E5WAhe3vwRW7Gsmg0W4ShxPvHeQwPeb0g/Uv7ygj
es9HT6q7Q70vlt0yWUxdNBhRbXtCjfoXHYr3ItkYX5A+mne4zfqQSupPGOCq7b285zkNzQpBO8J3
W5tN6PXByY8oBrWEgA6LtPTryCODIuahg3MDjGiNeczOVWkE0i1JPOKlwptuBJwK5UHKtyPilqol
im0R3b6h5w4k4PpS0SWGht2Q/BQbUyGylzbkrVHd4CMozeMJrDH6OEd7UIpojFZsNEjpolmN1XJy
7HSOeUCIidb8BzF0curInCvDNrF3vyX4gJlGe9TlHrtWiGnFlTCWh4e7ZIGgRzRoBUF73sZbOCDL
MWpDem0f90jm78k/d9vRFEWSCr6JtaK5pwvSnIHMIF8BgcHTomHQnpece+Z0oi8KuRcbLs4YK05Z
zE0RYQNLuTZEn2KrBzOayCAC3G/gYzgGWKcCYqxsZapHxLa8Szjtaju/tr6Ur7dZ7GOHmq75/8lm
VgqkocCJ89eeHA3IxTtvTTYBBm88L2+IASrHluoUW5EwAHeQf7V4yCVAUXPJrQbZ1MIlN+CIYjw2
KTsQjr76itg7gx3fS1tHpXKiKRoLVwWIpmVDKKTP2+L3TaI1BMz5iNmtg7TGtkIZdCvo/LtT4hoU
IYQcA95QFl6DoOQ8B8HZJosZKaN8L/LO80noqN3PghFXDYBfbGFpkC+hfS6m1LDVTxAv4zKyKt6E
semlOcYMwuXilOJjNIZbzif7+zbFyGbPnEmLl3mMP9qogP9TPy1PuQZMmZsebMxcEx/0OeAT7ykn
CPbfD6rPxjWNZ180dqeC84bEdVt7ZUMUQ8OEuBW2caqX725Likd543cI7dVYjrWRWgoCxwUdvQZI
ZM6tvaCpNJpuM5v+2ploYA8978y6aUshWXYjV053bqeCIlX83NgeFX2zUOOrGn508XgJCuPMr/JT
V/v5bTl/0XbQko+V4EEOFPn04WC9lGtShexA+tR30BJIm5zkbFT2qRVXkHGPbJlngtN1qEaWMQgZ
irJ7qJjj+W89nEwWCHEykhO1Vz3C2/lBSlCxZJRVEoh7OJUT/gbMvvqHqiG2dOFJhMqUneWPAg41
G/UzTeNqNg6VGwfPo9QEgBz3K0Xwo3RpmC9ot+ER1m4zq2CiiDYzACpi/aqZAJxgfoK1Y7yecW2P
cfCeriAthlyME9u3ztdFtYP6ykq2dXCp46HRrbAJaOr5c7atQ02BZg3SwZwj7BUSoZmYv7rHy7Fv
tx71thfAcPROsjlZq9nkqDABJVHVM6Z5eUZjVZwCPwS2Do6zmOxkQc0wr30guXKNACo5TrO8dX2D
ktbdxYLR07Y9KeTnUD965Siv2RhJ+JXkQJmdco5fYmU7HY9jH6/Q3f6KCxAWQmAtQO4QDiCuVWqK
ob4vvOka2BKDmukEY/Xr49OTvGUp58MiBsRW8/aY79JE7pybIiOYieGWZt+hYSOH5pRQ8OCRA63T
1sfNGuitrdnnP+n2ZqqeN2j8vaNToMghqvGSZ4vHGk9BgJr7mtAZIrifl8jF/+NG48mllkUEfWTH
mFoIOqpVIFX2XV4fuaGTomAMkYd4pg5VIAiOs8NTW8xFUN2x9iAuhxqc526IwyebOmHqLSU8sczx
OW4CxgpHdWtiqYbeX9UnRLpgYw/56VokYBv3cuTCTQo2XDKTf2x8wt5Wx69HvNY+EqNOuIQ2LFfu
eyjgl6C1YTslILI/xXKhwDdQ0uZCJhFQg48o0OV6f3wgbZ2xm74pClHHig81EkG4RJ1hIjSChudd
rksPCssix7nbiYBy/mEpj9R/isOh4oVqXbIJgN2OIdN3a651Wr1YJi26wsgz7dMKC6SCiChrGqHs
Qy6US8OFITmhHyUggI1vupw/f9chPqLB7Fvxd114clREPpXAbW3OJKETrTLJpJrSpNj8vCtGWgz6
rfXO3X1ot14mtBuhf7vimyyQcFNNM/esbIQtiiM1ButANyrR0uenPc1PK3DmoZf7mpZAvfmEnygq
ZmMIlEoMxf964oIBBs/PpqWL4LVgOSJnL6yAeWjfZzi6sHE/GdS/07rxKHvrp4PKioLHgJPathT7
P/QofZQ5LAitUKrDMflpeNjWuasoQakrq39qZ1MRRZ5gpKegW6KVCw0B78+u1tGguTFX3J7F/LcR
loqikGU47fndzbQuzqYnszxIPCCYU5rfeEImoLxM5wsKNp6cOHTgtePOteHA+l59CfjxS6x2qPMD
ypO+/1PcqYeP+oOh4taf6xxuTKah0QLx2xzGSfcfwMh8fhzO7F2+kqtxXGMwh7fpUmXfpJvFOuZH
TJaj3HNgOUf6/7YkhQQKcXl2T6yffY6x3YC7Fn+BqrFWln+I3PUcE7mrWB0nvvm5KfCCfog/eY8c
Ngm3m42tC8BR+urMQnJn0JeAnLvurVxywwaRoqKSmlBpz4JC81kRWUWrO1KDbCwaU5gDc6LIwFGZ
golvv+5WUiOE9ZwoAseIhhX0WE+KbmZeNSeUcj7rZRilDYP9Yih6Txe7W4H1Qh3KEg8Ya6c/5sS2
2SmDef0A3RP89ZBLFs08o3O56+tQFdd0l42cUr/spEE3H1tkQC/XNt4NMBgMHY4Mh2ZtNwwGtQvK
9OiZAI4F/YGG23WE9+v5hVNXqRtWyCfPLcg/gtIyMHUx7vNWWRynCOe8Bu4TsyXEUaueGun9qZG/
4bQ0/TDDUWnx9dzwI/eXmhpKYhuCAIOQ5Mp6k7ZG53DSNeMqRx61xkisArb+ceN3Y+gPEPzn+h0f
yxcElm0WVprZDSyq1235ZAzxXYg6Jj32ADtqzlPMovGYPin4hQIsZXWl4lx2Ss4TGKaSvd9/FR/q
IE62mEkEF9Nsfsd9XK8lNZT3NomHYSeICseFwwCOrWDyEY8hGah9oi2kVcOVhFO35jFmsFwQ1GRp
+GhfpCNfZlwS28PgPc5FzmNznS9aOcQDpUWCfjPGxYb9rfueO4aWTjxTtRiPInGPf9dO2a3raIkv
qcISGdB1qSlbXnWy6rFZYDnvr3dO8YooNxbSParYiUWSY33b92/rkPjKiQ9r1x3wWriQk+HijJpi
BZNPMhENKeDCv6euo1nOvqMU64k12B7vgsz5RYr5jJCYrjUn96r94vjZ8aBtRk5HdzuE2LJgBWv4
2k2NGqfjzzMwh1IwWLuHPWEaUmFdyNeBObqBcics7v35pcBnYWCCPbrcknrGU1HWxuXgY3fkp/05
gDhqVGE2IrPG76v2itzO6k4moghJ9h+w/Ft1Dz5d9ZEALU8W+APTGYZeF0SWxn7oYqi5mXBlqMYL
shjrHs8PqPkkGLjifWcGXj5cCFZhxEGqtB5kC0DtcGXC7Vz1Souoy50536QeoLBQR0OiEJQkxWET
NzFm27nJwPbhxBLzMC2aQiOuxwolWfhomRAaOU8Q6mnjUFXvepkAUl8psendD846fnaiKNISEcBR
sHs0x4s1c/vzaF6y1Swak9d1H7QmCLaDGkqnxMBO/m6OtRE9tVq2s6hBtJtwZwpsRvsq3zYjfNSg
8mCACyzTlWQ87o/2Q8BfaXkI1R8pw6BjEtiHG/Ub7+8kBBtYi/ZZbsKFkTtybiRMjutHLNDmUYgP
qs6UmHxuHqqVrl7HjzMyf3K8akAYFbz8O/VZn5Kp0EGTs4DYkajXh8cJ6D04jN85i1olL73iX0qb
ywoQ6NNzbrSCK48D15KbaB2NqlnlF3uG/UT05ZiE+E2t1Q4ASKph/rF2uyx/iFPnJ69wgYazOQQB
GnXM27KZcJG6jbgAZPK0FuyV7dWsHxdSQOMbABYK1KjARAGChAm/FtMVI8qjI+xaPUQuoCZiG3rP
VZ6adGTeBJ2E41tZQC6nsK9OOWJoq2FzdfzN+HR66SHAOGIg7T80esXRCEOg+uRZOdaHtXlEIFgL
z1aaFtMYoX/bbH6tBhFFHWL7SOMstYn6vJu3Y2Nm6UVy9ViCGDNUgUsJz9p1FdIst6qGeXe560bt
EzODgImiKKnUx3g1GwhD7lt1+K6ascjkaZMBhYr4++CUrOHe/UTjmhgz3646JMCb8lTg6HNv+6ne
+32fwHuGvRZuntLt+zD1tWYSNnCnuesffzbtEMF9KoV1h4DuqnvkULDZC9fotrqRWDzo/tNfCF3B
9qvoOwyeFFBiB+aMyTjp2VGsAzk6hZP4iEXWAKO/6G8ovjXthXKh1sNtsqj9tk6CaCfYx/4x7zVi
72CxAw/dZZdvPVSQReXahLmlwQHzGKq5H45+QSIjQlb5LaWssSXN1KTeRH7Wj/vnjFQEszrDimNp
W0M0BKFYbglUKWSVXrq5XKaKG3Z4uHGLAziur05sZeGcP6a2Y4N80LH5h/weTzqHPivBieokExhH
bMvFrWWShwTJLZ/Dv3iXDXHYDuvkjB2fyamJJeiKxgo/YEUhphOvT4Q0aklki66mjSW4UlB/kSvr
fXgEnnjQJdOTHyuawTSv901IGJw8UhxZdThSVIgRdtrfys7y+2knO7LZN0sld5+kbQJwyhT40uLG
177/hS3J5y2LFv08To9PghPgQMmHfLaRA6btID6I8ZCNgNuHLIGEPJyvBKTBaKmxM/66vw0SWHHJ
oo+HOGCLpb2h3D+YO4237U9MLOCE7gWaYVPsWGjlMYWYVcNZvPUwBSWLn/kLv0O6+7qCgEmTBILG
9G2Jsv9x4x1gvo0sVE1awgGDxZ9BWnuYomnr9/Oe7XF6VgMuspybT09nUTcAZzweSeMA2H+0SqWx
va0x+PoZ7bYaiI2753ro+buyyrdQ37rU7Pe2Z4znRlfd+N7wILFAYgkVK0X0eOHAPek+IbH+9CXP
9iokvC07UuRit8h0ZMjb/V03LO3B2E5OLE2P84PBa7ApQtyA3X50Yvy2reDpONHRgpMUZpm0pAL/
0hfTtnoLkzyRQ/FvZ2hAzpXZYkGKczL/GRLzibGQoFfK8I9LmoCUCUWPRZtYuL5jTP1KoUQWaL5x
8BrRMiZVPC06XCDGb2fB9gUtAqjjVtHQpDOvvabsL+jiEcpH+7lA4HSSYmGQypiGkl2J8tj6zRJn
8dMa3MAHPv0n7DcUKKrAI7B5A+TIW37FMrfcyZ/eQBFUB7UnYBVHQKCgpKV4bdrfW49yJBKsOLzc
DzrNYpqdxGmgwM+5sTePs34dELwG/dUPCdvoBfomzM+j3YvM3v8y4zWXWO8Ps+iT5HfR0vMtGi6l
Gx5ZH/VQtwALzeZQXndvV/qd2YWOgt6bIDke9ViHpCziXHutrjsv6l09JctLG1s/QCsS2QxSySCJ
jMee4cPOBMqb6Nb7QvZ9UEBCKu5lv6G/H56ZXRmU/Z+juBz8BqBDCrSFoF7vdpn1HV/JVA2UF+NR
JjmT7207API5ewN4Rvu9sKS5IhIvMGF5syvaH2WK+BVZT5nHJnkmNQHaJwNgZqeFmiBmlGKnJ6qJ
8katR+OgVAI39caCO4bSLjs+nmnSErKHz8E5Ib4vZQuSaPSuNyO+zIrdcXTlRBOUm5M6XtyujFvm
KIaPj+vcozRH3jj0fXYxpD2vR0qds5yrhoFjnhUPOROqhN/8C71XLFyAwUArW81JD1TYQcHga1xu
nO5kr0UbEDa8/SBd+AHurOfNJhkk9oR770GczNbClEfx6F0XYGQAu6w5o5uCkB8uBkbsOtPI519d
bLR7ZiVqW5brAgFsJQcKl9rokBSTuThBfHTFHxyWKa+9sDv43JzrCpJ3+KsICEyNwd+0xz24m3s3
/PQMIZCIxDZv6eCYU5k2c8c1kzDocuFo/jQNyd3mG0wkHSHQEDT+/xxlMQZIWCYYRxGD2NCeHTqv
R8BRFXecN7oomfdTRl0SzsclYxyaraob4BDXg3+/5I9FNW9RvF6djOObUbap2er2CZuGX6Be9SMj
/ZtuGbVt+ds2+0ZY9B50SsXRxFRnlbKfMZpS98tyxRf5p0JOyW9XWVfvih7dI4v8aR9+jEVxmfu4
CZRwXWp/BvqvQi0VI23KJGnSL0xikAWMEDQ+0/ObY3IzK5mJyYZkBTRdPIBWCUrOQolW6puUcb1B
20GvDkJvjrLW2Q8Oa0IMOOoa7+czfE7EoZsz5uSiLGH6kfhMxJwKG+IzvgURK2nk6QpJT1td91Z0
2IjXqJDmoRBTfuahmIH8u7WfYugmfn6Ong0Z7sjYjFn29hHiFeSruVJKeVxIOhVcd9T0yw1OJxkJ
T0jYamoB8F141V6PJOrCSJR/k5Qqb7vDObF+43vOn/WbCjO0lgcaXoj+RFcLY4hq7rJBW2DDEfbl
ASY1Cr9E/OJ0C/MR2kK2VdOjAMeMugfVTo2LgntuMn/JgA/HjyraZa2jjvAaj7rMG6CAepCkwUS8
FcELtFh3ZEVquvrCRTQK8bm0H+9OwXpnbPn7Wpk4Bbo+blSRLd/UY/y/70/VVni11kI8mtKDXtmo
d7C96J3SQjrMClBU3OstzIZeCGlSIW1oi59difkbEl3YdAt6xbd2zR4jkIGrMWkvcllOZZh3yhCd
R1ZXhmFqQIP6t76OvjQmIfCt6s7iLxY1q9yJDM7VCt5Hk0gbqDHuMIdnS1PcZFyI/xOUqsL3xuv4
f93bbYQowzBDSIsjnXgyV+bH0EzAigEjXNndMylrpwcQdZ6UZtShhmCOvQcDGZPrcYKkW0T5kgUy
LNIUt++IdugicsBCye74n7dExyeYJqETKMCUFri2sYuTjQHLl/fNZEENiSDQoWkz+12WWYGaTSuo
rndRYaIqBqJUER3hlIQ2aDVnn86EKTscxgzuShexMGwtPPwidaXqQok45ojA2uUg+MP0WHDT9adc
z5B8RnjDAKcd0nQtlomkWrmrLH5RABtFRiJBK+yJI2YugtuXc0zx68TyUMldQ63fP3DZCQ9V2Rye
+B3kMOl3dbgjRb81tJw/KkBMGYsf32GZqyVPbtS36T8dInPgNmaWTqYQrBe0P8/s7+SOU/a8py1I
pDjej+xzXfxBFZ2JjE/u2n0ALacDO+nvYRVOD6YBh96RX3bG5WfSVgS/aXH+yHGGbgwm30vXZOg4
b0wGkfl7gJ9pT43q1ztW08L8cFZTm/DWj/l4QveWjLdh2MVfvhkg8WTn2KfNExwFW/WGpZx1jeMU
67NWDQm0UBszDgWlzHKuuZxCGU6AEfZMSF/DSoCWhb/C21Ki+aL4dXsDd6quljeWjitkjcWTzA0d
UkQF0BiezymmKouputnI9VBFFDOG/NHHqg2FHhljH8UxOKB+/LrwfW7BgDZA3lmiOto82Fzl1NDO
xZLGFNi2QXYQi4Lp0DHHEvT8FRakjwdq2py/dUBu6/bQQ1zLqi7SglkK+MIRuGqDISmF4k67M0C8
k945I3uavehnBjBdCRxjnxHvLb8t4XtKYNtgZUNgQUSo9/Pp4Ljqo6rWiN4ScZEksWc1UxZHEKhO
CjxFEwy5VTjvH7MpnDOu9mGDf5Rzkgft2FGkpNZN9dc9YVH0IjPmESvsMguliHRR/VgxnVnGCnB/
UENrjHGzXzNcw4XBUPWR6RDVCLT2twCKIdrMqU43/tKms4ZHPfJ0IoUQ1dHsvxhmRLoS25bQqEp+
SGIQNW6LNdfwXDEaVditp3xi8JoV9stK6zCSqfmiXkgsZhATc0+LZpVQefQ/q9pb/T+/vsdw6w9+
LawtjfMw/xQMRbrFrxTYRDkEXioR7JkR2ie8rTYQ3NZwRuMwIUmFH8Hs5XIFf90zS3vUJTXfSWc6
FOX4n44IDXQxZsq2SboMPYWEhFdhEo8R7odRfnikNlReVASIqlCTumswl2d70jKU/9Yx1fzJTmov
aXAPZmmOzKSrm1QvEkQmMjTn/g8q6QSrlcR/268I37XEleqjgF08ZL9NXGZFANNOZMOOcSgFUmcw
BbsBazWZbah9xtCZY6jLqvqojUEhW2gazZegasfVijY3A52hZNcfcAbyzzZi7Rhp5DsGJcTaOdVe
7G/WqcgNAk9go3RpC3vDffuqJ1FJSWYrCizr9p4t+N1I70HCZ0SaUos5oae/AP32oUnAYswIVQX7
2pqDVZ2RS7Whw1WSiq5K2oCpA20h3SnZ/b1cR6xShg5hM9q4f4PQcMIrnvnzbR1SWpFVB+533STH
1nw3qkZ8SloE5Hz2CYyteI3je/IQey2mkgu1nRryMgdIPJrIBoxAG5fe0SHIkCKm9mgy2VH/0LGd
xq6K1sdA7LuNh9wTjUNvvNZ4eeX8m1cn6uanGYoc0RamFz9mrQfjL3k2FlN/DIP0Pv7i2Pj8fh7k
55RvAW65IYo9S82to3rjqBlAB4jH967guUN+5R2uQ7MXG1mJEw5DVrsQlFLY1N/F3VF3ILPuEi3C
L2anOxZMRC6avnyjRXRiuYU4meQNjFSR1qL1nMWDdAua1d6k7kRD51GuXKrExxxTryy+uo0Fve6V
9u4vw1/2svo7OuES2cqxnkSyw38wG/Drl5ddowIl3WJqdoMwY1i4jbun6aMs/7Ny7iLyj/aPFGRi
lVCrNaoS/yKXiGuLnjOQoK6l2bO4UhVn0JttNCqsTaxUr14fl51ftJwGfR8Xd3FNiRx333WiVYjE
J9n3tNJsvocTIclbhixjIPl6V3XtFypS1V1f9rluNDN1NRB1PMu315SqB7+ubqi493Cuac4XKPKv
q2ocjlnOHk7RsZo8sAVDdmfbPh1veuVq5f8cHLQHQOOANs/ZL9rVJmJHV6QzpV4gwUU0CFTLdOiG
l3anQ/bBSZMURjhwAQoZ+4RI3vRGKvkhKnEuIWtSO0NNV8RK/p1WUtHUTvLBrO/+JkdxZshxySHd
MPA0d1WIefs99CJLyjPV7ts9dnCl6L9cKaRNiv2j8kI5ND682IT2x16LhWv98Pv5Er2AGRqFKkw6
d5etN63MYHriXiI3yJk3s5JHCWGBYu/FcjWLm9RP7Fd/g1P7BwZyKwfxcl/Xn3A4hMg/e7eZiqtd
ViX/fNTdAubHwI57dLzEx9vOwuU/TbX6+2G14ZnfE0Gl9LcSc6rzEFLLW2xgL15IXpubf2ZqaiXW
5k9sqaBztZNP/0UHuX7rpyRIwXRQ1cwOJgnItoPQ5pfMXuT6R2v/0OHmZjW46qhZEf9fv+/sz9QM
QBe4wiKlB4pvoNDh8uZ51K11Xj2S3jHvEYWlNj9KlygXNj1etsBP/kW7QwPzjYRMo2kf/eoNs3hw
BTllpjLiEDQA7DwwgBU3dN75yQVmE7paBh+IQSiltqEikpJSsxA9trhBSSc9S4NvhR+cDRGAE6HV
7XCqmhg07Al5gODvJrsEgofNT8Mhn/fUN3wATl+uG/URPJcOLQRTwg7uiyoDi+8fbo0CrMhbVlLe
e7N4Ap4DHQr6FBL7jNFxELDC8hVWRlYv27r5YlK24pT2vg+ggK1PpE0dUGUfxkJLuv+NH9+mnJxR
C7HFDJpJTxq3Va0/0azQoC0EOaZav7fsvNVxNKEsqyYWXNfj6tbgzlr2B6wyaodWwvWk3RvsXXvd
C2PSKrgZ/+jRx8HRB50+/KBgm14qJXI0XKWCrOYvnzqoNCmNfYc1uNEUbzFtmX0UshWF9fqraXh6
UFHGeYDz1Y2pvMQ8UVNxkRgFvdOF+UV3caqMIDRmzbNjw2hhyFOelmSGWGB3vyec4l9ov8xEYWl6
MlE3Ukbk9fLU4uFSGn9c33tEg679xuHqxMvJ/a66vYjqwOhxbnTR992w8CgrVmRXHMM3SwPUNb05
9O22kTYAr4rt15WCCW+147dyan3aoSem666V7Pt3CKMPOsdJcmGDwZJ6DyTwcUn2bjQwhKSXPbQD
iRxv4xmPnwbu/onjKJ9YZkXxJRhw5UBn6U+d3foanYp5W6q0u7n9KKAcGn5QpvlKMLzdt9EBf1QQ
8yorckBaUsIT8uf7667dI/s4gGLlpif8/4qF41C0oNkUXf6Qe3MhFV/1XVNJ1+oj/9hwFvu/v2qe
WQzw4OukKtDB/lo6Kipi8iRDUt4t2fEY5Tk26Da+FJ9DROzBVL1xUYbWLoxRd0W7Zjkc0xPpaXL2
SloxQe1RgCIqcVPE7ieVMsvKZ/IwiOjJi6siy6QxKhpM0wKDGu6vXjfjI8yJXzB/pwyV9GmHBySD
YEV/LoCCAfANGuIay3CUEQ5HU4uKwLPXNrQv80xVI4l3BHC5pAsSYeZB/U2YLEQsRAbty03fV1HQ
npmazWRGLmpt+BFSbXywLP/HNuYKRdbAP0U36b43kJheArVO223pIOUXxVRAY+m4Oz72hOvpG3op
QjNHMfNViEUmFUFC93o9SqC43jWv2kxb0LVnKUlDK3TN9HBvLlK8z0fkoPVw77k9BdUZ6/u5R/yI
tRW79zM3OyKx6mGkZswiAlr6j6tJYnEYRZNRSAyU/v/MZvT6PDC5q30o+HkwUcM78s8o0uxMBEWI
FuJnK6SofrYmESEncRsP0S63KlGSBVisx87IO5xR1OYRuxvm5DGkYhNQPev3S+dVKNcymVamziv4
JqlgkQvZL0/1ee0TW1ZdbuaQohpiTP3tyx4wbFHjoV2mZA8IBib56XefJ88x1SC/q5k7z8JWjrDv
8cJMX6//3HbajknXAUSMBOgjIFOxVJOGWW0Vsq+QMGWvTylfq6xKiaCNc57HdIGJ0+6QDq9H8QnR
pFP8rKtqJHrMdY/PDftJf+pRCIvUNyGrTuxT/HrXnKCMoaSQemKJi1ShpEO9crA1Udrnpa6RYlO9
ByNFAkoFlFWzbvfu8bDnV/5kqqkWGX3x5pLd+fAd8jae6t9XlQafA3GPV7iiR0pM+eGKfUhve5Fr
PPdfledsW6FbWHOqCTovcH63EplGiL4XkYM9YQAKLhz8jgobwsgnrBFPlW4qlB/f+7IEVhWVCa3c
Ay5A4pocR7J/h6uhpQz5FchMDos/3P8NKPiAMWgwKKK4YWVy2nJ5v/rOHmNNAfa+tTQSSaVW5ZkP
1ZF87+dz27V6w8Gm6rutCa2b50RG3CExl1Ev3iWYLqnIhBe/1Thpn5UBfkT84GTBxMiz19hKNBSi
yCnvXdpo62azepTzS8gMnc21h69E0uIFnsCQsOhNsq2301EOV35cC+jsh2lSFtw6AStIzhI+0nlt
Np0b55l0toyEo03UOvNssgKQahm2e7g/e71ux4C0LF1IoCqoTzA6M9+EsiUEKG3q4Z3pPKqFhACr
0HtP1v8JSBnw6kbCh7GXCBAQO6l+mo43opdbfAAKtxRzJz62pDIU4AM5k3GtXZZcWYqfk1XDOL1F
RPaONYaYyfsLsApJ5ZkLxqDYEivY/lgf9o1CKxhwHIeRuawQfHxeXLWKMy3iH/2Fka9rCD9IOQoI
6HHl/Kx4jVryCndhl3vPSnhn7scEap1ONATCSAatFNXn4+8rfOojbXiiAzNj/G0JtgEvWgi68+i4
i9FUa6LmJi8+5WmM2ugZDUv4Ok5lA3UMO5dfOs36ugU5kdLoveTcUSYiyQei4SL+JYpdhGPERMZJ
3+vVGljF61C7u2bJ80T+sKzE3ZKy7X26hHvVj3yVtJUUIh+uyUV49Ugd9SJNSWMJXlzmtMTzgT4w
Y3DVtyU12EVGSi4H+vC9lX7o3L0kcv1G/nx17G8yHguKZYmDKpVrQdOHEhLSSmM7xXtRWzeE3UKg
037E2SELDTKz/2VjamX2ZPhpOt49O1XEECxcmuagThPS51F4KCqBYy0FSHkqDiHggeci1g4oD8aJ
qvRnVWzruxBucOpKyZHU6R6dEEoO2e6ZF8A1KCsy7AUT/NPjb+fLBIfPolSHhKRWSTsSm0SsZZjt
z0BvreV3CmXyj16lFhqOIrdFchp4KboMmrBmkzdLYh19TEy3BTfFkZ4TZ3OddAJOL0xfXymhr3Yo
7B6apEmU8d+1Of8lOZfuDAJrp196LzK58BeREyNuZaLEQnYRj8xTkkOCUbxV/934ifwE3lpBkr3m
nLLJE9m4VzkfcSOdgb80l3Wm613ow4rW84RdkOeRu0sOuogoONXcTVZBmoZ9I4TMy5Yzo7CH2UmL
zF6BILdrQPD8jl64PxxC7Z651L5hRn8BSBGZmvJOGR4Exl0Dm+SJUOw/jr+EUDxy3GRPnPSwh+/G
2s/1gyxQcUI0p5MmeqUF+k7vkjMtBWTCZvPj3HyB3cB+9awmsWA30dZEOkPCALU1SNmkUcvUBcAd
QvSJqRNpNv4l5QCNaUc1vSf3UUS8jrFbAI8/dACj1Qa+lHskiAWsXyblwZ57cBREhrGXoVgtN0Bw
ODGXLzabrskani6STBllJ1y+FV8KsbVCbgR+CfLTc1okuycU8Y9XY5qogLyk0AkFDI+sFUbKBbVc
M3kTQ70+LmV1bAvcgR0/jeBofiWaB94mk2uyA9kEw2layrAxtzFwFNZhEpun0/IATdjDM0jEJN+J
RptmuNOocKmERNs1vfxjGSf8l/o6G9WHtbC3q3I0v5wkFTEDx3giMQe90zQJfF9DUdThNjl0fsu1
332WPTxBZ0YKn+h14z4PppamX+lhoG+/NH1avJ3YPIA/vitakZf/C51engKHbcYCwKntZLuO/pGS
tsAxSj5cnlSl4pWJQLqD2xM2Ho3ucd/SOfWkvIr2VAhTr+dGMgsgpXHqsqNpzQwmZlgSqtUFfCJO
FHE5sbF9L+EZKlneM7KpNjWxV0MsFgOa5GP8aL283Dy8t6D3osULSKU8/ZFaegNPxk0QtSokvkon
ybTUnEkZWEEYa+7vo5GmwsvwdGgjhYxI7Uk3BX+s1Etp30lw5lMXWaqgT4od2tXrspA0wLVIwdHh
gqUhOIDbnEBlRSb24Ea7KNHjQ5P+liOA3q0uSulMsO/tEzlukZBg7ZaIhqzZXRq3a7FebWDDb0/b
FRsGs/5WuMHJP2pt9PRri1j08ZPYY8tYtrEF7JzZXrfA2xY93zHR3Z0+CbDM7JkKYFA6j8l5iwB/
n0y20AW/vSGyI2dBoKindjSS9fSMKfgFyIeLcny/9vEXhS/Y/rB52qYRP7++ZWy3ZZ16Slq04El3
VzhjNTFk12hn5mb26MLtNZ657RUFcs5qRVpd3GWvq709hg/coDH0gWfctVMcU3tR96ftwHvSypKc
00LHdw6AlB2ZYnA8zQ0xjq6iaVTclphVFLAhl41VyCw9hauF3oHcjmU+zmXfYMNM3WOe+fChFit2
Lu9XjQDWN/MC2Q0iaf5nH8nkuDjyxOy/kcDVbnZmf4Gy3tAsVVMSbL/4AgHq2BLNFalwN5LFyiyv
OTm5sxLndMxn43d+B3z3oX/8XTzJmoxqYQ3FBlxJfY5OHbeozlTw81CLxb81gZROI+aXouvvQZSN
tYPuvn25FzWtgO9t7tjvPYS/EuCFci7Vt7i5Pz32EMny/CjxrtpzQJ0gIPqcO7J6U74yRcvZdiQV
Kxoa/uQ500WNCNqv0Qoq4JGrRJW283hKA9SJN1+XHMy/0ajtLsuA57JpfP9Lmfe9/1h/mftMSrtE
19QIYeDbqHC1cZCda9fIgmxN1fvD5+0iJi7UOdSqj0cHutCOfi0U1ZhuA1E2g1+CGvmnHrgUUcTa
LrWh+ZRjGnc1ICewpwR01CE1eLwhneyb2Tiam4cF3vPtvvhnaIzTQg760XsfazldgY8ThjDabMD+
VEt1SLvrUcQbeXhxjW31rfn4+krSqrJCASYmBnetXz7uxnBSA+2JmnbRnkn3hwa5oWTk52KHc/nS
z9r9ECIirv23Ee+b9xkTMIY2LrIzMxKYbgrtsw/jfu3mTaEg61eKguNNH3gnUSm7qJuNHz1CLg64
jQssI2WWFye/hjZhJnYUzB5tUuidaBZi5Sk9zmU8ypsqPpY2BktWVIlUPjUlD+zxFx70timBByQS
FbKA11iMwjArUqqPMPYYWeXbZhTtYaR6qDihTBIEu5srpEMMAzDuDD9YfJsDz7BX/6EqyDHZfbQn
OPsi8fc1aJsEgneULL2W7iFFjJmxc7iRAb06O7zKlWOapUqr5u67TNpW9vcdRJgX1AUY6bFnIv3t
WfKVOetXQbagF8yxcu7NI6YypsL9IxcD86bAj7w9a3r1keDawCFXJ+W2bWuO2/nVcShQPYe1li94
bfpLET+NQysnnDmwKbJ314VXMGbrIosnOAfiXRFZjBWFEQNAKGodFy+DawILdA8/M5oHooqHn5ny
0YCnpokR26inXiHJCrKJ6QLB9pERKpmwJ+4bsd8CNADlTAhW6VKARQjt1e5dfDrJu0KElCCcorlA
ozHx+RXZUyxHqEqJhW3Sw+CbEhx31MwtdtwdpwTLkQpYCrg06KRq+jp8HjP+6Ik3FciwbdarbsIP
oF1TduaeTkBFArTrS2LXzHBj52jXBYRgZN5T57eNqKHx/3tRCMV70j6/a/4w9u6DUn2OLI9Y1QWw
+byjMPzLlTO7Uzmd+H068DVcB9x7g4Gb8A1ei839C3IWck9dH+/kgDuT/6aeuWm90WhwM4WR4NIg
VVKWXoj9aN02PXxB1iA5xqAl977bK8DixPOTIp1Bb5AEoiiAaj1AD8txtFaTa37oYi2ieUDpm6gn
pcgXoxs8XrPhzIiYEAxR8rZdQ+a1sPuXO8E64I26VxqQPG9LE4kJja8fz4XcNG6llh9xTWyvsvwv
OsxFK1UXR3sfB/IKHFH+1TAfetOxUxXWmoXR4bMfu7uPDHP+PUu4CdjUNlOikCe0gGdGqIB96dcV
2vH2GnkPeuB07CpjAycHVmKSEC0fJ+T1rbH90q8lpOTnHxDYRP0zmVsQXNSt/DXB1DQEy9Cux2Nx
LxfUJ/CcBfb7N5KLgklFg2+H+D0so4HN0rvPdIym67zzsdQWX404UJW4Qlwt/sZMvyppUQ+32EkL
s9YAmjwLG4m165ezhox8A+aMx/9BdPnUW7kTYG8FZZ/mx5DSuGNlvNnN2KxK5j+KiwhY6Xg2BCNI
LOM9au3g01CrWcWn3O5xAlDJAspRWacRbCP+kPqRo/6DYIfF8/h96tUrAGtopyPp0+vsz9+OR97T
DGpRd9/CfpNOwLGaBQo6DBIlKMA3LI7l2ogk96DlWhmoKFdBBOdCm19MYwGRpzl7svcHGEiFnW35
rA+hJaiUypSc6Nw5If9f88GXsbiJmYeus2+gfkafzWf9ZnvhMMh58mRmliu2AsttF4AaHsWSFe1A
ddFAzsgyfgW8/mJV4mnabDSNrlsXGok1FBmD+aJWPA/haVWmjv9dM0oz9vnwUjHhv6ASkL/ve7Vw
2WElYrxZIEYRTFizElAAp3DhyWVXOnrsizm4FLUIfgyROTqv6S+xgypUWbWhWPwIQZSF3ZfUesdF
WRw7Ke8/j3/kfmKbBo9+xWjJsgel4zXSArtLFPH3Cq2v7eHDMYq9719zfQd7ORnYoRI5Wo9Fl5R7
/QqeGsGqxbNBkdUiy6DhNEZmtVrnP11FBLkC5Rk/uCc0ULESd1lGt0oQi+Oh7obwavbemc5OkRHy
qQmMG0Nt6KAvNQnSISKevlpiDQj/eDFOoKAiUlc0lwVSJJovRSi4zmmS68JuN5mXEjKaR6a40FYu
Cy+VN0MRCyq1M2aAiqMsjjCd2hdxCXxfSiDVQthwLUSK6UfqrDllTwcVCizWUZta8ruA5wR32Wgd
iMxJSIcqHKTp3ooqWQg+bWFsGs6uESPagk1uiMEjSkmSYEbNDHP5EuvA4MT2IMCVZidtCokyIcjA
/hS3Pij+xb+jDm4nR97eFeSGv0ztFgXih3t7+9rt2Yggfy23qpFR6iRjc1N8UnxdnPCkUdOXsNp/
MW87OPu0WN/PGgy+yCjtbuKCgyKvvqLq6l2ne0G82gbSlmwvBXRAG6Jzj/oiUfNOT7iMx7GvT7JE
5oJ/uswlDM8VGPi6SZzpkEy+VCX1PUtaJ+LyoBP9lmk+jcVN2vafi1XvbMFVaP6DN+vTropmhh4C
j4qAegNFOPsNgpybIPkzhHdnK6zx+KgRmDFVtF/llCx4a5ch1F9vRTo5PWOMzxRAaqyp+BRHibPL
EInBD6BFOqSymY5AX9Sv+fUS51BhR39KuzXLObFwW/0Yh7p5y9ywJ1snxDLrVki2dTlBYtJc2fKn
deZmYHWQqcmrKWT8Qom+bmm9wrH7b2cIsGgoH2kzg5NurcVM72w40Pw3WtOTHP6wBviXkS9NJ4zq
1ApIunOtCvs2HY0xTTWbgNU7YTDJ3ZgIIII+rXwxzVNbLfnOOs43NPGTpViAMpSqryCFKN0gyBgo
/P2+s7Zh4OO2HtseFakLCd5cn1NoeqEwGWqmSJDoT+BDC55fRSHuoJ4tnzR+lyLFPkniqRTrMhXs
5MrZ1D4NTRwKBrFTj6WQ40i+eKrpbSUxQJ9HB5OhFxbhVkFK6Fp8iLdfNbai1z29WbQ9ECXWWDc6
6dYw/dGOiAi2aG5dLc5xFRbG/KpJckf9W9jjjiaUgQXOxFxzqOr9tUNWFij5Cb1pA0pk6vbFkHti
ooXPM2vKCnn9WhmepcSuWKX2A74TzIA/PUoDp6Lwo6Fdg/QYFAaMHx9c+5bGX7tqcW6kdGfhwU3W
eJkbXphmTnZ/qr1eOEDyid1IUY1HrNezLfSdSUPD5KIq7iUXvlPniwHrf2v7UPKi90qYAGS7CFo/
i6vEowtSyhYyXisxbRQMirxZRYqiUcOnVz6qGMiFsA8djgS14vrUzNwmX1AnRu9+iahMizL+PeWa
X+DYA1UI5KTCT46NwiEqhj4aPWWsZOphm3Gf7OdlisV5+9HHMWMfKHvXFYYUptFpoNjjJk03FWbc
NkYR4nlhdZJ+0emp+LPmTlAt6h0pKiW7hNKbspFY9NQF2+Hn2ELl79YavIoynqGimK00/8bAIghN
33TO+UvACxgaIzSfj5atpzFCpXZzexRHHacMcho+Bzl4szeWEnMsGiXmpnNYDRgIvsK5QRDcmEPi
Gv3BFyYbbDAg504eVDtJt57u0kgN8jwR48gbAT4Brd3yJp2O4NLRzm0i4MtgF5x4AGc2fdq0vsRC
2um7dMLpsfIhJReyJQngdmuSXavtWNVoAed8WXsI66IkbNCNxVouwWz8WfeKVFfMg+TLNyY8RVf3
iZRnZbgC8jln1YzLvk+jYakgjLUU8FV8LiMNaxnG5HbPYAXgSV0D96vcVZZLKRsgel8KX1DLXt99
FXEpc/kOvFPHmcN+alXjbXQB4kkKUcQaQOwLYkcgUGcywG2xsj+ly7MVePNKeI17EFjaoLhDJbGP
WM5SlJgDHUFotjORONlrLmf4tR8ZXlP4gA0u8xyatbaXTc4015fsIOumc29J+9zS1yMmzkHvHmgW
4Ri/GHIk9pWWdItVrTNuIxNKkcaryJOeKIxHslcjIG3tC+YOe6TJZQNNy+KA9MQ/cJB4BW7Xc0xq
J0UZhn0na02H7hHYKuO5072naqY44ZB8WJns4i40f0FeSfHU1rLFaSVtEB1pAsOsu6Ip2wYaNNdX
nhPgCtGScQaqWx6hDeSVnzjI4Z3fmBpTyk+9LLqSeFV8lGL73mnL5TuPgRq2Wbmn2YXqr0vswDL5
nMXcTs7J3NiHyRosYCHZ7ULZK3XX64L4sBeJapi6hsm+Oibt8B1cy7wBvCTJAMSo8Pf6P2eHDBTC
/wM2n2h+KFV3NOGIhA0wrfyTedBySgtL8uungUuJr0zZl9sIaTd8bU64qhdPfGDDWz7ceKtgVy5g
81PeyhFDDLXNt14wP1b1K+Se6fKRbO1y2yk4r7Z6kKLes0N+qAl394gyMLQN6onhMGei+LEgDdxV
4jY+SpuuIBZXRZ3VlcJSYftVJPjNNTWHz5xLsuTmOn9VLg0KPIaNafeSlQ0vvEICeEPygKFiluoA
Zx3lDFFj2JCV0oP7WyX1N8jL4rf7nqj6Fxclq11gfuWoTdnmgjC2H5wxEuim9UMvk4pY66NNTcTI
+RmhCLsbmlEp2pi7g08cMa58kNuwyoPwOT+8W/oSa+gJNBYBFsJK/gscUC+D+yIETN3hdOuKC97A
+44GlcOqk5LhbnB/9QHbaDQJqvfQyRLeD7sYG5djW4MsWlhDbqmbtf5G8cis5zS0LrEf0HyP421f
/DLf0wSIcsc8kQBg+NR0RTvZc8vAZxXYdR3m+nblpflv7rtkk6KsXzJ6/6UuhfcEOUEuLfn5Q7bD
Z3E7KefllE93knAQFhRHF9xq+11B51TgXKZolo3/hDDQ7supI+aqQscf8AbPOYPEmZN7AQd/gjeh
a/BcmKqYdGAGEC5i09Mw8eOma5bWFDrvStBgan2JisKghpxv5dgjCXTHu3kQYNpwkbQ2Audx9+oK
kI2DkA6TwuKPeBTcn/mYm9OZRLGxLXMcgq+TF24SeWr7/6pRKTqqTwOsJkO9Jwvz/obicOKwYGxN
5MC9arJBrWLDCoAEKFUni7+gfSHi8X8VDRVjaUKSefnk1RTkDM+Jf/wu1RfRm/fUeVDBrG87OoXg
vRaomFt9fr+BOxYzEK+Y9eX/MJsdP2fC/u8bfWfBeUIvtu37zfv/opkzL2QuqPuqGV/qjtK16bCb
w1U4eXhO5OCyLH0dlJGmg4sjLlhKM0pu/TWdtIgqUNc/H277AdHzz4xaz+neZBfxw8xS4qJsgzfG
88wh7WFz7EveHqxYX4Nowp+s0sQ6dQIVyRKh90ige9QFSEPXkLv04wjthhQY1AMRJ7PZVT9Odcwn
tWqOo84ptxbmrsZh90dDSBRZ11j24CPf9OL7RmPUtxj7OxZ1zVAqCdD50ATNHTGXxZ7BfFY69VLa
c+++Odq2a2GKfZkQp4Lvj7ReJVXtBfeZ0VQa+u0e1GmyG61gUJcfRutoHD0cOCSitTJxnZNNyO0k
Q8J9V1yIID3B96RRpm0Ga2ib9vZMSn5jlC4Wf0ineElivAviN46ybkO3fD5Kz1dcCFst2CIqDFmy
a7Lr0cdTWy3x0SDOVa/e44mIUTM8XCN5/RCOEPiiY3DiKhFAYRTeE9LdSle0lRRauiTT7RlJ7bVd
3lrp7ihBIr8P2nYtUyjIZfXLTrYFGimWmcokxb4/UbP0IZ3vazfyG3hRxyCqRhzJsnNMd1oHQQDU
Y8XTZ638DEfBwiNqqcTsJcW0xPK2d25PKbu+24YzHgOoSNuIFt9zbUV6bMrroOG8OZIv8OvQczMw
N6pWc3UJm5QJtQLJ90p8A3bhVr+pjCGjrUBxjuV+6d8JaoSEnVUWcdC3jvyzLe0hV105VTMEK/qf
F8/Ob7Bg6dAQacU4GDowTACSV5Sqag9QPpjk/jXXFQIxyfFWtw0l9gMYQ4zFUt+AvYxs1UuBdc5w
DJLjEyjlJH4aN6HVL5UUYbYifDc187SaHPOX9usex8/4EPnCgNs5qfMpiSJ1DjAguluJe3rEy+NA
2pv4PWvd4y+4GWHqd7MoC2qdNgO85xknnqzsKK3raF+7hH6nWtPE7+mSvjtWkrGk2IssKosimVPK
biOWzqCjByT9AT2320xNckc+ybnw5Og65QTFZZxTZKjZ0jZVB334fbcL+VIFrZK1TuWuhM/0PGOI
yBpG1pXaeVX7zIgw/BXVAe0/mYOa8bEthruWj6fYeaZeiZkUR2elqnwOtfOBk2oht0/NEdlmAFfw
uBWRM7TfXq6IEJpHvYA5r2JPYnAoLWhlutN9of2aA2EnW2o9EfAL30WTrPy7y288zwtXbATugmXL
1GGnBOjOxKpl56ijTjh205+2/fbf3DA+LmO2TT9jLghwUUX5dd219TyuLzqKtbSQ6Ep2bKY7HVVA
HH5qYEizmH1wl+0d5a9rf43C7pOuwFjP18u4nqkP4V1WoxTfHt0B7eIdVCgdRmoc29x1+G9KGnOz
jbCBrSTnsFc8ELWnFdPaNE1aWpkYpbmOxsPIz34kNokdxMN0+vp/LEcOACvB0a9aAxriKhtMgcPl
OXAgoM666lNyzWe7RLHIKRN2UBhsWov5LWa0vrckvnydNXiBEZDGt6vDtuZ+MILNqlmWK0bftVb+
qsxxX++GNWcRmI4+nHBxckG7lMNIF1dFOKL9Lpb9cBE3dzZ+FLr45Ga0c/smEE8KkT/WcEz0+d2r
j7tlSi9XTxmj62im0x0EeNyavbByMgQ6k9jpw1jalg8LSuVm7R0xVXZ38Og7S7mYFiZMcOAwAWyC
VIb1QJgvKrWN0t6jSl564OsInNB+ZcMhpISZQakSfDPKJU4qiDTxMNn0EkhedJiawN51t7N/PYIL
J8/fgSKMaZhDDkuE316gAEzQUqd3rqmgUMHyD2TaG61Q7++cjyoKCUwL+zmoe2eHXJsSY82XlQAz
V+aLNcNXba23YQ6EO5BmwQaDCFV9Io85CXSTHhK51l4F7vzzSLhPhI8NMCmNWO4YFgLTgqd/S0nP
J/khQj7QKfxRJ3rLzBPXtQEi47R56pNdwQGrCi72y7RpMOcupKBHp0At9wwJpcyR/64rIWMLAh1b
NuPjVM5m8NwNS8QKsDHxu1SoO98XAlY+96G9a6/ZxVWPb3R23a8pUG7cDLulkb9YE0AOIf++AxZ6
DQtRXc+XEfRVO7ChwnzA/jOOngA6y6RRUJcPQmhoCfr7uohFWBeXvZL/tByOL0wWdIGJj8pTIyCj
+h21WcXa57fl92mKP7meSrUaFQThTb/qjlwrZOwbIDGCw5sR9gDOUqIBXs78YuG/47ReS8DMOmZl
siK5uRSYtmEJ4VL6610utUNciPOtgtDP+6geDNubjphXV/6t41j7uMA2QkRGa82/PToThsnXpkES
dvCJZt0P9FaG6DAt/WBJKlzV7lOz5Kxyk3bE3109Z5VEKTZ/jlRNM6PfoU9VSH0+jYEOG9fr+M+6
fkCQ77v/Sk8Q9SRxdUrR+bkULuOPa1a34H0dv4iP4w6kNTRa12W/5l+QGac53aaMCgs/uQp7GINL
87wa610Zm4TqROhbngeiqW4t8E6O/gDgqnPDzBJrTmgz9pTIp1WkMOsrc/BEp6p9LrJxPQn52fVg
G1pKqq8VLLet9T1EHT/1kMMoK3m759RDcOiofsLsyyr4LK9x+EoMwGmtguUadLydpRgzPJ8evic7
CspHM36vDj9T8X8Bq6p5nlyhqczz8LRL4kxis3pqiG9Tt1l2yuZt896BXIi8KWiyrT2sstDtU93d
noF9bbIB65ee/L9VThODgvvT0lj3gwp5EEl223MT3oF+xYG1QIjCxFKgIyyFoCLjeESyIayYc1kw
SWMa2y9Vn6q2ZSTuxAHhUQt8qoCvPeVXTsi6sckxMb64KfUMa4uCSYNICpfBsG3xRYnqepdQhD7f
v0VlGRHoV/Ecm4kYxeMHa/8vwauO2D5I8Ogudzx+kJqmKdwzgm5IW7vDTlyFVEOQcZbMXfmsO+Sq
dMYUMivSSB+0haC6TRsL0Nw/HyhEjbkjWyA+S77hnOwH850fPR9wF8alX+1jDojRkC22CYTmsK5X
bw1jnhkvTFDyfD6oudvhuI5cggZSomiyyKfNpB+rhixGjI0JXprSWjG8viUpL8UFi94gFQdb1Hp4
PDgm3VNpmHv1nYeDubepiIw5d0bI18iOU8HVmDbz8eE97oOHdvNzvM3UWiI5EJPmcuTuQ9oR760e
5IbZ9nGFtukbxEiEfH7LbpNMbiYk1LYWBUmhY1n43+X5W5bhSeucMC1rDciqfJhZiePyW5RhlhXx
42x700Xg+uvjefT7xRidjaFwWzUz2KvShUBLBTHyUYJV2oljO5zwt7p0jEvy6pQFSrq4+V+fZ8BY
Vp6MKyuxbQcZTI6HIy2f8wLzcIAEeYkZVvo+XfLrb1KaJ4kd68xFDVN1IL0g9PfoPy5jQxwXRFNP
Sh4wIHhtQXha/vel0J470HXYx9SH6mif9jixLf4XVxHZSiRH0o3znR2++jOlWGdJx+6eB6M6zMp8
bsiA2qEcKBrBeXd6tu7kEBRZHHNhhpDY0x779MsF4+E38dyuplpjKHqFW+UkHUo1XSiM3Frq/btK
V3Gc43hpkpQiEmS1S40wMAVk4UyCPZJexkY19lOdPdRLZApSpQONO/bGV+WzIVMnIGHOPxRv0/Tr
Di/hVVQIq3a2Z3XPA49QqM7ROahTmSn9V2nG+xX/pE3eI+s7oYWVdNmxYRoqOQi1jeVWSCUzxljW
THKRL7NVoSKI5FZ6L7yooarz6oj4GwGLAwlePnFmz940M5iz5inCK55tWMMuk7px2UHl6zgxQFQ9
x+PgVMPBO/IMIrfYJF0y/RXJ7Ev/lZSxYSNwgJOnhewba05K5EGT0A419K/N3DSXfR0lvDoQ/mjk
SraXzV/PkLpkej/h5OOi89Pcdu6aQOnLIRpOyVGa5lbSGjVj3FFTo8rbT7M9yCWVrhKwgmIaCk1I
MDe6XQL3/OQCQkl1636JzPs0MYRTTtiUByVEmoQo/1fKCTp+m0M6xodHsDjBrhuYkjPVcI9FLb7z
unIpaiCj+DwB5TyitnFEQJBz1FuzbnxAe+BF6e5z9Dqsta/s7W8301dDHxq+FeBpBXgbbYV8T9HI
VQWERZQTlc6lELzFu2fNMcV/Dcbo6/pLxDwEzNB1TXdhLfrAmLNW13cGOlrg7ru3pd6OtF/eM8tY
8ODOdFP+SNsKrbXlGW+759DfAtYuXpqoReLYZ3A1KBC1vSyJZ/p7fUfLiQkvFZ6Y1DWPSOtUX5Nn
h2VU6uxh37ehQeMQJ9IwLplt275PrFY3ePSvQL/ZUSewLCdLgG60zZY5DA2G9ffqtfi64jsqjFmR
RO7qov1DYrspUiaLPKzDyBMWHyxnfqFIR8+2ueGkq1kMYa1C+cIrynZ7qjjll2uTCS2QGEGndOb0
LkJjtauB0dzseQ27i17BkzPkmS0qRH/9Q2hiRkYtouEsbB9wb9vBlqQGJwU8hy9nqF1VH4kBwc7Y
eoPvsVt7vpR7zPTHZjSfa8GXz/rsjPJeBDaYBMZGW0RzWoMHMNm9xEGNRsUDWFQNw0HCXtyj7UzP
McZPd0JPAnr7Eg31v0C6tfKttDi8YSXvrmaukn7CJFMIEbJ1jaC3+eVgtuF8t2MRHyeoBez+Z76f
iqyvOF3hUXi7f7MX4QE3jJrc5p7c2KZSPrWaL30NxFFYAknjiSXS8JNvoIXgGU7Rwp40X047gMdK
xrLkqDQMbdPlnGGyVMLi0/SpKniGiTBiNAp9N/+korR6g04mYMvn6mryYYe+ZEQMpwPrdYtANttJ
S4wrcs/oO5njvacPrVEEWTpjFpcs9Xsn3yVc+wqMxS/zz7H7+x/IK3MgfSJvT38SAkA39NLAXizM
571QbFXvvD5Cj8dNkvU9IIcqNakalOx/Lts71JacGqOLiR2vm0L3x11yHMg5RirnQq+y9XRA16RM
XMab4hT7Dv7gKYv2FtgZkTX3TKwb/8vrcHsCIVnWemOO6en4SOfFcEgqB/eaZBvxwt3hF0tEWFa9
p18zSJWBmN7cekq3mUqP35mivqViuej0NfU/sgLND5QFG4GqDwBIx0v68vLfXgZjK01bCju0fcaV
m3f7ZZA0yRm3qrPqAiNJZRRIiZEQg3A9cBx52rZxhfnkMqo5fiwXHxPMxGLO92KfRculPWvsWc1J
1/d2151pUXrRja9lJt96IhkTjeBWK5ZXtxpH8oD4PUlHu0oA5D+UKdOgZAYLNSZ7H95xvFn8RWsU
O0m5RhlYIH01HOGBJ9PJtBDqR6uq2hUF87JW5WddbbJdJ/ayUVVSltlkGynl3eukFAJwHiF/xydt
dLp2ovbbojRMaYwHcVEUKzDpRHh+5uZiOMniI4JCVm8DbnSu53GvN2Dgg6lAquI2thjMROPLKb8b
d9C02bFnn9Ye1st2Z8EAM3cMMgzY8/rMU85EGlSscBzd6OrWWEzlYsXPlMu9gCr22ZYr4t2kf0J4
i3UyYUv7jHI2NNSANw8GNAeFs3ulP8kBHMbQeFk0x0YjTzQp6tnuokEajc9H+J6ONnrsE8/xa2Rj
V5nVzj2JP7agzZnifA7fftV3UeWrA9+OnUvemfnqNOb7TkLpyZjsxKbNfLrC2A7A0xHOgJYdV3Ea
J8Ys4F2ih/HOHe1SCeq2lon/2gFPAk+80EEqh2okBnhb+8Pvnrl0KztN4uORADMuiP7uL63TpEdN
1zpFShuYFYsO6neRLYzfsiZcTSAQjeOHbMQluDCXthKc7xtDpzysFVc6ALS6g0RBCg7HXsCJTgFe
F8IwpgC18TScwP1S9MyB9uWMMtaP+GTFK1CRLaRyy53UQTjlEABRgpZAhEKmShZyaBaBAQTJJ06h
R47cH6mL2Yj7vb4U/j9rADDSm7K99CjQTPFcurwV3lrBmRE2LoXvOCrvMhyxJxo/GgtMGJ30mgAj
+QtZ5GngH5Lv4addANHMHG/FAYwKNhe18wjhTS466kzV9M4xWiOO/DjFW5+O+r7Zes2qjEsofa1+
9smJ3ZPiYuSU+X5eOVBjR+sMdW/6L7u+KjwaKyF1zpeI7h/G0ggsK3DGAjx9ZUvHBp84iwODTYJX
8o6aPRU/+bXs22XCi/sjuwwJPu2WEZkpbeRANRVzuTSImi6ZwTzqUDr0bNF4RnTogtJrtL5vmU1z
kGZBuwvBhNcwtspIHS3ao9vcj8Ffm/JGI0XCyOAaJ7LNowPSXFojp7OcqIFzcE7dNiG2Rlo5BEln
STUeS7FmPevv93vD+Z3V1NadwD3qr3KDyOySaDrRwdpalyPImCVVYhMEeQ4u/t6spRKHtfMufMMW
TnTQroQ0720ySyhWGDU8PxH6o9RNf6jIVqlMaI1w3rGYpEV3dFwvJNN1XJoyOx7NJu2dJTiUH4Sf
qvCpeKHVKZU/XoWcWCD1d/TtgKBfMDzZM7Its4HzFV22YbgArQccO3sFyFa0zk8oifMYEJ3yFZGB
Z4X/djXZJn3KXZDQrEE5s18k+dhxQNWLz/9FL9OJQvLPClUC+UcMSBQ0NXiI6AqDycfG24k/Mydh
BOdAGnJ7XVbA13M9gmLEaFVbpuZMNqJxcPGLk1K3Qvd1Vw+kQs6jwYxmni/eIZSpGHEOayfZ8QKn
0/BGu2i6twROpTVk17LivrVn7dKsocH5ZqxBkS7C+QTOUHa7oGN9/5GXMwJptZGTtH5zfAbdZehL
16DQlQAiAGBnG54Hg/EzAIOlFdDvPuBmKMwrHiJux+zJEYFlX80RdRdVtJWYHh8Retnxa3OAaHP3
2vdTOh236+JK0F0syu7GV1yXtcvw6R3mULqIVzYWCDmwV1tc8HKt5taZfm2S+Wkj0jEs7tOX5vam
YVXjRjOUnjfSbMfA1vrxHDfQ13FqxQzwlhFdE9xF6r7sm7DOgC0Q3o23N4olyKcedoXBxK52phej
RE7s3XiH21fUaWWrrmzNFJMc7moMypTyOMA+pIarYOpPpDIZzT3NYN0QJwNFqP36Ul1UxRi0WFQ+
MINrIlQdUfggjP+oQSZH0mnNmgVuuVgZfVVEIkLZ0MqDMmDtqNQn7OktQK+5s05el70HbVh4somN
TBbDtyR2pwOi4Vg4JJirB3a5bM1ENwPII6ySL6I21ZnPxyU876SWA4d3ZXt0KLx2JnTsfNcxHkkd
93ahPSsW+4tb4GkvikjY9fMiSXtts+ppvrNmSxuGmmJpoHjYPQvqmT+pkzWjZ/f0RY7H6WRlA4Gv
H79xKhthonHQq2SeW/bQ0Xe5HumPqYeeq9eIJ9nfdy/A/hAoD4P4SpoHphB8+JhMlFpkfn35n2VB
0eXHAFeuksLEtnzYQylR9dRiEt3nxqMgbT6SWZE53n5bQrbu8cwoXGOHsGf2Z0X+sWxgqXp0TxiI
9A5KzWVYhr8M7pX5e5hSE223xvfs7WPJdPVBawRwFTyZjzqv41wuQEwmZB8dndtY5BI2ys6fLOAg
AdnIEM46XCtwKFaZD6ABhoFqNL/I5U6vuXdVO3VOk5HUAnBhDD8w0cn40NDzzPc1PccCWDcRE6pa
noSu7uO3jSEcj3g/JcE86DoByq3xnPKgaVpBHxHIkSanuQSoF6+oIT6E35wbaQl/ah2BQnkdti5o
wusbmaYMBUUQ+EMhAagrizdkSBHSP1QL5U4+y0mkO1zT0dDhVmkMlMycyS9CjZ80lSzvkJ16Prob
lzcvXrh6ITBqIqdSKi9reDq58MnCSJ4yC8G9DLYVb0cPhfVGKFGfxMlFp6Xjg/fCeJqNWgRDYZU1
DYxAPaLcpTDre3nxlQ/7v2GsiJ20CJc+okapmIuEIOEpMurRc6U/x6L2KI/QYWkONVC9hF6k/oVW
mx27ChHXgyK0ItKqmkKdXPfk+EfUm69hRWVdnYxkAdn7ENmADk6a21AX/Q74o8M2jcOnrzhbQtGR
JmqRskVypvddPDRCQmcGvcj88wM1LnofBkek39YNoFox1WlYbVv6+UGvMrB3ILKB2GYaONVrJPii
H5FzYfUmoGGawDiM8Xz9RH56EAwaotyThnQfgPp4MT1UD4EAoCwwAmUdxmeAxTv8S0Y/JJF3jqji
tVPHakEANSdRWdOSYLTUCNrDagXKrebR5SUIYZlNxWtmPLdOPzFuaCKEo8fltawoRjcT+tj4djOc
B51hATiDE/hBGF4sNHvvfpQuy+v4W0m9JeivhNBcd/ePH8gv6MJGrrBrwBZl2UuzMo7EcjGrQ4fE
Q87EtxLgpFF4DoV4SbC2r3Z6aTOCAhYHod6GXZmRrqB8HqPFKGj3Ga0BeWTadTleYlbBGV4Mb83M
wMDFwKO0PRLas8M1JVVWGOs8qSL9FpBQTtee/CyNAsATtntVRFlLNgAgmskw2Ee1oqXKhq+SemuU
89wkNEHtPDJEs9rXE8Ai5Z+GUgacnYlRsmVqdkoqiaI3M3a1jaBnxjqdDzq/Rt0Rva5SUxBfDycC
Ny11mRsKKJq4tEklsbmB0umVheBpvcNnqIroJWddElr6VTUaR8GRq3tq3JmCQ/ekS8HROAdUFZU2
TFg4e8XJ3/vTn17uWUhy1TNmjOpV4Y6D3EQ2f+JA8+blNuM3kw2t9Z8ewHSyphn+4hKctnQ3jSzO
0U7NzIUNqwJ/7pjBPGMN+vZE2vTsp7AQffMqwC2vT1EYEQrGIFBRpMbHGYuWSDIISIyGghjFZEsu
QRAfttq8oeRRi+e9oYb0t6waSTrr4Fe/H6PhGNBL5wfYcQ/O+8ar1h0WtkpR3nI2ECYV0w8NOa3Q
kf0XnT+f1xgna5J3vByqmuq5NPux7RuR6yIwY/X5RnmopvunKUsq6mWAkYby6nHC4IWJHnDiZieo
9PYdnF9zxyRUrd0SBpmORgSunOs8VanQzQgPneX2gGZip5jusYq5Ps3dMYLPH1k91BG9qNKe0f1Z
S+xUxF/NOVzT5++oFrQezmJOK6uq73O1X9R3Mrij+wr/6XxCVmcwG8GLEyG/VB6nttPdliSx1RzG
W0uVRQZ9jTem5kKJaq47tUWkjhHeKlyE62xi4KJZ3cMfhTEYKHjwA1GWP23v5SOhUv70fu/4zHaa
+Q1JDsSlNh87cJRIwPKaWnR7Aga03grzLF2IHniaIneZTFSW9EVdk3UshMI091vU13x7m456Aqwd
SeL7BpW5k6Z0Oczx6DYkpuiU8d4Z85e2R4742i/FCZBzEy9XWd4v1Xfj1t1pqkK1FhCig9W8fnD0
6iUNp1eGiiugsohOFvEasakxeSFr1KGE7dy4bnDduc+MfiEN/BK77TsxcFwqIndyNhq6XSpcfomr
i3hgKiOOPwMhUIuAMFKYBMzFb6hdJq09tXwxNmySWZ8zouv0RjEEk1Ji00lbN6FRIVXjHseyDNpl
vO1eeYGNQKQbZJKiNQ41gMxstL5nFM3O60KI9j9WtDvoRWZXIx6it+cp4lxlvBPnVTpbofm0G8Cw
m/eWAg7MNRp1SyRnvHpAZ29gI5xnS9rQkRD9FMGITVibRo6jH+JULiGM3aTs+x2oEWOdnJGLFopB
t0Lrn4K4/GrJnyfCUeCI2BlqKoKr/llboPH8u3yidfXC2ov/TeMDRdMWNrKiTATmEpCooME2Yqlt
ygiphCzw2fZAqqo0wdSWoS+3v0MY8bh3sje64F+0v1Qf7YsXJwCfJEkEBSDeqVm5/Kf0BIJDgXr1
L1FNiuGe0BySTLg4W6vKlLISWRhjoL8Zi7SWc+iwrksUr0ftaltr1fGIfwdXHuQBYmWBBjy0AkKH
rnQqWpUgRCINCZLUgAIh9DVgLBM23ybN1r/cOM7jB2SUAUIsRMGUyn3NPqo1dZZdEfZInjwmawzo
UJ9tKNx5N0q7+lV3gMwxSYJJrLuTiwU5fqxE2fRXTuWLkRNZSemajY+00diX1uizIj7Zb0XL0/gz
PnRsV+j/ByjJwSBCnCqYLsQF+HJCwsmDSfWaCPaUVwDZHAApDz55p7Y6Y5CGCKa686/5tpVa3nKe
fDczEgqD0deUTR9IzZn9zTXPTnDKWrDTv67w2UsrHRLaJsUC0N4FQq0CWKzniqEI0zKkjrP0JNIj
Ui8yJEtiFC6tISSnqaFcUWZaKvMKpsZcj8dQX73pXl+0grwVojDVLpZEyY3/nfIx/X4/J1Ue8HT8
BQQfnF7Io9bY0mPVYJQAEDzbTJkn/5EN2dtaTCc7bIggAYrCPi9jf9THXrcbh64k6ROVkfzDci30
UueAp/J/EXrh0V0jua7u4T6J1GFmVYGv8YJHfng2iLoxNgBFtOS82OKOBDG6MhLQ94zlPuWFpWVK
Vu/UbJKmrnsri9GOKyRLNzZ0CBNz4PuZdIXGAKF3bx/IScOv0pW4G3zqLLvHWGF9QcAWNvTmh910
d1A8VKkay2RvlY4UwKZ/S1og8wsP+rL7Fq9qvY51tPFE9IGKD5+6M2VfEuZnypuQojTOiHQ8eRrd
xInPa2we8EFpPDCTUIb9gycdGPCxx8Ii4KF+4g4cW7gCyDFJauNOkPwJiQtTIyPb5ZOk6jnhqR49
/fSeuC8wHBOWGUqyJ/tuwWu8Pt3okNhOb/MzX+N1cqjCFaMJXLUNCVvHY4+pTfAcvYTY1FiWnOuI
9/K36CJsyPKdf7cUghpANL+HCvGpH3JCrH2wAqRfmF+ZwXOktbfp+p+L5eR/1YoNtIEEqeeEXQdY
ihYca7zSc5376CS+WkzB8oepo3HvYIG9v9n0ht+PkQAk84tKK1suh1Nx54fFVIItwpy4Dyd5GWKt
ArA4+Z+TB00cNZ/t5BpNfJilgRvARQ3HJQ91Mb0Ua0WSesJi3ZSYZ4XR5qqtV9QHiVtLc+O1y5ng
5UjwUu/YB4WgS1hGSDDkT6S3MQjvYFGp4kbGfichzLt6mMTjmEflu1sM83XEATwQETWuYPd3cUxi
QZNtuCdFfgqLTaljFk6U12X8IZ83MX7SjsJ+kRL2hM7JYA591Q9+S5+VjyaaRC1yWEFd34gokUnK
fXAb8seRUj2HVmbjk4N44yvvuet42c+Q+1zjx4biSWuvW7PvnNrWfC9JrDtKVo+HyE6BEUrTLuD3
E4F/JIinRDPgCMWWhLidxcPCJui0iYB62BeNMnOyou8SeqMIemnYZTn5QAJCW6NLBToTJXqTfwPD
Gtvh/7XreOFfQO9GL0tHgoUMm3FXEqqj5sq2Mg7Jo5Q5nY9kH1Ud1l4LAQGqVOLB313j0eB/zPuk
T8RjBney+h6hdbnxAq6szTegoNEQct7Mq54sSGoz2ubM1j29U2SrjcaxLf296SlBE0d3bLMHTQCD
X6bjIq2eKONYpoTQAqJkvW9R/b6M97Uomtiv9H4LI9nqyV+nWYoh9y5RV+61zfy8nEmDK7p34960
xpZMVrXau+SMgzPKyWO9zCq45UfMfO8Xnxsjl+6NQ3cu8/muPhie+wHnFtyBFvBJn6wCmlSpC8ly
/K0SlNC2FIcxdzobZkCCi0E3ZApsvDvhGo/sQCUWQVTGUUd46HPhWOyFIvmIlaAufyjgf1YRTydb
Rdd6F/rSICNQtSNKdUJNQJeJWBE3LaMFlpwsrjZkmJm/WhMo9rm1xVl4B0eQ+XBRsDlu+5aaz1ke
8JdjIFqbLp0wUqLdieODrQsLk/pjMZOOnficagk7rhYbewBGCIU3riorngzDPklfLq0pBUqTvEyv
n2fmbhpTc137kpnuXuWT/dtwH6+WzSCwbJws3DUO7qpjIwgpXkd2XtfX2cu0YUpMCMXTQdjXIqwz
6P53q0/xAbZce/6IUmRhsyE+rjS2oHH2UG4lx/D2OxQE5zwIy9ACzygiDW6H+MLLgv0y5TLLGDB/
cjYUurnFSInMEk8yj59JF+X1apUzmUMWt2pga0UjzQMK5Xj0O+U3VZ46hMidhzrMy124Ciq2tzAA
mRZFCKcEcYoEjvsd7y85AEBFRWlG6VB1lwyvw3kxl4xCiSjuFdcXp8TZ+wqQurMOnYvHbLks3y8B
2Bjy7YudjJpxteFSNAj3lVjFVbN37LAKy2dcPYD88txTFQeWBn1z6RS0IfotcyZIFVhkB1WAdpSL
qTP7N9KAYQYVDVIfe+LomIiSkghsyVAMg0TRujLes8OPBH1AN6uhD6AdOCowAB5fpc6aKuJqKife
jzBQYk0HTvSKKoptzd/3fa4lZuPUzlxcO3z5Ta0sWE/gpa8ws8QckXr/b4SRzASUu4P0JVg7N7EG
lHiFGVnSb5VBuW68IOeZsBw9DD13E/tc1mr6axAV5iQBUI4zKKjkMbYIkjNPT3lEHGpvkoFQba2N
4DU8ATX14jBAjuBJbuKovnqV1yw74AGlcormCfQht45e/skZx1zhvZzUMurp5Nslz3UXkf7arjAv
1YV80mekqYaW4frFwNSGoS0kV7aX0zjj9RL2EpFTgaJhkzCdeHZ5rhtpsyzFx7ASy+FNRkZ08S3u
v/OO77x7RTWE7Ig3AmrUFpi+SXXwJUNMHdx2JZ/GWtcBFBgH/Yfp1xmMwFnId9KUf/OpU+LuOYCX
4Q5FSyuypEqW2DXuEU1jZy9g6s79ntycryF79vNwZstcuDK8QWnzUwsE9W51JE8PwWFIw++JAjXZ
arWhqtAKm/LSGSjQJz7bBwbSI58Usm/VQzQU8OSvusJM0w/59DdO2URODk7CiIer3qs3RUJxLD0d
hC8NTncPq/h8WNa03x2cC4e8K/TsYgudgfckB2IWi2d9qgEhpNQd1aAdL59C92ABDruydhY0bjEC
UGURNhmw7Wv0xULoR/07Mj3Rngug/muWCZ+LaHiKMA7BvCn6sEf/uLJxvTwljhXNTsHfUGilmMiO
lYgkBDa9bK162kxjf+IEGi1/MCgqIfj+hvRfUke0HAVRjEanlZooqQevZJup9U4uz/GPqGj8V1yW
rKu1ehZ4kecEYYI1o0O8ZIx8TUPXjVtVLpSLZ8ok6WOBNuZM/FL36vmj1u/pMjniBNNibXVllM8D
1CBJLLvZUoBhsk1S96pIBu8E7h+eFUDfhafnpiwLc2hKDVF24il+nPUumfzP/9Wa1wAkCFEeXquL
yB/pjkQvIAgqqwNlCvi0QK75pRd9EHzuNYNxQyUoRg+InGWV/ecbslrod9au2sjOWxxqzM9SKk6g
mC4CjSkB17j1sd5Sl17dIPgIMIKNCJLJETCGKipqs/wcwLw7QQukHl3RUXo8DxpfrPSrWsGCTqh8
Iot/PphXPDG/AggVFHZrLoUJ4YOLSV1x9uW9CpGAtlL2IpMUm/Rc9qUL5FQqAwL3ak5Jy9XVBjRy
45Xu5aoswXFMfMowgrxACM8FQgXGqwcDp/RNkqcr1+0A+uCqpzS5i2Xhxs+E30w9O/wFqnd2ZyPO
84fzzOU9h8Bwx7dMqHlMf9Gkch0zp/sWv6dHuUdX74GrYYI5G2hj4V3Ywjk2DQO6kklmsjExh2Y5
2zWpVowtS+yg7ShN8WI2oal8lBel0Sg/8fypMG5UnvaYX9ASV22cSCyL2YCjvp/ujxf2u6qIUD6+
v89CzxwHjW0BaLSbBJ0HeNznTdVV0l2WxpG5y02D+nu9u04R3mWqDOO78MjqSG1LRQmHm1FwN5c9
OCKJkxiAcLz1WcUC/3Q8LBvGSfsYlGI8Tu/KtWtykhhnt2j1zwpdTOSa10pvMhMOGd3cD/LeEkMH
afiClNopozW7i3LNpsgxPoIYNgUopdZZiBMQr/Zp3zib8iUHT5ndTmMDA55PplOcoE333cg/1hmh
UBzeCk9n7NMp3E3r+81IZ179X4WKzKPUtm+9mZamu83/UKJBjYaiBXvE8q4sCfVYWiQuV18pUDAN
HTIIii8QV9sWySefPOL/iLbQ1ubte23cq7ZUMj1ETbvOSfN/UEhJ40e/QcVMQgncTh9v3XRLItB8
9Wv1gMUk0bbyYt64DHaUWGppJ5ahJpTPjudq6q/SrI/a30NAzGy2QNAel4o9kfasUuSI8//b79OA
aSH8Mji5y+JsLqAQZaxIn8epje5zJiK6GmKYtOfj4Nmg1frEzhm67mYCs5CcZCgiLm5tykvAoZfG
kDadulpmSVQoev2tQiof9ULQDQkesM4RuNM/+xj7Taucg7DxmuqaTbt7lNMz9rqiLwSZiyexlLpJ
gpz4KOmtebMSPDwX/hfPMBuppuigoAhRzg4bj1mkV3lksEZjgoCToPqsb3s7AtPGuwH1tyRnWU/u
4qiaeJsvDtJV/EyLyn5n0gMuowJQYzc/2QJoSUSttlDmeHKHWGNtp/JivpgFyaE5/GhziUgywcSh
YjjPvhCVI7BGf5T5RTHRPKzGn6XcF+yEehpHmoWqNZTOcT+O5hl4B2GjzzJNzM+Ctiku515LtHuW
oUew7fQjphll5itPwuHxR+PexxYXTRDwRqtU1Ivdca5XW2roIBzYKPh1l29aXVedJJ5BL1ELBYsH
PxY0DsJ+3amUXunxgUS8SbdoQUZv0yrndPpkix1EHRtRtW41rr0SNp1ena9MPcvcQYwcvflkXMUd
+EvZepRONdxXi5fuvo6hHXJ85awz/loxGmZtIN9c7EoUIDANOKBCq1Cvqa+I6lg4tmupTqjEJvPp
16Cxkv7IBFEReezUs9KXEry3X5pbkYkTET3bH5HdAeJFsmKXU9P9NQrSIqCDdQ9ZADjcrJHZ1kF5
M3lF67S6beAT3HxkbbRBJManWNc1I8k+cHgs/hJoybdUpvK7OmE4XFT/JGDAUKGRNAQAEiDYWZaj
QQAckFotMj3+tNdUTdmrr4w1lnYcM//mGeqwpn/0vgroaM6sf2AUqNt/ACQ+YKK2O67yN4mW55VN
VL6XjseMPp3Ov3l0agtXz4nywW23rPyaxu6Z1lvj4VAz3Ve5EIaidLy0PotU6ip7T12ssCKfzloH
cTvtZatFOqYG2x61ez3yP9kPujxRZSlC36FIr7wvp0X3jDA7b24yshLNagahDeFzFFcxz1+ELY9g
TGBeGGh5310uqiQJZPIxl7gsh/Dxs4v9mBrZTRBDK40hHa390dGlZVVnimF0iW/2CZm8/yiq3bVM
jsWY6YxTuNo/aUlo3JS2tISxCBO1M0QLg5tfsrXjMqd1qOhKyoYCqNS21Bq8YZwe4LZJBV+nfFEU
8gkriqvDwrZOK2dJWrnM5PNezlowMA3ZAKichi+k9Zt2cOM43qS/KycOXXjIl1fvlS0wtiVbAtN2
0oCGcjm4AbP8eDDaAgeUDbBoM5VSe5SiqYdw5qRuMGaAnkZl8Ke8PACPTx2JhRvyJE70hdefYIwO
A0mSamEqeBNtdLbKotKGIZjU8QtgeVhXYCXmQJar4gbFAaYVlstfVE8q6N+/xSQwxKEu9UuEHn4j
Mv+9zYi+CBFRWnK0ZJBw6pugjFEhWphKhdXc0Ja/9q0vtoykMkUAW84gPKcx7uaoBHDdFR0mH3Ii
eom5tJWUmlQxL60AGt2+yGyKXhQzcwjmFbm1Zo2FlPYgU5LqouV2VgT1R8ogjA8pjL5EkXI5RqD8
qSxtRVi3jKOmvocYlhA/j5lrRghpSIB9G/buM0mBo8tlIPQn05Jn7AoXXxJdFvSNKi+1LmUlWepG
RJLynEHF3hGT4uwr5h3s21AwWK0/yAEaxo6a2d2O7xdZ2KHzf3qOhOjTiN9DfrGnG1hlEvEgUdF/
Pi9K5n1U0S7/x/tXlWRRM8y0s3L3uUP+6GpLZAzu26KoU/zDt06B+ePFQy7T8bVkuZqfQnKQPQis
cIbFm6KGixJOL2AQRAu4cQD3nop75R9021UzFVVqedEvNB2Rp/yC+tcOA+zrQpJYHn4wcriOAwlH
ZbGaIZnvccqGCzDAT/7ElKGq6Q/vNH5yg2TqPn0R4FLftYc2OAh9MsDBCK4AMVqUtcXQRrthv7zs
fGueB23N8euu9R/yMzPGGVIWFrF5ayhtAZ8hkrwTh4yUXGRMlw0y+DXsBQBhfW/cTg5/ySWL/Hq9
3EPv9EG9rBfrWv2UxNRPores/3/Ey06QcBUhejw6WKMNT5XFudAEcuU8JjWA68bPXWUNDjNt2RYG
FoyIFGB/UtfWWZ4oF6Ze6SBWumGzxgzq/xUij+gdf96dGH5WUYzvWAvosEnrPbQHK+WRUMn5otfG
oN59jtHshL9zWcWLldnE3a5NJ9lGTruheZ/dWTStOf+7HqWgPNZOqDrIT8XHcBXkY8Qk4jGx0VCj
JxxqlRJYaTM3t0Qm9I38p7XN+gIJsnd8ywXPeBUqWPXvUtDhqMZAJ5FdZ5H9GwmysGJ1nxbOwgXI
c1IXNHITWAnYhNg5PpPbvI6p/RsuU9qbbRJjq14438XhffhcCO/LbvEsT8je7SWLoJWd2xJUzMoW
KfL1U81jY1Ni1pUR6fU5ol7vthrIJOzt62a/f/EtXsuZW8raV0DeSmIOV6GxuUMYPZreau9KlOXo
p42iMy2vl1H5PswA9DWlfx1rXH3sjJSMx6BEv430Pou0rpvA5JX4vDD4yQYkJ5hq1CzEw9V1a8mR
+x314GW22WwaryKLU+8jUxN5Fvm7Z+tuYFzrKLc/6iIpydK5n76N62aI4n5XB0NfMAz9T021qmWQ
s/zEf+QZvAeW5PeVuxJiTe8rVigwNFyABdGZaEPIy1V7wvWtAvUtsaU19UsMiMiglTPufPsk01lX
yNuvdJnDahuKqqimO2aiIq/mpb9mnAVe2WA8M7n1CPw2Vigi+T9OJD7cul8jiqdQ1w+w0v9XTHDO
LQl3Waz/ID4exVlHLADAjj29gKuCSWBa+jkBmxddAubmQigg5RY5ZW0zgSJTcfdxz2UPk14Bfv+P
jUN2qVv/v+IIDIhzixXE7Nhp2Cq+PuR6IYSdmbZGFA7yValONNYMq8EkIz5dcMrjMNNDhcHGxvD/
uuCC/4qapdASmvvshRM+I3s7yfyi4UuSXq/5TbbBpkoSEAWIsVx3kt8UMM0Mz3djhA2OckEsYS0u
+YJJw99BOcanwrQGupQZWdud/WXGFJseyX40Gmk3xGCcpmPGIjZyAHp5O67DvIxZ2X+jNLR9dP0K
Rnp/O+sL/JTe3bAwCoXbzGQDt+UhQgHolfueQ3fm4Np66QzNkF6F2aB9pUOx9CG8umVH6qwxOGFT
+80I17uMGEII6BRzMp52MaKHxGGc9zDAlED5GIeilQD6oLzTH/2aDxkatEbFc8KoaCtYxvp38Acu
njOXBtB3R8EJ7ZQDjPtI2mrwM3Pa04zzl5GYKqjR+DWpCSFAJU7g1ErvpWJ4pRbcYKd/9HAbN0yW
u651EvRfBGUCBXobJreObwiasPxCWxnVn6yBD2EXpEpDWczPoxTfiDsAX436CL11oNGHcmOKYw38
VQC08vJBanZjfVvfReNgLWVTpD+kRABcnfUZAzbfR8Nc/QOlCqCFmlkA8W/HqJ+6yHR2Owl8FNfo
p51z5X8ylDNQN5+wsyNTGDZUilsJU/kYjEmi5s0KXEsmP/aIa8xYN2V3HDfB+wolv4pb64NPy+fa
TiyWr3hRlDm4DMuYYVW+e1kAOm4TMAT5f++UIIPIbTSx5otpF01pJVzBtrCbxtfSHZ4D3IURiBYs
SDZAcm7xD+FF3QvKt3wxWfBuDq2icoyMX3oNDlbyEKDAcD6tvPAGfDe2euvqh6yvw5P1NqSrzd1H
1+o4TZvaAFxr7WrWlj6GjQzTGliALdb22Hu90jK8LiQKv1dh0UXrPozctc4yrCb06SBTL8V6m1iH
x0rCeLY1e7Bx/T+mjuK95pZObTGSHcd8XHQOi/YIjgS/DwVI1WoOSgfun5jgB+Yra7FqeE1AeMS6
4AJrYFaw5iEhJkl9PN/8gn+yNKRTG/E5o+agPkMMp0+ahOtXVzbv/Ey5yPwUKuRRxmCbQFvgTfG6
eNxi/FNG5SiYudZPcQXQViNez3jd3w9VbL4YVGtY5Rd5rKsRCY25dWopbAjCl9iO7Fsvg8Sx4xAX
3IFjO2Oy7Lbd4vKh+8K3wexElvYo8tSp2BbdArDEe0xMZykd/eFDmxODgiSIV9Pi0qBAlL4JSQfs
rN06O0BsN+tn/yDQFi+fzUXk1VXzfuwTS9lXa5Wl8nKQKVqDckXNaJIMigFdAUoKTH7lptyZ/w+4
B2XcubDJmmRGEuGaoU8SO5YBs3lyNqMwg/yGO5s6uyHbr8fFWnJnEJ6LuzXKgcHqQRGbyFfmxz/L
LZauq/MfCGzNluWUU5Pt5sqP/v91FsXMrykfFbnrErHjg8HvyfpYsM9g45ZdDq6E5u2HuofgSrq0
SsVdHTfvSKZqK5UMGaOHypycwClIhJ9ZA8LgOiZMyNqe0GiKOSE6KqSgMaHKO7bvMBYnzDc9wdP4
zWDXMSkUXp2H6myBZO6ZZETtEFoaZmvBX7F6WsGeS+HNTvl/3Ru4N7G9E3dH+6AY9KdYQhnetFTn
maQd/5/YgZfsL/sLPZgQ0NxevKQI/6eVomNmlciNVMZMzIJ3LJswcj0gYpjzN4pyjGYhURcW2/Dp
MpEifmBwNQK3Pj99+BRGq1shxc9Tvhu89rM1aqnzcTnNGrdmV2jQf/nrnouDyjNh9Rk/ig93ss9X
WAh/YNBIrTpIbD4DFLNJVaVG0WmeJZ3KZ9xRBLeVPd5X7PJ0q9oLgGfroAVo1vcBPxE0ePJylCge
eltImZ3f4KKWrhmm9mWDsvfGhZQwP24ZrPjDZCsgpXkUD/sABS9FLwINAW4riEURz16cDUYXDqiK
j0loEVpLjTaIrM+R2LQhxhRrwDX+gxswWGomITZZUB/1KSx5Qz2C0NPKYvk0rRPKUkihDQMGNJHE
7b382tQcAI5yaqXatFYtBlRwkyVlCAhKEa386jS+QMbQo6LG31hSyIBAFkuWGdFzGJ0I0g6ibcRf
dU40MqQmBE/0xSYmjlOP3fTVer2iJf26Wk9dLgHIIwa/2UwQuXJrrkPuFob5um1Q2pD9EqGcSuh4
ZM2LnMKkFyTqYzjrOY/znOoGH+iGsjD3tfBbWZUIJJMrnFoCsMW6mIONr6pXU7KLhaZ9M3ygQPZZ
1Cb51RXWiRzFagESXDvU37RgwLMUWEbQCa15wOYlCC4T3+CQUCcGKQBErOoxlIunwMp9WJiW13p4
AZ/1Hkoi0aOkscgi0OmXknphzsA6v8lGliZVWMmCKaUfOi9XFMwyNSmGdcnBNbDlqUoR1jq+7Wx2
iYq/NdgDUkl9KDj8xKiyE9g49YU+nD868oygoXHJARwKS8oceTyj/tXCvBEXDeH4bzKEgWNrXA/0
eyyD+drxXx7Lahg2jg1rw5k3337gDeV9rkZY4R6QPZCBoJZn7xJrA82TgpjfHCjujGUhzqxVTGH8
e4zt2QZPthoirvxpfjSNH/hARxXFVfax2xtauGqiXItS84jYwJGDRY4zixQHCT4lTEmUrU3V42/w
EPAr59Itmn5F5fs5quXZD7bTfxK7+SFrBb0MIvxiPwAE7K4twbTVlMluQTSyHu0ep2rPxUC3opNe
/zbWoss1LCUMdsOEzljtMU7bZ9L+HsjX6VIYFFATadfakVtFDAnQldVMCsmcie1gBTEjaUGibhTM
noSyqbEQ/9cLBLEmiIHk8nwMQ53fXg+ByCJMHn1ddgoeoCivVpxSGGUlOHx4zKm8Kw7g5GBUsJF7
e4drMlaapkiSiEKl0FmNSVgOEHcGGqzKMpxVIMWKFUniyH3QhwH8dpLZH5v/+im6VPrW4dF6w37C
1+wON0uQXZslpiwixu+9+g0E8OKS+J4wJ6LYpNWJTKWRIH6VuMkjnCoM9LuzmzXVzxiBzdOTSJCs
D7cJO4wtwk9zVHPPbaP+azSUg8Ek1vJ3PCJwInNgkuE2oY4cx0jDyOGEuMSi1d3tq8zKHZQR21Vy
Z/+Qu6I60u595zsrNpvsKQBCMEdDppv5iN9qRl2atJ3ieWpCL1P//OBlolmOmlg/n0/DV2A2Q86G
GqEV9J13bcWb/5DXYvIcdv1hhwwdYDTXGJyNf6Vwm+RpWXUpQV4uB9GuG7iosGGp69JaP+/t3rEN
fuzmB6wuIJDYmor83EnBJ64rJ4rvVPAT/e7bVl/votZqVbUBp1pOmvGrRMR1mB2cTETIqnwkWrIx
wBabRbQdnCCykZPePIZVhD40kGZGYoKT7DiFeHH/uwV6hj+DGNqsV1leufM8ulcX0rt68CQy+/d5
7trSMaF3WCdDRmkobG3sFa4Ss22V48u1gUKBjWLjKRCGM7cGUC317f1mXV9uR6RI/m+exo8pk9sR
8mYjAJnlGh1o9KsGzNOj102Ks6qP/Z/t12X2MJaV4J+xk66tLESLOogYX87yXvYgM536kJHwOQnl
J5wpfFEZFDT9RRkocjJ7W1yMWx7yl10LXFH088LNoe2uxUloCdtN/Ln1LA6gdMb8xX5d9yKc8TUf
AeG2jvQFew2SLlLVV46/dBVl4JgvuxWsP16xkXvx9HA5doSk5z4JAboqPw0oMyLVR/oU4z/FXeW4
rhsbKJWPKMleZVl+vYY+hnVt8OboRlqQomVzlSnfQxgkfBdR9pKYLQKXsnPO6SJppO/gnTZ9AQmV
gPK2oBx5lG/6+fjRzjWvXiK94pO+PzxFul82iLIaycyWzdZ0dVD1+zuyKXmshGG7sG68C8mPj4HR
vyCAB0fHNg+pPj7Esmbat+7dx755MRITfZ1rTUs2QXAe4KOswyQwST9NvUeYrfm9XhyCHhBBr8Ik
aYALOdGlLwKUWN405crk/4Q7mCiTVqufaPfG9H5P2MZyO/TKfd380enLSVILqE9LXF1c0AnZ2mdx
4ewul2aa8IPs6YI1I8mE3H8EaZ91mHelgl2k08F6Mh3cjAfzCwwu0YBOd5roaWZsSNfh78UU3d9n
1uK4NuQUQu2tHIEUeXDrhk1k9zZJDnu2ewHT3zqVHYS/pQAxx+mICBgoKXmGgFUVIz/YHLhMw6lt
2Vvv6K8mGIZ9BAZfk07rHhJZy446YTApa0Dy42MeG8jw1pd5r/2B/dEU8MgQxIuESLM6U7DZV4tE
RscSb6+ctoPZEony6YbeOXq3tuxdw/0BD60rYAk6jDtQBRCnABy2KbaY8nqGVveET6EtZJ+4Ow4p
e37JadTvDwupW9A3NJ6WJFebyMHS2s0wYEQVAfADqhHHFJHjw3ji8YXKJBpBG7oG5Xx9odbUg039
lWy4/RolHqJyXFF2uXybzztHM8RoksR7ojzqTu+PWqUBugYSpBfLzGxBndzX+XS7Tc6yNWv99Ni3
nipZT0J38FyVLgOCzM7mlDMx8eLCj73BqKgn9w5T91Cj5vMt0m93WjTo4SV18368/QwPmjzjQ96s
PyqUjf+zPy3tj/kSmNr13iTBuxef/EhwpFc7EHkMK8dUICdRmfgtjx9AkKqqG7uwlH4x9lJ1g7J+
Onb3OKtooBcHfWUxk+VLk6SMHAZOlR3pdDI/vw/oqacPwdimnuCRzdeIx0cYwALYtQtGIFp27dus
kfaAp5HxabyLYbnWME3c3iO5a4PQ7Wy1s7BpuvkREJ6ExOVngnNOeeWAlZZ7S2cVdi3/1CUIkfQJ
fyLY2sKJOIBbhS28JObApNHhws5GwHxCHTtt9TCUXbO5YVRwo/+bpvfVJN0KBcrmyt8W13qM5XIv
mdw/+vjuRrkXIa43VpvROY44N3rHrBm2BP38LyN60OG89o37OgIoS1HclYfk3QMk0p08yvpzCVHf
sTDzDFZ7DjYjs30D5wZwV/xFXSji2GfdgdBQ7hr7DCqbWcUo34LZa+9RZtf6VnmSUXhVJO3TnMnO
i3+5y/cmKtBb8cjoX/b381Nqb2EidAd+3KWYUOfJIZM6yd+RGJjnlipbHSgsD0c0X81PkcdH5NcM
VqQksv4AQWsHWM4HPJyWykLhJDD7xufbWcoH87T3iHGGz1Yotcqc0Lj/kW6qEB+agzazzVlnPnSc
F1bRIKGDEHjkBe6oqlswT7JBKUv7PgpPpZypD0u6xbcpQ4pgeuDGDsfwEgGBoH9ijbe8/8qqFPku
jZsGUMO7aaRn88Xy3U6P6hFZmA1HXOfyKFRaw5wXJfoX5FH/ZgqFgAmoXBKeEHJ+JntnwCKo1Src
FcjZm8aAZ6+JlJ7i6TFQN08PIMxvMS1R3TC3VjAe7n0UAXLrw1qPglaDEovcMEunlORH8AdYNInG
dB3BN49IBHeQzNEfQbez4oTDy5pa2bEFtSTPcL0aVZ1wPGIj8x7Rnqq7B4YpkEAwvfcKFgNB2bYo
gDszfvXrCmxh3UnJu6fgFUi1znsbqCSFq5SbojGOIl4bdXHHAR/N/RLlPBGlkY/VDNg+gQPa3x3B
YLlDwe4RQx0gD2+5zFyJ8gZ5HMukxCbdnorHQ/FkBcfUbCkm+ES2pigJLz+NoJqCkgsJ+jdzo9hL
K7B0QbaEX4EexlEo1IfJeD/dCn7iRbbobFa2yy8T9kolbQyzVNWReoA7SQ5AsWxcBQ+CLm+weUJE
/iXLXTHa4MRsqHuiYgg/CwnhA+Q+XEMeVT8C2e36mRAwLcPefKwvcYVry3c9QVVy+kQ/cNvfFlMq
zj0eZsum9XmUysl6b0lYc3IDbobQYUf4hOFwOgj3XAi0+2WsTTSUC+UUkSdXX+hEBorUqGrd+j7p
65waIaERvj9bS9xpOCsS+7N4037xl5Hy6qet8aa0lBG5pntyUGDYksxFS6JBQ9Tym6hBalxf7Y8W
6XUVf+ZAtJpkpWq8czNydR0rXu72YAjKmdUkmGtvv70gvqOClrMuC708IRqs//H+3uDOv1spGhIE
paipBviqXrDLMjzwdwJ3lXse8nFyMQR/dVcTFQJfDbtpju+J1rKzklhV3zBFBYK/7zTJrrEwqSFk
qIGrWiN2Vc7P4rKSB5zIVznNm0vImbgLES7mmZnm91kklbewnqIWN5Gy7TapEk3FySs+sE1YuAI5
jwdCy68a7R+bSeW6DdCtet0A7qThOOKLCT/mqfC1/OcEFLuDDiaOvHRBFsB80Qqw4H/Qs0exLb89
mT1T028Uoox7kVjAvKuWnITJA/6M0NLItt9Le9+mLkvcfeyUKq9N+irZ5BCL+44WBDHJ497tGece
EqB16TX8LKVZ191uQ5Wd9xRpX/Ao9hkZzpNTBdsEzCXvm1bW+Pk/1D+y7MwT7TKgZybbFcxHyL0L
+X5qBGh7nHkc3moiicEKn1U525BZQ+0cIhrrZZW/QbxPEpTP/uEIEdXLLJoEzp9zPkmlttReWulS
60UKmy4stj01Joc4TsSi0ZIHo1Ea59crt2VaHW3U2ddQBgu+VBe5BuGtSN+9SMKYQa4D6zYMcADu
h6O2NYqvNdqvxrI1hGQdX6XSnuWp8hyQ15Fl6T3OCSiNZxoiqgqMHgbrEi0gQG4Op0hzfzSHv54o
1xAtTgrXRj7/yi3KtcH/MUrQkL48SJuOeyg0jzFsWrC6Pn3MkU2iQQTf2/U8AeR1LUs1RsH4yBSz
ViTdJ3pgsYjeRTF2WLhF6+EIobzNiyJ24k+FpGbW/cQwz1i9V7kUTTe41j5dIsLKyxZLt0kVJEX+
46qi+gLihFml3rgTr7Kv5U23EXtAuQYZm4QAHECZ6G/iMt5sXmDrckf8kKfCA6VrKNM8fhCIWtxg
dYekK4IYuEnpo0K5e8RJVggcA3+OqzXooah5rc4b6VtQMvPmlbwsTVVT2ue1HXevp0PH7SnG0yt+
tjYMP7XLqojXa/QHn+eNp5ZU+msP8jAskkCwfLDvMXDyq5Ghel1gHkZx9S5Smi4ms5Q4JLtPRyeF
f/m0xJmBI0m+b1MPCyUl5Mpo/pkz31E5oxVxC3SFCqtWYs60fMtVvNhEoPb8jc57H/GVi6DBoTKx
nlrmChZv+n1eKtOIyyWyPLHiJJJ+fQ1Kk4DnJHjb0cSaaHdBjqREiDCgwtZ96+L3bFTOoDH4I1jQ
Kx3/Xj4ivw1xk7Et7SQcIQFti/cqWM9Tb18OEzT5cqwbWuYjOIUGNW8fkJlV0UTMfceVjjujSWn+
jcCx13ku6h/jN5JFVsV9a7oObJUYcPU02l1j1Lm2O9qAZhEf6GqgQ2BZ6X9njleUivwaTCw3l4/v
DtJrvVEmFFNF0LGrSQPcW6lXHDiOWEL2FrLXpjOfi5d2Dz/X2qVw42YtM5TIWe2a/W4fL9ZcVOrc
wMTUNC0sn3RrKtzC47QyCznAh/xJdLojY/cA7sLjXUUj7gOqEZ2nYOTVgU9HY4deKq5U5bjXcw09
Gw5/YZ+ZLD99QJJ3kkMY6M9KyfgrL+IOJpwxzIRYzYyFV7S8wnFrC9R3se2h2h3r2zfjDxkI9TZi
pJOKCLMScUD1dyQ+EmAPu4EOOz4idZMO7JeDulRrO77SuF2CSNHwwFEXbXILlCw0F+ZwlW5EHg3c
jqWSDopcRWprA2uD1CLnVP74/KI9gdVLFac8vAMAznOULlblDzVffGGKqGhVmo2smct2BJnnLuxz
mIc9wtFVhyw/ned/2ulm58WuyQMONit6V9R6yc1B3MPQ9H8QfPfgnf5l23J94hqXjXyz4sMMlSov
oJvevAiMjhg9yj3Mw5VGEFHNW8qZ9d9ilXuV90EB717BhXkpTrKI0lnj740wzAMtHJiLTVgMFdho
NIVAi1qfMfq729iWkl63AwZ5L2fAx1xkzFdCT88fooj1JMR31gsWhMLfdSdQyiKR8utnnpIRpzc/
Ea3F6xUUGvLSVHZ6rK27UVj6b7Db9Hp/9awUWhWA2bztY85ioOgz6Sz8x659BT4W4wJ/wy4YjEDX
IfQ43sUyl6eQOiYviO/T8bcJ/3BJZkYN+JDvxSNtun5nkGhoOu/jOu+nu/5MyJeL6Y6oZFhDNwHK
897baXIgXmmIqSaHkSSInQTfIi+JtZQPhPkxTHNDFtvwzzC7Sxs191HYbqw//7k6LkaOX1heUtwq
5BLLP4HuPkkKoMcvt8p2frqPO+P2tIJVwsd9pQMfwZn9Lb6POFaTWinSVQLFROKHe0r6VXI8sdDE
2HVLADIh38ZtR9Kif5Ns8AMA2Sb/U/fCUvwC1+p7aUk5i5T60Zfxi9UcpNnZ0clo9lYjNylXN0tD
Iwiyl1dIgpiaq9cxiyj7iS5itifphp+LzLe2yJDMN5qF6fQgQIoU2O6Pz4GSLPWJqCMAKmZuK0j3
rAwi6hvT7GNEb76afKO007n4SZn7Q6v2565nDca8H3gqm+U5IB3FfAmXyUqCQPaeNInCURvoa72w
k7ePEHnGPiE/6+y2lDoo8t9+ZqsXi63aLUEGAJIV+OYhIn0ZvcdbIGZUY9z0OgmVHfELmQ6Yvyrm
jLD/KRuyoTEy5CH+RE3ZSU1E6FRf8v5OSNAXuMSnsOmFvOSui5isZLnQCW+A7Rkl727DynRlwUO4
5oeEFJv2PhQzfmf2HXGRhoI76QVYO6ml4sgWi2xL/mS8tsKKoz2MmUYbxbJRw/2CpPa6kce5DGlH
WzRNf6MGCPQ7VBy0TZR8B6yh6OyhSBhk5OteeteSbZUC7OnQL6tml1asvVbwMyEicZmyHuDnRNAT
lX0BtLKcX2aSJTz/OEFRhZTdLhWbOkzGtNThyT1Cxsn6zTXhBz6zQaojO/eT4lHHT7tvqMs97Y1V
mMK6ps+AW0cQAQ+0GDfBmXYVsidUw8RlpilmOjg/wGXCbTEwr5s5nFPpB4BqXZZvaqU2l+oDX9oX
lVH2q7UuXOX2RAkhDxv2XTx64EQsujIeK8jN5I/mwymxDVzHobmNndJFhH/7vufc7PYXgQRmaAmu
D5AiRuLaCsl4HRucDXvOLtIZWfCss4i2BBwBiDHGWSaVbX6o/YmRTWbErnf1ImfUpHOXgvrv6wfz
BySZqfkB2f2gdOfMOLiW1WeSYG1RGPgfwZcIu35s6xzQsCG56gMOkB/sRyjvVs4KtUnC0+rF7brW
0dhYIzzdI8SOuC5+vvtKfg6tkbrNOmnqBsheeFf7r2kbimB2fRdZCuzBzE7a1izxBAL5V4UU/Rw5
qn2u3+Dst3yyi5crAuUR8/y1xz8QNw5K/MgPCXZC2sCacFpE+zc/xJkm78MheDnrv3Vrit0b7Y3I
XXHeCEhnLsBiD+A4hDRu0m5vvAjWwTDxlMpm2QFj7gkEyi28VbXzATBwaflogG4M/x2jadgzfMvI
7hIUwOXR8u26+ne/BTe5WGvOL+FBEu8/EOeJx3LxtHvYJcmW9J/7sBcBeJQUUyTq9tmRpAQgfFoL
tgj9v16pdt4a22Z8xPAKfPFQZZUFQ9dhL4myIlSnltxkPCABvkVidultbklMZ289uiqxHS1jkQhi
GWkn8/5AiC18HO368ipQXlqT1z+n0XKdXLBp9GKXLDIhxroEXqc4hhyazsv0iuuuEaH+X2Empncj
jXtvu62oWG45n119V0QTxPDD8Wx6NUpPPuy+18e0YFuKkvJRhfNil9HW00+zfwrcpMjRctXsY+3/
gJQJd5D9BsF9+ierMyVt2M5lLjab9sCMrpz3ulr6s6DkPNhMcaZ8rcD/+86g0fb1KrFH4TtIOGWw
LuxEKO7Gfm4S9in22uvhaAuJqgOUcITh4Ko3IdbGPi1BCD5pqDhNJ3kIk20uNwV7y+QDxe49Dpz0
kFreQd5wjXD6v4Nv6zb4nC5sbmWlCQm8QvrLfgHTue2SKFPahJ5RFiDWLQCwzEOk3Sc5lLPeUnJf
Ykg2wcYcq9TZiSHyXN85kFwy/Ph5vtz0A+a35ULHPPfmCoW3slLlY1u/a+ykjpzMoIbvBqBVEBB8
CCPqQ8iuVBSFSHGESvk63jGG/yWePcv16uJrANLBRbiLWrqM3KqwAvGwr4QqOSwNq7aWBrLURNYi
Vr6CBfCk2lQ6eVm0IVc6b/il2+DxRctUJFp4rFkxewi8j7YANWlU4WOyApDNRYxbvf/Zhj2UmPzN
Zs3QILVVN0EKn/ddRl+GtSpnyNauEHs4nPDeuN8DLltW/DtiUVkzbNLDIj87jsn6VXFzm4/wfKmN
10YgTtMXNtI+q0T5igADRozMovx3CQ/WIWCWPMBbCn8oIuRIMvZGaUeJV8CpZVvrY1apnno4qaYx
DgGpPxatcb1in55gYRnx/0Nsz5vnHt/UB31gkRr/ZH5dXR/S+u5i7YBP+o5tjBmDEv642/PzyL4t
iLkfR+4QV9pOXhmvXY7ajn4iSoBh5jogr2HUcqhFCL7Q4L7Iww0ddk5Sn03Tn9GarbjreXQ1Gy+j
7FJbG6OROd3wb6Kpwz/5Ql6eq6MT4zY7GStXMbUXx2IpO74OWWyJKPcjKt/3W0rwsigDHBnKzQHW
7/jPonoQWj5fwN/6TSo1M5y4RIlXRCXCXjnOsJrugf0NQuxl2mGZ+QuzPL3tonMKQUyCiYqhcKDx
37VNaMcruh7o4xf2sNbjl+/98Q1xDZQft2TS7Z1L2QrLUzgU+OOtvp/IQwoh/jQx8oBBcUpz3Q8e
EyiEvEKGfdzqn/ZjapOAVMuF2uMoDxyVBFCk6wylksSf3XqPnBOQaH1U0Sboep7lxIh7e22vVDGD
bkWKIVCt2FAPoXMqFZf7tp2YM58JwU7EEgQGE2Sd6tTbgqUSSkMwCtuALID8Q5tgUZ3wYr2U/ihv
aVH+qiLGaDLHj0Y36qi74KU5XqDLYQjGiO3R8oWTlE2DHFRz/lxN3ZFOHnV5p/getz2qxmMyxCJ7
LazlfEDLlmfLAfof+sqzf4U4eC8+EMsPytxPDHbEuXWZrgUT0A4WfUmiutAwDJzuIBNe3KJmzn1w
1JvNe0cBSt/cdstWbITEPGWJMGBe1oG7Fw2YZDgKaT2SVLwvr5Y+5591W0/ov9x02KmEsQtpw6vC
8USvHlvoPGzdShKZVe5eVBBApRD3/tq/7JwGOG+B01TlJcGLEJDcThslRHnSg8gxrbFyW2Hzlu8F
Fk9UNcfUzs65ysbUjGktbjlQIOUCB9rP6uSMZOvoqlFt8UsGA/bpmE6RldS+TemouGeNUs2DZsUw
MYwjhVbtE7tMKPNpsmRuXQzxDKSalcghUA952/9Hhuqoc/sH9jgsJIGdQ1mwWL3v0luQ71LTIJ3e
MKgViUGqpGcSLSUqXaPfut4HY5R82+9Vil36mTbeuEgMuS0Y7XDs9x6f/5y2GNu94JqFADnqG1+4
e8mGFF6Nb33DyqAisneHMffZPGruJeGuLz80It3NC+WAZUEMUgyM/SRd067zAogRqe524mYGwIJL
rEPforVDro0aCgTank+wwQf/gBoTpxEt+gwJYPAB5nv0/6WeDdUvXhYl2y1FjqSs5FL0FM05BSOG
FBQBLi1Sln8QauGaKKiFiFhwJKVUyD5OI2U961F16vpjALpnrapmdR09vFs/OfnEQUreEy8Rf3th
gMpN5EFDCggA8LahilB4kqom2nidXzuM5wEEFHr74SCvhekTRDnWgLmcKYdcjwU/x/niaQWGaFMN
f118YEKj1PEIOl38Tv5DNIpJGq3GFB7wEg+sdMZ70W7T/6Q19SnvzAB9avYvcJsPK8jyMrwl3Fit
LtC0fdCxKq0m5KiVn4mgUagAOghdYNRdMgqXI+dhjje99sZIy9y3jTTiZRI7aS2VZEy9aMPLOOOA
xcR5cKR9uxgTE7d70wIhPItGKpoWVmBtJ2mZYPDpfZU4wks8PxCJOyQ/t/X6uIFJtRUeAjmSugkA
HPMlggrhbzUwjkTEA1eqhGdkS1Ib/kZXt6O5RkmN8Tf3lCYGcqH87LMS7HxL1icJnEpR0Nr22e7a
JcGiiRLWxnsLqYUDS7E5dhOXOkURth/SlEnpVND6KW1vp1q06yYygbQSIzGTZKXycvaRuHKIAN8X
La8hL/VkGIHzl7WN6QgChgMykwIXfuxpJGXVH7OqqATt8YRagg6QfU3d/AcaS5G3JS4OkAjR4qpv
Tj5t6BeBgnTwzpgyRR0oOhPPhAxAgeYLgl7gU01oVxsuGz+Tav3ufl5hSfUM22QUqalsTp/+Ykev
y+lhUcSwFIAFVVPibHHTCKNLU3DpfqXZPbZE2rAcCC6b94prJ0zZYiiN8K9zq5EhCblY/4bHJyvp
g//bV4wWOI+6NSVHLWosptUwS3qh5SxW1pOTluz1FhkTRydwl3JrpUV2cMAxBJrLHWSJFj3VS9ii
S6xKe6oWU3UvyLYW/KHdQNjIy03mqkhHGAbi2oMLGulo+0dfPMgFQq3kBBRtp/+T2FpQrjEXsaiZ
JwubX6RrUcZlpidnk1UfNFXb0/kHLucGS4D25zl1n5GQNkhYCMBGcf2clFbBfeYYJePr5DO3BSFF
CEqMQxtUmFvRx0/yBbkYmPYbaqGlE37713DNT4HPfWfdLoBHTo0d6bXoZpXDOyYZk7wP1ywGPWVq
QTRoNj5eDT88+IZhnOdAjy323GjFJ1OCrGi/JFRy9+IHVu5axJ8GE7UbD23vucMkllOh0xYOd98F
4MElCcNbJfM4UCdwSUvNdjqRKxWyQ81XIy86wSrfN+NKY+QJCBrKo8ybPl/D6/dp8iOmR2TtfvhV
8vwy6Smyb+1CDJdNHi+ZExh2s1DK+ebPGvbQN7x0KZ+5TKTMb/elNXSZ/TFEpA/tmr9kLA3F5UIr
lDGA9inQS923+o232AA4NFH42aM41ZbJdYJ7JEuhAmZ8TYssnGZXQ6ZWGZOpu9PAo80nzrUcp+iI
9np0urnnxaj1mDAUIOw6T+Ssuad0Cvw2VwaJS2ZVfLwW2LjnX+fzDGHTFnfQOIUvLrtBJSdAvUeF
ECOF1LxcgBuVZ06c2qwupeSfEB/t2UEffyDMQ32Tbdt11Urb2KxtSos3sQs5gotjN/pM8K/TNqzp
WkysfbrNxdOQM2j4iUVnEqxdIl3hFQKrONl8eOJwS0YhAHV0yjAdb+n+IqKIvVQxIUVktEjI3OUM
V+T/gDFFdIRhGGnmx9ZW3zTV4RmEKxVnPbnouXmjmSwmtLhSNv+WJWotJBmS1gR4KqK5KyVOJk85
prNTXWGi+1ZQubXxjNQLR6beA6SBLlRmCiCxGWtnzCxvDNkBvPegxuFlLE5yQSfvZ9yeNupJi5sJ
PFkAMC2dW0OR/ROD9knwynkoUAnUTV1SjPAr4XeTPUo6diFaB7uo50RLbAEzmrZ5ZvwCeEukjna/
bJgguuAb59hACguMTgNbH15HcevArlDZfYzGynBxJ+8L2Lvz9D7sp1urHe2xJRP3OUyfT1f6el7W
dSKI1JzrYWF+YhUcxgyYxKrzMnViyDs6ow9thS1npTn+PXLhgxSeMiAWgoFHxnYlVM/XPS+wTjdY
SFkH4LeF2RJg5ncqARYsdDhiQcjdHbgjDIKQoyuUz93v8Tu28rTWfzExtma8A+Jd/sN6aWYFKukU
gWbcM5mY/MjHiCWdwsxje8NecfFyk+ZIyibiLT2glxIG9BXOhRYmo+CJ2tvO4uD5PZ8dUr+Cl5gU
jRdLYrL+QYoHYpJpImPI3snS1ZMd3wIi2coVjCkEvRjgvVPHJdxMXhWf9GBkkIWvkwwI9sd2iydQ
HcGftfNL5TAiUgHT8w4mdfA3rRInDnfX3GuxnSnDpz07vb45H8J8k/phQTMVy+uhIWcMt1KwQhai
Ox+QYfwiWKDegbp2XatZdjgOx1pAvxYl7IxdpiSbGVSDM3ciif6cYp1hazuV/7ha28vdIvIRt7sT
ujTkYkhXj3VwcCTeUY3srt8rbx3niuUAhvrcST3vtgXrd7Upsd1cE30x5TQr2khrI9icFq4oTBCN
N7CEGP7dFA1QKxCrtFZdGOblMf4Fcdxk+hxg/MtUz8Og3no8Sm9iqz9ery+iMu8D5woTShHvrneU
L7ueLJ0uMPiQICqaWNNaf/fO+ZXR65rq2Gjj+MtHFWteUnpROcN4zvyeGaVL4+Jq3Ys9JGy9qZ3z
uiL3g55eluJjRT2SlAYRjpYTP2BxNssJ81JL6ogbsmIvONrocAJlxveEaxeCkeI9qxxjnUScQps5
kStfe+2z75i6RGc6hdz2a2fx3PYa1wfO4oIwUkqfv1pj2MeyRgyWemcGfRTMSyXoaYs59RnN8vWN
X7kj4+BTcSlr281PcapXNmwZ1LOQtw8lrwhmFwhOlVWWEZDWbt/GVFrUoM9WjeUcG7avdTBdmT2X
H4MVykbm1n3seoQOPdmt4t41Ctbnp80ZWcjrSGS/tCwNoDN0AD9I3WNFv7uJ226wODqGg5etPQQf
AkYMi3jeuAqCMD1XHMY3SdSwJAxtOs2+XG3vEPTpPz/2GoBdB77ZhWNhRTa4SoX56amd+CPdLQzd
GR50Uf8a7DaCdjTRJaYbfBfYN/TWuU04yh+Pd5ZIRbbVTQlVgc1UanUl2//Gs3g7rcGtx1cqvFH3
EQgg+9WUVF9Uxihasvm2BQdvKMS2hGh2bYTp4ACH94ZVGAU3wHIwnJMPzky1aWXXuCss8WBkly8Q
FQ7v7WkO7KWWZ96lYyUf64QX83hzGQMruQRYK/+m2/aqv1CYjFPZ6BoIAGNrtpAQroDTnD++oVEO
9gL0U6v30YkKVkJEosffkH8kJ3WydR88hDL/kzx5Dp7xzUkE8dmpyyIMEBZ3J8YjzjedjrmQYpJs
Tcun59k/sge84raFlA9BN1VKAUf4E+u76XRWzbYbWPkWELFbfPR8U8KcoSINOxos28Ymj0Gc6wDC
LIx7fMMg1MCOnH8Jiocv8qVyXm47uGmYMsWI+xHE16Uh2xXkcWoT02NOHZem9HT6DRZCH0zXwrop
O0hy7k0oTihFBfJPQPbFzfLctNpRXw9fuC5FXKbzPTPAmgzO57i9ixX0fD6sfTAryIo2TLQuOyYF
iwq2CZEIyuCCjMUsHEhqiutxjLwloBisWiXIiuluw7IhpAxY+y0zDjZng7BZpWDGC2navn+eLFV+
kh8UWKi6SOac4iEyjtfmig0urEK+6VfZ/MKwVTJsG+hnloNCg/GWKIOWvYH20cJ+wadmhSG4GTh1
BHCBCbPvlnHqbuUTSCwiImniFevGY5mwQYdUR7cPRdOnOKVVO2RPn8rcw9yZye7q8h0Qgcv3YCNQ
kuTRH8fo0ZHoXLWsrlWAL8OR+sFPWdh+zFLO5h5tokAB8wM9DmtKqjDixY2nXmmMYohjMhUFEngc
uuEU/ZpVRfnX2bM6dyY/sSxiGgk+0FdUiDa3jm8/R9LbcNmbI58b5ss5Jk9S1gB5LCOh+bB9AmNs
l7rz8MWhM0LLJV0nM6ltcxlAWmy+jxtykmo548cB2Z8oV6hIFEDqrcfy/jLx5tl/9i00kZJYPRTL
eNturSRwmUV1a/1Cqr7MKLaHI+q2gf/hZeqflM1w/kNS7SieobX6xyyYc/wCnS26vZ4HEXFJOfEO
pWWLxeNafZ0juDH9qzGliu4feh7iFLbJMVypr4knz5pJURE34kGSsfVGpRBA7b2tjCmrmNLBPBzN
wyfFWOy22jjbd9+sHuTGyeNZ0V8r7aBzP4PIoRQYqLm5Z4bmmlfuKtOj3p3cJ1+od0HOcwMOwGgK
esSkO4Aqz/lS+RnJ18ziUf/CcmYo7SaNjRQnDcMOxkeX2Co51HO3kyA/QLkFPR4dlc8wx/fvuUu6
v/UJL4VhpzJduJ2WlzLgEwswlayIfhd8hitmKr2xN9z1P9/NJtCkQvdJTsv8CAVAFk6+TY5Beo6N
v08F1XR4H+0weDUDs0AqfhSaWAvVcewrtscYtwKGKbz3TGgyYdcOVH1cE57lYbQ2kjPDN9tm/HhH
mm4KXMQXKQxuvGMwAoPxHPTcctIFo8h8dtfbpolzRzzAC3QUBKRuyZGMP28yhcvDxnt0pvunn1ka
kt7oXuvrNiEd4R2ieFawP0EtPSQXYMwOCM3H4xl2dng1rE+Sro59lODVcub2lafRR0Cn2eVIrMO7
2OqW+m9DmW2zU6osDCOWxnpdHtr/w34f23+981Obiqin9QKjxC097VlVbEI5XfrpY7OFtStAUguw
9cw1U+wWjjvrGOH8xVll7c42pvlrwao7ofU/FQuvLaGaGObaj0ifTfpaBG3YvAmqio7SftQ2wVcb
AGxwzvaFXYhbEvBAC1GlULvg/u3qF/QJrIdiLmTv04MQGKw8MoCEbG33vfxu9epBJOW2IKaFPxtt
bINl/EtExy/8Mr8gXr//ShGXIlXuwgj5VdiJaJsYCa6SKbjg7zgQdYf/WgwRjGVWv9P1O7VKv0Sz
AvcmOme9TWzyBOWi4EnsLV4E3pV45DDNuKyCG8Zs7Y8CtbqBNVVD1D58/STkJEouNVXk4H5Gz7vJ
q5fMvepVsBwZvyw2vpgkQhGBdisDH7lTDfW09DgTTGg5WHlbxDgz74UtVjeNRIcFZE+dCoHSs0+M
xSDsMH+azrQkK1iO5xXLVHdWyYhbA0rIqO8k5XU3Ye/x1w5Vr7FY6uZhIxAOFyam48XoPVGk3TP3
qT6xdxM9FxlydEPgc81RdP1aFbiUiTLJGVp9ZzXyLrMa/lg/3zmaPc/9SFEIKp+aRFFRhPYLHIgM
9eu8RL6sZRyTIGMTuL+wtEy3AggbZShZNVkn818tfS9B8/gFATcaclunCXkOcpZbMxoR2O27L0GW
KHfpwKwMj1UhpFE6KKRUge8MC4MMFFYIrbCALwMCHaI7vN4kZEsOrD1dmihdSfZKJaVAQN0ioWkz
z/9k+N/wHnktb5KNsOWWavmw5e74ZZH3IvzG8KNYl2SbjC1M11wGGtXmUoPvTF9ZfYT3cJYwr7fi
+498BqJiPSHLOBp1M1d5Xp/hW0kTYFQ/BGGd/K+Jz3lh4GjC7wD+OmeCH4ozE6o0U+vV8Z2v/0od
zCbo2gDNQONknvoI3IsavT7Xd7nGiglGza3majiBJ7Izb32NUg5EUIiOKE6opuzm01kOkyVDTNNS
45/NCLmU7aemgF8hYdy6zKY2BWTopZHzMniVeOH+x7nJ2nt0c6VYgy6jfVhQyh/+28TBxfXWEvt4
tzqwvz0HVSmWZfYNJaUETiTVkHu3YTuQSURbS2vJd/m+Ft5bDt63mG7VU6DLpI2WHLUrokTdh06k
HxfHOfXbcy3DbechNd0DzK484nQr0FVGS7bh/41uMI5/0TRf5HXp5Rapv4xr/sj6wq7qF+IL9b3N
ZTndemzRZ/IuQ+yNbhGzwdFvcEHBtqiXgaM99VsGIl7QJEzFSehoXiByUbPSoVuEC8aspgAoHiVj
/jLXHlIiO7oetlUDAWgZupdkyYQE6xVKKmpd6jKcXDAGpK/eJ2Qo+L64Ik+UxqKTz7miPtzxNnb4
zpx20MgNG8SUCMrr80Y88FH5S98tTTtWihWdoukEvmaeIfyQougUxOKX8vTMUqdrDKvYmrk7b+2I
AoR30FfCW36VUe9hEOIm7kfipX4RhT9fGp4olfRLN17GADWn8ZgcS8Iu2Rfbd4+J88yHAPri8yY2
4y8sYsZhortTVcrU0B9UPdJkbTntETjDSRCMwntXynjzZFcsdXCBwEpGwOM2ZJhu08v0fZtpUCcJ
sYU6zr1QMSTFmsCGzWmbDRQfAo0c4QDblbGMurLIf+MLycfEClTlRuQUFSZ3/AHPuMtxaO0cfUa8
nsdJ2J6Di+fvA/dDwLcqXA6o8FMOn2G7w8IuqbsoUU9UmQkKa6qy9mJEqyrPfOFud9jWxiIM/kcg
P+sB7R+Ek19XPwCoXfWnDzdxFckVa6sf5e4FlKhdt1Qy9LcYnANoUE5b76+lKVM7C2mFuNQCdg5x
Oo+nmNgMTNEy730iGcG8pyYfe9yf036+wxWERrrVcYR17jfjJOWrRkGimcrP0SZmPQLxmBVz4q7B
mI4Qujtvx2e1pRMWEnKSf0cPzAKZfCf5Ktbe72lRW1tgeRCxdDpgsk0inZivsc03KvLWwJ4Jsg1q
9Nt7UwdAh1ujqpmX84hjeqBRffx3YjX+aBWzz2RpFQgpN7QrcVE5VK54kD3wCjm4DFcMyYxdKNVW
DsjE1ePmXdy0uEHVbB/f50L7mmtfq0knKmdwP8FrB+Obc5sQtLACZT1+lzoo2AsYUxRBUFFmJaGd
q7MC3Bp0iyPu4lGTFL4+zIm8zH/sMIgOuRJNm5i2iDjp7IJL0F7ORLWVMF2llZjxpTSYgPpjRBUb
j0domIZiBiHrQnbLPowe2i5IUKv7+ornhgIe8NHktlBK83ap5Y3uCHaBq/3yMU1L/IZ5IdFVQRjE
EoxzMBUw/ObGvxKmgn32gAcyi0WoT38wKreIgOskvF/ifibT1TDxEyks5YTRvf3N6MHjtCX9e+Su
NkLCvrTLEbSDOVedVLs8iIqpYdqmzlhBUu/iAXtfk9HevBZhgopzi9GLGhWpaekGEZCqLya+Li2U
VFSEKdDdHW63VcEysrkOsmCuzysVSKFgVJXvtyuUyW/LEa/p8cnBNGdufW1OjeRjoXftQjW8JOSk
Yh0ZpU2sIE58a6MB8UdkuLvTh+LtlpWNH7ECfqZy/iKoHIB6JOvumxkRd2yBixCunD2vFxAdzmen
FHQrAF0Ud/ypJEUpOjaC51Pnta1sNHkrtazSpOmbD0sjGpg470Cenlvl5KAolqViLoNRYoAZ+49q
WP58xugiQOHuTS/ykgLwZ7/SDXkyqCesB3KHgz03UFRHoO0Zf008osob+AsPiDa8U1A19b9DY1OU
Z7FzrRYMoA0BAASLQH6gtpEUjE5P7rlPbdjBXIpGIWkTAi2IzRQKmeyYmC1nlePL3m0MDof3/HHi
zbLwPyNdVlCKbtCQo6l/z7krhLIsWl9xwtPNNCt3pGIV06srJu0qBWnO3gtI8K9hhyec6gAKQ1ai
tvR/uXaJySQEAPPu9Dei22cSwZlUeqVust42e5bVWB6OM8WUWJBw3L1C6Euix4OVmF7ckz7m9+oJ
RoQ53ZyacaNA4EeOow17/HkUhWsvvBIQNlhtOj+PANPYG9vmxxtKCX7+pnCvXx7kGtHEgzDMV0lF
LoI/+ZHy+t8TA19g20yj4F1gbheJu+KUFkuemOXUqPxWaD7/IpYq91wyZWXg1QEugdaVrlsdfCsf
yvmi76rmEFCsAowc3fGlpMm1iRtw/uCYkpuH+46vMdiFGHc7aBRPXcX39q4duMmCFHYHqzfywL5p
qZDfNYLtJACKPol3TILD1C8U7EIWOAFA8IT9r3yhvotkSgiCW9mZ8hWvwJAo4qlDI2Qi3zP9p9Rc
glw57X4Moujw9cpJwtXKwHxMesf8Ot2fQgKS9KJc+/gFg2k7uLvg6JOptqLiRrevq4NBfbtTvv/p
fO6r2YpQdxFgyib7+1+Y5w5egqnesj90SI1wZJCVbZYgzXzMeNrxiLpyIcVRfF9NcbPPTJrMpFXB
JEuk9EZtlfP/G908y4JLdrOkWSpzosA/LuoBbwi6Dx91LoOrQIsI6b7bkR3jJXWe/hY/UpuS1JwE
ykWaM1YnFiZI+e0sqPJsgOp/uyWb2K+X1caPrKbJlHAVoaMIVgBkxM/lBq7Fb7JDLOZo3O00a1/S
1iuNLgt4Od97RCaUZ0r+ruO6IApK7HfwFdZBBku/M3qQaUwmchpDTMMWwsSqN3MOCXApQ/jhnPZQ
QFbLI68mhzjz4Xp7sLH0HXfeY64P9JfwEvQDv6b83QUtlgGudSKNnYB+YD652H9te/IwCmVnReJq
0SNCNbRW2WkYdZcrDE1x0/Rl0dapOCUe/4xs31i7GrF1DBX58AZQ/E8XM/o48OePB12rDQI+y2xO
LMqIOcCwvReiXKuAucp9/8O8mqhb02PYGFSWFJhZcixuNlXRdzmw1KAFubPrPRcHzhjP1w92Ddfz
G55YUEH56Nj7YSM0R8sOPKwYcgtASO3vC07pWtNNM4p9xHf3pPm/2E1h3toIgYfQhLUxEDrr5pZJ
UqunmhfxoMjVZDeoac8I/VMGykSNI5rGo50EoTd2Og33+E4Mm4YfSYLJbiWAYp7SiMBEXlHL+WK3
8vdVH3yObbI7J+d8R6rdUjnZlvHawOa3UCQn/z0OkkJMeo/74sjn6KriblOcnOd3NR2MXmhhevaM
6mF84OB7+OsIoybvZm1K8dVarqCA7GLGr0p+e/VS5cscGEUd7TYVZrly5Q0GN71WLAFK8EO4MBEm
+qjYFjqiFsfQjr6XqUmiqpOev3x41sQtctqVUlF6K1OLvv6L09yYxrDu4jzTgAZ0VBBHFxt/Nvrk
xKRUbJ+npajDcAhas+kb7/IqrfIQkO1L2/sv+3WaChwDMQklU+DT/xUD59SiCKI7duAPxpLPxM9+
wxJBOKCY9HC5wCR8Q/P23IfvjotnA6CBYfCsCsnjy9Ocps6lVkpqBtRX82xnE6HiC8wChspVgMkP
eyV29p17TOnm8Nvh0reVXGPhccX+b/fi2NqUZPGn8t3HdVa2pQkLUDTUxnKq57AO3bWqMk/yvapC
7oSzD8YC/LNIymmkNjUoDRNk6PlMeS/IoUD78UafmszsJrLOtgx3QISXQX1bTD/nrVrWz0fXvGhc
qMYRKveegkQYcqW/qJ6wGe7nERfbiHYni3nhmaq+m+Ur0xUIbjeVTT6YJgSsLJzS2moPtmwiBHb4
7rD4cQjF/r5Khe+FDdfaEpoyPH+mzZ9ClFF4NtpklrffI7JAuHiEAnAdnMI5uw3lGRGnA96b3PUg
YQ+w+bQNTADmjzj1sBsUlFxNVSyRaMZnhjrU1BMnVjJ2fMvjlUXR1km6UKhYjbXiBZCSX6zPaKDJ
qx0zIPzx/XDfiYJQmI6y4/AsJFyaEjLsXCsg0RrdZaGj2DtqMWmNuxK4vpEB5RD1uCuQfErUFTsq
wOecamRGGCz8VPpuBSxSQzQGqvHD/3eq8jExYcCtwnRkxF1xgaeWwsygZSDHAmoqbOh7W4Rx/PFy
5iSpZT144aSeaKaItpYrlt/ihQH42X7Ln/CZr1B5aKvVVbXSW4iJjCcAI/xpqT19KCydVePla7gE
48/Uq1ub20aDDrEJxKj3fi/hi8JpAJenzPmGq9OKB11RlTLic2/fkn7WW0ohn6wEuLh3jW9U6xp0
Jc5iLcSEFI5uo5TSJxqs6H4lrDZnAmktv38pD3w+Me2N/hqPrInMStaVp/dinQM0IOopiJxu0ypT
9qAW2itUvU0Oh1WIL+rzE1D34ax6fxJg4Vlt9o+YThcwT7AwOBW7HKiLdyLut/EB1BM23NmZOdnN
quJBQseeY6DDXX0xX6h48uWEFhYaYFIO+7jlXxHQi7qlv1ebd3KyxUSQ1jSbTmehawwsYD3QEW2R
mF+v94VrGWfKp9yZ9J44FZWNFOEkVwobppk0Wy6/IQ55UqphdivnLH6EvYihdVW1cfNiG3Z0U9RC
Tni7g+bb3UjE6WBrMdeSUuRSQqK/AYrB8OIJEMtDY/88e7yEvbSM8sOrNTadQ8uZf9ULGxKPPDig
goNR7SYZD8IxUQ1HKJdFRSP5wB1xF+6Ix0gg4E9WmcrlJuIIufMOqgVkGN7P9wd1QOXbXJwC6n9S
c65QKBhq3mwWkWyzf9plVdZLB3/arTc90/k+2VANX60WWbgKH0iA7tvI0jruHExKwIHqIoRWJ+rA
1+JNyfYpjzS6IoL4HSFyRnDH8kOs9aLLH/k1HdM2PGRUpfdY7XzEXCJYGpMs0d8D2fI17NG97kcm
X1NbPBZxua8MF+2mSu3q5i+m9JJuwi1itlzYF+OJPnJarTwxISmOxYf95L41pfyK8vqtYlOWH2jk
FOuvlnLUkNB0nfvwnbGZdVes20TyoC/o/MKaYmEfLXPPXKTU5U34vlMSDzWsCw4oogVKtJu1Kxfd
Z88VI3ZGXWzGnEiXPF5q/WBddMsSOOUOTrJDpyaTNFk88++/ZQTIIvg7RpTV6TskibW2yG8rEWH5
a+epGui1nB80IIEgTMrQQyYKNWEjJrdA3OTu/elMD/JyD0SNKL3FcIywG4l4M+rrNKYt6qWxonx+
fuxHBKfdBebUiG5hOJ3Lh+/NVUnjEl4erh7qqHq93C2eO6FU8iBSoJ996Ezxn9VWLu7HOLWipcfu
1Fy45/5JxpGFMVrSBmi+HyydT7qDCsGAHx5De7Lv09erh/l+JWGtTDAuIiP9PBDbm+WkwW7n/rRl
5NKLN/PYEbXXvzEIzckn20D0HD1w/sDzZNpZ+z9pfvgV6Jhm7JqzJZRkUXE4Hl0oFBtCQjkWUKnm
Uu792rfv+LLHEdNLt9Z/coyolzStkZadhwaJZzcX7UUmziuWQKlD07p+FFNXwY3jhTP2aD23h1GB
alpxk8N6WXt7TZTUwepMng6fu6HXYyZFTnR9p4Q9pQVjPQWCG6k2yqHan6//gOI+AXlEXHJQwj0i
R3qeYYrHzTEdwwXY0JjcxcYT6qpdL8cw/u//FyMQKk/PhYMtpapyRA0lI5LkteV0pJnp01xwVkj4
NbqjZmEofHkVTsUMNmEZGxanfMG2ubz2ndNrMZV/HnYNHDdad1BZX0Hzgp6MHJwpSqfO/pvqEt67
EV0k16NYNOFjUeVZXQ2wb31PvEOhcARhzwmx+CUAgOKOJmUsgLoat4WMSn7/WSWht/ADi38vvuv0
rMACESshM/awp2su7a+OXHyXoPypIaQINOeupFSmhmt6Qc6X/u6J3nkPsuPPUn0B7zzPPGAYL33G
ItV8d/9N0r8R0HTgs1sGFAoyhnRSvz90vL9tVSlOGfjl+SFI3s45JnAsnmWDPdiRpL6LmcGuFYue
aNzP9pM7VoyPaNraERATkryw7X7np/+bsn+cO/u+byCJQCMRmFXG2eemhPfTp21iC1Cp0E6L/D72
kBj1o7ho21z5AqgUItIiph2Sd/mOAeOnSwGogupIbazNo1BaeBMISizKozyt0Au9u5+XwhamrQnw
uo9S1BG2ZxD6FFEDmz4y3k79840/EpyGdvH/d6xv1R5yCtfSpyYt8sLsklKGw+NZRPxeQnVL56wI
43lICa392iFCksEcaZRL1x3pNPp/A64r1xjr3RJnLLH/0PhflTOvlJl5NaUrbHbGegVg0JF5cb/t
d+1ubo66rIKs9jPH4wYJPKx38QFy0GkXvwB4yBgPkyJBGnRLblAyFwoohLAuff3GL77i3Yu/4THD
mUDkbGk/H3siurvY944D5+VBQLMZ/acaEVWJLOeuYqNkC0ogJNrIfpFJ08VGqXUKYDj06kYkgoCc
EVpT0Y4aEOnfK3KxklLrD0OQaH+axEUlegHEUHbKu1Dc8cpQWntoTdK5TX+xyKobTvKDc3D8xLZ5
/ZG45OtvK+9ARN4KkBImv+vnIP8AhOwWgEMqTXWkgZMU95vA0bUCd2kDTJSSEOztA8L0VfpnU7nj
3jcotl9HqWmfxrF6cUrw4RyXVceaJ14FBr0PK/lJYmv/TNCQ/Qec6nqOoBvXFQND87dgysyojo6x
jmSEcd5BisZCrIEyGG689a8lfN/Xj2hq16GnEHFvulPeTWkMDyVBS0glo5fnQsgfTvoEfcv1ICFP
cuqPUjFTdntQyr/haCO465N9H0IGLiuXDP4W1OOlv4pid1QcXqHI7blpWEAceoD4qz6iOhAuKHUN
GHP3a6zgGz4/yksW92S7ExsYE62OSx6glzEakDC3WIe+QaH45GD8y6lXvEwWxg5cLB10IPuUZ8oM
R8ZSM4y2wv4c+EGz8f0T4Eezv0Lw0LtQPLLyuxRnN184zTCYitC0W9i30sb34OkH8u083cCmyy43
002em6X2olkifzcy3mJGjbDf5UF2tTn8DXIMkR644O3PaCLHg1Tz7yS6i3TlCUY2UDKzzdBhn4+s
Da4u77Ek1T/ccjwuRJoDWS0sTR1lXF76lR2ZaD/dwA2dwDJtEjzh2i0Be87jbfohC063zazukm82
QotmYCG4Ko1Oq+O5cnYS7o+6hTC8k7ldy61YAL936Hob6cheGv8SW22Zgnejht5KXkyieTqiuLik
M6wKtG6MXDzy8KGJdZB6yb0837YSQEKkct6vLbc6DB4XTK4/bSweFr2+5boDL2FiI0M5mBjvMCXD
iC7vrhbJX2HlEX+FpGXePzt1pa7vSegbr3sy0fKo2PkQu+qEhg+vpmpq2ggafCiqTjiXcQqD+puA
ugfGa9/Sk9QGDXMZxI6eZvagCkhRm0s59sCZhKPtF80ekYBXe16cBDFCNmKrXT0hc04r5oftDM+Y
KOSWWDL4gaRTsyLDu/GV3qkQiDwnJGpwFzoK5INb7VhwfFg+KAD0BBD96Owa0colDUlfxwrqVWHN
utgRPK0yV1d4s9zomNtrzp82//qbD+ycPKDQd1rCzeHJ09RUKRnBuOFaTiQrcWv6KKL+p9YAmJBm
4viWq3MCSG2RGk64CD8pjaFuF64TZFWgaQi1LR3NCbO4Xs/1QDetsMwcOXwqsEVVm5TCETvr+mop
Im/6MkNYFr6Q7IIy3UHTXhWD0gdLJ+Yl+xhEIjS16hpyNEo7HHt3bhc3HYaIQRotWpJHhKB83JQY
s0Sq2nLx8gXyI3YjS1qvN+DmTrGrjDZtC6i3Scjz3c0OLFE++PFTD9xb5Wxeh3C4IR2Ca/+w+Etz
whDcgCZx9FeIIPXYY+YbAoqbunQ/HUcXgivqV4bIOdPZD+5hJAZHyvMo2esMXvCGCvEtYzmis+w1
Ob+dKhKxjFrRacaStrCRvAISnSA6iajNa8qgbadKz2qoJX5QtQNsvZreAv6FAH2UtNlSa4vhJMV2
6fcmmjCs4rp4+Dd9LlSgYmzJlMKmT04aZM/E0Y9NfcW0fNL4UACN/AC7hCxmUptWLNSLBoG4OrBH
VoPp+sn/fv6b4PvtJKuthaM/KsPIDbLrSEVsVVOhWAY1JpVFgj6AAb1XR5t75g1CnXA4QOSjdMQ+
GIozyFQA2GvW712FMq0NV01eo4znRPzgj+5MIh6Ij+MeGnS9lFA7MLoNazXpDdgkDLiS2tfeLdha
nUMNitDV2BhoXVmVHdL4smfB9IG5iiaZvyOY+a1wWRLngabJxNSdPETch1hsSGmK4jRoktYG4tMy
XNGFtLTce+jK8e3XrXV4kgdDpjlpxTwddwDYT5GIZ6o4M8We+oWGnd5oQ8/yftuJI8+EfzB6JgGS
tIpO73T8VuBXfx5V3Gl4NVPmv2SCyt34V58T33gsxQK9X9PpMcnuSW2/WDao7CVVUqDGYrN9Shy1
GjSAG6hrHawZYh38v+PS/nvo+EsLjl2+PzrtwIJ6uPc5x0xVzTiAaAlwhryiynCdiH520nTrDq6G
02S4UIXBv/m88svNLi7+rJ8PLJzR/JmWvIyG6ZXIpYpK7Zn0tm7rSXfockUcawl6tHtzYjsxPbhu
pi1QCV0Hy4+D9BzJqk+HMFWszPH9/VtLCbua9Y+Z4B9KBKJzEhmGtANiq745TNcIksYF6hQWoix1
UUzYV4C6SimWV9MZutnd/ZcfeXSXX8IJiekgth6zknlj24k9yI0+NNWn3a1EceaQ2Ty/FF8q774q
Yf6GzUg5sX1v1juhDZSb3vHwAvVAqvDaeLpk014hMcnPdJ0vJhflYa8h83cVYR6EXwkNyXcH3JQn
HXbZj5aewbrcukiP120sYr7reXuJwTFK7GVz/DJMHb1UO64F2L+xarC0o5+7ODE8xuPZ5l7QKMwn
IdHzrZ81vJHOwFnLYFx9xlD7URa8A0oqAIjPxwNySFqM49TKPu+0YgTXS1wZJyqaDFMgWVJFT/k1
BgnEegWZLRDbHX/cg7QPP9Pm3HRMgh6WDWa5gH9ni7uh/Z+WwU0IoPzXc7OFbTn1lMiThReg3bp3
vi9jfMKZn2ghrkBdgGIITsacwHjscx1EdxlApu9n1XJaseKk/T4jYkiqbl8jgtBxU59XWoAk5aQ7
ela+QCk5Uzr/YC48BWaIpVjrBVOYQLyNgPl/ujhQap/IOU8hkaN1L8/lnXNl67A+ApUmJXWfdxir
Nvm4oXxkgut6d45JtKAo/kIkeZq110Coofg1/GD3Y+gxrzEtyoEB5lVa6V4ethQOC4dk5jcy6sVU
0lMBLEmi8Ydt8p8fxFssFaXbnpGvCvqdQmKrqtzM2KHkohnonTMYJudghzw2DNbbcsDECaXAE5uw
K5fFh87S+ZiMXJf3zNbkAPZijQtavi0tLNEiGcStkhb9638awJN4Eh/4J72v7ALkPsc6ZaehKslY
/6B3ssf7nEJacW8QM2+WhE4qxHITDxRtwaYSTyu0I1mzn6hGTdIF3nMwfwBZz+mUPYe4riQBvUMl
mxfdfnyRU6ZtO+45yn7Q+jj5wlkf4mqcNgbtIFeFMd50SmO80ZFX4kb6d7NyHjgkdBH3JHcll6q1
yXYaNPu9o4W0PrfamWV5a5x7SYWZEP8+ifiSEl9EcEg9NF8E4Ph/jKu6AV6KAUnD3HnFIc0Ew0S+
XUAmiQWW4hI2OT3T3B0hNHu8hOwBzbOC8sUxY18lyuvdWu4js4VkcdP80dtyWuFcOfLqbEAp+73E
wlUHHbQEzqCbXVo76ExU/d97x4EumKAMOJKWMShCUAa18l/h0hAPur1woHOH1Wq0SHGkyohPeK2g
zQ+RX1XzxrhS4sev1UxdIIUzlSenBEay9cIy/Nc3H8mbF66rW32ug8Tc6FMkN9TW78AhBoiNbm0b
iQQBuY5dZ3BJHY0DDndlYZvR8ah/anXrX18werSV1yyRitiPOzQ5+R4yXzoooJ7sGFmJ/Y7U31we
FwXG4pGp43y614duK/Af4SAE+agsgddfz9bXH9nz2rF4Y/6pT/oZ0QhJTl/Dff/pXu/D1uCisO0u
XSWTtQWHgzk8hY5iZK3B6SB+5OEPGMb2b2G6igH4HhDR3iD8HaIOemRmvx7xAYwjN5OGgCQbNZs8
WccKoWQm9poK3L1b5eEwgqU1ytjlrCvzSoZyxsEXoai5j9WP+hOEvHB5jWvhbcRWvjLdJtS2G440
ac20mTcPRF2x67CXppyKCbV9odW6PJfAqttXeZaf+o/9Q9qZ0cjJbw0T2+cy+oG2ArC4naTmL7+e
NfUntkYqMKBcor1fFZ7no5J9iHXL5ffipodJxVS1f/+e1+JJ+ARI3LD2esdp+cG0N6xPdmLc9ABd
edJiowiRVTTkc7LSibbPp36HIcg4GD2xw8MINANM81Vwz3xJPUniokn5hIFuUl/FPrQsO3vaALdS
LL0CkWsIXdbFn3CkCuAZoXTdnCWAz1VjR+ioeSCSsSIaNL/B91Hcs//oluMkWCl6Tk7tVolwP0lr
hHr1OHHVHjoEWsskzuKKbT9SWY4+N2oAMJuhx/jIrog9b0EVOPR7eiLUANctuz8T/GJfgKsO2eSR
2hdXg1/ww8HuVCHZYEP4fRWQocazvz5uNsq53uM2LOv54ARjywOk5NAunW9fC+asSDUy7mpL1IEg
hqnezs3Oac8by4BKTeZAs0giCVLaJ2RWmRFAfRkipyEZisf2ehpnE65Pqvbn3Id8GJ+98icaH/YF
WbINO+VaQjYntct+aXQGwCQPwkL4Qh9c7YDjJVNg1dXNyzDXLlGtr7PX8Ww63lATBTjqP692xtC1
Q3sFgG2t9pGa8k/m9v8Zkw49Hui/G6gCjK0MZy/r6eT/P/iKW28ArsL3s9KiY9it0Vx0IaiGX6WH
WQajxP/2WPwAWu/7KXmP9ha489sj591rQ6sFGABuodyYkIjn/XtHnWdn4EWg1nRX8dXMpFM7KySA
iRUGcV27esJ1mPh9A9UclUGk1KfUsSCoZ6lkeboTCzcPMjO7dKQHpZgJojNCGY2Vtvc1DIdV/3lB
LvTxg3K5+sf/BuVvfpwxYRt1UuGATuCARaDBWFK6wUFUEKnRRTNLOUZydkTe0dZbrBY7aTO4UDyM
PulPmbWLuQ10Novj1RaxJgdO1cVJDJgzYrZr++okIQxUQnyvLdNpB8bleJkrcWvJwJBR0e0l3M6y
ZnNw27LExkwdUW/jAU3Z8G7KGloGJz4oMhjAaSV2smZ0bZpg7T4dyRiFMaw47ftm/FpFtKrAAV1E
MFyZ0cECESM+g24XLC9euBxnHDFXdTn1iwog8L402TZr3ZdZmRErwHzqRDWLSdN7XBtnHU4ftIPh
E9/fekwCCesCztLHIF9HUSa4+1VSKcJSrfLtbNJuHZYcB5BOg25LwEusbe0WFGS7XiVuaLlnHO2o
+v+I6EuWBg8hibd2RC/YGevl6f4cZlhT6Z9lvMLWHX4vPCgbCqysCYfFjkDipznhGiTSTdFWXPT3
AoyIM9lTF2xcEH/GkYQz7YK0fRNxfP0lJopJUlpM0WiAAV7xD6swSq0Iot8K4lwGh5Su0uIRFhou
ky7leoXCZGglJLhZL/nffoT1srGkc/RM/HJSkaUexFx68hp6nb5Mmm7zpbbBIYOEAXDm5pjISSL8
a4Z5cMRVK0ZPi7OPK5BhTNR1pTE1IVIEWfXJCC7N0J86vPj1KU2Gq9hHN77QDnkxlp67vrvXjfmL
IuDWr4lzc3foun+UTtSqHvDQyzMkrzrJhMQCtWjzBHBMmLObIUbQ9Kw7Uh2cTiWEztT7BFs4KHMd
FFocBDZRH//2DXG1O1zT8EdHNVIn9KZ028ZblS30ziY2ELCNhPMpcFixf/V58PYFyGO+jO7E/VE2
ww6iu/FU/ftN7hkuOhdwGwH8gPMY2gUfmbeoVTeg6Cj/zWFQ32+9ARzm4B+x53ep2wG+3yglCvOD
Ob8pvNh/bMrMCSh7CW1zLHr/HEJxvM5jOzDiUs+LuB/HTUW1vPAsWy1/MB4V+AuUVJ7JyR58C4uM
+fIooOTJR87lD07sm0QHY1b5TAmo1sFB4BOoylQh/TxCsLPMIXqqfTHcErFWjX28l+afvxR6MYhP
Ks95HGufQnAD+gTNBCMRcTFY54vQLBh8+w8X1HBHd30cG5792nab1Q6hpYiI7Ja/hflkD8ZNeGYV
cu6evzWdBvGgnfw4aVIXYeuKNuzTy1wKzMbY5qKyNtOxbC/814DtaZanZ9xSkhniGlv7CE+U2Uuk
D46mfLIkpF77i7I4ATWyez5bpZ9+h2R9G8YuTB+hMDvXY1D8PZt+q2alrnZh7xz84ZdovXeq8SyL
uEVgtuwaGVIngi2lRuS1y5N9csOaKv8lgDfii0Wk5Z+N6nDJzKMbcecubUNORrV+vtBq8WgKNA3p
Yujuv0I/kktJcvlAGxxsbYevil6nGy4OCiPVhQn02Y6CVTcK0C5AlXBlbCIlO4K8VXmXFz19uwI1
yKFd3gLRT4TodWRknDgJM3g2iwRnwb0t/bzDEu3x2f43WynR57bbyoAC7/1NYalDocoDZXpSqHi7
Xm0q6XJnB2lXd+1cRJVzpsBATz0E8L9ZDHh169y6HR07kbs+fWxYbd2AtUj9bFNrGEjUBKXkUck6
tazunfZac5u6ebeN0lQavxI1Mpx0rzI+DbWq3g9E5Ri46HUjbf92cHedwQQSQrRjYUgWmYCcBtLb
Oeulgl0jv/JGAUNHHuCCoOeUDBy2nIRNoDg55znCJJ2VPUfPGCBDW8yylyEmoBCihnS8gNt7kVsy
7PfSz3RnOnAw+CGPR/ouhLnClzRqUWAsoISNY17iNlGIVn3vI1T/5KsY60rc3rzzKQzN4YZKiYac
chJ+w2tfUMgKXksfYU48AGYhzLkzfR5b9vjVt5eXdiLAQB/w5WC6PNm+a3GSgY2L1kOmjoCdX24T
bl90o/cZKv3n2VzGkvUIT6Iq0jQ/uMRkfRfWnicKTrWA5pmm0vLGG5BL2wI1S+O6cELDwn1GbCYd
8AKadThq4PqYanZdNQdNWuZ+GfHLUwiaQCJlIDrwWWoKzCnF8EF60YsZQhplzZxojc3KjIkxGW3P
lPOgTTPznFtpq0oFyWBPB3tFnILd8lcLaI4k6vEk4toJqSstG2Pa0ra/2TaYqwg/wLBpOI3cyDNw
/YGUuL7uMwlTfgrDu0Zu4JEX81Le8w0qDvRuXH/VzDcmMqr9F5j9Hd3MX3yB5Ki2lndNOvuR2SPz
19ikzBf2xMQMEzJV49mFcSzbvH6clQ1zpunV+rCqdLmKJtEGOoiw6SUM23n60CIwTviFyvHo8/oU
oYmzJpkSiW6AExoaZ5o7Ftthvcaf76Bh5OjS/RgVytv8i7P4LSdDSR3qX1/NmdSpFhMmRpbjmfcu
FQFZ8JGRUkkcjZMoPm1MnjkzUjXfG4Ea5Rcy5UFWC/kByrKSKcBtt/13115mOQ8Pw+LNR7PgRe3O
uGyami2J0SDa3cbWNjPwAlH/8wSu5e7RRg8sEHLC/e2MZrDEbbb8C7pg/LGWEP8grG9n/4zFMxBX
fRIHfW02C/5dbVHDmhmqdlrOg9oBqCbt+uqcPzQOSeXVQMhGIYH//AZ8aToyj+fTMykNgVj2t989
4wGiWJUMyG0VB8bBapJ06sWP70Xb2SJBQvZh3dS9vzVjs7sQFZjFflg9SMnDris/T1nkNkMxKRT7
8YrUpVcTdUV7QRQU7axM/weSTI9YeZxdLxs8yposxHiTn8YORA7TpDiHUI+pR80WQD0mhc8N5DPh
IiX077cTIXTYCkBDCvcA0AzyZ7DYRzmBkQH/E0UPi/7FFVv3Ag++0il0oErDvJz3nmSAnxAeed/D
3g0nCU0RGa6t4rugTpOnYq8LdAHhEfVf3StCz+hxX0J85SjXNKF9ReSVdxcWmUgzgqDpiPru4ovE
Vhw3wBVSpLadlzvP/jj3a0ne1YXlvJLhBpoUN74JS2S+CJLaSFrd0ossz2s0u3sF+2AZbFS5Ebdw
AtRZYq7nzd90y5MBkK+jgeNMyjhZF2yvDt1m28rmrTpCpVo8jlPh7sc5Q/AVnmeCicVg0Dwmhjwf
Sjx8bhYFaiA61ksfJh63bnynQfnE3Fc+R4hp8noPjOx0hONUbE5P9R9u1mBdPCq4EtJsqBiPgrFQ
FbjPbMvOmullfpZQfVcR0KfD7hq+cNvcvD7vYnC1qXf7aZcYqySfHmi7nkhmgyHs2zUZQ2OXMfGC
/TDCSs8othKilF3n1CzgeQTYLqA4x1AOlg7cj0ujTkRRbteccnqxkxQoyvt6jYSI2H2blP1MGhgA
UrYuBZf0lUfihRNs5enZ9EZGpQ7lnQCXx1+C1qFSb9Uj3+0yZutvaTL9J752s5t1MlGMsBsqqmM5
mqtFjls8IhFR2UDmBtwwlVEPJQzhswY7w00ZafrAmGAHDP0ymmRmzr+C3UZPCzk01szGKpC4ISyz
OJS7Yw4EDczrZ0istzH9pwZ9ebmzS990UBS9TexU73heNcUvetWiM6t+f+EcOzi7l3b/BTfdMXPK
rVwv4wjMfeWoGy9PBIanqxYcdXCqK3ekTKEgs6hawGSWJ3rRXkyxkCQH++z5lyqK98pxGEqrNgkt
yy1+LiUycxiDqbERJ2AMrpGBxjWDVr9s9z7B34iipF6uwnpYIvKCp8781V76BVbgL0Os3Kny0Scc
dfjOpF9Ofb3m57LOZzy61asyLFUrsmOQFa60Z5VvWy9vNSuhahTePyJsm2TNE65iM/6Tv5608sXc
U4N6xSvHSEAMG8D3PQoENV7fCBtSZ+dTMJHs8kwLyg+ShNJDgWNtVm/Pgqqi7hMLeWiWqGKyOW87
p9njw2TxKrybJ8TG/eO5q7eN8+BVVlI/bAGskercSrI0EnvssC0fzwapzsDq2XYyRwGIzgKJJpY8
4+VpeM+ONkZ6PBFquDdg9rV1jwv5y61ptcN0yJG9WzbWFPP7DKbyrDnmvuG/WsRYV3CAnQosdJnq
N2sL6RvtfsIFNEZADXUpfpKRu3z579LtALpqom9CsjN+AZX/T8BjcXaYP30/3yuTa+hk2GnaDGkv
reAW8Sj2qoBNDuO75NKFe9JlmQLqMrBZBghLalmaMUETUEJ2S5bcTaGAgjcPDMyfwwjhBzVAKlwY
NpIQdaUk4HHkQwGMmU6WAl3Z8R3TLk2FRfHPU6irw+7zlxsoYCnJ4rRs5VHv9jBqDWRjn44RY/1I
0jPu+DbDNkbN83/m0FfQ/dxH5t3jRO2NFg8vg1JqBXS56d3clkRLBEVKNN2gVF7oHdCES+LUSBQs
LrzSN+cgT2ZDNV96a/4RINmHWht8XFhuvJhUpUC/f/BYequZwXcnu097drkikytaxlPCnphHYC2O
2eFiuocA0t5xaKi26uQyl0lXkwy156NCdvZAzIX5w8VLBxR48f6VEdv3EnZEJzyZF0AQOAPThUe+
ZmZXICMkr8odwqlblVs2HGZIgHawjodL07ISVESUE1EeB1w7nX03KUFLOpwT5+nglu6j48z6Fabs
N0QdrplJsxcRwYvlvhqtAtkxwkFzz1u5z4PwJsYXGw0SkrHnugpvG9OOigf79Mhlhr/GADh0HsUe
OcW8flvEO3ust6omLDYCMzoX7jjbUt3uAU0dPZ2UdXnlm7zt/b3Staj5wm5J/BfzYPS81X7fLn/s
CDoCgi1cYjUkwYUsaO1SEIOqRFMJqJFfPsYbHdeIctlLIxzOgqfjpvk1HKuFVLC/KILGbO71ZQrR
7WRoYN5GXuR81VOY45TygA5CGD3HqBEeOvSaCXLvzUfST42QpEVy/xhelJNAuZ+11vSzsGpRrxKv
aBjHefhTboCBGp5PBZLlxU8ukYnCWd8LlK8ReolwsGuInipVgS4qRtwAmPwS/e8EHE8LR67ZmoGf
YfDgs2aeNjgAwumZYHagyW/ss6HdiWCsInFU3+cJ69WyJ3nQZCSAXvUfUvc1/uwbWBkrQPRHy1wg
o74vSaRpM5ld/8kl9bN4DutD+nbEcqEPFdvoBUknAY3cAwGUvND9bE05SDdfEQkpZ3EuZ8AnBiak
XqBXSC3WoGVXTz1sN9k9bD6uWh4k/5EYOIVqeuS5qVLelCaMCNi/tqO9qCFAzcGXyunFUlqktFvB
L1WfzKEFm+2ACYI1sA/8G9D3dbi8ecJ8CDw/xmlMJAJjQEnaHdu1Ha9wITs//WKGe0QARBdC1NEy
PmCl2qm/mBu4DegKxO2NAXrQJsQu5SlUBwEd+/jTm00nCH3vIBhZhKJ2Ni24qt4LtLfpevErXN5v
FaU6gd+TUz3VwrYXFVY4vmRbpp3VOsb9QKo3Ug9iv+yhIAoVX+bLOpvawZuCOFFRZMT8Ek2AKKSC
wS+ePWmUwA2yKUs2xOpWpIvg3DdtdjNliAxIcGXmOyFGjEQP6AYX8DUY7Bqq2y4tifmo4FsmKUMg
BEffTMRwjEU/zkJRibIAffBG6RFcpFRtZm6xKEGzMeqR2EHHl30jPhbeanRgY/14uKPlENMMy3Lj
RHuD5YWkQdJKPftznXypRF52o9JZaXNky9GY2VQpjC61MHYdA11qRW5TnBScvOSvjTfDMhfqkWgm
q9xPytn5U3BjxO/9v1QYK9SOl+O1few2ShfxIAwjgWvf9xReYpWVwKxDkUcNY9WZtK2Ej7lJGbwA
r42ow7c/13VEt6wMl0sIzZ6DYlDOH7M/7uETLjUJkQ/b6nr6zX32vkhTwbmstFQFUGabGo3MYB2a
FHLnrfH5UkyTF1t1MVYF/42SMtrPStNU3atp6bEpGV2GezlD9LFNTQ7vRLxGqEsZoz7cdrawdwhK
UFtQzJEJdDBGhfTSRVj9zXi/o8LKivJb8/PlCOE7K//i8H3fwkoOaQiVQI1Ee5HAEWmBnXDYl3v3
zi++S9+7q5Q0CWwGq0bqPs8L7IPlq0Wi1GvdG+AcTqunGqcXdieZBtEzFGnArt3chEFpuxruDLWx
kA9iUfKEjqs2T8n38j+FmFjlp42osyX3rBrnoY7FJFkTZyxVhHRPC9X8VZDucjBZSQlPGYmkh0I9
qgBX0Y8Q4QnOW2obfbxbhw5IkK8Huby3aVI3lqpaXyhzLkmc4+laRqCuTgNKKotStbSQFnxv86de
0xoeCI7LO7SP2/tlA/T0GLJa2KFF52OqP4KKQf9N0WlHupUOiKc7UZ7cpCM34pKoqivQNg+N4sqK
aHRaeC/xRlPi8NthDY+HxuClr0pIrTm/jWPr1qB6POmq0t3t0X5wLbsd9pS8+smFjuCXCHWWnLhv
hzlf4EepTVOZsDeSwz1Jw6wOlvx/w/ZXOlp/2wE0ctR7ISc1v/fZv5/rNpDMHjOwi8ilFKhXsVR9
zobY+m378Zb9AftMEYupOHjapwfl82H6A3A/dnUIpon8oiUT2LGHXatVkBUxx+BCvvE6hiT9OJ9F
HHGqEpb7ed0uoBHV8dOMFUhtOym/OW4XbCKn6YBO+x2O5O4xaHe/IItgKlXjwhXVBsOYf/6HoSHv
r+vAwBfCmHx2obV3Vs19v+gBils55gJUhAqcZiXCu0MQoDWOcrN8XnTnDVtB7OexWs62EX9pzL4V
BGaLwwbj3zltkCSbGN5UmzXRpcQV601VAE75+XxQ1+KqKouVUWdgTZUQ57Fsg8Vqp2PZsIz4mRqV
ZTEu4EHFnH9Sq6ZVL2X4LP3q8P0J6/sLA8fHUo8rE2l6cBQ6hg1TfS4sA1hi6D6bwvU6uSuC/0uN
3UJjfbqUUJsBxU5AfI4W7ldkP0Ok8HkSVNpq6Tjo8C3ARFoY2PECUB/GCZCSZLmwPS+tN203Qrk9
pntGQLGnXDUiKKV368WJhNg6igS1gsvyROJOtkc3ItadqGKFQ7BsiNqYuvAWd4k1R6KX7ahLQdT4
G0cYDKpXj8q/oI5046pY+yTlqzu92/c2kpvcXpAuBFFlkB2gkj4pFIGHUvYCfVdfFLqjqmwBbn4Y
kXrEAOWtMu/V3VaVJ6uo0XJnzXd/eWb1h3oDocKH27SpOcHunLtjsSnU0NwyU526DlzAIPM1Id4+
UskcI9gV3rEtLm+dg7CMybAQVhs7zsIMnTCYfqObVGwxDEtT3xbMthgpnYgQItSXMqvN3ONeq1c0
wExMx65+eTkGddUY+Nn3vaLgFDQyalU+LqTPbuyNTr0LLgdAbFX0jy5H1OP36IvdiqOBYSjoZ1q4
s/HDnq/UnQWI3rKlQF4X05pdypZTvrqS3TAk+qYpci0kfgLxk6sRPdk/uvmDz9jtnSZl2d6YNt4T
2IBlIKk9GTqW6DvkrsGoxXG2wRtCWFoz6o4qE5N3fH2k24Q/lOIaFWQA46DqMQiMuYH0Me/iCCpy
MpJaeajvQT6Iy4HJIUh5J1apWNNEUzVA+KbjcnUQhOiq1m8FXGvUTMK3E0nJzInDNpHoC75Irpo9
krhJ3KbWl3LoOTd6SJUIJTnzrbnpRn6y6DMXJrrtWPNuj2au2cx1QFxmdQT2qo9yPG571gaptFE+
ZEZllp70UZ/YPL+Dn2jfsLmll0t7O1bgcTV6Z1Jm4p9tM7aqxLDa0jIlP8IKqe+SMwowqintZsAb
3PxH3Wpm1O5WFiQiCaKnCk/ILFn787LWOW6teOF4WsAoofrTUhaA4Cum9fBbO1zOD9MPuj6vGl+h
OJS1DcJh1qWKqHLiiWFEgMfKic6Mb6DZRX4GPMhxMxzqHeZfXBUyG5psxHOCth3sfqJvvJUGWyYj
aVae2r/awywtTUnGTdjhFqlm5+xeDCPoBW67PD3O5Ka6C3IwI5gOrdwh920vzmwiGblNCLcPs94t
CAnNUNfNk9MPGwVE73+PjiRqaTR/RMLALH2h3evkCwAA8NQn3qsOjeCGnPySmTzoq4TRzRIo1pPW
dFkViZlIyJVMcM99xM/Jb7rB6Xk1IpNd121AeXmFqadZLaHkYmKua0302CNp7NQwr2RlIiYp6npq
Rb6PJjV7Fs9K6f37W1Ij5bWW8tdsHzozkeysXegfSqm+QMPQjMGITfxGlQSC5KljZyWMtMc2bMDm
qGGAMuliMmVl9RkeIuqv6qNWSTZtCPboj5utgefdNOggz332aXdcUYSLpyRus33EqUAVCkSk+U7G
PaIwR47cXuZscDJBlOnSy1suNPnpoTcKgIJNYILb+1GtPr8frMa1ADRZjOj5bajMBj8wGbp96vij
Ovf7v/JVotCwxoUIykFu50x3QMqpVakZFUzBp9ddQbZ3EerfjnvUswsVS0/Gj9sElA3GjG6VRi1Q
QhaqD+evcvHbXAauh5of+Dw6y7nR29kP5MLOLSgE77rLZ2OcdEdXA3ggkJ+4xtN3yQDIiLxhoZqp
zSRcHtfmPkGv7TeURrNzVjTheiO8zHFcQhYwjXtuhWy9pRSrhkve9ZEbjMSAkIZRi3RJRidzSZY8
YbEm68uP/v6wuJLRY8pD6tNJetahL3/C+ULMxeIYYz7F/jzbdofw/1WaxRSwHaNqUpsRmvQmiXpY
IEyc+0Ql7pTX+NmEHyfQlC2qASPcKZBnVV/ozQRhbadI7DCKkmyssRXenY9JPYZuh+dsyZbKeTYl
0fJF6q0iyGDlpnhfILrm4RlCjtZEJPZyBaHyqND9dP346p44TO92jvYqpUmr+D+SJwKND3LitRSL
QExSgXAqDkA7+MdRU4EhGXWOaGm9y0MQfxOfZQhUx5AJ0qInjSmJVsea16H/zLqRPWNdugviWqdK
SeqZ5aErWbulIifI125k26xIBeaebMx9fgwJDSU69llmUMSOb+CZsyrKjNluVNAut1LlPjaZyMJu
Pycw49j2lQRnfFqzoxngSBs9Z8Yjck12xvv8MLfJkEi/Muj+L6nDemKm9TlXVgDdrWkM8Bx4UvJZ
f/CWF9Pta1qVpNLJMysN3Pahs6MbXqtWh2OIyxcz+6dpp1xwiMQ8VIDUiFhgPxIecsM055rbQjVe
Kl8oV+el5+eBer/uI6BoslKIfdOXmfV8YQvVi2BcYgRrsLvYEkE5NgRgMG++JFNeUmTbI3REIUzS
uBFDbVV2z60AXGi/Ql6BNrnW054WY5DNB0hpDeDFSqch/1focAN2jPWgjr1/cW6GzYt2aQMOwZ2w
DKcmTzbuZl+T67YnkULOMH9xk2sy2db5vGKfOUmjYJJZOz/iYbjF7Z38a+2w7RI2BQklU9oT/z18
D5FG7ImlRh+92YWWEVoCKe4D4Ywe/SK4dFRyl8aHcSm6bwNzqSIlhZt0ssKPEgVvjRECuZJzWR4H
BzFrHbFK4fKqZKHMI+JUHkJWVBmpSOZ6DzDC3IxZAe0fIpeee+Wz4S4l9n1bxjc5rUcmywwyqRFC
mKIMw89hStV0ahHcFfED7uPgi1uwEnma4xPIJ6edT+g8NLTiz4csMTMpEC5NHL1YsvyGSm+zSuFj
I+zEJ6ab/BHJ1GVpEkUzYcjx04QwBSrpF8MXJWQWd3ApNn091xQRLfVpXKLRk6kBq22XbxjSpvOa
L4NRkfY0sD0MceSKvIJeCNTjkzbmgKr/h9U5oudDZ8DQ6hEOBz5ivpx9ii2ttYrkSFLqzB4ZX6mP
67naaIrBK/6M9WNGBsagpXml5ICQI+jVyETi/2gekTJpZbcV9nU7OrtIh9aN/x7q02NBNe3xhbI6
BoEOmDHCvB3KIr1RfTGmyv9B9TMMYMvjh/wYbgPxj1Ki1LHubR8ve3W0/77avCAPULXuCZXIoSDS
NkKc9iP9Jv8m4hGHysURHklTMBX05aLpNEuro0bqTzi1ddn1mKBWoAuIIvamk22NfXyDGMeTtx1A
RypI8dQdd6q4IXJ441y/YyxfVtl91PW2CZ05IvLFWJncpJ+EIjE6ZgBbPHwsm0bIgH76vYhk0+k7
0CEmpYRFSIq2QEkzJlvB/aMcYiLu0EdsgsSMpzy6mrsWFfQy45oH6YmiFd2chuYx0OBW1Lc2BlSn
Hk8pH7ENOBd6Tw22MDgvAgKh8w2mPbLBTj3VPKm6bllHOScv4TEnit2Zsnnmwmo1unGREZLNjHz0
OnXboPeVLdeZ6S9sotxUid0/0wYCH+jEWe83SFr9rKYQFtOUHrT3TkPzf1sE/O7fTuBJT6Q19QeS
6S08T3x8kCA948SYW9vF6OlntkpPqRHpQRvZ8MtNPnRQt3lCs9GSm1xt2RB7QA/hcZA8oaprLCJ/
qTr6YIR8Z3W4XGgbjdvjfAbTpmx1leSWbCuZT8jacCgtGYCeuWqpNBw74MXlH+NCTcGDg/U8pdUd
Iw4ZbzeseakgDsLfgiDVFveVszWA2t0e1efVJKIti875sdNsleNf/BNiWVjRJL/onsKHkW6xTWI2
3QGrV1kmVqHkCTRpCyToklofLHK4SHxFGvlCskwWu1zXifo4NFHWkJxF+kkBHeE1dW+Ngl8Z9y7B
Q+ZUniyFmJe2aZFN6YAsl0zIOIefaIHxOXm5e19LdMBok6wId6WxF6OVWNcQiGqSkt+fsaNW8M9P
NcNpcqAkjBNl8gpSxJKEnh6aN12aBksXSRAYY8FhBaV1mi0AxUKho51Jf23tNjQtjCCyu1iEB1Mq
yPU+dqk0HuyjGDxHXNL/0xmq8HTgjYOillYhue786lRLAZDxBm5lYGTuEXwB+r7LhFQv7l94r8cY
oMLZ4mHrO8F4anezYSCwNZHSNYHine2RwFZVcxT0r0NRSB0HT2gJrxcBWBWaonWiBIv9fSVKjz2H
qGCM8SZ7soH1cLoEOV2rXx5x/DFOb+YruBMK0K55buS2gbpe82qu9d5IFtERrhYf50genru/vvQk
PtJo85SCP3Bgb4oc2/Hejw9FJP6nussVjSwJssGVE4xefjw5SQ70vnk+VrbNCrGxpvrqMoLltZW3
hVmYsU9d7oFzWUQxpbAETPlrXuhKAgWk06K7+p1eNtB3attZGvzaDTwGDlBroTd9N4G3ACShSyO0
dX/73Cgiz9YePR7Pac5wSH4h2UoK6Lr1Af/SjHJYrBl1fKe+U3yzueR3q4sTQyjUzGu4BDgKHidK
91WPJ6GQ7QXKVO5cqTYbIEy6y2e/n9+CajwJQFUKqzM85QjfgayLUPtziQfG5d/4XJag8Fi7DCF6
hD2nxg3QjTzmMl7AgUAtKn+c4fPlSFnetaBroOn45OiYAIF27AgE0T1WJffwN3qoO0ybSSMh7WFn
v59kjxZ+sr5VF79A/hVshn0buNKE7yO1Y/6VEd8yETDpNdhMMSGu0e5rDcQt3V7JNDAc+UG3rczv
xh9YWU2MrgyvzWil9sK2HQkpXwVqs/yaQS47MsAi+e3DUIYVFy3HvJ3k6akowu52cBa/y4Tl6L2L
yhx0WoAaTI7AyqLqo0cfkWsy1K0AZQYpxCik959M63Rm4hBPf/vceFpt/G1AnGlh/YU/6jb1nTPX
ytdnm3RVbFwBXydeoQgVPtv5OOLXiv0CYCIEU+GiqHhNcjshLaXBPCy1MC0AtOLtVZSNTSQhB3ZP
G0kNcO/5W1ZSITfRZ2ne+MkvWdym8pxFhQzCGic62/p8cdG9uaQxyHJNl6pQwQXsz3TrdtqjeRUn
I1wjCE39iSa7uSYk7T6mBl7/SsDUdDr3zAXlK0yZUBe3NHiNqmjQu2DcdPBHHVzjqiQjobHQxieK
mFv2Ise1TK/sxnB/Iu7YS+QDZ4wzvvv+p5Lc3UxEZAO0ERTCb1S6qkp9Bfju7UvTPyoJnP/i+/GX
rFAva2VSmm7VRLV3WlxJ4E6sY6ZkmQrJ4aSSixAZG0eCb+q0+8Ri98hJGnZhYGBA5rpdb6JxRZI3
X1QQw6ZINxURq5EzYDffa+l0l/hBME8qCu/9qrJNsJMbM7j1IJi+cuYYxbSgpzN7OBeiXd12nJoQ
jEMpocIVnblsC66WEDH9EnXjKzmYNkO/0L87Kk6qW5/A7vhPx/t/hZb7ZodEO8pTBbUB7fZRDGxz
Koq7IuEhXF2mZKGXpwwNMCcUqW0B67DJE7j395IbEYfMaxmw3RzCr6CcC2c89oMs6SeSMWt/Lzyr
2DkgVuH38Z/2H00WapdKCEIJyhWOrnyAr0O1P6h9KGlhGGp5x93doQHht0JGyJ2pkXftI1r7hnFs
oLBIQKIuU/j161evRgG3fyGVZVOG9QbOqkiBmvrF7xxQ1W9etuSkyjgRI4mIciVChH1P4XjZJsk9
B+isfCjk8igctHIESkrYi7WpFYzBgV7lt6CeUq6mg6RC+ZkmhnS/pr89T58981pDXPYIHaDenZOF
bBeOXnIEmgl9uoV0dSm5eBnOGN8VyR+jbGdJsgfCnARKcpDVJ/OyvlccFN3JMGtqWtdqNfI8UpKU
/rCsuN5UV0vGptyvb7sr3eGjFHBDY/xT0F8IQ4SnajLRa7oS41F+zFTc7/ys5bkpl5a3ZerhswN5
2XFruJkURuYKPUyYrZjZCoO/SOFYp52Y1px0ulUz85TDFTEmi/ZZy+7jAbGPI5MJshGi2OnDqZrU
peyVMGyGBxqtkFrnNXlA6f7JCD6ojL5p2djeK99oW+FwHTsw1cnr2CoV7Xa3/zLKwQU68s0OGlVV
6LGG6i57ZBmACR2sY1/FuNCEytXVvOw8ggw6/0RaFbzX2ZCOCfrRglYjCtqsTHk4PYwPThGd0441
XO9P2YRS1ikIQvjIe4beGF/LZmAhpHxejXcjGUI5donbyVx0ePvboCw0EFG7xPp8RswzRsZSDj+S
tOacZw/mGHZmlid7qfrxSPuFD2PqBArdT73lPdS/LAhpcKIHG9Pa5VcNGW/mx85xuonPKbHIBUCR
/1+16RNQLg2SL4l6v9vFf3DlK0njQefZ+v8RWKQoeezQ6Sg/xQDNR+vFBReNjmqJjKV6vdQiGga/
8bdQEjkcglWIt1Ofe8CQvsbH7glNqhbtqJ8CzD/JOiwN5oyFQg+vfl2waJwNk2FfKlRsNbs5iLJf
a+42SNl2q7MM7KwUIMR+UceTYrZn6mDa2cV3Sm/ZTNFaEcDjzqUWI2AyY4i2JjdlAlmgfpw3DS+D
75AQnQV1EPHkv2V5xi0x/btTpExnWuDVBdju8xsko138luKXJb8u03hp1FNCIXPw9X1JBs50+y2L
l4br0Rhot1MYGbakn4IM3lMwEvJrhWC52SxNwsc/sGj4kbykT/tpP66cmLfEGMhEnuB38WZ1BjBp
wc/S+wLaRqbdrQp7S6mPnXH9oSpZ264FxvTGUAq+u0mW09vgVMrV6nJ9X9dWWuKWyCyy07r9qTCI
feHCZg6G9D7nyDo0qqwwkWMNeHrkZONhWJQzVRKEP+K+aHgmQsPT9vVzbyhBq9huCz1PSy/oNNiT
vL0cJkjF/k41M+HNLii4sqD5GqhjDCLx9szl3maG1G7gx/OVriPj4ywfgOX9rEcI6RaGxcF0DHEs
S3E4PeQDFaBg6st9uuI8EJ+Q9PeBdUGJn2V6EVUaSdiqRtYS/wGAXUKXEKuboA1jQBynpuSsJQn9
7dB4GBdSEOdY6ehxSb7P0rKsHQzE6xoWGEI8xvmfOrZlNojJem9rFwGQrZxxmPzv/YBN5H54Z7ol
K2wwBvIChdYVyv56vU7S4B0dav3WIHOnhkSVALtaNsy/W4N9U/0U3aW8eitYNxNHMhzIe+Pom29j
8vlaLciWPdhV8FaZou2FADYEELKRE6t4ntTnZjT6qRZXTuQVMFrNSoZfGy/cKKoAGw0ZrpJ4tk12
LCQx/a2hjDwdJxs+i01iVvEQC6sxreiKp8GlIFJL01jQ0Uz9XIPCLlrfgD6EqH5zXzhGR2ZeFRiZ
ocQnxHP1PGFBr+gdO4FJnmaP6hzEPT7KHhA+GW5gPhaMziuOO1OxGUwMvGBXftF43GkeBMSG5xPw
TImENFRLtyazgrcEWZt5yIK1N9swbpNSdzj98Lg1Yi0ge/F573ijAeDfHyboT9jVKeSAvRxBQGfV
cAJtTdxmR7/CTB+JZdPGaiuadsDtN+rdeI7BUk+BbDcDnEehngK6o9pORYLUbOjcvbRfBmAM21iZ
encYHdwUycl+MraWFgvUGjUe5ZhLYaPoSIAIqxt5l1ggofGWGoTCO2VpLZdSbnwmxmuuJnDsNjOh
01qTu2+dAX6bFZAtw9k3XWp2gwiF4l6rGu+IW3iPaSMcDLoKJr3DomiDQbEMnUQBFJZvpNIQPB1b
ujHExme0+kMM4zkS5t1asnnzONNTuZXJds0O8FwXD+3BAzJjIwj+Tcj/Hv+pDqPDTd5n7febnURa
gYYRGWHMP8Aevs+ZL19MHQ5NIlIdUIP6Az221Dl1jG4AZe47qzh+pgovHMMzE7iMS4g3Y61JD6v4
XGaY3LAlPmGzG0BXpm3wkaVNtir/jcOCgkJ/3e3y5Bxzr4FjW1Eb8T49qLFzbNhh9xf8pKa3u3bF
jXUsM7uJ8f4jAV+gaSGRuUo9bQ1C6qEBdxb8u+k3mwo7th8HiYBjdq8PgEyZMKRT8qYfe3EMayKI
k0iVOIEN7cvYFqltC7csYEfb5kwaDKK2u1zr5hhiaQyiI7bNFXM/0MulWsnGAaqt9Ag2eZbHovju
9KCOfxyHBDeuWv3QXNQNOhLSvvWE8GKi5IdIYjn+B7HDrx+8ATtnloHMjnZYCH58EHL3VJ8Ow2xL
VMdK1oaxuzfoW6gSatc9yS6VN42syfVaa/cdh9GEmkE+xFAwqbprmBUZBXOejKpbGyorVTxEfDzo
WE64bGeny8FduduVFRWIEMGhg4z3B/pGulrwLO5Y1uDIsXY/LGk8cvRXSUfE5QU8kbEZNEVkzUWw
k3NzznI/kMZKDybVhNaU/cYDmPF5ctll/LEpmh0SFUSVbKcV9eI8Deib0oIUgpaoNmjnZdncTjrm
W7HjE3acA+rwSReWE9tRT/uCIOVpWyf04nySsZKef5TZBE9e2+ahNHh9Z3qzeetFM/Ji0U+xJGZK
qsQkBd5pcERU0L923XdTscry7GfOj1PExOdBruxBebfRtdzTUyTKcrUhy54U+iiu7MTqGok8LQHP
ZjK3trtDC+juuqzWasRnKcFq3dzfUss/czponGszBhnATydNK7v6uJQzOvlVUM9sHpo9YtLbAICC
Pm6/Ijm6OlCgEjtr0ejrdfVObra5zAmoKi+LHF19oVkBGCjBZF1LAz5oZeBq8hIsfUkDk2xIfa+g
rP88CjRh//Uuu3+IClLJydSrp4n8w1YZ+Ogd9QlKXcggT3yn/atZoUmNe0LPJYfybuY2OthyRfFj
FcCSvEkIhq+Jqut45gRaQcBbI8Rf/BcXokUh3Ho/JifuXshfPCKHfd0I+1x38O1xCcNitZuNxQfq
XEqidLOXWPTgAgH6r6IDOl/1eG+CrDzHpO+uGGOp2t/sG/JEY1J/rgbiwINKB21IjI5aB0OpSqwU
tvYtmKoPSIuOeFYeKh2lXi1BObtuC6P0BS/dx64j0rvyeeYrwBzpfhhBHXzLoTYE8UhCV+qAKrOQ
RJopHnRmC6XxuBvZO6jBqj7/pKqB0SG63GUmjIilZ/mE7ivCNSm38Jzwp49xrMW6iy37h6/mIBVT
JaeKXU47wWQv0SHTHu/E+UWJYmQeAuEeEKEB64YUsxFOz8G/JsdovGzPyULAz1ln6iJ/xlXrpS6w
sLL17dP2BvpB0ASsXIZjndEgHnv6qC6xfp4ZQEFSw5yzU1TdSPUMkMurYkDC0b+Hr02x3YP5zDfM
O9SlrKiz5zLX8dpLbk8HEtjv42ZLaRweCVm7JbUW8Z0vmQhU2p0Ed3SNeZjJ1amx031FGFzuhY+W
1QDs+dfcrbCR4BinWbYTuG3jATWNB70rw2SdHgiMPSyfRf7pLzNA76iPk758RQPZtcEYzj0qARhm
+tnUONmz00+qPwumUk59PfKFn0N/UuC+QkGwfZHvnt+LXY171u68arTVquIPUx2SGj4Md4b9QgIG
C2GGOsrnP3XRLEQlpaS+ENxVN7zTgwSNa8XGrk1uh6PFydJOUdQmKjj5KhmdKkClWC/hJkwcLpaT
d/YOMy7gM22wHEzCTJJZw98WM6KyvTDVHp+VulqYnS7PUAZdq6wfg4l8huNVzNS5A0339yoEAgVQ
TGDCc7ki+OiiJQ9//7nWzuKmV/633MmFuqNBYqxIOO/cLM9ZL/9apApyJflN9wIlxjCkVo4iTUJs
/7g5iZTlWiViKu1oAz6N65pmySpWJJo9CVcilD8gVomaYJCSizo3aHDsPsVTrMKOE740SPvphlW5
BU3zkQZqkhVmGhYr7nyQATZU3U6FGgf0PV0fyRCmU1J+kYKIgFLjtC+ak9Uclb1LOyuWKzNAFYxn
yU0P/Bfznv8NlSmWXbPvtz+aKPlga4eNRyQ6H4QUucUimTAwAwDHsBA92b3nJStlCmnPh06cxNX1
n5njEbfVuZZBnIXTXP/63P5HjxF5LlOE4RTjjqv4HlkFU4oD1+SGnGrnMlYulBRwoh5+vJXe019X
mGo3QxrI79egGd8guzUNDQ5aHIz3AuzFI97PgKSOpNvitIYag+ru3RePdrJt2TXL91d2cD0PD8kX
ZzeLoKMAXgnrYVInacIthQctKYlV9bpDNc4c1PfzUKTUatmh73Xy2Y5e2mOK0Aco1xZODw3Y4HQS
bFsqsdOOC1q5UxzuKdOmIGKWXcL1wqED0VyA9FwneV1Fl1gJ0BDRabuXJQ636dG81smRSqVABGql
h8Edhii9Fb/z8zgEQnE8MbZPfo95bWz9O64Bhy0phBV46UrDQRI8iWjh2BPgihPUnlYBQ/DTEgxP
hJTN6C7uSUArv3aYGHjDyI6iTe9qESI464yD5pR1OBvahHTwBxtjQLUwZRLPWlQ/MC9AFTdF5Jbf
vm1gAFF4R0Cvdd9oStbXIRmRczmjX7ndCp3upuiZTTI2wb75VbI8+/wKZZwAqluveWLfJJ7NEASx
zDK7czpxgyt8T9Qq/TxyjcBujWcL0iHUjnvurLwaN6hzU6fvx9Paox0rRl0Ph8pHgByuHI++WsF8
okpv7fYbrc0uqOQdhKpUN28vgoOc8TP429lB+rMQ98MO32FFRVO7b6G/Zh8JCgBb5SUKME55BVmB
px+8TbIQuUMRVmyyerM2HwTrRR3QPERtyyn9weNRDpuwOG9B17wQh4w/Igd70gBzYXZcENhZs+ru
0pkAebUhh0cpEuufZW9ypmCyIhg96A0vFYGKwE/3X4RqHaqV089PV5lXB0WFbHKADEYQsxZ0Xle9
l29eqex6lvsLeWfy5isrz47YKrUKbew9C/8AI7wV93j/JsR4xDndRWKHNJOkaIVmCiqByb+73tE8
tgvjRw9XNVLcMCTGCUjXRPY1eG+UGeDp50h51fQ4MQ52ZpiGsygem8Hbzxbxd9kT0ORc25dHKO7f
OB78GqcVoffjnjlDssYjDGZrVaBxxEKTnHHfKgbV323IlWbzCl1Buliwz4BhvNjkqjOl6ini8IRa
drzfwtWQmcpPuGSdOj3vH2SVha2oO2GCH5zkRtO0E6P9/x18sQQYXZklpBq10ZRVWy/9CEy56/be
HQ/YT5dAyiLu5WJmL80KAMUsx82SSNRGG2nRa72WGVg26Ys4lVvwHsYolwo7GRlj95wTkjAQDxte
gcuW++gLnVGJ/VsKRQZcWEWoSaQ/DFgJn918TSqoroCxFyk3M8Kt+1HdXMn4SS/hE8R+I26oDegS
SobO2yzkt3ulugJO4OnLnezmDg6Yj43MoRET6WUE42JrIzSMXrz+TXXlEbVjo9n0w/hJ/O3ZJ5Ne
8WiZT6ZQf2oJ373rbnEPxBxy8ADKOYAttNjzWmel/w7Qm9XbbHWYM6L3+lMuMG8k3Ww/EQBVRhYl
PKBcJUSFsCWZ1eLtNHW3kE8GDeuRpqPCcpd6ZTuEl6xDgVga7pUN1U9lK/EVaIY5JlAYW43Wx5R2
cnWidlJApNlunlNCUNTyTERJ5PnlAwCMsn8Sn6+BQS+u5sg6xrC9h+R+r3GiMhk0RtplxQTdNS9T
OkXWGbWMpI1DqgSJMDnfsy3P+1VOBm+hHHgXwQDgCurt2dcU9na96vzgGP4YwCpGLBeyf9mf4oU8
K8RcRiFVWNv+AezLBvS9t1Yxf7sHYeOcQemtVnHr5nvMAfojPf2cGs3T5Dba1MQtLv33H5o5trVx
xu9dF1850LVT1O8p5HHFZhffUYJU/iQVSl7aaz6EuvXNu1TjewX4KdYOaPICkO5J0chvXgaVLh4X
XhcYZ9GwZbPgvL8jiFuHhTimSGpmS6O0NxjU5nQd6hDdOzw6bfBjMbSfQ5uxS9NRtBMVxK8/eJ6J
bse1Krt7H4Tx3a4a/pH9dMk/Qy30Uz4XWWGXElrFCeXUqhxBgD2sL7XsTfbYaZ1fXXim3KOrA3DO
ZirTDahIQvZCORutEAcJAuPlovS3o2VkgiAuEpQ3Ev5zBbNOT4c8vZ9vDlYS5a90f75hrMMcubsH
OOuZlfit2z7SOIramGaW2X/trWHRYG4a2ZrAzGsD27h0R8dASHI6RFxQLf+ZXmULa07qwPufgtdU
23PouqQvBXoa/ZVzTp1gx0ESwqXrorPQ+S0WLMq7qSz8F3CNWwwwxeOqwuRrzKPCZt0qVFWsonc2
AL3LE9dIbYZqA0RIqdJzbj+2CZQcCk5bcyLeEQbEekjUhNYwEwE846AWnqXGQu7hWjloHQ/Y3Wy6
dPGg5D7TG5PbRzatcykcDUS1EGx0w+x2cD6NEtvBkjJX6B1SfNCt2vjDC7IFby8nwe7hekyw2uHF
nIqGy6O9pu2tTGuR/1cjey42GFsVjoNo3GwEPXo3ig4w6JsMY3tvuYHFqlodcF1vxstk+kVvt0Q5
IfI3H795rJNF4ZPYzAcOgkwIMI3l5BiIN2vW9X0M7gtRZAAaGcmv13+0JexfTQ+D1yLxM25/6gue
sEQlwLSediK6zJ0yWecjDaSAf0Nb2u5sRFJC5eOkplxWHASuF80eNeDfZRZvmkRoj/IC7WM2Jm0C
UlrJp+WxW8TXXMiT8fdVWRUvEfFFZ8k/uVi47Lss6Dp8nCZfg4GN62s58Oz2wudBHlzii4tH49o/
Ng0EMieha83k4MlTDIotZfZCurCMczYlB3R2//Uwp3zYnBzOzKqRaYmwsBpnQiDs5x5Y3PtPuNv6
SPJY3XV0vJizlM31xxrQpj4w2RJEe6gbMWor2A3NILkIjd+8wSfWSbBQy+0kaJzFxdG+WXZm4GXG
mr8QXN9p7g1SewifkTbGT4MQZFW63i/q/B/clTKySW0pPnKy+XrE8qJgheJ1lq+nUBrswG5UYPAt
8XWTwXU6ypIWNcTQWQbY9YL4wYxBJz7IVUnJ2PZRCCT2ZLUeedlYyBRKfpSVocQksbGjKhNcZduX
PgMLSQxp4v+/jUdYXzjQhdkPnOFqQ+4zrxU2YNYnr3vOCzEPfgL/6hjxcHcKoV4UfpFc1+uGnv9q
fhTC6FT4qgH9n9EswFz3qRI7OShfs3G0+BIdnLyHeJVcBCzOGlav5JXo8HDzkFDLFcLS6SGNh4Fd
rJQ9eGqHktYvjaWiWUWljvYIjlABxDQs5mJ/XdWTUJAIa9rxJ2G88jcMES/p1flcoAs0UFplc0A1
CrpPb/IbYluYNY55OU8BJDZ7FFjHNjbHllHs9VVPDyxDI+NTWqWJaPnNJCmqV21sUAUCh/cmPpWC
QPTcvE5ghvJyrOoHVkj9N3xH7pjkiIbJDazQIQYo9VexsJiM4GfNagegRzR8FDl3w7+2zBwuE2Me
xRkpd+Ux+j5L8hGbpbJnj5Xw4/56AP27AwUCzI996mAM7fNVoldC9fLtqsZemJ8S0oNhZB32cJKT
FMB/gF6zeB4qzxP/tJbPyzhT+sMhTZa6fyaYy30nB2t/GRKXc97CcW8b+7x62EHhplBXVQdnqN/L
anzHonaNkABiioedOvzLqk+pkT8DpZJL0oLzywNWYi1+7R3wjCUf+Uu2FE6KOfwi8W30ZpW39XR7
v6JKhGoa6Mf++dYc+OkSnr8I45xsYfizJocyinlur+UUTDh/vh/sfpNCIZcH5/7SRYtbxi22ddjf
ZZ312LuhtoXsZ8TYuO3V1f9uoBhlOLZYi3J/DfMQ/TRrrJ3JS7lHZ5mD6IjOU2KtLw8yuSuaLdH/
M+BYZkxwf7idhRps+HAXcjIhZQ00T1+1SJLGETOp61/jWyG4iWlEKfPoRh7WhGlVWXfRyjNtz4io
mYMYhZSwHmk1ljJUPa0VZQ3vpHDGvi4icWUVg/i2qoD3hhtTfC5/wRCNvso5nYBsWmVKwfKB/2Co
5fqzBOHtH9AmwJT5xxnE2wsYgYxc4DiiWne6vOnW92Q9XE+5NPfCCtvCMwZtrj43YxrU6dy1++Ns
jUYimLY7LDZK1ykIahcSLMGCB8MrOhYsTOKiXH7BUOEIxDZwRXf83F5z1fWntccNEzGaeKXcUKpl
xq+3nDjs9SStSxtkZ/FSBRdIeWsiawVcQa/svf3UuQzSxhlXq1+jaf60BmF5PqOGPHm/AXaSk/0S
wcenMaxtaTFYfeYsjW2WYWziiyQRhm8aB4mpDe6EXMt5lcHMKgPoV0ujqJtTQPTGG8ttsC2ygXti
iVzPBeh2BBqeB1ME/QKb6rkcoFaiXC+KK7JI513/jSXkKgVFddYy7pLkSH6QOq2jLoIPz4AJ1xFS
n4QmJyOWOwt3dlVjitiQCe84U4GIFCBKVegQk9f937pv5GviJdyuJ4iTFeyCYVVHSCeKSaN5oURP
LQPMOGjwSn7tLl57nmeSP9c8e8GYe3n4EaZVoX2jviiWTSA6/OARH9+9NJAHS9a4APF9xxL6/BED
QYEOKBw/XzeEV9rmy++bwdLGbMHGVx7LMX5y5ilE3C726je9nor9UXAaBmMzccDSrCwXIwMqmxKr
OqTxdno77Kpv0ZmWJaGQ1bHRvQ/8KdvmptnPRgQtVUj8pE4/ktekDNY+HA4xi7BqoIEa7iqs9dp+
hl4M5XzzGEx4NsRA69eqDML5+sGMb5thb5ueg5tlA9IP2CCQD9SLTvtSkieSUIM7Qv0mV2JjTfkk
PWUfdVbe9/HV2mBWTeJIV/A+H+jH7w+4hE4qlzVwsbSNSTXHgDjV0L2UHQiIWezn6si2kG3mZrN3
UW0w8djpoJskQ541Quf4PvSWln8uNbIM801UV3/4vaWKy/lVRebS+UADlRtRtOLlTQWRHq6a3iP5
EChmsdjKuJaoLdIG+eN2fQEAiLW40MumgRKA7Bp7/vHf+GQAH1IDHdx/TjeuiYwuzduy602afPwi
tqSniIY01KH3J9bOwf22b5Qw2AGCleZq0mVzRdfUO7kXxy4JcvbBL2YyQtKC7PBa5Vm4ysIBSQF0
omxdXt6l4sSmlxF/aiY6qyln7e1DyzpdhldY1vsmAixtFrfC7szQkIX/QFMi1vSRKKxN+jeMJDcw
4AKF+7zX6RkmWjWhunciWhzuYiXIkN1x++jORrP+mzW2ZF2rJbR0pvDJgSo74WNdTNF5vkD2KCAi
I/GuXhYO5GtU2do0bIHR2aYq2b5lJ54dY53R5bQ28uTgbCyxldPcCNRnxhm7qXkHtah8BlKiaXeB
AP1Ky5aEq7mHrpiWa2qxEjwMK0O192j1Tvd5jUJye0wBV2h0L03PDoZRFxSTesCFDBkvDmyHe6eA
zmnpneyXO3tSgpBKQtZproxl7ZSON3Wb93Nd31Y+ZfKKLp4+IX8vjSVtkG+0GSpGISHqv6Dpp014
8b9sR1wltkcmgdlOtVG7WgEEwOQToSvM9IZGNFkRlzRTuIffYRefDBR9vb+AHptDtGwnPJTvgyJP
nlXubfu4ctYDPy7yaj8n1D6t7AN6OnkceZ9O0NwxkH4aNnFqL11TWt6Zekh4u5cEckxbTpX23m1I
oi18o+yyfz36/kFUlAC5BKW/oztaiTnCGdj0ih3XzGWcccU8B/jVfih9Fxh9syOhuCDdJ6/L4FcA
0TYgIwALOEAHMzxcqegIcVCBGKUDhz0XtkKJlYhu+ztAwhCp/v1aVpjkQoH9zy9bCUWv8TwetB6K
I27VM2bpj1aKkpgrR3cb9FfvevccC8jPzQzsWDY9tgiq5yS+AAgIEjGa1F3Z7g4TA4o/r7ItQB9Q
qlA9VijX7DfKvwcINWKjGZc0GmYTvfjkoVHih+YUsBfu0lbFcO04x543NZAWRyuq0mz5bs6nJcgX
qbOgCTebsnBXNBjCnu8riKX64nCUW2WGyQbAndrRhh7dsVsHdNRLykXAWkO7SkWOnTxIfvgvpcfm
wTwjn0KnjRr4lHC5BI77Rpv/506OknYbxdIgJ9tuZPasocZ+dbFwpYezsTxiO8b8vAOk3z56TzrH
MyENZAcdpKApCQ65qw+nIBvihbmkrIUF21mHWP2/QODp6U8hP+qC6LZRSO3eQodjGKvmlvnh20v7
lJSx9gcd+65CdM/G4d6ODaVKscxcSJQA6g9i2x6xApCKXtPHQUARECMpAUUHari/F5v2Jwrb2p+H
5ksYiCRkM06TeViJg4hs0n74th2A4b1p7gWKOgIcQRewpcaCv2cXJ4a18mqtfDAKsFKnZNbJyQqx
3ZoMdwxqUc/JNSC6rCKs3ZEzNhqkqwwUo0EBO+V9m29C7dSdM1Pu0XlXM73x5xa/PeBYFEETdJah
2qz0vY8Ke7cCepA19S4P5OtlRVrGernUxabdfJqQDMlsciKBuXixlY+SFlktbmofTb6X2KJYzFdn
VGrDR2t9NSiantDfVqNjb589arlmy62eWatk4yNhhbE5qjEJJmiprOz765hHDdC3287UsKGdMkv7
vTmAh4WyHyDNvQlcvUVFmJd6toLXd6MwxUpt8VNBgU27oBpqsgAcvUlNEERqPylkZZgtTD7UGsX1
og1DGZUUFX22DevH6bZO7tURIHw3yYJS7KL931+wykz+vfHJzuMtSYU578irS5ISGNvvgnXELO/r
EX+7w+FLX0YuTjXniJ5iFfER1iyv+2uD3XxEphla8uRxLxcZ1krLF1d1qxjmDWylW3RzxEOExPIQ
V/0kuAehGPxKu+9sSwWJBfkD4Prvb7UVtO2aDkum6QsQiFJy8X1/6R8ebKLAvfSCBGFSt2vde1tM
gDLAxqIFWkLxSXowEE7r2Zn+SrTAMy9vv2ICCzBFf9QqznDO1vcQix2EyIerzIKRH+nTeisjzNLj
3Bu/3EcaSAl8jIsjPiNLx644tOyiuU3pl8tXzXP2Ox784mwNPWruuE8BKrcoqzXHVJ1KN5aZHCbk
ZVd6y7vmBsPFtgPIndG8iMB9e4Y8F0QkIgNcDwbuhRPdPs6nGdt1ihaCZSQcuRqkFI4XDJTICOVO
iE0aBXVLtyJ9M7dDfesGmZwI9yHn2X5/a5BMGKO7QUEIBPcK7dYK/ZhfuF6xbgyVRNEK/rsRpawk
YY3TQC9fpA8U+GI2JSBwes37XCuw1sDA0ImVWgRbwCYNXGZaUkQR0n7+gMCM2RWzWjIpcIG3rn11
pNXhUpVtcS2oq480oh2h+i/MT6RAwv24RUEQVAZqwx+JdwvouBgMZ2rsHMrD/hO+3aR30Ne56LzA
fUmP9fCwKXwMSfpRoZS8lcM1uMEg1KVsMHQBnLsretq7AbWIZ9JWQx1IYHBMBRz1SsyOMLsu+Ilk
TWR0KzFIkVMXkOp1JnDlenSSW8T3YTvwoE0UfFiLBfwQovV3cuVSrI4dpp5kxzhbn7ANqZQnIjCU
M9J4w7XCONjkgVly/wGLbdZa1oarhw02L+OihtHcwNXYkqGpQ4pdV4XdmxwBxY1P8c2yMKDA6ON+
MWJ7BzhD84UDBdg5qhN/U3f+Upl/BW/0CqjI7bHFfwXftriJDjFYFnouqdO3/A9cHxfUn3/v/M0r
f1KvHFxlykb5MyLUK7IHe0uWevw5sLgKlffYRdVzzDyXIASP8GLit1AAIr5ddel0TyNyRbxq4u62
L1TrMi1L2MPQ0iEc3DIMbcJgPLu2qYN8hMMZyEGq3C1YTXgnMq1r9nk9/m2I6sc72fXasR6oPxO1
zalZhwmvi6/aW0FhFkQVm7E52TrLSMM7pUAPUvkudlIrM1v/TevcFI4jqxej9795JMplp14DxMHY
IUyQt9Y7UV+L3OKzzRHWtLBe9yix2+7/UnE76tAlsTDJREPR5oWCN8MMiaVEcPsjpgtdSNHN6pSH
SmWHiZQglnJ/gwKXJr/RlLctj+NwobkCOleZGhPgUdGPk56fMgc4NPTQBtMamzX5MPZzFHb9W/3n
FDi/Pn+z0UmhthS/QJQflPn/vZxvAS6tS9w8sgq5xkWCRSmjcVfzowfaFUjiflF1lekBejkTQLf9
CdHCG+F6fVcjzbs7O8dP971lJUKGbGtMoM3FUXI37mthoAxUQlR0RRACLuVxDiEFQxcdGYhrZCRP
lK5otDJbT/s/MmTxb9O3Z4N4mkCmQOjxJW9Cz8gQCNgQvXpsncwYMWo5TZaQYowwBBPJQPsTU1Y+
ajqrwuM4qFYhAg2isSf1jihr6IRJwE2J3U2EedkHaY/fzek2LM2rX0An3Nd1+ovkUXvfB/mdfyDh
dzUwSjIs22utxB2gyG6B9h7QNki8+exE2zOxidHqc1zDkEuHJx/aGvROoHnppMON6Azj5IcfBUWI
a7wdnJhg0ltQm5CLNEwvPiKaqpRTCZA0UPRU6aWr8aQEwftKbah82t7UmtsUWIzjCwcIyMGQuJYw
GZo2pMCEDjEyb5nQYm0yhzuDVzjMaUEFdFYZEFc+OUIrrdhTfbjypMJkAdJDKwXTfTrQFTxARwN9
CRjn2auXXQo8SixATf23VxMd9M7pm1W6ugMab0oKnxO1UwGlB95WF+n5kFh5bJxEQC+hFD1zR2Ct
iQub2Q5s/1Qqv/0ylwwZPLR9IfOGAHwAurrOPraeeyMmP1qrCQAVx/mJRALGR9thG77F7+I9jZqu
fuSGMd8xPlgxh3k8nX7HXfyyenGksSue3n3XgQaPJuulrXxG4YLEsZAk+X0jCUhH8+x32UbpXJod
/L54YGa7x8IwMJdzrqTvHRtS261D2O53Z+b7ZYcWjpTZ25Yib64BTDtqCIp0aAcsS6SvTp3bVFLJ
eDBO02xC2w+81Nq+fq/lYOkR7ISba7Bmv1YuRg7yDCsSq4Kih7P6GKuYfjDPbMC1VPPSrKEVFeRa
iCT1vtpZWoSl89YYSBa2Ux8FmsMJxrQYCfZ1cyv2/8x34SmOIkZbCR61lGP6GewUdXwon8iERIk6
T5OV6tJ50ui8xRUW6auuGarVjci2KoVbPik1faN1wa370lSOsq64sNVx2v7xUGZNgju/zm3XCnMN
kFUT1k+DGqiWyYbfYR9z76swfUv77hG2o027GEgk4o6olj1TMt04Sa9d4ujKUXa3tctRamDwzBng
K1rnc+W+pguPGGrZpkyyCB4kbYKiqyAN1kCL5DskTOeDbYTBasJ1gIDLFoGCy04zQwKXb5OHKhFR
Zn7lkCo0JVrTgbTuGcEDx7zLd4X/oLPjD4VYWX5XpQWqKYajON8Cu0Yi/bC4sRu5sbfy/6luDxHY
BKBvpPjogT/Oo7YBosnFNWR1ZKEwMlWqXa4W2vMeac0tOv+JvmyJHYKvhJb0vuJj2hcpf8T4+4aH
LZo1+yi4acxMELoevQRSJO5IlWrTUSndd49XX3mlJWdtcEAB5frjSIjWmQVS8uPcWTy2MKfqHdRX
fOfD3b6siQOj25KKhinZklGR7dsFww3hea/XnnTLA6CNclQmwtJsLggI33ks0l0V4cQ9w2LGzqhS
e+DXWlLUpgyidtLbS7rj4TJJG9KUX0qIzOSFDKYHlc4AU0bRwoNCPf1RWPiQtb/YWjnFuzukTfuF
QHGsrvxzlGanLu9C63DKjq83pOynIomktoXTW6lOk64NQToocHaH8CDi1OkRoMeYlPZFKMd/QO7O
P8cpvr54+bQU4Q+5UBgL/4JSElKByXKFdxszTUawvIBKM1gvjUjHSDcdQXvRo2Py0BcvVG5gFckq
x0uk7FsfthDkl0nQkNye0IOfnXustuk6FMOY5onUwEi1YzqNVUmc8aCDLibHhodYr1770+o1xwj2
bB1xN+ltB2GEYQxe0HLFWsNWkb5hdRV0MlmVT3oCwDPtzPvNkLoRn/Gw+MGpNWxrT0QwX4WLC9AA
uS/S46NeR8V04XuogLh7KSrpsZm7RFzSwoOkgbmzu45Nkt000dMzqLUB4ATkDxspLj62tIEqy6Ue
sE5PjzN/lhgSySMIrlxNa7LKNMIgx3jqYNZ/2qLeyaiMsRCcoqaCwYktwCZoG8V0qmfC3DM7+GeE
hc+tk3VGrZ3VygeLNFtDEZ2uv3lRUSgTu76vZBQ5imiWgcJl+ZBlsglqEyeGWfMd+OR8fUY9zgS1
MLjgzmSpmYHceqI35ae2NNpBXzF0qYzS0+rEPoz12tvz3sinbvozf/3EenABMREXKCzz3EPfaMsd
Qvw1TgIbXQp0COE22w0YrWNFYrE6ELl4Jj/+i6HlRdeW/vqy4qcdotdbl+UqlpnYdSBAZjrcOw1k
QSTs1/gcUTLyqcGQqyXFKhZM4MPzgqO1SFWxEXThphy5KgQKNekn5ayDrJh9VVo4qjnJGPjFhz21
JOTFU60buXekT88fSdg+jJbpFoRj1EYV6sn712xjPhuoPL46ZOf4XYa/4SI1ooUy7XNEgumq663q
bIpwCfTy2+/bah9vVTtK280FETZQBVOP/FsyhpvUZmqAIoXzcl9RsmXeR6yGTCXA2GSI+wtnf1cL
qokGHLAAddRNiRzRci0R4TNUijKgA36tvhnKjqiJvJpwOp5Q7ZvCbHmqtqIwSxypYYP3dbZGBxJ3
D+BVloub7jC0wEntAbCjLHgJzDO+i/caRJN9znNVu94KtO8fG/G1QB0zcA+AIL1adzna45qd3VK8
bRsUKI75YujXsnhMFUq/fJI5essKVYXOjH0ZMt2kPpdI+Z6EJnscHAc2QPGU1J1gX908CC5Gk3c1
nxhK3jMhL4lQWp9Orqxtuf9OUe/GcPxqZgzCxCXto69kFJ4j9xO3sw/hT7FZE7b4l7y9rHnTpY3m
NDUsRNsRFJnq5Dr0TGurRnyE/S8u8uXByNHXnP7TH3jnxfaFOgg9mPzA7v72AXKq2oWa/kkzezab
CYvv/tmSS630SDaF0VBZYN5sQU/0FadjwGFccIdZjdD074JxEx1DPoHcYPEmj5LWbmisjpofyle5
oEVHmKX//m2QRMdJrkZqqyQybYqNcRzKHKEyxxIWXn8hBXOHtoEmYv/XhBKyp/S+I9Vg6GhRVC3O
fK2vThtMe9pe9/v7lQLi3F+M9Slh2zXqY6lBeLz5wFFdGCx90EN9706R0NCXXahOYmtcpPNXVv6C
UB9h3+Ric+O8JccQwoX7GEScXGI6FYDZtxPz34GAg7gYzC7sQdG+pe1dinKEdl3FwtOJ/bh5aF5h
qlxfgG8MzYxkoXBTFMw4OPRjcvd6adxsNuuziHaAaHqf+T54PVx6/8E9OFc/M31ZHAJuRMunQLWv
j2J/B6y/kazgBHxNXU8JODGilMjK6E9wS+ZpThk4ZtZuQySQWv6o5ACuF8jQmfO58KCtPHSpTxHq
3V/ZZziaB1SwIMxK6jGIhtC+04c11GTNEyAKlH/CwoCvxg4VPZBw+YQzJwszyTm17FrX2yoS8rak
H1JT4mOTLMp20CDLZRvuNZxj72xeNkTgJIOYYmipTQCR1/orAFBQrfnSK5HbL+R8LNpDWX0HtaNN
kPdw1w74XWfM5JebTupQda5iCCytHqW1IdnJav96PjreM7P2NrbjlxotXiIn6+WUFnMRhZTxNZzB
hwSuezDRm8hJx60SFO3jmR2DoZaQy1+aNIjAV8RmH6BB0Rx5ZQkNmXV9y1bH8lPa1W7usfnDC5Sk
od9xXoAt3MuMBkzCeZOIuLL1heHNM76cxDVYf5yDGJbT7uoJwMjYjWiD5G3fcxv1ab9FKhvM1jdd
xoJ/gAa7HiYzswUJpLKTgPKnfYr968wYXLhV/rHNEDjKymQdYNQD2XtQ0GwIx5yBmXBbL9kNK8eN
uNhyPeASVT2nncDI2RXPyfiVvbTif8SKHdst5cpuUdH+znlja8QreBVJDTxZn/pKykDGgbgXXi4n
jWrZIWgLtwnUF3aUWtn2fLtBlZ/UppY/TRp1KjIQrVDiKCV22NeDzIZDQyXmWa06z093MKF2DFYO
r3YUvKrMcb7J2QjdQEHbjxVrDIfyONylT5QqEHJoEQjbUSzYIcjywIsG33WW4yFAPW5a9+Ivd/k3
EU1qMUTEhFMR/hoFm8z6Dl5K2lP3RI7M0QJGnHJKYU6KVfugqnkNc1UMotNOQs3Q6QQias1efVWp
IxW9WiMPc3XTVO7ARySWyoTijjunYe/ezDinntynp3KCEtzgiOa6NYIMIgR+z2fP2+a+mVjQBQe0
aEre126Orwhr0UmQFGnkzNVJlbsnly8RBkiURLQ9/stI1j35bTh2YwqxbZTFOjaaRbapVLCN0/+2
tmD9PIZ8ojL9SoVLW1ulPDCC5MniibF6d2WUd71Z4r5y89K16xWdtWo6MVKtAt29cznLlVlVe6CX
ZTV2ippkTXmhr1zUU4s5Op1VErXGxN1vs+9KxG1qBBj3uSd/EC6uxIwu2BJqNZohGehwpfMLp2jX
Tjo1IeFXfGDzVtACrwzt13J8XK2jWnBiu6b2crzEh9VPiZ0J7POePRKHHKaa4SbEIGzqUIH5iM9e
84Kxrm/BNooxIjusJE2BR5oRsQ314dHYrijWzBRahsK+DVgxEZW38hBg6YN81J2BOH4sLK5B7MZG
QKPOJbrsAWcC5waUHOP0aFQt1NYexQKITCfYzOlrT21GuRgaRJvhrgseJb8Mjg4P9/WRPz2sIn4G
wZFml8QX/0Rl2SDWMZwNZD7h/kQYC86bTI55lwyhB9AEEo4WddVnCzLvZhMCoIgJor5jbO1eh5yF
hVg0dVvhg2jARfA36+ivROtDBCe3aglF8zQuhEv4MLdSHqs9sIL2g3UVvZd3QxwXxzb7Us72PT28
7lMl3wX9I+mI6Up9Umn+ySmwlD8zQWlJPvct1qRR1zRXJLup/SsLNJRe38/4zr0p4w8ncQrN9jJM
GHXilOmNBmmJa92BO2p/B36bi0y1mhpyi0hhig4Cy4epRgGhrXC53v0ArOX928mjnFpCjZaiDLzU
lZZaW83WkHS6hIEVmDfILg9w96kx5Z5xD/pLJ+HKU+2+pI88cncpWXX7uZ+qbXbVKJHqFJksoRjW
sR6r9lnMzp1hJVBQNsm7vrXxmpgicnRC3jdniHRjAG8KckwJi2h+5qlyKf80W6QqeAQhFBzdX7H/
ORhVjyEH3PJNoDVoV3kQrwLvmd8rUXlCl/9c5gmyfPCv7Y9sAslBDVVJRL3258GygtOa0YqH/dPc
AzXl9MsRRUj4J+8nZL+SlXH4CQsI7oFOeAZmWRLv5BntEQU4AgBj2h2KD/elcl6yF0AXFP4JuqbD
BWLVpTovZNqRFaGaT7s1GH/tkAi8Ls9nR8JNUAVawl2S7VgGzqVfq3oP4U4Xe7d0zt36L1ROJoit
gF7r4o2B5hp3uZ09Lv0YCxlh+AURQc/59KDoTI4+Uo0q63b+hsqBfYOXhPDIHt7qMQq0eUINCzMs
5hw2c2dwPgP1C4Bs1nGzbQRknpLwLKngQ+wMwk7n6piQuveK07/51/Uu2jKtmDn292cPDSBXl5bI
5v7Vllzx5UxZT3n/A56ssO6lpCiYr1IQ9+86iZNdRWy38W/wqur0CYR0pD0CwRdnl/0h93g0EXi2
DiRNXcFr4heuP6lNMRNG2Q2TEEYtd3O0EC5ZeoqYdEkLktmp+I8oErs+NWW2RtXdJw6/QQTKEiL/
XQUKT2Gm8gomcqzZ6NPS/d4//JNwVOpFdSCNygB55qGyqfZ/B6MP5wRVE8mb6cxYsdaomteUdTyT
hpNiSkJ8HCSwaMXrPX3P8qSfbd5hOy2OeP6T/GTQ9C1zQlJtkz6zUK3StK+VQ5C/FucdPSqk+9pz
TtbaJOq1ZWqG0RAWE4xN/0XGOIEvUfgExiVHUoswMhQ3KMfrM13KI/uwL/y80cBLZUkGagcoBq1k
Lnns7Wqvz6bRmIJt1W3LRMs/90SP7Zihnoe5VR8D72DAyl8loEee/+pidkneXP7XnfnPwiTscfWu
RZMgDUmnHWb9PTfHb+2hau7CE37WyKixmccf5WF9m3h/1T9tPQ5BzbMW1Fn3mvhKB0sB7vnlpEZP
12auJPjvR1nYi9SJrnyKOAQ4gUlFnUPhUGxMUcbimDI+oH9PwUCfFskpTMnD8DQ6eAjoTK2BW7GB
BTuAa7t4kRvJvK3G/GJHiBZOJylFdiDKGzUMZZTkRHDIgBseqS5hzoWOg27t65ySfChBtdsqMZJU
mL7WxBLALQQNj6iE9MccpI5vaPLL3yDnMmoawlLYZ7QXYOyKFkiWgznQUy5GE5g6xDmG0n3OPlDv
xfTXG0QMl/i9ilcR1uId58U7nUYrr3RSBJ90Py+fLSJOkyzn5prmrvgZkcgrBtR5qSBvNiUmxCVN
pD80M76b9x+YZp0p382VFvrzr1nvefTf9v2Ts1djRCItGV0ohP3T1AugqNfd/piRGGYh6Sc55AYb
zrFfD5UQOqRBI+mYziNxoZ5QGaBMjoAB2GLr8QEq1qW09EpXQQbxkc0ZcZouKOu9pxReO53VhBJT
rRhzKmElOydE60NGA0mCdwXgvxN+loVsU12RBMfxbXJwHkoXePYM08Dt3GwGKg363BfueBWAPZoa
SITKWdNQYAyA091JYMNWf75T/pLjJG8tub0KYr4BHchdHwEafftUcF+glPd5pmbRPPe5oKMXHRN7
Dn3shHJ20IfOkhQ7YEfTGTXFb0m3JJGA+FbOzY9VUtiVpkU2E8isMvELhirNXqp9YUi+29RkBoju
25Mn3t7OxiNGoTFlGlNQM98A9J3KkFEBirbq9UHnEnCPRzKkLj65N0Fdzrq6SUsnWm+itpw2Tv0P
lpCjWfTdbmGxiF1VtTaB+ujJAOfPN6cNEY4OeDVf3y0M9pdN8iRXuFtOUxI2nF40DNWpPoQoCFkn
QHjueP/1OTsrk65GpBCqTjF3I10DHoBhQkKvbYao8fBTbsYgbY8aisnYj/w7SGhAoM/JSgDHrSO9
9cvDRMpdJra0VHxVOPqTtJrILv0Vkm46Mp7q1qarEMzxvAC0iICoDXJUW4n95WoiSmI+ZMDky2hn
EWGiedPogNGfEv+mRNr6bn2o51ih+z8FtF45oBoSRvitPYmz42sorSqVIDtQBJYf1fVbHDN8aeGz
4odsSY9qAkrKAaIqstkAGgYjmbZVSYkqwQi6FTUJz96R+hzyv5oywwF8IxVxtBqW8iABKJ5iFXIT
HZEywn3sHLsa4b+9uI98un1nlvgCSHDSr0L6SvWjgVwljAxsIlZXGL31Deeakf8yTRZBwGcG9IJR
SH8M5WXaSa5FYzwrJGyzqWjXaiU+GJNBaarEkpv7m1MSve0ETB7zAaF4MfDqg9LuldC3uyDHSneh
HNaa027nNoenEXx6CPQFXDv0T983Chk93jjgf4CX1ycbVpOijL/80xgSmVTr+VFUsGMMRNcH7RA5
KlYYjFY4KLMmdoS6Pw1brc2dqpvnmtKOgIh1cchLjUmucjD5iVCO6ey+nHIQmePaXOfStdYF5hPA
NfQL0LnIyPQ7QFaWVUTpPQxXLTJ95H9u0zfVU4Np70da1TFkBNsZUe/sR7HACMTpmrF0FuEzzSKe
PrIcSddA9bCIazEbw8H1EZ7FcZuZk+Vr0eQTY9jW7pdd403G0Jj9fdMim1TijfhdXwT02oFK7a7o
XVlk+ufUvkHWL74/6VyIftZ6ceaz15O6IKm4jS5l/pOqbRrM7SxlqFqHC/FdqrNfdcLPm3f7tI5s
avlZBz8QaUIbMBW3bDJj2Lu5K6y6rJx7e3KAPKIoOUhujaRn/Q1OvmwYJ4k0verC8PpqxbqJPQPb
vr2p/Kre1vPQwhiFFs2W6y8UxvGjG1eMuMfa3H+826NpYVQihsw0ky6URqDxCMX+UgeYw+FdXJlY
YFB0UpRazOGvCQkdBBofjtXmWNoC9Q+W8IOlRuKnoyUChDNNyWZ0hqcb7EH42opQFhHKQ9cv/rnA
dvjzAyY89kNB9NK5y1iDkrgAFdBYqoaeVLEjJ4N163Lfd7nrQo7/o9aQzeH6qnb9w7kUsOcDpgVX
6yc9cNF858FO3dB4X9ostTY84b2n5SqV/WG/T5y7IK/hq3I3vo6JTtxCuOiT5kQXMRli7ZLulEAR
6dTRMPE4rnIDZUvM3sL/rycFTpxZaL8PJVateOK8O2MEfyvzugZNcmaKSsjjTY5BabUfatD/u8VB
Fw5Wyl2sjuEKewt912RZLnbIKj9byQaqo1AFadotDQt95dzEXH7zsI3OQuQ5BczLbQzqMXOx83ZG
+e1opccjjbwG1EtcVBFxqgMr3ECJpztK7ZNXYUyoUs4AtL7UoO9ObIHDWztsduTRflIw97ACOCWn
rsatevfgOTsdNThVBtAO6n4ducrLP7+Yf6nxTPxRY7Evb1jvdQHbdZzbmySbfCmmZ36qmcTWPR4U
pJwQVgJZvG+vrz8APV9hKtABC7DsuJ4SK4XqMF7+ljtOFjoN+4rkQqVhiUApnJHhw3gndgfbM1gR
AdygNDfBn3gKH+odqDYbc8nNrpF4G2W5+d9rb0JTkd1sz8IXu+btpEgO5/k4cwpEpQfaXJ3jwjbY
het2gmC3p818UQZT9eVOZ9uOHJf0sTZ75UOT4Ppr4OTrdVByvDzGdx7+J52B1L6/LzVoRuDr3jOi
JAmdeFusjzldfkypEPXuLc5HwvMB+vrUKKMIZSDvy9RJ7xLMWgtXwLY1f4FCX8wh1s7tFh3aj5dc
vi5TI09NOx0750SHPRCNnRy/yhPXxp96/CufHbLO+eG6OZJBp9XPUNUNkKDefXFI32bx50/jA+ks
K+tKC1uTE4PHDSOYytU6GVcQ1g2TZS3FJbKp6Dy1FkgSPSzS14CFiweg53MCJ5fRTk5KGoZrq7uk
FYjhVh0h3cHRXSEyr/9BGyOepPw9kTsf46kurT7qHWDhY2nAOL4ecmM69BQmAK4YmlOVO8TLDMX1
vyI0hct14jtG2baauJ3IDN/4f8JBM0H+V8jpl/nAOj6DbfPRRzpK6gmAOgjXku7SC7bb1mpSP2Yi
9wGznDy5wdQpT+lCFN9Byoywpp5ikWaFhrqfuGPVHWdZeA4FjpboNEZCTExALVFA3vX9LZU/o53X
TiFiGxXyk9vkLrStKzBVW0h51E31GRPmECri6R51vK2nfxNiioWsdpVdeSsb4NHcUb55SBYXtPfx
6BxKFCuHIPYLJz74Ht1Ry/5q6EtB4HIhl8JK82gYRoHArNsM4GQ95lR3m3mqMcLPiiDEkEZzS32i
EURilU5z4cMm2SKFP//vhbDtM+NLnKE9qW4wusCSMli3fiIAxbXWFNy6RySwTYI33V3+aJzHUfjG
q3HfdPpEoZOK8EzcE655fJmLTIdfJOkZ9NJvhRaCK7MKlLVEKdyNnbWf0tX5aXwKlt8chpZ5CUKk
s53bWfM/S8nXg37OPfLoBMrjMonj5pZF6A71zXTqhso2zJcFhRYmMa60h8k2Sc0HT/uYE+Z1wHPU
HbPVE4Q2gXspP92SjiA8ozBViF9Iy1uvAJeomIEEvcaWTeDL9TZDvAj7k/PAMZkMxsb4MBJiI/8A
XGrFcZL4HG6GPTZzmbu/c9zPrKrEsYLeM24pIpyGTXKcO9XGEWZT3Pu9gK05c6fl2ZfwkMbEeMql
+kRJGQgLEU2sTjjeMCG5MmC2eaON1S1R09rUw8AwK8QSQnbxREK9YEQryHhl/QMe9YaTJtYmr2ox
G61WnKVsQFoHmzygH5KEGEkNFBvzJl9BDWGBl1jrOmRROfHNA6VSJ9EKc7vMRO0MXOssAMqGomvw
5XpNL8lGuE8BPtZNE/Gm4fCUpnAHjTCEoORlgk5oB9ppPCfayEMSqSVrE3/5cpeqJGdylaatgd5p
jm1Xkqr0fwnwMN59My+aZjRvw4PuRrEumgBm32ssfS+xu4AWaINeidqR9fTywHsHq7f4yiVJZqbx
OomnHEbIcmG07KnfYrYb/uYh15WrYbMstSZ6ze/SOAEmWs0SU/cebhPPgKxfh/1tXdsHGtbnuiUF
p5WgFKj6wljrL0DJt2kbC1TCcyHSDUNIU11jqVHO33olbGkLVC65tRpL1knAwHfdtP1M1eN/VLw4
W3Lxn2WRel5EN0ubopYdDx6RkE3XKMeDZt4K9RvkgyKLCAori4s2vQHuuSdxxWzlkBy3r/RJ1PUl
jpL79ob8iDRJFCsZZsMmBNywMvKEC0iYimIhB+kCa7yc9U0Db9WW/trYcu9VFWUZ5ePZuhbpSiBe
WOPgS39sn8RzkBLF7gNJDVKeu5kwF0CKZ6fshxm/vLFFfg7i/Fx8Pnk2LVr4F5Ixn6P7BEWBc5kI
MfMecF9IMg0mqT67g6130wnSv9C50ihBvuQeAaxgqzhnNMxzBzIp5GFFhMj5hgWWDdFcyc+QGyBB
Esl1/E/aEw0NI5HR3TiuOkkckGnrJNzWUT4tqzFu9UCLAd4u1ZxmThcVEsi8W7POXmVSkxj1AhZg
zBkVNX9k02CEta1nlkDCJ57i9Qoy2Tg2mZNIww70v3Vc+RoTH2vzRbC9vDCnz2Qoq9XtlVQ2pySm
xUNHl1aozvuvptjDb7JXNqkw0UtgbauLspGX/mBz3MsJY/grmaOooXYdObz2NCYjOfxeuVbWtm7P
whYl3K7F6nHRO8N9P7vzaf9g/G5+d/lc9+voLYDftId6mJn9HZLio99HIjZ9l5TkFSIbyQXpcPc1
Lhq5AfQFL6/Syk4fwBM81wAA5rO9mDG9MnZtA3ie7sqp/Nx2oFTOXkpiXM/Em2jwH1JAXfmWH8kr
R9gyr1yzBCZfdFLkFFkDRlIPcnddvvWOKcoPBiT3hjXR04hBQpwdG08cPc1GAz55ZNn/8dfV6Fdt
lTJbfu7jf+ulKuO2G0bItHb5Iu90OijPfTncwQMa728FN+lH8k5Mq2vo19MJkGfjNnubcshuiPSG
5ROlRgY1jyAQdQzodpHDfcxWi8L1ZNYinvgliUSpu0D3oeZzova0OaD8BVZo8cgLKIIc6M+f3R1V
ORa2jPo56uENnYaLzBxciqJLvQhiXykYszZbuWSxsS9hemTfmt4A7mD935ewVADhq634th40spWC
BIU0D71VWjoGaTVW1x1PBGhiXUmG+u1KxDv+yYo6PcS4cLZAJpob096MxKntjREldja7Rqd+/GQE
1tg/Op8edxGFonJPEXXQdGJkiovTQpqy4HIDxaXZRv/XL6cOCDewKcRsr6+Lwrg0uor6FjBtQc7w
1rUlFWRWTvftFWCRs8R5YAahKk/26XIMW50BKKlyWxC1fZAFrlzwGw918llhBp9JzrKWQ0tvBTw9
EbBv6PMvCO61wcTfcs0SaVIWpyPBq0ZtnZHiEzPLfL2Rhkjgr11g4L5yGYomcPRzlIfS111vUZWh
v08U/BUw0qh8UxX90qWQHYSnbeHaS6jTP7gNp0oL78id2n7XUGf91efjQ6pmbXdlvhHiejNZlDa2
CvT0rFDdQbqx7GApOJXhzcF/b1mycDWaLh2vUZCyUt2+Evt+jfhS1IGLoAq3S457jO3jRtuI1s7Z
wqWulRvY4gOnIR7SINxu0KelCnsqehQ0M7KNDBtXFELKjDbHgQHQaPk78TjAeQ3gIWg24jSBfVp+
4Tyqx9RwyTLg/xuX6SrDK8sxayKwdTSHaUGf3aFCRJI6fdNN0gBGzms7snmcKIG1toSnVhiTFRsI
2Hm1MrhFr6nu+xvhIztNRxwebOlVkho5KY65W2ZvPmucWlM6gDY0dfC+h5K4qDJ+3PkZpDy/cxlb
m8NOgPXv26jYzq4Y0ukbhvm/2y8kc6w5RyIIrWNHAwqGn/55KPMEDLMC+rTxjGeEaJOpNbyx92rS
AMBWzg4q6f/b1Hb1RjsKVoc9qKoOC64iPowlGFs/YSKvNw1J3NAjaw6BQlpd8Baw1cXAVTULxdO2
9gnnTmzJjf7efRzYwUqnvXNb7AixvF3fmSTEQMU3JGXjlFINcz19Ecd0o/6zeK4iE4ftzNGjAbZQ
AqFHTrA06lA2501wt6tnbilDefEpIYd6ndj/eeTdsVjv6lvaCHzIZbNPTMk8PcB5AJ9nx9Sbqo4b
UGDqjp3QxBzZ+uXzzuYRhMYzsnPBozWGTTkFGLtN53KZAgxi32wCQk045kGiXIQolUdkTD/Pi1rQ
EUPCk1X24/SqYL0nq3NjMtTdck/Xavtu3FGwWzC8GN0B+K008hyAy1buKcZP1VduDZ20QCLjvmun
L3C+diYcz1NpSLxzBKTz6kLEd1jVNJwrKlSsNrWz+2fA/iS92F4Y2RR5Q/mYS8+w5JlRyXAL/2/F
uwbmoZ6IOvEIgrOd4hw3hboK6jdAWsEkWwjZIVOa3vclmiNIQp548iwo/H3B49uEFx2tgC3AyaDO
r6wQW1956Er3f45oYLVyF1u5rW0a+jUF8E9UICaDdLYNEv2meC4XnWdnn+ECLcXJ31LK6sjX/dWF
UfQngRTuQfFQUdXrOVYpv28bZCb2IjCdCjBLYKjcIX/c9AH1NHW7NT7ooGEjBzM1RifuIqgHSVM8
2I5PsHWpFqDujp+xKnAQggF3N93T11r1osnMxdRl76S5qtqPZhdtuwvYF/JL4lo2fvYIpQzIqk2p
5QObUkU00fKbRV2NhISh3zmgRvIYDip4z0izZXleUq6TcCLy621/n6t5809osZ3gUpc62rBdbMNw
ksb1cHjMVtnBAA0auImCsUT0GqnDu/OjTTFzmu6GhDD6t0lpgbNw1XvzR+ZTGhk442dmZNnHNbg7
3PpfvGFvzLE5ZrI1tqPrc/V36QmX4wL7JXeTp2lTB2M0HtIG9Rz95nlXN/FnJph89oFJ94XTglxd
XuuTNHRjJAjwKyzqBgUX8w1+A7PKLJEjN50Pt20GN3sLCaxR5EG7jX+et1XornerPzk5t/bB+z/O
Hx2Vh0gZZ/tuztpAPDXxMiy7uTWgtJ+4YPeiF4jmiydfK8R4lHBqpmOXWrKGikIB0+aSh9FEyFNT
PjVD1U1hVcrQJ9it+MuT5O0dsCDNKBtCRpwm37fZ4CRSpu27BXmiR0OdIUFsK/kB/wt9ITdCyUnv
XZMm4Dz+Bn70oMsWfT/cnMBIIN4HnXJJWe2jv3fAspoCiJdDi8YWGKMk2XZPdVoRfg23Fp5w3f0d
M0PXa7VP5n+UBHLpHSYe0Fa56KMvfx/18LgUvqxyJBcY5zk8cE3GgexxYQTPqWmub7nFZcZostBT
h2Iicd8Lym0ZJH8UzcLFC7RcZrCPgKBOeI3OHw0SeT7Opu8KbbEl1TBBAF4wSpic+cCkJ7E48/lD
YMDl+9/t9YjTUM+8LrSQ6gTKRJkLtD568xpr2xWC7kU2FzgcD+V496ZUJawCXIf2FtTTm5qe1ezc
7SIe3nAmXYA2aVNnw9GXNgDV3hikl+2p07jDPYz4xNWKXADYdLSWcUmreVo4H2j1DrRJOokcHzZr
QGDydVEAcfnO0K/2Y4pZvmosTaWMU2+TRCcQEWozwcM81uPcpC0O/+Z7FP1zCTq+GB2T9ysuGCNd
/HQEZ01IGJgOn8bkmHl1hIy6iHmk+A8BOqoBDnSG5yrZc18kgiVEipXSTWFStw8SMKPmo2btnYbl
XbeVZAiOebKpDztErADSGZwRu51OCdYWvjYGDcmV/QQswuvXJRYL39CihNqIu9O/AJ8olJWML3Fx
UwRipviWrS4brEAhByFqhUekrk/3o97UwIyCO5yvwUhoHgLX+lMgo5xhb/oU99t8vnWuizTmut7E
nAOzg80TVNWkMNEOf2hRMJYpj+vidbNhYADfeLqKRB8IeC903MzrtqvYffPKk8fKnCP0D994qF83
JaevFrqN3VRVhBOY+LolndrNZGXPQ2y6Tp4kzTbWASq72PF9MUgEcr6Ldll+Ypdvhw6BZ04g6ZY0
mHkVkUVf6szkfvRbVf5SHsoT9uzC8Vos9w+SUsDuMTfO75D+K2lp9dTpmcxRz9ncXqQ4GKtWPqo6
ElB1znSUZUJ35aUPz/6NDQI4Ujgh8STSIu7JhwIUhb2b4tR/jciv0nDk0eKDNZK7kLLDitygsK7l
1QpUvLYt+f/mFF2yYwUgJp+ZgnVYHJajlfhcgKl80B1PPHN3JO0kZmb67+v4RqJ9BNBTfuO/VpIv
NpybjKg/oRDK6NLZrP0PwhUJYwda4mZStPLJLOI49K3jhG/WPdgi/GX36MWmq2/8aRgZ8KJWsj5E
vwEHP9pfGgoMdxuySMqNKOwnjCD5F7SAA8DzAbbFchCH3uxgfhX11FRg54oCI5z7AIOURTtXGkOp
pDJk0B0hsyWT55i2M31L4s3UbyfkDZAftCUpt04ZN1JZDUs6SGUyVouSKX1g8n93M18bmVDG1+Aw
BP6fskjevh6P2mxtzH6aVlkErbuaiUIBLtGMvHgHZPXf00VKzELb18VDmfeQOp8MzMJA7BDA1eUR
bRlk/dLwIz04s9JQ2xHYJSf4IwT498V5lPvO0iTTUbKBp2IVfa60u1Cx+LtUyc3d/TpaubCx5dun
2G0l81Z6+0qJX6Gcvgba9ilD4ctF7AsmADRgUmR/Ok9XQd3094cqywSWBRxZ/j2NtWEXRKvt7npV
yb021noamV5Eoq/OQtzdFXHi/ROuWHeg0/+RQ8Ctyf435eaGGWddrczlSkqSk1zJiKhaFk5qhgyH
i79T8kEgXZgXpnKktSxClkptuQc0DlN/l+DWEK1gL9Jc+HFieelskz7h8sNLoWCjDjzZNMTeR+6q
V/01uYJQ5R9EtFiGVBLIaE/hZabO0yQ2MeISbh6gc3yrttYhEyHlAqe0zu3FnyYSEOBGilFDr7Qb
upLkssNXJAwgZP0ZzBp5RRuzMdU9SJu2vZtTO7EBMQUr/vgjRmd75ldWousjZzNOVwmwG1HVMRqt
gaAU6ZmOOF/cjhWo64XcIb/TCMoZgRDD57KxpLZrncJRJqp6ag9DWdbbVBS8+2xLxNpWQQr5AzS0
ZlacmKpb5xIDCczVnfzvLl9Zd6ZWWUmy4HEZoUI7I1iDe5yBdmb6Lygvb4Hz7FfiGVWOI28mUe0G
xtrt6JQTLDYyPSJnNmkLtbo+NZ5iBT4FVKEQGmWYxgnLp6Q+Mr+jQWBNygZ7MUNCa0/Y+4xAdB/E
oGgoAJ6nO70gy1jqZ8AUuE2jF3V89QwDvLNaUJHG0ioQRvli2is48bI93sPljab8fPb3knZMzwv2
7Lk1qNauptDJIXGQ/ElfymvFuzAFMjNa5kRrM7B13xEH2l8wffcrWc8BPpbsqq0QThvqAlfnIM7P
kNeFkuHowW3nbwSH4lwmPVflnSKOw/rN0/EzF60+s2cvkVpblyAfXvaLQvTJKiVRiGOyx5RYCo/2
gr0PUdddL/5apTjl41NJhrZ4JEKB8Eum7wAQQInY+yub3nhIbAetLfEEthvXBYhmMCFFljL7LwXE
fhm1LjVIpMNAdrTU+qHCFkseWBgrFgIYvZnM/m4833sE/V+T9vugYQYk3JkQ8lTCpYeJ50P5s9J7
CAvxXVc82t7lAakMvmmSrPG9roAiacAg29lAGhF+MDjXNVmMSjnNMN387QX8Lmw5mTgmgsPJJ34G
vyngTMMWWdb38epvJjUHBJ3Vg4W2ZalrBg9oDO+JplU59BE6w39XUu/jq3PsCl+AWB+FezXU3Tgf
IaL9dqqbgKdz+grNtOrzSwHzyCkuX4RBo5Vh4SGYcpN1jbUqr/saqpBzCfMH/rWMb/5g2RU2KWZ3
k03lMtHrxaCazOtP8YuPL7l8rxDOgyL8aPpjYvHQOiNFeh9N9vGjBZcdsHK6wYU2+rLs9AkOelh1
WRSkWjbNxcbowZmPraTE0dx2BpAlBau2P1vZBkot+EWoti5gLn6ivvpziqLcJwcbHkLq7tCmWO3I
td5Zigu5Pj+8xcHrFZNHO9qj+ObJzI0fNF+vWZgzKAbGZW3OS+zCHykVzxCOwoAt1deOLvasNSwT
0Yt7ejMuXad83HfbwHWnjFR13s78KAKCsewpOGrGnXeg04HI8DYoKsbsehIWGRHlzcKXkAmprxMj
EXsK9DFKyzcg6mggYZg5Tehfl9xAcWUoFlu5szSWbTGlv8ywMFXP4cfQEWB/PuyO8aYFFbsyHiTs
+yhL4iTsMvQVYwps13T3MiheK+71y4SuLFNJP4c5r8CFAcigGTzm51JzO0rmRMcZluTFA9lbUM53
eRQ2rY3EGE2YrIV+IhLbAiePmqYzFRInMb/mUUght1EMK7RgWn/3czFgGj3dvfspy9tPZJr1eULD
AC8zSBhKP2Ifa3eVPGX7euPaKuhPq5G8JFtXUOSveCERYE7xQOUauWmcDvLWqDUG3BVtFzfdwpu7
tDqzQmNo/aiIeYAetSOMBC8LWJy6OuCeV06DBPMEOD6clk5CZfcaqJ3ahHL+IuvEXb//P8n/UkXJ
2ex5dzVo4/Btbr5z7r9aYT23Ed69Xq+wqyjGmQDUy2zSqDgeT4+KAgK9kcwxETtsghc1P3kSdo8G
ECO5lN5GFG4UwgGjrh3JbY8cwr6ds3q2UaAQ3mRvNzQ6jEVxwuG7smpMMvO8n0IsYq445eIeMX8v
HGb5yY+GPNgwuge54Zm9WUgmX1e7v8awWUK/uY/a8vcf2uXKLdvCsCAof0bEez0kPD6+aTZvtnS6
8qcGWBu+dVUqRxzHLMDlyuuNZdBYyHtLMOnJ6pqkqZo4l3Gnb7f/WmicCdIwVkjOsryO0HAUaYhh
IMgOkeiHlUh7v11NprYF5r4K1LOma5+yWa/z2XM6SDMI2Qf0DPTrcZfosRBy5BpCGN356kAO/Dfz
3Tdbpj/K3yZe3b2igQdB1jRQ8gwPXYr0mRhr1e7pxhk1gsdcxYSZ1ZGwUZ5tAGMMGi8nscrAz4if
Rpo5ZT/AkzQxNCRhVL9PnUaY1wa6tLbcJhf2a7sveehh0WP0VsWZfL9w4BvWmyo58nKjvZ8J8x/I
pRfXeKxGB4lMD9v/EyT+aNwItlzLL70+E+TTQT8J/88dUhinGCVRw1KnDjPj/i5NWa1TnoX4qqxL
qVuvJjl1VCfZqiv5rj4CTGHYbVne3U5yFMQYAF6ujGpyt3svPnF3dvUKTaIA1qL7VVrGi5mxwjnI
KJE11BSQZkS9vvpNOUip2sD/pWmUP+Fzfws6ocVqlH/6gi6tnxvP9YwXtRNoBIOK+EsdA6l/m8l/
3xP64OikgGb3VKrWXrZbj1Lv4uw+jiW98/RwcP3v4Lxj0fsmcDgMhAi/CpKSyds54+k1W3MNXh2W
SF7dLqoTsCUpkCFkDXTtX6+9ofKCODClcw7ebXyVxJl48DlvK8wjNt9H0DbgwRJIgWhoDo/Ke2dL
GKD19jc1Z9/tUlSKI8wnnIrwiwrKresn6xMFP3NAHDo9LSaz0rKxmrWnQvbTyPZk58Jml9kkEUDb
gRSiFXUmcFSX0L7Y32TWNyHDlOsJK1OacTx1FksnuQQDduEdNJxzRObA8Qfh4gsLT3aHd0wfe8Jk
2zzza6mbNGSt7SuZXjdQQ3nWNaojGB+xY4MJrtrQdZRgbK2A8tMLAZlITszflOvGCyX/y7y2Ck/t
9L3U9Zwy3Z5oaTHoYmHCNUoHL88A1VPY0o/XPc/+NGqn+2VnT14lppFEhyWjZFKk6pqWmTpeTSl+
7JTNbz5gzhLVw3hLmaYx7FswjfU8my9WSCIlEOKWBvG8hgRCoaibkLte4FAatFxfSTvothOxTRAM
MLZ41r8HEwUhKB77vLAY8s2dy/1B3+A+rqLjiS/Zh6JM5RHXf9XPFilra32etFhGzwd0pa5CP7DM
yCBbR46hEYFwd2FtiTQy/d+r4W3ggtuRAzkb/4FX0Oeb9U8zn4QzhJ4mNY6ahx98CClLMuVW3Ydx
4F7sa5nFQdXTuKrxPAgkK9j9Fvp/Pl+zzp+Lc+0CfMbxpfBkXNTI8QkRpn5w/yEUuptnJ4lHNWIp
wgI35EdksLKkA5Lv+AX60OzUfbr4vIbKgYyX25Ddnu2vSppDbUnLgVwY9t+w4Q/L3OzF0YFcO0Ws
4sAy1CmvhpwGJL6iswvbX/lKEDAtjCK9ZorQ3Si4cNn+B/iPF3ntpYtg5OtFCLE8iW8UyT2SVtdg
Pe6RikX4+pA2G5bMqgqboBt6DofXHInvdwULXXoDEDPZvBZNHik/EwMDBO8KLlLPj/HkkyNk4620
y3jO2IGj1luiisINo7STSWJuSRSCUh0jgcf///5B5+/kOPVOCZxjMevIrdrEe7hxTAaX0k/cer4K
FGU44mU9GvUslSr2RBhAN5G5T5Fyoee0xl1/QMDxXXkHKbHdcwmNxyMwU94CGYdYbrzN1qiP2ccw
L5z/tWPcVKTYk9dR3mcMRyomp1b+2zJHbpDiHCDVYQFTwcOCcdfx6pJsVrbzuuQea7bXL9YlYWqj
6UKT5H/VZjBxOwxQGeoIBaa+zR/pIF55P49v/bRqC4xl7lCzCVtXh5QkNT3MTo7lYyGWWwaoLaHh
EuJCwPoFyDtiOBO3lov1Mc+tZa24YVAo+XY4MHxGRn3dI7BpZgM5BkU2Z7a1ILeJ0Z8FoIpHFhDw
Z5d2T6QHMNgaJpVSphHqX6poienpuwmDwKkneHeTWb18KOa299SBTm8BvBr5BZ9AUzgxSLVZzMae
1A49XwbONWxd0RaRaugmmDHvpCgLMVBB9GZQwvLrrZfsVcubfoeMwOMq0g2bTfF0pg5nVwPkXQzs
P/RvlD8jFWmVhDTEsqq/7sRv+xazrp13HVpDvxxNEcQZ2NT6HC7oZHFwuCbkmWnFe1suDcXPtryE
fV+9pi1l326JSASqR9SjIEJu/72Ve6osMd28cB2DE8EpTwNp7ooWgHe0yOSpheqHedW0ITdu9FiX
urkm7wxu0aZKyEn9fG+yqmmF/QISEOOdkxU5uNVv9ihjB2eyhcaAusJTTdBr2SKE+xRDm/nQMGbr
AD5n9hz8Hzi5sISrx6DQR6qCYXEkT/TLXNZdDMYk3HnlzwLY3PxQVy5RuSBNdoSntwP1jlPMgu2A
7OgfynWP5XBVdjO9D5rGnHobwKbzHUcFMz4ocJoXWA9AGMVPOTKIdzvzWXGaJZ8zvDSV5yJLzFuJ
H6RAhJzffiS+d9pjxcI7nh/4QAlDbh9o5ms81dJt3GW6apVTelehJM8YhognQVct0LNehZNgh/Ib
4YG2pXMm32GmYi3de4xW9+F0nJQhAYT7gFUIxHXcoOUm3Hq0unz5n+mliuDDeXBPE8PQfKSVV81a
2pcsSNQbgMp/PUY4sa51CDy38t1pwDpztSpTueq8JliuSsvxxMeJfcjEebgO9WgSI368CsKuhYE9
f34AccURMPxFa7wntUzz2x9fNS//3PaVqD75650Ko2rzfcQF7g12qwMAW3L0VcWc0hu1efYFdXmx
QTF9go987qFWFdtDZsvptD9mth6x6JiAx6Grw5b3QZ3zpD9TAuEWI0afTXoovnVftB7Ry0oX1ctu
Wd3/I2FVvL/tkt3UAlRByDm90jwFHhEdRXcI7tUxge/yVHw0Kvvm8MvfKCTcLs99GCH7oZAcy8JW
QJLhiUu68ctnXVDvaKAJBJMDEa39dVcYWHkY/OvYdy9+3CBOnExOR41nY68ptwohuNFDxCZzQVZA
TgAsSniGtfyo4eEIqkMX9J6EOrea34xM61WnCXeuGcO2IXKIqLpdbtwDAzG+rEoRuUcRz+K/sFF9
blLJB5lvWffQKuyPE5h/+28qlyz5b3nAd3wZSbOORhXsYXH/dMaC4OgGCzYZyJJcU1AqSKf0SjgU
oAjym6EaphkE/h0uzRK69f1nd6Az8i5ZSvOL7urYYWOmXCUWGMLHCjtvMGDlF/0tQJXyzkuOuUWB
+qOtIc/XA+GoqaX21IResJrdvGhBLQbRIE3794drQPwmR3NFEKCa62IhG0oHL+Vn+1sHtU8igdro
lP6NXS+G4nx3GBT1IHgFPwwurX2Z1wcLzD1VpHOL3wPa9Y2kJ2e35CO+J62yLnLs86O8ViTbGsA8
tlRisqeubJpT3V/jWDqLtXdJ/P3E51yq02VtH5ZEx94UlCDfY5IskNBGbgDKTSAqjdZlcjDU4fpj
/uNYkNLMj3pLNHSqTLvFeux6NP1cvOvqRI/6UR03VyP4TEWGQ4yP261ONENDG0BvQiOTWUVR454c
YMHlPSVe6sVtYnqx/aC4+SQjFAjVEC2QrvD4bqPBlFm0gnI4ZXqdlU6HPQtgeloIlBGp1/kwepfa
ZsThxgFZANgOeCAQwcjEzrukZntLe8JiZ99sxCt2/an3ghP9uJJ/s9ddUR1JF8phYeu1vaybtcUw
hpvfPHoRp/ItVKTqU3gLs+vOObXXATu7f1cjkQ2MsaxQMbkUIyH6a1guUoT4MbLTUUrptsyW68OA
1lXxCz3JMhiUAIabxWgsRACxmcdAb/kd1iREZ0Pon9mL/L8ie7/TP/EyeFMC32k6THAw4LjqQuNI
8mHBENBeqFRb02GwUWbjhfdWSV3GV2nDZDWHDc+ZDiitt4t0lm4crd+GuU9sLTpR/D2z6LFBEkXf
+9cYdO0leCUHdVB9Mv3AWc8S+1a0rUseiPTJLBmmxTsnvtFJodhi7olrsSnR8uw2vJ6pLRy3QAFO
uVsX8a7c5OnLweRzAU+Ca+SB0yoNd1Jw9QHBe9RSJeIHoCHukA0FzNQHrSK5VAIe6tq4sahyPLUM
phslz2A4su/XV7YJTWZAaFAsjnjLKtf5bYbBqB43RDgN4+EvIMLI/h086DlRx/KsO4rrDjKRmZtl
xdw7ioW/r7dfMsIpbqYD4fq5zy6cpLUgWdep404x8G2BvO/9POHlgwxjHIBs6EZuwOF4MMJbQS/l
/g2DJ0icZPXhaZ+0jlB8t8J0bjl4JeIU8923Vq0Z3JpzL8HHCbNjQiqKKP0oyyyXI95kEVV+2DDe
ICpz2aqLVg2cnOgQmeW3ukSu0H+/Ga2oZD/Nc39MvIUiHXb8uSdzFwu+NPPLfCP2iqjZKx75zm1Z
P3f2LmPEoU1Gnkwmubx6BkQOuAdvTBOhnAviz67vF2lB2rqNUb6kzTghMbTAHX3NET+K6czY/7NZ
cuV+9wgAD0vyPnjvf878n4tWzlyMcO6knr4f9ZjNdVJsDvRl9R+ZnkZvth+APlyvMT60CRrlpM6z
7eCoJMLUPpMzaKEO0NepD2iO/ZpvggsnyAhbEoeevSdY0vAhxzlHHlH6CciUla7BBCZrLP02CCY1
c+miebbOBWgatr7kYa/J4us2w8xQjn9qVIhQ1JVMgIon+XKHdjrvtDwe+6zjPwdoy+FiEQx94jt9
QBoHoQpki9AEHZ4YPCe3+sSnDnrBt75FCfmiNEEHW2fP85nnSRqF/3QfGTeNzYuqP8mIzT19IDfV
c/UZzlKkYB5RnHm6Zyrq+o5+qyDtRNhAGL3mh25e6qS91Iyi6PvAEVJyEKOafXIeMI++oGvJv99J
YTCwA3ktYyJHyDeyg1HZ6Fje9T26w2qFtP5q2+TP9y26oazxYpCw4JCygGtqdSReghjmTS+G2bWX
teyQqiLmcSStbjIj99WLsLmvhTdf4fy+GyhaTcbq14A0dSILU7vLle0aX+T05tNI/FU9rgZjx+eT
dEguSAeWgHLZfnLQWfTtSMZo9SEcBaHH5osuT0m4gz7PPTvaaXwWhxkts9rYXkoc79XqRQCNEzVi
JiBLhSCyvSvXmJPmrFIOO9I7J++EICJPIAngYrmpv/L9ax0l+EMM/iGxWC0ZZEhN2quMfCyjGdzz
ZJbIRHwOjQQf06jJ2MqJJOT9hpBgrhU9a5WeJzJuAUeFGpHwuRYFpdw4XMPUR+YfEnvf/J9BW2D8
5F6yarq3ge4TDntfdN/HcyOGQw9/Si5WNz02SWfFCrQ2u0qP6+q7iwbBrU6d60TWlnVFqrKYgq48
AYtNnXXaph3xNoIs7jq6ek4H7ojIa4HeqNMzAm6VvYsstB1sU0JgjV7kfvDJjlf85c5Xq6aIJJUi
TfzzfDhlYg+tLGyMEsYTOOFLzWJEYYJCZ57xwR40fYUYx9RE/UWZY/Sv0ApZsz4dlKw7AhputxO6
nm5maWAcQzjaLzP2EU5N1Nk+viV0emZwhvY4DKH6g0xtYols33roi78V97NK4QOodhBFVpq5trFe
O0kwNpv2wU+iZ5OZoBP4B3bPINNwyXQkNBPvau5wSmNTjN1KDjcw9GOZiogdMdWMUzLXPeF1wKYw
m1Nz02nxWPGFNfixakvLoV6IlmXHIGv2dS4xM1wYWminVk9N+RfZDkjr32FTXpLuxcv5PBiNVA5f
KHCcxQxAI/czKBJJPRIynwqrDHcaKF3jlr2HZYz+9VqqfrBrt5oVTtzsMXJjimcfu5rgRM9xvY+b
l36N1TsdVCHoqEsD4QJW4k/P6M8QSaKsBMnwxZtcqvymVFmRo1AaZWhrOitx/c87GepHynUVOZIr
qG94l+2Id97nzF9fGAQeG2Lzdmc5VH/tNb1HcoChFm/ScKJerSp/ROzZazuqbIidoEM3Txe6C+cm
8zW1W0FvRgsbI3AJM34uMoTvtxRbnFVXeSYmvm2yJ5cNPfvFFlyoNkh3Djyhw8rN6Yb61p/G8DiW
DI0B36hiBoSXC399KQ3sLr3UJ9YTTrIk12qlbKfdMjG7akHjFVs3L3o227idWAYvcp+qeGdIKC7t
hrgGtEFYaZl40LyLUx51gh84peTECgheW6t5Pf1DqecAuwgcRxqV90kjmQS9d+TAmclQTBfzM9ab
iB4r+HTz1s33s++JdPqsNOtJiDSPlEYmHyUD18fnex+jEKiiyg3QnI/XPaDSdclXQzUit7iYVdz4
gG3ANhfloeOV5TkHYd1vpZwsUjCKzzLUEguhPbN0UEQremuyeyAnpW5eSJfu7PTbp5tkWIaMTNdO
nyrneOdt8UFQcfyKaFdPdnuRSH+D6zzYylwYLvPgcjvno22jH46E9R2UsCwVvCX4BSDsEpV1mwLA
vmP2TJTRd4vXUlOGX9xx60eK1gA0glcleyNU8qibv//vrki+Glu7pAQKJ/SBhhonJaXfOBZu5SdH
PVGRjn/+6EOPBjbhTYqzJDDAgDaI8VNu1z44HsVFEC4itfUj5XRLmnWundFmaiNlRzSso6avHdAE
MaGJWwv5fn6xEup3ZD133NghzbKbcUa4gL99y3eNj0670Y9RsG11Poi2/UkgjEINDEXSD6fN7PYB
4Ks8qMbXhoU2THnBECGXBI7EECAYthNmRd3wcc6RqIKTOHxkYsM31k4ou8aS7Sw+tIlr384JQCsI
37kXNkY4d6c1etTsAUXZ7pccOUs+q0NqDEcc3L8zl9Iei4vo+4wBWVcoA3FzqjAGLKKk3QBWOan9
Qe052mCWqlLx1AJ9LvySKqdDwOL0KaoZ2RFaKg6dMkRM6ceQS12lFxIJ1gIAKm2/toPbkjznPKCE
9S9piKZ84U+rz5Omd9EYf1CdYqRoqZU48IbpnDqQABsBQgFf4lHwHfjQOqFkurz4YcKUCZFv6lPt
EbghnT47O7ISlEiw4zSviHhsiio6TOBLbmA4OVXsW12oibf9JMLm3fnlPb/O8nnkWtDbHLYoQthZ
HmtMfv3AgPmykxqmmaVc2E03B1jufqDVGXXC802har8GUcyx+XG5+t0AWDBnBZLkX2rdNpEuUOxE
J1mEivPoKOzOADd+DiOLvDOaP1wfsL0XZJbfTi/h2pTOKVcumx1rgTEgjQdlyKkWTXJw8TCP/IcQ
Z08AWpqfgYRyMNt4tv87ol8FIrjcugTZfgsHlfgZtTzdr+dCjPLQ0XCjc60/SCWXyfSshpQN9Amq
2R2vh8OYth03wxpRh/qWHKJxfbE6dCX9uPpsSa3VhI4WD/4HhUCO63iS+pCI7svwvGKb+FyzhAhk
nU9JWSVCB0TYz5Qt/0RdKue0aRukG8b04dqZ3a3Zv2mPgbPRNOKU2XGs/jAerANrhWKDq7aRpNUd
XGUX02oPYefUVmF7DQOscCli6sfg1lEZWLYIEV7S1WX9s+Kr3I1nTuNTLCOPl1yP4MMWIlhraBW5
xi6J9BGpbIxoA8zXplgpKGa50ap7FD1etriLb3X777NUqNrbuIjtseIrwke0f6KIr+FBkBpJ91pZ
AIQSZiNrL6bFEYHQeVRlgKUxNyNBeXuXmSqOZtp62VRflg/idZihkEas1z5tNZYx9nIfTLZe9MRN
cDvuFshZOw6q83cJHxfOhA7gJgasDctp7bt8+BsxSamc2Rc82LZ66sDGfeDRzzYNHUAb3L6D83sB
x19GTqGghF4Ov6E7NnKEoDLlgzJ11UOycB2UGrTcfeOxaaoNlqM061EGIL7hzcA6Mt1Sc+D8t05A
96razbzqsO3YKKFOgcfv4kEVTe2TKgN/o0M2WqH0wd1kg1gW3T+PvpTR3QGGYzc2l45TDY2a1ZV2
/QJifTpanVUqjjYDZsfn/+6LHib8UKqYE6FNypIEgv1ri8ndF2w3XW8Ndg+OuSotRaW8FBd8RrsU
MJJA+a/a1JHhQ2OXhFF6hHvyUmWx3uuQxVhffXWEo3Lo0zD7lPjVpkcdfZVitcG5/Gee3W+mBrOH
ToW8SyMTlBeCyLdx3tBARd3aa4SoCn7Oc3knVIrkkUI0sG62wU2slhaHMOnEO+1I1iO0Xybs5FwH
PVN06ueEqYAtVcKafXyerw+jIvhHZnLtoOwm4G8HWCj1jCkm1JStV81ME0LfEO0z2jgXX/dycUjQ
/QWRvAU4I3kPKsy/RGO4F29FuxMfk2w2836oU1NK4Hi2AZ6Wx/PwfS3AVCX4p5zyverrbo93XbHk
oO7ikJn9VZyOFEB0Kkr9mxsvTH1hk6cxqKq/BOeh9Dzs2/4xtr+G4M0Q1QlnvXf3rojsLdgdfnlh
se0/Zhuxr9wAKtgTgH3ois2nIOgFW3fufzGe/Hlt5LOGIEk0bib3KbiXTz1r5sACZY1HzJOd3qZV
WIRF5oFFYG7qzQyvTJW6tpTgiz6g0Suhp72xaSbK2UDXW4LI69ITXSV2uHwNfnJXENOIASgLxTJ3
HCnXLCSV+tbS3JZXbTAB5GORbh2owroHJfrXDPE+aHIQlMM14IAjfK1SvJ6RuLM++VVf4TawdW7X
LK+LhxRu7W+73AFAd9pkB0OG1RkH2aRnTuIDCP3jM/idNI/2xKz/UHEK03XR81IDUfvcTXbnJ/Cb
XKYB0Ril3woU+afthMZo8s+mGqvKH/aWUXvn4w8bP7fe7sX9uX4fE4Yo8jJAAzC6PCtNc0uulD8x
9q0iee7oFVV7jmldhWxugJri6dwmYNZPlwYV2pggWNQwnrTvwTrtnRduWU1WnAvLNoQEuCfwuDx6
Ru+79Z99/gZO9y0stGWdaKgWoOWVrU3Ug2uElT6P47LpJE4PaZe0CF5yRuXEDezBxkJaXtmF4g1T
LZxypwW92cqeo7cRq0fMCKGaw0hC24IgT+8QyWuugHx/TPO6KAV0LzsLHLKm9fSXlqFl2lVKesGc
FLTKJ2uJ75xrSq5QuILL2FdqNlVxdS7KIHcIO+SV9t+74zJFkY1K76zGFatDQF7ipOVs2J27fchg
oxMsVFs9c1Ij7YwtLasXr7Zb5ix6frbOuCldas3ZS/Gel9tuMBBoJLQGKhll87mCnqcMopZW6ohM
7yCG2gbI689ziIuFbBPjcH4Dpdzttk6pA2Dutx2gZgmIrcPYLFmQA8O7KtCPsloaNbGCykUuO+JV
SNpItOC+sPpeXLaB3r1Vp4fHzgkwnsI1N3/QSo2h3NrMyYUF/qb6sutX+iI+gv93hRztrDabimcS
PWZsgUaXMKCP9zzANSo/Wl8Nvje31oKmB6AgN9SS6zXTasw5fr0jk4YmHhipyyPnf+FUA0AVPPJZ
UYjTy9an7YD92Lfjs9tiHvEykFsf4BCGnfMN/3d8A8galkDPalAEBk7LvOzpAjA5k0QBvKLa1Etj
elA5O0ibXETKsS/o2+CRHFMpx/RxvOniSEo46Z6G3o7aQTj61Rh+GDCRz+rsDSMTNu8Vtw1GHsep
q89J7LmQYKTmW4Xc2wx89xGTDpzCY90robs6kMtAtws33crAGRwAfq5nloeYP8QnXyEWMYRwLzPh
5HoMeTuTGEaJx9E+ryoreRmVOmil8MitJwOyyGeISJs57hwQmkck1L70VfdMDxFB5fYvgJqSu31W
nUR41dNwKYK3RUU902bQqTcDjPpJOOJQ3Ay1zAuNhAtCNxaWN8SgjqQa7OK4OCrklt0J9yB14BCL
l4GtjMSFyC2eBWgW+9NrvbPmhK08BI8KmUHiA6GdWtZaRK2btKL8/8se1Ej2522bzdZJ95CRSPX9
UKDxYdAkw0ELSbUHPPZJP4MSrf5oUaiEUPi3KVK3JginD7e+jRJwtm/o0hUJFNNWtiCy1TxciTpm
76NKSoyUalqeovBiHndaH3KDRYImtcynzA40MpOx7L+z2VO6aElMs24FYKwsoThV/YN/ovwX4nSf
IpJl7ovmytUWYy62FDypTC7zLcpzwKxVmB4ugAirurD+WTMnQnJQSFISavDm45trzbW/tmIXStxL
F85TpQXFyUUlsSVk+F+RouNl9uN2/qjixMK+1VGhyCXLOovXkNDFk+S3j7NOAK/8ThFBpgY6qX3w
XCEqKh0IpaD9Tcc5+SpGuL7i7NDxcs2yrLuS0+ERUyiXwhiubn1i4+Ud3cPCYK6DpNqdBzBQ+V9i
o/qp9ibAtWnuSSppuNTqhcVYXzYk0RKgf0xHMks+/HmztoTy3ZQM/IbaFy4a8gy1HJuCpaefXyFo
P+Jr7zkP6zM+wXOmL9OkGSaMSQuTHDVp4awaEX2/oMYmrA/XbFHEVTrT1ZM4KkYEnQVMS18ZcMkd
kTtC3aFbm9V0z0kxocRR395MwQJ+Dm0LIood1QloAId4IpFfoj6tnJLYKxhpLWJHviCJ6qCusNpU
xrFGzkF6bsGPpNQrmj5ckwuZAMqZCnP6eFBP5WJcD/uM85t3w2TWhErrgy0bV5LKaNRLzgbEU3tC
HSHFm9m1k85ImYV9JL1dxbA77OAhIY9J9mu1zSzluaiYLwhTE6XVOYSB5tOI2sF46Vs2uDnrt6tO
hDLmGqT7l3A8v+Zgpdcekgjo4N2myYZKbthkfb97c7EM0P6dA98LJIWq3gCT60YWvr8cQB3EFAWB
MDvhLpCB09CPqxI7av9rTQntqVDv04RYxJCmYIcjoM1hku//x8V6poZRB9746xcMNYIWD9sgG3Mq
hXJItAnXnNOC+aqnQwEkDVmW9Pw6PK4eL/bF0JMjry525aYXvB8STkmiwv8lufgdkS4ULeh93oST
uKP8z2RAF8a1Zf2fn+xP+Xkwqe0QE8c+n2oPZGsHxE6Wio64S8mSscuFvIAFVx4sORXAbwAvugFp
m233idG2uhRGeHKkxABcqHd2anJ90m5UYTwJR6XFH0xbq9KgibfW7lH3Ag7avRbqW/I23NYGIiA3
gskm3WZbUWaWivnwY9PMcwMkQKSyNW8G81uRcoGBDfm5O7QcUuTx4YN7ICxWfBOibYgwDZXPTYmd
7O9tC19I0xTHltdUp2JLZisvqsX8gRkBj8WqVPwQmoZj5VfHToDJp/+cWeM/Q9mdisC+JeGOiZmS
gI0YzeeLsMNov7mYs5F5CRBmrEUEe0vpbiaImBXoMPDGcd9+dAXtiUuaFKN9iaJkWBGSKUIo2nCY
qOHIU5DG6Jk/YmqGqo8HMICqYtTt+WF00p/k6kFkwDHa2coWRHOvjD9AX3KFMVhG6RV38bmmExmP
f4ZYn5XwB9InbebvUdd5t3+RltkXPXABVM6TG0PCZOSLJgDPONGIH3mZ6OEySMzGwyFkoghtIUXI
isASt3ZDhXy5mLKaRWDUCEkLHzRTQiNRU0vk3LxAAjhTQgJOxM1BvEJTqvP0XIUQXrpIBbSr72uA
IeQA3ZNDfIbtkb2s6hjTZU6/1wZ5mH7gsiRKjfsCsrpdF4cH5XiO5s++qzBOFSq+reKg+zQV6Z1y
Zgg/pvwS7/+MnWrDeKBx9qDzME7dmma5inb2wVd9pfcKVTBQIjotoYQB6IJHnUJwKutOK7UdyEGU
27rHydEbJh+w9hXAn9MRPCsKHI22yUwJEl8G3z8CX8pfa4rhlDfIfJJFMqMyYFJB3PL9hXjyM2MJ
IQTgSv42ejGPhLHRa+Wwi9FfZpr4Ldro5GVjRfWPPlcBebLIb4iVF1OCPQJJ4tYb/IvYn4wAilAo
R5DfEZkoaDj3wVhbqhxhBeAtZVUNlfDyfjmuSoyomUBhX+nLarpm6xOKI1auLDm+G4ISOgHzTxBO
i2MBWhLPoJ/qehdOEaxA8ElEQXcvejiS9N4WeEN3lVpeQKMP4kyImdietjjhXpyGOhlSWC31xxBa
tPrpdCxWt4yspVyxhd/Le1vhhEzzIcWvbqOOCtfyQKSmAqGEIZ+d1/hdq0372hAwBmzwERL1iBwq
nrjl7tdWgCREw1rAjETSkZo71v7i8yCB+t0YdLdQO0tseCf0rJAHm8JdzGExk8uBSyPxuOrpk4Uc
WR5iiji4tEREjhw2F/22jtmgBRhJ8hfOtQB8Pevx0EMkyk6XKphyXlR3C25+0hbtAuZdHQDPUTQK
WbtmV6ikDvnpYpSf3dGoh5BwtyWtCLy6RpEn7upBSd3k+iYP7+bDx/flTqTAI/9TLeJGHcdR2HGt
i7OLEGT+NEFDeGZzXcoIYa/i2YgwEAekoxgSz/erVlS8IAPX8HtB+YzHgh8hvNbLVsLBNh8svmz+
V3v2A1spVQqU3ybwqDSIASjE/K/v25cTjWXhlrm+1jciBiUw7Y76t/K2766q6ESP36ljMMNogR7e
s8GBqTartIZlbMi3hk+yJtgrs6aRp9iVfUdvirScrRXjDlkoMUBQ/Am5URafw2SaHL6jCy88r8rA
Il6PZUMd09EtMjTGEizffNIynPQc+quZ9n46XsSTBASnAr/10XQy5S0ZfiB1AHoWvUSAhPCoz7iu
wGme0lsZ8Gnn0qBMwwCjzfbrkip7O1fw85ElyNnuDPiy9vF0SrUlix0NeeDBmcmrZNj8fLwVkBR6
vW1zTb74rkvvRNQdgqk/a348eT6E3HfnHbiLw7nRu8fS7HZgE527TLiuTuB02EdrrcDoeStRdpHp
G2YHBVB4FDxX9yv103f4IetkZEqyEgt4SoBLILM2k2nTRKc6+LcBmB4OCR+Ammjyz19vFuFEN3V3
smhwc4yZa+Nyj52oPIZl/+php09mXDgsoaEFPbVUlwm9rysQoozr3AHG546/KLXcDrKmWt+DeyRA
clduVjKdnEGlubMEqvw/mv/hXU3zgfvj5KxgJNy/URzVzPaOSkAp+tmxdGUjWZu6+A+2XNH4LWdD
vW3pje8RoqR5vIvsGYgNP4MTejkqqtZqxwVKlQXIB3PVWKFrxPfhT1RBs8TE/aAwwQEHuxiFNEVJ
LYYobAX6X+JEIvD8YBGXUVe6erZXR4xpTC53b16SdGFf2+QAUTC90xB4fT7ak5F8ogUo3/S1hDxm
xLXA/KUCWJoOUyxxfZ7o6viMiQbitwdo3gyOmH2gXUIbo/de6c5Vl1ekoyJkeQhtNpRgsJmnkQw4
YZTmDvjpGydmz9MUGmjY6MRy28rYtKkZtWgJQO80FokoPzX25z406mnM3HHoqTBCsPf2R15MW9pG
1t41AmdPp3WicuMtZkE1Bv6LecrQKyTwbJi0cQPrEK0uchXWnFIokYOedn3JNUsNZ1LTkhukt/lY
kk+D6w7XU0kFXWVUJyf356BEF+y/Z4yHvR8S+INsVZECm3Gv0ycRor4ncm8NLgK5twtCHY6HehWO
3tASiBrG5+SzMLXGFq6ArtYOYUjqF7cpsQY6Ugn+PBWU/qdcG3CM/gqyiN5DLiJpTYqwVJ7cDSNM
82BEPUEnbP/1nhPPVw+dEYvr7zZ2dTKwB/InBCRXR4yxA+Q5aQgxwMVyB7DILerKqq0jDDOX0JBn
Xvjtw1UdYjLIkxehN2eQCswyEABM5ROWO/dsfWg2irYtvWN7m/ODWpFNzdA1N46rkEmwF/9h5gIA
JiifdQoXuxTIWC9udfAyufzQ3l08ifpUwzKemumk3e9mlaCitUCIO/j9fC7lDpXow27uh0JfMtRJ
/jU/mEWjA4wgSn5Gr1tU4t8cgx2BKKFsjL8AvJlUPrEfMGN8FbbBqzR8qzx88HuF0iVaBKi+hTCh
3ofyQlI0UwvSf3ZrgP6LCAGbeRiFoW5px4S6HtAISj2cscYjXkm8IloQWqW9Pav3lOKE1Yxyu/zW
X9dFRyksa8E3Vk1qkEIyWaBq8tS/MuQkb3J7tsXgFzkwqIf7BWvVGYrqwHkWONbiBBOJbp90Xg9C
nrs1B4yQOclyJRxomafpBprzjr5+mJ3nK6WNPuSP5Ye5nSGDTruI1Ssto7Iwq4whlav206T1lZug
pmL8NvLGe840kPylhg5iZ0n7Ge18tk7LGqW3vWUOCl2ux8mD4O4BsBr7/yNSmRDm33Dg0HBp8MJp
J87tALyS19Bd8qHXx3lNQAOS2MewE4Umkp5h9L7nvzVcFDO7SIpM3ReITB5zQxW22IlpRvdgOEvJ
TO8y5ZmsmuqSiHdJsdUolAXtsdM37GDDBHrzwH+mItyc/bCM8ZyFsnzC9Fhxd3nwOiJyuyJNebXd
C9/XQ1nVadVL1cj+mWVOjVjiXhnqz3ImClF2nfuweUxwTah8GE72sgZPwrDAJTwyJlLIxr2CPiFn
M67ZKG7+b6caFBaLC0ywdnMrWyW7jt8jNOfR2ui/DZ3DHJ0bXvfnXXMTk2ii6rxYgE2bMpoYJMPx
4ZVWnWX5MvlYQ8CngOzJtRAbrw4X2KK+OPgnA065YlBVXg8YZWtHhaRpeGbMd79MVCnWmlzjAZ2j
RPd18FjAAFhIaIQnUboO/alS2BRW+mF3fFkrhcRxmva43tr4YYQvaQE8OAkejl5rbdE3d9Lj9Mq+
67YasGkOa/lv/DZwcyNYd4ZDrtiTQpXvocLcrWtBbzXmzzQQrrYP0eLf35qktMN0MKhYxr0jDBI6
zNpyGJ/n8J8p0y5BWXWEgA0wlEcnzRJNDUuuPgBy8vbozRed3t2qeGTtSBhTi+smZK+u15SeFs1T
4Vc7O6o7LnazayZUUVnKs6PTuR4uNhz15mg/GR6/k67FzCzbJZYPiS/8Z1eqhybBQtGD+KU16KBH
DpLkmzw4kELTZCVXfjo+bL5RofMntMAVxTrn0GxiPUk45EuJiWU3xZOBw4M9Cg/sNl8Q8S/Pe0kd
UIhNW2b2jT2lCrmFsfJmcHbFSb8Lx5ozKBqjjcrzVCeI/eLByygpphW7EJESFMOgyQ1nEMuYjagL
ygIYFHV+lhlFuPKo1xyrLzZhaEhZg5qUK0LLlmbITlb7L3aFDGxYQdHFQgoImIWWPsHGnYaFv5QC
Sxz4+UtkGVKjU3O9R0bxHtKAFD6KAb/KSRY320gXvUPyXNEEvRMWX/ajh+srZRT4EhRCi+epSBS3
qUEEAUfAji+UZTB5Z+3ketW9XCu/UiMdBpF/nZR/Avvsl4qd6f4Lj8NgcpSCE5ZNvz1RQdcUqCOw
Eb70NGusH9TvyeVmmu7638e3RL+eXKRndChAgxPw1XR1Zzzp3lV4jLO7Mws3Yg/Spygdlp6fqwy9
5sPHjPtK0XYEszqV7gto8iXMNUbg9HsG1b1lDtEkUqdH0r2k1Zmi6Ip9A6XTIJT0S68ll0VBqhuE
4Ct1JJxVWy5YVVfXe8NlsreWm/hM36NcHoTOyS8eSkm+MyviqE+XQDol01sorC8olM4JGl2cg1kg
OHepNcit1aeMCthhMIWxpWfn6GW/z5vooMgNU1Eds6uBtYXB7EqNdhxnPXp+MsUplm65thdfsIZa
Y8Y3bnHCbJRARaZu8Dvy68WTL0d2l8h9iyJol2s8M6xdKDgSw09tW1/U3p0dpkF/4hIEyXH+AtpU
bLxRJSZY1CZFyWp3RLCphOan7zLaJnjB24Danw2IobVvmNSJreMG7pVKKGPk4RMhUGLphvZvsbg+
5+PVJru8spiD0k6xm2WhuUJ5jXbeMJb5FB2Dw/F8jWh8ApoPaOcpPgp8O+Ne9TioRYder3Y4qFpi
urh48TOaaEziE/Z+2LZxsIVqPUnDCJXzyv6an7xE4XHBxgCA8+aiLfZWsSN1Q7+8pOfvPtY9VZPt
14EIh/WhSxOlmxpeOqveWVcZnUB65J4LMQ0w7pA8hIjkOVZdhaa1TIDveFccji9vgp0ttTlMDyT4
tEkwRJYgQPKQgROqWz5KjZQnl1oFkKRsTAAXnwkjGLgUdkN+zLF/195LhYEMaop+HC02HNPQi9mM
IaXQ1XkZiXnTf81MraPtQ5pZ2UK7vSrdthrLwVNT2KqRm3ZCuIjytr0rDrXSqXD8Iey5WFRkpwM2
T8eziLNeifx3u5Dd3FDSlpsj7RzfYo7V4Hph0NSMqDi55jB6eGUgvb2xdUphL9detDWhH8yyXV1S
JvKIBWN6ws8M+lB3K+36frVyKZgFnZOg48buSZTeeGD5Ua+GOGcu2JJfQ7nAuUipfFvYE/hlNg3w
5vqWzi2yq/LITQB9ngczx6ObmtSCXJrjoJM+wkCIx6Q4Epq+jmLXAGB/FMIYptvL5C7ksGHuaBls
oDk6fi+S/pbHx24dVBjd9EDnIN+tRRfeu3Q/YDhFPx9iOmCJC2bMI0Xi+xLkAWIRo4aBRXMq+VXD
TjM52hMORH7EV3z2XQyxsHvuNefOyd6JKe7JkSjsEQDkztEofIY3XOim6bPZKVU1wehIdKpCF+75
oqOgulWehCnSJoQQNUIvWiuq/kDxFgwXlYKW/6Mq6Frmrik8r8XZHCb53Jm46I8cEbFPWUdaVEVQ
5+xHxUTh+ACn2jrIyBknlBVtIkGYd4bgo4Gt9+bjsQt0+dGhiBXM3dSpumywDSc8DQP8qCAAwpI2
yvlIM9g88VhZUUAPowWx9ea0jDgg9iUZm5hMP4pXxNPBKNmDyV7dpJSFU9VofBoPncfP+OzBi1dJ
YaZb96WSPiOcQwfzLL1ZfbU8ocl/AdbWLYNCJ7Jxn5jStHYWKBelSVbSyASqmR2taFfVgrm0g6mo
MHRSFpwIduqbIPp4wbCw3Yh4yTshozZ4JT7ve6PAL/nwi6QW3G2qiv/8AhRM+NZJ/rB5vc2XXeQN
MOGdh1Pk4aGTQ+l2dJlD1edCAClczXWSyKIzyBNDhkecmsUSe4l+djdFSomk4K8oKwgb7Cx92ZsX
R6kaRYebIUxFxHSvJlPQmqc9hdb328tubL/rVT+X+uV9UKbwVjLyyWuGKMMurPLcTfIC7GkwFXb9
L1UTijrja/l1MZplOnozUVDPixfh50FKRM+J7mhPHjNazeCEjcZpZI5IgvDJFZDnw2la7coURjHT
ZQB93QlTkAGDCqbCARudGShGJQ5TnUGUlBlZ9tXc4QL6IcocB4dxiLTrnL1kujxOS2XLi+mKdqJN
tP7dYkb2sD9nVJBuoJ94HVUMdDiJPv4WORsa9/Yi6+FHyuuqvdHdhLJxgWm5DAiAGiaSAudPqxie
UlyoL/EE82i5WjMAQq5a79NJjzTk1YCb/0fHDxgzyVbLCV2TF4wQW9bA/7mjwCfRmHzi/ouoV8a8
xVa5SAtkGusyJGH5iaIwbxcD/vPtYL0YLstsBm1yG2648dbJ/ZKjdKB03JhOCQcmiIZUV4WZrFLp
sS5VcEK7+4d7Tp8m3FJOuk6slfFYkkS7zY3ZQaS/qvrVwqRhqik6terbOYziZNx1FKKdkkTF27Rm
92XSksv9VVC9w+vboK1gjbh5BSeXtIhpmFgW0V1DeavGv4k81vK0FPzMoIk4tTZQ2j0Pve4EhzBA
pRBaV02OvzCQdeYYOWNMP9i+SneVCXd+/wlDWZmhIn0cw2M9DXiXGHxwl0ONfLy47xSuZigPtfo6
Zp7Nm7lw/taCzG39s6atfYtje6jFE0xydDeEjhSlF+Uxn/AvdXjwQ4jZ6C9StsYad9mi7zz3m9Ql
62ksEzQzVJcXYc6bds8R9aFYgjWdC/F/l8Hm8F3ffy282BDxmixNsh9Ptr8vaNY0DAI4Y5XABT4U
c2Xx2QgezRc0/JGDHetenwxIPOrETx6cZJ1Ov9/JB/r3il4Dq8EjQfAhui99h8urVD7h4Jhh0M3K
34sJBo6RYNxzhmJ72hzjhIEZ5gf+s0sVBJnGwnTK6S7yIS4JWwXAmO1gbYsSMXBxop1Jz/0ZozJI
iphK6xErBgKqP49JuUBgzIX5WkZg0v0Mc0XyCJ2vkTqtp2LEeRAqjLLmihfjPCR6UsmVQQhBr3f0
uf9UHroppvLxSNYKlFbVUAh3pEoGPyaiblAZpBb+0FVlwjf3HwrlMsnz/DUg9Cwz+GNwDazDxoCB
VSVgJ6F2n0KRtmKSEVDmICh7OFsl0sLSp59avXD3K9YxsLgWtfkhIkfXSU7oLO0ssKoWrZJ2kGum
zb7FS3Fhm1ZNCsN49scRol78WnVrA2SdAIhjun86KMa6JkugVstwQNyPYz/ElTRHOVmFEN5/DaNO
UY7ValO1MrXeMsOiTXHavAFnWGWzKFBPjbz0iIzGxvDKNaSXTfkNgbHD5YydqqTLG+X7+iGkykxZ
h2c4HyGtGwC6L6s9NXyW4iGzUL66jlF73w+zUSOzLRf7cdnbnpy4y309sC0NLpnuBnitWXlPkaGY
KCuTZBkky4I1xL1YKC+xOAVrAjN56vfsJ/CRcuduWEG7BgPRNSlj299P+sE/yEyRCyFgQDE2ejHf
kSR2g2ngo+8V4p++yrovwvyVjXFurGv/n4JNHVPAcP4hftSzir6YYLeoUZapA4kjsPvMuPH1MKqO
ovPOYTZWjNuyG4beUaKsSo8WkYKHfF7DMWEWpn/mWtlcKN/+88iOL9FfROL6/iF9pDcqAoNK7SuR
Mvg4kZtmBJLf0BBUABulKW+sQarNkLW8xTaKr2T8JznPAVLYkHuq+/O4lDuNwMEsRWg2K6REyuAh
au5eknGVSCJZKrvfRxEpiCKcq61mIwP+DuTov4CePyPZkAQ+zsGpvExdPHAyL3FS5u7r+WayHl3s
edrlMza86A86M2NEabAs7tMf4rlYemOGpPKHZ0u60wkuLlocPGPOEDgl8jr+ieCgqwxQ//0yaUPy
zYbcvZk8mrrdIC3BpnQaZMDrIUpDsctMGxj6hFergV04iiSM3cY7aKngn4wLPdFuIT53XIZOdUfC
UhcocGkf8iM7wMIk5J2ZTNjFLpJIIi7C/GNneUxGoW9b12ui7kPwZtuo3uOALpjzGAu8BQmvDGMh
zr1T7+dl0RDZzSsFGdSr/XU57UVZuZfgmnB42PYC7z5x9rgy7PV/xcnCxGCCxh5Y3BmYwvpnosdK
+ugnIXdFSOAEp9k+uDwIPbj3DoHdWJnItoBVw0Av3ynQhFtMn4rXUJKp5gZb7URlUYztNyWExtO1
oFPgHedmFjjEo6Kw5ME3B0TN0iKHeV6KtRRcaM/jW9HdIfl4YbXLbMo7iYaEC7GnEvFb+qnSPZ61
FRlMDqclj+yiDCBpkyn8PC6mcAXTfsZuaQ8zx0AgyATm1EqajaR5O/CSc5SNbPWP7py6tvnNP/If
RlvuO+ZFy7wQwvJoyZVgfKhI9+q2d3StQeAMUwKERD+JTMpbeuoqnfzH14GTzKx+gw//6rPn14X0
/WFmAV+dComEKoWu98maIY/hSCPQ8NKiJ7pPzh4canr83vzaHV485cuCTUkb46N841IkCN9rkc9f
D3508mWi5PD9HsG2zs+dCMfxcYNdNvbqk2LnkQzuDlw+vGJWLHPfImz+EV5OhrpvvB1TCtCLcDUh
Vb06y4mINVwT+lwUNfkMExeOHufIbn/LyQ6N6FmwmytJJQHvtDp0V2OBtwOku0jOH0eenNN8bufJ
MHGPbn/47UBq9R8YygOq7RZ3XN+Twf34J6NJgiSmz875q6/f0OfvRTAmOsLtWGnc907ngEtyZaV8
/7AHVvR1QY/TSolbsFnrDAx3pMH+V7qcJHNty3NRHIIzIS9yXJdReC+FzWvd5CuLOFF5LZS9ZdnD
y1o+QRdWOguKIcypXo1je6GjBOJEKNm1T2jPvHGrSZu6rLiAYf2pdK+WHsprU3RFn/6ecjIjXoty
bphhEgUE0PPYuT+mra5cNLDoGBNbuzNMPsTiBn+izsuwp5ecmVtt0CIs2yFTivvNj34veumJQ62X
3C69LJFQUijG0oGzYnq8yYhVLuuXjS3NcybJNyKqicve7kh3tRXxFRAevTr3XbLvNCat2UvsAiMH
M1ZAIulP4JPcMlMcHnBFS8I/zDZcBe71mgUPC3LdfVzE3ulSzGK/ig84ws9tuHJZhQW/T2Di5zb1
YAx8X58safxNlkSAOjnKHDPsvXuWSjmK0qrcuq243f0GZ7lF5r06YjMOr4jFoLmgoHGCOl1oQBxt
dJrjBRBjM3V1kpIT2XYUvuSzQgBjPwh5/V1NUV69YFYJZGdvNplWHk6EST2Ipi8h3yGwt4ryIzMf
phTKrt/X4/nu9TCHbVF348qUZqyQN9OOThP3GsjcrmJvXFdPx6d7QEXs6J8ij88BOJMJAV9n7xyr
sCQDIi1QLCO4NArv4+HqXNauUKigDhjMMhQ2GI42Vm4cI4BVaG3B/aMRe1CXYOYGut92hCf0PU/u
JKgs8KrDto0n/QJrDTxSb7D0xcHuQaEUk6hXWgokD2RW11kW1VVnptkUMdJw82LsjCfc1hB4+ZFQ
897CHkDcs6RRfKH1yWwSQFcsf8ITLvi2ak9z5ud3m3n14y0efJTXwarwKVPthZqRQsidb+sUy2al
8VBxtvladjtKxPWbFYYGsy3i5rzFm4LDHdkHEdjaBuRM+BwVXtBcGNF2YTdnqU+DJyOY5pbY0pJg
4ZdbKlfXgqkn+Yzb8mSmaFYqi3JIxuTPk0208obM5YzYtNALewI6MaMdgNrd++BPCpVJsb6w1yyK
zaBWcs9c4Zz+NuEGB7E3Pi7+XsSWHb5UexiVvr4AAMLkrErWE5/d1Wnq/iY0I45aN/k5DV6sUIas
EN1Da+j0tkjxdZ0S1fQvH1ASGKb0UQ+d0BmbrS971gu/skiStNz9B/PArzHyjWYPFEuV8VoTQvwL
cEOno+Q24TdO03DZxhso+dkuLIB9XGyGAmNE1MhSphaXkeDa9n/ZhMgbup0f2qWw6A2QS9gm4AT2
m1r/SQIm0m+2uUINwto4tbNhfogmVbSVIi5eE5lgzPxVTdS+NaFvUy2r/hn15nYrlFN4h4UkQfYG
W57bjGwSydIUQ5gWqdYk7Jv1QbMDegVzgQM9WxgxrqXwNC2MdBBJ0XIdtZ8Zb95KBEH8q7cYScHa
sgOZzcVDSDsdmBsBEwcuAi69g0b5NTXEmXy2J32AtN8nnMKeTdoT1d911E60dnTY+E8CoQKHAFvb
1Rudj/58xn9OOvaOhqF8QGnmVHe+Zj+PlUxgupAeGF7gDkdOiVZHj7AzNN/suN+RyOuRTWz2hbtU
hvVxcIx9F2xMnNBWJdTfv/JzIdRsjx42vWSY1z2+3Cb7qPahNiyRJhjeHK/FrjODA0Y7xzkUqwCH
M/fPr3n1F7NeGVM7xFsogzUp3r0+PIoL2pqXrVCz7/YQWbpIdieAlWFJqOYp8TinsLiiL7Cu9f8f
g3c/zdDAfXI/pa7USRq97x3qbvMAtnnWHmPUzmWG+uWRLwILtXqQahRQYrOsRbnZJiPxVK1eL2lh
vU36WMVptpqA0mOXoS+aWQuQybP4CbxBcvrDUvIC1Gz4xLeJqjG/8MMfpwOSM9ojKvbBoL4BgooN
ZhldrO3stOJJPAJv5nfnkxx2eN2Dx84YEdNlqH/HWAIVUJJiofVu4dGu+aZOSdbZEC7sMo1n5bGO
SbnScRWtGX+/09K/Llq/ULOjVKgGZShF7hm7c+iuLbUzX5znCAWHzJn9WkPn4rY1738DegcvgRJQ
Ti418zRij2V/cVWsDXAsBhK1b6oDPCJynov1UM99TyZ1cck2SH7jUMcOSa91SExeJX7NVQTOXDnp
0oeCycifq6PQ33S59QeycOdCRDHeIqhRzQRAOdVyxW8oV803D1juyXC8BEQDflPoN4NsZoBSPMfe
duNaahaAGaTq7Cv/6gfpLJUejqUXeNVyIffHTtEJhFi8RKh6d9mPGPtD5RDV30PQrmKLkQloW2Zn
roxXeLETb7Qtr7VhOQe6udPfAzdhRDkIXJ5H5hff/crFxUvlwzHrhHVb9O7NDWYfC25hfW5cw5iw
TJPTkvqy038ecnun7aDRpfZPdnW73Aaz9a5m0qmuBJVHEWIT9LASqooBr/rC3A7827WTpdcOfbO5
SIYwqM5O0llykC+00JOWzcaLVPH4ozBF02xLd9aig+sZxI9f2av42fNfAhOt3bBLoAd7hihVPauj
Fzv6koO0C+qc+Vcx6ircDf1SREDBazINFE+VAOsi0xeprQycyrI7wxMsRbnrzt6l1QppEx7l+cCS
6p1UrCtyH2+I1FLbuUiQKAm+Pm37z6Ds0CBGOLiPuruPJPM53rqe/hsug52wqKbgp6mqyxmNFQiK
exkZCiyan457YAIKAkQtKLQzfGTctMStqzg/yuwtectVzW+nc3xM7XK6WsccufqZHKewCEHR6Bci
CbJBl7qqp/cYKPAzSI0oN7mm82rDBZG/vaG1A0d2D2oY2QntbQBfepVtdpo+9FgOKXBs40XGmN3p
CdGmd59+EaR4Zon4OohcVQWCQZbxzOsiRyXzO0QmPrbCDR9Vm1SmJtu1ofkjIXBwviUp0bYKAox/
mZjAYrrfefCU3GV48nxzxDE+tn4bWos1ck+48SH2lRLm0oOTewvBoKiw+1wa2Q0koXPP/SwE3Ug9
C6ENBFPTJ5/84BHIxOOqZXMod6rmnOpvnGU21U3cGvwvhZvzKeASN04MVpYAvDQPjgVmwGG3WBCm
m8QEoI76HnueDybdt3iWsqOEo3yw/9QlvbBqQivywwdnjz9I5UHsDz1WibGcIlj4E+ROfYE/n/y2
NNMiRpuK5P2hOyTtHJe/BT6B4D3vNJDnv4C7EAsHSsqwL6quS4I4f7SjwMIwP/E+wMtMaR21acc8
KBblVJl7aENHvEGj7slFwaXFr0G0Scy+Sdowjx4tHM0FW4mtGbS7UCmo0P7uK8AbNj03EZ1GI0Te
sDSOfd21d6l3FApOX0kitM6EK5uS4wZmNlPo/ytsB7QS20wLjDM774lKPC4ytxWg/ZrwdLT2j+i7
IQJiiy0qLo6WYqsxg8wiwucmSyIvv0fjaePXz3M4nbo8Gbaq0JYrn0NbfIuu2A42V8NMcVioZua6
VYlsRe9F7aKSpQIiuV3sPkXzsO9FBfzVsVOHkJXVCfNJzgBtlM4JU5hhx9E0ReGSEakbXgqXSDHr
sFM2hWtJ3wpHvaZimNVCw1LGRhb/c5GtSD45YDo9YV6Fw25VTEqrtToOIEosSYJ6KjJtz2w+DgCN
6dKLRWsQ3m1N4JZCDOjIAvnZT+Y9c71sWyrlQeeua/5Kpz+Kf9ePyLUfssFG99T9iUem1CDToaS3
zAyEd7tFXT3ePrm7frUQ7MOAYa3BYXrkn7kNomOAfSqp76L9rkDWTkH5iaspd4LEHtsvsj6+1rDL
/84W4LQrcA7ykdYN3Gg2RTDXN1QecrgKY2jb8ej4/urZbQPwtuY7Egn7pVIXu6tTdDUdkESlWO40
ULknfDyhDymIeuUPwkXDDOSxmaJ1RDIDrol3nZZIKV3IbtnzXQnEx2bHN+Xul5qbmVQeHkjFp3AJ
uTRk3GxKYpB+OcfFQF1rUOUb3q/sF7INCJHDbqIsWJkTrojHRAa5tMtqKjPjpsz18J2IQ3x5lEid
ueKLNrXo5tmAEo3MUkb2KUxTwlmVjvJ16kDTuxqC6FXeGzUsHB0TWuooe0dVhlFlkguiDMdpfS8z
HH70vdcW+Cnifhd09LXSTsTRovbP+mXYpgg9rMEsfx5nQrOYtje8d9PKF31nD7dLsv+7UH6WdcgB
ZENzy6HOxYlZIzK9WoEBxm/yuXIQWlDJ86NZ7TVNAC4zeDwa9ipM2AVSVwhxjJu0gyGYgvSdN//c
qHbK6lHfEnPR5rE19hfWkMVqVnONcOV1dcKv/zh70p2yVKPhvq3Mvz7nPqhvNhqXsRo7iW4LruLa
gMbcYVKC2RUbODVfAjo7v5AoJsiJgKp1/N4lXDzzcW1uftof+MNm91IWWTLfjKGEuVzZiK9lYERT
LTORw530VN1gea7DEmgUETTD+GCOfV8Da5/fjqa8BDCDBuPaZa5emiZSZpzCTKHwJJb77UaFC0fh
bx9/AvAzsxUnVJyIvM81jqAjXsnIEICAYe+R2dATE/izVhFO+yAfim4tPlRPvBfJOX7Kw6xWrui9
YEZxBA2OYioQ7LYTMWWsx7UHWAya0/3yklepcuZh1mFbuNaROw6f+FsZgnvyWI9t4lptZZwYAh/I
lpP7q/Crmz2HiakvnAvej6Q/W1SelMpH4I9kfkscXTgWL9kz+E/guvVGDKY3Ou3ec3c/yLxsWwA/
EAUY/19Hoz98pMcSBT6JRVRex+AzAqmbjvwKrIC0wDSv07MclI92rdXHCjk77dvfXnlpurQtwT8Y
UJSvd4i5w0DrX2dqrrmeiEqtJoqkWPrfsKRO6QAdC5GMHxysZwr596mEG3shcwYIhwZsOFtR6x4j
i6vKxOjKT1Bj8yvcmVNnyj34XcrJtAfGmTjQTbOrRSnLM3jTagbzXPFmD1yCKM9lOJOuZxIfZKPY
+5H05/IgJl5kAQdMP78VuHQggfpl+V1+qELyYWLU3eo/U81yttRVJqh9Qc5Zhhz9TCaJogSSoqME
V0uE6oZS1E/EcEWHXKBiH1re3927TajuoC9p5vUBc5F36y0SUSIJywnYofezVKNd64GziH+tAG9d
eASDZ3Kox6sKnNseoK9XmZqHedsG3QA77OQmkZHMKzCPnE7sw2528kbjlPqogIcNgSSmlCJXJsp5
HGbmkoWJK5uB7i8H8Kv8s/A2WI5JfJZyocB/QKrkyl3r4wI/fq29yrFvkJj9LtUFPHZySC10ozAw
9jWP3sd1xL1ZcezIivABwr/RxvMoI88NjjFc+SKWBOgQnDmLqm9jMDv3gXBZm8VR1VRmCzWVfQIz
LEFW3CMIK9zP64Pbqgn9ykVMHW87sQTjpjvdCy7i/byuXEpsy01KKzAWhVKyMa8YvjHwQ22Tt+De
oWgUd6MjOd9LVxHxnVsjPFzCUFW2zEVGAnFfFlk9ePAqzJ3c6KYpIuVhdFnCxKm7VxdJ8wF+UOti
TC29jXGYRqwwKHqkhH+lCibH6j+EMfsSF7ZBoBLwEB4icVO7jhm8lifpYHkAwwuvLKdurMEzoUdD
akTRy9SM/h6YVvxY5zFEJPTOCtvlwP2WxOS/nGBF+yZ71wLHYQeuPDo4wGf4UwYCRxJTi2DeJQ95
7E6YRtTcgiQBiGvLSN/0ve2HQUqyBQgPvz54Q8wnOw3/PK6APMhmtEnDcdDD3n+BV8fGyAuRqX0Q
im0Q5jfx+5RuQs3f7Co7jCNTB0sfBpdDp0W6S0vOnCptPlLZO/YluxJqPY3UjJRk3rRZn/PKx029
RSBY8AaneIRyOaOIjWX4c05SeNTITEWBDMa+6+fuQBnrx7Hag85uM2N6yDmlrAaemD0BeK2ZBGjG
A8qsBKJ05U0Mk1YxwE0ud0Rf0CE6D8Rs4aq4jq+sMUcyOcNMqP7UwAeNHswVdEcq41nO837CW/WO
jm0+t326Dzdqc2wS0Sm+zgcFvcxaRsUsLQ79Q8Bc9raGdvmHK8abjmuLD5YKLkpwH68/sEaKCvaz
70dAPG4LJnwt51qduW48dIB7M8+rpBo+WwFFNHEyFTAkYxYzW47h3yDFHtMG1aK4BGeCNKjghwZy
uXqz55T0FjAYiDWydfvvtL8Beah0GCIk89hPPuHpKnmv6/6NOBolpGw+qWhWzg2uoVDNkI9CtpjA
NSHJWPWF41o3yz7xL2TnJ5bQ092y/hxEUPJak+otfhP1z4wonH/HwtVMb1l2Lqua+ZvAkvFDtkDR
4UjPrxm8d2wDqXh3xjNpJkBNTybnpb+3CEPjiRiNJ/oQFJKAZ9Tvnx7cxeXpNw8UKFeY3lpOZXMJ
B8oqXy/f8nXAw/vNWX9eDeaLTYEaG8CFuGMY/ffja5UXpIJ+lhYoN3Lj0F82aU6nWRhziT7OmQ10
4pKRqTnLQM9h7MRtJr00sKSmt0WtoeursMKRh2QFNdx12dGi3xf5oGJtdRp365NAxeVWgR/QFAgl
hZk6RtwnY7HK5xwYTgwCOi8FdqtNFmUCsZp7z41e3nN1E8a43TXy8wsBIynoZnslnJGKNLdYNmXD
vkkipymSES2F0jg9JdbXKnFsouUiwc4CnZWDYQD3E5kB89J5s/NBw0c3CnHTQStTPAZpN0Ku8Oyc
B1QduoQpRIhhuFejeFHQpFfamviqdPIw1H8CJqU/L/U6uCSRhfyIFGUmrlxPgWTLaQIM2tB9EpQL
vwmuY1z00nXSH0vWLK1BRjc6bAmNzgyvqaMDBSP4eRproKgsa6Ls+SGREcjcT89DX761/Gfy4ATI
9sIHer9OJLrc5j8+G18D18vShPr5/sXHIQoorf5bbH07hXFjPuElhaiJQRVops/8vuw4e2gyN8Bq
E2t7IU/oWQPAfNvx5Zpxn0mi7vkKWeHmLIUkLrTvsT6jEcXrDqGR0nk7UBwpsQCQDKlyuvUd3txs
JDRGJWXiggg57OLC1xLXWC9HwPOKbFjBiclUmNsZDjqcHYwtdk0mXmRoWbcVAVskJqkAgjuCIgcN
xxpnR0O3Rj8UdchbnOsa/zLHTDSP/sQm13yR8yni9ur/ivRR0OyapHwZtW6jdGWbLnpCem2abaVj
Qq7loWLQN8DC3a0qIUC9fg0KhN11oK04GUwORyS8Zlx9Gs6MpAomiIq6Jz46muNiO9Zgy3bZYmNO
xq33riTmA8YegnIxd1f/NmAHk9qRS7btK9fsEj44loZx/+6KBBuaAH45Dz10kwTyQ1HZqYoO6RHN
5c7jHrG2B2ZU1wbPmPeEjA3/DlIg8IeCXMWG/ZGvG6SXIzWWUfRLlUvxjhMQJwnglA2k9EQ2OcNK
Mv3hqbwFf2XOGLRTLLYWDuJGHcll0wtTe2Z6U+jkHphUdCO/7R6qIrV7CJT1c1hmqIW5hlmk5Wc3
tgNNa0Q4tdyneRhihVHWFG0/Is0RRZtWakRKn0IIJQ2sph1a+q+QFLhTMxVTU10gc9CMxsDtM9Ze
H2Mgge17SELzO/f904ySM1k3AromZZu+8aZnn3Fzj/zBv7akhdBFTXBnDFFpz6S63hJBrM1E6yuu
gES9z9SXeWC8np7TCpwH4gi+JVqLKAgLJTk0PwZDTKChhtU7ryZydoYw+Clbz2NfjyggcG0cekhn
uvo3hI0PdyaMSx0htFfc6n04q1dnbvhbjDYdPc7lll6hjyCSDJg2zYVyMyCDqaDyFUIjpuGPpYkv
UOlkCKyTu1za1lpJZbA4NYN4jqBOYfN726NhP5cOs8RRbx9L/hYjc9zAkzeE5PnrJCfF4pwCwYiz
MangWS1Nw4oWB8xI4ugKOxYLTt8LvSV6pYNZDCX1jCcs20EhqBr7O1POL5Mm0Aw3Kt1jn+LCeKHv
o+vPTlMILWvOwCapfhNCLOnj61MSYHvLkiaxAeQXOH3nxYvxc29+Zos7H6yvORyEZJPtv/89bi3J
jYuv6Tcr9ljepmkLwvYhuva0KLmNlD70k5mBh3SgRmFChxVTy/w42ZJM/2VEBc+4zA5zVGIW/ysf
jj8UgZsLiL5LDPf5Yl967HlyHZc4MEdzTyK4tU2QGzKIPdvqrBb7dVPdQgA0HxVmwSbxnQJfI+Kk
tXxNBVcJYgyaf5dnBDGJnWduoPwPpU9UvnULxlGIeFdBxSuOZliM27HojRPmXG8ZnHGwNrh76SSG
u3WlTtm8jEoHYtrwnoZbscG7BupdL6N8gxWFeWrkVzYduQsEggWOlhQ+UHKRJ+329yYfAwlwfTc5
h08XPrQCVsINDWmMuinQ6DLO8uXDSWGBqLO0wjT8OIdTRAdOCj0cgfR09l9e+mNmWJUJcfnJuLdH
SRF/qemtcE2nR4ehPRnvypLSx6f2qEPJ7Er0q8aQGkMCXpueGHU10lNHSGfeva7+nvTSndoP6qqi
zpfGyp0CgG47KWm9Huqyb3ialioTlkI+auJ0TN9TEtjtEWZVDtfFW/pw6pXzChals6/8pUX4Vr2M
naRJ0YA3MS4+yXKWXUfJu6jH6MjfqdNCT8slRCW7PnYm60pMwP9qCFxrJDUnR/LnDlmbK4dyFbze
GfnDUpm0S8SWRthq1LwkCSl+anFgiNywb5RV2F3rf+uP8S7sjtxG8woxGuQhXESoqYvmk8SvdeJH
Epr3pBT8wvgDgx0ezR2G4d4a/oFO7HI+GaPJljg+5ksFOX5q6w3sk2/+X+2F62n1YmblX/XYQzO+
EsrAw6Tb0YBB6NIpY1qicpDPusQgvAuH3NcTlN4uK54EbLlEeeeS8fYz0Lh78BkGeJzDj+Efv+/n
MSXSVdLA1aKENjGSW2HaK0nm/xvCUHTwZcKaiksxBb678NFgy4LvNl7MhAbAx8V+vGkmvk0DR58W
5VxM3O3QOLt6o6M2k+bbUbRwYjjEIWqUT1yjK5AlyTCSl73CzO71ARwCHFJwZTnQAcRhSgQIfv5w
BsRVL7RkwSO2/uksdPJpaA5RNy+/CfML0Y0bVWkD0TARuT1gKrULLTlhVMMfh+OZnxH5+Wjvx8/0
cY+CjeanKepDoRxf/fNCvVkRHQ0ApN8qoWN/WsVGXd5FImsjFV3IwJzz6IDjXTWf610iQG4YOGcy
6pKD8Sz+UzWDMT/1M2XvbP2S7AlmJbVq5Ik2UFKKgfRJ7JLhqvYPi3peEfeQecUKL8dKrwVPnBC0
nQb0JJK9BdiMC9m7fY6WMys+caaSHPgjToZ2JPsPkux6ZGehMhY75z7kgT11ERgystQiXl+Zm9Hj
25WeX5XDVz2oawj0fkIJtmMDZ01PVICFWtxp39rQhp57PcK0ZFhcqx4BpC53OQRnhP/ZC9zjsYuR
LcjBVIznGmJiP+ja3uZlvxtySeiNXrBbZUIiSJhnaZuaUVZjXLqatchtpuN86SsixnGkyPrJX+WF
ZYP1sE9nionwu9hY5o5AQVPM7qeGULq+9sl/EtHXlvYrZCpBTQEWq5CVsBbKfZbLO9io6p5YI8wm
+nMVUn7Ds3pSVaQ0WTXlTDDwl3szB0NZyLLlOlthIVXMiHl/K0bxzij+oaWSC8lQQ78rVlcg4jr1
0DTiEXaYmW+Swqdv4SZRdqh6qa587nd6Kxj8HGUhxozfY6Gv99Qu7CWnRaE7cdzNwjVmZuNJaeBK
5E0fcM8kSEwfiHliBPvIxYkL2ZdL5YShrHOmrvEVZGY79vqlex1ZW6TKV+GCfqQn4mlJqb6h/bhI
m/oLXPIcLqVAp708wwV8UV+QXaI0h7/T3sG2Fqnfkd/KzKyPHcb8xjOc/I0ZW3kDC4BFOsfuo133
QU+EvlnJX5IuQ7gA1TZ5txd1CxniJClSYWfRVvLm1QXiytv1u3UsIeCtKKmrFRi0RB5FjUaPNrhb
x2kYt5Dw+ygk7YZjq3R7RvC4GUwvODFpds8WWrw8ACUSRHrZkr7ukwGskkFYWHpA8O4a2C079cZf
YNwZ+2ED4qHPGbBhGlCmHofmOZvzS9RpTvuyv/RpqUrSUdDJpGU6/6rUJ6LkmBm40d88LtJ8I1Kp
HY23onubK5ohlHLUnAt4pjnuK4dH47969sQpsC5PpVslw9MPyRDzKLcJqbt8/yxQpCK7wXglyoBB
rB9296A+SKyOkkjRz9kLSfq5zqPG/fmn+2JsUqcNgqfYRW4P6PPtKcFJQvfDcPq3QX8gVUlos18y
WY9DjfC9wAbleNBalWCAw6qRPxR88Qunf+gLhzHrizLQnKANUGJRBDga48EkKcKes8ejF2p2/v95
VJ/8PciKruRy70Y1WgKYxowiJhWnr3IJZPhyO1GWtJPjxjnYQISjy1jslKvNt/q/2S+I/9Phn5PV
UbE1UYveQVS6ymrfZFrlB0t9rhsmCxD+jKjGdhCvTyDEtc6mfyyxKAfzg2JEzJwIwlQdLT4ZHP6Z
k55QFFzNhQd1k1IlNgBQNiA5cfKTYNA/l9bVDa68udP+eKAuaBAZjMmSyeIuYuNk031HM4awqxpX
l0Y1wuBHDFjE7C9l/5Gl7S6TWnZ3NMOj2apKOvcbt1Tj/EuMmeqwLFgGxR9HDAfj+8xxwiRKe86i
gNjmtSH3dyt35FCqGJ41fW7rbH0BRZZ+6DnW92vX7Jn+zGF8FqPeYXxaDXNW5Aq5Bj7X+iWdF4RL
jTSrJHXk9NuxmyrN/NRdDaxlXRkudWiyD0NprN65QAPPD2ArkFCwyo29fxqgLFOhNOvh+dviR264
W/9NNMWriCHQJaKVXEkbXLFAN/rtKKUMR5znRRZXyc0wJE7Uhwd91v2wOhVwl4QlU0mTFOZYijZc
Sx49q6g+PSgPxDIPiVIDf6qXnoSA+oFARLiWd9M54kFcAoDl5GB66N9dTI4J7VW42MatEXwJcY9C
/vjP3c02sSrybF2hGc+9nVhFR2n5u9SwOdVxaebeGy8I0+Fn1C/qrGUd20oS7ejvPgaXQyL1heF3
B+cG137dwPFD4V6qaJ0Xmy7mKP5OpPWl5zv/2FY0CWljoJ2GabsSABjLOgiAYFP09fkR9N6estrL
tSStQLUubzVi1mw059H6qvH3CQPif+il7sVwi/WTi/mSj8ti+cM9WN6PP5xIaEqDg+Oc1EB+iSl3
LR5Fy4jHutef2Ty6Zobfeaje4z+MtgA5zGVbk1A0viyP0mBUSh/68zU3g+RgPAsAiiiWPHo1VLvr
tJsSxQ7+oj1jVKhiO1aiEg7mhWcmX+feZuTTx0wWoGObLeieL9/oU/K0yJxdKG89ECz1J7rMOwhZ
RRP467QAbyr+9QmX2J1SgexjRr2NONmzOIgq1JQxto45idthyWSds7+o3CU5CVH2mYobrg4h8vWb
FuHkQdbEyaa0HPmENFEmQXGKAQp6+66EjDKaPQSAAL/mi+Aw1iCDxN/cj12TnJFaolV4cox2cF7O
tLY3eHiGsNOJvlUMyb5IVi3rnEj5JMjny3TqLmJdYlCdyPKwlUqMxbZ/l/LQSt3KrD47romAsuI6
EHmiuoIPs1bmwBpTfCuY+9mjmZGqVv9n5pmm5mzs6ZoevBbWH/3KHHXQzBxI/cHX1CzT5bfQ+9N1
v1zX/ATd4Icrm8251hmHskQqhHg8kscFgvgKM7dZiRVt9oHuYPY3h7eawDEOOvt8Xkt9A9cYDIBs
O1H4XSe959KFz6Hb+O1oMVggAwOkuyr4S/c7yTIh8toCER4QyGXovYtQFRyOAv4STvocvjrCy9zh
Y1b2AcmRl07IEUC19lqZI3Z8cuoNUSb4nRpJLOTljZCEJg6j31bnVQTGuSHl7Oyd8WD1igiZ4P0t
JeXQ9Tp2my3HOeTik+HjFrcUNSHDMkRnlPqBoS4IIfaHUsOX0STXTeCBdu26BU7NRo5Rai1C2qa1
Zu/8szXeeFiZwOGX2946Bbsk9ntXCqkbVIKonB1SAXATbVjDAS5cAgJIaLrwlOZ7SzTh0JRUZ/nY
qA2AqLtbdCDxExn4LZe1G/4Of2Ix/XDIn3AvTY7WwlP2LCGFiR9wKPg8A+eX30dLeXpbwcIkW3iK
xGVfKy43y3ZcZk90TqJI6JVMoJj63TKDP0KsjbZaH63KPdytLKG71yYSm/su1u4JQfR87WWlOMvu
9N/iXUQRyl+bR9QEsG27tayVkIKLLjuVPXfhT5xlsh1GZp9+vJp3MdLadFiMfJk2wPkREt2nCxAh
9r82Z488QGSlW4v5iiWHOkb5Hapl0SffEPL3Jy+cbUoNtd7Sf5eC8u/wGKSGE/sCDKAlTWJw/3+M
JmFlFcniaq+WpIaB1niHKVdBXJuCvoH9yKUfMPdLUp4+JR74PSrC8KfdG8K2lPZ8buuWMxMvKHzE
eS2SZH4+OUsti38zjGZlfCIzFEptLS2YYLgv0sLOdriQW0t/3TFeBlZB26tPRmMHM3JPWnU+ac4H
jcTI3gNpmPFayq9mlEU4QhjKXV29FBMUF9cl6bFpeP6LB/cFLLLua3mi3AMR0Lyv/cS8lbI0hojZ
SVHJb1qnee4edUqks19PwrCWgnybJt2MywR1Y8I9u6Nm/SXRCehBBUOHK/p1qsVYJZZUNK+XT19J
qTbtockb3jvsBF4tayfxyXs5Coqf5LH6jnp4c/e5VqB3LqodlZm1f0Ps5WJM/I3yzzprxOIouOc1
9hLPv7I0mWwiw/Dm9Imtcm8Zbq0Hd7rACQxD5Y9CFYOTImDXqbbLgAfjb22+Ra+9HaKWAvcmm/AM
k1EYj9yWRXDoDo9RQCfYWLuJpnRFj7oOpQttmIaeOVdkYdv32v40nycrGjPRu3XeJdn8wOHPLDdr
kXg+VD3gSPIdHwcNHDJE2fIyXaufT6v/NAw8gRrjxGEMvSPBI3Tw/SWVkzGqKFxQ4rihXTIs60h6
2lCj68C1R3Rmjn13XkuULMcBeyDZPRPhLxq20/qEOn9mfwe5UEkI1UpEO4D4aBSLDwECz5NFM+6v
e/PsXXajBuXddB/WMTx8nyL0mOvS2Q4enwKcdFuIUVhrIbOFEavKKGiTfgow8l7+SXWA5E8ZBp7i
k/E3SVMXzolzwyvTZm2iu4EXdcScVyP0XdHuPs4SlUqsfIjlZV09+VCzdaaR7x+jISATdodtHBjO
xIikr0sVOXxvg/D6zjET2xDtwUvpyDwLazJAHtbXQMQag0D3G/AKu5GYsFrLf7Ut3mmyqfqdQehQ
7H03QS/WwemWQ5g5uhVXITOcuJoMIY+44WxkDCGNiCYXoE9KlQ49APQnUioPHiXp4lJ/EFHFTdBb
hqBFpBCoj5/j7k2E3sRvr3p/E/fQJllQgumaybEiKEoUrDib94xHCsRazk+sUZNHz+a1HVSLzKF6
72F1HYK3BzvD66t3EtsfnE0LmQ4/QhB8girnlHYNBfUuqUxiXEATG1Kaz45OdHKi9Ij/e4+VBrDb
6f/xUol3Qv2I7jRvZuLReYHPcd9bnw9gwf/XL5mYOrO2Xx5pJNBszOBJkIG1jeONCYPGH4bs0iX2
VmBhriSWPaJV4waiSF1xxlB7zpsOZOAz5bkMvKdvAHmFKXBkBjBU0B8b0e5TWj7XOHTocqLR+oZc
pIDMhaf0rvJmn8SKFl5g/iI33St+zqxAtstBPf9s7GMOoufw5RC0VncGHddmTpa/k9G9Baa9RQRl
w/UT4Bxfc+I+v6aW+zz5ZpddfRsnfSr9Rzkj13sXM+69yC0wmtiJcQVpluw2/tk61TML8lbKPoYK
EkHmPUiv67icAZvUnu1W9mCVYPESOWNLZCKfTn3CuY2jSzsYR2XtxtgMyArQPHt3ck+rs/mzIg9R
DgJXOp2IcTSAAfFWUFaCllTS6JVr+VoIxxTeSA7aYMaaAPIfkASj0o9X/9GGlcEce3cIec+YQlEH
XaFJE41UWtOj2mFNjbdaUkjkeUR/LFUr66mRzPQ/uyFt81R8EtIIN/bcIZ3RjnE0i2Hwki2PFWao
m3aiwK6szji8gVcyLiNIvoX3AhZ6lrytyXlaXy2LjkCxgIeil0ew9x+vDn4v0Guim9V3Bq2QNSim
p/RCqYskRFsr5aOkbbKWgmSmBcWYhNe1xijbYEaNIDfhZP9VvHb9svKISMAK+I8ciULIXo8IIcKn
9CIeefY9w1oHQqdK+qpL+MemqXNPskJPKytwKrthzrtEV9dHHWoph5djjZyj+WHIZFU5vHJdF7F1
vpgbdKjOJ/Ob+xbEEel/ffqCC3Wby4L+TtOSD8bTYWOcyZAQ0kgQxKpcDZGaLo7DyDwUoDIsGAIB
/dUWuVZMgjmHUW/yolix0nTQJpkKxcHPDKtg08tvJEAnjeSHH3S1Tp3w/xK65DUJ/dqdqs3cr16L
fKQeUeSz9nq60agFe3V9i1Z391QeT+Ega17CS6XFG75+Z+RxJItMR9iyuBqAGjNnVbQ/1Bw/yEZA
PURRhaJBdVqregSLq6j2jlxgnzyOAfiEfzxcHRKc9X3kxdxGyWaRm4P6Lj6hxg0nQCHa7uGKeSJz
9NDrQs8Otj67z/2EQgPc4gvg8j5eYEZJH9/oVnUvaGk90suKgYYavpLAuFj1x9X4/jUoQ040l2TH
ex5J9R34WHGb2Jl4/vmCsHydm5OFkoOF6i68OZ5ZQbraTPK34rWtohaL5imMYwdKxumDfIS8aULF
JtDuRu5J7PoEuz0YsYSMmMr5mXwX9g6Bq/HOf3JWxHY19S1qGw6UOhwym/P0MKFETXKeShf0mwJA
5USg+SM6/6v8RWXDzze/aEcodOVdRJ9/L6yFwigT8OXnLI6aEWLnbwxh/1ZTPiK3SvvePKBDKAmZ
tJuFX/Ju97yB3HCnF1huDwMfMjoR4tDJTXADeXvkMasPdMRmJIkvSgPdVsOfKozkWwWuuxu/1ba+
d2DWMW/QrWvXCjnivLvxDiNvpQ8nbhRzOX5rQLZrqCW0D7ZJ2nNtaaaR4CE3nLxFuA6gM3QdYW1x
3oHHdqg4AafO4LLKj+ANFn2tV/MitgAPZRVuJ9bNfdXmmmzL6pZDsKANjoqxVEVGXevapNBlJehr
DXdlXMzR7ZMjjQ9aKb1poZZZI+RWqLwFbeNaoeZW8/DXJJLOIX5bt0QjCj97msOFxNgoMjcobllz
JzIBSfkIIhJ4TZXInHZb8OclKzlZKZQN4fY3Zb+J6RlHWDGR0aPVPgap3wUxZkN2S/YRtdFP5Ct/
vK55XCcr31yZ95BwgiFLQf4cy0iJSsFZ3O1w07ez7IKBm7a1joCQSrA0SJPshgvHf1REQL9LUqDs
L4qMa7ypNPGQ11Nw//i6GIO/J0tYQSwdSOVxovoZVEAemt/w86YiK6LmVZXjV4G2/NeimvlmBwI7
HFf3q74RqQj+mk55/s4t3/L6UnGCi9Lv/Jf71RKTW6s7wy8GlynLfmVWXzfMPugeVWdW7pKKvFmS
x1XGz+9fNouGIwmSNL5ecTqdyedVE3x8rJQ6tqOqUlKulF2NyLT1wkORiAT52C/zIjkwsCavchqc
KOch1/Al4ZjW7fyX+pzeh6iXDK4I+EgWDMjHQtB0t1t6TC/f8qsuyF1ZNwecRWbN8XZVmaIpp04D
y7FRFHCl9/97AvhdxvWjmBS05I2qw3LQWSfj4n2aQhKJJYdpdoxAXMtPDga6FlqBq2LAfdd8s2nH
885lblMnwxaOrk7zs6Bu1x9lbmTDG3ffXC6hDJSrga/kQl+XDHpzQN90aMFfYGzmCL0Uj/eogNb4
6Dsc9lZOIXHxnFmXm8/tFRkMpEEV7xS8sJVlmDfwr0cm7GnYwVG6xdx7KLtWNFsELrdb3XET64Cw
jjPmrCza1ESJtgyu5sThQuQZDsM8UFOq64clAsrOUwDpuzWXEgVsnBjijMfBFgF0F9YVlYKCBZqP
w5KPAh1ADzOOdQI/DXJ7gICKiAeCLGUBwd4+UcUvDGHyuTbyMhP0ilAudL9b1KLQMkFPx3w7A2Al
U9LkgD8mYMTGEFPCjUEPBvem0YHaw3VEAWEDrH19wbcDHMMolKFpG2MMmLjUAsMjRVFBdgo7wRqg
iMKto0vytAHKOgAQwmsEO061G4CwQRuuPL2574nNCQaBCyAlOGhQUZfwAdYeZx+vcbO+BXKwjBFS
0JRUfQwbGcdS61n6b+lujLf0sxT5uyYRuJxf+n/5ElLVGVx8kSZ9XpXp/g6aOc11w6CNL7xCtj8M
C3pADIDtH1HhyKfSmwyvI4Qaz3XEKSYlpTcpFFfWhX6SgvSqnNWJRMuCrMWGs/aRdW6ECJ6KHhz1
vCvOnNmsjlZJdT8H7h1Loyu5Y5FjZIWAzVAqdxZXV5c+ObFPh1lmJ4zzAlCWs2eyNF4jx073hIfi
MW8SfQxr0QnJuXtoC+aW260Cth0YgkfBJYLprD7Xgftaeh1UZIHBJSsp/1vsPQvi8f5ciV93aUGp
quO2WsuHOTWc5qClOLIinnZR8jNxysVTCGRDjgyTlzAoYohRIvxegEXQ1hmJCFCiGC8LMOcmqnBg
TJNv1Pk9VPeqSgC4R40C3Uk4q8hUH7Ia67+8ZfdGmG5TCWnULr4DCzqZWXIldJMFgXBOys0OHSgz
1ryqRqeJG9jTBXavaWj4rU+7EUrBhVGKDe8KW5rwwxb0fhcJY1RIzzu4Tl94tAInKgLUb9wzIacQ
8wiDbBc8gIAm695ajC13WapJn0JWeBYrOM2cIYQ3125hEUkdygq77f1CyzE7SMNTvKsJWWluqiek
mZJTcAYNer0wlgtpDWPeobqhSzPJrqWTHCJqvM+LnQiARwL9O/kPelE5LSY/cnh3yW7o12h/CKzI
UWb1FbEl8E4cA/BhLvq12WX1FHk8oF2emxIKzulQYKkjwExZq2H23dcj/uJUdOz/XyI+64p2sSvC
LRh/uxLW9DAonhzW2zmplgAyNzkshutGnxcy8036HL6rgtkfHjz3g/U5eyPDyc2UgtkgDGSJJAVa
fcaK1vhmHkZnHascZFsZjcsa5lrw6+k2W884jXsR1AT/GtcSClU+b38Rb/G9d4KqAPznPF9u4Ztr
DTyiVWApW/o6EEMMtvrR4e1qnMpPcBDBD5xE0ssV8ZAw7yRz9tbphFez1u+8ybqFr06Cv481TAzS
K4mRLJTFbqKM452TGrkEuc6T2Birzox2Ul79kxzK2T2VpNIIgidJPkofs/6/kwAchC4dEwkbbAnO
POrHRKFsXYG8dWUcf9Ft8skDetdRts4MOD2gLDZqBziuV7fgEHeK+J1jbqH5kb3umy+I5rQOB+4J
BeE6TB8cwCo0G/OeGlaA9qV834Ef/A7ks16NEFf1oiYiwezmgBHKUrvq9FE6wxLW5I7UIwLNB4sU
hSCFdV1q3PcAfM21lgG+JxkWrndQSg6LiIS2SLqK7QALprs+jC3HmbxMgfdIZ9NKSa9cMNmZhF8b
mweocPNFKjxkrOcsPsAuui3q8Fztonc6c41FX+4q8yWPBlXpGqkhOFd8LO87ECyAav0NFvLBF4n3
VXmHvEgs/itCSFFz+D8RYWRbAM0IgiK6v0Z/4UjjEu2bE+oD5Lq9XjWEHN0Oi3FOcU/V+w+JOfgU
G2s515/fw8lan2Nmt0cULf0CycwuVrdotBONB0vRsBxYfYMENJbB0YBBcQY4SFBw5/BoqYsdkNNg
UDYDj+ggO7984aO2un2C2MNM1eQU5yTZ9UZygWrkPI6H8XYnBYZljWwXDEnLmZ/aT+i1Sj2Rmkki
/S2sNex/CsXFPbkuvCMRfurhJi7b0YI6glX+WaiuGkk9BoDPGcLGbAfVuV0B7KJrM0wZhNz8+YLd
OnbmcHs2Vc34UiMyKW2L3K5Hssw/Vm3Hb/bhgk61KAVzRuLx/M8XYzJuRVLeRbgEGYJWApzpLuCu
yY47H2lMVK9yhSihTP9Wv5W6QgJDLdZ70Dl/kdkCML3lVdCkuAp4ZCx7gvRg2fnXMvQpPM7qMR2c
Ij+lXHmXS1FOpx9Et3gKHDSmDqrtyf+5GDaAKglh4o+pWpJ4a/5CgWPIpqcFmM4IC1VzUt8lauXu
92CtjNTcdtoFaaVMQxqyxpuOzxYcz5aPO4cI0MqbbAUS/JXgaIg//qjQZSJfabWyAUd5jrlRYW6r
anOg/EjdsBHw1KKzQsCwwBrfRCsPAgIXYOCIaURPO5yInU14spnmwJ54ZkraV5JJqgXyMWGGNtKk
pyRYhrWWgr9ug3KdSBI0QSGdoZ5OmVeJMjMhjkoKIxvHl3vWIffZBH1ISmKWga9C6YKdPBwoSo9z
mMLniqyW+lNyue+wx1oOTogTjm30MnvyEP63JEKWvyWzkBOhHoxCli7YhHj/oeQyT0jKb0jt7JoZ
/0oWg/ttC+LTYaHAsj2/caBrvM1QtTlWo3V1qUw0LvX7NgMz9jiXorXGunEA3iLvP+6UN4DEgBC/
5pGSsmfXE7bpvZkdBqkd9SAA2fimJKEEMHeETPTaUupnIWXnbKlG3qCQUCxOpfO35si9ybohnag4
oUkc3ysXqLiCEy5Pmqv6NQIWBSfKR8lqG+C5+KUdFT4oTBivVjUpxQgDy8G3FkegXfo2CAXvY7Xr
Ni/OgM2A44TCGkvCr1vedH7PCrJS2ajF4rts9rOfkFLsPiIlvEPecpOraRcwVd8MKChRPcFXhsa7
n9q/IWxVZQ6xuEUagJJp95V24ZdJkI98HuRoKo4KJoXmKu9ySm9N7n64WeIsR4BijLPivEvrkoTp
OBjAXbTqhlJ0jzfz8vrYwN8jSfmGSf9sR22ttE3F7cry8vGhxEKSOu24DaCt1QpnZZGnaVSCAUg6
4Vqx2oHxArBzyN/XfDptSN73nV0E4RkPNSyJ6g1NXINPYrYOWlNYRODGaaOU6QPGfLIiWHsegmT8
WvpWcVvgsgBwEwSX+N7z2lcGTmjOXXxN8noNVuXQJG/HNZsZQSz4hm/9OFIBWOhsQhrySnhQDVnj
ev9qROkaRdRZ5TmcG5fAw7MBpiDaRyIrmd+KUBfSfeZxCtSYOXHsG5aw7SCGCzdBRCvIPpJZTb6v
SS2g+7FcazptUxx8CzYYzDfpy7gPTDfkeRt/Y4oeoJGe8w8dnNzYnmCxxUXzZTrMbuXnhKP0JZ4l
dd95dyab6RV9e7YVcC9Hlz9nVbSnOcLHszaruTryigIKfZgIUkkeCdeR23C7sdK7bqTl29Eg4kJn
d5XmzagBqxQ5jYwcqFX0hId7h6fXpH3DTvJmaf5pdaxvmPn50r5QFO5KYskMFPKwyN8QKhXWaly4
DfosvwuYXw73WS0shU5MzrjeiZxhLBnypLKfFMJpwfIbYU5WJka4C01BeIvjRm4JNIiFpIoBtOj3
WrbhTWIYmb701A0FMw4LDUC0D/BYDptN0sVWmGT8/DbBYIy0Rk8KXqWhxgBcGLvZxwLWsBi+b3xJ
/+ANwXGSktZiA3s0Vkhvoxjewb8e/+iGvVyPfkdD1jI8iHrOqwBaPet8QHnY1NpAh6gwHheddFNC
qVwlHlTWXkDwwB7QSg+4YW/UXFIzUhOEmN0vXwOLsZHmRtfa6MePMSbzwIMC/1mI0BYP4juf7u+e
GMuJItxfUXkAvQHxkYzo645RXV5CVZY6W1mHuP0BKaMZehBxdUQT7mqi3vInfm+oddULLS1pTvIO
L2WeWkpQuPT4Nt02pp0ZEN9JcAo2eAzKj8K+w/1HoUsrl134h4jjWZBwwDvtkPkePvKMUZzXf9pl
KZW3u4jB6Fly3WIaNUreNtN3fxcyH5Fa3np88b/azbZtNYCCstPc4/uiiaxWrKy173PMJ91wUdSl
6jWJyBamcDm12wxGI1NivmuX5o333X08m2fx8kezHPavZa0lhexSQDX97sCYUgs4ifUKOsVZoXyW
L5S7Nr73NHU6jMCyqUp4wD1knT2PlKd0YDDjrAsSPZeM8RU9Xpty+WQI69XQRhgPFwMNSyMNewW2
2cY22nv7ScSGLpd2ANT1k/UsJk/DUMN8Q2H9LqibZbTdLNz5Va6qNRwtC7emURHQdeatKJ7NWzAO
wHWuVvws8wn0yQfgk1pVsPskq9AkVPHFh/zZXb4awdEr0HPz/CuyxBk9D3qWuOGgtdvSkRBMgmSP
bH2ZNavO5c398jznyfhJBpIZCF4RFRtTqeR8I24dAkqdcqWAr3WRVI52MZhD+1JgB64GX0glBk/3
9aY4CFmTlV8MORItUgpkow6tbHNu90be+f7sTp2sxMDKm/J9XZI0bnJ9vTdL23qdtHdqDGBtVJTQ
nakyw23+qw5PYYqav0YGfvt64vNxGrYLOc+Rffi4+VG6nQt7fyTLE4pe06gU2TVczBluYTSVNY2a
bxdi1cADWwjCyBZND5jrJQl1B6vlZ0dQFyE/Rnz1W0Yb9ifczhuXlg5OnE0mDgtpQeWQ6iocQIoq
jvBh9qljW1k+D2aAh5KshqmEU0BiVjZeaeN3oHdZMvpGVbJ4YOVdvkAWwC80ErEyGNQTz1EH3RLv
Wn6R+ODiZfDDp9cbr0DwoD3mToLtVlouJexpoMNpJMzkGyYpKYgkN/WZ6VhE1grrXpmnnxPqVTpD
WWBy+XusNpW1k4nnlu2M7A/oO+G8Y5oTeBSN3jSIQprTMXVEg0ikGHwwIhuXExyn/c9O1SKI2KR3
drjev03CIQV0YstVrKnOc9Esg27e/OR1u+rmvSkOrfQzcdLUgh6I29QfLDKMGUM/uvz7Z3yIKTs0
UA+fA+5X9Sn4JV9TZZFLs5bSwlMcYTkspG5KLed6CYmneCEN0b3baDu1nqZznWfw4mrpfoXmuHSi
WlAjWogweMulSMbnq+4fHpANeogDo4NpT6BEZDrJE9iFClcozFtWr8wU2lwqSzbKcKNeNzrkwuA7
+QtqYJcUiBjfsfYL+CJiMIyudx84QW0M98LaJ3P6n/lLCcWdDoEnEiK2L8WlO2vFV0ARVOar7Ndp
jRs6jaPF7JoZkfloHICwdNWeal8Mvx26IGhlRon++ODMyBeNMpjANkwsGKqhLmE/okfyipYvO29H
TivEa9rDDLaofEQsHYCTLqaKPXH52HUVD3NUfyhKHHvq3xBgGcv5QglraWK0/ENvEGA6m2aDIDxb
ZN2zGevZMpAFQ1vJWZnet192+xvcIC0whIQgw7etSv6tPhCL7QdQBbDrw9w46u8CUzBFwBGBKRav
G7JRwXjjPAPq1NoCe/D/m0l77vvyS2JLzbTQwIgdxYhHg30xbeJWgt+OIJQFTyQp+/jQs70jH7Nv
t4LlHkbM+NENTXV5XTyC3fzE6X/tLTBv9eaR81XIrjNg7TiYi1OlHFp+ERAl92j6achx2y9lfHQF
QWsdpAfJ6C2ZkpBkb5ijLXR54B98yv2KYafg0jGaC4lNet3VAGbtmz56oHTMOHFVgqqZ/IU62wMD
4pZT6lkJrMygIR1b/BrroVT1Z4IRaV7jOlGDjCWH6+onxrYg6YiJyUVRqV2yOPCsG8xlv5ZWZ8CW
+aCHwFtbFknhzdBMckZtHysmfOD3uF8wC6uKx8rzak/wGN28lZx0l92PvpYygZB+J8SiTseObcwb
LchzcIGtK2Z8OR+/frPgILaqz6nShgM5bneiaVgmj0o6CXub0w4FVPaj8ct/19KPmyAiFoQmTWWf
IGMxkOahEMjAIzFNf+hmFaoNrUiCnh4baG822XmTPb3NiTozwd7maPCs7dk0RmvxEUtV5cY91kQv
0gjdoFrNF55/hKqTdKBZ1P33OqFvuljVNJMTz/og2Ld1RiL9cBsd9pIex6+i3F82d8QhtQsTDAsh
h0Dh+l/reIMALc3YRkMhYHtxr0mCP29YUhjdIAa31Flh+k+lLnXGYIbdt7ZOc+iXXRkjivSMjrq4
x3iPhbuRzdGftkHHtreWVO8Msszz4/IXBwpu3CwdLc+9l0lO/6K5Hmd59Yp5n++a3mEdg02dSvWt
IxVc5DlgbbFAD7G7r65VZH6AIdPWiYApeQ7joJ7akY6WgS5E+k/VkLon4PiTABl5vqX3QjdYHI0T
JeJq3PjNOBfNNcJuo29jPjCcwcMZ4Mpgw6ambBwlxeUJrrGl4rqPEI9qvwfeYfnANm6NEmtxZibr
XQZV3o11a+EzqAxXnO8U1dJABG2yhQTe/t61eVlj23TVDgWGH52XD/OjmszNgvzUhahoVgwKFL3v
GRej9wt5XjAI5o6tfeggxLGqg4ogjhl0FnpeFXxSiIh0snyTMDT1b3XM8gotpV043+6cAWujvuJO
DhqlHINw98TKuG9ijdoahtDxQmECccjX6HtP7+I9ZceLEA9JMHR/v3T7rR14thA685ouaqhPCYdI
THEWyMKlv3oz7IjvgrbAvrSFLYgBXL88xsgJVWYzvbDOr0z3nhY4m08d8HCQjf6sXEoA55RhX05N
+BaMGfCg1MWstQs9Ivk/ShPidyWw7buf63eApqC+4bfMUYBQpSaWuhhOBUjdICnCWjXv/lFUjtEb
QxvR0Wz7HfILTro7X9/SNMgfiNOmTgYqBsQx6qasTlPYL6ZZxWcc3F3roDamWHfC1qcFqwZJXLUb
lwmE4F07KrMkEshpkpKKlVsy/fL0+wFsbByBbA+w6KL/+1mdtoPsLXzYWXt6aUE4/L/kotq5zWwX
9vDc0bnyxOZxRuJk1f8aUkO9/E6LnOg0dZFEIYi0jhvVzddONGlBqJJMwhant8qjL0e1C+T8LaH3
tNHBd3/zhcQYAuZdoGtJsqMUx4hCXekz7mtVupV5YDwMk4Nfj3hgL2R8AJUP8/CtqflUIbsRUVAK
pJmOm6fwKBI5CUm3jyBjv6J2KAj4QyBXGZBYXaLG/CBGzy0Hb0OftDSmlMg3fHkIL4Ox5PtEi3yI
cWw/3Wr8PdCw2TQ/g97ESE+a+HmfWiqPINrydSQRDg/kbBfEnoYvcvbnMvki2ylhyEX8zkfvXv5W
pM2ijjDZexzCQz8EVeMHIPHoV+VVxsnjXomCEqBN0Gal7UNFzqf52fHiXsutA5xxrrbfDCzC2ZLl
EgEeA1uLAjnBaJT+x9FE2pNOQrrPNk3PVt7bSX4QiEJymttA38nO3S0NSoqAE3fPm8Uejys+j+IQ
ip8QFhkQkgAVoRgdsV1iPGqSVrnCTXr8Dvwokq1sbZ8la23RxtdY4vXkH+q3fmFwy7gPY/XjOQ/V
Zx0MjLCIBdd79jNeJ1GDMqN9UhfvSTrlI6Rgg8Sv17lSJUYXtjmDHWs8t6RlGp/anCuxWx//2sjS
CBxuvrpskVvHsxg4cuhrZKlVUkXY45tfiKMtBiuHxm14H4SzCreTVSw3vspv2WTh7FNnyinEOTyN
FjROiHtv6iurGxphlspLyszFbxCJE9zJTAKLb5PqgYm9rWfclI0oUKcHFB2ENMH+Gusn20rThR4N
6BHQwq5yxxI4HJsrVUEu4CT3ekidcmkmy2lnFlTqnhDbnmwdNSVrS8ePpm68IrzF8sIoFbbT1C5l
lZV7gh63vAe+wpZabkG1pFGLvST+kYPxoQhbfXMvztFdKKLK41iQ7Wq8On+Qk5CimqiK430SJ8Cc
dc8vW6ZU8Az5an3G3Hq1RDbglti1b6MJqJgqk1I2cu4HFSctQbMGPrwztn3LHM3/deUtSdg0rfI1
YphRRaFMfN1IsYrPVhklsKjPiO29KV4gc+sKqHr1A6+qMnJ0X9pdSdcamrQFIMkduVWATx4ihK7R
OHkaWGkWUupl+Aekz+v6RQvblV88tr1px2I1HjOCGKA85TlpOj7xjsTKDNWiBVRVzpShJu7oV7Yy
BcxBmRPaNA+4q5jm6uUld0eK2fYlitVJs+UnSlYGenA4f5ZXH9/jgn9Z+/cLZTBn2Xifsrf/o6YI
EoDtXLh+y2kwWXNUxBK7sqAEPXTNKckb7pWzweYii+FWBWBXYMZMuX649lJdDe5k9J0nbGdeHAXu
fH/f1EOiTQ2gNsXLhG6yR23bRZ3Sduy/+RWl85a9ePYlsJsZCYn8kbCEhNAOUq6wXCJf9odfQ1b7
c6Ex6Vo1nVi3cofFg6LRd2X0BbGK71O6ECWzHLutGMhzWz6BOipnPJPxI002Jm+9QI31N3K52DsS
AkGLkxrgorQhRc4w0yImC4UQ3fmBu+gi+VflPjlp+uso7mBndSC/szdTztQFemzY6nAmVpnfHipG
2AFEjcw6O+h3lJ572qWh7JgXEGLY3bO1VRPVPeZujsgeeJ/fLV95mnwVXTLmTijTGZUchBXOr6dy
4IRt10jGDODyySjTGky2NwgsA+sQNCznL5LEX1k9ae5MSPw3VLJp8uI4/TKNzon7CZYOBdqaT9SK
oii+ws8NXYrdZh57T3zJEhv9F4/vgXFsz4oeTb+sjvBsaB9+KQVdapDk5JlpY29qyeFTq2F5b7C+
zDOUpKbqwE0B5pwBN+gHJ6nckXMtl0vEimmV1TG+Rm7gXe3Z5Uu6vRT+aVImbwl94leBcfyWqZp5
dnUATtvuhok2GhWQJ/JJUQQX1VhVUsO+xkOMjNry7qW2WH4pqR6ORnbmYMNrEhwmZIA8tgyJ3Sps
J2Pyw+JkBlcqFD855oiR/0343NM93IIUA9wVPFJLnBc54oDpf7UoLhnO9OrO+GzyMrtH5y0ciNoH
ZnRr0Og7IvAlxkCh2VmYAQUYBTMSRAowL0wq4XHmkHcS2H8I0HOxqkCn9dHUw7Z4Qeuv56VRSsYK
IFYbCi1T69MFzNMQGiHus6KK7w2BgQH7vrpisN9NUKCs3EpeVgJz5uTeHuRrInoJG95p2KJ1Vans
vVMWrvZq41CyVuRykskXQqc4PGBTxk4xRdDiYakAHvnDoHo7QH7AQJDCyRsu0OieE0uvgo0evzBF
U/DWcBTiiBg4DP0tupqRP1uSq0qRfUUMOVfbMEcBHzoFhRhT37JBcgL56roM/AryKA/TYXV8ArGM
yfswPLNaHHjrzvUQQYuabKjhi6NR6aseFK0M6cz1IWZuc8C23+38HKNNg0bJ7S+c215Yi2cKHgNJ
5efaJjBgC2Jwz5v3wcVMDnpgtA3/eJFF4R3pi4VaWwoUK9GkTUACQJGxzBPqQbhxE1LRBUO/8sPn
qX3sCZsEQ2C8bL28d/Pilzf3Fbhwjq7q6dD4EnXa63BwPmXnXzZpM83r/b12SFo6BEORsYF9q/8n
haKulR1RcFX7JeGeWs6nqcWZOQP6UxI1W7MtZbdhPtXhAWRUXhsF/OFwBYlZUz67Mvig/mZuWzxK
Syzq2tCMpbLn1C3kKwBNaFQLYldsvsV7P5ScycyDnRAC/Sq0V+TodyLQqE3OHCaXZhHLxO9yCoad
qyb6RtYO/4tsSwV0aoIqCDiQZSp8Nq7G3DyD92GA2FCS7SLEdhbDyQvmaDYTnq2odhuqMxw7MVHF
xipnA91zKhuAYYMd5H5rrwQ6boEE3k6D1+3FR5JESxwyeB6SOiOmBLmFGmxxT4Ib+DdUeKxVR+dm
i98mnvGTtGCs7tne+X48PyHbUV+i4gvQ3CezopsfrT++f7UZKoc9yzywU9OGZPKuV7rDqXeJS4sq
OeBIAYHzIGgXPE2rV9hvm34MVPMGFmXWI07zIwwM+ILj5BCGkCUkHqlYxGv2hCkTdGN35cfYHgSN
/yWjKZjTCoZ0LWnWlrAUqyczWepxaWtQyd3/qFMDFmxrQCiVAR1XvocQwhhfwUb1arB93Ysa4ttF
8IrVPRXvBO4l+Z+8hvk91L7omXHBruyMV/m8C4HSUhoLqX8qFllaGEbeX4cAEzbRw1xuLi/sCSJL
XKFkm77ygtp7P/dK+RocsSl1q2TZPbityUHG/FgvjLH0D7l0knT8oxO7Ec1+mZyU2OZcodwBLXJ9
z1Bvk1dqzmnZMV/DtqW4gIoF3souHRmepANA6OuS6qxAetsm5gcYQvTDhA5acQf52P4cnI9uY5qH
07SsrMjtQq6RJKGXx2NMjABvXOQ6M2pHjto9UIXa3X/WsoE/qx9XE6FeED4sIssXd/O3RsWTuz/L
AemJvbq9yG2tiAP1R7wNZMFuXM91TJ/9Jwpv7ZP3K1mTOez02tFdp/o1/8+o3pF8Smnv9+6F1S7R
qpo7y5v0qaLgBGgbcBp2yff4kHeRakF7XmXGm/3n6omNPjNML/73nceAtmlRhOnMj9DkB7YWvP0I
i3MB7RyVvFkHZe3dq6lnXq1+HYk14OqZ3RIntJboFilwrpZA3C1UEnU1iBwUWpwOlw1h5O8n927O
8sNh2365AkXixaZfhmCwzvNsDwktxe9Abhe8RM4X1rSx2dblMkpvc3IUeRsCdSR8q2RWk/nmeIMT
yCjEPoDNOw77ak7zisauSX4c6bRWdmaXlGxjkYQOvAlDCzM7OjaJZ2/nCgvnqlP4c9xOfeA0361N
A1yZ7ezmHRFoTGHSoOhOT8fOVTlDUrCEc6Y5l+ElPbJjYY1g8XS95p7mvWHBEJW7YGjhSFYXJi8e
oxe9cF/HMD+I5/doHi1ljC1Tz3Fp+/eJUI/Otv5IZPGjt9NmmdDwihjmYj0RRjQruddQV4Xro4D3
pBQ05dnlfBeXeZq/eZ9UlaVWlwY1r2tmvEst8bSgkEk+ocw3JBKNK4nfzn0ljN3uaxXvUB32AAwF
rkRYju8VGTts42RtJ2/ycbF+GkZ0bfEybsosqM4QoJzjTjh7n0SpcYxgqGfzVJkh2MpffHbibsEh
rYjGa/NAKpvWuCtxrekstHQaQGttznVd2xRPMxABwinyhBkl55DGYMMtfYczJTw/xeJJGTi5rEPt
8O3MGxmj7E5J5kYF/O0PS4HNsLLpeQn5+/EG93Obi4Ug6DBvUXt1mO+cR42q6/wcpD3ALEiAhtNp
mASQmOPWYS5MAraYSCioQPIjZlPye1JRXYy8MgPWS7IpbCI8uRRrv8npuPbkzwvY2T2ZkjhjO7Bl
9ZVOD4X/2QNP+uWlB6PdUiVjk0+y8Y9w1GjwHzWjykM8cspBuOE91L8qumIrkibBwrCjGjguL3aH
iJZ/nvJlxl27BO5U9uGoY0hwSgMKYyIRxmu9BV/Zpr4CQ3jjRshY+H2ADB4Qf54Wc/+se6J3e1vA
ejj+0A/IwwR1Fp3RjlMw8edCTvCcvdmOESajCGZfnanSVtjueTYdVmvMA3/5kotsP+XEAavkX9Bu
XsouAKRIG+CRufgWejX/wuiUSUSVXmp9mW4S9h9Zz6aOgdIP65lmJ8Ev4lBWqBF6aDV1TuUTJRga
40mxBX3AzsLVQmklo/ucRAY6KXyxMyJz07azMpfd4ORtsg4MW6k8CzCoY3QfZBReLqIgq+hBdbl3
CBd2TIeKpnXOl3ln5zdWB/h1Z5XrvIlyNAnCcdkPe9PQaeZxI4lPBGPb/KmDDv34M9pVBwEK6NLe
BePWhfN9BmpZyPmGGRzwDtgw1VLxd8vl5uAfv0tPnFdE79PoVLdxNcN/drziAGRuW/JFs4QIN9B7
VQjzXGUtUqpUpPSEBk2ped0m+owyD6Q7Y1aYP9CVlW0mYQ4g7/6pmCL3voRqn1FFbBcOaejNvRvZ
vLZuqilODq8irsXIvfNXPa8URqNiG58Xv/1tU//sE5QVb96OAt0S2m8/GiRgg+iwR7XrP4IxArLJ
jHZeO2LI4FAMpjDg6gQXHY2upRJVTKSVKNoj/69st/7yaNEBD8Iq4ZsIYLpL5oTZ3PyajhRuGXb2
qvCdv61SYzix44HZUiRNHdEG7ubLjbrTWymGjMmW3gn6IU+EK43a/FhFYlt07gIIvw1bdnGnXaI3
2gan3Kozjp+eydBtBR/6IxzmLJ74dJsS4qw69gneUrmISPFRb3hqiAwgol0z3ss3Z3GbUqe4V+KI
TSSV5fKC7Nzknp51iFsVhkHQq5lLPkFTakDo1t4StJx1CEutoYjkpBZSjaevpWx09mBwc+4o1VNe
XhOtBlBLEStQiaRPpXkdmcDzBGLJMRInMmrhpVZc4SIlnTtZbr4GUsjU/dpqPd20Txc23iI+Ner1
q1AsQIRrCIhW5owMYjvWyMBj6jX/4kaL+woHZzTG52A5jIqqL/l/Jph8q+cd4hHVNVWzNbAkVghR
imjAI55C67NBv6YbkLDOQnFxTtwuFrml9hUGDgmvLBmFyuucBYWok/1JigJaJNVBZa7AorPiWvSS
R4EGa7732mT32PP7DJd3YQCnGwlmnVNeHJIZKsodEJ393QmS/YmThtx9OssVVSTukeUx7YeHTI1a
36BLNbi3rFfinZc9LudgtqMjuoYKtNsap40KhSctyX/RR7xyn6Zs6GHyQGE5mw6xgQ4zBMRZ4Avy
bPhTLa+L78nGVozb33iEQPaLgY0CoKXhNl+ac0bxG5FkHvBrrVeB8ebBaQcBZVO7IsHzJRBJiMZv
hNBtHLs674CyKCiTDIZl8yvZIaRyBrB8A+6uT/xYnIJ8LDsnkn9e0Qm5TUIblD+7fyUz0abtoKHw
qse8kbl+Gd1EzV0mNeWAjDvstSaE95OQ/lm3pH6DUiFMQHt4+4NBlESvgNQ1S9/KjnGDGDjMiJmd
d0jw84INeBYi0LCAn1/Bh/Xty4aqsKqibeAmiHAnMPP8Kkw63cxPKPMyF50b3/IMRH9rGH0VnNrD
mYIgvgHN57Q43COipE+o+QqFlkrfO/0SSMCwaSrK7k9bOT3rmyIl2H1AIB7zy1PRT4BOzyPtWMqs
g3365FpHjx14NzGHz4v3G0daSX9P6txpUTaQESlHRsn/1sVqJuMy7he+A2xJc/kbAFS3J0yKbB4p
wDdQnglY9FXgf2XP+EF1QsXgULsDarLd3z3hWIoDdvSQ/hSuJ2E+0KJYqyJPlAGIWHfKMVCIcoYZ
GuU4mxB1pXZc9R7v6shNn7/GGH5cX/MKTyl4KZNdEZ8NfI8kXJ1OoD2X8LacbERhxzXHo+4opx5n
W49liwrhoOxXFOKv07LYJFh5YL7It2lY/DzqEScafLSHsqGXbZy9Pw06fSThdkNg04Bd+7Nsefyi
WNgSjCREFxmkVbAE146r7UyLK4j7ECkkcCulrSF+oCntgBnnWIyGtEGN19sOMBdFvmG3K1Ellsme
YSBX4t0sZjbhLTKXmc3RwO6sYb2qJQABlkYSWqCpX3NwNCbr+tf4f2z7MBaHZNOwu4nBkrUF72TK
rfLTsSwT0fL1CUj6f0cNmzyFuMgEkHwNmLBiILHz8DXV3kcfxBlaVv7X+QzkQ9ifzGFVzHgQ/b77
O24U4bbNHoTdiEecA7C1OXLICt1yNne0oSI31xmO+E1czxlGhnBwJirzY6+bQeZpmHi3LE4Hn7qc
02Qix68mLB+m9TtM0I5JGUepMepCF3jh0db99E9A//99fk92lcxQ2DbGCau0WzInAGQD7zoGdIPo
JkOyReFzDXsEWWnXDMQV2+m6qMPRWr2dNXsAKNjiUUsZZJWGcfEJVtICRzmBO9s788LXPMwuSXZC
RCTedwjl6Lu2gG26t1hh+oiaWPDKckgINF4Flw/Do6JUxP9tae2WlVRcXAMVGfn3D/qgCj58rlGR
w3cYgFl31md7qTlKbEZogi7LPZcsT3Pk9IIjHVRfowYJzRCAFRAv9htxL4FtQWjb5omWM+slPMcw
j9TCsznc1D3125JAsgaY8ovkXc/UvEj0S/oFAxNh3NxfPHmbTiqJo1bzJP3hHihXBlba2fHf2QwY
B/l7yaNeoSOCB+rTGHELfawYjF0E3WOifAVW0/tUFimefdf7IvI+RKIEZ168UuSNyPRSXpqU4bGt
As80wjFyVnWBJ/AS/17Gsrdw1IWanSHrY4TJvyZGKbKo341mS4dbLj1jMCdscOcayf5gBGIr0lRc
brPeOd4SZ58frcw8L4ebt0bVAOCl+48cYRoyZS1WrN+/BwuSbw0RrauW1RnNzfW50dYFSVUIgcie
H7oN41aWcfyCZWX4iBQ0mYvFZccCgdF1r0lIynb1TdvgJqYXXUpjUpkyeTsKcFNjgPJZLDDOAbQ/
RNIhwi0vaty6rgpQ9Krw521SwgWqpsjzxvZ9+uoWCxqeIkkrfEu5wtbVsC+QgaaMlzubPnmeK++m
5E0xf9l9GyvB0SJwTV5NF1H7W/Pm6jsWEiu8u0PdP1qIocVAJei5ufDtFKzcKS+9MYEI6jYomVWR
3+4B2Ks+ifytO6i65RFl8VcbG5M3sCUUdVumCcVUb8w2DV+XexNqraskAALL8Iq9XGu8+dzA3cR+
+R4cx9snxfsxs61QWlkqZMjovhfeJooWImRrhfdOHDhPRpnKLRbKIM+oBmeOeC8J0DcV8Ya1i6JO
i/vyStqcATdtI/O9nN+ooOaS6bG1N0sWQOQsd1RGHVVpPvFZxyXcxcSoDl1uayI+yGQk8Hqm5wrJ
NZnrrUTHSSo67aI6rg7mrF0zQAup4VbCMZ0XfDDX5V/ntURavfOJcQaM+vKq/keMVRq+pMMFZ7xs
+tFQdXl2WGE5NGDz0OsFjnYfGhQElEs5hoF/wyuAu4DsBeIelMRE0koDrNFJ4fI1eN+gYRkoWmp9
HwxUmq1mg4yBdyiicailnj3SVYqSBww2YdmXjk3LSrMY1hdYM6UuZ4CPtiZarFsLNZ/bDPiIn5NQ
AVvi1STp/Im2do0Yx8gB7+E5uBLlY1BDpywHglE4Ni4CcVLhxRTx5suVIYjfMBm107jvsuqjox/N
FvRyoClnYEAnj91FHljByqNrRroGcFEmyThzQmJFHS9vyvnwqYuUKR9GVwXvCS5JkioaZ+/Wf4lD
RwwintZtYP8HUm/UY1i2GtQ5PbCA/W3ddGmEEgjUIIcAe7SXs6vIMZn9B/ha42F917ahVCRtUD1x
ILPC+s9juvBa0Ad7GGEjqNmKwtJXrfCalpyxgmoCsFii2WCxYXdkWKa+yU1lmdMKP6s+3zXa/OVo
56fFt62Kv9RJ0f4iF6gvs3gOOf4aO/fOP9IVQl8EfiQXdwM1E7tYoqbgFd3D1LDtkeVGMXva7szN
nf2VFdeVJqDIRLEcN2yIFPpn/Pgliuky3Hgna7m5C4dqDOB/64EqS3MIf3TzR/JFKdiL+jvVGt2t
dfTK/FcDaOfPyYaHd8pNQLRnE/Nn4PQIqaXTLUSOfiDRZxOHwfXDvBE2o1bi0FM8QpQRCxIN959h
16TG0QwTHflRdr5JCVBU6b0DSnn67xDT1+0iqsbJzFOXI6Fb7XEviMv607ZTqywN8sUGE+0nBXVx
Ey5/7D7OAWkrpod+XZGm2i1jpVq2LCsE5zEwJSGaqnBLZyJdaMvWjoFv8agWrgHf9czHhKPWkcyi
3m5a9PcnHDetkifyii/nNl7U+9WrhFnhI6wDi56dDVgkrTm0nelf9MqJm5jmM5o61i3OWkoCEETY
wC7Mn8ESN8htNkn1YUwmOEECo9kUxQBUB3p39/yoa/cvJSD6PU5S+rjQ+ZoakrGVbw4jNX7IITNt
w9iMR/bFQDXDYnkcYBQS1W/PfBfykcGViQ71olC2xBvHhaj1P2M6rI3C2aFHhNCXM37c54vnXD9x
RhZ64L+Mclpf5eYI2fRbRfNElkNKM1lPUAthIPonMcHGIEK3IujL4F9QvhTUtJdWxK5dX/ydhBnV
2hYDXn93tHIEqu1pm4/LW/tNN7Xv2hz8l1bR1oeVvc24xj4GQUI1cjwOLkrawCTh4UC3dAB98sD/
JtEyw10edYf04a2OSB7tifie6QHMcTvTuSTtA4OAY2iYaQ4jx2hac/pOAo0HUgulxP1TZzkF8Gvq
p4q+4+J7FOp1ASnb5o8Ss/zlhcxhM53niiUBwh842MNdLppzsCLsUtrvfpExez94XdaLCb3vcsnn
9Qw6rEiHubRkJPJE2YR/23sDZTbXY6hxjIcBNqSQkAsKuyRF2HW3tFeJNmBIy9+Kp6H2JL25vuHa
g4mfRj+gWfYZ+T7sNRi2ZjV4jyp7IjU6WNv5L8NVrNgCXSF/kY+u/iOg4Fzg/xZZ5DOX7UmZf+qk
i7viNmO77Whad59oH/oh7vWZT1c+D4z7mR9LE6YlDqnV6x/Xl+KfKJo6kkeV6ItrNExyJDglRpxf
tJi20eg2gpSlxhUK7VZOBbM6V176e2zWSQgdlau4LuInJE3PGwYondkhgRRsL4lezKv9bKCL6pLb
sQr6FY0pt31Ay2u/eQWBAp3N65D77oVqgbaVXq1a4cthP/1oLWpiaRLc+PHtYMrFPnlbpXyUjmX2
Ixe0yaQhHoILWSd/ubAVVh8vhVLqiNG1j5/X9yQauTH4Vw/BRY0JPc8yFjqXEYzgS+AbVNXnecSE
zgG0kdUbdogAXqSOzyPIZ9imx4X0XQvmXz8ZdAqfGp+rH8hRtxZDxu1eubYe3iOtpZ3BcHF0z868
N5O+6wGb+hioI/x/VWDI67JtwxE0rNhYnSZzFD0yPBe8z+Mh81SUEruE9tIhaDT9IEKkGdJd3KPD
Onz4dvtCVVzLbxXQnbnpi6Kf/j7WTassHblFnDiyq6SLuU2Q+ZTrDDGbJTNEsmDLyL0swjJ2k/dk
GFA0jONDKzHr7F/MwGvDLkd8P5cy5Q2XyFKwCKlCdPuixEPelUPbEIXPqMjTaE/YRLjSGGHcVC3m
oMXLYZPDMC8ZwXCbTSnOpYPXtR3Ah1EsVAINdyFusazYLwsGOngNujiiW5z/mAEMJ0Wq5o+uQzXW
M0OcD87IvUtIToZqz49zq5tkGU9I0VInHrpdFFFTTlciTa7MtWfP/d3/thF9cF+W2E7zmgeKI8Ja
U1wR3mAWGg7Bx4H76wloiwtIj+vpcbfbutPfo8byfBF4uz1eBh/h6w9vDanrwje7ijtRmG3Hsq5Y
7eHqou/f9r98JL1Miymum8ptMlea0Z6p+gf+8Z+OZcEGv1ylUB3KwQz0idGDY1OVJ2ssrcE+2OJX
FNaT/LfUFnXlOH5IS3wBYOyPD1BIDy4hBAKxY1J4WCjKlrW+2jp0tbRNm7reND1p8IO1cY1rkyI8
MjKACZWYdaV0nbXGCe0uz0nBr1zul95en270c3D1yens+/W9MaF/HAwRjj1ENvMVua1CVRWKy+m0
n88eTCm0FI2/Tkif/OOpsQdJvjW6uvm8OLWuTMOSbR6/ZC6qBGtFKap9+qTKDp3EfrI+3yjsHlX2
Rs1x5N3H2GWYW/009oQ0MfAeQct26tCzjzs+R7npGpXbeFOKGZA7UV5CpFaRZHGmPbaQFtQtP1pp
VVxeFinsc/Mpn9UODkggEk6QUCsS42EPObMz02GWJVa3PSSXAwQShd+ghm4PJ1brc6gg2JUIgWnz
cXgQ0FZH7MfWpabFP7wKL0bYfnQOJREfEK0LvIsPJ6gK/7jSWYI3Rc8EbR2lX/UzlnO6XBBFPjrG
WpiJ3aHkXdXxUrHDz97FJaDw7AWjX8+oOvdaiz7hbHYjYLmwIdrLQEqsk2DFEYWJszeC59wnZq6a
8nww1/PYfm7VdNThpZ/Ckh8Z09y54IVqsJpuEvKRV4vR8lppxIwIg73LtM1pKJm9DXg1LQzU5MzK
JqWVhqliD50qaFO8E6ITXNBtnFdr8PQEhfj2UVzZaWzYWzYKYWVqircIPZpGpbehgzy2qdHPYE/X
1ja82QkB37NGSMZ+GxEj3MAom3Iepo9Fsgf1DyHeB/pUfg/y3531oXCravpo2T6XvAdulEkmgXTo
g/TwMT1SCJuND3tOPa2R+Ll7xDEAmkfzkXmz+FWWt+4vJY32KDaNQsXMutve3qjEb+SF37zR9MDq
kvuY9FVGfliokRoD93tzm7m3D27yZEtSh7BUTFqKT9Sa80LF1Macr3CJzbKg4OmIJqpbIQ1exBTE
of3TbE5AJYBhaJp567rD1hgzsNM0+0It/vHQXzeyZqoLjfSjtbOYWv3XuvoculcxE5C/fOIH/48r
VEXmOBUOspIZGQ3eWrhXq/R0yrLcqM2LURVTWrPpK5P4TLMIThf2pIucmHDHyeO4BZ9GObcn4FYd
VBjNIVcGJkR4d8RSY0JMGNsuQTzeHFYhCeaTnCj/MPk17OzFcMj3f/4yHoA48Hb5C8gOPDo9+HR4
UeyC2rH4BjQKGgd4fmt2UsVJRSlBr4qSBYMD+ty+CKE/zCelT5p4MJsoXLJ9RBqdVIo85PvlH4f5
f/UiPZTJvmi+wmxBisi134vw6ge7Mq7mAB4fXNivrzmZ8BrlJV8khxBFc6R/q0/+0hwc0z8aZoA8
sDRMlTlX30EgLhC+JBYsLlZeeEQ2APs2H0Jk/M6dmKo2phRN0pLv08/i/g64EhJ3ag2rYXzwJl/3
/wVipqamVY5q/N9x9tAT7LGVAykNuAcwRcnf4rPZArW2O5BZ5uryrHifIwsEO4cP9ymNydzGhx/q
UeVnmB6hW/HKNxaVojujRmG1Fzho6H5+nUNNnP+/z1zJU/qkxInzqiWaNy7DgO6bf4r1o6WGaEw7
aYEW43n8yH09/O0O2nuAFbjuKZWVJLf4neYwR2tK3c5OueCI3V3pPSaYdZHjJ+OPbr3rZxw5nrtU
9dpy0wpzPh0Nh+Yx8kTODqnRH2T1zOb5eTJBNmaGJCM6O/lQa05E/1VZzm0lHau+RVvbBMBmyZnG
BjYkgFHO26azOOuuMLh0+jl6p+qXE6edFTwGSaQfi5yc6OMbuFEERnTHW1wU4Y5nBp5WM4waOp1I
dPdFTGQ8Fd5DJz3EDSLrMmOeKXcHPaurF4x34dcQojyioQ3YA82VQz0M2GAuPkiQPnTduKmmJxNm
BhTx48pr1G1nmjwQQWqYcg3Zc94Akv/062xE7BVTUn/qtoDzeVY+KNbJqVv8O0+vLto7naaFSNiB
+R5kWC612xGMscz04TFgUKyHN5H5EPymz5EjPS8XRg6xfSldzenuqC0BNkmg6BncOKKimIoJ5A/I
HZxsf2/xBAcMvSfpe5N/2GwpQUzJ+0ZJxEoxq1LDhlDSl7l2Ve1bR7xEsYOMwn+eL1SasvQYn/JC
+/x/qQ5euctTHhQTIyWaf22EmhOJarMbM9jtFZ78JJSTzPLb/qD0eD8jc8xO+2Jp7IeRrO1DFc1m
HIhT335idTD+5GzrLHEuJ4f9tdZz+rxmzsMULJtmm/aJhVOpMNILuOotJnGdL+OGachrOshu5wfe
18lvSPVN6BFTVpjBqhr2vB2TAiJ6dnAxkkUHoFcFmYiTGRias9KEqtU2a8Pd2Q6GWJcNRlNSMr6n
FCYUAX3Fd4riKi4sPp7O09+R2pr2ACTKCIQw54/pHR4j5v0IqvocxPKmbHxTcaPzSZA3zZIn9Hb1
5u+Z/KBo5D+jIHmCO8RB3bF9gMQ2ZG/EODyUoUH8HsDot7wETJ6z8PEvBlwLjxxUQtAznMT+k89i
PId67K07jpmyBzk4DFsokf08uYAAxQbffLB0AmkOjAUQsvQmTcY5/kafK/q/6gO+pgcjIWxwT3i0
FXbQAKPbpwtPEFUq8lI1L6TGDW+/ZrH3KqQJTXmlACaqalzGBEd1o1PhPr4NCzl1XmaLL/vHWtnX
f6KHlVokBvudHVJlEPipQPux/PIJtxgnHCkczWWlSUKwdeCZEeLEZe80rixWZzaL+pwViE1KEwXb
52ppkbG3XMa+AyLJdqlWv1q3bhD8ePCA2zTZPV4Op45G4nY+OFOSuEf7S4ROfoZMR9k0af4CUw7k
n25LyIiGEZLFe8Nkl0aa2585LZlF2p7aqTsZRe58piLJrQ8uJtbUnSpksIBRGSW4BTjnXot14rWH
jDknOR+rOE4grPd1sxEvep7vWFhM64v8pwc4MWR3Zkf6Md3HhcodOs7CH4+rsvXtzISo1aRScigl
cBiZhNH64mdvbSpRJrNBUR8HwG/SVrP24lCBHlo2MfjXA78BiRGloQ32FYtj3VbG9m1eI0o7L1l+
lPQ5/3Iw9dGg43+gW/mGI4mrVUqbTY37nKs7h0QHGDxdo0U/5Wk4zWhKJop3U0C9v2HsRdy4qxwY
SHgPdH9Pbw+Jc4ygcLv+yo7/OjkG+WvB2JazJy50Zy1QZuyvxJimpO7NDPDxFPUAMe9vlPTEoSgm
/iWBdj7ZNf8H9vPhl6RkYgNnq0YhvyU3IWo1QRLi7Y3FTdDInNEBwDwHSciC+g9CKhlDh5YyiIpM
6orXbzwvONvoMOa5Ensj2euSiJKO/YTHAjfhpHRHot5Ufjm0f6WAiH6/8T976o78Xr+3ERKCBjL5
7miTlRi/SasLNRh9hCcpxcBqyuyKONmtVMV+2dN+Y4fLRIPEaj8YJwqMxtTzhsCF6zqd6EB7ENr/
ANPhbGQoCtOOdQBc3satI/L/LC7UUcLt+HB8WWj9GsyYGVGDV0wR6ehwFFHgHsHPv62Y04293jPT
o7yz+FYMHG1CK6OL9c2Ue1f+pJBGBiDVMhog73Mhb0KeH6SddtkVJtFyvMpebV9FHflefc3LhTx3
dt/4/zpsCfsdM9nrbkirk/pgrNB4CPOdbOMtehe3PZWxOSnzfRLWLIK8BxDfORI3effazKcJECz0
L9U0ZcDE1aueDR0ci6mol/+40vEpYE63Cs7dK3FN2CzRFbzEpiO4/DwYNRnT/010w0Dr/8Jlr0G0
rSNjQXtIeI/Jao96gZwtp8sYmNzNdoD9li8WS8b0KMQDp4n0uGoB9APnoNNbjsaRLdMR0d87SqzE
FHEv8ou0ORMqRaMxixcg27XilNeLuZ4VRBlX9wZ7H15zXHYdI3qGAScU38Pn9cqbUz/XO5dYcyi1
XlXczWNYS925rWfmM1nRjMxjF/LFtqbuWN8p6BWTWTj4jst7oAYZbEFOKj5rk+5xCqyQUnFhs/AY
Yv83DSdpEHA87LNFf8YWxt+ISXTJZjoUEKw6CoTvV2je+nKGkfgBMszEdIYSzOPJD8ZkKCZ6ZMzC
CKKZIcaZ5TOzMUT6dt8PGPFgI4p97ZtNWDbrjjO6GubWbA7W3SOpp7y3TCo3SUClGi4y1zLSf8xS
vEoR5WYomRDu35MTzyU8j/3La3/zTx8WELvkFdmd/cNEGh4S0LxS1MYrURY4vmkG8tqz64oFC5Oo
6g3j8xEQpkzIQGfop4KZzGBJZP8sDoNIxYXBPhFyw+EcNu0+g76ctf5f9IJ0wl+SmSYOLe3Z8fpR
i0aDr15LrDyu7dwAVMepnk4d3wQOz5D9rmHOKxqUczfCkOmkuAlUchGcVKQf/Vagp7fPZElLhYNU
L95/6FhJvyYmzjsgkCemVGkeoCCCng6IXpkBHoauu4kxd+cHOM5V+3yxjqHfR1x4IpB2qRh9J5+o
45pK+TEHAKkb0zhhP3mpxrTF/3S/XyBJBOOzS2lL1HBqB2V33nuKSOBYqSddXajyKi7g/gcTMg+e
bv/JcvLWpUzDdiZXSKI/PTadaQj+RUgzPfoGUQZibIpJS8fcpFuiI/ccnQ9InUh3UTZg495P2PKi
OGnuoZCYcJOh7YXkh9EBHb3yMGQO4inU234u0TUTIpd+3WveBgYl8mAdp5bDYe+DN6A7MLU1JXS2
JJObJQthjIWMOJ/7XqZooLDLhwhNtxZ0F9DeNOErvQ5kVk7Fn2vRgzgJz/c+dQO/4qHOn4c2+L45
JZNyL4Jvkp2N0ASYZUQoNEO//4e4asq0tUPGDW++rLRQmWG+ioccJNfgf9YfbqPfw3cxDItdCmzU
bcstvbS63mFxtqIc7bXFJHmr5Pxs4Ais8SaBFzWJABvDiLYOUQvGv5j1cvI2E9V39v+yAhZne9BY
f/uTgPHCbou52usvUJooeT21wdbTL6X1AqeKxVt9F2cvHzsQrlTzhoeGrlU8fj1i/YXMx8s9Kswo
SPa3XLphph3g/VX7TaAVZWwaC6Se7hZ5m30Q+4Q86hicJxv80YzVbg4ZoYIbMiR982ebxcA07eA0
xM0a/aNcKFqQyjfanI9cCmhEjs1pVvruHakvwGpyKaTNfld/TOw8ZDAKeasTmfngZJmsTjx/TP0c
z7U1rT/My9o04orYoRenCbvLwZmIsnfaFbgVXl7QFspg/JCv17mC2gdGHXuShcNtBN9OXx8yj3AN
niFp8EUntm66dAsxt8P/QvSIr8fcItI8vGlJrY9MosW9Wm6fsD9Eg6h8WXWoJQym16ZDr/um1Z5B
3FVOa+isaWkrY6Wd+AzUINfXZ5o7IzNEd+x2iBwJDC/sjo5O5uFP9hA/fuDdF4RMe6IborNRIxvQ
lYIYxEieA+8A3FgHzIvbS8oT+m4ARlLLrTH/htQ8wnlXQZb4UVzyPKxTCCOfg7eSvYvt5pj58v5e
/Y8CliLiWo01nv6Em6iGolFvWIjY7aA73IsLKv17/wP0H+xxV4KVFaLefRXKpkjuYDi9eMJdHmps
WdVRhya+UEgTaoMTwMVeVrGnHQMKR7v7jACoR0J6cznURBsJNsm66xJa0wR5AKZB+lYYBfYi+yut
PdZMmLVAuOV439ONBfjSpY6w9+/1+I8TatKYnUbgwACo7l/+ua+rQkblZYMJwlr3xkGLTkOLNPdE
/m038DVbyzCSpOwlg1XS6ULMv+yH5J4NrGhp22mAfbuEJg3SnJ2yyNH6GHfpetoAQ2+s1lmmi9cg
BpXCOUIo2veIsJo8G4qKuxBRI96+Jz6yDr/EXjTIT5vd8L4giEyeOVLKAy296GBPsJCbk0hd8jiK
kPqXPYtQ8Z02gHzguNEbCVzsk9VvIAZkc6plmBfdzaGtEXQpFeoPnftwszDOBnPNH2ANJgyZuNQc
3SamNChs36Ch6nSkZi51ueKeMqWX0b0ZMbXtHKoSomlPgnSgVaIGVigHW4F0nAStJuqWuwz/zFgH
47kJYk+hXulBZEytMRz8nmtSzX18WVrjugolDtJbmefc+kohyQ9hdvuBvFQyQYBQinnHUfcF3yPj
iIRggWAILiKbImzdDNNb1xyn6hHelb31cLau4GsigyWNqmP42ThGYBHPb2Y2CVOqwxC9poioRPLm
YD3ZPfxod2ZZM9kNyZivizWcNvDoLG3+AszxVvj9G0683uEIRcmJ+PlhOCdF0A071B/sVg81GPBb
5kjFf7yAgQvBmSeABlQgwuNhe3UgrxMP1VSV4yzEKswnK83IGEzoR6atTdN8zAJBlDaw6W91iTJv
oVwRX1HRp7cIPvLU98G+hX2eMzk0IloEkcRfPHsABU2d9lUWuouINEN7/v3YSiFR+LX9uuuOoLE9
W8C8BYoIBcmenlKodkAnBUhUenq5vJKRLVEdY+4KNnFJ24+EX6EmB5ItvjDfrM31VQNqRSCRG1bQ
YLVdFTi12VXl4ATPZtjeSH+38SCsZew0A4EOh1uEZ8UGzyDE/taNNFDrBGfiI6klrTgLLn4m+DUf
i0acx/YlDMEZybsjnw1ZHhAu6BoKgL8znqhv+jKrUG91LOdURtcqMNVMEKpsrgPEgWVEg5/k74T+
p2UYHBmzpDIPwh1PzWUnJdyZidIR+DoTkziLhId0pTxsRsCjjZZlge3XOFOCXNVEdwGzq4O+tian
sAokcBlGR/bMNNpc0QUuGxeNQ0VIewfy5cqIzmZqjAoN4ndRG362Z7b8bF1AIS0GZGJPC8MPu4X2
uKUEYNLgX+c+3Y77WHrvQZhCs7peosQfOtZOhBkcGCRrCyJKuuhWryi5kUwqGNdG/yeYvuwiAvRD
hlH5ZGPaPwYJmutniYDJAAna7YHCl4Gtr4c7b7ccGlIvL4YpP3YwKxlESHz6ptcsr46/7SWlZrB+
/KHr+q0cjandzV1gtJXJChjTBJpIIes7NQ52o8peHLk56Yp3DccU6DDBX+rdt527ZcnO3FAYgRzr
uz38Fjv/q27nwtDDVASAsS3E0M4gFoZ9JIktXY5XhI+hqZgPub+dg6/v7Orz18tuNKuPjSX7Cxv7
ANyLOP7odKr1GcMVoQeNcaE95G1DNkYpmCTaTo13bDQirplyORxBzmOtsc48fC7gssdAqhwADYyr
NQ7733fvnkafBNepQ8LpZ/F8lZ1l/Qlng1BW7ybVRwxBjXrfZ2xloM03F80lki6Bl5Nv5EBqbgBQ
ZtYYHR0GV6JMDwoEZbcABWQuO0+pXhyQ3lEzGsPvGNFZcdtAQUd/dmpaNDKH0PgMFverYUTodH61
BhEjcaPsvCVw6UBOEfEwEp3L/479B9sHbh30aBPzty9LNi+sgRl9e7NcUPtbpUn+XKZsEJ+Zd+Q1
EMo63JzjqtoyhzU+jekWLy7uEEoHISVcLwRXpDQF1r2RcA75AO5nKLJupiBjAe8tMJUdgsVVoELw
YjS2jAWJQcpd9u7JAwdKQhn4iCky4rdVIQvWXScfVOTyQhh3MUlAxObUTggjdgLRY9UAYpe5jaOg
jrhirfrvD73OR0dbiWvmN0Ham+5ki9zkAQ0psf0N4OrBw83K3AdDjqMsPE63FYXKwH3PQF+n3QxI
PSPVB7Gz+5IoJhjt7BgQTuwR5U3bU4ToMCpKlIk4e31g6gfA041gcJHqvoar0wPEnPVBIZheMawX
uzXwKZt5zIf60YGNswrGYmeLOHvf/S/h4FuX62bCX2dsSVWCptQ/aykPanM7sMwdm2qjKqDcZetp
xrgup6Zkn3nevigel7wuOzXaH6pN63l/QwmmZeQEyC60ddwYdlZE3cGJAhFGzxk1FsZwWZnCS4Vv
MRn5mCaGVJ6j4P6VWpp1RRWYHE45UV29L7UlkeFv1gOn6uCoPR5Der9RltVmu+Uk7bwNVh4lHtau
2leSpbQ1s7kVb8wcQVn6xr8NXmwCUPhm/99PEm0saKHXi0gANKvDbtd66/kpY01k9kz7s21UMwdY
G6RwVnxBfWF8CuyX84Y/n456CNRWdzolT8Ns2xenlqtnJwUFTC54Uo4AlRsaAX9DEdsQZk0ANw13
okCU+uT3mlYaSLVf4Uw1XIZRGhckYHCuF7OAoq7dhQZ1eIXxax6+5iEdwhMM1aWor662WshTK5u3
jGj/gfHyyMrNQHp/1AS0HgEbXSqRhM5IXD65vjBzQv6oRhXaQB3WtAtVQnEsEGJVqbg/zNArSOcf
wZPrxnfx3JXmlRrnIo4McWEZUb3ioaX6KIhc1ZhOVRB9GKshyigJWIWKOfm8AZ8BRdirGm7qX9/2
slrSAAxkHU5WFlb1gXyI1ibhwina/oxQzmTkC3/Ikvg0Z6dG/4EBoh0XX+uquHJ8PVdU6YF0jaGi
Jlrm8QWnHEV+YW8VS1kMnVQQqUaqjEM8e5ZKvHk/LOwyA1zINns8idtntguconb5Xb6buNRI/I5A
1ohT2ICL/BdqarGVIQTXHGh9zKHGjBq19BI6kMy0XRBBZsvKSL1ls7YAYTjZL2G8MYLFndj1xg5s
qpBT8PgGGAQhw1OQ3o1NU1LzjuWmNQOZ2KlNx1c7A2iIw+LW6MGJuEaNAIqbbuBXLnQIhmN8oqiR
6LAUZ4LR6oGfycrozfWpIlBCwu3ILdPWtpAsrLeaaMFlIS26v1l4yQl4lJcenKjEJ0zxC6LTO5wD
pGxBasGAdibn/0jCwvkxBUqCXjih09xWsvQo2uBLWzvisogNlMEGvitq8/AMUnHZMqkNmzLRYFCE
AMkmZOOHhg7+rVy8kikcCyJaPq1BO68a5eAsAbHDTcb0VHZyfaLfvKW0ow9fFKkvDpgMkEMZ5Rw8
Weu3ksNy8CFuuJTL/FeqtY8gcTAEtSFOI0viGLlof0m+OnRDpdj/uQBZLjXqR84l6eJBx6CSdZ/v
uLYWV0GrGczrzJvuEP9QDvtxJTq7aza2+IOKUDnTw+GtT5Kw4IXGkGgJToRSQOVbYLQzfJKVUB/5
z0raKml3iwawQp23avlTCWQmdFvpZRK5lH/ED7uU4e4PCgYewSjV64keQ6cCcQJ8u+Zj93OvvyW5
JtvzWJFnLZ0xZyEfEUoiGvlmfL475i1sbkVi1qtVErIYTzO6fultnSntyZOiRGYfOPUJshlc3CzL
uecZtJ+Mk44CWG36TrbKUKySqJA6soxjbMhGrZgfxypzaQM9xGd7uBII+HzI2/ghSKN3+umx5oWS
3hJpfdqmhI06uR6qLtpG7R69xFZgoL6v+Wmt+P6jhCML0gjSOxSSE3Ro7vADz+JSCeGeNiBAkLj8
tOnlWpaZs+ySTvCpAyp0O20aDQuzDl1pLJwf9CYPyMpcwFdRCuRYou55lpFddA+/VsgRufGHonL7
ypZU7SRp+sMHHDCAW1/Hc1CBfJlrZG6gDJeqYchssBzt/6szZliPioZdPHqq6tpe7DTWiu1ustGu
BgtqlEv7netd3e1dgnUbM0P+YR+owbVdiMSo+gvPEGgjam8YspTOA8iL4hTq5FVyYdOplyAgUZZ6
TtmatPPI0Uzax4UEgwRvQ82bOQc31diNtQMiuA2L3wJt/UKNvYxS/CNGBdhbIu3GTeid+eH36lOp
z9Lr7oZS+y5g0hI9gvJqp8miRv/gz3p054fAGYee0jT10SQ2jNKN8P96eQTZ+iqD8utE0fK/cIx2
p/VfMzGk3IcU5+wM0HrbBWLBABsaBcVQstwHV1YOjqhq0nRfcbGP1iQYa18OEeiXaUgpKfWJg9b4
2J7IQuozlOCQwGbQ/igCK5r1SRpdKQKQqzE5s+nc0dYycnLSodeBQ27OgcWyjuEftMDkWsblfXu3
6cvKkZgs/0zG7axVzXx/v36xhNFjZ/pi0oYiLhOB5XfJ/h13/dMue01ziPXknceVWLUMsi/v9Wkn
el2N7lNcni/e4/DfMm+wiMu5wAHScG4MDjPjYCo7+TFziMdEAXOV7KUuQTh69AGGv2SqNkMWa4kt
5ZpGGQa66jegIrPuR5sIDpJEZh29QuoEl3HqXatVoyHg4p6MN2syBS6TrGDco0sdHuRlQs7gYZFl
DYEuDQ7CnB5gFdU44J+niaYJcHso/KE5++JftquVkELZnmviHrVFoRbzDfQ5cKZ8E8hR4ry7OfGo
RfVmFEpFrZVu+1WclWYb6yh2uW3pianqOI+sUnDy4/o9DBWAekdNPwosMyM4zEjWtaBvWmSS1o2f
s4j3HXOiKaWKicXMPj3cTi7nrgd9SOY7UKSJSRAwtmqxpWTv3H+ysZFUcUbLZ16xGgx8VZDIQdyx
R3DBHBqFbg0Jvg/Yo4ALKmnipKuksC/irst3c6Gw9KwPOusrbn3OX3RiVYSa0DCeZX4ZnfZ4dyqG
o/79onYfBURrxeCaCDpnAdIy3WtulJoqp9riS2MfRJ+duhko8Eel2Y5VcFBFrXi9J3onabH3Oi9c
AAH3dmlvd9/6ZuJ6d0Rs531FOM2Y0TFqUbDCTsvT9sSrixiH5L0iP+cnHW0oVvi9vnq3J23mYJDD
5mFLIeTkbyP5yekWC9QRc5wM0DIyQ2KSwkQig+C9zz72r7HASao1cpgZVb+c1CpZGgfMkAqqUqG/
2olMXl8H/zLe5m1ghNnXDfBVpxr+SNW9COhXUcb/fnBNNNp0RCfheRav00klr8gNig6mJ5VL9Shb
fOyynKbij+ZnnXRBAWGZRd85c3G1xbJCEPl4vGsEcz3Ke5bjvhDV/ne8BVvJH+gC79AW2Q5gjVPJ
IVt1vSVMz+c65LxhhFIYIg/CE2vaHCCcMeKJ+kJhLzLjNOhAmPApB2FJ1IWjvfIbJZg90gnGPgP8
W50q7u799VGBwJkIUL+ywYfHB0TBu7bQ1F1qTIGap8iPiqGCuoeCkBThlTr3FRgT0xmm+rKomIK/
bXwOedPH/wRcEuX4EOxduINQrK6UgsrgFHfQd/bQ+OLcWfN39gYSGNK8XeV08NrryoexPM21XuSa
sq7r+oWlg8B7PR6jGlqHgWOCJybPb+Dw7qPkUBYGlWR/+4w5QkjNL9tYc7OnKz8UDBn2jWePl1zX
Si8Md+u6Xx1FxCgQgxrBLDySj+s21Iss+6RSFrw/p84M7jtGsoerVZg7SiFWPNdexT+HzFzOPh6A
6YASrDeYCWIjW+vbNgra2uu21lG684oixkHoGv7AtrriH1/M2bJ3JinBUs/vcIVLgVxdvroM3CAf
6eRJXEXslxUbG8aGsRavDt23dD8RWV/XgjQgzI8J6ZH9lFvalaSJEkgzhEy27eqj6IeYqQjBEiHD
spHTQFlfOVXZXzhA7TDQxTnpgSEmbGiTdTTL7yGvcIErJxdPzmSXzu92iguHju4AFJPKenjUawzX
ELI3GPY9oujrxCDoGIMUH4byrcuLN3IdHoKpqEXwrDL0Q9uFafvsUCIUNmAjadb7gdNGerGXKU51
rxkmIdoGWnv2sEF3AuO0eIGTKsOr9caSVDjXwJQYVNaUpXgtQew3KyeX4dAmZVHgSJWh4DwrwQS7
eFJOL3FrkbGyq61M9030AYC5SrDjoULv7W1++B0jVy8fUsdS6RDIv2DaPbfJjjBVwhB9b98151iw
HPGS/xkLG/TbajDBrIscgjpz8znj/UtC3ttnKh19Hi7QAqMqSWesxFnXWrnC8HzLwoGVFtU9QkFY
uxq/GKKltbJH0E90B2aILGwmaHtwoQJYLx6nkVhWqbZp921VdGAeLGXzChkl5/kmMYRSeDYdGTXK
OwW1VCIA3AStcsYySXmlrjf8WlFvd+PLZ+QeElbTrl22rQxzn/XoRhDiD6G40krA/YX7fVofnUOI
A2syq2Mi5OzkYZHy3qstyVd68CqIkkZ7GdrT9t3jbFxSUaNmun2JmcSl1s9jQWlGo5RlGEHJWf4/
28yC1Mh9Wc6fw5/73g3Ne3Ma+zdu/5H0YI3xRd2SvccVnihKf7yt1IRKe/acrBUSrWEvMjEtZooP
sy3F+nDmhpPfYuNhI1VtHSxFYr7ZEOhvLrRIPBRcOnyLJw67OcHdjHh5ahk43MPa43Quts1AZRmI
bKOeM7gHrWsxe8YXJEZWSwMH23FfbcvLceCcHhxStQFlGZzXb68dOohAJJrrQMtSMiwmkdUsA6M+
gBItW/vfHDPnbpce2jOkHZHel2bZiZcuKwhT+UMH/H4Zjrzywvjq2Hu7ufH+MB0HLwGHG5Zd0s76
ngKJJzXbBmj5pG/aQAJNZpez8YIsGTjhwAt2kCMYjtaJhvUGkjbC9wd038KEWx3zAenEcbXfTV4/
pzVoJCAwL/iB3NppYpxq8NOO5m+zAcZAJ6DdhoqwByJHuIenxRNEd0Q9s6EKdQoojAbE9YEfnpCR
us+ys28iQiYQ6huxzPzvGdrJqQTH05cuBwCiBwCTIWJnOO1A/v2BxEHkedkX3tfjRBCuHh4ZzXas
CTlsKXNmNcgUTZuPiwBk8d9T82YWQtn8VQ3woBSkzWZDW1/GrG9Pbnlo2PdcfS6QC7QGzuRsJOV4
pry5g56gg2dm96HXRzxX5wljxRJnf0DO1o/pJS/HW1gy6VN+UolfbEfIsLjuP33S+CfO0eKc29Tt
vHblow2QFZ8dL8XGJF9uX/0vJl51M7aSG0k5H9BTOCz1Ey+mPqBists4Lpv6GHRM7eYECJbkHRfR
kOo1lupQI4mjc97GO8BCONbi7x0uJ0tr+yQdZ3MYar90R45vtYhqJXlH+ZwxKsSa18P6ZjwBhTV7
GGyn5QhRTrf7wOtMnPo7gMIv4/lMuM6Vjy04GVxFvdZLIIo9J9vxy7Q3pouVH6BU3JSiYyVqysLw
UoYu4+m7QK0EIyATDyv8Wvs3LQ5tV6gT+nP0zqTDuMjRkO52tzxDOSqK6cqbJ231G49T3XTj9xKX
hdz59ceeZ0MjUIOXx+/vpNrStgUeHkPAvt+TNYEUObwywlGL+YgWZ3/Lfn4Atg5JAJyxQGSkYYek
xk09QxGsI4RNQXvzo7Bh/OMb2EsVpjmXGukInFfM3kxZhChyYBc+n2FSkZmwdEcbsBWyJQjqptFx
JSLDUelGYCSgwG2PJygfCwziQMWJZXwU93+g50Rc/j2ttPNhtChEp1p47w3wWP7Rpdrn7lnMTOuz
FG3een2UyQg8KJFlnvT4iedOcuYCp8jDltCHd01cad9LktKje/uJ+rDj4swyoAAS/+MGBfoz/IuC
TzAsmVqzeNWNVK5K2PaLA7/atgbi0ilbYQjBdCev5atnsJy09ejf5ckFx39XfaiMhAjbu6IVIG78
iOZhAMJZtnPl26LdwZ6qp0bQgFAH1QKsAjGn8FXOE1F+cdLnmRfaX5oI5xB4kG+IAwvUMC4dXFon
yOy4rWFRth3dcozT8Dl7ZsnWmqY/kMsNOT/6Pr/TWaPn3yRtn1FSG9U0Ui2gu0TacIcVeczjUF5O
3yktauVlWVeCc43iDO1c4YZQscjt84YbZ595XdmX0Y69Z1meOem1FDmSWBpcFOROzqqTffL8gyY0
d20lnORDQLcFxmzsvtLmRZpIoJHuq7h5N/ph1LXMMFINYcQMT0YAIG15IIP3sovDCTrv8Zm96vTp
a26W8q5GaIcqnCrTezNQMC+UoIY3PPbyeBT8nbr5QtAVmCJBtZvTqNiOB504veqfhHnHSzOFST+X
Wtsee/uSa1H0l/OhWSn18aIFw+HU0NbF23tmYzKZ/VDOXxPV77sL83YD0WmdcNLUTwGK8Cvy7CrJ
MhuX/GDQurBCRfGhhsrimUt4QE/jl3l2NChD8nqd0GTAdB3ADmCCg+x9ypWrfhI8MpiDoM2Uqne0
a4iaRbAzem0Vlxj7Fb2InfXRx9FQyBkClBRAaxqYfm28T9kh3p6QQx4GObq9RXGpGxZSbNUhrzhx
K5tPli2merpbt8WIz0YgdihUIe5vNT5/Aat9lDQ+MsvwSEWMh4S+1gfd0KX7B0by2sVbSRcB4dRV
OMWTGwVy+VYepoxVcuGvRtbeWuYoqeFAQkWjF9JCEkdRibJLN3awe4U26W4ajtfq5+eZyzq0AgHY
DQJJ6mBRZ57h7Ihfg8PKs1LNjUe6Pr0n1rOZf+DrcQNclacxcMZ0FvVYhpbTHX1sp4xvcOiLieeY
lB6Ixqxbngl8KkaITg1lnQfKlP5IZCm4t5e/d295nsRZOjj5HK/hN6szE5AquoxaE+kXgf5yBQrG
b1hF2Os0TEEcBhsMY1/BSW0/C+UGM4+Iv1X4KgvlHr2MTNacuizOB1S5zIPb+E1bd8pfNDRYhHrl
FEZCCQmQtrXr1dl/hBx0KQdFp2Df/p2Iiq1AmaPGVEk4CEE8XAwHrAtK4NGzvYVoeLlYCalY2BIg
7nPmRzTEclM81VkxD/l8DaNLn+xtCi2wTIB8sphcah62oAJ1pmPeY0qHnxUNpifrCE9fWi0U0d1h
6VXLScR6u9zIoIQmucqzClK2gYiG5andEBPRLWKu6VL0eM7X4GZAAonxlU9A8QFvErBnOoxN7o5G
v7zn8N/Dlox9RTNTtOC6ub4YgF12UiEC4JuQqmBATVzT01+yhAhoiirTr1uAlBznuYlQSJO7aDE6
015O2atij6cEMVzCJngb0wjcVE5WNC1OwTanasb01DcNeUoV7Fy66ARn6UaeMM+VZ7P37Lti2k5Q
jJxgSdtmxrFe37CDZ6LdqiJrNSPqe58CdXCefuQ8NtN9TOBovsDxQuRRcWnSjN/9Gun7Ey9Lf7AD
VaNg37zwNhzF9gGgq54hGjT0MuMvMFOwMJ46F6/KtPwyD3kltLgkeKZ2imn5nOlcQFqsUwDYetr/
AH7USlGzlIhMwEoMup6ZIjYyR/jwTQVQ8E6xHyDl8bp+f4DZ2rU4ZH/RDtPgXdB6i4bg15hjHQL2
HPJ6Dv2o9bkKQcZhuTx3ZKakrJ5WluwXrY5f9zv4AoJi42l2iPHF76G72BDyNJaCpYs4AHB9g1a1
DdUDxDYbvVaLDkfuKei2ml1J+Tgulo91yFRodTiKGC+XlS0tkEbU+isrDC8UK27Kl8FXztGQmf2v
eOI+ID1EiEwptFCxyRW+FfWT4mHwqspOd3Wmr/F76BAP/ySE9rvHNd9gNN0qxz31nac8yuq+J9r0
VHMUy2+RKo0O+E4wj+qkMMF4DUR3hgQm2WEplRJtHTcZLBGiQnglUi1mdfYwvLuZwLLLQgKhe0r3
BM16N9Y18gq1hR1V46OUCqJCi91hF+NToRcx673TIlAXu62Y1UQYO+uOCQl/Y2Hz1T7xk74H0yEl
rs/CUyIX4XvfN5zsN70oY3cSe7CMa8AH1llVSTMKy1imLwWOMl6B4KR3h0pPDMWrFFi+k4UOEvyR
V7ukEcZaJj/phE9m9HIcmLqemXg5MhAcpS5Z0UwaiG0gLn3us4B+8EeEZW67ho2t0KV3x3h5Uqor
uJlYJ3fNKTy0fSeFWXMXrcNvQIPj+r7aGPeWN8gRAHyb+lT7kPwNbAwOl4nSKtxxiwJjnwcYI2WT
j4TSkvo3KhLs62BlyKapN3VYozbH27HCmuMZF7bqfLRu//BwUGE4m4wQTYo1gJENdfClweIU6Jwy
8Hv4x4i/rn0ywBidWgDoinRMHskWsgXVBhKz50F8G6nLqIwAWC4pGtLcaVEzMjdiddsCgQ4tjBdd
6B0/HG18GKIkwjBck7p5BTYZseIf0VTuFxY2ttmwr+/9K30KfIsTJeVNLK3BJhexOhznTAKe3FTh
QWvLj9oGdo+vFpsp+jWvf1fB51Zswf38SXhbsAx2n2DS4uzcYugJdWFqoFhj14XDB5g9Hs3qkIbm
OBRQeJHZ4lKgknjKFXAFDfnZd2D3SkJzS1dlUA2ycyrTXolGFpMkxCr84F4auhCTDuis6yjDkMow
avlA5kFRR94uKtWln+Hf1qJEx9IkgTOKRFFDDV43zjcFTUNVMhlTd/Y5i4xxT117vsBEod27Ex1c
hI39BkZ9/nLi+dZBBqyyqA5pVSa36Ux1ioJvxaekPJyTFlm7pjHhowJNhr6+Xr/CqQVsR3MVLbtf
f/q2u3rN+PfooGIu4Do74M64SSchXT4dkG8xHupkUUxVWcJuD87zLYlimJdOjlAm2nmxOSlTr9fM
N7oiDLkfxTms2p/YN7Q43/ZhOCsdQITzdsA4U7dpR5buMjJNmDraGMtLK7SDsg5utAWb4zbiyrJr
W0mB4+k89Ok2sRdXYDBO9O4DU89Db1JHrBiD+bFxIwSNViwjHriXKL5BSzoSenkHEtIaWju1lTjP
tdvH6Jyqip/vcHFns+RJXQm2MUW33WBsyl7gOMv/doaQccyfia47jY8SENDXMz5O3nRszauSbX5R
0ky+pSN6Tymw4EUJMtPp1I1YC7DME2Ks1H1YeZsBbjMGhWWJ3fdi5BBW46s6jCQZywAiQITTpMuq
dEQaZwcfImZT/qNyCpbiO2tGZF74wzF9/gAlG/7G7VXU3yXSqIILaxRp+ozD6DMG/1UocRS5oxiO
iRwMw/vve5qARzTntEZ3lhu5qBtcs2a4RERQluHguV80hbGC9JkBmBb0YOo6IggeMekh3VOA1998
htFy29dC0/BAK6wcMIAL1KGQrPIShcyTB13vhsSzhHpXT8L95jHQ0MjMPyFb9j2ADb/XlDMRdZ1f
pIhXBlw3HhcHeDzJXhdCNt6X+l1yv7yOPdoi/45jWiO4TIqX2+TOa4i1y2wD+C2+nPhmtsJpbCHO
o5vpvmiKoXA9BLbJkTc9CTJxT+WW6WzyDm/bRkYnAOXWfB9QpUfpJAV7uWehpsdpg7uaaGOY5NnQ
ieKgTOCNNhCs+gYvMQrA8c8AX6apORlSapK9wIrANEv9M9vv03kkvrmc4lVazzSug2gGE84Le2po
/CMFIS6bTr1j3xmzarP5arV1AH6WvWgLuDd5IEotpZFfaHLH1zLujspuDqBbTGI0ZpivmovaPqtU
FV01VpoE//S9e0whOEiGpLm+aqA74DvOF680/PabZzMqVZNTxPOIdSN2Z5wcdPdMx54XAyTF96c4
wHvUUnh4wvk1iX/WjezrqO3GLu7LH5sDqVtssKa7MdlGwTJIvcIHXBYkzBnThRaUxzDIry6dAThX
dLPbMRs54m4bzOxjyIYJksslmhqPeq+3rxOlYlKDW9HC3r6Fa7s4bbaB1W+29SrkrvVyvWEfH8pl
5PXO11CHAmEJpQ97s28teFucp6EZ0V2/mhbfV7nZ33g9A8oCbkrwTVVhyH3WaX32Q/Axb+IY7Bdv
RAjSGn4fHNqeKrEM/b9ISQrdbHTwNTXI5nsKtIZRop+y4IPwpBH3hD/RDBnX9fmlJbEvxno0n6jM
eki/JxePkVKPOYDcZTWay54fsQaJnhg2LvyhnwrqTP88Ek9u5ECUGxx511B1W5DfRq1DVUjdFxvV
hPD981sHrcDIdqyyozy4BbGvdRXhuvRRWXnpJezJHX600NUdIOzNdnI5U8tn/vgswW2i2PYYGpJv
ZAqLbhaldaiZyWBvYpojBK7bhxkmtE77GGPl0+dbSGrYPOBvtYBWHL5wAKOMwWuVsnjnEEfTieS8
knZSdIoagoS0vu7X5Y4O5a4ybfRbTBwYfVzdugt5zGpe51VdVizGw/cnoGos/XBaTRZVbeJZyQJi
E7bFA/Ftra37cEnLJ9bFTjINh6ecyzYjy6SQoF1fWqLiWWL9ebRcRidZbJfdIAcDxydhm3II/mAD
QZB/diboDwj294tWZ/l8jk3z+g4mVq4Rt7b39xzsn3bxYQsrB3zZb2LPU/Yy1kITsV3pc0hsiGib
/uWt0QW/SYK++wkyoDNfAzQi0MNGU+aPJkaF897nxWDfyvYp19LO3aUmNhwbxFDn/eB6BzDkgamy
4zGlnfwQa8c8soy9QGgbAyeSUFhzmTVOloiXOiX34sxt2h4GEe49umY6rdmqZBwfhUC07Z0Joni4
H3ilaBFO4I2XOLN5fbcNFbZJVeI+3ODCH4X5NPaHjNeCM8pb0/KiUa0KJaywx/6NtCAJH7bYhpSw
pU1ELv1NbjvH38RJ7agmK6oJhUcA/AsJC0UuayKw8891rOMK3L60Vz+e4Twse4uPm0MEPcw3ezw8
q2OMdv+kOSAup8SKVtZneZ7zftYjtIenxkHQLh6TwQnwmFrGAIb1aVlZuBAcKFIISIO43HRYVD5T
PXOM3hptTotIE3WuojFh8iw/FHs87nU0+ww/xNzu6L5whxiFr689wHBywx84VgADTzHZNOph5bT5
i54WgiiToX3SafePhQgDcZEHviu+LTZv/u1EcIoUP1Yqa7hpUTRCEkWNTNKN5nEDhDTqjNwMao10
+LhGTM4nASG84QtJvlIgpDtU5BurdcOAeAJQhEJT2yLbbEY0XGK4XWyz9y2obw53VNcdmAo8Ytro
8zM4BE9liaJj0JFPJc3MrEfaa6Nz7b1iTc52QnU7ssbAR2DN9GnJ/gI9iCF/liYIXwxELb41KXye
Ppa3FZt6FzbrMP9Uvsff9I/ypyMvWwZzXrXkIH94wZS/GSKz2jF+Z51j65pATHzMnq5jmnjaIk/y
3wMlVPNxqPwKdFojquV2G846mXPy+eMnShlvp5d5EjBIuK5T7AVBr1bZvouA8iRBKnwjrYCdAYoi
GA+7jhWnJ3YGBnK3CndjlJRM6ug6k/5KBy1CCSuN/HCVD3wGn+u+Spl0tyvh8bQob3HEdSNmtycq
Ob60SKt3BBIfXG2+ETYqGZQeFlT6RO8TXfimVGcEsEudBZcVoP4TV3Y+9aCPDyLVItQkKiCWFlZd
6aSPa29cWxxA81Ucca+CW58Q8ZHSyeEmLoZldVmVONA5v0dU3q6fy+UWNTS5azOFVgrSdCOQ9nMh
/8pRFc+GmeK0oV+FhHGf7BDdDqGDBlP3tFMFHNE+guzIEb5ujfMV127vwlYS5REBflSrcYdBBLeZ
b+1it1dBjVnirHzEMSmZt4a06ag+t2p6yz7U33QV31e3CT/NoT6VwUCI3sQ18xGbIEc2LkjFfZms
jgzH049gYCgP3bUqCZHJBMAOrYawYrSIXvLnYPdGYERypEPyppeQ8BvNCfxNzhVfnVewWEo3ZnZT
tz8HUMWFzDJFh390L8bhjZ6REdkMJSFs16wmYvpJ7o3sjyQLMwtMaAfKWt3TT8E2QtctNuKX9U+n
Plr/g9qqQnVOQk2rudpKZUt4dq5QOEVoKU3FBZYNmoee10bR21QAjEYn0B0TU7CXZRQBkjsFbd7h
fBhnamoxSkyVchkVs/lwwfPyW0QlMdoj7rpx/wA6msY56rY7CxfLXdIfDtn08LZeBPDfEP2UFaeu
HaTyTUN9bE6yyWbdD2UAZCVdFkukOaKgdCM9gBhcznA5fTfZVBtDl1y7X8hln9KJWWj8nSURiHAV
CzB+3DVPgeUPKel79XjKWYq19wTPXT+HbScqOgZDi+GLNM9S5o4egsmCswQB6sWAW6YLa7WljNsm
Z3UHXysBFY2AsGpBTmQCUzsB7KKQhyMM64cOTye2Et4QlggyWU9DGINmVSlJZfeEsTBNdkCGgu73
QHRG0RLPhYlLgTXRon8LxPIG+MOprD25caop1WvWIEVVVMsmmwWZW6CRBPW65RKZ7gAkaYrt3q2r
+p6KOqZWkXrxyWE424QMCebnC59JlLjBmJXWPnyQkucMfYah1n+fYz9CzNeH9OGuCWfkPFXoRVWL
G34GMK4kS+uYfaUwI7AlWKpiqxRqtP5LKkWbbjL0W/8l2CHzPqvv+xGp4sUrw1UHZg8uCpl4Ep4g
lb1JaMw/QUrD4w1sIlISQF9642yJk8csFTOIi8Mm0Q68QMS6dxF4wbWAIwbveOY/Whjm/6/oEVxR
EaYJdPS2zSDZXOvdL3mX0KPaL6/bmSZl/ooHKXOi7IPEf5QVnOwJDgRHAjr6xYD8Xckc5KGP3Bwh
XMf7gM1buvI2VMBEQ4mTP2pcCLG9nat3xRykEvC8wzQDWiJsEC0zHOm48Uxq+fIZ5P8vM2Y+NR+R
hUUZMT0THqPBxs0QOwb2JNdbHllVYWUAcBXruuPdUnJRM3uZPfus25g4VGQYvul9IVgNigrrqXd3
jx3bu9m+aBdVINB/PDxXtLnEiJvLazLhFE4R8/UaC5TEDmoBkGZuC3MVoiNxhttSGdssrEbhLATk
WQXysHhD9L01qGwUwvVLYDcXwNr96+iuS5Dm7peNw103gWc4NXNZXxBMAr+mMMl/jz23jo6SSp4p
fKckqlVadzazpfcDEeBJemoz0pefYuy0I+ceTbAa10pQp64i6p94CRHBqQzW79FN3rnf6tEOeb1H
lnLHc0bvgo67Va0mvTT9Dw0VIN84g/Ts97FAEBG+XX/9UDBD+efd4B4yizMkIGmc6iihJDmH/UfA
E8pMvDFlHEBKrU2c4a3vdflRnd4mue27jkmZFuDK99HuvD0pDZOwzMu21/vFrL2+Phy0X3Vq5EFz
8ai4qQG6SNfouRsjE2oXxlX07DKyWq7kSQT0lMX29JBtP3gpnh0dA4WJ1pQI8Msn2AJ1kuQ0L101
e406hhMUql15n4GMbino8zsCALE09l4qlMDb22v2Ju5rjgHpmPuIdCV1Z68zF1ssS1AvkzGNDJQO
3nWxocW7m3W3lS5UoxuvvWMErKmA+VART0HtrAmUPx/ZVXer7vxSxtTntPkx3V2nM3Ml5stjdcSR
AgKgJNG0/iXKvKGf6cC+5vw49NTCQeGxhWwW/cvDEz7aB8l8HiVId/YOBLTs4Z/zMtrbIXziufHR
aACrUc46sq1LcmpQNOJHmE51IkLaNdv3uuVtHw4dyoCn5o3q3mlX7c1xLUCN30e+yU6niQ+FWDXy
e/DspN/He1yMhi0Zb7oaqvLY4rQS09I0ETJKcJLNuUEstaheeINWJI7CGtEW/k/tc6xbHqayhMwM
hherMgOfOOhhtHO/0SQ4e+ZL0r/lYM+SCG4nmIkwKhXGJBxZ4ugAWSTwVegn8F1KOexH84+qQTki
0Sp9VDBxR3gCAz3wE1qBIz6lmMpYIROyKFsx9RcsoaIECgXPMogeZIOxO5dAg5p8ZzmcS7oG7KWb
qSF96le22+MPSIo9FpDxxqiIjvDd5yKibeUOdPs/rJgHmHPQRCFJ7NEv7+seu76PC0B55szvqW6s
hxiVBef5xdRdbA4ki5w6p/yUHQlLlYmAOO5DXPaiNaHLkeVqq4npEguDjHRhiFmZdmJFG4wT3sTE
V++pr4cX6TzRuVyp6TyswGJY28t+kwLpo0HTN/DpWdAWtIoeFa3lZPfn9ZrnAp7mrQsXFbRxUcxn
SuJdDVfQ+zBiohOEFDqvoEgH0/lS33IDN37mpTEU8wQ4w5mMMUWqAHuWZURK/XVPKef8m3FEeDZc
lKuNadlV73gEgKkCupWpUJTXCgDf99vVDK655sHTvJN5mVDprkif4ypN62pugKIZkI6SYS/9X8qN
npv3w8bVcHe+Oyhkjxq+nTrlcWs/x3ormmmeBaNMzFL54w8T21C/PgVRUGEY5ACYnAx429RJvEIn
lCwV7c1CLb+do9qiSKk+DvV1sRIcPf/Y0ARDAxMTZVfmKHVf8cBwBgGtYhfcNoAfpgXjkrWi/OuH
LvHdPYdR9QRqWD0FC3MdrgsKzaBtisHZsPhcL54KvNAKDMCxsL26Gd107gwclO+j+3Mr4ZuvfQAZ
9lxIYP8WgAmdV/CqVTU6uUsQhKnUQlySCT9Yf/W/Va/PIto06pa+kMyH1s1I7rpM7NtcnD4quUaU
1gqeasK2UJ5Qqe3vHA90YTRFOHz5lt5oUUIDl9VYxyb59fgVzuWbog7vyxDNIdZaSY79E6o3hHXO
EMvwqnNQehaWXgMMt7QbVCGUMXQ62Ny2Yrd9XzP33sCViBnwZnbNd6DbvDawh8SYPectQ8ZT3xlJ
c+Wk0WYwRJjs1bkWsMdkpLkCkKbn9vVxqMcOWueuWhK+DIeLk8GIdvV+ZzsFtLMH5MvSfZvfHZBH
0aOKLzF8savqX+mNSlG7IOge2jdJa0IvjsUrAUs48LwFZYo0xMnDhK7cr7LiiQUPLTERvhg8rkg5
2azHWHsMvxrqFFaexTakHgJ+4NQZcc/xjFL8grNV1YskwnAqpZ1Vww7rKA4jL8ep2D8tE12hgOHi
n31mwIB7k64otImoHj71zM7OUiBOqGeL9Z8mJ1WgKPsZ9S49SuzK0q05ezEJkrSa7ffM+UIG+oHr
sZiRp/B4WBFzDlqu7aYcQxbVicF+azKm18SdZN6zBGMcTRUhsBsOxNCCCquCKgGK5k/corndgAl9
3eVot6TPBONA+79cUVgNocp/MhFbT2k0uQbVOwAAOuC7RVVGAgcjWF+qcJV0qp3N3e9nYVsQ89+X
1sU7O9qhl5pOIrXunCYNHIlTA/4Db9yw239Ez1VaxMJ5NDlwwXHGKNkcwd/lSg1lcEbKP/girXFM
rkrACwqngcqHQq8w6jXDMZjNU17777DIFHuSooJtSSg2uVhaYH1NCiGesBcEMxafrCnNL2Ot9PA3
BTlxXOpb6wbbiaPx9vdT4INqq7AAKnDFU3x7MxmIIeLxSYsypSq6K2jFRtzsCbgHb5V8EWauQBM4
XYBHaRHeosmV/CaxsgFC51WrOJDuD8QpmfKfoLv0s8gjqNxkT5GBbx/oUUb0MaR4YW68iwOt4SWR
0c/T1BNm3GA7WGLqzce96uUR4XUx8f+lVI8V/TD/HltSO/gW70I9fVb4+3jkiGI0cWO7N9o4ElME
isRV1UifDcycpE+ByO9NIspJKGGpZw97WgpLhgJ9FAoO7mEhN995HLW3KKXHSSpzwAiAe3NnDjmd
PCjx8L9JQww6aNFyY07b9mpfN2HCuTqYtBJfG5GL1xC/6qjO6vMCt+8yUaW36JHeta98xr3+J2el
zGJr1zPdoPLhfroD7dAiME6URNceZDDiIfGgdz5OsQFgd6bk89YQqQmjbe0wc6UsJrMG0QAthETb
Dx8J/LDVIl4Y8kk1ATLmNmJ6YBxPtvpeKLSj34pPmZbMyxwsnNvHjMg8cGoQ3bRa6BZqaoNxNgVb
FbHqSti04QeffdxlPvbHU72m3dsEnJyTGnbEKXzo/uN0CvQS3C46WBUh3MEw4x5L/7qPbtTO2IP+
AmA8gVr3gnNTTYx9IO/Rz6fTGd/0UzzJCYUQa35stu5yk7+BRCfyrtSahdTqi0FN6BSsGJCyGpcS
rT4XzJJwj6HPFMuQt39faxV62noFNFRb9neMAhWJVf0mNybVvoDlU8RO/9pXSYNKmUxTKi8pHklW
73QzDFSR2uft65OQAxsNO/u5sdp3SDJ1YTIoDMjrYG7ydXB8fpi/iBZCmMkmWQ+U9OFAsxMBrb8I
ySwy7STPmxnxK0xLjN+4aGTO3xpSs8SiHaf9xctVMUoX0h3svQVGKs4RchLkm3d1BWk8h5/n70iO
Eb4H3AzAau5qgW3BKs3uPlzui6A9U0FRLgCTrUK3JNgKkmpKIxDeq7JRwLNfMfgD4v9Bg/JMr4r4
AL14XYT0jWPOGYLp9s60HmVFLU+MKwKfq/L2DI4JVH3gwALhDd8Xkdbq1CL6gtJK2zaxhM4gHuEc
IjxbHOTIYcZ7McP6iGOYfkMxYlRV/AYvv0slDOtFv6BZMmu6wDpznopG2AtWv9D+AkOUP7LX7IXE
W81Zangmi/GRmUrUm7SjAMsa71hycEW4NXchXvn8rV10DQVgv2hzllvWxNQhx+Qsm5+yArIMfrjA
BX0NsYnziV+O26CpIzczRMhQZ4rxg2YO7/cl49/dBAFPE1fsoLVNFL9qzd6vwuT6cI6gtCXQRJVo
PanO4GhMdUBlunsDEXiJlHB9hiWAmto8AOP5SJ2mHfMKzhoZUmYEdliQWxmbwFaN3LI7V7wBZb36
7rKFn/TgboRNcmOQOTK+50euacPLAbE49T8o9lYMif/54aMqQlN2V6SxM1mWx3B3Eb6EuUo/+T4/
RzAOr3qlmR1iDs4Kjudg748Lf57xMggu07wog5I/G+1uiMOvPp4Jz2/FRuxp+vCA3vFbbUe+zRfA
MptAY9W+kHTMZnQjVv66UPk0wlFNZSxCmLd9y9VS63fIuaMM0WmhWHeXEXVxTMOd5e862e3YWCV8
5C0T5qkt93dUCEfdU4TKZClEKd5Xs2ce10E80wl4aEwGJHQQBtsqXjgrksyBlwM4Wb/5g9ffl6jf
1dtlcK8tWXTKVdi7ih/eAyWL/9bBFi3rBFpfP2S+jFSA1BUSN5w71jjYnahsnNljIf0ASJ5GGfu5
JCyEt83lLEuJrFmA5j1hMkv+4VMxV6RyaAGPGs43ELHLtzR/3z9f8MRI99WgA4YT9Dy7QzdGn0/X
X2jAqCac26RptfY3WPxfwyfMNEXhceidBeRa2h0AwtY3+RzaGAeiOpRG/Y3xnNPiDkbfjjm0u4Lc
LzHERUHTGwiBoUAXkGfRxT8bLaIZjl8wgwA1/R8Pb3drKMLHuj6oY4SdGW3davsznb40a7+fVCAz
k4tFzFi8ozBodB5XV5FxW83EYi7ORpce7m8uHUwsllK6EVchhuGh2VT3Ct8hBuJ9njI6FuO4WCPA
pkEasKTI2SrqTLanGBxhcUymnRuRztGmftmzXP7vszTiwf0otQGlxkuZ4BMjXjGVi5Eb8/m6QnLv
FVLyA/NNGXejYS21e+HgnLjZW4q8Iaip3Z2QbXzBCHClh7weWIbFY/FdTsPcRBBdQfDUgghns/aT
/jmRuKOygr6h8w4TcCcnAlsTzIDlJy3wezsDgnyLkN1y9t4VvYcLzm1ZtJWKn+SW7mDQFK8qL2Hz
yGDCz7zAAFwKcFmieLlIfTWr/vPO0ylQ6VTiOFue9Qn3IsQ8YMbxfzCobsTs17cuaO2PSyGMMCYK
chXVuT6kjfYNP2e+Pypu50U8igOomoUv6FsQIH3aZgGZ5JGMa+IwbNLLBkXAMnAc01D4YRK1qYs8
V+Hpf+Tz4TFZVzPSUm+1qZUOItgS2oMTBHuwCgjrui/bu1PTumC0wPw/df5p3IyFnJPHS4UaPIXU
cVy8PpBI9bp0IY4NB3SzEWYQ3N0pxtJs3rVOhAuVImAH12EXf3JxjAyBclpxZJ1aPNMym29GGPHU
lPXU0LOpFX9tqb+2vRMiXuDgrnL9BKHf6tuTDX3Mw3MsX5T6tbZ+cFHq4ZqRYbyfCvJLeUcg0mVH
2y0Elk2wFPPMPWKI6cSROojicDgn/zh69WVSPJiEnhLvSiB/FR15LsLZGn6F0GbMiXbuH5Dm2znn
h60fyX4xxJhQnZvKX92olD+uVuXQRCnU68O7swjO43pQCFPWNIGszkCO6bS2hbTIbqaukEq09dAo
1s1R4w3hpjSMG1M43wSdIGpu1Pp27aCQSxWYt6UQDEKc/j9Wbbpws5HPPbAZJCSR0d3F7bxXZJYx
5/S0zbWovHoAXg5EnLVYkPqyLCZ3YI+ycz9FIYqEBHhfV1uZ74SkCdLOnI+kkESZNRj4OlA4DqoX
o3EixrqzxAKV1tH02sFK6jsbcHjnOWwgd51fkMer0SVYv72/Xnh9kYnWaiOYZ95FGuPbb9xPPZmp
+s371mKZatDSXQAePKRZrfWLMtmNWxRb6ebiPAGCD/E5X49oIimAlXrxvdEApswKaE6rId8vkf9Y
f/PU5sM1zXAqJcwXe7SGYOOca5q/E3gAokkUAUigzSlRITuFkGTt+9BGtV+JINI0WWddccTcEyzX
868sKW06upvG76qVmtIDf5vYooUUcHBpRLgyt/qiH2HmBpw/gTmT1jj8kkcVa2njfDPPRJ0YJEdQ
tlnHIlhiwlNYOY8Ph8hXrgu+UiwJSbruxWVm1pU1zJHicVlox9Ck0nyCA0O125Ru+lCIqZxEdEKD
BLaITde9o/AEGucDhuSTsdQBJDSYl1nHsq34IDoPManpyCSSTE5XrbJv0jxVRW3jVmF3+69cN8ve
7No7Ixnjwn7pVK249esHit+RRaiMJ7TOSekpmVhN4fB/kbsK3KHKpLgHDnL+pdPH4Jt9NA1y9yIa
hK+aUupNHZ/VVSbbkUkS3o1A1Yag83/k9Qjy4HeXw9nM64ALsQ+QlL0V5bXkjhMJ5RpidKp8aucG
T4QTmCGDOYYPv0e5Y1BtvHwkwXhUDTSPmejCUXBCJf7jMw2RgMmjASU99e6Ev38GHM2UQZy7UmyX
3byou5PmAvNVOilCDg6ibvIzYAisyAH/EvSf6dNjeJiDVtXz/bc86OsXakOtEyaDiw0slJSxny/8
5DZE219upE5EeES5LWgVi2YipkEJovZNujVJGrtz8v0gpzshaep5fOjTCkvnzahkQvlYeSSeFdOj
slo8TgzvfFokbM4lDs3456xlQyUiVPH+4vV5USzVuPhA6elxTB8w5WZarfPG291o/LzsyJ+XGviN
SjmamoAHC8/2KBkyjQE/GQ6CIJKTQRUZF6Jx65XJnpC0e5/gmiSnd8lQOMjhEuUBeaMevQABIqsW
e2JxJ+atEtBAtxZBG4oM11Mf4g60HGfqKfYEWHEip5qrEX8UgyVt1zwQuMwzmylUTvPcSCUzNUiT
5ug/NdvGEJTvTjsFT3HZQLxE089D2KHL+J1uYGpZ7fIdc4/ouRXmVTjkcJszC3GYwozw0a7dpdfI
YY9nveivWj2fVlzRwxVPk2jjdzwUFYQnMFWcjSjELwO5aLK2yZqDnHRzf87loVcChrEAbYVZEmlu
DGIAyzdwybTfXUoPcqt5KshS5aHI/edVxkrmE6tByjMIbdQZwD3pfBrRFeFqTkHIKTOAvyDSupf2
ZDXkzwlcKZa/SnPtGgKyxpQrgjmqt+gU602KcIy1p/AphAGStgowkhkrnrNtl3SCtaHpNbZHN+kE
0Beg8nFnFSDrXDTWGCjMaxmj2M7TaZCdB6VmPWl4jmUNIKiA6KBgjgFSz8NiQGPPqI4tKhbsZyQW
xRK9Goke8qvQ0TisUB8LoJPHVKw17gROJvRwU9rdIbk4XfucpF2+0i17xqLp+1XAT1AcnrURM+4D
cKyFYO0JplNoVsVFuFfOMumOUO+R7epmKA4SJBqUOiwQaVfkvnqKZ1uzYG6ASdnFkU5rctI5MH93
3bZ5uSIsyfi34kQxRhE/Mma7ZDe0brvcVh6qCHpeGZ8PRfaOMqqly6MMssNDUnYirxycHxwjyOfp
umTuwukfq7bHTHz7/fK5kpfz/pEy1nKzE3eg0MIPOxb/FZXXlDHkl/unHf1k2h+95CHaGIeSdO9H
vHaA1wKqZQFGNRXUsEgKB8IgCCHGZRPo2/mnRAHFCGvhEE/sOgd88abB5hoOIDa1RxvT3qfWAymt
p1ZVoyGeTUktMq7nxqJoSc1OaEL44X0kTlOq62pHGxzGOFlJkukHVh4OUyPizZNirIwxvXLcwkqx
MKfxC6Po5MAq6awVrfg3Xn4z5h17F2ubDvRMrGug/7e81xFD6VmIa0pPLNCQ3h+IUrO48tGZqTAb
xsdM6kO4wk3hg6lmQVNWk9spkJrRhGRCz3Cbzw5fZbEShDnlffs5QmC4nrZ66XaagKqZFV8GB52i
QymcKPuUSvXGzTlACZZ6EhmIQUyg2atd4ev7B0Jf/j08u0AwVPYs530JChHJ30LS6rOzIGfC/YXk
eRF3qxy3ftScsB8ToAOI+fcv/4sLKHh+sZdVCRj1nRLJrRrRDxY7B5Re6UXD9RK3j73Qv5Y18MVk
d5wveAHoIDFtD2ZWsoul2fc8GT7xMUmFGELbHimFSqtnLlAycA1QthAPCahQ6cTGCvdwHblCRcmZ
017kG7iCQUGbnaXA2OTWiIKSOqIoWdRBHhoWJp99j+m94OOSQfovFcx2p/5g0G4SC3oe0Ic/iDro
kBKqk9tlw86caBAJoCAf7G3wmdWgukd6poDIIjvWZzG0XGxTJmokc+GKusDSJjHkFXrQyVx2Kv8q
95ZHvpGyHD8LcT1SzmuIhOkO7HVuoiEy1RSoHSdnQ7vWOGaWq2TZD+18hBbYwY0+aC5MSzpsW7xx
EXys3V82oHsvj5w3pRKNLdXu9bUUanDu63Zs8KKA6453nv23zFlbAq9thaC5J8O0z1LIFrH3kMKz
GB9onYb7T4NIQOxRychKgckPNXsKqb42KZu20gNk6b6NyCzSdSYYHn0eYnzYm+qNgWQ9trZu+ZXE
dif2wyrDJUWoxEZFakisQ+ikjatYlSyUD4PgQ82GJA3HqRoQDLvPl2OyIGbnv5Apxs8qOAHbCPgA
1UfC9APG1VsLM4iWHDUbqmT21oBYSWfRguD6mP7z8XabFoFovG8xclMim7k4wCSl/y9+OBD2Zb17
EDSaTLWaffbBASHp94WBMHW+ryEbd0gvGog05qtXvwX7jCb1iy4cT7A1oyn+2hehGghs+VDPOVOp
cDKqo+sl/mILtr556eyrwoIlmZazTu4yxJWFfkU9A67d5xLdcEvn2aA7xmL8xP7PwAzH0gBrfcwK
IwYt13doYMxy6oWU3zacKzcGJS3EOvJ47IKiPtSLhs01i0ubWLObSZ5DYfxMKlSbaQYeNIymVaIP
lNNjGUMKGK7jONKQqrpYd4O7IYlfB9U1lBHyE5/5VtrWOosAsoLBw7XaCI3GZpOb8XRr2F1/whSH
bDFuakRVW09q45lWUPnhAT5yTDzfqNmnmgR0k91IQ+R+cfwOB+vIc+Xom1A9tJ2YF/jgrHmLhPOA
zRvew6+kRWaXOn0pKbCIQfSNbhXR0YKidrYp4GetROmHoicm7D6CviQdgoc0J315taR0BAdYg+r3
65LWL3IlLnKTgDgBJ+6IWKKggMBKwbBKW7Oo8prHfLLzSUuGw8FXXaW08oYE04Ei3O4DSTqsn3kh
nLNN2zYFbhntZJaRCOiW3JfliUHA7Ghmf9J4JRlI1aQ3QUltWtZQQdo0Gk8gMr1enPPbS291QV+i
Q+ezrdM23c02ZRV2lifvXq2HURVAmIvqDVTTkaemlDLCWhc/ZYGpr+ToYXeuEc9MQjBwHO1/oCxv
2L67gUFuxd+yUpnCoXKMeSeCajPlgARCIuPYod9VyA2kgXgHBh/ZgCIVxk2mELLlURtziCkBMWE9
Jqc59ziiYfs/EKa7NRiRVR6FfJN3UQor9R6KX63HOrcs+VGKeGk6YH3A2E394XBKZbM9JawEWLNg
rOFPoD1Rf/CWMigbn8Tm6yzESjK7ZxuuVOTV7ld/vGGQe7HWW/WZ3xF7QL5slwSW7CAyTQvUqzh3
ImjOePARGURsdp5D11bTwOMb+z8OC3AtIq9xbT6BSw/E8fAf525FHYwv0N+4SUfPP6XJYYPwYSXQ
Llpej0XsCP9T/ZY3Fnc14EJ+k3+Vme8IZwvnkCY38SfkXdVIZPLspIqYo6vHvLuUEFKKHQ8m8npW
lU9bEAKdgDDViILWbsBRVAhJHFc8QEGF4afXEWjVU6212zUEbHP+f04gMJFDN3ozE85OnyMjGYAf
TZrc64vdDZC1LgNMV7iB7VmCbxJl3kU2rEaYQNfF7SYIzsQYHHRawQc01UM/mI8ZqOF+yuyZcDJz
9YmuhcpK8nDTBR2bkB2l9v6fJgU5QhdyZy18wyWjJbcSXL1RAc8nfmws+R/9/E5V4ImjiLwVc+4Q
+m4NWJbGyodapZxmZ1wL4u3hfmXO/8ZfW2lyudy0ZJWTeiUeYeT3jFibDALwZZUx8yT7nLuUKyy9
GTTb3ZdwU4QEVKl31/U269aB0l5o6LO+Z8PJFeA2ty06hrLTkup5rqf1fdAYKuIQVcOR/JsOpSim
wwfZjELn6jY144jA6Q/pb3BA9J3ki2QaGATOauPiBAd6bz8Y//VFiBepLLppoC9v6SsmItgshezB
NyBKV9k1O77QowCJc4hw6i6okFEn5YbVAh6ueVi6uOyOu8f/I6cpU6bsRJefq/Gbfe09e5xvND18
bdnTOu1avzd0KdVWoIOV5TfJxQLvhgJMqOTRzI5q7/Vpgk/ngfiUNl3X8santo5YY/gtZZfgQoq6
05FNS8zpM52qKpHJq+PO/LfgHddbGYLTzgdFWpn43EoS7tx4GXcySCvDiZEiaWJy3V4hXh11rsTP
XJzNuFTlMxqcQxmM7R/dHjPteEReB1Gl7CKptvENCKcy8/178Q8yltJQFCoez3P0eEGuR7Nxor0o
QOAKu56rQ5RiyW1H/ZyYjD4osvLBBkPfbzM5f4hbd/D0hBqUNC7SBj9lt2h7xddEdyrtCOaqWynu
CP1WgYFPv+gg71paYceZJdFatUF601lhHv8pOGOgLkZmTl7Em+d603NSL/79Z7U93hkBWDUlVGUO
1cnO9TEbq8cMbuANgMm08pM5qJ+9S6bIIFuWc1j89AyhaJePoJ7j4OZ9ExkRguOKEs7kmUkx5/Jj
HM8fXNuYrT0w+lNOmQDC309gJBWXnhSKA8pAVUmAAt93oR/kkvwXN5UQ8+lPwQwR0kj7Atgr+560
unL///GUfuiqbmAvmdCAH0EvsF3aQF6uFnJ1iQgDt63OTq9XOus1yGZbAM8uqTXzMon0f6KLBQkZ
N6joMb5RrbriC/m1y+JOyOJI5TN/mQjAgTTnWNfa166Dd7xK32zXANL2bLYNzYJ7sMiviuYOH7NF
EgfsuF0FxajVefl3RApL/EsarqDh51CqZXY+C8BTueTEk8UnqLZiTVO2SE5CPvDonYeNGgNhJoAc
+2JjHZoB3kCB9CENsauk8B67TU1JHhsIDBq+zQXnkJfnpakE61iq8xbrDn6rySRIDBzipmDwr3Ur
/0sWFz6p3Plc4uzbyLJK9XPK3ZGNTKlF8RqFzEH59vT/jkZn+oGPuB0w/q3NmE9QzeMoB8HGbKf+
Qmqa4dlPsuwjJUy/S2E2VVY4Hl+Us1jykuf0JTsqPVKn8Y9CPYZaV7HIbaGXQTGmO//6eEvvtxUX
zbwbmn/g1W0gQREklDIYU8VJoRVAL2pjdnmCEJrtbT/HyJI69YcGQM1MgrR+dL6mxMGYef9uMK+C
QDjM6rX1SWwt0zycoEB3wnyaG9g6fY+I9YJ4aPklwwX2qEHcWJfw03ER/lOb1k7EpCvF/aF43PxR
BhWCtquma3FXwXTTAS9ixjkuKhmq6As+W7mclFtb5eeXGrHg39g0c0oqs7NMKo5yKY5+sffToyFk
VlA7qpnQGYav55qMkNZrLGIe6oOjUWQwdSxT7tBqiA11mFQXSnq8xUSnPGgUYsAFf4Tsxkr5/yjP
7aelCCLF+Jg3HThMyfleMc3eJ1CSOXo5Qm0Aa55PbHijXpwmzaaYcnkp0Uw3PgC6d9/179Qo9c6W
1XHD+zsbMfL/gCt8L78WVc5QE9FvLKUdjtTnwbPDT28fzVELohvZ/KvGudmav93O7Iig5AILim65
qn0yKmKjFFTyQHHj2dnxEsvNphjmo/g++6N7/1Eb6Jox7GE8UTr/M55RSs4ZRShg21kSXpEARQsp
+JnOX05MyTn0J0pRgTJvfom6EuQojGFTzuc3T6vBAndhadrJanVcUyarabBeZ/3PFxpuyCEQ9TFu
SPa0E/8t1Pi++62aVrQ/sNdyV3xh9gsynZ2cBLVAG2o6wx8Z5kBr5Hv22aYmdAOv64/U9xHvg3Vu
hDEX3iQZ4WsyRPglUsTmlFuqqfpXzYRl5kGtEvTZNinV0dhgYLdF/GG9At+PcfWN3yfjGTs5GjEO
gtv8yGx4LIGV9vlFNIW6KQqkhh0sr78zwAidLkCYiJiWaJg19bQLKjuqgU3/jA7x5x2Uv3mpXZ8+
jN2c0c1i4KufEjjH2TBJ5zQ+/aU2d2qr5vZFXwo78RieQOqZvxzdhbGj/WOVkXatYPUbUqPfUcIq
hfAK5ItSgFbSnacXOLs/hl1OD6it6AGm/kok7NoMKrISNhxSyYrk5MFkTVPxYXycDecWmIEjzwEO
RS2gYtdrLetTIFVZjWvpS+SI6vnd8ThbDYvr/3R60eSVyZLgUy92FtCJiF9HBehaUkjkG+jbx0vX
mLOD7/N8GgqAxgDhNvXPNcNtfgUONIFjDwFJ31bDmHhN/EKB8ZCZm7WFjeN6kSsBaMg5BrACN4sa
zfz68Zw448rXNaJ918AWDasdIaEW+C/EaS4zinhNiCaWH+5L3ZcijRwTWb8+T4SHsC/c/uk+NqNk
+l9HcCJhL098FepBLlbmYDtNUcJyo7v+uB0b7k8Wsj9DKPE1n8Ux/LPBCC/2fepTYuNuYs4ha3ST
FUfb4eI4sznviewoj7jSvxaivFiGW1DAWnJwbTByF/wnq9sqgCI3eiqnHAQZ5lF1SSxZfwwYxqk/
IE7phM47q0MVL41+3kCtffaFsucRw9JOad6ZmVv81v1lVM9j24XCcKGfVvcTupqZZ4c6GDh4fowQ
QipdW8kGtOIUTU7vO0f6NVz8Lt7DUhzAw3ms9ywKj2Bkc0CeJAYNDB5oXMsnz0+GhW75pgDGNLGe
zTCaGAhtcyWTUWF2aWVliapfVnmGmYQmecN5EX9Xv2E4OylQDrK346h/P6zeym2hwQ0THRv5IzLE
L9rTTLKDfizuT0mUb7mvJ8PBOSOhJ46ThChkbSSPmIngqrkkoFxFIWeVC7uAxG0Qj4Fpc3rNixHR
lQ2zs3oVIZrCh8wiiwHOyKLH6TSSO9nHf2cyhx1XCr+Yaw/St1aqqgFRyOGsWrRvghPMYbLAz4Oa
xFcD9EJhx46qXje5tN73X9VPpwF1CRfN0BCdmF1lyPRwuZd+OFUbGJCWaH2RiqgwRBbn8EpMkGNB
EpL0DEP9pWVjs5XD6xLYIA2a4bPKp3I4aIHXxlXHz/Sur9S+W3Y3zs/nJIyNtNjoek9da3tqonpA
Q++DsT6yGic4Ijidk4IbGL4LjFcI/GXt/rv8O8PfjpOWvG3ZJQLeoqDXYnyFr+s4fsgxjQ/Es656
TxA4GtxUPlEsT+XttRmwriwOJv2jf7MCOG0QQEulcnOLZX9mFA3NORygsWXPZDVZW6cgLDD3pGL1
CsJ97bllDBnl7OGPpVW8ILud4daPdont0MZmfdszFJ4sjdbjeEaW+7vX9W4YaUQPk7AkfEHXFcXL
WrYkLZsumN3cwM8ILpIy5MNGVAIQNxf71UEN+661V5TVee4IkhC4EY90mSZUxoKjVNpc7hHsOVZA
SORPNIFd/FaMwAkbO7TsA0HHryp+tjPfv6ifkO7xriqnV+IKi9o5/jJs+EEnHyxdW1tQ39//uNb6
NHDJ72PYvZt1Rwn44z7AwMwdw3HpwfVsa6Wi9AVaeRpvlHPGoSNpfS3EV/k9jWJ0Wt3VEaOzZV5b
Ng0yjJaxQTbCnufaIPljPLR+ED+siSTOqt5Z80zsRyJSx9wItVNz411MyUTG2Zg9aC8RnZ+wK11M
v/PyBTbQyjDpCad1vaH6a8C0cGFpdTyMlfgm+KcHtNGwPZEzKyKzaAJ4xEBv1gQVJjka7IApE1Hy
7SrqMsi/N+J4oIz/6/jKCAQFtmoOJyPA0ACrsFsBeJ4HArKS7oaPVLJljXte3rzb1huopYqmCypt
hGxrQ7NqrLN4tEgWVwMf9PaN45rROdDSRQ37PpJeObmKZAbrFPG3SLTNALVRKiGqHDtcQrWk20uV
nNBHGgHMt/DyUDXkhABVSyToceeKMlSzWhJ2cYFdokyPk3cLhaaAV6ErC4jv+dOiZud5iJqNTgE2
WzBiaXxkKcvPFr/yo+ei4xiQAQU+1IkDzDFi7ugvnO1pJL/oazmjTzpfrDXu07up7px5F6V5bnq2
kqCLVGuN8ta4JmN0/m+ETLMNbmaN3A+DAyAJC48K3OGHCtTomEt5ehDhm2NR9kybkdvDwLDA9aCP
lDNo87xreYERkUxO58PfWNn3H0Vjrq+U5kJAjxPemje1tOQrA7MdgiFOXrK+raWZiq6lp9/phHPH
lnhhzpfPVKebN1hAs54ZHGKwWjzkO3SgIMYaN2r/AVpozeE335wHHih0VV3jGEqqeCrO+slWNfCh
LjObaHqp/tcWRbgfiYey0wmnmvxpi1wR61oRxD38GlHGAKw85FTzBqPpsKm21J+ITU+k+jQknOgR
8DiOQl2faKPQ6VQ3VINPOXQopdsRO/X8a1vbiD3AYVIkAep0H7Oa7Yj+zEtG2G2tfJYEPnLKtAFa
fZrbWfUpOjm3LkDJe0Ub0YpHNvgErwTeTeuciMXoEWaLhL1wufVBDb8ZEcT0t/ckfxnu5P7PHGMs
050W2z3mBC7tCMYEaTyL7jHUFqgujjL7GVxSTwNcxwnDjpXKaaK3TgviPI0eV8FVbHTj7yFZvc3W
Dk+NTxSSTPKB6SrUK3KevmbMJTudtl2qCkOztqhFjC/o7ATzOUjxWF6RXTAwryy6cAeZpSjUUOJG
dfzTwuo5SrXqrJrtzcP6UHedNOhWuszU5n63x93R1qZHlOsQipkPR1Fd2JangaWEMAxVkQ3heTgG
rPFRk+ljxb3uKcFYtfjxaQ9dWF5krQroZWrzeXhnP4WbaOxdKSiNsVRjKaT3iLRNaDzsOwIOBRgJ
9nQQlG4OFtk8coEXy+Vhe1sBiNlgiy7jGQgUOr3dbsE6m2OKcHMHOj0BU5vhUWQRzpRFbkRPIuu4
wVZ+KaslKzYRK1PRxBDglTCGUsp5gHpUi0C4+65ZRrzzfBSSAcMFsMID/IeGXgTMH1yYC+qWkmaV
MhGtJSofxtroPl4Zv5RIeBQDvp/JPzNCTZIaeNddvsnx3WYk4v/Wu5SrZAuSNX+gu17OZAjsGNSB
ETzo2eBgXNvOGSVtQCcGekEo5WFZBTlGmbeR2IDhp13V4APj1XoES2btTmVUCXkVAnvxfrmFGsCm
gJ35xvU3pHtVPT9LmtbAYkdKfc6MivoPak3kQIm4VwLbPI2Q8aa0wtM9kws3c/hpL2SlteVdH95p
htE745+C3sdn9E4/rQbVZ6HiQqQ8a1WvRhjP33IE8IFdidDcMcYwlL7aeS8qQdxQhirp+juo6vXZ
246oyJ9DQZ+OzdodGfEc8CaVklCjhFgRSEfBWPPfEWYX25tqyKlOEdhe6iR/W/prwBWeozArDaub
66dPTGf31blGpEq/rvNTqRuWkTQTYCbew2BnZRJCjwQaYk7K4hgkoB7ZDE+uxBQMm7nKgm3nCsDA
3DBt4RzOLOuOXiFltRwcJ18ZThICLLRuvDL5pGsFhMJzpLvTHaN+Bs3IGiQ9BeuJaudggrfOF7my
/SIvKaIny74g+LsutDoMSpi7hzASoFwb631J18gwo0OsLBdlpiP5APbLy/fuv84YN+IqKSJFJDqg
utL+YR1ighRx1GqvhrHQIbDXb8Ft3ZQAP72xFHAtInlOhDPhMvYuvyafILv4b2/uKb9gA/xrtPZ5
5QCK2nJ3Q0v804Ol0ceViHnnkDeD/qdFoS2zJvhXCl+RNpCcO3qtydp7ws3E2/H8zlQfDAxvLCSJ
TEcMtwY5QWiL/uoyyq7XJG9J+XIQWMltGUwyrfmSKv0kU+Jw7HM27UNij4cVJCBGou3h+Gz5dIBl
324Sw0f4BTfsYntm+VqKNUYnzVtujMfjukKlAKFvWyPkHsAUKh7UDc9PXDAxgfI9kIXSUVogUX7+
i49NnI7iyF1zCpWkVB1f5JM0SX8+scCCzKMfyENSnGfig8QEEzs8EmEVXIWiJO4cAB9vDYMrpoHK
QacNG837CWMxtRSay2gztu0OFUHTNLg1B5BFmwW3gxATkXNjnvqFXvq/q4FQ0lzeiL2ZO8CUSnwu
O98yuDb+Lmb09oumMikewQhc765vUxmu8S3cqXhLjVevQmJ7OUBsa/OZyTx5Osp8fvOZg1owpXrg
VJaOCW2c1JgtPKzQPqnRFEFLN0oKRfBhZGITyLG3E9j24x7A0bZf914w4X9zVX3XGvdTobZ6iFB6
QE98gQ0l1vVrIeBtoLKv2cL5A2U8TTISKMMz9nq1qKvZskaFQ2FS6vYnlYF0Yi6kJsTXf5y7+fSD
tXhswrcHV3Z18YC+yZVpuQeepb56Ms3/mnLVgKwAx3fYeNZcqiRcHwb7BH9ZPNVHnzEBThGXQIYt
0mdwvHOqGdqGyyMummneVGL9t027FprY0oV+rGREjOfC/QVxdSoq9mqUo5M24gAzvM7fmx0wEUq/
7dGLuHJfc6Al1OTEpYGTzjbXWY68t9CzDRL9Qg6QgiihS4QdmlH7y9NHoaqG3VOy/+4eyhMyUOoY
fp6zdbu+OsC2sKDkP8KxfFxsek6bP1M8+k8viUDJ5wGhvxmufWtC5lo+hbcXjmr0m4CvcNX8RA7s
szXlHLfgjbHX+bq8UOhCrP96CuS7WKUOnB8VMnluT00qh7GflSieJ4WjifO6anaSwS7vTbnEmIN1
GXnALVtmbNVRFQTqN0JfVXgYgqeJt41GEb29Rpb/NF1OR5VpV8FD9ZfZOIzYu+uQkhGxs+OeQys3
jOjE5DOag0//9SG5UQg3HMluQLph417nrK5qd0tt4VAOXoI3zq76bPyn555fPFR55HHMMk/2i7zT
zZg7oR1clyDswSZi0bplqLLD30UiZY34mUPIr88dxFIvbsRsQyzwJBCWa/Z9cSyX2e3VTYnRDx0N
G8xb2xDJG4evJ7vcMxbDF9srqZr0Z0xLXxQSmYmBPPULFIwi8xebCsl/szHdkvBZ0oiqzsOrzZcM
ooDtW8DKxMcl96tA9wZupoz/JW0ECxX2kU6odmre67DeEmuSwg3zCdLpQGKNKI72InkwmTtRxy1e
4pgH0aNYizoZaXQjOH8jE+RnhrnasYr5DCtz+UfpYlxxYXsvGr6Wnn9iaxL+8v+2Ak/9Yb6Hg2/F
iK5p2K7V0lCMLTZ4xQEwD8oa3DLmraxaMmU+qE2l3H+wkSc+KomRR46MqOdKPFv2SLlQVb40jhUG
kusJwUYXezGVbmPI5xAcZjAsHXG+ytkUhCgF0c+RV82wa1gNDKpJU5xAvDsIvhsvbrcLBKbvJIcv
s+1HE8Jyl4zkp+dGEqazG6HPaDvnowPHxGOyqjelvIR5o6BjyrQLOrgpnkhcHLWnVyylFQo8WAU5
o/ljZaDA8gCYvFxn8MbaljJsocnCWcFduPbEmSYZd4nYFHQwOK8VXlKkBIAETUBrr7uZYCShTULu
kKhIAe509tao/ML3FOklBjxkExoik0MnE8bKMWI3lLV3mqRUMM2SnSK/dgV29zjXoe8hSHDLN9z0
3wBjY9VnITowuVBH9hSmrRtmouwfhbrmlgOFleXfwWi4hvYAqGxn3zbayem80cCXJk4a0SeqDX+Y
gooAQNFVwJYbDInAN5Gq1UlZ59GsxvYRnQ3S5PSyC/koIpR75ngWfElbLwbgoYqVjN3Whi28yYCf
m3bO19p+WAXyPomel9JIlLlz8W9XPZsXR/SypZQ8plR5/ndMUPl/kiseOU8Jwos5fMzn7I7cFKJa
s2A1Igcaf1UkkoUXJ+Rt01rQ08wqAucAkHnYQte0hnkceUxX2xDZVzwvn5fA64H7gDp7wziPsYRI
YDT0y0h+JNv0+4G5EVSzZz3CSeiBZt9nfD01rhnX1B/LPNEodawEDg6bC7rlD/QTRfn0ro4Dparz
POzboWjcfsl42eGY+wS4xBkY17DcXyxnF3GI5EwlwDOgqNVXwDo4H9e6D1I8v5mxc19vyUnZzDjo
NnQJAJLiRHc5OWtjiIGNczruLXVw1BI1Csoo/AXbX/CV2QTn4jHxPWmJD/FGOf4+9xbymJ9aA0Lc
WDi9m0aEYwy4EY71Jbo2+8x+ISwnjkHpe6pCbE88269/vnCAvVIvf0eQJtnyGrL091eTr0iN4Bbu
kRTlhHtURiR69DLUgE72rcVwEH/S+veFVUM2Ig+Zl0kcqJp0W27dAADAXSm+Oknbr69AWKrgOv1W
4AfQ1bKES3BEgUoa5n/gaGFv0N22HQP3Pa33e6J+b7oIi8kgBdEXysv9EQT6KgubOx5oiJNnbCK7
iVPN16K7zUAJIZH6Q5gE8HI6gm3CHozhZH2FA0rHQ+cgJSSF1DEsn+32z+ZuSHOUIjVZvX50anS7
PMLFp8kQJ595h64ofmgGFAZej0w5btHPfAfkb0WRy4tlO7faqYaB85WtneHgAcWmFUAoZXGfXl0a
561EsFUvhmTSyzU7FOKMAlHRptd93CbX+71X9Z6Jzo/+LgK+vNf9CzOr+Dvv/1YtQPCgcdcb4Wks
RPUpnEnmnnZTTD68Up/55w1AACuzAQtEjVbI11H0/0jPOqMFKPRGDp/dIZHbhhM9U0UrzqK2zS6J
C0N2E5LCXfxSUzy8MhrsXArGyKWAXWmzKR0N2DIBpoP4g5YQKRKpFEWgZxDNwaU80+Ntdbndxduv
B28zUNwsct4L5jcIPkOk9WAFgSfUp5mqsZwDIEK20SI+7TaNqVqbzbe7JgGjhpB9EL5yL5jXFLMq
o5n6rAQBIZ+4QpfoG5laywFm8N7Ci2d9TUPuaQXOFcIMhxp06gkbitvw1vNtT8cskNsQr0reKWeS
Upc8xd3p2jHWrZ69kJ7Pa6NKhH1zVGiYPxPKKVRQfhOpWS8nJkRFIXNc1U/E2ipmcEU33M6YNdo5
pcHFv5J3KwEU+JwhfF9QdINiGyPDph9yuiTMiYE13eJxwp5Loq+c555E0lih/B7olsszVLylq4Pi
OmKnpFwDuS9zG30lMeSzu/mtt1DhGTrwtB5ANdqpZTAHuJI9jIO7NMcqnFkxtfEHleMoyVqmgd8y
Nu+a1oTB/QK0PqkIcxGiJUybp8nIyxdYfk/tElMnh6iLZ0AuQmYTK+m0CtOWmF5gKMBNnXBYEdk/
MgPw/oAb/SU8/kLliHImgL2RtcRgbeWJrNiNpgt8+pptUIVbsd4iUsarH9IFv9kvLuPF1gNktJ0X
1fZ9MJ/I6MCpT6xYvOg4tubktI+WX1qiDIN2dSk6F6LGLDAoEOflBOqgSQAUjDAUMju36gNGSY8B
fN0Z/a3J9G3AVBFIE8QQKJctIOaFfiI0MckISs3uyjjNKc+mQ1lu0X3bHbY5qD79ObZ7hv9KxnN6
X/fy2Hh5j+Dm9iwdJsmWm48KqJGlwBKNzcLy97vy1qSQw/b5NzHNeRpIPAI7oUfYeZWz2ELbgPiA
6ELt8vKl+BD02hb4/mPAw1uEYsfNdWdsCXLt0vJM2gmpM45F1y1POP6XBeDa6o0EWgckuNMccGUK
y+aXatphLHH73NuRU0dA2KzQ2EbIWcp3jiSG+X+CPym3AJs4TEk0yfL20bxrZDPVtY34oDoxOd+c
LOyrNy2o0YaQ96HXq7tOiRykMKvZdhQCLi0UhS354p0BS7uPVzwwiMyJ3DCEXx8JQDkCAm0aHwqA
HpFf1K1uclLd487r8g9YZUOop218Iln6DBtMAEiPfUTf2cOVk77/esIbXY81+1SdFijlGp0/KTLF
MBYTZ8E+wlfLv6S6BUKsASsbWygv1IlmgHEpf38HRvt7O1/+ixPQdAM90hvv2AbHeA0N32rLz7Dy
ZE/0HbgZTD/9nkbRg5/wX/Mxt3WPNZNTWwJX73DAFvb4ua110DkFiQyUmm5QFqUkNgp6Y89MIQKz
O7I+zK+m6Hw1pgCTKGk+UrNWZ3B+MK0DYZytPWE1heWa7yzuacAKC7XmGoSOl8sc8SwJWhmsUBic
6DNWO5BmzWlHTFUDMhcP5l1j/XgFhaD2o708KUL1f1zXSIi1aKfvxk1iohd9cUiVYJNROFbggf1v
NojcCWjGhNKjlEOm+SJasslcDwIee8/Ktj+H8TmoI82aebUK1uossWG0/tpehK9o28LfNJeAnxto
cl7hRoBS6Ld0TN4vLAEBmYjjVvw/oxyb13GUDz3G/SdspmPRFh0qERUjQG6AF2rYCEeugPcu1xl+
ond1ZHCYi/YO+v84sd+q4qpc2FewZchGZUoFmf5h5hkfQ/Obef6wr69NI5qu7gZPQ6bzSEFiglHk
xHW9Q+8SEienNsCMuACtisdqmWMwKhmJ5403C1U7W5L1CMevAanT761WIxcGZq9AzgTz7rzIXt2U
wulXFWJLMZhkdjeT9bBybYePGzV39pKQY6QtoUQRjq/JqxibSH26SbYNoDrBOKhZ2AQiDzXiudB6
RbFXjgYiQ7unCVHoG/pPjLSiQ/JlkQs4zCaUfq21dvQnhob/WkDq4LvFv2Wnlhsr3yQYMHe72tWH
OeRQexYgcqYj6uKzsEYn9GX9KSPOnMA78CF8zgoa9BCtf2RvzdFaVF/gC4ufaJY/d//1wP9tJIr1
ru8JsbOzqxwXfBdEjOiz0mi83iCfeR32DbHy1AydC8dkJANoNNOTBAUuuy9LxKVVWKO7LPAXqabk
L07OU3ZuFvU5RcAXe1oK3zB8edwDJciIAh8qVg8lRKxkb+Ns/t9RBGO6qYgshFQ4Bb4Rp5ELoKHu
3WQk330uPfXg+3O/0aWavK/Fh8rrMp2Z7afrvi1grI9xOpMnkn/wz0QJPQgm6v1u8gCVI9MXCcma
ugokCM/tE528ZTztlFB0FW0MvPQ2GCr/nJM3bN2hyxpCmudGbtdQcYM5iQfB8touWbwEZH6yoXs4
RdCTz29cbFSFXu+GXQCuJff2ruzOLPYRu1wFYQ7lOQ57bne94/v0DQqKh1PJO2tNgMJT3dVs1qjz
CmQc78fX4Q2zKCaS0wEXL1teAVQPKb5Tf8XHr2MscprqCl73cuIiw4C2PvOHeXGXedixjmFvS1+y
ZZAetfVpGQbTEDw+mxT/gslOiCf4iFvHcTsxXhynD088h8VG6//fjYSp4D5snDtQwc8/8JE0ZxsQ
hTobqHiEkeU0ikv4qJvosgWOAw6l/Bpi19HbRq7nZUVs4ldvQHdBBwdkDrZTdYRMyZ9eJnu6JPMI
L0bXtdxODwHhsVcowW3RjhJqzwEqV2xjwIdXlQNkYVJwp6WW/jYp7MbJW5rgSQnkcpmUX08Pm/uY
5+PUonaop6swScGbudx+jnQWL0Aev/LLA5Nc6c5Jh9OZWNTwhRkIOnnN4DFh65fFz9fRnbyARVbe
nyjHmmbtZobl6JT+m+tdUrtmIHXxZ90QnEnVbRW6Hgl7nYAgV+C8qUnb8dOd4mawzT1G2i/lFCqS
21+LF5cFIdmo329vOsxWiZVd9dwP9r9agGBWuqjQSaC+09lZ211hajz95fT4C1DHJritcM1JxFyo
fOdy0LZudTSorOslG6e0C57vMY5WioQG2lXtfk+p1bPlquAnWfvndxFMRG5Dp6vcapcmkXZ42NN8
epknbxXQvuKHpq88fVl/Bi11jcM6i07XtnRL88NhVOIQlB0nQn3eOn4i/t/zgg7whtS3IH+Sot5k
41Ndi8WL+j6KM8qZ6PdtIzwmQTDfTssvXOYoSVDRUzRm9d7owukNInXGyIBLT8SRZCGs3Mxgyo0j
DeOfhtj0/IgyHHQHXki8lw+E6CIe8bLxWehEjv0I7Jwne1igXP0/HJ7JpiGKFvPqReM1plSaLUMu
1jJiV1VCjO8lldo36adPQ9/x8WC5avx6atxmbjsD6Jzk33bPEOBe0nK6COSR1uU8nGpNllazbpZ8
8iqnQ5zN2nuSSLM75BYybEfEfYzy9tgrjzaMnGIWLRD0w//HAX86iywpv61EksBFNH6vLENPXCFT
SBuKJVLUON8WSSCMx0gidd7kOVj2YxqMyTl28rKeV/FgTxVHLOrynFSNpViCOTFt9psjKLfFQHDR
z8Z7ADM4hh7x08c5Ejczh2zlhv0ZjvzKG6ouYG+80LljUSq3HIZBOM0V5zTdbmUntHbJYMZBiPat
jzhqOJabTZZuPoI7GmSA932vHGHxjtYtWuzc8YbGYNWbzAaRU4xIZ/O66glXeK5DSPfFLigbOW5G
l+xJgTfZlChjYg9zIVXXCC7ogjmBHlE17cQNT3+1vD9TV5OVS3xJi2aIFCHAJYLDCFD4zDJt81B9
gSTYTGbvNHygQAUU1rEBeIgjwt5gtcwEEoTC0S8OUDsU4LNobdQbfH3dXZkWqP1fDG5HhgUSqoKK
WWHZV/qLow8qEccNbBaFOdhlfMFLbjSQrBrJdBQFA2hmcIrX0+JYdxp//AZG/wlBAAPN7mTsUkrr
KpGmkVqUu/Ukgw8KtsmQTxBp25jVBruVvneMTXQq8LCtV5ujfu0Qxut4Y+U0J+J+JvYsaexbK8uv
BnqsPRZDzoJr3G8fnUbMKJp+cpd0EhZoyht6ItILVVylrh+Hn0tstEFtinGTr2lfH73y+64oEW02
swUkLN4I/FKT1doMQLcW8yIpR8xp7b9Ag44+PD7XxvAFv4qc2RmPHb9w+UFLVHm1xQFJvH62I5GU
TW+nSg8Bk25OMJi8sY7vtrhLhVwR8i3CDjL9VFdRDwgH17ggEYDltBgIxXqeTIGPux04+NY7IwMV
8mz3IkQkG82EwTg/z3Ppn1KBhTGVXnREHg1v44Inu2Ts8xjIfzR/7hOPJxNe7R3is+ZkELHMvIFa
DWtS8Zj9hJh3Qz05iq9fEUH/6xVKGp9FMsBiPeEEoWWre9DBZbn/YbDTFXMBYcrywXFVeMcCm7Cb
FEYPlw1+mYNssyNLrnSGpkqYk2GKQUZAU1a7cKu+RHDG97C6l4F4ndwTIzuTK/3WyYBTEGnfj6Fq
rKSmNTV+aAr/Tay566a5iVd7oAofiVAwf4ta3zVgc9rKnjNw3rm1oRvleJOcYA0JPacjDJV7HGjx
KSopE0QXTev75lekKLOi4BumTZU2DTMISYZPqw7g3+1q64D7CsxLgRMKQNKW4AMASPrdA6dZvnM8
yAiqq3zfYt2zqXGQFVP4F+kNu3azxEs4eH3Rkik5OL6AUUJ77kj1C7iUqRVLIQuAPuiyrnDHEzrt
t8dfe6QNYh1tfWduKwlf8gz+IoWWa9xL5r3PpxFAvFeYPKhyochbBGg9lmkhfN/Q53My3e5A7XLL
KO5nGKKIll9CeiaBnID7dpcgF0QFy3lsEDppOJXjdogxgQXxu6Ug/a4RM2W30QwodKoY+36Fmfqa
x0xaMCs8Vak+T6GkYb4yk63wsNEt2dZS4t1s+Pv9mpMy3/RyHCDtG/wyuqMNG6X5OAFNn2kxaJ9r
P9QUZ7EOSucS43l2IzYQkCzZ44yzw8MlZzl6uccf0YtvAPRS+rscDscH6ySrGGfEYoytmDbkCLA5
As/MSOwtPlnxdv1/69uJqplB4mNnHLRi9kIsCyIKGNIowoEleJCPytqz7TDIXvaMi1lZ+UYOtieO
W+vVVyCSwxQWxD1s6PCA8VNlmSB7pO33bYgMOQObd3OEhzDLiudXuOlhu9utDiJy6zlvkCH2aUEA
+LbKZH5VddBGGXV+HEfy/4RL7TdrTEh+ct9EjbE0p31mF9bXn5BPysZMfWXuL5YzTv9dqNpImLg6
xJjPavl3CNItV4yGkTuzDqeri/dv+vlgzB2Bl5f6HE09WIZPjJSZPnMVMsUJojmCm21N9c8lu4fK
p5qXNDNLZJLMng3vLuD6/Y3PJbn2RDvLomtTN0W3H/9uhG0TMs86WlCUZGN468TspU0yxIa0QFvR
TQDKqc20jMe2viC3IOlDB0yUX85n92eAK8FgJPwOhGsZy48uylZKx743+IrTn4DTrkzP7QK43/BS
fI3nSnILWhR8TA9GYftfiDQlTuPONuQl2fCeSkrKS/HAuhlL1seNwrlUEPDGp5bvKFulPsCr6a4o
o4YGaIdNne1JjJ2s0whfPkMqCMYWNenjky26JqIqYN1340YpjTyyWOS3u6dqBIsQJ5i+1VCYTewY
U3Kv9pSWWt8fDJV9TE3LFU9GTMmdSrmdJK78MG/7fG/q5v7eMZDY3bi/AUGnXsvTXjvRrBQ/2UZg
xQGAgI+ykK1ANPLPBk6Hp4TYRIax4vWiwzzaxcrm6c8USUffGTKBHUSKgkWmMKZTSx4Vwl/6vEAV
28x2T9ePAAok0hNPUkPUv2vsOe0n8KXmdakt0XbXbX9EXKgkJyGpQYLCmJmsGcjouN33KyhIdfzv
gfPqGywh4TqVIqJWHnOjh0L+BwYvvjtybnsAbM9SHVBtYzQ3oUC8zG9ouiLfmkNYJsx/pQ+H8Ojr
jXBQHGky1Pbo6i0nV1WtanLUopXDWjshLtIzbvsqwjy05WDGDkUmgcuN06FKZrr9lkdrvzCJ1wce
35yP3BDBf2e571Esp4srKQ3KDKRf+3HLkJnTWUIvJzuQnNFxvAdKLfAuCY0kE8VtzMFp6qkZrppZ
809N3iOuAQhLwNAGJwKDLBn58mLfUJeJuaNHUUQuIQsbcM2U5uP5zebCzZKti/+lYLuWleaTrWMK
TEONMHHJYlDNAB2GfBTvhvSDmLryWMh1mWiCUtOIhwKSzphAjhaLCE/rsvmDGuhDV2XfWGElPHuQ
SGIWIkgQVLjxx4zMZa/DNJo3ro5WP8zNa1EPfeTwRzzJJGEiLXwJ4NLLCsRUZg2pUbDGVMVDpwCP
ZnBDhxgqwxlT9dBC6ZdKCQGZ5EHGXUygklx9kgDXOQ4oawVWHKlOyA47fwbpXBaJrUEJ7SQQIzVx
gHLHKOmUTDVt9bGxHz98SIpofvTcUDW+sL5AeYs4SCXjp1+KXnZrEP4BxSbq3Abz27tgdawEUcKx
rAf9kxBPjCM9s0M5CN/8hkcGRIT8Y8jQP6NZ5j7PdVPFe1czhr65MKYfd8cC6vuvJ2LgSdHRhMD+
VRaOcK2q+mV59cRvp+r9hClpyMjg7qFl6x7Ds+VmgeFUZCKxjFVPBWnlW6ffixnLLudec3UChzco
CX3YAl3FNUSEAOeAWKJ5kNTGh6E9XEvhW9iOl9hPW4w9+Zy00eSGPCqQR2BdI7bgkln4h/FNqDZj
26WIGRQ2yIcin6IrWCVpDpmUFJptnEBypUYvff0zsdpGn4PyY4wyowIyEKLQ6a8KNd5wKXS6Iivu
EmQGOq237pt98tS1UGlQxDoQIu7iD7up6fWBvDhR6Q0pN+qEWnNWCwmnaHYz4tPy4djfUP1ANXQu
35ylw2yzl7OIDRustx8AvHvDdXXIhHeBuKGmLirYH8gXwZ5acIGamUxnIRhRQnuphSgG5ha1Xay/
9CLw/5m0WB2EgKTSDDNA163ng6GVNLcahusXSw/LH2hvBDSVhRRwLmzgLUjdpdUUHYN3Qwjsn4jD
dond47sZcHewAPm99evyXzJtKSklMiNbc+ST/ls2sv5iMVradNDEdG6wtAy7E1xGbUJ1ABzP1JZS
OJOJJ2tFqxyk+HOWI0PamP5fxGIG4NIOnvuHBpbaDf57UmlyBC8QgrZZYLr5SuAQrBW2JK4whHrC
g7MwBm2BgzmNgxwag5f6VhrNZVtLZqMrcoLR9eG+SggDb82Wb02jzEMUprvDskOD0Gbgjk8KCRc+
/QNM7BE0gi2iM8bJW57s3HzlIpkdXMmHbAWH3mbAzcQg6esTgC4iKd62I5OUC2dbZJqRy3/dwJ7G
EHrIOcCQmH2CDdiAYY+PEB2c6pohyFm/lbLz2aF1lsEdTHHh6oi9xKYfkuMBxTVAE91JuSVibWj/
PSxXta26dcfQKEy5CGPsDyz1yDn6kQMJHoiOnM+2RLu71D7/ZMGse18iF7fHH2uV7gBMQCuFabqd
LG6syNvr4FXRRSf2wsxtrxmLm+HHxR0z8xvyFfuh1NxcTHIxTBkxK5ZKOaQ4ibTQrHDVmoTprFSK
msNKYzJ8WkUW7wmrbKSh6GcbPH3KQckh8EajbMTCSwT/GoqYJNbOH27M7yIJAQBwEsG4206g/Y71
v6XKGQNIUyijYD8pO+w6I1EmlbHZAQJMmMX6MX8orbzFE0zNPcZOMKukUssPqBQPouhonQNBkLca
VzVqbWy9ZdFZtPvnHjIsAoWAAAuhrpIfBIe3EBLAUhBaa0LDxK82NNAu1RegkFAPAenGf0akmro2
Wd4nM/1FfQYePcgRzHCVtu21DNDkiovyJPhfevvgqhDtUViNVfiAdiUbAc2K+CMC92BdrIPXhNtV
lbHTaRO4Nux1PesS7pvW9f/5NKe94mGKoxC9K0Ej0vRWPJp4g2VS/+fa/jgbOZ+G/ZKmEvP9rqda
p3F/WF5OXydOEkuDMnjXCT0hM5cD4ZWu9UTGQw6b4Yx+6IIVxRNfG2gFUQoCD5gxbZHfscU6UA/G
42zTu2QYn912uqvQBJegSpUZuTiHjpBq+bgO01nd/eOupRXEQ78hF7yB3WhGPfFY+XBOeEDaMrgl
lZaLV/hrMYA8wCnqu5Fc3q55vuttNfCQgTjhIvJJT1ocde5bp/NSpA7zoOvW7GWy369/dxsqlk6W
s3TZV904AgXM6G3e1slzcjH12enGlF4pDgYg7hcvjtEXAEb270uH5Ky+31eDgdBpbDKn3qO8OKUt
zaM433D6ygvGzIeqvwGr6grOddYGSu2N132Ov1z/jEvP4SxjBEQbm8+dkFxYhM4f2i3joiGT+TzQ
qafYoYo/7bKU7WiimaDETZfDW03kU2z7G0M05cR5X/lV9R7ZE0enZhyzmEixmAHe8gIP3pqqlCQ+
wxq19JAc2ilZCJCvnHPZkb9idoOIou+1IuSSZvDGQBUF/YfPeipiZBY8UjyGndJQtXOI08fSzS36
J3gZQ5zEDLuZTJBvsTHVBMtwJ1Mx4Ygzbq/O60+q9OAdZ1lWvUXs4uFmO7N8DU60LFoqXMzxkuAn
TW0Ny+UHXpxXRI/ueUS34G5HDY6lDnn4vIJgiUpshNIlm7y9t3gmJ+gH20AOAt4hEV6m2NfpYCE6
+BgwVVJ5RivjJenaoFQZMH2Cil4/5awx4mXZMopYTExYUUGQoNwZ25Jje1D8bv/EHC6wU+FF6AdL
ZrPQ9q76eZ1tph6xG1Pvgmf7EtGuLd62iXRC2yT9riTZB6sIWExu7t9XBFveqQUfQbxcA+3xB81V
JQkkYGJIOapZ1u8cx0E11cNoA1rn8DqHOoEPG9/RBjOHWytoLHV/7ISI25HFSclSIMJRkuoERCMC
uqf6ClhDO4R4ECaFhqnITaQF3nA6FA5/t0xno1baG0miLkVL13vUaMVfE5A9V7CHbBFC5m0AXJiQ
/mixbGm003COzbgH2XsChREEthHf/yx3Zx8ZEeTIrkoGSq5/uTmqr3Y2Sygy0oUuvnQmuJdbtidG
wC9rKulKc4eXC03mDgFUM74tAyl3TzMWIQ5WIDQQQQ6UpXNNOGiNW4pP1evJXTibImjcyzLMRHeu
eyiui3XtrPCCQo/P+bPXQMZNLxAWzI7MO/UAnUspat3r6S5A+nroDxbn/rIRWm50+u+TYIiMT49a
MZT07eH5bCkJZBG3CKqmjzuQHTKLkTm7IyaghtaAjgXOVFtHWjnmvVoU/W4z8DNErUINtwtS8iDp
rPWXw3sjcqBmdULuNR1fSuKQue3P98Ec9539nzwaoqm4QFJtllG+It1xWDhdgC4WBqaOe9CLV/F5
IRRQXlMgMbIetXAsl7hg14CprI/SwpUHFbEFOAvXeRYolFfxgu9D6DqxmMUKHLLQ7DqzFc4yUqWi
98lVZmMxG9FV5x8TilKLUF+NgVHr51b1qFB3RtbjHKqjrXAdbGJzr6PPhjoaf5IbMOYLH4hKJGwO
JMTi90QfVUwEhIYvXYl3qDUGUgcdBrZGg7dFP4bY2y/jD7lYgoail68kCsv23nY1u5Rko6dPpnJa
PQ9vEfqR3Fhah5i9dRyVZam0cM9hgwg9MEbR8V79TEIJQ2oLj4PaGuUmO1DFxiESl2su9wIa2NuP
IYz0s4sNtvUGXdPxqKLkmsv0eEtRj9EhY02G4r4XHE8uitbT4ROHbs2pcSizGA/e3aOrQkjyyYVW
vxZkdH5Wjkd85rcKueRiV2AuMgj1M2+JF+O7tpEuWop134ouQ5nb8nnTkQ8X2+e6kO0kPK/+RLS7
TlvP0RKB9Frzj3PcuUSnURTE0sMPTlS4wKq3dEu1TPnhCvwsb9ViJFrEFbFxP2nsWTsg6XXpC8t+
FeBJUKG4C3ZReEyL02xnQz2sy24FTUWAupj2VMs4k8v6NVMe6jJhBBJoR+6WMfi+4Q7o/CYzj7df
8GSnbPwpts/BIt88nA9gzPZex2UBBdNj3Xa+IpY3viFYIveJPkOVUFEFGk4nHWUHifeDnXJDfq3d
Q2bjF6+cYFaI+KguO4fUKlMEm9WN50brLrUDa6IG5m1Krdj4nAYysoeXA2Ee0rnja1KB5XY2/Wuu
Z7N8CNcVLbVrOGXM1pMNEW4XGD3ZeXjmc6VLR8QkpeSfSSN+ZisUce2q2GNy6uNKtQ36ojW/6meN
59c6mLHGMkZaKwZFTiWaLjxyzx72T3LnIrMigKPsO5B4HCxlS0sWD8SorapwO6KSdY5j2vkMXUk2
2xpsnpVHta0YJnEK91tUoa1MvaD0UXAiNUu7ebq0ZlaQjtmbvjdFwvkqk2H+Imn0TqZhjZjARS1n
ASp+p4ViufiIzHN/r9WFwcuTdmE18Ap48ECJ32T9WMHPBcYlnG19jfSN81+Ukj/JXm7lpvBMRoGY
H/OOC0zzfCeaegQ4IB3gVWzt6TFkMkY1h/aQsLOTjOLqJnOseOMgYpRMIYkReXHQ+i/J3FNVneKN
ajZbSFYSvasA5sf3WValAPd0FGRQcMGvcnziV/GPbGHgD4/SjqBBlodQSc6S+J7+JwIjjJFZnhYR
m2d5HfP/npbiuI4acBHoKqid130FeHuuxBReLhK5MbBg9T5mJ4jkh8FGvxbPpvZBQ450g/KVJ7qn
rOnVDvLorktFzplKwXHqMdv7bPRlXht76TKhAbmhnZskSqASKex0tZR1BDpQn3Z1ZS/eAx1fKTT+
sWzFzJmqWkQH3iR1vAqElQ1+/cciagZo7V8CTwntLnxuqfivtJZHOi5JNolaXTi4AWCGukd0wtDQ
d1yrkasLAm1mIlfxcvCs35+R8gIoka/F4iWeM8HS3wc/FX0hOsgyj0kk9xBjehT7zwJMzYnBY6lf
OyGSNvtjWN2IqcGWyiwoAi0KbFFF+a5+gV+20VNfU/ijDt0LYOalMNtttGJIeGz4ufoBYV7wzR/c
v5w4Hlw+L0O4ywn1ruStdylJeE8Qd9FSd+7WriJnojpHBzgmJvNUQwoWd1aveqrw/PP/ritojPh1
vsv6rxxN1SoWMtr+04zQuRE3gTsPaIB6qWLpc7YMuf8wqOl3r0BrHDmnhwb77iQ+uHnk1qhmsZQa
OCa+7xSRSyHn8+gaD/D1shZFUzf4GeXV/Ye97n/sbNaFWwTC56F+7+VXSl5KHE4T0vtWcc+afBqd
d3rA/ulhMMnHOdlNNU5rYlTtw/qzLFPy9mAU/25gE/PHwXl3a7ShmvgLHP7+uVI8z6mrONFgqIbG
ZAoZ2U+MfPV4FBiaYwnNYTyb5TF2WPvROC0bjlL/HTKxtBqKwrfV/Nu38/RdYN6wXDS/3hEYf3j+
HnlclM2vlWtj3pWd8hiDo+EfZbzNETS4TpdbnLsSW0HTSm6MX49ny1S/5osCGU7QFLZ9i8oX3qjR
vea5p4rswllfjxwmv5JmrNDgY0rGeQEmAtlTgK0HDWfEZXMkBzdOYwO4Y6FGIxEpo2Nw68eT9Txo
ZSh2XomQY5CROLbwq6cq3iaSM7f4d7FTfAinJz3armV0t13s3m6lKLq94FJLAagrPYAIzUzw30yi
HWdFDO14I5HnK+kz3f+DSV0BSbEOi04CfnSvXs+YIbHZY4EDPysf2nyfTlPbAuj1wftfyynEkE53
4NkAtQixfcLe61yVwwS1knSrG3QbHBRzoxDym2Z5EWyBrWImxC01GCjGSibcay7fyks7Xujd3oZb
09W3QCUba0+n3FcyYkC8H8O/u+ClvIdHQVc4/M5s09E34MbwJZw+/YaAva6IVRSUNa6s+Lu62xUR
BZKlj4Kz7mfbdGOydMJqukxYNYrpevJaH1LQNwEtVabJeECbXU1GvTW9Qn30w5p7GPkQkN9d6ctK
VLU1WCGbdF9o1KCIdKYNCJLTrbMWfGovXooktqFNpM2+Dv+vD5vgsCMd3GlKgfjiOiEgIqvV7y4f
fMIsD0cv68njU5pwecrsTND/Z6OvESDF4tOXviVLnKs+/w2XipFCHgYQHSEsmZt0sl0wrUy3bYSv
HAiWkMkkvrtorAe3o7zwC59QVAgO7KSIOdV54RqE15RR/EOZUGm+hj73JC7G6ywf1p5KQjcn7bj2
9V1eAPEpYMkxtKbDTUKfDl4i1W0YEKOO2tvwYA4J2hgxGBSYOo+tCnd6UhTl9lHovCkcM7QZe0fa
JXfwafLiTocvysPUXW/5YtDKEiYp4TbvoDqHxkSrCBBME8FQUfPSTWBNZ+o4PuEzI9qxS2RLKzCU
jmWHZTG3fOWQ7ngSpYOYcjwUONQ7Lcs/GEP44Q6QwrSSUvnwZTAud82BSEWS1UGTSlyYNvMHb9m7
wPSDSuvWUasxi7/laAv5zL0mcxfz54SFo8PKURz/aRKnHVEXiN73WoWNmz3wc8m+s06jGzC3Myys
yppPKwnhUSbXxypImaZ6OlFFt+CesAcPiYs4T5F5pedlOGsh69UqaOe1G8C9CtqPJYh69fPDy9R+
7F3WTFpz5N+VkIVrKla/JXliqIpj9MCE85YQkZWq8zdmNtZEzi/NvsJxFL7quHQNA2OwTMVzfRY7
Cj1MXEjTLgCVmF932cpCTTNHKwyYGTrLJiaEjEFajD5pTah21caH94kHW9Jj8ihSjY+n5d+8gpye
K89O+Wzyr3RtwaMP2U1L6JYAQkhmvu55Ut7k6MkT/0tG84qyIJ2miej61HSqqmaWZQJ1eIiBD11Y
LdwFwQKkEROM8b9HsjKPyLq/6tjFEwDw54djpmTSHnfOigXvBHwQWXG7BvCP7UfrYKmFEpmjcr8J
6RTcGYmoFt027dyIhfIIf4IejCWqUvi1uFT6ROKjzL7RA1HUeWFiSBCD3M4abRG5TtebqpaKiLjx
Y1u2UWJggu8pCLFrBvGomYH8QDO5OnLbNlSEYhE9fDMoZI6VUffxgBJb+nzo6zQB9kKTqjLtVEkf
LFIEomYt5D6HrjeZ7bbe5uzKv02OPHqdU3jguk5GKNV2B4uMuz4FppRWmx+uVl+hpuY0tLPqlccB
4bgETdZIi0IuaGbMWmmOr9LLE+Vqh3OdhNzE0VdX+P+BRamDdZoivsg2ylh1p7IHLyJmUhAVUi9o
Nbm0uGYf4aeDZO2Z3hwjwRukMEoGzGTRk67cuEd+mo4uD7pcuWhyqzh/a7835XM8Ucflxka4K0aH
owaU39VKQP+eKiG6ImBzhZ95UBhOSyvLppi3q5/tNaJeIxQdoJDLW0OE0GWW8eZPqFzB061Y8CaL
gkFRPD4Wo7gizow9xPoydNy3FMTewNBXnfZ/etdUep7I1L1PqfZ3IT82yqTlBRnVV6yiCisWO60C
BUuHN2lJ00p+6a8FejvV6TK6l+NqM3C/PLKhbT/A13Wo1sBoCXIKWYxwhAHx4Jx+Kl2czeYMGC9v
ymO6kITcu+5wlV15uOaFj9Pcb3fb7GSqEBDFZBDAEzMZZBc3dLieBKaoRVMq/CR0YJ7SBXHO/x16
1hn9Q+RXOVDsV6K10THqfmKwKR1ruoGHjfLGr5uqzRTwDTNkNDE/lVCwQ6/YvzjqWd4TMBGbOz/C
EsK6bpms7BaIfHgNXvDUVYHZd1uNtn1SunhnUCrRQfm7amo8VocH0zcisnIob5tlYXoQqGu1KREt
2cfDp8WV9ouVqkb/jNFnu+lUA7L1vhcR9nu8fdCYOUTy8NIHhUJMu07WMkaWRVxKeXmi+gXyTd4Y
3Led7vIn0340dw0XWyjWbRfDyI9hbgwhiWStvVtCXX9a2WGWcHtbAMbU2I2bcKQdw+Os+WeZ2vBT
ichDLyIipcIeeTXiZB/Gu3VWnYaLsiEZGfL/jgEGZ93E/U/TKjNSfx7LWqCmab3XLSiC8ouV3/0g
jDFanuilZAKO/tKhMvsStoATUqvuwuIEdHhSsTr8uEJ0FUT0qkwiTowKmphYBhetZZnOejpm4Po1
7/F2u53TYy/lSYKRpOirzGZTK/9g6ION/h04XVVgOytMm/9jJN352hKhwvo9T6Z+ZRyWH+VS7lqG
npBRBHbQ4XPc63nKmEBnZAULIJrSo2SAYdrzBI3pS3K8Hfl2zdo0xjmQDClvuJTZ92a45hfPK8EQ
5CvNxJBwleqp239paONrbLlBeMIUXIroCCrn+eA/Olqma2YMDA51lUqB9bN6ePDybxDpaVgSq4cC
k9QE6Z2dSQd44Lhv1xT34OsaCCtwq2P3OBJuTHhc3gmR3JMrHSRZtKlQV9RG+Tv4u5mkau6xvCDy
s052/w+1d2TH6yX/j0duSQOuiPLAMqJOfDywwjOYWg4drOwNpzExvDF3zUivV66AXT7TQkByP3sk
6sAWdxRqtxSXPmyn1rPbFkwV2G29g1Job97Qwf/jyWi93fVvIDynhilcLS2OUaLv87YR1C8wpMFL
QuGMuB1Jrfu2jeAaTnUJbNSQs7FStHJgHjxFt3/3qIoDiw12FSNQHOxBO3Oc3X4a4R8MKn/aURgZ
EzyjpbHHntFyrMdS70phqc+LF0avbSKOuhchnQQ5ww02gk+cxBwgdpSvXu7wjhBtlZNPOh8EdVe3
5qeS97+W1d0fsHFc/+Rdb3ViBcY/NlX5w+FKH9l/R1c8pniB/FYMF4pCS27oPW+lmk6zGuYn0153
YOHo4Q/hzD6r9ZgmtbagdvB6bSR4AjkKjvmXHKWxYD08UVOx3MrPIB3p9jVmzXUVj+s1uPbEIq6w
2C4jpxEaQxqmlOLJ/HKL61waLpn8niqTM9eLWlWXrABTcqE3mkDK+8DVRWGfkkX1ABkYrM+bU13E
Xed/HbzA/28aUx/blt35JkGMVpbbCGEdPaVlIHQqWLfdjySW9U0F3p5tiCmjWZ+QRls689PE04el
auAiCQCeahu7IyE++VbBRlxHaFrTnglQarM+FCyqNi+NtB0Egy6JVCfOoNB+blnZ+ECL/0cbsfZW
yQ1g8qloF5UX6c1YE6+5frO1tkcv2Xq8MggSShrXF8ml3aPVyWqCjulo1cqBYPIOdveTzpZS+na9
CZtz0IaAj+m9qOHQdReBYEdSsBu1dzAcYE62PYBR2ZJsEp+JXWhwsY2+byVFQmmGyuzPIOVbsr6R
5RtU6QZO3oB4N8Sn1PpV0h30zz/xbFJThWph5+pPJPqvxIkvJ9vrTgPb9bwZgwzqwegDiz5bg5VA
RI7bDpthtCGuCRjSYcIKmv0XaHUiZ6YJiaxWlDi+ULPGvRDBCWYTsSQxNo0JWvzMM7Czei3fJTxa
cniHQf2gWaLL9tDrxiIYT+y60J5Nw4KnEGnHbk8+cY5NKLdLR2Q+wLvZYkItXbhMt7gUfSfQEXxu
SMIZnbb5aIvv+VMHQuW/2GMXZ1P1XFatUzcou4plnshJCr2a+wpCadKCVD4snECQQJkxAGQE3Jw+
X/0GL3w+apFfnL8VCPyA6X31Z9mRXRYmYQjEGTy/zIgZavLCbPWiTBgQDu2qbVKI4ktBA+ZjajZm
fAIeCrB6kqBnES7y0MudoyrfWIs1ixq6FSc0obNH1AzfV343Lw0ISIkG0eWy0TWKf14OedNcPxLX
YbdqNpO1Ppo4BMXPAXFoiDVuTMY4GzfBjnM7iYG1Ypq/BIDHJgkpS789YmXbap+ZfW7hl48I9fTt
ODuDtkt3C+LGQwr9r4+aU5mNQy0A0RmjI+ogaieTsDhEbrtW+LHocpbszYVyFQwNIsQAhAEkxDSJ
1UNuMcVkxcS6HR+sKZzegPI/B1sL2XbQ7ocK8Au829/VFwo+ezqSnk+G+t8Ub8dpQJUSjqymb1A9
NdRmIpgXyYH2lYh0YS1CN5LVblfdoF0gtUy1+cGEpGXHor0E2CuG2jaVTsBKi/lvjipUGNQtk6we
+7V9h7f+j+omB3aE+SOMR1gE7JK0la/8ZozmIeL/XdYxvb7WwCZ2fYXR8S89H+LiWL0pyULmPvP9
3FHZxjXwJOEggpcAFz6KAfW/vJtxYQqpWhCEHECn25cm02B7nuObGf3TpS3pLG0cgacGKJk5j4k7
+/bVLvd8X8HiRi8yCpBNWfaiqVTQBis3Af8WDfOfxHRNEIsBcg6x+HyNZP40NBw3jjGPbdVwi/a1
NevGYfErKO01/9uSGZF4zpSbcAW0KqnPd06c2vchgh30/VnE0C/0bDxf0nVi85ZG3EN0r/Wwls1k
QHX7DsHfXaVbaywBnsx1dFLPpa4YxCQ/AHDzFPJsZ28Ip1r4H5rWftNeNGegmAo3+IRRhAlwNgMC
+jVMxcU2pU6Hs3BSpliO4xjjpeIoaTBETpxP/ySGRwDimQo3i36fL4ck4X71ObbytMhbgIsCX943
i9e6RBC/SU5tqs/glNYop8QiOpynvT5pl0Ohi9l8QpARQNrHslYTYa6eCIRdTnBMMR7gbbeHT5ed
xzbZiHkKJ8MZwkx/oAbEEOLCp/0x63KyM4/mu/dDAf/TaILtSwfGfNzWRsCmPR/dQwLGydCrcnQz
X9TZUlLLG0JR0/SC108ot7lSgJpkpnXqFFGS7WskOEylrrCmi1DQFAQMrVTTT4T11k4e+P2NMrsn
kZRtFfatccvJpcPbqbJuEFsao2F0oyPjgYDSDGXb/OeQLIn071S2zbpjb9rRbBObLpErM1lLO35Y
wPEb3FQjiNj0euAdnP766HCblPsDwWTANQiUSpMnDSHMMi5grpwD6H22Tjg01trDe0DJp3HasbzV
s9W1+A4bUygZ8o7jvFxuA+3Xv2P2WEhP/p5AI476LmiHUWZCeb97P3mwihB1u9kvaZyBzcLa9JZi
yjlYG/BbqGTiXvadizCCezT6dLARzwRti1QRqCDBYz7tq5IYoDogcF96IJw26BbvbHnRnNH7oK6G
TOLrq8BKyfozis6+Hop2IQ4NZ5zwJOU3IebBstsXIsTx0uM5E4zlEpn3/CI/bP3RIpddSOPqYZM7
CmZ5/AEsexI+ujxmFyIHhQYrCsPEtyuL5uYFekqI4mFOt9zD3u7FvAdCHyipH/ADU66E7E75YYTj
hsxFtXFQO3MmP9TclpSa+6UmIUN6k0tU9UBUP9eGkOffj4nIidJZC6u7S7Vqvl5Ds4bs2HPAvTbx
yK9AuHibsWtY4zDv0HMYCtlitFoNLwf+Ol17g+FgQvdIQlg5/jIaG2iSAVZM8E/7F6zy2qP1FCTu
ZUYJqxCz6nxHO3ETc3oJzPBpeg1sEMoqRnKN7m5fGeWu99P2fOEhViK3fh7Jv+TBHW7eAjrux0Lv
nB5myetPppU0RM3/L5wUyrEDU3tyh9lEan4o4a8ZpyOADLSSM/SseD+zw8Y7ft0mpjJVfZ0+GVkP
4CkFgDxUqyXjAymL1fM4Gc2AH61oCfxwI1uWniQX7clTCJR+dVBkzEWUxE6sdOmqQ2feuW5r2A6G
hLkClUTYFmqKwmYw7ELtR/VDt7+DSXlSIjzptUVOPJNwqztlNq+w65USLEeAEVThzLb85MmBZcky
cq/ZsgJEyJZ/q6i/QVOYZCL8mS3JQ+cfoRuFGYabewPaEZiXzSJS5zqXKPvvUTZj9NvbnlQmWrt3
VpjRi5/OPmwfHSAH4fyklY/m2YuwvuE+ms3x81Yq/ImCkQ5I7QWcFNPKStxdMTE9DFYDxUArxqgx
wrod2Jq1IvbMxMHhnpjMOqOlKnIJREoW3+i9gtVG7uLnKwRq/xB5qOekw9n9lTB86WE18LkgFS6Y
hPb7J0pIToUeBjvYZ6FsMUEGuw+W0WiTcuCGwOiNHxWjH/OA8/5dWgmlUAGbBgxPrjTn6h4kvmpz
HdhYiVbxMHu52AYRE7T9xfqajGpYTQX9OMGxKDVm7MawXq7IWeThsPvcYSyFexasE5CTFgKCjxDl
VIOuQm1sjLTkPTRXztyMjnxRujLTfVWZkA+VmEc1qNOX4Qkp7oHQmaBy2g0C/kZzCrBoJPuFQjbh
xQAV0T3cQAw3eo3qU5IwMVRJmo6B8TlqybGgyS2+ul2UaR5j4CKcS9YWHiSVFPnJ3vYMLeAltHJA
J3A4EolIDihxXAORyt8ubKXu68PxuyuuwH+GVxW7SGIgkb8cvB6eet5gzJE6ANI21ca3T7m6Isny
LtH0CwNXm+w3gKlFW69lAoDdKKBQOqf2ZnZewH7RcoaOA/Hc0aLqKoGQ9wO8Yoip5tQEULuHJOx6
rZhdzWTloUWLPn7EmiZkYvuo2ncL8jVJ9jIkCe4iRa8dx6qinmNbWY/a6yOx84IMpcqa6FdWeGRB
6VDLKIM/G/1SInEQOHpSJR5Hx2NyxVY3yM8aO9Ku9RwMBUUS3bJCbeXHuiII398NP5UyH2Jf2Fka
0uV2XaIBCdWDTC9B+UZBQr/ueQjDtGrioelQDatf//CWbpLBimgYBlY0t12o/CV59msq0cXgQcYA
hNzj5lyFGlBNmBA8ER5WswyXA1rHAfZTVX6C1dQjX5yPPcYZpxT3nMcy6suop5BuvOh058buasCt
WjpMqS/KCGBoOong1D/61rfrUZk6wWEtAos97bM50Ouqxmh1nMJlSl5WAv8ARFmmjJLZbRQmArjw
fO46VKZI5sL/kT7CvAJrbYjv6Wi2IxuloJ/CICzkIxahpipzpn4Gb2lvz8z4CbXMAQIwB9hHS/3a
HZhNwxKky1B/KTSaDGWJF/dJzUbDazUEHehEIAJrf/SWsAmA0AeWobN5IEfrrZDzq2FZr27bMU0E
yLgjLITj0+pK50xChhEq6wdPdyUErdFfjwKsgAPlplePoblNKQKSqEAufNQNJKCcwZtxJN7FM3sg
ORx6TmbaKYLOtskUiv+3xQvx3os68RNoBBMbtNvpreuUSSVUI6cJuHODATdvGFww7EsVvx6vAYLF
qvcf9R7bzQJa4q9mKGt9k+quHO66CLxZ0yPvbQ/fjJMmLfVcz/9+hU0FX4OvLxuf7vtcv4wlVrVo
x3VAeWNCIO7C6dEbwn+ZAQLcyz3Lz/Q/qowtNmJ4yTmQfCYA2iD/Co5NdvcTDpirZvlCExElxq53
8Dc3VgbXWmoqfmmspIsK2XQNNuOFkOCQ36/SIbr2OzEUDH4lCAWQBaXxZzr/LqWSyB+dvQD/VQ9a
WTw9WI2XW8uRCJgQckd+UNYtB3wDxho+r+NyiE7Bix/BTivTEZbc5QTYYL7cbFt256ubwSOqo+Vp
gJMj0/k/WBhJ8OrTtHJQ6+sxk470pyYiibNhSr2TKGjsU0Odp6H9UIDmic7Fv3zdQxfdcS1v/pGJ
52wxmrFnWurIL0i4yBZ3acbaEJbfBgax55AnNA0Dn51GnqfZSAXpuKlHi4BGehn/myas8HCJapJD
YIb13P/ee10gaZWqv8/K3qRw+EI9njQsAo+7pNmXEYNeSRcTBR+cFSM5Piz8f7K2zJm5H/yDpB/z
+UFQGAtd/m6PTGTLexFQVBP9bY007GJ2A0Hc0NCDnynNq6HBBPHWBMLm7CBwv3NUmz/v01VYhgis
VROvGi/izIEe6ZPqTdcbhi2bjLhyTz0n/EB0JUWWepMoL9rJO5b8cv69ZSJIlAr83RhKQ/8cdBld
MhDsKEmG/moQdfja3uyDIy3cvrF9GlR4B98aYYtovVy60mf7Xe/9ryClBHTB75LSOiR/3uuTLByP
CSFC+rydpOdv2kFE9qqdSiAUfG5vhNFyKjM2VXJRR7QI0FAPgu3TfsTn9nG0Vc56lL654xRurK63
mxZDWBJvpyvcxRKnmVp5cIRplLW7UrrG7KQ1gwZB2UTe58ML4UAIrufKA0SuOvnQOuxGutMM3BBs
20ILW4EJIR/JRN4qA+xmZ56M3kZoYXBZ2ALnIUW5mcKdOgrQGITh2uJnqO1gol72x97sjVCAqoRF
FyyoWyb74kLSbch3wSTUU9igYr78/HSrhiZEufpG+YPbCPQX0kG+7glUlTIv4a3G15g8Dw1BxGok
ZwLxlYsZkWFubo3UykpeyI/YQk8GtVT702XlHYIAAGwYku/gSjYaNEUtosqDiza+cTxfXRqzylSd
MGEJCZDfkWD69136y1LLd5x+G1kfxZmeOfA4b5+EqXxFjS/t1eUIyDxlNBygU1d6J3TZIu4Cvgq3
rVeUOR3runU0GbNWJdN/Wi+/8I2fm4MwNLAdxKqVpBOByTjIBzH2UI9F3pJLFXVR15Y4ysOHDZyH
jgFzMZ3Bh+///nEPLbQC7fIBlLQsgAgJAqPgnhodjd6dNAqOBWrV2IhtPqr06UfaoIKPof4L9qkH
4TqQMuXx0bp18ox9ArqXA+c1dMOmZV1Rl1IE8bPm6+xSz8g9xOk/GudZAhRk0G7iS4DL6iv11x3b
5MVcMHD0WSRHkwRxTn8mGxGfba0f3ms+FXc3glK4KAP3fjSU/QccMzJkzcYf/9utCMKTqFJdo5VZ
DNPLNTlPkiC6D2MjE/xQvNGl+PpYGQMlXsvyMlxXIYp4qwSkuGep/YmEzZJAweQ574ALJK0tQdxN
87jRftJFDvEzlg/YMexDxK0bLNttRb+JPkPnjRGQTZorXjaBaVRevpo+9dJgWNf0riGrtaM+n0iz
ucDEu4srPN3AaPAroUonaJQ87Tkl94H3a8pPLrtFzRvwAygxAd2SlIOhkMJK6o4nRhAKUl6UvkbM
OhS7R/67n4WpLpxkdSWQqEuARfov+JM3Nm3inlluaQQZmLpAT1sdGPAtAu80RoAkWBBiTYxj9+LK
xZxBCEa7AH7gYtISzTwCaDX3u9HS4wZ9JJYcuRAPCKMAZy7Ruca7HnERNkZnrqXsOPrDN5gw/4BM
oCkG9Rjqg3uAxU3GkSWcW0bdBCIOJhaA4OdtdpAsk4nAVr4g0M4CTgekYZDz71eUuc6utCI2BjDD
4xsgN2ufhZEe/8Cp65cA6AL2On6HED10Avrrhou7UM+W1rJCtl8s+RKaU0bvLdtzEBsDaRDyvYic
LfkZJGi08JS77I/l3Ys7pWHJ2cQ3b4JQ2YsZOyioU2VdE7yIjdVgyEhkLlGlNxgVEK5uXmpqKABW
WxkokD70Ps26blfk5Nwh+XY+MIbSMQVfFwt56r10XSU3bTUgin0tnBzWSpXnBphu2ZZ9PSKd7aCS
46yg1z1uscn1Jv6bjGgp498X7+X8f8Z7A2VjZFBM4JXRESgBS3xCgxM6SGQH2ygEPF6nUCfPw3Ik
IvQwg2YoBnurz7S/TU9K9VAPpsoRpBc55ND5VweVs8QrAqvTeVP/Y5L0NI4m7udeTHmT4+zWw2mI
2GQl38NaLjpiLqMIU7DFK0ADYPvUh2S+Gl5371bwRbR1lPg9xvfv78eeX//xG0o29ii+bhwem2Z8
hFqfuIEg4A70NqjUju/9QnNKoPQ8v36AypsR5RaaguEX1Bu6AFBLiqCk5B5yjlkzuQLjwPlkTVaJ
X0vsK/gRa6xrz+iTn4mVFZ8iosB8AECe4hy1U3nNyLM9ehAI1Np657zbuTKX+ozBeoKeWOzQL72r
h77rzWqB3ha7G6ChY/xWMbNe4o6fu99Ey3tGBGw7h8mBafmoVnlLfDPeR0ybY1kIG3o2vpelHRGX
gV3VeEyeu+1KIAcMy6NgLyp8BA76lwVPxHgi2QJlWLnYoZELGVCketluqY7X5asBm95o38Gl1IzM
nGy346XhdxE1o1hgrxBoTzAveFohjjxBWaYCJZW9SLv5GJe0OYkP+9BSb8ZIWa9qfryuXh3smdJF
9lRcxL6RKQ4uwCNY0dMTaIxe3AuxnbcHAM/WAk62uzfHCVj1bl68Tq0XqFxbhaUiB47RODL0NX8g
S3jd3kHYVxfrSnXC+gP09kghVedsfmTKwILTEIh20qcRD/OiCSAnQJfU3Y34biyByX2LBmlIk/2w
oVys5rvCZnpRKl1oO6uHgwqzCDQzy7QwWucQ+Ju360Qn7+L77XocgwhWn+4tE15is4LEkICG4nqK
JxOonjP5PdhNTAR3rPXcbw9+xfBAolJupfYASeJ/pSCvxXgAsC2raSg5MJE2R3GvSqfGNNYtf+Py
fABG8hn/uQM/mTBPfSdlJz2FxOeLBQrtz9EXYYiE2J8sefP0c4QXbKczKpCh750GC4O1kWHvVICF
ZGQRHf3oGsennjbclOel4+qfJfaHlL0bU35p8ZvftgxJjLFx3PnlLI1RlCeyre/4pI0nwe0g/kk7
LxkZMUOfhoghHzPCTQkpvRHSRMn+RbRo8Cq5ObK68cjGCT+8g/Br/MJsJTJFlBNUYt0Qh5dp1VMy
Uya4LptS7+0533wVNYGz1MRp3aJa3iRzrn0qFu3IXU44C/0OKXNia81f0CZmWhvR83gTFpRrOB4n
uvU4gG6ji8se7jSGV2rPpjffctCyCb/OflWvdJMe3zwsL1kexCF1BioALXiiv8AMo+AzSolbB/zB
n2ez/9clMH7kxB0MgrIRvjKUcSdS4gCzKlbt9omh7lHKCeoKMpuPy4WzGihqyrsbu9U1gZyyl18C
5OqllLjGs8z3ejZLLsBCeDWR1JYHichDvh2T8EgkY/xm/XfMwxuh4uT/KWADNyYjMXuBpmqj9dR5
DE4tYmggDEKJnkWN0tLY0Nnabw9ivgXOl4QBseUQ8oZWnaVw1H9Nqzgp6RZmpsVLsNArhFp+AXNs
nGfwz3swYW4EzVyZwr02NUvmslWGcYggnL/9LFdKSS65j/PcZ9t6183D+3jYvHmu8OwAYEEoT18d
sCbXRNOQBVybdIKH52fIzegq/MXvRWCY+bBYz74vvCgO+E1heuR3i3Z58zDKT0PpvsuAWyhOncWo
h/3Op3ZxRKqwJixohxZtVnRJ1Ri4Ey9lhRCen0FOVkpPVPlLNH2vVKiyi6cnZtM1S+hfC3nmVsUv
1GzO3J9W0sULzzA1gKOuDYJYHWzh+w3ND7X6L6OU1O3R1a1eOJt/v+ghZCn+yXj+YMnwDxZ5uvnw
UIxZGkiK3p9fHfwLn0mjLkFaHk7RNf/APvON9EG/NG7kZ3HNZrCjOgw24nXWV7PZ5aMd03iCvXbF
l3ThEt4ZPWvGiViXrL97vP46C6RPEKuOT8OTmkwN6vzxM6HC00jq/QXEOInJQli1TSldFcUv/6Iy
1b5t++jkSaLG04D5/OxIYfxQs3d1p4p7b/aFA9QL+X6repsF4IZYsarVGetr2oIo/ycYZvLJ7RcL
tXtAgmRCh4Cn/PZO2ncClckAMB1twIVJKnkdW2FYsCYJeQA9gS/zqJDh7k9aueKz+B8bPNZmpGow
UE6Kg10eFlJA1VqieNpjh01GxXKG98hfDcCLge+qaUPrdM6YWv5Yh/g6aSlTQNat9ZcJNwTMduKx
QhMNcZZ7/AyxKOsrYDja9zQqRWpCsKi4JVcMxtAl8u0QikI7eL+P1qBSrp87dT9GPcXxGUNwJVFh
cxESwVRpuuqwqKYA8ZyYgRhvUAaD2dm219+L8ftdzBBW0m3SZ2cgr1dP8CtwPfiD864xwBmYudIM
16CIQXA8BTqM0VOoBCfquChqqUgA0LS7FZeW7GkJMuC4CY6nc1dJfvTBGToYTTwPIFKIw2j3FWey
n5dd7OUJWQHgBUmW2llYvKxJMjUuVXasWmdI8BTE/SybPFjg9uVuKHNPs064Wp5rKwQu6YAcJMjG
9oDXxs+3SI7h0Z6PM/er55uJKxzCnH8rkTzJ0GCeWsgFX21YkqrwQDc+ObmqmtCVbLn40naDv8fG
nnceg1+76xHVYx0qwGvhX7c40szZ/X1FB3OiuwoUPQJnUTqtJOzcc62XSi3DhqpxxFabKBtl36t9
AC+Dbi8akUF3WJwG3dHz5BIhrSJu66f2Llu+kHEt1ufBYZGiCMzJrUVrbfTdDw+J+2gHAhleK2v9
oyPmTFjMfuWKQScdDphCEBOCxJ3R/5ItwowjzclrLdZryVL+UwfimxFsB8XE/gRO9EtC8PwxeJls
9AGWFsAjsnbTQ3VCfLAPK1634vgJLCpiVzvRtoFWMaLMGyuE0GJQAeRRl8mrMRP4Dy09QaBTenik
lN8aWRPzYjGFXUFpKFzKHoQXRu3sqz2R8X9YzeJmRpFgcNQzYp1UvKeXDDOdyMBpUObJFYr+8DGZ
XVB3pVPjfrP7YjU1veEWbChHc0w81nYhLPQGrTJJTOd5ygi41J4PNHRNOwTZJKeTkjVvBFVlZ/yP
aHaQXJCjOU+0+dKptEQvxcBmaf4rmxZLlUbmKtjotNdAww03+wtDUpmS7LTxeRPFLroGPIwcl1Gm
J1fA3w706rME4eD1V8LAaaUjvJSPa7SONyzF7/ijZBFTWaw7hg+FJVFkSf96JG+1jtjv43qrazUu
CJbCqhru1q9/Dft19UUm+Zcfg14u7+z3OVxnyBZ3F6IdFl+VFDFK/QtaBfMRUQ4a+3RSnuGwzrE6
T0SRCghNbbmCeOFBlNxHKxn1choJak1sdM4EJwt+atUtL+jiLqkfnFSvzE2xpVBnlxRy6Z4HazMp
j/k+2Q9ysEROrKgQrv8XDJ/5Yx1ok0KKhG6iC1JDIuBydhylRvJh2iQw6l89xEFQmvHK28Pta5R9
ZLzwmzOUbySHwxpIKzR6QY/GcxiUFaVAxogAdnWbCL/bW2Sn4yzaHa+opxsxXzCZUqE7vpLIszOi
ogLOvVEuFhT4ecz6/W+o+qfeG0h+JemjN6DJqrHJ9OB0gFS1XZNWL0nqgI4i9wuVIGKCEkTF7Svs
6zp0ku2FtXHiVMSZhB5V7xpUrKcuyM9w1Ms96QxuHYV+I9JH4tMMV0mqYf2nFc1DS1WF4kSQplF+
VON3qK4owbLJTGy4P4kxEMu4fu5+Ybj9NGoI0xS3f3A5Gn9+iwgdetHuFyvyt2l5OYhjHYvrFaXl
0qcUVt/Qalrc2HCp++0DY1Y5b2SeHhhRwH5psC/1HEGUXCGav96npjdatny8Z2WKxGnH1iT6gw2y
gnNwiVneKJyX1p0In+Zx8DgOoc3t8j2Gu36g3/J5j/x9Zfx/evhmJlXNTNY03EMOsDl3KuIYrXp3
YAsBfqc3gM0WIzKcfho/9bU5IBceqopkXGaNNUTzK2TiDftPiCTmVk8kh+az7y7SiPzl/yiqppdl
oqSXqdTFKjiSgluWBjE/vL0eMKpxbNLAhPLNRtXq04qWAX+rKmDepuvlQLhoQVt3moBedkrU15Cy
GsPxasONVS87Cm77TG4E0lobbFrbVBiy8Nc9W8oy2y+Lb27wBFpKntoPQUeJ8+S1TL1OtSfwtLsv
FSUtph3TpITHCBWLGZQ86YyUy+nk1+6bgEzOJtrpo6u5j4OgEkgNdZYPT2u1p3pM2kVipGx29lVB
o8UJfI3Zv9dyo0JvyXLA9u+X9JPSKhjQgsfAhYws9dQWkvoIW4S7PorQE98U/8LAbZ2M/iYqs3wG
QfNvm0cWLKlZVXnd+o03I2kT249au89gNQ6neVECH6OMWHEm8PQ3yFkmXoFGHdIlPouhGYJKDa5M
0pUkbkFHzn8QX9lxx8oxrYoZM83zTeJlsntd75tCs5H062tocH0QhabJemn0exKyorWfHCDYDU65
CMBGMswOo5+b5NykAQHCD89F7SfZiUql4j8XzsdZF3x+u2wm3BDEodTl17kReh4iOUb8fBO1TaJx
mvmUhhi/iA+AVNcgSvjyk+IM168S6vcsBgDkltsVm77CCFT2qwP04CIPkmRd0Xw8+Z6/V6Mcy+4d
SYnK+JgHeXlxhF/K3wTVwd0QsBxv3j6me5mnE8fVZ+irZJGlobdKWDbXgib/yhYwzjjhL2iVytqL
0j0NpynOGsRyJvfgLjw7p1lYeRCY+4Xy86Q9KPikv8IbMPBz/MQDN5d/T1ztT0ntwHi17KtLYvIC
4jc3AH80yP8Oysy0j0+3vgIxsuBm/UjdEREqO2+4gtHpb+U7IOkTjze2TMeNiHfxIoD/k07Af7wV
u1kqhcBxrT07virSoGw9HHL5YKc5+dd0Dc4zukl4VYKUmla1dJZq+YnLd2OvYb52Ix9wIhvFaXL/
c30uetQU5Kr/iN0HWtqup5jKczAMxKWVICTgdtoMCIZF3VPmd3wJDoSa1igyqEHajbzpIzf3bvgy
TPhrtZ2XLsC5CdZp5XeONMl68bUMHNNXH/ujWzv944cTutB0NuL/9lF+uR1MpQI8RP+WJm/J0ZKi
YC+L2xJBbxUVXnW9YZapjoJkISZT7FdnsXMgT0Aa5iZfdXSMTKWrTdp+7c7BP7JK0HQd3mpKmBnT
Gi//Bb9KcVdFnkET+S/4Ub42pkCPJAHOVFK0/QAgKAj1CNuZkvqN3NFCAQXZP6oj8zwHBNy5Os++
A4j9s6WD1X+AZuxkt0J/aShQgZwwW7p70duX6OT7/nYd7eqfjfhFjHkl39fTxNX6sTVN+jZS8881
Jc99b/lZf+hexlxth55Ru98bH24iT/tsNUlgaq5LJBIVzetRhBfdWdBCC+6GNU7eBezCjdzljXuA
ve41Nbtg1wH+eoNcxIX6QBAS7T6kDERgXcke72xexPuPIx6b/xp5xDyHT9Ehx3XPeidyX3aoU9NE
71JlWJVWPmFFbXAR0TR5Wmdv/m0S+U6jMbqAs5T3gvEKVtx6xNrTtF28sEmqArjppAWnAmZQrn1E
tGf68boLB71O0e6nRS+WkDGtlzgdzZhpbnfjGy3W+y8Fi4SKDUFRZ0IWRiqobscQIeHFMDjIK9gC
f6sRNNZWv7wS+LD29Bw2Din2cQ60UPcYpQ15mJc88t87ZQJMUErPEBtUayj/gFhSlM365P08tYl2
iaEdBT5XPn4P3E2FsFO1xeU8sXJpZe+GETa0GRPuEP/FTtLtfEWEy6KhYTHHveCcWtXSSBDz4zU3
BXsfJ6LXVqMUWIUThsrin10Z7hpUaYlhzke3WlkjECuXknbWaSQcfXfs5+EPMKNQpnZl9fBulzfR
gXzPEb8X34Qjo1f4nRqwC4gzN/MGN5XwBn+VQoLrK14iple1CTbe9iCvl1cikcTAqdd5aEqGqdAa
K8KhBAsa/4tbKCncBYR6X3AsUpqiwKSfMYtm0mnFOdKQWj8W3Za8quqwXFsiD7Xi4NmXJa8PfqJ3
R9c6El/KU0q0EMGsyNiLcEhRQaBfBZpYrv8pxy+k21PtXvVRaXKX8G+lyFRdz3ZI2gKkJMZUy2+H
TPxv4nPyt/TyPHf+29Z+21AiwJ+al0uHhLshTSUKDZXriXwzkxKLhx4pzt1+bgkJxZLOGQlPCK+I
vtfwYwVT8xAZX0hkPIkpzcT0sW4y8Ap8NSJDWmpBjOp760uB3kH78uGNfQYdsCwW1N/76epRLumw
4Hyb0A7akVyoj+dlQQ8OqtTKzsoubEvuw+ZW8ikOdzijMNO0A0DuidsYuHm0zQfZJnBPkYX+Nzsl
bIk6vhEtkpTzGSgjy/zKbWh5n7f33MSN/X202FRWaRFGw8gpMLBiB1vCfxFyi41DVQuldHw/RA/C
Seh68hejTyQpQ6dcwXPIOXekjHSZswzwyZydfQcwkGZLD+/OIuPgBo8PI+//Vtuk6Cvl2BFLiekY
K4cxFulZzRJ1xWTsXQ5y+K9PAS8txj8yYJ5EfFv4A60KDk1odkkU8uodig4jHdEKYUiva2643+xI
OAJDI0cJBLxMqgQncdo6kRvPHgbuUzLhYFWGE7IJt0wpu4z+e2afgx6pzjILm3vr7SIsrSCT8OVj
b4/V+jyfrfd9gcePWk4uR6ejeKypsj1Z4zrjhyepKJe+r1UPWB980cG4IlwKDkcv62Q3WqwSqQ9y
bDDXedP+gW1ZIxHoGRNnTGPxDB+/vKvBsBhWR1s2lipIi56PET0XaBHb9epB2+XJFH0XCOnK93Lf
umA28Bc+LbGEs76sUPqgKSE7XZAyl4KD7cQ9kIwNm0WZ7PUB8YBFyBw1YxiM+esKpFdCgh8VWJYD
EgCkEtZ0QwJUBXDRjItlsHXoVTuHNfCmPpDTWFXgYmJdKAdZ1liByRRzgenMMB6L00NHF33GWqMX
dBBjXh7A1zZGYwTHbFbvFkehSfLSEddgVtnLtTEDT4KQ9bO7SlmU53HSwjZLdE+zsEHxJ/GCwKNl
cooCC5NpWGs77DEdDrX8BGVV9ujRjzJ/DX6hSy087AafWrpoEIt9q59H5pmWJGjSLG3ZHYuWWFmr
T36mDEoPiWE1X6aGv+KdFHjJRD7L0aXW0IYN7vXcNnGARHQZ7wb1tAxMF4eC7ZxiL5WZ5Ia+9Cm5
PGFE3avPJjEoxLb+5i0o1EwK4jtJ7mpesgtoyLjAPaRP4OatvE6xxR/+kgqbhhW8ok5pPvA1Apib
kPTQjsvlqBLdzc7KprxAEhGlaM87rc4MO2ziyN/TPMLP18RKOWQig3+NE3xvTlt8AO5X9WAEP84S
pbS8n3KqbUftIx1lbeQ7NjGE/M1qJuqxGTme++iRRir24LOlRuWJu4/zXCSobXmmEPs3Vtax9zPH
OuNGoY83z6Dif8TH5pxKjv56qK0V+euwx7RD31bQLQQILeKsYpGA45tXZLgs29dFyXsKsByVoB/Y
DqfqP5Zp7HGGbrhHWq9hG7MZv9R/Aur9zzsQ8aBfBERCbJmXvsRLWTYyke/aaq2SMuEVE88XrGUe
sSC+Yz9nst75mkMe2YjtsJoZdm2q4rTnx4NnVOvFNyjIzzvhtJk6SKnRS2Z7muLYitvwpjENPR5o
nQ3TGIaSbLKrrJn1GLWYVVzXP8/PFxbWFdoyYmqY97kqHWvWadRFt2FsMfj84iybXtkCBWmOUAGt
mcJze+b4uTKcMZXOGuDa5b0GexaLOpRjBss11L3zaQFRhrLaJOho43V2hf5iEr1hxqjYoQd+3XlS
zl4VGkmZm1QDCglkC9aPHZXHQRjPHj588C+AUUOayYbLFXuhJBQ6tygdpiY6KEe7fjIfznncywdI
CIAMPpnZUnvqsefOK7QBE/U1h7vrPql3iKqT6QQxSUDTiT4u5QFNf6HWI+spCR4LfPZQzzQdGE43
yD38VEy0j0dHqRQCb6O87rrDC1/rEZcUqvRAEfIXZ+MlgRtbrMhLLwSEDvlyjutgUtBIjyO7L7Ep
dfnX+KEVDTXq+RJTZL6RpHEuzcuFsrZ2fZcCn62e9L3NB5Xg6FNvHlmCvnV+6ZXaEUo9991knZKH
UilFUc2fjQnrJZMo+sjFqsnIJhC4upIX9CxXZfDAaN8irYfT5NnCbSsKHBjOLI9i3FHBlSyxez4r
oxr25vlKRD0FccGOfORsh7mj+zXN9WckL1C1DRDCrSUFXsE78Ov6oRAtayLHOnTj0Gl6YpOaylhJ
kUyiJFOz58zz7nSRzHQJ/8/z+mLSJ1Axvh3apufWzSKnlzG+zv6y3hvD/a5HZL4RFQesHxVWO4hz
QMQU43XbPM/az1MMAaSr8HiwaWcQtnkY2K8uR+enWY5bkuFHobK3p1jLVO3jf7uUs5HzZ9RWOQhK
NZrpFg25q0LmEfA0rmMKujdMPy6adev4KvHn+WOHSqfd09wNkrBwAnNo5xg5wHBoy6If3SnvipdW
4mnwPn2InkzK8C8A9cnxEgEInBH7rnH1b/Kw5DcX443zF2lBTT2GUxvl+lmqA7j2uYecBfqEu69O
inpylW+JdXIvisNAFL0DD+bmvxKdlJGbGMoqzQzGidRQHreme7JU7zhg0xF8kdLTdfDQvtBC7sAM
4inrN8c0abuVX/9kz3WoSNZayGYN1qpJsWlMlGASuMM45f3O4GSsV/StUlM6ACbRM7Sq5d4wQ1N+
pWAtLJS/L0uqRU6e4ufHU9vSZaQcU1cgwdI0k81efhn0Ql+64Pla7TSLN1jWBsVZOitWca4Ipzu8
XnZ8kZXdAU10lcfaYrJslJLsNvaR+217cT4NTZesZnfgSeyFq1vdDyeXN3OoOKP7a0ePo6cqaIF1
dXXgj0IniaPowP/z324eNSstatbOWTRS6t/dGJ+HgmgZIgXEiD7+wbJj5DevX2kKcv03N6ZgXHQE
SgnGhEjlSci04FTgIz4TtYUtkmYE6pwKd4s72aUnBg3gYHjHgWjxMtFjwcnH18sT+uRYuX4RDWu+
C60FQl+r1hIP2rc9Pfj1GzgSv5RV2moZlVB2fLWjB/SHphHTcHvH9czU2TNFtyH5rKvL8L8mx7IU
PAW8d/tcyj+/bR8JVTgGvj+qPNVFTeoSl6w1DJqGMpakGsQujGuLY3pulz0QqyE3JsyDZKbO4udo
itD0iROsfE8HzX98Ihpx+V96lnPS3dD7FgkusaOPwuevS0xoPJBAe48G3/XgD5VTNUhRIJdo+KmI
eUjHpgA/2H/u6aZ4XaORqPsOWaZ5wm5HOq30bn6BoMz49EJrK3vx+sjCFLvd0iS19N2Y69KwkJ+e
VYwC28XHBQ8gNrF2lNQwxUy5Im2VT/C0IlLe/wTqxw+pKtTa2cNPgjMiBlkyuFMxwQX2DCmIzhOP
dojSNBM6iuM7qb1MGo6gWljy77oz32aFSMC2fkKXiir1XDuyo1VVYo3/heyqtVYeqB/i62vl1lTS
+XbqEFiVxTl+6uyRsIfuYHMLZIMElLGkZrQolV8MhtBgfInQiQs9g9QLsRbid+bnn5OhcBKZKGE0
/aJ9gf+td81F0zWEWU+R0aFKh0VmzTK9fg0zTndLyzPlsB0FVGF/+aLtY5fXIdz64l/ZOK+EvGp2
4v7Qkym7q1X4k4VakFlcYrfsJk6GMkqD+vtjHHyhsBrExQUOdVHPqKpcNg+nr0Rhj7xqPZn46JcX
g9MpGLiuRVo7VE3ZDvmzf3kMCjUUVmPWO/x6cR9xdHaDZvnwFhZ6kowRSb1xzzm0rNjEc6fPmSpZ
+itqDDyDN8Ug2DBjapbacL4/2o8XtEWJwqcJ2H0ymN3qQmxOstbKbaundODlR2NO96oVDx4Czi5D
T6ba/bDJGJcfeQvG1Q3UgwsrjTVbc9elaxz/lOOA9KcxEjdLULqh7svmiqIwbff10S7+dp6CV3Or
TSC0e8bwWlVdh6jT/XS62nKGPH1EPxuJWWo6JvOJIXcO/zZdGtn7FxBO9uMjhJbuIWwR1KidwkSs
LBopwa03eN2D7/zlJ+XFCx4ZtpuB4RofPEInqdQIXBQUVhWG5q0WrUJutNhXjRl8CNQrGuMbGwfX
nIOfzro0Y/48x7TRa21cXOtuXlsDPv6+ukhj0ayOHqFXv13fNP1quG3QVoG8B5VYueZKJKsIcG0L
MRjVXsH8+TT6F4p6X27CROIwaWFEwufvhpuB5EYMaCpPq4L/M8o4YXYegEVytQiT7vV5SqiRYpvL
mB3GfDrpIgo/uZR2+pFfN13aUu7+RKOg3HEIG7sx6jQp9ilmzhMTVqdlu2YnSl9GtLfb5kKlN6Us
JGyVWBkWV7op+f+thsx7mBrai31cUrVLotrD0ldBVT3mrA7A0BgXAzk5iivlrlZj/AZTc0w4BD+G
DdGgKqmnlR7cH8k5HQ3fSnrxzGaoQaxk3l+UvJGaTaQusT2fKRZKvBtLlawRnCASvVMoATg9is4P
WoEJzC9j48avVjB5lV6k79/R94xgP00/NnbFuMjOAiZXgJgOUFyJUyX++QsDGpPoL/ZiBLFObz6+
deMlzbWV1Nxof3e3Ly2BrVnThW1N8PaIMT+VGX0tJWLnBdwueKoMnPZ2seiLm/u4gONJjCDNlNWb
NNeBw7yrQp6MMFXpviFTqwgLKZrRY/BLJmLx2YeGjHks+ztMUhJtfXi1d5hR1C8WW+vTZ4guVad9
+TBOFAJUlga1CcBfU5m+9tb1Jyp0E4INUpQprB/K7ScfqGFVUDIvFZcuTdtHfzLst8lrKV7RgyCo
P4Awsugk6msCtVoRoatWqz4p1PRezWEG17S+vNSvh4gf/kgKzqJWvuovG4VcZcK8sDi5n5Q/bKFQ
+xbiqZBblixINb1DN3PS1WY/FBfVl8yPfuygOVFnN18I52ZbjhMAczmPj9QYi1uJIl2anbt9HPNc
/VCYggKtOBIgli63XK2iwg1l13sl6HElUrV+b5uhSt5G5kj6ofAGamfvJ0a5OPN6xFrAS29F+mzl
KQ3wQP0z4Qnph6d4FLZrc71vXviYzCiNYTCem360XzGeNpCtz8oTPOHq9+im1u5UsZnq/zJvlvvF
4ZPhCIIMYc//x28G4iJgmB+obK5UBwafCn8mACjPYJ3ENB8hKi9x0Wd5ur80U1AuliovFTr+aMnu
s0+cq2+GrLUKfSzOf1RnHYEfmfSQ0eoDvMqJdnCjLIcr0k2p6cztbMpKVWogL5m9nvpG/RIM0Izv
5j1pmxnB5ZlIcPn9MCAVrncZXe+YBUvveHJAvJEmkJXoBi7COZ3yWbWHnvsdr5peGvhAjek9fdgK
eiyQ/eIyF7qM24WqJXuRZCrlUBQ6kbELJhKOXxqk2Glm7tlzLntDkti9YbsjjdJXTIECms+BeZMP
OmOkagNdEmVeKbxV6ez4xhBlUopcwLTAMGoyBfdyPt7pO1YZsJUmU5Y+ZyZrn8H+9+zLCoDWsuGk
4prdkG5SGCOYiBLkaKfEGXec/7y7ec5KtaE+UEt5QDfwMPvuewWAJbqgUeADrxyzMJUawHFW6GaQ
oUqz8nNUWcUkNXuhzjzdoE4LVAyOKC9Uolmjw4xgo5LdvdYY2C+iZr+0SJ1lI/tv3ZMkqJbsnB+t
S7jmJ68v5/HgJrVJVt7WIvDye9IvD993d/uEux3BwtNuuuyLcdNqi6lZxaQzb5QPe2RQ2ewXRY8L
hkgFz/gcPkaHovccFNh2IHX3uQyTLJcUQBuM763/Q2DwgBapQ8eVp2exTbdZNwej6z6ka20xKqQa
bSxpcZ+owRAhhgCuLlHQk3NdXbKLEFxjZKIhUcBLeDKcDOakuNnoV6/JYLQU2b8z9ysz+k5liiLd
bzQKaztq7zjSrUJVNT2TuGq6IzD6rnuuxybSfG3FpsLLbhFeZCvwCf67upAKcaQghcONDNM57MfZ
3VTyYTS4mcLw2FfXBZowaUpmrwjUidngQYWVn7Cn1uxxcruD6KH7ZGkExOlYZvrI9rRhULeKM7XI
7LUcW8Xl8fCOAII98Wi+iPvZYi6H/R2CwOGix13dE66JQtrsBMxRj2Q9i+D1s2r2ToUfu1vdoaF6
Q8gdIeqDyZ/0bIhfHaTVnDb4puPcP9ksKwots4P5D0tZxnycZGWdH7RCxiSnxsw1JnRx1CHpKDeO
Z6bjY5LezOghHX6G2eRPtMWWZUr7YlwW8kR7sAqkSL/i7uY2UhLRtI+xGXChObU1PQRbv2Ub61eL
57l6foKUtjbiU6bVD4zspnvRPmycCj58aopoRn5UXbTG+O1/4SL10kW72P1BP55qKWKzRN5K2awk
nz+X8ZJZvMp8BW6fnBadXVk/N8sW18NAqjLLeE6KDitFjaewTjtmkWv2TUWCfd7r1RNQj5v4dYvy
kLhbadxAGIYISHpCzeX+yVYsp+aGIpP+YM8lOnMX9sFxZ813X/3JKGsS2JS/Ds/X/1vo3pilM4AJ
FcDIyK3BFsasNe8VOVQmAgb8EENxylDLgrxpCxAeyNS5pomgSyBu4hkFrTk5z62pox5h4N0P3KFr
koUKHPnaWgPvaxSK2i8OOIplZnv/9P0KCzC5GTRJw+lr7Ehf1VTyYcpYH8pJxlaJbR7OD/ikPBLu
6r4BNCZurb+Zr5QLi2EBlYLp9EivdD6SJW0F1VHkcjUvUVa8rQDQPINYK0Ph0NBaIlscXaPHV84R
imHyaNofogCDWTQVd/R1luzzKVeaRLC6Jw1eMUC4eQ90SEaX1RgCgM2/tqlNwAWX5ZKg8Kq9lbDl
1KRaE0RC1mT3pGB40Uh9txbMetdiDEArQyPJaJwlFliyeN9ncCUiwb74zUXRiO5yc/QzOS4JUCcT
8qI54IwjnLQjkLCgX84yzM6ENOca8PMZet4f8nlgIdEfbzY+iLfyLq5ywKJTLfBJbuIBmieVuOqC
tejqddQuiW7DXE+C/8MrvVJw3+7TU7zL4+afCOV3K/YAqvoCajDVGEHZfFndsE5IJC48zEPGh2Wf
wE0zjaEapmprI+l5+AWKjhXGXA65D79kxtAmuR8vhG4xWTiLLUCWD8mxu9XK1E3x+0ylHzH0bbrc
hcfoZn2yVmswbmGMXE9fJLkSdX2Nk+6H/qQGwDw8c5THF9y5fUS+vyTZvlBqrHNCQqtXFTwb82jX
NxlXemDyCXp17cB24klLyKGu6Xf9gX7KzJXgyLXUsOMUt3SJENDYS5HVcZI3R5bQ2ukHzRwUB+Y3
edtx4O604s3XpcipRHD963PobGhWsnzvGsiIiy3uPUs7ry96mxTb0LpCTZbQGH4ge9A0fyWRlki/
vA6dI5Ms6g7gsUsvGulxLLp8WHIMISykEP5/wNNM3rRaPgJOFfd0n8wvcCTDi5lhDAb26tQw1mdG
gK6VW0nEoCiXaam4HvrNu0aQNoVawyLjO2jkAbpqR7nWCOKihU8BRT/2LKwqOwzLf6640VZU/Jql
NkEv+cTSBxEPudSsTqP9njMPZHuVyvK0i1ilg2VGTNkSehWOi1RSIzVZUrYYtfmIRC9a9x5QvxpG
qXPPTClXjLR7zqRtHP3rc49FJbg3E9OBp7CB9HGZX7lVSTSRvb/cEUgZQbgThJSxAzi7ozsOTpNQ
qELYTrcXaB56CaNobnxy2kMNsdirigqcPRCQbDUKxK4TeZdHKH+UUdy1C3WzbKyUlV65EA6T67Ie
7B0YRNkha0hti50jqj4wWmwuCxromGyuB+WVjQlp306b7AgHR/zT09/BjAVpzMRPig2cX9LrBoBe
T92nar8BSdinyCzNzHU1trkOF6W9SjFgXdnfLJ1+PYroWpqLrMnm3v1LCtrs0nNNUWoqx23hNMFf
KXg0aEEw2lT0Nlomajy1U0tILXu4XAdjUlD7KpXtZk9l618EmSWUo8BzAmoi/f6jQf9i25Of9Cr8
FRv5hxwRrr5Uw0LTt4xRRJjOUSljYELAEusC8Gw5G7iyw4SMneskbnbA1YtpXiZKCxBLyxRtQC9P
GJD8XL8XLXGbj2s7x1UcoRjkOnhDnfKGPJS62uX+Ng9gdAx3TBeveuLS6kuhzsuCo1HMPdabPPvo
s2WIku+f7ATjc4Ojjz84QXGUWm5kWdOOIKZ7MkjcMcsRXSB3crpj/0kqERJXLuLnMWOr4ky9F2hR
ihrlbh0H/TAD7C+ZPK29YZnNxDm4akD5Sqi4QOpYYYeferkT/fra2OQnbeI0pmVVGmmdz/z2GQqK
ozC6o7tJwcn/kK0SG4Niyo9foWhVA4EToE1eqdVgdGLqEL/AHTfADV9qT84h032IM75crKG23efo
LfphE3hFgxZQ9HxmyS8+GoCbHy2+enzHSN0o98PY0dLQTlH7bLcMN1s95EJ1AU/LlaHdiJqjbs25
VxOUVK7e6lujP5I7qhRi5agpVyjVxozw6vY4vmlWUqg7Pq7KI04ntaYwP/GUcIW8ko4UNNiYCoAe
pJ/WJr8MQciAL0gLtd+QqAarc/fRl3APcycHK89ImwyV1OelBN1H7S9jVJ4jrQvaH4WD0KYMLlbZ
6JN5LIFhKyPebjJImzssXcC5j87yCp1b896lPgHy/HWKUog8S0DO5tC22yB4o9az8iX0LacEl3ps
kNMwqmGk2Krfxa5ssCbwcacsozg14tXEvUCougFLlqR4ga75av9TLa53mwK2HJkth0NslkCteBg2
s/hg3h/zaCWWSkWswYKDz1pIWPuG/ZXJWskNQqEi43mNhLgIKAN6dywqWBn8uefW1FWpSeDudxdx
AhzCEm4cdrCBdDzLDy45PRUudsE84xoPAmarxUMdCZ4o+HlJ3gili9M5jyK5GieJSHi+dQccG5my
SyCXDHK4lE8vnaE8BYEa08XW2xipa43JUR3VT95JFVUa6eDNqjUHF/2GKnw1TGuJjXGyy4Rv4d7k
nhy0PmrsPZRdTQpw6ZHBKvzwuuCMObYnNblJltjWfVeBRcze91eKfK1U7Bm5p+GmYFvx8YY8MXMX
T3CYcTgdXCpofPO5qleXgBNZZn56SU2hGkKushKTpgtYj/LAopvVM5EBO/rw3W0Gsqlf1ocQmvIj
E//y0tvOyGXKMy4ISaGQY3Yp9YVUz49hP5lxT28paYBRKbg3KhyA70//Vdk61ZiUaKtZKmNRbxVZ
SzcO5TE+Is/CdF9vTPNQUDyUprzVSPNmX2kI01yBmAPfHNtrmZmk6qcSU+ot9/gwqGBn84OhkzA+
9TWfqYmgG5kigOQPEK4Faa9pHXatLMk5kT+Ag0/hFHf2JvuH7snTZQ/+yT2r59daIiW623xxEXzF
scefhE6zZ8G0XwN977VRhLp9lU3SMfP7MW8D2cZYtl8gq8j5grLa/Ve7bd0Rq85uBCGtbba5Miu0
R/8IDNRYlhiKxThu5zFsrvpAycpozM039yYPIxW5gJH4VscI262NojopBlyjTjbfS44iK77y+eMA
SctC7yNrCD6QFeG4xemzTom2csMHbRb4GxLmQ0bBZVzq80TyjqHbg4WdN5RfOOt8zOfJKCmUn/9b
DeDhHmJp3nhIoLtT3W63hTv/PKM8vaoPlgINnDailow+eoJ1PjKzU8f6bhIyagl5EoITfIn7TFxB
6XIaicYj3GrnXEGRUqEx1T4Uo5oD+X1oDObw9eh5xO29EOdzMvkjDAAyWpG9MxxaW8kZO/Nsxf1F
WgQttOMGAmS/naqpXd1w15XVRw2ds1gmgdjxNImgjuirvUS8zNWyz0foEmtbKuOp12lhG/IeXBi1
bkZ/kNRhYL9do/co23jCQ7e+0bTmP5MTnQrPTILNCNDG/3xX1NZPbY4Rx5EvsVgZ4Rh9OLy3EMsU
j8G7f3chFicRAwjWiizRMHHaCq60BoIGSv0SgCPt8mNNwCFz1Q4/lgy/iF34ET6Y2h1Vr7+ENpyG
HkTdYaxBgGdXbBjohrZFsGVieAaMXyJrdMVhpUkj85TEU8mLF2UgScClCKu/t03NJiilLbTvZPdb
McUa9ftEnDI+/V6o4zLFFj0gT04mqIKIvU/axZcWh68I2AR4BWO6wATQ5oqtoiQ1TKqzMKmdnUt9
0x97WkTTbqia8HN0K5cIZ8NnrDHiY/dfZRq/oEq53JQDERYb60snAlyleaulQOt3JyKPl10UHDw/
iDbCnu73VIWlDsyoBdP7uKwguh6SWy4oQ/6OhAteJNMcCdxLW2Cza2jGkhZ584kOmoL3I2BhCz1g
MtPZurzxCXxzVUop5IfvxhNRU8+9fEmmZG3nRqzSN3XNJZ7rJNtvldGX+aeh7g+BOzJPn7LyWQB1
onmNIXpNl5YFv/E2+217lZAb1f3D1TYyce53wgaKPlHbhyR39aAhg5QFrN+lq8sTzcrzCwa80ZqU
TC4fiE2DkWvaCcv6o4XPOBoS8iNM5qj184xTWnU7F7RD3OcB8H+iYkVGWdiY1ST47HlwiJLND4HO
X82EZ/HQ/jcMNCpeNmi0gYfHI6iCtVtTk8s0bQnQBkEPEcQzQUZ9ss/TONeg0FqFGGI1P2VmbcX/
QzOIsTFWtco2afQT9bveHlzgBcSN0TqRNs1iE2zvWIhUMNCyVqcY7MpIVZymKKp+6q0+1P5vnPv4
94E/C5XeArUxBLP7FoUUylyOq+nArL+6BQQlofBVMho7FBYar/Zzv2anP6zhOatmqhoFuGcL7uKm
rETqPpl61GEXl2Ao37JJyxoW2zxLNgKmRelawWBVbVOwfjY/9UzKbu89qEv3RQu8o25XvQn/lMIQ
RMqPZw9fIMt8w+6KLG1ZgwoqXeXfJfZ83CvIRw9cyHFVORxreyT7Y5LQjavJJRNF7nGtw+vqv1Ut
ubm1QfBz5o6QB12wfh0dff58qQTd92r2TGAdF2sOCDA+1fkbJ7VnjhbPIb3kPO70eo26NDg+5S/A
AoeLpZxOH2EKW3QJAidamzFrnHF4Zn5CbO8eITgA851Mezwr4aDejYM/vp4/vJkYdL6XtyDP9dpz
ZcOVqYsiJQkJE6L/mPr3z8+kMR1dOPtJSI8hkX//4LQoLtaL97zRW+z/Zmn9J4PhZotURmjvHos+
j1paNHbBIINdh2n5ww63GmLGDV8WIHWaH3F/a6JHbTmWYU/ZKOOGK9UWPq6IBQtT0xQEl58hk8PI
m20RHYbR1Gfcx0tSkmVXnmXj+vYXKB0EkR5Hyqo0ObxgZzQr1yuR9usH4xx0VM0q8dOB8FUJvrUU
aljFWvWyDGYHch/HzyqVdA2iTp4tg7bLPbCAmApAX8wC9oN+RseVI+CIDbcmUP6Ttksltm9YJOo4
3KMdrlpzbdx5KQXOMCYfj3XHI8EXIMULTX1oJZrDWOVpJfW3ucRVWop55dG2UyL5XbHpURaNDVz+
vS24X2u2vantG9mAF6obFhUD++kJ0kbqRRw4d03Ms9MUebFleRKgr1eG/RXVEwgZnm3Fp0jNdfnc
NQS1raPT9e9t5OTeAzLuTRo3Us5QM+2UOzmxHxTx9JZqmmiILcaJT7F81zF4fpfTWVZkaceAQRXb
cddZg3WW+x6s03AOYir5unlEMZQDxDueZK6awamSRwX7t3DVwVs2moEaYa6r1fjdOm2ZP4Q3JB/a
97Bbq0rr1KHQeYle+W31vQtWIQN5PAnBjfTp7DKlpjhEmwc92pnvFradR9y78yn8NCT5cyMlmJyN
6oHnanRHlvfuxt2szdqP8aWyFHmABFt3UJsroeIRo2Is+68ot/CROlK3UE+iI8gx4mAFeoIkKQ+2
Jwqd5REqI4fbgnSE8eCT6yy1HgMO8hvwJbVxoHtTtt26BsYmiJQwdKJFon7oYesi7EWgLM1tYwFb
LdP6zyyerFJ9eEQzvgpKila9XL6vigBP9e6mVZpi/SEA76SK2xa0Q2S7q+vTA4yv+8UQjMli3k05
0Wu9mou8RXSD9u9Fh3HK5oOJf9+ugEkE/ijIv6nhZ7Vxrq7g8Nlaz+50WnZHjshuGoY4zWrQz2Ko
HiYBfBt2FHVnvh9JbneGHZljf0HrHNdyu0+17kLlMKomOS9NhLgF5kdQEu3zq2VdIGTqZA9cy5D7
DdBHhHa27pNbxHyu7kiBUf8GBloxtuSlHn2pWCsVXZC1aruMQuWPoLIGNSXsEXAXhUa+hnad33gH
Gw5IudyaYb4R17WgE0E1+xKZpml71Cm+DIJD8ng78kHRgmdhKWWepQNLfytw4SNI5SZRyOoFxuz+
ZZH1IvIBmAJcrhUbS4TdTgjbBMVpCmiO22do/g6G0EUueJK1KedltDuHbHULf4QnKpC07mAPqBHC
OogEW91krYkz7W4C9RsnpRCog2rFVPhLZH6zEHhWUyXt/dK90ru60fPJAuVTUlNbhRGCVg8PcuNy
/R7ZIdysCWxEGUFhpHd59lqWJ3Mjs01J8nDpInyXF6gR7CawwdWH1zN/7GJAnIbd2pAY6fmaVoZC
wEje0198wOvezoTYoK+SEgCxLw5D4C+no5aPcCTCJgNOUOi9e6ss2drTW+Uzy7xTAG/6jQFY7tpb
U4An5W+qzYp5N2a/8NeyTdwh8o3DSDs7Uy7EossVo3GN9zFgwt/JlT5LZYoPSDejhwUyQPBQLw2C
ltVf6zust9nZx27pl7Vnn7jOtvDVVSGuAygdTixqrUSb3qCQsUvReedRJqbH5FoBJfuIwC4OI9eG
BgsdTenqDG17stsvq4Rhwg9sj6IoKlKMqB2sIoXetGgsv7LYRdj5Bgzaxjq+50QFmngsqHIISoxC
BBSuVx7s/MGN3tyiUaRqsTnKPhRrMG2icFBsPGHXtfNXTANg5ocZSfg4PBCTukuq3KCEvboP9PzN
SIoEvRgSVDTgXpQCCfZsjg6KCPPmVzJZumVXN/C93CIqACAxFvM1dib0flhJCH0Vl9QN04vJJ/Sm
wm8lRfePDJhZ6WqvNQYdvs581WH+vVthY6CUCJEJYGOa/B354sIqEK9erlkCNtnaT1qtbBTrTu6e
b7amFW3Exe4jAVBz/XwfPxgBh7pK4YJDwp4y4QFPS2Hr7Q429T12uhfFunXEzZUOlLOhGVepGOe4
F2Z53X7+iqR81nJe0yqYA9SnTl1dIVZwJcz6N5otHuwvT0MD4d9y9vcpIAHIUwZz8XW4i3ALcZA5
YW10LasICA388crpFzXTfg9o1L7jl94ICCBwKg8PMPtaKMImUwFO0XJhmtJgiIXYzgH9DYy1naqg
/k1YpL2zsTykMaJg/TEP4qZFxR/BzhOl3qk58aB7iZnmtLviWD87cGhJRPIs3SMA6JoldubZSnP0
HSQ3qcxT+Th0NKvpQHSPGFBPvLMM2xYH7IiYr+on/pKMu3vnunevO8lFziyqML8r+FeBJb1jQY5+
m5CLM0Y45fDl+7RI/MrMDHQ6UBQis/cRnytk/XDEwBAz2vPF71h1prDqqxqILIF2MkkCXKqBcAyS
KFMF5fKRah3DcTVyuwF6XVXEKgwBt1uobJalHhjDdeF561c6YE2k8Z1mCWvlGi4GIjLNEydl3yvg
k5V6yllZajds0JIOLclR1b9+BDKkHM2Nvo94IDUO0ThzGjsO8wZT/4YDzKWVBhVBUVYtoA5fNama
AIZlmLCwJWnR/Vc5bDeCW/hU59rp21qFhL14rHDoOzCYby3KesC2FoPia2uKXV79JFYVjdjEDigd
Mq0Wu9yZoqGcVui29xZ/nKFmDQnw+ECNt9azPDK7tBXeL6AmBptLUiBI6GU2yUi6Lq7tuqGmu6t5
48lTFeLQltyEjrfOsBM1majuUdV2eq16bZJyX55GAiu8+HF1Uc9eN1sPv3TCcHY1rSbCw9O9SAn1
aHxDxmENfQ8y44rOFGCTE4alMnW2V89VYSUmHsM0JdBTx7p6aUe3DTLxgKvPu2Fjw0cGzqS30a0X
3MPTPUPvqGek/hwIl4j7BCW19QmB/Nu8mJOLxjpYxV5wWYE0/Lh3E92eAvbw1vALI3WMMPBqtDQU
D0B4B5XHzm5f6OD39qFsiQgGOGmp/ikKnl9nL9bQmkCPpx3nmASUd4DXl8PToZjRs4HdBzSuYW51
Vri+ds3SZ6i1afv99uIdubZNaMrOG3ispud6mz35Cedccd6EhmIsxnPfV+7LwdJJz6b/zWUyMNac
w66trfJaCvY2SS9PMhyf5k5ndgdPILUm3/0xZPcTAd0pnTle5xKAm77HLRNL3TlTMgP+HQmmcNoJ
nXKRFm6Bop4TSOF93JVypz3imNlwBcfKEwgErRjEPSJGIV98wEHTDjILhmOEndYSUo+m+tgVxca7
ykHEgNgrWzD7ZY3htucjjV2j2NEnMvrCSchXiDQpSnmHjEjfXR9SlD8NzWagF/B5SVQ+nvvEfqJ1
78us8CS/uhpzBfIvjtVf0AB5wyd6ylP2UkW1x6ss8fK8ZWgxgRaWf4cR5RUeBEDdtddg8VeXMH1/
EhyK/5r/JZ5xmWUyGON4SMOxOpO5od/16Q59Nt5nCEltOxLqCiNOWc37HYOYuM/aR06U/VChcLRr
6mcIIovCsup4osUaW79YNRohG+Sj9uXIjK3mX+E1EJ420+igNrkubAHntPHtlxmutfUU/K8JtL0F
ZgvKHf3GZuxgFLp7JaNkSpgn+Bp63CV58a8G6w4GngSliwNJAmS+715Xb6jXF7J4A7ThUXE+D6Ft
yb+LE/4uXIVMVV/oTO0Kb49NbiB4ufNymugQ9wSH2RpmJE6VRaE6ulSSho7JgXCv4OFqB8L49Rdz
3gz1XyirTsCesDYjFKzPvVnpSH6oC3eqtGG4pNjbghIu0k/PBERRGBBLAMjXwKnFCpZCsDcLtxsw
TyICUho+4f6mjQytRPMDTI6qfCBBgae6PixbMbM2dxVK3auNcvRdfGseTf0E8ZzDz5e9A1hXwOup
b0JHLqm9eSUaKT2DTSdaxPFzfwWxOAwg1ACnbrcc/Gy6JUzzxT5bbnNnpxINNTpLwkmuR2Q9kjYB
CRkncnyjwsWO/4eRzkoo9theukDxF6obs5ff07SnBA+T0dVCkt6/IG2nhoOPZNWYcHKB2ohfLLjA
RJg40cGLGbG7iVgC+G+zPpg4O4FpujZRi5wFP6hirJ/99wd7MOyZPfIN4SVI69yeuTuP722pjfxX
kOlC/bNUTL9BBGFvbrfbb9JIzQX+jSJUNtACxZ3UytQGhQK0tybG4PAyuqsjiHCeLaJ+Ju2Y90+g
hlYAqCsDnNChQUy/Cvj3KvALMBS3NzQr/+v/Xp1gR5woSIdLIA/MWMTm9b4Utr4MsskOyv8uI6eD
B8dGFSADOPs1pGboQB1wdtw1nEEFwVY7Yi9DKAkvvoE4vRrhXWt6pWqX4jKe2j/bRbHcGoaFMBzk
v9PhO2OnwRIg4QpPnTAB8O/n44+peKSU6i0isrNoqkIEEuUxrYls9MPDKrYntrAiaGqrv3KfDGMi
LgvGyU883KRwhNMnweKJag2x+d9H5Fv4fN/GNxpKPvFvi1PthcOnBi7WtleymYveVhtwFutg8O7j
e8eBDA/zwBHrZ1QAfKgrK/OuCSJ7glXIwYkHk28V+la+6Owo1Dx+/YrekSo7VGP2mlZ/vNN3YYcm
xz6wZL4uTXifHAfYMkdAZkiSW/0CthsgyencCbSYQILKH3740ClM1IxGJCa24SMJgo81Cr25jBbD
1AKbARhZ4jriCGLhdlVz2tG0zZByHf8V4OZeJ8KOja7AtsHSFP2B4jwVKHBYhF89UFQZYnwAd2Yt
upBv+qZPZAT1CkHJXRQdKphH2anQ/79jn9hoFIubVT6ZMFSvCzqhvsT4V6yfhzBQp3BkYdASbOJl
YBtRDT4KE2aLAamjngJ9Y7sjLyme0PcFU9LKu5qaRh+sEb36d5EB/OfRNYFCUcyhtnRMv6Wlc0nr
+T4Ev+xjggh2MevNu6uVu/MBNHWM7M2gSgzvdQvxphNyqzR3sQxi/KE5oFZeZ/iDnA8ERw7BbGus
0HLfZO4tkHKW0Mx7ysLxMV23almv0fi9GBmsNx2ud408c7KGn2O2j0vrNkiqdzWkzkInUjTEGClk
CxfgIeXDiPQ8TIkuyG3R/MPsRFoxeiNl3F6vHSlcPiJ6/qaLXvfAbeLR1GFBY5oRKjrwOmuyqUsp
XCHtRONGxwpkeK3+CFBudzlUmJczeq5aVjCfUkeh2cIwT8x3VGSvgvyB9vaASIbPXQLtURAlkixp
nV54xoA/UfhXF99KS4NsSKRmwnqdJKGz1iyiUmSPIKGc/vRz/7HMfIMIJ41/4L1c4+CMrgUmERYx
bzdKDE06f2THoHsFhh4r1cs7s4mfDAqTOUFAbDwRPXlLaWLuW9YLRPG49388fQ55ExmJ6BZ8obt5
3rvBVFbMB4Vbcjyr9R69I7BweEDCs0S3gCdKKb9r/MeodWtK5vo/1e7RpdPvlMldxmh63lyx7YVS
mNXOMSC4GEzdXYeB9CQEOAY8sK/s4+fc4LzFYh2FjfdUVvba+jwHfYfjQAxGe+7d+InQntUgBu3G
frZ2YJ++voZ7d6xdb73yE/GkMq7Q08jTEDERZAuFD+kql/DG1YxIBvQAuFOvPZ0eBLSYvdj8pTHr
IKSTKWVSq8HaCixbf6jTjcvdTmIpxvqDTyWq3JHXF2g5ACmDSdPMfDozPIAQkTxj9UKeLG6Tv5gR
Jg7lZhR9YVDi/XkdzK1m8L8P+FX1TY8AT5SYoWlezCOgOwOskv9oW2OlldEEOrRVdA9VyEsFFef8
G/GKTGzW63KQLqWzVSYEZBVvWYqS5cPWR56ZBWTrA1eRRPWSQ64m1CC6ySgAbJsfa6xQMC53IQDY
Zdi+wRsa9S765NpnSMexeLv6Cd7cLeaQ5skhQhESHv7YOPrqS3cZ/R4pS9iRTr+BF/08ozIVq+E7
Ntq3InYkLnR1ToRsT+kHrbhMsT6EQ6EuQEOluPXRqGZaR9s2XeB0MgBX6YqyGz3RGtqHZQ3c5mm4
hB+bpZx8qmUyVYtw1njk4xg8oDKUHvBe+TCgA7KpMlmt5076wPaD5iYxX5Y8qP4Q1Y7zA5Zr2TLW
/R8wZ+Acha8VgFVKGips3nEqSk2xFz2hwmwUmC8aoGHFT5b16W+O15RXTyRhcGxAhSzaZMstsB0W
n/I+YNVVxqCZGwqtA4UoYHAeCwhelsHLcLPrEoy5tKrtqTvtMUpMSLF5tdh6/noGpXWSu6ejse6L
UQ9y0niCpNcDO2DAq0xF0Z6P8sdzoIiytqiPPaxUf/h9XckfdKkVAQ9uqO87W+lQ3Dn/N/9sMeJP
dkVLT61YnDolrFdqXiVkISeb5BM3B7VRj5Cr7VR0FZYqux5KchJom5ckz82tPd8a/hjUD0lVH52r
pdIc0RSG75fjIbLpI/K+3kEeEmlzFy0BG1jmozisUk/5pCLn42J95ZLzvBrGz1MurCTQSHgslF6z
IKHj0jUg+EHvSbbAaDA0X+MLNnRGTzxuQVPviRmuDWm5it9ffrQzLtBLH5RvN79d3VJUnnvmNzUu
TzEoAVNLgQHPYYx8XbljnGNbu09oRljAlQG0LKD89XsqAVfsV1K4u10zQcIJMkBi46sOah+dq/Mv
WOHR+YVvDu636Sa+R8rPrWwzyQvlDm21KsSiILdhwSmjWgPl87aekTA3hoMqfalcjb06CCWxJYZI
IPj0/CVnMTgNVibZmmoxXKL0bYADAdwY6p1tx8pHs9eEOyS1KJDMJPDJ3+O+s+SEiMjiNryDyy4Z
Owba5sUPZ4kpW3HtSpt9XpNIe7mOcyOdBli+Y3/QeysUGmS23xQklZNdEkfxbOe6gocE+1rNQkcM
zAwiy873teDVu3INUpukvkpLmQVbkOFBh7FzDVRDpCOGWchTgGt+5lelGl/ZLHDM8WHxslFY0WhP
ra4vPE+6Ey82eTGU0W14ysY8KO31+A9SEcPb93TzIWpxQH3+7cntXRfQBzuDFrTWLI0YJkmiS29R
GuKBTSFBIZdVeUg1pKb9WWhsfzxoPSaou+4zs6gaC9JlO3CGyOCxF2ATOt+UhGCz+Z36dgeP1Ugq
j9QsYTWfalULadM7qZ5aFZenYLxY6fFHo8Wso2uoDKA8myDEpnHhAmHIgONH2x/0yt7fX33IoiFY
FtOq0nA4F8NAhC2pffTSA7C/QM1CcDhDnKpPImJntBCEogh00GmJQMdZX1kCNZpsbWoPipWgfxek
Y7FK3ISjFLKsbCQzGc1V5625c61L/dVUs+CrMdj6Wwy1OQ++HAFMnFTaOPpnHnXoXuQInKSh0df0
h5l9bBnAoAnZH44tx3hPNWD12KBF6G60LtZBEpsKOKz+MqadhR5YIWYHoXn5wh00ctl/FCMwScpQ
HG9B0zglOoTOQ4zXvKZE9MaI8xrczcUG5mRZ/rn7afXqH+8VPkB8zAI64XYbV37Iw4fbtBLdmNlE
dExJ+0ziNbigCbnh/g5xgdZ9jcAdcUdpXkGDASdcTid9+EKJAYd1HndPDd6rZ70WGvGuDD97jsUm
Imh0rcNY5DRT0cBVvAWNX44NJFpMJG9YGGpuNU1vcu32UD/fCcc4Y8atb2+jhz4jm/Tv0i4hpfMX
b1pNaBszs4pyNNccIJoVX3fQxg0HXHI4SoIuYTv6dXI/TQ9nv2XTfkYqZJ9uj8Fxr4WgMDxkoKRb
sUXKtpAWQE1Tuv9PrhlWfOyEIu2mU20KE9DBeDKWXxFq/jU1jm0eN30oIbbS4s6rI7gGDWotox/V
ll0T19Mer5dO3MI5VxDrCzYW3fqG21CSptUDve11amVx1aZNXAKAemRIGaQ9s11QiEPaqf7OOtQV
3oPYwSufBD3S+gBOVSlWlW1kItYBjUBMjiuPTXb2EInjl4LSaJ09fjm/3pr6/g0+BkBs9znIQajq
y3MxnUCojBIrjbDJWo1rct4d1lHidGz+UpKMcWAU9ZRkgz3WeMfJv+NvUc3eajfAjo2EpZNsx6/w
TsWP9MD1RR9Sb0j83B9BH7joxPjTEAZMwMFJ7JyVudQRrbhee+G5vSlpxgHQ/0lMST08uklShCrP
ME0jWtsm+TuEvCSe0vXHlDrdkzqbsIWq1u6OKeOaUPWvU3wbl00TgBfaYmepKQ3JpisxzEH2QM7r
nLNIkCIpyrbU9N5JFlc+o3HbYhV2gv8/hVJaVX2DXTJciHwb4jh2V2bRf6aTG3zf7/rtrFjgBZhB
w8pyfyfthzdPbj9YgtBSq7lx+nGZ2ThsJDgP7+yXcJSKNvmU8YLIOc9EutZzhtNj+xadcGtl08ap
7yDKpcmUUKphGDZf9CRla1/9rTyXzk0MrCZkoC4PO7dE06O7y9JbvMU5N/3y6fNvBUG1kUkLztrT
q8AdqeKIK307791AYmPzz/3Zrkj9V2/AI7NSE6QJu8Hyipn2MGSk8tTT5QWkEn8PLzoEbuvMeKY3
Q301rCn/yQEM/bH+QY7NRWYTnVT+47/L2aty2CClS5HAfqthH7A9eyDAFckpPxPwW1SPwUwlEDoi
vC4fq9Ha6QjLe3+tbNMc5oJL6HlqhfNUcBNvjo3oTYnFoqPz3b8ysPV4UqNcPBfqgxNjPGJLMpBi
rPrWz0LNgLvUpVyu0cZWHYOtUT66O05yna0tnro7lN4xugtGyp3oFQmrEOuIecesC+HkM0zzRGss
qx27U3UdtvKVmj6cGyREo9Shu9GBVpcbNpD9fgnedZ+Nb/jCfCyGb+LF3H/BFdCqrZU6i69Mbny0
mN8n0KyCErER/WWijtRG7KdSyKgCUrgYjou2dq0QLbrEIGUbDotIWV8qH4GrXZEWv28nl1LVL2+Q
wrddjCe9XRUHYYNL33rrr0xCEnlgWqsgkyIyrG3geyCy2nZVGIG/Gja+PUSv01qcnhBrvK3LJoPV
vzkHNC+sRPhdYPZW1QwQtwiueZM+1lv09+hhUAAEbJwi9bGVX2aNGuiByenjjQ0j+2npRCTv5iMw
y0q9Fpkf/Xhdvwf+lDzsdJEDZbcMgvHOcHyGjgInfmNCiNcBIYqyq31iJI/PI8xxY8w6Q2tlMDSn
4Vr1V2BGuGL2d6EtzK0kit61n5yihoeEo2TXWgGeA64mCb/kACUoJjJHaRnaZ49/VnVNGdii74wL
Vwqh/wqrLmSIZBFFzvMPPglOb6EqykszpNAA4ALOeNAWc28/hUz32jOY2anfrwFJGdunZmSC6rM8
D3C5SBXIwagYnP6GJ4oSrjCHXS7W1geQISWF3VTmJzVEmgwkYCEhMLO5aOG9cI0y0Q+Dm3He0RhJ
obBOOTH0abvMLS/fuUXeKJUqbTPI0UocuaIxIHi0s1L61a19zweCKCeN+v1iN/UcjDcq6p3Qm4NF
sitQhrGx7e+SlIxbzuUs4F18DKz9BfRsws2eueM1294EF77HOHENllRJWB8RN3itc/Z+0qdLWq2J
i57yB45Wwd1qzTzdAKMpx8fS2zhEepfW8oYzn70LHTMhna5ihMsBUIkmrFwAL0TGDSu6RpSTDrvN
KXjhIvRC34FztTxkm5AaCQDva5NEFhYVoyXYGV70V3ngaU4KojqHua+otexLlQcnT0THnnMlJ9l/
i8LC2Am2KkPkABK8FEEiJUosDjmEebF0W+q1ZB+b9Q/DwhwU30hABS5EXOx7YOKlA7AdrEFYDCWe
z3W2pGYXYAxRwvszPQWviCAlTThU4wHbmVo+AWPDFbqgzHfzcMBPC5tesAixvcsTYoPP5V5Hf+ar
QF7c5V0Gu8gSM1C7sFqbgTvPqXGdVk2Dt+HVLKtxQ9kxAuDYlhEtrCkzgLJEdkljUMA9mou4xmDc
I5wcy3dBpI8jqAEXWo5befkDvPyavhEJNwl8iZPTWNp1+lxK/K+eVsXa0v3PmLm3Dv5Lcn6VJC6/
QKhKDe+kmSlk01sRITegQmBz/bG0Yadpn6sIg7rxOy2T9bzu0SsxNQWC4WbCKp6QLTrkKvtYMiXo
YOsbbl0CDv0OceZH5/j4z/5i1EUr/5kVGwM/9lDiH7sqoM/WtVH7+VxPlTJ9KWro/BSpAbUoGfUC
XWreOU/cExEormJhuuyvOlOj3FnQL9o+FJo53/anvhLrxLBnV+Rc7snyuFWHXtmDt0/iUkn+VfeI
RH5ClVLFg9n8pbaUUSpnSElwdQ/nSGFtHJ8KIicniz6VB2E+yw0vXscXmb51mrco3j6QAmlQFQXw
MdckynYgFHZ6WagklFoEjOZrgdtGMfh86JZ07njegUEpe0UY7U8ZgdmjBTsnDt5cSYrAjnPSWOOG
NYFADj2gERxxcZcgNFYFAqTkE2NLKnzf+eW4eFALEKKmakeoynA/IT7yOSv40sDB1M295FNvi9Wt
nZmNUVOn5MvVBuQTpDo8i0OXvzJrWi/SU55uDuol9ATjS2a5SwFKSeoszs5HUReOsDXtrvPmRzEp
8miiFO0/bNYn7Ch7//tN9+Na5XN+5h+dNaA/8OGeXbAD8WV+6qTpN140DGg5aCLw3CD0l6h2wiT7
66bPH3CKNzpdgAKLK/NWclaRbYA1+qps5AaD9BnzbYSBrp3tg4EkNQexOUm+cfXBPi/Jn//b+oRx
S5J7T9WRUnizhfbQ1UYG9ni2jOlHKQS9koWWO72Y4T/x5M4JVAgbvjhlwp0C1oAE9uLcUGYeR7x7
BIp77YKYCmQLNxEAJ7EDqymGm5cvZrwGF2kFAUYG7QT0i0CxKEqXXdOuHRYZ/WfXT9h4O+FMbVPj
6bDyY0Bals22DOXiYpm1Qnbhf6QAN6ThWFHJzogmq9YFXeKTJmBb+SE+uOSfIptxZBo3En/a2K3S
cFqwglbGP9AkbSucMkAeMUwr5RVQvsGwqM9+fSiHZ/DZmQVRL6aj2O2Lo00+pJEm8l3dCxIHojEI
VpnsY8dp5A1HSA9n06VO/BHG94I8JzTxwNJcdyZ4smXNq5dmM1bKspkRLnvPtW9D/WPEHGAjFNqk
GFg+K8foBWBp+jIgRndei2j+HP+ORmerHwl51Q/EjzYYHEzWp3vdLazrGYUmd3kazHY1eObeDeEp
QI5XdHeCKedx5n/Cd2gkp9cWwBnBk+TjCsurE53Z24cu84r/5eAJ3ztkc/OFA1YmxPyfi7DaN8NJ
Y7dKTYz5vHXHNXZLOvTAIp5F+6U/571w3K2E9KfigESptpLvsAk735rI4yewrrQas50yoFHWCq1+
0h+wVwJNQEnl2+ly2NOveH6yWZ86Y/giFUnkhResCmQlWIOuZsHZ7zOT2KciZE1LVlRRJX7oob0v
v4b967DQwVmLAkBelXs4zBXb5ADSBeYUoVUBkMZSk+kZfMWCyMifG5e3MH++AlfZkFsguSeGwr9M
gfEifTN+o1eL43pXHd8sE3zN8QlrNR3JcOxlRKfizS9AM1jLTSfKUz/W9dU+W+1RebqyQFEJ6VjY
F52bB/8HxNT4ezWsd3608L8R6It9kGGi+/5aJwb4CAgKLC8J0znPqlZuD47txNRkNUR2xAtZX9Kb
joHcw9DfhRj4Nv3I2AZuhKrp8UPSJLe4pWXFl9WlNEBxvrKda5ypmsXBVhJVu6hJb+/IGTUT2qkH
SqRh+q+1+njz0g22o62X5hydFWNaMsDQLX05VtqAj9gGofzhaYIMwAqyNHjTb784pr7HhHtmWAXb
fkqUSrsCGxWG+lYgo/0C9xrYgBQLBvMryvvHBWqA8SCyKYnHy2jfOFwzD90mT8nIywzb+IbfdqsU
E0fzkS786aslnb3RSNXx/mZAq9ieJm3ykPwGgUPhtDd5+rB3BUqFKm/N/mmNfKp/dQH53ugTYcd6
dtRmNAUTmLlg8ZUO7Sp8SDuiFNX9mVchH729pUmqAHaJKCiPsFfGN6jpGj0ivylmKMZnQcg2pRpl
gHiOGSFenYGYYdJdqh7jMpKyAL7AULHmQguyMg6w2cVM/O1Zd7kFHL+OyKX8IKKLn93aRVm+1Iuo
9pkH9nQpbp1x4grjqyo86hfkOi3eRhHVP2mxOIaVes34P8ZuziKG1fEXilFvSpN9CHr/3sQI/9PA
qeIfFoNJ/9lMZyviMHT9wCy9QIhbDKczRZUTbL7UCBHFNeRcl3ShnmZN0/L0LL9ETHMLNjrFcHIh
8iygQiolZNbRT5Iov6bHp5LXgdOYVIcat81UD8+MlzhWBqZksITx4SotCaDYZ68mDXhAcPl6Ktz0
/R8k2/II6xYzramG7OP4k1rjVJoSBL42Qr/SihkMGtVuX3fy5UeqbbfYQdp5q8ly6aEypfyOrsAN
JnTfuW1DkyM8URKkVJaw3+ABsPPFUD/5C76F/6LlNVv8l7pCqTIMVeV7+q0XjkyUavbllo+l/Uer
pRKmqzY0S5y575feVg8CXTaS5snu/mKKK1zWBiPNKlVyZbz4C9VDnmUbrucNoGOFz2+3WbKA6fxb
kqxzqXL3BykHrGvfyvhWo9FYvDTkx7FGEgkhVbJm/wCC1we4WdtEQxGbKwn92/j18+KS0H5I9ImT
GxriQMqlBzbq8mtkey3M9AtuMsyNWMQJzktTfVzO0FtoQ2Qi28F/0e16sof1yipC51/YzLCUx0tp
XPmV9eRof1rJ9TMCNg/7HatSGk/99TeHn7cvyR3Cy8npOEvfLUzKqCkCn611x4g4j/u2pgb2VEV8
/pKr99DeTAKwPucLJ2J8Op/gDbZqY9LSn2Q8pHE39QPmM86ld8BUWCgoVPEl7Gu1dE5iRgFIHdfY
CIxCSGGTQ3xiq+5TbkmF8OhOGWDA/d+S0lTEVuMI0EyzamV3lHs+9DXf2+19JFGISV1FIOEY3u9f
ssc+v80o6ra9DBIXMSTH6mQZNW+JvSMUNcj1q0ZbY7QW0HtquLMSGtf67pPar7O1Pemf+lVs3pht
101iJjGcPdBeuELPYhEq3nRP1wBHmpyqhs7gfRUs6nlXghZK2+1oOzSaUEMn1GmTFXcgC148OESE
EGss1yzCjvIgQ3Mbs0IrjpPfXZMRw7zUute6nuT6ZnVvgnNHZWxemq97KfFnabj7uR3jLtA0s/BC
5wPr8TzX7/ZoG5XoXiJR79FVT/ar+VkECKpRocnLOsKm9X1nuvdWt2KqUzIl6Z2q1BQSF5ziJxDF
1bpOYdslVsT8Hv3v5I6Isv/p+XFAf8eRsUbVzjgiANP+m6Uv2B5Pu8VIbiS5ivpIaGnbGZc5GIUa
fWgvGDdtWliZXrJhyetHduao56mmwmfC7Lb05reeezVNIMLk3xTK6hyHZ1h4LqVKX/Ddht+66SQG
FshDPLibaT7jxOwpT5rpakdNZiYMJqU+my8CFArRvsB+2aW6+zup2Fr2qpSQPQwVb+aQwm8OiueO
PPDL5MfR+saz/WQyHcwZoZfHw9fCXpyfWmkhJ0jee6MnWFCUdP++zfTucB0IgHVq0nKdKOfe3zLw
1qhueM4b2YxKl25jkIuu2EpPDSHVZUlmsfkyCvsg03cFm2VbsXGc31+3cMA3JWWMsYZw/QA5Wu5p
CfzS2GvenIcZLCEsuUSwuyw0jNCtH469pp7LTznEbfI3u5y0NOAMLnTWmOYb3KLBosTYVs/uWWBl
azklAGL0YZdXdFXCHMVE8cSa/fJYaBMFEU/1p9hQ9mL+1fLaEzKQ/R0p3QXg+F7rfkTyvPUnsXL2
/0ICuYqZMGVHaxlpAc5UIZ5dx2D2Qxafr0YbCwjmoxL2ubojGFKnfs2EOn4unQXFQhsm6TH2vPu8
aPttyeTLH3llpSTgSvP9I553h/PpmMqFVWzbuUSihwZL/2qafIT2aiJ/MUj3tbiO2XTapGyB1o/d
YnrXbCK6yADQAsH75dbDE5o/s6qC9z6kTUcZBAwb61bP22z0tZFouiHN/IvHA0xAvXEA94fIfH/G
biSUc8vkGKTOy00VRA4xnLggUNpNQmZcZGcvnGGcZ5SS7G+J1/UYrlv7viPdF6h9sTwluVq1OAuu
k3PsJ8c8nHRXttWQes8m+YrS+32Dl7U//Kv+EP7tUbT8MfXUVEuozMmOe0hCrGb2ZmJzt1IL5z63
1Aw1OeVLGbKJisaaD5/B8wUskjoB6RBHNU2LZxoe621h++WSeGpxSiXXYqIjU75X6YQVurkGO47C
tk1MJlRC3aeV7WRb4lPNGiFSf1e7CBoROdgiQBhk0x6NxH9mjOMx2wNw8m8g26QiOOuFEVLS4Z+w
INzfqCO0iECRTQ1mszv2hP7O6GakYu8ze779ncaRsYFHZVyWz3SHcjlTkNVhqennKOMIT1NeDuY4
jFwmBPnfAjPebQQOszSx5ejf65ju9U2C70fGsp9im4rn8pN8gjVhO2bTWq0Jg+KQ/+T1oDlb6AmP
vfJY7Qik7kMNMjkN/bM9MDGCMoxnZTQKPOGL6o1rkCOtun+Z5X1rKPJS/hEMkjtz49Z3ys5wT6yD
Pr+33/C2Q8uSOYrcKZOfES/hYVkPXdfImUBsWAbCUzgI1Yw11hTj6y2CbwmRq8TIYMPweHrrPZAz
PFc/XuXufQV5QK01oqhvjykwgpsMgb7uA58H1korSn0wmyaEvm4Aar2Uyp2hpli3rmc5CiS/hBN+
hLxis8UCp2dFYkp9EcrNaGOefR44nO2lvlBBaPCDUVqxcRmdaiGTH2T6MUPQeek8Zb+47/5tz0p9
mJ1I0DB7GPogf97lrOh98dSvzAWTPmQ04jCscriL4h+KrzzLjHJb+1JVzq/jVlDGyo7A8N7AqSR0
do5B+bJxFHNmwkL+aFBrNqLT5H6VTM8XrHP21dU+XWSrsD0eClCv+To7AE2FdxN0o+0Fz8McITbg
S0WOy2APUGbpvIT2fYnGI30amp1LjfrEndIGj7kWrQhloSC/j3ktynB9vasEdX5hklSX0aXvI1YQ
gSRHdTWhTZOTNzKG2XNxP3q1X0TjSAZMx+HErQQ6sLNyugd5mkknjdv3alHL4qmU2PoF5s+AKUn8
ILSVVqgfJ2TpfBmFNEcBn4ExLmO4BNtl0aGnoBexpQ1VhRhMQvDRljktskhX3Uy1fW0AWt3y3xYN
rviGtFNK8aX6reCgCYdq3F70uI15En68N/QEzZYASi90mlsUoF2zX2rdB3jJK/l7DJiB0/8pbQUA
OFCXDUtzZfiT4YoscfjsqzqPwC9evhTZNs0ZGDtb2l6qCksqCgUmaCmBDflD+FsdBwK/mp2pSX+e
JLmJ2P60AUfIQsv7PmACNVY4VM99UPnNwosxzNjg4wToFgUo+Oww9vAZMPpi5BIky0FQvStv6tm2
a+aoelO2DHt/1GlVITC5bDisq8HvdoF41TTD5Zbl9QThLM1wSneFxuYWd30C3C+s1Ol2t9vD1+KD
yEmmoaIX4BYGWlnmCwjDhBbfsCJp3xGingnCj3Cxr8vYy2PaHCAL9faUkxojPmq1adCrJkUm9nAR
++kFD7xCiwkXgXRZdXZDXahkmj0n+o/d295pazAT1B4wISkdBw8h5r5qUP0AcaCY02hg8djDkKQ+
4FQNSqW0W5qHvzfesg+T35qBP7OhMA9EvYofOmjoRpRCmgrqDyE6KqNOoTKIMtZQnz+5yYkw6OBK
4Kj6NnFI7FMTtp5kpYThTXWEnlPLXOOQEGAk1aS0HjbBpEcyF0u725bJX/utt/D7AawQHi/6S8Oh
DWkoBtAJuuwJizvtAD1BehkEae3XIg1oQWseB6DOM6enXEkF40jMMLnQyz9frkXQsTQehlokb3rF
8Q2repFEtEuXd+wH2bWpkoS6WZdzNdNXM+wwiUIgwBgD03+W0q1CwjOkiApuilUo0nNbG1eoqTSz
34iuonchVV8rpeaT0B23nN5qmugRB0HsIZj4S/HHsps7boBzjACJpwJIyk8IAvGdKtSr9h/nvAm7
5nQz1PEN7ZOuLjZ39LoWQPimZl1WcJ/Mv46wWVgYMT6Qw/M6EGT+KGkzM3e0d3/iRCf3LgOKgMSb
nNOo0YRFn7OpdTZNngfq+LbSus1o4PD/Ws9ZN2jNIrPIM/9ccJkI7O7rEKQByOjyDfL/pwKnXoM+
4qnRCkzcBPMhdy613/AxxH/TYwB5ns4d9QNBHZsJe1n0i/hwxDkqq1zfzF1l7FVpFjIll2eJqbjj
yCn4CiudfGjVJBYWtuvnPu/OHR/RPXgUNF2La9Ara6Eo62EXG207OpRbUgrudBCUFn6Ph6lAflih
IeqzbPrhlZKRU3rMLf83UcnDCEsdLWk2xntqLb3c9ke04wGPE1r/Aq73yQPGFciWnPmWPgiSV3lX
Zf0PlbTCroGNhFeyM3V3MnFrI7jNBVh1b+KVHBZP5iEcE3inBN6Rm3vx6JHl82/9W0Q9/RpmOCDz
LtoBwWLdb3EV03Q1yGC+AzKyRw6ryfhXIk2OGEC1fkt86rna0e1LEpievoT0Bb+TSgwTdaJahYP3
bnNuHS1yBXwAL9DSfvtduJnJcJu9CBLd4OWaDFfj+HtIUUg0Lpg1zis7XuRLf6jkvHhou+pMzCZ9
mkhLpFhHuOt5RORGaGzsm7VVaBzgu2Gupv+7kFpoT6k1RC6YssutbI7uxPRdiEDWGhQfPsrmla1u
MXVniwS3XXRyQvdVHCCA4rw0dc6ztWZrQAwhLO7Yf/qC7wQNIjVuzk1MIR3j5mjyRJ0qZvo1T3at
AX6wFTrc2SdgF7P1jK7KDgseXaaQlfIPC9cYbQEjTV2qPBPo6tKdkhVMmsHOK/rZFQ4/kMicdefT
LrQLmoExf360KbWVGQaIafJ4IQqX27WbxFLssEDulX2t+//2dUpP2JkTposF3u/wagHp/Q3l8qVp
2oNgcasFb9g1chh9rD3A0FF3E5+Htci2RIOSyKyA/wfefP4ECR4vu/cWpEANf7pYve/+t91eoK6t
rxs7eU3EBE7SjGG2Ag86nBUE/k/wjVK2IamG490VHTst91qSmqGsZLVdXOuJgzmXjDlYW/Wx/oaf
wYA7OaKHD67jMhMouvkrL66UrK4tZOMl9iMM5bEXghZ/6pwxiqBg9m0umRc3KJFJKXjL62fj1eFx
O4IXGjn5mDS4uhU0M+FcbfLCP2WjXODEiCjG9SxQ796Qi6rOkkspzMe7smvhYy6FiIQ61ApBGi7h
+knTapd3NsqQqmfrK9xztI+fv3wSDXQy0OXD9X3qXSyiVQDVkPmo82UsAFCnLNURghOkS+CiMHKb
J1zjfPCjhlSC4GB8oP9iT6OGad+Dyjz33aHwkdykvDeNyxaTGynureJcIjpTiu+kMG3r7v573+WS
V0l3NThxVgr0h50vRJmLxr5IjE8ILY5AZ2zQHo+XQdYw2uNW3FOtMgYXOocq4eKJ0XleLBYb3QSl
PsjMjNvs+UAJA1oNR8xzL9uBfLbSTOvlCfG2gFHHNrYx3/+5ew6g0IPyY/yqHid7TLnGyJJfX5+x
8hTFA0EZ1qPRsaYbGLA5ghbJvFa6Gt1WDAdwLHNIa+SizlkCjepvjn1goq9qwcYdJGbGxDJs0RcB
dfaFpBP15qecZxkrShcuKGOFufeadAiPw+DPQ47k436moWuZtqj2lPat1IPaVSHsIH/yxlef1wlo
1ogo6ZRhMQfgcmn4KphGMpkk1XLWl4OrZ5uQz097L2qpKxylSoCi8VBt3823XNOw+VcTE2AK6N3E
qmGoYGVD71QG4tq48kWfPFKV5hdVOVBqQ7HVUQmn7rGt7f0Z53h3IdTGlnHkYyTdvN5NXm/35m+E
vJ2fV8vJ6IKJcrLE2tBZ1F05rtq6rvthDx6CoBxBHLA+a/UajusAed24MIMOrS2Z4TesHA/+re2D
WyOG3wuvf6xbY0nThmLkshI+/ahVSpZO84H3cqZgcmcEUVoLPT6IQDt3lGTAbNsnq+6Dpe3pHPNO
uHMDJaRtBzqKBEYia/3iwS9VzxDkGUK5qEkhGbdTI6cNpphs3gsF+liNdiBSBBSRrfhM138Afh7t
XrJdG50Q7LjdQy62kvtbp3IO1Xg0OgeflgaECPluLcslQ31LSj4qrloRZpfhVvXzOVj8F9NseyPq
mos+rlYooGq3u5zAcdWfvSQzo0THjJCpX6NP6sLxrMEHKATOvtzSJ4IUrhEr0qUBh2zv7bwfdOzJ
zm1Qw0EK4NjKrBeJOpTS9iWJtjYK39qQ7S9mfyPqXKRC7YZH0IopSqGpEvgymUg3KZEeLRkbnbsS
E2CVSbiK6OcbeBiS7IutXLJtzD5/9gCpe3aTv44PKkZyJcHUy8XTfpJ6VFy/u6+sdp8hbizoN4wd
mR1ZfD3P54UTInlQ9y2lMJqRahXS/kmAqSmZMoeg7FRNJE8y9iR8Q6F+kZJT6xKqyPpFqzfZ6oe6
spQgFlGtR2QGe3TEY4q2AX8XYBpaQooRKuaiRRyL9yH9ZL0C54GjV3cQ0+eQL5dgjEDhqZBCvJHl
buGybfxHUOb9UXS28br0sh3LSJxti6c8DK7LQkezIB1MtJLTsv2GeIZWFsRRxVmuaLhq6Dd/ej4r
RbnKzJEmV5KtT7s+3dQznfhE4BltcSCnG/zJ448LUuLSg4znH8bZexX6UxxKbzEh/8t/fCDhSP0R
AOrHG7+cQvRE1hIJuil8inlr4irp3FFb48qsFMctn1mkd7+BeWWXm4JcbaMauhNN9S6fbz7WINjX
2HjReXr45wD6tq53c/X9wo8A7dp+2XDMoweAa/U8V8vN69ZiIGnziuWQTTxe3KVBAgpA9qX539U5
uyQosPZaEUrGx0NtQ2m56vXZ1M3spEzRN6ExrhzI2QmFrSvVRWdO6XWPJV/OxT1cjjtChkC3xCQK
2jiaFQH8vovbm9JhhZ4oR1szhAbWExAANR2XjCkiMSp7V4VZUROsLxxsKKYzf9YCTKOtB/wHPdwt
gGnf57CeKPm7uRJ8pJuncbQl6XkQfl8d64oqpvmRSk5Zq3D4NjenRHXK+98uK+NP8zjQFGz3IRtQ
YLoXSztB3Tzw+RTSjVsfi0wjBgiahLudmehkUKfzZKY1K2E3wjzv/aColeP9sspaADxzg46d9ILT
YAslIv4RGgUKjwQtNFfq+MH03urIl7iLp7ILGMIUpHTp0O5kfFSb2fPEJlhTzTEz5e2XBPxPOc60
oDs70wE9zKwyPXenxvtQVxEdZifr2qgWGZCDpv60fNcdoIkjnO4XbiFaLqREczUC1d51RWsmbbkU
pvzLwHxjBIuTGb5NRXV9bqjhgpdDLRHTCDbm5boGJ2shTYBV6TzFk1AaHUq9KHHs45DMuH3oe2yE
ijiyHV1Xta3WrfW26M/xxiiB08iumBE1E7scXnDTDvaffimcjoeXURDIrJLoZTvBsBAiEytLgwRR
zq9bqPD65mu7mNg/xCVExGeOx80ua3LZiFs5adGfsbjvQJ7xp90nUD5/ANrWezLof4s8PRFBDtzI
t14fSaoBShdOtz1Qt03hJdztD5mmTP4Sm9Qw6wEH+XJJUmAYdSx+CxPJeyMYgBIeaun+HUGk2P5E
aG7v7N6ojn9pjfDQhNviAlf/PVcMRkBKXJQmfW2sh2qsjabIBs+JneSRMdfM9aq2AxJeX5cJwshH
RLWLWgi4dclgja4pGTzgDUZWjNhCii9zydykX637rJKvwpn+foWplB6SNHXMnToASBnUHr1va04y
LKDvE15b8rOdH6lcELQfh/m2PYBWtO3YbW+OeSMtuYBSwTwoc7LRltlz6WPf9k1dq6W2P4Q91snN
zJaixCc6+xYi5ximtLsv9PqT1FX4YF6FbGXQOeTwpy+j7MFLcqgSE2+do7do8iQ+3YNMQHmRrQeZ
ldwscBNv46Gle4TNrkaYGQ47Fr4gmj1r6J2TycPiJ+SCdCfiCbrUmVl3N36LLKr7lgc3jeIqOFGA
h8RpOuykBaypfwTpw8cVE/OmMELIcyv1YAmMUe0wLNDCVukvYcZaPPUcZ+II9DoQ+JcOv64h5fng
41ZUj8TM3STJ7XMAWeZ0Lnwb45aDfOTBIxeg9ewnoe9rfv7zhsuUQIdZZoRNGutfYtt/q540fdKO
m4oz3n2JAwDq8iwL4NyXelJL34lhw1IRUkYw562C/JzYKnHMUrUUXXCLoShN7kq0APhHthBCfKzJ
LYSJm4T5wzCK/0E3ITdOAQWBk9CiXUr1HrOUj5/28/boUlm4EoAokTFLDJmYeqHF5rKi8xCQZkKH
EiRwMmltaxoY/c7cCsfT7hDASpLtsn2JvYTyejYKEIJYO277oHWVDEDmN/BOHoM17df7mrYDZ3Dp
HXcp9+qJNXMnIg8emeGoNSafHy6Ca3XHAv8WpCtTCdYkjmVR5GJDznnQuRfjhj+RELoCK+PWbgTa
18f3SFfWTR7SPpPY95btf6cYpiFeLX2eldKHYGY4gWEPhunGc/m4PPmGSHjNB662/LGl3t7VO6T7
1dt32nLO5Woe9jZNIFKUL8Z680do3Em5E4Ks6b4dybhgg/LZRr3cw+GxwsTYlsgKq42tbn/DDeSC
tfzpcCDTCm15DJ9vl2P/yxZUUdMNCIGmiWmKhvRgp9JsGx2NuJ4mH9n1hmqN2HzgxXnWysuKtuHI
68NScZdd4KbCcoE2P5i+Okp6Ltpe1rxnFlf9WRkW6kXPToet9xg2PjLqUj7wAJxkkAEnDa8m1ARu
dEvSnvWu5zA4ilKAZx0V+9YoTIgaea5xKf/jMXj0EKKvC1eLkaaMzhrU3f2T4hiMzj6K6sEmo3Ce
YNeZRNLYfZaRjGa0mNOudmvibROMRO41xu9mc9VABgX3tgkMM0pLX7PLLbxdcW9PIMwBxjt5CGD/
l8Q66d6BBpC2v3NTxfO8uvWa5V3mUFxm4jC37TgHuW+YhEVLz9anJgbzB5zvzXiEEYis+0PjqtSW
yDnrpNdTWeG1hPeBOokkyWWfcPYaNIIXG0XL72hoagx2lVy2QrJcpHU9Pj5IrkMDtEttQNxF+VvC
zmTbw3mZpKzIiArlUwzrDpJbtrPGHgDG3eD5bGIYaTiTT0ZA3XboMtcIw1rZbZTc1MnzsZG2TgcP
eyj1Zw/RGhEmZIs5V4X9U+1DZli8EcpNcsHuonxaTFSBVWYWj9G6ao9GsLYqegMqlWuS0BCmTwgk
toAccZ2WWTK/XP0tzb+bEdgxkcf8ErJ8n2DfVI/n6AZsAnJfisZQyuMDrI9IDJYtWjeWQ9T9aXRS
Xa2VUbN0EloxTEtwDrGHk4h8p46tbv0thPfy+pX+0mGV+BNTP7woHMra4oTs76pZxQTn9ph8ppMh
jjwDGfbANHWeqNXnP5NwhwaQluKS0F+k2M+zMNuwXBxkbQuLLw7jTA5UE4M9be4HINV+fZ0y4nXT
Wa9Lgw2WIryMEmVJmi2OW25Q+4tUqv+fPiP5kH4+lTV0BMxjT1up7kuFpHd1gv2RIg/2xHqnzhmI
WoXzdzwf//OVpDHtzucwTz8c7ONyY2XOhsVbQFbwet1kqENtiq7OYDkXkw7eklsdnPDoEGs93Av4
ZFtxLo8z+Ou0QM2p6ZLeE5WtyIzsLUYm6zcrKyBVix80HcWnLIA0Zoizp+yg30XRSeDDD+DHedZX
zm3/bZ/nqhETaH/vUvVpQtceJbzxDc65JfxxSKA+J4R7WLLHAOANq4KAX4jyVf/T7Ro24sZ/da/R
qlV+Qt0tO6XREdJMDabQbpCNxkj3eVdMskFExNndyTT91Z7YF40ITDdA3/sXqDur9o0Ad7mcobx2
k6n1fjv9AEnLQki6ruJc4MQhntdqDXhDD4tgvZ8j45vMo66vp97DQWxY313sS+2lcG6in7PFpmO4
Vq6DTyUN8JjPepYXW0M2YVkUrRPkEJALfEiJp88QPuHIy8Ku7HX7stL/kuYfvYMsrBnIR1hM4OHQ
zyB3slkop64tfUSCqzVV0XdAgE1LkaSFgjFWpbYO12kM+zc8bvFPPNFE8Iguh7C+Bcu/T6l4YXAT
FolMTiUrBERfBU2YnFAq2jWCcGf3lk/1PhIdFSViRUyiwRV02H80sBd3x1Ru4stxMA+gwpanXRsQ
XM/a883JvbvHw7cj3Md30keM0p9DI7CsJjfsORJgMILw5k2F9gsHTWkYatFfmoF9vQO1+QpSupdY
y/d3f5OwQ97kjlgYlTKxQBW25E9mA5wjd6Mv4nQo5J5Oc7AriDCBXmFnVe2mSKFUGBjorOnRvlnr
apkckTGeZl+rq7whODMuDh5vON6DmzrHqUZcesoaji68NGA0yMxiluM34juFRVsGUDkrBszFhyjJ
PNG8rRT784fJpPOk3CeT1Rhl2aJl8/lcYVtfjxE5CL9x4M5w4ZGUNWL8F4913Nj8Q3pPNeFE3WJ5
A3KEBBbjiDGnQDNq/KN3kufbIrAGplG7mLNtoRhNKXboDYUi+uqy45qNPKr2fHJ80UePMVapG6u1
K0Gy7RredHGmpbdOA6Sc+DraI6tfjkWJdQkNB3yQR+vAP1HHwLsmBltWaAmfwEB4xC2Ds2eYPOIS
aEL3SRxbceQNontqyWLsfT+lyhkx34TtFbPLiYZkIULSUQlExmb3I1JEne4xZLCXnx3EEYC1JoA8
d6HYlrOQ6qxuGoTC+PhJnnJiXIQM0RhWnu891NaoP4n9riK3Sq9qqj2yx0tRe81Is4a9keFhrkYT
SyrzRI/2jB2sQf54+ogs3TFhjYWFAAxV/Fk433zBCizvZy0+f1oxQVQFAfaaylTQY5tq7i8qYd/5
SPpiJr1bgW6Tbyu0oRfbW+RWAOXmt3s4Z7DawdbLcz1nOcJSGR/Abiz2G9JEeIDOCPwRhNMBv7jK
QMeqrME+VRBP2KKJafG+3hAcNYu2gxGjsEFAL2E3gPEk1DnpduebYFbIogYFPWZu5Bxk4IqTKYtl
pUDerXW46/qGXw3fDkNZVnGt9T3heN/eu70miTPittY9uZ4kacGHmw+yDvVNuqG+O620d4ncPtCC
g7SPy0q2InJS9IVF+PkTckaXMNaL1ewrL/XqS+xlThdxcedRDJxQRPk6L67XRU43eH/9eW6Jwx0O
i/5lNmQZ1kjv1ruYg8v9wcYf/YQora0Vx00Cs68jjLHwqPm/eaCJo9w0AnLtl2yXsx2LFrvoV2Qh
dWO8ZuPfjboPwdRyqbJDdhXHmahjDQZDAPVCyG0geEF85rUztyjNEdI0McvVb0ZwUcnXBDTCrMOB
HgFHqyaT1zaYgbGBAqLHIsMTD+4dcv8mWAAwH4T/s8HOtqKLeogFSMN2O76bJzj7ELUyXKbknzHx
J7e3uBSPSyODDfHPPm4aCIh5eZoA/HqrYcr4YAkX/wlAabtEJiB+nuq5iVU0ImWac1bCGQlKOfZ+
DNDN2Vug4KwNdQJ4nhIUUMUP25Mv8jZkNr3R8ObdPNVqzVw5dQ09FyL45utxF1xVQ6gExYtE7x3e
Usy0ktbpoX8s0+NgbZ/crh9Vf8XjdGNVB6W/olpJaP0yW4NFC4UQWfaLTuFybTzRRpltbX4D48OP
05B7E+De5geZHaeH9ia+QqNLMe9P14fIqWGA/e5jmcQxjGYcQ8iPWc6lDX0nTyNBZjt6iIowsEX9
oYzluokmYocv6bDM2TFLzD9FNcxbEMLXLP4g/hSliXk+RhzoiGvDB8tbIeyV+8r6kmyoBXqo7EWn
7ksSYrQbqO798qSj8WBvfTDP4PnDNi6Hi5+fN31nmPiRaRDYRhsJ7OeVantjGrYHy9cbQ54mntFb
EbcSU3aKn6fETU1WY0f9b4PSS8KJwzq7V3X8drAQtWPzycJhLoy1muQiHjeAvFv+enOT/S9OjNZZ
X89cS5iEZv0gZFg9eqAboDVbSTdv1bOr2D2q0Kowd1bO5jMNCzRylo+dRufZUlyBFIJmt/ELoNIf
ulA7g9/F8Wn25/ihtdgD55A8Z+ZOr+97ftaCmL9NBHXcvBjV96dkxhF59+L0UwOZt7JjmkUMsOvM
/XaN63N2FSOVnmuCQPTV8fjIYly6rNcuBXpytre8YtQH8jJI/xat7BzjzpXc/vSRg5iQDVDAJV+t
jGcmNZPDgFfbKQRUjgVxpaCtvRQsNLyIE1eu0kLEl5xY7BT0jMUCYofU4o5uyzNWjsFGDdgGnu5f
BxJBkXNq/4BJJnZ2btrgpOhdeCGvIKqgPz5drJWdpX5g7WIUfPDO/51E6I8ZpBjJmYKAq2WfukVN
GfId3xtPaNCgjcrzFivX1s+Hs7VJcWrlqVbTmCs5odPclGwNNl+FVW7Ws3+82ez3Dog6WCy152Wn
MGJRvp9BO7x0A2CHNLB7gVjGRokXAIfbuU+ldQrCPR5p2+XLIuW5cu3pNDo1m7Y56eb3RURSiX9r
MGTIQbsPnSJAWEgqTIIU65+Kn0N6tGZYQpUY7sgv4FtLc0n7UtrxbSdkztXBU6v0gOYgEWxOAiNZ
sYnfYvwgtjXc5t45JkD3dPx7lS/xnvip/f57a3/3EozRn2tQhaOBhUS1aRIS2ujtAM0dYmsEVUpo
+38iMtjPgknWov7MfQBjgG377fE8rPGnXDDmwtjTN6fRe8uHjITlzU7m8NjVIMNzwHnY6HiJRd15
Pz8Q0gCBWlWrzFgTwomkETJjmMEpJWCIxSHA5cO/4FujSNybLqCquXIgB7yWZmSoAh+yE9WRM7Dk
z+wlDSC8GAH0gH3SIaPwA3SBj8Joon+jtb4MOeHCfxhXCM7L1GzKPPWuj8gfGJmLta+kTVk1+Ebq
pMCXcxsSU1FqI1dsyuQrBUMitmRchnZIvRSngSZMd4k+qrQbLyzQt8/b6lLZ7i2HQ4j4qZM22DTL
owyRFr7Y5thC7uvhuvRV6b1QfRWBaUzRLaca/NacqN3ptEKGVgM4abG84kICwUtqdXbiy+O79jsn
2XUDzwG6jK4kk+p8D9QRcvoqILT4ofesJqQ/kXc1SE8iP/jXQ8xZw+jNZ+XjfFHV+JleVgLRknPo
YBk5buxnF41AciTplmSiajtAGQY4/VLH+WRuPgeGKjDjed7jM4UvODzDa2CHmssh5QH2hgoxhXEq
I724CRhr57aIcv0mMGbcpQJXVpEYkoh5v9YGQ0dpvx53PgirAvHsWV/exOJTbRpGsEjv+kqy/nxd
vTvkOfyvG1NnXh6oBgDuFqw1cVDTDvUq0q5wHg/qzpHNr3HISGaQFyY6/iNRlsBBsIVfEudVydlk
OqM4SHTjdCDvhruvjxGcTzOkDbnPbuVkc222Ard6YGOpwraNeQ+YddjCNOC5kX6JshPM+6TDoV6b
gX7puL5M+/CzDOJdGkGURu3dDy5lLnyvdQAsLOHw84o7vDe3jSCf6FqEoezCRRSe08FuJfrWBQXh
hjhnbqUB7HcLlI2m37ORPFHSAVAxICQMECsvDrOpAGGvgYdePukjmvcG9M/0ffBWXFcETEQTAdAM
j9zEoTDDsPo9VrGzAyINmFO2Frcb1C63dcyl5H9xuLkjxo2orE5LAIrOh1Tf48yqyZ137shqOScU
+df/IhjMrYxiRmjSYrsQpC9jAtIaZ6gScNWiOpFmUFIZYel+EyT8g8oM2/2e6M+zxEJXZ013db0y
16/VvbsDtToqQzz6RTmjNtIxQ6gNqdn9eg9vaa6Zrt9+j3LVil8l+p2lFkqvZ2L89hEpouyNFd6K
DAfDy2lEhyPWR0XVYGGHTeWm4xw2sfqN8ER39SAIbH2dUQofYpYdVKIMQUv0z/UZxeRJ4kaS+Nbi
oiUkH2BCsC9bcEsRKRoQiJLDH7MAvsE+tLxPSJeZzCbRuiH+hAth3gMsstOXNVQgUYsJtKK0CEZo
29lyXVmF3LScHklCbCSw9lZ9oJ/Wl8Yl65yssnowRWMq3W7C3WBoyd97uH43CjTLWfzOj2+CMb1V
w9Sbaqyy72RjWhZoLvou1og2pyoCXK0j3gykX/umuDqxVxa8ZQe3J+/9SvqOon6Zijuxyp9eMCWZ
wIOvMZgFnq6QI4J9DYd2sstNaqzuigYh2SKc4eYfx/Roa0eMAKylpERppanit3lXAQDQKF67HbR7
Wy/F/ry2TWXGnQw+LBQDDQsxQUipvUMDp8SgOeAsVpl56r+uRO7LnGB1w3JOUTR4PsWVm43z0zZ6
4bJJD4tFIKAx6T9MipXQ8uhonKbpXbR1LbPuRZ42V0WTfK+Gn38ReFtiaxaLqO4s5LaFNjvolBoZ
dXjuWSFd3aDj/P0P7D3e2sLoTBWu4Sgv60xzEm+Absuyz9EQd5JeEl66/JmWFcV/n9fUuUK7ZF29
s+bU+j0VZ0A1dycHi7SP9mpZjmVR6QuUhzj/H3X7HvzlJWW6poiIG238deoewvZ7V9R4NGkG0zpG
7NdLPt7feRTBpSN83T1trZUZPLsQJLUplMF52R2u++HpXN1wTVIOpNJfYizQCf5I9mbfW5fNnUak
70ACox0vlILkaqm0lv17+hH9Eg+/Gd7rg2gZ/XdYSwnON/TLcirMh2L/f/9BEFCvNkrrTqTKOX26
tpGx1Iz+uwlyn+vfvIc4NHyYI1FJyvVuuXyJKF1E7Nnmem5Zu7pFEhA2Hiro5xWzbF8fL+yzxdvL
lPl/BiB5bMQnblcHb0J4KrwIEE7IrvxLkv8RPdSyJqZ9Oh1FsQrsEzyLHS6uTgXejvWtBA758l1J
Jhat0GA77H6x/ZalKDMvmarlcMGLJjvt8npNfkeMILuEkAjV3hYnZN4oi5UAEicFbYY7uOCHylwP
P3erwoMoEs1xu/b0iY76nzQLOdr8kK/atGY4IVvklRF9OaZQPnbrMghU4kq/qVJKYGMj27k0dMeZ
RqkK0f3vRt3sAjwLw8PHXGRlCMVmIDHdJbzfJCitngQ2WW6zatnT2k0CNLWyhQfGFYV3LdeCQosp
Vq4GRuMWincZlQ9VS6M8DpQPCIyTEqO4CDe12kjEgNCjQ7S7HMvAJpICG7cwct9AHN97CNCE9IgN
KOYFJ7yyo3HIq//Ac2PEer0bra3I/CdD8nesjJaTXRTlw4kEiFnjyr4lE67wnG8wryO2qD5BAmtJ
YtHCDr0K9uav6eJM+KU1hH+gQrtIwo6ThVy/DJmEXo158PgRnUANLq0SKkXRnUKPUUNdJh9rudFv
n8x0XS00DwKgA/EV+G5zICDOkDJs5DPPIUPY2em7afZJPnDoXupH+zT/vC3hrVYYNxCBbt1dvpJT
DL9QtqUB0OSf4C2wK83qoAItIcJejJNHl+wiO/kZY664uuBMGSzVMuDxpXZBIEd7PCLa4fCy87DL
WPv7KKZOa2aLS7DGBCp08TSfQxbVhfZkNtH3p0CCs0X2fCv5tlnp6ZnENmt9DP+yLOujb3W1b9Ky
tod3xilFMHzHISoS6mzRnCm4/tDxlRI5t5yXEx+SL9KMkA8JKOMHEr8z8JGHLK3y+Y6nYDSzYY1h
EHPduA0G5bqaPkneymzdIle7pwaj6mmGN4DW0WywM8E3QrJMt9QEvmQ0nRqEdW62iNwDqM4kHvTC
dcU6kjKcSQYguc+CXXhkpW2DR2X2Bm3WcYVi3h3e4IQE1lQl+1wmGJsMdRtkCEwSZZqeXyvgZ8ee
L+1fFqG5TsAcStxBqyKuqqMwVJ+nC79CjRrgE4DoW3/aMfUprdNcUZ5a1LidpsbzrME3Xx+ukR73
3pIgT+XMtRUohn30K831spnh7VNnzZsU3g7aOc63wdz8mKbfMhifN3lh/Zjqb/4eS5u6cxfrD2//
edM8RAGdKFjq1IcM68LqnNv+vRQDLoysUJeSWELQ3Ywt06mUb06ud0a6GaMMgL/DVv6ANi9V1GFG
wfJX4bElKkezcI0e1W5r7Vj18yk3ZJUHQraMYFuJdeoQraHafSb3EkKQ4G4oNq9VtSm0taq5hpig
IlHg4Gm/MEcOcfcqAz9E4XZA4J0BeA+sK0w6tFEKRWGfAzQyAdTiX4LXlm+RFoXk6jrH5qE5RSlX
Cp9DG7eWqaLZxRHDmwBX+MFsLRgz7apGjEkaEJmo8KtKsc6yqPiQwzVBlBwe+FVEWol5I6Jcu5jz
6RDXk8IrDDAVav5leh0zCFNgMSq6ESdg21+oJelIYc4YCyvoTfc7kRxglex9moLf8dk4vIleHIgl
Ci1/mu3nCr0qv5XTgMJPVw7FPC7rH/PH3oZjvXKj7Y2moP33rAXcUdwwDK8q3zDyPaSVws7Z65fA
kCEaO8n0IEHQidiEYhOLwr8m/93xdeqgckKcxr7Dh6xiKZobNxqkhL4tNG7/CbHI+Rn5Si7A5REm
ArxmefSjTEzHXfFNYvMF+CjcN57cJMjVUYMaviX/K2Awzu/ofxzig5O59aCUl366DUczuQG8LoVC
xo3NW18J3hrCgBWeYHzTJ0jm/mNyL1fUO8/lk6GBvFNzgzsL46ZNmpuhXeDAAK+S9AT2wnWxErF4
s1pDj+2Y5Sx/RzW+fVGUngg99xNazjSCa2Z8GSzk8vqAktP6JZ9Q1wSgV9pDB8W0d6BQWb3aIDRp
kwexmfODZe6odaxgQoT9gA4n+PwaMQ/ziXkT8/Vj1k5oryNt43fU7vV6DjwuvGvil0W8J0HjuBxI
hsGyhToXIhUUHyIySLmXzjJp2dg8KCSVhysHuSjNlnSOqHJU9OFa91vQ8qtca8eHcmowbt91i/tw
SsGoaFV0tDWYwAdJclG0RPo23Wyn/Vt+/8zTsvedRO8tDbmMj7m0JgSKWc9zrIL+gAM519kmu8JX
19v5oYX4YnplDSEJcdk7Url1SJ0nmobc0LAtWwyWwCKs05qat6g+twLmp5nB4WQvLc+NgoTRWR3R
w6+BIYdG/XKow+GhUya4KSYWR2iQgUEIkQoUnDdv8Wgkn30E5MRs+gS8MvXA8GFG8ZQCYH0wtnsI
2eDt+HA5TeSC5RrfI4baJ0fosX0EF3DQIOiNMu+jufGg6bgt6gqA33alY/UNf5CRf90MBuGkV0LF
eFsLXRS24NN+tv8gNaYNZTCKvlGyIB+16JqlpD69EXqnE3bC4fquVzV2AMYhOBVVq+IknzyjQhjQ
GK/0A+aF22uPP16pFzhOvOXMy2WuzrBMKaKv315CfBlEKzIfCqjJDeGifhA1soljCmitQPkQMXYz
+7Vrdgr8GFIvn3aeyW4FZy/hXFPM8dILNUSBkL1cJZQm0xOoH1u9DNZgfolIvWtMjbUlsSX8EArP
faWuoVrKd8dNYqUBpOjV/PDnKtaKnXsP4cuv43o0acg2928g5yAVvaOMhL/lEY9miSsUM8ftOKB4
JtdMeQ6TwfHL2REbn4pmoNQaHpKg7Zev2Qf3NTX4gXf1AqbBxJN3WcYUMxzI2rH2gEjABKmEN+Qa
XvpbzW7+ju9kICMHtVpsmegUr4XHd9s2zxdSmJ7KOQV7N2KMeCH55+/nWrDb9gy1ZwPghWOuaUmm
eMdfmhwJG/WnQLR6Xvjqx48P1c+94Bd5o5zbNPFaO/P0kidLEKrTiofwWIner9TJl6c/Qkh7avlW
71gF9TxF6LvRlu5ZjUREgBkXcz0t04ngGnTwFwX11LKaigoIFJldHk2D95p1zPR/nTP7bBsov5oh
OTiWTxMfm8US9ls/KwzXk69/usUbVT2vO48hypwyfWpF799CVIuEdp7QjRtdQPsXoQbBEwFfsW22
g5r2iiZJQTZL8MJg61yG8tqvMAXyIy6rIlisTo/NyaD6fJslzOF5Jc1/o9FLUmzGOGp6lS99X3q2
l2p2HgDgcp1AbgmroUq9eAaemlV9KNK6GEHJnL9XqofRx4bX+q5q8dWxSLqcjGNApqLgdoK+iTen
AJsON29eUjnyFvg2RHg3b2itSeoOf/ThkQLuHADWBQIe9sXlAVTzUw7BN5XaGrlPpOcut/NbrfJH
dZDu/H//ImggjCClFHlk29MA5zwnWMMQxDPkDmwtitvUh/YLG7WIvK6e+JTlm3S/3tPNRJ07jT3y
V/vHXRocgG1g5Ph/QBcQSvfH0fln2LLajZU0R1Z0dB3dMcADSsM4Ed6b099PJCNlff3u00p/m0eJ
eBOXLTvMdooDe6JcbyY9ZLWFTDRjJMGEGOzBNr6YLSpiZrSunlMXiLsGCcbmzfiW8M0x8neY3Zug
fHc/PyVmK5HcytIeqbyY2kRc5jQ7S/BH/8stwASgV0hA2zikuAb50BzfMGHuwCsB4ac3HKE0A+VU
NxikNP9YUQQ65+xzMtCsPY6zDd4sz191ZEWDuCFhyrVVq8nJQOYPXNUQ8rHxwk0R7M9pAtOduCBC
w5JY4CMDQxm62bW6i4aQHSMeNfUtP87YIH6tGkmp7dWaVBtL0GP1ZKOOITlZ9ePJyM93zqmkY9Aw
UnvtavU8fnsxdRFXSJ8OIF+9Pd8NvynVdWkHohvmxiZ4AV5BW5plC38MwvjCMuk3uzlA3wmWfhxb
CLmP24le8dK+rtoPWfZJ0v9BLtKvbIcpoMeCfl7QwijUZjapDLmEyhRDdzilfZDqX3/l+0wI2YQi
ZnNqfXRR4fcfwnZIBW43yoVL+Gj6I0ApvGTkRDqjNaY/7a47pH7GLU8RYIreTnBl7ApgQTB7lP9z
b7s/Un7Gx3X8E8d52hOZGaOSiftIylv0bUgqdjlWqd7z597yck08AvzWG1Zep3Rq0uVQ961LF6qB
3CZbejm/8qg2LttS2y8FJXdQGU/QdBpnGV4yWkNC/l8wrtsvWHkNDsjH7k1O8y148g00V+JieL+n
hs7FJoY17QSnOJ0gxrvvi2AEk4wjTcayRT8xyMZ7Sff5gTzx2OXXFolOAnCv68vAtIdyBBzsQ+/v
WwkkoJxLnpmvK8KwcU+GVdXMIVsBPP2O9oE3xgJ1ZgZRqm7/ohFkR/E4+qnzfZQl24SdO1ZCG/p1
Wrbovk54bhPEOCH0F77YNa9wsrMIFeEwrg02VnLkX5/a01PMusa5wehaxyyBM53Sjh1aQWUIQJ+6
TwT709JM9z0i/cb6+csnj8aId4+wd7pF3H7GjaVbCbw4Lc5I/nDdQOqYWl4tYDYkVOkM9A0i4mVy
IyQo09jqQGg2wrHKDjdTMSa0lXqkv/hvaKmce36oB1wrmt/z9ktjj/fLD2tImtrupNXdJ0MOXtKM
wpNhj570AePZm/AawJAEw1Yu1bXeomWNiYDZj+2Y+9GWMKpi82lqzbbfNOdv6V6+COHO20iZ0I+t
NNuoabP1yTIA0ZGilBR65xK/fYGJmLh10XicPwg9woAlyAXUgxHpY0xUeluYqu7fRnxswbxs7Ywt
pji4sthocuzuWl9w8Bc6RCT19UNa1M6UrMpV53HYpAeYpAI16aS+ZF3gSqvS7a+X3kI6fjd9C6UX
Sk9tGj1YG3reGbMFjfXjYeGNjfXNXSn6ICuSYgiDvTlOq8iv4Hr+wghgIp4uS7IMniTW5jAPzlMk
FnvhBIMSg4Wd3frHK/fkjC5Dly87RfkkB8bfWRCYxOYTHe2Dqabyw9f+4vSdTzK3/hOOIZdJcS7I
I/t+cEliAMg2yfNRza1kd7kE909FOljOkxEIQP4BTWF/DrLSQ3/sDXQVOT6JrXetak4cZOutPWXL
ID26o5uz5cflZXMXrULH+a80tpofmqC3ZQYkKJWmak4rzl8zJRLXmnkTaAaBsbm3+YmlxHFkBUzb
FnpRLlvNiWRKezVNuKg/7Gsp4oWi7aYMAkUI1cXsswEjvmQCMNdBuWmNSYtYPc4/jyOHepOjyazU
WwMVzLE8r45iiNHSnOVRIbGGpuheNOaRJqgpTDdxAzSZVrJ1NM3NVCuGScm+xlUaak5xkjaq9zSw
pd6VinW9ylnlvz0KkP+ceOu3f0bufB4LvJxAQWxGXox/UTN33VvuXkbmzP8KccORiuZUt0MLI0Gs
VbHcYWsK59pjj5uIGGRvmztE9KNjRlharRrcbvEsRffODWB2sFmgguz9O/JAL5mckbRWbtea4H/h
gtqL7KghAVecVoBPqNLS1Hb+JtTA04DB/dB/3yltt0ZM1LXqQNlEYTIbLX0KjSa9w12SIN4tJbWX
HGIrAAUwaHF0xwMtE8Je5btJk8IxMLEpTqphVRFDAHdqAVrT4NPUYw3J5rro68xv34hurkr7UTlo
mtjQYpoVRPMQa6E1ZN85ipg/Jop+LyDjEI5lrP+nrrTtO9m6wDy9NlG3cZZDy+5QrGXB8lLBSwgX
6zNsiGYbfxP+cNjEZA2JsEQxGWyxp5Ky72eLrHZ1oNNEbYDl0VYalNiHEtNLvXTl+wM+d1ReeGrt
F2ssmMjgIUoLv5hGf+HPTu3gUY0BVR+ybkILfCqlgOxb8cKjUJtTqsIhIcuo3NgaufyD+aAEtg8i
oq1rLaLGgoVVq/O8OcyC5pTBvAjiJZ7pAfcS7FmxMlCWd2imcoqspeVe8917vjHzTvmbZkaPKFWs
pO6IUxZVwSs/61OUbEsX+Ut50bTCFt7zJWBCHt4Zt7HziO9cF0wsnxtuJybA29MQ3XNF19Ud5mqK
qlFnJvjlTLIzvWraRO19Y30vWwzzF4b/XBZ77e62xtmPNXNUFAUMF3NYD3Gm880c6K23ypbL4y8X
oOz0ShV22eZe2j7RHJWiT/geNHJ1fEatsb3f/Y920/2sLO2tvBiJh0lIwz3fvupLkcF5olAr8HQ+
zWOVeUHCUtLyZWtZ8X0pcNq0naPHpC1n9jXW378hZtHOfdI4kW0qt2qIqnA0q1FcT3LNHRaJrJlk
z6Nu9raE9NfB8dN+JsAE8l/KyzZT23A6Yo4rLY8Omxag1obdJBdYiduGamlEEIUeb2ZlNisMdAlp
ieHAXCZSflow+FIXX2ktOew4I7eYnfDwALHiTwfW9gEhXIJBnZrsSJ/xtLt6vb+3Hv//Sm9OtkFz
NSzF4lh7ghzPwtBJHvA4f3mHtqWB75Son5kPEchijrfCf956eLbHB9SlKYtUM25FalSIvW1tZunA
KPipMGdsbasuWnIeLyenMjBceidYbzp7NfcsxvRfMHCmkYh/y9g+/ovmr58g6YMUMD725mPiUsEE
okyXyHFw0biZfqND/TxaqJxVkITzYsQadCDSbHrwUyISMrblK+/RlvKm68lVvwOHo5yDaorfjRFo
NYsjeQMHiW8RN39HsucoG/+pQRuLxMLaASCZKI3DBH75qR+a4wngr4pJG9+Ht+rFvluUGxskxDcA
/4dwF+XKIB+M5L+J3zvoRM/haQWYOqJo/RuoZeUvkLyy7XDM8XY4BoEWVXdhiCb9+8OERu9YP3in
3zaDt6Mh4DQa57SSTsgNmNHFTq7qwGm0XnNr8lxGiEzw8ZRJYMx1t+ZdalndylLXYVDsBoY44zAF
0c70ockz4Z1nIt5d+7RjElVh2V0b23foMY34jMM4kAsoixGzB13Dy5xGh0/bdrSRftPHaXNQwfaz
0PK9XttTaC+V/VXwqivgHh+CpqcMkZ8QxGpo0vN04+PzM5w9lXZOQob/jm4Hk+fGbZGQNz3jBsvN
s4WF2uzuQ206Ham+BdrJqexQfr0b98d/9C4ReOyHTyX1k+ayqCNPK3nGIcEa4KwLtxCpTXNuxWz0
3umak8is8uMBFx4Mtgc8oVlqxGlpzW8mxEv6gBDXGxzkIZshp90gQHuKMk+D0W3FAWIFyxXCBVSX
WZLH8SiR+959ZQSvwKcZpOZZsusb0ZXji57zIvHBlwQhYlIYBFZRyroCgB7k0dCk+jIox6iV/vEb
BybZ+mc0fR/0mVm+9es0PLmBAzINmV+TGb//+dp8ytipSWfmqcL3DepVsZFVEO1JqmskYpp/YvR3
iK/GqnXGYpS3o8vWVoNxXQtmDIuMOW05CNh23FtORFQirmdCejezZrKwHSHKXDIgPtEdhCajTbNP
cJI69oSkSbVdnAOmGIaBHVbOFTfl9PGPWC5c2j0KdYVy86RdmE8gBiZarNm30F9ylzu7eBLiUopV
j0C+AhGsuW/yzUWE917MQIf7tkU6s3fg6cQMGS9WjpqmsyMW2t+JXNqmz7+NBR1/vYMpIIEmuQVL
KgYwxvK2ImTudroPnEWM/7/8Yets6ZCcCBhlw2At+yMaK5v3FC5RYFSMmr2ccd55SdbpHSmxXydO
s3+oMamK4fUt3jVf75fskOmDKaRGq5g6RO4GYlokkGzqaDiQxoov2lf7bjOp0CGejQGdWTZXPWZW
psMOJl+xzaxNkAiZe5R8rAhSFpMyTvFAPiyeudnaymCOy88YXYMCYar9+pHuhet/yXmcqzUsOSpK
gmDf9saQP2ztRyjerZvu/woLCE+PCID70sFio5x3U7t/RAcYRHEzw/7yjQ2Ttbr82ikUQBepxTMV
c/wPtLbqv8y4vQePdmOK529KytNl7BafCrQYlnVmEtOeC5eSp/dJWYuxy3PP3P3wYLgrrEXtX2a0
8rwhbB0A9s7iPwyEYEUPvB11sk7uSW3KlE9dZ7QmqpjcsVucCfJiWA8PlQI2/7PvOwtobb8pprjz
MNaJqRGI9tuReniMbOurcGmeJ48lLLNmilWSBlbV7qfmDZDHYex8dp48TxnglvCffGBzkNpop+n5
ceCNTAH8c7pjzfTkTYayLOynZetWHeTmxs+xDwr7iRCdMPBbx3XK2/RSpNpKnULGbm2dq09Tw6K/
7nmMd3P+E3KCDXo4zbpcoVpuf76H5ewIT+PKbnuFVmlB46p73tAsi43L6kIUrZb2w1tMWT4Eocva
90J+7p3vnr2wakbtaIHSaSM9EkOC5n5NSbknmKZlTGk/yJ9spvUHVqeRQmio1GwHl0eIXjS0nCyS
EMVd5JWRwwhpeDqTtwfNeMr63xqcRQ7RopD7ivygUCeIvS0ehyJmitlNSt+/K53BJ0gHjBnbKsmN
UJEg8ury+xWsniARAnhnFfxgr5oezn6uqWmx53wuFzmGsTdrmMw2Nbmc/o49u2sQy/L5nEdNM4+K
u1UamAtKpD2tB88ryrl7wncTkyWrtgMTe1x9ddvxPT+c4WcIoWOAwgSsy7JftGQTtAjW0pHTZYj2
pY5YwRk+lz697EsX77V5j6cDbPq11yXT81W1dnb/SyuH6w0CYBZD5S7GfF+rr5AsCPSFfg0EAp+H
oEpdSs0w6HTc/WYxG2FyXaCnTA6SLwZUvVAWPeKwg48k1gGTzSXZM9TrBtVApW6sTPvtE2mtyZe+
BLUCZAQ160dvHmbVhaN7oDy7xsLJCft7D5YgGY6/yz3WX7T8iA3HIPICCmfJTnllEpfBe+oaaaCK
tUdof/yTowL7TpWPkUqsqVAVYPlF4XfQfJbpvt+xRg5l1KmrqUFvutf853ZRBiEn9G15fBsDhfJb
2BFiDkIXCLZSXZ4tuPKzv8aUcyOYtF+L1BWV3FCQ+EFpJtn9OlmKEmmehrtwhvvfmfxRQSoe5LEZ
kp35ddngHVIdqYy1ca6d9bZvTwKou0XygFzV6m8ugvEL0MzIGrGOF6hvmwgZnbQd6N+/2WscQQUN
/W3k6X0HJHnBZlbQfdRdirkFryHmjLRykD/4Ile74iYDS2Bgpx1NzvKG9dmEPdrq7BT4dqaB77hg
pNz+yehxKWCCXgjuXgmxByAWLaAmjeqqoEqwkYcqAKKRER5FxrQsFvWZmwfinMctOXD+8tSrBw7T
O7yzAg1zaP6cVy5Ypk5gArs9o0QWwBwEi5nGX8QhS2Nyqskim9wVcPHp+N3J5UKS/7JsfykWLoKG
bYxfJYVDKDDxExH3fmgMqV6ZI3uQCLiJ6YORDl8UoZpe5WsZYnsjV6jHhJ0F/6kxj6zQoKP6Giiy
3GiAUfAwcq81oxBkajHufFRuHAv8ZXlBczpR0JENN3/KEpMcJmlShw7fEVF8vYAL3kiF6PGlEdRD
cLnIPWeEK2I+l0bn9G+YDeZiGO7CCQrGNF3krqvX9V/Kh/HEfv+Gmuyygch5ucjtp9IgrUHmqUB2
p2eUi6CKf7kiCG/3KZaLt3nGb0E7rRYP4Qg3kar8OzPsncBlSKshuh+r012Qjkd0zaqlZLWTnQe0
n448jHYPmcftWtn9hd33nYD6jmRvqtSYAI+iN32SUrd4lT4dQyjTloIVLV5Aru8jB83DqonSEBS3
+2vumBxrwvb/Ais4ISk7DvBB7Esz8Od7HkP/YeAcX8RyY74ZNEtdlNFRh238i2VuPTQ5pomCYgbk
46X0kpBPr8DYzbELgfMt88rXxyyvzVJrDO8MftBigTs5wrE4aGR9Z0he0q9vgqOes2WqdSVLLYMF
3j78IJg52lOM7rsKSgQjq3/jYM6ZBhO9TGHOznnsFyBc4ZrOd9Pd/A/pUIBLYrarLyK8aYZt/8ds
SsYN1xjiO7+k7HBqhbweCPZXa1jvYUsJlD4/P1mHRYDNUd0s6cIdO3lkjclxxvY2zdVVwY35yphn
MIxc5Q4z/A/I7S7BLfmsICZhStHax3qJ4Q5DkNkPioMVPJkLB2BzlX+U0eWVZ1yrMfuXRx7+M3mO
KbmY2sZX1WDGStxoemiHMDaDIrQD7lYsAmXGAtLOTI1WXU8bZv2pAXpZ3sZlhP31Z27PzTx5p01K
WOLgPn90XjbkD87Nw8TvacQ39lBfdNYoZHbsTUqy0+n8q9ZNsdYycz1n3uFLFvQLTnd8vHesZtzI
NQjBLODz1zdWXBnBGleK+21DCWRmQo0Sf4wcur8dzlXhbfPf/9Ye9CUFgX7i/9wGnF+cI9CJgOaU
zQC0/NMgFPBVZtRfZEikTUQZz0gUIbcQwvidM1Awe0fB6aeBayIxEdHQKZYfHF5SoPcD5ZxCSpZ1
8f/St3Iqf+2CfkIs3To/3GiM2OU3n7aDA3Mr4Jo560rSGDGZ/J6FO9p+j9rSFuUtKiwt6VcDbziP
l/EjbSYWrOhJ17JjZDNF3fjWyeTkRYQBEcjqKRR4vodoZv/Ppvn4DbY9/oiFPMeq0dOeZjZlVoCn
Ue8qqf8xs5Y++GxqjAlsoR+67jvVvb5PJ1GMWtAi+XeBTJf1/Yk5oXWr1ROk5dGF41QQJL+hCu/v
Zhu9Jhpts3MeVfImAP+8mB5tt2Hp80/1FY1wl8L8VGT4MvRkOgyPpYbIuBj1XSty1Y2rJH5dE4+o
HFqlyNFrIUyR/FFL8gs/uO7gYK+MJJQi47B1GCp3rWKgX2tsMlMwv+PLLhm0DBdU9juAP1H807QA
7iJOaw8egkWHFIYr5mI5e8tYl4XpKBYHfrSIYdJZA3xjwnVMrKYmKyhgUbrTRif9E0GmPX6AYU42
w2mLKrOtZ9mbjGHAwMu7buM9qAZ2CT1EqO01BpvpYr4og2GnfKrA+dkt8ZRZBpID0Lblo1Ir4Cng
o/6LC5+DaJPT1bmgVruIE5fSG4xvxz8mYkoe5UA/XpkeQFuovxTacQjY4R18P5U/7gLHD3WBBmMl
DgBnAEG/63/Iuw5glFI5B7fg4XUEdnxX3trzRxys81UrfqjB/ZKzIC1BIXmrxuP5yxv9THPh53vn
SA3EXwyaj9n4XGUttQjw/sATidm2KAolzlhfHttd26KmGQf57HNe5JDSh6cv30fFC1/8sGwpRyFz
tdj/OD1MfNq5N5/qiGvVO/DcmRmEVOamgoNUS41RuR8r0FC/tcUfHcR3I1OAOlLyArBY9HM7HGAC
TbRcJ8gydHnEXK6SJjVhC6K6ZAx80DaIWbHi/kXx5FvXnFHu/wQ7nv+XzKZ3GNRw88TSImW+2+89
st4e9UUrYtZDyK60ks86Y56qxyiWS7zSCKQE00iZRgmBcdVqC0YRAo+ev6reGgTBK283+voSKkFF
NXUO0nEljk9arXX1xHLdFrm7KFEZu8PnNfHkrR6Rn4h8xDcES10MmdKGUf84/3u3r6BfVVGERehD
85K33cJ8D0d8Npd5ZlDF2Il2KhPcyoMf5KM8oBHkla7FUGVuhXelCaKUcT1WJ5FJhncLoKXiAyIP
Ql3VyJMCAiYb+BHrvmmjErInpJCTIyXT7OCs8jPsXb9L14TNIgJLFeVe8DythfQDlKC1Opp9pByz
ZQTk3XFPjtUaVf7jaQBQl+zBD18uTXFH2Q8AhO5IXSAaZqqn7TT8sWkOms2vx6jlSXA5cJt0itVt
FL4nSDXyDAqhFssI+debfQxpjWkLLCqhOEIoSWs3gsZ3pLek8txX2nO9B754Ic0cTjZHSVblEV1j
qmE4K3S9c6ACZw0EvAYGgDgy+6Iss3Olet/W+jwLQCO7D4iZgzpTGIiEn8GMYUHNS07GNKcSY9pa
O76GruNZP5QYtWPwcF6uziT+jLxNGfT3YjHSCHpQzJPzNhXISmvuLnewTi5MMnj1p2bkxQ1/gE5+
6xHmUiWqcLHoDu0eeuR7UjZE2X+QzODa2tbenhfBFAQyf6//aSWc5krEwtkLCr08I3M9nLG9C+yi
93T0aMjVgK4+GK3mlKdo1ckIQopdT2LlphDXb/DRVYYs22SNQDfm9piWwmdBPpeeXGZ5z7vc4bHb
z/IDNgO7rzfei0M21I+iRR/OdXEesibViAddxYeA64N0/LT4kg7vQATxqi3dsapqdaUC0ytLVqFK
+EJLSTmw/wOXbXfCBfJWlvO7gc7+/urksiD1DUm4Kl+iulnSZbSkNSlM4Yd5DBMEAEAfAWwJYwRK
VrzwDM08EMDWJLJcxGlBqh2IOrK1ZOg58m/ypT9h+JbbgXaToXaWVQJXJMcvJ7iRHwHLUZFHdyv0
KYlV9qkGIrCL1UpscQU4hjxrgVrxHynqAy3DYkmlWKe8FEGg3HiUee8J80i450AyyE97tQsj+VdH
jFeJ7kv4Xj0Dz1IsPIE8heSmOME4YlcSvzepYZYtXoYvqTe/Nf0/5kl7L2mpSs8TWJIpDrEwCXn0
FbzYXgmB8KWDKrW8KEc5s/0veZSwM8GXxtE5xP1V+TBujQJ2RBVRnk5AxqqJ8sIyz42Ty6m3HjPN
YEB6Eo5JlvnY0EzwhSO4CPBWuJI0PuPz2JARPDGomz3A2qwjqMboSxsfx5j8F6OjBKY0saxAHOhR
iZT1wmg8FvHveMc3CXqC9EVjXxrO3LuWUBwsqMdlHtjzZ0u96mbZkEuvDpV88t+AFjVyD3faKbMc
tov+Wwez/8wgOs1Kl4MSN0EYOF1EoMKxQNZwf5cPFQre1LvB/JU35TmrjBgl58XUWIpIzBDPlRM3
3Ah9w47TJVbUscgMKFGFZe7V0RjLjQKkwSWqpEnXgd6K1ACl2e72WwOWISHHEei3rTfKBKOOl284
42ZTLEQI26WspF1SvnT0ub8QnsRAaksNb6bAHMiOED4HHfKxq6Ub2VUyz2CAXgrql7ShdBg69TW2
8SLghilholUEtqOiqAS3INPeoNJrpClL+CUVGopN4mJ4qxM0zSlAHjq15TvO1qs5RPk0hmhNE/zQ
6Ke/XsD2b9eWJ1awb/ALF9mNWQdb3XQFH2ShO3aFpm16CCyno+UV/xLr9qsHC0pf3sBW3+EH2fwY
B4bdunVjkhnLfpnus6ZBTcyEoyNrYE+uJUd2JkRtLGT40REBWxgY9a9OLqii0QcY6FF/GGtoIsDZ
G9l1jcm8ZZNcFogeGiO3Byo2EmXX/OuflfhDjLMNFKxF6dM3Wyk4ROpDG5UN2XFGWAbZRPReIdP7
TLSScXl1y8fAMUWxrH0gopqyW+S7ns8UZpZf/bPAHUdecI7ntUn3IIIOvzZNRBueIY3+BWz/Oitm
R5EE6Z2EoLBAv8UWOS+mho5mKU4TDEZqrSRT/BDgpQl9KmZ3YP408/fhheUp3x6CqzCO6f6T/N9E
fP0xLLxzi0KyeEhpmPiD5c3dGMsEkd4m7TKXncRhULN1lSm6Snx0gNG2yNdqePne3yJ7tibuZl0S
wuKo8Ug/STdJkHVstwQ/YTZoFcNkf1PdFL+rMX9naAZAyhpwU8lJ2IzBNCPP2f109MRashI2S3CW
MEtw5NBXo4J+QMxJi20t8znbjccqZy6P7ia01kFNTMN1MLEKNTiSrWc0EMPWhlpUCgT9S4rlltk3
h5jrCUwMxeQU9lqfY5pV0PtEWQ8dTNxh2CpMieKm+JqtgtDS+f93RK+ygJ8xNnHvGZIJsYGi29wc
drO5bCvYDEfR1kpjdBbVpLNYsHr8U1XAK+lhbxaEsXbdaieczrqfa+MIb3DdcTYVkUmlPt9nZhGv
Q3xQOf0XOQoio4rZHYxxErv+r9vqnAJtJ8QFJG1gDye+zJoZYj3s0sbs0nytJQb6PhY58tVNUVeq
7BZMcVrANK8iZC7Wha58AuCBDcz/5TscETZ5EoVzN2Kcba/jZG30AYE8zERoYIeyps3h8OhRmYUU
nmErPyEYOKivuCz6MrRAkUWIdZah/sHkOyM4A5CZbwjg6zK9xWd2vUckGoxrWFxV4isAUNgtsxmu
aQwuu4A0GA0I44ZlHlp1SppcZBelHZQ1DGWQqbuvEGnU5Aee46thnqbNqZpMsNPmEIFwGH6nl4Df
NXy5L0C2dMJ+pcVckHgHbq9yOIJq7mOygQE21Wo/9aydiWFxvYoECzs9E7py0KjcGl5gjEcSDKIM
ymPPuWSEJIndZ76eY16mSxVT7Wr6W8zOywtlbhIo3P30eF/9wLEUGLDGS/VvtD9UfC9Ktkebsowy
k2bRKyDvr2jsZ26bf0G5DdXy2l2x4zEk1y5jJawGSz0SwphEvre6ixERbFnh/bTVZRR+6VTi3Miv
BgPUlT031kUr+Yi/8kYvD/M2NIbF32hZ1v3C6XQjISGP6eW9Db6zY2LbPVAUEdTEDjaaWH3ZHRXm
OWXMxQc737rhYsxZV1LmJDm/90ehtCCr/0vgactPJO2KVlMr0QkjjjfvzrB4ZQMT+wazgoqud29Z
d/nrk1hq2e+kFycWiT+3muz8qao69tkmJo3H5qrkXZI1UPaQByBSYL5JKQuQNnqTGUdT+ShENJY+
NSa3YwKBOzBcYa6JZuhWN35h1zjXSfFKDkpXj0tiQZ8JX4pH+V4dhPKUQSROVH7iZVZlIh3IM5Tz
qUFqerdtyKOZcCmZiCy/qmN0P54a6ssI9M4LxfOLNHzMjoircSvJlxoV1kFocHtnm/Opnob+6mJm
UhXwYBC4aYZaNbSrNYiCX1UhlmbRfvhsP5NS+Kz9b+Kl08D7i5b4tkmap6STGRMRRSe0nMynqaj/
PJ2ZYGP+5VLFR8l65rWhYMonWDeHl84OTVz6e/Rq3BS/ef7xFh0yLWw4YrXCH602l3MBGzEnvAD+
doQGGiyqnglsPP7yBmrFFaWJEFqYdl9EatuzEPKLqCaa1/XA+ZXxTU9IEAXZ7+TqUSB9r/2VnPTj
eNfK7fWTjhpd2yn61EEaJ3vDu/CqwrXnMPJhINSgsN2gF1lH7tj2S6VFKPUX5gq5g7L/R4/ZssJh
yOPkc+/Ms53jByeqlI4X3Wq1fmXKp9cT7FMKZesr8HDSKG6w6eura2dHlbmqgTdD1RDF3rX45S+K
0QyR2MXEnXmqgo9FUvMyxIfTjQMz0PzAXjQnwQEne1syybtPeAPBmIikHmfeYoW8ueKs1jZPgwNx
dzsYJALPz+z3LammRql/A/XLS43SIL6qM7HdTaSFr5na1X+rUXCgXgzinWcedkDQ8SxRC6JE6NAu
zEom/SHUtx38jW2Iuv/8W+8pmC9WL8nZXnuuGqNDlm34xM9I+xfVT68dnKGTKPaplimO46FgxZjV
iJWjPVLhxQ6/oBdoPFj96EdfhZ9p/vdkOzAChTV0TBLawjGZrU2iURv+0xM44EGkcYACcQNicPME
fcY/tlQ6H1VuYCVrk5mTEHqeJ4LND/imOvPMZC5kKIDwFUan2HVEnqn8i41hGIcqZQdAnBFlCmCG
wZUSN5nl/gdRa5tFXezm1D3x3rSZScPfFDRHk8QtKKGh1iFzbcjQiiOG5uaHG1hVwNcz4LTdOCmb
ORQ4wonOJybQB1f+yBHQnShNcgzP7RLnoyNgLMyY1XQZqkeHhEuBQbv28CV446rUO/VlBxBGNmf8
koVjb3yzgL1/aNE6v7Caa48cbW9ivUyiTBBBo+oPrMiWGtiru4R9TFlTFd4p8rHPies41esplg1Q
pfNynj1PTJWxnnZEQcu+faU8w9s0WOr5Al+NYX3Fd9UYa4CXMvgmh+UPKhz8gGWO1diDxzThw6iQ
cIz770ySzZter/P97qbTKCytqQ+1CoTuspu66YLnnjGVVbbuuml6ae2DxsGrtl5iBR9DJPay3bRe
GrNWDvA1oaT4UCfDHtNkeuSYBtGNXrli+8UIPzBEABNc0FiJqvKBh6/YLaBJ0bmzPokXHqnkJ42V
2KLZgf+jdIkm4K0BFAwXEyQ79/tIi9C4vLgNyJrULaJDrM96a6NtT5CvWG/kcCorGTO4L5PHWPPP
7xEghzWYGyAsKdBXyfH9FqOnFK3EmNF/HZA9RpuVkL3AN4lI8BwSecX3VrlN4rn7WSoyYioHhbcL
9E9dwG+plmUAzJPnm4bsLVJ2ykh6LDEpHfbc0PFpmP24MYHZZgaRAWuHVgI4YFb9j8B2EsxnVl7x
+glp78zwthoesYwHlW2Whg81KcnlKpYJ2k+L1twkSMK+KwHyhdV3aN0D/o9IfRAcwZJcdyGnQaRp
bBkMYkO57NdPPJEe6do9ZLjqSy/5bcD5O0E133fym4lroD2Ip8MrmC3aA/nYrM7kQgWkYjRSpMAH
vVwqO2AvzKUfkPM8qri1h1/9wa8p5V0RoIc9TtOd5qZ6JgG2ppKZVQyePg9vq4zAFqS+3GUcKsK5
eV2IKBWaspS2CbmkQHxZRNjRF/IISvmuOWc0j6YPupsLl2cgxGqfh+nF7NmM/hElWWU6w5USGLeL
ikTgVy28DzuRCcUzbcsjT7GAzOcwkaSJ55o3HLZ+NTibf+oUrUAm0xKHfRFqZrNWc3fTHTAPMc7o
BC0+KT+NbtyEmamLXRPkFjautYbYqWNqnD6fhnSA/IkdIg0WBEeXDCRXvKV8HKGXjVfMXsRox1l8
aIfG2rJ4BosplPp6zoDqS7MVgb1aYf3cgBIyWq2YaQla64lkL0rEV7P9PV8we66YR6blBYG5aTFS
sIY2EOevppBXktpMKKiszKtMK/uwdoV7KzxJnXBoZdMJcMF206+qRuqhWfjmSR5x0gycyOtpyx6K
85zUPZzSi5t0HwM/FyDMEQVGXrLh5dijX0wfMewKq6lyoCWBU8JMBlc1X9cxqFZgl0DiRkBoUD66
jN8E13dYCWKPqxerBI0jNPVXrre6KSd4R25SBSuPiz6sHqsiFJeTJDjPQLQ+Og/flX7CEmquj/Bh
L6e3XUG6PFD6gNU8XuDWwHtKi+1jI2Jninyof2qVYDgit5HuaIQHNxGh8/tnKhGGG5ioDd3iFTmo
aER3GsLxh+tAdtdtuelVAZGjdPQBpasuDWE+ZTL1rgUV0qN6S2Od7ji1dkTSuZcA9h46ZbvkCmW6
ELhAl31+anLtekmnt4PwQtCFN5k82aofbI3Smi2/5q2QtNSIxbUy+MnMy7hPiHfYjB1Epp14tOHf
NIBPh2JX+Y7GdsBwWFWp3X5Js/o0nBKv7+wASWpZFXPdJRHLB2MN9no8AwKKuSHaFJvsfQlYXZfh
VoQcApx5FYCvRvErmPtxk/umYRmKhjDNQyT48AdUx/HOQdonyb7P7oVx2nIItgCX9yqJGFxUylbd
4glY0BeNmLXsrMqW9PhPOwEF42uD5MMQKncoS2PjbkGFGHPGkresDlNMn/jqUbf6LnMPExvKVyWU
ibfpIapVCsY/uZyG05qYoCB8fo7DeMZylfyW7QGpyds2rYh9Eyd8c+WWTiqgxbSC36QWjA/S9zwS
DAwRkujuMdmHaNSFegH530KAbt+sUrBvR+SIglI8pvhTJkFYT29GQ2Ksl2gz5tAlQv6ja00cEvnC
Ioq8mCENvvjauxpKyVdEQOcy3Yyd8iOhfjAr41OGv79QzE8PdqdLeYJYMt7WJswHaHz3kgqt9uN8
hO+2frRe0UgtITF5RdLdVmVYwomv3KeTU2KhJvfVjP0o3aM2l/uTSDcdjPjzCj311V95g9cmB+Rw
nhGPFV8NbGpa+tr4tTcC1xaO58Z3lqlwuCkZsHfCwiqd6CTUQBRGKqM5qxj/dCVLB0tRTj1wpTFG
7euSanZpesoCmdD7vaUD8nr/5gbtmuphZTKHb68ZJTTeyieDaRPGhzPVJkI3gSFyEzfj9R2lCGCr
mvwNaG+GtyLpRiM13AGqTO2mQ8pmqz8BURz6rlXneK6EhQz4hCnAbCQGIRW1eYhCKd7MQ9mdjE+k
O4lOLNA+EjWyGIiViYAkM8mjQCgDQhZcWcYFlX/TVKkDTTObrwO3nNNiYrJVBsqJsLSbcE4PjBVD
ZOwk/Awlh4e38r6b84D37WBObB4oDxtx/IAd7wXvfVDUjrph92gugrUBJUYVgtKF6L3WegoWKH4O
hX0Iy9buvkhHyB2kse2IdItMVddqVcGgsdNeIxxN2WcfxyA/xZGIqLBIABcVai1OSRFJkzN9QB7j
IbHj49zO+lkQPpU6alwN+XGjKDCTfSeKbm+qTlVIrqAWZPAr3lBjBoj5SK/ntKyhSERWTr2Jz0vP
uvbTbUgdpa+rk1p7i7nGDKeCnNRtQBdTv2MV8Ks7i2sVYkDgdMj/6pSMDgRHINtTOprHNerH8cky
Rf+3s5o4jQfLo6/yDgxhiUwyYgSKH1U3JlcPN6iYKHka/NZSGaqnaFK1zkGYKgxxgOgK4Fv5ZToe
jAL3JtkuYvgq5qSvRxBiCdxlVK2XtM9T4/NcxyuxOSqFI0XmCM90DIizgh1CkyecuCUKHDKlUiaY
BtQDw8U/V2SPIIDql6i+5QSiuufjDChcpduf2RRDTSUQldFZdr471kWs/ZR1x2lhJwMM+uIYb6+F
vY4L5CC8HjLmTmcWWZOOOCFrItHNh9lUD6hK+h2GDF9WSR2qiCxndIgbBI/SZsVyY0HWUqaQ9W6O
tKsaVCV7J4EEKLqKeSlkOTOhM9bvCkL2qBH/FG82EQ07Vd6Pqv3KCiPuDlcuVb65ilr7DsPXHbg9
SJvjgos62fV+Ke9vSlWrDaF2VtfiGxkbaqnAjbZedwEmAlzud+s4DD5R++Q1e+jPoBe5q7dxq0Qu
AUNCc6I4Xnd4o7ADUy5Yic/JNi83TPFhHUKmSlbBJZGht2sbE923B3OFCnscSeo+f8YEKdBMjfdG
qWzE8tAg2NYN6CADB+Se+4h502TQHse0s/COeCGHH2eD2xVREXc3Za2RrZpC/KHqfRhmrtRH+K01
fHQnsnfmAE082rb3q4JpHyTuh7PHBkR9xpkklHmlNwiiv8uSGquVzxea7AvFJE8sO1kHqDvwubuJ
ymb2VItT/vRkhZ46o6vwhDA8NFHZHii/bCkImdsWUa65f0dYzGR00ezCeznbJ0A+Ia+zccAgp8+r
5IwnS37kVew79HnRBcOQzv2EsclllR87+tCMkkPCHn+LvKZMCy6QbzJJKlxL6tDi8Gzl6s0ANq/2
CLg0u+lIyWKgDU/GPHtnbMnZ+3QFXAVyP90ArppcQ7HJz0/R8Fe4pkpNOlVh3c2Y1zQWDPCtrwlq
Zl5fbjaQARPXCFh8Xt+K9v53pFQnDr7BmGp3zBSvVpAR3F3zGPFwRbh3MAsrY2gNJt+pmgEvlG/S
FgbcPOUAUH0xiYnPyz8pkCIKXeGsgLWEf6UAU9gl+wZsFZ4+6Gv0UzQ90KCE8cFtgHgm2rxsiBJX
2lKvaSnueg/1D9pARpl1NyKGaS05IjTBlGzv8gI99PtHDfoAQaRtb++a902DhEVaop0jZG7ibL6C
o2oXjbbQM+9Pc4VPYWearbpKa42r6gJeV9DUoxUN0/YkTkcxp4493PMfJTMZgizIysccN3jmWPQo
/eB0FtSU/vnSUFHBHXTNN6Osf6FIOA6f4yn+ZtyMCqUydJamop3YX9SY6Bx1o5JNO1NGZGiZ0Gwv
n6KN/Xjc4m+ChkicP2+nf65D3+GiXcF248e0hp362dM52W45E6y2eFdqC0TJFk2T4x57I83g+ZMP
QL4inhF8DzQgAAQKvjV8zn6GTB10OvNSewQd+mRSZcWWX+myWX9T2vNioEPcoq36ZpD9UgVsZySp
OH9Mgg4Rrxt30Mrpz3Dxl3qFKezWJLQFOJhFRdzxjkjcWTA39LgF32wlWzNbhIebmtGRTQU6yxv8
EVaVPUaiMzGvJbj6OyW04J8M5UOEITiUa61yCvNgOLJMq4Qzv0B1DxfRvAhmKicpFF730TI8mSYN
tQFYLLuYvi0BXnGMAno0iffyHFzGeX/tNeCTjp8zW7Fo8QYk3eSl6nBbSyziEXnMNwI6DH/Ak9/3
a9TD+zhgEHkvgYM205UwOzVaEsK93cjacxtfv+fc13ApE0Wwq5WSY8g8QKBQpTETZb+VtRDbjQ5r
6roXBzxpXWanMCsoBCz8RiQRYW/1T5EF5ySks06llsTGcO1ySUU7qu4LsVeFHV5lBl91WQO2JRtR
Kecr5NiW9i1SCQ1/f7LIFqNMeSulxYPGwAGcW2u+guyKfNLGWZVlw+aNVuB8YwhqD3W/NTqOUvqM
Wkr1VZEz6RCEiTBPECY/QsYVwCZwD3zUDk8kVEsQunJ9DKPSdhYMwGPi6WmkGudZGnQ4HYLRQHQJ
Yrl3btOaFfn6Jr9RoJE+M6rzQqk4RxOh5JfQq0ulN3aHgaeAxjilVK5Q+Sz6M53polPSX9oZZSWU
jxU+iARnTFuNayYtAyqOeE/6y4mBy17czMR03AKrIm+miZNhbeYARGvms/lCYe78+gHOae3MUdna
Er1QaTIL4jU806ayj2a6WMHsAI84AbD1cRgS4Ubr/pX/CGxwjdA2tkQKd5lUJAZIPVdhGjAvXeaq
VeEWetyQUu9AuAfiBFF7TpJlre2HmyysheghfeutaTv/UmYlpIBmeoXGN77uCOEEZE9/tCB7SCi7
9FN9jKB6SL6BVunVP6TkkxcECma9oUadiGBobYCpIfSSnfjEAdyc7OCqihZ4BnLABvouLZUfRjL7
wkMgrhhw/3UbLyoTPcJ8vvFT/FoFG8yqW9UBFNY0nWXtwijZim5bSgGKVGGCKamZ8XUTwrS2P7ZZ
HDM4n1t9wb7fuOMgVaQnyQufKLoXkmUsFedMq73gUl2dpuN4IT3zJcwLyB1zJpCEBuJwA9xYJ90V
eZJQ+fm7sdUdGTLJAlbsKpp2QfDOAMmSRhHG0l/iCxUnVUm8QE+/w0QUkKZ5wqLNed3unDVc9iPk
S9KdHXobavcfT+MLYpJ3HoRyEim7zSlNdxG2DFD8YAzKmTxFF6N9OM0zANTD75HH+QeYBwxKm6NQ
uZ9aiQTFvg+Pc20pnkKfdh32WQqxIKxCHwiKoxTi+wKADp2QsB+XUAw7tdA7/LrSExwiXv3vpmcV
HOAv3Ps4zOzSnUdfA2fVRmryupJMorpdtcV+BlApRaoEm6IOvzpRNoGfp9U25dTBb5viFSRyB9GZ
uaMOLJFeKa2f6Uy2QBJzmNopFKKy6WucO4NUaSWAXaZcepIZfRmLyhqmtwwijBHM6REPSNDcby+L
FwTk/O1CjBC9qUGiSdtenZ/S4mfTlaM8ZDXbRALXF7yiCoX/O2hLg7xxdFRHO66OmpackmH6cUeN
g+pvMJymMN/TsaqhDqDtbqAa91vd1wdHuEZGbhIgAWOcVFkIrpjsC22UORyHXprBBX+dPnMI++rv
TZazJCfRAMZWPfnaqCfNcy5ab/bXQ4WxC2rnjyMWy7DuwIw9Qzyc46hm2GOIGjnmriTNKacmwknX
n3dlI/MfWkECRfCSxrQGOth7l0+3WRByMLNyr7+Eqp9y4rf0Z0tlXd7vGzLdWKL2tExuhVYKIoUS
yeR5FywUQlf7Q03v306Z5BS5lczsHmp8QLpHQkr8I5UTU7UW5s3G2X2UKNieO382xNjShEftmbii
O8105uZeumb95rYBWZAkteyKh5iiQvQvrxkwHWmFvRUcp0ykb+V+K2iH0MWWqA7hoFBYM9e6ySJi
YJbNNZas5/ilxwur0uOBODZaRaSbGDtcMtdboEBTUD1aqKITrbKFAmH02zNVXCWooeDBhqWsNs7p
8vmPbBiWPpUu6ngSTqVL2SyN7Qh4uz4l8xX9LjoXoJC5RDiN/1/krwdQWpgdwcWqep6L1j4sEjvU
rni89cOmlaf605MjR+IDvg4srQHGdQKGDhenG2UIh3kyWng4Po4G3Fje8B1batWBrb/a0ctNhC1V
+lYBg0rY30a9jyswnlU2Mfvbv5659f7e5ENYYmrWgQZGlrPBxeXW0f9bmQLxneHudbGQ04hMCuGH
uMjyGLW9LwuagMpQijwATOWegq67pBX9ZxDlmyaX6DQarD4ABkJpaM3L7PbsmLk/RkocdVB4acsk
hfagvopzbf9RSFRAXNpsDLLV9ik2jhI6rHmn2+SL61eL/BELaioXWBWNEsGTpF/K63spRQ32G5GK
0LZQ6NEgP+0JurfKS7pTe3cGe4kLrc1TXNILk36cyIVXVFRPp9Bz5fSil/7FBCgkmh1U0gW1sEz3
3Lo2W00KmRzPFBcd1rs9irKa3w+QHkiuBKhLox1VfuHeY178HmZdoA4wx0IL5+xULgwstaoMb/mL
xf+t0UEXChHUsQX6LH0J9N1KoaMr/bAgR83ayUNY8hu1h7vb+8hqTGzN24T0rJhyLFx+y1uoAlfp
yuL2h8ns1ERsgy+9o8ZBBygvbry1JzugIN3yYH0Jh1Cbbll9OuQY4cveU17ueTKKT+RVUZXdjqQ+
htnwXhl1ty1iuHAmd5HWfsjlFLgqQhjRJAu+815yh+olnuBAyG+WT9edxyaVWODqIPW4n4oGO2ac
qst4TSbZG1JNitff664gsqFlrwTFvK5hWSQ4htc9qY9X0jxDzk2MwKR0WEJucyaLvcZfjpoMopHG
8yfvNJsR/UacHhZiI4Xg/Mj0E4s008ZbwyTUpNBP01Y7S1pN5+IxvBKANqKiicrMQ/YNoOtiwKGh
KrVLPkUHiQlSyXv7R2LqBNe0po/U5+2h6uur8GmR+sYsOsA7JLe3nR9yjU2Z8JWhxduDqWM9ixPX
XOF0C4bv0KbSfCO1vzjX8adbd6mwqMC2GUsEves4sZQAgJLe3xc8FniELp8eRmzakqcDKBW658uX
FqSvcxwG3q1F4Jrxg9MM3q+5vK+LUFrvvKEx70grwc8gaVPRamZTb9+JZ48toYYtABg5KqIn31eh
8S7OFaFgWugYEU/Ep5h7a4JyYi5Lt7ANN6aWELQUpMV+FJHCQm10+Xmw3+P+sgXphdYI3lKXQ1y8
k76US4TUx8Wm8bXQgC2h8xqmW8y6akyN7rvge1vHjwxXSa928xLtjPwiS9W/Ccz2fvkyWPaUg5sB
bv4iomS+VQOAO0ZrvLtmHSAPyuBwWtE2aULEaPfoW5OpeBza5pu/yBW/oTNDZyVclBXxX4HccQSE
5QSsmeJVvUDu+iP+hMkPGBwdsCsIHiLSZ78PokGDRUBqcNuydP7k4nqtmleteZIy+Y7AwJ/4qX7W
2Q77EtmJ9hv5locHVZX9XtJnKqy1LIohGlDWZbzrMJtHQTYErJT8GX7ZRMSTMactZYXGdVToBppB
vteSXgdSUvxA8w72zB8Urp/uSbfFSwoO0RMwSnCxuD3lXPtH/oH6dXTfuMbzEhau7QqIpSjYTS7J
TOTl83bswi14m1J3epbi1Ct1LMg0tmVeVrKK1oTTroWTDWUFMxSDGCpRh9rtzof9wm6HTIrNqIph
Jm/BDzVhm9sYi1t4f1Si+P6QE73a3NXLhgwn0trrcboL4tHrx/HBNnrJ/AZuIAFwMxhB8V0iXTc8
Sm4QtYznr/pzJ6xL5JVHeek4bqCcNF7igT5mhdjhQqdcGat/hDBO9NMdEcrYQJz4bg7PzXsub0hK
uZ7K92b9wTZi6mN7Nw/IWW+ivBi8+aUmxY1YN7Nbj9UxQVmeZKRHi8os4IopsB+gDHilDPS9mpZ5
vfPViL5KY/4NciLAFqNLSVUJPScQgr4VEgIhZAp+aFNrjHxpGjvdcxovpI1uEXKiXQX8bYEX3BV6
i3dHJEbC2nfRZ88zV2miUaylNPBDdiawNKsgMJ/o53HAKD24ALTSLSSldnQMwoXbJpHyd2fjjbIn
sEaPs24Pv6clt+tNpqoNw2vdsg0k2dixbf3R2eEllPRWThYstaQ7j/bhsM4Zp7isQlihVVQGSRFd
F3I99BH+DM9qhEuHNv/ivAlUSbaZhPkbrdiMS1Y8eYnVVHIKjEwP4Ts4CGg8vROVyL/AQF/cYNPR
ImzLTLB5O1ubWEsLrBXntUAL2v8Wc9atabL/NlC13jxk7bbJIkUml+8K1y0ARjHURoDvrDtzh149
I/7GxsFAfWmxeLo7yEZGX32bHqOWQZdjXiA/heDm9FF4+lPO+5AF/SYAr7avAMbSs4GOAEglxOLr
E+Vqj1gWmcgMyklFD8mLNhJViEj0VB0uHo/Ehjk73dobK0dllo2LlgXyDkeNJMJFKEWwnbfcJ4h8
ppz+JuX0jysLOgVDKA8oigRAJKGGxpjiVoxhwezo4vVHcYvz1I1BDwIPy/xY+es1zWcEjYrz9lVq
cqACYS3WXXmSAw1br/4C6iYLxJBWJ6iKbXDsABrCTXqo8PFLw7Fqbk20a9Ai9bNr3JFWeAeSX5KB
2qskE+YjXHLDGapYecdjS2NomfI6KHn2hTxeEBnZTLEIF6MVMMuj+5KOLGkPgk2QecjUnTKfF4kU
pX8fFXL/wv5XpDqa9Pltmq9zUup3Y5jvK2UtJ55nQtkmYlTETgx9YRqapgAh//COaMCJCjZ9ao6f
YrmV/rmDjtdIG+qJec9MXGbzrajdwNwrgFPZ+xoSTMbWXSo8h9DX8+2hAZdAPMUtiYr+Devi5jrf
ZHGFDOhYIhemx3HhjHEDC82nM/L4z0+XDxgdAnzqjDlQgbVuNzvkoR5ldcqYKs9trlwuBl5YkIvE
eI7hUMVhEzOTkZMBcfqLs3nqqVimexVebtnvcF+MMcjeFpR5O3BuvwQ5HNCkL13ISbwOQq1wcONW
E8YW24X90E+oKhB6LcQDr204WP6SiFfbbcdHMktcKnharjpRH7kJvhQ9PXmXDCdIaNAK0x5hYYm1
IzWw7SJATAGE+JHb3KmVO1uwcQ7aHGqhDufDOknxtSOQHPTlKPC6cw+/pQs5v2/rw2AvXXacVnyk
IuVzuR9m34/tX9YQ9wyGl+gP9Uj5YKCdIdpybniItSnLgFigMyreNAJaZ4agKwP1a4/qffEVBmif
LDsuEciVMKkqPO00efg4gixjvL6nGKOSi8OnUWpWeD4ykQem2qZ8yHrkTygHyjaXJkh7zu8NaF0D
dD8jeIQSZ/+5ZYLUf6Wsbjtr2D8tWtFWo2ip082/E6VjXTACGM/M/hOzDtFp2mSi/qC5CHxhwjUB
oYEae0908V3FuZnGaot2Z0KMrTj8vMSFOuxO6/NcCXh8GKYW5FHWsGFu0BZUgN2h0PnKsCPhMkxO
1bR43LsJ+k6QzQNha7YQr8qc8Mgwb7e3q2Stg0ixslAdPEgkqwUcyFoXBS/bSuXjLkQ0hfkml9Td
PmD2r2cqvhWD/NoZEt+4ieHZbWYRx2EaWeFWCRLWZkiZl27DglPSpJEXk9RK7/VrNR//vAw8wh9C
N2ZCFWHueNzW7L1qyV1Xbt8yEZoOuZvwSViFNs6TDKdfpawUsYN129a9j+v4utdsxbggl+hoSz8a
Nng8pdOiVpaA7HO16Ql2uz8R2lE8XgGZ2VZxXasp6NKMPcKKyrbtU8XzdPcFSmpL3MQYZ6wnUCh5
1v64iJlW8frP5WU/fX+33/waUFaVgPZRZiI5AIY7IUhAvnxDFqvkuSOd3I6TjbTpmzcb/Ot65F85
aCZHjuWD21eERIto1amkw3ZK5MJcVp4oDxxpkbdW5JN3J6qKG0jJqYgFKj6w5pya0JfJDlD0Y28q
UdyoPtF6Cex169uMSldxa2+CCguIgAbjQ0BrjQRoxaV3xIMRIQjaw+bj2TKmhJznga+pjWjookut
r8qWVp3i6g1biYPhWpkFDSboEjHmSgtvhYo9ck/ZTBSCJu+jgvFbIwz6sY7AH1+v9RdtwqJNDdVx
vuT6gRO5on71+r5bylnpSmG2k6EQWULgXdGoqEIKANGoLF7MJ4gHMDHoECJd1mI2Hmeo3BoSFugm
6UFFq3fXBJ3NoAw113lOjN+qIXLMS55HKIOJVRxIGSw8sNce0lMyBS+XTo3NOJYgYsjHuYtoTsk4
JRpDInIbIf3OfNtVmaxw4m1BWdZFuA1n4UdNpK7J9yRsYn0LBNwdHmjwRznP/RU5ntA3cH5j5hBr
d+UAYA1xoo847S5WnknhdG71RQb+jTdY0Ev79x/J716u4KYcPk1ml0BWe24+hGjOZGM8pixUTtIC
5YaQX9mw7fk1vOYMhg9aaV0iXfHhoKuhJDKHlMePnRajJtUaiuC47ejillt85FGELdXdDRSd1ita
715JvDGd/NTlrMNmDfQPzSSEjfO18T6esFmdSL6hCbTcFT3mLg9TZuQ7lF+2g9KKhW/Uijj6l4c3
y0gjn58rpebrHeNAYgmnB7kLcPAg100gQj70hNWxCZZO9B8osmz7h7p14tB9GLKsb5KxgChMc6YS
YisKvLrO+IZfNbs+LhQ25l381l4XVhTJHokizGLftY4Nfcpbou0wXht+MGIe2Qo7EcTSO54DclUI
VJlVVD8dhaAM/4fWp5wOVTgksALyhpVxF4LXOIknwMZdjSd7vpkPKu0Dcp98LQXc4J/x7FDyn3if
+y7nlMvoYgTNX1SLDM7GC0AlcvWTNll4TaScfgAvzRCzkePbS5gSbVp7bBtNAjCKfz0N0XXI9ykW
8o994a0p/0f+mT3EWSAx9iNPRoLNQatcKioNjPH9i+DD7UrMH52hYm3hy7PF1qLJqBOSG5rVWV+S
ns0LrxJU9HigSY0uAnv7/WHN/5kIWlIgw5279uUows87i3DT+df3Qeuq/QMCKTC9lzUKJnRJTjHz
A8fuUqhsKPzaCgsz7SL6bIMbS1uvau3n5TOrqxcOtFnz11f+WtaBF65J0/BbhkSdd4Pos/IuwF0b
1Q5COR4VEPGJxPcxAuYG+CpJiEpuNVdkdxNiscFx70qsD7HMVUeOo8lXIuokIQWFWzgq7P80KXW1
w15jff9n/LT+I3LsGwHrTSBYo48CDKgVSFlE6hilcW+t2EGlmNQKGVrnSsw0NCbL5fNFWRKYLnmU
15m7HvYe59FATP1O54TvuHkPI3HRK7l0CuwwX4PPE8s46q/ePcrkw3/6YQS7ikCQY2EVP1u8PIdJ
kv21V6wJ8cuz1cfyPyW5WAuA5SmYhWHwgblD+hCyjYJ5edVlLnbQ9wFL0U7NexKaNNoGPm3lPEsL
dqXJMueOvXrVmLgzm4dso8VGTJYajHHHfziPrWKaFr9wqCThc2sPpONdJQMsmHspvYtuNRUrSrJN
SAe9zQtRpQPm+vhz04qugbMIYhzsYvHYUmW83ilRVPQntIG4Z96GUg5efv7l49qZhk2b0FTBaMcM
3f1m6msqBX0r70iy3Tq/qiMjJjNQmaeXitdcfQyPhHzoaNxtzzhS/MMJy9Q/O1d9PrgqXtEsxKHP
GuhFP8ZGJmqfD95lbOlH40gjKUqaPfTl0Xl4iG1QbtlWu8H+sThKGGH8Gxl9sLZ678gdCPOaHjhN
PygyMd6Yw5ouH1rRXT7aChoM/GIyZReo7jUQHaQyI9BxqM5KOMy3J1Uh93ez6PdCLG8O7GZY6wtI
2sWsXsk01aeUNtH3Y43JLdUzV9AnXsYJ+f6E2hONx46RDGrTrYIh3Z88If5AXentaLxNxBDwEyFX
vUbs3kOpjIkC/5LmIqckInv3JCyKuBfMoJGgxgZH0HLLO77wnG/YsU+JW7p1xSs7J1YFvNN5/iKB
W/V7+Y0rAfWBpenTHGk3Xl3gNzALrU4sW+l9Cpd7Gnbq1b0+JToUGEhBYNN7RohWyZiIEcjKs5Hf
KbShs8Xopbi4b4o20G6ir6exagtC6z6PU2yJXBG1BJFlmbu6M/hkcVgxDnY5Qi+/ML5n+5oXptbR
nslwPsFNse82jtNVAw+kdIQdGrG/4haYbZseicDCBsik5YUqmjefeLEsDRf2WDtCOFAJFd1rhBFV
Sdltjh058BgKpObPc9KLnmcWjfnGvVIWkMyLz9utgqPoaoQt41GqLoUXcj/dBYwwvG+mAbnebeLQ
d+60hs2kfjKk+JoS1JhBKB3FJ5R4u9hsedBTeL7NrOkB/TMWqokIIGBX3uzpsyf+DC4qniO+xPfg
M74mQfsjBddp1BnWwqKkvs9MFEapCxyEyQItIVvWuHB6YHoGjDo1WqMRfCXkIiZHSLqWF+E6uHkY
NdmJxGDiBzD6Z6+hchN2vXgGyhAx8anhtpBZVJ57Q57jgkv17GBitZ6QW5MEDIUnOLid5LOsvf9E
Obl/U3jaXLbsSiaDKVk4MozPkwU0bhZCvHwY+e5nelEiVF9jujqdYAzA9cz6twgDk3KwxXbBy1hc
vs0L4XPO5jNBq4sejRQrM0yY/hiyRoCplGtQPsNJ1hNrpt+z9RDqOOY4dswVXURBtsSp8Ssj/Jx5
RruRbdsZB5UQfaDXcRzixKdOeQLRmFDaukIB+z2DN85PMaH1rpMUOwovsK2A2bAQQKJu8qHOZ8Q7
lZ2MUz/qFz1KDBNiLxo2EnMbK14XcHDZtTEZs1xP6cH7EL0/QghE6PwCgwxuC7lxX2vw0/uWeiEt
Wqf+jsZ25op+aRgWK/2SeNl8erXcMpGtBufpvv3jpenWOmQxMOleKPbWQFxvzJHNw6pUFaGfBwCy
toCxpc3lKGNvDQg9xIATezr9SKkHC7cJGO066UVy3O9NGTJNxFGFJkmtm/GbNM5b9fKAjrud3FZD
fRfHKhaEFy4prjksN4E279EFkovV2qJ4+yIaNQB/IjiaM8eUfy8XQVZeB4lEIw+B3sqMO0/UCWbQ
uISrLG1DKqSBIifRZBh7DgNgDQGrLffuV4FFng4T0ZsRJB8Sw33wRtLSefp6wo+Q3vBbkUeU2F2O
F97CB8oKIiRvU80Ta/fjEXw5BTVXwIKridcMv7GOtr3Z87hVh9pzuOm+xmmpxsWggmEIg6FPNIn0
ozW01hQuOs5/OhYcw1DiRRFuvmWTgX/nBfz4XB3WFoprhVi4McdRvs0lHelI1Z/G7tdRyD8IZVki
R5vO6Ixxzp2jErIl202cZgrCebaat2DDpA56wgf+m4ukEsktSvILzNiwxuN2uvvzG+FaccGTjymz
ZD3nASP4zUnp+ErUapT0fu2MFBRUOZ8bRZJEZHGrXwXn0/m8Seb+wFirkVu8v2x8+kqqH02q8z+K
9AktvgeLsX4Tc8JjKOlDW7te+nSb8IguHmY6aYqV2UsHs0EbhQX3i+nh8SrH++w0PAu2STG3DGbi
72LuETth3WvRg2sdhHf7OSJgkIyPGdRVeZENzX+u89RnDk0LQInGHrJ7BGdCVZpWZGc+mGr3cgHr
q675TNNEOJfIk+0e3AtR7d3fLMGUrSyOLvdvCNxsEgidKZkHfs4a16pQ9cW02Yt6cKt477zwMrmp
2VBjcdWfZLGNo/DSmGO1LxOf0AgOCCwRTW4+9ShmMsi3YVzLZNiGCiNPDIQi1eZ7hDeaaOMdYBFC
kfau1vbgrYhMjg4MA0dLw107+XtUDRzK+B5Jv/LRxc4Og4Squ/4BUKrz91S5Fh7TTZc5TSxisC6N
0exS0qwZN2xZqKpfh87Y4iBZ7ZFRFRYYIVtSvfUWgzeJIxzthRaOcLOAYMjDC/MdTtTf/YxilLiK
8Ku2AJ0JPtVyiMnjgcjYrfVAfZAqK2DX/B74VEbHbZ1Zqk0x0UmlUcTFjjyrncbb0bWvkURVHP7U
oUl196lonmlSuiZOD5d1cHhA5XWSw1kJx6fMDXTGRMPGZOLPPkHfYNbXsJEbQmJ1A+4eZANnstHk
/jChHxdLzzLzMMlPmAUOgUf+0Q8Agh0kQvb3TxnhsUvWaDntIeUBFme/9l/km7EeGRUdBJSu/AYo
LTP+44PujyHAIu/9YzHWhxGT/cFcZAzYa6C9go9qcNkTVgwJr663sKv35CJEhDBUIafvgHmlBDux
uS1Kj4e4c55vAGH0sGJ812FxcFXpoKwSj7GsBFIZqiyzhPboP+94SKMopWvmG9xrM6w0m6aySV5U
mo9szJjRpqoDyUUbQiUAs+cS9o2bLUkg/v0n8hSyAYLuhw5iYmpmUtUZOPgwpNyCG4pXnsDAD7te
V0lVCLagTHP610TcrsTVPwc3z5thDGSefQaqUzxNBDVCxHdDbDg0prI/1isZNXLdNOq3kDXZYajU
8t/j3mHhm/nmxRi2WS93O1wxRhObGx4pdYyVREicK6bPDVEufevEx5qMoleCzD2Hm1mkBGsaM3vA
zsr0ipB2QJAPOnSFth0KuDHErivrDqRUa5axgNRIxXl/rjbxTF8MKLPzdTSli2wGy8cQerH4WlSI
9SrrvJ/XR/AK7AbnDh9SO+3jaqlvwTL2FP/Dj3Egi2p9vIfz98xvJlIY8CSEOqwl/5xhjXik19v2
TQWrhXeRAwCavxU+jujxLhIPkBol8F5jt9jZL4G9wid32dMMUG4lY45o7EN9ssILDe8bkTPNWgsq
ZEYnUHn3vidmY+R18s+42z9o1aDCxWzZjkwfZcEi14pXTMP0sjy/gCoLKO252W/vKavgXxYXGZSL
0GbklCYmIfDL4Mm/g/jsmtTPrZxPaqCoMm/6i8wcA3r6MaWDjOnjIJYN1orcJyov5pV2lx3UEam/
B+BAFEdir9+FbLlb8L8axG4Qqm0L3SQaSOFuR/ugMJNkwoWR6MhU0KoXySkatdr6jmpimj3M5X+x
QRQ7hXhl7IW6R7i4x2ygpLTyM8psXFkRaKsMUPxZcfxXgP5PTOFS0XUs3HfrTgHb2HVs72JMtZxA
uaGE+xW0h8xW4fMmGQlLuxhGH6Pd8oDPganmnGnD6yC+C6sk8NWJTyrwgbCcjzLZKCiWjQxQ3lD1
e1+DANb6uS6R8nziw1uiaaFn+0Z/VbNxgl/P8hELxbJvenbG+0MxatuNHoABZ1GYo2SdfRlfsY6k
kCH4shAhWsgxyYMcB7FqOAM0vt3yviQMtG8ktgqbiHL1phByfnMov6/S4BUQyyvG250o97GTuM91
x4SdWGtlUj+2J5rWrm1g7AY+IH1QInTQx0+7bFBnwjIA/UKXWM6VpMZfzvMuGPP36n2MHDSGCwRp
KRA634njfFR1akqMpftWZKdtuA0hcIG34EO4UORbGGbwJOt6+OWavQ2X+NjgYydJXJPOg/KNneL0
DmUHspEu4QLRhwZseUuoj0amiKh7SMvO2pwk8tp/qfihdIdC6HB1+iLxLraby8UeJ6nkwGNfZiHa
vHFW9oufj+usQ1TtgauLAMtwbxrleJHqVH15EnRN5OVWa7MxWd+Mtznbh+v8v3aTDExPGtn0EFjn
xceO91PK95xz46i4vX2QsKqdQTZnezHnNlVt1HCKQhacZpJsrzZ7QnjUTZxK4CRTJHlbj3uJUV6c
ahRoq6LAFgutCrUy66V9P9vjgzCqvTEGgShayAgfylLX7obZ15mIOVmBJBsHdTSe5BxXUeI3pzx5
2xx3J53Q0IhkX2umwm+D10kznfQ5ZbahS+NbmhmiqZOnfRV4hs4wxSwvoOG9pEIVypDWGJhH5t57
DYhwjK1O6T3arp1lURn6jSke0VbgD2PeGpudm4PWYk0MzfjhFlbts04aUrvghp7CwchOOPgNJpcW
v4ynUybDT4Mm1i7TVejfzm2nCIa9FQDlU6V39eEC1qb0AqSFA+tdOwsPx4MIiUAGyJ1sCr6RhDZu
wSm6LLPnWzgdvevKyz6o1zPyeIMRFQ7Re6mWW1gWB2lhzl6JdJgrg7y7UZlXrVddu0YuO91ktw7d
beDhurvSAUDKxJekXOKPsONaSmKmMSp4XsTpNZFb60aRHr4klRhgFzQQPtIhTReK//1GyoFGfTVX
fyebngV4Mar8Imh4HRcvNBkKfehm3ccv7VsIUoxpqrhwalpSzIrXuK19kxj30dHa4dB5/Gqs1kGk
vvWP+1BlHc3oHQIQ9vCAhIe5ioiJnHE63Vklc3v9w6dgqgVNaA2/rm1ah4oSDL2vfaErlmtIlHpb
G8WkdWft0KIAYjRxf8zHTPAyUPKoCRehDMWpbLPoiPfPUPwrxvGO852mtcCMekkzAgWy3FmBWcMZ
bQAqCazzBwow9db5yDgAU2xw73C6OuMxMlviL2OSWEa7ZSdpy2TnSnsixvK5npSedvwmDsIqKxar
3YvOcylRbRa4pUuCXKUIo81AFLWLK0IMxmdPmKcNB6MwZezhiB2u4nKwcqWYcH78g05CprH5tQmR
LSIloRAv3XoV8KloQq0asYYBGNRc5tPpJ/xNWeqTf6bMScH/w9DS5XWKJLbM2b6ct8Z1gCIv2uq5
p7qzbfAKBHqoZBcMAMZuqUjfLZLdc+44CLzXRDsZHLegOb5+Y2nKAdMmmjIdWIhGqZkkM2EYmIxO
eN/yfGbUQwQEqZLGsfXEaNPWkNQh215SJF+ZMKgblzJ1/N3mfREbu2J7wAvSuRUD+8wwCj0QxFCI
uXAf4PcISvdln8TmmjXL6Fmzwt2GFGRXFOXj3dDZO0BEqLb2Olzajy0MOa4rHkOozE3K9QU6PZfM
bRE8LmEBGty7+QyL/mKvQxtwWcslFePvMWb8DBWzKk7uT39eKl7yIPZ88QAPEuTWXFgUia2Vq6Gf
R66HC2LjkgbDssIpqj2VWHj04FkNOUap+TBqzeePyxHsdYhx2Am10xg45aS2loTBFKQeSORUxnMN
XeHMP8Ixv3RBEhUHX3SfUNEfXqwkR5Q3GqTYaTw9bfpn5gSwZxfWy9pQ10k0p+7n6E7gDNecpgXm
t5MRDYjmbRsDlGfAH3KPSHsPq4hOPx8SSAJwn8OWGV7c45riTehJtmj2Bh24PYcl0Z0A3WHukhr0
c7ot/aRSFno49/GiNpgNgYVDX9U2dny5n87GR9qoRMOjs8o2P5lB9VFo/CtHOrsDew6ssLnYmNpP
drTQRdnKC2YBhD/lKY52e07wfNaceEnT4uyUskAXQ9MQIqHCtzyRT5ZOTpuDSxr6n2b2W9i5FMzv
6Xq4QwRQ1r8AFa8XKq7QoP6UtUQpl/g60c+KeZfu9eDBo2euHNWRREouSSubeOMQm3A/UzdqS5Sk
G/Ph3iXog2wnG9tSdq78Deg5zww9Qbz5BQMZPydzuiCU/sW59gTt2KPYojnnoZ4rvRGFrqo+TnDk
OduVecH3UOxBIFMFH/Eu7uvhMR5FY17jEuDH/gUvrNdP79TX3gFsO+l0t9bFVGRvd1OTeufPH2zi
jXPGLUchHxGso28ZIEAWKM9vMI8eV9BmTOjts2UFfX4DbJURk2777x//hY3g/qRcxmCTLzWmLCzx
AVB3ePQn4amLMmsZlQDfEWoRdU3HbXWn1HKkP0SaX94BRCXnz+Iu3fn+dbSbFV+Molevg8qRgRT9
xNP/lFDURgw+st/A5lh8cIjHgYKilQYLyPZqTPu68yaZPbrfKa/ym5szB2J2HaKf1dR81vlVzU3D
zMzRDxfYwrMJTswSkdh8QedZVEPJ01/HHJ/WRgJniTw+MbVXaDZS8FyQ7vO+BE9qMVCnzTx8JYPf
QY49jkbgj826rmnkyWy+yGT/cVARHTk9hnDeYHVqFpAElNZXqmHb5XqY32HJEUNl3smWzxcPEp3l
iTo6AMmz4Q/UqochjEE932MUK2WcSNnALtjkc6wWYmMucqNlWjANcuR0y0cEE0UKHM9cMES+Pzyv
gfeY6HVbVWqjr3jQnXupOYCb4TaEsfylNCFYQwYjsdahvnHV6PM+R4xieUnKvPTcSY7bhTriQsFI
gTXgAzY7b443XnqukMSCUjJwMlgyYfllx/g4qQKXEDJm12ozLes2COifqZuUycvFJpI0lt2BFWqc
TaoVdHY/3sCUGnjGV7qA5VoeOI3ipr+2QVqSluKZeCD9zR+FSsjq7FbRhgERxiDQypuD0x46qzsR
579fIqGDurRRJ0SZ5RtUf0SzfZnYTptGisyMA+ISCUuK/g/WEFHabiTV37+xsoaK60BsHT4VgO6X
GQNA8UFvyATjCxUW36zCwRDA7E1YvdyoGScCppXI3QN12MXXb8fbUuFJ2c9ZSCnNvYHBlT/Zr/yT
3FweJdh1sAIcEgxiI54kiQdQKis87ly2PPIWogiOa/0Zkmzt35eA6EibOQeyXloNHlRB1weVLA6u
9vdgdP9fPNUldA1adkTnkuveQJo+hjc+f71CIa9topNlzC/BrXkoRU3uIHcPVOA2hqH96NOX6ReI
yDoqFKQ3bJi7IB8rSDDygJRih8vSqGG3KAMe1vDaTXzLMABjYhpJFeVNPEl4RxPEj6bgbhWqniXp
tfPUzlyYq9tVmTjPw/Irw1B1UEOUG2KAYVSqCGyFRVro1QnmUL9cMapyjLDRDJFOrwxXt2iGfHpV
Bci/TE3Id2OI0Cjbz9QyJFQCSJj42zj8ZQhEsCBrLm35QA4FSgcIUyW8hBgJBt3pISIXnvucG3MW
kNuVMR3yTJPeg2ZD357ueMbNBnjqczSbcSoOfGKOcH7LtvvMGPTYeR+YyXYGWgJLe9wy+3s61CqG
PkJ20MQq9gixwggCQnfRY56I675V/h1pWTd0dnex7FqHVPzXtYR/wx6/pIp3axKx+p/CYsWwFAOl
RhDz+wdHASUXvqrj4MPBR34LnASYWKX7huewiOQXRuUpeg6/JueVIuWyspNIdn03T+nelsFgosPm
MXeaxgokOwTxY0S5c6LrusMqwbV7ss8/ZYTKmZmQMPvw0gxHeEdGBHkcDnysRpv0ZCEqTv11AP/X
Ezek3Aw1gMb7dwe0OHhIcpMVTLbffts6kPwKzoNSMdgw4Jl/PS47qPwahj8qEpxQtCcLDhcO1TKO
KIROWXIwmlHgmyx1e+PMpkFv6FSvkn2bRfD7r/XUjeOuysntw+VtKverO9R6vt0TCb6NfLOBumcE
gfOUKItk2XTf3l5UzkdXs6Q1XL3ZucWuYRSWONwmtMy3cl0Zq7jl+zEEAVjP/O7oL5rJ9eJPgY33
G1CDO80ebbeDfBOkbwK+g8gmFYXn6uXGhHTSweyocYf8LcI+0344WY3sHvxVCMMjJieCZoWAmv4c
NkwDtT3NmxihO+TjDMJgzfBRf6+1wYNECccx+09hiYX8y50sq1wjbdBHkRBG7flS5N1CHWi0w4xV
iwF/v4M67nIw/5jFk4iTOYFD87D/47S8cnGMpHmyPsPrqGbV3tLL586nwK1XQV/HcoFEXXLAzek6
O2s+91tDlKJNZpIEFdBJhrMVcJJkPlhOCIcjW7svTGBTPWR+9NKr5sSQDO9IIh88DjG5WIUgt7v/
k1BSdEeVyt3rb9CbEhsO2+g5827Q8Hdpuir30bYDvoF3yFpaux8wVduo4IR/z1xfsQSY0VcZEXfE
wKS7bDgD906s1dWsd+EqhVojv1J1NOG3EsP5vCcc8Z9kdKsN6OwzEy6vmBvia34nEYnzAn5k7ZoS
mk0EJIQ+4B4UlSSNFwfUrxyCQZzUTIL1u4w2LZ+zVrP+CPjG831bU227EFUnRcerxNf7/ME4WhAK
VDb6MS7VSRMoi7ry8v7UPVZocjbDGPoORN2Gj5UlzbvwEZJehsRYG/pQ9pjHJ14H89tyKqX4kV5S
xKV44M2xeaXmb0lcl4l5yS7st7nycHIO6gf9r+xXGu4wzik0IgR2YQ+zaLl0wX+kRWu5L6lxwjc6
x0CnbcnZ4DnZBMS2cpOyMlLUjK6N8TZ066dJZLOpDTBllgL5lxVxcQyQAhU8S1XuSuvwBOjVz5QN
5HmktFATpcG/VVZFyNdhVWZFlwgyZmLPW+YtHWFaCt8HD+BmstkDRkugsEXvmTx8eHxGFP51aqF8
MBmsMIeurKElM4b0Isq8ou5CAc5BwF3gTsI10gfzzDd8s4evE5ZqI9seXctaoJTqVh+z7Eq6jVuO
BDjhXXAwFJ9MmrnatLUJevQQvVIYK4HAEoo+K1xRmdLrTb0wHlXwoDD1BC+Cj64qNHi0pOfTZ0mm
NmrMrqvu0mazS55UL83lSSnmMunsYg0fhMkPa4zJVpuY8QUvOiCXQ+DW/g8emykUIRz4OxLd+/Tl
hb7XA8XOnbc/s1h7GgR9zYf44bTGjwKndxjYd+9lHf3ToZiamyuoXAE0/zZ8CRAZuWLYoav/z2Vq
/VwYefbYCn2FGC8iTp4Bv4oxCr5b2LmCpu5TfPGGUbgR6LsQo/f5tzonkEBnMldtX3sEFCtcj93v
hRUNr4QtIsV79PLuCUoyZjzWsoKd3rH/GtpnkiEZg1uNmtJMP8g2cpNARGrQXC9MusnsIWdBDcwl
SG2whgguiLm1XvBbnb1li8skyXmQGLOUKhm/c/TfxtwHuGdzBhTBkGo1H6Pol5rdGvoRv02NQSp1
YH5F2/8DKGunUUQCcFBIj8oEdYmSHCnqDJwSSAvK7tTzr2APWUQXhwGQxTz6M8hnzeSj0Jz0u6q4
eS/p5svonOpL1f8DKbZ94WbPX4d/hNNxROw9N8kcUEew2E9rSMojohJ5eipnZbK6WqsLP3Y2MKS7
/wVVBSc1vyTkdNQGFscc3bx3CuJKWjUyLND9ZZMdY4Klj2MJXCd1Bbw4vb2DWk89D2ohyy/PfV4q
6vx/7gRcihO5xkOdNk7bvQXv00ysNOT/hCDzFz5sFRPbJWHII/W/C3c2eLUK2rhH7scP740vxvla
tbqgro75xlQl8EjDM47H04/ptyc4+EbK7o0XtFofubKl68HLiWla9hqKYPZe5T49aZ9lHpd+0ugK
WzUWtr8ypcU44402IPWpamT+OmnStSsaiqaSYtQ0RFxyj+ExgTzkZLTomqAiaux8klqZsvbb0NF9
w/QACTYcVcsLv8KzeAzm2rHTAmtXkvGVuzoRk8yOb0dAKLK7z0oWZogM9v6Idw1QYGGcvrVaoTxL
S1Y9bjPUhKnsp8NlKRvL24RmtA8q5gp3TxpuoqkMm/a08oD8OjpOxdWGJZY/sjlb2r5RbxYTxX4A
Zx6GjYsQLGAC4pgPNu11RnmCkwW8DqQGKkLJvCjZ531XpYiDVAgmje9ZY40/c8TiacY86wllB6Bm
ZkFcnFGQt+h4SFEHPoJYLrfG0tsjCwCrguPyzmEYkuGKLSlGa21n9HuFv4MHYPO5DRT9zmtIB4kp
rmylpTNqGGTDYuQPIWs77V4IJDrtB3eHWfw7JmxTJGKCcRC02la4IObyQ4rnu6Yrz2tNHn9RBhoV
Jrh/WKNC08ycSFpQqIKQUGNcXPrmH2sAwy8Ia4pvcxC4TgnnY1vBrDmTyu7loVU52Kjma7EVs+4o
oVdVNEbFNmWZ+lHj7d1bgRSXD+/js09RmpVDNzQr7OGJybTpBXV+CMuTij8nYM4AY1OkGsh8Jx33
fn39wcLVwub8jJys8tPeEjzi3/guZ/HjZk4xxTWNj9sYmXDP0wdO/ApZHQZucTlRm2OZHb/QszJH
GGIqY+LVDKywnVx8E8H6K4Sp282bFt8PkkzRk/4QjMQqF6CCUGAgfbTbjXoTFEYgb6m1hv/NS7r0
ZPdw6EjQjtAHrFvrdaZDS9dlxnz8866Z7OzbwtEDawGv2MEqKGGqdXmHCHz9eM23nRYi+rFRdXrD
IORTa7w2oVBkpME3gHt1r6CHjmTWILUCcIzJ80Pvgi0IPCetr7iHLqJuhSQrX/4ijucU1/7ZAsuP
+WrnPCFTQxBY/eXEJpNhmsikiA8VdHsH8VYc+BptxOs4UPAoUyVvmXc7SkJgXBm4kF+z/CEpsnXy
b3/7zCS6ILS9Q0DoCA/MB5pahg5EeMUSLF1qY89M0Y5jAu5ozr6vqXJm8haif1Pji2viYbJtKolQ
+w+9C3A/YqQCaDCnXiFBdp1Q0B7gBLRELMf2Kfse1EP1cXKM1ZdYoVTcUNUqlsDqEU1R6U+YJ7RR
xGbPxHMwyl3h6fWJng1yLJunoHKAu3yIn0dqQ3NmN3u7WpmR5229GMutkxTz3HXjmIVssJrmpLL5
NXBQ1ys2GCIIJZfPWQOg7UVBRE/O0d0dor2ZNVQ7m/Ny7br1smnkATu31mn6lEGYG5Z+fZgFy84Q
xrADTF3HbPBZzltvSGWLOAFA+C1OjkajZwgnouebTiFys96auy7Cfp+IjAEGR/k5EyS8QJYm7ZCv
0LNhqhkM6iVux3WnA2AY9ctm2G+gXoAsuALd/CRVGvX62mnsnusSWto8b/9VzRKakrsXvaKDB2XB
YDDjBbmituSoSSoPUhWeDl2iAmqzGHLqHBnrX0KQaHTIEvPgZcQ5S/6jSZkwNznPyHQt0uux+6dZ
TDYerhGz4jW3GqrStnhTTZRaKtb0TUKSwoA1q1eCBG0EMy2uoHVThPNFZmPXm9xC0sT35Gb+NM2g
vMVUCFxZ+fEU4eBn4pFRCa0tiVZgsV/aJ3MluMGqitHn1tPFqjYL+fzMhoSKZlbCB9vEE8ANfUnf
4TMAiyfIAcbrbYImnz2faSLx7Lj4Ltu0BtWbtL3ASCe3gU/NfHdgViP63+wMg5/LGILO5sysYJd4
waTYYSj9SoEhw5SQRyx7o3nY5EQZbBzwdB7/b6qRgiRunfaiuV6nkIWpIhjcdSCl9dDzmuttN7mr
YMatQQcFPPCx5Vh89GTsDDt0AzHbEXCnU9u8vqoXDBRmVhZptyOxg0Aa7BGnc9rm8gRgN69ClEpW
e35gH1aleT05lhtCLfdEU7/SHnOisHKHaF/a8jz6+Ih5NnpDUMVXXfD/7sf16p4iTnVJU6vuGaYB
m3svLtqES1cSTOUY14CZ6M+A2A4C300BxtnxO8QWL7ZwRwRJ11hs87hfgCavCMG5EmWws+n5fhYF
91OoOh8kYjIqz9Zgc/rtLfNCM/cNK6PDy1ct5CQnOEXZkvcf2vAZaKkG9NxceW1QS8rmUVoSz6pE
OTuLknbpxIiTQQBa1hPOTUe0KTJMufAUXkdRbXlqLa5KuUpqVoTDc39NmwJr1VEIv/WmtHKxW86m
ixtNn//deP2DUIWY81xfbe9BaWqwmNTsYvsssU/xuel0d8BYh8RuP1BzZLsubfK/MK1dagKxDWLd
/xHbIVUS6w5QFHhBtYlBe8TGpVlnGBS+KrQ0sZfGvbhVBlvfjH2NwLsLhYVRVT7eljgMA8uXJM7z
WewatcUvEY03uSXGATakKGNn9Fvr/2koQyRhsWvkZQp1cyM3Pgslp4MVUfh/939PRU9ncBmJpur9
6PU2PvpzzmXXtHYDBmjZbg9MNHpOpii0EwiX16cBUBShLsNPSlC6Bhpfs1WABrrB1RT4N6FtchWV
E6O/VLFzaCcVRQ3SsX3mqBuu5sJXM+O0AP6MbqDI4TjGYxGjU/VmW/ylQOZhQJUzyt9iqI/TGEjL
UVNu1cNr4O1W1DH0ryhzkB/bLAGZ2IW8g0OD+lTzb79rlV9HV4xc9HhlsdphHYzYgdhDSaJM753O
mG5TXT4bng0nVJtsGWVuDrPrbCvcqHmQgAzKoZLKc9HM0xXcszbwIw692bAJQWoW4Td5epAwj1pP
ptPY4oQrf8jmlnbbsy4nn0ulqxMMBTPqRST83HUKLOpQPDn7e+c+/dhWSfrnHdXq88yV8cG+WuI9
hu9k94rkk27FiFiXvd5wHMynqiqW8XeMoSL7TyB2gKdjyTDcwz1Adg5AVSxrGmeDG1IaEPqsXz2I
9SmzW/XcXgYqE390NFUBoMQ2ut49inCUgvQoblAMeN2VXtoFkawg6WxNEddz9TRu2PTRuidSokxf
UCs0ZT/4gL5g1mCCA54BIMjxccCS9fcv0gZruDx6QGs3C/R9Zu6sK+vPbOHe0A1haS+8KYD17oq2
vwgqtM14pkdIJ4XV4Kq/rx7Ryd+cFNqrSPDikDHgE4C29szFbIyyvkP/yOO7k9gMsY84NYjxWvmz
i50paHHEfCiZ4AZIHDU27TbY2V9LGYUDhF5kwssQQHs4aHzC5RJsPmSF3iEWJ5lgHilltfreMT9l
G+X+skBKgcYS9ghFn5krvcspnzG9pY3luXmTPdsZehcnHopGHscl01C91DCr9FlChFGUrulcDL5l
q3+4idhiJedMuKHLFJf9fVeqA0xxS5uO4rN6hB9Hy2o8y664fKuWenHdxgfoLvA4xGvz+VxslmKK
PVPX7FakSQ5uNePmsJ4f9pVTvXMNUxqdvlJvaU2Yb/YKiCS5uHq9jAzt/I+113hzSV3MIwcoYhGY
3Wpjj8aHsQDvTBheN5QvML7j7b0rQ2vwI9jqAzCKWwWeUo0VcbPSXfaypS1f3eqBdwhxdAnwFlbI
7SvbhjiX2kxEME4fNlcOcrGBIB2Osl8t2odfV9IO4BMvguAQ8EBTbfp0Ih9nEnIOgmvaEHwalNIz
Kv2fY+BD2Jq/L/RMDQJvnGZ8OTvPYYhZTPvO/P4QEkmXyFks26Wo1dRafQwI79omX4A0GYIOBrcA
O9xNG6yEbpmZKyInUlD3oxNmVLh2FK61hpdtisWlYTuM1iymaMnSRCGl9TgYJ68VDAENDO16Mz5G
fANyV4B/6Px1+gszuUvbLAzdAiEUDMyOhIdHGyDqwosnMO+eYuR2tq6q6TWewk7M7NhvGGyUv14+
hmd4maRmOGr8hM9yOYmHHTdJV33bCuY8WIpWkmF/vxAZiL05R/ayW1QP0kDEvRvCURwd9CIKVhZQ
HUZiZ+TdT0layAwJCBcwEA0c6kPJRldExyPNPk94Najw73aGxy2/BEeYRJTo+9DbV+jJo8rrexTK
8jumUmJTj0/heaqfhPZrsabRnCYyBH1Vfw92tZzpijtpyNS8DUj2FGSJfgZsVLN8AgxDzreGB7T6
UJjxmBJc6wgvQHJpFxakaWSXC5xw1zIJx+zIYzQr4xVI9v4/FCFo0eRXCSmAMW1NqckPs8fVOJ1E
yvtKhk3Me0mmeA5OHNvTgvyarCmmwFwd0FEpfRu8mzAXQjhAgltWOiJmc1Ej6ZWcxaYCHEq8brxS
QFizRGopS/c0TfovG6/PdMuHLaLfCvPP2qyDXs4h4jwP7/19OaA++TJQ/XN/mZJHLb0F/JYRtJit
KAI3WMs5rR4Z7oXlJdxfB2fdz/NqHeLQvWfK5K1sreUQnVN3uBHq0yo4dPbWZsnxnwyvqfbzAZhn
/cOWehV2LLuZya/n8ybjGg0//4kzHOMN6UxwO0u1hyOe3k1xtMxh2PUjnOl9AL70oLmkb4cIoApE
ofVMuuWJYtLxJWH6C9B/1cpu/TqqF4q7kSqH/nMguW3DgkiT9SJHnDV6aYP5ftOxCKeV3Dj0hNLa
KGkgrf5WjmF9neA97DAmid39z4PkWcdViXAPAnvuPnjO4Ax+AWN8WnfGWzIxfDgauAIT19oXg8r1
kaimbABPpx+80R7OMwAKCS/ztchDVsSOGYVwlCWK3C3/9NaGaSfAsbnjLQWUREH/YQXfnJyLffru
WIjfWsBs3jET26QtCx+fVgjb2/Q2kn2VW/14wqZBrlgD4QMUM+sUAReqlBEhG+SxHGrhLWCiFU/1
0ux+NI2iWD/QXcOextk7eubNFQHKDyG/0YA6ZfBfSEIqc4ik1ro9vIqwvQDGvMgLXyCCNKAw5ZFn
wESGYbLttDx7VFGPygf0sxHBVgDoBAPov+MqXXjUlKzMkU9X9nO1MfMb5+LNzfrDClZJFX6mVepX
v9J/n+0jGljC1kExZn/qw22nDM16q7kctNGIbRjG16lS9b74zJhkgClRoeC8fzWViCpQzdbdHKAt
Y8LtTK0LPuQ94QxsH8UN93V/U6ohYrgHE/vTGr7eq6LoTmBjOK2heNCWnM8G9Y+/oFjkcz1WFI/n
kzluStc9o8RD/a0UF1/+6XY0friVrf4ap0/psiieBknI21GiN94CytO3A6NI5tXikqUPLBjDRxrf
g7KHziF7SGwW5CdBelSPLdgWxNpr7VPqOXh+E+TL08DdgeqroHREUHWzjxCLMZ7NiZ1CZXKaWrcL
pCTFAcP1TI0GYJDmrtwa8RHvt3Xj5C1KS06KM3SB2NAlkhRgreP4yVxk/J0VgHX6DhBqUg3uNROF
TmhCTsgb7TVDJdwLd9YvO8wIrMY1y/h3w6nAvWNNPF7tszyQXFgNjlytqF2/GDR5TzgteZ2PChEF
fIfr0eUH7hUPXWgO+q9rbrqZIaWT5aT95pqogcopcdsiet4/YXCJEZDdYuQJnJZ1wGFtIy3xEDyN
xxaCmyY8zPn3TKUUGWh1QpzsggbHsRjUhbjCB/Jckr4HVz3ffU35k3eCrqEoO5pCR7zXxVwZt4Np
LCIxFBXE4b0P955p+qhcFEh7CJNP1ocsENiM18eNUc6Fsn4XsgXNTaHbbKRd8j09sVWYi6/zI9l/
IRvmDiCW0I83+XveRSWhbR+2NLvFFulG24iZ1Sajpg+5CAlMu7XLi0ZjioCj8eid25X3DatbWMCD
ZWCa3TzZxk9602mjciotMdYPbiMeCqChvrZ1ZhE1CfiqoaKYLvT+qgw+NaFg21RjnWg2cJbGWm1h
pKni3276uReL6gq4SMx5xtT8ckZJVtJqObiR2OFLOF47bbx+KNIVDuGSuGmhOIT3z02/INWDzE+V
Q/f9cufS9zd3LzVxhKb4Zs8MpnhCoOBYSXAL2LWdwyv4itsr3HCpsr12GJkqnB4sMS0H6zyIr1W+
PmmeK/Mh8UJjIxOLq7gfii0aTzwS7LOajvxGz2WZneFNHhLmy+Njg0gsmnxcxAew0ADapHv+jyMz
HyPplWfwANV7Hcw/EjQJ18OPl2cU5aEzvqOMgkYJKCYhNXBB5h/UVhvybgDZd5auJSjvBoDax5Bo
SjczYAOO00gcgn83HNnUgSenUIQOIh/Kz0F9X7qZiYZBcVfM5V0+uNG/EwkKIaKJWNZ8HVUAgUXO
SYlbPOLRQ2IH/jrvrG6qV7qbWxOupYrU/J9ab2AQYaSWn2al9nPxL+X/gnRdzwsKdniFEBykVaWi
3oNHQAuQ0p33GwKdc53P5oWeZL+ySl/HQhMXaH29LYf55avvczyyJQ0WOm1WNgMpXAAFONfTEF2I
8bVunGcqJJDg6EPZAM61D2A9XgS5LboSmo7fCe0GuaV8u+RREq9temM5ulBd+NElWRc2EDr9g3PT
nYIfUELm5yn1/JlZYdLqAr6CQ2OQedK92ePYojC3pJ60UFWQDjWwru32xtrP9CKlQi7KYtHHekF6
5K6+7pXOvMtXYeg4bakBupppM7c0xIQ652gqUqrNcLylXgXKabsSOCRlIk5A59/qihpw4NT2ebCP
VTl5ZW0C0dGqirWB7Y0W8U8elWZQWuJRPtSp+696N1AJ7RQ9kdA7SZUiGn1fcgus3Pwn59UGxGJt
1aHl6cHyEvJ6OJgYcAsGR7vAimUnXZk571D6xxtMmA+dUEwd5OwZMHXIQCDfrwsDUmnBHcOcd4bM
5RVH3BsDOq+j043cuvOMN99iy53TMW8H1a5CaGyvSBolbgMv1LhLSFXQcufCCpMJBxM0CVdtV9O8
QpruuIjA6Z4UxzHtQfMShQ7wy8C3IfOSOYaNFJzoY7fhM5PoSx2+6OoWwENB7hH9S0GPpA1nzgE/
UxI57duRAiX9+ui6+4xjIRMFKci+aqazqbGol1I+1o+q3QMHzlQ5VK5MLIqO7t8TaFJWFpPL6ra3
FSFLXhvxunrlKe2Kw4ywFQcecaSBVDcFyB3gMc4/58bl9BqVgEXraF+v/Ovz4WRdbWV7EtC70Xw8
fvO9JOsKzJUDJcZFLEY5+7uhYbSSCFH54e7ji8BAKIQPbeJGQgwtYvfHzYnXqPDXbRmDROTEKcPB
9DStmx5/i9OZGe+8Hpnl+VSOkJRvCDG7ZuoQzqvp4PE6xc5eLBMb7wcQUIY5cwQqAZbzLlCRhyfs
22E8UThNbfguUx3JD03tuRgDDchbNwk8S+7N3iUTfJK4/gQeWmMTQx3ZXZu/h1UMPQAk+Sfi2wU6
kZbNMm8KSex+qHlLnXklBpw5gm4IYb3C8uvAMHtx0JV1ozz2609yB1q044CkDtZ1CRLFkTx3B54z
IxTLTP6ztA9w1QUOTkx+wc/FNRPwdMCRW56DQm6EGl21GfEskJrrOm3bW35Qsc1NuTMHn/fmkJOZ
tuMR9ucgV9nFo078v5Oo7MA+LNnKzvKptwGMteztI9R79cFes+Dmh8gFhe0eqV9QNm6V8pVlXype
JSi3WHNvw1TGFBkxJ3uqDmSU063JUq2lRqasmv9vTliNd2vL15VYTPwG82Im0dcMklTXl/kCWVOf
DnXbSlRz9odzMfPsBYqs2JEvLBJUCjTh/RGM7ED5mdueY63Dx4AYYbd4RSVIlhex8oK4+tzJfV89
R4LCO3uNWghlIYhOGZNF3l6fIxiW9JnMjEFuNdwH1AtTDwe1knfJ37gFlT48MxO7ewNkATk0JK/U
3ySt2Eo4nSs8mYoKsYI/JnmHwkdtPwnUFxpH2z4SsN3/m79uhsdayWcIqW9nih5leOAd+4bkH4vm
opri7W+0AS5w3uS6Fh7ktaVoQ8terX7vVOBwFVrfGrHoe4IV9x7p/efY/w2Q85KlPHrraeSu5yJ+
nQAR4B9gnUv6MXNM017WUWn3JNVjoE+PSQexfdSE+AVsctQZTD/jURPaB0kdkvqKIRoPn9auLNJx
0zj+1Z7WsojLQwCCYNeh8iSJHCQJ++iNsZ+LlegeXsqBFMmHJRx0JrdcQAnTui7pBv5lOVaZRwHj
JhTKBQ2U19MXf9eyCXgzUpFTcYQbIPw2CdaJcZ1U2aPS1EmiyY+Oci8Cz/eyG9edc1VBkTxWdwl3
DVru/J2eMilN7d2nEJlOgATpwZSfaXqimbih9ZfmKWcqQfsb4StvsTf5zcdFx3hSY9Wu/cI/B0d9
5QbtEY8A6o8qrZg6C2N09WoJXc4ClnwjW4eYCMul8d1o1SAVqZnBJ68VYNR1KmZsKOK8zaaudFkX
Q40BNGdWK1BOZ/LgtrF8MK2VjZY/o5wXw8kaU5O93bCenIrfp0PClGru0S/D6d6FzSLD7IfczwL8
3VKUqVLg/hhtxd3kX/cz3d9FtdeqcUS/zwbBJDCyKh/ny84WYGAQKDEUWSazZU2Ah4r/PVN4fv4B
jAt/C2lN1YNORJ47SZKsjcuSM9F6F/os53qKYKTTOzYWZQpI3U8gpH+xN5JuR/RcD0c/ZIpmG6f6
ZcJKEMQjfFiBne0dge/Qhbt/k3vyFkAfDEgFs2pg+Fvv0Uz5JnbA0x/hrXkfJ6mcYUqKB6rACMgR
lX69PKTV93RPVIf9dQagv2n0YORvsS7KdBPdFpmdUoT5StDAKl66PzXGEGyEBWWW6RALqPfigMXz
ERr9crMUtHmjWL0szaZR9FpITwngh5XhHROyJb8iZBxl5NWyb1B4/R9rFp9x2cu85K0V+2VcFxPU
njGPseDZuWpNkt8wQn86pRJq8pGKzLUJ9YOidnIqS+qQplkjydpndG/RU2WCl5+vNmpoCFPSiSwN
DoQQRx+7JgzJe36SnCDPbub/Ye5OYrlQwMQ4dbtp7uK20HGtzRrEAHHhhWplvlwoxr7hwmJ/M+Zm
BCDnLfHQPp30tDXZzuPFozOPooQKKmVaPZxkZmT9+95vJVrSj7nJX8y4+/5k9cRmcn7FcInOKOdh
HILnPqEw0OvohdFkBRz2bfuORt58iTxInphYqXGpNxMTTeJx8RepPY+9ddieKA5Ro7amaRWQI8vM
uYeg/PIokacFVlb1+gllgNg411QWIOoHbIGwNNLyjmu/e1oM0P5QeiQP1g0NvWEZCczfmOnkjoQd
N5FaEKGuS6OPQxUbYDFampWyxUmYEVliPlsQWk//tCLCFwRBZ5VxUSmnKphCYtBKoO87fzgvDU9Z
KB/o9Y1g1FDIsDdMS162cvQKDFqY+W1C5pSz4HSji3KkBatjK+AdZ9mQVLzsbtpmP7EguD2G3LTL
wyk0eyfVB5VeiQA+TyEvpjsHmPMNfgFP2MQ45KpyIFlyPNcFpnvTRhZ9/NpMbdSro5ECVs9i9/n4
RLwMOcJ14TnYuqZd31uy7ATCwolNWSuqeQUU5emYuKj0NmjD6xuUmRA9H8qEf11NYkRjySAitR6y
q+BMCyU1AxhqOSdc8/b7ouVLdr+1WUzgFrbidFp+ZxVGYaF+qupSOh6ZkGrW2axcnWURICR+sLUI
qAXFsPRKF4UCIl8Fxkxgk25Q+CnO3nkGgChvKJv6x8CyjPGGwF2ig81gGITDhvtE9ssTQJMym6Xo
wQLXn7gzKV1t0xcj5dIT8HsV3kqJqZdCopwVrPdeEsRZuNGIWspS3y74bP68oVpgiPQgrgRfi3o7
epwVmRyDResfLj2wj0DMi8sgpS4EuV/T4NK0aXi3sKNAC8+jFYYQJJ+t8XNBYT9mCuvc+tB4Cenj
57tmPLTjgf09Gaxz/bGLd5wS9EqFwvvWGqYpN/+S601g/PvLFxYzDAoLvW5fXKnTQJ7h7/OOOpK+
8RPoaKph/3/DX6t3u89xqIqDN81sI38+gwJX4/07BaD/jrLZRjvzoVPFvgqE010/2DnBGKUnYe01
IStPRct3xY1Z9VZ21/usqTOw8sHmbAGRQok2jRqRWqcP0+jNRVgrLtc0OOx02dOav2y32qSROMoo
kqeSsC//SgzQ9BKhnOyB3RJ0KvBNVZtU6vrCHZUL2Kog13Ii8//u+b5BsUBDawK1LukB63XI+Iz5
KI7OrhYmef5FAzOrPaJ3oOV0cW0IN5k4BNene65DS0tHZI72BGmyQkFey/xSE0GcS9D3WyCgVi9y
3hrtOM663F2Kyji+XCQn9sV2tYh4b60JcG/lkpevyHsQkgD3u0NWeqvg3s64Fm/GQ6iN5tzR1PwG
AS0m62t3OwgZCgxGgtxq1Y4dP9W2Hu3GKbsqPJGSAC7SrQ0LBCoTKAc0Qiah3axa16vU8OWKKnoV
ufPrQ7W5W9dnoTqKrlIcSA0HRIgsC6DtTzI2SxiUS8V/PdZIEkIyFtoxNWAi7VEExnEZVbIOtFj7
G6bhwDLLeuLG1akgkGNRpNud0L8mwh01Xfk6PdbhGp3qv1VADDfpz9fFBufWXi+EhahHe3sTwkbX
g1LEPuQ2blmkJE8k0jRBoWvbQAEyqI/p3Nl3WFUBKHAD01XZ6IKKUCcnU2Tpw8xnDrSjWaeGsLun
Mlns7RksH2/pQNMuR0Y+WpmVt92mCWfQkCFaabYYCFYGjSMM4CXyoOil44tZ1Plm5y5MWl7XmHPH
aPcJwFws4K8ISIkCHpPkC0puF+jNIR1ZqAkT+AtNLeKlm3jI3zL5O0OqwVi75F1ZBk2fSC9g+W/d
o/uyMVcDh1bRclzedO1Dnp1U+1Ibe4GFHeDAdnH+J+dNLj9ndVHlke1e9h++XN4cDxeHY92EewDl
roP2WQkQCaTOLP8/azZEdZsNaY7Qavm991ow6pKzkWNEZE2Vy//8n5OxA9GTWD8CXiKpkDKizc16
Guky8JVk/gnz6PMc1Amd6MD0MMbt9bd/kzHu0aN+TyGZ3qKMmnusQBMIRGWeVGxq194Ohj0t3YDH
E51falRWo8VdFJ2/27G8j2wKXyEhzpUY28POKkVGBPEaxAJJ2aBE0vuA8sHGEAsLi4ha/gmexUzx
xdDrmGEJ0Qh1e+Q4AXcNeXBI9oXzhbGWxjrI/I6w+BSPWgX2LEAeh+0OGyXjI/HVS5Wfjk+aR4hH
Nfih7hp9Egu28DkA+WAEo9yopsZII5fTP1hlga2MUBCmRvErWQPGcp8nkie4hbLCggbmevVV36W5
eA6pudqkAYi+ps99X/AX669GQ3LjHjNnAIG4/4MLR9qjMQUCovCLKvUhPaJZIDa6wPEIKT6DV8Qp
VDfaun5zPenWeNCmp0WfRh1NshazilgUU6uGAUIcCBwO6PdBunD3J4hSHT8bEMtrOwSaFD9n4Fv7
xPmCvS0/k+ukGBriuw9hGxtDy4IUVSDhOrpkIZ2Zt3iXmjAz0Sd0zvb0H8i4nwhxL930IoOVfI76
LPSrcsq/8KuBNJC8R+kH4++y5yaxcMIgBg4Fl8mKdgXLmcX7PvkIn0tEJJi7KR72DCLG8mioL06c
b+gtroLIKXzco5nX4uNqoGRHzQcg8HOFNOHcQfRRlVJGdGF3AOA25+ojQZYOsJubg4RKeumoJZOa
H0oqR7rt2rYLJWxDNi5cY7O9X8jZV40DmD698X2hIYcGqDdZEflkl3QNyQdiaS5WNaTsvNuWW1ET
EhRqXkNqqxa+low53o/DJa1gUdiRUx9AiCrjAht5RDKIlvqGfkF6pZqJaj9oZ/XeTAbUKQOlo6Gv
aqB4A9LuLrHF3hh7uBacTXkLibkzt1uLiG1hEF3342cSBBN+693qAlTafVrThu0LC3vzRlGiR6sr
w0gU2XWlhFxhNpjT+9xJ23Ab+IBwcIm9fZqc6X9YsQeXmCgc5Cqqc21LFIrl4o1dt82JX54y/Lnv
0dHupOYob2jMa1/U1pR7GZ+zOHrcz4MK2ILdWLEWXB9MwJph1frcreZ+jrWllffZrAr+Bks0wy3f
Pa/yg9lytNP1ktP0CMy+pqvnm5C8tjSkqMsjCC4v6JJ8+lII5irDQKCJYZHoN1ZMaIPMml+W8iYQ
WvcsFJauTHKb/6035JEKYzLrqrRlX7x9apuFt8AFO82jIlxXFIIk0aUtI2JLHR7U43FLSGiy7lgq
grQMm7bYr60DZuGZ9I5++znkm9PYf0uWu/gbTKCXiemvkC+kz6KTeUpuU8rwCKJeT0N6tGZTtgKL
oBG3SoUC3RJlZtgmhMezHqlaTJAqoT0JAHnOL3Q12OuWVJuJEibV98jOj2s/4T5ZxlSHofGxRk4c
tR9DOG/lOXGjfL01nmRFyWgmL80ZvAgYbi+NNkoKiWvuPLGg/i+hLahvXrN3egCV9RmP1oO5YkiU
Wu3h154AQCO3E10eu8R6DHR0JpGxa1H0qOdu/9c3VxD5+HNefEXKjm6VPIm2ij31kvfb5/3IqRBT
4cny+1kunaTroMuDYWYo2i7qa9ijznnJMNjBFqURuMd/1C83We7vsf4BeQspouoFc4DfsQyc/MSO
DLXx+UGf9erU1JbX/lC+3Y46NtQJoWk4PkrVTlN2eQrdmp0ZIVjWhy5NtfviOiVkfHO0KG7Ux9PS
Uf8RlYV3Bo+hU7LUIEzWWeP1zjbcGf+oR1mMfavfUz7Tk1cDw3oa6M4xGpMlD3amOY9CYAm/qx10
3AmkL353Zk5QS5fPViAAmLJku9K8V0ulKIthvszPpbZe6X1gSZ7pego8r/0K6ktdRqoQGlwO3cgS
izqdBdjCb+mbcexcPVLcblBT6cezZU+g8GmIYBWgul5h794W+FRaxN5sDXBQy9YQbWUxZ5AzXN+y
8aww/v/BvmxkHJcL4W/38YpmdO2cvwgXfaXgY71OMc2rnASAjmqK7/VS3k0iZLRFb4UcLfJrC04M
Ss8u+nBtzijC3Q+L5F+I2Wtlb/ye4SpHrWFCVWITQHM5paLCu21BSYcQJ+rmAMQkU3EBCw22S02V
Cx9AsGAMQEkk8Snl1znoo0yVw1I5BqXcLXLLkz9k6R/JzL1Lw2JjO1nFXW5mmNP5B0ABp0p91HWF
NjjyT556Y3q6UjDmhm/8rI5N1iTvqrl68tk4liCQz3FEwwdeialwmA5TqCZTh+WKCWlZeVHKhrKe
+EYgyDhhFWXwjWE46RRdPbNHsv6e3Qu1g7SNhj12vMDb1GyZxWLFer5d1QoYUhYFLqmC1lLppePb
gQnhVNcJ3YtJoiL/fh+AaSBdfP3n0COl/Kt/vsbvc5PdMgrqkMzBO2CS2A/5zbsDFmUqgOfza8yY
HGsOsYyenTuMcDR2ygmqYT7zE2GZNkIRDjudpfpAV2fFNFue36PNyxeXr0/q9EB9BU37clc6jCLb
vagtcE03oaIyLY1Vtz1hbWJP1dQH/gt12Azal74bPFZ1EBNEwsq6JuoE0boR44pCt/VVl0dVToQT
piSdMqSrlwHE18ITGyuG+NocexxDisTIunckdv9HkUvPdDMs2InlH+aHfEYM43eU3/zGIv90mF3o
0JrYOwOuGrisG8g8cbYTN1rt1dh3TZO2N1+nKXbtHlUu/0FbbZY1lxOD3dL0xCHazDiCMTxoQ31t
q35OeJlQKQdMiwRTZTtNSaS0G/n8HbB7NFJ5ATmzEh8vRh9KHNiDfA/lxiH85cq1ayhzEbXBYCno
GZcM7QRdsonha07+CEeVczHCpmkiUJGmZL+dI8tjbB9xZzeExYv5XspPZg3Hmv+a/uZF5BRp96P7
adGtix/kELs6WzXssBlno/DaqLG2P4Cval2lLQPrQlgc+BKwOLN5e28OXlsD1RYwoZvYLccLy1lB
ljSWvSfB5sGu//JMFeDfwyKvIJeNdQPpOsC9B7GTy8aay7PpB9VaAwUXzTMdGhjcfQYAytpWm34I
2aUUFSiDesvd+qJU9PH39Gznz+SPpd1mcBpKxqp3PNvvAS5PYz9RkyLcjz/0h7vFBVMMqHCQB7/P
fSyiG1VXOqGEonwRRRR+rR3vPlq2k5KYSdwtCc4h8vLUKc7WNwG1FRZo9otI1sBWd3Ll/00/Gqak
kIM3GR2ye7kUfU268xbAl405XAezpklOCtyvIdbEOgLvTCsmZkeOk1DsOQp/8YRCrGsZt15zdEA4
5QbbVYbXUqYatv8GjNjbwe6qexBB//vS5u9BidxQVobFYnM/sBiI0NpLXlvWQRQkUq/eBCM8rBB7
Su+yzDhOrXFhCoNLMHIy8UN+3c37AyyU9p71sHvHvA5rdmpIBJ3ojrj0K/aueOOp+9z1E2s+8Ht8
FGK7dOk4LAIY1y/xHoLyqdKwthk9pujT7C9VFy93An2uKivkyb5lAkr29z5Ui0fBt0jsf79tubRa
6PpBC0CFJhsy8+7zXymQOezPuwnU6Xjod3pAzQ3Q2WgXJ+aGAWZkrO+EqvothqYXcoluVG3UoHA5
CjgIJqf1f3aaV7VuT680l8E7fE5G+Tu8bUIum0YLtbbXmlDIp48UBQ4+5w3GdJ/HOC89xXvoAR3k
FXm4muj2FS+RqTrbmczjkB+XAryEGn/POjSt/Er4+GVVrdgXgiMsL4kcl/3pwACkWYq7/Pt0JItW
2PIUC03ofPeImsD9TogR2cqkqhkwYe/7XUVnp4wy4E75mSq5Up7gQMIac+9STWB1w24mTAFB2wng
xicAztOfY06BYmIFds98E9n+pdhRvod6EeCNdQg+jCQUtWBIhEr5+BygSxG5hHkJ1uemJwsJBb1m
ytyrWfQLkxrztcYUwjLyZp5gnBNIHkKhDcM3pNU87ghjb0NfddQn1WECoeg0px7eO/5XaEUgB8CA
vm6JUy6sRGLY7IYzF9kgaWAI2WQdoOuNFbGsoEwdDhAWh7DCxGYp1mzzeKSTyFVicspeiSjT6oJl
izx0uwAOt8Z6oBFjiB3IS7ddh5rlH6EhSqPMNENNDBbcm3ro4c3ZOfad0cx7SzHKaDTpUBUyfzTN
UbmMlnqE6tGxMErfZOCg0MGrkUgIsDXgqEjph3mGLeqRk18i/conJJOT0dNdJKA7jfhCUU1dUqIP
YsMij9bv3+ar/tNoipudP8CRanhPYUZLZaBAdeGYpFfjosc1ZFB06MzC7zuB5bDlmIJWGa23vifo
b1buByqsOe51/HMdXhC+KGuxQLw4BJa7xkTz+rgALZAJ7i6YAicF+G+SUFsPH2zJQRyV1ksI9g0q
Q979cWgX/B1uGJzW8uNVIZzwDEhS445RkvdznmIxgg7JE56y6s8X+OstlMazh8DlEythqBnplNYF
Ajwn6nq7KlZAie8sfnWpAdWR+1kPu0gCowsBgeK/daR7pPbGfG5ZD1hLv+tIlcLgMUBZFSL4mThE
rCAOfdPqIGXyFiXr51R3+iz6WUsE7ObiIiz45LLBoL1v4PPxika3iXe/ouahZIN04JLbZCyxbxAp
KAfABNKTnLb3DY/LiFu2vlHhXuOjZ5Y+lhI5jOgMzS4fXMWfTphGLAy8ZJqaIDohTSLi/0Utl0lc
kkOQUnvyEcVdIlvnGKY8VYDHHkxp86ruwxH3b6kFrYau40ra1Ge1EjROKD/PYp5SPQdx3+hPflyh
R0HSfOvrJkVKm/F/uUwI9I5lWIowj/FkMUca4c2fIKrCOKJu+mObMxNTvLt15RKLWtvm3/TcNPSX
c2Ht78maqHLBmkTaWBxfW2GHX6FpAmvm70Vx2b4lhpJtVqIM/JS+Du4dI8FiL369/iE25Zx4WcWr
bbgd5cPO//u/UOpdSog8Y79tyz6MisMt5woBIcng5Oa6h58YgLSm+qsbHwIYpXuXzxR2Trm0Cb7G
M1pweWAvbDb4zHnab3l9MSLNYMp/RnXnGZXIhUqSH2pWsyUBMJLXvy690jwHN8Y7a6EbWwJxNyKI
vzk9cZrpyxn8MQRNxX8ft9KM/BaJrv29rtQHmpoLRoK9rDLpo5BBbz+lvvSs5fXpa7s1kmfIDX1y
Z3F8bGWvgZCcpINlA6YAum6CO7FXO7ykZBCgJbaU86VfgCIo2Ws1oiHDzmj76rV8VQRwbvDwbU1Z
casvQQ1ZCUZ0cdHpeN43r0Ej13kmaAs2E3LICVwCEiDjMijBkKZk87vOrybIoXAbr3hPrN9qFKdJ
sTmNDgsZVrw4CmYFF6dqf/Kh2ezwon/8ieokOacvoK2l2Fb0GZNIY7SsDwqP1dFzT2FyxBPFDHhj
c487AsQC+eEN7zvqOaiCTx9FxeZ86aGVRtbPLAEhZYyOaEpkqO8vPQFUu1+x2ES3rEVNUVw53iQU
hnKeVsjsc2JOkICXwB3lsk123D/WUKxHRdOsPSHqlbIEMGQVlTQDOm9heZ62lsdnIYdyIhmAlC5T
tjwWf1WPWAmD6vViQXLub620lnuQ/lVRPeEUKfpAxxO1p96R/vkRw8yuxD4hzfbcg5fO7TXr8IOq
J2ykzp6gflpJgWksMCxM9pZTPT8IUKLArMimh5NobtWW99PgxZWUYlIXZLufdzZyAQoMZzhfbqlK
O/BvGJ6xToPGXFjkHXtvb+pxAO3HTRohjKAdEcRiwn+1/G00tuhiwbgLhS7KmtGc1is3mA75uxSd
lP3KMYIklbWL0CQiu4gcai3tbR8qZplm0qHdH1S5nJ23QtP5/Qb2vq1+P3XO0C9Z/4f+36shzfhi
uapV15nD4qVNNGV2PyuiOh1Jp6l0wWrxqPDQtNYVz8OFOCNRKBE6AC3A2u9KW6Wn6/pL54v6BIuZ
6x4YVHEGBeOgdUHPXLQYI2s50EoaoC+emlpNJp/x0FF7CCHF5Rm4EWpHavusl7bUk+oi3hb6FUoK
3QLbtioA3z9UHty5OOCABFVkeUHJuXIfd4Tox9TtrjPb5zeupaW3FVLOVspg3asAX2ftI1iSDyrL
PlV7+L4wePzOhtz/rYW5+LVVkm2kUc9lxd8nn1Vt8fNqdHWhjAoYdztWPcKWqh0VAIVo4ytZxwzs
2oixgKLBkwAyd0Ka9Idnthj2rj8cgGqkfr5gwo7MPqXvCCn5n2odnv24r6rsAbhlUb01KGY0sbVq
o0Il/nSoxWGEam9dC/Vf7+GyKlPCuANvHLTK3KfMKfMZSqbYQ6oKBUnvoe4ZvY9MvNwEP/TN/Gd3
cSjd0jAojLdKWGtbA5LY8Ntm5wMjnNirIY34RapGxMDwZPY3/50swqYh7DxQaFw6Hb7tUPAe0uHN
27fhxwKA4V2s2lGTq71/cLR+J3NVTEX5iNleOi8w3YiRqOnFodZbSgxdDPvDthQaffauo832uqSJ
Q1QSilGB+0nWdToQgwMEbGvBVddU07IT6ZE5LKMD/w75WdiG9GgN8nSO5Tm2yvpqiOPWtqteqIav
5wMpTwHiwqds8bvLjJdo4kcckkPFbvB3M86KsGscn6EOzTtUH65GWIOqeXdPVub8YnuP0RvWR9l0
akQ0YZA7rvdymNfM5BltlaxpsW323OE09Y/sxEbnTCBT3wHsdTFf++TJcC9a9NK/L7y41D2E8Vz8
4LhavXzcNwu4HrylXA5arIvujOlPejc4XekaOiSP2/tah4xhHR+LJrk6bY7ax9rI5nZ2327zYdgx
i3CblovFq34G3bRbwKtC6dPuiyEM4LYrwSiD4fJOKZGNetPmk7FOC3zYiJYleYDm1lFxs57Km9W3
gtn/mTDVlpTskgXAnyqojpZEJqLpzgIos48ldPtM7Z+eO9eq4mn1adjw7Fwhwi7+/LmTaqpemeaG
QLpdJ73Ahav1knlED666pA9UEQtCFpxMhdVJgUAUDp3FhwlgOkMINu81dQAGSklr26ekD6QLGHKI
i/JFVJ8CO7VNCAXUUMluzmGpJN8+UfjOC/i0CraXZmguqF3iFWQEN+QE2soH9n0Q+elMvEXYYMlz
u4BMul7ON2hRCkV2/X2HQ/UNeDAOpgSYR/XbC02Ls0PTpUOPKEkpa4pm3xgNrQ9QgD1gro32rZ73
xJCzS1GQL+ImVbW4fPjqTfzLZma5zU/ZahzVxaScsIzAE4l7feAF1iCLGE+UJxznDFFrwqvncUch
QoyhfjCRtPVS/5AGh1fnUdjlDesF0936MQMzyXOb2BJw57t22fLpBXAUnauwbieVFJ/ejjVsD4bD
+1XWQBL79U2PayTvBgeOaE3i/mUkiIwEeemTsrskG5TVjnNgJmJo1wznQlwS0U7HpR+5xfbJ4u+i
71QWGPL2KMk2MbRNj3bjp7Egb1+6AHbQL2lBdmTl38mGpeqbRiWVX2gK8cgfxh/8GHcHsXd16XaQ
AUmTRFv2KYocIsx6wCMIgdfw9gfAiNCNy+wu5etmt5aoxLQe7V/UYgmaaIDjWOz89hOpLvB66BTp
GaaseAH0enXXojhv5cp5zfpGsCzJvCbrd/doaVnvqOgxCBCG2UD547sZXefP+D6O4nIkuH4TE3do
uW37sZppSuMqR5+ekNnx1YgF/nLSMdP14aC4dhDwn3fSSh4V042L2g2Tj7eLuqALfHE+4LHi/BOd
GUzwX8w38h13TewnQx5eUGpjta+YXxyGLySze6fIJVWNTgcEW8R3bc4inctWQi3GlF4ypsXAjyI8
F9XK+OSYy7SvC5SycAjM78TLUlitu8sKkRsV5J5vn6TzyKOzto8bxVSImPe4ZE85wanSYGfjNgtl
SJtegAg6e1beNP3vyfwdmLTC2cA6YoDYGh5Ngp6Ie0m57Gd9iQU1Nb5YFmTg+VIEsWfxS3QCEOXZ
1AnXTGKVaUcJeSbEI7FzaDvQ86gxdDS9UHJboQBYiv8aK21WWNj5f4ZHkvlapDmhE3Q8dowAMslC
MleNOv4CVAGyoM3BVlcPL28Oct/W8S7chY5jOPPiQeX+dERja1NF8o9+9eFAvf8y6VMmb6dz3bHu
R0878r5fInqv3aFtKOTlsTiEs2eMOi5KV/gGj8yKuFbTnpQk40Opt5bZs6+kX2nSYqscQ+zG6oIJ
Yni8nsJ380Uen5trUIzCKx5ERTLa0Mi9P5SasDRmt1318qhBc0Z5+vc1Mc1BhQ1kme6fBr8QYhXB
j7uvtYfQG1D6HelD1Wut0Su/VJk6gtPtyL8Z+LffaPu7SmBDXDIH506x5sqA3uFWRopm5vkbW0Ka
lcliJUBgNfTC1rkYYDFexZUaMVK9GoBOoVNUkI3/RdbfDzLab3J+VNAtRq8EZP2gf+1ZuWsg1yro
mJj4iutEQhbzeuW7HYTDNTL4emq0lQyALxf/R5PPMN+BORM3o/wjntdOHSDU8zsZno+bhNQo48iu
vEJITKNH6WtxlUNCyhP4dAw7A7wiYTLrCAz8ZUqLXB3a/MtZ25PjVGnw6QwYxLsmKVmwJlO75pC2
Kk/FhCGBcKTGNHV54qILhR5oXiHmNan8vvKFKC6OuLWuNowuz9ckfUW9o9gt5c+WVBau0EwskUwv
BBdy9Zhp96Nc+Fs3SmNxceIUAgmI4i+nc2U+LY533OMOBs+snJi0pL2+GSDI+S+Mgl5uFXXR8Rjt
8jlQMEmGDOAc95I6yXeGua7CqGtiMM2kSDUscNbOk588bPoe2Wgd7cTLBjy5De2cNivDusYz+MDu
x2tajtX0/F5dCtEggQTM98R+Dz3CYS4rB5klLO/45Km1CigsrRfQoNOgMmoBqRdffiy1zqgALhHK
FLbcNKZXCE+jitex+jLgVo/3CTk4k6qoix5DSO4uJy2wllQBaBT1AaVDAYlKUMczxt7F/YAi2bZe
CYuXy4BbV9zKz3wwIj+gfX3TB+vcEeaBRTk6y1pZZzZhwJgL7RYhQyEyxPHaX98U07Up4+mTIcGh
3Uis6ahBN/2apCJUm/6duCeU819PDYD4zApVKbFcgMbOyta+d8VAACVG8ZA3GZRjYUnMxvGezKnj
TZHrEdB8mB2ThFXR4LZJ01SG9fg6Te9H4AjnLiWhp8SmMqa4FWPvOLfeX832nuB13Kq/5W1528ta
6eJiKGZAp+PqOA7usvoQn6uuz2+wkw6QBtQIKQ23/8M1skiMhZo05gK9TaNejFYKmGggkRu46sKZ
axpOUsOEEiW7wUX63a/rhY0/z+uwgQrm+DX/dX2zb2SdIWL+sJ42nHsUxkmocDePYrjqukBasuOY
0DnDS10Ynx73JFy121WeNM8do+3u34ge8cvNJsW5mS4gRKElOgq44SKKFpDdhFRALbyso0ihYNtE
XsWAIkgjCWTlwAC2ksPwCekPcBF5SR3kro3M86PNWcXbLScf1G03Jq8iJ0HOFxPMlu/Vh3C8LbQC
J0HqV36+W4YJ+8XrXuBQjjDotrI4wOZmwPE0ivsc5GYAI6l1KTNa/mozWlmfnio6Pv7H9u12Xazl
J5tSfPwPz/U3dBgGlaw/sCtJ9il9GRAbNke94JtMvJlPBZF+ARIB0+1NHCtCmzHv5YgLACM2CrMv
Q241WEh4NEQ/RIwpPjg3LTUXnSWjgB9rqKFB9CSQ3ZSK26GG/zSRsl3OQ++qMq6I/9pTn4ms+ptW
dF/FWhIkT0EpDre1BxbXnX5g94Sl7L9dZBFcUaYzCVtugcv3kFVEeQAJnUZahvXgc+xr4NYOoRE/
eaAs2ZZENB7BGOxqB/aRQQUSDrxLmYChIIw7OMgi75dXWXR0hBZr+EA7fP3z8R4Hb8V6y062sP1R
JAwpV2ktKT91bLPHpRJv/zhU7QS2+969Tme0qDXorkBBE+LO4pTnSbuz+xe4VX33B4fws3E1FfGU
jgVXV89QwAxsh5bxrs8UzBWuMfjK7O8K9acxaRjhtj+soflqyc1LtAUF7qw0bUgytp4NRGAtYUgL
XDn6XGe1magJRW07/pnhzFGkBXmU8naOi0tyVETfK6j90gz6tLoXcKzTqSlR84ZhTLYX61StGGOM
9CEG9/iWLCwMhvz8E3/2OQ61fcJOTj1DqUhO4ral/Nt23NvxAUbKNtJyFCaAtGvN8w0+ULm9pe6v
/UIHwDwn0m4OkFGb/ERk8YbIRYsNLd3NdWA/fCTDR/gE4svwpJjsqez5EHji5DmADez06/XYk+wu
uAPUiarLWDu+RzH+D6uHrzR3wVIZtHcS8PSLZtZHEgbmmKjP0bVEIFGuJMNmRiZos2uZQcYlEnGy
pXgJIjEfzOYzSAtd0/5CGNQbRJDar6UR1Gbfom9CnGKvQtbRP2Qhx3hDWkWR+oSQ/+NFW4sYfA/u
WkR46jKsDG2nke2Br4Y971j9TblLY2Emw1ZbV+m1GtCVggVReXmPJKoOoAqYIaMOzyud0cdmTH6w
YiA2KUR4Np4MPh0EFcDdJC7GRYspknOpMmgyNMD/hynD0VKhcIcRNbtzAAMgnlfz/iv+Zm1Q1XrH
gptKy1oTg6Xa5eS67NYAZ/tnkM/oyk75Bm0XmHD7AMSng4PAIu3Za4nz2CjwZhnCiW1oln60Fqkt
IYWGMOsnk9HbV8gzVLdYxfP4+9MZ+DomeHyOSoqImT4VTy7c3nJpJtCWEZwPPGa9amGgiLWuAD8K
O51PyUwV110v8T23pJNAywAhpeqfgKtwwSOZqLpuQqVs9KpkR91TFBtx1QD7b8hPZUSVStw6CIJi
8t3FR6FdejDBH7hSqVHOIFpX0iVzoWD87lmbAVNXj/Yuzwit4kql6HiXKgysw7AVqLYMpkvL8pWc
YTwonOueiZt0tYFjCF9/KqmhSc9B9QcIi236vYc+Izq9iiHjlWZSQI8fiifSvw7j2ipNfVle6ezu
D7zYKQZqlLgk2PPqdkncXXhKnF6rsdBns7T9eyHqBvU+qVgPeNqicJ8FTaA1fdj7i/bW57fz2Mpo
qUO2gpPN+wpraktZ6oAi3fqnGqUTwdDn6iHi+T+CfAPTM72HgvboCdbOrTNwkDI1fMLCXPLDBgbd
SC5DNRs5MfFkobeO1Rugf4k0B4Xb0dIKDx4QCfDARVYaFiwjnnbvVIvN2nmtKBUfx69Ipvjp9JVK
lyC4ZUegwXHaFehZUzNYEwCmc1A5D82K+vEMOyVdCs1oY2hyfAIFM5RJGfV0rBE/mVRXMzGV8H7k
e9RA4mr2P5pRW6EQPVUjFiEw/AdNLjbSBtUacH6hbD+e6U/gmTIwpMMV3ECareAqhhw9xVadEb8d
N81ExyyTqOisZK0p+ne3fI+iP/+TsqPu/W3nygRq0t+LODQwWImrmhTAXBwoOILwkSVgXbMxTfNm
lUpiOpYTRoVTk5ETpaUcnNn/XD8veAvYxKSBCAWobr67pK8J4dsYr34ODQKc2CP5cQrrMrQTRwL5
9/2s8rRn4o+ECz/6e3jHHYSEAQVTf+34xBQd58rUMhQWkb4yB+xq+e+4T//tiI1EyjOEiq0t+a34
DBLqwgFMqlwTTXTvE6/aT8XNZaHshcigvukCzAjSweamzapMsnB96oMQYfSOpc53OTN1VJGWZ1ic
bndXh54chWlLJC4wwGm2NanLr5SN/FwQXeqqgLwPAYULo+alpTLmqLgiIK0T6qtqOFzYkbPmIZLf
55wl2KvJAJm4+sqrkEvUJxbrpy3L0VAUosbtOItr5Ax92YSd9M3Y1P1AyUfrJrLv2hg+hfIfYT54
HmWoti5l7DzHOaBhh7unuQSi8r5O5JVOrw6EVAD7tYhSbIoKfIRoDMI5JBCm9TFn2yJGEwrsB+GO
uI837mPqz/AOCgsLrizOZTw8X6EiM5vofWDg45wm9L6S5xU0VTvd/kUnXAaysTbERbByYOExfC74
iDWkoAPAy+2Jwh6HWq4CeN4OYy1FMynE09e/sUiETaObsZ2DJTBWMri+vXiiIgOYJX0REkLJtyTY
T3DKlwKxUgUmpCoL6Gx/vyM6mlNkvFy/2sbgsLjBkgsY5X0ad5yfgSGkk/evTMpAbFRQ1bQmhsXn
/XegMoZAKp4Rq7iLAX7LDE7abSzw/m3D/bVgRnh3VFggDEVBWnOcrMrm7SCWyEhGn3KVFzlVdWv6
KyCDj6DYZHBSDgdw7ydcPKqCpH/BzPoujS/NulwtZjeDfr5Fb5lDxS3exEKMC9YuplTPgjiK1/Nh
Vm/qsLaRriyWtnYoZms3ATqpv+j+IINDIcD6w6IaG5Xo77SGSvGv/SXD+pHTxHhxVSGqaNUL6D+a
L5DhNtyW3ZPuJzh56GaU3LLOQcly4txDuIYHGd6eaSyCMdiErhW3QotxKH30ipud4fYLAoEfyjM2
3qmhyEeURZw5kJJ6ivPuyhK2Q7tYmHeNwkTYvvmC4dMOYmBos7WrxjuGGd/jQ16l9d5TPBgxsqSQ
9/8Y0H5N46Vt0/1WYdWFRihuB4x9XyE4J2Etwm4Oa0DjlBJK+iBb852CBYz1fwEtGDlLudF7rbg4
PbRHYDIlW81Syr6G+UB+xiqNAtQF+x46rw3IHBVTzEIw7Y9bRVGVaHLUXVrVCsYOw5l5sPN6+7Hb
mAdAEuJyvBmB0jfuL3pRQziJKLTkeKXQnK2eqkUuC4U7+3P2auHI10rqEwEndPwo4k8Gno6dvrM1
bf5cBWiqIN8tPgjR0u5KPqYEF+0keRRV22kepCPfnIH5M7CWqd8QnBCjBWejTca4WL2qsHohahIL
UahIWOfIS+dbZLbzY6mTGEt7y04F1SUGTtVbsOdRnwofOkKIDxp0mehEwvRLUPiBHvpcwGqz/f7M
hGHTnw00oUr6sXg/vSmlpFI7hGO1RaQWNTkdo3aKjejzwcxpFMyTochyOjZ9QOWB8uBXrfP018/d
mv2yalHRuHS+qfOm9DcSqEB34zqEIqA4FKnRakGN/wyvnFYRKyIM6RT/KwhUQRiepkhy9D1VV8VM
tkCUMbg0f94jC3J10T1CjMtRADz5pjCRA1TaLQHfJwoO0Uo9vNeKD2KJLWkgN+j2zo48wYEJ/JcB
xBDXNfPar2GTJs3Ij0FWLN9ATuvIDQy9YQrLVBS9COS4lTEGmJWcHVvyZHmAYbmPUqPZMAu1Rjos
LChjCZO7nvm9S6mPtxM0n1/vo6fP/ab6OLrWOdtdLRWiGwa3SVrEQa0zIdvUQutW7tdspmH8CnNp
pSVdAH5/qnO/9gsHbTWkYRd8cYcjmKV/xwNq5721vxbxEPo0o0fnCEGEHwPLD9MHrXY4N7PNIPzY
RGqzahATBI7tp9MovIefJf28g2nRMj/h/hb3770wu/wBRa42DUJoquBEC++XROrZk2lme2Bh+jMt
TrQMwxGlzJw76uL48Hu1eGWx/KHrypGhym3PpyLw0BoOwG8YOMomKm9Ym5CEsrzFrLJFgRyFg7x4
VFYthqGzFEzl5oI+ITDZ15BVFpAZiYz4PNulxczkPnto9XQ/ynmJIhN+Dt3BFZUQ30V0ENgWgBTb
q/RC9972wiirtkfR2pag9nfP2Xg1R6QmaTznBYpLtIG7OdaJPpp3rlcvyzZKXuJ1QnZ3RcKNQes3
deVC7+7ads1aieByKB2NRS43qSB7Lg3TN2eRdxOUYptMsiMnHyo9p2ly67Bw7Y86ASB4n/Q5pFAN
U3zOBJRbVXiK/H8GKAwTwPV+nXv7rTNGHKMMvPxX25Y/A6MqEiuEX3+OOcUKfG2bmks4v72OE61y
4VXMoDUTdSjr/M37yhsp2wLYG1g3vZYxWWJRX/oIpX7ijXmGfHE1hhBjiB0QF9qvO12JxvpoZvYq
UZwBH3s5sI88iEhnSFrikkUDmh3XJ9C7eLCFfMS/g7F+XP3YGKamD1oSJbXFfLNi0pbt10wPLiqy
oB6xQGdB/s6L9ydEfUzEp96TqjNXnEn8CzwAzVptN2/2aRBSlWkYhUdXXptawRJD0Qkz3aHluVkY
Xn/rPnoMF+gNQqzwJ0mY7+NproWOquJC98ya5HJXGzVnmHoXS90K5dzYf1iV+A5AeZNu6rJI0vuj
pSjlCRHVmbPriL49E5nJNpjr15g2z7Xil4l3cxswGoXG0g8xRecgmn+HjSaHkwCD2sY2+mpmh6wP
Uh6U7CQjqC9G2OkR3sKzGSs1GAgBLVEItZ5e8vFKFg7DwUS7DmMT61zEb2HtzoxBGIDW0nPmy5QU
UDAZDsHMHw0QzyX2d6r7+cYVEfYMgM+NT5uxYTi+g7i9MT8mSyvUPaEjn8lRR0YHEgM9886loqFO
49crlLLDpI49OLpDsJy3AETBvcKTPIqBDxNE1b0MVNVmjl0LDctPT8AzSQnACAnoA5bc6TMHX5rv
afEqyYvZnneCmxD9pumAW1HJnIlC9Um6borYc31e+Z1LpYh25JSPDUjk8ccUx7/HcivROQ1Hn+1h
XX6d81dWRQTJYJQEm3tpsE5gIXD8gscOX995zqzGMCkOe0iNewEGQk7DnUELHHY0stbZmg/8c1mB
S29AeMjsKp1PJOWokIoHxcMnS50IQEvVxcHmCCbQVDUUR8jIejqDvQXwVePEGvuVCbQxehzuW8lZ
uGnkyN2dKtYsbwQbPuHxUoEG24Pqh+lQIO0/eaMUS1o0KVCabt+CZoYigiDoK8EmNKrq5PZ3H7zs
u8R7hgECXSg+3PN5VJTu6Cn7r4ADv49yF7P68R6J4NlU1xtoHxtLUc3Z1f7B1sW4X6UaDOLe63iX
IILNb0JbT0YwcPg8PTXxuVZTkZ3vNMX7PAEhISe7kZ8wJXIrVK6zNtgdw5myRK16cRIVOUrAl6zz
r2GaVQYLtITwOzvPH6D7AldtCoxBA/htYho2h4ba69P5Zk3hYd/TGVMF8uraJ6fFKerE2vSDJxPj
YzPxMf4wIvSQBfocRKkP6ej1njoiRsVDAayCwB0aLePSbUw8kL8lG9KmbxdlrKPmf9fF/nRcX6Ie
27vo0/VkzJkXLFYNYeNjMpHEE5zNrwVV280B+sYfF2ZYBHdb0S7gW08qG0XMRvaKsMGDNmkOj4XP
YVn2eiG6xiWJzJolVKrI4c3Ox6KlpckGcuPwBFQIWvp1ab7zGGV6NXY9dCk1H8fZKsWHnMuCdk27
PlJMBTcGn+Li27nxEDPCmQSkvk7vrhBrVUh6bHN9oMELRQSXtkfZc+y+6wshXZD3SRO6xi4bCDMQ
aLxfi6cdeGRBr4ieNEz38V0vcQi3YeB9sv+kwLxoGBnP4ZzMcoYo8tWJ0RKT/OP9cSLjN1vgn8HX
d1/OcFTacxZLDo8GL0uw5nsMtRlZrgoWxPR3f0/A1jmm50ONvXYZZ7zEarAlp6eXnLHvMHifm0Qa
kdAkdHGRLoV5f4u/6Xt+WljdFnHpKdsvBRcLnyYDxR1ddBQfjNHmR1Pi3KOIeBcpGyoe20NrVcp7
tc+v06mXtgIuue6r1/4gIkQ781vobxXBDnAsv2f0PTqJ3JTygGgtWYDo1lnR+RVL9LOG5vGKiLJQ
2dTcIdguN9Eytn2zyYtc3lY2iT0SCDDEoUeKk2J5p7IvTHFkD9qsUAXUAnutlFK0TvciZwY3R6NS
lE1kKRnZTje4vbZJbFqwwJEmPf/5AzUFdiNI7/Ik096z3OLgNB0J+O/VHE9FD5lTNXWsfU8uxdMr
kyrjBn8mDHSESbE9+tRMQswtSstHVezqjV/YE8pZo2H1Bb9PEpZhctn5lJy9LVrb5S26qvt0msJW
8pJqtLWrWaqAJbaCy+JT7VALMUhHFL4ccgvpoHe/NkvgDHQxqKLtDv/37Qqxz9j39sDwYwAL4Vo0
qHca1YCcI4hWKEvPHVWvxEYpeksWhwcUhfoZy565dfL9CAp2eJ6241p2jxSI9nE1L/DvK7HO9TN0
9wVDsYaX1yer0+rLA0TLzu9D0JkLwUtBK1TexymuYb0mM+PDpmIOSFB6aEVmf7A2u5BEPg6WPjWB
iLkbInVwt5/ek5/NrArN+i5SwQVOItSLqXG9QbR0yu0JY//PSVlPykxeU1CEYrhr36pAr/XGjkNG
FAKfCxmoJveauCeu3/+oZ4JcdJm+ffycxnkBNqS9dzCo29EnX5UpU72FOnuWorhkx+p80Wm77VI+
x2YewLCEdz5fd9HtBEI8wP095cWKg9J71GA6r3+hobgNa16Cda4DV90Rhn0Wah9TV3NkC8GEhWnX
YEBfYtPRr68eGnLROqkNmJVF39asXbr7pdvrLP7ZKjo9LGJjoybbAntsa6EQHEUOZs57aK6Q3exx
fSi0sHqUFJKH3hbf6U+KGoQY9Na8RW51BRuBkPaLl4/WC3RsDVFpBBK4uXaDlZkxuPcUZFubfRzm
Hu5xJCMiXJ2/0pA/mCSJdDAY9AKjlp2GNId7JynChF1uozWgLNqk0+onCxoOsf+BCsA4p95VUF1j
cQNbEI1ifV7+PbVvD4wclPqiO1r/zUZwRR6X/WLr6pCjR9ZHC173NT1qLFf+DHGZd6cI0emZmGic
f1ZF6NNEcfED5JvnRvYlD4HjvdZqk9Ld6j8qILbn3chcr0iKkxza4Uxestq5ivH/10buypgFs7ix
AfacQGvcPW/WqZvRG3UsmURtZT/Lr3KnFL28BallsB2TrcOSBki9YBgTf+Q8s+FTeBgYjzmnTfuS
/54OCRdECCCnM1Hmtq47MF9MRRTRNGLPMPSgPVzylEN7+TtjSpLWzmpWGlmUHCThPBleTxlIlJpY
bhTCBcGJetlHKCJw0PuQaxIfxQrKSFcOIRlEZz+yJlpvA3Q3ZQYBf40U4LMpSTNmnTqUYFmLeZo9
FFu/I3N3qxJvCnYZ7Yvy49fF+K5CmYPcYWOMBTfewwtXp04vAT9DjdkjUZBbueTt+JHM3EYLMXB5
nM6bwD7Q7MrLrURkpjspjGmvrcVVHSlXgFQSso+6q3W1WcZWcIJn193E2EUrHK7CEfTQfkdEHMGp
04dhZ4P9pNATSuIj2IErKaMQcTBDQ+fb1PXSqLqcJHGvxIAM21QOgtQD3+GKJckigNU7MsHg0dBH
vhMFuPLsZ1BJD9WrINuGadYw0U+9eJ7qFKSqzwbUfCK9cyL9cema9gXKD1ek1l9pBKFXaPUc05Yj
73/mb9pnbql441EyclZVrDhicThOeA8V5kAFq5F35OK0210KAmuVOC35CU0BAcuPOli+MyvWOhia
7YE8U6+4W4Co2uRW90oJeorlF5OEPuJ8TnQexG3XdR0KA01v0f2bIgJhkclHhMrdcrpr57sT4cLC
aETJhi7bt5AQ4Hhg5vLaAsEqfGSOHM5ObXiP6jg1sQojCWcqycqsMyyRRuke8Nz1BfORvHCczbxf
e+C48I2We0tFqQucRozMud13Y5YbRUV+vi1iCoUCiixp9bTNM5a3jTsTzAGkOUN9MD9kcgtChIHl
U0jjCv3Ceggp6RTpzm2RzNHv3kNT4JUexapaNftEEbXKwiFcX0kuU5eO39a5szn1KEn7QaLpRWzM
UoQeEhFH8T0Uzo5lCI94C1OILaAovVPvg8d6xznPv29gh3nrWSPD4G8BeFQdKvDUrxoa1Bd2FZKT
YKR7/tGj5u8upGWSuFkUYKoxCm384kf4+A+rubTcM76rOd0QHln093a2XSR5z15Vb/IHng73Dfip
789FecLg6NnDO4EWInLY6a8cRpxzAQam2YUutRFI0ekR14RzK67D2duD5Fqi+dQEmuD7SJ48fX6z
gUh9vQ3yVUVPfiJNv0FgqOji3dkq8TzAnHYJyF6es0UhnsmjTBEu4SIyP1bQKJE5B+tw/m5xfH7N
N7ZAGlPKgSuKZBYj77X0qXwqBo8iPoQhyDf721ZDYrZe55X2Eu2xIMouW9H7fM+RkpnfKZRF45s+
QPgNNYFsqEeOvoZ7yzSyfTAcwmPJeDZHD1Fwp2Up0gYOrHPD8UeImTLZx0BiiAW1y/GoA+QeUp0R
oWtcXZgYHClm6Ci9sRyZ/qNS6bAjkArWdxciq1lJRlwKBCYMWlQz6zzKpsW/MSydxBOhALpbLnVj
SoXbCuCeze48Fe4JxTX3lQqg8EMJUjNX3ofhDCTsoW/FYg8CV/p8UHcJPy8aEGaeUUyoCAm6Mff0
DeVVqNZ1fTJtIaOyfndMbQclrPrYNRsmiUh6Ee4q+RfFWs6gJFlMxdCWTspoJQ6xKC2DPreWlxRo
I8T8xdr6u2vYDyb/BJq+ckJnD6+EY9mMs4fT5qH7dCP2OpRjIU2pED2x/vLBWHOSZvP+6iP7f5Xo
64qvYKPHd16K0UwxRqqKO7tvEbtld0R/aT0bWip6gK4rC45nJMxTktvd5eGnj+fr1NRk9pAUsnCS
i4WyYXtWT1wwj+qyThLPQlkUBYWKRFoPba1tdR5zJE1x1uvB33fWUgllJIP9RxgjF6XfwlrV7OKN
M2IbH4ZEDBdVWYn6e7f/ayAPiZkZWNQ1mWC1FOZ3Irpk25G8tBP82wkXis3Qpk0p7bat5TsjWDUg
mmirTH/J8X5kjJN4uXlbvLy7zhIKgWN6kVpoTf38hHCtrXb2GSntqsQTw9fIwfyBaZSWHk2PD5qb
GfbayktFgu3sD7a0F7uV9IWQYWxf739lY1i28iRrPjtQumNJtpTOd/3lcqE2BvSKq0OTjT1nhF9b
JevImxFTkY8FZv8l8nEW7o3WnqkxlXOSrw6WuO+CF5yGVTBRsv1IRni0Q6yACDXpXK1IkwAqcSIo
QkeOvmTgHSN38sIISPeuESMfrkRzzwnEaoTd3p4/o9cCMLnaDS/PMMH9m4hShQ9jN5aaLRwOQuEZ
Oj56+LqsXuQnfjpKm5Yqmr6RW6MN4jh2Eu/pHRTsLQGfbniVmM9gWxHnZKyUMVzi5fi6UzdiMFsF
QoDaAQovq0oG73qd56OAr+ocOyP3rD0qdjus3HzlS0Zqq0Ti+HXfd0a/egrPN5nF5vIJifOSV+pW
GliBE4VMyytswBRVyX5MqV3oKnngDM0anF8A0Bgx6RGGOgm+VX2uOvS7zLopi+VpK+VxP7hATFQF
5IQ8/cnVd+uvD1pvZV4PSs3tTtIkdO2MyfD98PzBFWIFpUl57BFJ0kCeFwc6jjosAe6IAGunfjbe
phu8TE2yRq2aDwvKBZ94OhLXA0rwgI5WmCWPPo/KPRusNsr2Iwj+Zo/LG9qvSXL+x8WLcRzn/UWC
iBK43B5Vr+arjC1F03Cs+T4kYHO7USN7X4KOP6rQE0EFNlavymgXYZO6+aRnnbEBa4cwrd7dPWjs
z+ruDd2vZOS0CBda5EeFKtjRdNh8Qdtt4phr9ob+PW628pENrBy5PqAP0I+rAtLdSzO5BufTKJn7
XROhl8XYVNK7filxTQRHSyzUM12eGzRP0fZtPe3+Bo2UtclAZs1n9/2jr+POLmC8OWLfIqBy0vvs
RPAFQlrov4qq0H8Bp2WvJTsW3XR1p+8KlwIbAXGsCy8V9N+PjMTzg7l/9lQucjn1wcRzesR33AO4
ZPOZdOZg4HTLQh33pDYVF3z0WScOEVcwQGTL456CIQd7Xb4uBMai1TnVyPEvBWaOdtzcRM/AS3LH
WCEo5VlGDsFuLdm6WdTRKTRvOZrTDfd3kZlZOaVWDGRLjApVUEWzf/IjVaXNr44tVgcgjGSMJTad
PYB4HhYMHdOPPjYLFW/M4etszbDIXpfelQ8HCgX2Y91FIcHXEB2o60MNilhRtqdxexvP/YdjyItP
CgiAK8z3Pt9yqtbvFzqqHs34InJUvntdPNXhkHAORhiPOUEZVVuqeAYzSxbzSW+dj5x3OnjiE2V3
2KwZ9I/HKZHFWKFqoyt2XhMM1xEO44OjfKP4ArPdRA4NZ27JpMzqe89BquKERr301C6fXTTg0Lwy
4lkVsvSBcUKWCchkcO3AjFCXObMXCxEQ4K0yyxF6rkRASYVQ8ZIiJZeXR8ohJX5191Km8xZWfu8g
Ye3ubiGCBi2hTDvx46XIYq0m9DfRNnBPYJVcOmb8Oq5bGloyJrhp++WAMZzFytBxqGTGxFA7SzEK
7LehiJQcbeqdEUHR+qwcdcoqShwXK1C/vba2Dyuhe8Wj9TDje/z5yOZk80WFiaZzlEq59eLCTom2
i5EH6jgsK53rDV/tRNfKUX8e/PktnXeCImL77vr2j4mXyaRaS5U7tvo5JUpm2JSxczfY4gSdEFRL
xZbztFRNUBYwNIGkHhpOrxYh4FlOaPSOJ+nscvXyK2CF1Zo8dziNz/aAvSAFuk2dsE+o2ebm+zZ8
9ie3L/PwYVLam/KxfMpSO8vz3Mrt3MtK25vPWlz+H/cxdzj3PH8nKeW46zKtRguhtcVv3qGEYccv
/E+UIAAblgClnJVKNVxC09/W4wzGR/2BWv3l/M516qz8Fzj0qy5u/NjGbjqfY3LWbWY2E2ZsNXto
TjFY228OiuKRWwjiiR2qwkrodSaTCbGNpzwd6GiTaEbW44knlBHn1ehoR1Oj5rd0FotgGtk69AKj
0cOU05hp2DrcEL7+M72jogs8JgJPRhvhx/ifedCjzVmodoWffYgZr0Ffq/rRJzVU6CuFIgUjU+cx
205bmsEBchopaZaAxwTVuvlk2lo2BXR+coDOf1cjZ9zaARYrFvtS6CD/5JEonKNJ3zWPSoYnOAiE
4fkYR3FPaLXv9yXrpnADXu9eeelGaDL+k3P54yPhZAkmLz9poTgZyjkuuVC2GbpfxBTZEj65ufUG
NFuwjniYf7zAm8LmnDlH/Saf3KwkEQXDyK8Nv1YjsfzUEX9fMcfZE9jUYYXM6Rzue9G16ZgM72Q7
mkds1UW0yVqvC+cmRQ96Y3mmVKzPijc2uL+Ni+QcTXMt9hEH1KLkDlrsh2KZ/YS+0RhiMuLb7Lqh
2TuEfdvJGMIt7kdy1rLCrhhae+SXUQtOLEFSQhLtQMqSIBTH2153NvHinLHYq99gnag4HXZcreg6
g6jt3vqwmdpZGg+mBG6iXAEnFdJagIXadL4ZyTvRuQfCE/6flLtDR7uxko7CeMmLTbygIJfDf9cE
42lL7WpbVDACX2Mex3b7gYUeUa83KWxWFgrxog3rQRP8lPSHRnHziiDqiIpdSpheAIUe3KaUl7y5
JbEnyduh3+L4pL9+kLfJ1DvgAY9NLokSIxoVVepXbrBeDBEvOssFPDsq2U0+54aqZQVsV1SdcZhz
4WdA45HmFVXSyml4qDWXawJeWbxqaA4538NuMG5E7/S2GXYkEB2arrwtri8E47o4Q12/vlzuKUFp
cbLHDdCq4MSuK7tNQQrhF5783picwuSx7PvWjgSXz0FBOW2BsFZlfuNrecc4eI/JC+GSR8xxklTB
6dN9eT8+Xiy1AmB0u2Q3A4ormR6akqKS+K/lDr1VJpikRulghaaf948W/bVxPqkrIVHVeNPuPWp7
FgY9MPE5ZP9aat0WZcvgkDUMeKU+L29hgNAyYNi+l/yPcj6Z92flshNGafmLhbppQZ0X471bmDTO
S8rfp12qc4SSVGXFjSMydzyUpgkCuckzJ3Spszl8DBMPo8VKgEU1/puiH3e82orFM3j9do4PoUZc
eaHx/QZypwRtW5BRnHjyqpnk/+iHREpGHMD7zeG5U+lcIsfXg9p5/IYgQq7Gf8u+rDrsDGuRj5KW
ul8/abS+UqCWDl1NK+HigW+azZ2d3Oc92VEI1ycdBvov6aojx3xgiPpWyoYB1FRSSdYoIC4oTClV
YCfJue3BOQLFECc8CV+YlKYrpM3q2sfW11tcIZsL2rhNJu+7WhTMgI7IXalfjiys3m/CbdODYZpz
CJgBrgAuMEuv/rzxd0w1LYV84uMAqKMf6Xi6Mj9xBXd+mhIQHkjxBU76M68jOPEE+0rlKJsi1PSb
V+fzW6hb9x9vY2kNlTrTe2gj8BdlqsnnRgt8WNtU4KtsPfXHMkiwXCJldE2FSjevnn1E5jSWuNiH
dktBs8ucFhxYXCVQ4HCPIiysxiw03a5xWkHxAt0lWoGQUDjFBi27T71rLjYLWP4CEhR2C+UX+Mo1
SuuUcINtEtpV+IseYtJvPzQFUXZ/yocUeRsGZRq7g41k1J6jjM8R5qrZakoX4DOmbbhAq3FNMNnw
HBxiTaweIb4LT00ZApyBdWzLa4EHOxlz/0Ku+7DcSqoI4Ijy7GB8b2+6tcP7/BkDIs3aVt1lq48+
O7dq8CvBJy8vLXVpET0CdiMSAm4PrlYTAD6PdK0sDDnUbKFz+TR8piCfjnt/1k8Ko24/c41m88VG
Zrv1rVOSZ5om466YPYYC+c5qklSMb/YqX/bQ5SLQEbiDe5t3U4+wdETZNOUFpE/MptssLePqANuu
Gnxl9T2f0B6Pl2MB9trDGyW2w25+edCZtwBxMGgc0yCmUnkPtYQ8clconqhSRX5/nVfeDnApkPSE
R74gB6DEio6CQ6mazQm1/qNa14tEF3JrCFcB8AKFDDZobox4rj8NuNdDJrKSqBIDWZwDXHzJWaDT
J3O1pLF3/APh9XDqkJHqGAewcpgfGyca0XXVOkAzpezy2G/uccpAtmZEjSHhOJeXK1SBgwqxAjuU
91/0kCGAE2ktmwAXcbLglip6l2sNzGJFo2hoeVdGsp2WBQx6XgwE+h0Je5m7Der5bAfmHwZ4w8jE
J5Ciz/uvr7LtWWxb9JRcaSODMZK+6SyBasOza+2fxtfGSPeyKLC/+YE64OulXvikfPGpPtaArA5z
sgXApmASTcjU7isvv8si401vb6e/SJ/MHEqiFg43D9fzpx9McGZNGyhW9k/FY/I1WFH1RQ1aYR48
KjEvxzjmSrs2l1y2ACP1JwWH+wzz5UgrWa7aZLTyn2IlHRkmQ1gph0zE5oNFK9pPya3r4a3hTL/Q
mTdTLNAiPBiN35+VhyMJcOItcwA9g2ONPhJp8yPzh61QRBCCkkVkZoq+Omp1BBlkoFbcdTk3Bh58
Bywn+YehbjKBJ36d6MHBGaiEGPV4zthQDwpPtwNhxAl/uE5EACdkkuySGDgoseFp43R1I2tAcCHa
tb/PwXFWpVGz95b+y5bsdTZFjZPre2owuOfPKbN0u0u+FxfeOqucF5HTbKSQZUpGMojx+6Ws/x02
XlVmHEde+t2R3I47tAlKgpZFIcjL7VtCh0tJv9y6wl1KKUEubb7UGLlE7TeS3B+ai0lXZm1jYd6Z
SPTePzYmeueqOiGSN2j/G3z7sJ2MigqRn4/0yIFQl4chiXgCVHra8S/4eaJ5tg8M9KBQAeHGb+y2
e910NJyzpsUAfy5D9UnWMIWoh8Db2jJPTsdW9GfFEWZFvR5X6p8Bs7p5Uu/JDUzHcs/JIXV49Pto
76BH5M4jgiODhUdP54epIEZYk5kBrS0taicXXYZjG4s3io29OoyY+g5Rw04/OwBuffosZrdQ4rH9
hMRaoZPQ2zNtCTsny/HXeH+HOz0sSrFRVj7cmWJtmm6S1a39r5/EmeFGa6Jm1o4koGjAT/TJj5hS
P5zBsZ0V3begKXQy0xrpyB9q6W9PWw79vb21PjIQRawmZfw9f6nXuCwD7cU/+7QxyFxsd9w2/uOO
57YgOAD54h7vcATbfnncB+Jzd2hVuuzyrdPCUi7dByAIl8gpaTwhYL7/dtQwjy0Vw48HXYfiKaLr
9T+6FCvsN2sc7DcwEq5FcdOU8afDyx3q5Pg7e5ieEUXB5K4jrKnm4rnA4d7yKzhjfyFrbt6QVqIp
V+FFEcD7NEdJ/cUykHBxCfDlQv2FClUfRbrH5Y4xjv1TktNS7qU8h1Q+jAD4uRvyoT1rQEgXylnb
FciwzMnBcWKyUp/Icrz38xi2KhP0WxPqCZP+W7xNRgdJtxH0U/zZyAhM7Z14G/VpLkGemvK1h3sG
6LN/4wjeL+oLwlndChGOw59k3OAvptXUU2ozPh5F7uBRu3r3tx5b3ENl/m+UK5mgOVZ0Wk6yJlfW
mX3tjbLVIN65nLWe+k/cij10/cLXy/lKskCu32DpBLtBBEY5MJqqHT+g0/vnLt5G8SncfETuk9tX
5kGr+O2gXcz3cGyohBwZl+xdZhJvHwFr0jX8tM1cYWwdF1att/JDZJsxliT41QLCv2dWAtJKtl/k
Tjb+A0SUEu9ADQ5Trk3OzMrpmMBM0LV7e4AbH2mKOeGCGYOr0OM05bPX9grH7B6W2gctkFzl4759
yCsi3CpQFhZciH8VHJ59CtEZbpdfN3C0+MsB7MXBxp3ILzy9y4ICRIqNaUuos/V0GiRiD5Zp64V3
HdPtGwZBcWuWRuuy3VDhxYqyKe5BBYcO2Vc/QrirPrLEPtfFQ4LCwlhqb3Bg4GWhqHSOa68Qdmbg
9EL4ejlKmaVVoIJ6i0bzVF4gyR53S+dqfSsie4XojBTo98Jx05Iz4ksBMAKilhU6yLrgWWdOLITC
pvvLmxwDLq2x+4pQqrNbic8L6znLCXK0i1SzI0Z9MR0HZWix0CRSgBmn5pEJeDaDo15dOXaMMjO9
PfKUIBpHLONxJ7qIKSdLtUphRqk+3Uz9w9hlX6S0beNXa2FXybGXWr3yeYzLQtd6Ma4CU6TPouz9
bs9M7ZUiH+r2uoEMGUoLFWW3//en+kFqFyYPGfJN4TmVcoIXWmRvjSk3cozubsgVyzzNYkFvralR
uG6oqa4EkzbOKNcqnqgdcDDIeWX4It3KHqoKdabIbRJUgNL5khFtASGHJhoIkUBAKEQzSv3qczOG
zZAlbhecjnlbxDWHQl5nrk8LMu8OqUceAL2oVnCfjyhYkAugjpF4dO5o/BSKE8I9TbGJGSNZwTVL
XQfwvBbGu9H43KYhQHXHw9i41h/WHfyeTBONgSahaJ40Z21dYbzGUwiSFdyFNltFg84qnOpAIJ6b
YFLBA9Cy/U31gMfdXB9oMfRgh502IebsGWqA90nBsiQc/7hH5lDiEk1ZQIBFIxxFOpe4Q4ckTT21
nQVBrne5S4nM6ECgOg5qNaBT4FCC4dGoIM2klaSiv+HpUhoGttsZeZkm9FNN1BSYB4XRXri263vP
Eo2q/sxmDleChG1HKxWjvTLxYshMXFecYwE9FoFSIrG/YmiVb5BzlInpUWDaMu2KBzcEFXDajqPR
o5fG6O8HW9c8sIUkRYkiyawTKSajb2qWvghd5PnFohd2U7c1wa49A8rDYQBNTIyjiqY6jINqDK2i
G2lwYJx7KSnSz6XJpoYCFnk4PBi1e9LimzfLgsV/jyB3hNAf3JYR81XILiTVTSzYgvVAQCp6fjCB
uIE/dz3aLCXcN6JbpN0FJvS413jAiKLg1Ok09Egs6XErS/T2wgfAJeQe+g3tzhcSrTlhQmA6HRr/
tJYmoUfGuxTHqU8bywRqG/+YmgGpB5uCVK7ToVKIj0nIY/IwyhLn1B55RY1KasAwbVLw/oKZ2YPa
hYHiMC6wAaaYVfMic73hUjSGYvd6AC0kYNmI2A/n7IYDXT+MNsT04eCE/JZ6EIdZuX7N3pyGeNKu
XSCkhjUkyiyp+zh+LzFnu98l+Dt0P6yHA/S/jO/1DZTBJY3PhrcVpYReTUHG8c20I2MtJ6fzm5HJ
IES5nR+VQzWIJr79K0xZM4AZ4hABkooosSCCYTBo3lzsJ82nUYPGMkdqtFalpWGB0wXx01O+zYPn
pNBAC6hbLJLTpC/7sWP9rkxQ62XaA1UTcdJxWPkhKSOY0CECR6mMb8Ne+SVBNozBRwgWOYcm9WXJ
jcyS2jpOERYZamnfzsPkc0t6oHmrQRHYBvVA2LDZu67bh49+2EOTZiCpP9lIoLZGnQ9r+hr58dQO
hrf+uqFhfEsSn2gT6gbw9lSvLtxTSNVjXYTPO7nYyXyaQR3BsVqfW9syUjAdSmviSVgkRCAV7NPf
qhpacnj/l0H/oCWXUUVR8SybLHkTGudsbYgWzlZafMzz6evcDku5Gz0OhwMGGZ437E2q9pWGNZb9
3CV4MzQvmCnr8tPbEAWdHig3Txv9tB0jJEZHui6N0CIuNXDziMONDQenaJOe+D2pa705Pz9H1iB+
IpDCaJhp1RMNDZIc5+qcwjLIF2H43A5rArKRpd77eGJWt3vMdSkakO3g04Lb+e2qlBngZVO8QpeW
j2W8BbT+qpuhDZKLt7r4LFnFDW9m0mbsCwZhDepsxnxzXdvrDb1blVtIJD9oLnO0XFxx1kl+/U6X
SlHgDWue/ZE44VEwgXIvi7uZfd2SD0v0yUTihCdCjUigzgzBfJdH6SjpBjxnd31HyRh4vSVcgMBM
2uih9fuMKlOoGO5ZdaNZeQywOZLNsYYyBK+wTrADaunLD6oLum48y+oSuU1LpkcYWsxAm2udAeFj
7rgqio/IYpXvVHtBRkDnU0gcHE7S8WmLLNFu97OTKnI/8lneT4/YvjUVTNsdV7JhQgFiwkt4oHdq
s7C2fJ/e6Fc+1Y6KOV5Zs+TCeAEnI1RJxz0wkfqhke/nVNyY2bD8S2Jxh/DtebFWpBH1+wMgh8+J
NhD8NdTd7/9bWx6ZWjsoz6ZZv6ldpD/XNnInaS64bXf9aCcvK4q3AOh8FlqJgMUlUyKrAVVL9c6X
bkZMycRr4cFk/JUoT7D0VRwFo4SxC+rPj69Q+eyTU7G0lf1LvHUlOiZPb6hKu0FwRKCeoWyoi8fT
tdw/aDYAIUvDcF4Mjy0Vkz/iVej19aFHIlH8znHmVHaZ4+PB7YccAwvaD0DmQpi+KzRE0vZ8aW5a
vqQe/7LWlFJbQUkZtbE4PjgnRN7u0rktEHV4g8IWeOs7gkMomvK0I+J5kdKdkviwVZu4hOByi6FT
0wpt1GwBt+FiwpDSSsnk7SzUSE0M8643h17QyXEo49pPhhjCG/UmjP4KKPQd3b50t2qVhD8tTfuk
da96Ds2PZVk3rSvdJ5w1Lv0eix+lFr7VKMWjD61dQtquHwoxKmS7ANrlzeyYuFvoR8zz3BxwmipS
4/WopPB7GuD1vt5wLFwHCfKg753ehEA3bRb4LCszngquQk11b+ZlxK0W5SslonXUcibERHLkoifE
WOHu5QSLa+KDi0NBi+vRjrE3NRQvBIcX/2SuJcATfux/K6mEde22e73JNxNfHG0D8z6rWO/6pm3Q
ek4PylPQMYE4zaQiQdoo6bWIocazllyoC9j29Qc4arkPRXfu4JoFbsfoh9tLXmSE8pYFVb7gtygH
3gyLX2xIBgjnEW/AtCgrESyvuZtHIuIF4ceiQMPzhaCroWPrbOpnCeawJKYxFw89pr6MncsMbo95
PrsRpnFfWh+qtL0aprczqnpMuGXrdvDaxwEoRfYlfF5gPJ2jpemLlVpnQRGK69JAzzdTvrzDbuV/
aZSg6/5WFRG/ezqPTVVkhnLXNRP9zZAB46cXlYHo9R3e3li//Gsd4rbApZwJkIdTpRKaDZa3n8EU
q/EuWpD1BcmIvC12hn6eUElG0I0nSVflrXMREfMsP7AIvlUccWKBrdFOpCQPg9tosyct6DDKRuGk
VSDaPRPil/7Az8ETCRrrhuLPnMNkIVjrLkp7RMcGAGZ6vCF2TzycoGW7/1GIPKOpbWGxV4hyz+wd
VDTL6WtRSXrgsiv77FeN1lEJjvbIBit9gRI/M3+D1C49IieJDAA4AuXtbc55juqZVEvt0fv5VUKB
iBe6VfCI4yXGd0FqDsGnF2h9grJvt4En4qav8ryISIQPjYOpvd9kHtrMqclgRriHqJI/3yr8pAtW
WlrMfVKySeBnP9WMZSzH+jdhitlhAZHK9GAdlJpG0A3GKdiz+ZXhXkuhP/4waSa92XvqOQSphgzs
IL7OYRXuRt0eYWWf2bivMOL6FIxpmBVZCCjfoJe8lj5KhJtLusa6KOlmZ5Z+gp4WlF67eIMOT2fF
N7JqaLWo9Blt6JCHwZt4ldgQMMn6f0g8XpHSeGe7Dj+uMUeHv3O18jv87cycyIqh20kjYfvPBMjf
u74iBqCB867JF5JJ8xz/fBRYDbCo1cQ+xYDuE6mm7BmzOwZjFHPRAAftbCL7hf2bVfh+KpX2EAYe
VZBz90Lk/wqYBIue86JxBGZQPiGgoFhpSZQIu6TXyG6AncjGuajOPUzNsTwfnJvF/voY0lwyiFi0
UmKrxnHlnsPoH0JCp1oGu8TdrT+IoCuMGckQ5FYRYDTY/Nl79GtNS9xHXofokCfhB90pL3HlVodL
ybNhn7rCxHar5Gh5IrrcME6aND6Pe8mI9N0kbSBTfOKYUFMlC0Se9U9ShzGWRjfL5TxRHplT0cwt
GTSjvhQZkLxCpCA3PJDuDsoBYkTDIlC3S0aZQlFB0C1srjWfguIfZd19n/WGlUDWF0blN7GMJ2rN
lU9O1Col+cAJTv26F41qHVyySeKdHQWB6hVyEina+Irkxqb8As/XzrHYQGFLiEZyTgVt2pIxbaK3
5VWCkdYNJ654tnjQRMpWCBo/XeByXFtV6TRREOU338rKIJrkiEDcnO65dXDjkdpHgl6EAb1SsnE+
RDdqRM5k3XzGZK8wh8+Ld5S4dX3zFaOaAH9BiFkO2YGxdFzhjTH9CeRXjhi+MdBG33iFhfK60xUD
yR8gAzZJPL0M5HfpnZ38jWfDipjeTM/qjLos/hAM8Ff6ippw2mrM7tOf0XasrY3zVOOo1ooZxSu/
OuHhda/9eTLrHFsVWNRyfDUZsMKhKLiL7nUcHDIrwUT2mlJeUhSaAvAfIN91YNQjDCjx6XqCvmnx
Y1XGBnae8tBawEwSEN0N3Q7bew8wEpH7i0fALNfOgovwPd3LdAaXT6nMZZoXg9EWO6IyGByNeZPy
noFrkXiEhuWNBW/JRd6mmOcM/CnJKs2TqfsySYONTbbJk6wl0bZDBY0z0Fg1OIyjuuNU9rwSLfJX
jZ0thsuOa6soBI9uwngm76m55pVduTVaVgPiJ7HS+n4yPgpV2xI5KuBpvcLHTuOPCqK4qF/3bHaB
aBiNF7IObHFgsaPOszeQxzacxIgnSlRid4zAcR2ldmrNTdTwkmbahIU6w8hErokdFiU27igObYVB
i7MF3thm9zKOKcIjJIc9NzV5pw1WNKS86VBfnlkcswjL8IbMAleRjs+lPe3WKWwM60q4o1JCPN1T
GY91yWVR1iUvml5Po/e1go/0Z0SZ2W/NddFXBwlmM0qLD2Kr6Lo+4Eqm9tlvcqPHvm8BGuZAg8vM
v5u51nML7ofyYKHuBn1FYDipvmX+FegNssIoIYbricQhS6SMvo0Q0Pmyvll5oKYDx4rNvVfpvISi
5WxeAkAcQlWruMbFbg+hadG14xewrF6c7R8ymkKXbIBrrJUz+GSiv9V8giVNvZZ1SsB9zMG1CdWz
pNAwhywi3nF16H09aYeF1mquVQau/BNBWlWAlbUTyx9lG44YDelQyR1QLcxDW3ix4WSEEzQUX10Q
qmyoUXGS2/5E3rD4mQLw4AvrbNXvuL2mGVShhXAzYcQX7VDmCGE9JRq2j29RUrE66Z24j6hJ1yQ7
2SrBtU04jbGc1ldzims4JdFDQAGhKSKOtAp3YS7gVGRGmVK1vJKB/HLBVvMDJqdMTrXrYtRWn5dA
7yXpkg6X3YByzcDxn5aXnlSott2A+LJX4DiMYsempfT7SXeHJQjoZhJZF6Akq0zmLrCwOl80wQc0
SOtasW2nSMSP8f9s4aGPZQR+pveawAwazwUYrbLHeXZCoJK4dhqRgmD9GmKk0dE40Ae2jDQs2D1r
qaktX3uhK4tqoMutNFKB7Fj+ZT/pC+UbHmO/M0FiQZVCKnRSZnJTYIdHoZUEJfdY3dklfEva8nvG
mF9r9en61VM0AbooXnDkPDfY5P0v7mlk0oe+OJ53NuuSMwlyR3i+wJ6r7/yBOThAIYQxpHtJSu6K
FtQzQKpWNZkIjQ4XMT/GQ7rtt9gio1OQ/L29DPvXBJxoOSC/PmC3sfOoXnThVsLrIWeNHeajR+Py
2YR7TwkBxi4M6Vi/6r28/Eq9S+ZanG7x+Zzj0VRMKcCSbQbFNVys6eNtuT9VBDIWgxWfJeYavdom
BCbhaonYcZry0MClyV+YJQZ/bVvDHfLglbYan3sTSP5wctwUyiR63RASZ8ke9ct74MjyalfnqGPS
/GyK6Gnwt8Nl0i+IMqH+i8JRpnAPn+xMljRZmh7ArpAsw7NYqaXNFPQP55H6BAZacBv8Un65oLDq
gBa5nn5JDBjRRbfPf6iX7X8TDmoA0n/CzK0WwsOuSOHpmMxkhWU3cpJfKVJb37mfPjaOT7Y2k54X
PcxUpBoqkbe+CNa7D+Gkw9h0/HJXMrotdHGsCrulvY8g2DCTcMvePCxuVAzDdSOY0Uc9qNYCP1IQ
EB8ac6O9USFwILB28SFHA2sZ1BJ0e+uRhe6IOx86/PGrB6TOdX/zPqBy+VaBAfbr57w7vEC+pMo/
yzJnyiz41zZZVTUKpjMWKAYtV43DvFIAyY7iO8HIaKkq5qEUhGKhkbYw9O4Lu7LSrYryVz10kymR
yhZX+uDIIL3/eoJwbRnLIFsPhl7D4wxKSR+PNGfFw6qrAkLOJ/BsDw8rsnCVY/T7D6MB3gDF3dv5
A3x8cElTvTSDc5pmH+KU1FjBTtw9NIZ+V/6QgWQ1CRSAiN3Ux4dOmK19NbsgydQZw/pW703H6iGH
qQ+VZz8ylPpRmpZu/RGGvey+wlzhOA1rN3bg4WcPqewWWyAP4J6Msz2jEKJPfaJZT/sVaGTOjRHd
c8nAjVHVzqfAtjPogbKPPdu/9y4T9CXhsUfgE1X191uuhMMBa03uuZ1J7/Ry5b3Lnj6+2DR3iPrn
XCL4uKQBk/2TbaQa3vXm4Z7v3uS1gIc4x2nQDxC2S7VhOObtFENQYVep5plEsa/T25H7Nz1/Honp
okgGV5oW9XxrkdhxldxSn3I+EHP3fknhEgoJ/+1N9spsVZfWcLma9IdPV+V56IVNLN1LqFpg+tk/
VA/KMuCPaLzwfiKo6EIj41q/fUc8jXP+QUMYYkSDS7KEx9cBzzGNMk4Vxorp7+IMikw9I4z+bLLz
JK/0WjM+UQ1/E75xPgtoiPYdHey2QDVFaES3WsosqKXqmsVeWOEWb/HjRpnGH9lWtPmcj/AeZR7f
XkZZBW+zBngs/82A8KfEnlMJJYleVgmKN3vrffny5U5aFIhxhstmEqPSuuR+JDa+gRMZcjrA42Zl
DtgrP6KySQLu0kX0Qn/zmTt5PivmqIkLKHMY5GK9RS9fxdgVOfxx6Q7ZjfWqtI2N7Q+5MucPGnFh
j+HdQbH/ldYbMHAyBojf5XkNCwzVaCKVr/w1Q7nvxCnKQkqijxB1CYiuzkPmS8xleT/TtHiQVpnG
MqxgFu+krw7zIUsnuCjJqTBmuIp2WJAIuouactWJiLOi2ty2fKirQnqm3/vrHQiccQpjnlY3cNJ1
n9Zc7rPHR2kSJ10cFDNhBJ3rp2TEWRXtlxF0Q8CnixJew68RfI6NtqjFTiPv0eO3u2fU1nxcXbsm
ev1qmNK+fvNiN/A00zXuwKpCVDn/v2Pt/8rTArlVy8SW1rXnRrzBq88SAkepJkdieT6UE0o/oWc7
7s55yEBzlWtPQjCkqEFv4ZmA1HFqjsaSVWllwEqI5lJK1vHImEIWEaa6+8AdeATAuYawwlNXq7Zu
SLImeiw93exWTZtiZTSxVxSloHRaivgR+Eb2v9AGEGlpU+/gjFJ0G/4jIBo58g5fysirMLxVkmKq
QiRav/kQjrz7xj/Z+b7d3AqGhdZjkodZebsjIw9k76tSKX1VF4zsAC30CJgIFyzudsAqcJ1L7YYD
MI9E0i1Pp5E+p5UxpKjLu7IBU8NQx9izrknJKbXcjI9s5AA6pXstK0F37sYXCieU4OnlMEkKrt+h
IAOAEluNTSOw8CULRuupV3NIAHiWR53vkewzo8JZYOtpPn3gzYYJ2WHhJXpPIc5KdxtVTqKgvlwd
AY8VZYeFfjOoVj9a3v4rDIUB58GitydNIVaeK5ufU9Aqk/gqE8t0dGYBEsrWcU2iP0933/QE4Ony
gvSMmZYCob+45JY9uVxXVNp6kZK2i5HOC6zXqMMllSWZFEOQJxIjEpztvQHiUXopsA66UyF3/QUt
ZOsy3QF3Z6dUJv88EZ7bcCXSPRm/8O1CUk4/7zFlZRU+ta/0RPEtJ9jJR/qqgU93epeDMXyfapK+
Ki/y79ejLfYHaVMFx+AYEauFYl2Dwm+ev3d+ScsgsBxmSoxk4LTKhmRXhcymkAHDnl2/vBh/GQJy
xvAxpd0voPvy3c4pHKZZrQNmgN21fOBWJPxj/2j9CV+DTEnjqRUTDgu8s7oxuTWBhiKc17pYQmo6
JPdwz9uhB3fsF7HpJ82weM5iq1+o9m0uUTr6BQrZS2g+5qKWNyvWYN+dY3prFPq11tv/+RxAGZsB
2eCRrFT53mCkBTbmrw7eRni2lnx64+ulbfMBGtJVIei0IZ/8wd6/LQo8JoUXkFwTkWTFn9qzm7Fe
H4+5sBY8boywMwqnyFSAlWq0cxy4FeBOLwVzyczj377JLt/KxOxwf79M4RG0CwXrzoC12kp3NjKi
gwTN55lb3SEX6NcjepPsBjwyi4hDNekKXw7k6PCxcuIb181qqXFfNgNJRDsgj35lu0pCM5LIPZYf
LjMfkMasMV1b97se5B3vXYNap0q9I5mvivvOsUG0CSSLm68GX/9FEQect11mLijWshJwb8ZyY/k/
oRvDoigvFgNskoUw5aeNTRqgDlGvsg2fN2qt5+J+neBaY/jCTWodfCzrI7sDNTaGF72U+NJsQQdv
nmNTQC8qP0GpVYbS+HtSP+l7C5AYW2A/+LQ2JNi0FCJRPmrfMYg7QHpbrAjuComqmr0nHvX+zBW5
4eeFp9yG5W7c8yh25Q8YT5bSA01XIrR6/MqxPDpxbGEJ6xTBBhtHxfCHn9ShIzmX2LkNimi8ehZx
MkaAfQW3Gu6WBaQaDd+d/H08XJGsvGN0dvf9Ae8JscnYB6xW6F9Jw15+CjDPNv9MUBrcHjQii4qx
XNYWBNz2f3RQzsnc4EWjeDgzTN8KU10XDpJtXXZjR3ZYs7jQat9p19VptracP4nfUb6xlb7xh9pX
muurBkzZurY9ru/GaDOpJaQzy+4gsFdhtvpU7NIkMY0GSNcJ0X4GaJ4sZ3+w8XGKadFjYhD/W3Aj
Tp6s/blq+lRCuQKvly7iG2uCvT+4Y4Biy6hSIglJ5HQtB1MDObG8eJtgB1cu0DvNAAU3O1zQhFWg
IETu4JwYRWBpRLoGytZh1/sqqMsIGEbUemt2Cmxa7r4VCuqcp7wfzTVFmVMirOBk9x+BlxK11xLI
MrD5spmUup23rjt6z2LxxWPT3YmZa3/Mfnq69mX1gYpqPYLkgngUHjaAWzSfq8/SD56jOlyYzxBe
7d1eqd5Be3/A9C3yrLMB13lHTtCqNLp3mTjAkjVLDgr9kGbczA/nFQoxeczfRKDthg1gJ+ROOFUx
gXFcFniWT7OB0Zb2EIhsI5kOsrObYwwzQIax4HQEezexiREQtjR1u66Uhgh4djimm858adCFXxAp
9WijgfjiOIs8jCw+RoQU2IUHukO6LMTr2Thh2Le+3C79IDrEYfV7blOeMTPfKSAObQpudigVKXd7
lh3hMfrZrTjyLsN9Zp9HM24MVTe38B+eewhn0Gm8o0R51n1tBh1Nuhg5zfy0yNpp6v887GdMXFTq
EGH5mlIZQE6Wh4Ai9i4zXTom9n3j7nTZwoTKMeC2QdGrwk2Y9D/UDvzOJ7VmcpQKQ86AesLbJvvE
9fnKP4zg3Pk4SNhlHt/7HnNj+7RA3SCntNrrqbUicyVOY6HRi9FiW7vu7KYrHKhtGbkSGWLP+TsP
o6uL9VuY34fbQ4e4XO72zI3s+KpoAB+3SNoVWJVKwirYpNb539ou/HhbCpijap2ODlL343nB5Q2W
M3sILPuIq2BKknSQpoRxqgb1/Pj3+DIxsVUuHVQ7f/kniUuu2Au8bkoTT4itKQuA+9NzTlJTMC+2
3YqIc6hEluCskrBCju60cghx94JBSL4k9vWCxUHG9ShlUKKPbb0/YonssmUI+XH/j3Q9T7i9U9iu
gP1oGVCySawBSxhM89UwlL9u6QSQC/UzPWJnFJI++6VBXRVbBd+ZEiOz55pVtubQZ3BXYpMTbNwq
ghq6GE8a3JXbPaQGyXIgceGGg0jDeG+GAhojI13ksFnZjWVqPvyVQYPGSq3ScGvNRiL4wGMpAASB
p4ayHjhp4juveKbtS9YY7CsTWinSb5ccUdLU9S7OIdC/kN0qPBPTWya+g9xZp/Ds9SZ6Nxc4krU6
trul9zMdXMWPSgOUQwA06eY5c8yd+hqosSY7VRY8PBhYrFYUm8oR+U6zhAEo67h9EHWWoREzlwQC
UM3NmP2VMv+of2xbnqw19i7/O+b4S2Qs7u+atEFUuo+6nx17JlD38pZWre37VygmvH9pBmlFiq3c
JRzSLqwRTQhnQB6b/VtQrpJiuPeOLVDIB6aKllLxwle0wrzkxc8g5aB4iq8M9ITvvcpYk2fIsXsI
HQcTLsOj7HCjwIOwBhRDGvZrqh5X1NUviwnCNPjpnWr+haTJFHGFmDHVUGgOuoWdLtmWAG/sTezJ
/qNlfx6ImQdKOkib7vmXxN1d9yuzL5JhydNGKGmoVaNKXisDp9eVh6YqjhPccfl3A1V+KqonjM0j
rwT2dnqqLM1orZeggw8796A/pSFGz1eezdPgJfV0l8ozZzp81ZFI9VYpNjQ6BG8PEF+QbRMI+M5W
LbjcNpMR1o+1SCWPzHajj7cct8WYThKeCwHZWW7ylcalXYkosQxhm7uO60J0Yd92UYF2F+4C8Wzk
oyP4kaIc7WLhZVqzePV2/9Rplzm8bySCP/X/9Z64/76O9ZPjyEjBNJe5T+lqWbjoD4xemvGyaVR4
HFflMdZeHmPftyeAp5aLhtn3OAhpQbu+qzXFM3hlT43rKU37CIw+h3HwG3WcjZU4MlMcyXTPZm+X
1wJ186mYUAJnKmFhJQ0SBNVfIF9wFRxewra4GLcE713AJ/5lpbNNEEVDHLKXWjNsdst9Pz9pjSd4
5xYhncJmE7IJatMaxzkF8Mwt8iBLf7ha0fEJShVeJ34hNr+8f3uaLKCBOMNlxxYjVD/A7AxSq3X8
lAWSaNskAy4lYC3YnNBl/1hH9bOeow2V82K/HmjMHfYP/sAIgriZ7SXwnf2+oTQyVJsnHUkumaY4
K2OPiLni+MkYlxI3lxh56E99d8SVYX6HzfY8175tqrOcVtJE1xGrY5d10qxs5e2xHOAteUoK+HTF
GZdg8sEbiJY4QcqrPMJxpFIUGkOSjy5QW7DpBjjp0pKeZYBLFUDgKFuqvkW2LlRcPBhAyIbD4PMZ
HN1pHHqBXCJSby6Zad9zBPdPKURFatdIVinBNB9pvfTY8deyZp4PFTRQsVsSGE3+JrvN/9yg0AFp
pYJhffODbYjtaDhLxdAUDZhT3jpeYJcYct2MPb4mHurhwIclK576RDYy7yOqVJjCKuRYAOyV/zHa
D4xq/bPHtqd5682Zrq87ozdoE/zzp5ujLYWraph0slwlmZlwFHqS9u+o20+sIBBegDklmfYxu533
iNI4GKzuJ0FxLN5RqWS4EpERkhKVee2QrT/1FPwKA56/hUqKsHalVMsnVilBnxwPZ9HR8HK6fpoI
Hxg2DTQdh58vtJtBPDWvkK/1sLXsCIVRQy9H38JhjUdAJu3m7I6F6oG0iGZC32KawznP8xoR+kgN
Q2tW3IO4AK648ig0m6GNBQ1hUxh7h5GcgTISIi/R7Ws5Q3jWuGTZ0hLLZAJmVtBpSRvBtGweOrlG
S8aS3cJujS74foZiOkkS0fwbf0Cua5ytXxFEM2tW5iLQv6wpVtGARl+WjxKH60vTlvWn61AnQSzU
D8f6cNMekZLLjFfHjACt+72Eej6alTFVU8eUlnn/UvGPOGD9/YDUs1STPe4EJzsM0sGBubXS/gEe
7Bj/eZE6RuHNFCZCIEUi1NrVElhr70Jy6K2hri+5RecH7Spf1niuvwuTC55gPFzY8LNk+P1VBN8q
soGk5YSRo18Ro4AAsqRDAmhyapz/lsptxKH8NI5B9p5uqzRcDMA/2Ztbas+xmDkrPoh/Aw4vLewn
Da5pW31+lvHM2J0SKhMC9fhg3WavE0/QJj108q8z81ifJHu2pfq7+YfX41SLJBBzw111rOs9W6eq
8qjk/bOpph36xAP0N4IOG2ekLJaL+VUFxIJ9/zfBo3vpXZSG/78cewAtIEh7IUHWzyd0+0bKhC3v
AWUmo3u3eDOT76D/X+e3Wi57ikpL86rEwlKNrN6XN71D17/rEkRpqpBm5CcMwnoDUl92nI0lYTRs
EIFFupzL/TmoOT9UrtpZfSwmEF79MKLnpnrtg4JqRm59ZIkme6zLVuhwJhtzLKtj8QSGgIDPsnKL
8EKloK18pFpkL4rZd0/IwLFtHn7j22Mwth2iY/h3D+NWiNYAD+1WAXerFefIGmGnMj5S4yaMD+lg
Gcn4jhdOJbKfrvyRTSOyQGP0nPs0VE2Sbw0BSE9oRCFCv98yD20OUQ8k3ctQLc/732h7i2yR6Sgt
fIpSdDRRWaWoumkOyC4Z2UXhGN+1c556cKNY7EC31s9ozDfePFinv4kf69xUyg9K2WJHWKelZEQr
80YytNWbWNp2D/wP/XpJEhnbQ69xEaWBPN2df3URQVi3C9TomlKJTd7t5N5SeUS18ZzKlF9Uzqy/
m3jbfuuUr9MuXL5jO4348hefOo1AAK0W/RPmni27D5LyjOw4b1ZG/TeR+yammQqcayBD/i1DPY/S
+sM4cmeJ7weZdtweXvTQLbgRYHPE2cOHMluhTFcUQaauh9IyPjVc548RfheXNPYa602QJXtN0CrT
KXOyOc9d5F4ghPoJ6f9gQcpOvg60i6yCTrPera7o1FQaxp6K3XIFzsQ187ppVt/3+1NIWBDqI6Kg
HuG9G1kwShL6W4Z7AMDZLYCjVo34IMXCH7ZHKfSlOvsA658uTD2B4IxeNCaFNsa0y5+cd0zdV0Fe
F8lAURZr/M1TD847BsDu54BXoJlbAVmVhXAJRx9yMG49o5gJnTCJJiBmj2RXCXum6sRQkfWboCvU
SzmGCfVV8A/FlnIeLb6y59+l5WLcE/mIl5SXRdwLqwzTp+9U19mUCQs14AeFlboVD9v7Bi4TVMqg
4THo5Li+duGXqyQXZjMfGCsZxxRbKVaRr5UPpdm0z7Bo2avIRQ1/pZEtivyyG+pU2ucau2HRjnjf
LcMg/PttM9fHHzi/+43KUTr9yQ6Gh7zmMx+heufyKZy8hOA1fVP3CRyDyRDyT9zx/j5ty9I0d9bB
kclXaCuIuhkOvDbfJgPQpIWvaJVxDeJdJuH37p382sRzqqQskcowL1McFkzRR3SqOliuWzySOKgP
fVlBbOM2Kg6dWQgFGqHjqyDeuSOj3GPl417EtINn65va2XlCO/xcD3yjEtKxaQ/8nKgPvhpBffXd
oevH8kr7ehQmwpxuF54sL5uswvlSXA1UVdnqc85+XVCrlmLi/aaKjbEXtoPykgjbRan2nS58tq2q
ZRyVdE8W31l2aReRSHdf06nDXeBGWair7/BGYSMb1IyoDDwXbOF+4nkwOEhrMjnkYtoRfLczhJpD
9i/wa+qG4IIy3qUdzassxaVaRorZaMQeLZ++qFP+wCDwFAyp8/4vEr3ODZ/ptEtamQ0iLncV4CCt
0fyja7PmbtoNzb9qepTJIejtNNByakkszksIxlur8hpqmNztgIQcKITWFSr+8XGJjKRitxs/ewiS
Y5GFVOm+jpL+VGpG9obvCmJBTn/OA750iXFkZV04sTMWr/B06qkn6P1Gu/SiYkQs40wOk3h45nhT
njF67BotrhFaUFnmuM5OECPV2oWorXA5jkvl0DqtAH+TViXk27P58mowR8pFTMYQUPzYL9jXtgOe
m3ak+9JcyOvTY9XPyMAtqCU/3+1fEWX9beYZZFiqba8kfsqLMruJemTJBkK5RydFKyZgruwXKjEa
uIikYc/UkpHp+Y6lu6wgwPRo3i8UAb6/PHvE/PuP7qzSACZNXvGeFrBK9CcKpHu9jEETBxRIFWu+
BDGoQv+2uXk7qHmLPDASfMcvRWEPTE5zarS1Wk5TT0EBaBL6EQcIjSOMywHsCQ32Blo2tRa1eNh8
jh8RP4C31wFw/5xurQil2Ompv+WZYGPnkhX2vlS7saz2ZPqp3R7OFyaam0NopElGDoSOTG9qnPoL
iitue/i5NvARhHKOT0B10+lnG+9gDItQA6j2eqKLwCXD232F0YgIwrNlICgBsnAOwAhFA60vryJs
k31bcpqnzpThAHjg4KE+rEq6CfjQwnoEwJSDmzHXGTyyotodVoYjc7q4rf8k9Bm8NoWC4gKeVtzJ
XfB6ZG6A+7J1E06To/Q446i3ktb/Eyg3SLaWSOwRX2CLoavbVyi4RpC2zNsNrARFbXv6I43Lw+pJ
MTnElcRpe5LKvd8yJABPKVN6ldhqxXzeCt68yAaj8v6TFiY3LxwyepDoRZEL30McQJUTqGVjVNsZ
4WvYhyRr4237jdp9HpY9/HKanLjoX0WNvH8SvH+AZnWCx90D1KcDl4xLhTXDxfRT/hvvLOzgIChN
HlMxDMA1IbvKJBULj0kTgTXoO0KDF/LrbVgEbpdGVaqTkWPrrq7iWiTZwpmfFqsYFTgusY7eSVL0
Jhn2DXcaLKEK3PSV3A+S8KMsriurrxSCKAg2NxUHbSuCR5SM2ujtcCNWWVGTQKYIeWskiUMKKtG8
ltC4g3ETVfTUAvMKHYejNtNrgvK1qmWJu17Ewo9ZdG+PQw82k/YEeF+qhwnt81vyOuA1cbO8ulYz
YWFwrNhhM521O1IcWCXDHB3bOHap+LxC4a4265ArWB+g4UY0h5rH2dquSvq3ofLgOydnSj0o3oNu
6B4UiTVJdYPFfJPe/w5ZHHhLAi1N3cwmsBhAI1/Z6Gumj8pFKFvF8c9OlEFVIEyz08CPLVWL8qE0
jg3sIeDItJyWgkKSUNaZGsZVBQUs4H1e2Kw0sMIVumG/mDuEHc09+5h1+TkUReYr7Jn2hDihG7bf
cBiM6so04BtVuEh83Da5zG0ILzKSEpDpI2qXLbzWm282surPIuuAboILMi6Y26vWTU8CAaukaWJO
fgRfoMldIhqkB2HJUqfmg7UvYQO0up8vZhkIZwALoZusr0ifNIwsXlCe5Ogxlpa6JNur+CBfs242
875xNT932LWt2i8CegMjRojeat1sYA9vSQs+QD8Arfv+F9AYwxA8176jhT+NyLQTn38IV6EtvwHV
bYV/rdRy11XIcy1kSuqW5gMtG7nrlyTGL/ptj31g1esNxHV7tB0V198Nou1lwj/jB3yVng5u0Cwp
O2WB9OfN3KVXacCzZZ8ti664Cc0ui9dwMJYygsgCTnFI/9mMINCBCDsuVNwfmLYeckJR6Y0jCDV2
FwRJLbjj0rIECBrFNk8BywzwpBW396KOFjwZJZsmA8mLeOwtJeuddhdiTWYH1xTrq061d4vRves/
SH9dy22yM5qtKlqGAqbLgK1KO+xObMq4zyc6IygLWb15ekx1zyUKP+u/od1c3/kdb0Iswgx8RyUR
7sbLsrBNCi19dPFEHb6rO/81VbajJadIR/fhDwK9I40uOVLUVFmx79zNMNqU5Amtou0ho9qEkAqD
d5xy24yy2/z3RvytkC8AmDNINwov97sF2UFAwyNgTXcHXDEto8t4LXlmPQ6jSQ7dm5vwtPy/vGpx
8cQd8fpTcwGlepeio7jQEJW/r9RNKh6v4vWTw7/7NVvLvTCSH72edfPZyE8LhSvBhe1so9ZY+387
tPGfYM4VRcl/0fPrYHfPe7KKk8zQPQfU1UX3Cn5bcfhjuKsVoRdWigE3gATc5m5o2kxGwveEFuM5
VpMv6A1GrGn6oH9dCAwen8Q9SEfB/Pkis39E32bL2y1B7ALyRyaVmpoPLMgYuHB3RAX1veykcIsk
lvco+mHMcXg9lYW9dqEmmnWBdZ1nnt/jO2cuVEnYJ9hsmkf4xNLuxK/iydOEHzVKJdeWQCc3N8f/
mSUPMiLxTgI1W4gIMKTQdPGJDpo2IUoPs7fyRU+s1rjorqeWVX+CAPs3rvSq/sOuYYw6ZKFG0jsI
kpyvUyfSHQ7x8+dSnI0CmnOFoCfkGH9UtaDu/WJU/658ozMOrefgCAb0AvF52Ndg0QDXvEaFNNmK
jeX4a2dpBGmjIZ32YvVpIbCegWntzNGD8ZVrsOeIBBWCv6XRbOnW4cgB08JtgXiFNUO28EWWGgjj
YlKsSGLlIgu/QhnS9/2XTMBvVkOS1gM3Cf/AeaAHkzZqza2TY+S/bIxCdgLr5uVxfF1+mGyN98MX
DCpxJKk8CfIBiFJQCfFjxNe5ogxLgNng3+zGo15hjIpkU+raFvgW7/tmCa7EMTtYICo5llmi9/+j
MSXrMcQWoGIOUdbhRgFaJAK11eGq/8sqXg/DS7rol1uqOqrLPgLiuiREZEhLnCyineDLPh/3qP3t
PASEBiaSnpTCatWwqjHHqDb72hWh6/LngfwRF99pRp7WxkuvsIP36oKHghgeT67bSysAkU72913x
xDCTBuMWF1CXizK076YkzL/oOB4HPeI1rtYISWLnCfuuHOXXCgcM+xHOXiH2B0Vf/eGZxUu2rxiA
YaoPcb+o/jG8cgmmBMnl9TgU5caKgXTqFYq69n0qNbiEUv78q+/L0V8hmaAsY7QNMKdJLS1599Wg
jgv0AjF94VhARHk/DuRDvGq/AlPltOddxfXujPYBlg0DV6Be+mu+HpTaZJEJep/Nmf24+01M+8Tp
5ZHTZCSjNExteQq451+LmpJdlY4NJPL1C7A3RQHkRUf0nERr/riFC1+2YwgmH/ipeAU1T9ifAEAE
SZoShZDRDjqhupJHe5W1jnFOMFKKlTiwtVMNfrF9PIeJjKLyvTd6cHvDg/LaN60Zfe5icrRBNj6/
HskJ7mR3bp5/LUEemrQ8KnxS86WeAdnFBtIffTScoz2gQE2ErMvIhnY2zZIpSvUnw6iI2eEGANOS
NBfSjcTBjM2z4IZYsyRjKjBcvY5l7jdyW6XZd6Ey2Q7JmWBt89Yhrl2AW54pzA0bOVcn3PY2m3XK
ZjApGHNgR61CjWBvcKaDH97lBby58gYAfmyHhklODVPRTi+vDzaegXRi1yfrnINnUJs0ozzNbC6r
+5Hi7ZjSe0ksleQV5zzeg8tQLwtYZb+eByBbXUQ6Y6lbUiwk6pxcBcG8bCqFA7phPvSRprwSW/PG
ejyWCdaZYBzc1Vx9UrBBB7EsACYTRVcSon0CraqraZZJ40AA8BFWC6oQQDI2AefmjKt8wCLNuCIW
IoPqIkyNrce9ukKy+2FOwh0L1A8M73pM5+XHGjLTHhVf5tsmtG+fPG6eaE8xVrNcaw114DSpOrMQ
+UaezOAc08lDR9FvvLAl4isfmC3L5lYZbdFTxCHFTWumYcyHTOD4GI5qVr1l0ZjDsHSoWSkjDpfH
8JCbX770K16aSf4hXTExURfJ0mF5wmLgyzFoW7VRE8mjq4VVFWd1/N4S8l330xiCR3n09r2l75LO
qj4+LX/htIQY6PgffVQMx1XlIR1JC+b859seX0wA1wHJrpLb9enL2b5y380j3CKwaw+lO3eMyaMK
0dSJ6Rv//RbQnrZFaPYJ67UffADifkK9WkQcXiXQHYAC6lxVg+di5DN8ETw79rHA14uR+3bBcptG
Yru9VvTtZOxpaQdgkq9a9KYv+7/Hl+0Q7CVvu0F5VSZd4RyJP4gFd6S9UrWiGin3OypajxeF9ISz
eW5eMTc1eJUG1VC48rJRh7ik3iCG/U2mN0amFwNtn/ni+hCWLVbDJVTS02lWfGtYpM6hv99utSVT
4sC/HAdkY3eSqqSyeimNG769ryiuVhSLnsEw2ktnUY38mPs12Z/AeCVWyXW31QgxFPMn4rgwW0Tw
o1j6uEkSRInO5ZmcgRUu665zww3QQ3TSXcJmFMEFpYpL3haAB/lI4ndHd8OgEjJSbRq5pWgXCynn
wR7MHOthxEAwH7w4wk4zyFdNqNaY2NJzaG9Mct6yEVepOyFIgD8+eaMXxkJfOwvSHEr0GdVw6ClL
HEJLXxdHy+fvd2NQiNn/8SuiVKzjPzctf0/WIXx2TxySlad4Fc7SSqE8OSgVByJA9S9H1eXCcAmM
kXy1wfw1e5bEOtCYTwYXuAO4YYsnsDcbjix+wDgvEd6LZwHqCIuGipikgxW1IDEB/vrNZC7W/OPg
YrsvFB7DKhEpyNTIMiDGEseFJX1FgbFpxY3hUeuUfalIqT34y+CmpjqGQpXPMu2O1Z3TLrKsDewB
f3C5+1nVYC06tov2ZDDrQPLPWC/PMafAft6a9H37SG2nsf/kozhmL61mscS9QbtgESJgqUc7OEZJ
iiryMpnj/0TOK14JpZkkoX0ehwrihFwUL6ljNpFc76fDILYjDNe2hUwcl7YwWgE/GGTz6a4UMzHn
f62demppKGplH229KF502Hqw+PjgIqdOA5/B9umnDCWYVgozJ6trOhIqvPyEo9lm0YJTacckJOE5
TD/BMWNqQjvIYNqhoz+b5Eo/Lo1SBpKjvBhsCJASzIBb0BJ44v+m8NTf6QeRmrmOJZc4/0/Lpgue
/Pkth/Lm1HDiCqLrUbIDgO61SLKhggfnmy09nualbvVpkq9Mu7kcWP+hwNO+i9YFv7ewuff0lDHa
WRAPg7gAE9Mg31n/9M60JGfhGrtV72JxWCjMerDAOm/KC+NPmTp3HbHzszXi+m91tH6FvzgCi4DT
a3o9cwPC+zRMrScsIV2ZWYX1WKAnOY8WutmAfzEQNY8MUsRCePYFEdyuzvEvFjUIMV0bEU7cvHtT
UAdgwOrhn40Ypih4w50KCAkhB4+K+PrypDFMzh5NzrqXZBtyJ0gd+9zHzakPkIk9+LikXWs8VZ9j
tLOgARt73NKK6cC9/KMXesN6jlNRTJ9DLfKyA4FTL/fbBosALYxRb5OK3HqLTZ6G4MvuG3bXvGSG
kvU4XbksKxqwrNByvsLljerAT3fChLNb5OLkmml6wgJWk83my3Rbrx0ZaHuixnsRAAkt+ac9P3Dg
wm5cJ55VcEa85gR1ARNZ17r5B2q7K2mUFGlMbqOcI8UwCcUpVKJ9mt6NnnCdDeiRppN4Q4g4N4zR
pbghgwVm52/ZT2DGs6yVMraQGSpJwTzS/57/sSSJUpQ+kWSmP3Z1MrJqW0He6H2yCZyJt2akzMVX
iZV6SWZ7NTKKMMOiy3Ki6gwls0s/7LAdMwXqsZm9QQuOPz8SPzKeM50XhM4pKbGSjvWo4kOMiWth
RL7Hxjmttqy25pukdtUEDlvvaTfV7e+LayLJrJSMzygCO9aSh48Y3nIxkThTfNDsFtjO9X88PvWM
s6nMGlEhR9CLc/IqX4gFNp8oww/MH1/Uwaa0Okye8Jt7FS7lgPjW1ceTglbu7r3qBF75nqMMw06y
ikJZnY7tDiWi3iRrxRCNXVXZrrLT3EWU7lirOqyDNFOmtsJZISETUzcugGZyY4uJy+c5TgXg+mnj
PGBLpuHLI5fNSdCb37BCzp0eZLP1Qo6jjjJSOHlnp58s0BO+83bWUl8OKyiafKSci6prcnTs7ddQ
OiOtjN8BV3K8buPkzsYQ9xea5PWxbh2OVnB/w/iomMcLInd75OCyp8hiy0AxqjNsCkZstD8o+p68
tvdYwOlXPM+5oBXZ1CFMrMmc2OMXrk30g6tNSQf210Yc78wh0ZF0wj3RzfadGxTOqZzJgt1iCFHb
QhC7Yh3nu8/MW8LnNkmb6ZqfSHXBl8UNXGaHwvUNY1dwag4VvVDcCvCst6ChJnMNKPRzNsIeg7sv
a/ydNtpKCB4oivFplXDU1wnMmKmXQS+u+U8SFoSCksH6+SQ1qz9xAuqcJp2uerpMIcNodd6InYTx
Y3aQbge1RTdvc9sWPUFHWv7k5xT0XndNeIk5iIF6t283RPaDyAuj9/zIg8Yvzy1Y44i1P08BEj/1
iGvilD/CsnFvnaTwaTinKKJG6Poc7JVRUmd/OWTKMqD48W0TEbXLqXnQ77sujcxkB9vjokZFZH3N
j1G0tFBgjrHmh8kQqHWVTQjoqhNl3tQrv0xFdo+HRv+2F7+4JbS+XeEov2mgKDOql5qy/mwM/y32
1Mz4m9ABdbmz69NVHjK7dGhFj0odzg3ZxsLgIha0lnxTm8PZpJAoXbYR4HZ/Ywv+cQDWc1XwlJo+
VYqbZVPI2AMB9vs1RNoz6rQekzRI4QMZJ5gPqJfnzvlZKluo7kU2D11+KtAYUDTuPPyuvBARB3I0
v5dNpFe3CejQ6N0HnwefPKmANlEyigRO5wEU1iJuTirMPqFe4BpmUX2ys+qzKA4jl/h+DbEbqZEO
Jyk2IXLwaQWXzWzxWIng1X8bI7FfiehzSOm6bEdgMIckhVkNGBkP/iJybHN1IY4seS7v/KKVviNp
sKqtKrjUN7xi5UTl5gcoZma0exkIPOFInl6aZUjNimmUJr+6wOM5iBt3/XElDuK9Fc3kDiK8+hTi
DGI4yav1pK+EksEgEWbdKs3eU1mPVNEp8a0t2Ppy2fFTFMeyZUEnuVOU/d2HXKqysM4qHpo4HgB4
RGK9Rd/qP8kGGrwz2CTyB0GeYY4lSecmY1js5wnYu/vHBRAeFO7JvGSuQv2ZuJlQW1xrhzLY/DQ9
4FLDP/nzhe7iNv6yTuKS1UTdIof85MqTzFVNTmCYJdjU8fcYRSxd3hHqDdEtG7WwJG+DwR2ozTUC
Jw3DAyEsvUePQpiMdch3PG+6eYtYoaejV2Pv2/WmXrwmDRG02SDaDZ8Gd177Zk/7dd4ZhDV68jap
GfqNPPySrYU/OS3ZLYU9I5K9Zft30inqoWD1YlkeJTBuRahwi25uMKaJS66caZdxhmlCSmJFjQlE
pPIlQ+KNv55fCoFUOTVOldJM8VQw4hGIu0A7ojqY6o6Me0301R2OD4egniGYp2lkWnRkgE1tG157
GK5AuttZ9pe7nr1q6nywvZyCE5vl5qsfxptyCykYboszs2FRW608ym5GPFAII7wlSWXRLi0566ZI
WauIoPVtljCz5KITCLAcQlcJ0LwyFnOikw3CGNqELMvqfum60MHyCHV9eE6cBVCFF2SRSaddCd3h
/gpmc5y5LUie9FpSEzHIyCceU5ogiW/j6ZCyeZDOXBEEQ4k40y6kHstSUrqDBww2zDeOePGppuEk
u9CoOxFXVa7v3CJWAlNT9ucsKNeR8W2/qfmFLryStuZqE9cqEyenrnOzN3jPzs7jH5PJc3XOUL+9
jBMPR4E0oENsFv+3/RvUPxqf/kAUeuAU6GGn4EzOzrWUKnqx7ShDu6vIs7lWKe9YsP8sqOHItD9N
5FIzt4Np9Q3Y9GOH9W0kNu4MovnRLzYjOnmRIvSnQ40lKnL6HjNmDGmrR6taKuO1Jv7s9Xk6yAdz
sLfCxmSZcGofcZvm+g75J3izvmmzuefWeKtQGh1Gy3hi/kO/0Zwow0ZQ5FgwYbPEDhfqC66Vy6v4
OFupVeTID8SCWVe5BpM9GpWFi+CGKgV6G3DuBGbvcppJ7a2ekrxNTP5Gpp06wp4PK2IiR7hmOceN
bdL6xFJcnYo8ebce3T1kQrdW5CyiFRrQ34x9xFZtSa7OiJoZJG7mqe9sd2HVgrPwY19hoOUQs7BM
gOoDb3vahMRRzbTx1hbPlu5EKdTW/rk87m0dOt+LNteSpwoFmL9ZDsI9UbNfVbQHX5m25ZwQ2+Ou
rMUFU/7dHS4UakPazU5AvfL3GTLyhbazmX17H6nIUTgxIVm78Ig8MQrDZVRpYCAca3Wc+8Ow93ji
FmQ1g9iCj1/aj9EPI5MUsHD8F6hNMwU8XOYgkllRSd+cAsuVV8FWQzktBUhgflweUj7pzenxsnuR
NYUYycr9V3+JmK9cUpvS8QbyxI/D/t8KTp/K590mLfjOY1U9FkFNeiqSw5WKZpd0QFSehdPxItWu
bGcR8mzYRF0gGKS/FGi4TYmskYTq3nM7Qk0ikudNo5lXf/8nl111+yxu9pe6mtSmofo2C3fekiOY
mbVoStfJP4S5raZx/WHa1elF+J6SE7qCLB+VJsOhPrI8w2Fqr29e9RokS4brbja+r3ZMs33FPNVp
vGnPIPzOueO5oOSqeYTgGEX012yUWft8oYJqS37+mX0ypvJtc7Q4CSLTs7KtU93+8M06XQFk4Wt0
WOMUPbtbfVchF3kgvTIUs6j6yjNftfhhoYcKoPxieKPerwhGSkFHeRWLYPbXA63xioumXOr65mkc
m07euPW9wphqSmpUsGXcr2nU7+w1ZEaO01y2La9KjMcaQyZhSfQO2IBzN2PJ+YbguELCpAyC+uSp
ii5vdED5eFev6WnDswpeXNMBVsp9WDCbvkc8M08MTn71fN9WM5ibzB3fyuMfO5EeDrmjWfCr6VfV
8fZzcRSr2mqLCodw7iIyzBerbpcKC8Xxr8PuUxgJFEDkNa1m7YWB216subxf3Pv4DKHtwespDLmS
XL/qaY429BobTrFM2XV0H6FhrcXYt3nLxDOaCu4olDQKrcbpm7faG3TfG/i6N9BSbkPT7E4sXF35
497ftom6IjB5dfZFNiKYSm23fC8dyQ2tjOcgXdYUazT3MMgiPMiIglnKRe4N9gzxWmblnpIwNDtb
WLYpVicO3WtXcYe9zHduNe8bF2lfFE+RqFOeqxSVTLOX3eoiGNlG/kokMatyqinqs8YjC2No23/r
gk67ELsgqmGyk3Dbkt15+HNxAVM+TudGPdL+KJWt8gSD1icH0b9n3fXX1300/LRfwz34ityXidSK
SP7TnypBjwMgbXPUIa67TKm0bzAAEDwp/SGT/V7bTnS9m9uPt70m86OCjSZzTyYbdM6rTybbjCLN
seNNF8X147W/I1Z60dpf1sSoWG9FsRIPLsBp6AgRTSTMJc+vfBPI36MSdshxQRniiOse6/99TbMl
J617rO32rf931HlnZVGfEpDgthpbJ7KDuYR3HFyHNjvEX5OWghCSB2604Qk5hhN3gXZtjOQ9W1jc
HZrResS3g4vjKcQIxBwkZdnzG3vF0iBtHYJqY2oS0yODwu+jwwxjXka4zwlKqiXNaQZG6s+xudT1
pSqZ7s4np6SEKcttuTpWw+cNASDQNYauy9QFUEqwjqUo6odWFiCVgyuuuhwwuGSyqA4hRbKZ7Xq9
GpgFzhBDEtO7ttHs5W8vIvVeae80nUfEpOdQC2ZbXl62xIxjoOGOEE98i3hHv3pHWXbHWwjNVCHv
AuDntDlM1aYyXTuqS38sKWvW67MLgXd6+aq6eJ4lw/HgGgIcwAgMgSL+bD67spbzRuiA6Be6+XZQ
J/t0va0nVXqXfPeZ8y4e46G2l5eEYIHZAlSXJAPoRVi5wi//RnDCJLEOIQACOS0cX4efo4lBHXvl
6rEMs/KYJCbCy5TIbEW9G2SHFNMfDyN7X/wc2PYno8KKxt6KRJl1L24zpAB0wAkXaa24FKKJOAse
zCy0/byqdyAQaLMlPVPHMfx0fscYpH1iuQcfurcoc45WyIxUDwgmzgYDf0WiHEez7UwrwHk0o5Wd
0k2YNfDI2wjBwuzntLx/1fcI5YB1U0a6to5KlV9gtBfzChBWcGkNdRfDQgpmcUeWc7J5yu/l5bCX
irxrkZgj6oO1SSMVEe3nrpa4q2qYujSwvG513CE5YtlQf9UuHDIsoVwPLiWbAhCXpmqhFKGWxMXX
wSSfcudQ1OTZp0HhQ9ylESqzTrL2oc9agjSHxty4CBb7rc+RHbaXaoNOQftdtv77JvGd5ThuPF1j
vpJ6PVqBL0fvUKogElPuqY/HMANgTKPcA7Zu/z/LqK2DGe8Ys9xIrp2wj5R+gqp0xH9MRUnStYSs
Qv3jIlh/yQPf87qLd1EqMdXauBwJL7dEfdPn69lK/TBnOYqjfB+ezhek+i7cY7B+aXdZ3gQgZbHf
DNio09yezAJdHRz66NicGVPoZjwnGxHDMYAl3AxRrPjVRNw2UKP/qCuxeagyI87lSr/JkgmOWuTa
mVAA+VWIe4e7wX6sRl+RT9xRJeBDSenmsD2guOGL5Rpev2yyvk+QVlmyHkRaKEFrrB6oDCpkMyIA
vWnXowiIeE1dOjtJeEbl6LOB6QoBWU+ufgffUMR52Czm5+1mArtei5Ad6k6PSuSmKhWD0OR09RVw
Zt3gwvYTwAVytVGBojZNJkoNaS/10Iwo6qHKnSQJ1HgJ3OUys0VqeNqxSkqmaEww4ilwrtz/8IgD
YKBMAVgDZ0m/RtEde2GxvCAemGN8MtzzcNaDDei03bje9EBG/vAfuL9ueN/lAAbihNUz1D7r/2fX
J88K7/RaME6N8b8elLPfOG6mQ0uDZWCNT60Hpl+9waFToxf3zRKzQ5m0UziwOHnx5s7yOHlaWBXf
+bkhVYOAL6erks94uczASMmxy61kq5unL5AmVQOxOkTrN/T56re/wV19qTZgjj87HL/W98qab5Si
1zV3nURFqi7RqFpWG+L2Qk/gcJp3bGMT90kvqHmxO2/5R0Ce+PWLEueNmyslXZu5rWokYZaiBJAK
od132mnJBEypWaB5xST2Z2TrptiIWWtt3e8km2JVMr71khUi1woLnoyOLS7hVWFqkxiswHSC4MsL
O1f1jAurhA0LZOCHWTIo4sCg/wYgNMOa6zmdpH4qSk5bXXnZmxyE7q/EzIL8ql6XwjH3Op9kOL+E
8fY8EsZ6o2AmSvVXRJ50Pulz5JeXaVzo/lUbM4qXcX+S4xVG1WMv0XtM+cKEdRLxVEoaHpE+X4oF
L5DBS5wfkYuZXj0pf72NGHxLsRfxCRIg1R2iBBrH+heRFSp16mTbrqpEdkwfVzZV/LJEshaJwtwy
Z2C5m76EaxFJKPla4z3P/Dsx+Ab2wJDZcO6aXj7DaspI8O/5kTCstEgXirFpL7f7mT24ueBAlzGt
iC1xPrNGW1Rvq2RK4OoQXZuJ1EIjIyAf6TrokLZse64RYVBDXLrUSY4ViL2liSS9+ydBEUsQSVbQ
SEd0EYwD1ofUsVYug2L61STxjM7d5t6RSkC8VB8fki92ptRRQWmUp6Sz9GzC4FcjW2rJ/JJrUfOm
k13uDdBmIcgyw5bNmJxkTL45Jt4Fr88BCtwRTRSwRgVYBlLBlAGk7mnSrAupb0c2mcKBCG0FB2ac
KTJYBpO+3U0eXs/8StgfbuF8+G8szfO2Z691aJwC16wky6KTB5PKh6RYK1jaJxXDkf8JbeYUzINT
np7pCiSJhqg9hC2au26Rc9pVr0rUdhzXNwEc/uX6jXlXJgFE0i6Mamd8FZ5HZFMCVEi+SRu7yvzY
eaXhRNQ1tnVV1ajJLezoWLPoXCEsbmPOj1wUbC06mlFx/3RNMIQkrmf8UisQdWgej4HpDa3eLjwx
rjMdJc3RGaicMfnxo8fOI4lYB9jJXiwoCkhXzqMQnBpIGdH6bds+ei5s9Fo5alf5bCPs2apqrWj4
CioBTvelaAsc1WEv6Dv13X4/tGCjEFjiXNsarwQN61PBVSV+DMBH/i+qguIcXSXRdAVm4Zl7uf0r
Zr399A2y01ZGAefFaNoxGblGdLjMv1u8kUkZs+tq5qWrAzONFAqVUjSSzSfr8g9uxPIRLKInA3kT
sU1eisg7AmDwG4R6QigknoGrhhMmDyfxBI/Cpj6oLhYzOLia6v5k8W+5IMZGQfqzwFC0pb45fvtD
UEO7jObILnpiUQFZZNTLD8QSYyE/Z3rkfX6xPoQzumATZkQVUiOcfMAdSEDqTAItaWwxvi3fCxPT
mnoN1OxnfCHNphKyAX/GaiEnM/Ol0Dezsh/ZvZdvhIgkMX1nhrVISGmDqYaErQ0X/sNSxgPrp8Vu
mFlAzXNISsYDdciObMEUaqJ0hTRLJ9WFFSiL4URF8fBAkinVK6GRA//IfSiQlocgDLKhHbuHb9yt
LDx3KmTe1/q9nuankqNJpU9e/5EUXRPFY0z0SzGif/jWbHLABQqszzrgctM/cGbznYOGDUdL7dEv
WTRH6Dbaj5QMcVSHVnVG793NHwXoB2Kj2C03F4K8kZ4WOq50EYQ31okG5CC+juBQg8Mrzx6mnSp8
K3KJehNemNaRxyRNNwLtDqMqgIUd3f9O69JHHGy+8jj0bzMjmriQqGTrXyDIUaGkdaW1gbqGIb6e
lbqisTFT8Tjz7mLmDx4Cc96KdY5mWM8PuZyaj2URS+rGwCCgftQCSRA6t7t7F29k2WvkzvTEcv17
clYioo+AwsEI7fl+K62QwTsx+m59+rtwUEsLKgEsAMYhFAMXiAO9l1HFEfZ04F2YlXQ9JWIVr3oy
vi340EUi5MjjKfVBwmiOyBY6DwdO6biAPTD/yWERHoUZYSdALgiE84gC664Y4zvPwVcr7fw4GLCa
ASNr+PcSiyfFmOAf0kf9HO5hl3+fzT7TjDbDaIOwSA5s1p0zEtzPGgEuys+LIgicTLo7xXvsiAGm
q+SLK6k9HXVbHPU723QnKzpDzMR95gofm+PmjmEBKUsyC6jPZHIvbLwPDFqhEHuNAZ7qlaTw+44j
3BINuSYEQhjBLlVFmQJnr76W7jUlqshXiMQ1li/QNkNtZVlRrnqApbZgk0vosmCPxpW8/Rti4kLQ
vu+PIdDFMa8HqOi+43FHvzPhTKIFmDeplUWCORTg0AJZs+AjPwzxL9LUn1VW4JV3iRKrjYqJAwQx
5P/umQ2/5aFVlMhlOIgrFe6A8F1tkRqREFiDPPI8hTmml/k/ztEaTJ/DozRjhAlkyK0/ttzdZAQN
IZcG/IfCiZGVE362EwJnQHFrjefnJarlLkTpsPEVUQwJW2kCZuWuII2mbknNhF07WW+LcVz8oLL0
MO6lCZX/hxyfsfObDiSU+qUy50u/gExTW3ucs6Gl5i2EkBRzALqvXnDilmdcw9W+B4r93/lW5lgF
4IXHH7K/Z2rxT6MjMAJ91CC8Z7NzCoJ0kZkDdvDJ1YLklYnwTUo/4iGGouPqENJlbjTpv+EioWiE
8zTM9U1anNFRFX+BVUvpnTLFeoMlS/7KP690B4YtQpZfQxwaAOwWFcz7oa1Q/SM9xvIuQITNMygl
uumGL9fW2gUWYCsDIAWtUsS0eVVKtgiAKEllUcJ83k7lo34hUULo4YeGaErGBTD5f0NkeMcZiOHX
O2fAErG95EVWNPjW6UwdEjjml/ciUvnhrgTcD2Eqlsqt+WRq58hpZPHziHUuvv+HQYWPyG+Mdi/N
E+eJRT3efLpWBDc6ruh8h4fGFwAKBIHf5cAytIUjIb7Q8t7BqQg+iGd9+83rzD6q3f9NLdCHg4dr
BBKYOUjKdqTYn/eB9RuQuaaykUZT6gHq+AxYqV0wCIO4JWnxa+LFJAS7InEpgr7kjn9Opk3k7DQs
Q+1AAwJvkV574cirSDAqoqavjmIxhulnKHjiScVWrnSLGC+1ClktDcoD7g2OsWI5t3b5aE2B6ePg
e8z3g4uO5mITIoek2zugt9arKVQRalE6Ault7Yn4powD3HTv3MP5lT8kvKaIY5ZzgpuNcsAPaC9p
RxgLx1El84my17anfcAsYjtxBGnWldtsCUMGA8C8L0Yt2deqXVsupUDiPCndfIJBTNHBh9x5JTQ+
MiikT+91aPcoD92WqfgT6qH4qhp9dC1qeVxpq9brm7x/kAWcWSPPgqhIoRRgwTtIXmM8QIQLd0+m
juDALgBFfkTupzD8159I9lAg92rkmCQg6PleXybILg1b/ng7p/+t5o0mzRbLfWE4Q4q5pPGLVz27
TSO1sihsukVfCaakKo6f2aRH27KtFaJ9OpqXR66jt/0/DQ7cs/dhBvcjrpjJWBBVfpUGXcBosgqD
TF3A/K2WJzcoWMvBbszYtTwtUccimZlAWmrVFMlpt439+E00gWBwWyAWHUQacHEogcLAN0Uelojp
7uPvNCBPOHicVEllOESzgY62CowK9qUEpZfBAQC66CIaaz3i+8thEOrihcSlsoOqRO9wGcmw16wO
y17Z0qh0WEYsfkaqcXMjJ18rW7M/DmfzsyTUzsJ9SZ8+qkn465WuebDomzXsMzwVZNvW+rYtKFe6
g5OGCuMBMfics3nYTdmsad0zXV09XILed7rKCzKFPW4kIevyAShh+ws42pgRBk+BCJa6CWSzADFX
8/0p6s+5WRcRVyH4bGDwl+hs0VGPeCbBNHSNTt3S8xoBtkeWmMv2M3rExkxJMJI0+nlSxb8JMGTC
jrGbEKq0WM5tv7WEJjEtg88CmmBan8ehZ+ZWaGDpDdJyoVy7KDJdLaHatOptfMge0bIqdjCs1F0M
1bLN0fKfMge9sW3lZwNZN7u1bemzGGx+uZiKmVNyOIDxUCiVOpRjRS3LvWBD8UOLvz349BjAriPS
oQmUNQ1Pe3VZvMrkJVUCKfmTuTp1h/JTrDHcbrtt4/tiZ9jPtvsI6g+SQPPsUXge9AgMgCp7aLX8
tr+iERhPXbqYUVyuWpqbPz+bJrhEi30lpBAJqp2PIpspfIdgUlYN9CgqraLwR1OYA9HD1trTQNEo
hIGiSDuI3Wsj6qiKNu3R6cWN7748KDBXO/6ChhLeQKbQZMpnH+PuVA6KPcVqPRYQHTX5DPl8hgxc
DhLzCqq3QR5V7jUwIrAqe9tyLE4sE44KCY9STbOL3abeSTnQn3mKwP35/iTuDagjnInq4svYpJHf
OO5bY1Q3uAoQD0p4ThsxRblBG6N67U3zofXRMzwIlvk5g/oCP3K1r/9UH1HPRgq9uq3Ta8REapg1
NDzSO3ekC0d/gizhg3JK9G62s0DqZlU3CqrUkAKqcgKfEdcs5oIJBsVDeo/IBSqyHt3VP6jighUY
cxtbvGpxQTw31pDh4VU7bUdGATO9H2S6r6SCwsj5TIStWHrduYzRCu4NIEF4ryCoq0MUAHPSGYdf
1pPMsbHZGiKfuucBxhXjxT2uyejvPJ33F3dKyFtUtEfVWFPpdQa/fGIachGCvwBNs0glAOBg7Wav
qWagKEvke7dsTLxTLI0z6sLOzLuZwjcTMCpuoI773C/exRpz5UK7LiDGlrA/eFiBFsaMlHk8iemG
BHqrgXgMmATT0+fSEBz82sfIUNx81BPC6wPqsYeH6l39zwVDYuENNG/ouRIm6qDqozt4uIdFyV9O
uEjpDWkeb+2C1j8a61b2UTgF1NZUKEhxL3KuCT3A+I4/Z+a2QJp6dOjt7bTo2xVdGl2zuP1CdGiP
xN4SR4qXCjwjOcQvnZ7rGM2mXnu36Zuet+L15bsByFJwmdXAnkkkoSit0j+vkTgEhZB55oY9qhPQ
9KPziJb+PDsh76e/TJDvvwXdfaQv4bNKXfE62lMA2GBHf6pKlw2wEzpZ5H1NLDIt/AZhJom2lqfq
41GQRO1lmCTBR6qEUliMGnFVIENl+8HDCO80sVnaVzmacujnTmwHauUHkCwC1xw5W8F1b5NKZz8y
jVkjuwgQSZG+QeaP7n3kvc8gzQOj7iYsLiQK8b9EjYI1AYQXm15mX1xdVUtS8lHOt2L8omRpSwT6
IhWgq8UANVxkvWlDfueg4CSZ5cic8HU6AphAbkW5V5Jykkb79jxT1Ib1sjY4R+fB5TSMVhOjKY2x
58Qp/EoyOU3z2je9afkgK0UNSYBvlPbO0BNlfGpinXhB4Ki3jL52FzZ+kj94dh1Qjx/0PEVXZ63+
vz3ujuIc1tScFKmkg1nh6NCmGReSKj6czVeVpztzSc5ol+Fmh+x6OfDuksYVk1FJwWw6McY0TIhz
8UYm4kIKxu6Sgeu6SfY/zznePpyNv7WH/kxpxknFqrHPGkTgNVMmvgqHZMfs9zeagv8uxZv9R5PX
wZ9mPTiE9j8jadwC+ozAxNrIPl1OevcFt/1J5q7w7lFl2hsQWa/wl7iz3VW6GvvE9ErDghCxndfH
SUWZB8Hyg4Poqwrq5CU/NmwZZyElG15+kCs3iNOiB2+PWJFledqPGVfIbacZ9gSarnouDFmvfj6M
XR9OyFGKfuhe4LSHv72EHhSb8zfrqQC2KuNfp2IAiZmIhGy7Uqxr+Ssak5lvseU6XYqbtm+i/ssX
eDcIRNLk97RWPBtBLXd6hEEUV059r2eoZ+UrgQ3Dvrj43hfdXY+oDjHO72uEqdxtQdRcbu56xItF
AG9DgV5C1di9IuQ3sxJAD6gwW9MPBBfLFNRB5Zlq0UXWI88p+TzhRHCIrfMmkr5HToBDYIyPtaDa
l8K+qS9Y/6qOFooGWhFw9cTHA939TMA7cuO6EhEK0rglfKyfh7hu/hD0v+P7jzremfMFD/WpIMdA
vKmmkxJ1iTFs/kvBDdllKQFGJCLlP3fkXfcFptVW80lzOWXcj68GXz8Isbtr5UIgmhTKVwW9R3la
EhtOqJj08wFbmxYUirPaM+jjAbaovySZODBkSz52kZefT884ZAlJZtmG9Roh5FCB4/ZV90gf/o94
FIsL551Z+S0taiiQmlbUCG7tLeexF7jR8QVBMf+W9rVp+zaRQxe5bFWeocil7Lqsk6qyytI1XhRx
JmtgCV5mr8NcClVr0NuSob/qH+cD4G/wpC3ouBqeZlaqODY+2HHSb0AHtKOtZnVomydtJqDT9+dD
M3T/NaWN6vAwcdPnxyoNc8N3yVIiHy+8j1+QECoKMZkRLZcMEovskfCQeWhtGtZStsSO+x6Jk6Un
k2h59xmAT77O8//5I8QOHSGFnQYAa146YcC1IpEqXCGtXvSMd2pTlOBgZGbj5mBW4qWUCgOyvQ+e
kc0ipF9beURqLTQTRNpoYYBHYtu2KTdIdpkb6+ycal02dDGlOYpYvyXVIu/pMguVCNAVTSrf5aj5
gM8jvSF5A2E7dmOv8XfYk2yShMEN7PBrylMtD5j5tUBi7tBWHcJOKnOHbMp/UZqdbA7SphA4amnj
BwxdikvC8xBKbiOsvmPayD7/QTHow/O/wNzaTFMsbxUo1xtrT5rzIiMMPLXr6wFVtZQ5aESvaoIe
DxmkEiWuwuJAith7W1g+WUF40ojjCmPGAW8P9+Hilrqfw9wzZJ6KA4Xrv8eDkfjZEbvZmFbepywu
XoweNqy3pf1hKLMe+lgS3afS5lJ1DxrFqv8wgaLKvs5ij6WkflLfEravjISMWbQHcSW0u7zfqgpe
MWdHcsMhnXZhLQkgiJ4bv/6Vc2AuqBkCwZN2KnuSQQd2mBRDwRHIiy7g02fj+8wOisZOpFH1fuTp
Po+Q6T8jEXtA5aujShD5HWF3WCrxbVeV4t1WwwHHtZLBixezF9NvOgpo2YrbOIoqIWzrwTrSFLri
xS+iBb5vS8plk3X2bDq6mL3hoaa+8rp1xmOYEWHhGhFEhn94vypVfB6Wmt+dmWjO5x1oIJHpf4vF
uZMEkX15VqNsstodB1AyVpJJNPraS3wX1cf42WF0J3zUdMF/5cBksb+setazIpLyWqWmsfffNvS/
Y0XkDbRrFOEqy4NvLH7r38FzywKUiNeUh7U6vOcgLMCTOESBtpMIDLKFKy3cbkjhjZ3E78VVhrz3
Cm/4klWrG9g72YhOR5QJJ7BLBKSD6IV5I6Xxki6LKNH+peYktbIYzJjQrgjFOOuFlfbrXjlM5NBF
G4NpGZM8Z6dDneF/K6bi+W6HN4HQJSr88/lvaLalSTzwNt7ogXUypAQe2LpmF7rimPDBDN8+a8lB
1eagpbn7UsaUt2Sa+bTDV6dONaJiEncx+2Z9Fo5VVhpRysoAGS4uscB4hc+oLKpPbX6EyngCWmYi
OrTfWpPuhTbqu1iyAKp5zrNUd1eikUyWSwiy6kp/FlbD4d299/B+qfAgOJ0r0iX8PfRetKUb+xsK
9ejfTgUZ9rA79u/7SRHpoNfjEpWr7w8LjSgqPUitxeHb2FrA9gwE4chfepoHNiqhNuODVcw1dMoy
zWOgfLjH6R3fkUappJvGt33S1T1I6C6ORP41yTuFA3U9wA0Pu1LixxpbdikV+8p3rKs+hQbkfelQ
7Um31dr+P66cO33uom2+DuoGHCq5A0MpHJVXlAmdf8uOgqaN+CpqVT8noe1dieMtKVeEkh0Nu6bf
LZbW9XbxOEEfO/GAiIp9iKjS6Ym43naiL+qWdw7gQXbvRZ9ZNbIt21nwXazEgP2kVw5WCikJi7aK
xih2M4YjSLU3jfclNgK8+0oSvUQa7ja96s186jvI4qXB5YA66N/visAcny5kn9xw/MYSfb4CuDO8
SZZvk2OQV4rX1VBYWW8hqVlMepU8ijBrUD1l+Ap92P3ANzyquvAU9qv7nm4W4qB1YKr9UtFHODwI
dn4T8Mb0Zfeolzf7bG8UKRK3SbFM+FE+VrdMkPOnZerIXTFstyLLbMVN36ds101GFQA4tH4PWvf9
16d6n/PlayXimrD+hJIta2anGEcskMQCH/PTQPqI/sVtDz/7AY1IUsmNtjAwVE4mQxIhyzhg0ljv
nrgJYT6fFzCV7OAHLDrTvSlWYygp9lVrOLIqJw9ABMBH/bm3JAmWn7i54jGlhdHL3aVD4EjoeR2+
+VWEFlAIN8f7I0mJ8x4x0Lt+p4ZV70rhJu4hHjA0inoZxNQIgAdV8XgNcOl8paNSpABU5Suzdc0e
SpBzvYDwgorMGJ9gqDTazeiCAIGhfS/v6sMkwyIcEYTfpP7/VCpiGqvDX8375nxIz5WC66ytrWNU
Q+cvUS33TisFClAfdbnYv+Qzsbfpl5bkrR4aIHxxO4qKhGlBgsOZpZpVlbd8RMsV4uMvFT1MWWtL
VqRcQbVn57+2uyzSA5I/TUa3nCkVTKEOi7bJucUsRTmKmN/t9aEpQKOKJSVZsXOOuY8zMc5lSWaW
28rckSUG1KvN/fOf8SsvbY4GJ0axrBDETOIehiOThgLDzEDljBJrzLdjcCLGb3VG/1vPBmK/UBzh
0kYS9PsX3b/8J+Mb0LnGzytqkOXpfnVKfzEw6tASQJiplqzytA/iuCOVg0vYM6JJucpY4UaFl/cE
oxyX1McrsKmZmblxdc6mRu47kJNs3fOysSxIXAzvvZsCB1OlQsXOp93lWj7nWgzd2ahHAHkgvTa+
oq3t5UuP7rwotycj4XYSWmUUUyNiP8gFb2dovbi3SAolbUxYgJ/QhbMKA4Fpltc9N9pN3zUiDTcX
grM+6pHAoF34+U1qhtCAU314cPKwtK58O0jhjatOjWstIY0zGCjRBIzUK/7sAO7790Z9/CHqI7WL
O4keEI9yTGHA//CEtRm1Ba2qrXtSfuFUtEzWsOSoj1pWadeuk3kpinC451kGEogD923f222sB/Q3
pUB8/6ZvVkf1fzvtSeeoRvCteeiAkoJ3NwBJSuUWmvFuwzQ6YiIbpE+ZWSjLw68X5i7CRTmdFfNg
p2fLUURPZJvER5mZPubCD71hguCYQ9ckR8p3PtWExCrX/FmbI01PfoO6cL4duRPclZhn6cETBF8/
i6FjbhG34lvZXe1Ocav6mbCA+a/EOgYzQuq1rIF5T99iNbu2VuAI4cz2webnxhFlG88MoKCNkCaX
DapeHLw2LD66VlLubCowiPSmgn4UWhPEOCvd+tRMTbXJmuwcXnAKJUanV37dRKPZncr2jPmAZRSD
tN3N2rKpYfJisK6D6L5TizsJ5X4H74EgxVZGmC/cxg4iMRJpsa9J3K0yho6IEkTrBfsjBQ3yZgkK
W4cWRBTT38N9COtZaG///uj3839Gnaub0qCVm6cVeOrYZobfvVd5EWgKtfC8eJyT8TvANqUy8iFJ
c4n1NdpEcw334EgZVrHMmHqKznjfecI+ImkeYTx5U3lJ9DKtR4/TlATIiYHFw3a8Hq1ternPVcnT
ocunOrQTD+aZ0Vd7Sd5lcNiylaTqoFBDu67SHNZTQCPN/8wGRbBTATwQwPR6JR1IlwaVRxoCBdkM
0yUlt2u18pcnmJRaRRLbCrS0oQ8ZAx08D7y/WiPeGmHlNxAZCl0IfmGPYKgatOepTG70RyTdZX5f
5ngYllw7ddrTP13dOvGdknKIhlLmCyEEu96GloF9ZJbFUuGAu0sBAx3crrU/6jsIF5QwuAVsooQI
vTGy8agaDigBbX6kwh1paPqn+P80DpCQZ8rhG73vMZ8pMy8KzYlPQuWcqD+LlMEEeZ8DnhMYF2sH
zADE8C4NimgJ0+ofZrNMOihTNywJ/vdXEzpTJh+VjYqwnfWB80YO0OJlHyfornWvRCOuMbYB/6LF
KK0Y/9E043regxxNLKG2uYX60nYwy+U+SP9Fr1ZDrEmQg7ZyT7Kv0m7QyfOEDcw4cIxf4kAWLJaX
AnetukxlVkIJALflALZGx3CQiLJF7KnIvxc5H5X/CiKnlsTTph4k9q7Svfgknp5vriOTdOK/enqv
D3Y3PoIVRKk3NLnUi8r3q1MWZzOatHiSHM9KYZREbSm8rDLuQMOvxrsdiSvAUN23exQdD7JS4f1F
DnLdEjZMUursJlSJ5kBOPWXL4bAYFgksmoncs2efHgqxrYmy/IWnSaqHShEw6yarODg7p+57ogh6
1kJEqR1jbA9VjZzkzCtqQnZkvVm2CIbmjSmA8PbW18Y1miDjdjvjYP1szVuijdiJkhF/GfnLzfWp
a2fcsLWzyb6hE7RTP6yvD4HFg8IZLnkBswxPSimFQfUsMs74eOnVo1pYYWmqBVX26NlIurXpoWBo
J7iiKjkz2HsX8lQV+b51JhCyx+AahcOdzV5vlS+M8spbOyPNngRnI4+RUJZVxhDxlImuacLRNbq8
nXjmtOyIz2QhxLqZRRUjHJ+SzWGjgHurI59+i2I94Dh8UmKMPXf5FhF2xR4BmBGqQg1G2EDWHrLu
o8p4r6Q6K9UdoAGZxR7pJ/yGyDeCQionycK9KBkHkqZGkDPPQvDCnzfFsIxRvnoXzYP96KyhRYcZ
e0S/2rfhMZbsxrw1vx3ebw1DNS6p0wBdAvl3qkLJ1HtT2piEga2+EIO9GLgN4kQSLedfLZFhjPfw
VZSEpZ4hsQvBEk1oLgmFvCzZdZcGVnYOEd6ASgWXIKgURgXsKHmHpXX0f6Udkmfim1FA6IED2QPy
FlaoxH46srHtM2KRKO6QtkqnKrpJqx4PwN0VA/20JY+zqzlOJwidrqnOz+EdRH/Sj/ze5QBZlbJg
0gFRuf5v9mVu2WXwEclw8DHyR5P/wgX05M5lLejr8HGKKSb5NSqAdh3d835mI92JPSlMlYBotbH3
SFW2L5rY2+wLk/L6soQ8egdFmLXXqQtXDzqBp67+DrTmRVoDRv95mo0rjxzOl+NBQT9RhyOGlHbe
hwLBV5cNF11UMku50ENcle+fBpI8klormAjQwj0bN/jeb7+b5DX9g/wbWwe7IOJVOb7QY0Wo6jYz
IrmI/7vMV/utRb12XG0rKoH1Io4L/ZZyPN0FAVgze9i6NVWumuQ6wacAPz1BoMGjZK4EMr3opKt8
6TRB660VDj07ev3PR+S/QLJlAmhAV5+cSokOJenFkb7X2NLI5LnfNX5CyfRS3/5p03ElG+VFhTjM
Awscoo5Ft10t0r+gKkuDlbhqNzfe7gI0Ism/I1PWm5Xmz7Qp2DM/KGH00WuZS7vGljpxuMQ8LALs
7efXjaU8q+KK5WvS6YHokn9f/xPQMTrDHw7QErqNalqzec4HBuK2+QhbxrhSF/rrdadQ6ZQPEgvC
nOupe3zIyitC0QNm0LvkZRM8eulQa2bCNa6r1PKzEEuNrHta5tsQz7SLMttxsZSgRPNrWHC8zwDX
ZyV9WwlvkNA8ZwERIR+zfzHyGj9nKmT40TWJbR0YiOTyL4wx2cbmjhXMcPCU7GvdinpQEg411tT8
DGJYfQ0bbiSYhSTgxusM7gYil2BpmvwFwku3ubtpRtLkR3gCSsZkTkBOPsNw5ujKtQBdrGYDQqmg
azq3Z03yKMB4UA/KsDeBDxokMPPKNSUEZ1c8KYePJeg7fsMSc0N5LbKdrRhsPfhaAgQ6TFwQRyFW
jpfm/ZQanicmKLnnaZy5VVI0CUJzkKssvw9G1hkFPmdWzWb1UKioD2hZkcDWBLrLgudacBtnjoS5
7qBZAUCbZixbRLSQxUk9EFiIJICOhAq0R3F7YqwmXxSIXYpRjyhoP9reqPuwZfc7c2lcteequF5r
cxH26ygWA1Vm1p0aqo44P2OXFty0uI35/Z4LEoCX3sn7W24nxVZrX4KrEr4sFxX0WnrPzIdFBCok
wsOzkYXqLfUtRPSQXtrH+yHWMOG/4pWK3cR4/ATXHWVQmyckvLJQonk1QTkRKRvi0XM2xMNT/vyv
g57v6qv49yp7utchuc0CFO4K8iX2NWN0nKznjIz88d+yMkqV4TQRL02Qa0aWK8JPZrVrt/h1fDf4
A2tMg2unC4kQBvjQwSnPfPJcV+LlOrLv3WgW//ECmwsXHZSgltuMNT7dhM/j14690wmfRb02iA31
Dl1cO+jWmH3bLWLkyGE9v34ihWA/A2j4hB9shYA1MmEvlcOTR7eizU15IYfa0hVWxDHkRS+1d42v
jAodDX2B+fFydK5NfELP7WmApE72jhOVQWbwClbf80EsLay7xTC0Wzg6cA/5lLERa/kPI7ShYG54
wAUCi40VKduoAbdm0pL1/C+fBEJik/3ZWDt9fqWDWl18dZdkcwGELaYdvNuJDAAn4zSFgJ4psFkX
u32EOCQmI8zHAFYckczc7ZoyIktAsHDoo+oxsqyvKJJZsDOA6dbEXlpULZunmVOY2NK9XZzqz4Cf
H9DVEY7zCo/4pT0ReSj+R5FrdzPyggcbi2PWlENronBLNQ33M++lH5g6aNsOcWkhcEQmRuzDUrb+
v1B66dpCMJ88om7BYvejmBQRdvqWNsJTDol6YnArZHRYdmyYBpCc5MWwqL4KffPN2fwQUtrSV0IF
5kS5DbeWMd4GvYkiAW/612QHpAcPn3GMSJWQrXdbidsarhlni3v5hnK3r2PTEgLWoTp5Zbwx5OLx
NyEUZfLRCESfKYyiZ9cZdeGZalcqtvtB4LVtoskJZ39gUbP3lPX5iQi1q1z/sXVgkYpbES+VlwhZ
lvZWHlsaUafz7mxBSe47rzrwujdg2D610+Rd//eqyT7WZ5PTNbW3MzJaqCZnzs5fQScQIhAm+8pT
ERkIhWYW/FXyeVX5G01+oGybFJclP5TXoXh2+7FkR4s/P+GydYMq89tyeFGzC6WiodHmQlDp+P+1
DvNMxsH0H8Fv5e5FtuHoInUVDwPnukWBCZ5rv2kE3FUm/HlDuFu/PDtRpAuXqh852n+bDmVoMRK8
wLNJWO/XdIx2fqPop7Il+YjZS9JA6O5llNctpQ4UNAgp+W5cdlZUxf4gZsbr6h8p36KzXhTFX2UE
JjW3rH++mdcY4zNOjVnims3TF+5NZJ1jSdP8DmoOfKAeaeSdTGPz08QRIvxEdKNYAk6dq4w9/wzf
6HtK7L5Y9bAKi0YTHmhkhcmq6gIknM/j+9ILI2Ya3q+nWalKDFzhmebi+LpoddDdFRJRiTnEmnrT
1E+WtDtv5chtXTegL4dEDE2+wjeJ8QioENP1EqFhsTHjlwhkBFw9+atjcV/d3G2FHRB/rkWQTGVF
Ry73iCaXedel3x44e8M8Lq/SJIA13un+Qu3EOyA9ViAf87UFmEcjoRjkPuu6Gd1SlSyMlitBflQJ
DQXHmOmR1lPBuPgCMNi7m6p19uokUJyuq5yc79+DHPBGyqCWxTZEhc/WV/PG0DO8Wy08xxvUibTW
vT3BvB/soAnCbRWLW0YI8bVukXcIYSQUt3N3lOo6Lra7xt1m31HYvm9fHN65Ju8i2RVJAeLimBtr
UjKJOxzdomRngCYEeEq5jrob6BR5H8UiU97hjlhwghHrsr+mn2k67RwG/PnLPe+BodGO12Tk0p7R
6v4Gz0+et5jda8hvbchFXuQTkqx7l2gcf+edilgyeInnDvcvs0oXJgcQKopuIe4cl5XhS8YmSgL3
YsQzcT9Iizb/Tgun0UIO6pHLB2q1HpHYPyO3Q85i1v/RJJbFNGJMefwxpoW2RUGcqHaIDwt1jQkd
qEXSzzi5XcD2SqC4p3ZrP9roqvduG4cvaAGbT7q3F0uNKsu/pKD/qySpnOGfUFdiD+oLpU1ArMnG
BdLxmCGlycuUUKaIiuTUvmEPCOGDs26uo+IYQdrorwFo7RSKCK4BDORRVYA4BH8Vdh5TZvRRn4h2
0CUu6Jq0QEVRzNnKAMkrkLrCxgujCbfjXPb/ulpjZ6lSZPaRg89OKWF16HFXfbmkJyjw1JMP0IuD
u000n2FC3Zmr1y5nX2OfMzoaoqB9vxW1Jtos5u+QOdr+w4XVgF8oJdfvukIXaSvCHqxVLjOKspZo
eFar3r2QnEP6vbbdLXH4sXlQjljGdSWktI315/cmVZvLDTGV44inyOEvzEMWk4wlQ3n5U+inKmu2
SLAE1RlUjSQebat/5YmKp/dC395hmJuYT6kU+EIWJAR3CLqNajqUTXFzyOMzSA3Pt6lmxxw+aJCl
R2Q5doXqzmqbX0w4I/Bb7nBpSGfFzOQDw1Mh8bHS5w5IWhnnrCsZMbkunwiQO8RBGifZT5REw1N8
7VXmsbZMbo4TxVnjYBHYndQgW9CNgo0L0hZrYgv30gU9/+GRpDEszAw/AIWwpZkHkSkb2pJsePH5
BsdRrCcl0QqgOCnAhJJFUJAGK1Npojtx/I09K7BJyjj6YOkwdT4Req1OfqcdiOqE+fOCSyJdQLKI
BU2kfjY7p2YqbbM5t3FWQVhjKZDTcLduJNf9pVss/n8t1i+i3vOQhgpqawmQFDI5zVpWeeS+TXTH
IeeCbgsiGdafFMc7OKWVkd7/v4cmp27jRBLJ+Rbh+ZAt7fLGhCgAGb9wqoMFhfb9+SFWK1yGGEZP
ZCL5pw+qgWMALTaLMZssZi9Q2oeXh3XLCCJ63+mhAXkGYC4UeLZpHTYFZj2GgABc31Qp7KcGYUR7
AH6ccqhYytUv90G7UiBZEL+awa6ZrxtEC3LRTLZElYbkMKv0PWoVstZ1I6RIgFizlwYq1Ki48Np+
+WaacQ9RtHG7n3hi7qzut0m4bvqQo31cC0f3fIXvaMVfhObMtxoY799KfPRyAsmigpQnoFRH9bgl
hQktdUMapxnWjkH71BUHs5S54KXeIkLggSY1y61UO+IqjPWx90HeuS7TX5cK8lznQb0lkgJzSj9j
/spwhSfKaZtGoHKi4GLM3xfXc9wmXJtelCCXTBuTG8FPss7vVeYwyYLDQc/q4HLSTMSfWXVbnKd9
qxgPxCXaIhwhwwoSWtIBp/su2/MTzvVfYVsW0e37ZR33AcV6A3fqeNkqJfh8QywVBkRrLCr8BqtP
pi1ZQIV4IVIt6NO4uEpS6plLDi9MVmv9HxSeAemVdBjn6MBdoxwT57rlLTG+mJ2Gl+pXfdjejYnI
ktlDEfLCCnKefHA7Z6Fo8u5d5hZIXYVbRj2a+E1wxCpvniBi3Q8jKz6uZSxlX37rCs9qsmjM1nP1
KT3yqfmzZPTaEsxikDNLG+AWHai5Z93jMIBxO0pSqqdJn4glY7PJaATc8yPElesa91vUv2GF9VkK
GHq3RiqYvrxMJMV2ghkAgGTQHC506lFR8Q6g3RxQd+jYLftbVkXn47u8Wse/dLohfIXGtwyWz9S+
fVjaAv/8+FXHMkR2ZxoYoBDheuZV+UZDy83Azz7/Tpenxrcqd94dI42KDn346NDyihE58WHhBhNl
hN9qiGDOOqFVd78snektJWRAB2A2qk/8eO/nimYXMLj941GJt/cuVpG9E1SiayX57ROKZHzvnSMO
PxmOpuFmtKFNHN2soKlnXail6z312UGqLHd9CSABh8NOwAE8ZpMnEivtlVoV3P0OzQMx4YjKAtha
hoL6e3Or4q6XhcVJGOO56PfifNnWvwjRpgOAjY8kCqiCyorCnaaEadZtE0uuYKDkJttTaj4Y7dIX
WHyvHyu9qCYNis96g4iomOzDtFb8jW3sFEz5/HhfDKreI4Ilaw43QQdcgiXkEopATqs8gV2gOMq6
LXPE92qKdwvJ+zf2kju8Zar/HqdeeBGnDbWia07mr/Gm9pztcokiDqPbSw8XvbAtxlG96hRcSWjN
FrLchNsYXSXTrEPGR9HRYiB6qDdvK16E8BS51zKH/E4tKyDN1ZprG8AGhhACVdkgzhgv/EPmtaaM
7dQq7yXeF9QY4tGiF5vvckKO91B7zZxgqYtBXpgmbJ97CYcLTdUT5/2fKabMi31aHBEAMh45Kx6C
6t7oiH6KxBOeTDK/dk7OG/W7Kb/pmkiNO7Xex3L/bhNkZ4PAdZ+9JvaKL9lollBX5EyQYqH16iw1
X9d/OLtzz38C5Q0H+jZ0xMVc0qcyjN10YK+LqRUnQnYCa+u3+t4YqRyVyKcVWsMYjCwHt2GuVUZQ
xn9LiELMTK5Q0AW60YmuFhPOeXsoZNwnzibo1q51pYeU654k3uKvdJZRnj40jxGEZavNiVeew+iL
PyJJsi+W7iMA6lb7Hw0WhEfv4IYhJtXsc1smQuZXObKBcaTkljGY6FznQ3PxNArdUK0BA4qJEpsh
mnQ+gAIlQFVSWQbCkyRrpUNsPiFP+xF4SX2qiAyBM5uzTeIMkFouNQ3rKhSyZStXNT8EB5E58wXy
hEehIJR3lqSve1XAUbsKB+bPZ98p3P6pwtgLzjM3NV4rufDf7EHWJ5KtBs/XMCuDo7Zb8K60GmXp
RgWbaXqK2MArviyu8boGNyR7Sx4C3BmqRDbZ4/q17/97paKA7oTl5Qt6UsIR/DrDRWjmVu91p8WO
po0O0dweQFTL429ecsRz7y0D7ltiKDTmKjZpGQZEjbi7gu3Jy/aBTjixq2fmKJgmBUt9lzY4JCRF
cvuB1AvUjT+yabqVWMDfwc5Uzoa2QNj2v2wOYIMWPbWSjEOKVRRWw5HF9d9iCtzFWvD5RhonY4+J
C68XCvNVrcjjb7Uxd64QTnRgA5JnSP05+BTxKr16x8Pd2WP4ZaubrWJKmIZdUeshQukYqKVZ/BbC
I4CzJm5V6OXdmHSv8coCnUeqPApJE8c1Re2O893O9jtxrQZWiJxnCqqTGjDwYZ+kXMGuBwsVqGpa
brRl4NRN4ROG5UrSduwg19GwBvMd9R9u8hnmH6RLkmr13HOygha83zw87cnnX4pSmkJddkUHPbbS
2Kc9y/puhMeLscd6lner3d1vNuYGR0j1MGleZ8sZHpbO3cD6LR/JG2JnyogxjeGUBYWB4DK6SzjZ
hl8wdivOcPJITPb4vUT5A+33ZdkF73yCrCq4RICJLb5vPAYac8f4EK4JSomxb0fyOTQvHs0QhbTI
PQw/zjP4GFNflwGl+QC+xg2RxV5rcHmZZDQ27M7m+7kl8t/TTKkYoAS9nsOdaTMfygv3+aSdclcN
dpHo5eDoK7D1lifV6wFYqQWQlgIH8zLVrFfZ14w9O6uqGneHnJ1coLGdpmMNi8oOeWLvknLUXJZn
672KkcirNDloh9JhRvGUj+oMM72+m0bK7jfSlrhmqvQFCVuoa1v6S56i7et9JK3jTngWxpGUZmbr
7B6+FHpoDFDTRf45+QU4l+jSsVAe9/iFC4MFJrAxpHBDCxVNoLAchc7mNqON9KqP/rS4TJVvOFfY
ZOt6y9nyGikKAO/QITImY4L89UTcfXYIHX/lUtFbtDuX++0kL3I9vs9t9MSjnW/aVcyJ/LOATQ91
lE5tY+c/1l/U6Ly3cMJ/C0YubEKP9Ki5z49KzDRZn6CQhMW2SDpfqviMHN3iDBJ7wcOBxjqUhLVK
PThDpZHgyZ/rJTeq6AgO7sAS5R7m239r0ucpyaoKTCcD1iWRkB5w4wSq4OU0juQWjPoYs+7z88jc
RHdMU/xl9XKPdhjMkz6TJjHGmugvOMqFICJ8NR9Vk4VZJFf1lY+7vk1vHCuMAO3o4ebZ4GA67KHG
c0Z4Qrv+oIp6eVL96NLWUCLJifuDP+vaY/13ZflJcTCnYO7GQn5qX6qMBk1MCwHLIx0pGWTVUHqI
91yTlEZYZDcFwTvK5QjBO7/4ocxuukcHc5C+85xL7O4p736NEe2F/9tBrlOPcgUGZ8tGHxGvVe4G
ntQi3eleKynLF7VxA32wNfIX5mxO5/0nxpRp+XfUKNWKbUYoOJPRVzTP9Ktw69+0LBtHVW3YOHUt
fpMnhmjDFF/P/tVmj/BqlniEebP0tDEHNEl7I+72nAI5phDOy59j0PPh8Ss/0tknyEvkQgUPkmL8
AzYkW+abluQpxzlxQJc2/ugWKBJiPRvv3TzjsL+rUEloVKRdtkDurMJ3Kcywx4dnxTWHgTdhsG9p
EH7oVzakumdxWOgBhAGpryjb05P5e08c48JYvcItGaQpQ1hEs199p1CuofUr0TnFNkEn1MpDu9VY
O1EDBgjrUjKYcgkWBYJFgsOQsLecqiSAHfcFekutyaYXuPIs2/phcmo+jDyAUHeqdejlkl3+/EvN
QXW64QgLJE1OLEndCzSr6dQAmhJtaz2JPx6K7RWy0keGeJl0o2vN0J/i7g5zRWJ9hcIOiwMEuavc
5VixlfVRRL9v1lF4Ym8UUX9hhfMApOJEdqtkf7Bo+Uev0lz7LkD8nxdEHP7jFTJ2wHnbxVtaHuaN
ssmNBqTVn3kp4y4JSh80ygL0X4kptqz+6Tci8rAMdJQVcPNnHOT3ErhM7kKr2LmD98hFrwBSwqUh
ylHJ9JSwFg6eCtoPgne7/l4QPCw+LIpvhScoAsPPQGUQ2oa15NRZwlExZfRttbCxTBwUGJrhZ6Fk
N66uShXo/GazjQ0WIa8wNOzwn/mAXJL+qTFZQz6tJ24htx9l1HGyN6p6Ny3G8I3kuoFxR/vP/ePK
pAKdwXacokSCN8FyUOzRSnxBOmE1zgQeWuw1m86snRXomGF+YJQe0Gx1zjO9CidmRYO6vmbgUbkO
IvqgvAUY7fzkeP/OGS1B0IslrSY1bFrMNrCorDCJ64rXGuc9DMimac04MslpZ9Oh11nDYm9RKSsf
2S23j4CS7LyASFLo8r6EK6qkP6bCuqBukxsKfnZG2wwhwM905rNeKDyUxdhuhlnUq3D3Rej3aqfH
q8Tj68hYcpNHjxa+AYMG15+MF1n8X7AwIF1eFU6QBv3U0P7FXWA3ySS3vSsSNFQFgUOm1vuZijRX
f+TeXUc9szNo7noMtqcijM1x+em6w3zbbfBgTzBl5MzLJqL2YjixWBwpw82wmHREbwr+Z1HCALKO
PlsZ5Oz7B5k6vUFu1s07JVMFibAe7tzGauhtJxnTQ35mo3gf7rSKbIk3oTJnhBGVeiBmj1KahY4Q
lNNyTwfdIgfufJwxdxBjzY/a6RAABll7noLlRvPwE5CTIq9QUHxthrmV5iB8+qzeznz8NSCslFLU
dj+PFd/bWXKnnpeCgBWWdxAf8uwOy8aBvcS0BGx8CYt4D6yOzxNQVxAYSQXDEWbDEZckIcbKpZ5R
25YmsN9kdP9B75eEXe+4a2rYtxih9PaYs2C2G8zTfgoDEQQ73tAxnw7mHymg0sGDGGYmrsQur0gC
mF3vQGreoUty6mhN/02JwnHLmvmOzztTaFkzk5PoIym/nHGjGrromm4DqAh/+4Y6ycqBX9T6VRev
fer7940sqG8VjUN+fjKWt3rYr6ZlXZ9UnsvH2VnpDRW+Jo1DV2g8KCnBhWpkf1nKlZz93h/rCMI9
khbGyfA2zLX69fkz1UoN2GJZ7VT5Cf9/BNhMtTlDlHPhQwrVMslH2UHobxe92T9kYCcXncYT9j/Q
MxN2vBWxjOqL+Cz4U0m9Zs7iu3qX0eRtOpTbsrS23Z7QnTgL20geEO5HlqmIECAG0zMeEi6eW+GX
X2+7X8okJZxvC8dyZzWW5790IH8ywVjdpWCl4YeG6Wb9/YeRynZZyHBAXmOxXn65qW2qf3hrOKv1
7RwS+oDWRh3Fvl1uTvcwHJ+uFu0Vkk3Iw9bgCnmJawbMuKydaHOTGLj9a54b6M6VtkO2CK1FNTt9
6aOHyZdH6aQm7v4+XcY8FX/37HtKjKuPTCAW561vauDtcxYI/n78qmvpV2aCQYq9t0kTFZuAqA8u
feoNAYVync7nr8M6DsmxW3KJL87CHVp1p/OxZBo5MWkjtOkgZDAG9SEbjIl8Uin22dinfh9eWPD7
cKB7BCqZxUzBdVhS4ChFd7HUAMdJ+nMNI3sNNkunFsZml50sdJ9NOxmVi6RYC4qwHBth3xVMQPhz
FCAP+vgsHqYmLOAgZMs3AqQnVjILVdequXWpheM4QzBQx3Dyd2MrEkfX/VQD5V35W+Gyu38mqS8A
PANn6T8ao7qJ7E7lv04ZURkoeL0Yh1UsoE/HgBy4OA4ivMuKVh9bN0wp3Jddo+b4BTotXm94QdYW
zdwR/0bCdBxwycLrbBQDqCc7jcKCPwx5Q+LqINl+PXENDlekAdrYjw4QshQr8ghAwqOCWOLK55s0
IhA6+yVyQUspGurSAVl8KhK9h+YT5TzumgCEjSiajrQFMdP6lDtlJsc1X9y7KSXSR3Z7URyjjLvU
P2RWRFIazE5vn3mP+/milws7zmnjUvJLw1MiGrHi7hfYQIZMoy2SNw9nEcwZFbevReRI5B7G+7rX
yKfKShwXFMX4ZShRnSiPeHgORDu+HvDhyE0dOlKY/XJIRT4QNz/KWOp2odsOWiLIKwWmBO5r33r3
kyycL/PL/JA1A57kpEe0lHIPXFdF3PqsEQ4Bl06GGPYGk9MvpCS5rC+K/etpWmXCabY68vpcJpGA
8QOi24rquG6+N1Zg0HcWWDhuqG1naZfN26fkYJmMrb3mLsFM/tSODquvKxejrGCp77Ue8HiA89Tx
pcMFhY4WxA/NggNnPp5ZXAYvo+9j9X5VaQcIuJhX0EdEci5qQ5ZtYZFNX1ftkq535aabCVoALT/s
hg8BQPhRQ3KeN63M/mnTKb0rsFL/WgfeCPeJZj+TnEKK5LnRMDjSVl/5nRFmKEE5KJpNEK2JNwWA
aF4pUanyfrZVluV6FHuLguyYiseA6Ms2Gbw4zHXfKLjdtCts6lW+vBebhN/0xcUHKJA031Ffwoht
ImQZj5rohN3nPf7jr9+68E69Yj3bL206QkpyULUiw2P9idBwy6BDvy2PQlKHZD6tTkz//0NK4xsW
B7XX0fiv2UMRf9O1pbRltAiDTfCJC6Tp8wDUa5bW0FwddyTY6U3mMycc++JYe2BFZHjxZ1MprSoM
sG1iEu/8btgCNbpZlFzzRNmU0HuvHETQMj8Fn+m2NZgLthbrQG9+9Pqh9kTeB6j0hggv2hvJ/Tr6
ac7X1w68hr5n5psOxuuWNaoED1YfYd4ixH14MywaMr/FMLAmgCkzJWGbUSPyumS2LjQcuTkwTIdE
ubOWXHBaDIsofmRkUqkHRDSE1iaLeMmpsqeNpA5XOPniKOAruikxTdVKRO+6c+QQhFIXs5oNvIve
YliCIXXEn4/MvxwR4qIhuWYWe1XPY22rAQ808Zm5erHllFvZl7anatqCi/6oYd5PhpfV5mvDVTVl
9h2xHqNciIgTNbRQ8QyXjiUD7T87UHFLin2oMviwaN/0ldAibwEPfTi82AOTUnTSK3xymbXgLGaS
ZbZLMZ7k2lbD7PgrF6TVKu6cU0lOe9+TsC5/c++WFlEjMBQPI7pYB1JW1jbkXba5sXDNUuSAyxM/
CqOmMXTSFA9tQ50ldXO78o40NWUNotx3L2Eg493IdNaKHjRF2lu61jdYi9oytfHeoDBlzFcT41RY
DcHbzDaNwIFD3daYKI4Fyvy/TC19ng4Zr0DXRZsnUhmvE4httOO63CUXH7XjKYt3M+wBrv2qLnNT
z23M2pVl/e7w7/IdhJfnLtr2Fzl+0ixjd3Ve1jAayrB3COCS6Z2acsPxipYJPxOtGoB9G8hdli0e
QdPrOUJfg68ONL7ZbBU46qHdE9sb+weQ95+XxxRkUoYssCjHxwexqFFYS1Z3yLLgGENEtvyG7jOe
is+UrSJBqmLiuG5bRWxEZ3t1A5e3B3OPqg1EMRcNo9xq7ZPMMJp5SYCRzd9RJgNW6Ct7JiKMOCHm
uXXj9l+wotGjtdgtMT605uQa6giuszCZ3uh71pE4VD5NLnDmczB19hCma3/s+kZos7VQr6OJ6Zxn
UNRNUlTvO2rynP2Y+7jomCFaafm24ynprvlW0Juh6mUywnY4seGvZVJms0t1mAmwxnq7aZg2/Awe
9D63jJm47qEnt6f43ZXGcpFIpKnvOVTa+dkfFPOzaBqIv6MUdlpAhEvq3FhKvyqtA8qeHDyMQIyV
LYeLLVO1lR21sUKiIveknaJ2UIA1tn1S+RMMXTgScb8P1oFYdZF9TR6HQYJ/qPjyp4vZTOH/edaf
gmkk+3P5e3YVAgKbUSjsKoU+GQpyZQmzi++c9uWnu0tf0YLMQ2vD3314OL36AbrY/2PtYNJq8Wve
tDx4IFv15uD8oROkeGQiDNkuRynTpJijCME7yjwKZSN+OLxXFXEFcIZyiyKfYjUua5am6sVecBsw
/fmKKgkflcA2C2e7uEkm6JdSTk6k71x1pFzAdK+tBRL6a5USyLzN/0bc4xVluQ5ASS8fttUg+IzH
UbgkFH6fbMhV3R6xeYhyCE+yPFQPj62laVXMwjLfH7eCVE0ZxCAMh68suUy3goTngDvEE/1bNtle
VpNRJs6AeSCZ1JpOLREuHNOlhtivIYSIPURtbicXWxQEHRX9YhBjQ1+YptqLB3oYoCI3PhoKpTEC
b14TPv6zaRGOlLbMfXwf90H3emn/udGcMEt66VEBDVhdEsgH7iacQxqa11dEW6EuKl9V9T+gKcq/
fzFOCAg++ErA2FlhjlbTu/YXYtHlrXaa3hZ0EOn9K5G5Zvo9BAEH5ndxp3Jo/gPx+WicLXSvo8D0
w5V1TrEKu5nx5qSsPDaQn24W52TlJK+vAmQEegdiu7FqtAaBUu8kE21nsMG4GdrOgUSqHKvQGQJY
H+/1v/c/gPcQ15EyVKKJwe5Vc1A4MFQK5e5uZugIgtPbZTiSdx1SsRGjdKz2KQkDWA1KiGuR9dV6
OEIuI30ru5uFiAkL/RrOR8aRZB+7S+a/rSwhhd+wJPkQqlfotIO7pj0R1MnxC5cpyIMWP+0Wt0HF
QjQgVZfWDES5/h+liNPnzV1G4XHgHhTe/hpQYGcgEylvTTWOdh41G6IpsWNa6T+0CFi32/42K7TH
FUcIWRZjzUsn0p2L/Land11VkzyVRo0islV/XE4Sx85d469fjhD+qNzn88j2yYUIeSI3s2vtzeNm
9hDWce29SOvfmVw9SPh/oJD7OSbXmg9zSnKQONvdD+w5OkuGcf/sDtVNbS2SMsOEVGxyFdAwF1dr
PksYvcSCQxVVEHMmlk1JsmLaYx9TpzncdC2GjWKD/010zKmD7nxF4E0nGi0Dz0F7C4hQSpVYZeYP
nzVJMqMd8SSDDS30/P5HZ//P4p/eqQv2XviTFeQLdBG50DRg6KEQneR53YE8nc2CwSJTFhMoCUYe
Vm8HXDfdOzy7R4QCc2bw4KCYBCQ7TyN1Akk2JQqhBMm563eZG6aegwOnRSygeb/QJ+kIU2Es+L3m
4Smw3cfb3I/SMyDoM6Ne6iCGdmCP5HWK5trxTtOnt+lU+eX5Yx3N7lDfxTpwHZicAZtLMfbR2DpK
ihfm2sZx7JpMvPQy85UnLAoDxx3erUbA4o2XoWHO6DZuqys9GyWaWG6Xjo3f2QuwFdeZbbuacO+1
19xxxmIMi+xhLHLCVFyYCQuDrrcXKblCfxInPxrhaAN5N4Qm+EG8yxakDXwSaXGY5bhvU4CLUhd9
Pd64XUkLb9oWwkq5BwcrJGiUTtoozSU0bU9y/6jKYCy3/2+im1sxwMi78iXpr6s+V0rwvaeiBEnb
uKDbAPHdTs6tA5S2eB1JgzGT3Rtb7yVr+BNtB0gtSa0HqJ8vAnGmeRhFdQ96Zp2DH1I2+m99HhVo
37Qv0BLjmnNgNGuliGEjG/gAFbjUn077VgzaP34oE2jADudSRN+e1X0fxqwPFoCDngcSUrjegOTQ
/0WD5jbg9ryGyIEnfdxeHeq0tdhL3BBoeGGIqZ2pMG4ComH1JzN+KMqfemA39hTj/ijQXus3Osx/
4GKwzxypg974ui0JRRSRMocPGqxStitVGCWtouL13GrQ93oxdyqEVQZz77OkfM5FBzFjvZWtwVwI
2Z3goH0IheNsG6iplPDhdTSKjx8y4bEA5WLglw+6ZP3tMG4iOYaET9p7igMJR+7ZRrFBBK5Cl87l
zGp5do+yZuX8N1qEc6uZ76hETuR2a4WTzFuBv5IZ52W0kjLDXrrOPiCwGQHlXM/z+qzo80pCbWEx
41WRFLmGxeCJLquuTg9OgUxPACDHGvH+qqowr3ISI+zup4N/3gHgpA1V0qTNdmiYB/bIwCLfNrAM
lFyanXZAM29d2j38X+BZRYPMSDfM4hvRifeZSraPvVKbb5P3qbw9DDWuKwYB3XvuIBIqcwocGAhK
p/jRJWId0DeAhwgWY20XzERmD70Zbk7QijVEJmWtb7uvdxvK4dQUWLXZDYm+2DSR0ZzF0VcDIDN2
sub4/OSg59536WafEkAvisjIhLcL06Y0RnCdIp2ihTPDb1ySvGfWi36QIjIxzOzuQPSq4o8fqsk6
R7gCCStuSakJm5JtlBN/I1gg9lo+kfiI5UsYlzK3z/nfp6zF4IyDiIPn7D9cMhSrJPQ2nOCdnPSv
R7I7/Py+g8m5zvaM4f549+QBnqNxm5XnCTU5dqNw7Tisx62VPaj016CbpjkhXAW78XgsNcW9Btzy
PAEcvaDBXQZobwc6aU0qELRM1O665S9YcGyXMkMy7IiSW4xrK0AcD7kMqRFjNDM8n80KBsJ1M+jE
BZWbPEbuUzm61N4bH3JXzJPaDxQq4Alm5yTP5SaThdeL6PViLHb7u63GopdrX1wSyg3MvoGnXMTx
CYMD7GiCT88/K0jgI2lzBlUwJR67EVxRkbxKJ8PzP0+oSHRrlTBVVAUEOa3klf0CqYsduTv/Zz9+
4Yobpihv7+qUAOfuBFD3kmRm0/HL8XwvpF2GKVkq5luZqE2ChQ7HyVLNIUGOUkv6eNY5wwAFX6cZ
U1Z0/xctpA7VVCtWJTK1xb5zZxj669Q7ZndKvcAnErUyUll6VH0pJxP4/H7y6v1j9ZPVRyKdXioM
oJ5qGkfDfgN4pCmUqEzqi89XukzMWnZdwAb9BQSgmMGpP6bT8M4WKl3ig2frI6fiF6xQAviolrLW
ymoqcOq3IdkMfl3vAVYJWvcwjWUhi1+aM6O00cnIjDZAUW5ryvPMzM9NO5Gw3GKj4Fdg12IS6P/V
+hc8Bw9GPMnaYkseTFhzCXtds9VnDw7sP8dHyMkVMBCFeZVEnz2zXZBSqDC/YJ4EnkEtml3vGkbR
G6El4MDHEklpZu3c+6/7QvAVrIxXHj69Pfam1x4iVDev5Y6xYRwGFkYjm9P73P7YUP6VrXIBu34p
RNfmvtqbGHDkUqsaLTKvNNr/K23mnzmJ4cVupCugB1CDQETCFAggxMl1hEV8TAg69YU/idsdYUrN
xU9xQmwhzv+DcWNalSkVCsO0s/LOKQmreOttKDeDhUgzLLJhJn2y23IiHES4UIRQyDv3xRxyvM65
KlBVSrgz3vvN/y80Ir0IjxQ5/2cQqJTEXrl3OeusPEYSSh+U0Z/qwnEnPgO4d4z5kFsNrfL9lFLS
C1xGeWx7K6PDUMxfA1epyXKh62DDHI4nngsNBbNEoI3zwV/npEiGM4I5ue6TkO1XTD4ISBcZa0J+
QNTNEhJuQtVE08RCYK+x5nRF6KmBJTUxBtsSt+RIg6vsHXpLaEiEfqYIcdDKAWADAi70n4qt/fgW
T9B6QUc43JpTnH8PEtllDu93wxrHbWmaTkczsV7e8z3LgZDWsmRAYiQKJTYwAq8eJosMY8sNXHu4
U7RR7UjEZ5PmOlULP69kHovBsJmUTV/k/c8HXfMwyAjj4sy2TQW9UF6cFlzSHfZkUfnw2WooKmmj
z9wfdoImbNwSIvAce3M8QcEzMLfL8y3S4n0o5eqQ9Bf+gqbl/Z5cwOGaH3FydCZiGFtCGL/pw7Ly
kq3bNHk3oXcDZ1RzQiG7mXRC2NbejKBdfS+WGz/1jM0N7q7cVIG9rVHJWA9Yv6ieU3cyjPYaMwza
0iBYDY0DWXb9aPSMtdkz5tg+mzR/m/ghAz+cBjsThtPoSPvGaO7VcACp5Pkob+w3VVbiG8QCN9a8
KcxlKuNAQSgnrd98Xa5vOTwxyb4r+Qpv5InKg3dUOMahENyAFE99yWodvWCw8b0Nzg727JggMjfD
PXscWnxvO5079/kI8q08Mm36vJ2zzxKS/wMKKhpcn+ULCkXV2S2nvom4LBup2Fdoq4rWdW1+NTIl
5+dG4KFGlLfy6F+GHfzvYBw+22gKgXGE58N2xvcEGhpoGkfuhgYcCT+WWFc0e4OT+fnB9GioRvD2
CC0LFh/xaxW87Hotk3/fUqQLPUN7W+k3eKD4VSeMDd+uc+tWaxb3VOQUKSLKb3RYKEI11t7u3jBO
y3OQlb6iul2K7IL/CX/BaNPc2zOJHR2TAX2kZJ1iBlu8AU9HIdSpv3CWLbNtkO9vKiMdNaa9FZbJ
+1BMiYe9+FOIOrWxqqgJvuk85ec/TJtuFwLpoh6yvWdhtqa7ooisiGotaLTY/0XCxo9mBLhHaTBi
qi5cUUjs54UyObR69RAIntzesdKthR6jZzMdMt9bi4oqIehj6BSxi4DOZ/05MmCX4s+y2QczMH9j
pwVFsZvB6e8bzudR89+zbqZ+7m3B+82UXZ2RwPQkfAPxv4GzJaETYF2S5eOjs/1F1T62t0vDVISL
K2P01fFqUu9XnizJkoY2i8GCuEUF7cQ6PY3nWsR+BidfA4pzkkmOjxi9VqJiIBqu1/vyuE0DD9oM
8Xq+VG0JVtsSMPl6NKTV+LSeXy4zGGkn5X2rxL4hhQau6yaKFyneDl7ZLLzc2iX/0bTT0QReiJqs
faAqgqNA+HG8XxlyFQkof7q94uOIOZL8p52r0G5vxH6kM/U1DozY4U0cePOf4CwgqYwQD91so4nn
tMTTm0agmrbJrZhf8skcmD9sQrFxhr6qbGWSkkyMYNpSZTSrLsHLqod5bc2LwyKFpt4nfsoQeWyB
q7HUJ5pU8n7NqIZ5MBbCqn99spyAG3roPfrtTqeE7+ynCyy8UrQFliLBE2r2njF1ZrnZQYmQMVfE
FBqsZ0w0GricDyd2LexP8xD16vTEr0vg5bOvfEQh76QUjte00Uo0Tc1AGvr1z+80aT6kOOSYxhuK
SIOYylJtRXVllPR6E2eDuAy5y7vOJGxOyaE+bsZI9dLET7HiskKxJurDulxyiwxKlasSZBiXPsMM
UoaUiSzx+BYxWKLjuArKgt85OPSooj+uR7W6zlaRH7CseU2bo+XZwVnCOuxm9JYLZ4C0/ZybA43P
NXPQS5z9OgHheiAtsTooiHVjPuB148mLrmeb1OXQ1kkE7lfC4hl9B+yidZjHq+NZBE0IgwnsnGBX
fiWE4T4MEqLdAUBirfZMmQGTFcBGnXtcdVbqP7TQtVLCQpY5h1UwWVDUKqWqM4VHeIel+ud/VFrr
wPZGdP+AgMzVpK9TcBA3s4j3OyuKH5Hth8Sv3yTqQt55Owp4e3fRKzDixXFXihqWtVslKyJ1IcBP
CVCMefXRm+pQbsEKTtjGsCwb3ACJyUWW0zdLr38m59fEEHjU6rwOY9r4it/ifUiU+Xej1sg/UcEx
okFu+7sWEqH+IgH5RlS9blxPARfGA4Oo1S+XJtfAZJ6wktaeeVAO+STKuifCNBRYMPAw+Z3uxmjP
Rmp1vls6CXWmdekFqt2CN4Nke+ZT5QEFJqdggZiUEaCKyJD6/h91HA30dm5auRFw4J+nr3yuxM79
xl5Gyr+ibjTaDt6nM8sZL98gc7QEvCWjgocbaVYcQdP+kA2iirJ9bUAqumANnTRvT1ldJLIGjJMF
3Li+11xsdXe11P0bR0sSWO4bk8dEKOrhrO2AlbmOuPgB75SEL+u7BkKlMhOuQCw2CasSRnMYtVtE
JgpnQZg8ftVCDH0uRmABL2yC689I1dYDSVL6QIB9DjEKldNGIBWmIbZR79WT+gjLS1Lehmb3YPZO
lSDkR1fnnV+SPLUCHOOwt0nO8qJ71q4UrBgsFaK577zpXYizxpNpwLnsnug/PwWr2jfo3WZUSiQY
0LWanddO73ZXR7d00/iB2v/hTu7POcrIRtdZ0uuiRyCpY0RGAFz+eI7CGQ53Ov2+1GKXFR9qnuRf
vpbGvhG3xS+LLk1+44S4UJV7iF8st//YeAu4/0fzDttuaCQwwESSvUbSQegU2RbDYCB7L5eRgUSr
cOJy4QFJwRylg5Edu7hWMPY2+00I+orFHtuncSoS5MEqg+BIdQKMKuYLPVXWfj5uxx+LQGHjeDuK
HTTuRtedFC55O3Iumi4jVx3IHm6trwo0SXvibs1R0OU/SOC//gqtkVEetgnM80YfPKEGabOyCcFF
KWDWF46z9hscswGK92erDmeZdnpbpdLiBGxnYW/PcExuempvUgt7mxkFw3z/5WrTlZ+94s5VIck8
6hxgJdhZcts+GRCCSoelzbtHGwby/SzbBAkfA+1dh6pxgMy4renFWHw1ybsKuUGtqmpP3XYEIxL+
LM3+B01f421kDp4N0Dcoo6xPLGErVPySskr9AbkLKEZmAERvkpNShhhAlKaPYwCVmbMIqADds1Od
VPeJEtgNCwBKLC7d7XihfZb8bMxghlJznX5RIhXI9t8cE3voebUL943EVzBbQfC2rNVwruuQuta3
LYU/7HIHKjmVeAvDdV4m8aEgvs5rBuqnHhQKA/ZYfGSj/DQ+PgRSMfGhmjgubntBYb1Xxe1yKlUc
TQeYp6l3XOdA+SE87xZ6Y944Ki3xHcZ5oO4x+ZXQOz2XDkiKO0dZa4zThNKFKZdblGuqAnGKA8VO
/BsYDUqBQHXz3K7LK3OrXO0Pyct7AMTeAKDDAf13IQNOJzvpwyUUs4O68klWfhgBgKA+unb2gNcc
RkQw5eVssGS3kkD7jWLEURphAC9c3qvTaWcMNshiRrCbqBGRZ/C0OgUkZ3uRV8BkfruikGXrmsKh
3h1GLt/8oWg3BV9sPa5XLBS8NzSV/Q9ZjcEp+EAc/HC+CIlw0h3eNhUBnIf9+Bah3N7o61xnBJr3
lJB/3MBxu7AGCGMQ8Ina6YMGrEHEEwl1nRWHFhezQhxJQTXCZnsuLi1k7pOqYFlLEyC5ADwrIPIY
6GFIODfu7tqcyZ1Mnw3o/5ktPd9Su3Zpy46VipVW1YuJ35Yy642GcguBO9dqvqaKhg9ahTS3YrJ+
hTRXRHtnYzbNYEgu7RdPEH4MTNp/9mnVuwpXL77KF8tJQkdGvZFaNk4zv19mUIm6rb+MtjG6mTaO
qQNfsESgejUmCCb3YdgqyR0DyUbsbnduQWU+riPR1LCe0YDkQSeSDhT8ioq1WITX8z/eoVCbJyF6
XRI+AUz7PMbdwsFkhrIecCBwrcSHFBdl0RTZ+rHV8b9w1d1OjrlxntL8iYrC/mqvPGbobwLP890/
y3UNQ2bzx7up9ccvIzUb5akb7kPetRJqiGk2a0O+fJCIB7jhb9LrZhRIQvl9k6tw527bIntt/dqF
4hN8xQwlNaTlRWo6/8rPTNqdhIAu8JzthwH6Fpi8m4/7lmspol1l6uhuCAjCkydcsikmqnJ5Yrvs
CtX1dvQXLrebuaezBwTbGssRuUXCxZEZOCHvihyiXKa4Xrp7NuKqbXlZG++IpSGoCltLtIrARmPy
n3l7EcxFigpYd35ymIvDSLz0UxmYWuZo9bpW3uAxjd/6qCp8/LX5dCwZG7wanQnfamIYpkh4brfp
7z5TUy0pXCRWpX6TIIqnwKFX9KeuOpCZR0mA3EwXUrFY/icVkd+VCA8D7LIf3a4CdZjzeBHJS+8E
rwK2wuZS2w3FwGttlx1XGEQroTw2RVGCbGMi7pZ2yOUykSGzZvwIlhyLIyw1YcPhvjYSt2CwzmJ3
tB8o3EFQ8gzLbTkZ8+gmTPbZkTFarP3M+ATMyGSaS2ZMESmH376yz2JCesIUyXUoyUZRijw6ffV4
qO/msRryibOGhjcDGscxvXrqa5/CH+mftS5pHbJw0oSPAl2GXsKD23dxVAA8x+gbwbd5jzB1ZQIx
rrxwlo0dEGvJytY4prXsK8kGijRLMG2sxaSKB/QZxC5ga0HeyefdFV4f5hNgWgQRN5x5TmkkwwVv
tB/LdmocXhVZ7kA8/fzLf4FnpiWn9iNZX7SJHG3K6cIrL1haJ9ffl0tu7FHZCtXZUM1AvUFGiDfp
kJpr4baspM4OPNeQGdiWn4kq+02rp+MiihzkzIMqJYL02sFFhj16fcHh2MqwrdJgn3UXMpncdzPK
lcxQFzzMBTcMJrLDVkw5mg89m5TjLh3LNszbbzplWBA7CnmRYvpQF4F1uMD75pt71DLEZabUiybb
14yarez22QC0tapEo0Gp5RQjswro9v6IyXByX5NgMJK3cWkw0XXJXbnH/LZvfu/LKbgqGpfUWKrY
mzKZ0AdFuV0E/iHhdkuNL0YKKze4EDxykuVshNzle04XAJNPBqMZ+4+0BMllz4elUwJjtubenIxp
s7AY7SEDzVWhatGa+mMaIeT7Z4g6707rmUiNfVZ8DARLLn0S+6RdRZb/NXkAQfNlG+xLK5E0lLdz
KTTrhRwCHwugxoA7zAfxmrY8uDu1IMnKdGwJ7MDLasQTtJBaBj7X/K3kpKo71C9/g4mIl4GWdAPS
S/xsTyaohpGdmKcCw0aL5YR6E/rlI6YkoB5azSV94S3CAwY0uXTIbcO50sAtNHx9zPLnACc2lJ5q
kborl2MCf3jcW1dJ1tsrvvS7Fj8XuBU7HjtxN4+oLKv1cE25t5+2VPAJodGJd8v3RvA2CmwIkre4
0nKBAk4v3sViCpUPfa8F41uVoUxRaLo3247VVukSeSQc1x0zaG6knHrxdHzzz+ZbJfEElvizcb6w
fajyJJjjYyv36bjbnAI7OYSquZcAwcA7X7unXTT6jxq9Rd+pk3D34chxfIy7nbEyeDgTNFPOVeF+
CKwPp9TCNovSEeN2f4E2o7QFULMjnr/jQOdfM+eHszw1a6TwhHNKjc6uy1a3YONxEgwrC6usrU7b
jE2mejr9G2rRiPsdmXBddVu1M+8qnWdMUOEb5Hr8VHsCcGsbSu0KjwyuhD2iNZO+buzzBOT2ALPy
STcKn6wbW+V712KnbX60b9TKej0vWFH1IPHRbMwSM5r4o6/zMrnkhm9Qa1KH/273K6KsNE7Omqhd
uYf8++6eTz6lFFhdlArzw67Ai/4zBfxxj8VjkM90+2Gua3CLgvtFsc0mXTlbiYt6N4zlmACv3e0f
1WI7OXPq/UC/QiPw+sPJy/4U8AqKcktLVeS8KurvhNXPJzeNhJQuk7d++ywTuBFZobLe3uaE7OQ9
8G4+8xhLFwCbkKZv20UPi9Ya+eXFAJkn9nIvCIjuFefr9lwJb+7H1Z9ePv75p4zioXSW2R1mNsxy
5FS3ooLbgQ7ZyH7Mh3G8qXqdaJclRK/pRIc3D74QUjQlK3fTwwE/5TyWYW+WXjJqWApgE9m3O7a7
8HvwpHpfExGFFGlVl6ZDObhihpY/sS60LjKGrmItYBoO2rckqJ8chHYf9zCmblMpHSjysNqth/E5
5UskYp3bw2n0eiSzGIEtf7rKXu9mOhxiIIOoWkfTnvIZvqw8DHBD+334ttRFHcV8WwStBOzs5RTC
uyd4kpr9aMPhMHHA5I/s3H6hSDr2O9dF/gCVKxJVFZf7LytdYkUdrFIlK3l1yddbaeKdqzTYfZ3N
+DhVIjmNxwqh/ygVnxV/9dNritgcMkYPB2n0pey+jjMABTw4vI5F0lvdpVsMmNQM/g5A1aRvJXW5
+Fz8mBBnAJ+3hatV6++pou26jswKtAYq5cGNWW5wVcWs9H/t1b0PMcSR0rprI6E3Fgkm0PbbGjs3
MWPziPxbWJlh5YBHrf3KUMysYdtaYlkWnzVeG/CQGCgyxKfBrSn+wG1Mf+MRPm4ZMl6pYTRxYElM
Icjppbqx0yU7iPicf1fKw1CbK3KEMve3CslEmJvucSfy4rPUmgJhgkMuIQMULJfqQktwsvx8YCi3
csLtxkjXrp1apNW0tk6NjTKcnX10XJBUdgzXqdItxe7WleLQgQwO4nrVEVDmS9id44Du7lV8+Cdu
noJI2vjHenazckflniDNYzckseZw9KQ0tJ/0mytMbaCoYhq9QRRdgjQhxlQaO1ZgyHRzcQ90ldnG
eO6FMvEp83AjGuBt9H+/cdipEnh+MYI65K+PEAu3g8RaN3kCHdHWviEEazhoAVtX2R9OUjkGKic7
3UtWRWXijiy81Vq8Cy0/kjvNqLk92w+6NQtgHovIhEzdWUsPEFsBj+GxiCMDCduM3VDtMfFmJgmq
EPeNPbnt34CO+zqGXehRrrzqINI4diWoPNBP65YhAZvI81KsIPkkVChlWANc3KcTy7fBw1CKOUA0
lltud9calkrmSBFjA2Qcug6g4vr3je9T6Nkb14gxqvoubGggiMSHXdBlZksWbw8EB9Ou20EXZYEC
0rtYarWHcmu/nzZpm19gvackj6U+2PkUtCgUlthaEG6JHwPax3IJtJGobd6Uq/hjYNRFgoAk0dM/
+T5ldoW/mZQwPLFBddyo7maVyM9Wy0+7enBA5v3GKQu5BmugljPOeaButE4wBwPIzp1G+N5XGYCx
J83MflRNGnLO5Uo8fJRF+PFMnO+cO8/Kzy7y5tf5BmAW6SqWWE3ebAPf/NA+hd7Xue7S87AxdHKR
2+x9h7Jhg9HAdb6B4XtXbs0kyh7xsxH0FTx63dMuc+C9C9uU2lY2dJ17v+Laip5pjrJ848LzQ2Rh
xna+s35qak5wpZWebYV9+y/6yhIbLBHa2jEa8QdGyD/XRyQvEx8WruHOxMEhFQ6CbGe4oigtaboO
c7Bz8jJme3/t+6NeXeWItgq2x0KfMktiHHUI/zDCrpyJfpoJPyzeAaEWfCIpff+I7qL1X1PNPBX+
y9qUpj+lWaAoLeruW9HXzv8kxujZfMaqOKn7qJAT5ZYThcs1Z91HB4gr6ajldXPcNVeEfKNFLjjZ
BaXj4zgR63KdMc9eTmTfrH7NorAyFNc02Cr1RfTtcJS63D+w3+UsGQBueegMs/BjkDeTmkTM70IQ
8bSdKbtX7RdcmX/3Hnl0OAVq3m2ha7XMPiPBCAe/eF77/kbLtxz0U4FI74BuiXSqIanH7fZRwL60
ulWLq0Gso9o77AtrfGQrP5fV7mG2RTO5icsijZZvPyt9+OQK0lxyZLMlL6XJLIj3A78YrwBn+q+W
9dz6PudRb8dFdHwyuxTyRfQ1HqPktACCJrQXLJpqf9FRzKjUWR77swQ/3lqivmMS1MbzICH5wloo
008PEvRFYQbT0m06KUotXdKce3faM88enluKpohGvMcubJRi+bN9KX7NaWgXGX0AL85+V9JM3afA
n2Qp8yCXnp4JP6x3VbJXZKjQBIkWkeh+m+KB9iDoqh3qr/t21NZAHq93c+1edTB8eBrA4GnnDIJt
AaJEzVif8MKjv1Wp+dWSLh+fTKkCLxMYGIMIGdkv5Z3TmFDBvXX+ExdxNHRSNhopXexSpBadAaiB
0qemc5063he+Ju4j1S6mNWXuN2k0MdPLkS8nqt6ZvxGGolnhjJtHdLVPqCrb+v2X5FDvw8cct/SU
9xlkLrq/TsYxMDlVLW7mFUmEZNn5TZ2Jcxt2JKeI1U36wiSzK2aZbOoeWkbOI7HMilj84adjHFJm
Vd+m4w45sQyZG1k2chvNP5ebzJ8YLQWNSnvNygq1LyRtSGbkmyDIShrKtiDC2mQJYF9k6UUyZyys
MXPjDzjgCZ9yAsp9LBkurTDZoBtdx4aIn4v/GGxmMV4uAjGfBpEuWthS57wQV90WE0mYyUi/13KS
oYKtMlTKUfDB356c9wDy0uAtc3mNEi0cFw1BZP8dKFwly9el3CIf7Hb3UqG2adLUxPjl91iu+S42
ka8zGPuRRhk6yVJWAyZ1l3uaeSkC2oVUZLb5DdgM1SLhXVPVLDKcDO+AuLI6jc4v28kJcNJ4hH+H
ctX5AQV0jdPcADvUGB3Dj9khXzl51bjWD5RCcarpIHK9ZC6iNMmIN/nktl4OovdBn6IiuqXAk8My
ZVqA2YgSVC7Mn64DKvfzndRDcMlFyGtP+F1YqrMbIl2ZJdBuPiu2zUvIadLqCtWzBkU1Mto3JEP4
LeeGW11DtdPjIs8L/g0W0NngMOWZ/u64kgP3+LrFvMAIKpQvpHaL4dKKSQdrbpH79jtUh4UJgK3/
sksX5hYLpiopZikJfluXbH31bAtGjoBZxYvZjzviJm1x3E9ZS63na4lAlvhmD3viMC687A3aPZ9B
xVFJbBWyiL7uVVcrG7Zla+rKLgqXvVRZPStQi/42LiUAzQPgo6aC+Au8lgjdidvUnO88981i4mRX
EvFDL9XlEu9LRzcICXqKVoZ/e0QX26DF8h5RGo0ZfGO3oHaYpcmtItgw8Z/nnGhJbqog1DV+I+Tv
JLVxOPruTmh9D4I9kM3lehOytsAw6eBwaRpFJsvEOtmH/N8JRHMZ9CpV0XQ4tJTDnt16qGyjxDiu
45pdi5DUo7sUfDzGe859VjjQxVDf09KFyPUNMaw7XUuGfSKJBrsnqZaqhUIvKNmVd/t39AsuYw5s
q/QtzvOODNfsmoCj31SjFxE++gTxxOPwI+xGkX8zjpCMj5jLkVonRIABiRoT4SmFXP28OYvm5+YL
BLs691zb0GoS0ODW8mEwuQghU0JDiaClwocix0wqYpmyJSzyEc264UCbRYdgvcZgtsR4RB/tybaE
sZh1fjJFPRYTuQbuTYNltuz6mJyL34WdtEV8DEVQr51itS+k/VX+hMAY+Kz9d+61Ad6wXXc5ZAEB
lWXf+SJixTc+fM+hfkUdbtq4BLBjAMCQvTbGgboULB1R0PnltMD8jEwAXI6nOn9XDS5XPXNqR19k
FhhtAAMD9EbxBx98ae1rcKH0BfO0TiBrfQOwBfYCX8V8bODeHruthMrkF40hGnuPej/pmeI6mu5e
uARayAgrXNppUpFXnjktEeiJKwKtSEtqWE/fV6xdspgO+TJNotubq/VEPnQ6UfNH7y2BOF8+vImU
ONLonsTFJuOD9Zi1xr/2q0J57o2oF/uPYbj078cvG8/KZH/fbOid0w+Mt3QjgmZWjsNBQjo+Uub8
AJ14SKvmk6OMZM5/kAbx4/v0zyNnHdkKEvoAZp39YZxtFxqVuttRc2knXrkPGjvScSwk+9EYU0vl
tbMb7P8ATxCnK4go5Arfzy0GbaSAMrqVIoG3boaU/BT5LmwYYXRtpsBqcqGNEBRql1SHO0vurnLp
m6l92WH3eoIoxXTICW9UuwdVtFarehh79pFpemeVI0b02xdPA6eYyY8crnSu7lf07oxTN71GNBpH
mDT/1AMCLz8yerOkRyAA2265xnRyh1SJxF7/XwojeOD+XfZ7YXHATlsUyYFlFavPUIodkJ67IYhy
J6uePnJRcUHTiv1c+JsrIKFOnsBbSmsSfqX0INXnyzYF3ipWcWhDKv8Tmb1ll2TcnqV5oQ1vj3pR
huYCrk9SyWUQ2EFdTC2palyc7YlFnltu0oiEPc/IxYwuy3Boglsc5YeAQcXK/vE4tQ5yF8YiAVZY
jfvdsboF03miRIb6BINo9V0mqu7kjta7FbIO9E6judxBSSQYI+iuM0udkaN6GiIgzadWYsiNXgir
mgYnoOo/9SS4ilPF+X1641fEEXFdFUxtFFxL1GRHANg7onOreGgXMgDQlxWwAC4vH4rGwmXkOMzb
gM4/TaUC3HhUhe5FqUOayggxvpEZZ7IHQ2UhPnmiiST8fC69oSLYEJkXpntyBCHpdQR7K4S9LHmu
lJzqB95/mo9JfBcxwiDaD4DSchcMAekHroG3IYcgxPFrz4Ov2eh42qDEoMfhjciG17hPpJi8nZuW
2yg7q9W1mxqLZhb8hR6FUe98vgfds4UzU4thnn142j0TTkpX3ThBc3EF54TbgD2NRCrdzsjn73JY
QsNkZfgR5+vtz3dBYL3mBJxsmmFqi8aaDsgMleHBjP+nv9awnxT60wOeW+6l2Hb8qq1s8FR4xeeP
fDqcM2ocS78AYkrbGHDoT/k+a7PgmH3M1q7cS4tXSmQqRypiFSewee5lmVSFFLvC8WkTMsRYGfY3
PYqqZ0eO+LT/36VPTeBOZIzkezMvRJkGL8xDioH8NmjWLdaLVgCn2jxhd2ncwn1a4QhnKbYqYvsY
Qx150t+xrDSe8OiML+0QLy0irwD5z7GcEr1xEZ01vl45+6JuYkmaLxXG5NrSp1DYwIlkHJmDSw7A
qglG9gqGrTk2KMvHSRNLMK+ea0tqzWLL0j/PcYTiquqLa5OciGBZlsOPL6X5MwLNB2kmkiEIURF8
k09Z5ape/julYpwgVoTjuJOU0A6eFPOXyL6jF7UdqWPzwfb9fcoJlXWNGFb5KaDUAlSxWXYVevst
2x2Ur2mn85WnY9OZ3TbsTI0l8iWT+L/fVwXbENsLBE5GfbwKobgroQRCc7o2keNZgpr6FJG/l/OM
f52mAcWWeYVKPLlrd3ybP+w+roxXWhWQW2ZKDrKn+YjoV6ihq17NNp8EoXnCKc9I76rxem0YDkMt
fg6p4pHdp7+CJJjp87YvcGA+s7fSow2WEnaG8Vb1sXlUKCfm5/oZGAKCOtuE2DVko5wkQDG0eKbP
DAJoztsXPpUrJY64B6zjwPYQEMXGPdtsh0VwC/+tt7CHqbZoAg0TOZLfK4npzpOQafSwbvwmoHJz
3vTJCMgUYtxpdsytsHWHrFzMwIxHb4qgEa9T0owRcE5G5rPcQo15vDhevEk3RhM8Fi3Wj7IKvldM
frOfVJf0CWfLVbP4/J2WkTQ8/XNcnceVY8WmD7ct6mfHhmB+kajPFUoQjiIDep3o7QikyutJZcpT
yGZ5shmy9lhvoSshiUrDjIR1lMWksV8OwESSxWNBiv5HhwdslKvGXPV1pRbCHtBhtfU6NTwvu3v+
SOQXwlMou9ZB5/u36/Kyn2SMnvn+mXKqE7Dx3WxTZOQinBIHL/Ls58eLn68EO2vvn0mxgFfp5oYq
HZYEl9akcNfq7JSoja7OcPj8RWO30Xb22NVa5m6QOJH1A1eQxyTaAETAHd3e2KZAlb6Ts74UvB7C
m6WoB9w1L0gt1v+9oLA1/639YTwBiHJXx0FJwzFOIz5mNPp2vRbM0Y+4UOUXUZXovxY6A7qv6vj3
DPpq8+orkmBUZI7dlr91c7efAdmuv/wBluDOlh8p+DrjU+A4PHV1Bf2ytnICtvbftn3xiEaCfEi3
b1Q/tHU5kh/Lf8v5Uisy9ZZ3uaPcHcUsPrW01THeelzDsOaT9FbaHKseiiJryMa0DUuiYOKo9R9Y
zpLKktFkxhtXRtkCHE7w4n0+Oqj1g7PQe7xDZtOG4UuOo8idyhRxOYFw3OyN3v8HkFISjsw4jleT
TI2aTnoKH1APNpvYG9kq0sUXeSQPtVpmHiQ48hHBS0r+l5bp//ftPyf5mEnWCc4k5qDkdif+dh8y
MrftxQOhpvswLsi6qq00jYYBy5DrWPtNykBIq6+w90x3yr8HczMo8Zy/vthvBdkIpohMBxtDyaVH
wxKP8XZfPr5RmbnzFdyEYkg3wDqxbh2Qc8YmYI9PA8m2U6tuPyFLX9DujDvK0a0vAY5Qvkpu7Xmy
Q2+0ONPXd1woGLnGVhejgMUy0LlRQafEMzvgwDwbgvBdRKhhpqGxl0cEA01Jd5a7lhcPShw1WWsM
rW+fu4jfWZDOM8reJbMqRjPax+jIgF7iw0lj4hzQELH7Yqef6Ds6vMPjeeaA/AEqstN8SGNbsiRV
KD6/IEXp9YQEEVv7ZpADikcv56gVco81qLZoHvH3hrC+xry9ItbulnRbY1qCYdniyTEPyQGsPIzk
qXbPk4qARQZY1JjJRaLd5D9yRfIcspIhMDg+iVlaFMaRdgx3DS9/9/wpZuJEGIqhbiQACCMlKZqa
oW2pM3D+quBxgkSb3JV3o1d7TzzDBEmQnZmPycKu7HNNmONgm/NdKVx6sd+gtLh2JT5al7ZGcvnC
D6ypn08Y/2D5l9R7iLK+KzNuptKq6r1F/I5M5IkxXBJfDJfH4ZtR+o/OuwFZXM9ZvGx3mLz+yX4E
ZjM07DyYY7UMtVGtuZbxpJXYNDVkxO4FAxY0UW03mncWlR0+0KlPzsWpO0U74obPcTfVwwJN87xt
gNbTScg/x1dAQDGs1amkgS0eQgs47bqpWMGSIhZgBt9PNGrwpCD7hFp/T5CWHUYZBrFAIXVO/B7a
BvDIJyZBZ0oadnKR4B6P7A7Ntn+Tq7B1HNOn8ZF3lyBiSg/gvoysSLocOstyzRnXwdq5bv2SEoK2
YJk6eABLfjE5wWjGef2b1SKVlJ34QJjsh+NqOK69A53fgDXXqxyzVG76d08KIpJ9wTV0W4ZBogyT
Dr4lq5S9rRMsbStqyHWshEr9GXBb/o34+2d2FNzXYUBj1i5K7Ncxy18j+oHgElrJePcPoSZz6kV1
gLliIT9PnbVv8cC2KqmiLQP5Ic3VitVZxZGxpcYUrEEoTecjpBSw+l9oFKtOQIJldHXaVB0oEayb
akVSF1QNt6gAd01C/niXDKbdtzhDSgtp1QpIX6Hg0jmMGHAuzWFEZBS0LLN/hgSvJ0ovHc/u9WQW
bfQMkFTXM2ez7RG7U/k1wnAg4gEVBG3sEWKFgTeUXvs4oXlP8X3ykJv1uUQp/fybqJJehBRnbzOi
J20uJwN2HQKEtgdfRGAe5p44VRJcatyzmWdE7eY3b+poxscdwYUAToMRXEKxk/PxBmjlDl1VlFqw
G67bWgQuZEeXQzdMgXn8RoTENmOmMS1ShseKghYi2hWaNdLYhiuK0MLhib8yiNjxGxs1fSyZS5h8
DlHUluoy4hvfFD0ZYlwxtla8zmv2JyBZPLhJOI+VuMCSkc2h1xU/lX4vv6YdmFOCRwoQaZWnb4YA
G87rXwsyI3sI6SGWfNrULwp8cmzYSpgsjBzFMX4a6mRqpkXVqCa6ILMPS0YCvcSpTskwfuptD5/E
il219s3h0WZP4mMFmsaHHlPIaCkOodl7PbU0y9T13CSm8TWh0IEm6PU7DlcTWBOq2X/WEsebWhy0
lCJKaA2Z1Q3mafbbJDgWrAITaHtvNkBdjmjIjkYUgSt2GebTcPzI59EZvMc4DxLJsJFnuOsXlK+5
V6Rx+giS+tYUJDc/U02HAl3TEu0I0Z2LRYQfmsvhc60xXfg/ZvfkugHf4MeYhzCpFrTuSsoLFrmE
gz7w6ntlzHd1GGA+TuFrwp0Sw69s5U54dNRC7h3eUxTbuzbbB8+t0kV+29eK/WcTvCwLjpCDzmgR
yTiAUt06e125p7Nl6+hHCeXKA/hZr6tyem22Cg2YGW7JBaNiVviBnWgDZxCYRezKmXKp9jMFG7Qg
wOT0X66zgeDBv6HRZ+u3VuGT33j2pYeLVkMuWOOC8IEuI3gGLg4ZUuLfJP8lG4GefG5Enrcrjhcl
W50/XMsZsMYkMjUWVEUscWZmP2OCQcyRsXKJgvpS6nvhn5oA9zTRdE9hiihOIgiOwWdbspoTE4Ob
FSFVr5Z1QTiMkE71zQPcEAiTM/RRIE+IXiv3he29o3um4hTKy4ZctirRn9SdJxmxtGAy2bTy5x9S
lVTGtOT9cy70m2FwpYombh8erZSZFpRX+Q8edZTbCbvSBo43ENotEqUtkSZGXxCA2s3fQTIosIir
HwZNFIxjuXeXV7WAiG38rZVCSLk32U9A4cxBw4cNopADumdaC0V3W6fIwN6/j+bRn/UZjCTRv2gp
0D1L9VSuNvEVlh0edz9f42MWOR/PrBujLSF9hl9af/La8ttbwPOyXWBUqUXJ3cjOOp41o4Lt5d+E
Ezcfzn5cMJNApYAWZ9bOvNXvGCVVIGqPS2fHwwlQDb3pSfotoZ6NcMQNb1pIS3+RopQzNa7xBIXE
L+8VUMSmTIuuRcX53cQz2ng9UGX3UTGAwdxONmgIzjnQhtzJx/gUhdoEsxudzOxrW0xwj9/nOfsL
OUCGpesXoVXhQ3ypbqvD7NGa7ov3nANdSzMxR9pcetn14yixJ21VM0cleHbSXvs6Iv/fwkJ3GOrv
+5LjrJrf9+PNaGd2A65sIxMvZMHvHsBHHnJpTaGs+Lc5xlrLL8lpKQ7QSWSM5JnQFDqM/KA5y8//
d7UQboKj2RZ7ipV6yycDs8zsoG9HoruYoJ2XaOupb5PRUaXO9LmKN+0vBZjzKKH/XuLTgDMs+OaY
VW41uoTjMcZFPuFpLbNDrCD/3T/1cVadX04cdsapbWJ0VdRzTn0W1V42uXyTQYwdg2voULAfZ56U
4kUwqY0VcX2TJ/e5iPzLbdb71uQ97jvaARfNYNh2GLMpv0vBv+OdJLFTlsW1qndOYIkyxVmrttVo
b0YcTSTT4twykeQj8iUge4aYQE4wD/AbNqOfhzk2CzACmLoDGlbkphQByPGjgXE+xj/8dnpjtzE4
nS1C5k1AZu9UNxQhtAYOhLFwkTsUOVAbeH/IvDM02qBxEbc5RzsB4i0Cfqqok24yubcEEySbD6oe
LSyWQl7WXeQlADIHhbQ5oh8lsCsNFBCzppcmAqmENhDY6gjLxFUuiiRcpHtODR7pbDVEb61eR9es
gz/LTjKXseV0tp2tLxZPRoqNYGsn++6yp18350wTtXNx9MvwTSK76QILwgi2seFOKOq3rfxl9cHk
/uPkI/wW/wyf2VtUzq/xlHHJk3EUd5wRFb69AoJNuc9esIQn9GcDscNDeViH296vhmccPGZUhzsA
xtRHCti8s2UWL5B2mpCYpkkaS6tjckvkkQPplNkHorL//oE5vbLQwJFOH4aIqkXnDG7DuuCbwd11
i4YydRBbYce8pN+4nHbnpbQV9TYG0N3eaMBELfk8npAVaxV6z1Yv5rbUmguCr0HhBPoBHwcSPwLJ
sx4GCzum1F7DLhvBLtn6TcVIzpUdg3IzFhJ6Ptg991O5yruKDueRWwFMLK6s3zzDL19tU1aRQgpg
CkjabPAipAK2MSvarln9an+Wy+m+p1TO/+umW4DMAs/KSNboCbmC/xjASMEKs51lQKe0p0diRFla
EKhIk21hVEW84Q+m+JbA7uCBwkuT03yXoV8RO23Fi8XzIFH5kL92dgPkVJ91jzjXNo6CvRN6aIbx
+xW7Mx99Hsl3eBFnGErNYoCTzt2ueJBCEdhXAgy9cpjHShMSSkG8mCwABKqtXneIdZSYsVqgHamC
1HV1QYVEKsXcYDD5E6rrtnZ7/LPJqE2SUcceRUohf30XhoSSUx5JdHUQYjiS29918sJ6eMuCETj0
CxZKvWAL3WMeBGTctQeSUc1j+txxwu1dGqs3hUmtn7EFtJiLdnwZe0o4+sH26yxbf/r9djmeWOVE
Q8KUa+iAMYkFPw2elvkLwPGsdvoLQcAXaehqOTDtnOuWPjpQj+JbKb3vfTvLQJcFstNPvLYqvsTB
TQKZjrx1IzjsuHh9dA+JjWpv4yDG+1mY1BO3cPsXrqbz8Uq4k6ijs2L+/RYprKM9HsmtGAEcAv4J
6rCRiDl/sa/RW/3IEcnfrbf8qFOgH3JEbiJcish023EI7vJi7H4yay4M5WleQD6CWOH3fQjuHsF4
DA/C5eLZNAmbzZfq+2tXKJXL2J1VbgJHrODa3w10OwMRFCECX3M4Bc08c7jB6EIxrBuwfpgO6lyM
XlRvzLevJpn8k///t8Fcl6KXGZKQjZuJsLrLrCKu0mCi/W7bUYDO5LJpdhxlKqaDA5horFglF7+9
honKTCjjKvKN3vnViDbSXxs8KUJpSip1CRTmGhh9z5iVDvdTc+SZvEq94LMfAkQydC/fMImASQdL
CjB9Dh5vQwFU8qr8MD3uIt69BBbU4jfF8ZRMSuMuWXfShQ/UiVmdNZnSDEE1DK2X7OyYbGn1n0nV
FaWixzKsqRFF3a01GPe+Jc3LK8cSmf5ooUNk0UGS3p5l7MKc46EkPA7S4jAQF7DqYZUGsy9dN8c9
8fcppcCwJ4wnFx4KST2bJ0kDgyIG7REE4ekpB9C96Hq9US1OtMJgQxTxlZLL9HqGQHjV9rju61zz
JHbpwz52+kl8HhYScAHbra0VECmaUSRIZuqoAU7w0JL+As/rDMp1XhcxUX/FAKN64d9EXSnPXzL7
XAE8hNtdQaMxbiLUW4D3BUxVIDm6B6Ij0K7Jgd23eBX5XsNVv7TdWdljwdlnr5YQeBcWeAiOPIny
aP/RUPWnl6xCq1VVmOE1v/tPg/1/ufF7c4McgaEcRhzgkOGbmO83cCPrnntAX3eSy39SYk0TiV+h
PMo0ylDcYVbp7ByH+lOjB/BCDAJfzgxbxAFy5qgoJagJ2zTO/CfR/SvunDxq8Vz69Dul9o+1PcjF
CZ1boJOMggPbou0s4ldZnkpm+QmO5nQ9qX74XiRns2XIyaJU7uVws74AqThFg0mTEh6/nrL8N91W
R4NJLVxstlzJQ2h08irBBCHg2/pFxlhKpWS+uhkCn2t/B8HoWk0e1BzgO2V7kI/cop7jgTqSHJAs
jcQikLQyPJN3az4eKMN0o3tEC3XKJTDcVjYYeXUacas72K6lXp/uC9WgZcfbnYi+h3GQFEac7Yse
Hb/OxvG+NJh3Ezookmao2njM+rIZINTe6iz3XZk0eepmyPLs8HVg8N/9L6Od77KNcIeA+bhDnTVz
JYYDyD6m/sFQrjkvi6mBILuu0soLm+Dv8ezYZhc+VNjPmdylaaJVm6zgc3I488fg8CgGukJVGRCJ
sammDk5n8ekWzHVBaZZjm0nHiX8cea8dOhtrMyFPgphJLK3jBtqBY0qT5GrswNKnnoeSKl8GnhGZ
1/stKsj6USKUxayEoXBv+jpYpX6rh/Qbj3Udz6j2WM9q5T1Rm3UhluwPCJVtj9mk4S4o0eZL3j9s
tbRgRzD6St+a7x6s0+W93YRHUYyk7N2rYjP+AriZZ4FEsUiZa/bmqafkT6cvDVvhbHmZdBbIlIMv
bGE7QdOwRADEa1HOM2pnoAvFplk9tkpiK7U+lTAPYk+glI9n/1GjaOdJ38qvrUiXX6Nggj0479Nm
csLKRGlwvBiKDUe4EWoWd5zEFc2e/fp8pb/QNTsmQtp12naou3RojggP6cDueKFlAp3XwG8vJyT+
anHBuOgSyHn0T/C/EFUGE33eMgnpsHm5RdzjjY6S5MIlP0tWhFPwQ4oiYjHf0S+ZvK0u330ApxIm
HwNS6sn+MtrSm+oBevSzDYKxbVOfbh9KfSPXQIoweTya6GxVvgplN0hlac1j3DwrXfI8M+MSyp2j
IsjTOnt4zvOGz1ik4GgOhJeARu4v/9a8KOIDQpZUAVpzX7SBDYIjUohEouKiVQUOCGtBY9j+Ngib
1gqcABLLtrFOf9+ybFDHkpRQztxheA/L3KPIFv4RYMA4n7kXrI8BHBW+4iCGv92ttgH58CIfwPwC
p10UYzY6S5fzdvYFiEgNLG3QNFSZ9wgfTyE338PWPfDOX1u40NNZX9bgZBdLc6ljHnnuXmeJBXQR
fNZ7mFGMklcp/CUGqluzJMRkmgXcyj8dX+1ZVIaZZrU+na1lKS3jUNxC3VhxDRFdfQZfRcUduHUL
KBBV9KWA/m4m/kLBYkLrQYDTevg3TAUfrPuZWWnXlcjEXw2kaIJbD+r1ju0CT7qj68LfpgBHnrRl
OzzPemjZBy4cB70I0r1h0/rhG7qCGkUvZrK31RLBMNQV22Br/eyjI/FsKNgwBAnaJdh1Wfgza0Hu
NM4f//1kYlzNISYY5TMakY2NBle8oFbB97vpqhrcSNXJkywkrbavCC3xVBeyQyjNwoU3DesrPiBB
eHI6hpgCBHMEK3PMDv26NYeW690LYPd2yXNJTTFMQNmI+ASXNajAn7/GRsDv82DuRkuVYAjMF5n7
WNesbWn1+Yf4JCnjhmcrS4QBmoe/xv9nJkIWKhFXrxvsPfu0NZIaCHjUEm6JsXItklbmWGMDd32z
L0FWVZkJtUnbqUxaEtQ77xp3/NzdekTxMII9jaRrTB9cjbRASVTA/SegZ6AZ7P+25DygolXeE49+
m40QaVWySxuBLOA8vurNEX/0XFPFCA88ReMdOlDV+RCiDPbm64LRPiAoWXu5wohJX1PlFjwnsMxb
qr3nAPanwlXUNd8Q9HNdUCQuFuxvj2A7C9x5sp2WDbt9wQdiS0b5bMTRURZuwiGJS33RnQCp/YzF
Q8gQVzZcA9D8Su+/gvVd1yBbuOQy8xrNLhXRJRLusHH0TpyOIznxe9b8iZ5JlZyxcbAlvDcXmI3F
ncHahoPdqfURVzRyWMJ5Fo/5wDAeCFrcrcuVffHc82hfsL0tsKBzTtH/nOKZEMyy5U3ZgkngHh5l
yEuobykL6h0+O0FXLK9jkLt5YOThX0SNcIK79J6pzNNDlDYNnsuHY1h2LUG6yFrqLWEM3kpoubqS
Ovd51NyO+98iI/s3rwn567TM3yo+PDi+N8hC121QfULBm0kTsu4IPEShu7mrmAGMZzx/F5U9J9Fb
cagDN/EC0fmhNtNUkGt5SFfQcKv7Nb3gfrGfKgiJFfmlm+JZ5M7Cn7uzbChO1Jjxzm42gIIK+rfn
u1Om/+6D20jBgHtbEw5sy8u1lJoBF7t5DnHA6vIwvcPtf2p+CrIXlIldyVKAfVwOGDffbArD3XSR
r8Y88ExMNwrpbZmQBCeraZw+kyfDJtsiQcuc76aMtr1nWbsVcto4vwj5VOgz738g83hIUh9QGwcu
D86Cpd/Rqw3TLjQZiSoIhmBdYizFLEdBLnbr/+QCC2p35hSRfzztrr8snryCl3Q1uf1uoprksRR2
7tILjqKDbszIV/q3C7WDmhaQAjjObgD8EGc4YPUu/8nkcoRRjILsifDGxpeLB1+a4LYn7tHYp7ui
ACRkEok2R7m0Br04Piu+5sA9R4oGUyAD0fU+DUfCatlYHGTRS7kWMlj/xhF6wHZWdGqiKU3Rl/So
rBU/rIaO9lwDxy5bgx/zmieEfDhpuvU7jAfTr3uW+MmvXRhwxWTLFMFZjLHR6MvGI0BTeM0yjMpv
Z0eDgNffCF9ymtvW06cx65btHofM3FHS3lCIMbJ6Ge6jZgb7OskJFvEJZrfyePPpvKLffl+z3s8z
H6x53r0CX7URtJ++vlF9zUP1SQ4qjbbWsBejKIVMyPDW6TlDRpKpenyDbs5wQXzjIELTe0UZtcnp
aSIO0lXja+YeFwoJ4S5x1YnwSnbQeXJJyY3GVs3M7RodemRtOvtsmvprGvAQ4KCXYr+eOZhM4Jae
P/YAOyg2bQbXBfgPgVKXV4hk3awv6NEP7dd36Nc85M0E0qmEzF2cdmAiDkqIPeFj8UFtoBD/6eQu
7DBmzIKNaKMyCvFr2oVG/rV0kVYOMdnmovRRFO2tW8v5o1cUyp271keCY3+W2Q15CcBAHZq9bFkE
E+7XDEoIx1pM2R0mL5CgegaN3iP+OAgu+VT3a1SfmWRTp9Gufe4J5IEmoM+9ho+cS1hsPAIF0GdO
W2n0mMC29d8RNN2luad9Kbil8hczqY0/N0ALyZfmSOu8E0OA1eMF2lyO+4y5gYAJ+rd5BM09qR6Z
lS6jgO9XUqZ3T0MQefDGeImviXOn3Ycwx3lvH+09zFI95ZHWddlz5oFYrenkgGX2pxdVmVeEwZ67
OkDsKTr6gFvgd/IHxEBsKCioAz6ZghYGMe0uORkGpCD/eC3Ma39CWThZ1EEvNfGUiHAAek5ox589
/u4pPqL10bbYVtfsJYgF3Veoiba7NTBPTQrZd4he3HaHsc1ZPUegRIn4uaaox0vHI9zyevy8t3Da
8gP0lCiVcCEHCdkQxbEJZ+EwT5LxAUL0PayJuNNxZNaRx1KRkJUP0WcxDuur7EYkDX9YYTXjG5xv
mv+aInAv0C2B6d8vCLLNfvmQ1QNZbPGSu3aBUcWq2h1W5wTqBzjjQppRu5Mu+rKzO4jq9/TFMvV6
fZKxMZtTNmHgULQel5PR46c+QKOFFJlwaXGUwDhCkL/fvpxI9ukZWG9A6deWgtwgiuQetcpzTORJ
ThfydZ8lvndeBu03W+clTu7q5JLXTQEzqvM0Y/vzBTqS45SACKJCuPVPgeW5FG0rgwRQYuucG4/c
Qy9QJ5pSbhpElP+xLMPNVZVyyn9F+wjvqU+X1jKspdKWwQm1G9iQI/sqf76cxAhOB7yfcwC/szcm
e9koWMpsv6o9lkONofy78bgYDC19bRu57ataJmf4E3t9NvZckPlPVZX+AkVplUspZCShhto5XTgK
vynbzrTnijUx4EhkZnvOSW7fBu8YntJ7F32JWvt1n9VvPbjil6CfXiul/6XAHG02sp2ifWjANyzP
Jb4JyyOiqV4TzH1xnlkdkQ1X5mlSkbEo5NN0Gp4awWHIjR7CzR9rSeVEfYcbmPcsZ2dLO9XbAgqW
li4E0OA+MIoefnosPHFaOsNmmnzJIfOViEImyXeKRwYqKRgSbBi81LDvFwKyEihybaog1V/vQV8p
aP0GvzjIz0KHxkEFyRp6pf3bc57QeHCSN7TTn+b61bcTepGoLdnkSNhmRaH8qpzCMLlZEq4uhFEP
5bas043TSLJolfmY58z+SOD3wCTbTuI00sqF5UKaF+QSZwOYP4HemfPFEumkMcbIKwPnJunMn0LL
KhPt9NJ2C7b8vIAOn47IohAxDzFA733TBPVYFk5xcI/u/+yPbTISXFmg1nUYGmgBKvPXvKf8NJKR
O/wcylQELHkAyMpwR7SROpE8/Ej6Jj5/yvSsRcat1RwxY7osrVVrcbmHJoKssN1H+XmIIFAqUlr2
QrkB6NqFgJSb9IUsyG60i+yQCLr1QiOI53ca8F5hIoh/Tp6eWE+QWbS8GiZhr7WbBxBARvJ4Lw2J
bw0FTqaBc5gUrj2W3MGLJXXXZ1qHKbAbih7VDYZ1DRkzQDGgIGvIoJHoKSFzLBZ5MpB/I5P2hD9y
CHP/qrTc2c/iOurxjjuVBRBqR9b0BLFeOr9knfiJGXYKr48XUMHK9KP4C+rsw1hb0MAetoSnBiVc
Rcpw0vvN5jYKt5sw5RpBMQO5p5eng9DpdIPHzAJD5Qfq1Jrsexjyut9322ue1xt9IfRg5E81CiJq
f61fIE1PVq7z+V1OqbZd9xR2dl86VeQlH06nK0hATDQhOwmnkfT+w0cMg/yCLiTZqo2Vj0I8PdLj
xWMrSy0a8dw3WzQWKdodAqw0npMYqafn20NQCsjst3yYoNjWiR6oibDJh0NXaWNjB5XnktHKzuQm
zwKxeE4kPOmG3GUQvBrpzFJo9xGGaFCIzyjq5TrpAD6BQQa9XU4teqX0sZqPPfo1Z1Huml5G0xVx
OHltrwJa79bnxWguGp64jHYhi5dU1uGeQrJpZ2iqrsNosuJvs4vx2eOK6skjZhvlWo6XwU/1E5pQ
3wxNwwlUOakrXpzj+E3+fRv5K5xvVLDeSLI+ivzxt86j5uDfNOioC899ihf1s5LKB4qujuZIWemd
xh292x4nmSGHNUYMVvgCxdNaHP4UQTWAKf43KCdJdD20o3OyL0k2elW9e63DnMeFl8oqsd2Y6qWa
OnD2YbmppBBkTiMu/8J3yBu8apO6TyIBV0GqQPAX+J8H5ykDb9Atkm6pfImgWzKP9GcV9XZJMJ/J
IdlidlFm+IODvyoozIq1O+JYYexlvwZK+guxVZNbxHKwp8SBWpusXROlibEXtv9Rd3mOj122r3ov
ZNIKB5QAwQUDuFp4yvv4rcqAzqzwf7C0bel+2RA335cW0+3fkG/q2zvt5KFqt/j/B5BLbr+LoQVR
VTHly7hxDFh2Hdpp+AGoMoFMc2IpmZFRbrwVeRdkVaU/vEg0G38s/sv+ZiKuQSBoYrAhGs0YpIqv
Djgs0S/HgpNnibfDyTgkDeVxlrspcYtlIbFOwDSnRc4FNqDWnMNr7E0wIQWh6K27uxX17h0S4/jd
LuvtjUkKT4riDWWALbf0hq7iB4ZOZJQ/3czpbyi0AzNkzqDWHCQMrRaD2NF+Snij0oL/hPFTTx1S
qTiOF52ZX9UMPtUAt/iClcihG2wY7Ql/mHYZG37ccrXjwYcVf6Oby9WufUPaC2fjFrsUPknHLbpa
tBd5qnEd4OgPh3ztvJpvUQpIV26zjg3Dz3bXBbL+bggJAai8G1CqYjRM2I6wjFjmXYnjBtup5ST+
jigbgRhadDvMfkjRmGmzf5YuOLnIHplbKH0C7wjHQ0j8+17mbyCu9AA8LiC7XN755Tr6Tba7awa9
x6ju4t6Jdm5a9Yud8Y3O8z5qcv/MjHmYnYt1QDnGbUtX4id+y5vQVCeTgLrYd2wSMtp4NHMk92XB
ezSPUEO99jTFQ6VegiDfivpRcMP5SkaOVmx1NcVP98Djqcym1tQzb6JtOpIEKD1VPKT+OMQP1SS9
ViQ6uSlvyxRx4Dd1jlJgluCmg6jujA500GevwuslQXtudml7E/UdcVGdpcXrLq6k3qg/Eys+BRea
MLcGvJUE+WGnRZ4N+DnuRvX2dIen/0r0/NS+pRT9BWBqFAP+cie3ZTLwJN+YMdwBnjrlJNBS9Hma
J2P/9RnO93U0DChT1L7phQo9Nvt6kI8/fXB2EwaQl8wElnBSpFCAMlyEdomrCe4Uhybkuy3RWL+Z
K4kbJk06R+YqoBRc2JcvKEmVUkOq1jR/sGgRO1wCR69AHmwNrHMx7uND6P7ZLQxqsAf9VulzySPf
dEUjaPXt79iBvwwt14rRKVN4RK378OLv4mDWkZ4dGMjQdiItZAdGUHZBcyqXk6FXkkyHPwfyY/jd
6XNQnr27CPtCQjOF30tvamK77QlOhXj6y+HZ5WwMmTHRNA/LaiHRESEAwTBvilA2rEUxH38rylSZ
jaMMbuPgRbUI+9rF5o5eh2by3lzRfemnfn0mvDRrihqbnCsnmmLjmX3Yi5X0cYZ6+TXG0JWax9Wu
eVy8RyQs6iUK+76UW+KpUSsTX0u0NbpfNV03NfNeVVfp2t2D5yiSg/TFpjP2eEXSrazMFmJylNOC
1qYJYg9HgN4QtyZCwio03FNwK9dvHWLQm7RUSj17uXI2n5Jg3tijU1eYG31eGimK5zKJtVxWPoE7
63BrvmRjqKv3KcYspYuq1Fe5oe4uwT5eXRi3nDyhD3N/98M8rJLIUXEpVI2I2gQY4iZaBWBKOxgg
CwhzYNzA9gqSzqX3kfEfxiDa3pXT2tcRtv5RgCELSkyPMVTdl//A+GCggkn3Sm1omwcHHeM3q6mN
1kYvMl8DYitqdDSkHaT457Ib2leu2CMquBK8/8yj+MV12Wjzc7eji4Sq+t2qdGxVkqXbPj67Kqq0
wcEZ44IcHSYcjf5OCThYXsdCGg8PIFIY8+Fn63pPMW+6N7lGqL3/0jjxBpHonOBzHiktYLsvbewg
Dnl7IxC+qtwjXfuk6VAlCKnj2xDQfGzB7rPpfXdl2FVejKwjzssy00lTXQQs0wg7obIvfWTYS/z6
vodj7bM+tjp9+ZX+y/yASHhVR5JuPnzo+Bzf9waHaj3tbm5qaWZvshYvFhoqR6K2KI3TAbWPEmcc
nEsO2nqogJc18VEtZ8RMr0m8InexZd3snR8j5wUCYHXVKvwvjEOhG4g7PGxjmqgDf5Ec0kRUuuru
jBzD//0aPzIyCswy6oRRjPh1JUsQwGoGTo2UunWGyx8T9p0EmAGCsZtreCvE8vfMMCc32Fx2c+9V
fHu3oYKq5eSfKUA3viJog+JTDjnChP8GY/CsyOT2tC7uoa8S+Xc60l2/a2NXcTuCCTvPU8Kf+wd7
rHX9bfxbx+KBF585AH3Uzqr8N9Bc0K62+/POfPvebYVreVZZjZHPAn324HgNPFvEuKWfbD3RJbG8
UYsyeZVAEzVzvSOAdBY1KDUqHsdoEySR7PHb7grMQtMmNi+KyzEx25s0Y6Pi7BBowj8zIi/iDCYA
3/BXyyXUzrm560MFckLbT89DiiEblhq3Vagke0sbt5PcdXCcuPZSlu/oGmStuF6UVGaIEJ3EZquT
7cXrcBuz7y4iRIQOzAFabp97qPTVF54Q7OkKP3tz6cCXhLVKThd0q5wNUu7Ze46CC2W5N1hNDvhC
x81jjGRwLH2hjw/opTyTO0Lh779ho8/0T2tRIDPKuYeTDg13ZywPebHuvvkTChWZGuotVtq+fDud
KzoTDGNkYlACR13kjwfARB2M7LACTV6Qq7ju86Vt7SWb36nvJpk2/iv0cvc6/no0VbQvDQ1hvJ4p
Ml4QM++VcKp0IX0CBIKw2K7IC3B+Opgy1eqgYSmfnqUTAC8fDzXa9WlBn12MSIck6AEhh0azuLFw
0pTINA3L9I6eS0TD7L1TKzJgFY9GUu/HT8to7U7V+NNEEAw7VTTNoJ+FhDL+TpVHyfhUFZcF4oOC
2vQ1547rK4pIiiSrmUaRDvkLamoURvAyUTMysU4OZ7SCoCfS4lhp7CDvhoO8Ny/FvOaWsEerYKb8
hcCtLvDkhNFe3qtNr9mNhqIGGT5lnnuvfmFcv+FImxb8u7K5Xot6+HmOTqmjejwXkKNW/V16qHf2
6Rdn1/3Q0umvukiWoEQC3be5QozV/UDaQmgOTypjDnRcOAL0f9pRQiWiIeGM+sWc55czLQftW108
votOCFFlJNZhX6aFVbz7m3OO2sFFALULh1j3PzgK/X9U9BtqyD9X4I4kO2HTMxdnYVuBiaMPEj6J
1xYxlivE7TgezyQnVslLnMs5FFZaplt+KNWmcrZQyCmZUhgvEHnXSHY/hBAPRNV55hectVNh9YGN
kbwmtuWbIZiL6tGTCB1fP+nMiD1T0UsNy8qMYcPK/UXHOZb/FqN/FwD2t2H5OKq3ZVVRMlkc0JoE
2AnZ5WYlZcJ5Wvn2hdaoy921F/Q27hGKMow3vI9/jpAqTXvL50330smI9fUFr5YBSy8dBMyHHs3e
nkiE/ibHlfj2WobXhp7st7zri7pbq892D5cTxM14DimbOlyS+ebEX9NmMFsh2DeNdhtKLl0xnI41
XZitp3FQRgSpuBwupyc+w0Cse/YYjRlKRdlGwMXVIhi3lhT6VDr4oKXurcjfkzpAZEUMRAVsrLr/
6rX+jh+deqxqbn+iEgr5LVkgQ/uV/rUIViT+GMxcrSY4r9kLR3gC+21zaHPs+1MyjZ0KpGvEvkm1
0zK36zGihqB+zVGh0bwZ/OdrcFxfM+AGaRq10YTMtAib3qMAfUqjVsEThdIj3Echq2Qaf4OQ59sZ
ZJ3z1yke4u4+M1P0Jw0YZcoUbl8BeTP8LqtmEKKTGrk37EASIsV75ShfSi1lNmLCdZ0JDrnfy7is
pd/646PCMIhNBSY4oA9OGQjNrmoIx7Zx5RbWa+9Js6PQjVRanr+PH96VY14MOc4gnCtTRomJbeaj
QlBw44TNSKcvD4KZyP5Yd30kUuANKQld0dUrjZ1+m7qIvUAdzbgl+VU7fTBJRGEZOeQMyIBdkU1D
2u3rAcjMRxLTJCGDVVYLR+XIUvqvg26pbMG8KWLo01igXwYmoWlcuU+WYWVrDpWH0qJgO+4jNkDW
trHmPV8fFrxroD/G53+ogXLdm3CntW9cXkhhxVaj5di7ngj00kCFaOrUhD7oQiO9hUzJozM4oxpH
hH7PWyAptYTDvCsJIiQGz2V+fZPdZtOOgEf+Q2Z2+2sX4g7I5jihjdPKQzEAwvqf3mLrucmYI9kn
DFtYeWQ6Ym8ZMidrnb1bBGb71DObiUet5rJiOsWXk2r5q5yEJJuuc3kN0z6TQ7NNaCVdW5jnuqWP
6YMxZvVynF5+0sLGh6alC3WL4N9YUsFeCFsyieuY7ILG+ovDSQ5nNTO7Iaz/vYMwGkhhSWUI8zjC
a8Ddv1yWsFCO4/OmFPusNs2tIsBfPJT39yftDCARUonmbLhEb5CGtRIklk5/VI/9drW3dJ8yfEWi
QQXQlPKIovP7rWpxy8KdUvhon9R+ADNFP2T/V0qFXUTQzpMvn/wWbZNc9VyuQtIV5RgBQrUQNMuP
Nqy+qe8j30cLGAK3ZdXuerKJtYWyaZFLhlC6YTasdOhI3gpNSWI71E8Btq1woT7e00iVW6IUBo1O
sBWExMunrm9Ub5Wj9j0wI3u1F+g8nsCfbBRSjZ0mjWilPcgbimHBJ9RB6+R6Eda+gZaP9j+OYijg
KleX6P2pOwt+hZvMY9NeQOP9RFhmdbdEe82Z8YnstJyfNUg8PbfOrA7YwmRdDDrQOCbEDAzHqVom
BDBIh6xdIK+3DCECuduvfhJkXz9OGme3aQcfzXAxnE27/QNLn8S8V3tlLbuCsySvAav6NE1m4P6H
GcTshU2rO5vGtfF3JFlTXluAIjcc0uI3TUL7gwMZO3Mg6fZGw3ZooOfr91TLWeU7or07rXdqXXYy
ykeSP9N0EJnYOjrBWRGoNXHPa0xrLTpEraAFrVro7f7KE7OziJBdvEP5khELePCggESyZ110+n0b
y/CJIppopyPkpu6WoS3B4k/flqoTnmI3HD5RqzOaS9tFMKswndwCB0GmDuKBE7ptrYEKx+qYgrIw
Dg0v01eJ5hO3PpFbiFpI/fqqoAv3IfgRoSqFemzpwXuyYuMKWjHpRNMAtLaxDzWxFI9BrOfDb//k
2Kz/oNo3b5XwSCpoYMzZHUiOzwDFMEqCGKBFWD9ige7LNldjWBvpMAMFZwD5HtJClqS4sXPBMmV8
7/YfzViGmHB2uRll5PyH2RgVtuiGOQP87TVCC+MLF9J6QsZQbC7fx/TwM7HgIdGnK4JV9OzNJWl9
1F9Ab/sAfcCbLBw+CTE/x2Ad3pKkOIXHYGS6QTPFEUGdZFGP14YlCqE+RYiz1y6i1XLe+acaaM3M
GSSdppl4Iwh4TUL1zhBn+4v8H4wNIQ8WQEO7LAfPkZw2q3q2c9czBi266Y6aqjEXMbq0FiLZVGKP
+aejIBhWqwdS13SdalfoL8NrK3UCwsLiGRP/+1M+f9Od9e1oBK06qViXBR/WkVu0n0J5l9devKvk
TNUfyI+X5OtUh7v0SZOF3HPuOwYgjL04wAYDpDFRkXnaIcWY0sKx8sdEPuwE0nokxCMTbQkv9Apk
SxvouCL3pkCMYE5iyx4DWwOXkNNfBH1x3aSdht1NpMfIeGJCFjZbHsCrA5iW488M0VnsMcev7zwh
ZbXcFXTO3xRUzxcVpDFaxlQy3hzrp4uij9EdErgb/j0Nf3aV3qNzLKbFVWA735A1ZiKJG1ByzNO7
45axDJwB4bQRlJh+GAonbzXaC9+D3lFyGd2pREGGMvjZBucf3fSKrEGknI6GKDK1T2OEtbXTCeHC
rabl8G0s0G7jy18DC06guFR5TctYw73DhS+hUjm5Iqm9PsYeaFnK1rpKbS6EGuaADrTj1VCCilQe
2Ko6PNHlmM2r5mLHcjiN+fCOp1rkVRFDu6djWHUOCUJdtWgoJXozbaf1QNUNaZozDn9zPmMiXEwK
wOFntlmTfYuu0JbwOolKPWkC8yXoHzSsOkhmR1hbEWVfGKs68OZccN2x3bGD9IIZ8ptJSpNWtmuN
0KwPHryaWUtWmDZp1gcSUIkOzG9mQ9Ro4Z2Cp9vWsk5O7W26XTn64FuD++IYegKhCXrN4lBUpqw1
abMNSpQQ2CD1/E1Pougul6wmGZeWjAVTYF5h/afyoVQJABcthlOmuQymQ8RJ+/a5EZOu48wLZ724
EUI8KwCvi71KqxaabfgwWuZbgDCE3GacGfvFU20XLMYVQdCZV9CR0uk7YCH01k78+vt2Lak3LEGy
qbKc+h0iwhxghzQyGf2hPWYQz3aPS52CfvRw9xyUqt7f63digSELaGapDyGw4j3NX8LA+01QPFoa
V0TwW4pn0wIttCDOIjwin/MstMLM+ll7gnlf32TuBV82PI5GmtAtBu4ix3zmqQdpToNuMFZdIVRZ
VXaq6mhux8pbdNcscyl0Ep4BLUDxbglOOC/l0hfE7UJgdQws8FToj4dkQFwt0XJ91GQ8hkW1BeQW
3OxV9rgXo/U2gyG4XLLGZaLCUiPiqyeGrJwHVYxvdEwmukUbSO+nwcLCu6cMA8NvTFQ7SxCv9dxx
it6M9l+I1+ES9hlj1A2dLPmCfQV7CmmJ5nYofjgOOH3I7FGzu5s3IW8iuUF0irhydeQB9wJnUkxM
wOYkeaGNEq6Mt0U5SGXBiOsoJU/ftkRZmhVrQ0fXZtT/VxIZDVVTAXxnkD78BXui/0oRAoXtkEgY
M4vwMX0uiEw2BnANnl3OR3CQAz+qzvDQQCsBWBxWFcHYN14jCp46MZGpGTTRbeQA2IHMcOczJ/hU
VKJbaDj6DsFLCcvHXjtC8BpMZBTRvH+DzcxsUamF2wHfrzCDTP28si/ZFENpOI7wQRrrNDWWAjc7
V+LXQ4pUwh6g2pIaUG7DoaS6H9FUtBV1smAtpds7Ek0birpfToM0eVqa1QmXEpi1zt8cdyygVhjs
QZHJ7r22knB/hyOnk58gXb6jYeohD3fIizyGiwm16K+cEVtLqg8iu1ipDeaUC3vc1kd0JcYEvvTd
H9LdTdQlwxaDHU8TW3xN02z7pxajzOaOfav9Suz8RJ+Y92ro92j6b1qAKR1j6okUDSUUeQm7Avj/
Tdd8xJYihtylGZWeIA0Cc8lZPqk5i7CIKnHw5kv4N7NZywvkeHXUyepxp4i7Drr0D+ST/nMMGDvQ
IWSJzxNLbhwFp/RO0hGds9mz1+TJmqGg0FOi7IQCdziEPH8IGPM7aSz3mVSV0tuuyFEklEYHsHLL
TclpG/W+jLaHDaxohQfTIL5rsHc5O/5ELNbtQkjd1wKW5p+f4Osjwb5cVlqn6RKWBgj91tmAAeZJ
4mmWLB4CZk/ymhlHxuks26BiLBEJhvlJNaRmDP/VvofYkNauqTHkFMfJPpZHU64ge0A8nBoJemZG
SFAb/ZzFa5XvWdxWG4B1MmHoaHMAGW1VfDWb7fM4wqxaukNEmQV29G5+Y5SAnh3St6EKYYjJbimH
Pvtb22KAR8ePIW3EZK4StyynBiUFm7uq4BbYJ/wZv3jy3UCHjhH9l2kzqPL3BWaiZ/8TA+f7XBNM
z5tkZiOt6YpA1PwpoNGs/AWXDQWVsDiexTfZK0iDFuokmjQ6LjOS+lvFu2M+XhPUxzlsY/yBNW0m
UeSK7BgxrsLmVKTa8U/Zo7E29VgZR7W+pF9ZpTCk7YgQyphDilDlJmPNDS6jCqjjNGXsOqrqT4Ed
1CS9VqurRUInaYx2AUaP84cJIz6FMJp299a3rkUwzYxeqZgILXxGmkZmMDntJbliq4Dww5DWP6vf
X+Tmmj0EKSSUSRY7nKeJopRYT/0sPY/oAYApj7KHMnRnmQ9SUdjeknbLXfVNQ4Gf4IAMdYZwdsuA
wjaP+PqoVBI1OmqBr4jGxiukVHTL8mpuyyxS6Dcw25+IVhFvkYxePYgFvfMX355gB4jW/JIfBMW5
kDDJYTpBsZJP/M5BfyFT+75KF9UmvowHF4c2V+rOIBOWH4Afz7kqtkim/2pV3brXUmFR9QdJbGIW
FidT5xpCYPvKTPwtYMh5FGbfLgfukLyYJ4MY4zSnyoHXygwQufjPF2nmypeqBWNkvMIXYiUpjb5D
u5JZB1eyUAq0910+KhiokO2O8Ifj0BVHFzlMf+HtrWWOeG7OxDoNwgDFzsSqMAFH39buY3yyHFZl
8UaxD7NMF7ay7jNtEh0kXjIQSvCJIfFcPt1iT9/5etl2w8txlnb8gJqe/G6CblxAgztwUf0310s3
5MN99qFQ4l7z1JsD8qU161KIWoo0Ez8X5ugXpRcRiQUd0trI7UR8KLGSLXgjkTXMF5Lwc9Si/dc4
k0Mc3CD5b2dYTERb2jggjjZ7QCelwbwGVYFnnkGdQ1vlWcNDwsCIOZ0vBmcBB7bDC1OB17Tb+k6E
iWr5LBecEtBn5S+G5AZlUL3ewucv9hz2+kSzLA0O9FEoR+fmmDKZPUcoBMqJJadzY2/RoKHL/LpN
LCkxKewF58sYFb930QOOH6MYCBKL4qxsxIHEEfEHVncz2bG9zNaGOGZTxLIFwITnPOubqvWXMmO9
iTb8YvtH35Me5nBHJ+4m6KfwHZYNKI59vF501AE2XqA3mo6lVvkxxJcKxD6USHU2zc27xPs91FQI
Q6/hgOTw1HPus2DaEQ1xkHe/fbokg2oouu1NpYyF/AZk1JYw6suP+e4WTZj7ynNkjWwLUdJWQwwe
a3fMm9NgXsoXa8Lxd4+IZWGWmgk0YnmMI+gzBa34GJT7sjyd0zSDZJ0kZKk3RLZIzZty03eT8tTi
416l5izBiMbu+dEzMdE2RVNr+GhQJTz2T+eLW+qzBncjUFESxyE1MHTeIU4LS9oCZcRYSyRxVQSo
6LYtb7ybhG/4rw5NRfamsEOzgkE4fYrK8JjUKjH0KT58+hl7IEfy88qUCHGGUDZcT94oAprExfhu
aAziFcW7cdCY3Z3m5+2YbzXw20WTTQGrgfGh+4chas05hLBkvuFoxV9lh2n87Rz+s2mg9CX2etGI
iwGaO9ufzLrZaim3cYaWFCJz6oGRNcTB8xxOFuXeM5cHDTZVQ6CjNtbQNTtcYxTzLX+RuOMBupZN
mTWitYvLCV+tlrPUIzdS+cwrq5rscBWvB02aWK/CoqVAO3te8Fz52dwJEPuW4paNCkFSpu9HlqJN
fh/jrBQD50DwN+AbQujdckUa9+gF3+61Cjh1PWddVEwQidqmVYp1RRyHPx2g4HYPfGxW2V5KRPLF
xAq1Pb17wcahGAFQZhJq6WulX8mt8l7JAxsgyPd1hxvSKMJ9kRzQkkDzPbNfXpjuQCWExcvfHLH1
CK7shcMv8dmdXnLUCEURb46NXzu9UkCnQCleZOk139hJTYm+e4zBb/2Ws1/2oqMcxS5/iQNGJkLn
wTy1KPmdFdRT6EGYxBn8VzVQB8jB/tU3mE8T/0xEqeXySptOsAxorWayiah7s/wRU6mAA/I3/ZQG
6FGVUqNcF5RkohTcifnX8bJOlhEMJWfcQ9R9Orxz7k9gt+Ivpc03dKVzmG34V9t87yX9q/sau+XJ
JmH3XUDrOnl2bwknncm5iN1pQOHPJEH9kzprtpCgEqHKFnTRg5jTV0a/9/7IZVVLI9lqHybLFlme
faEVYztU8DFViOLf0AIprujxqV67oZKLNk8B5YXEf/HJfkY3d57bDllXN9L3zNi8MlQhfRA2BR2Q
KqngTRWwh0cUBrnCDjEIIqyVkAwuHpbf+z+XOHJJ4OTpve5bk9sNbMladr7WvmlYdx8iF2w/cV0b
+f1RIrDogOYPzvHuWblmCyUKzlb6JpFoQSnqYYYuRsTsAcHrQ3C3+s/ZpqEJHSnqvbdRTBUpWiST
6LRaqGAoxa/tGWFG3HCQ55LfA8Z0FNPxTl3B986Rf5jyFjEZ584ONCOxoepe/4ytLkudXJAQNIN/
HLpatlBgot9gMunw1DWl3ATXiY/Lzz1nyzFB+L0tQZ1UGJmfbVpOQQCYT0ZGSVhHfIFd4vh0V2bM
k9MVfsxY0YoFIxYJww1K0KCZCyEneActlMaUfFtq9X2A50IvPpAb+FZlNO7VFWF+atK5/gCWeBrK
H1Gbl8qW1vBnD1b/nxnVf3xnQL4rUjc7NdyQ9EZHl8nEW+tq/Y7YIkqROL0323g6s399ZgI934SL
LXQpHgo83bSXjJPDaO48xQ4PGFJnxUDDevREoF9eQgeedGF6VbF6w55yUfgr2NBYAcpzc7giFsES
siwfR/Vq1MZKpxdojm6suKxakZd/M5s9d9tGW+LQtKHCtpMgMiQoZqy3KgczXr3+zoAb61yF2Urr
Ogaqmh1VTgxCLD5jJnLQF66itcs1iN6xnx8GgXSBmjZSP5eGr2s6z215TEuuq06Xk97V0l7PWh6h
2tJn49S6qbkhuf2VTxkqOxlb82AnpJ5VLbo87ag4VwJ9o9f09aUZCmlXoZYbg31spOVxBEPL/5DN
ki52OCq9a0PY+Y2OVJIoPrEhwvzxFXZxSm776NVvOXDxhnt7DQcD4oEK0Nbtbiz+vuvOzph0xbmG
MZS6O7oMJtP1v1P0UDfbT5xH5nSJI9nUvpcPl6rcwysgbc/w4TISRjh3MYrlSaQvZdVryohe1Svu
ZKsr5rgqHVXoIP5t7ZY/gf9/QDKfLap/8/AL7UANU0aHwYyQmCUHZukKZmmERrVTRX/4QiNlFDoo
aq2Wh4BIHBVtLC9Ng3fT2CIkYbpNmceAS16vYDj6/dZ0XUTx86c+sVaZlCm9NLqtso0Bz4mWd0SC
MM2HgAHgoaEeUCaWTCp9ktsvVR+8B8EqjfxdTUGx4Iwb4ksaO1G0TvjZnshkYEp//6ALTuBzAbFm
823MPnA4q2BWy1NExaCQkBdJ0msZsf6wicSuI57DBVlxqUF+ElNTHYQb3np0s+mQArMaScbAXHAP
EKnMks5VnGFJ+0v0whWI+3vsl6eYIlOO5lEYhhO1mCxu7y/w3afQ54cgYRzv/+YcvOwLhq9DfUVs
QyZ646aCYVODabSUH6EEnU/QCYi9kRZcoxDx8T3PK+gxPax5InPFa/AN6BMrGw89Nb18fPX0jDK0
gv91cRRdaBowfB7YLiQHytqLCgwd6HIa+iS4NhBh+KDvZjzVQ/BqKcaQ0FJ47RsuaqP79w7LCceW
QiAX7JpaGG/nCCC2STCOJa7FN7Qu1EGRtZ7xnRjAI6hrzvpsKdN4DOsWF6u/As/MOh4C7cy1PDk4
s3HWk7TeGsQPwG52UDYklue2xveEk6xgHRFOe3eGP2SGxJ8SCTI1XJVNB0kvK4GeIYFUePlHev33
TY3/Q2L9YVtE8LuJSBR7qdBROXz5Kb7td03pOW/GajkQqSVzFTyaejd2QN7Twii64Da/bYlGDX4x
2oO3jr4BtFAp0+JwJCQ8mGUdCro0Vnz6q/jw02Bt266LkdvSNPkh0Xl1t6fQRJ5cEVzhei3Kdo3Z
ct7a2X5xlcKKXyVsIChmNREsKFOo3mXiGf8lEesvNSUolQV4/0H4wefLBia8BALu5KphoubIShZ2
CtGauTZ4lxfDffURhHwGFk69hV4eCwRnf9CXQecDAfhf2xz4S93cYcc6m50fGxeyQXfe1VW1TUJX
8Sneha1VIpTyM9sG4Oek8+m4cLQyNiPU4X1DAszABsHu0UomEVEspEDtxo+Pn1IxgkLvdqr7vg0g
Ab+fZRqgMKKDTLv89OmTqA1NeV4PD2+i+oSpuEuhwC1o92d8knt7WCl6+RtqmnuWZr/vG7F0LAH/
R6goBgFMHr/aDnI4uTU5Hkv5XNsWqlMdORjgYr0UGtKq6ODsrR98wxMmG4N66fl7Eklk5vmP759L
TxrCzMCRiW4Hcb6dg0BjO9L+8yD51k88BBwsTvDgFCg7k5xhxp03T1dqvOBF3w1q2IyNQUedwJw+
uJ9c7rC83/wqXWtcisLJUt7+cjd42DDKumOAWg/34KdxP0MtqcfOxmt1ij4UCKQu8X3T/wHPyllw
F7Kqhzpy1k6WjH9fDbeV9rkG2JRq2dMSYLqN01BtNGf1mtZd8aa1UKSM62Uj4amnoIZep9GptNac
x76nto7roq9qY0B8e+DcAoI9UqEmwCC4x/rohY3daJnN6wc2UXCa24yA6b3rTTqXz+Jyh7eMiaUD
csbmpBEVfZytgPBTSmxStmCoiNaixEv49mHtJLy7ex7FQdyy9hqDGjA9wqJf1yRP5S2yNIXqR0Nl
oC2h/KO6sDn97LxqAREKhAvV9EK4pxSvcKUOJ8Hy/KLoifaY2bVl/mo5BZwGhSSVIdRE0JQfLBEP
BGncauY3SGBb80zq1cFvYHbT+2kqXxyJUTAA+LFDuLCKrGtbU2IUkLayUPeJudR1LxgDDInnwuAA
swk47DIwem1C8plubCtchePvumhR99dwwZ58cmjQD0vgwEkuTc6F5yJXg7c3tmWMcLzt7AulxLph
8SJ5CKnryOPMQCgOf4de63TtH/gXNRFvQCUMWq+n2t+IOjNovXdlP+7BXPw+jUAB/ZYRwIOTYZjH
OIJbXXN59oOfxpJa8A7bUkRKXOoB9emYq8BrM+Ck11duVUDrGxpiNu3u3zCajO3YhNvqoIoOCyX9
CgjvxyXSSOQa4OE3bYmO2+XlZ0xYomLi8rh0At5cLwJPFYC+UO8Wq3DorIAvIPcffZmvhmki7y0e
bBoB1xIesdELD3oH20IBkmrqZw9jc6WsQLIH2b2WiHlbxJvLULhglwjOEiX1THVRZ+eCktcNrmkU
KdewZboW9FPXMiZoYVpQ3rsD4x25FWusK/wfV2neG8/4G5d7P0fQzKYKlc3jwVg6qtw0Vl6SbkO3
N4WclkXmVECVZwQxefOhhl7ZWXz/cpmGgRAT+zBB7ZyMRrcq1+YP99rIlFofcH+8JRTfQweqI2Jf
daKl7e3j2gK8dLFfytkfnzJyMjKXhs9sxdeCxrv6hq+8V7/jK8fb7A6C6kls0wh10Bsb6Dndu4aY
4BEMuDHI2VIOf5nhgVOqZS/wDDyHjUfn57mhdR0/GLKWYtJsva87/l3GkNlcckB5CzPDkxMwfZiz
SauGO2cyolKsF19Id9mMFZaU3DSBwuHi8wg8mSVUKb4jYgaoRVVruLzkwPCx8G3tiFSCeNNb8pO2
voNvFf9Rl50f13zLd+W3XwPDBLhyK3Mwt/SRYTSYbwLAxTDVbk1hcjU+YXa6j5vBOIVOZ1aC9Z67
69DBQY0iSWR7nWhEWu7RI2Xcu4q5qRtzFL+Ve7t958v+hrE6+qpwCjZzL5nUzpRl+M/IKW25i1el
0/1iFLq4pnuR0TNPKwuXwSlKaU9kQo4nMvN/m2kL4lbmie9QZXcUVb1f6P9uysqSXo63pYLv9OiK
1ntpD8liWMGfyzXY4S1aYvvxpgepK5VJbMMgjdTXY2LIxY/Td4eqp9WllpCijmmJrIBThtXZLQRG
ZREMkXZQk8qGXFQvPlJfHc3yjwxKkOtz5fDq1K/V6k6RnGx+n4+LJluH1Lqp5VxuQblHmXDhj6Dx
9pkO/0aLSAzBjwBlBM0VVecqIRRLmOPQJzTMH0iLKuissEFAofWLcz5iHsbo/Cm2phNG8GtRbjWm
b7dL8lZ/+FNS8tXJm9osI7M2s4+9UmqqE+pJkxx9Ks8BCz1DZqBV/b/VYUhYXOr327oiBUqYXNp9
5/rAfk+zZtd9wE/jceHmzxExbbX1Gzb+n8sh1/Zp6zIevNZ+NLYsMqrnDYRXWOhE2t0iQQbPBJiw
JezbnrSp2FOpgSd0y6eM/XNOATQ31z7c1jsZghDz4+xY5B8UGxyQjHTj6bo8I7f+t6lnOMkRODng
V5KnWrmoJ5G86+zwjTF/0ZM5+djSmNj4jrTgNe0l9bmUXR1LbwESPScQlsFc/cj5xPXCVVrFXM2d
+Fsyn6Jhih6qii1N5qx4Vn1RIEp81DlJT2hg6xjjQdy+HT4yeLOMWd/qQR7YIupNLKZMwfC43GdP
6ozAGP4luVTtx6AXXcLwN5EbzHdlQqlwPA1tvtoJHbkGyX7/SVZQjnPnRNdZuo5z8IU7YivdjAJJ
+ilA68uuPQMcTuNXVRPvg6jflg+sUoZ21Dk/tj2BiLbMPon0LqJDB0SX+T0BKTMeD4gyt6m0RHbm
MZ/bDgoRyQwOIQOMlXBwsZbWcWl4l97HrXbnA3KxYeOtkzJ7hMJNUq9DAkxU9A2p0XqLU8apKgkv
9WwNhA3UQrQIdmLrsXvvVlumttyCHdj+gMxMpG7BNb24Y1nsyMnRhRCyZByEA6ii1JPIc/GUCLVj
VKkE+oSomOYpd0xbYLqJmkvLkjBXMnRuToynfSOkxzFTu2aWbLSCBbcyoj3Kz9lfz1jVQgOzMJCo
45ch7SnN/rFa7xsGsjqWhINcqjeLHwKQgHyMU0fM9Nq1Xb4ZxJeI2F/SMqf+IWQ7nh4ZpXeFCE6F
M44ISR6eGaCpSV1Nx360Ed/HowTBKOZyIx8OSY1OuTEykagUT6rFUtbrWv7RmYmmG3w+OdG5poI0
K5e/I4Q6EMKV5QmSAac7evBpjKaX+fD+zT/ED9oY5dar5Y1cVVu3w6HBoPH3rarLFZ1jF05Z918k
qkU9L92uZ724msaR6NjeBaTOGi5cssiehwbXT2sW0hR1JSENydIlpJR7AEatzqU/pFrcwN1aJMQb
vNoJkWcTQGSe008L7uneTYfHgWG5CTIZo7HYH62d5FAcHjsyf1IJbPe/W3XkxZGF85qVVR9+DKMh
KohvL0MjoPqcjvKcheFbkjpdYuaLlpqx1Dg843ZvjK18bvZq4n9JnxQ9jpGh+FvXDOgT/Fam/9yr
uNs6cs9DfwheOhYe6gvqyW2D2urv6+llMsILHykF3wmlKgzYDFYhLhn6ck+uR1yFZyQRe4tKxdOM
YoISvOXRhKczg8096m8hrPgpqLukbNTPTdOCQ/4suQmtGTD9fRDiQm+iYSDFrZ5FWkV3OGHg82hH
ELzv7HUtqIX/v/TabkXib2djaEInTffEwatSn/qpLdxD3E20U8Xittbxz8NZfowYK1HzxepN9Wb/
AwEymrcLjcGq5QZqOHWyUmBV0If5ksiRqfeoSrWDGCsFW371xGwI+dg/4e79TEeDkh4eL3f1z3Aw
ug91bJkUZ5jJfV3VtZCVA3giT1OldFR1U7tbzeTajXLzgcSijF/+hLqUbimzIfF531n4rYNhfPCp
6wp9FM0KqFHhLVT3U8yBlIc+ZTq2gA5OpBUyWC/ecJecIHeFMznCkn0elE4IqZoH+fw73+wYOHsn
/iiXReC49JRTFQCgHmDgKzrAbrMv2cuSblHyMLibjJOik3L811/S9whger7PPKcAAoNt3GSvoaGU
qFJh/u5W6WqstntRSTZj9PKBI9I1EeeNabA5lMsrw1HubXlrrZVKXpzNkLR8iaqkb5kl4x5xptnZ
NQWo9nH4P2yVqGCOBOcOhZhMUPGdBy/WI3PIH0qUEbcF64j/xcFbw6acigG9YDQfCVSEzHc+FAYA
3mqfkuCL23IAnMk2MEOxSRdX1T0R74/IgSoQgYCSJ6TCazfNHO402IY07YhF3dYg1YvrQPJIoNaL
hObx6VozcofgRXPV2kRVI4Qv2xdLTiHsEAPlf1FSKe3auSwv9RD1HsRIIra7N2uVFXTFPkPEBjqa
1s4Hqhm2jQuxrLNrIifvwO6G+22MsbBjRxnpGW1vgFjeXiEknp5wIbyjNokavprmRfU/bLMU86KU
gJt8/O3xcXtFWl8cM4u0EGaY+iqotceT2X7a1faXGmt5BkaeDKmgOts4Cx1BhJ3QHIhBP4XV8r06
jMpXzu1IqHkgW4F5wA+d378Jmu4ebvth802DBf8y0T7dWfTn925cJni0xOM7IU94JQohPwlNuCJb
OK5vJcTZrnX5lSXomZIQSnX7nqHKW8tO4EJQJRAG6dXrU9KsykrAcIHtqFJHberfinlKpq6KM6XV
pwmblKD41aiIYFBoWIkef5kZL9uz8Gwb87nNH1/eXjER9Cg93Bpk4NNFyzzsRbD59Bzb0Iaod4HA
sfDVMcMv0Z3s8rL6Dmv4rc8BzQb3BQwjc+hDZ93CWwnEwCRvGE5U42kkYztIQlJjMGpA3Xzx6lxP
Wx3gGhq+4DsuvCc6Mg3E83LyJVcqJm1MypVk4vxOslRwgcruztK+mO7Gz6nYsVFbNV4tobNVYfDT
yDzgIa/cgCsdK5o7AVD1zRClwV+rZcploCOG/amKvFRtmXE1p7vKAD3+1vIPPO/lE1KP2/39c0DY
IRufDgYyI/MuKFzJysgg71/rdLfcXt0jGLixlYAgpdUeBq+ZKr/4C73llAdC7Awd/2VZrH32asQN
KLgToR5mu96NTfAKo5K1BtPeiTf7SnFBCjqtRQ+jfVkSFvl/1KzteARx9Wz23vOXHLM6+fZuNMzK
u+jp9jo5Wf+N9TlcWkqKgp+VO+GRPZMeiUydc80V2P72SUqeJpVcHpSnD6nKDw4tKwihmVc72cKt
G/MYlRxM1xNKZhk8RdvZ5lVCU64CdBlP6/jQebwQ7zh2y0ibT0cYan+DIw/6yFYFUP17zFG46mVB
s3yF4B0b5lbaKnM2M8xG4ZIb95IGJSeCE7ieZkZo2VHdmzHG8Q3dQKzp4NlNi0DG/0yfpbBTZBAY
mTZOu7YsiltSNlW+jSY5lDqB+JXPF10oJAgLGcAF18XGwRXottfoVkPbyy0jAx4goM1nums4RDha
udOD9zQIiYmE+ELAPSRTagyHeRYcv9ZAx9RFR5v7WjmxMa3RHu6FTxi6oD2Vzmdjo/zrgGa/ntf5
vlUB6harV9Vsdm2DD7eH3cS+4Sed7ILBzpD6+1OQcZkTwPHvOzwd3Rq1426njLrdiiCc8J9MVdx7
3ClHu5SrCQInniiM78wwKLEmCbZlI05x78D0DmIUAbSCfbciI+etVhSORxUEsVeJ1qaIg/vL6dZ4
T/0wXr0hlsiJNJNcolIwWm66ZvwSOVI8AS1Il+Z5wfqk9r8IkrvaD+Cxh7WmeX409pHPPM2dJVbW
f5jB1Pcbim49xuS8dK6yoNh7aWshetlqD6OiBRrDkxRf+K/64lYRXCNsROv/9j0r/+tesIl88szZ
LbWqikJO04dgOs5U8sNiPy91mR0rhkxvODZKTXFw9r+5XogzXkFtDmndTTOHsf/ZdKZiGk4HlHDY
GkDbAdBhrvbHvEB6wELGG9fJojwfcpxsfYjV/Z2vD2TOXfsq4bMQLWdUiuM/RVwXjZOQ4BjnS2eZ
LVJL7M7fZivQDiYX/rVD7FHZDky7ppQUG2wgnpZNtlf6iq4C7RX1jNCP47Ff87TRN3JXh4ryQKDD
JCGRISxuUPcF1nnlkBXOaYgk+TrWNPsToBzosMwb8/rMGZK6pO/q1P0L/0eOxr3MUFd8Qe1iLyJj
UbMhOJ9TrUl0rgdgl+zndgma0iGzBogUlWP49aY7J+Gs7AkHDEYjD0yOHLzXrkZi8pxnpGQcfV28
z3UO+VPRXRRTI0QB6HlYIPqG7828C78L3nrFMFvWLb0pKQ0VgT2gCbeAhGWaNzpV8kMrMC60+aGQ
joNA4pu2TI0aYlj/uWYPjIS8uifQxqnntzPpwe06tudHNEXgn+12xCbU7Zi1RbDMjNTiGZz2ssug
yzH7wrrMrh6Dc7HKhKSxNjPRdiPQoRsSXc+mklwQ9aDQoIfYuyoYjSiv/GZr8IdFaKV4xUw1a9gV
7gJxHDyjVuLWesvAg7EZQHuCt+6AmonN8sikXZ2522Qxe4Na7a/SRa+ep1gEirdoDoUCtQ9C6Tx1
4Cdl/q88PCUArOOAplXSLyLLaJ8Xw8OMH46E3utrp9ztKn4ekVgXPn7sbLRWJyE8CJfeSz4p/hD2
mB3N2yg4O/DNrJwAYsYkWyBxvp54x8TQJU6A7HjFd0fTEQrzATEV/6Bomx6FqiOL8yxWygd7Juzb
Uz4PAW7xFTOuOQwsrR6sMzeRAHGhpwl1iipAT556EJRUnm7KV+DEk1P/3Kfov/e2P/r/Qh6IJqQM
uVmeS2xBpRJTCdbG45mDNDBqyupzsbrzgH8CwlMBn+qxlQL32+xAkzvSxyKYFAfohZRTURUguvWO
ZX1sHCzniRU6fTUhmhRwvifd1zGlxM91ER19lm6ojS+CaUQfiy6yLgob13WaRo0R+WQbiE3rSJB5
L2O9tTcOvZ/N3rDWE6izE6CE3BD1QwuWQe42YMXgxMppN7mk/ifSv7MkReaB3pvzJKbYtqJVb3RJ
QBI+mfvHChI7hpEQU03OvbcDg8S7exUpQpuq7ds0p1OZkfXkDF4xZ/aBrgOye10wJ/mhJjOAY15b
g/fyK7oZTAq9xRIgvQ5DQL9nRQ25bZkHIHq2TrJYGgtnTYxXnPoaxhy8/xrzoXf0zPrC12587vmV
PzCnhSom1vFyIPSF5qF6/G+29LvDXUoz9PzeMC/V2Mbfa42CHSJ2UohyhYP/k7GhwBab1WyrYZ6H
Xnf6WscFukI5FiA33r0maa/KdpkxrQQqmcjgY0wkqKAx9LJNP0M7/n912rfs7/uFT6Ky7gI+SqKW
s4mc4kGmUII7kJSZ+nVqBK2v7y69uO1VNBLESSEjaQ50Tpg2VGLkqNyPh11IWlIMWybsGOTy0Anx
UL20tbN8wtlMItTtI+q3y67oghbeCwJGBQJ3H3cjIRJ3gUh7etMV+EiwwuY0srp3l6wcFZ45zo69
1hER0GeuiJGBaR9Nl4ewqRBLzT+yy30/aMX5Jhqd0XyKmxVhg2XBDq4M0zI2ub7XX99qPeNrAJQ4
29amIL0PjB0Qz1hGANsM5kSLVC19uwt0/F5/pkIeszLlmW8QvuHecbcAlJUu77Aa5HP5XJr0d7NF
GEMLHYjfJhbH6xe9HKG+hw/6QIjy94Pcp6VBeIvAlbDJRzrG/RSXzbBIlGqkgjSeEJNVvOUSDChk
/5C+btMuGcaxgCl7RppabGrQmPQEYdwgda9piUIS6AZt2ej2WzjRd4I9TN9BRuYG5myCob21WzNQ
Hu91VD8WSWEX7aFw5r+NT5VH5MfyhRkTEd0GkjBCcCwFHWyLClPFK87KmJNfDYQ8Cm4UewQ+5YmG
GeH7dFqhAQ/ltXYjYaqqORBJtzaoT7Pl4LmRqGuJUdQbHMoWPt2tCAlRb+0MjrS5OkGgUh103gEJ
uas26PATHGjrlooRaLn9BDvQR8yIppvhOrRabC6hFk/rYNVRpTiB4xMipmaEW2gqNMbjmC81yzbn
xonAuERIQM8iaiWiDT/bXu6ovHiSjC1P9/x0EQFuxQiH1CU9IoFJ87PkhHnC+Z/ttnafZq33wFUt
yAJSqrInGyEf4LlgJ5MsStayShOW4oearbFsTCbOV+To0+12YSrfOpDB0UkBVTLZ+TljKd2q8gvI
ytjS68oMgbun3HZwqoGFk+t60NQc/ntORTOJfK6XGtuNnb+7kgqoUjxt4Fzq3YuLCv56/cF2o1l1
XDbWskJuKEd0BxTCVlCAKVD1rkShc4hbGekzXEl+mdi0uoPdCOQMpGV+Xax4SFMn43g3ftuUa4jd
tSFBJZHfdd4TA96kdnpMacNK6czLYLNOQXFFJhbcvzpxhG2Ju5WqsOw7ayvtskmYtf2/6BwnYz39
jx8G5Rspt3dtzCroOxkRSBajEKZvqy0hqR1Za7tWobnBJyW7NydxR3qFLFEXnJD+MD8gQlJW6wX9
1aJ33cjHn2CpO8P1ocAboLlhmZiltE+DPpVfd8TO0Bt0qHRu/NdpsT94xNMKmcoFjWZbgGZI4WK3
NB5YS/cbelIHkQKrxnAuQ7Ab44njRDF5+hmsteTvAXg39r0vxvzqk2n9F6RcjNUTSlgITRjoZf0P
zGCU4goo8v0bslXviik2Tt8li7dluNgRhW4z06a5ekQGKrNMsa6tIxrOnewRY5R2AdtEdvVqdool
mgidQKt/FU61akJq3VQL6m1Qe9+nbit0SeLW423MkAj3toEd+o4hj2lw0rvSZo8qclksGeKFil/v
P5Mvb0t1moKWoMo0lT1jX8uBmvB77uTEt6wqnTEqumWKoM2Sv2BcoF6EbdX2gAvumn8gda6D1H/7
RZP1jzHyVQQvrKFWPk7ljQvUYxbHenJjUE1LxAksxR/G2u2K6D740zcV1mnnLmEQbyHrlVAVVEb+
Loe+Z0XSrYoVYQ8+TeFfTQEYbhbr+EyA34vdaHWogJGP9ezyYCWg12m9g0InCPNSlCVZabJ3gRHm
YwaSMEBQYuR6QKAIgwO0CZQIWAV7FMBwQSXBMbLCBwivWvlSDdZYWhyJsolAzu+KMO+TAdZz+lBy
szJ46iSeil3GJ020nSbrsLIaNiysncKap/N4ksT2uSDxIDV7yl7/GvkHkk4ZeJy3PvCM9mjRrtSw
RulaluBCH+FBMP34H2h/IYAG0C2TFPXU4QlHRYJmS01T7hOufzsjAsn3cQsgKFUMP8hx9xcVTVpF
fF23SGcPWAmPRBCLfoTEa6tj0x6kUSqUh3RL44gU7c5hB6zOxk8jZNJbKLh661lUnHW0+5jBRQwA
tWxYZxVI8cVFboSuwlanIyW1n9Cy/X1xwLIS2yg4bGa60wYTadcibzXx36kfkVwo0XJ037+VbtGs
E1iOp6PIoHhZufX4wBTxmJa9sg37Q+htt99oIfZOOStRG9snhZZPSXM/6PiI6fmunrsDtinXgnSu
Qa8a1UHm7WeNwIjV1NfGuAT9ylFnJO3Pkd1VLWNqHB9x2+AQf/MWBtW+APMKPSsK9lsle5Sh4sEw
6HCn/4I9G5b6tHai9L/Prg57vfoEn/BsFt5KMr7/4I5lRWw1Suhf/Tu3SllASVUuPj5GxN2EJmpa
C9BxamHjdOsAAMdkOPfHRVI/c3qsDs3E1BgO7a9nqit1Rq+KIOO6KmJ3cmC9y1PVH98LqjtXQh0v
DnngX7iQn/JB4kHiDgGop1sfhl+xoYgkfz72lafzr+vPr4tBkylFOsakzisQ9tpT3N89PhHj3wKv
XfZS7Gajp5HLOPMiiAZ7dQNrWMguusRgw52k8KA0V183ErnbzkaZKO/kfI+p4kBD7RQu1+VGLEUR
i7v0kEEycx6Taozyo7ODgCRJ1zyTr3b9D18hdpMIGlulSrFnwpHmp+a/Wt6a1d4psLHiImnr69Q8
uWMc0/5j7nOEkyFciwBxX+bknEGcczescpwypA6PsHvv388mUgrTI3XnxInyuf/4RlFaDZQMxR7Z
ip3Ju4OhLQM1Un8mTK0QeIh7nr6LZkx3MW4nu3LYtwPkXEm76lqz+o9OLEK3V/uyFg7l+96oZgP0
Z9uyZZ/fJZWcSWGCqwVu/D9+tbJH67OnZfiZeQz8bivnmvHEmPb8Dnz/wgwRDv6iCiHAqU3PnMAS
b9zhkSnRKKYXPu3epF5MHQXJFXEGmH1JZt11cjyhtC2p6RnpSIc/YGCDQwslSCVTk3CydjusIt7C
BlWJbVnvWbYDPe+UzxjDqH3vfGEOaXA7rpTrQyRIk/Lz/ndVUoBJaPoazKXci/YrY9LGnnq5nftE
jnpUhkCDntiRQXpelkrItSieyC3rBCyZdQb3S2Huw4F926g9PbXk9IW97fh/th9RixcvmoX7eEN5
g79WYperTBdpr5YtRWb/d6Z8bsN2WULSVHz2sqVO0lN74igFX/hTLtNpQw4fJ+Imj9ypwMU52+J7
YoqAm31xboJahashVNxC63V0mn4Gl2Bewaqfab+KHd7xZ+jUaRElTwsGaFzdVoyQZ9U5RTcqjBnU
Dgi+Z8HQKvtkQF23+VEcIvBP4Ddi0Eb01W3fMdJTqF2SQyuNgMJcL8cPVW2dBJAsSOgb/OXLeV7j
LREUCLJ6riZ9aRz9imkmubC6XowoeiAXnv2/OYtvhPLYIY0b40yehlXduAD6123UAdR6yj+2xs3y
wOSyczoKdpJrwgvAbXUCz8Pu0ANiWXvMGK82PjRpXZ2w75zPn576rBNjt74g4acoszkC81AsUP+n
7cAamT7C4qNdgwYUw3YU6tScZq7exY2/R3EY1YIoB9ijSte0F62uK9un63ck0o/dhJbDNaajTcFU
niFJr16cH02+z61wjDNmt3A8CDqUzFtzaoZFFX5z76VTZwb6XcEkgl2cthYFzJ4CrN/ofHTF9iL7
v0j8Fb2TGI1W4THvFH1OWt/hK5Gl7ml1QS46E6Lf2Qm9s1/JZz6V1OInVwvAX8O+u8dAFmuKliqK
lSdD55xRcbHX0OqvtGHeCyO1QHlhOh7zsDa2QBjy1JLa5laI+dNYxZcWMxSb//xxVto8xAU4S6YV
57/1Sf0g9WWKoS6tytjqk8dl/tzbBpcOZatG9JmYqJ8SUCWTqbaYwF77cfmt6RL2U09/d68WrO5L
U0BytF104xOzgKzMYf71cvyToRruU4qixV6Pr3o5wYkZg0kyVvgLUbz1PLUnzNgzKqPAYXlczSNM
2TSl6K0LkkFxlsPcI5qYBLGQFmaiiAHRbgLZeuVforwIeuUbXZCqPbNIQpbxL3Ipkeb0PVXbZxKr
9U8F3cPcNSQuOvd04jRTeDbdrZZI11uZvtzvQ3EmW4RwvJhUzlC5kRBlug95kSVtLbWaNu5fjiPk
VK6DTjrZ7fU7VxbZbYcde/h12nlubh5slwWsYpSMuqidF12UJBNmlLILF4t6cCMNERFkUCQN7U2o
uO34YlOSI1ee9dijaUI8Qrehkh0gyjEgNag3x61hJ6QhTqmIYneRFJNBBD6aGIlprfti3LEYnRW+
tpjzkkb3qLbpoSNjlNcrYYtgkpBSfdwxEP997XnaDxh2kBa+12k3deGhbacyVH8KTZ5ytCMMcbOM
0iRTqe3Oy/7c/4eXexgierZ59S5xVG0OA1k6sE/9nsxy8sny7GyjHsxY8XrAy1W28RMwHQsCqagl
q4fxtDi37ZLICsayMwoLd7l5QTX2RrgpWNkiswn+avbI70N09SeS4rUf31lrqnkaG7C/paPY4BRd
VdrzHNP/lRi8ycAbvb/t4rS39Xu1+Ipi3hIhe8YYIZRQGis8z0rXKXYOHyBCdftC7RabHEtCWpDv
mxzNBW0e/8u8A1BkUj2ArgcvUznifanuLelhscaSYEiKFfe2Luqex2qJ4HJSs2Wfb6CbpqVIt64P
de83l2xvzHksh904C+SZOMyHlWciIP6bH7vzbTKv3BjY48EY/G7gCtcg2embRLz+p05eMaUJjyFc
/OT0y738oe5MMGy3ox8Dlf63o/glWNmmOBQ4jP+qiCnBLpx5HYElmu5lBT3UZrtGW0U2bBqhZPLF
m+RtdMdZmhjuoUROul4QMUBOISTIPvs2pkbUl2YM7VWPr72EPBrmq+XZ/8WMWVjM+ObuRosK3SR0
HjB8b/eC4K/615kgZXL+1B1+nQg7pFvl/2UOaCN/cQFCQX/R76t3SsK7dijB5o5K5JqzqIdaV+iY
zpGfKqB5OZyBq0LeU6xiQ/Wf0PVZbNfI669APsrwI/4KHSwmavFC6BidXne1SwdnWyo63AIx4cjn
KJXRNCjXr27/3qWXU/imm0EpcvpJE/N4I6ceBMn+4zrfuYE7exAfmbNu3gt2YTrMIVQMxhVIu6dt
l9H7hRRyGW/HkxZgDTTu1JC3MDFAHPN5M7lEbPO0h6zC0G+N7eXHavOTwSvp7nYU5K6mYDDsQRRX
T5HL9Rq1eY5f9yiYdplWxq/hYhM5on66JgFz8iaBIlqRt310FcN/SyvX8p7STIlaRyfIinlSUA1+
PUQtlf6O45TfIIMVsGdgL2UPxP5SJBHzf6h0tERXWKkd/ovKwW7lquAVKM6B1pkauPZzYP2cIqAA
iqGEzr/7Vxj7+FhXVjgpUmVcI5l0MoZ+r7WOhQtotQpn65vg0ZOiRGG9T5aRY4DbtRFi9nHdaKuY
oaSnLwbuocUJNyPNCd6ZISutPMLEq+FPrxm4AEqsA6ctSt0exMZX7p2Qf/ER8h+vEkog4BkJvSid
5JciqnunSw+UZvvKdhRN9duJvJHRKt3KSsGgNz3JkkTphCcVChTO4tZQ4qlK0inYaqo+iVndBBgQ
zu1iMJAHpZ2arZHmx2yXN/7W3Me/nsRDmInFX1ip/e2lLjCSAD81a9bwMEbFhsHr6MtEnI4HgLuL
AkGJFSY4t5Fer0NrZyuKpJjOqGjBWqnLFPjYj3YxuzUbR3rVUR+QKOtlQmS1trc3OIyxs0rEo/iz
KP1Tk6zPsm1EHsI54JcD4nsu/TBstE2debO98Mglj2nGlZC+jiGc44lH9GlpVxQDH+z3ESZTbVGJ
dYXsTcVuo6K2l2FYkVAnu4xH0TxCZQ+rCDApjxH5/VynNKrn3/f/wwCzqs/f/U2fJ5vC+oMC8GC1
ZrQB4/FjJgIrRs4d2Mh045rJ3+jXLSoedthkvdXj5424AbZcWFFKUcjnAWcjJUGmRwzyr1rP9Al7
ZWY/mQGOlNTlgQkzSsq//lm+ryAjna+w4HaaB3TlRQINFX/uvtOIzsIPUKnTadmSicwj+a2Xy8Wf
6S5Wng8cp8yLOIDz6X0fiFhRc6tcmswXIeTBoXxsazA22dbWfF6QqLmllBn0kx7EHgJq2hEQn0Sb
F5TVVRpA52Yf4sncwlEUa83KJ43Kq6EstwlpbJcJWWr1jiHDQ8u0dmTPxs5VamMsdpqo4nIx3/Xu
Zh/c5zP+h/ZjD/oXphEuDJSj/3OvT+IULc0RyNVoDtRxqoToII7JgfvHwsxtZBFKBINzL0j1B7Z9
Np+hxHXQh52Feh7OymaD98pUaWcJGLjE84UghWciaFdmupTadyKIIIdKCvxe2F2M1BzJBrQiHEzk
MJlwt3tLOtp1Ab6XMdtaYzWGyDRjNRyXI8evj3M3FnD1COKHoIGJvlFu5+YzbM3bk3NqaUjfiCcK
9W0+izNirMbwmt3IDaK+eJTfwn+eAAyrU27A8DBf4FYqRcdLJ3OWgtEDqHOtwtNQ7LTgoVu6SUho
LxKfwX3fYDyE/CifTfDvkYgxI9YtDEsuMEwVnZlyl2WWZGHFvoH87Yl5kXfz4U3YQjDconz++nK4
dKpGu97J8MU/aevzYwRkRGCo1TxzmRdtSJjI09Um1VrBZmg6Dfv+sLQUIQzQqACV9rD7HZ3a9uvt
wouhioJ20WQ1RglDEPurx/Dlxo/+g1p+h2aKukydP2tX1fytArlj/aG99CU4CzArKscAjTUqByDS
kFjch8LuyCZPjW7vFVmC3w4rynSc02e3MsakRh7a2lJzOrmUEWsB0DKHD0UbO2HvXY+qGnYXeNfS
HhQ118Yxk+so+JitWbRFOfwmMjg8r6TlAVf4sqILJ0AYV21Y6pl/Zx7ZAEoKkKcLu8kkknxAyBtB
y/t6P6JWI2xB3GgPTo+yR10u7xy4BC1VAclWsDGO5hc2dmHR5XLLfv928FTcxTwd5D8+hVlculxi
zfLp1BiSnVW237V0E6FBvz6sW3YwkSVsZ9AMVdT94LTEXYJDtS9+hd6j3vw7HQZPGZjCOxcFn5Mp
N9U1W1/jcTD/yW9Cvz8SnOlDV6CTVvB3qrD/kQk+lJj4OHF2B3vfcSxrmDas7dG/AWeIM2iJ6RKC
BUYWPHkZpxyW0aAgNtRV3FZhfs55+HGffjB+e2K+H1OJUs2V57UPtpltFONvfNIDPe+KOBP6Q1gg
ynZE600O1lH03X5bb6IFcrMyuNYAyAnd+GYpZuhbC2hp2MiKF6ZfzsJ9A4SQeuFRwCX3894wHCrd
GlzMNCQiVxaHG0kOHnXO9SJV20NaWZ8P/VTBv7vsV1ihMw5+HxAmIRM8XAuNcyb3MEXmILicCAWr
Bc6VsQESWXdLNuaLqgmAdeE4Yu6tWP7e/nyioXlnWfJyfXkw3BdoGem58Sy4CA7s3ReUrTA5fJKn
GXnYSV3WLR18q556xDylCC/vK8Q7ggTnSpF7N6TgVggiT+BOcSCA/Acay2Q+c3qDD2whSjq0f8qE
c9Hg7faavTwKy4UoPWohO+32El/9JBFtc4F9Lut2Eev+6JM+UgVV05szlf20idewXCsuD+x0bmbI
aVZUGnAr5mPgAikOIK+/e4WN2O2dTy96AYoxi7JhJgMovL+eg8OiRUWQQzIiCZMJRUEciJ7rEzAw
NE3o2rTv6tB0hIeDGBB1bsndvrb9H0skZ80S2QCuNv7RzzcyogPNBpsKiX2W+taA59dUZC5bEE4P
bv6HkaVxd+fhhmACHk8pUz4mIB7NoXF0lktutta/FoM4VAa4scJO4q0+SCwzeCHj8f8A/UhEvs2E
XzlYrtV+5SqreZkZs2BeoHh9EONRd7gKKfIbFdnSeGDkOGODh7ZTK9DekGX2TGTS9J0o7LuurPcM
nKOu2Pp7dFVZ9CRwCWWcMHEYtzlRXUP2OKbtn553MgnMVvnUzTUZm0ltxDgSlnv9YnsPvXz+7wT8
SJskkvHTCLij/XouqWe/WoVU7H+uwZa5oIp5fJbejjkE+8XMac6m2IZj7I+A63a5sUq0/fB16hiH
qBmlaGy3aRft8amV3sUWT5cxqnBrFxx1hZzovqD95Q5aY7x/JhpUBNBi826zfigG0Ys6zcqGH5bk
3aDyC0ZkeQqTWR/q5HIrAq8c4t0ZgStrETmY2xRRzZkcpKeRL23E7tXA+xbwW6HerzcR1fOCPcuD
aRtzfbhPttiI6sYab0LsxTBwhHI3MQYWutLcSUJMClhSIoLuVonM3hxWVF0nT3TtGsx9gD/gQ/aF
xF17mpbKAg0sp/X0qg63ypjtNXMfO1jQqEXF9kLlxJCEwHky9T7KD/9HqyC9qtLBJAq+zNFiw6Aq
GhPtnQR4kcDHCTma1CND0TlBbwynWBIU2U+pyc0BPXIUx1Po+hGcGvMXcGOsnnc50d4DT1iz0zae
lDFVXDSdLS+7G3vHkb7tGt2J3GuC9XRUWyExNT4XNIDBZfDc69NI3OJNmgI87Vi3YlbN6uHQP2J9
Gwf2XBW7dhKtqCOnM72Sav1PjL2Wplqr3RIRWw3CqagzrqO9O0gv2ZWJBC+1FbzoDs0lx6ZtDbS2
8epylpYjMk0GsV0BHKovkytzew8iaGfBBaGvuY+JV2EH4QH+pde0CHs+dRrY+aAKBaX2EVqv39pb
8mk+XTUto5TwuEy6Waq3SWhkHRth09MQltigQtPosoZU5G9kbeZHanPiv29hKN8+NyOM7o99gxNU
jJOo5cwp5THROd74drOfK+Gfk9Z65hP+6GFX9PSBa6dc4RGCIVqkCD4qZGtOQsBRL4T3iNyblEax
rIFCOL42b+Ospv5OG3a3quskFRdGpzBe7dP/RgRI3VqaDKIMQKMKPgIdkvpbuxecgio6YKcw41FP
xlFtRzh+66s4KBTvVl0MorNktJ1ahMfkxLNjy18kB/CeNInQbGHnU3rpY3mXhe367a2epbj3euBn
6+qWmLfjeFfarBV648jgOgn7qjV7BmZV8acNiE6fBeloPO93biAO2zB+M70+OvvfIHcw8qPD2jEG
awp1BS0iRrTcoMNr1fM7IvvucWHBEOW5um3IeIUOd7Y3IkcvHDzg8m2rYm6rA08sxolzfn9oySMh
E+yqWRDD+qnA+FgGGGrZa6zUOejND8YBMBx8jhmYWOUFOTVvWHFgdqaH8Bs70NzoDfYD3TnkEevy
Pz9QpLxACR0iEVLpFydv4VczrIEirjbEMspRba+g9OOjxI83Eoh48I2eW5N5+4aayiitkWfBHtdi
7UDlWbZtkGPk8N4sHznF+H4jQsNMgiVsHhVKxokY9mWagBsr5QwARuc18xtemYQP/NzTeFetESUo
YWFJxhjh6oeVhVCuOgP8Q3YfBVgTED6ED2eXTV7WA/4lMUQh7mJvNQP2AJZHmGFMywTL1zz94oaU
dwv7miaaREw170BDJxmdt/ybB6Xm9VrFEDwH+a7Qt9XNqHDZs8ijERUnzIVWYHmz3e+d2Q/itGYJ
bKdtA59k1xc8P7cDxwr16yuKq017+SDi56+Si24akGTBc5mEuP90+vKWnJ9Wc0puuOglozwUnCHM
Zdt6P4R3JsviFjUmsdIlEysHYeu1CixLG6oBMiyEALe2kDDJU8vLaVWrOb8Wa98YuRSZE5mmSeQo
Dhw7ADsPSiaPDmI3xbpBpnjWT0y0F/IVseZQ4Jy74soDtYEnlt4TPGwGFuwiqD0byCV0RGAZF/43
VYd5TnK1PeOzObNJvpMLBf937jzrlHn7hFXQyU44+G8RlaDaxevObgjz1HTHgfMREt6xjUawajXy
Iqof1kJakIONx/1zLgSCxCgFQiNUX9kkw8PjlRLgR57oEhsTiCj1SVIG/POkfyU/KlrEvchox6L/
7hWvMj+3qVcXh++Am21NWe5EcChYhUGu4Z1vhOj5OubdiR/J7+S558RS7+QFpTqqgxhSsUiuoPOH
W9ZHmIj623HAgBii++pBCjVxWAf4G3UujznWfo2uEOdpy4hJqx929FAWHWIOjqjNU5hw1eksL1bd
8Vl0l0ln/Z9sy04+ZpKUmcagZz9gcOfTFGwpxRIe4iMDnLNKryAU7M1+2NtDuyRm7UbokR3UZv3w
pMs7MhhuuLgKEyIX087VNzfruM+6+7fiCSFcCv+ni7k+OYk9Cvfj8JOlTVj58AUX5yTBuV5RCeau
Os6f8qM0zb722lspVxMriderZoiYv9E6in6EMjQMq06WN7c0A0215nj8mkhGoupI9MUh+dA/1gXe
VD4CjOyBP2RBk9Wvd2ahQ1fEqBB0LJXi+ozHSUfdD9g87eQCMIIC0OEtUlMzH688tSLsZ+juVl6I
wEbm7Ycyfa9ebSXFfDgcWPzQL7Y8479Vvf1qFJCMlQO7TsjkzWe0aZqU8grEqe+96AsZjqmF3eeY
NihRuPj+29pTG+EKGFvdbdFyZDcbCPjx99gHTp2ZnRfkga0BRTkK+nK5ldX2cVKVdRGFDDgIjHoO
pK2B40TEM9tEuT4oTMJ/S2VTPdedqrUGlhHeuNI66DwIR2LimP5bJ6DoYSggOunIPgHoe9oB6p19
HL7+eQ/z7rqCq4WERoVvNFEPoXATCU1gK2PLHJI7H/ze5eY61X8hNcjwJWCtVVXyD6LeTKNvsWru
Xpyi7/c/ZY3TKqVMvZocDFbw8XtyM/XvA2sFLrHSRuJMKh+tmsQV+tTYhfvDSvHuYMffaMiDseLj
cRXtHh2DiIFPAjZF5RrJmmhagJ/ayng6YlCRPOJvi6+BZwsl/HfCrtJS0SaCxB9hNN4UcwJg6w5b
GhxGwgaCMqe3yw0+ZGU0hxK0ayZWwz+fxNfFqJW2LMr6cMAcKzTI9VQadb1s6Ozt3owtqSwSo39+
IXgVcXbqcmvU6M1PrWn9xHjlFN0x+irWpOwMkiQ9ybWexGRUxaDNEGWF91sXJFQjJ0TF23lJR/8X
saeRkUzQrubGbB/itFurF9Fg4K0SQ2pVotYuaV8FQnoV7wfcthdgJJw2b8XG3kzui3qiRr2LOM9n
D2vr66Wx44nbDKKQmRVpKHUq/Q+/5ETm2bJiPaKz8miRZCXrEgNu7ffgjZ/Dlw8X+tIdLNdJIjq+
gbdH6Fugvv4RHWoTmWOfLAmBxIuVqZKibwUAyI9BMPkfkJ+NJ8Bfl5lXhoLBhQ3wHxIkDAJw9I2e
x1Ty4fPSeIaze6YFqtN4iPMEmubQKVIkF24iS0X9ujjsVYzEWsNqi9LLt2Tz+/H0AjkQmz9kNKYJ
mb84HFnbA99FO7TSLg6eKB4GI1TC5ZGcKf/ixjw6Xuq28JPPWg5cIJAzl6pY2wmszQei2BWW3O5l
FZDjuO57obQYy+9stO4CbBEHxdx+aUMH0rJir/amjFYUTQQbnaoza8PNhod35t+BsDThzkP2ZFN3
vN4Co4JKbPidPMBkMyhldMV6TrktD2MZv9/6re/u+1mzQTmuPcBwD5bsI0T5v9Joa+LTvpSdjGoK
D53rcGI/GpXI8wWe5m0gEUGm8ZyGHExYzuMhInC7f5Rrvj89ClNHq/IS5eOyTF8Ir2U9mK6lJZp+
4QeIhctUP7PVG+NYLRBj5XfGJxzyaKoJMoVxoxCZlyz9AU/2DfAaHvK41m9+v0mW/ip96NMYs9j8
yT+02f/sZeALhPf9M5Hs2lSld0V1+gFlQT9tLoub903oeBc3WviA9k67pBeM6wWV9MG9CNOkHtlq
PdrT+FVE0ZX2CDvWuWibv6UpkdnZcVsaOk6/e+vrtW7HC/ZxlneNOrfprgXB1fkfmSdupuubA12+
77n1grv5WawYzozbEUccaZMCJb7xGymqeS/AQTNz0dQYwzxoPMQOOpMxUc4Isr+6la+CcRBECNY0
Tg6EWLOwgM3DXCefUhtHi0aJBFw3dkFFDvARyczZiKcxSN0agDbrb/nLhkHs1hrkmOOR4tbGpfiH
jrcNh6HxZGipWnxLUP8s4Sy07n7t+zywCVoTyuKFKlwawnK/HtA9KcnboF1ji3mrnciu/7VFFeRG
p72fuAmaUPghKgjYad7YggeXTjn9jqFFQCqM78YMyAeCXMCxHKZ5OmHTA/hKZFYsrJ/xu7NtIAUB
JJu7YNpuDOv/iJCrog5OfTKm4nvtScTuckx6OnkTzL/PdG00cxW7WSBcCjhYHjSf0YAR1J+smVXI
oRA+V5dFwUgXw5CBwq8zIHj+1aGLKc5PxCF5zkTR9FFuW+Ph8TMzHCpbLXeuZjZ/IFjhG464Aldn
mtqJQ+iw6zBkEHSy/Fd6ARNQ/QlrMA3LJ/KpQ74YJQkBnsjo80Z8BESm5uZoJsBeu4jMukBwZLlt
Sj4dd1n7b08030JbcDv9rtBcDJ1pa4O93s1JZDindTs2FxjjJ+U2JTVJRcNfCDCvF1btpEKRWGvy
aqrbGVLtnX7QFWC9wjtZ6zPCjCxPrM/hzEqJDSNogNRfiX4QXpUhglziTUlMu411w85qfbLBw2DE
Ax4f7UBVatQVqWH0HgO4EM+MWj1aT1DoiDW7N4jxmwxoPkpY2YXXzbJc4w8aYqMjUPia6747Zu4x
MY9P4aIiG1o1ijAgd3BmEL9Yu2/JMXWIAAotq7bxyUyIKkbDOr6fxJ3Xvre33bA4FwDPmAQJcEBj
ETvn4yIeJrMGAJSncCslllchXLQbO5a/XjiJIVcwCoK04w3S/arYXlvK8mEuD61FpDyKsrkKUqe/
d22ypIqwh3rLOQVEOdBmxsrHM/eO9JNAqC397bpxN2JClBfmXhuIeO4oqHPtDZYcbc5U1yoBc7pr
N3K4wzm1iH/DmZRLClhh6WHD/d/M3MddKU+rqIY+VEmEbaxNtdvozAI+sQFyrvJylEFmn7S8S6TJ
l8C6Auflbsd+2jA7UEAYohiklhJi5Ba6B+70pmr9L096WMpLOljM9OfmtTqsqcbp+CXT1Md5jxg0
uUKI0EOyLKPN5VivibGrtyi+HO0UJv9GmxoGiGfCbG26095Pt4Usu6VAiiKbj8Qb8RMgSkv5VYH0
uiWzjz4xGHquMXn6AGBC5YWFMfJ5ILWrpCzLV16aX535n6b4GDYfsg+XINVrkdf2PkB14IPP3c/s
wMQ/AfomemtZI2F3txALXVbLrO/osPJpNFvjMK2XyFfnXUk8x0Nn7sFiuswxc5u266GDm7AEftJc
bXVfA/VAmRGkYz6PlVgVx9g9RkcZoVGs+83LSmrbu9r7Txw2dG8l4xPqDiIw4MIbk5ZFohGxX8Ky
CY6EDx/Mx9PwOdEI+sjW88v6PKI94nsahtULy2lWRx/A7UuAcCgJQRIRabWglgzojeaJCkDcZy3l
IBGJNP6a87DQJo1zKFpF+GIU2YZO4I9B0jm3niAQfm/KIE/YJi7EzxOx9X9YR5vxBHpgn1HoZFC8
/INlp+pICBOxD9lXLqL/+cHYk2ZRprrrnKSGgf85iy8suDmMMfNGgQU4qmrj8lFS+Kl9KhtdviZj
NoTcmNkrx5EouS1PDJOGbgv4cHRVvhSQmhM3sNkxP4peP6hSe9wBBCLCcSATQvKHUlwwVFESwx4V
yTOr29x/2s6COr3n+EvWkrnB1zbTVS8LZv7Q3C7Pw1ivXzqNOwDIqHAL9UFg6xI6+d+0b+jM78Ci
vbTp7uXn7yT1afEcXIMEMJOSqnB0YU/juGA1wt3LOxxm3FY/YF24o57ja7Q9EkhyUzruKssXyTlJ
C1RBxefRxPyzkoNGohyih/zq4BNeKy10dyG+4XNll69whkfeEn4/NKRg/uvH9LyquDD7N1stBAU/
iXvDedA0+uQjLxuhlfpXuJ7IuJgMO+N2ZQe0/DLmKRu1yShBRqFs35U1YS/SzyxvwBKuOds3xtI7
t5MBDOf5EWAsit9+06yP68DqkraiOxxMPZPXqGc0VWK6LDhRiU4QR69ihIySdz7VDyY58fjLc0Vi
PxvN2CCcx0QjZjO74H71H23LuN96TAfk6v8pEayrSAqAFe4do0/WBOltX1L9CNY6aXumnxLyMRKn
HPX4x0Lg2n5qa0Krhk+p/aWmFSmYRl0kcZK9bwqIa599/VRObAjKQeh6m3zaTC28gHXOQ5sYh8AJ
ZqjY1VqnT0KaX2Ab/HFLgWTscxcLCWBhZnS8VmSA18gA+MNGl5ET4/Rfog2wt/dbOFY00T36a3M+
GS83akdzotCFHGkbmgOoHFHj9DRMJ1kQu7UrjB0VV9IU+crAaMxIyNYAfv8ok66SLZEgI40VZF+I
lTy5Lqc5P3TAKD7EilX7tXHz7u/Zyji4i1Z+9SmaNTm/hlSHGsD7lobv6QZoEvffVDhZsm/v3FyY
n4/jNQupM+lcEsPADVuleB8uy6c6WDIjxK783P5phdabWLdm2fRxuJUlN0WUdJthB33J41FxC7Tm
kxMviseyXCJYVEJ/NNi0z8tdFtuhvNn/lKX0vSOTQkTKVRTJDC8r3a/3b2nAMlWNXcmjl4rfyQaB
BO9CmZqB4PKfx9RW6qKwi/FEVLRAW2mUYxgpXQBqS4Fzrokcze4yAktdlFwzygjSBVftt5s6XFdl
jUeuG6MqoeD1j/04gLQYYuIyYd41xmWs822r34Y8V+1DUuDeXSwZ1yUX8J+O8CWLLIRqbj4QWQYS
HBquXqX6gWdJ+5/xcpWC21m/mi17Lc95V6pIvKqJohTmOAU6mosxCRJlMeo3ZUhhWrW+ktVqgIU+
+i+qtnkSwPerVK5H4JFDOfLddWhYYR3tCT9l9dQWu3u/owWXL+ruil6UsU2xweiKvNg/uJJ/eQ/S
dL3dSk2CX19/xJDTTyMUX8x/14MHmzbgLKWvYJskPAFhi9p1jkBT6HB5BZ/QeFix+5bRAfWzT1Fi
ilei9p2MLfgGGvOIdrnM5wfeIpTGKb+S6JJHHeRo8P+1N78CXu+dr3tSl+v19h0lzDgT3elsrNCi
li426zr2WuQcLjazq8nnRy2C5NOB/MxymLFuo2PtqQvJByxXIOb7O4KA9ax4lzhPBd3yy6dZjWUg
Ua8nHZ8XwKSgcnuErbSlvTdnAUlJUQwoHhstXuD0UnubYQjjtc9X5//1frA2BouJDUtgCu6xOJsR
+4RY8T5a9U6jwha6UVefs6UTKmeK/d2uTwV5sNAUbZvJH+phWjw/Nut/jPrt/uv4LjEbsBgxZTy3
xWlmtfLmflTe2Kn3ayWAFP5Wat52Dk9sTb+jhk9ZzXYN0kmF2pOAF5lJWDKr9ee1RGpCEppFfizd
CK6s4qxFRaKf2qgsJVc4xesDo9QBLTgvLiq/NDH2/T9y2yGC1K80tKjdwsezPzYUmz6Rfmhe+eA0
lI/+1MomydVvrOorHy7AurWLOTWR8hP1RBj3VPBXkoM8LeYoFE62Gms2HNRY4rE6PelWaJ54HS7i
DHlcHDOkEu1W4igFRHO7cQnq3tMkDwCjovFhNeTgW3wSS5W8lHb2uXyEH+L27xvsg+WzyQKQKviM
lPwRB/Vq9qXES/b0KUxWuxFO0S7ALUfxjq8nK8m0u4YtoLXolcQOKk21YbnxQxa+F9kZfNcfHftt
jbJzbfdZJhwhU1vYYrX4vlqpmkEeMehUTy2emDMUUxmgZZ5kCQCS3wnQQQUTyQmmj25i1NUDWMVL
R3X5/iuH3m2PBCs0Qvsx9BvXa0FD2PNp3S0s5Yn4o8utTQ+lbL1ZON9dSFAog7bCAIbhkr7I/2YH
NWvc0AoO7zJL1fUaedmrbPrhPJcZ+3XN3ctcp3eoPmxAfjm6u1vUXtI0nj9v0OPxFR7T9ORD/bYw
w9EFZotmUPYZxJpmJqS9XkORiiMwPzeZw+LxbKSdMfjzJakCp1dPVbORihIILnIdA8AfgY9dMkc7
ZZYxnrV5pWpu/DzrVl5uVEeztfr7Rt8vytNMgj4xxEWRoaaelY2ccVt8Cs42bIXf9ZhIwkUo9lKv
9bwW/AkruzU1w0LwOw6zKx5Z3zUGCrzfetK2XEm4SUISPPTXtxmty7XsJc56d2awLGCp0ht6/zcn
Vw8Db33tL4QbVzvLYJVqamaD0MWfaBvdn471Z/OMZqwDzTqRONBqm8ovHCjsop3uWMIBlQXceALl
PVyXvD80OCVRLsWmrHYBa7MVpetQBZBOPuRGIoVlillrbktloiW6rHgkkbpFY6bGi+woTsnmepDo
yYUXnPlB1/2N9CsfjnErDQcjvKOBn4L05wR6XJorNRgYfJHqgfIbOBFo6NE7nq73w7vrezCATMYR
bx61fVWdG8b15Lbl3mbESx6/3DUMSuWD/Tczbn1CAHlPKgW8GjnmuWEm7ua52WDCMXlWs77NkPBJ
vHm8SQDHP3epljb20Szc26iEpCUj4hm/po6IOag4ZPrtG5XAEMJjB0US5F/yUwygW17j7TNjlhl6
A0MDzXq4AM8ImDTb8O4QhX+3SPbCBGdkSiaqDSDBdffd3s4WmcAN/NZ9W39nSlkbIuweAHavUIT+
EQl9AoP8wMIRwKjMu0TRpnpqd6iTIi0dZTtGPYcp+1E6HJT3Ly1hC70k/1sgchFDbQxJb18z96eh
aJRACmThDfqAz+T8KP4+sXlI1dvfyoYJQhxoVynBIwIXv2L+i2wze0Ba0bMEe+P/4DjYHRpP2Rpa
A16I1JmYdpl2huka0f2YUkM/EvTwNdbS4RqRiiQQdwBYMv0A8wR5Cgde8XeXI/HgbdS/j5aQVuR8
QGUFrwNhm8fqg2UNXjKjbB4qckK3hWOJkRT+SLvaur2URJE9fzcJkici4fpzmyMbRJJYoRRo0kjW
6G6FsvR1u0MBQC7TvuHGqLWGaxKYtVlKclgUeaPqymLqjap9J4LZadsKXj6L48b6w8Iosk3t5lkB
Vgrsi3a/hOuKPsmYsvbkinSw+v06ETlcgwtwxDPRPqG+Ym4J7JmaADe8XU97H8Wr0yrniDhZ1Tn7
ePNaycEj50s6Z5351RSjH5Rk8eurTbsDrEZgUP+VitGDLIjJLiYKR3v7QJWz1ESpBK3KGjKpIFXZ
9U/YyzMvUudl2o3v2m1Ri0Qbrj83DRhHWMTHSGDmJeiVLo09pmCa1hVDFxC6xbHQE6KAEZmEDhfC
5IUowyGXU7y+Fi5xHZ/272hAnO0RGTUiyGRR+CbXAQkc5hs+wzRgBesp0E7Ik8TNH5ex9s2Ppz9W
2t1ILSeAkCSbD+RMXoMA6h7dFiao68ZYRjUFwYDdmAPui7MdfQZBqlz7Ag6abtANRAq6rW5t7BaM
yVFf61SrwJ8bJSbpNmT44jRHxLQ053I8cwowQx12tlYwpxXRO/Jq7ZdS8Hlss5qJDCrUBgp6bjVh
Os1TgfcvztALAGVcFoLb/rhFFBv+XWTP1aIpj5Su3WHneJGkc/bbw2OdFY9IHVmwBeGmnNgDlRJo
xxRX/QvwmQhUzoZSlSVheuxA/B8cIVZ1IUabqDwMZKQaf3FeUyo7tFdeS8q8kdusy12QEhZqcw4z
/rK5MaIv8yywze/w+GuAYg4jKaazsoz/piqevBw8fodKC/y7PYgfUlbUJqQ+NxQZqahuYBsxteuu
kD0Wx5MhYx7D2oX1OM8l3xo/dJ6IeoSL1fdgAKxrQkvsgKAJ53Zhkfou7hkVvwPO9fqP0xlz1h62
eoJkMdPgzQxWLxRo+7d8/13bCIuVX/UYrtx1PM3WM/0q71Wevqg7t1bY8L8q11gOQYrl5dqyw8c2
ahrcnCuCg+tHMH4MPJCE363/4A6tpZu/vuUEk+GC6sPJXLUu7i23lUoDLad23vFY50Z32HfBHSJV
PDeWJT0QNOxw7HzG6WAbo2KzER+Ci8boDRFQUr5eGyU6SlWaU8079VbdTHbN3nMS5viupIWunC6v
zysy+O0SRPWRsH4LpuPXeYMJd38+GpwqsumwDEMy7XO6tKu/R7n4ueeOvB6kj+fYlxBBCicUTAJW
vdQWhxc3JeqHd1ZGSYI/+iO5kO0PIXeCAw2o/4W4J/X9i12s+FHoGzmhGfRpe6xJUpy8JKEzQqVN
2TPGhoaPipuXAmGF0pY/m4kM10Nb7aVce76TdLmkrhTRVTy2tlHFhi/ZXk2VbBjwHT0EOs8K52kH
NtRcH4HD1XlQhRw1EyGCL6Q8OnQDAMTjj66brpouKnJYoEUMD552ERqrjhYL7l+6wzQHKjE74VQ5
tsXyyKhVt6BBRsHenBW4VFgdSD/l/L4sTouEKGl+2b64fo3MniVnViYvfXUwlJ7TtyGBm0/I2T3y
9991mQj1pYJaFRUE4aVLaGpJq5tHJ+PHfrBz7HVspolHNgb+uaeiAWiWl7Ihz+HeVeXWFYOL2cQi
O/I7/OMqhmzVBlO3qCMc0Q181FeL5TNrMRq15z6D0EK5UmzrWGl9DAl9Uy2BEIUQy16X6od9bH7l
wwFUwKCy1xCwRtLJdEXDLoS5IHDiEwM9gTxZI+ChS2NwvYSQAhs5D1ZnkHV4TQTjrziZE9uP19r2
YQvE0ttDrtGvk7fbNIxAdc7ncmcbbd8PT/wwdVqjbhh8DP0oZAW5XCVtmyfVnM9qevmWHCwZ78Yv
+ji4Iu1B7vW9wPmiapxidbOY49w6I3omry6zVAoVE1m523NgGv44H/IH+O58ne0VKqvV2vaVKWwX
hFoGQTQKH9ZL4uRq2fuLrMlgw0AhmVgXISFf6PlLtqOvQj4SxJn5OBey/xoVft2gBtQT8nreHbWd
h/NJaZrvJE/ZbOnd+dBE4zA81NoPnDxkGp05LoFwz0mLwcZKFNan+Bg38fqUaGkModotY+GOisrZ
tNQbyX93s641xjLMp3gIvBZH3144e72xzyECRHBExS5juGtJsOgoayPkqNlcNdgLWHA5854GUnsY
xrCUIDKtz7zB7W6XwWXDXNK9Uur2NHcLFDlvLxN5qi+8xUm4rBpgSLtv601/c2myWG4WMNGtf2UP
byhNnZeK0b35Mkhy4MhGCwgmYlFmh+0EtJsE1/XEUZxng0Qj2+XQh6B3RwtBRbXyrYlZR66u9s3W
7A7nzz99aa+BDMyIvU1xIlJTHssZhroPvMMAOvNg1AmpSdFxiEDJcBsfN78XtsOrJYjgDP1L9nO8
2KKWHt8TZGkqf6SNlZVTJfxHbX5P3LJoIBuDF2xdwPc1e93+UUAcVAen+brDpu81e9/FbujxFtPf
/ySfueHpvSRZV2xmk3tB4zbCMJSwosdu1z8ipGxp1blZlE9JBYc9Ft3bxV1qchS5gnOvSqthVird
/nAV/eyFecKD1p/uFLDHuftUGHdm6jakqHFFRdloisPHx4KpZhKs64SJiC0O0A6/jZX2t+9VhISR
rc+K+5kvxLLcXerhANrDNcxes/iXbDGFJLoNOdtzFgCmvBV8IacZcLbHAtVUn/Eg2msbPkCU1bqZ
fJZVy9W4ENZVjbfPJbRIpf89FRHUk1/awM0XAAuRxTI0xq+YCdw2TWAX01MTd2MNzdd6UCvziSdZ
0J9+dhhDPktjsC5wk3xRIUHnH9x55O4iSvUCG12nqQwx0z5Pm+XnuzzqMaBy5P5QEC9mxwZgSwn4
rFITQYR4pYe61uXTW68sT5xY4oVNXWbdGCRmiCAhQu/LocHyN4irvOHTglnpaEBzHn4uNLTxzXDv
SQIZUlrsj6Wk/B4TLs5JpySGKrKC84oEJEINteJ3Fp0XxsitH4MhhDjIZk1vp0mr1kMycNxdAodz
bHTOL3pRZPLQO5DCgUIPCtA9zloKtCTQcbr4L+Y4s/lY5LA/1XvdtiKRzOlDYQ0AaM11131pwe2c
V0rpdGM5oOcpNJ9l8SE19cRslSyffilTz2L/yWCTENYmd3aK5oSjXYk09xasUEJxxUVovbl8uR91
wv7xhFXklajatPK++XkcK++4jJwixLzi5I+6+g+OZg0Mxl1Euez4/6cW6v+LpoPBhiBkFYSYK/bg
APYHzuubC8OpBdVwsTOJboq+HsWAY6ys5ii3Agp9AavJG92t5VQiQsEu+dacWiEDtAQBVvu+tMfS
QdtFkIvUrSQCmEPBCBblNtdK0iYP4HGDrQcRe4iJ4IrywGkrlnDhhjrQH6puXfouxklIxj5FZd57
LPk37/msrK/E032jWglL91RwbSUT53G0nZ3aZRzqdklzV0R0wDweQxsAqGlwhyup/C/a/k7mriq+
xsoBVqaJyTG+y3NMJJNTo0ZiT94DPwGZFIyRKHO8eR31rsma7vszvssExx6ZBZRxjE/yKJkrBz2U
FYdtVeWy3u33DqchI2KAChDq4TD47v+R4RPDAlfiam0flH9FL6/gYOvgiL9OpOlguCEKYHufgI6q
hncoER+Xt8ByAl1yWG+vbg1SZgR74Z2lFhmxSSJhQoTITJWRLAUImUXqM0qn1YNyarZcxJVme5Q+
QFvxZtSVJd0dvLm9TLhLbs96M1UBLtQiGqHEbyjV+f1t6Ek7qJGpxDdbmlWTqx0Ql85FVGXGZapQ
Hgy+Am+FiGrxtdOwgw3ZLwgWJp3uF8NaAlVAWlliUL0GBeEP4h8f6SNU0yjRJJs+EgeR/Y1dPv3I
HqvItrEU6lzgEFbvQNJq88DF6Pdr09y+jJIQRdYBoJ5OsbAyjPbNLLWLw2kvPEz7qMiggOK0/EZ8
X+VWTd7SL/ChagrbnFgsK/stgOJ7SEHdDAuPLhiGJ/i1GdR/SITS71vexWryn+OrQDEGr+banVR0
526XGc4gD5P0KIH4PF4tup7htjv2viuW+BFXGXGcVKKUVxDL8rlpOaEPHEERmtHnRvrvKttQEu1y
RZfb3lMuUUExnaqUChe3SK89/D3LSShwEa5FpZX+KoKmuvlYsdRcl4y1+orPMAcG6rHFPayOiMcE
CxQkWNoDviJAmexZCa/jEv5Qa/lIs2Ft30yWA8jHKuJrDrOISLTjvtyHIDWnqHMxa5gOLvtZPucM
gPwWvFds4clj7Lkz6iwPiSoh9QNtHE9Z+3z3cMd5RHjJkXPjKkjBmdtc5LIf3jtRCU6373XS1li7
PJ0UzNX5t+h/9vm8VGLvddYLNSvI22lIbkZnSh/6gDbm5gEpArO+kKScSt0s0aZc5pWLq9qF5Si+
evSd5VBxa+3VVyFY2OnbeH8IIsBjA7MkJ4USTz/nMhjZOfwC9x5zQqHJ0NK+lVo9GpN8N86dJ/1h
VkvhjtCbgucSH3VJsL0xhdOYK2yd5mOtNHqpDWaDvMjSElkxgNb+Z1/gNcpM08IIqNn48fcdjj90
qO19X3oaJ+drGesn1TyuTyXWQzBTLmYrBPwlxKCLFmU/tC1H+C11YM0bTS6wQVgqXUhzXhxsWHui
bTc+wfz0cB1idOu5ouZYg00GRcb2PY2LUreZ1AkZyH45OSYn1uwfN63y6hUYjyXjr6RYg4g971O7
1RK1OtVkf7xU2NODnrsCXO/Cv9m/AvOZGMxyWeU8z4npeTRKbEPv4sYbgAMUXiD5OZxVxN67QKrX
PLhIlO3wGhUGrPmrSS6QdhB2kBhivWpEEOZLIeuooZj1//09V0wOF2MBhWs7nKhYqbKvGfdeZNFW
X8Hd/hz71DM2uYkKPfMrUWc13sPqKG7Aq8Vw3hWDDv5TY+GoV4RcbiaIJ+EuNt79ExprwoWfvoNx
H+esL2ASHIKyHnbNRgUqpWyIJZeVd9IJ2ip9DWHwixyagWrAjOsqBqjpubkjFXF1ugf0lLLSef/Q
AA7JqiYYjt21JFz7SaxcD5Qpz/wT9tKAZ2mBzs/nmHzuYlFQDWfuwMkY6a/MxGEHOlVKu4kuF8Cf
urqm93abQ2ESJA9j7P4AR06iRl6PNH1MkfpVKlCH5xkrIDSR0fIKA9dPahAAY9myvCIjKsMATjdj
XPl6TI/dth9iBnlft6G5ayQDDZWvL5aAVCXkRxq4DP1KvP5/Fm9P+ykkovrju4dCQuq9a5IEZqIV
66QBQrkyf3E4tgRcZjJHMD4OL5sp/0rpkAJX/h19resATlhjuKX7f8Cm2psEZfOM/7ND1EaYn5Mv
JLc1MUvNUnVh0vOBOk0r9FL4zBPkSs0z36uqT4Cw0cnkU9pEMVZBhIsCPUowDsr19BNPBBNw0O2G
bAamEuv6kJfVFWX8IHNYLdHnFj+QyyA9MDLizHPgQRzFS7q8OsNVAjy5S2PErljotZDri9NAwHBM
6OSYeYeRrXlOFTV6svXliTdCRlHN5njgGmq2XN5hoecWKvqcDqaBAHmtuGVDDb/QSxNYzIaAaaDW
j8Jm9I1pB8LwMW3RbECIhYGsa5qMikVaa2QeaCQ3tsC2MJ1Eki7hL1oG8RNB53hGIuyEEUSBGdN0
1XGJH316C5WBzYBrKfV/veZsOx1smtAZueo1g868b6Ole2eWFKdlKPDyBpaVJ+ddeINAKOAkDUJN
/BcsG+L7qIOxFh7Lof4aC7NfDEDvk/DDT84FsODcKPoBg0njzFb6kpwoJXYenCN1acJwQvi0/OaR
i7CrRyu+LYRFHWPgZaxxfsXaKI8GIWotrOqNg6kwehjjC2YitmeJOuHNKpJny0jkmLeMIX5ltNtu
PJFfDekRayzD3wFuiUQu7gX5ieGv6XQVEGWH4e9OHMBBxeSnDhPf63Fa/IMX3DWNdKojqr8NmMBa
znnsiJoLyI/OQc00uzkIzIWT352RbrSAduvrfBmDgafIzrLeaJxp7JJeHxk8G/Wkv9jLt87Rc/s1
CnplOskmn2KIH5oXh3vSGyfM4vVZP3CuXS5nLa919q3Cr83RU4Rbo5DjVqitS0w62312fZ/7KFIQ
nIzzZmEObRJNChTWRV9mjiryq/MPyfcujydKq6zwqs2hkutVniJpQT1G9NuL+n7JeoZ2diKKUu3D
2wTb7C0UC6itANE97IWK3IyPlsrUiRW3haPVHO7oWdEQFbiXs7jY2NHlaYc1lPtzdilWsiuToeNP
gjvc6BGfCEqPQONSclEDjLVW4t4b/0jSjKFPQOAZSub6Xk6GyL0AxwcFsD0qPkV2bi8YwmZ6SW8D
L3dFcK/SkH/DVX1MH97pJ2EydzJCKkFiqwL9DnuQgQV8FIX4i0eoQ3NlWM8yPN0WCTIcjq0fCCgz
TkmAMtY/wGbKm1kXSLWGjBZabnNzxKO2gxKWk1zISm23aOJEOEZYv0Gk+qUfPFOSbwFHY48GM9do
ivOQwXZdoFwNutTYpRczDp55P8LvtrZFpwzLfPm9AgsU9PzV2IaN9Y8nSAF4QgmapWj4zFmo9tSx
dfMqbcjHFw7FTujtLE3l2de1xJGlOcByxLWEDDQRf8rzv6aKSbb45ZO2F32GfDZHlo9zmCt2wujN
afgwasZ/0cQ/vGZvfsRuZgrh5sJ7EI6Kv+6s9dRzIpOIChtZhdNGZ1U5YJiLoaqLjqX83j4YSs+H
bPag4SbnRoQ2p24Ct3YWaMqqdVGqjY75KEtH0P+47ZGrk3IYPyQ9W1Sn4GNEv4Vp07kpFHBoOgs4
PhKJcXCtLBzDzJDmk/yCfKDM9ItiN/NRFcpbkyZeHuUTrgKEAbO+XYZq6X/EcyWnZONsB11MfESQ
/x2lPqNXRGSbwxIh4H/QwoahmRKDauU7uAghF/ZgvaKgmPjmNPQdcAP4/2Ui7V/XnHby+X/lwvBp
7B19a12Egdr+M9D0ojgtkG9kZqfVYFTIngJfJh8ltMwddMz0UdUU9UYOgo1dqg5Yla1F9baZPeas
FR1ch03WYQEtMxQb3/npc+HXhN0dS5hF6r9rVopBeiM9lqIbC8V38OcXc5rXimmrqifIUZ5kUylL
G+ItLCxYZEJqRn398d7d33uWx/KWOvxQX6bXz4rczbqmaWB2JQE5rnyiG+xy8tGZ9z4NcK64dX+k
NmccjIm+GK8wtguQcbJXjDPifNgg4/LqE7VnLR97s8pImeScnwUgATHaCTMBFCzjuH0jEiVHhZ7+
5SvLhZEIcO6E28HWK1Q+JDonrNP0FUKsFVVY4AuNxOfr137j2auQw0t0G7oXpnfo/2VHwIaXQc6Z
62MJQj0kfveBivrs6OuAN+lu5GIJRizTk4jB4xNlSFc4Z4bU5mzZdZmeB3hE5M6GL8vu4WUvJbk+
1lt2j3hJvpFkGyRt1eUGksPAraZx9Gmzxvwew0GWkIn0frib+NvH6uR9VtntnFvRegO67xp5+pLl
zJFI2nTVGhXR7Wq8l2JoNeM65JQvAIrpmQZPXx0XnY3oo42znz1XrEBh12ol6qDLdPnsyntb6/Fk
0P5piqG/TfIGtteNn4d9Kl22gp7Tulx+wuNmqoznBejIVhqZMuXki9AP8rweMIlsq5HPZ5DWpkkv
VGg+9nvYJz/MlIfwOcDgeEfYIc4lfImJThVsNJez9G3Ng4+LnffDJIixEo3PQEavKTv+fM0WsR7O
a4jtYuCVHIL/x0QrcaJ42RRwEgbgxVTHL9pHou42SPURwEEWY8/2vkmPZGHgR7Jtq3EEEUpj/HI0
/nD48HdWAzabUhiIFQG1eRPIKEuN+ecLBcTAdoNyl/NPzJmia1qq1JtlEF/ngf8ukpnWXUMjqOX7
shWfkXoXiMAAMTGJMpbksghkNPqGnlmXNm8+kmFwUIvI3Sw52JefBPCmyQSRD5KNJ63Z3t+aNN2v
eccAzSlYF9QdTYJV2kN9rtdCqG+lOD8SCc97npBSNKCzJagjwJq8GX3y+qdEVLm4C3zFNTDoNxZ+
yHqdnf20HT9pjjMMJQXJ8hvPmKkx7zCjxyv5HR6/WbFaCAdma5W/U6lDTWboa97K8F3sxqNIhcJ8
sAWHBdmMjYjiGqgeSwuVpZ0X2zFwEtLSK2jFA9G+LWyPaEd9U8qhPhitdms58ik4Z9yxyJrw46C/
lVe0qfCmq5+6fNg5QT2zcbw+1D2PE1NKgQxootvFF/E/D60xqpqK3LGA+7WXU8pYWdPjoEmcNm5Q
5nyNKxQTwmBWmrupN9RtZLF9SIp4D08M+NJhpuBml68YVZ9T9YtcGp0ouBXaN6n/n4VJSMW/ma2a
W7Bcj7Vi2vYz6ZYSjtnoAE+lPBDIJjaZfqLsMRFwVpDqPo1ruhInFvMmu6M1IUDfz2fDDagy+mvo
VA7vl7J0u2kUPraPE/ObKalZIijHHQB7Hd7fYPGvKH0cnr9rYYOSpX7I+JW1PfVZHFmjIVLSSWSJ
lNtXZ3Q4uxaK612eVuQak4w90cDNrmKSM6ZSq9YWwCIko5Sp6q4dOt8sibWsMNKd6oZBILfG1cOL
7cte7ebC6pIKgRKdfIGIfY+8fEcJsJhrl5wXSci8ax9hkkHvUz6meQQ2C9Swl78R03oly+/iygZz
luyAzZbMilsEN5h3CPAxhT/yMLvjB88kLiFpyILF3amuIPlOSibxG5C/66vqV0V9IrSJc0pscIR9
JIj4FyjoQ/kMmLUqqqpO+Zm070TS8IIfKw2rrqPqErBb+UaDfXl3P5BnDFB4JFbUKefROVmxn/fG
WVayyua3xCXEo+hzWQaEY7PelFWrXUmrJ2LgBAFAWaWVlbq0MVMcwbj5lWD9E6CUsASOLauS6NMy
vJ0RRazG2UXTl3Zr80INP89GPevtY4EwGTmG++DUxP+XYh1Bse3kDdNq6KHqoqFXWE9J8dkDMZ19
smZYWL5yby2ecAZj/qZHk5VDT1UMaN4yeZbEjkUH1PBNrWP4z3Luo+oDAmit2NWjIm6DXpbPHsxC
IY4GawVVQ4eNUsqNQnP2ZnikVh50aEp5HzweqP4gyuM9FJYDJxYfeofTWIYJx/OfBuhzMPTC7L5/
hHgWbkrtVsYGHSuJMQDMm2Bmvi7KRN74QvUk8AP5oKfyKY70b5fOi7Ue6UDzalI8X3fYiLObr7BB
8wfT8ha9RtUM0Shzabd3EMWEmIt6siWj8YmP9wxLH8MShAuGmChgwbtK7FAecE39oVIHbuZ9rvJU
TFSGhB21ixUJT3kZY7XRYunXVx+U1xVCrPuGDuVM7RTA5vMqgjcLJjkwNEK28ACjQkSfck+/OXTo
3Au9n07NXU1pTjbLv1mkWnLHccCAsEm1IlzCyCZWSqnjI8P0o/nt+IRlUjpStC6qoBR03GIHvIH3
zk1A827BPh/TTgayAReg9X2QCA6Ek8ITsNJY3C+qvLzBqZGt4HAlN0ZB38jn9axeban46UmZFIUQ
nednMnpm2WZhWhihryYLR+8wzr96wMAcMuv4iy5/n8Zgnvt6gBxh9A+sBvZv7/mX/AVBmnVXUEjG
TZ+psZjZwQnDmQwgdzNjnKKGuBw21WKzYx3WPUkOHPHf8Jc8mM29yOcGpUy/2wU1E2GNE0aaw8+S
L/08WPrM43MFDqs6M9xMC0g42AHAWFRDEO76vYeX28Le5gIxAdo7JSFLCZL5MA7lgXIlztzq1en4
nltXJ6UsSy/KUJxW779cbzbzFS7jTew2/WekiPu4APZ0BkYkTM/r52ibipZ1shKamWnVMjUSX5Ju
6fr2eeG0sOOM5LdM5GqtTWUX96QdLQWU46vmc8ft+KZalT6FqdsQ/SlnomgZ4rTjnYKi1d8DJGOD
HMYNB5SR/Giq5Vch//OjXBm7eBjxU4qmNJNs58p5TskgPG+RY7uaVbUuf8A6tYhsnoScYzlpjGVH
GNA2BTH6E/CLU54PnmoBbosIqjKR821NMmMZTZnr4qaGsTUonrQq3dtE+fjq4dfJzBnqOpF6HCjE
EPrVDYxG7v+3taOZuXHbj8sFu1LReCDGLHzTNCMhoTE84VQtVEeV4z+kzWYTFcq68p9qOMvLq1Yn
Gsqb+a95CiVI8AlufUEvdwv/8tbY/ls3yZi0dfROak+QlSbi0KTS9xL0X2yeHu+92JpM9KP/uNco
Beq49tYSNMJnWZUbMStc3X5WecPl0MpjJlxjGL5uzk3mBUddKAjEj3/2+pseMWx8f20nYc5yR4Jb
v5Y+cHNKW32/cDhGzDRi5lZC2n/T22tJZuR/stiia+s7x/A/KD1Cqr4h9s5Ffx7Z1Oo6OmJ5fh6q
LtU6AMIoLTI4lD4bnPfQ00Toonn4pIHGU/NumKVvAxXPkkMRyK8i3J1yINkaoasKxxQG6X8Qw5Vh
VhitIyRDe0KLR6ICHdGqZ5OcUpCg2jPYw+phlRrqCDz3B7fzwL+Op48F88e8iTHN9sdnwzpQa33o
xI6So3u8tcQ30l6qZPVrbw1LYrxIXOKshnSRGELIoP1V/8ps2kM5z7NZdcfLPI8keWsT8NwMlB1g
sE0blIJu/eikk0IIzQyhRa3M4ssR+ePt7W3HkOdlnjZxacP+wb7sYwgVAyWGtfluzhSbQ1IYVa+m
JN+qiR8B0x+wshdolV+/ByNTXLiHlNjb5woZY0PYGYRxCro436Qn7dK89M/hsRk08nHRVovypw8I
jZ//fTN0jDiDpRI8wLN0X7iglUESQc2y1HY7hqGTW7ieS/7SAgsBsCKi1pHdSv0PE4higm/IZ47O
CSDQA0a8ZBFNSCSgcPstzJQtwBwL1hgvS2i1YRz19NpiPZS8EQovakOpzuNr7bqqH+Z6i3JPQd/7
sdYjYf3TfPbSxgmz7PGSZzuZ6EaAAH2KfqBu8zr/fBKhqK2qECS7dE+aBFKM6PigewRhXz44zFiK
U/IpJK1nkjJPECTA8+J1T53hF1Hh9XL09gcJ9EV3ADa4w1ZR+QlNQtQBg10mqzrJagjkka0LLy9k
hvznhV3YyQMpNUpga0vs1vFPJnnBuZhYDKJ0N4nDugC44KCYQh0FZY4SxRy9w6A3F1mJAfzLkcPX
R+IgGX8QIeQykwKeNIpFJFlCrbaYrG4WnLbiUMI6pSxEB8qFbXkRvjmv4vAEFTxflrjnjTp4nSUV
2NKSCkO5qP9sqmby6InZmu8w6AqT81+j0yJqQwvKwsDrY5A0R+3hSVRMw2iIUYHurzPtLJg9uT7W
h9FjfQfMwL8OCqG8LglgeLsqgqdSrdNYEyUyd8UCUvL6LqN6Qfvdkum57Bjn+kw3NRH1M7YQfQTM
JBudHc/8dvOB6XUtZF5bh8s3AcxrHI7COh7ivTcg1FhMtGl9RUCKZwcu7qHbClY5t1NyCJUeAao/
J4xTu36bUgzcoDr3lMXelLr4HLzQ3gRz7hFIn+R2asu6hyAv14Vw0mrASH+oaNC4c6vz+EPXYVlG
VnESSinziZNrH8y7bGKHX6qZvTULVtSKJfgTh8ox/DXxVHvPowKHdkr31lKF5dTNdZM+WVOj4Iad
QiBqp7Jxp7uM78H0vMDSr63LPqDoga4TYk4ab5dldvlpq6NaxcfQ4jzNxQe5ts8OqL3/AbZfy1Kg
5f+ZOh0ql4g2/Rdowlhw12eb7DRYo/usF8EvB9FQR5w3rKt1SkcQzoYryOUjR69C6cgaKrionslf
JML/k1FCcRtCKOmC+B/OzBGo3o9ge7Ogr+JfQ6hzaL+o1/o/w9H3UeqaFJaIdQPw0ab+vUs69XeQ
yk8MrXIpTRf3C11lwSoNG+LaepYV6GfRcVTgA6QIG78YEmr3rimldTSVnHhtkD7IGgxxaca5CAaq
Ktd8EOh7iemYrqDRngJ3Bg3e6BN3bOrc4AraRxerJtDap/+sq18oiHCE2izLWd6IAh2Y1CiS/kia
+xEcCqnRAt2ERW5K6J/ifbk04+QRAaRDskTdFgWZRsL1WS/snMnRqSSMutI1P9VZwzieH+Ps7ere
IHd401CYURfuozRwT4BeqpmfedzmtJ6KZqZp/T2jA89LozzjORSCjMV7L37wgjprxY13vh0dwsHI
h7p1/Lm4giAJTGvLpcCyvMv+7YzvcbdGWIUNVspjnqtZyzHMEopXEnUJSMxkWrenZ1KrXdGRM3V/
JJqe9BJbh37E8Gpf2MEQci6JDoJFIevP4+MAlqpQT3x9VsmQ7iVC5YsHV+Jk9ZrlqtHujLUiyLqO
e6LYcfBkGPyU7XbPlhNBjGGPdPxlhRpTo5RK8SzFHpY30DCxQJ6INBTDUt5Ni5yhdjtB9rcrYI6+
QG4jMXSCHg2ivMcYsfFuO7h+mrGJJvgZpqJ2Yt3fKyAF3X4/b7RVUVZoT1jcu5C4ngtQWHYQq+67
5Sgmtlg2eJyAuHrG8Q2zUKYal+tP3bYeTguuUgIzRGxPNggXNdAhb1gY91knlbx51/kjsXz7nJUk
sgiGazENoBrZv1pbMh11ahRangQwXl3FXc0fXjN2qRuA/j31/438byfM8EMB1IFtu4N3P9uXzp53
1BBlBhwJ2zUcAYWYnLWPKpMeb+IFOEVichpy9/vRmmSM20F+JXM1fQlCjMqU62WsEm0dgBn4rvyS
EAKb6EaU1fLioiC9yaTHmAxq6VVHn6aRiK1jqFTCu6KK5ACiZZaNsTXK4Uf3r37WbRykZEdrx0VW
uwmMqlcz8VPmHpcd6+nNAba2/sWEHDnIx+r0ctGdAMdKrqb7rBjXyx/wP+3WKmePLspuv8LO6+Ee
mmvGBUHSpfphPTaVqoRV3T7UcDO8KYHqxHWgvzLLc9jONGrGEIaLmA6OJJSce1RCo6RD0FAN1Qko
IThjIf2qnfZSkfHt0p82RqQs8S2pTnMltEQIIusguEZQAxMyvV01xKahHbTEsOvOXb5SLq2PxeQk
GpMqEhfS6MQ+VPzSXQGgXA4qvTwbGlc4ZCTfVgdUIgxO+zzIZZSpSWAU+gkXeF76yirFBAzVWUil
repFZZRih651OZfEekj43rVec3ah4jrxUw2kTys7n47PLQ/EdrTV7Co1AXKX8L3RNgJ8gfp0rp6W
N+LWBAZ7kmgULGGPnBObcDsYX9G2pF3RDXKseoaKUwzZCZ33Me9zZFx7ejyQSx/X2OzJzaq1MWnu
21vWjVI96y9kXCcgmGhVkrCuwhlLgguK1s0eK1ZwwQso9azESvhDX0OFW9RCNOhELxbug2J0b0AK
ZlTNvc0mSVMho8mf0HMUfohzn4LsC882V8tvSCu/qLU6XLS6MnHh4vr91spdd41tnU7YhC1ogZMt
9FGO7idr3jc4s8LrGCvsWDnWJmwvz/JlEM05mK3Ks6Vd5izTtczpHR/RsI2wfMVHjJTSYERbsCFh
WqQASZdq4VmJX/1JHgKnGAexhBn9e4JKqM3ogm0jFvJAGxIK1rT6ydjRrjoJFSpkKYkpb3MEPRgD
K7sTF/UdgAugpGgx7GcSHc4JPK5QkscaTpp/WKK3d32Z83WdzLch35ivdBCv3ZWQE1PxZI6gyCTi
TOYcWOchb+GPhCiYFDnq1y/pv9lzgAOBLuHJq8FbkyV4u4Njhjbq7eNGI3qbzzTXJ4wai0maEzKT
uhCFi0Z9vSQX7cYljETk5/IJoxsFPeaO3tKX3EgFoD8VGQ1Eru6bvKNR5o2myX9oNlaZd0JxIw9K
6bGh+c1AKY3KQhzz5j3sSenr9hg3oFIXDmshWQYhETpj+p2oF6b843F2q5kfYblDfKRHeibJ6Ufr
TYnOJlzDojZhvFTwLKLXhOI4s3HnayyXzTLQ7S4Fef75Uwz2f8LJjbZUSYslMjpP5UJUhqpTtyPc
n3lry/rhKp4YPvCGGZSfUr8bA6e4xyprddsGeRjbUPcpjYQ4aBHsO5416JiHkLi9ZU40F3ak/lk6
3LQCFAAJyGX+0xQm4G/PEz1uQUwGfWCZlLfn3Nxm6wW/XCTdS/Q6OChxc4emxMgC5MdFnEiTIRu8
PUrwUO5CJHVBvWSSx8OnuDGW9MJGqqcOHrcnubqpk9/7yEk/y9HidN2ZYXbHKwolYvBUAu+cTuct
92wxbWwyMw3QOfUXsA3piZh9AcYW39WjUv3VqUQ1a45zV9Tqkoz+/D+Ut/5A2UUPqJwE3QeA8rcF
p+HEd0eKNcs2mSIQWYo3zMjPuHuDS5TGwviCe5oVLenep1P185szZPYvex+PrTJ+O1ocF9J3RzMJ
T5yecey/NR3yWtPb9JGlRRUl7cNkcbiIY3Uynfl99AW1KPcsqNyA+JiK1+kasIgBQyqLBxq2ZjRI
gZicUBLudrDXWLwbt4pqyDUOsn8japV6TiSDywXwJqWgRR0WUa5d6YXHYNTeOSf1B4njd4KHhCWO
W2Mq1AU5QliCdI/aE4zMhHCokHNTvlORB0dDJWWt9UoHGOzQQHugb5lzo8kszybn38o2biAAWd7j
0PvyrjYFt/wKpdVPy+uqLaM4Lu2ifKcZ/WwCQZ6X/yhWR8gVNdF8aL1m5BV3Lk3sUBHKgdoTN6Mb
u1KS/sJ+sncWUJE971ChGapfmgIRzCCKpEZRIaOv9TcBeXKyoHSOCn9awtN0GppPW3ESu0SM3q1V
G1ArYRGAonEqpqyQwuemxJaLQtkHrnhHQKjvhd6nLehyWW48rHb4R+PlSbboLMCbHmT04xU7LgSV
AR6g41rSG8MQ7rH1HV8QyDYRq5LYRdumsWx7yh0oTQcijv9oPuYEAIIQHdjmYiNzOrY5ca4V+rEy
17TuzZ5E1QhRglfHpqy3Sl3P/UYQyC7CMymCbMG0FzGGXQ5dRcMagYrcJDn84Y1MlKN5QqaClHWp
QQiuveqLUCV9SgRJkKM+Kwd8bBMD5ZBho5hbqoyT2xK+joLNqIwKxezlkn11aTMLTNk8EY3o1rC5
5TNsemSPu3zOd5Jw2vBKVDB7uIiQYvaJjJ8tYcWryc2uDY9uca4pG42WKlWSQuCc9/M33Fmli4yY
0bYkhUApjjbHdy3wySClGqb8XSCJBDh5JNFuEk/hCfLxEwAkKOGT8zvv5u7brZifeRoI95Lzp1ak
NWP7nsPRw4alvwJ0sIhS6dCYm7ft4gmwyeuKzJgvaEIp/Ja9n7YG3Sm9b6JDohG1+2jiitpJc6hS
lKLeurFHFGKm2x6mMAzxTfvNAv8vHQSuhvRT2jozbek0COiqI1CcXxcwJqyZxTMKR+OUiS3loYUK
qEryMUMagU7DrZTEv9gNrvQZUk1zzBnplzq7XVv4RcORdwUWyPHWWDXComhGJExGPmw5afUFU2Hk
MyGBYIeWRziX+UVIPPzE+QnXIX3/m3Ww9EKvn2YJuOeimRBliFbGjybZYp5sZvyqk8oJh/k/xtvz
UQvGNvP/HmnfpcOqe2n7sI5Wo/jYSHyz8a2E0mOFVYFBmpN2IS77eRFvftnEAZBY83GiQHcP/NQQ
Roj22gDdbf06J/eIPmb3gY3UbddMF5Q9jN4p7Xxe+HqCY5ZVCF8yPaVRY3tJ4l+nAdlwkPZQrRDc
ncuBBlDTs/CUbCxNTGRnW4AqH2iGyz/Fk50fgNZq8G4y14ccAHM/cFFld92XuzuiNOVkvjgTOH/C
OwTPqSInRoO9sLCkQsAC3jQZGolP/RSBvEUp+von9j6QGDaHzJPDipK1GlIlSyp3sPOWc0lYkEVt
i8jN9i3UTdYkeNwPYKjoeK0Uk88zQNBdO8VZSoRoPZfpI2DaN7boI5geexu8VW0cvDEDJCBBhFoz
cxobOvK6tUb64rcx9w58/VemUXuppJu69Ix+0E7JY8OlIfItoZzFeAe2yCdtQPoLe7eEf1V1LnjJ
STHIfBBO5+SzFNFnQPFpgaele3ASAFghPGejBJi0478lVwPNBtc5ftG+g2KIJtYnGusVClOO4bLq
aUln2tp8r7pO1SzoyiKSfaxNeH5ZfCoDooMzzPPs54mLaqBIf/Pqv6sCGyAN6dZgsEwRDzEijCOu
yVmgasI1uswpdXsxJ4DVhytg9WaUV9muJXLtqZirt7lac+nAlya03mF4EaBnsOkQ/2Wsh0vhMoiH
PYj1SBlEIw572vk9c/YxLhrH+cnbt+z/mDgQ89PsOPm3yLzXuwI+8Sjtnxz/Ea1IXS4VbDFuNwy+
BfwCO8c6MXozIeNuOdr1Ip7ombo2seZVn0CylXajZyCnBK/abXPUPe/R6QDMPzacIDErvsRLspVv
K9WtcUQzRGzr6aIYTKFUVcpQSQBO7IFhcTmq53kVgAqysc3vh4P+/6aQNFFbotpuOBe4o+jlOMuF
9+x7wyZNtGNaGt9GMkPnHrVcZrZYUQc+3o9GuW4P/amFzP7cdz1tjUmSWh0FHjO+v5IHkaclV9by
Loge6iAFaziXumEdShleHHhrL5h48RYf68m7cT889tb+3Sl8T6Osi3ADER7udOJuhs4zLsvIJKHC
Cgy+xztLSTiUKn6s+ZQeKw5L4giRgyJ8R+jcvU5iWWoEVSxC+ns5J3ogCmjDdsb/m66aXLPm9RqH
xGUZkdr64Z871jaE6IobnGWH+sFtzqMGmrQrhzI6L5pSF9LyK0rAJKT14EouElLw36yqFNpk5IZE
f2K4RjSFqf3FJpvtE08rnIaVrszMTneaip3n2nqqLzPlIaGDsPVZ2h+H13nlqU8fuyKjq2Z9xKLP
o6fTXUkoE8PHNUyRPd79JJyx805ScOmcnUEHAxFIMGxIzSbpB8Jr7mFFg/e9RE2xkPXuzKylmoL9
n5VW3Df8O52m+b1g7SBlWCouvE9sl6wcV6R2GKvY8Ly36QISFZpu5FCMu9z/t8Dl5e0C7IYDvf/W
o8nMj6h09j8NmroHgEEs81vP5JPeySwh8lgnVvDVPWMimgUnX4V9CYXMYsmOD/IvrkWrs44DVPPn
sNzs8r3aJMe/dbHPwY4+jqwIEhw72M+V7SRUr7L3jPmmeZlSIq2r479dkUChsoqUa937xQuJz30f
BtaKx1NtsO2si1Zc4qEcVzcOIRO7lPsAT2yvyQftUklp4NSrFksZLaOd91o1y3pA7O/qKZYLEwKe
KWQjLMxrB5BXtn5rL1rPIBWmmmHCiPAwpsWudlyxQw7tcD382xqcMBFI60WsFv/D/JSnGd/D6OYu
UQyQA8KFAD+gHdESUzT9v0E0EhjfG5XCHsiqAgF4p+WjlfyfAl0Ha0SE+esufWIR6BBLmfc5dXYf
NQAVWd6PbD//Iz0bnjv63uuXgXqBkC3zyPMCaY/BnFymm0ZTHPY6pc5HevbLfO9IpchKRqNojXUo
YIqRjcYK1KJsgNzJApMuucWhuDtZsWx7ftJvfGwN7TPRNM9AOtWmoHGJ00v8mff6aSkMcWSjpLSJ
Ea+cA5sBnTfaEgEc1IokoHBLnQLOHkJ7Qfy5g1HE0H9HE09Me9ADzHQqgLyt/4k5tsf5E1YP3Ox6
dVkMboNMl0hMDbUegllKBxhMiyj/g1CWh5Z+cN8tyRkafqxneVkqgapLe+zJDZkb9d3iD5rKwHHE
QWPIcV6neKr5ai6pfW8ki3vfNptRx2QoBUlKt/1FOdTGqWVzIbqivrzmaGclZGCt/ogk0SY7aNDH
/8e7GMefIeR3zVr/FPJy3/CyjeWcbmez3RNTSmOxFFZ1sG9x+9n/eSveCdNur4hZSjpcwAzllvCy
gwLkAcJGVXPGwTuM/agMKFvdRLvFpd9n0zWRfamABJ7MBQ5+TN57ZWGzDkDbXMHZM08E98xbrX73
hMjpaUywuc14GPudDjGzpU3f/b/cCeg35ssIMdRhhN9n9EycLEy/2gvQDd5Z4KrZuaaocttwwF+z
ixwovFLieL/skIkIAtaZ9cqRxnyfW/UCWuOXVrQCEM/QsVRv1u5RTpvwxjyzlk9LMsofuQmB9mfD
lPH446QRhD9HgdKXWUzbSTI+3o5PeOcIMELosI5kzEwAW4MveTcfzHt00b+tTELtP6panl0Tmydz
vuLu81cfOKcDkQ6FZyO0zvKS3/qFZbv00ICuHzikTBQd/aK9vkvf1MeTjgwt3GyK/bZA6p229IQv
47b0XMaXTl70mEJ+HGaEw7Mc60f7vxFyta0T8jbx1qqmmc/ATw73rj87VUF2vmEEgoGwCGAEJeoM
4ojmzqoJ8TCyhwHzv4n+arVXkfMXDa0BYV2CBHBuXmuZoaFdf9rn8hs17IfLFpg7DkOMLbLhTimN
vjfH0AKWgZQYaRmC7+om3J/w2lrcpIrg02p4ZYa5zSoVzteip0lS+eb9GbO8Nav1DvqZhGdMWr0j
bFDGekmEc/oASyoDukqrBq0Clbh9N9kgKe7WfWxBGmU85fpNk9IKfQ9bjhja6vKn5wCkXy8/nuBI
S53olnUNO9F3F57IV1Ay4pWHMeXVXZ/1UCK+nixYMi8RbKbKBWPKMSgcoNq+oYK0j+1f6wla55YC
bswwablErcr0JAd4BKtEuVvi6fwtJ+JILaB6NCUBNDrrxANUkA+u/gxzxQDpWeIoHVRtz7dlxBTX
LbaJy79mcwjZtlzjKsEY7NIcogqGVso2hVI1AhLOmsZEOo2dFQDsOX2hrAK0XCbZ4W062KbPQ6F1
1V50imBc1Mr1Qs5DwZOuZr07ofJWHNWvAZjlv2i/cwn/e3ZbN7ePcQVeJHvGAygkUYsW4MPYN14M
veE0Vuvw1UXzwhNYDLxF3cBSi/Z9V7cQnnXu8L32EtR/9IQNsvT7Xdy5B3vtgFuvvQaUw6DX5fhb
JQCRtUHh9UzbTHvftPq1ALCx1kwlXxYbEAZaXmKrfW11sj6L2S8lbfLX9aK21mHA/pi+6uzN10v4
FOHLKDRPMylEPFjTMbLvfWcj2eMHhrlgOn1LgPm6PixaAlTYL91IeyJAB2dvFt9uTUQ0dduWrkdw
ZPJf8OABupXEvw3sechKsibk3TzGJmxRnxttsDbctVhOSsPNNXEDih+V/uJ2IYwfSs17tQLfKjSn
MHpv8nyKBRsy2fV2EGyf979Wvg7L81IH3O4vImbjY13kQELFNbOvDP85qntNISXejXPaBHCwtHoG
XbvI305D9LhUOgAyh8NyX4D+fzpIzhbpD0wC5rWpzp0JSkGjy66Q+zv+bsjfqnaqH4a06X9jLVSL
WjO9sEXGDEYt6T5L7flacMTn3dux5PezVWWRPslIuZuJ+fzJFYmQUlxE0Znl7yAWmbjE6001oUlU
n02bkXzoMUEsJBFcNk1bfusWuDRQcsQIFBfUOpbN/yA0PnJIc6ypSURcga6SZnpwV0Tss+nLLdxL
N4NEzGlhbapoOdDgiGIJ6RL60ELAvmKZmdvtvGJbyPU9qBySpA+AX9egG3tbiTcpvF/ehZmztIqc
bQWt4ts1rB7gbi+/DvNcn1PSWXn3xbhp0MaufTnslJNHkYqv0szyJSlsHAJiq/10SWcNMKkNihej
fOSPNlWEBh4Bmu5+2bgfTwMxuPwSfZ4CEum4nXJB6JRF7FdJ84CzrNiD63+oa4mOt/m10rmFvnA+
hsC9zrnut6I9nVaLgE6PJg30aZHPOc+Xcw9Ug7ZONu6/NwezC7CqvLyQuYU3D3ybccrCYvQAJ/hT
vVsoIzjAWCXhOnaul+ooUSyahMINgZO1fnPR03ZALsOMua9bcu7Ere6M8vITVhf0sIme/nAhbKMr
G30v5OJmXmonV/UFZFQzLSqCmrCwhJyGweaREbz+4eOPRgpCVU5mSkxu/Tw5nmi/U6l4ckvJDyB5
7AQv/XELG1GurU/Cg0pe5DsjOcIOQrdLUtwz2tsrMDXkEbXOa40jAh/YMMNb+oJonArqLetA9RxI
MDoKBfO5DDpGiD+5VqBbQOins3VA5KXk0xq835bcAJnNorGz3daXuYi/A4cmSXjL2D+mDAFaB+BJ
imhYmy/Xa+9ARM35lWghelrskuTG8haokJcHAR6pVw9EdxwvhejJZEt2HH6wXjzFEJbf8yNfO3RG
iiazV/txSh0g2LmlVC3JTJZkRklgSRQjsgJNm/D8ISvUmoxCI3OVNfEy3V4AGJkrxqxnlPRScQ7u
iGl0mN7V10Nr+UnEjMTKnteXXvCdZVh9Smf2SFLm2bUiZroyVhgyE0RRHLv/z6AGOMEog/IR3TUG
hCiT/AOmfZfy8bevZO/KH1Z7NJVhlpVp2j3MWr+UvM+B3iCRqwwwlOWq6vMx8g1hvKKIaXts4Py/
vN57x5BVEmkxY7iv7FVHXbatY1etAyrJQWzWwTUVSWG/c8VnY3zYqXcofU3NkZohDz+7NWepkK8h
qZlis/HCHjgQlW/hoSWp+IPmYEAgFTqKvPTmiJFoM1/F9qPoOHZstKGeTaC2NIXdD1luFbTIp6uj
9KMWcdVlVIjqPuIh7UC8HHGSSp6gn57bVv8ZVFlwGRxVp0wVe7Fpz5GrhlAKpHT6vVe0Fo2nXXm8
scl/OdfzfCKDeWJk8PtW8V9GIvbjYVWrVFWn/0cqpSDuBtiYsXeYcjnJ+iw+6hGDGjwIe5/7GtJc
1D2qm+07KADwUF7AqHsdonw+/OO0ADeNBwP6sROHR5+a5YNEsxU1RLYI9e6zi/F8sp3Eldv6w8Or
LcpBWouXeqXrN6x73GlgsVGNhL+YmP205FVVhOU7ay2hQgzP5o86Y1k6iC4U0MBQkq5TTHgI783t
r934MQJAiqcF4GV1muSrWeK0aFcsMfOdd2XtMr7jYdKhi0KWk9R0svCkHK9vIN6Dvy5Co3gt2Nuy
BU4t5opKf+d0eK2KgBuDvyYWf8FxkGj5fPy7IguMrC/M+oupWr3aZA/Cnm27TFj9CT7Fch/n45if
bxXBdMglYp97gk02MkHIfLRlxWxxsir9D8Xibded2HyHs9zpc9Rm4lKe3mvkJelVAVKDXJMa5w6W
OgZzr50LdoAwcExdTYy1BXxZyzVLCClTE+LTKOJCO8kir5FL6CcRSxSOb6nRFcBe0nGFvdjvS05h
hBwLalhZBdbP4VlIQZsesDcSzeih6UZ+tElCVDrawcBbXbHPp+k34HtyO2ktIGKYTt15gwjT1wR/
1IRF36/Qs3Y1txXkT0wnrnQXeeSzZtz/s2cMXOXtSZ0983mVPMriWEKBnYFyVPeLUzWMORuSUBVV
cosFYOHGoVtvRfP6kUQR1dGveKVx3Vd8sjSjVHKQDUl8q9zAATsA27HbeeRec19jwomWF8at5DQY
ua4fp9QjvaYyiOIL2mkdWv3jCYZ02CMUjjN5UT4YkNXMasv1TGR6kqX4kxwaiLbVwEbiuhQ0WxT/
Mq+zO/RGmaBgmKA5m0sNgdoFHYMwVPzw1h76A2grg4Jf0mGW9P9tw9fXIPENgG7kZOP8HEZKOmN1
lKHXGvrLWH5iTdqvogOCUEo8Fh38HX1B5dgcwMcTVq2BIttMfKdQ5xNR2RY7DogYdsb50HGZV9SR
dUvxd38XBtoxrcVSk6dgErW0AzdQJjsqmRYD/Pk7cxd9tLKhQ8qvz/ZCdzO9AUrUMQ3V0vWsh8zo
PC6PoR25tSKogAeekQGqn3rQonDKK1sLdSU/KLScF5hEUE1r1/DaKUfnKVomS9Ili4iY08GdG6UP
7Pq0nkNlBDyN/W/Ku4ow+gg70xnvO/h0rQdWdIwlDN8EfRv3JkT6+gqlTxzn7byFDjMnKyV9/ln7
S7MTY1pjO0SAKGSlxwlNyGAMJuaC6dpfM9cdHEeUwDNTDpfUnopVuqzyRjHCV0zGwTWRywPv8uHu
wahUFLpYGaPhAWi+7TixiA+/N+10eVIvrLVJMbqd7PWh6YxGoFYf9VhejTZYm7Vhf4Ja4eDH8NNb
dqGQFKB39M3gysuW42dBjim0efpIKNa6ffsxhv5JmbiPHpWmPa0dHdZKkMDzcHwgFtkNQzBk8cUr
5cR2xsx7uIw71d4yZEKPcjNM37z1d0K0HsJ8m6FVr7nbfEhBubLkjSp2vkgOGqGLhk0RuiiZZVYK
WzNlPIxezSfLy3tZSEDIEGhPPa4B7LbD8ucON6PuHRMlNTxKj/Oakc4yXqLYtItvQZUavVsHrJVP
1sOaOo7p/AZdiu+Sbh4RBD+xlVbgwDb+bf0P1gkhSP8SrP45jCye3DMmyx8+MObCioSBZdXPq/ja
yhqr/pLZqIwsAxVgpybt7h2XGQlSDLozN1l3LPzbnbkDuVZlx/O2JpcHdOC7PsiF2OL3ywl/28OZ
Ue5AhSC7NWgCF+yaX0OW7aLfmcFDlqcXVWQCYOIgp6j3ruGfPOYZ6gt6dU1dkaZHC5abm0bm4szl
heFLqMh/1UqJ1+tM9GsF1exwCJlKmBsHfKJRHPD34HcW58BWY+27pP2SlOhSkmFlRrrm9Hzsh6i3
/dqPHw3mEJ+N+QgC24tRestpPwe7yxtE2zEIC7dTcQo4+mZwBMitX0J1cRRdOCo717AJ4xu0Z+p/
O9RYPOn6nCPD0medbMPwhXKWJCWxubKPEbMzVSMw/2AcV650hMk39gIkZmeLpaC1Fl3w3tZeDhMd
aKBGTmPob/tBR1LODOEZbsoa+Esll8r6FPMzBmvGfUvV68QCMSA+LU1tq7U6oW1gux6CpZpqb4FT
itFLbt/5V2UmPZoz58SQR0HEO6xe6wcdsLzEPf/zE7hs/IxRIpVeeTFnkeYfUoOBE03Q2DgngVwN
V+0KUOX6HT2jYg6q9CnsI6CGkkOPvYtRHOltR/lhiFakdpuIQPnlbHH2ImoPVBnpzfVRvrFhKfyk
J7OFO+aJ0ypwLM7sAhgmmzK+xvzfkSBEBnJJx1Vuu/6+eEMZYRXRTJ17JgTRDTpmAEF81n45AwV3
62FzlBMdRiHcRHkReESQNApQXFAISGO6llzQ2veK/J8U5RYtUwRuA/pDZq2pC7iBLmehXmbgcbUu
S78g+Jt8DjtTJO23G4u75pYqubkKLCOPFET2oR9yh18kPC1ojZ2QJhbl2caXpMgMh2DwNJnpm12Y
AX9zFcV+qugKIhrCNxbDilG4K/cAsN/k6AWUkHt+ybZNWWhRa5ExlXf+ospHqVIu8TkJH9tKf3gD
tQVV/AKAl23ifEPRm5GizJpKw95u19e3odEFNkneyegYlnINkLAs7E84hiX7H1S5krj2o9c/RII1
h5BqQyAwEcEK8c/ntbp2CTzwx6KsRQKjjPqTIwozMPAaeO8KBhuuI5SLjseaC2+TH02oBrFpgKXa
lS7zA4ecEaqKrBpkfUdfZqSDMcmOYToAj5qRbarCe06Wt2q/caokDA5/7Ry3zX8uxyD7zLx0XaJN
cE5nM4nzcOynfUzRWI6ruaceO+gVzA9g3B0D+ucmrz+gJL2My4iNX3ue9gyqxDrQkyP36v4k5D2H
fKyJK4+gihqDN19nrzy8V3AgMzMUHyraHm3mWwGt2e4RZxEsOFbuRumMZuClz47obRZvuLFOA4QX
Hs63nk94Wktb+qcuaHzB6eBhAwhhw9VTv2+JJMJH7dfnI/UoaVcvc7QUxeUc362joDDundPtAEoW
9OChn+rIGu6F1qCk82uv2axJoc9R4Hl3WEeAIWeTKNCVNxkQ8DDud8WIfG4Ov9YDK2eQnTN0+o9L
GMexwhjDQNxxxJRjzjirejp934d3rSYAj+ZJa024Au+skC+eIx4qP+H4+GTrSEGWNl9G975ZZp2J
wxaV1JkzZOwhNZ4NDqIqTdNi6GlWb/I4AelcP+njLb7SBLYkYzJEHcf535hAsdzp0gzctUnXtLFC
OyRr5jktP9M5MVboX4Je8Y2o806JF0QviNjrzDWnjWMqAemw1U1K5R4ZAf4L/1dV12XbVLCO4YgI
bwMAWhmBXdq9d/GLzekQEpnZZb/3SOdrGsJg0YGHo0G5Ld2myiG2BJklhW3+Eg1lE0++FbUJBo7k
qQp9HppAzYUQl3CoBWv6ERTq/WXrpW+WDDKCWbbJRaDEmU7nZpsbbAJRKYohFoiudgzH/vqbcXIF
5pXqVEFjXDjfjp8z/qCRue5i9IIkFN0moFb8a3MlInLU9FSrOemRg+sJphBkVIQMfE7IHwVy0Se4
qczBdEVhnvLI1EM6/cVwQBrJ7h59QFbQ7IKguc6SJ/X0PIHCypGgr+4iXIr4jkZl7d4VKMqsIWmI
nGG212C7H/hm0j8G0Q4/kWaTG5GAAHTp5i0VXuE9Ryj06+zf3rug8KhMqo/B8uQ5jZU6Z+U4xa1v
NC9tJPajgq7tU9MYirPWB7maKEM7xZVLMLhaNpSSrlQs3L/t4a+iGHPS6tg1oWokRlgHv9iBdWXX
NJg7lf0FiYEN3Ost4tknhOy0lPp5m+ZY98yr6teNgqcLyvSongoQB3eraM5xIcSWw+2wbGHwTy03
hu7qdZMPh2VE2PtTBwvD45gjhEEZMrwNxWIhRrujlICAiwwBzPgSev3h83hg408npjBlJGymL1mH
SK2BsDEd+ScIKJ6WFX9skdNcSESqX+V3Yms9wwv5EPy2Riyvec4qiWxhaeCtFXHwbX8SYjwtriwO
RcvTQWpXcTjVE7bT3gFJFCmjZPzL1PIibHpMX552Vj21pVy1FoGTGp7sfoQAZwX5065Sb/FL4iE0
diPabXo177ADM0eKpVBiDq7qsAd50Y8VD+zpMsjtc0dx27u99BV6s5gQ8NVOWOri4xanAI3XOGHx
LIlB2e+Do8LAwsZ2sXsD5T4PNMzplZbWBK2mKeQ+lFdOl7/c0TQJUpo2/HmLFN2o0wfbf24HC5vO
SYtSKOtepa2c5IKM28MMvEcqR5kfybCoOv/r/IT6Q1fwyZTDH6Xq93+SoKOiwP5zUVljKTR3QB/x
B6Ys5pLHisRB1Z7OSeFK48DXJ1TDIENMmx/zc8y+ZXKM5rUMt1Jlzipr4jTGH53HrihK9KYXMraE
nBq0XjA+gVLij61Xl6TAgxOMQtTpAepb16S9Xsj5JNtNNsQ2ecdV4agE56/IBHDDDVa6uACsiSa6
dz4HBpb2bbqanhsZVLviqUzPoOhT55ixYREaUiAdBMP2ANvCRInwsvuRmPpnf1pmSL0t6lMoHFp0
71Rq+JvWWslCRsjyeVKNJh93JZFfUM3dpQ48pqpQkwWGk7kLpBo4/AO5aNOzYmJMHVIYm0jB5659
bJOvkRNlEeJSjL2D2x2am/EeruaYEWAppL+1aMqqyIquE6hEA7da1aCQ6lJ83DMWPEf/X3rU/A7O
XCnQ4v8Is5a54YZXvkOUj3spDcdGIz0AezdSVha1DqL/fQZpUhAWXwLIS9OxjgXnBeYdCcQ2pu5Z
1a6rePUAXPPF3y/dx/eBRHbfIaqWFfZDX9NcxhYgAqnBAjf0xkh76nn+zC6PxesaPP/KETBIxKRe
+Kai+xbg0ue3aMPjTOpPvUtz6n58Y9Vuxw2Uj2+il6m1YWQr+xS06NRlYYe75A4V6fDsgE5HExIV
72qvY4yo4Pu4esQ1KunAGJnzGy/6NIvVba3HN8KqNftuNxpVJxdhC+OKNUBZ8lJKzUb/99+MQwko
+WwiYZ83hZj8pcCqHPtTqIrJGvUrhuIZlA267CCCRbvk4m9b8X2+A05UNyyMqfSE1xu0aCzdcms/
o0Wx31rf56bKXv8kCLpEPTEGQRUN/wmqxEpVIBEIexS0YJ0AfMatF/sPv1lgey6SJ6n8KtkuObNT
RJXM5RStEYEwyTQpuL8Z8CxcKSgFKOFZzkAA4xkzeSzP76xMH0G73ornTUHixx0uD3d+BAlyMlea
IExeaXD9f/+dJ+FWO3q0E9VtlFW8RfAYXCz5nBFOs1WOsXrDbf15zMzjnHABdw3ijo6i09zkBY29
kVc6Krd+D9TowYDLHBLfPYbdIhDnwYOSJVKTLW35h6Wk6TXJ+qTE/PG+Xy272ECa9dsoeZ991Tq5
HPKFVnpxGxgxipLdCO0Yqw4hSM68DwGL28BpwxnIDB1senwKDhRyS5zN868Bq7nM9KUWo7HlR0Nj
J2taheVwOkioma3aZt+Aq/aZ6BhsAvZtsCVGLfFoYscNKzKYVhhLKyHywX5QzaYUhSLXfMhfe59E
KYMPJiiVX0yqYnYARsXnIY1ADYwE7jA3w0tnzOI71oI/c0RnhEEaa9WfEB/s+EZItu1X/KcHKXyZ
7NVHimGLPMgh1q3gVy9/DT3FpFrsy3O35QETNFCI3L1TxqXJYGLiiW8G8jf7Fw2gZourtV1IvAln
C8Qsr5eLAJ1VVVGpD3akMlMf4s6d57W7nVclIqsm18v58UFLhjCIVH6vSXW2pqgDQTRGvXyQ3ins
RkBeraZ0mLLbAArGCQ/V86ZQhslCJP9+Rp/E3I6kKIhburSL99HdQv38ILEslbirgQE/PtDi6S6Y
12c4aKcnt+vgdiKFFALTsGaw+Kaeu+jjdYilZpFfbP3oqzax3tdC8/x0by0cEjuvSjhefkDGI+IB
rpCY/nUN6jzmpEaLa/+Sl9WwKk0ODZc/XNa3oqevAmF58B30FPshDUfiRkLvgI7k6zK5UiFJ/SOV
NV+MjZrN6/zU9LSgtQVvqZHoMdFP+PiHbKwPiG2b4Wt0w3dbSZyW4HUDN+ZHDzx3Lvs6C50PmOvS
1GXG53vhBXAKhStwN/riYD45eWk/BVUk/m9+D6ETU1WuQDLZa60zHElGtMgRHLJ0FfFIZOoe1aZR
BTYMRFXGFZ5nZ/KNHs1rl2BDi0Q9QDad0thlLZft5Y8lhKcUHCPgn4lNuX2KPio1ZcxJsQYBCEzy
9u2Nss20C3MejOFEfsMBOF0I9qR9kRzhjkLL9jZF4pnM0gDDP34zOauajR95UHL0RBRTb7PtzdXq
eWcqifygIX6owWbDOoMCeVpUA28lBrJNmtB2JLJqwLuU/iCMPYRqbc8JVrGALJMYHR84a9C6eo2l
mOZ9+hf5PPYf9mMQU3UgID1MohG4X+A8byZQZJKxmNiII1X4mQ9E+Fbu1lR+qbcebDjvT1vCYiod
aIoVW1tJc9qBar3A1A5Nb8z1ugYT1N83DDNR9DJJard+zENgSHmCO4ZNX5/dIe64EU3H+mSfRPh3
WZSktIKzlAH9b8LOjjR62EGthqL0ewf5zSsdOkDsSUbPAhcS+8JIcBBeu/cZYEZa1sBbaiYrdROo
KmXlC0hhDJaiDeRE+FqQHuItklkN3GFz97UOPAPq6Y9CfjqRsuTj3IvByTqo/zA1ZWlA/3UvnZTh
nrt0JbPZaCY3iwn5vo5CxVTdc7GIh9Se24BiQTWyRhmZwd6SoHnRJRxVNFhCJl4SP/IXHcws7/E/
mtBrt7zjZm66crMUghHzrI1/bI5UkR6ZQOOIKBILGe+DrxFnHXLN5jpRCiyJy+fa54KtkQ4FUz2p
LUfkarFo7jRgf8O2giTLjXH3vkDxIpWJ90Fdqx/MKHoHTPccd0v4D+SOL3zU4QMpDQDI6uzbx7fb
aG152jctqXP0o6Od9pwCZ14NE6PQ5Ic3zDsfKntrz7nfBI8QeFwqaAK0Z0N502j/CID35hgIeKFe
HZoQIVXxL8tVzbq2TwaBLF4r49xlucdGRI2Yleb2s/wr5t5S5juKOOWNIXlZUE4HkfyA6jDuclTg
+U6CR2glI3MNaAM2moAeN/kFBYaXoSJYZsE/gbL+kknpTsXrlG70JMYnQgoTxm96ZvKy4KOSIpng
QWBw3J6ozZvon4vJOaTdKVJrh68l8LCSPJzWfEeJuZBGcch2XxTBlfHBO0KkU0iDMXtLAUTprkuf
0SQEG0NbbIGAc0cbjaQRoQNpfxWfNjNIzaDvYrB6QEG8QI26yrM2nnPet3YbOuRrIrI4wiD2TIsm
GW/26zPkwxIsO4dy8Gt05TDBis+U9VPFxlkf0y/76QW9cEl6Sl2OUPvpj7tZiCb5rwfEX2mzqg2D
ttraVW2faWh40hCDoilUf+rgZxKD3Tud63H4CLpvLY7jVQGiKWkwnN/zyzW/r/jf4p9yUOo6FlRN
HM0435CT2R3pk4tBWXvQkkiDsBQ7im/A1YdJppCAARsktaSK/lhzxDSIrtKmd94fQFVSOhzUDk9B
E0FFelVXP25f5kA1nzeYq3R+/uTwSQwVdiLUMjn/BMrhk0DA+wLi0jS2ueEQrmVJKOdzj03xvxYJ
yAmREc9aBGRzxGY6GNy5YyQhNwIIlE4Mk4k0qFnMoBzgNg81o4Eh8j67swm50pggoSsLei1PpuMS
vAhG9s0Ct5jewBx5iQYdc9wmjer35sGB0QhyqG6CvAN1l7esAnupwcLfftx2hfMkbHw+7jgO4ZNA
VyCCBpgNqNL7z2U5sPJixtyTRE2kzE9PZWwnzpufmd162guhWuSrIyOmIaWNc3Mcun3L6Qy4CxKC
rnfAPuklK1SESIwCqIdH/ln4gG3U/YVDKPvZgRDdQU81sPV6wYrZeCutiw+T39mdfzIqfrbpyt1J
3e5YZp7BLTcsqil8rLj7FrITxOlQHD0aH5YwBoSf2wFB3GVAMs9H0rO/Ql7tb7NwJVpbwLElEk7s
05QLlzx3lZdCb6sgnOwglKo1ZjrbXct8+Nbg1qdj1TRqDrC4zMps42X8hpZwhaw4xYYYrDH2fvOo
h2wgCpjNt3eVpfrbEtidWLzOGAhj8CTbdLoWm0CAt7PZ4hCE+aKU6ZOvvUBuly/IUl45XX4WvtEH
1YvJ1beQIKmc7UOjN60JXgUkd5pk8M7eLbQfcqEy/hETI/3nyTqzpfrcCcAURYVsqpAllYKjAOUS
gbAVQ0OKQdzJHCrHWh2F5tOk9pO1FytFTyLFdanySwp9E/W8UtWrLK5SB71tkEXvWHd0/Mqk3ZKm
+A+q+0N/uX+ECdybvGVhz4y+Zl6FT3zTpfLOs5xK2CmiJcun5rIpwaqy/MALlADb369uN3IHD1Jm
q8MJuqHa0dhpqPDPi/INxtMX2oS79ebOpieB3jjjbUSwKT8eXn+Q+K7zzYcrf+jIY0hSJx7reBfo
Bwo1WVDyAxr9ez16gwqIZsrJq8zSZefw/ygN1HAKLJhbYLe9Q4Wey68cldQ7VxG9pz1017rNc2vo
8cqqG0Q3SHQJqOpEd4AFTl1OfYWDJJy5B+XMQFUGhIQ4A3HaU8pMQw7Z2iu1RaD1WdbOGxe1FkPH
f7nEsrsOdf5aM/I5eMwyc6H7uBTEqMRk0Nj5VJqIAjUb2Y5GSCQlF/+8YzPx6B4dt1qLMZSAcjZp
e6dm2FGdsY5WnBD0+fCwcIelz2vC35fY+g4YVDIrq6nLIhtYM7SlI/EL35gM2dHYoaqx4SMEQI4H
PupDl8MRKngjcFQ2x1XkRgTdxUYQWVY8ohhjIzdf75hWQcJbFHFFNm95hghWMxmhrSvDz5WUH2/i
29eWU7X5IKJ05TiqOzOn7V5Bn0F+7Um+AUnF1WYLf9kz7MyqoX583roBT5eieuUmUF32KCr7BUhy
Dj87sCDPgTk2jx7Kg1oLtLrreD9VQ8g+p1tk9bs8IjSQqyOBxOHO8Byyjdog2gDbCsuWG2emXO3P
SVn27EAWtIzru5e64Kl4/vRogl1U4YpngUOYqEfmg9oke3BuLbjRIt7twuRislXZbvWnESee+tvI
k0V4waF4NlFmVRQo4mOm3bagW9Kcz4y7TgX5oF7YlDHYgUIWUnJh2CI9800TijFukdeCbVgJtq7n
lbIDY/Qvf9ffYxOkoloCa2VTlruXNasCVfJt2e68c3LoEwYrm5ripuzH1ZEVtmAiKbq21bLazWUZ
KxKukGbSfBbjIJ13xwt30D+qqkKFa8r9inlNgFo+gGu27fJvD36fcwifpyVcdihPoF4aoL1dwEMK
bXjJj+MzHVCjf8JZ7QyVcD5aCMHwwGt+vGfdF4EJ3zm1E26DauJ/2sCAGnPAbS53EyHXrOSKupWW
Xkggaqy7dQpvoVxtv/X+u8iLq4yEPoUtT+zXpCgumcgTfIROnmsLfxeCHwmRacwE/Suot8mcWCDi
T7cnnfXaWKFNkYrWQj2SbMEGOdtod5DEp7mCgHc65f+ikdBIa5T5PJ9JYj5taeYKRAbV7GTXu8eF
ix8OKzW+mZJLOf3+iIIsFDkewcwpqVbLi94iv1UC/f6NjMncdNixVagLYiUPH1JbpIUElm0DkB2i
LP1NFENLOV66WoABKMnM87PH4y+aGsjSwiJZrQqTDwwvutqOoNRJGBg1RYSrrLSz+7oiW5t9EkZ+
IaGwQfaXtN7p6TdXLXRxDDnS+gP3K6FQJk90JuwVuD5FFXUtr5ba++IHta/NkM+vrpG9L6Y/5bXa
w8454q/IHzjzfHVOoFsaiP+fXuW/9HGy4N2GxjSNTnIgizuOypVoaLJSyrKXO44cNJB8SxtPhiab
7B2iNGruY606FYYy+qdsf5VgnGw0I2YuxrjeNtvkzdUZ7XUPWvpNOyjA6Pn2yM37wTC/XKK/8lR5
lAJ/aYURh5kVzf1JSph8vWAKVLnwjFSO3BR9O+cpsfGW99p/4DvfklSU1E8HRB8Yeq8i0uy+VdRu
xgHfqVi5+w/UsF4gvDYgtj2xW9U3N0AvsSyjvoxryXB9lBqwc4lf28U0q2LNS4Wse+JeAnYr9fKg
2gm33XQbLE1vtw7L26FQt5HOMdN6oehlD/59XoK3GVh31YS7tZpQmc8JRgs8iSpROTkEjf+mM69A
uRNwHj05GVPoJW/Utp1qSjnM2ZWy3NbEzU7b7qwLNVcPITQIrYnCs5z1uYQYMbsnW+H7lDZ5q4Wf
ZaoWK4G0uV7gkNxFJiCX2UvAHMI5s4q5o8FHHpdaNxsEU7Xt7nldXzv0F3PtDURehCF6Qpq3O6jy
QH60oLmYLXGawFPBs0uV239E0Uqt7XPONq9BD3uDgWEsLnwKuFgNpvzbvM9RSa/Jvj0hs5OSSahU
MqUqzRBHN6YySQoKbVmmk94yYWfMh2pLel+DJd4u6yO3i87wE2FA08rqMpI/GUWrtoweUSWB6gy/
8PdVnRLpqQemYEIcidJUj1oMVzaeh0F5/8qhMuhEhZh2ZZjWeYDIvEMCieaJK12Q7VICNBlBC6S6
T+cxH1CQFDviONipwx5sblok64jY9D8Eo8+liZvRliCCiIEeEWfjm957hAM/iuTnteeiC+mArtTU
ut4CLeibraiMbWKgllAGgwNdWagnC7UmT4bhEUgq5Ed+UfWSmDhl2f0uQwbU5MwwqVGgbcXHHazE
Il6NK+9ae3JOWaclbHTmYmgvE6ejF6yNGRu002eS8mRDA7Ep6hQceRNjXa2T2U4APTzfpXhkwRYg
5gaZLsdRkon+53PMHKhUXWW5R7VbAsTY664ZcvAbC1oPxUYrcUtv/K4Jb/hkWNQI5wtRInixBmKt
b387Gsut7rdXm116850dzdVmO1n6IfPxUHA7YWbvugjaMIYH/oW47Da6eMq5dMjjakUfA9r3cdh2
lnBJiNqWTZakQNQtDoaXflSj+9a+ulAIUuD3qlqKMp3GWgHnJ60jMOYSygFUyiTYcvHskZd/A58j
IB7YimPzhMBLNSmjAhz7t/gMI6RCT1hE1TY+ME7KMchGuj+35C02U5Tib5cQOrCHDfRLF+Pdd1Li
uSA/1kTkz61MelPy7UrtZxoorFcKPOAAr2qz5gZ2XzqDgsRPlqe219s822Do5ZEEKygD+nN9shhJ
svsr3MoO4CJcsshqn7URocKzPoZehKuHFV16U7rrhTAgF95w3CNcgveEO/j6rrssklb0+GEHGHrL
5/6wQa9GZapokkZNEIDQheIbvH5VRXQ2bnYpOJ8GiKXvvPYixXXvjeYQZst8TuYt6n54uZ0XmpmF
qKYBz2E7TPFXwOkRuBUPp57wkDkqtgg3mNK+7f9sAGFE6mYi6Mx2goVKIBbDCdtAPVPeRMx83qzd
sH9HwWneC5U6ugppfPVI7q0k+w+PLU6oS+Tk12iNmzikiGBGPvIYRqq9pW5+N9MGxXwXJ9MTASnE
oKUJJ70gKAW2KD4YVhlk1JxWGm3onBQaSisLpYk+SNdYS8di4NVPbXs2Zam2jPIfnNuMqBZbrOzs
dklGczUhQ43AxwSYFDTmGgdV51r60u3/OM4oDrWhvME6PAyiAxoFsW/AmWtvoh2Hnhaj3TDU0k+G
Spylsf0QFdZCo6pQsyOT3/Q2pcWbqBruw9pq7HbHFcNRMoU+mCnv7aXqdKMXkO27rynupt1kNeBJ
ecsbthmRItyMVun/WUfNUuOeNFnoncVubojNRxIcMzP+0PwQSp4JXOxCD9RJ9pReNnivc4jGJ0nG
dGP7cUNIHmZ7CoRlhsbJ5HfUYvYQQUHVVewYNML0BLMq1qbTGX6K6UcIPxE1yTzS8ugfS+NZXEce
mR6ELfj2hb3gvm2dvmw34FEPsWMu6Rb3H4K+yxElshHuKW3/GtaKKwKkVnmajcPt0Bl1Rt+2Q+w/
oyrJaMkh33CfbdxfbiRQHxMScMM6mW5vlhZn7KnjqbKOAp+/WKruzRuHt1f6iwUJ6doqbWVGaelj
04LLpqfbb0YqMdOJeQ06IYg/fs5ZHBS7ktzPrgzFz02PSuOL7XIp8XOTI0mb9Qa7C/o4Q2uJ+I/m
f9V/7aG1Herl8E1l1WrkscaiIp6hf5hkT6YRtK75FTZBvkIXFkS/Zbbwnk7c1n03x+twTParPKAT
dMylTF2mR6zMIkP6tFiV7GIn+o4K2FveJWfYEwvBugpfK4MJmosi2CqLutA/VmHD+fMu9426JGkm
/xFmz4DhpYVGJckXPWKqik0KluXw0ypXHtGEZ+MPfGlzcrpojlpCEmrg5bkUczPEriW5iqvzoaWP
h8immcIwUGmeFl8lC/LBCV3c+V++TUdL+tsRb9SLJeTSbcORyyGMN84I9O8s2SoyhqBaoHgJaHDD
v1BlA7k8ldxSej8gpHKruK4sX8rgOwPXdWHRB89ZLV5ForHh76ReasbOg65+Gg5BsA7vmJHjNzSR
gWmm9DQj67izPiPDR2FWDaI+6bHSLNl7azPSZqXTIJAHOSqcpPXh1ytu3p6jIWLmO49wGjoVjXJT
MB5caZLM3YRWaT35jZ/WMq/u21ddbrCQkp/fj2SZ0nJTGolxS8CawUGPRG1OEXuGO4cpiVrVIuLO
w3MhHxsQCHr3Gw5cph9tWxmTlSAu+6PkhkAvV17Q+MByHYilJheu8M0XfGhvc4uh2BBPSmlezJaK
jgmvTB7ywgkOFnFDbum1M6u+4UDOT/kKq4WCMVRz2gnYLX8P6RRyWKv3bKU58Eh5QzmaZrakffZw
EZMTJP2oNuJ8ioKLeWKhf2S1SVAp3zZ0LHuWApBwyknn1SQT9r4zXdr1HflYgeph/xy4Hk4bI1WK
UzCivnxJe5g0QC9Y1zeCJLJSGtgrNQAw4XjhPEnbnVRh9Ca5xi7newKf81CDYiQw1wzGh7NH/Ra2
L4B0fvv26eJ5iVvZBHEXeDzPy7R79MG6kcgsHwyoW+2IT2uL9d6xBBkQdNh7cy1JNbIHysdurLPc
w/UU7f9lxU6CYyGkQKikDLZSD+P10jX9rcmJyPIyFDeyfO775ukJgb7TQfs9a+axzp1NsShoJFwy
0MQf50JsoxFKrOowZr2Codh0lmln0sjwAvrJGEAc/RpqJv6NNapIt0V/OhE90uT2CEBKA9J9QskJ
/+izv/QkLw4mbjcPmStKaMr9LzElw+i1JgwKjKJDgD+Kemd75xxD0nCxtHx7FicGo9sIX06Izxkm
1v96bZfX20uVQZuBPQSDjMOF4UTvHFz2DDvAS7fO2rHXghYj2Rx01jpBxU13R9L+IO1/ZJ/OCbS4
ZQNwdSvdGREpGdiQlbwFGgmyvY5+M5l/GqFv/nRzXGcC8gEEgjmE7fciBydbD3+UOg44gq/VfTvF
aYkuAXV2Zop4c87Umcdz54xYQ75VeCLUQwVLa1YJeHp1SfIAe1tIYKFJ1hH1OTUUa3g/nBcLN+5N
i+kC2oyiAV0GoXegn2RqmvCrnNKKI7Xj045pTHivrFbkZDtcr5hFFP1jY71FZ0zQ4LtqK0Ni4JOD
na4CIvU1CDHOdzcJdeU1yIHCieIRk4fLjaNXu/WRlIq4KhMFjHPqwfFGLLwcYv7vhtlU6b2mGPnJ
8wi/842F1+3cJaNCoz9Nd/9I8FPIBGFD5gEcsfuLTTjhFZ3TOM2OJM/8JjWSPvle06rhIM6i+tOc
bqE9PD1NaDWrIBExJVYte56PWS8l6zhbfZPlseRZlpE2ifb1fBXpfzZ8BIVWpKZN5iAySCb41pgP
n//Y2i6/juMOBNFO1NYtf3kVwzJTc5qoNic+pQQ9n0C+1ppuLW510ZEP6RfjXlRDZ4GKT5OvAsQh
WuZ+SAeaOQ2CsGykrgMHjDovjrygPTrQL20+8sBafJEJ9+cSwOwquSR5OnM3aUMyq+/PsRx2pr7W
NT47F1nduYBcmWA9APWefV6VyvID9a0qPk8FiwX+nQSNm/8n+DfZe58TOH4ADm4F21E80tl756MV
452cWWoeI9f72gQlSohJI/tJYZxoMC6UMsF0aftWm/kRCu1XojOMkhO5v8iBtMbxdR4P4ddy0X6a
wOWw0TJXbekvOIH1U8lOrerV/u77ZmY4VoChiPICRqLTYjeBcApRnpWMsJ4re36r5gzOXUXiByFw
CSq+Q64+HILMc2B/ddWKTvtjaZFOh0hNxMqDChNHJXluwLVVQYHL21xSEiaZjFBa1Fr9I/2hNfOU
5vtbS5nedn0T1dxunrGolxEs4MvcxleN/iFVDgIvkSq2xKfPHRPKbQP9ITXSSEpdhjTKfBQZ/KoH
xCf/+PVwuaQDXtcEak90GaiJ6plKpUlG4CNhh8AI5MpFlfyG4ZLBxRwYgUPSx1fPHrK99x9cZ/P+
b4bllakKg2LkqwaMyag35NccSUbwpb7wvXN6dfLiF5N+QyjAzH3RMQrJpH1+bX6QDloMcRMth8X0
z7qkDDxJiCdhR1sYAJygrtharygQd4/7VbqAZwLH7Rer+R5qe/+zoeECEZzdsOwUd10iX7HTRg51
GivoUs6Mg43N1+6qpe8qfJvxr5Zn5/fnPMCPrI2lvd6IN82fY/HjDmkXvlUq7R90ak6CfVTR6fR5
xPXswoRcPC8znNJb5V7eHAnfkHG+vla/DFx+K5G5rJJC4NIFWV51ZA1I9MJO6AdEGUnzhMNE0z6f
Pf7cnfEGE3pbgjgqur87QHqUbhsJH6/bH656gVcM+dPQ+NRDfKpJ86VCZ97hoBkb1VV+fnbL7ad6
YzIfQTmEVrXUWhSGjeUKX7XGFW/d1/n3O/Rv8PjP5LWhh/sPwXnm4f2U6LXH1qFVrbyWaSYtQsFO
KRjARIVE/H6bd2MSd3Kl5xrm9PM1taRnur2n9osreFQrXmybp+jFImaMDwpRzNqojpzldpWcuhGp
pDbxuBsJXBHKvzt9J/2wdLq3sxSFkFrh3rrbmgnBALiRMAhYKL1412WpUw5cHHuPxdiUKS3FVFh9
l18WJS8H2o0r/xGbaES763r5IzadKdT97rb9L6blbgF4hCpGScBGz0yNqDo3aSMeESVGDq5d3BOH
VRvCfIv6zRUOPG+zUm6UlFvmwcm9tfI7Hmm1UttGJujLXh6J76Jiff98dAWARG4rRJLVRiyppay7
xHiCitAIpmf3giiKgdHNpfKtKNfbb8Nqlrj4nHaCdzD5tYHA5Ok4R1brsoXiKb1VUT85s1hkQbwP
ae8vEeoumw97Orjh3xxSXtm/qI39axmBXsUi2DlzNBKPlgYAJg5OFIfRV2B+ntSc5uB8bFbmm4Kk
zmqJZh1JV1noFB7tGb2wDBlSQmYw7s9JecntxJQakKcQryM6N9mRxyt3bS5uaajnYg017csfkus2
JuNysu49638ELXBcd4mHVi4TTw1rVISwKCmoA4xAAmfO0fcAzkyWAQUubOQsZNs5S2xS4jf8xOa7
GdRgJ0kPvWlzGz77aLNBuoL5z9HFU/xPlIxETcYQJcHglduIbvFURQocY+PfIWvuWFT5uL5nMrDr
9jo55W3RC2mp8QTDZEzk22wFOs+EqSRoXyETNjEhLC9uw0vFzdfeLhHRjbfokP9VE+BisOVmYDuz
36fI56JdbjBf51GSz7SY7SVNavaIQUNu5Bo8Wu2CRiNIuK5fOeUpckU2+xxIZh4hhaNLMuSyrOSc
TgPSPPjqzSRyVruAoJFnyA17rz4A+0qr4DeVHs2TTO86lK3dubyodzWgDiJQ1cnBDPv72d4rbWng
ohRDrOCCzyxwUDOi2D2FwV9rf8jrJulfSapRB0bQwaZONgnO1rvPOwz+OaYJ2aC4UpPy8mlVLlBK
wUxT8c9YHJhognobjYSzfA7Pcz/t5PP7CzJ6T1pERrrdg+7ItMoKf0a8TrXQ1UEBXSlHfkQDu5EK
8LTKaSv6fLV5gjXdHinA/tsMpZHkbxOFUVk7WMw8plLEMeh+3J83S64Z5b3zdSXLdeak9KVKtjH2
7RQLZtC8G0JXBIYSio3JEzb/fQ6e165v+uAX79RMz35SjwerWy8vW65NtA2Pmj9+New5L/mgiMjF
SeW6M2vk/avxgH/GRI3EX/VcmRABcjI7OMQ/CVfOB7uC7F7vxVnCqZ/jDysn6MRY5ZUF+0HJiQ2x
IXHCObx7aiUI//b6Ac6w48sg04V44O79Ni2uYaXpYj6scNzMkrPnfbSlK9uYNwkZqBZ0Z9zpRv7P
bsplrrnxc23EhGtn8K/mPLXhZBr/JDHYFNSjxOGNuZxThYJvwHkDv1m7K5AKTDcLswVNB5IOFmsb
riC0QeOGnPZV2R5hCnuLTik9usZLaeWVgxMHQ/z/yo4+7P2YGuecRrCzX10re6jG1ojVloTPJemO
Oyd79hD4M6ruuRql+Rd5lp84xDcl0h+nhsEAxGASGe5OS7zDkoP7QD0GGj0M3+/r8fcqO4oWPvsO
FI/IQOhTQ6MDbwkbX6A7FBHNQNX7TRUjrUqsoqjwX0yvNUTROKlJxfoZoSIMpwzFVz5GkmHQk6dI
ozgQ6G6S8m6DYmL88yEeAly1zMq08QBvIxwZ24EGf74ZYzqBUBhp+is2cp/bdZ1CaXKY1lluNvNE
eu8/nLWx5IINxOmCu6rGVmYATTlXedlStw4oc0P3GbgVw6bPuER6ZuBzktZ/uLtti3GqMzNMClqF
mBl2/18PHbxhEC0qWblnehLwAdKpyIL+kt3EkaDge1xQwc7D2SIG+ssmQBM4uF4kkqVqKqpjqsXh
lawWJykOCMGauw+YQqgR2SKVP5iAuSGV+2kHAduT3hPY7JCCsXxAcx2/FGmskshOhxAvmCJC/JPW
O8KkunaD07CaEVyPqB5A43SLlpXAFQP4rSbvSTcWFSFX4J1nnrAzQoE7t4rIMqa/ylhGnxvVpvF2
fDkK1WO9GSlit5ZOduG981E09AsI9AKWxEJaLA4vARINUN9RcEKKFBwzqrd3re3O4RjWO6Mry800
l5L6efBo9PwsCYGT5hvwUwBJEA7vtx7oUk5OFr8LtDaq8DOueMrpW4qEVuNLPzy9LbM1ita9fTtr
mF+ch5kaskUoqEKN8yDqsxscpGy5DFhTOSuzD1IzFVH5uiLcBYeN4orErZMlCaqztxPeChGeWfEH
lmCRXpF3pfaGl7GrZdj+i6D2efbxfUISeGu7NKZIqPkeFYV06BM7QTAYmVg784DfIxjTeP9icw2U
/4YW3evfVpAWeZp65idIlIEtHCpTS4d0zHKy085AjRtH3FmzngfgwiX3z3h4R97dUO+uOJnolxAZ
SWcO1ADhvmj9fTFQljFaousxDzipLem0uQ97i7YjznDAESRJ+1L94cVciZf86sIxhQDggdcHT37n
YZ9/n06+j/OlsXZYTJA9Opm9rU5Mi4dliTclTnCTxmgtxRPbzcpmbBBO+EVYUv/+StyWnruMbRD/
4Ev+2s/bmTIX3rn17PH94YWu3rh9LxEC6A9cmGes3AkDhuEfcLEshvZIYh4ZmwaTqRzaUGKdbXOF
lJd+yKewRTRUcso5D556EBqsu5EWGz3GFH8NbFDj1z7NkibMCiItp0gY2QpMAlhEyVt8ayd7DvlO
XdCERD7EoABh1bZTehQnHifCiy5pF1RHtvoljklMH1VVAawWCJSvRxWDtSS376qZGggxb4ebA7nQ
skKUAjv9hjKmne3X4aEmQtrtJnaVe1ozQj5tBo261fO3zsdhcG9Ezpp+5Wqas+Ewzym7QOEp/ffS
Ad9uw61CyZepOpAVKr3LTnnJY50JGagTo6xa51sC1oQKCqise0YEYjevmMosHciiFsk6SnvmY15D
YOKz+A2eVKRgPfou1+ePOiOxYPdvkSH2uTbmMZrNqBLM+b0BUx4htGs5/OW4Czv01PhuiJ3is4AY
Ys7JsNYvq9iiKuEv+/XXX/PNY/8eRFYwNA9WZjjTu+IfoKaM/AGe5l1zRWl0KHMUN7E+JHF7L2k0
zHW3b0Bxnc8b4XfGi1j5SwKZOGPDNAbvOnV2AxIKqI4NanhXUgtSZctG0uQg7lZNArULpb7u45tE
ZEk+ABSc3GYdSlc5YY9FQ8zu361m9yKoAaIqRbgNixheg6wAWGGUrns3QS66talFf7pn9Gg5hvAq
2C33TpbeiujDjSZoJhJvFd8EyPnbp+Ci8TsGT5FyZAEgXWS8LzJSaB7d+t019GuRe1Z2K4MYC4kE
aVb/FocOIRjfaNmALWZDiLMT2cZB8T8COpR1OsP0Ey8nUr3hHp7XPc/HCSENP+CnXJ7JcHLvFAjE
AqEGu+Ri4l7HjHRRvcTsoT0WBQ677MgaQcuwR/9wIj/+0e49ip0459TtO/uWXxOhLEC96nYo/l/8
C4HRhy1DOi9oclOwezmEt+HWDP/BGonZKWE+j6z9JE7lGsIGIjhf2O+8D+tSjYQGdAfApjkInGAW
OZHSLictkyxgPlurldkhmIgU0OUaqxjBu95NKp+lIqxBlNuuNl+8VHEMTRa80WJciC7YKfyoe9kV
Xq/rNSM7KqL7QHNbCj1MPeTRrMNJ8EG4x+V0D9gUOf5+GQ7Rop3TVEsG8McMn5rvZA+P1Ssq0q8N
bxGXbTgKe+Ie1C0qH1QHXv2V0p8hJWg37kThuTxyazH1rDj+ySN6TVd2vtvhB5kkx2dPrmMKdSUJ
yXUgEAJ4ygbkMk+fOVyANjlNrQffZ+/S/bWYAQjQPEBbyPyRW4aTw8JKHkE4n+ubMuoJ3ht958q5
dt8q+YggGgTt72dK8P/dLeOl2r3iEQKZ/OC6fN+714qjKWxlLoeauXCi7lrE15nmwd0x0057BGyH
avIEacueR4zvXuPDISiHwMqwYYU+QDtNfsFnJ3JP51nglXLYh44YgtlhgSKeBUhu9FCERWnmu9DL
lBkMXTrSMcAYX01iYoTd7wcTCTpa0OGjzO7DQz2jg4qBZ/zmWJ+/IytFpA2rMs4letg86NNizL41
8msyFDWQo/TpQDEZw7p50CC/oIXRN47zA6eDFvEUr7n1t4n6M5PQ/tmhUEYBNtNA6G7MQLzmavwk
1t2/FR12J4OiW9P+l/WGpwoYZd3rUDhlasaYR5EKUyfoizQarhA3ss+1x+G493CmzKY4gUpjPH4r
Zt2GbzmhswlUhwyqkSR18iXovuuPsTM18ymT/sCTQoPeXFcW/bDf61Toni8mRbLd+ycyIo8ywVI0
LTQ5IDBTcKSBAiML2H3CP0XLLtMuLa8jrAL52gfAhEAHUi+EIQVfqjBxDL4jwQQxRfMvUpPT6R+9
LYWmHgshEPVIgcqCDl5tNn5Zy+TKZyz1acBLuivtrV5Z+ADLGW85gaCnlaszXjbSVTnnES/RLK7z
bzKbnxR+nC9Hf6BHyNrcqjDFbMr0Nn1czgbrOqDSknT4jQLAIbuzJtMVneILRf5nPTfaHn1iq/Tz
3j1yI2hGBCw5I+6tfaEOHVt54yK1jfHQJdALLm2SUdNSOYBRGm7kPkajWmyq9jU7OzYWTlcQ+lCD
nmiSuWO4sbje13DT8BukZV5J2cDjUoNwRMc068BBpqtRnOUG0zW6AVAlpUtpFMia+p+Jj8ttKhKf
E2jqcQJBwpPQIHlI+EjuOpwjtEo1quCrQBmS/UkPJJ7Jy7x2P5HWbSL/lv3Au+W3jxsEdYpU/AzM
g8xKUaxotYHKluoxtmMM8Zzll9pgkM2GXDXcatdXHTIS1uQTnoTirFd9zxNXu3iKo5tO49XmbvVy
C81sGoMmCY2DOK2Z7TaS11PcBeVPa5TzSxJ72Nt2hfM76ApHUXvzMsB3mckY3oWBPSoNUYqK9y8n
AYtmz2tzRO5XPsblg+dW98TBZN4SUt3aJn+c6Fvo7kZtnm7MG7f5rqCt9gDXFUEJaQNv2OiKGZ6h
ukpXhuM5WY/qEK3Uw25NNuOh71yBwVkziV/2UWAfB/5mTOlopTnMVYEycS3qGLxkr3n94a13yn57
iD7m1f0FTcaiHT2FgxuDA7Z7j+YtzRsk/y9NuGBcvH9pwGKrXAbOjVaw41HrarLTBdQRdkBwbaxY
PteMUJ76+fBHgjz6tK/N1Q9/C3SdcKSQoJwOhuCa1/CJWDnAIyVw1RbX9vmlMXkOrRBkRjm/tY1I
v3ZODmnxj3guSsI3KP4z3V+32SA1tD9jU4RkRNbdHloydOGTZ8ROoAF3tGhGC6dLlzMlD0+vEuCK
txx/ND++9rrrkI/LjDTquqHALymY2fmASb0A+FZLfuGehsOW5FrOIJTS0U3Kmsb+0rWPOY2G+9j9
D4zX0FiLs/9Um6IUmdBvclMn5NWmzXT4rJqT6T1oFmWFpSEBXAR1xAzjJLaHQUDRLWPuk/ddIDLm
p1vc0LD6rc0Br2xXFFEEb+eZ7T10BgJKuNM8FaWRfeRzaQh9kZxGtVlWvqzwuQqY6tkJi/3BN0ZO
BL8/y3xfWpTIY3iny1KBH/hYueVEhoRAYf4/0ed/p6J4jWTJHNSXbb2gK0vURBba4gfUDgI3YJHG
Cge2EglJO++Dmr5/421ASGARK2JJwkGqKoyDvpYo4M4e/niNry6SaeBAiM42ool4NyTMghBfJZIv
lIjJq9RKhGJ1tv3fjZTTxua1zSagJp3sv67Fhs/KqvQC3gjpEWOMMaNQrA2LaAI56L1fn6ertfSa
90+yYglJYUTIVzr+c3NzvsxxvrmTBzxkr3vCWCp+6MzYHj3tolLo1q20x1ub8KnRPrw77g7VJsgC
1K0Vx75WWU8c6iXY4C2rPTmJ4zFrX9LEVMZK7Oci8TgU02yeFJ46zCDhxANXS3KZ0VNS4XDuM8Ns
411X3W/lGvtQXR4NatfKn84JqicToxW75GEyoedwTUHrAvNFT1Z190O/DNHchwR4J2TvGFqKQN5m
6/BhVUgaSC91kaV1nfdSOIGgDmO+zL1YkUZBuopRidiFJyFE8MgkArEwoa0eKNWwD0d1sWq2yq27
76tSuxynv1c7R/JUDcWlri6qub2Q4+bHc2jCRP/lEP5Z+dO0NOH4rTUrcfVzJM+zE5smnIEU6dWH
7mEAQ18T6JGPzYmruOZfD5GBEb078OZkzu6UWeTabLpmq3jOkAJY7d99BcVjPQn1eTVaup3FBSLA
kJCbdc6Tecpf3ewhFg9r6FGCwg33GAzRyWEj+FS7L4YZ4Atul5x8QYtUFaBxKhwQVyN2SdKw6rly
WAm8CyPck4wWNGWdjwKQbmj6hlHrVftzkXnGsrXcqBs/wpLwR2otdpcrBOoDi170DVhFp2Pp9DHx
SXAl+uTVqqOe65aG+IImHY1IsCiNUf4RBtaKhj0tvg3mxu4g69X/TwafAq/Ucs1dVL5rkhIYiR0g
qwytnWa5raDraUzny7t700MET64CfqJvXfqwpy/aMCdGp80QcUnMt8yQu9UOhxCJhBPeicsTp3Cr
KkFlcEiBIbNYReAZmOoPIM8ksDf8xReCX9qKGpfYRxyUVmcNGBcq7zHQIyaiNGu84bJPfGJZw9rE
hV/xK9SW267Tk9k//azu6YzhISI7BRm27+2L3egEC3Sts/z5ZHkQGp7aYVTUv1b7omKQza+pGe6w
RBd14SSvPkvRCWP+ExUgyl2blAR98s1mFdjQ0Xtk5lg2nqUt5xQhiyrGYqhscpWPjGRHe1RSZIzV
/wUSSxfUAGU+Ik+6HImfuO0odsSJYHnGE1xqdh5RKa/2ZzoXxd5dpqbnBcrKcSeq+fqXOdLHyQYh
iVg/gYpyyjgKVnziFBclgDqLPifQQQNg3m141mjz1s4ZAsatNscT7wR3TLsf5QQV3dkYr9KR/FnM
q+PW9tkBLEOJXE1GO1wyapHQh4+b8xXOKeg3XAl4niYuirEZMR25vWnVbQxXDSkPJMqTMYweug6t
oJDQXjx02Qq7gGY5xKYRL4oanqH7KakkZFlB45yT7oijwG0HOGN1+2mqH6TM3emgb6Odc8JplAU6
ll1ZFzv9o7YgBNsb8R2duhY2Gklvsqe3NKT/qoqJUphz9glnfyi0SH5eC31i4+972Uaq9CqGArYq
t2QAydYaRudGzfMb/yHcpA3f5rz4G5YWtniuaNJh4rD0RIksm8az+jy9QkRoOpN3Ore8yMYeNwTy
HmQmcqu/Sh89HsVsUjazS/X8k46JJTeQEBp+VbD7meTX+0jksO9GMkGP+U8vifNNvssd+VJ4UPn+
YvG+9WWHIefZ/F2LjTgKTeYRkMGdiqYfmUSEG+XRMmVQIJW4IE7DXBOZmk+B71b/z1+SHjqV/7vc
lVojmg3RXJCmgD4qT/5lWGiIJ2N3LUJPgcUoFS51h7Axl4f+sFLwZ/N8NyIEYmmrPGcF/XpHIiZR
FC7ZtBnLU+EMLdkw0SLIqwqLqFI/J+ZLIdFqzQwA0Mg3R9EkyCPI/wVY/qhuw0kM773llyWMxqoM
cj9tbEgCz8adGR8CkHlab/++KgQ1PgQg5+rScOTAQF5itj5ufUZCLm7+m3c8ND6DcQIJJMKMYJ+z
pX+O4wy/ol1UFOj4VKXHp7M4QjSBhPfT/pqTqCs3BKkjLKpdQEsRVTHVW/sNbe/ESK7NdBJLduON
tP2l/nIBhLBkPIfUvi99o2yhZYou1m6iuY+LLpTpU1Wy5zx0r1B+kDoRkUKzQsUEW9T3ts185uZF
LZKgEZbNB4sUrd7O2wwfzHsI90+T3e/mC94GR9Ob125E2WplL4DASz131bKsHPDXpcI13aL17EqZ
xLduSUgFkSyKXa5bZjDidmHhTn1xKMAvaxZg6udNxJTlL42wHzFfRPTRrYThqUP637OtoFIG2h+Z
hYxxWzVPybVRkMzBE5KOvD/y8SPkF0efNX1Ui2OBQ+WqVAk5W4/cOcVwlSX1hICb9OhWHyLfa5Jv
sEOsQjRPFeQE591D+FeGQ4rLFDegZwOzZ1ORqyh3xp1nCScaNCd9EopI+cvgsRenwD+Cqqx1Aajf
w3ysk8sOmyP5xcY/y+Gb1FeTPZiImkB/ogeQdbEW0MrN/irgEkEmwbOhGPmTb/ghwMtKQJ7lJdWl
bxxEZj6xq5xU1GDofSG70Aagv3iy41/r4DuRQ525sPLrtZA563XSUyBwOPjUO5TbwZKADbgJchis
93owuEnxCVcZAvKwxcFV2ju1EtiC4+n+Hbyz4NyU2Qp5CEe41HH/RqPRv0I4hAztEXqVyBgCGolX
ySvfsl4NzFdJT2o4zXSS/Nm0nPwPPUt6RTEywpHWUe7xTBS+Gf4NG26uke6y0k4xByTcVLjTRvbz
V0Hx+o5OQQIE5+XzrWJ9Q0IOGZE8v/TR1pPHpx9piAEG2ApMx/1U3QXzN03G8Ao6B+nvcQNEMmQj
jUFKyxkWlooV4O1TN1L6MC+HRmtbERqH6aiRo1e4I3mcS2yxTDbV+R9sH1yUbP64qB7Vt4bbexNt
lTonl1TpBfpsyfaStPAp5VfLwXXjFa6OI3BhfeWA3IM3B7iOGSkJQZGeRHJaVgcxn+Tb+AF6OHox
wTIWHnBqi1q8+5Q2e5+vx4O+bpa5cDjEXiLpPZxxHO6XZk2/DvSpI8JFa0K2I+XODJZFqiC4/Tux
leXDJNiAfWnxCilvGj4pcMqkB5DtQCBdETCLQ3Zg0wBaX79R9phbZyp6NXJK91711enhNt6gOByf
6b0xf9CoHky/mSWQPBwjVtqXzfngYlujtsFJtXd6THzKiMv9agdq8RU7nG+06ehm0zGfH22bKaTB
Aa4uvI9lltC8WW6EnGeAEOheFxow27L84AcAYnnOZgH3tOt3gy2GldhmSe8v82XWfLDBl61C//ka
nTelj7jR1vEY4UqPQbvfU0jurm2WPwHQO/N10g/9Kx81c3g9rsB3py0e5B0ozzOlAf2WGeErRhx7
vIlwL35vao4oWz8glbbkDxyC/nUpJpE2GHj5wsx565PCVVp2c+dF1Bg+sqjoXwaodbC4v1nvz9h6
wI8iOt39F3WPHV/aHUaUZcK12tYlEKQpYDeTf5N68pAGVU+J2wXyI0BqqghcXlvyt4+q/ZcAeKvN
PaZCwiux5VZ6G+8AiXFON4+aWqHviNzotVkI7A1n5Jbimc55nvYVs9c+rbwthlCpGvLn7zEI8y2a
whS9d6jPf54VEjcuWhGqIK3i0/Hf05LqFkuq6ZLwyiZnmP//2Ev+H1igh6yCbUKVXwPbkL5y7fRz
XaYm3yohqw9c7lbHGES5kbOlqArULAwLeGB+38GHyYcqdWGdj4mvrpILRpEh7KHCP6uC8cW8HudI
NQoQ2074A1s/TQPyhpopklOwh6cRICI6q+/j5wOehLqaf2VHLG+jKKDAf1Z+1khYzwmOmV5ORwVI
YQOFRwkJRTes2P28h1oo7wnBRi5Ny353Lv9Wc06gDLQdxclfV/veRI4ZMubiAFFRYuEND6g5lIEi
guwbS7EjEuXCKAI85kGEDV7fSPH0taQjHJ3TELiES2/xbbzAI2nmI43Ig8nzunAwIHWHkuyOmgqW
KQCQZlpgZgitTQ8GSVovMWhFT0o7775TlhCfVTdWqFKV9QbQV/1+W07G0qkJ/PB7S1phmsAGXvgf
3EgBrtYSjj5L9g8mr5Sq7g7nwSIVjlJEBy7K1UU8nihJYbCw12Ab/WyYP4WL8K9+SkG3EjGgkIAD
uqu7+axEAYwz4lGDLF6xPPWQ255GeiUQtw1VSIwRkgiUbB4a/5IOuJskcqU3IwBTCrV7HeO9QMQ7
I/CwzCn6BI6JcJAQgEMvGgVvK00SItUufXB3MDO1S4h/8Sw8ypAjQ/XQ1K42o48aXqq2yZ7UrioL
zIgYop8Hx8rg3NxsMnlrdwRZJr8QiAqJoHkFHunvxOe+Gjy2gcN2YPxt4mrHNcyBA/0IAIh2zasX
BMKocs7WbbF5PLTT15j3l8cOFunxZK3UHw0FGdtzVpSTH3uRf2frFz8uVQjlIeNs0C84R9fFZbtF
Rrdopd4X3hOPoy5SVobj8TNnolyTcPNqMoOMIP/Dj5zVWUE0Bfq0eK/HXVrkRTZ0404vpqTVJCnS
WcZEckfu9MSP4LWuxapSmz3dGnn1y6HztDi5FNJ9ST2sItAldR73rkEZXnOOmCuqbn0Ty4xCJc1O
DTYIkCcERFt73HLPrqb10vuVTlxcIu0zlfWbSw2HvapFgNfyA5JihrldCfD+aOa8pHTQU4L+RNkw
7n/7LQRRqBvMcJf7GMmQPMrMK0fqxE3PW88Dynk9JrVWVoDbgP59zFYt75E8/5ccBE4jMZQEsfUz
ZvXi8EgCQHf4mYCu9rjNgfHkP3dJ5AtAs9ZqLZs2x7It5ZbPDARqhk/RhhXLDWxz27tLkSJljTKk
zQk5zqzU34orpng0F4+xXsgZOU3vPj9k4EGTGP8vy/2Yr0QIQE6wAXUiD0nzPEiKbCPv9MUMoH7p
dfMPVENtyE1fey07pYr4/13BRxYNIw4wMLY6coiW/iMo12amjhKfkuU79oTq56udf4FZZN8Mnkiu
7BkwvMZyWPTQen6LaeeDKqX++o5UqOC5OG2KSzLYcBZCGKx1cVKuM+hBohPHDcqpCpNLczlOo7BZ
QNGf4n/hjeLJUByS+iRO6kiqGvf4FxwyGn76yIVdt6ZB8c3cJJ3v5gudTx1A445gZvCiaJ96qhkq
TU2H+m4PLRg1ldIrfXKuyUsiNuMznjMpCnlm65nzjULQdHOf0qrL7+NLUW6VEq98ZcQmY6nloXeC
BErVw1tjEIMN/2RuANJd7k0qj/5uyF9yk4wcy4pdGPGnWqq0z0L3XXSrxzuDbMQesbvwP0ew+cd6
Xu29ILda5Nkx23+PZ/9N9GJsAxCylj6zs4+4yZKmxjtGdiMXLAmA+TB41jGmcN7GDWg61CFtFZNg
zv9lovtILsl1z0J2FrcVwcmBUBJbflbh7MUmSbrb3kmIClhZTgYrQv75Fux6q7dnESal8UAVMSWc
BltjIAgw9guDR3jZdE1OvKrSmN/bCCPETTXdP9GbE2ZxaUQDjjuOTZi8tghmMIKGSHPsOwYbJq4x
HQbN4LBs73nbw10hrhl/GEuz62p8b5D5ILflINVVJi1CHbYfb+w22g/phdnUhExgIlO5B0qVceJ4
YBUu8OECI0ltZEaCAJh+fTA/UeMxW1zHmfrr/WZDKt66uujG4ugGCiibQdUZ1bbjZQqcVsqstMhF
hllSvNep1huGJm4OJCKI+q4F5pRJMoV2P5/ZMeAj/er8vDSKo3zC+P98+R6MuERAtBLbG8sgjo/c
6mbwZkCy7yoncSGdz8C7bFXluYOZYs1tDDKXPo/tYRwsGbEX/6FYw9TdRfNviNr6NlPclLG3MnR6
M9G6Yg0Ys13jzN1VoXRc7wegGJ3fV6QR0weqQOO4zO7lJbfJpt3JtKoXPbkGdIgXwkX+kG1gKpVb
QcuKHmmFG/i0axGbQR9l7TvPU4AfGQTGQQQfsmVCmO2oXWUt/3Rgamk97qHHf49UHm98J/RVwYuu
9hCwj1hBuVwI7s/2PcP20f4DBFhYcdzixJ/+jS7FmeEZD6WQZZvMt6GvCvhSWwL367E5e3XQCl43
fHPe0kvByYzhqUoTm6A6w2XFbgVpm5m3ts6XPZ0Z7IWMpLH26AdAS0NTlIkvYC3iaZ3sF2dpDCN4
XEub8jAbODKEmu2VoPdeQGB/iNrrflpTckr+flPrUgkKr3fPpbh+wMq9hbvu/XyNRzUMzYnqBFYT
IFdJeq4/FQSko2lo+u5TqDzGNE9KU4eigASkzooIYt2X1lvnpx/LE0UfTP800GDf0+Bfa+VFfH91
vVVShGKBCiHWgjrT7pwASWKtoZuoA9D0SZOBwlwdyiWIViGCL2r/Os3oJdVzbvODj+r4TR4wYAsT
jMgw47uHqY/SQ6H4FOwMDKXkzKDmmzDAwdm05k9pUtBLXq1zy/+0e7597lhVxpnfx9DWyFntdGew
38tRvrBgEAU5oCWByhPVrTyiGp65tpY4CxSeDXJCW5uGL6N91VNx8O51RCSoIJihHx30IxWHKwzE
+kMoh+3T17Xo7Ac88Gp0gZi1c/+k2mPLAufy4mpyRx2+IEqd3G7hy6/2vdGxfG94mjORholLBx+t
ToHr+813Q/XOgq3WCrfr5vTXdzEL1qnbowVA3aNoNjoFH5GuL8qh8h1+JyBDc2iulrsFXUcqSXHq
PLbyXzqcitE+BUVbfpc+nyAO9bi6uuFswoMeP/ePYLNmIPgNYmGTqeL96g+sDQGZ2pZMRBnWOjH4
/asaGiNxwLw1+MTAkTyVpAbduDKSl5ftkBXbXkKGJH6eBhwieWVwGl2Ydp+XXMff5eQ9W4ynkjHn
F05Y8NPU5sy3LLOxr+OefqcSJtu6oSfoD/tu1GfkHz4ZB3hbnORavfmQo50fWr2qYR+GNhsqiZHq
tE3cf9K8dMJpOLP68fBJOnr8VOKjnWSVHlyFV2rKuLhoUV+/dNW+wsq4F0KSu2xDOq8rgPSIyXv5
L+6+V2VfXocFbqeFN/LRNKZuw+l5pNa+9AaHBhDlbYXqIwEaVGGoTknaxH6IIrgqn3OR4kPvP3mk
ViCaxP0SmKZczCZx2VFjyCcTwnqNG+K2T/4EOsiI8DOs17DD14VB7+oc9FvisKXdTVZ8ySTf51Nu
+IrrE5+hGXkl0q/jS6X3BtAvshLqB8Z07RiMAZWpGzgMLSeq10ZnmyCnrjQMhV5W9QvpmiTuskPb
X4sBbpwqUFpuSYHYZLZiYLOg82w+UuHyq/SKU0y3W01be3CZe7W8HLGeMrjlz6kj4MEp1vqILk3m
e+R01i6ScZ0fvL+gFIXgWomdFW+5U0KTpHgoTFFw4e93nSxNSxIqmbC1ElaHdJkcabUHsDmMJt8Z
kTctk9JzuUcvooZydgFnOGaBDK+tpB9u5g3HQxdZDcrc2o1hB9eFSyAF5J30Ezyn5hLnrrWZmcCu
0dCgzV5RBrpAQaFpC95kRECEVa4FhCpgcHncQn+kLdlAKLd8+TSlX+9PHVwqXRadqKVYR6/dUaWJ
+08mCqCULImpimMTLgtZ6nxelOgiLH6Mrmyn4LXqIyH2v/f1zs69bmoH3r4wVq5sKvzdVGCuttXm
1Ljtx7eT5Eq3c1835GxQCtyu+UcHzNZNGzfFeMDRkQuM8s9IyvMaYo9ATXw7uMHdA41g5N/fs3dy
w7cS8kxbpZXbz4VxkfdYWjJ8L171Cy4YfRWPtn1kZooYX5gNt54nSvW374YsosKVNwmyRxJf9QdK
AgXHt74P0ivn9Z5ee68ARa+zDOOG+cZWE3Yw4Rsjc84AK0OZW/WEQydYvrF2g4SqwyTb9oQmACIP
z9bLxLIR9YLhhrqU7P177U8HwMdtmstHze6ryE66xvJxjBLxoFZ8gT6Q/WLFoGWikxY/BGtihCId
ERYcuDUqEYVdmgSH8+0Ngx3Ni0DTzEALuQAcoXj3sfQXiSDMNXcqOULNT+Oxbn4LgpcZrVvYX+eE
dNMyxu3DVdQw/vCwr3ixmwACiS7sKyS0RdDRgu6ze5d0CCa1O7rwfC/9pmkbt2GIDZUUk5flg3fR
6dGSeHYAKcI5T9os9V1e7gCvWymVa/cG9gEKzsPPaj5tH+ExtxcjxgoDFpOLJ/cquTnc5GKehcC2
+/FJAF+9GFePAJfLr6dJ6cA4DW+Ekr2R9lwmmgOfnuXqKnoe6S3FNQKl8XJj6NJcmH5Z94wZ7DMi
xTAAS/a8Mya7kJioQW3H/6TYnyZpNBYWWt8VM7X4o/kn5ajU6F6UdXYR3ap3UvVeolkDHzbVSUBr
JmBd73oMKrmJNnwB9ZEp9OKwf5Ic1uo0WG4Mk/0A95m7RFCnctdTTKkcqGXmNF88N417fYrEm4fh
N+GZExcOMWQC5t03Mg7v+uuwKRtZkZgX+wHaSRNJcILnNuSikqod1yPySW/noWLIWToQfxq8+8ZD
kF08qQ324f1R5AW9Keldu2KVc31qFMwupI7pK6lOmdQVmB6ehfyPgEhxsepQqx1F8/w4rs6hfikm
hrwCKDO/JEGl526E/EmXYnZCyJBZrqDBBwm5NVmLIHuUprFaHq9u8Xp6k+n1ZNulblL59OJmHEsT
Yu2qZxIcApNbX3TM1xTaNFISAb0R4lpHTiH/whzlgQ1xoINGcBUaXPSDL1EUn5XqdG0upgtr6a7L
TP2jaMgw0HwBF+HZ5CkXiUdQApzBa6pYl7IBo2nHh5WZDxl2cmbjlIusrvgMjaemdc1ty4AjRmtD
sTQODRQPGtMwpQtXzTbxwB4HfmL96lklwgF/CSNo0+rbk+Z7OAx3OGtiJRsVgZKHkeFQO0qgTf6M
L1HwfUOZJDqyy9UtbzN7DOYjbPZh/y7HNfG25yN4OMSgp6sdsmX7eTnO0yLIwU3YiYhEZdl+zrl2
BnmjYJEh0YdqgK84izO0Gkz3gBlJAYUPUTDFL7Xi9kdRn1zleQynRu6ZlL9Nv+wx3j4MT8E4wkDp
DFjoC60F72tQrKN2xKbux3mSURXP5z+KbY2i+FvINMLrHHCW5zXrwGtGdbqVfTZdTzFOkr7ZjF+T
4Btu0sO9BD43TbZH5O4Km6fMWdfyHnnYrx8x3g6n8ma+a0PVY3qOW/JHgbaNk+0zTgiQZ5Dohvir
rnHAyFMXXGdUqyHR1KDQGShdONzTdaimwRRzcmyHU1YqfB1r06Xwp1CZ/jJAQbY2bO2bnJ4ntDVg
+iSufPMNwDEOmLDEhI9P/dKmZZF+PheTHj4l0YVXnZUlFwTgzTSq3nWGgtI8rUeXt82Ur8KYdvXW
qzvJ6QqL+tO8TqpmBVrpXn+PIcACuf11SQ4X79wKHz2di8d3SJdyVldAHVRxIk3EOqiPwmvIATic
0KTUkjBRcx964/+JpQbGcrVYXe7AIa9WzaJF7ltCHNRWENPpwyG7rcW3VnzfPRYpPsrfqiJmd/G9
U3/vUHHZiFxYmmR42J2cqOsn/ixw6L4rIYBWAhK/MxUh7ap+X1KGTUWFwipDioY4MXwuJ+GNlm90
C5H8Ea9uNrUPDFjwK/V6l7a3BhLpWDTlzBLMfWKl5cCdcvYuCs77hxVLu9QTjITSxa/WKb+wvl9+
2FVBhQoBhz/0XrrY2VyqSKZTW0y3lN75Vj0GxXcUSSUhjKwjzaNauYQBbluHwGGuctLX0wz7xE55
PXyMVDQ7RN5oiwv29cufAxyVbRj02kCNm6Plqa2QotDN54S7NGed2Glqm7+UZLoTn2m5eS50ZBLo
uoIJWB3fkj+6KyOOVU1YHoScOTTWpkJNbe5IZVXHAtcwKceJSuKlSzA8QVrhVfC3jFkktvzqcl2Q
Eb0mi1J6M2ubCLwUP269NS7J9wa5wCzy3ZPMU7EZrNDUPzHtFMFXL2CEbyGpw677lTeGU5rO9ZrJ
atl/pbrBwWnljllLNis7z8dVeYOAaIUD+jbQs4w2k1s9q6l32oY0lLKOelZnAAJ+JRpOeaG0SphY
00llluCaxXzHnwoindW3LszN97B5KeaiUBKnqx8S/alkbjmVSMdQaEPfedyx3zYpylWW0ZxKrN9V
S2UE/4LIhhNT6iaT87xgjWyeghjSkqK7PawxEIYaK542QJNtl9THuB6tRmFus0R1RW8rbfuQEvtp
XWGT75pALaIgD5x+l5DnpaElykunPFoBJQFJgiBvo87ykZjcsZvVuDwTh2Lx5jCYT3yyMUUspdTF
X8ewjXOftGrTLQY3brxjT60L2NOBFHaL6BlpS5kwvTH8yXoXnLrhfaaXNEO80WBfj6EYEYOxRaeu
qDY0XcH9iVJmvGbRuLiJWx5EFz0J/M5VGrOX/ZAZKYoByzvoqgn3NJQrpqYLzc54+ufCT5Vcr6Z3
SfevbjUaf7BSB0IgWVHCzUf37Za20maHhByiQYF6zTY5NAwcF9Xts6B7h7pE32rbT4cerSnUiA/g
uvt6ecyrumcQvbUy6huOb0QvE/qz/Ue5sVium+dj07aGJ0uAHRd0bmorIhrPvG1d3KfM2gtdMYbl
pWly1TZR+Q8/7fTatXvEJL9CNjBO25E20aoVs94erb493pW+I++fIhSyAM/Vg6QrL1p/GQT4ULE6
L6S1oTPp9xDPPWUKWE+QFKbgqmu2LhYuMhSqGL2AUK9iZGMyc3iU7vjbKfKzefG6okvVBWy3kqPc
TC6n3BF/o9WyBtY8z6ZELRoFhu2n81x3WvyWzRuobN6j6EV6jJo0rNO4D2xdmlAjToEqc9GOB1p8
45gY+2wi2QuILGzIuoVjFTjWeMFqh3zpJyq5+IOidK2dDwa7bXO7jRQzhjDou6/6ed/AdUDlmCFm
rbzaxgsHXEPnmKoQ6FhCu9qz+7F3bU7pxtnO4cD1RTG/kEzbvzXReOYThicRAW2n0DCiyOYPsZA3
ywDdDGLkGB/s0XwBD8iqdXjHHPe/aUUxrhMmzUIYD/s1eTKg2c7DXIRK5u8AVLSfLAiWEnslRn5W
l2K5+zLSQmE6gAFVgNINba60HAWpnvLmsLRGLwIbFGhkzTNbsSEo1phDrMCcQDjFJukOyIOJe3ql
WZiTWUvYkkjNSpHFSRIP5UpS4i3s37KVuVClZpIYYdMp6nSbgQytz1TfJG1kIvBy2N1+G7VcIGGG
mIEbTaT2IHbmKbi7DzwdMQGRFkB12mPuypOkYAjCEQkxmX5DQLrXvevnvB/AMvND9/vU8Yiod5mA
8/EEU/4CIeuIEVfTppn3IdgolzLSAcM0UFtz0GQc0YvQZf5K1GzIJqDxwhQwc/u8Ez8WJ73TT4mr
Da8DZhH+/ywgharfA+mJ5oA+IEfInKcM8iE7Kfi7N88vE3++/ex+wlDGfLOjS9V/NpcsO0QBdJ7g
caMBx9QZ3bPRSGijOKYUlPSj/89bs5Tg4bVkkQDWK3K4mR2rEMReJRo/InkpXP23IqnEoMqzMFK8
ze5ohDI4m8AJyvxwTZEH0cHC2ivQs6iu12PUljP8tlsIiyIge0K6DtHc45k/M+pR4+8OCz1rOVjZ
21PjcU3fi3Leylpbng1N5tt7g4Q5kZwaoIFmmQg1yT7JVKls7CK9pKMDyu4z4vxuIkUUl92OxxVo
VKSORzPAMs3n98MBi/RUuKkdtGmn235KlT9Jnh7DB9rI8cj7kdgkbtpWA/jtVsNz3oIGhdJD6j4/
hgrghSdNyRFFecJ81CedaNkNM8zg9OEkMIiqq/xoJB5R7Qcl2I/FI86B5Kp7eAEQmW4RUfJUDtcB
9+/VuM2e74f0+KZsDIku1taeb3IjkDv3wqe6RO6PpDiPYcJ5RDc0UvVv+PhYP5dfiZ7/eY67Fo/p
7MXb21K/mLAkaV0PpZPhD/TVh+YtdvIsHMmxxcsP9m8tq0y5hs87zzLkEnmjYIy6GKIvP9PKWmmN
C9Tu5wYK5IcqEfU5YmPmhq04mvIiuitFAhSf5AIZnpIMdo07OPudbXSDdnelXrgOpI35KTaWLYjW
lns7W+UvvgWWzvT8WrkPC6NnkbZf4OTcoiuBEluuj8e/jKp4oC7lMhCjiQ9Znzp9eCDTV3RGwEPl
d5+vRup8VkQ2+Y9ICfFkDT8Ph6oi5EbfaaNc+l3OXSxtYH3sLJ/PAxEEgEmN+JFWU0DknL9MRrvW
JxJacPz2BnZCUvBouO+MKiYRKd7mDaqSKv3yN3CSf3ACvqvwFeDcV/HSxtjNo57/JOYju+rJJmAW
8pGbFMig5YAWrNfEqH5WORAohGJKN4nxsnLCuc1LMP97i5igCdqq5MmO3QRkuwh+L5vMfwpjAUVe
z6+I+oYwJ5ZjZ2Eg1yV0QKDOSvm79lAZJo4w3pzipTo0GBka/Y+EmUv1CzMyvgdtkOryo7DMhSLr
yQcykePPkGYRlZHKUwVoC+9aR1nfzNFRZgYXTvwLH0lMKtgJg1Ygz1q17pEBX7qrWmU5UOlHJya6
O/U5DLBWean4v70tfqqtwZJAiRLJXZ34TfrBuAD/f3EhgXk04KNAJ3jMf8ine+1bxsoPNWpszht1
40qaKdXwc5RlIoFME8TnDqyDQsYCBQrGW7pe/svedu6ieMnaQwk7x1S0uWFxYWTsYuC2WbBPXeJt
Isp4NZOszzhvyNCh6ISIeu49ZCW4w3yuvdEf/9v8cp7fEuoTcvWP9P9+B8Y5298ViiIoDxSaJosj
vu8cYqgaZqu03Vzuj/PwCckQc7S15aQOZYP5tVwHZsXIPxLklG1zHNBq780+Mr5mE0dfeb/i8r7Y
StdRzEJ515IiDlADkj+MAPAEFQ3I0DEDyTRhLwrdwrAOBpb82IMmH/GSHXd4h2yT1JD4IfqgOXmn
O1a6AU8QUqQfNUE97XTRz2tcBAbN4ZHTXcWE3ulAujngQNVX9g1Mn4R6z2bDZkzI6UoHfOEHY3Wa
FKKotPDfUuw9GHkBIg4Zf4EVhNqSmn/WOnDEcpukVysxaUyE5F77DYmZWgDjgT4LSuVkASGmuI/u
LozjG/7lYoKnc4vOgiud2DmTHYb7+CMuCWyEeRn5syZSlbPBrLDOeuF9Ihh5kiUCr0Lx2OHJLmV7
dXLoxqossf09J0AT7oaCEB+Q5jqDdaX6Cm/EbHdOx7T8qNnJavRRHNLhTTNt4MaksRTZUdrFbmPc
tPGSPlymPg/1HAVEF0+76dw/NN/V3MMlD8t1P3dgX3VVnuI3dZBBEfLurc9XgNO0a8k0XRbBRpCs
oLpD4AMp+LIfTc4CGJ8TDYXmKTiz7qeemp2tRy92vl2EbHPjKeBhB1iquS2V1jbXNWzY37u7mSjj
wLbEiwIwMCmVqnc2x8obj/TsSxGD4TbugPK6oDw6z5iAa+SbyrDa4KMcNaayUDeYlcOSFgtHtqmv
EHTakTWLzsS3jtmw3X69KZDv46/F2rqWVaE/l3yYlUtCZoJUG8gwEsL92b64mKPv29CXElc1JpcI
Y5DOh4QcaF8ppZsc74oxZPDowApnUOBY6YqroUVXCKDCb9gJOPbEHFXF11B1cJEk6eRFzDs0sWN8
rzc3Cyl9xmRmDRzJtPokzo5RK3drRttqCr0PfWV8Iei8QgrJDR9HtFONy0R3mJavg4bR3S8L3fkD
WGISFIHeHXIUuNK0lY4qlAQvmhi6ExL35f/N8TDe4jmSxRO+DKkPepFUfWf+fE8xPr5OcuNhGpfA
aGNQ9AmvLfiA1jx0pM/DH4wabKueIjS2+L/iTwDVWVcdD5jRN9Zti+7UPzvIKLbjAvqm/pLoT0S/
ut+ikqpoQ2ZdenuT+tOC8SwIUzWR881ma2owZeE48lh29qLw90FPP1puqu62ozOOM6FkrFSGFl7j
ywg93p/b6Q1fmvlFfaidJmn8e+1+uvyPP7uQtDKhfG9E8oLT31uuYNJaagpxACw0ZqmGLu4s1kyW
wOQg2iTN4nyoz5v/eQEfQNupZWCBeIG1jMJrZTdYPNdLL5Wc04Ld2Gz2yksaTd+eGgnDbJdnXc8n
bpSZbkQWqz98FLLBAAxuNRKDY222q10DubTKLI7rXy+kk+b8FUHVQGWDk7L1IaN6seBwc7ggt7d9
53qwCCWDqVy2XsVHe2IetE3DnUpvRrUrfVp/647q4mtoJ7LuvtYA+tYCx57YVDf8v0E11+tiZoGe
xZJoMlfivZDJZVIiv4LvSccsIKpf56CJVA17e9XGvCqMnHmC6kWq6oplNdov2kW5e1ep7GWaymMJ
Y/eMu7WAAVVtJTI7zAZqoUl1AeBIetF/i5NCvnU9z1KDpbGleTvO3DSVVvfggGt7LFwcwqqppu0p
ylRCgCftdDvVBrjVem7vEBbrGV8liksb1ECsI8hcS0SB+YGC5mRdxeOf8sV+J6TSG38cBFDdJuRN
yDhKVYthE1rKUUY3yePaSLQbpnu1yKNLwUzc8Fo0GtQs7/ehMbZSrV85euluzTmK2fATi7C3qsrN
/lrAYbHPCTWDaDhpa+YgWMkLSoG0/evYMY4Wr2qfSSamM6Y0Vas2nRUeTUA/w1Svx7jR4tNPDL2Q
YqEMOrRqK2x4P6sopGCULvaQ+RJ5AimJLYoVFDRysMlkEM9eajLEuXHNYNySpQuBW88XBMgdCIfL
2dDN7V8YbDMATHz8acCBlEld9acHTvGyNh4AhpSF29UclWn4S0WHsuL9a5wx+Y69/+kMzguMG+7o
ssbt4iUa8LmDJ9PvwkL6gQqcWZosUWSU1/yau3vk0oBf1lY+G/foB/k4MqFmdELkyvziGrfmTZEH
Hub2SNvkXtgl5yq6iGpPHo9/xp/ccDr+OPlu4Iaad5JzsXst0xI3k/bFAXuY2MSxOsY6QgLbqpcG
pJCOWy1uiR9Vb110JCICzn1VlBLVW3gCRLetiYzHcV/bch4aXa/vBaNwUHgn5yprf/gnup6JYcpf
DH11tNsazOoCxd1ZUGIctvdpmvNQnEI/jY5H10MZ9ojgNQzRoUxOP9QH18lZ0a5HhcXZwrLD5Yd3
4i0trMjWExJvNsojYNTh5Ux9TKllFTn7h31/IY+aAElkuXv+UXndAcyTJMvZPg3WzIqAGnBK6jXX
nz0aZi/DMyicXgDmD7IqSBkrLRWE5u8QVC94zYcK1eAkJjXK0TrZnjxMYI8d1ooT+KCSYUR+hwyd
Lu2R7ODN0BNhnaqSMtZGzQKP/c7AF/HyRdOGq1CNutWMaTYGdIEzcmhzNpqJ+ris3sxf5+3di4a4
W1hFqmmzH6g+JsmdKB49GfK+JFco2dkxCCBLfIZZH2md7fjX3UW20BMd5C3TdOxOaSV09o43rVkI
NfzcLscLscBevc5ufopM4FSMChykCpoo24szflRLDq1czD+WxBaxkF3dECjim3yIE2ANL/wWS2Hl
PVIHEqMfVBi7TeHQ/Tf2sWa7avrkB+fFC5i5z7HMdVqQwIIAW/oodtJVUWShBaxc8v/3O8+nJAGv
QvZiuWa3nnM980mMaMqNR2/GkaTcU5w6KO530iV73/raXJtC9GnDn0zzhSY43Odt2L/yGuBwBc6z
j5MZ0TNVoDN6mvWgxjSWqOz1he60w2SZJiUMEQLugQ11o4zNser/LEhioDcn+n3+EEuJsYkdXQ8H
v869eb4qSaqhjJvPD1t+nAjbAOm0BobYY5n301c1b0KRDVR8g79oQZvJq+1u9xx9GGl2FhtWih5H
AjVLRVU8HX3GUz/rgqGb19NlmS8RMF3MYkQ+dVLDLwfGJwptysoZJ8fi85HLzPHz3BxG4mNeM0fe
6xzdBnJWF2iyK3tupQpxwRyK5O+dFFc/ymlElk9Ssjw4YK5TguUDaHJbpiDJMOnwc0XrQG95JYyf
GNBdbE2E6MQqX4UF96/wfz+uWT1of9gQV5bu/465N+qv0IXWwEbJKSAao0ghdzoakG01tYOTvGqq
iPKcV/olq6b0sp6uM3mZq45fQCWdgOgKSio8qaebidQ++37PStF7uhWgjcq+O9oWIuDTD9CHSz44
YwFynnzn1X4GhPTl6EeM71JkF8dDlgR0pPb6Bo4FsqGO9wPE2m/iX+lgyDtLIqdkAc2RiZhs+wvZ
fdj/+pUc5l8aiGv3/fZLG4XN2WhGFNGlpe6SHbJDw9rDhC4mlL23vnoDUa65Yy4zmtqgNEw7nB7q
4+ykYIEPWHlrCsY9olJ+RqnrAed20SfnX/EQ2gB5UzWAbU57NRJ9mjWACh+WxhCnC0jA4FETbe2R
qFu05fADY1EnGvTmGnhCsMA270G3K1XO3f+rVGGeByEnDxOBjDe5cLC0n4mjPQgCaXYjbhaRFeVR
Z94Qf2JOR8XhCHZTXsco5vuQjJgXJ2aAx52ZndYQeIozgLitBWh/Frm/i53pjxO6kVEWOpU14m0U
9B+7pp25PYgaJI3ACy6rhk9izCDJ4AP63Rl1bRwUcI+dUI15MO/3VbnHL9fqgFvUILsacgDc8LBB
oMX9SWRFiq2Lv8nUOWTDzMhD1KXVHMv2tQ5NhAwA1m4ubjIqJMqcze0jjUjrM34dwt8RhKsiPU2M
7h7+yTpGClcm9QGvpOW9VRmz8MuOR31kKSMVuuYLogXas8uJ11Xwzq2a0PipWorpC8jYkkRpL7he
a2W1YamdE3uxtnfMa3Yyio30eUZsYy8ZGtdjxJlMTaiRcwqG0I2IvMG5Q2XFsqPIj1C4FyQhfQ/k
+4Kukk0+WuKaVkmsg/9Q0NlzVWG0hnQhw6NGXSbal36CLcBj6lk3x/9SOKy4ANxg7ahPMh8ysoQN
vwDtIeJ0aZ7c4GqSRr94LLsb2VKwS7oJnEpKzs/jp0g8A5OYe750ka6sRHzy6ZHR3LUSX9gBCVO7
gwno3q2OFFZH0khFhYJpwottln0T0RtwrfwYiJy/b3mTr/BzniHRkxvh8YGGEd/mCrXsyTQPffbm
C2bhc7Gq19d5xbtwvSV6BklVTWSM8bo0gnqEQ4SSgEHaffz0c1MivG1PEkvEo980ZVUq2ueX7uq+
JF5/N+rAplmWCRyDLZdWEql1IBY5Zo4Q6IhyDzKy/gYmNTDLTkuSfHTUpU89efI21jl83nFinG/M
bOZ9Tp+GwmQa+NNRdrQpViP9gZmUBVgJxmjrA1BdKYA8M7BY9gK5jgYbN9xf9lEmfRt4AkKWlPoi
EbMulqS4i1iF3IE2MU4AIATGcYvOc8iSDUiBqSbcXHZ7A+qlC0opXsLcDr3pOlysshNnb+B/rPU4
OBLoulll0+Hdu/6YxaaiMU32fkFTunFxVNp8JXKnM8LvByJ+WwWr5oiIlGRzHCfZo9BTDsxOmv9Q
wS7dWF3SsiSm6znEgw65gTJmkahdOTzDjH7DiKA5Hbo8QPGTIefn5KUFLESs6/Gh434PQi0Wb/Vk
5UPOSopr2S1JeOS88g9OYDYTBgQqy37x0UyShMtn0chOja50pP3E0SlpOMX9uDjMunF+Q0OXIhKO
niYzFQPZzC+5YprhcDOGrUo8hEcJevNCt/sYbWE/8cwYLBrNvpUp6RulyW6oEFVJPm4zqgs4a/tQ
szUFDkQIJ10H1VqzPuWooMttBD1MdSWyubwMleFi7sKaJ/8y67tkxGXOsx3XL/SP53z4eWYF3TY8
M766cukRXP8atmGRjUS8BDSsDe6cDyj+98fUnOX/Rx9USy/PHuAzuhL3oL+4RYbCSPitA4mBpseX
qTFt1P0FUE24lBVjDGHgsXoZVHSBV45ZAjNJXjU7q7Tk7knkx6sqz9Ye9xPVXLE8pgx3VmggLy8e
SJ5hBqXk5BLlB28Vi/dR9qQVoltE2A7XAr+v4Gvtxwvh0bFPPUKme5st2b1XONgpRuD3JTp2u0+p
aIUUimVm55mg2z/xGa4xiaCGorAAhyTcTYPp7OdL1q7oxk091BApqSCS6YdR4pJvJXeQ8N5tT1ON
dgmxlneMLtOVUDY31WV41DUP9o6X5HR1cFJX2jBiPZfQLvrWik0k0dTUzs7TjRPbvBiK6LgOWsky
NdFTL2RSXZGoII3dtmMOZ8Lc+EQDOtupVlmYTHJlJZxzr+00pq2OiPMlQv50op8LhN3EqiIkmoCp
xGKMcSsFlIyE8F60gPt1OZ7W5S2nwqavoAUcgVi5PTxzfZX8f2fP5gvQ7ahOf6/MFOjKZQKNnBAe
yXRxbg/uo4nDJMV8R/ZYFa6nWYsR6ifkfdafY+O4fAzoMP4roxGUX30RWlCgsRXcT1b2TxrqRCrm
cbwQrRz/U7xrHy9Qar+hU4KEKjxz3jvgK95xekJ3MocaxKjW+Pgmtz4LJQy3usDSxJW7MlPpYeGq
N3tC2vd9AvNrIQBGHLnv/O/d8+sN8OkG/Ju9GpzIr8ycg17JaMOVfgdAke4xtH4IlNuXs4Y3DDKO
9vpILXjhhFMTIO+4K49VjanwJwbLHj2tQ0JIxnMFVrezGuNYuRq3oXign+qL69aHx+uX452yfUeY
1/MtYegfn3IVG+or1T6H4sQa1leBYXAD7kVminh0qrVNmDKBv/FBQJA4xtvflCDtgntANwdSdcZg
QnCCbXEUnHDtQfGL69AJxY6M2jJL+mGb0j5HoLKr+VRSJnolhTEtOa1TIMRiOcu+eOSauj465Qfz
A3IxVevJLgZhlz8Ovrgzcddo3C+C4jpSetzWPytY0bsmgHeZjXsg4S5+LEjjiQj9uxCcCQFi/4Z+
O8JDgvbMU8oWMXbNpu3qKFfeb7pRgi8kyGu6Muto3lVYDXMSoaPgZ69P6WadnlH8yRQmRhc/UxFt
bX5KB6qFLH6k5VdPYgHF+GaxHa0qeF2C4MnU+VdybzbJu0rEmZzgMCnTU4IwyugPSQ51EMGrbTOJ
RYEyaFl0/6udEsVzwWkNmsJDVfl7+uFvlF84mQy9F3l/AQQMAvWtfdyVmKUhCUmi2h/jkYCIHraB
qYx9zi39huWZBLJr8luDYdaoinXa9kvS3tvkmOHR9EUpChpUpyEqO/u/Mpl5OBg8AOXFQE6QG8iq
OjoqP4D3TpYHFVnGlwOoMv7hVKo0EAj2YZTItfl1ogao/rrN97ey7BL14O65IIUH0d7JsnJS8CkE
zhRizkXHrJwoJnYR2OGBaec0Q7i7siN3o0VRkFBgiDWAp8Pp6brcl06whwEMZJ2xBLWnuz/Gtakd
pKECaJMcFOeCSCl4kZAct31/S2NszlmWdKZFxMIfoalxEn8XDLT1Fc3QRvoalP9UvzuDfXEL+3ks
uyMl1BsN4HMWfwMqazCsTzjg9KcHa3ySzok6JYePpelaD/M5iAGlVuvEKciNtuOAYPwP0sE6zG6N
RhnKZzcWuhkJHG4srpywEWvDkLNrPEE5inlHT+bYnvmk5tU5QXL+jHzqz9Nhgsfq4AZxp7VZR2lu
o7n6zrsxxbn71UHGI7Bie/Jf+K6Wv6epS67wbxlpN55sdhDRJPGkLJME2/x4zUCnrH22mz0DL6Ru
GbqvZNzUR+ydY1YjmI7gjJ1zwSs7LtvFI24/PzWDemY2UYNIvOGSKklHjKZFqSiJDvC6/VIoHhiJ
WvVsEeDgvymHfdKcVR6U7943R2KaV2SGpXQ6il6exk8250fpPB6uzXp7jruGAwly3RAX5ubTNHYq
V/yFW7pKOMtM5Q1MXKsz+sbPF2fcMHRi7p7EdQeoI/spmCkvuQ5gsineUzMobJ8zZlQDNzoSRbh9
xUK19irEPt8S62o7dsr/qfyjpmZPHXE1vXPs1iLJ6omTwAPgmHZzJuKaG4chO3cpT8hTJ4pcN2io
FQjaJajWiQJvvinh+ycgYmd4Sh5o/8NdlK4Lp+JHZu1EKwbyBntF/OjljfvsnZ70LMB7qCdGQFMz
xGbqSEvHZqNjIBhc6ISpH9+uqSmY/UqwLrWaOqTtn/OIR4HydAiQiH3LpfSAOqqPC36nmPr22GBr
AnatVLhPpQ8pzn2cJtAHzR+NasApVP0DSc+gQSHJxvHP4ebkuo7tYMbrv7xbwf6m1EqC1la0ILlX
V7jEBsNfhnP4OMJ1NUmDTCm7Yp1GzH1I6yabpG1fmyhfO4+D8QcLoT6XLamlh0gw9yNwQUfXmYld
8oswPT6N2MvaaAL6VQwAkpHpc73YzjBDOV2SXMD7gAyIfLsAcrc2N8C45gGsrK8sUMccvz83jjf4
OsbuVdht5/zNEgY9W/UJuRrvyKhaBn8q1eFtQYnYgNx2Y6mJyUNns3rmfpa8XlaNmLrh11juJGMf
3FYURlrG71p8woAokSoYX6hVkwePEGuUIbFPwaGDELVFRyhmt639cJ2WtbdaeQaoXkFhMeRoYoSQ
xNKjjOA+s7Kq92K+/zRLWT5QYE4C14ASlVx4dGFimG9+4EKWtFHk4EK7JRlHZTM1ZKPov+wGfzUc
XYcoI9YmuX21y7PV90aJxV5G6xHMl3hKCJEUe7Erc5dfustvVOyHVR3n775P2w+ZljwzzbUsjcvy
HDhcqCh8to121ntWXnxKlyJP1YKWB4fAS3skoYJT0pjoOTir1m+eORw6avm0zjx0IdTj6TvQgtZ3
kF7ICQlEb3CyahGsdpWNqbak6UfLltZ1WBqDO66EU4lPSb3G8oDQJkF5icMXagHgH4VB/+y5qZQ5
uFin6lIq/LMJ4w/N4bXUnFLfP0osp8Yn+ymBljYvsvJ4hdimGXFJJqTIRXPrSrTDwskWfXiZddUj
//NNneNWEgo0/QXBLJtsp5ZXoMRYCq/MceKJUOsXTzmSVcZOlmA3rdxF2U/8F1DPiarNScFqZWUX
p5RKvdt+BBQydpRoKRDhNIcu2xnjdP/MViTqol/BFcqgASSFpTwTTrqRuyEgTbZMSmxx5cPx65C+
HuC6rik0M/AqRkNzTomzICkPHscG7pepRUsD1SljAykhdJ4P+yRbQXmW/NCMglSTv2Ab8KmTtRN1
cUv7eppC8/BAzZ9F6hPRrrtNvB9nek2plj1DEeI0sZ6BcI0BDvNbNpnhfhR4jMPlw1jqkDI/Txo5
AG4Ohc8X937ZYxz/2hZN91pfe7mg31bxnuh1hGMptqzukaOv0H+5fzPkUKkTi6XsCJiWTLSn5T4W
qW8rPqWw8XLaZLDDZHoqEaHq1vcHoSnbSRTdrWepcWxOqWd2cKjowKLoJ4LuSfTdx6MIAJbL4FI0
iD8Or1ARlwJ0hFZGN244l5JcnqODDVmtK9IA6/5JWKGCbzHF++yX53/0CeK42Xfzh805cRIP0rVX
dKEaGFjhAhUSmGLd7VuLUuyiMVFDm2bSUk1kPDF02YZs3Zp/9yZ7hgQtpehq3Rmnu5rfQqQd+23L
kL6O9xUa9ISsycfwHA7S9Tr5HP1dAjxINQ/jbuX8PYgsT3RHQ9Bl72XebO9VT4ECd0VHSJbxUgFR
JQf9alTbYyL2rH+Nrx1yDWHK/o6z8vH1rNqndOLPrY3EZU412hIlbgw5lzpA42Lt96+Lenno6TCT
SxUfOXJ7X5l9SUSF4eiEWisiGUEsZHz3KKSgm66nja0Bf+l8bYT7HuGKtsGSPEfHGQ++xiTIzMl2
ITPc4JFo32zLWCFLCePo5FP9XXDVxUPBstlbo1A6sKlwhY3KCSLkPDYOMKF6ngdtn3fbRfizjGVy
6WsVLBq2XBQwT81s+LAdGcJq/xPJYCImGnFlFWIl612nQhKnSQS/60U8A5P5dGb80wzxFZuO0mXs
X4QSqJfnZq98J6DL6n4qCxhQYtZLktI2haCFEnK8PgrsqRYCubV8TGeIi9m3KbR2GTceY5Tu2m7d
0z2mwQrucNEBXd2ATZY3jGTloTKUopKdl1FkcFaxx8fIjK6QlM6+C3wW6ClgOnBveLv0bBj/jkJ1
EKyMU/mCrkDm8WDmOnC3aAyBQT5+o1Ye6Lr0WnJX+fKnTWEZEIxAfR6U17Lu4HKSRsQTjpBIDzzQ
iDcKKFsKWS/UoXCT//hqf23OYzngHPSJhFLnwupqn1GoeFMKV+2TkS1wMkaFxNqGRNpl5GlfmEyB
TwUhW++eCyJilhpfmCRPnSJdPv/BB/rwiruytdyZ/bs7Bq+V52dQFzG/2R062QtgWuC5bG1Q0IZD
VhXHo/k/NL06HopfVKmh0vlrTdZrdi/LQ0tGx44PWww0NkPVx4YbWddNeFeetIq/tCaOUIpeeyZ3
uy12JuB3sOd8abHtAynT0wmjCTo6/RwxNAe8pqsUxWMCa+TJBjqwUgGjiOwicBz1D9yrumoEBrvx
Qr9W/5z6VGZL7Bc6NA+j5Bys5LaX7xl2lPK6gwjFy4rjs1cqpslKm6CiErTauIlUcg1nLyn9wpGG
GURrSO1DSNnhJMVtdo6JTCF2nZ0RFRNzJmp0vPZyD2ek92yvGIaQYJlFVVRjBjDFkOWw6ThnHCs7
c1LXAylunRl02XLOBzggPQ2IjXIdtnG4WUCs5uL2TJXmmZMHtJJzr8f3FCO9ivz8e9LU/O5N+gwG
11L66O/8Uk9311gA1ORIKQ1NOheaMXhk1YC5jrlcolGhAntjzg1NPPAirhLOxfLEEAWjIfwygW2G
sCdmlvH4U9hq6McOLRL8+5LvoN3BMq8wntA1kGuQxiGlqORVbXyAHb4617a2FNgoo5L+Hrj3z2G+
OpJ77bTyFxG59HiIfuTiHmAbbcNKzORkVnxeGV9pI9LFo3cqBrpZFA6mlht1rsqeiGcBJgWVQcsf
5q8ByltHEJ5L+8w548bJbIuLqufuGnLuJXPJA5HqUEbFOH0d1/OR/vban05i8P0eI11LA4ICRN+a
ed8jZfgBKfJreoLOkGPGChow9FOqcbrF31pwTUFcs3Tx7/URHiszLz99b1iXaPt8dcLNKYNT6Kgw
ru4aafEOIJ+mE+F0LEWAjKs1BPpUDGc0QlJwq+o7TUmTU3oRas7DOWfgpW0g0+v/Iba/W3ZXFiRS
mBqbaSOVjJz2ueMkh5ubbuYGBzqORO1fYJ/CkSDN9Bz+A5vgdrdExcAYu/b71EfHKLEIWSIvklKC
WVkT9xKkKw/DldkqzSSlnVtnLQ+zBhXzrWIrSrgS77m+x1cATqXyHBi0C2x9a7wT3l5RNP3M1SOB
grl2z4fI9gxRkRgyP33AY/v/+fj+TIsoZzuikfTfkvHs5eCSljI49s8K0LXkoRA/1Ykfbm1yZ3HZ
rXD5asEPGUhnxhTFqUdDGUVGxFRIy+o6A5nF31+VHKUNmvVafFf1F5aH0WuE7Sz/nZsTBCUpg3H9
lvlqjtXQNxAsB4jgqyhCiVRW/pbn4AHoQopfXNCa/k0OPpUN5DW8GygjWa3h8JabmV8Bm9EPtzd9
2m0v+hlpNGMyseLMBlBChS24yG/ZDW2iKXIjIu8GjHW/1D1KwiElEFuMhzY/1ML/49C3LuPEVrJc
uef7TENJgyshGlQMtkAuX4dy+73Gk142sL3/THNbzdRaYdtHt3KhralxlAMnNKO21GauZEASeGiX
9tL6oXzrTEoE2s9FGW2BThtFwXPoweLS58qkhZX0f/edW26EYbMyLvIuxze32PQjcrqn9tTJyGfO
hdjyQWWjI76e15/MQ4/58BZ/4CPd9/G1DZkMSnvqruB6CNP9aUoxNaNCxsWWjcVRK5Pa+SUxMX2Q
AqszVnKT4NmtnLSPtLercvlhdihb0vVbeWtDYsvmMDnkZTy6RkHv7lqlB2dadshm7+dPpIk21STU
SKf2j6LDFoZukNG5IAjKb/hy/JbPylz0chX7Bob6QApjvReHT01wSqoB29r09FCa712rnXsURUj3
m++p0fEwtbJntBFGdmUyfqD30lWvAs/gdV7SUqq7Yku3/Vesee9QVfyizPp/euoECwZMYQ47fa47
jxw1KzknVbAaJslxLrZwzGJesXiAPSvEUJm0rLIIHeU59nhqhX8NlZK3yZ6cYfNm8EsQXsyrGBgH
Rl6sc4pJ4FP7SZyEx8IxTOzQCWvY8BrgULK8HMVu/pxNLYgNG2mVsuwe/6a0qWLPQbplo/zGAE0G
J2P6GF+6L3TYlExlEmEJ+jayo1rwYh/VFPaT+tcirs/C2H0EZBHVf3wURjcx7GdrqqZT3MHncWUM
SS9Etxf9TZ5ZlQnrcsGJrNjuEsb4IwyLMGT3DjuB4+1uhyKfwALpgxEHiB4/Qqb/jXhsAEWtzqqR
CSmKvCIH7Nva61mlUBzrDg/7L5C0ZSC9dkeB2eoXaEw4WNyvVdVVQYYUPUK/ylxXzZfwrtkEMijL
7s+L+cWhPGQYxozucl8J5zx52B0MUVhR4XiTxpviKd5YTgMPdoCyABlv8/1fxJWo1h6wv+x0jlE8
+imcJvVjSCoSgDF0x8xM0BunCyh9p7oD/ggg/zLBjdZmg9G/9ve9iRwzhaC/tn3N3wyAIq7vrSvU
CAOQmCfFuhnQB9nT7sh4uu4FVGNz8u/aAiW6BxjAMOZFEnkQxQAEE/+oJ1ZuGuAfbK/b+8el77go
9xMw6q5N24ccpMEU85zCo44Z3qVjqaZy/z1hIzOzTVthJGmMnn0sbhqjlJPcyJBNmJKeEpphfSva
9Vl8r+AeBD9JtTSfj/3pSZluIxuDJt8eM1cqJNqHWypFVaMYgGSPiQvdsKwZy66d5efIdjCaRwz/
RQBnwq+24lttlCy5NldcngqKAEW8W7E665NBT//xjNagFACVyamsO1XIVZFVMYd1g4UAZCOZaIXU
emhR0OV8z9KM+lIRyKsfKGje2k8g0h+/GLVhLB+DLYfQjJJrcUO0ow4S1eGJ1AS8NmjpD6YLfvdl
dKhLTLp1nDrQ57/pCacQRLHNxdO5Cbi83CunBm1yJeMuLaVAUV9KM+zsk/csH0PrqBI3NlBTJYQt
/I2crmZhRaNI/75y3yRkHRXPte6yO6EUIAa6DSihxlpT/BzE9l/zmIw6E94bLUK9QOKxcDIAbEao
rO6Sg5+ehYE3asBQyuWSka8Bw7q6VoLcuLWi1XWEZHQddQooRbn1apqM9XqwVYlIVkqxB0f/HhmA
vAHXk2ZDxpE4OYxfqH0KsMJa/JfwV8VCPk+zbwy8XWPJaovQZOXKSxhWAYw6sVDWr0OixNHmQuOn
G/VtaSgPQepzItmx/0ggrWRcUnpnesfw8vP9J1sIdBM/CXzh1I8OJPTcWX/SFlc4BdBPbRz+HCYG
4P+CU80oVO7KV9M5Q5sNKEz2TRFBDZcpzJRSRTDq9+Fy0I2lwL6GOBhSsB+eXxQChM0ESn5SRiZM
RjQV5JLdvdtEZA7+mLLs//Q+ppYsVZBxklcyiQvRmYtEtgrJwUKvOwb4dQB1sl0mNTkoJxgW8iQk
Fe/hQXToh9y9hceo9RIQVlO1FzQZ/5dL9i1gTNbGt69S9alxDlcnK8Y4ZnLUnYcz39StesSwsjIu
ZbxddlEMFzBxKZHkF90Mhbb/r/V9WcvDPVWTMiratkP4KrxoGoXfKPY00U/4EesJJKWqLpdqT1WY
eDugeb+g1yZhpHC9pKBGkwfo0pcW2IjNn29TDNqLBGICe+xn7Ubj0N/WP3DAzL2v3l2oePyT1YsV
8jcwHDWFythULw7gvMtaw799BJoVjB0I2oPVPebF0vnW8C2mYJU5GcoanvEWtjlqqwTOXgZWJG1v
y1hhoRwOcEmzswjg+4rQzUmEBc4L/KghPNzsXV+dNFhZgpN5hPA/hxwoXMoAACxPh4ulo+TUsgev
2eqW8wBfdf/ETT38ItuScYKDCe7BXc+Bag77waSU5KCt1IXxBA3XEdiSOiWikDca/C3sKjwWEPfX
sbkN7pujz2nYXraR7dwVw1s419GAoa9+geK3juJ3vhi7CzjzAqX/bNA5v5EkXCavgd9hUtMJYqQU
McZYe7VjjeUEar9rk3csYL1hTpCk8I0I8O4mffy08y7v1UWxgrlvp+jkrViZqIGhUqOIQW+0JV60
caKcYuziFg/xXyYSqkFQzxzpHJOS6uI0PF5fr/iiP/LXMruUdny5aJ2II68AQxljhR6ux9xOxSJ/
KnA7CxI33Pb4Z21YyrLCYhjZah1au4eJBrg9qnG9FesTxQmxaoUKHA3QffEKC63d7acBV7/auzRM
pwRTz+99UsxHI6JR42CP1h80iYSVMXZZ18CwObtSV+K2pmitra7WvOuBc8nl9zRfuIBuWy+YsPET
RyU+BcZlabAyIPsM18GHOH1QqfQ37xSNWb06hS9LSdqlrOycqz9qiaZ6xS+Efb5NT5Wz6dtBjYFr
Vne4zTB5+3LIXJccT71p1xbL1qEPKSdPwdbJz8OM2+1cF4gj9wnivd2sBkqn22fblPX5XNB3awTo
U1eafWlBVd8PtfJ5hIbuuVM2IlfpUiWDqlmabYznbe1vK+8k489DdkC8audc4aXRZoJfuNLUNo7b
fRH68xtxqpl3AZrhO0NFVZKiPCKpHm23jbVlFCiqlZ64N12nAtIXpCbhzgUR+4lf6Y06xyT8TPTb
Eo4GIQ5mhXhBVFUGOZTLSo31UuMtl+sGwC2s8pdNOQjn6K4MddSGGvQATIJVcKvsYUCMjlrxRtCF
xe9+/+Pbp/s38MxcHnsfqMI4uvKqVnppl9dE7Lzah5C45Mt8wai9C18m7S+wP2/nuKD1G2ehMsh6
ms943FKkebYdShqJRqhxcBva01IDm8GMgSSDVh21EmXl4M4hnuNcrjdmr6gtcsKA3Hy/xmxZMsnm
/wYKIOF3AA+n/3LkgVZjDTB44K4KcvEKWdfVvZ6jl3vpFgBZEmiC5jZYaX7FeQNJ2zP1RG2oM+SZ
Mlf3psztEqC2j8ZyAOmkizKOo8/S1gfHWG+9cPs8W2C70Of6jyeYJZGV0c8lVdhYjXA1rMvq/pkW
sawz0CoBpbhzJNVJd3kBBwwaVQa/2DEqgVGTdBi75ASW9aIulQOH5SogtElM4wvvnzEX3ZuNLkc6
p0q6AdpetXapYYS4rB0DnCqMz8jHDGY2kxeLb1n17dfi2jIepugcJCqYzK+ebypvXd0L9D+LBFlx
HRk3Yq9xKV06YzewSPunbxRI2POJ4G5x/zJgtdydcRKjSEQGoVidbvU/unWGJu+k65cFGlXfmuNq
27xrJ+3aCUryt6J6yZ0C2mO+kx3Kre+GC8pOuwxRE3lAUVzhh8wdJ6w6YIR+X3xxrKizif472UFi
CdHMuqM7E0kyaK1di4rmeJU9pXK+a0L0Mdr6lXwqv0gY6xsUi/qqJff04Q6qTvP3ZwkjiZhuiBTL
0EfsjnxVKI0MWXgTHwNcFdEYX6R7xTswN2OCF+MAfweqBzJ0Lwc/sPi7j9d7rgCq+7cbIAG3zQvP
QukQoyzFduFKFbAnWN+SzvKkGxN1BMYGWysSywCG8Cy09vVL0vlgsK8bbeURojm4sTPJfqQ7zBet
cQGfMmCWWPWDR0gMsfCdmf/c6NA7wOY01nRrCqPy3FlmVtZsbf44oHB3ScRyPTHGNUBtqIV187L5
Tn5TZ+hDmUwBswL7R3BhIKzRAudwkiwwBgvKXz/1HKtnVIsizM3JPO4SCmGRBs/92w8ooirjr9+n
zvf1cYybUCbRwERQrSpougrf2qp64lNngIZSYupm6sgCX3Q1QaFaOHF3dnxHvssoIePOWxPnIvCy
Kb1ze5g+p+GUlv+ULPuCJImOSlrK49j7CeDZsEemAsehiG7z+Om4oFXJmeboZjAGyDKQ0RgcuI5s
R5idbP3FyI453nP8D0xnhrq4T73dZbf2vIuWDMWk+vWHK4HfK0wERcvawZfKJKz7rXcIrW3Ku4I9
plXLZ44PakuIRGlpf0FlmFkFLxdt1ZU4B3NIAsCTooRnYZ4TI7GIhs0YNU0b7U4Z5RC9FMT6JGPN
Qfg8lMjGT+q0YnOjxSnLV8v6gIGYIXPqLnTXuyDmIJgwUYF3347befdvx3yRFmMtXYeHNka7x4Fl
KSPoOZM3AJamRU42edz2W0Mfjks9xMs8/kQROpu2//4+BA3beDlc7HGQfDkSu8ADXZojIp5roUsE
EQpsqnjOOTA3QC8Tpg1Pk2RU7gjYPdgZnyS5HPTxUyqrzJrYuulNDezwiwvlbucyYfK46oAyg1yl
OLNVM/j14E00syIpD+fy+jx7Jv0EOqSWAo+ceRw6ofadgU5BfS4a7AEeKWPJCKYQbl3/An31gdIQ
wp1TYpNDoxkLcSt8u1f4+pEdSOK9sto/ZekSM6BL31yHPiwzo9aWLcUNs2todqH4g1FcX5fgng45
EYpF3/wjNYWc0YTP0waHq/TYrBAbC5OTG6l9gByZM3JZHsoMIniKfS4Hhg8ubfNPyyJ4KkP2EusA
sZX/Dep8dBzlCtOiNZbWH3vMjEfSejqxJb6V+2fPzYU82FxL+CZQwY3gJLv35MfokRK+kAw7U/5i
p01l+1FcrRuNIEJVa4ZNrgsMAeLRe3+6XqEnM2BkDLdj50eNNT1tefxT8orHHAnZ63JyRJ99NeC1
uRKBQbJ/KlJ48se2Iuhg4xdSNqtMGB1jT68STqpMgdnarnXAtdgGpdADwPxlPCNAcD/QGRY8TGYd
/E80mBET0sAXuzIZ5PyAfKUSAfwPMIHldZro9YTmC7mPkjjm4l7mMIySLCgHnnEBSVXab6YvaYmo
J8HM4XtNisjrd8boj+l8+xS9CWQjnUNMediu9dTTmf9U4xC+5+Rp6hWSqZuI1YKQMjkJ5aExWom8
GJ2m/kNKq458YbxgHiZmSj4AiwXTjd74TaV5IDh3iYdr2oq7FKUNn4M1ktABh+IkLYYeN52xO+iX
+Ori0ATGvNFg1KozvHzpOdDRQKB+fm1sNmD6GtVGqdS8UBP076oCz+gEU2fiIndX00MaEe6LNUhu
D8b+jEyppFDkMxsMX+iApw/TDYX6pLOoltsc1S/fOBEA7hBTUEKlH9nOvZ6Zj0DFWuYhqKAxNTvC
tkW2VzM+p1qZu+VV+3LFuSQytTiYSbTREmyK1bCma5ZwgO5ETiIITYa0Owlxge+kEJgpjG4WaMyT
OgutImEdnRqnjPSYUMaUS3d+FKY2oblGYoLNcSMahRkxmWqiRJnBX+0hKf+ov5HRnNlFR6Y+NF7K
uqC6tnrnHSCi9gpnSp/HgXGWOzmTUkoeUWEcLpLKZV3Eqztj1mvBxVsrR+2FJfm1EtWYI6haamYn
fS46A8OEHZqnEQBnOuqTweZnQXl19HavJeOKZ8acUWY9GarClVfZpIsbLnPBA5do0mQQ0oaFlCP1
gXee9oSl4TxfEJ5Q7ISwKhn6zgrOyTz/0CYuKSEBUftK10c5oBQ5v+vwglG9VnBBlnjQaqYpUQsk
fCPk6/lmsH6fli0k+IEq8qXOGJatBQOfts/0+NivQEcpMSIhHVoFQrNf5LfFRZgfWnguMqlym8zs
UdncCNSYO2nxrxIZX7pMa3zpKE29EhwL1cleeTz52jUOTYEavbVco/6w8p5v0oafQa0zsEYQq738
LWAMA/7MUek8CBnY6IxvT+Iw5PHMzuJ1JGX/VKSWnHhyCXdzG4qI8xdV3uxPwYpX7I8d4z6cDO3w
jk5Xw03w8r4pOss+NDHQ5LsXzPmZo0CS5p8cOWwiKSCPXFjyOE6Y9jLfBTEUxk/tb4O/8m6VOjby
NiOqPpvxj86wioDpj/TzEXwM6dNTlPaGgBjV3HuoyhGlPunhPwvVoG7dvN2MbnfD0EkslopDV/4L
yuSWMCxiaBeHscnW1I57eDCU/HuRw3ZkQCmSnlvpxA53OLDk74xv0QIGVg5BdDb/2iF4P6VvnJO5
+B782CtNSfKQ9+EfD5SkBooQ3RUtZd5veTnmYZpy1I3o41Q3NaAQECinV7flBWZ7RPOPQd4JNO84
O0KUVM0f2+V/cv3U4HVZ67TH7qJA0ilAUZIXhL5FGeIvGlRBuq95lkIbwi3g0DD0fvtvt0KgWPVc
JMVM0ZMShRL2Q1t9pKFm0QWGM26w28YbamSqu7o7+lQKNgEZ9ywskPRs22r04uneOFKrQe6AdcxI
GrKbJm0hcyCNx6q3SUYhRHdiZ9RVGSAk0CfN7joCEEp2pXmBUEBo+YCEebvOnPkBYlgCSsAnvmGw
xjEGhoPXyCNFP6ai23+Mn9MIfhAX93MfvSmqlzQkTXfQl0Tw47Bb/5evFmMpbYGip+ucTh7qMH7m
TPamSfnGGEg89k3Qj8gHLZLS+NLgS6ufqazoD/nSW5wzqv917j6/NQyqQjUi2M9O6fZ0CestkgLD
zSjRVG++Gk4fhuTfQUkip3lyGFzsf+ACMYP9GtxzzB2MeLvbr7vh3wXD6DM9oHCTz8sSzvv2D0Oj
Bx7/4tUP8qw2co4LfNWyPg3WBcKNjH18U4q+M8pMqqUhvLJaWEaVm5YLxoCRMKCdA7W4gvHDpXIG
OvlAuotuQGORnGJqET+0mPwH5HLioK6LifwijXeRCVGxKmigjzwDSlN0+UGoW/yPTuNK6+2bIy/H
FylKXQ6EGQtDmGzzuPCPK5ngVPyQcUxkYOBI140PyJAMm8Q7XBgsxlfzeF+TyU4rxSzNcuV8qwH5
kPV8t8oQvR/nur+IWgQV1SIRvU142B0uGy3ZHU4Hxwen9d5dHu1HG0xeRY61hcWha0oEpKW0pLMI
Zy5cUY1FL/wUmPAU6/z8oc54bK9QE6NqftRBE8g1iFSpz+vtq+HM+Y7uGKAAS5aA280t4iPXGHRp
ol/yyaeCY/a+UJBC3WFoN8YLh9EIWVeO9rA4mM5jqpzNExYl6GZs/flQmoLDPHumps/Qq/Iqxk/4
lIuJw27lvkDnKCjMuWD1bfE9RyJ6PhA80Erw46shfmxMHFH6zdHWVCDSdDp2U36Oz/Egkxkczst4
V+TaqE4/5/DLzXjyfNHuZdJOqdeT6fO41AjtZko+G5qOzjtOIkxY6Stl6zgd5r6xlvFNJDi3Iwre
hVnIQ/U21/A5KBs0VpPlyK9FGCnK2XlkC56nUzbWBYx+LGM0z+DpQKphYHSDQ5Ob92yJe5lDH/bS
WbBUQ1JZ3Bv1Jtg2Ri9Z0qyPTA51BooD2Er+AtuEwoaucOXQxJbnGSubBzIt5+LDu/zV7XCbvZZC
6VAiat2wDPbNfqQy6hrgS3yIfAGvQZwewDCbWfSvWZzFPViRyw8iZGaZ75Vqvp1SxhlwZsf84VY0
XoqJHCmX0BjIHoKlvvcsDeXKUGfcaTuxbeoB/xief9fdhW+fXnPDFlnHGmsU819cj2zomr49l53v
ZkDBkdKl1HONIqXVIPDOL88s/O4rG23Xgjvfvj0JJ5FpXJARTODB85Fewv8mpYKJff/VEvgfpUvS
YmoOu8PMWb3wFfwZo5uEraISPZcIW6D0EQwaTeHgBTmoJQg0L5S7DeeMinZ9xlrNJdi4TKNt4x0E
cK43n28FuD8ioBDItqENxk/eiyZML92zuFTzUUBxeNj9NIpeQcIHX6vTZ4Nlv/y+Vl4Iiib7ca/2
FiGuN/K6dN6JA4pJ4Xsa2IfZ4vsGuN9YvtLD3R6/Ioi+D6ElbNyoSwB5b3EI3nZty4N685lcGC3b
4BQyyGjYtb3a3BWk/ts7R0NiSUzvDJmNJ1oWsXDle0hremFXeHX6lycvgQfheT6ove7ByxqJUWTm
H63agYYiQj/Pha6cVerA5Wz5H6AXGtvEfNEJitN0g/0PQEav6wJpUCo3NK7h151gh2CXuORAvpH4
WIJNj/PW96gtYyUOVH4QCMSEo3fDRi1EfPsDXsRF5aD2YflmzE9acirnGMiUCNdElRQwUSvEK/8H
QvwljLo4fw6BxO/nO8LfXw+XT29qsRvF/63TRboeIl25qOKFlioexImGD/aADuchpa27k9oPc8g4
Z1qDFa5KgWwKBcdPZzkxMRVeffvSw6O3s4e/5aGPWaOPuu+jw1VYS5IcdoXgH0YleBBKPAoYG3pH
0HPkM4ZUy9hXy9940dXkOrhKVly46nTFCVq2mBLym4DVpsRBvAOY3HVdIgDkUm8QpMfxbNAwV8Eo
JZimgYWWa7ENuaAda9TTDEFqmxUttyEh65DkbCr7Cc99OVs9iCzshiVvCutfPi92KflcOVuiB7UQ
OGFKtDoYUiyqYiOi4ceU/qnHLcrtihj6sXc5X78IR8PCLHRnvERfvCfOJzccBpcMA4rOnQVVE+RH
fOnx6gHSRvE8e0ez1shMG/pr288vSE96VEsa6ZOFc8hHcPxSdaSGzsiNuRpYrIbUEPbPRZuY+sns
2Fuwkre2UHDsZKLINK9WGzOrxUYYJQlQxxlMB5WfOCj/ce+FmPrTbZYs6qVrdu6G6qubOjb86lJi
fvdaoUN4ti3sdGpIy6QxKLLRCrnZnq/ySRL7PsACWBAOpQPSNSxExgsnJ4zw9wEDLXpwmadL/QeF
CiezlrAKJFEGKiBuQx7uroo3x0wpdMxkl3x4fmTe3TJ0Odfz08NxdijvWrCTiT6FQkvzkf4oBVUX
aTuEsuiRHdxWFcWQ73+QMM+1JgZLr4H+RpniPliqcLJipdzGmzo/alwYtXYvME+6wD5r2JECmVzl
y41ATfaKT/OxYerAMjfxi8Nj6YgV87oPf6GuwEdqUDaxVFRiR1WUoA41/wdnlRIomRnr4M6hE7IH
lwGPF1CYVTIQe8ntGTfuYUK5rJb6ZWnDca4/H0f171O276blY4OrmBQ2sMeLWU9/udM7T14AH8L5
fpVzKvnWmSS1T+RQzXLCoUobEDHke0MyabjZk9s7zSI6htYUyt8TSCjuux/s0rtxvYAuIoTbtCuu
kAtrZYFHuZYEPpSQlbDvzN9Qrwo7FdPPfIqekl4je8H2umGJ2cLuUGAfIB8iDwa4b3jI+nEiDHWC
7tsR6p0trNbrn05iEE6OW7hene2R5BgrByH7VwLyg2oWrc9EaZph9PwfEIIUj2hnHDZO9SXeq1Nn
1Gj6hUmuZ6E9N/+3oXZjQYA14xnyuAAUfOlMNaZAnajqHOzTwyi+TOT/80ch8LbXFb60dSEWnPxZ
nykvbjn2Ypa4iFqyFE+/qvwzJKUznj2OI+S/ksfQmC2pLLC2rDSLjsoYOtt1I+qtWlQ+lbcBthCa
0qn3S/rAFhrid6dRMjaACH/8dOdW6PPYt6azsGVd3IgTJPD/Qxemmc9NveO6xKLxGQqZJahr0clX
15XE0Owi1MnKL36Oo4eqZOUGZPGXB8JH/Vj41bh8hmMY4OGmw9plvB7qOJpPn+4NgdEh6do8o8L3
IBnjmz0bcMhjlcNs5tXA11Z5dFIpHDKn+9ZuZ2LvjcnWAKJ6zICE7O4i15nglRxOEtg5mnrRMTyO
IVlRpvp7gscVY+UXEwOJJwbZdvDROmDx6RCqGHb/vKqwcx3ZggMvYzIZaE+L/Jb5Ek6pCPEPkpbU
LgEIDZWW91gCJmdQM5xVF6cCZ/aK51uCgHL30jIeCeezmgQIhUmqVkgYq8FFlwp9dtjLF2w6aLRZ
f7F1FS/uHlXuW6CtWVBVWI+prKoMFAjoHOxlfG0dX7QJgHf7M+zM4vj/V9Jn73XZMaDt+cNgG6OX
401frQ9zjGs5CvXtBVhEgV8eKV5OXCh3kdcWrkfjTfXCOuxTXvSW5u4Sh0Mp6Y2LQsIWcoImBMWv
AXd791DP2dgEqFYAEmcdUHuBShzsCrmKzh+o/QLs3vS9afYJsn2FWVat4Stx+y2KKqSg7h7FzHxj
3+3ZLe3pRo0RPn5BnWAz4HQoi0y6vB5vy7ObZvldDh7SMwh9kY2SvN0wN96FSnqYLVuL52yS4SLh
bHO2OMLqQ97/iq7VAXyWjRn4trp4GO645KnwFxenWMIyR3IaG+fOjdvGOxdR0GdfparyQtT7BREh
ZZr0rkikxDqxXWi2JUSdsUxvj5eSR0jhWrxSKI3IyZBa96CnM5jTWoPXnPHbd5inUOR/pt+4OdWb
A0RCo59bgNoRB3OMcH+Ied9dbi7P3uRT1eTK1WfJl7LjE4Y9bF6XqU8hOse0TSaQW7rulWtTro8Y
Yld08eG+HG9QHG8JmI01GelcKnP/hit+gwEX0mKyKQ4DxXdYC70YNkHHIvy7cEohYLHZG0njiVMD
4G22y9tpF6TuYsHv0sbYrnOzpxZjA63N8BYXzn5H7PtA6BvKLAIQL8fOxcF6stIOp1l2K1b7DqNQ
ep2g7owePgy8CtpIc7DiNzmuDmFacwDRphgeMNkXHMw0MMQDeljWH5pHjKPuAyv/PPRDshzkbB68
nRNJ1aNmL76B/qh5gD9E8E6oOuAgYwgLwrKiyBTt/nyU9aFqe5CVyEPTui7t2FpQ93AlbID3O0ZG
u+j+spBCx/+1t4Y/9Bi/IQHW3kg5webpVIVyTNF4YYQH/rZaIjWJuBX/8IenCOH3u4MRbpIYNWlx
aTG3pBjCj0nhaZ6aU8Us0wjql1w+03JWDUyRn/9AzjFD1Ynu4bG8LQeLzubbrDJx50iKRBiq18VF
pFslJlO+wLzkpsMH2l49fLzDAHoN8oaiAFYau5+E2fcWYabusaT0tx2e6DHJWgNiIjJC3+6Mhvao
DX/170QZC3drzrlwFfZmJQEKm0Gk5k9QpT8nD4EQ1NyJucSSMkXVBE1r0bNfzUeAM3M5b5oIUB04
rER5v4TLkXIkSSDiwcDbximky1JgCyjD1DanrfXc+2zUm1gWweq8tc2b8iU9/BHrv5ImLUaGqFoi
gnJekgaaO8Pc2+eDCvo0bGz0bPjciBCKlNPX+L8mtB4BgED5JSCFyM3Jx+zekpkY2pANE0p/0Oyk
aRQUrozL/0/SMVPbYrxAXQUykqyPXuF/i0IeLGszVmbOUXwNYbAYN9+hQMVua4iY92kZm0rfvuKP
q7sGeWuz85894JjbEahGItLsE+5X2G0ZlIpEGhbVHiLqjkwxMecg2/tAwF9EuONXH5YQSM5ocwjG
7pwogOq0xTdyE4rhcrxjyTnAB/rQYfsVR9cXdoS5ZLWhE/YnYmYwwpPsVlXar9y6CKWscLG2UJu/
dNs5fxxsD7bR7Mi0q8u5uu7nVOtxOV9c+3a7LkuYWeEruiU9IVVUhwiB0BvJrOqwBP08/HBBOdrV
DIpJNlRhp2UUAl8vnRgWHI+FXusmkjig5b2PJj4ANW/zjYsYLpG+QteoyoeE/8C29x8gg9bpA8G2
KmN15Fu9/z53sO32+RZGdYzdqdznLABQlOU2/2Qg2YJmG2NJNQcuLN1PNtBX9IJBIiARZy4ZkzSO
ppLCW1gw3s2KWGDF4yshAffed++0cuCpvQP2LY5msosOeUkkjFpJeHvSsxpk6XE8yynablORgybK
oDhUM1R6RN2zMj2DCWDWST3geKHaKKzaV3YYH+Fo3gW4UdvISEx9DuVkNQhn0UssVI9dMWWoS+V7
0lLn/9V50s88UW8a95aWQjfA05Z6GjD56F+gtbmB8JW2DIDBQpfVlQaYSAOb5+iDPF+QKIuDvLOm
hDDv5V/YyFixtVHJqnMUwKC/ohCq/KPJVzYIWR5Q+YIuIz91EOnGyQWnNgorZhy9IZxr4LqgBSce
NLRm+V8hhxXIMUO3vd7shykjmRzzf5TT525CaYGRtJz+3En6tbXzEitxAd3phhzLwTKWDkY37njl
hylgzUw8wUi9u6CgezgiyCQ48e5R05CYjvi0XhKkQJyJy9tocwt/fFkVtzSONowv8e0em1KDHDcC
BYrcNI5Kc6R7z95a8cKA0aLzfcOzwtweG1kr5xkv8dVuj4n2fkO31wB+bqv0uuqtuQyZUuVW3uNJ
/QHsycrhB00WZL7ZdI+YSYmBdgajm/N7S1VbSWDj+yMe1QjGQLd11A3SJLiymd+fTB/z84lTu2xw
a5QJ2UbabC7pfDLPXVtrmKWkN55LANEj2izUag9ePZ+ihImUiaUMOt73joQC8TnC/KjQOdLrbJ7x
Rh6+lBnmkcsAfp5ykVfCXI4mJ41VxlcYNDsG9FEJbVoneiVRRBc3XBrZINgeL7gG6yoIM1D84wv2
wHN1Jl5jv14+9Z3GymGOTDdqyTYYYAnxpTaQuz2/gXTo0JxCqWWS1XRvXW+Hf31QR5oyaoKxDvJt
1pHT4LKalBfbiQpHoFOUauwlTO2ssRl2XxNIsZWXhz2NQTC7B9j2QvDdNsIHPdxuUZ7dAst03/3d
jqD1q7A2uW5ISo68zMfmBwtEJbcbOcJJOrI8TZy8VeCNajBqoe92WrRPppg6s7aT87eiDu28gZAk
hkJjTD5pgDtYVw8h2I9Vg6+OAdjNBbxCtu4s9XK1yoN0CuxxNyt87ai/zpVeeCCYDZLV0Xk9AQ3C
AafPGhPkujDxys4DwQlxmZSmm7VsRe06XVBTSYM+v+PpDOq38AW/qVF2GxG4JVZ7svMOvALD02bx
spymkMz1w94JhvA/8N52najK8qkC+PQziKxHDSHcifaEUldcFBTxTlfPzABmWNHiBYXPiEFy60T3
/g+twg/lkkLCfYrCpn5tcWYDSwU4dPNx56tIkMnm6BVP23SUd0IGa4JtIZeulKXrSRfimLH2Exqp
P5wbBTuc6+uQQ7O906RCeVFy1kDsT48C9GLkPJvl1RBGyvWAvBM6pUc2bgcKLBK16EeJQBr5CN07
MhON8IXstaH1I86yMUkD1GYczvzfzuVIxzJSsREl0RzwGbZTQOWyauNWfAuLs66cbJE13sDKoR0v
ANxWZ/9XtJrshXhlhxspFCExr5tPssfKF6tb6QXGYGrdrgx9eJqjfDTAtq2EW3wSwfGDIA/sJldA
00xwmM+AuVZ4b6KeXm1ZEGgtpRfGbqKk4svRgNOgeC+ZW+4BgHr9WtGcRb21SOVs7IwW7p0B8OhX
MRM/l7JKFavqm/bME4jw0kzGFL7w0sfvjsHt0hEpvKXK1lKkUWUl38rKdn94NKyUTJyVedMXaMRo
DmkWRK7QNLzLUt0nvutnh1/b+vPha2WxMRIGh4OLwnezo5Ur0UEa6CPy0XE9XyD6b7UnJF1Ynojv
8WGNXJLYST8TtIJtFh1fjZfL/ZZXe0ie/GDDQSnJ5v7xqeaLedaRI/yhtXWxn564NMZYlg3NUD7K
BX8Wd7u16NcGaq2q4gJB4aahSuT0pNzntjB1a1o9pMuYD7T7Qx74MVYvgqAmUODzbT4TLcVVCwCC
/49RoRZHolU9Bu93MbUXnbK7TJyJMB9FmfrGj2MHXbkSP26unsmzx+cxePUi0/4LeItZLCDLvh7u
bci6CDJbGu04BPuRSuF7gBYuInIXU6Z44Skd9PjkCOo/7RNTg4fvQkihocKOkvS51Bu2BmUo7/dE
aRhXAnA+TDEbYVuHW7hlQRfTgmONIR5JGnDOFGrsbjUTBZITMF9rACKRq8hAXau0XlFcvn19unNT
5nu+miJ841dcS+xZvJP9QZEbw4jbMlOMjF6pUILhtHPmdjEobdur1NUkLrtR3LHiwSvgyJM+QF0h
hN7N+/zY13qGEn6kRY9PoBXkovH/ZTQorlDIAcKjfLI+pFxOSopUhsGQaACxjz5UNR16GIWcMeVy
jAGokhg/MgxwbOArvKJHCnsHd0F6m2eai7j+aB0aZJWBu2KXPhrz7nfIJYEt4RrkgkpZVbUs727R
uhCKQ/3zeyZzPzgoNaiuMS65WtjhltEpGU8g+laZdcE5uTH5O0gSIV5dKbHZKsdwMXzcLqa+ArRK
p7UDfPeHDun0zYPnlFUcdv53ksxdSd+1AvMwvB1Nl/DFSWsVsR/d5TJkyCO5QZROWuESb2eHaCuU
ejesGZ4eo1T1Dj+/evam2/O3nroqj/T8qtrUuHY1p0k/nDH6l6BBpnIPvJ8hpPS26wN1QDaY4kw7
3cvblwR072sBYiU3LFVIqGiGTEpDRyN8nm3XgmT+dMcmm2zO2rZDYKu1XZ+LK+3zDhAhPwh/r2LS
nfelNi4CnJF1VkxqvzL8bKdXJOUuw0Sm0cjihsqqWl4+DqC+jiqxiW209jnEbeQtPbF9kl8LAal3
nPnOUOe4OQVl6kBOLrXKN0zW5capwXIk7Tw0PJIN5e5GzS3cbI+FuCJgFUzEsBi+owKg64ZB07Rf
cq1RC4eh97mM+sKzzQ5kCS/XaCxS+BBhhE90QlCZJ5RJqeZgYpsvp3pyP0tc97r1crkJJbDwZEkY
QpDWQnklqlIzFfY3B6DMYXe6c1yRoymkFxbqcVLowNGoQFlypGCtqH89vPjOcK410i/PullPnOdf
Bf/ZEdknIdBkGCjdjYVHp7MunN/RTn+JGDZLPuJATyaG51aoIGfvA4ZIxSCfvZqkRbgGJvynx0U5
ZCfu/JXVMNDYLvqWcKdg7wRd0ZCagya0fOx2uww8GRVj6gnX3FvCi+OP43GmScaEejTFjI/KNbag
qoikKPq0T1D3Q2VAXhzCkgGa1WJ0mf3+FRX8IyXtyUeb3JA69UXWwkwlwiRNqK1ww9CHEkN7VUrt
DSEPHk7x5QUAKluHy++xJZ8hggCj9QO9w5tWBx6xKUvoyq96UlAYGC9JUmoh3RQySYIlu6Y/C/W/
9LlbR6yXbb9fl+cqgHBIO7PjGekKEyGoMTbBmKKrFqKMMNhP4/hdwIEH+eHc5WyKTSP+2g64nLon
lv3zmVNqsGPXRgtd0tgWF1UzxbIfjhIt9Pl7BoeElVt9Pt0HM4cUZqY3LQoT/ebJBtFFQD0l0ZJU
snGXuuFkR4BnZNA6wJSlGru40cpj++It5UHJAbjVnk0xYjjbCLWmWPk3Sj+KcSQ+DZ+Ss05/0JVc
FCu8bJjDt2BN9H2R5YtlS3+3efM0hlxKFGBZvuS3TaYkigrBSb/Pv4Cj//ZaWOQsUrlAW5DeFjYe
BwXtFyFQpKXsNTCJPP36tBUjMPrnxWXwl5AoSlKIw2KrAidCaJYowdGw98qmBHrzEAa/M2cqN32w
PKLH4c+GRCq9sKNGyZ2i1kCMYoAhO26pZbmbw+N8seK23peQ+tNC9QyUev9Kd6iAsBTELGqtr98A
EBj2401UySJ2Hw5e7lnTJ1qY3fRXLxq4fXohhjMnbUJqihj5XeRVbbTxvIvBYUJmGD/hQPnzEKeI
hTxp8b9Rp3vI1fr/WJKibxkzyyUme2dUGBAAXc2DIMOP5qTklGYVLNAdeZltGvvTyB482JJr+qNu
mwSaX4U81dyiCDN8OioMh/3H/b6tDTKJKicVt8g3Uc5MgcqVfASDMMv8n8mfi7im/Hk1felrnrDf
r4ryXqtW2q2/hQtVpmEi5RsQCB7sgeiO7vzqx0zhjZ7/RX3iBakxNGmXiRuZPUbHbqlj3Pf7s98p
KfHKSwtitNZRsa3H6pzQ/aixq3OTH6s1rMxueb5SKMztyprZlc6fbGyIHUB+0VoLilUBkdEIvvlc
H/srwrmcQgTxfDHDFzvDvBsrGFE3NHHrdthKpQxr5S0i7j4VVDEub7P2zc9HGjiD7h6swzt7OmeO
wFBjZQlZgQxtGVj0WP8weKS4/kKBu9IoVAPCHPPt9vXtNbyvms122Ix/+SItpcIdBC0z5J8ggBQ2
ikrRWkh4GT3NbLwl6o08GBXfALAmlQrirM97mEi2o9xF0iTsANajZgFFkNZBLc3OEyV9zJQNlDx/
942i/QRvYG/Yatmg4/bPNFvoRn/DcmCVxcCiu2V2YlUTVaoMnWW+vzdFUckAo/KIW+7SemlR3cPH
j3c2zBzpmFcI3n+itCS/dA4tyzr06b82cFCiT6NR3GXV9bRWcrTirxNR5w4R9d0vtzPoBbYSVkT2
xdZGeKp+up02wC3SdAr7LJiBv67ZTKS179C/eaafX8VDEwHcES8YbNeWvPGdpjkkPld31/gQbwPX
xNNirtbZqMvWBVcoIBwksqigdJENNui/RjwnXGZKTC6dejs+I2f4eYsXNKbCzyB1yg6TwfgP+ZdE
MWu0Qcmewrafst6iNRZRVWlM626Gxn8ESatB+vl+P3KOtVkIy1rlgVEwavthAyYKnNPEW5QTpKQa
+5iMjEolr/KmXHx7eAM+t+k1eGJ+n13O4jNLIPFtLnXaSrAQYxdUvhCGE7Q+VmrAc6q0hBcGa8QR
noXIhwgFY4TsizWVir7BJcDJXZpLv8zShpfxEJSbWIHXHRq0PQSXL/m22RxDsyJbtArTKXHS1ZGx
bxDXjQZXCoy4cD9qFKHSLxAN6bvdSUNCPUhIX+lX+qC8ABEnqmTsGwBUAJF8m1FcENa6fVXLU4/Q
zaoX2n1gZj8TyR+9nCs+L3Qyrcju23rT7x9xO4DiRxokj+tZTBUJ5AF3UdesgvNU327RYXOlvsX9
MG1HzZjHrUoo94h/G70H859IxTUGjTVPK1H/3YDTQvwHIjR4l14TkV4881Eid/idqnmjzxO5yNlg
EkFvlKMchEp93xdsqG3qZXaQ3olqTKJmM0txTeJOu8tLPAvW7Au4z6mfYoSb7gtAnOH5mpq4a+Y+
OGOpnj4ctI2Peub/+BBpPY50pCcUc8EGhgDBINLyS1FQ6YgkUfGJCGwiH97o+Fuf81do7Zucasrr
9WEslE7M8jmogvol1cZaOvbmNT/wHrXiNQjijpSLeh/g0gUoGq0CqUb64k/dpE59DoClOdw4K5xm
M27++criEpI3tPEnJZ4NK1sJT4oR1R05PZ2k3XW7k0MJpY6FjmeGmvQzFN+wQ/I4Sms1rOSyVl/2
r8MTDKZ21UYZtA7JAiVD1VZxc+iQyCz3sVqJ4n0it14K+B+hhfPhGspeFmoqIgXzWiYdxX2bCa9K
aySLwwE2MADUo3pwB+z3+m1+yp/8bfcCPYoD2SA7ri1Ebfy9TL/CZpImRE3IY0XKi7BOe/Q0drWy
1+28lseItJAQjMsdbIuDv1BL93VZbyvxChTAx0oIRjhWXOiZ9K2iAK8qv7fkZ7vfzOqUSvESkbP1
a81WtPbUPJ20odef96bsYXAzPjNs/nPb0zGlmlddCW9RyfLfcJ8++cKnF3u03KTaseKf0cxyShvO
ptXbe7dWzDZaBl41qLzHGAdTh+xCaPcq3UmfsmevYKambinHbqimRBDsPcwetknQmbTHEQq1oOUQ
xy8GLFPFhJp98j7afiyehx8t2vwDKM9qJN0TMevdlr33MA2EYVCIbpp8mXxSNm0oFq7NYzFqQ/TY
0kSFv/lWTVVD9FEAh71OqVVC6PAxU65iyeCa8AxcZESqdS/H8bJmOeck3lbW2+I0FQmAn7qX9v15
l7C92WqJ0xieZDr2w3AoAaOU7zPQ3LwGCOkE6yLkunMax6oRpf5YVLidHOeXD2VMPqPoLCEP7yXT
xsi7b3/MevQ2IA21bLOHV9WYaHxJWCJbI5Kdt+oBWaO0b1bHNM4q+8B1fwV/7nLbDz2nEemNvzkB
MT6OWrNze2O2NnmwrZ9aJxzlXKsemMMOdhENP9sgqiqTHHow/TdN0ml9JLVrpp8k4KfyCAlxIlsh
EUlxrrRYjPPkQSwcsaaNQwQ0ifFKFX1eGAkR2skAvRdM4Z6YbJA80ibomQRrX6UrEKVknPhByBEx
zhZnO7kGWdBjRpPLb0N8acsvBqfsuCWDOOpJcs32wKSJavVW+8gmDZ5MAwWH7y4eARJ8reuz8ffv
bX4k+9IaRNLfeiHuPgWvWM9HbRhu7Ff2YwpmcWaJgvCMg4NWruhKm+EggtDkjToLIjYuz3aD3U8w
XXncF+uumdr7X1gCJYWwnSSug8q4MaKcfwd95g3Ebh+GeCTAGnK7dor+8AkYYDzDj6FvmSfB658T
wUH5p+3Od9ELav10AXshSCFuP5kaRLvme6/kPTRjOc3vzFU3qb8v15oPn4CcNavl443mrDGiAV1m
6VGNU++0D0u+X7dr4x4YDFDJ8PNgopTwzRtDQ9cbMOup5zZeTxyfXxqZ+wsOTcLdF6A0Y+EMcen8
UnCzYki6m66XxCi/TLpwpVFVy8b+jk1QPOzb93GToDxqaoFcl3eJpf07Dv65d7JOlWfys/qZT7io
6S1fgBlzBFz6YPKTueZx7T1Xwp4w1rsD5xS7udJxGOd/6c95a67509YNSqBFTL/W+7iwc1/5uTZW
oeWVRYH5E2Y+vH9jfY0GWs2urQrsUOh4apy1N6t7X4kEydwUgn5khXGC/kpEYTH9eQnFbU2FE9ZC
3JuumjY+NCWiVteWON0hHYmWqMIdfYoM+ymW0Qi+0c1t38tBrSP+iSXSoCGV+9pWV8UW99l3/WLH
QiWOuL+7FbQAkPX8r/gO64dyqQsuohDwRCSqpFpQX09gUy96FRp5cCxr6uu0v95Vw4DJDdLoWM77
sgnrtR10V/jYRb36QNryqwPlj4HzLKmbOpxSdvHOF3x9PcdhUUIAey+L4cLoor4eG+8FDSqZgDfu
LBfQtNmmfaL64fEzb7A+ypjrg843FqBbP6FEsbdPO3mrh80nSZvGpv8tNf67CNHCAtdADOKeCUMa
1aYLeCT71faMZJfcJ+dAywIdTOvnk9uuIeohpcC5hyhXShsg8+d6a8cgRaYmUNSTXrYGpHJbmxZT
Mx68J4e/6Q8RkIoDvdRaUdAFPiOSWG6XRQyRCm7zKP116uT5ukXJmkie/H4r2OI8HezDWdBj4Ee+
r8xy468HDH8aEFAx69gtXGziSXtwSp2pVtWSIgLhWzBsHXpvUsqChpzOvBOsZZkAJGSn+JjNGL2m
PTgubuyXpt8r0FrLSgUKGTNLb6Tplpu2wb3OggfNByyNzF+VTzS+dIILauOTEriRR5QdwlH0xdYF
RCmsU/5XdYYaGFzBbDMciXtOEt+emoqcSWEjfc5rrJBNq3r5TjR+oChvfM1lDrDNqp9+YteaCgDF
972CrJCLwxzAI2XLcyd1ADyqG4dRk5J3c0vCjFuHurC8joZj05rc/MuLDTIaY2Yjz4RQrjxSs1it
qyM4yMeLudPSlUUD5oeGmzjPENSgvWq0YPvfRYBA8T54+NU7QFsX1IX1J5nhkENSK4rbLr8mwRMB
gcKmYXNf4b7b7LkFx0p3JD7B3jJxlQGrEu6PiphB1Far7VfIuEk+jiCGiJA+KULelv0OFQ3xcZqF
bHThBjAKt8Ruzs/DufqdbtmDRa+ztHxo2voO3oBuxIgJ97Dd/G57lF9Ib+9M/+e8b7WEJk8PGXnz
vdAloZ17VSUlqG4c3yGXu4T+tC+eOvtcHXfrpa791m6cvKEPnEY8WEhKRhX2JtaonZewqjlLZ4iT
4Td8I/I5lBsJdnA2RRSE7/FM5xiDvmTOTmxgLEXrGzNwTXyH/h0Bynn5BLE/pPasTPLpfO4gvcgL
S5W6RcG6WWWcG6ob1blMzPNVMqOAwZv+y9JKP/lK3q5GdSzi75OGMO2fsfz8vPcu+75NsW3zHSZg
6oU6OtYL/WFZQp3QcpyjM7AD3DIZuYrzDU93NgjkUG3kzN+lSzd+UqzoEujkmZ5zYnAmeOZThy+E
MaUKv3qh7RjjYFX4glyM/BiBmJuhhDOVIaqZL3oAWm3J6PJiszVww8XpdVU5wjMIPZvFolS1EmzZ
GMlG2oQEgzplVCdx6974PS2+OsQzkzqX+OkqnLL6GRvXOPBz+Fg/OJNNEghVvFMw9C1WW49lHJhI
qFPfQ4itKgm70P6vJmuU/kyScXI8rm8CFGV5IopIHfYq7JyAQzrLRw3ePK61XwZEDq4tfng6XG/t
K6ItTpZJ5z6IJavJ6StQO1xan8HKqyzDrP6gGBVW6NPjXpJGMW2AnX2NOyNwEtK3Ltg6/9OtdwE9
IgsNafJ00tyEBO3cfra+kn5zbyvcF8UNtSsJl0xZOBP26KBR89dy2b/uf01duI+UbRQ+RXwFJa6S
UL5FUF4gIBSCOCYQs+NxNdyc775Y/cOFPcilSjG8t/g5//kVPtAWAVPcL2PxNdGnpM4GVhjlveFM
srSB1JJB0hfjsKx4ZJTlyOvipimCLjbblKaCH7jcMR9jd+GTSqykWc1/qrwh9MU21PPe4qgJS745
ecHGykGTcg2K2RmJWIm2hA5IPBpjUN9lCZBgY6SQjPKLxMrC8qObPJ49lDCCrC3QzQqvnfJA0sGk
SgIO8RAvKBi+rCsvzE+RRGH/QuB1WJ/a/vBymBJxnetd4VzJ8JWi0KlU0wK2xS4SRsutZB4YoVxh
AJ5tsY51YzMiZc2Ozl8ht7h2pmapvhFMjGLZ5AQkXKdx9QWsTQiMkj199Amliwf8jUKoUg38K9zx
ayuUGUZK6zl8VTr+FbYQQnwOWoxKtB24h2G1IcuQy0POLUIWYHt+gaqqdvVLW8hV4o8vlRocKU6V
tCc6fmkstOEsMX4kzys9sp7CeLJ/UdnX4cx2QrqNDl4nSXevVc8g6ujdZRLkTs3vftUsdOQlIynk
AgCfe9ETtHqdEINvQYQOGU/CHNTCP4AmuWLIPpeZ39zwsj7xpvky244zyiwp6Ih4L5BuBesQDxMW
N+wg1kkT1KbvrD4DA8t1a/YSPIJLegDb6P5EJqJ0aelZwu/yXclRivq5Tq5kK1ND3gbZQyqLhhOA
whO3jNTlG2S3jQQiSUg9gFNL6IcWcHfD5MuKPO03uFUVb13YxB+rGb1Yr6WMQN21lPOYZyCig3wt
/HF4Hu2QU7Mb6783WgWFXQUzFRuLZoyyXAGjYQCirnz5Kj8KiHl51udoUkfpGhGuJMmUZJN/F7F/
3GHcexfQzQb5feJIHOywYtC4pfyRB5QsdN4HGwpdg8dpoK19aNWFOoeX7bkV7uyu65uO+kFX7hJx
eyf+iRHOhJVZivFIoeYUCLFGMf3slOTClqNm9I/1EKZdEMcZhL00lKseMimWKo5cK7BcTXwwb3L+
84BK7pCXhOI1vlmZWjYbbhZibjzGE8DsbO3v3qHCbDQJsgJgvE3mk+47BOiAJszz90iI0JmRIUax
ZFSWycbjHGF5kp+iILzBHiyDpN7l+DIhCSxmUAn9d0/Jb1TnpYuiCXKjz81qAFK3TZ3ebHht7wPk
aueF3LfMMIDpFODv/g3oL9/3MHQT9lkDdFTb8kSKQZmlBugQyrc01q0KyPRnNa9JeadkKb0oxN9R
2dJox+VIKVblEXU4kCdYw52cJrGVUzENcjKiQCLfrGUfo/v//PhxUj7r16iLMGqENITcXfv8oOTc
mKV4nP5pq10UklbNqck78SP5m1kp79pFXk8jJ1y10ENOjl0LvsEyt/KZH46USPE/X0ePXSFoK2D/
9BKii5KpHOjleq9tAXrptdB5REd66pKHl5+U27nZm1XSzhYAtMsWJ/ZSfSmN/iZl3gW+28ELoywx
RVrnW1aDRIjo78m+Sb9104mLBcwZJmDWqW7mfOsxnkbLljp6fYSrjT4U4VAlkBdr0ty4Atir4Htu
bQfhI8Q9ZQi4cOSD2dH4X59apumitoa9kwWJ5cvPQz223IyYmkb3IUjsCcfz7coCB42kPPTEOQAR
uS5GGPc287cGUayW2OhQ94B7K4jzsbris9B6G+oHm8ThJMpXQlofik1H1S/Kz7x4y3qTwiw9ziBE
9Poui3tarAeSPmhZ/c6xkWg5DMGobEaFww5pKdBhE9qLmQCDrTaXUA8afWP767mzd4wEPfejXkXx
j+37OBWIz1MtIybGPr4EuYn9821A25KFrSXnSm0uMzWvIqeUag+2pLsPa0L+MarQj76ebwF3rl7K
uvvo1E89OfgrdAERsd/6Qp/VdgzwPiD3wjroWe3cvh4rwNOxwldou6kdzSqBNkY1Rci5su4E4JRO
1+aRfOG69NRtw9WmPZXscPE/nKlIWyFclMYcD3E+0CWGwB/2oZeiJxXkXzY5t40nA2GHzpVRlSSx
i4VKcjd6nmQ3Km/ZxHJ6yK9q2TiJXqqH5Vhf8oXI5BuZ52cKR6QYORNjRNpETo4OY0Y36x8ph/K0
BNfslllJgZ4GvBe6VE23ckNEZjH/I5mXprVDzEbEhb/FpevfcF+QrZQ/tvotezTu+4iZ7llmpbUi
gaccYdkD3KcUgDtD6NcQblNT95Joo3qgJ4UA5+gZ3JeIgsGY908poQIexfJ84Jcg4N1Zko1ygK+q
+Z2bn8NnuJfxShOLJCYLJiEmIaP7OnSX953bOU0P5yqQ0YavDzS3C/thK0wkUWyN1mkZ2KUGnKtu
iFiKz+1IWz6YTVGzuAy+uKbeu57FbPKIw7nGtJ2UiUxdajseqW+3m7LUMBjuqYn7q0WpSoxabVRw
2CF3t18Io4Z3sBrOBYtB6zpTs37SXPD5EWsiLpNc4Hn5Z8zzUrEKphzUXvLZAGq7bcNop4rjpDYA
ldxNzxtjxW/4Cs9I3lX3jgeWzXd7RscTm0EVVEOW5fmjYuuQd8Ng0eCyBAdsN6nOIpRTEtZihyy0
rQFHPl9OTVDf5RBcaXti6S7XtClN0Tme/prVc8AFDGtU0HwydDdXRIzUf5Iur/F3ZXOPPdghohjU
x/WDS2POilaxC+bvrt10NaED48nVLbAegXbuGug8mjrvpE0cBTqOIm7xd88G9tFfTQwEh2lIT0+1
4Q5BtgPaxvsWnMuEw5FDbenwSLkHHto7Xpgary7UFvZU53+pFRcmnLGOmvwR/lkHfmR/Q1PFSrqG
P5+r1q+kWtShl67ntZ2wqLsRJuQGHHy5WnUtSMe/Ep1TZXGw85+ZNHGQ/C86ksWLZRCc2dGOsE7E
Fo3RP93qyJL8Wru9A1mAph7jMojlNgk7YSg5tZKBbL9yCO+LLpHWM1JaioY92IkxR13ji5l7Nc35
th49EM50KGg+f38Nmmbn7jpiPPkvrEYPLy91VZZfwkUGDfc8rwjIvVf73maFaXp+TiUi/8HBGKvK
9GANeGAgB5oKSovAmk6qiJ9vl4TPSoxP2AFMxTl2GbN1PJs63Ue99hKsUKbh8YeiBhALF1azuu9Z
8pVn7o4e2hxu0Lg+dhcvqkuWpYGo+pnd306h50cm9BB8kFKSb/99/DpxlFyeAkZkWWBcqiA9Mti6
m0UVnCTKlav1ACISMqX8fvLL/xxB2bvdRk6ueGhTqq+CaDATMWcc9iwrnb1KW7tmdy/fm/v6xJEF
bCZxpXzFrJ7QpWKBN2vSP7IoLe8OjzaKTD02wLNOPsb9LrgdHzsgV5eNZ+8rcWgLOaMMGzHWhMFB
g4brSTmr80M+pEry1F9hhL3at+yi/LF7JWg0czk4uWjoVQrdn0NwZapDg2qSegc1DAI/b8Mmm0aw
52wA6vlIk+P2UguAs9wC2/FKC2IhvbAkNYFf6KCNEPQILLUAg4y/dJMDVagaxuwKWhCgZ1+uD84G
lc3tzbnNh7x9lVcchzsycriNmTkBfWT6Njtyjha9b0CF3IGpjFLLzV9qeWab1mmIpmY4XP3vu/Pd
6F88vnOpVfJ/p974B5J9s6bZvXDr5XKDU5pbWNBruLF7+oZ3C1raOBZs9Aq+qm/CClixhmHVgZg0
IaTPJn3kWP0CWaBNvYs72fEqnEAMa6BAjeBf5Ih3iM4er+H9StMo6hxsvbfobp2iDo1ndwNMDb1G
p3D7k3SdJ0qvcYx92pB5LgQD8VWqMzMqFqjjHprO5TX1Nn7SD3NFCFw+NPao+65IO04Jh+ueL4ts
JdXk3Xo6oqfkIHYef7jfuuNOqm7UPohUxKsdOOSfaO9y9Av/7htw9mt32n7kBLmqHbTt1Cwg+af1
mU6Ln4HIcZSM5t5wK41ZRKpVvjuiAbnhrWmdkefNVbqRXSPXgQPUzfeFf+2h55rplzydMPodJmqU
9SY55G58s4z4c1Ww5JyTvXaxtyRCfubCVLJTQpazxpO55ruS+GMN+RAp6/xxlgYYxQKttmH5KBvF
haxdyxja2EOCJXdqhlbrM8sIt51dsdx1jfUGuofnRJBn2qkhUTXr7/UBzM/kwCBe62sbPp6znnQO
TeARPHQ22yhAaSnu4LpUDo8pNcEc2QfzeZg+GtgEuhs/04cnbtlfdJsabAIrpeUIZjccWwcOfDd+
arCLh3E+p4z2mgMpDHQre2XvnJscehGuQBi97Tirhh/wHWJ5E635eJw+/Mll0HaRpE1roqeN0GPf
R1TENqgaLgK8dEe412L1dVG2oTEHyCyuvZ/v5aNH4NjDlktNiKLcQugt4382T6e7d3Hr9pWXw0Z4
Tq5lUn2yMXPOEqAb4DlaVFs3Tu9CXgRuAq7CVFC4XXfCI9+5wbWRuBa2rL4P/HrksNTNbq4Eezpz
ZHCSbaSVwRBLwoNsOIMEiZoPPBao6xu3Zn0mY/E5Or1dNJmDVDbhvUiMssaAjgdl4sC6nwgC3Nzn
yBznzHwZgVSU5rRLx4e/CvbjiZR/9LHUDDWwDEtOS8Yw0iY3QgcbsUxzMbdzvVZ0ePWsNsQlRUch
WEUqK2TFhy9XHA7iChStB0LReSbynV7hJp0U7i57FlMa157V8rBcSFYXvaoR212jsscrLtX38reh
AWED4kfqRmBj674/NOmrChBcAPwp1g9GIwoQiN/tECAEkVvPpuq8ItzyQ4qVMAnqKWEtvYdCU/N0
hCy1NVtgBoCP8BkjJvVRTkMJ5mIoxXpZ6fIIqSeoDQqTJ74RQ3Njd+akk7n+Gv0sr4bbWhVzTxLi
BxQHpnsPLQF7YJ29n2L/NXs1okQ7gl7hrXAquT87aWenfDjbvHwIk45HLpIhcx0v/w4Y80sdtvfC
fNn+RELPMk3zABqsDIcTCGX4OkTdJSLldlahoQX+4jBayPn+U1YF6tIMUnqudMY6Lx8CJ5pjRkSS
nIoNnLToIiDshNAo3/7B9mvQLKlfMU6UT9R+4bplYue+mxEZoqbJ/uuqXforIgt7e345NEhEJCkP
Ofp4zD44cFUMIP3oacNJlAQcRr/ssEDZ49NE9z4HpOhCJGtARphdu3G+bk+Q7eAgOb2cuFbmmDWJ
UkHgsB8/4MT12bvgD8mT32r2yLCLa3QwWZL30082DO7l/L5jEapMlf4AHJ+fPJj6lN/qOOKX7Tpy
mbdDO6lOL2yhAnDJ+Tp3aKlqj/m5aef/kKamVSl8QzuSAYzNjjWrAw5M1bvkEHiUQSLyYZ8QihYb
lM/lBB4fdbCEbif2B+LNmihZdN5wx7ls3SXmJVhww3YqIJt5KY1tTJfKZ/TrIq1aj0Yr2pBoya/4
oKoYzcNX7SOG85mB0+T8JnJaaJVEQ6pWXH9fDgRDCK9yMlMBOeXGt/LONbxWmiJCJkYE2KdvTcZu
rTKCTjnvF+dacjLOYskODi/JMXu9UTxTSvGKv9GHvHr/bryUPN0oYE8rI/vUpSZcaN+F16rnLK0V
Kt/pQFZBeAZrZIgXD3wMS8ZPLC6V79ZHC3fvPsfOyCUJPHTR7NsDEPxiHjpJzXWZIQSKwGUeIx62
IAH0GSxLt08G9ferusAoPyrMBJ0J6R/e0di1gYtV4GyN95l5CML2rjVkqZs2HRhTGkjpVexcOhGr
gJ9DIXPJqMwdttjLlIgHbBawguMeMfm4/5jc1s75//kcR+2/dRPIEFwfvPUnbosmgbeXT+YvHqZ/
hIk+57kfqWMlIcPvk8tZu/kX4N9o2c6N/g2ovnIpooefdxddF49sHcfe7GHd2PvH9I+68t2C+vAY
0Gj507ZhrlT27Yz11+ysvUX044h8NYSCTgORHWGKCLN5NpBDU2CTXiVTZH3VSSpn4RKgDLZcYiLj
RSzIJNY6ZwGBRHGIU692czRVcslECc52ESOaebHF3OJVSzEQWPeCBydpXJySP7qg96v+WkRaybbP
NqZV6WLE6LibAfVOPM2cxz2gfLND6w507kXK3GldTzm4CltTHBtJX+LPFbNkY2niReFsTBnjgnmm
jZcygvbu4zw96lo+4bdQKVGQPj+GN7D2Y2MRS+f3v/Nf2jEpER157fjUPjjoA26429xdEjJ6legZ
91bJ1mofQo8ptPKvML5bahmQu8Rr1m7iHG6TlsRroTIVKx1ajsnFwrcDVqP1MxUgu1GzMelcTV8a
l2x/P8E6/+izw25iYiHwkvvmk0RGZACt9Vyn0e2jWRNNojXWu/jyC+Ahhx8MdP1Lx7mRHVoxs/AD
XVyg/q9BTUVSyrvkCMLF7ZTJ/OqVmTGUfoZESNH0DYMUYcC9Xa7fQGOxYuqC55YUc4AILq278lhX
DwM9ZuSYO4bOviPNtVdzzPRLd16a8afJm3K9k8HaN81me22Ho+7wG8CDYjepLc6MjKQqFE+JA5J8
jxhRJ1YGCGCmCq6oZPyqvjlCDjQIIC71wFvJ9dVc6PHksDOjREx20p7tf3q5ga3MoeKinChNSaJW
qOitm9H+lEQlr0rrzyfOUlDCos78Z8ltpVpKHU3ZYGbh4XR9YK4bZjbzWFmmiMvDLwS+jVfvrOFE
e+fCJugJYsY0dMElhEHY1FzGC4tACwwyTf9n/H9yFDKLK+3AUpSBlG/LwF2g6m/Ol+NqX62Ud9pk
RhuqjwbaK2r5y0kJcT8+54lOh5/KyW8Qja4lQK2uwaiLwW7B5sstR2hq9fsYY5DfwZ3sPQuYS3+P
VM3RNA+snnC36QSJvBRT90RQQmHOQN8FQmG00uXnnlpnOqiEhXHuSFUkmghWxZB+kDpWd4OgSAh4
wNhS+4bO1Yb2aR7bIbea3offyBShKH4zMd0N6DukSf4d+3rv50YsdEesgWxdX7t22KItfB3kXEJG
ZCsd0wnqAXao36FMyz5jUecNVrKYYqArN6UEbygCFaCa35BCHSOpTDDHzrB5rgdnowK7GCthCLPa
Truu/dGtL4O046Cjxx7iQJKWBVudQs7oOCjc1syOAm+pLGqckwZbF8Ml1Kg0YEvdBc22FMttkG2U
ml63mPfMTf7jcSK9oQAo8i3nSqgpD0wzrJ5b/1GTtmIXkqP3M24DxTifleV1oN8CURhB736A/H3q
gvBFT8iQRSd1mfxmybLYjSGXSyQ1Tl//l16uzD5/YpNMH3YpzWjeqTnukCdXQfyqAN6DsM4DU9wf
SdOqc83ozVFtvnDzU/avZ1GF+cMYbTAJTQ3rI/MBu/F3zdrxR924du9HneeZFk1xLy1dXEyfpznl
AnV6PAyrCY+7jfpyd7URr+BMRUBaphYjlqO9xNYr95jkT/I5LfpIgPH8+cgPGcyLIUnG5w+/0jIF
ZhwTRMRrN7+WAVs5yS7mevikqlgC+qZ/70VVPKUyEH6+Pwt8wWhE0QHfv6CA1fEJQFik47Utew3G
I+gUTlUoG5Msa4LcY1LRq+tRlNgcGVeYMsuB8AH1zNWBQO2ugCBYPywOZoL8w7nxstYtg691N0CE
GsYiuOHvHEUVIgpF0HTg1iy6bJuZ7/OQdaqxMnzZgTuKrBtf0fioW6qguCQo1ErXcDDbyyCx7Qpv
Nvv3MyYPKu1VhwmpsXpTZz9v6j21dOyW9gio5olXA1mOH1bIbAafv9v6OTR/R+Fj+vICVuLWhnwc
008lCFdYCjku0CmDHwafpPF8ntOoZm+0gjZvX/nGShE00/2+QpvDp7D97yT9vyd2whFle4pDONBn
KTOk/HordRkhUCGrQrCJbRjYwiSBo/d7203EgVsSXwEsOH0rpOY3V6QzyVEcuDvYzyoVIARBpQj5
XK/qVSVKrfdGry5qV9USvL1HX1HMez1dizUOOSDmX6VFbxF4DohoMoYRtkMhTG6Go5KYI7OTuRuj
Fp4tWM+4ag/QOicYvjusIL0yQFGrTV3bZI8Q/Q11GkHGE4Dg7We7+WcB5PdFchTwMwzUkVdrMEHl
km5lNJwHhZexcNMU5fpezKmA4U2k7Jb2AtwHhwSJ13yKi0vTjh63KWQcj50j0pT24OCClv9tzhll
f+leL75e57eAX1qnrBokZjbxfa5KdNV7Yab7DV7bhkNvNbwQXLhmWCRxlMkhuY55OzkvgpduPzVT
rmLFp4nl1VWSpO+Sxp4a/1tBGmCsgiS0/b1+1eMaS2uuFJV1cvzPGbz4BGGAxyM6DWBXr0F9oo3r
ANZ4VYrsJFo1/a/rFtwKgYPSz36bDpAjuZ4ns7hr9GPzcrLw8WW6vmg90Rv45k8gxuYVFb0RdxpV
E2Wmda4kg6ApNHGb7BRQcoRDIYvo+i/S4dzCVA3mtU9f5VslI1ceIU1Ia4+ROqOTbMOHbTR0KM0K
Sa5Nz/JM48tOGoWDywRnltSHnsWWQHAiJr+JvY6H1NThvfaGM4W6eBZykdn7e3UU/+Xl6j5Ryat8
sv5jtR3imbC0b3fOCemiq2lKrSihVt5aUY6CSfmCDFC2WqR/Io5GO/C3hsum9V4VpFMjV4HkNiFq
8pySmz9TX0smQyGdeKeAPOMtYehovsGL0MWckegAfjEsEiWPc1A7q5d3NkvbCycI5QN5vJebXaFA
hNqKrHd9UWKt/Q8uD9ss9FRX43akFuI4mSUn1rowq/BpXEQ6rNWKQh9ED/ilwMVP4ORSx1ncTVty
2y+lCWd8kTQsBl0W8EP6qSpPqwMmhrnAjoLuajwive2hZDEfEMi/ETAuwdNYZ6E+QCjneoWi6mqd
aq2G5xKdorYvi8K/5AV+2l3lvWfNd/SyPFNJQx0xYYH6612fDcI+Ljxs+/53pLPtdU4PzATQTrQ7
Q84azDiH6rOLUG+7rtPvULj3UvSGsE0LAV6SS238wjBgQcC8gBiqHRjlCjZfomB1kPxGBF43OB9t
R4qk3yfCjkna98zekAn7H1JKRENfN7Er3uY9sQMJMb++iYAK/rZ579sg1DtChqDmJM57wIiEyR7A
Rq4GL9Ksi0lSmChBvGr2mh7wfVAKbqVxpQrqNrL64RlarqRfAM0Pa1ZzR7Ly7Of0xRadlZmfoGTV
MNZ8FBf3qdn3LbzBFr1v6Enrd8RfHk6QqCe9367Dbh9MeKONKOgPYcJLY/5nZWH4db2YqjaZmL86
drE7/s/VbN1A7m09Is91unrnTSjFkAFX6igdNMK4GDkSdBJKvvlGr2GN5SB08Tq5pianwWP7F0ab
ZsJE72NfubvraB1OF+gXNhd0JPE8X4qDRmGw5h5UjrVLNLxuC61HqDbrvznVvzLU42w9A/rkT4nx
4Qh26PnXKXj7gAaLkjWRtUAfR/2Ar5vbU0PW+9MwmYEE2Axk/NdXfSnVA58wAMM8xWuQqRvPCyF7
48YafvLXwV/i7bvbTXeqAUS8vP8a3dLKWlbUesapv0pmQ2Y6gRY4/cB1slxVdm6wsCTKv9sz5mGF
5Kcbh+OzmWyKwOiLQYX4VyRkYuodk7wIU6rluii0AxOT7yYP2RdTTT6wyWcTBw8okJomVnnk3Vua
517r67Pqsssc4g708qsm4GQSbYJxGEXaBv+MKhUpH0hpF8fG8PWkQky+7WqScF4HTlkmSPxaGDxD
/ehLgnyBGz9JKOCblqMhzEtgpU0IrdFpKI7Zo8GMkuQlw185E9lVHpjEgjnFTQUHUVeN279D+lw+
mwg9RVNVbzY8KgFkmUkVqOBrI8ou515YNQ5Dweldjz0J44oIsEPcpOzbohgNQaNfKur1shNY+07h
RzX9QaJnyR3JjY9rq5z7ARQF3ppfVQDC9Kg066dyy6Lgoe1bEtpMd2nCuagFKfq/jPzrlSU8A1zm
Dtkj8Jkphs9LFp8gr2zY8z5vSVMQCCB9iAFWLjf9pYQJnVd9EaC5c886U8lo+KMtDLB0fcyNxxxf
fL7y1vah9hBicdSUb/yVmTyrHk2BVK28t+tDsSwYo9pdzQqrJGuX1FLZUiS957zt5AT/froiZ0Zq
HYepPgUI7m6uCQCBvafbv7LkV7Wkxo9zE+BOCQV/y4Dkg4wIFKs66s9eO8w68QcNWwxAh0tf/Nv/
OU/uYOBLmv4tJ2pFWxh42D4ZzIi0bTFucY6RKy7oKf+8Axlib9VqM4wBwS8tG2U+bdVoXnf5nUi1
clmK7m1AnvXjuizdCeoAvMsRbveYUkOXMKrBu0OjI5yOTOcuotWQa257zHYCvmubUdL1uk5ZG27D
7Vr4ljz362TXjddsNO6ul7PMa+tHciSFKDuNmjGQUZKiZw/EInDL/ywjri8tIkqh8gicpGUR4wDM
MFFeFfd5S7dnci4rUoP6otfkThMDM7PMJNvFOUhlw8Ha/d8PEc8hwWhFCAUzf+2PRFAg1fdcSQxF
atK6OjYi8dfHV03ry51haWGdUc9WWpiLv8jtz1L4mfJoF3ghDu1UuimoM1Zzfoq3oYHJXs+JWaS/
nkRYja0fYKF2o7ynDo6dc6VfC99Qd+gsnnMP+ytaf9bN3/RXx5Pb/KePsn8zWwF8knlHBA+qop6u
ImN/DDIC7Cd8jS6aPuvAkAHnsQDVzhKp101y6S+ETrLsU17TIDLPXSRLbdA3ja+IVY6nAI371JMR
ogWEa3PDz4QyyFPm281TnCKeNDoNd2w/r65DPY9nubE1m2sI5uNaEVdtYNDGJBohO5E2ApSln0Yo
Mx0c0UmXR+B7nPfpD/2GZEDf88mZXYo4ilsu+JHEzrM6lOp1PWCzKe7hkeAV43nWpoDsKA9RZoL8
+ITEAi9a2/8ZSEY3Xh135x9M6T9tchp8RrwIdIq6ua8d4ellczWXBg24J0BaVQsWuOO8VHY07fXZ
OoGIlTnKS+3oGaQx3EckHrD58uQxzfXClyHQvNW6zZM48o82yM3KMKxrkp1EO7ZWvNppt4newaHQ
mGTZuiNo+dZn0ydqJUNmglSAveeypMSRRT1qencUKlJfzvoON/d3iAxJcP88qCSPGinshk5KU8WJ
uFDF3ezZgk+o98iqx9Yzx0i9Un5JFNIa1dsdtj/87kdpP8DnJFSTu4Hhk+PEv0xVb3FIHI0sh4hz
G86avA12XOcyGs0Uw5vi5k5WpuCHtFYxeIeIBdz+WoCF54pucsGkgZn62KBHJz4MqFXHYm8K5e/q
ldzeeL7h31f9lyZyYebbQ+oMijo8yd1kcUgJ6o0oLkzS0ukhss7J+yN0vYQz9weo2kmHmW//XoAg
hJC7dq2SJdZgRKndfUNDsffC2rarhBgana3QB0nb1LjDL8+KojSXc5wVqAg1AgsPSTIKu2vTsGRe
1F06MQyVJjYM14JMS8NoZncfJgH0b4Sk9x2sEqZxFhlhS8xEiikPHn66dFFsX/yWY2SdWF1/2kL3
cHIVs+fY0lQwvPvRrbZgoFhGm31PgpSrbtfuHt1YKwMVZE7EkukDXA6ogp+E63Y33ZIkkIdFxdgM
WJvqzLvvzfBfbkg3jbQtB50fVrPmSMlaXqFl0S0PeV/7sl1n1A3ZZpG8zUO+RHyXobyX/rv8mFNp
J6SLvdIPj73n7wQ76ibJZsvmYi+Twpwb8yf18T5Xss9o7l1R4DnNxAgzftDXrNSVNZoLNk/AZWXA
UAjumVNogMwZWBO1R/TtUrv7RsAWeybNIyEderzEPY8V83h/QzYQHRk9iWl+Yw8dO75MxyGayKky
IgNAg35J8m7ScQIwYZSKVi2+/N79A9MRR3b20/zZNCkqkC8aszhqe1fD5rXNtgPRuZ1o2ROgjrFx
FsoA3G3vFgcSS02iT3G1Yj4JgB3PXc/y4Ey1tiQklJj9lFvpBOxCkU56XmfJ+QO8MPIaVJEUCoAE
AK8JigCHu7Ib2rFgqohorq76Ou1U79WR8rurfOfxnCoKzlXjTRZUrb899ndclsBAopO+I75siS0/
lkbBYSQFgcamYIbX+nia0C2vWX+yodlEKx8UpYluvLSXnRqY/v93Nyk5U34m/umk8QdsdHDs33lK
nFJ7vGGTn6xy1nw3oCpUxnueq6x9QhKJaPTc+Bo06wlI/Do2lPvZ2S9d/HtpfE5t62ZSBHgWQocl
4hRf8nqgV4EfHSj1DZBjfrgYKZMtM+8X/6ux9myegV8NUo+3JDT1/Mx9lxGTnE8/WcvrmRkgRsmO
/4rAxB4qvZGVAGqRsRY4Gzv8ReDKfHFnwfpstzglucZ1Q6TcJgCypnYLG22nEatrMfly2hGdgMvt
UFvjsioE1MO+PO8bqZSD2jTX2hXCE0vxeznpMRNCB/NQYFFh2h9+l83TOfGs1QSwVby+Bd2HdnTo
zfNNzfVUkbppG2CfWcKcPaomYSBNrFC1KQBKQndEKD13KBSBtqgZCIak0P74Om6q8kGjL/AyUefx
BxEuxTg6LAGY5pnljboZqQSJv2pz1mh3FAhncqZlqn9BIO9yyqODQrDr2fnSGJARSYr+qr1nr0Xy
QR8+o6WdMuoAbvwWzSShvExBxO8+bhD8Ir84CEcxEpv3O8C3aGcZ6MpCCdsB7WQ7zw6uUc5sK3RT
2dHcKfaWZCMliVwGwfcf1zlwOk5MiO90817egy/LyypVDb6xNlv+qfO1JBRVuwPjHFdb7Q0WediZ
2kSGWYDgspUOFgnfRzejApAmnlDymwbxCRe2wgd3+9fhVgOxFQSSFY+HEeYL8dpQiflVDr8Qgr3y
4E22kh2WSxrU2tT7+IfIDZ2w/Ic3bIT9HekR4Qt5CH7apNM/WVL+6IhmnqIK5RfvXoIVhscRlhsQ
UkO/j6Jvsm04JfCNnVPNILQqAkPk0Q6ZBtko1y+Af13V9tfH597lObGpkjvgywMYDY5tErpy5aUJ
PfEdrk3PW40JMoKD4yS4pYyw8ZEUH8WB9u+XOuVgHKlKmwO3o4xRRskBEWGSk4O+oat5MrA99Vsj
hiv/4kOqaHo6Ukk9Gqr2y7eEBJNI4S4oeTa5jPEWbdF4M49X7cSA87dtX58rALrVWikj6nAWq2Oh
bQrNaqenMmTgt9bDWBgnoFRUzCBNiHvz31H+jjrcGafbHs0Gt4m41rGrwbHdQ2als6adWye8qKry
e/x0h8ubST5Jf3jHIBmjP+3yExD1W10sJvo+PMEF3KW6uqRC6nDXNumvuYRd5hQqIeezOxPyzeNi
rFh30UuWLgvsQk4udz5Gv+ttqJDUVTspRPT8Euqllxg1y8SYEEiFna9sOitUwZy1RXR3qBwXUWCK
iGEz/NaMzX/T34R1rVJvSEtPfa7qWagjL7fxHRCoTh8Mpb8p6lVDeY4ktlCu8EhU70X2KhLMDX1N
RF2HLZBJfTeRipMO4yNXWNAX0WyxOv1jLHCtC/dCdBokNg8E+zSSCOKclxAO/23Rc6ZodhyOyKHT
EwbZUGN9je305JZwlgjUSA6N+B+kPE0V0bOHfCxqx23Zq+e4fFksOeG58ei9n6hBKC92eMFuS7rg
p9YAeTdLGUQqMCAMFuYJbjpSjJbi3vh6q9n/HRcfkZMuLApUsil9/lpY1z8SD3rGdOTvH7Rl31Cp
ZdgPzdBesWeLZOKiuHg3wqqjAeCuY8ngaWx73EnF1en85qMOJbUMIE/opqX8tiF89kp5CPFHFftA
Gc5chvZvZ2xRSEBE7a3m8lk0jw3jx2cO6lhwFbMNCSyH5lOTCohNzQtG+1Zd4DEP4EqUK7yoUvP5
d21pbMm0T5buAjdAjdmpMx9l/jaJYtBDtj1u1a8aCj1qhfFprEda8cZTieHOm2lWeQis8zzTZle3
YGItKqiZI8cvn2k3wwxYvhNa0eYdBWGJq3rb5G+pmx+2gGqInRvrYWxSpJvfRNqM0YGE04RbI6BF
VZaObS/5yaqvY7hTNQyYT121f7RhD/AzGYCf51thfZ7T0CV9JzUIdOP0Dl+T6kXO8IwB4FvfwRXE
wB3bs2d8SvkOSeZZvkKaNP8DW2hUFjbqrL65/o+SqTqRlWkXTKyhogTXobGfPgPV+13RmhWVMD8A
ffv0RbYaX4gixyAVMR5wKMOPVQ4SLNXZ0ZdboGEt15vPdMsdneLBU4iyosfLHDmuBonlc79QNnz9
4woWsGhVQ/byv8aE5hJbpAGoHQkKF3Y+Y++0awbfddkXYjdDmsZvQ3Ck5lpDDMnb940wRU0TEL1Y
/IRpT7vrOUPI8xz3xZYXQLxth+XugDCoy3+ETD4H3UV0Y382JjcZRgdx0A/z0blcT5StfDDr1r0V
mpN377nAPj+xAL0yNTtte6CdlIq6llrOkUfgphV30rDsvZfIfhVzJ/1UiD7gp3bv8YD52gLZArxm
QA191LtvQjW0T21yAGthaGB7H0K6xpKsyVxvC3JVhAhRzsz8bG75+l5WyLmIzqlKvJu375O4HrCK
6sL56JDNRf5FdPL5yZuZ2OJSlI7kj2cxeGo+l1ECrBbM5QNrWXxqdbFiPSMa507gUz3t0LDvOCow
DYuynxaM2Vm24ln6eIPWcgEwCVGuw2ZrthA6jyEIP//e9/aD48BeCW6/0B8uN8rFg06L3JlE3Vmf
PxV4RjmeQqWSJoeaMtOXsilKzUPNvedAkC1tmuWd4oe1qhxc/ZMIYrRygjNzP9xjMTa5sAF83O7I
9ZdVrkwt8kTJb4GRuawJLhlk7Oiig19zhvNnbxV03n70r4hq6SpE3sviogxit9/wo1ZbNToJEc4B
KRjfopq8IyQ+Rm/ePOLU6v61qF+nZ29Shuo95cNrObN+V2R7wD8/9lzxDRjK2XIChAI+DtT1wI9M
thIX3bfF0oF3vWg6LrMMsVNE6seLlx4iyAV3BII5qShBy9uk9l/qgVtXFLsmWrlDe2okZlKaEVrH
4F3m/bOKGuFigdVSgyIiC6zQTPbcO8XJL3ktuIhfRuYSTvbmQena6C3q3KB0zc5KQqmxT7Rmz7y+
5MRp8+aWZR8+AcYC2JB+VmmCHuejtVfKoLuAONq7jAgnLLcAKbqE6h5t+33LJeI0IIBsGfXP+lK7
1eCAcBbbRjftysrKECJvBDwwsGPb+xK8fSGWZy7GrL/51x3uVE0PNepPAo7FjQdzIH5+7di/AMDH
9+xTnDNJ/4Aorr5bmfl23r3/FG8cV2zc0qFYNGBme7k7aT7aR+jAs1BfAvbkC7/BWqJRltz7XDhh
eQ6fGYZENv2No5NuiQYuccNHx56P+yC22MYkdr6cVgAkIUntJ+3X30mQttKlr2MVG4QtA97LPkc5
6mDiwFj/Na63njkrsvlHxz/gny9GaApReyJFn7f08awaNoW3GYgQ40rAJTDyxXBWJOe73EVREoEV
5iDxmNFgMbC7p/lj7CTfaLaWi2nLd9nUWf9oKOR4se+30pqlVpJBlcZZ0hLtlewI5mJnYb87Gn0F
B3s8Yq2vsafJ8c/k/tZ9oQU4bQWBJ/sPZWnkqf9ljGkl803by3vIL3bU7Fam2tD0hskQnfumyzZi
nqalKzNoRYdDnKHNkzE4cgWjbEBUPA/PJ8/KZEW00xpjaCtiDwkMCUKWG+Ww45ZRRAJYhIMLI6re
zfgcWgvLXlbWWNBD5rbkpi9AynrzeQFLqWkznMJpVy4cIuQ6Y5HGuUH+S7pDFBmh0RHBFJLG9AXT
tFppeSCUginfLirG2/7fuvxRPWa6tTfUd1o1dWzH+Z8a3Y3W464H0Bgi9s3+pPcDFkzFh26aEt4A
Ky4kaCB4jrezFBxh/DWaKgGVWSviI+PkpsOhvy6MhfMRypez7NGOffzpBW3+WDHr65RC138tlAaa
P80uFG+pWbvyKJr8SjyGPPsCeBgyXOspT4BvCAU/rdYQ4hQOXgBXNAyLxlmXGWxyQsi8OE/1frhG
GRMMa+WKK08tUuJRwLgzn6Dg8gm5k1gIxGIotIEEVaV6Gw5Sj+7ZEze0yM1pRfNVncMIsn1MY0Jw
ZM+L1wHw0ZvxyhpI/7tz1gM2LgspzKTJkhHkuUu4Xa+cbJiLzy2abS8Kp9YhpSmOto55EzRv7vbD
F7sIyYD6ykUs9SzedSpUeRnMrl6J5bdKPjxBXyT9hTzgSXFjb+/Ss8xLu9C7ciHNxAe/GyGKU883
mfuhB24JUasSp722NESkyqjsfZWXGCVj/03KaBU2w2YsttLKl2dd4OKEGdtJhsvMGkXrXxNAysQ/
3n8519YRmCkF8NZfmT5j6eKYf/ZURcSbUQrzLtgH/cxJ5oi86lbZYODkF4JwwDY+pCwRj9ohn17p
HvST3jW3IkwaN67r938r7UQXzK3gDr5NXkEWCYrLWWZKWe+vs/l7uwocX4uHWiTO9ve0AKgf/hev
6gCQjsHNHmeGsf8Ev8sJVmHePkd8/KzkvBXaSypRlgC0JRvn6JsyAX+Bu9tSjkPqUMAdrAYOnYnV
QfGuhAY7gxsDloDqPb3ndIzcMxuLUAfOIqeDVMwfAJKV1qBbU9TLaHLUNdg8L+6tsQPinUyw/7Jr
lGbfS/RjB5jd7qXyfrXxANgQOPFupQpKBPw6bxtl0Ua2wOp2vwfkHCFIPP63XGOL9OFhEeTUXpXR
MKHuQuI97VcH9R1OJqHfktUcpqBaifgZj6yHSn4XHgEc79Zy05UcXPfYwPbn7PSf9WVnRSuo/g5x
0qUQdAbv7ZRlImOUwktUVsh9Fcz46VH5Y5lYRx9DiE0ew2Rd4V/AFZ97szJGpWBReDQlbzryOeJ0
Xv+Z5hdEKarOD+aZWhj30qSe2lr+4+khrMoU/Xkih60HbVKYzC9tW0gtzzTq9Kim+NDyjMRZat9P
tqQCRkuuVb84fFuX8v9l31ZssaETJFbYm9Jo+OccHWlzp1Pp/VDQFWH4x6KsrL2dbpaL5PaUNpvb
pYcMj6KBwhD7XbsEqg0ejRe3x19mYs9g3QN/aM1zyV6d2TUPaSWA7yWSwdkAHr3Kx4lhKKH1pcVx
rcw7nHHM7myYXxqncM6dLRm8xe1EG/Fj159ab+IdQUjj7NQxnuJJLZ4oLUiVPSvLVcyqwRB23znI
XPVAZ/jg/wAZMrgkJTuJ8Exi6l2vQap9FQvAddJjsJFCawzx37aZhka00ownhHLTz7YA6LAPKiUX
77+8AN86+aFTRyquqxe5h0Qf2YWjpupkgbXqkcoA2eU83VE6PbDrNyxZS+pqAeyNWr+E1iCwWA38
hje5SnMb7OwmsdVv2zSGCOZC7Vzr5xjndkA/OV2Qi9/ga5akNCRS8qdrs4y7xQfJ+zSpPFe5xxpu
A+klrzzGBLFkaM8XixyuT5JvL5ZyWTWXl3/d+LDHBqURes5r9O2ZSQDlzWJrPpF6+zxKaCGn1PHy
Pqd1jRtZ65wiJC6r3j4Z+ca1/glIghXgvyDlbtucqJfvDhF6m456vgLM6JD4d71G3x7BIMIvyCBv
6UnQP+IW3vIW927m70ofOrOEG9hJbqe7gS9vwXW+jYFtcMA1ypmNrnD4VY94ulSn6PTvO8XlWh1P
YaL2k676GBnFD3Ljo2PNCi60PdRnxL8y2XaSe5YC4pjPajfdb51z4CTzUBDAJspiLIKZ22NaW6wm
uo+6+yHkONt2/kHTxB/9UjgmL2tQ4a2db9PhMVAdTcDvkdXYeUjbKpFz+pK7fSoxahKoUYppWf9z
omhICo9Toi9F/LmAR8JnpfBGK5hf0kqQHoNGPg1xJPcEJyMuQX4u7Z4q6Yg4UqnkfZFNkhZynIA8
Ui2rFxd5b/qFzJSld+r29EXIkUWjeVosUZp6NqGmGV2K/st0FcioF7I5u0iYjL4RHRK0KEC70wcJ
zKfx0mWxgOjRC/TY/knRsFA7Y+aLQr2Zd9E2pclmg2PE/fP9Kn/oEUR8efPmo+3b3FUHclHpmpP1
CHuFJsd3l1ufO3tufqklF0JpFYIXvMgVQ/zzo7s5PH1OpAhCKGuRs+MW9waABbf7Rl+bmZvYa5bo
F6hWqKCqXCGytU3OxUlcVN6qUrmDmiV1mUESK6ulmXE/24HogeaesphsuIpfiVDa08uM8cMUmebl
aab2b+7K+olQ/w6ASnA6h0DZM03kLQ0SXqGIMUB8VjEBsmN2dfV7PLFNVGe7Jz+kXtpEb1KSKc+P
SF6Rt/KeLvWHMf+FAQ8ipoA0uuRrDWfcZnYWQ8arA46WezBYyVHQPp1vjPNjePOTh728O7qTLoCu
ocLgT0oaoAAAmqa8P3wJngKKxXZq05cJFo4x76Njl/QGcu5pt6CVJyxc+Dymb5GO4vGPH6rdCceD
kLWWLSdU+SIXXHQgTfdseie+bLGX8+JzS8z+t4IYqUJX/+dqEJsBvesXfEw8kvieoHx1gW2lOYZF
29VLTlJV1b1UMXtEBmWG7eV7Q+ySv6UTWOulLo1XtgnyGm+MoP4HiSJnFUtnnwt/nNrWUF6aOigP
t8Rt7gypFFAll+Jr7qQ5uk5j9JVo2n6MsEkEDcXXCRaWAhALdyuO6E0JNkENWGZ78UmnvfHN+wGM
iPgRefLvITG/Cix6jBF+PZfcFmjO+qXvbsTBF7Sd2OPNIAU75ex8V97SXK4FAjm9FiifXFC2IAt+
0Vu/eOflC+udsiLbJHw3x84yP5i0jAvthCqD+IKzW5nGjKWJ+QvMSJry4qIJpOsBJH3yKthwqv+w
kNUx0jALr8YkxGYPQASAWzr0sHhwp2yxeTZkhv0DUMA0DESYkC4IkO33hk0QghJ6QbF4hKF+ctHd
vhT0pjNHHfk3E5loM4LVlDaxDYyMFuQqoQGDTAHlhi3TiuiPJ7KxWkxRG9yhB1Ohf31JleBfCb3L
oQMYC5oO1xDE/ucKUbNMAVGoyT8XLCb37pWC2s0wMU4r1z/M8dFy5gsjLWp7o5WqQ8ENkgQrvac2
4qDQYd93margWi05TBndeuiuiRfZCyuIbd//aib3+hIXdCLetTQdP590mJNi2RGsDa8sxG8Uwe3u
aq+vdC1MG1IUIPoU+m8eB4qyssif/HCGka6ih91exSfKcU16hOc25/kfXTxVk1Ic7mc3DzRSIqBY
JaWgvue1GU9BTeBWI800pcbwjgTkv6fkNQn7Bmcc3ASM3cb26AIxsKJiR9Tj8zypEERpP3Dkg1yS
pes9pAGj4scGrE1zz09ifDhbUFE4aPDD9TfUxOwiF2D7yM3RxK7kMRa6lbI6KyeZS4MvEfqIl/IF
C1ow9r7R2WoXcTGYTpAjt1Qa8nbRifIfIG6dRu6EfHIwS90RwdwyRIdMVQ4wYnbzlEgOZVhmArRi
uuZ+FsEhZkrofToMGGf6joIOcZcpEzvlcVklKZcPcSZY9KWEr1FDcHaGeIK8LCikBVtlGeDH0VOp
cfLjarpKKb5aV97+fLpg+Y3/rXaRcY2NaSoVhRIjUaZ8Y+eFuXD88YpFODyzrVWZkFIvPKhKGVgH
qWxHYpytrfteOQh322Z/wUpFC3VyyoDZPBNY6IguaMLplo8d9SfwGzHdSAAfrZtMWB11KHmZmGqg
Dmj0q9cRwBhGep6D+mbIifm8GMlMAb/QM8VgM0ADbiTpOK41p9THvgDXXid2nzB+KwjtA56YeXiy
+h3hoakPQhX8N7WU8iozyGstP5qeokR500vGA+9NQnfsgpHkri5CseM3RMlT/fyraUMySTde1eEo
ife/0dCL/wUIku4+j9uwqqmeaHgqgodmBx+N5BzW5uaKrVNKPnFJzGIS+mbZfFJN8Q843qlgoPMW
EoAx6GdJhfOUKB6DwpJkOm0HQVCiNeXa5o7FG3jWiKAOJfJFIUvXpJi4qLI+aygXSU3yZdgyA28Q
4X/s341UcxdEeuhJf80ufmla49OfiBMv+d/FLMAVp8D4v/+/9E3dQ3X7JCT00x1U2/LxYM5u6NfZ
7gu4SaetQmfnSEfodVb3pTfD4+VJ7NNEz8g3d1/Z1iSJ80osQ+cClZrilnizNMylbGkpxGoEZtPg
9CRKgGvpuG6KhM4+niJaxEXVCaUPVZa/o2Ts6d3V4ZEKLITblU5GayrDNWIhk+7vs8/eKX1YYo/I
z5CJ/NhioVASwVGNkvQpsByI9XrsU2CXIBxJ7g/Lzj9/MtYGKLi4aR7Kk0Ze4hpkGqmBEg9McSw0
aV+tbxS+7toCW3z8Ufr3nQjsKPvd/iauBwsSuF/Kpuc14U+9J6J+HZ8EFAhOI/iNaPsJG/5KmqqK
gnr/nLFN6fcuzdO+ZwJZSADyhfOXCa8wuKwkubQhLtrQdf7OA/T5DKRRbtl46uvW5z35TdbLg3EB
YBc6XGYQGq0EsmF3Je9oSxmSAapdP6mAIhx14WL8srOaRmaGMIrPLKIauswr+gHNah+ET2xarT6g
s7sVsy1nXGJy8E2VlG4iGKGcCeJA1ATFLQ/4PGQxw212XpSq0wuD36y2KeaB/rXa5B86CJj6V7op
xejywxjnsWnG3gD4HcXt6HlgaREji094wIn7/8f6FA7CsEMMtWThQo9mikv1TK7QCraI0Hj3t9Om
iuDYvJP6MWXMACtM24RUit0nvPtdBNN3WeCUuNnFrOxIKrdWozA0nVbfJMdevSo+8DQLRn/9BFOC
5bFksdZCeQMRR2bEzRLVtbiQqH8dwsQKVko2ThKNnAFJHdSbCMdMBR6sy2ciUDSL5x79sp8MHaU7
kncFQz//R1hEtNqZ5vZTi1lTHePOcCJ+fga5PfV4OOGptZmxPeKBP9wM5TY5f90dnewd20egn7ab
fhkUSC77bNXLwN2Hp/B1+n63nCugHxvXUhico2l5CI5vlBoe+0y0msgAZFPj5vi0Ifg/RRUdrg7e
Wz7W6V9IfJAsxpBFDuu0eClSQ4nUCJDfkawz3eF+WeN3NM4Yjh3OnQC/FW9GkM4IUoLpa64GUT0B
pEH/3NkJnFGuF+n5FgSowm9izx7c9mh6hE+2mOn0kdTdU7QGW5RDWXl8lsefGboaSMgh4BnUrXlM
RNNuT7N660Iwn4OLqZNtb66imdnHX9HjR3D9zulzzMrqcHONqFGNmup0SPRD/ewyTFHDc0DyyU5x
Rtdi8Ne8cIemummU1xjiMPMxgIOLF7GIwgzG9n/jK0q0nfsQ62M6oJAS9QwTQPV11YljwTHYiRPS
/ZoQ1mlajTWkNsBevBJf68Yph7FmwlA14Wsw+y3r75f5YCqXaOJiCX3IgqBq4GnDUhN9FdlP08K+
+OZkFoXRz6hWqZ6VAYx+iKkwZ3yhhyLAtU7kMyYbiaHPRK93L4Z2Qk8z5xm8aMJswMs3A5vulvVc
yFKULqy2zde7iY2hflevMTxh8DSr86jrIjT83MYscBNlPoy/W3OnLOE56Bh9q5IiKpodjz0wleFZ
5uh9rlbjGLfQiov27k2r88vq5aMKAWt36nt9vSXkwNm2iZGmurLEDBtwQNLT75otWg3i+ydL1FZK
d2p07ooK18gc3bRNBPk0VShH8WvY+tJgR9+EIIAjHjtALzSphQfItZI0tqCTd8/ss36x6Y7c/jwQ
zrfEzjXd2cc+XIhtKiycSg2kJrbNL4GBNwgxvOgO6guPq6Wvi7yvMxFlZssukRtgUg6Pjg9XKpo3
EY7Kf5hScME93yG/s8l+heeuOOezYegV7LhV5mNDC8JywRjpqv7yDHsDXlLb1t78JF8AGlSDlooj
WJ7XdM1oycfr1qweaE99jTeQJQzHC/IDxUdSZZsdGHmBDyuZIds4nvsCdsDLD9r6HPwShGZKlMHy
GkF+hc6dPhJb6qmcFf6hiIf58KK0WXFrZfI9uBhKmNnrxgFOsDcp5im1cJPuu0nxLyWI9lQPUSSP
pw3O9QLZ1rdusMZ7+z8X7i1e5wLPZamMLl3EOu64Lg6zcfuNwB0Wv/ihv9vYi0h7KwO+6UwycTgc
RZjxcEP8qzH33ZsuHW2Vymym0F/S1Nz/z05OdA2Lox8Af0Z4YFExZBNvcgQZNvRdeL7LppAdHsOn
b8Z82YQlHGjoyniEjEgmFA9R2vPpfdeVCNOe/EduJAleg0kxzZuTOLQy+lY84M98oE5a9WrzoUPd
ncuAPdPSSQqpOUeaB5otqIs/Wj7dS0OR9xnuY9DVd+h8dahWuQoml0K2zoSAbd26sPWGQCaUQbfS
cEammMDbLG248CalwKvhi4qE2vFWHGgVJM8XT14E3J/J3VaEp87WPaqXZU63G931w7rHlMDDRrGB
dgkjfJEB2Kipp0oARurog/lE7c/OtyKlgGL2hmF2bvuCVrWcrQq+0rUVLBj7QmVLGS59OP/gl2Rf
hwt5k2Xz4Qw5FIpVjg3H7qZuzzWXIl5h54tCqnubWYImHWuYUF1abSPYzacCcoMiXu0EfdZV1fHU
aNswA/VFFGJrk0AXqDv44loszlj9duKzGAqGF8ss805qXe/GgqRJp5aZEHwsw8ErIGv4AXA7OwBR
EQOBK2hXg1cEcnf7VU5D/NI90MVyXk2oEhwtPlRKD20Saaf//BKTVh3Wm+M1rIpuozIncfwaUzvj
ovmpIDy9KDu0MzjHPJregz0PEjQwAg04COFDNKK8NaBEORZt6ZJDbTVqqzdSrnZ+X17V1BZxPlFM
Jf3nc+NF3oJWTT6wXnqdwhH6vtmcXfp2cSPAGKl2vkTw3U9cHDqkN2AzuguS4lC9dM3PqhCAo5AN
n/BOqEVd1yIRdAxJCDONE87/Cdu7i27OWTZ5eiRGUIIEww93hF61SA1LDwTNo269dRnG0qTfP4/A
J3tkIlOKwKmzl7VBm411NS/vjo04yH2KupXO2Z/Cz/wukbzSgNa1N+ysaS73+h9uDVfZWqqFTcQX
oZNwCiFfbGJrbkkRp2M0O8DzBLKmYfD9Yr3pQHtzOOy4CBAIejDjzjcD2XlA1K90RgvXuUzLtHZ3
3SMnXgY3DBjqrMd82ObzDe4cpu+gRRsXrQMM9/n8ks5LPz5ZtcJ/DpEANOwLCgZrZ7iLYIA6ggiw
vgT6HyGujHc9N2AwKcfFFB+fzuKxp78Q97XVKuHWfs6a9U+X8VPKxI/CaZhmw55H6Ti4CB+uyf4z
1UWhnObA8ddXGkCSkXojlQIVy+KoKFezumcBX7Y7xsBbYr/b6sQsGLMYA/t6cFDq8P3YACFtV1c5
cntuBxn79qhkyeVrgmDCkXKp1W/bN9ik67CoXuFr+n70jsxmqED2+f79IZgW8OexJzGEPZKMyq79
1Ebk/HQ8kTWSG67cVsE2fhU+tdHxOy04XXRP+RQwYDVErO+lSg+1jpREpM3QEWH4pO10Qg/SVv0f
ETalzxlC+7E5ONVKPH/AcVnbheK2zWyIqC6ZSrN5zPduUDrlwKtNLGmahvI8yv75Ttg19V6kgpaC
WWhlspP2VHQw4bJAF0NU+RpPJR5fBpYLZ5NRHzTFu8Myk0Z8xqV554h02237CwlAjtR9TvTHq5H8
ANsVhZPgB11WqaRIIopY6yXY4/Vwoi0VAdSxPsdzgaowShtDkbyz+pYNsGlvVmS5D/O0hci+Dd5n
5yizdm8fzhSoWoqPrXGApC8wl6yJlB3FVKntzwKqnaHVhBZc4NawQXsNqah63SK17GmcwCQJMAzP
TOmUJ0Ze3QTu1CuhqZ9M5HzsGTLmmsdTdL7eIfoeYqfPkbKzOvldV8mKsxxmXZQogYqY2c/xF+oj
uN3X6bXvihifciiCLmwdC3Y+/XfVTBKTobeNU1X8xl+CzZxTy8iNJg1JNvmuXlzh/VYM07Dk8e+x
x8+k4vfQKB7I0ZBCqzjxYs7b/Em2sqk/khyhx8I0F2tHzb0Azr42Zkp+hnsXlbEtmyOST6opOHh0
C11rx+jSOzqmqgCPw4GoDJo53EiEnRxjaD706t9/5+yXlbXD8/0QPf6pxgNou4RJiC0I2KE70nWZ
QaX60y2uwtkxkSj7vS6u/8mSJCvNOblb0WOZT/qusLGEtbDPrgGO70XrLLOUHkNEMA7ETYNFOQm5
YJOJ8feaSwfDQ+8m+CZlY8OtwWG0d8QAp97fXeLMlU0cyTfNClnjUkd1Dd4I0+lJuTcuOkawse5Z
pu+DC/ZvQhbB2tiCOMQNrmVTD/Ks8iy9VqTZAGT7sxr7ayloGP6i7dSIGnak899zgFO06wVx+P97
dVlusaMDa7lYnoIt8uOQC/ggoxg4GTR61oysHHfJsOKd/y7UXNDV5qO4JYd4oVzK97RmBj+JUSdf
2q+jykd7vf7P33jkIXLnT4Wu94PZGRhZJZR0duuQX9sgovCsyZmPLiopYNvTGt/j3HHlwop0JRp6
F+RLE27gZJeSf6SQe1SP9kOu9NPZzmJpGk18cay5lVTFOaN82beHOcgSIz3bzARYXeolGdjpllWJ
6TBuvg9iVbffT+g+K2KXGObVgZtLYRYVyDILnaf68tCJpbgxEewc6hllkpJCfdKc8rFsFAHxJrOh
ZyIEkzxdnrxwFeU1SqAak6C/h6YQ5j6LHIkMTJb+3WZViXLAKC0lQPBEA9GXbexC5PVFa+iYHYEL
5rikx2Vt5jmGEIS/Zr32U0gshYM/l8YrVGwN/iEvFLKgrLE+7nLdTCClRkl9smA28X9Yzxc+8EEv
t/9OVfqf3rKJapGwNgNdRZlp+8zwAQtJGcO45u1zppw0Q7EMl4cdmtEnSKBk1M4P11X1yhPdD0kG
rToM2n9TwwuDUP/9ro1esSy9Mt7Yhq4XzvHbCm5hcz4xyofAzYV6Lxq7/z9aJ+BeZ0tXh3kJkG9W
JMGLFjJ1CkN5AFJG31IMo4zswQVEV7N/goLj475Cyw8uM1XrooLZXnzGuved9TRSjMM6odwXR7hx
6z8jVgaHJThwlXC5Dk0kdjJtC3KzbHIN1F43qFi1xemNBWFO32CkF8hRZmQTYJKOHdoazWLLzKu7
KWJtF8qMJZkgIdpEaVwfSPIMoMh38JtdZuJ+PuvkAYqcJEYZSeP+D+Ftg9f/fIe6Lz55KkdnKx/+
61sSqFUfWIr9snvLpa5Hbh2N238HrJOR1ZcOvuSgm5+zoL4vUVrsDP66jsOTjGKNjCuV9nfD0k40
5Wu2fmT8gVYezDEpXNc4r8MRJ+iCWWcWhVFuzVwJ4KxFMGLm7fwJGmantutavzpBjjDtiayWZtGk
5Hfqc4DSLHUaDEgZTu+cdZDo6X/pifYQ4vPw4A4oTPUJbq9h5cMnoe1k127JTP8TyoFVM7TpEJH3
mxpd3sHy1IsKouBew+hlvFFyiDl14HqC10OmTq7oqFB470PcILPxb+geUFt7efIDoVHYDQuXMZt+
7sT7tO2xX6hhP9nzR3jX8G5JTCK+yTCC/AEMebYL+w2AnZxatRWb7CUQGAJZJfjocZd3/asyMqXz
JGg4rARKTryVu2cnHsJLHyMvnfGp6yL8usSm/q5wGP0WFIY8Cnk+QRmpbjJe+vbFLGdFBIO74K5L
Y4Bd8xK0+eLzL2ps0VICupWUOwdpnUojSraR1XdpoOySn9vFniDnKl2qmZ824Eei16XCqroD1S81
cfjYZXvri7DzAu/5sueV088j/oCnQtCkPQSGh8xl6uibwSTP4JbMT/cah38Csg/BtdboSOE0wq4u
ppWLIxt1qAbnjcdWojlrVi8zdDEK6tvkKMg1n7PlU8oq++TIdjNYtVurvhwwF6ox3/14T696G8sF
p0OEnyB1hewyJqMDJn9AVQZfRQqQc1QXMJtw5IZDJIzW1PQ9PesrOVSFFPmSF/hbHrFje5iY4pQL
6WTvcDZ2ovjuV1y3c0hAPpcTBobM2r9Tko+i9bedC8aB6qV3WSHuKtHnIcF6zVDmdi0oWC/HDO9U
La9DGLD5HQqVujopvugPiXdq5ookVsIx9zkeNcEcjAWwtL4Lnkq51HewiYaPjeqyvF00ELbh95O5
3TWvp8dfMXLc0NN/TqoOe3XFGLt8mbsUyPPDjPthe9xwN9ufLMaLiK7gCKTZzYJJlL6Qa1P+0qVi
96DKhHPg7xRruzH/pMiaz4p5C3OOKzLs+eL8D30z6B0jKEsXnjMFzJWBq/i6HGF9ahR4zK6Ji8s/
kGslOgB10vUxb9RaavgE12drJFGDO/iC1y/SA05Fh1Do6TFGCFtkwX5xum51kxtTEvA3yXlZmMFV
BMn9uQJ6insmLAV+HHwL++mqP/Td3KaJxjZ3gQkkA2je8uco/qJuMi2AYHDjMwPvki5ooc+3GP5c
eODu4WSoozWOqXtEDWqzBhQTH9zz0gOaaO1Wqz9hKhxDWrnHUZacSLqO3KqJqTLbbD++u1AehWWr
+Ri/enibS3x68RtNwKLDRnj13j/iwiLacIwHDvVcOUl2PuWdUq7S80Pu9CZJiV4Vmij2OG3yeRZU
PzlrhEQDGLZXybZalGHlhDNPu+wF/MhAVT6S9Huk5YM6FWPZclZdbdc3xPn3ubrOZ6m68pBSs+6i
EUWbKkwHV4eZOHXwokCq8407O3S/EvDqDe7hngcJ+2HM4j7ZBaEJq73BH2gfseYiP4ScFpP0pFFS
FO2V8NjmzcIhR+TiZBFozXC2uu4lbtGZXX8DUmFtl3z3FD44psE2cMTmMzoCABdWEr6bNJa8JkPw
vQQb+FTR4yrKnrNi/XOVgQwxWm9VH+U3Y3zao/p/fIr+j6bB8g/IhV+L8pmuJsCorxpq6zkzIeH+
MHKzc4BVBfoDSM7j7KQFdRjcE8UGF86g+ioEvNN5V1KgOc/H/d+Ttv0Cq1cvppkwDgoJIIwgT5r+
l7SqdiidxnnwMh4qiRid1ZDuAoT+n9khmDWr8kgOQSbNYUenTWYx8qX+mxgUUd7hbu66gFNz7uqf
unzoz2B+9ARBxt+OTFlO+v8rRm0R5HYEhZdthyd3tAD4tyyfXwefXaHqTAACAk9ScU9oPtz1ioxi
i4OwWtoEhUp2ew6KRNH7HEMJiPnjq/jFKd07arPi4OnHXIh/N/BEFLKS4YhNuisldninCn3SXH15
/eD+Ws0l3SGQZEceZ3OX8yti0bpgI/D9pwY9EI0sRUuIzGEA9JsZCKj6c5zFE59tqIpBdbPlMENo
v8p8csqMv12wNee4qejQ2G9kU8SoRiIc1VMV77/6k+PR8qMr1ug//QctBtdgiwbon+PP+wPW0NG8
c4gUkJyQ2W6QT/aiOIl62SKbLEuTKQy8VBIt4wKiWejeexAAWPBC+dSZxP9R3+V7UhgfB3jPdgnP
fMAaud3ekuyXUzQARmWgis9Y9+AGNtUh2uWirZ6BJIVwM5/lrVm6oUkJnCdwi8ZrUhIyE0cEnT53
qkTbCsE6nHh0G+1Ovuui5uVZPfCZjJ5d4r1PUdHGP3xFF0kpfm/KEbBiOLxN/LjulHbKGRO9cEd+
eoGLLJpREHxOJQU44xO04bm+CaPHac1ZEpv+rfCqXRqsJsmyxK4QQk9RR8p7V7mchQwDXbTZOkr0
YMXlI8hYB0JnAIik46aMFkR0f9sipeXxcDHEZ6Nmno6rIrVJGIPAMEHLUp7A4d6mZNiIQ4VQwAS9
vhg5bjMyHoJ3w5gEJWAYclm/xWymu82wYS0QHcmZES6X8+NAUZ60+UrXdfSJUr2UwVX8Qs7tpSNM
p3qVcwo3k4jRcMeFLTF6fAEiyfM4xW1EDuzMTtOyXsd3BikHQCd5Fxuh5dvMxtSd1VIhtl0NFgFM
Jj1gkE8cV2PMUCOi3PyPlcnVM1IIv+IOfj6lEPT/msz4kRD84T/7IfayNgSzuXymzTcI8K9i2nbS
my1rmaQwqbOJhYTCUB8Nkg1YnmZ3QsAkHJr32Mj9OhfnAYJO01kkhi8vat7FscgwlJeV8cH+UWxo
1trPjNyZn6fvz/rI8JrVXWziClDb+EWWgRg/Rc/HnMK+JeWTQta7WQdctmfOdQVcjz7PolbbiO6I
lBKEpKEOAmsy4F+bOX3nQK6NuvJMs2VxkvtYvtrUJda7QsuBpXegjD14O36XfOx4W7jr0bRVxODK
OvLt611QHUqSdish/guHGDRKZYHKe6OC5E+ngYxROiut50VSZgSl74CuQTq53s9YkFwDYNLTTuMA
ZwlJmnHcfDxKJc6zYPsFr1avVRAmajlSg3xjtZSOYxsgSYoMlflkOMnbpyWWE2O9u3IY/33CSGR4
MKGUWA+dzFNvbz1DBthlzBltLuql+SFzgMJZ266nsGTmAWkaP/At+5ihMxLCwktWxVwl1JUSYR9N
KPGCsrYLG4G33/tHLYfh+HPdz8lJgFWSoAFVVFbKbawCkf7ap5rlE2wETZ65OJobp38FNpqrI8Vx
CCxAL8uZfN7iCnj3S2IHrjHaZWjV6THIgZylHxfXK2QxtM1NbtLrInxUXGofeva0G24Ff4lYaKM3
fg2za9nD3Wxg7AqfZchWR74VgqkboIwDWQ4J7pGJxLtojlNvbMu8f0kuosCcEroFaJxoDJZsOXUL
yrejxIhgp57EIH79YLuC0oy7uHRaUb/yFoJQl7UuCsxjPs4ZeLp5+Flv25FIJTOfQkf9zB9I1Oz9
tJ+/x9S5dGacOYYYdprInrnYg9VnCtcmCS/EV/K6yCjLIA8Wa4XtWrwSmHU5ARnSoPNPRdgZe78r
3ngmpo+FvmC/8dczfBTJ6cviGtfOLVeBvLDxuW/p5yisrYHnNHSrY7CzekMoseloQH4YseToyA5B
caN7I9qS/kTY10s2Gy3AIRkGIr7bbeMw3uWSR7xwdupc943EEiOoGjqHi83Oyp3pK7WPUj6LThk0
dWfj05ucmEObdkFZ+jZ1h2ib5kTGmks5390y2Om+wTOu5+q0sZn1wR1VpXEIGIJ4UduYluD6cWTt
BRnSWjUwXLd/Lb8MXMZMIkhsVWP0WEyHwlu0wMPy3jPPmBlz6eUvDDjcuFF9RxKnBKDKMw/ZHNvY
VL0ypB2SYA+2FJgwA3Y9rfHLmnKdzPW8i841Ney7Ojic8Ui+tP0IIRyclGcUgRGDxgV5jb4kQ8MU
jhaBTtxCmyY1XahVpuGmkfIY+GUB3IAJy5YXTVuS/YPIfRhhrGGMWPDNANG096QS/5tz7mbsjdxc
ihwuXbiY9zMxKRS38+OvS0u/s64bPFaGdc4BRbbbKmq0xlnB9zk2wF+5QSYJSStk9W2FCY3hz24j
+tO1BQit4ost3oNiknnuhuVffQHJK3x0hcZq9CWqszVCEFyaBIfxULkARmrqEwjjObCCTbtP0HSH
ffpu8bkPV9YQFzda6EVrcsiaQE3tmIEMf/JRhJ94GpAOv7qT2KQlueGk6Leeq2g8UdJumHtFgy1R
TwH46cl/QTEMnuXc1u0GXwUWApQDgHiHhWRU7I+nuONZbo5MmCbN4myB7/kDSqDMtqQ0QZJp8qS/
I79PUWKXQdAEYm/lmwQTRNAkqXIrgRqgIGs9ulbtjRhayQg35efYnhNRfUnKIOSXX6HG82E2d0Iv
6AecZy9Guu3JdZIP3J0XbvNMwugy9vtDep7RiyDT/JbA9ts1BHI1CfDzySq38rn907XhdbC1yXnP
hVhG+eX3WX9098oMmgwl6qdRbnTdQ9ljIpKz2GKVogUeeRVAMe2uVsEuSz86kdge1OEDMA7v7DT7
EQ9jYhrQJu5UCDgmxreBVfwvrts7hGN39o+/QTNrZsMktJNA+GHtSeEzlCOffAHtVXRkPvSs0fLJ
/KXdw577+spH3mJor32bGqUQ9Em7ESAHgaG7iW97mYz6u0iF8KSke5b8ue+UR/EH2IdhQQX5uRdk
R6ENyHWk3gc9LxNuC/3ukShZLKqryYufb6YMD8AZd0NhDDpzEL7iTIrOM0m7JQygOhVEQwLb3DLe
N1QIBEQyBF5TIbT0kinx/8mSccyA7wdaBtwGkzraZNMSVGQ0sShO3k10CdEzkKbYBy4pTszchuq0
jhCfE27uetJ1tlKdGX/Le8BcfQBnU2sXberNY3qxDUOn7MmxhTxz/1kDSw/9/BagI5N9a89w2jlD
wHdGD5W7NMtUKYFgExdeCb6kCamNIPMHyH7yA3Z1WBJq1Fm+KSyzUD7XgaYIRzdRAumE1IJn6Z5+
p6L6T6ejeDE3uwbROX84U8G9ZFW+jKIde+qaLg4Xd/twqoJlclx4tIM6fPXWlnFIAHEJOOrt0bKK
fw73zbVsbAdJ/yv1IZcArqWEUcMu7BqaTx7QXQZtA7g1qrZTE8t03ReqXHMwLlyn+M70Ni8lLWqV
4ivNiQYgy80138fRlz05dxhD02G8JFLBu908bgGpYBP9C1QmrC8WW1RimYmoqCBg7udgl32GgQcI
xNUNfqH3UnwKWIehw3r0YwGCTpulEwKHiv1tH7A9nlo7wtMLX2oNstnwguvw2Z0MPlCgWsY+szRh
FbnqdiS5QK6TTBxRONzoXhT2zU1bgINHlt+TF+3YuvxOppd+qRJ7zIJzqOoVNhBu0kOp+m1BjzCF
nplPvf4Se4/Mi39mEDTe3a2lshcfhJBT69WFB4Og00PlcZpUzcSspR9rY1iszq19m1FvvQqkJ37g
mTyNPrKJkMtoom3J0czDRGPugKvYaAVuUtk0E5VdJJUOyHbek5FrMg2ZYD3k9dWkvEvstAq+ReJh
HoKz6Z172w7TkipsoXOh52jpjuEuC9/a1bYWm0UzehTvqN7e2g7dJy8aaN5sEVHwYsb8uHpnW8Lm
+I9wmoFVmPvrjXRCZERT2gvFNERCKTJICJ8N4P0ZvqZvzmVgqP13LuoHzL48uowKBGWWMPuk2GIv
Uo7jylPnw8OFHgrv43iYEWQME2ZHqeHJ7BpabVIWkiyw9mUTqtGex+18mZM5WurqDfAp/JC0F1c2
KDNhS9mS5pgxDyC0CuSO79jb/rSWiQg69xeZX30e6g7wOa+JE2G1BusDepiB4z7M5Mzy0jrerTlT
m4nFfrgLu1Vxe1yIEbkdYCVbvxGEk8nIuFQLCafpuUEo88H5HF3j6+437jS3vOLEnBbSBNbTYla0
XN3Y36S0iiOOrBEk7MtSWtYnQMRAjJBLf/Mqqxnlay7N5tm/7yKQqsdRwR5yzbgyVxHnSbi0ZnfP
tmHIaqahpfVm1EiyroZfee2DqWpJuXdPBhJTXkLs7g38fGJTkvxKFEUreQ5S/1JCOiCjs2/v/HYv
Y/CfeaB0PexSh4Txv38bLwSewtm3fji7hwyanyHijwnm95fQi+cIIV8NkFWA2eEPrReJTlHmMvti
AesrYj3sw6FlsaOznHQTj+Cn97W6qXAIcy5fs1Q2o40um4WGdvaOoEJlwjlEVltejpKkSwtcs9oP
7fkvayz1qzjKaTBMpRkw2iYOOI9507lJViVxVxmbfa0m7Q98xHRH9S+V4B6S9237xa7Q4qn0nSvC
ryCvBaG2UyLNC+/dSOwqUq4zC1ZkRGA+J1nxNkJtszk3iMYJW1taqlmYR2iJ1HLXJ+W665m/kvs5
+nPHtf2I9u2gx55Bg0K4pCkTnou08giSjCYQnVcVhbChqWow+uAy7pfcOOJ7NdiCtvgVOYIo2tJc
wmCVQ/xahyHZdHlsIH/x9v5pwSnbcIs8ECRDfvjEs0n+GplhgEedYs3Q70g1Ks5HNiBR0B9uXbs+
LJZfZBoY7bjTnJWTkJj2egDeQJUxIRH700jXdai+6YeS2dtuhK4tQlDTPgc1ttd3nTN7qUtlC6ox
rhb+csBtk2p2ZLBEfz9H+vIP+6P+Y3zmnMkf5oSZo4pFsfkibfmLYkJF7hXjM++zAk8ja8xmr/7n
kflqOZS9QiHXzWCG87CK68i+XilebDoA+WQ264INIlOkItAywuoxI49tcTCAcQ1ICwzSkqGEDsI9
fl02TXAWhQANu7cfm0KBNW5OoxbS+G+nYtffzmRJZK0pfjjXS5ph/qfBNdihdVMHB2ku/qdUyZSJ
VU+tP2bdHspvOWDa+FDuKVAZRrtSS8uzsFvE/5XLTTd0Rb8EML9DrtkNvFEmf3SCMYtLvZ0E5wqW
RVs/9VXM5ouLp5BOJF0yjHsOQNGtYLo9RmOH0882xP4ud0ux8YCR0yMuC2VXVW7nbQ2R7xDlAkxU
u8GmHrj1fAvaxOetPte0II+GG4chXozRJnsepWtpV8uzu1ocyTxkty6MVvbpYGlcMxueOuqbUPdQ
TAKCEJDU8OBh5oHRLtDFInGONbOiWMOhgLDOX5CSIueVa2c06mr68MQDpaIScHNitvpzJq6zdaUB
TMtk+SNnwSI9L0NU4i1cjrrh6V129b+K7/25ZxP7uP6mer+sFOcsFyjwFZ76z5py2vt5VlrK7yUm
kQgJDZ/l0oB5o9io5TKD76PbX17BHVVvZrhoho4ofdYNLKhIX9+CBIx6FR3/CIZ3q4viZYMv0pRt
Aw7JKOXcuzslvo2wDLfY4NqXK9dYiSWLOgiTKaoQxkfynzW5T6++uEV833sMMk5OR5H4b7sU8F7g
5KN7JvloaSGmlWDvxw3WM9++TonzqVWZ0UjuXjDyg8qsHAexNyoB/rf09eFYcm+S671NK/yZxJtF
LLTqliZqSm7tvPzwGHaRzh75UrczEQvHYE7/amuFZx5WvHSi2Pwaz/D6U7OD5VjY7712lfaCY/3f
sxn8tjM3n6bhwwEG/cY7N0NUlL23H59l0hiFq3SXD2KSViuDX1UT3mOVLWsuMf9sbdZ5Kg7uv71f
y4grRt+HFw2DgUUCvqExuyL/HaoLOZRJ65RMslXN0Udd1r/jv3Gfwga2IdS66NMbVYvAbsR3A6uZ
Z8pb2xw71Iybs38bUCiWgSTHEKNfeBWQkH0c6smV9o3y6EzAqLJsZ+6n0tNV0vV9YcpPeprPxruI
WiVKGFOxsgpG8a52VypO62+UiOjOLFSuK1tLCGgaFhFmcE2hHwnLgLcgE1qjYJd+lFIuxxI0+3/Z
GpB6hBCH0wnmQFhRGzfCbRfXoKAKwEZin0umLDHmR5oFWJe23SaHVvQh/HTIGKa+5jXAQQ35wYZZ
CufkhRiDYeTGtntpZpXsQHzr8xdl08b+KvRKLiKNwUZcTvB+SCVMbFqbYKcdPoCJsBdmTiPyiTXt
n6kgs+exipuDdf12sxRINs06KTszt/ZB5ba7IZuTnlP+VY8feLAFipq1UQQJ5udnz5TqkODIMdez
wnMJgkCSQa6U38ZKEFPO1NeQGzSKFr5jYPlFAl8bITeRe/ZKOECRO9YksbPYuQt2ufkqPCi0//aa
lrRe8fXTA60NNFLqTaIPkJYk/mxxhHuxA58bKO7Jl5Q7lKybKsqZI5iov2bkG9hg2XCxTCPZUlmd
wcZkjC4rIsy8jJUyFpcfZ3jzdR3f+cYeBm3gLtQmTYHJrfgGDNJWc7cWcFHX/DFO7O7L00JBDy4W
uQcx0RxE69ozCJLgw46wM3ju77Fx/1CwPaUeeaB1FR7p5sXiOcup9Pyphaq4gPrHuOTWXJiOpWrp
jp9dfWbQj5eaw+X8yv8dMX7zxBrjCPTECPNGI+5wXgkpwunTuGuRuABSKqYTX1LH6es26ZFWPb9f
AzKWCmzDQOO8ekBQLBNjCn65+jjeRPQLi+8glZf2/UtM9KeOZabik8FWyiQDwWEwNoiR7ob6WKC4
1Znqx3E/2fZ+VvYBlKij+83+8JHlrUy87RkCohEZTiJHp4Cvcjd6hUFZSuigrIEvSSxjZrIpkewx
g63j5N1c0XS6zMu3AZ+h1H/8FPt0VoWtkIePoDHbzFyvSC3Amw+BAg81YXUvSM78lNxNhNpvqFZv
xL7p1WKL+4dPvr+hAA0eCvOUuA0dHqgNOnjxeoaW3cHyUdRFnD0d3s/Rhu7Pekbc8hCdChKrmDoW
1s6HhQEwIDab+U52g1CDEEVJ1JHmEa4CYzuGJYx7nMT2reWGxEJHNz1L5eDvCtIJ5rANBZYsFOQQ
rIJEokaOj6iIisg180YfxMhiPHuQlct5hAoufIN8gz725Co2/uwMDaggV1vNAZnnn6PxkQd7kfJh
iWT5FYU1k7DD+PLERwIpOuIb0SFFcQceAc+WAtersEnE83iI8KCrjuuF7KzrAjjv2h6pyb0zYPpi
igtyXD5jHixBRzRhGmAE5PIh7bd9dbvMndGQ2RjZkkSu+qDV6d7dqsxm+NfCjipIf4IE3XQ2UL69
7GUIRn3/VI+b7EY3eRXHIlyHC963CdnnOf9301r6381yEMKGEJBnsykJkFTnto667fnAWQqp0Z4u
NniYUG66as0t4E4acEQdjign2RrUSRp2RSgQqwzMzmM2P3cBk0wt+JzXZfLMaUagxrI14zEKgvhZ
XpxqDWJxyNn5WhFq4yxLXzw9rZxSVOk08BqbhFEhIm7fPXc2/YsIvCqp6UFGP9aZalFzHSywmrZC
gpmzuDS2XD+FEIuWYXeW+PD3v97ZmZgS0fzll8nGKVX3s/fBy9mx2LxMyjKaMKkFnmv/bSztiXWI
vh2z4w70OsaIoiZ5iCsKTQenOFfCC4V8OtX+ZgEVhY8C1JLggq7tq6NsFU68sgnGbV3KN7eTt28/
MF5ZqJN21lY+FncffGbYtZZVQq/taTLxeUM2c07IGIn9lrjdSn2Ujk/pssyhHDWlgRADstPkqGkI
WnY/DzivF621QWh7RiaTJLU5cxo5v5Br48dAGqbSQJcpyD0+cm++NGSZrcxF1ChPe5kzghTEsvCF
Sjql82y0wNTaKt8Uq8Yt8PeX8h0WL/NR/4Q9iwQD8hBBruYDRF+Hp4swQIoX17i8GTiRpOkYrr+s
QualSWH8c/hRTixrwDKk2tRdjhnPvVxUkxWgboHhSmg4Sv35ADMpcOprrGETum1CO8q+n4UMfHZJ
nSVjRw9nfB4Bp/LAub9x5Yso3/4SLle9szIVxSk8Dt7fPAKjTgfIuMCDYyH8WLNaQNREYBcDQT+B
Ovze2e3AOvD6yANfCs4hJ+51/vSLbhjUAAnQN804k0K0E/O9THjgrO+jlU1LYfq0RtslzwT+TeL9
5zhK6VSilDwIq56MlvifPyaoQMX3zXobJsk7OBYyfSXUHteDmgidy1bhwSeAHbEOMHcEBAMX4VmO
tuVWlx5nND4CgZAuxBi2ki6pf9tXuXCU2ZUTG4EEUETn8P/EXLJ5ltb7qesueJ6ODsyQJGpfAjj0
jn/PGYZppkPf6CKWR6W6BnSLEH96Wj9So/y8YfieZBfYMkKGbrbDmnipBxXZgQTkxFo8eHjae/Tv
mwhrgn+lramS0t6qLVk30jISpPOq2GAE65AAPr6C+9rfOWEuAj2Lldmy1TEkKTxqQMQMqEIVQkx1
W9QSWOyvOkAGxzjaEdpX4cXuwqdlEkFA9FqF4MJWN46FSDx8vPnCfdA6GLWUIgtq7oRA+1d3OKRW
OCaO1323AAZWoiaf6Ww8jMHTMTdZyzHiYYbcbnxiibABrjzH65AYZJclKuCxL0dRJb9qYQSYFFcl
+4voNWXLnLa2BgIiPXqxqTLk4qq7++r3BPyJWCj54uLOXyi2ray12B6MgseXvlZT9/sQvS4Oqf05
NPId0KNKf9BYJ8oyYa5JJ36/hxiwE+PE/3MrgIVyHe+GyaHV+1psZE/w55oO4lYSUoGkA+xAE0Cb
LKL+ymabJjPbkrN607BdkVWc0zfFUarvizqJfxL2Gi0pvaom2pnaucXl2oBOLK0JuoOjbJwJv4ih
BTVz1t373jYuHg89cn28ijhXwsrANdSpO+xsycDN5+DmuJ3FvbrzhIAduUqRNhMFOl9P4FqsDHVY
4zgWzwHQrUWh2ApgzMpyHMUws0WuKUpQEqrgOgkJ5YAX5wBGHz5sFtaxbekhEp6vojtyDHRcTu1Q
KUuoTfjxtdFvnLMMrmoFG2EVufV95pg9MS+YNokwTibX/dc5woURpqPHQMubqvQg0nlOQAmvbTi9
jZrEfRT4Cwmf6gaMhOd1IT+yk6Xsn2eK776SopxuTymvDCag7Wy5gP8nHvaMXgQyqXG+SQ+3Tlw1
w5Jg2gZFgmgB4vt4O+fi4vxVLHurbLSqPG8ns7D+3VE/d5nlU5ichoQuOWT9drMJW7m7wgHtr8t2
SO8JRU0F5YOgHQa8JFhNBHWtHnCf3JdUkyPdal6twhQRp+j1uPHr4ufoTCM5+qiKGYnMthSc//5H
RLPuBwoAu7q0AUjveGXiZI+yhfOnVRY/Kx3+VK/Glid7GffDO27xunQu+SxSwqVy+nczYeOZFOXM
vxo1mmhDcWeShju0eITdyYrAKFG5dlfPo8ySvkkzQgX3t8anGytjqOwje8uE4hLeF/r6UrYC9fcA
fzGMQksTPcVrlraE8H6xcYDMElnMbNMmVijbv7gq3NW66MxVKiAkOKZQ0YuYKfRD8krEw9bt4v6j
1nVJ7jLCscEDF2Ld5xr5vdX0XqCukGWdsXz/8HElTIs1vICtzWXNh6ipn56uEsAfddHRe5rw5h93
5K5H9nS4lLzgOHgwFIwJBcVkoA4Er0obuycCSWGfoUQtcFFKtckTZ503tQhY7L4WhGixFGkliA3g
rfCtBP16v74V/HR6WpLK61xbcr8AtqZCWHgEhN1X1t8Xc4tP8onrFYcZuvJZHVOD0v8bAaosF2fN
gF2Z8hy68aMeli1d7k/smpnpeh7Tx5efNEgaMD45DEQRgl2NmUnKHcgaeEuYHV3fNfx+bJ/QRtkH
OkWqVSZidHkpFLDM/zzLPZLorHfE+018l3o17v/vpz3Rs/cKBe1dnwm5sz8YQAFTOwT3FxLpIH40
OuMIQjBLc8VIyGO7DHlRiw0aWZkuGOzWWHc9vjrwbgU6pjadTvmh2SmynvoZZHZmhkAx2TU5oxKX
QU4CCgmiEp7vquxY9GI0aBAm9CUBhrO5w3/HkKwo1KZEOgspwtkvfuKqZivoeZj78OKCS30svIFe
3mmUpz2RPlmJDqevCWgMhON8mrS7l592C/i4DxuYuRDf8lew/3ZhWXJrtDkcMSUriHp5ZS7/7ERR
Yvwy94VHI4KkaKrMOPQx4PlePqi5BqVYKsMvgnoeoae6ooEoqyZh2DfsXKyaBHiFKdwL/81oFnXq
8wkECyD0bfrB5LLHSQNWleGXBeThhWJa/lI1Y8A0ZW5NETHqUwa85euxe2eYXIu7GRWPulurHxeX
85gRUSoOYKSMTtgVVi4K1YUprGZDJ8ZR0/LtxDmAEICiwT9BXfV8Lv/yQYfTEJn8TObQnJ+quEJZ
YhOVCL7F573XgSXPIl1gB3ZVO81RWqgNaV9u0byiattbZjhkgfFfLUuK9181lfqaz1LUbirxz+Su
UGbaYstj7nxA0QP5Ec/BoAK/JmKCegUJ32u/PN0bVnj3zjSRZOv/2gjupfDqvs2hp6dDxPdTL96a
Vmqf86v8DNzFVqetFJgLjDkhhcQsxffVxWWD0ao92TZUI70AqtIOvDBAQ3sXRnsFB5UHOoXDFCMT
IE8PH/clKIDtfN3pBRGa4h3+cfwwC1VolAWyBjXR/sGkxX26c/+RjzFxoCf4rJkqoLXcCYK+KTHb
SpUSmDJrcmWfEHxJmWib8FLlj7ON/5S+TsOclY24XZ+gCmy++i/sV73ak1rVp9EcI8og8AAzlAVS
/Ysw2HFrX0glZBPvTijO/RzrGfxDboTmVFToH1lLt/ufrqPqTRpV7Ar/TIbppkWF5JZXf4Az5wuQ
GfAKloDXuIKU5bjksxaBD1BQ9WwIXHev9zxIywnBezwx6yhQt84Q/eW0c0FACOSTp8BgRViqGz2Y
SsgUH8mtDiod+OpfajSdAR3srTFiCR/6YoutXKKldI52Gae50sk1kixg7is5gzBfrYimQG57gXw8
fygL1fYF5kOtxEM0qL1PeeGuLToAQl7u+XtrA1Yb3c+eQiwx8EgurmrniLnOT+JXK04lj0VBGMb4
AnpQSRowIa6JTcRz5W8LmQ55d7mAiL5KxBP22rGmcQ6KsPtamvVXUNQ1k7KSkcOBXhe+omVaB5gi
mCE1Lb6Pebux0xnTWARbdIZE92JWQnNujlbEL9fPkAeQoiiyQknpiwnpcPIn62eWspSUvjBHVh+H
OFV2M1K62XRTC8gQLfQGpE6TiQcJ7lXc3b9beic23CPPCMiRg+JpZgK8NkXVsXvSGCcsiWdHqcAw
g5WumutIK04Fml6uc6FcEvgou4u9DFYgBP2/NlC5QWwQ+hYI/rrBRTL9DYYT3vNa5BWdCxW+Et4Z
nk3kkKZWKKKct43n2kXQCIY9VqiPKdnMJxoHObQL0IfLVQZjJ1KisjCyjcsjAFBAHFfB9ROGjN3c
d8QEKaSbJCkMNLiYhJ6fxIJHtYQ4qMIHOV857o1QmSgej6Fj/duuzKUR2N0nsn5H9uWdYQf0pSGc
uu4AZ92GQw/70cw3HjsBLTaQEG9XgpC9A8slJs9/pyKuhcHFzM9VoEt0Jd4enMunN7Clt02VsBkd
Q8vfuTxTYkFHYuthMjmluad5cLpUy58CYwtElrRgZkT0xFkgfVDMWGZquEPCkezjIRTYvK6x6iTW
8P8S3sGhqaJMxyMULCoRrtL6PsHpv2ZL0wkhuVmsSjTxmaz1kCOAjuK4CLAf24nfoPaoisyVueJd
tvp9mrzA+zkgtjTPVCB1H7j4YFJ8M0ufdsKyCXjyzvX+mQr6r4xwXwXWf6K4tCrrP4Wpx0/dgEiU
9mbYixC9Xkzp21GWB9Oemxs29Bdne+BsRJMpP7bd4h1NsCno6f3VpXv3bcU1qn9YDJLFOIatUeeo
b2afiXR4314y58KiU47MuAda5MrD88h1j8sU+p0kWCmtuw7H//4Sky/FguMZFq1lyvj++vZF1YIe
Fkf22Be+RXP5jgAnhPQ3aSX3TexaXCs9rYE8ncQY49oCt7TO58GjsHJ8GK+SEo8SP2EXTN9jV4qT
mvPvY4n2HTonTp25rPW/x3xBN/qcZr9+g1kof/iCYcOBRiCjTXmQOJUk2/CR80SnaMsnHNt+s+rI
/la3TloJwOSiQtQKUhQBmGE5vBasVlCepGzNtxmL/0rZQu0F+pVKAWzWApzimccs6ZkWW+XCky/G
OlN3CpeppBNsGCxBMfFZghcGExHfrDE9t2JPc/N8vHOH2iVwK76OMNKwlms0dJc7Qpnjfl1WpwLB
Ox3T+A9b4bESBwtQa+TQH2ivoWYPerLo+3OSc2HQa6rOOKOhjBpHwL+UMYo2B2sHzimO9j+DPkZ6
+lx5W5FcOhrhmeAgDKPnu4lxPEJ84LFs66xFiORoqLrH6b5KJe/yKXvq12IthF+/kh9iV7koUEnv
DxiDEfhdouaWVhlFdNHgWvBjUTJjn9rycVchfwwBcB/IqEC1WdFNE/nwcQ/F2boCA9UAxG5W+Z/v
hIrO1QTvSlR8NaMQsiqa8N6Y6LLeJSH+frrU20KN5XHDTyXX0CNWInkZZSno/Uhmjifw5EARGK6h
gwzgaWjIiSWo0u9ZarP1KXg5bFpwofyjhV4VjJykJ4oAC9pFr2mdO8eFZY3u8pZvqfIZ23ylVFf3
bm8kchMSgbsaknGMsbvPuZNMeLzUwQBMNzKn37O93YIMh+L97YojYgOXCTFrAMZnK5aYbsuXbeeZ
gYvui7gWI6lUOKtCkI1BNtLywvf/HqyeU82/km6faEE5R93oFZTM45hDAkN8WZEHfqRJ5QkLF7tS
MwslFTfpPBh9c5E2M7kPcrPcd+jH1UMgRa1adOyxtBfu86pip3Zj90C9lIAiCMWFbhBw8D+f8cXM
x0JuPq2uThrYS13ICqD1sLOUFYHViLY0exF2JMG7q4FwMLQ0KBDJS+fUtCDYLBFoJGLW0FD6UFe8
0AVMhAOq/KPZK8XL2lbeQULHD2nwpwX5BW0CQdhdKa9xzvGVds/TlwJOrXtwpSl8fm4l8EsNsjF7
3BgZ5ZUO+dN2CUHdKtObRb1eYTrhx/Ydq6A75jmAZotenpdVZ/T3Lqm3IUNx2y0fKPkoQfZgi/M9
CLlyMZG1AuS7tbvPhhmuYQv2QiN/jj4QJ++clpzdenf/8B/JVB4JjuanWbuSoA6R3o0CvDvaXTPl
JVFefyYaLRV12p82yBcDUpt+1iqQ4lU2za4ZoHJMuN5ww1cL3amxZko4I0H4pEqK2wzJjd2wh5/F
MVEh5hqZyGP0tKD7khguZTI/sXLUw0dqmzmC2JvN5hdLMzHwYtJpVrOif+bROjsYwxZ/Gl/OMeDm
Ir6wfvXT45qHoFqiBEbsmbLmtJOTGqcla8E443oeH0nLpHhxDnN4CpDeL0d3VFqx/qSxLhK/53kK
JugkaJOoHTBSWjO8INlORAam3w+daHGurNpoqNX9Szbyzkscn78XOh8iuXxaDP4U11VLJLhaaFa4
3ddn5TT0b0+GoRopgNQhq1hc/905aC70Rx+7CP4WPQbycLzdseqGdsF7xVq5Y8+19MC1bewAo3gK
snsNb9FcNJavkCC3bSNgiVZtpVN1dccelfImBkLkr08vo1l1F8pnejYRHIxAkL+0/YyiQV0JQStF
0Bu3Vmc1JpJkPXMsncC0jiDG7GPtHsP5mL65+/nRd6jb0DpowXDOEbNsvbhQuOKTm6DziwjXFlEx
yT8j5HQGkAO1HYzwT2TMS/RYD7u9E30jobaEVFgAhNtolZSlRRpZ4Qv1xWNjBxrzgXUOBCgtOLjT
fa4DuNaDH1GFSjHf0XFPMdstAxWvODVJ5WpHqYK10mqwMlY2psNJGmS9MDn/aJu9YxbDxeQVARNl
st8z5Si/sWjtiNu2DAW+0JMmJ1hWd6IzR0ofkHShE0kdbOO01XysZ9WFTQDWSEeYmOdRgDt6IV+c
+e5JycpJXjGFc7lQvq0uCaA91Ndommt1XZ4Ivi2VZKq1r0FPijm1x8olXNdR92nAbCDIA3njM2J4
BuXMjd4cxy8MREbhjLKQV197edQfS2VBsVacq661RHOpTU72CzvY0/yJJobEEI4JsuQGNWqEts2L
H5jD96hdgoYgzLrBZVdqfPbb6SEnrmYI7AB+VV4tKX1luAWFHebXGXmhL0hjQucqzpCg+q90F7nK
hFhdCjri+aB+X5FzBQGqv2m27BrRP0grGrsGAmIgDR2M/1ZlrmwWtIKvb6yAppRp3mDAPXs0WxlC
oJbP51WzNJLU18pMM2yltzwvAAfLVyGD4nDhdGOu8+wszwu1vv691kZf3HDLxrW0DFWTdAtPHM1e
EuRhuGCXbFnwCWGwS5Sbxl2zA7mQ82YZCX269IlZ90qqIrrha5kSUelLQtPOe5rnJJ5IjCyApy/1
cDhXuTbxdITOJZEEO94+ol1L6Z0VT+D89QJ12NF/VK5SoXoPNKUqwVTHGe9LQHzfQ3amPiC9/zex
5Vn3bj7XpY0se6NZr+FlXMgbbxaU9nUxLHpsQaQm4h6R2iXe7z4dqQSLq0bRntNI9VmQnHVt5nFR
lQ6EVjeRY5oLOoCaZKzGE+ZL6y0u/L3+eYTxiE9fz8Fprus1Vi57p7rrthThBS+P8g4sK+nKZen8
fJkcTcBLnWjB6uKzw6eR2PKCDht142YO8G/J16WFBfo1nH7CoiV77R/EKAoNKXqe25JH+wHLQLLO
DKRXkuTKKgwvnW2n+2ChZ1k49UYG3+R4300K3fHTUyovjUlAt7HIZ+Vk2aWgNoox9bU1VPeqGboI
gP61sMmcx0Wz+DCHhu2WkyoYixsAB13v77v2k7yzfqL3TK8AW8MxfnXYJdGK0ymRWhFQ0KVXQJlr
RDFYSqvmWq0WTxcssGHFdeCMNeDd9qKjq0wbSU71sT5ahzPnc44+9RbxcZd11uqGyyOM2yf16Xkl
sVdBMf2vxCbiHqMalf4cS6ZqlYpuSZy8tAc2J4aGE6BwGMbcKUVUrVvhC2cwQdyhkeMwN+a4IGmk
LHef0KXWSy8U1RcQ1IfbeOl1HCpN0e4UF0M8Pqr9YQ5RsIShfhoqPoNW9Zual36F0Xzx4jzDpDsU
vGuxQ10S6BUF8oo032bgzsjEPrkuM6cji4EYl1urD1EO7+Zul7LQur5RFrpM/yDtF1scAYhQS1Zh
eREDhAazpMWVha3SVLl8S6DlHxKnWtr4HMp6uSgj3FTSL287dnO0GUVNYywV4gqC0+zhi60RFe1t
NCxeRq4hRNlZiHz4BuRlY+odfKpArM9mKYtshbDlRz/TRh/zQVjtj2cS0w487QQK+ejus1nf3zXw
BfSq24dIhRAw282PrIBvgABD6TiC1VwYZ6DuG6FClQzi3sm4wCBCOcGYEMACD/02y64v0bT4RFNY
1uAbGzjPeegMENiTRTibfKZWUuWOUlRPyDoSbgHIhySMOMo9IvXTIEfUeuMNyjeYqrVu4BktKWCf
iYOwF6ZojSsEIy2j4v0HT/oo/dteamjgH07S2BMaWpZkEohmBeq7oXx18Ydyv0bYsNKsyxkpgmTM
qokj8hXSyzZXq2Yge6WHkUyOcl6c7p9Y/DT2u6FjY3MFhcPxduA6M/Fx333kiIaa8mkQ5GNsPIcY
HRz7kRk04B+4xcVSVSHC+vEFzwjJHHAwjk0/rlLkQyMeeUfOun5XlsF5Xy/mcIhjavnN2tvoTjN5
m0GYJmAVw0yuqLn1OmbsR5TSATewsLJ4YMuuDil2rQz8EbBUOEezmdyXHS9nv3XOYaag39KgOCs4
9pwQkV+EPVQ+6RWcsi1h5clEpnwhvOflKhb9Fa9NzGieRnGbbexqBSO4H3KgleXXAEIWOB//2eYr
PY6F4xAjUY+QtvCBkoe1TaFQs9xa8mLXw8NUA2MqKGzc7vMGt7sxiP4gD1uxZkJbNFY9YKZtjMKy
HuzV4DLBQSOOQO9qE7a4YC7ycI52j842utGQFpR3/isqyUwo2pBG4skNAlP+pKaOZpKf0Ks3EQxe
GC8GcO2fnRKXXrN2LUsZDzLMv9VfKLqzkw6U/loVBfAzjAK8Kwm70K5kOaRXCu65stjImOO49SXs
Y4wv09HCXl16vLooMxRWNKWbwKkzxPlo/uTfR4WJ/Y0HL42aKa+r8LUMhE6LpfqFm/aKie8V/4iz
4PlwhnOPJ4ksd0u+7rd7mJeXMsjWeYAs9EP63/hkKews7d9fTF6yO76KhcZRjFki3N24z8WCE3dG
T9/XkQ68AgP/qekCaY4qPNrxoqVWmoPgd9pRFLVfOcKdM3xYXCq5eUp54k9Mfp7qiVHglHutSHox
ko1KjKhdUgrf2y9tWND8gdKWXi5yh8QHkE/EeuUSMkq+1sPJrOJsv/Dy5HXoi5gcm4Bnfvoual8I
dnn+1UzJdvnPIzfTHbEiaEkXP4HD7Wf0Ijsgu+qYgbJbhpyu73Qm0nTMP2u6MYdPrwrdXBqMnr2m
1Uqq9nSV7O52jgsrYw6kNKMKOv+dYLV8aiY8LzvgKxbSJN24jzSOYFzt3V82nf/0wIfYS3snd0Xy
J4olg8CXIaWcvBy0abbMYtvTQ19ZcO1M8TR7s2qV6hMEttTGaYjaM13OvRllDdlXA+6/fXP0fo4+
6CWc83mPv8BkPS/9WLdvdwDperHe3LSjqRul2s9HPTHxGJc6yZ1Dpes4mhUJOa68gHngDufFUxWC
uv//JTaNxahvwunvjNQXt/8QiplDZPjAmWTOf6IOR9F7aeXmP+aNfV7jpAlzCWN3YstgjMR+k/h6
y76b75f1VVLg3MoML9jd352B1rIe1KCF7iIpUVNSSXX+5a4BkK2ajGMXXY+W5eL6dAqGTwM2VIbY
bpS5bzzLGOMuBYr9GAryGFZMgC+WqHrs3HgsmvgUrWWzXk6nUcuXBsbLYlh/ujtORLClsNgcqUAS
z2RcoUznZyVFU1GyrssJqJFnpaL1JDynl4Vy1jWyVbkPkDseA/d1UVsU2hBw3QEhCVAfkG8BCFww
AquaExgaK673UWpHg+TcOgNEDln1j1nZ7PkUwHpJW3sEK0ueqi8chYbomcEQd5OaIawyUh2KY+pW
v5H309mPsTAWugIKeHkUQk+IiJ+63buble+CHxk/JrubQEjEQFSOy00uQH/UTQU/2CpmcuASLe9e
QvL2gzWGGkd+qwuoSvv2JRNpTUUakAOEoiMG8zdilOQUcGz3JFfjmGRPNlZWZarMCqsHlFBhTpLV
KWFzSzZd4m4be304d+vQlqwaWn07wjX0b/gnmGpNVsh55YG2SMZ2pkMrKzWqpoQ1lYBXBhtk9IUn
iTs7bkjbmmuEqqbcY1V19muto9/2Te47IDWnI6a4pG4dao7Z4jY0NVhizbfdlkYKZnxLpNnzgKWO
Zd/NQh2GD2wZitQNQh+4iTuuEIDfaMhxp+lWsH3ztSbNEG14v6vVVIp9tUwD+BPVEQ9QLcolHDBX
O11JpqE6UOpHuzDsnooU/x0DFwtFRe9XSL9mt5rJ4eYpnqndRFfGbv5QkbwuQ9hSF/3q0u6L12OR
eoOrCPMDA995w3ST2kOsWMPi6QdIBEw2e0cHOUUAPXtP+JKRg57uOaKsfocOaSF/a0L5o/4NhKqK
MZxIuJ3+2B6kYYs2V8BWCB7g4dNOS8D0eKrXMO+HiyHpGlA4K+RG+NQetgWlDPHYXMOZso/deuMQ
GHVJJoqekjosBxF3MzPmcNm6Fs4DGdGvkwqUEcbL8oWKKGeOjNNXHon01yGsexZFS9YzkcdcPn+C
SMOpVmH/GHA9sI+X7vp7aR8gAc34+iQzZPstb5TmwVHNrlhtRIez6r/gzgr7axZI82t2ker6MRz7
bYMcZDBLkfUimDyPK5iYiYMHtcsnpmoiODznJ+FNRuUT7meF52Qp/bParLO4r1PYV/X1ej0PhCn7
78WUftx6oTuUpbiILeHOtGWFfKJ8OHvsUoCPfJnvHNjjyTePCsmjzSMauPJylxHCoTsB57vtPMPL
ZfEDUmiPYM+i+YvE4WL80zBL6decb6XAfPkQI+0REOEIKFthZSkNbfwcfep8EeQcxMKytCd7ifqT
rVHjOW0zH/Th1NkKVZRnVarCk4s9R3KvuaunNwzfIPhoblkWCZAJqZXVEM7l8+nYG5AXAfbtNkNx
coy8nRF2xfM6mwMIJbMVwafNV/i1kFNnzIV7QEG61yyuqQy5YsWPrz4UIq/KSlkuh8LzU+b7S/ec
//Rcl5YK4vaFJlZUwiCBBTreI10/S+u8R7/P0uo0Uax8QbnXrWwZ/R+OL5CM5YiHdpwmYn4Sfzja
VwTsahAhJQmHTrPqidHhfGacJxiEMdMOBykMLCwsol3hVic4Ek+doqSbPovnREv/80vR6j/et8j5
hnKNHvUKjN/+jUupjvY/eVzR7t+7Y17jiQCGmKG7y/mtzuMaAYYIcsH8LC/j+Kh/3SH55BWzIdnF
8inZAS/Nzdfo2GKWrDwAIO40LrTnby0VlhfshChrcGhuKzsLTqMs8XDiKqHWDuuq3bm/FF7Ra664
AePPrE56CksLsd30WbcEdX4jxhCVPRQxzUbQ2iCFvUb8alAP33zm56gmUyQI1Pt1LJJuoHd2TjqS
Ms5sioXSJiQkjsospY5qg4x8G5pDLhgwQucTrBxg9L3gXeXn81mQ/s2v3WhrXx8sOXOuH5k2CJya
XgzIuqU9LpVm6kfFyDS82a71UTIXEcf5OgI5wafqHKiyxYGtM+SXFmKwkD6NbenXAmwuIufuDSbN
jjWyQEd+ptZw+hhlRx0oTxoY1eWLCQTiqsWV1uN93D4fuqz/fkZzQp3oyMichDbQgp2PAANZWQ7e
Kz2eqfslaMAsObABPQ2upNpK8kualw+Q5beDYR71jsXjuJocfleOTqv33THkqZojNwZ8eUJ3k0qV
H8H74ThzGE+ObybKkoSWxU98g8urIeY1U0+XCy6Lr7g8xxfpSfGpGREyZlrf3IB0Kqqhhbo9PxZb
CEok8bUDkxRx1ItveUQI21F7WnxVzGZsgOqziJ9mek9d5gcrY8BhLM5RW83fQw2o4wM0mfZlvNPq
x/Z5JVE5CVAxIuAGlmZ+MGTfhwa6BzA2pihi47vYD9RBOlI8ZsTgwTMW3HnWYudeFX7iv4GOnR7P
ZJRd1iXPEX3XTTi/AexsXc7jetnRPUG44nbc0CzPJccRoMmFY8AHLUzJwSL8/EuNboQEFoZrqlSn
wWQnRuwDVf/i2kWVC/j7SmFBJmvJp97PiTvuRO9kuzoIKRTQItO9oCvlxr8Ee5ELs/fYBXIoQ68j
mAQuhackEGKEF+g2iEdS8OmIoaBjtZxqgFpJpFK5x/iQI1KYjb99eaYM9oo5KKfYWCEJbq7X9Q9n
6MKSx7eaalkkh4xFmo7SUpQQvFthLUaMgGTHZqi5Z6oRU6/ao5qni3s44gay2efHiIqCjNUmIPrq
BjikO5LYlBuCpoTz8MZof9uRiWNP8MLcbFBtznQvyl8KewvUdcWPSTtFF+uKjABZBkc7yaFd1uHk
M0eNo/mtgnp1L0q81t3JAPI6EjxDvguFibig0L6UH94kO6d8tWHWB3kD2gaL1ibk4lovG1HoJtF6
Y8LPJiVt62xsbkgRs1z5N4lWs+DxBKLb2tbsSpQ1MCFnlv43m70LQZygsMoXspLHLIl3/GlpA/IO
b9AGFvOansW56majOvBOVed8FuqeTxykG0/6YcSNTAwtnjZ0UApMw/xMEwsI5+qq8O1CFWdJvnqn
Bv5D2QNKR+kuSW9j+6Uxdf5pFe6B0hwRqrit2a3A5BNhL6L9PBa3IAjAtbEVhQjhSRfFsG015LJQ
cpD2VMhtJ11WE0DzeIiWLZj04sTYqb1D90z62tocASLsr/ykyVt/BN+rruKyO4DyXMUqH6vJYpcV
6TPCC3ExSV1bmI5I6amyI5TYHOVSJAplswqaf93EDc6Fg8bQlEYrFIIM2YJV8IOTG7gFfcDppahw
IfUu7Hq2TL4RzcwZITshrXqLzX8dg8Y9atc6CpZ8jZ1rk0CrEFVhxUkKv7qAkF89oRmzcEk/ZZtK
3JJ2fD7alwYIGQ80NN+VQLEzLs+mkpl6WmlieJQRJgm63jKg/UGvXGn3oR5rS0XxrmU1woUpdLyO
GK7fOvAtJ+zFeqrqGBUq1gNGtMa6gYgfKO6OqGubbWMPjfBmnpWx+pu8/AJjbzZh777uvqBVWYgB
QpvFz/jj9L6SH7b1JryuCn3VLNN6KQC2cfKSBxIo6pfz72YeDd8YQ3unMNLNj1kupmA97hTYsRAi
CQDSnbA/F5o7ypGWDZRmCJwBS7an13ZctRAniM6H7NSEfgN4QgwLfSwptFzJ681DhnOd7U9uT894
0TwwyYqEWL2yrzmp4KEmnxvlvCncCpdh3OpXViA8WMDp5t9ffGL+v3qa3MxeEXMCzom66YnLyt8t
28AfssL5C8oTlaGlKtVTDBEX2QreiKORY4sRULNPjpFjomle59kVsMmm76fR30QH1LbLOEpPfdbh
jawswQyw/1tzqDW2hYZH+A6pTprhriTqY7nl/mffF///fiywps4LJyQdEGq6fP75tCCCdbdgQn65
9CVcAUSrISnhjFdx6ykdTuukuoBFzv/WgAWRQZMUzLiKQLsskWfbVoM0Gvp998p5AMOpHYt0WAI7
+iIfisDULhBpbbyXYMDYwLYVcPbC0yC3wynontXUT30tUA77y9qcDJEgD+elM1iWo4jDn//IUUkI
kgPWaokudAsddLKKWtpR06qstawH15+M6gSN9mFTyvupb4Er2BXtJLGVPGZKi/cqW5c26s2D2DP5
tRzgShudumW0ZsO0g7bRoWoPeIZpuRwrhx0J9hoguhVZF35sX6QNbtt5TWnrQc94SmR6xq+6Yha9
JWEat3QhbS8929Ntz0NIagwuiqB7/jBtMJEYCZBRiKEundTJIwc09yG/sjQ/Mtf7VeB4s4FQ+k6F
W4VmFMe+uuAULoJFZWqy5VX/WLn4SUk1KXBTccbyp5jq/FR4t2gt5DR6GroHcudVFUjmXu/U6121
wnAlvKV6Ey7P4+IiAw+DoSuyPBTUdYbPtZBugEN13eEUSN9xswRUTqJIwjL4ly8AG5R1dJlgKiQY
wJ6HDyBXFKgl3cHat3FH0WY6Ax7HIlaXmc/GDKL/WblaD1i+Cvpj8SqDQBtl/7z8yZ2mfwUH4OwM
GPqa3Pg4Zw63FHkBE6CThXxR10vODvg2w/7UJInKG9NX6YespoQ+yr+zgq3xT8ZDFE7vH3wyAcV/
TH3TUMKhUaArAtk/5rTmcm9v6fpex9jhuQmSJaOnxk2bTCzTVXiz85L5dih2JLKRO6uGmptkjOcQ
ysCAGAFouwxmAOBahSWk8QPSPjkYYhd73JvfpjB3c6RD87mYHF5FN9i62/N7Kv47KwIy/WqyVvrN
YqcjjsrZKanax+BjUHudLN4ihERx61ehOGsQyY3EJyE0sVL960ZVfzrNQCkuv7SyOunqYSHnH5w7
/9aIQP52Ymimtf0svhvtTd5mguh4MXw62o2UYqkKy4MBziYd3Vf27PcKHa2OBtuchZcFHBDCn/4s
uSmh1ZqOSfIvs664u+q1TZo6aZkRVan6Dz+WKAzfftP6kdIIve54PMkFrMathA0FwLMWONJu70eY
N7swfxbXW5wPddL6HiVEyB2KEtm/uRF4HlY5HROt5dcdGI8xV1Gu4G7xSNhC4AAXOhLPdHEn+H12
JkNCiT1xZyPtbO3CcBZpF/i8beClaTERFWZn/jAH1tXaLCy7u4SyFrsnd+JI0BLwTMvn9tn/JXj8
zC/UmOw/IPpLfgpcExO4aiOhrfnNcDuGM3T4cASjoNtagSIzYkJM8E8qS4qAQwENdSPMtXrbJBiX
YNmoEZAwO/DJZ4YXYcBw9JAunnNHF23g5GhvcpRHRiV5+wyHPIOgNpwgmxl4Dbxzb3lP8SAAhKJb
0WxTJR5U70rLY5OW6EHMeE52doWTRBRDq+GzhpVPjURlw0r4A6H5zMjkjFxbgVSrSPyQfG7ki1W7
amZH5P6UZoZPmc2LwihkYE7zciC0khYzLaGjmJPwnNDVkLuIE4RD/s/FkhBhIUkhcaUdxAfALO99
zOJ6eve4RpiLq3ldFSIR5zu5W7I7d4kXu6l2jBnOPyo61SkA9/A9gFK/GkVz1UVeVKaInLLtoW7B
g5dnth70to6/0SvQ0UOAeaMwcbq4Z9ut0Xw3zqiIPXC9b0pF4cHHmUmPwm9XcRgm6O03NFtwMw44
O5rAd8QiDYylr0k+Hb7oZaKSo3WhlgXmL57l9zfEzvwkYWEWbRMTlMWecq3QYBDVzTruxtRlA09y
2fK9sk9P3/Q6cwAH6Cnv+SSV7G6HyUvpo33XCjiA6hnvbhy0W+YebzxMT43F6jvrdZrwxhy/LQiI
5nKBeHoDLj9pF8XS5fdwpylOaZQ0nSqHiHTWGu6Mnei4lHYlWQB0vPviJGCRP/49qbZhyoEFbVi3
a8qZSXSDOwiVJXukmARxpArlBRY+MCy5HAMNmmSkLsbCFomMl6sLLS1zMjGSY3dvWDbeet9pPM+i
Sr7yU926avofckiNQd0jQBlU3/pf3dQaOISPY8mR4X7Z1XZNzUD4ulSm5QKv1p9l7wkwkZ0sMcO2
3UwSm1R4tAWIMnixs/clCGzOTrtwWxR7Z93NmqBKBdcikiKOIKsziS8ES8sgR9MQT/nn/Ls7NiNx
RTBi8mez+8s03rt5CoL4sLVDkJ6zfVQUUVTEOjTqllv/lWxqGBA4emF3ZjtDBkxpzabs95xCa7Mg
As89ckJAm1S8zgdjx5+z9W4/HegVLMk4mZvZbdO8+MRxaqfQYDJcpfIqkm+V+UslPbOW/DXcxrPo
N45w5ONEMDSK005qQ7IpFeQfyFVhQrdBVGizNor4I+NJoOBcbxxK8SU4ZwKISJcYjLlO5CZs8uTz
UUA7TF8wnsgSJNpVrqj+O7oGvqyfi0PRyZQNscEhDT8gkhjmbVMCP+q6Vqy4dAKsyqLcRIKWVCVB
XCUdE9/yjE3ylOjynCyAJ46vAF0ksFUxkgiHyPUIuzoUk9z9+eW1ojCJ8k17vgl8ce+JpmJsupRr
OIOckv8N9aPupkJSOpO4Jr2/vvfGEKPPYvOncsGmQUtDxUqCFWNlTa+ZVynU0dExhhqcHhi4VMbU
jUe3WhRBMw0zr5xUwrDcnAIrApMyo+ZvIWgZUrJCL8mKPWGs31oMTWJPw+KQifM6G5iq4c721bNE
affh8JDFV9fCAA/mSfu/Qmm0d7L9nwRPd+XCQNo5QIbjSDqLJhgv+GlAYTbdKp4JnciUE5Lzq3WY
pMElNPQI3GAe7JVrY2XUV1ck6OwD2J57hdDJctK9Sha+Xa3qzeQszHzsQnrGGNcbQ+nnT8lSWDMt
WPuBv7EJNwbpx94c+fWchsNozSnSuWNjnTyWUBDhRQVAOD4l+aCLnwmS4UqAAM12I91fAM0mmTuR
LtyPqTgMKau07ZxrLizQv8d5UAkUvuOZmnt/8ar6PDwDEaSwdYFf+7ALbrBi3UKd8a1/YMRWGxyT
RKK1tV8wG0NAavswbPDhI2+f2CcRRf/NgARFuM+x4REKfPMbzLeuEeHyuHraKm2IW68+hX73MxL0
KAeVoGjdVDg7D6PadLvEKtXGbndOs26SBi5ZdKq2CNqTG5ZCqNOgh0RaiY3PwlyovaPpfzshpHs5
jGU75BB8U1AC3qdzCnOcr4G3fwGuZuOa8x+40UnKfgV9jY6KDxiWZSwO14TmNNwX+I8ryzMoyiYw
y/ZDTODMqU17uEnBvmw+OZN6ILdJt50lukOPSZ2duJNiD+WGFY5+U2pJ40sqF1WXbaP2yk8/mlVT
j+BPEnssHSuIgpF/xBp65UmQPjG7MlwpxRza33zczFcNdLtbNWwlTHsbr+QqdUl1SORNFLJKJByM
ebRaa3KyGBfMP4Tmy28t0JtlyUSyyNLZ1Cdq07HgO181hlmNnMikD7re3odBfCfP8QOAy3M2r+je
5BuWTWKxi/5GdB3HEAe2js7iMCrgqQr3M6KksydfPQOVigNh18Pp0uYseTOcs/2kQyD9MSkjeFM+
XVW4pVUX+e542BIvA1fw8qL9kgTXjCYmzcEFHJ/Oa92SBaMFDTRDyvw/BjTJS3ae7slMI4E6b0+v
0k3C1Sul7u9UOml6XkKEViHGLykAJHkPJwu+5lsKXKDUWL8XhiHIKze+aOw1ZTTk82jlhKPDERLX
ADxLsdNvHB2lpe+N42aQ+/pCkoSx75LxKT2mJAufIgH2MSNFrx0M2ZLSFPxIrHke50UJkvBtmCmg
6YTa+mw0midP0hVn94QSZL6D0PeMIHWUXKp8/TgtbPsSGK9Gcn420H5Q+7tyipF2MqzJ6y7WBVh5
Pb41I25Sl+NI9pjVWAvOrq0iiBLYmsyGl3f8tXd8eMdPgaZFsbPU6ftuUbZ3VOwctJwWD1R6q9jV
2GeTmKGcaC6bv2UcmHe4l8RFA3DqBN/OFIj9yUo3T0RKyB4eMDarenIeaaXqI9lF8mZ94PIOYpih
odLp70dQ1kvozzQx4Yf9duBkW++eSRDMpXN33/EIkHJ0yHME8xgsFy0v5Kg2CoIjwySaEC8FVFYK
MMQ+HHm87pfkr8+qYUM5vkJEczM0yxbCkt26RUCek+VyH/oqEhxdAiH/gFldTtqeAX3IQjSRizBm
L39+sEEigqRGdCeABTQEBBFxGDuW6dBWEkwZNiewMe8FzpZaNSQ8sNsNG8Fqr70lKHKAvuek9efm
wF3dMBVBDpSaS2D8Bylsmu3QQNxg1BZhE2bg70EYHZOJLPgOLjIMHN5VJ8UbibiqIftMR7Z/aoBq
XVroczqNiQh8Kyv7+sI4vLyhAlxcCckHzGo2the2Z8ROIZ9+aDNqhiDs/ApK85a7t1jB4TtawUc8
ySKsGJLjNept0D+cTBX+hsm+FmYOJwZgaQ1xLbrI2d30FJVGU5Q+z1RLg1dmsLH0weAvr0eROo14
+PstM6SEgMeTsKAnew3FA/bY3tcXDM7PdbPlfEeg6Uzd3W5Pl09ig2QqanQ37AvHBs721vzKpCYp
qL9jgX77MWu6eESzKkZqh6TMYyAVFswmqQojTBFXMeiZ/U4hL3yJNNjBByqLjKCsKlAoCoRL8Zuu
N9L4kWLH4UN7aXhWJ8ZMstCFcUvcKf+qYvszfhw7JLxn39+Up2FcV+zLbNv4Uqaz8sOtP09i9HMM
no9rqM25n7LgmmXy/o1flgoV3unQGfq70eoZPqwUCU7Srh8k/biK4R0oLyrp38eu0HzEmNGAhBLN
wFSdLZBbupLFCYBgIoD1vi1X1wWhASvP+SMmIgMxOWHyvK3OD0I4SQGe2uNzSXpAdEsKcd+B6VEX
LyzG76phch2vtYYRCQ5rFWHv3V9TPoLfoqJmI3u42Rn6wBcAzdO26BD0tiB4J8lpbSWcxm+f2JeC
PV5oYSouNA9bTpwHHo9K3q1IjdQNfzrxGA1UECxO3eZY9YVZh4HPGTIHafcV/Mgw8AXnhnPZmRwr
pncRvN0gk615cmEpCj4Ynq9VNWa5I9ixcftnQArn5Xb8aP24QwsOPECnilyjhR06uGL2TJePIn+r
TerMlUMU8SuftN7w5TOaXA4G70cr1BT9yt1x73V6BBeQY820ZHZ6G6lZgqpJnoh34jl5c7negfT1
O3+FpCm10IR5v2WD7bEiSiFd6KNhwWMt7PvpvJecVN2kwLKC0AwY3lAqDHfzDWSEKqiSa1W1XmHG
ftHyO2lMgNfppB2d4sLIkl4bi1QbUTpCW1Jo4HRTtd1Bi5MhnxUKnLHTM5xPu4Yaf48sYcgAo4U1
utZayfkrR8Nli608l4T5lxGpI7IAnKGIbXBjrNZKni1q6sgLVC7d7DD0W67mhZuts+XgNvcxaavC
gCpir+i6yYFW3bSDVo6jNtltFjQ8KR8880e5mCImpbSOKdtlwmz35U95iAuFY1wy030fnD6p6BDe
nSOvCpoEeGDLjJekGS2z4p1cqNlBE+PqplOmhQQjoXaiZC8YXh93GBkDgp3UxaRqGU6G9GJO83W2
e8YK0wEKc83uM1wMMbq+dmXZmIGn/uyfFQXtpFFHW+10o+SlssyDiWVPurbLLD3aZJpx5TbhwTgF
hoDGWbfgQ7Ea4z/yK2ac1D2kvyLSMzgXzmsW+we3S7e5wD25hfAXf85C+qpKxBwgLRAN34lpcIOJ
poiPxIq8Mg09G7X0P5TpF3c06zQ7iXaAc9r8Z60pbn1wQow5XkV+nAhNX4kAYmXIwRs/wY8Ptxx+
0Iwa6YpKbjIgRiJiifIaldatDVmiqN6sf0n+rUQuauDL1FQ2Vg8iPx7gNgEK8RgUOegCGYVq718S
6lzFBnve3WufUGEU9oc4cyUXgzUssf0193Ic9llnoW8a+IoDekiERtNcIacFpcxdrHzqnE14HN8R
j0KNQ6c2KfrRYBgaC5I4WNgHe8zwU5F7ByDzUP9jEBMeyXbS2y4cCrbevhBw9hsQlZdAv7iFuVDI
jisYBY5IWU+fhidpl84sd9jYuBmmkfIDP5SBxEIULgY52VzXiTlWF0ensAH7HF4Tl9RP1PW0HRUJ
K14ZhZxJhiy2LlvUI8NyETakfhj/2vSdbeVP/VcqctDtZeHjIBDkkQWkhiVjb27BrSNIH7gef0h3
Bow60B2JtOd0jaHalWp3Gzv9wSJG5rUi7hlaoEesERSg5Mod67kiM9IC9KQfpCCijII74R+U5wK9
HADxmmekBetGZPob4oqT7f49vITY5lUCKmsXmb+dz6qjHgCeFZ+sPhDLxNkwU5JQJoLaLMUHIT0l
Dfw4ZYcGTEZdZBnQy+GtW4ge2QKkqScJn+U0VE7jA7yhKgtIoBmApoP0gbPMFb9wnPIHgHKB5yJW
+Zw5+yNJjowPwPR6aj6oKrX5vsNr0s1Ent7Wt5xvY7qrTw5sJFz6r2v0XpiwjK0V0lbifDvXvhSI
xzXn25cnPoSy2b/axLxYUZF87uI/OP0YVC3n8wOieteekVwXk6cF8Ps11Echp5SBgQFmNUqLngQi
5iPcXAfJuAd37/1cX1BdzWUG0eDhz7ee01EFhpNqjD/i3DD6509aBr2SAGAvJnntJ4vBcnl5Tm1P
gsbjGMNitK2bZRoHWZYPofXwgafet+UDExX4H7svTCzM3dc2wX49p21tGxfnvymapXROO6sj01pB
cEmfZqameZW8V96ieGBwEO6lgS/X2VDfWWPuyz3bG0jJ9B2cUTXj7F9yizqo2/K7IYWZ04B6jdTs
yW1Omy2s5pYmuBua9K1jyTXDyquK3C73iNQXbXdYeERRuUoGzT7V55+a/LtQkmiVcVu22FC9X21O
vHmxFKE0Osb0usMQ743gw/fRteWrxNzSstZW6cWnYi1ZGwgAR/L/T1TCWnMSO5DThewWuKRxAajq
STrvj4/adbxO1MGTt2CieJwQjIpIVlO8NuDGRgUpsmFgiHdysbRwbtwTlt6hK7/6GPMiVFXOwtxJ
6nSLAEB0I5dMTOm5UjQNqhcWOl1HTeowL2+lLysY2PbdfZ07iZmY+sf3BWO4jqW/4KfD+X5pPV9p
RM+JkKD3+2Bs2LBkwKJEBBI9s/Tp+FfZ2FjsqKnVib5PoV6unv3i0kptbGY7d3jEStYC0y7j5ns+
0+SZC+XjlT7uY23zNEUi2x4bUdjcjhmUFCTfnW7Mmz2/mBGGEBwIinLMLXt5SwpwlgZSEohQk0fj
t2nbdePvqqRNaSOSbiU7mMxDnk1ZC8Roj8SD7cLvER+aICsgsThqaduzU2H2nqoKgNUhJNWcJ6ZH
DLZJPs/frXDxfTVAfMcgyHbC2VnemNQEKOSXjJQ53InM2GXLN0uYR3BvQjr1TjRKH8ROkw40MUfO
FqFT3dYWCWZ0k7YFNairZnDYs+KRF97XXGovQS7S6/k301engjt63dE1xrnlFZODKA+DTNPxLgDW
PnqdTepYWhVk6ACn6w2PXCfa5CxExbXACy3VD6ML0XP/bTj3EFz1EK+InsSsT5xB0iOw2EjHXOxa
AeJiifbm/PuPIoRR4rP/v+M/vPCZ8UZAHFxK40rQqB5EIqCQl0dzXSOpYYR0cKd6UWA3zHS6A4QP
eemBQMqR1DvHUCttsH5hCwESTISOM/9/VQOnA2IfKYovISqEADOj3wtpGfArT06+gvCDg/guNECp
n3CGIrgcS/WPTeTckAgJDVVKHIge9iH0Hx9AR9PW6VHM2r3JN90aPmIkgvlBPvYp8kkxeo9D863m
9EK9PELtI0ds8hYCQDpAQdX0Hd/zs6J1F2ifGfi7yHAxoktjyE/NfEXmYdzfwD98DhX1oFrxh0kp
Lh7oKWStsDLkGmW6Zni8ekCKCAsvLcKhomoeO+PyRyoYHxYZsB0vmlcsjWEBKyv0p6/f1BYrXcH1
sNMuoSDktFExBPzaFtpYdn4652Dz9J5OvcsvPRRoMEPJxl66Uem2OnvVFKl6FmJjxablB9GCOx/5
3RhHZpIGh9Lc/XZrCxMRXFVaTEIPSAOEf+laErBvr1xfWMdBqwSGl6KM29i5vtUrNEBrw9m4kqIr
33FWzRXSNwnNULXINLEqon8LG0c8pyuJnbumC5YAtu8+kK76yrRL8XnMySFIWu43NJQzHGsQ32B9
ZqfFmA80utWoW7g64EqRaKs0pyyrrYe9tj/EVMrVEehzgEa3KxtpwmJ+OIMr1IP6ISQItG9xJljX
ZgQqdYHtzvIqkUipgyz24tExJWWsjJNp3rsBvYD1y8cIHVUaMw6wlUQDuyR9AUfmrI26yiGuRk8u
Bt5K5NHFUIDezOp9KvNsa3kRWtV6shcECrFFa39iE3RK+xRhumjtY72oXOq67eN3p4rOi6qbHHBG
MW0La7WBNAvKR/+OAWkei+7M49/TPqG4UXybe01unsmDX3BI7n7zI0SScLyGCaz4xfzwokzXWQcD
lf2+algG/MB8+4N7+f3YtvV9mxHcNebEn4LQFg36Bm5n+P+5Cl5fffQCk5X2K8Eqkay5AAiwRTAT
7x+g8Vo5lnu9BgezSfRGdIIJb1mfZWVdlKpE0fr2pN8WQgrkr4Efc1bZvztl97HRlWLDzgtxVLM7
ce0SNBkqtcqWBDxVii5PX2vImWTboGy/8P82IbcU5B78hK81KkfdrDHo2baV64MyRyqFz8wB9GiH
Dat+xCLCWRgRoRq3kNJCY9MMkykVP1uX9hBpqPUbFo8KAqo+UsFSxn9mk0fIUpZQUaEI+cNhws0l
IvIwULnlailzDN89TJjxbE/4jpbzPHBoLaN1KI9WUPEaPJS6WgK56O8nCkkdL6Yz/klehnz5tB9v
MI06E2zwoUy6A7GZMc8MAMKGcH6yy309QRULYlwOqMarGB2YrgVob2PhxJZAsAcSArqV4GH529rN
FaIad0lg36D6+MipPOOrrBbFVdxAT3sRQsj63WTHc5NSF6Q6Ll3FvkQ+oD5+rgiSz7DbZu/sutir
E0C8t7beBWM3k6aOCphinqWTsQ0lwvLkROhGwBIta7myWVi1aiuzgWTYYmPiPy02IAWU2ytpv0We
3mD2J/vPPhhU0T7fgj7xGibWDZ92+QxqwZbhyounoGNhKAnmZanVV4kHobDMhWomdsv1TueY+1Oi
OcmhKuPmZXu9H7gxU9/o/rK42MwikUMpXCHus1qaE9K/iysOgDTvDeyaWG0qPWckPXfHVnYKUAT7
6dsMIqWQs9ZEzxknWZxcAms0X5jZvMkuLK97gUytc/UV//bCzsd7o9QjFIQ50KfESkSnimPPG3N/
F4rjJo8jgiHfC9lagElYCBzQqqDS/EyfRaANgZbzsbH+qBLUdN4bwJNcP0EFIa7mURzVAGCCQar3
eXB1Brlzm+midEXmKp65Hnipgaio2QMFsnHAHyz8Etk2lbVS5oO/N6yoXD9bF7MWy3dTO23A0HDG
xAW5goQI5UZDz8h48rrN0yQBU23kYgUnsm3RyZT86MLpIJbg45rPthvukTg7Y7/YWc2t5YHhs/j0
5xn9UwTOqUS30/OwFLCbTixGgaS3lMHmJhTOfNlklR3aIfq4KZny8T1nnVh+XkFxIetFLByDxe+v
kx4CT1SQQUjzSXu49a+aRuzdS+Dnvn/djtzgWkJpHb2rnzpcv/+x9bluQvPz1pajJH0C3G5YnuUW
ewm3nKXxoNX2+Z+fNBPzEXdKGGaKBiudQN5ROglGmQdpKbolRCEUfdctLSyk/fKcPtv3GmOODDKc
XrJiqMbAWsX2RmW7rJX4MWy7TXpB+ODaozhi8kZi1L9hebctu1zqUm65Z/qYyom/fAdyMaRfvUXZ
4LSDuc832E7RWFvvLlNTZeaDsYUXWYWHMEytwq7g3Opw/rvctaq5k3m7ifXEaNheRHWuH2wtjs42
4TnK5Jq/gSShjsewWNUuzIZHvR8vpYVnPQQTtzjXHdD0lv9p+3IWFED3fji1jJj47vjirMtYNGeZ
CTxSvifkZtLOl1GceSCUQh1cdc7HNETGcfe7lE403squwhXLI8fYHmIA7IY0jiFDnHg7Fdx5ryZb
Q0GzYh6qQm+rKQs/zKI5+VMBsugrbbAGoOwyfbCX5CZi/Y6L0KwXhfBqBWWYtcibESvuP8K5hsJV
bMJraea9szi1id7Jny3AK184vjTA/7tyzx53HTGesY7Ys+TjCg+rqMiwL+sYOhnYqYHyvRpaNsl4
A2g9+0x3jPIQl9FvTaJ3AyPcbJ63QwjYLY80SaCem5yCSSRl/R34OlYJ4FUl4RHwXSLUM+m+szqN
cIz6rw8FuUdKj8lPMI3SFjC9kxfFTFFsjdjM1VUaA6qr7gPQfl51V5W9F0uA5bJ+SkbYdod2Udj0
p5JIkaiXyq+WHwWnHQAJ6FJYqX+TQTq4Sqcam+HvTZk35bxn2uewCs8ZxJMCPYtzQMsa/gqxOFl6
Q64ZnDwVqIEOBANpv9CjCt4RdTBrloav2chrq2LJPYPg3EfCQrSRUjT3erKVsj8Mv0OydYaSZAJQ
3bt0vPuWx4gza7HPmv1IOqtUu0kaiJpxv/6qRYetzfuan7xDDnK25PwcnBHyZlpnjAWn7HwFbwcQ
h2n2c+gGo0IdE1xKvbvyV/aSWHQjN2GW/3MJ5rM5kPVTvj0ZIjPBniCIRktk9DJadS6OXrzkRQ+0
JpL0rOqkCGTCzeDdX/bg3ogbUPt7/jh6pwXvYsQJgJOdgVtD6I0TwDjZVZrOIeoUebg+7bll3JmU
UdXuWBJcnhqQchouRZSvxWBIF9dD7TKdGPEcTP01D5inR2Aa412kDzjNT8Mh9+Hq2LLhFvPcSpXj
2SpePM6mLpqEHQP08Teoru6rnUQYByUDRd035/2DOEOyi/aAGDbdZARB/kdIO1mPv8WkCgLA8V0T
Aiy+0p7d4IdflHR8uB2AcImJsIpsOSiMrOBHHIVhC73e+auz0aRX08p27moCEuaU3etxVgAJxAYY
eMtOrswqIZtmiEHWLpDRZe16w9EiqQx/NavpfeDtCGiT2sODjdgpkhomk3HKZKPfxkGYkpFxwO25
DwSoVQElXrZBE/XM1rBvCxH16R9N4jmw71B2VmVu0803FusAfOMZT/cByLvCqbZ63nozKS8Swb/l
rTCj8eDBXO/qqswRjXxJhi3/3mi88+WP98jBoiGvw1+x9psawepX4bB8wpc2B7+96ABhRsZUdx0n
Pz1ztv4tCkWfu1Xhla5TM9rJ2MytlMGVWBpW/1IEu1G0aYR89dTQjLnFn7kXcc/evyEAvzPprWw2
ekjnGLxtCU8tN3RpgNUoPTDwELMLuk6BbSqqF3+KmsgQ5xjrz5aYEih8v1HTFMXyZIIqnI29taNB
VNxdik836O0kE5JKA7erhZnWtEKrjzaJvdtgvpgu/gkSu2GvbhOzXGRrjibT3o0NJJpQiQ6PaqDg
9+UF1DVtPn/8Gr9jmOi8c0tWbCNaBbNg6dNwA5SFHm9E6sNZ8d8f2y2iPHyxFvTf2e6WJWjNEZ+y
s7yv+O5RynlCaq7Znwio7TRXXmn+U6TCqxte0w3/fOqlyQj8pf+RAivghJCN9p4QsZNhbpkoudr8
axcTYghUYjpFt086Pb+v98M76ZWmTyktnjohYxf0t3BvI8KMWSx96PYlk3ZzNyiwnxZmCsb7uEWs
5WJc7CI1YSYWFn4QL5qWlrZXgcmQ7rCfRHLwA6v7EA6TNnxaCEamVJyXRAX4ln3UMi5V7gKHL6ei
jL3UCCBSn8eERpoHBLqoCp4vCtIFZ+bI85tQwrlKZduniLeeF8vHs04DfM2aqiEDbNmIzr0slnxc
sAZZcYSlAKK8tHg1+8xrVr8f7ZXWvCa+ZVOJDTuxYp4lrbnGfcu6gVV/2RnzISbdq97urNUfePjM
dFqdcPLVvJGqCxUgXHVkB7hiJDzU/VM+HN8C0ArfcqUo3/2ZdndngYDNrphgaQMRRtYjcBgLqlaB
rWZiP7y8in8DSxNIgK801gHrameJ9tyP1GTnMWfaeybVWwRE29Aicqdns2SnJZVOuM/uq2/FziNI
8TF3udaCFJdG/uvi306Ci1CTFBuQFmwZtXOq1Ayzv3fS+WbZINN6nR52AcLHMGCuON2Lf7jS8ioC
07YCi3wNi0TEI2Ol/1mM7y78k97h7jd2MhpQPNALuZlvF/n9xh+sD8j2lT/QuTM4Gxh+RT9PKbx9
w7lW6tzKg3BFnt/xm+yNEEcR9N0q6q1jjvvcUSfpzAjus6LXFB7Xv4MmWyNx9aNZJ1IYjFY1rZF9
80UWGDezYSeNzfaADMTeGPrBmSQ26sQFKZxOvMd4nn2tO4vu5np8SoHQ91Kxp01UdVGnJa1ZCR4W
Dzcc0mGETJL17bwHjDpHNjDMP8yqYDEeyY7X8p8jX0jK6q9gtBYYB/Onf2B/1U2ptzp0mbY/jJc2
OttbbWMg4rGHIgMm25KoQvwDmUkwl9P3MdgP19UZ2x06n1l+70CpqoWbDxP/m9F7izZbH+J34lo6
Pz0TxSTku8fhkQYh9p7tvnKuCwxXqQNT/vbzgP9da386q2Mt41TvSh9IMRG2s7D50G9dmJP9xHXE
idKNGEc2z5onUMB2z1kLRNHroCxJyCyETAEVmT8Dc/bjj0uhZD1Tly8qovbsjUA5WNp8bpuMEtWC
6NbNTNwMi3M+90AEfjCBsMlPcWZzGzRqtl9PAOI2mI0igmGiRtfiV8LRA4ofhCw46m7u3GlYmyHb
7HfCC84PKcuKwYsm4PLJveP+SsJDVR2EYQ5BwwgZPKuEB4kx5V6axVbzTM38BI4FSz+WwHglpMCD
TNnV7DecBVjg6V4QZvLhNxmSoyLWIJzUOwN+g/bedIacvuZ9iXcxFQvTKuv5HFfF9OgysHQZRXqx
x7qidZYzLlKGVdEXltruCVCOaYK+iL1kngRV60vtzw/ZuAHoZVdSpMnURvnrORh8VxIRD+jcRnhQ
z/hh9WpAKzH2x2ojGaP6LKT2pFG3nygZeRbFOFORYrJNGejjXDmIxGSvU89VdxVh0vptJMWGcF4f
6LQ4jo+z2q/Ue9IZ0HL90pYVG+2OyUrYmVCfjeVd5jsa5teXMtniqVg86NUNVUmqeD729yxgGrUt
nGdn6rJdWPuz1QZpwyts1AjNvGbOXsJ4S0bdDaUMD23ETXh5gRsuxo+5ZR7qBOBWN65FnrlsrQe7
CT7tHiIr009atTjDXBHcmCNn169i6GCZflrvnje/KS+aqF166QaUWH9eYJhJfCwluuBr6GZ0dzpc
tYGlI7rlJCHeHKN+HyA9dRkF66ZYN8yWaJnKpBErtrVWsw8sawQeci2mhwvBvlPLlt7V39qH7Nk+
fMOqOGn9mzf1ifP1b7qYGWp7vAU1PbVg6Enk6xxLxkbJUsfE0PgT2yoCuXVoibjfuDlvWyKeByVp
WvR82upvHB0dClvCiM/UflDeE+pX2J2smUyphS9PHGN0uTbcYimrGPq82e+zIPWixKqbIW1ysr8F
uh+9pyoY+ofoEto+zjLBqdjZXJh7FdtzN5uMznyeNh67xRP4438v/bX/D0Jv4MCCACFU0x7zwQrZ
da681cYRuNE5k+H7BXv9Vq8iVL30Yvev/I39CxQSk8Xil4Qal6gu814meNKRbbMQR83ej3F972zn
C/Q2FgcQ42XAdg7SMga8e5rV7XLov/af3PN9X9QKHQYGoGrTx+JwQBYXzGIy8rgT8SMj+XL0cPiS
zlC+kuV5d14DQ/fdnEYQO/Au4Z45v10TYszag3qwWCOs9eXeUQipDUSmbewLB6tDCqpzqkkb658M
xFaPtzlYWnymHdE6Ois0OKhpEpNjUAWWTd8IDrc3pfMlLoPyv8a8Q0yO3bu9l+Kj+ra/aVgc2t65
oN2sqlYEMFvf02oLgHriiju+vFob0EhqxegAgNKsiJTuMZhKrd8AL2d8Dv4AGr/hXCIyr9wxT0JC
Orpe1oo0bgyh5lMQb9OPmuHbRzdE7n9rao+dYfMg0/gHdYlyvcoZxbd1VU6+2kSBXZJ1xNjhFEHh
sK/OnuZP2j8IyA5YqzOaC1CaU9gmd48QNWrCMZOw3j8o300AE5scRUpf1T/KBZv8J3FcFM0YWvcp
U9utsN+6/tyyUT6ilweCd72r88sxJPBmizBoTVZqE1N2K0Qc3k1TmO3O+x7BCFSQjxuagBmG6KN/
cWgkXSX8AONT41vbSytDWkB3wbu+LBWp5GCylrh7BjyUpxbkoVj6g/QD2IHvZ45KzNEWsrTnhQ5N
0a4Yc/RuibC9tei7UE2vGqq5JNDUYRp6maW9XXvuRO/ZvIX6QAzfdxiv1MbKMBHSvKMCkvGLflyE
BqGpsJEGxKnCcg/vNnlZVe3/1OOVcar8pKEfj9POY9CbXOeS/EndbnXybdfGykc7X3bBfrzlNbRp
bjQN8UDR8QZ83QJVM0nlLwjAAh+qCrRabDLFjmPg/TAFcmH4MqFfixBD0Tv6cZEQr7tzxyzNajaw
1/X/phiptl4e2e21ztRfHuwiD3l+8afq8riDeI0nRD/ZwQVrCITkUqwADxbYHF4xMPXK/l65x7D9
BgcLLmKNMcxCEQN+YffywfoNI3Jt6Zm4J5HGxE+B5gTUHlmXn0UYIy5gF3GY5iciridh0ABKLAro
XHpCZyiONWmARPdCU4JVbXDw9BvQFeb9kXbJ/gFDgzGfKn5IAb+KtFUvjR5w+a4p7pnFrGZvhXln
rQQU67Rz7x2DsULg96wkVvVLJTFi7zviETTbuunIDggVvsw6f7WiTOXCuCsAUw4DMkAcBp9hI+X9
xn98MUTNtpAD107MU9PB1YIy8g2eugwF/+iurkfASLoheiA7NAdu9MetS+/ltBq/p6HaEwd7yG1t
8LAtAHgrhvgQnH/4hL/dw0rKNoHIE3EO05f8/auB0kKkfjfQZ90yEZp5qGfmTnhVlxBZTdV8pgtN
dNwg59jrenidyuvV6XYUkfdActouqD0ysitUS6hswrBCdvgGdKT8XmjtvEm26qMuGN/d7szScBMr
bMnSXQ7PwU4h1PK0lmXnSsGDDveILar0E50w5UmIB0ZTxyrD/QrkEN3chrIkYWBD5xzvGP10/NQd
O3Zg51avyKGrzK/RY77FCr6mhpQIYzCDo3PD+IhsRb2Gpc3ug4QNX6o7Q5nsjETBZz+src0XlJ5Z
Fr+KjnblxWkf/VYWtOz/2Ow6Ma/MV9L8B0Z2S1bWwTAG9gCjKOVximFNz1EJOYdGo/PHdv8ysrX8
i89jvxShBWpQDA4xlbJUcuyQZLFQFho8QSteufBZdzJPD+SjFGKPnPd25YLMp4be2hi4ZDk0q11j
80Ub5avXDNCim5VqgBqei/4lJjW+rmzmbcQ2gmIOILS7YBbqJSW1bjEts8OZN3h8/lBjlvi+hC+D
38qFz/1mIRl8fKr09yuVFWpxsUWrI7ZQ9K/zZq6lVkIGa/cveTk4ug5tPNaQFEtWsgfd1Qzz4l89
868SpxrAwM1p1rq+evuoiIXBto96QFruzqEfZ8TYS1My34id1WvUSry2QGe+AI2WtZjC87uctYE7
7+lQyEgPBS8flC5HX4fmNzPtNwJcC5yi3ozr+nW3Nrdyt2ZLJ8/ZW7nNapg2uRJrwONqo2HJJFTs
yKf7fDxt8IQ1KeIXMvF2BaoVEFOk4sjxsvE8/7KZSY6IWbShGiMOH01HK+cA1wWp7HT0DVUqEuH0
pQOWofHJiQkgLkGbS0mpbG0hBJdOQ6vZpCq5/BTVJNZ5dyq87gW2hFOa2EknlOLoPXfWXBznZnEW
Es2OOEGiveRXcVzeNK/VCECN6Ku4+4f2U1g+OTCHccDOV8rFVSAjpu6T5X2whskzsx3Zl8uFO2Pm
XYyOh8y2KLFLqdXbzVV/HnvQ7fMhP5XD/KByQjQZxITP5vO3VpHe3JfsQZUQ/Wk5QtLyiwI0LcEi
w4QN4XdQoFUUaWMBSnTDjluOShv67ttIwu9Or7jZoqN18E0ocbro/RZyn24YBWWUHZgwhtMPzKHf
cbPEmNzcOO5ua43KmdqWDEF+YSsCJkO6ftdsS2YbpR/CjsuXPHJM0HUtFVkqrzjIA0zb2kcfXdwY
Ef6AzDFTvKLyJK2MeivA7Khs42oSyzKXVg1EROWVRNsjxTFhpPvuvh3dO93C4N3GTugeD16EIdKE
LXc4iMYsj0kuKfD2+Cv8qBYXdx/pKo69FF/dnT4yIiJ8eyfHV1BN75oQNkNmRA1ddWMw8Ayv4ykG
O8QYy2ioi5cWoineihxOBjpwy3waWOSSDFuPkGpNBqu/QQob7PSGE6GTEr3IBDwDMESp0e5f7Yju
KJBQ/n7TKgkjQQqdGVtIr5iT518E5RaV8wK1Ha8JeVMDKOjjhYRpZ32rsFLVoUm4IBvxF63FFiUG
uHds9MSfufjd2DCnOsTPwHOcQGCUjBKMhrV+HG7wsXIJp5wrZMEImYQzc5DILbYDp9v8OibEDZ8S
A1EnUKxVDPHGpFjNk8Z2tiOCA7CH2jPt+hXes+9vRS13+2wDpr4dNyuuunWnUgrTzHhztTZJFupE
y7BJnLO1N+Aw+MOV8bNmLvgc9iYKMuRSVjG5+F2/monOvMlBeOqABU6uTm3xAOgcRQW0oUFwcA3w
6YXPQl2ti7XN6ucbmpc8exGD4rl6v/Wp4QDJhnBGsfZDJh7FddaowqotjhFRzcIRMSNIMPogIFg7
6Z56haID5fYIE09LDvmbFBuNTGz+zHOwZAsiSHil8+zZPs7TWaKKc8Ovr1sjzLZlJcwMnSqg9GaH
KSRTfctdsH6Yx+N1HQVPHKFkRH8Cz1xMK8NjBUZJBYa2gnkMcH5Ud2xhyu3wYvL+tXjOtf6dD2f4
tIFh1O8Q0gfWhMoPRP12dBUDGGGZOY4GUCqrndXkY3hbysIYbFzVlWYVR1cyoDA4lzxtWwcMkIJb
RWRCZAVSDcGYyhyAGgB3OGIaFf60ICijZMrVZBkLyLFaIC21txwl3BLINWTPyfE8/owiRHvBLQId
eB0DekCtPBRTZmNfrGGrtUnvptG8F/kMaanTYzjaHY/ghUToyGfbCt5CW7A1LHrxNxmfCvTi7HuN
k/MmddoN3AOmxqBQ1dqR2VlrSUBKpd9CT4owSbx132htfY3X7090aI9bxVxkgY7cTK9HyRg2JhmZ
mInjAflTInW6bfE8PKwORWlyNbvo0e90LJ5Sa/uMozB6UrCLGcUJ9uJVrY0jkVeCnCqvPGChFQQr
KqLHlviXtlewqHGFvyrTfKPG8AqjexE8or/bSZhl+xbQn593jM/R3SvxlsYPUEIs0qkTQckt4me2
QVcJMK6H7Jpxwty51fZZsARw7ih8pYmQU9XThWZlXtw7saPIvEXf0ZLaKsIvWivFuVWCFZxE6/Bp
YjThGoLmI4pCfDXBz/3DmD0k6m3ATIjVBQETfysIDy/KwFCRH3fJzJ76ZaJsoTtF8YTSHSTcLbMC
lGPMkM5NEJd/hWSE6xTtNvSZfTTOwpvg/j4oiX+B+p47RkLiJdd85FjcU+Q8XJ1Owu3DVKT5TMeo
71rg6jmuGIaI6bllTH6X5MFURg2jEQ+LZv7d6kTLjsE0TdOYISTKAujgPWMLrMHL4q/u2RvTousY
/Ige7DHJwQnO84+ljrAMt/6jbA/e98eylCSVnWn5Sh31GmZHKnM59W/ZNI3hGhZcU5vpZ/Bpui4t
tgZUIw0QCjqTCr+l2LEgratq9Y3ZGNvWxyN/EIEypGrx2F0fPlOfS/jlbHCmeM8pOH0uTciURHRD
ZwL+n0HC6n6+ULw2rgJsYTwgaghImDuPZcbtkMrHecSAWQ3W/1haRjlWJ52/JdSAJ6PATG+UXx7d
OuteMAyv8dC1IXUz4wQZe61brwg3mrt3Ks93lDLm/2I2I65EMtUPUfWDVrO3Yc85RXWwl4dTwx4x
3J4jN4V9fi2REEV/Li1P8IWl0wcunSvQP3b2oA92fn0Uv2trbxUwG7c1SqYLScAdUAl3kROwvqSO
dGax8XU6O4TEaB6VGY4tDj1ZtAth2RbVAPhZ/Uvm1jhnf2ZrxDvSsGlG/WV8x9ay5YjEK1WaIiJI
1l45ZU5JGd8CxqhE6etrW37Xxxj9QHgTQozarUc2+sKoKwxslEQCzxydPX6DSbtHTnFB8EmP0sSU
XUPQxtDT7iRw7jLpJ0V/dAbOiQ8BkPe4tSb5OETrn6WEFIWVIKLcrmERd80aNy1HalR1qGrNOKGX
zQUEHafOhn3gGchldoYOPIb3P1j7CNtbP65P9kTDuG+Jot1DrTdrW9wG2VX0VJ17qnPB76S/Yo5r
McGYbW7HZeBv0ZOeJZ3PWJW0oSNwTSI2tJ9NawhnTgmQiSUaYKm2lYqqPdM508rNvznhX1+RBUUc
6aQhhAcdJNWlNzPzdo8XusTGp+1xnD6Wre2qUu6FbEDHT64kjIze5KgLsXjy9l3LvESUuNl09T0/
+933boEptflpwO13UuzC9GzkPm75hqmVYkjpYZ1oY+/VcO5U1ALWnqIw+RRJyRgu7VOu3lp5Fujw
iRzTstrcmOh4NJJyOLgekb3srZp9aX2j9Fi2uqBT60RA/mofypDvwaKUyxGfid6ZBvFXZu8ALNtV
ikDCcHvzrLMKXXugoraYQtLINQr1tDxKZpJuZpEoL8zRXexp+tShsYwQ/9WxdPKxwCySumUgF4KG
iRtIieyNE/Dg2dM6WsE4Raaap27Ou6RWuTCHJfzbSzcF/iA5kTFTGhB+O7aJr39pWDPIf8NGeMPp
PH3w1Hij0gEZRJdVOtB/RN/uuKBdRjcDOYpQr9cuprvzU3De1lgJtplzuJoeUzNlyWAjvfy/QCja
eIWCTMOSS0LmAbQSQC+PbS2Xoaj+cAqdiNjI3z8MNt+6HDuLGaVwGY6OAQz/VH4AR7t/yCILeOPo
FTFmZ+GC+31FNnb7s1C82uzsHrIWVSrxQufDqJ2cJGBADFDIr8n7hJfsAaZ0mbHyIHXft/ima1HK
31X2QVeAuUKuuGrCIxONBXMlHM4FilIs/2X/9e4OtO1ZtJUyJPIQctZr3Dz26tXFmHBgdOfFuGBV
V4QK9BaLjpeQ/aVTe7/krC54iKGdSRQcc+GFABzh5sKxHtyN7Kp7ndpdOrBXZmmpNHASrMQT5Nea
L3B1VPjdNGWh0d5AXoG+aZh/MRB2v/Dvp5Lj7lNUbLqeZ3x7upaI88u7p/aRVkz0wgyE8cjJwxNJ
hPU1iAxS9d11mYzoFlRTIHhj3wbYyNW85Y1alLpzRxqm3tz7GnxrwWLwwATJBjmNjQwnRP5Bt5m2
BDl4ymYYqVaZ1AfFkdegrFohK7SM2cOb4Owy4wREI28r25yCr6egPbpOmwsOn1I5EmyHzWivc6rR
Y0ik/Gu4hPdwUK3h0VbzJinUNAm8Jr5gfsecyQKSYXxAZpfUpWMZzT9sgQw/2VLjRseLEedPKJFm
VHkr6PRlAFAvnizlENYSgsRPfEO9LRFo/FrfwV4V5513BY+4W1kLH3uCn2iHxnPKJJTFZoBOQifS
YHg4GZW6Wv5z1ldKrwydguD8byQNYQ3jkqSDxyEbzUDaFF66+aiXJrBAwv35rg7HhBnIhBrk/wPW
onNr1/8jftwK7gofwivgcVkTUPuAFQnzOTRSLbgNe/WFkcgdj+Q328pKXcvrm2zUvfB4WolnL4dO
N8iMosoSd6MvuIEMp9ae5frI8vBIi8fGp7DfQCVMCMtR2e40uQZTLhGa29wR/JBTKfXJ4fPsbVVZ
FbUq3nWZzvHVqsJKGJTWVXToj+i+0v69gfQXtagccwBhSLxvs1rmpSnFCr2/lP2Pvt7LESXWW8e3
hE7zPWg8pZYh60OmLkqLyufzNMgz2TKC1B/2MWERJqOmv/xMAmixzyf/Gg6yxNT25FwkwcdDb40c
5KBL392EqpXy/hoijrJtDZ0h5Yxn/LSW9sw9FaSjWmg3/EElZmNOKlkeeHQ9TF8ne4i/pnqwFYeV
cFKDs5NKNN6/uUn/0Z4S1eFIbgUKImQjehCe0dk/goTdnpdVMhcmsO7dLRe6CjN0SNt/EbGuZvQJ
Pg+o+fj2Mrvp65J9eLuzYHTAITCaIw9peoy4CwdDwjTwNZaplKBnDqV9RhMuUa5rUQHy6iV5hmEU
ldxcXxK0yLPMbGhFwIeyftyjHaqC+IhgsQ4oBO8Xga8vuUCKGJJa2dWZr9lxRVdX8N1QH0SLbmJX
m0eHyhPn943MhS4O9L9UuYUK16Inl64MT0Ad/J8FP24Be2C+s7aWnkyYOsLmoU5sAv4b4k0GhkJJ
rOV/dbgkcvv5AjrbZ/FL0RegAbDtijAatq52pfGIh5HUJYs2/KREOwkyb6WYK774Nc4Da2lM/vPp
9g7QoCil+6T8QtskaT7SV5hnB+Ma8HPPY8YXISez0bfVjxtJOm1ifGfegAVA2oOv09iBhVa4Og1a
QwqJo6rNVwRUdYTr6ZDcvxsQK6C369u5pGt8nFIPOnIDXx/kqp6DL/GRMGi9e/Xt4BeUChqcWbMU
WmuGlX0F1xLaJQdZcQrsKm3c/Zi0Kv4gfG3tF2EoWdM3cmcnriwKNijSSlcYAjK2pMHvVQSUV6Lj
tU/dj7aZqyZOy1hBQoH6RokcK3ZvP2Finl6eK/IJ6mo5xfPB72dmNyK+B0DXCMqV84L27wpTQK5n
nOOhlFOeeSWV00Nfxt+IMYjFbkKfnaJZRIWAOFoGFKqIpROaujkK2oI5NbBGNrnMjoExTdO0W1UR
CbTXSKm6yhnuCsaGsEA3k8eem6XONcD9FtpqqZ9kl/7pgYOCZmRZ1uOa9Wf+M3ZCoq531WPBf9/T
mAmRawVsHQ04n6Rt3Depyg5AS9BrvKtvrPcyK+QeRQYo4YTh5kCkVSxyRxbD4ChFIyoOEr+2ZXz7
cOc6y+wLrm7e/mR3YGzcOJht9/hTSsQSsPfAMm4XH5TuqGo5sEu0ZQ50lm4/PiYJDtaLdqM9mF/f
sOpUgPQYCx5/2TUox205mojKwGmKmWueW1USNYqyOblk9632mlU7HGyltzWI7YgFvZ2WJbeM0GOL
nMKGH+G4YLCZydiaAOxHoBmSYBh/fd+Vpn02mdKE9enpP2bqlEKjM4zGkp3hpYWslVLBf21isaYB
MqFkJNG+yYeB3OtjIt5f5Lllu4Ohtl9T3LJ5Bwjw4oysOHHhJ9MiM2Jjs8J31DviYt8YAN8LMSCP
vdw052bjMZyPLkq+f/ZjF2OG9jLjsh4XxA2EHFP2l7T+xILolJZN0xIRQYfUAzrNV2jnOMCkD2qu
dLq2uuGf9UCfKynKj5aCDgACpH1cT4zeFbFvI9VGmubxMRKXpr9fWXrVhmYSYuVeDhC/9S/wh4Lt
Q90YG5Zce5XhJG7LuTxJFNggmoRMXeZUFiTi1Xy3Cr6IHCrM8AD2cto7pKiTuxY6nGWgg63eq7GA
n8akB0w5S6iT4cm/+0gXEz8VXrxKHtKHUEBxAh2gT9gOf3RSP9N2Mft+ID8/RUq17fSbBHwOpWbb
/Y34MxBzEUp+SUBOOPuu/Dmi0K+8CJ7QVyN82NNl7uwVu76aRZRsZLs5pJKwTA4fVMpgIn5VtOAp
tL64ZtD0cj1d/eiNmbdfv2UsXTLNm9anb9TjqngNvo7wVgwnL5STxK8aGSmtjpujy0F+99p/a9U6
o8CuDiSwhnlwTe7WqeaLfPifKRSvhNKJm26YIRlIf8Zf7YZGSXtbckbXCU8/P6zdl4jrHZ83+wzS
w/PGmjp7c82jIjiRjtfX7Sk4ekvoz6Uz/gN+HGs8o1E0mQjXbTeJNNOYTSXvdXTZf1D0T6bXKgVs
cWXTBbVTOwvQhcdcwDp2/jEiifL0F2P/KUGGvu4oo3+8EWJdZ+jK1giC2HijOizwKXqQ37lCklRT
zRTZcUiaZl5EHku5Dz3BCxI6UqWxvKzo+rE6M967OwZ0FKP7JP0QhqjwXhB9Cfq0qaRS3q/y6nH1
g6AEFSkzWfpooEbh1en21fUAZhOHEFnfOCYU59U12sniEV1OLqP0TbVfmPzAnZta4GtmpFqrTEDQ
Llu/yMZ/mOqsel+uZ/QD85pBY3t6CCyQnKTvexhTiG184ijESduegzoROiWCrcJ+VtHUuhEyk4gu
OO24KNEV+d/Xf3bxIkJcKUhDSJg9VoMaKFDeYF7B6PuHBAYyie/ByyRRkJvXrOXAuVEVeu2lA0Il
C/1A6g93+wGmwLu6B6pipWbTb5hKc17evKm2PeonyK2iFyq98ss6+EElKPUYMRB4Ov/zt2fNT3Or
VPbf4x8VYNRfN4xoGTOvH1tTfzzmnslEZawX3h8PeZ2XCuE4jnJdhZ/NT2CeT7vAelz5c2Xgwie9
3LfrKS3JVvOFyaSzONV6DrANLdtqjb4BqrljwgU/svKgUg1ol+cKuGjVpa9nN8Ts9VpPNFKEVoza
Q7p8f9v9g8QMKMGR29QxOvjug4z534uOMYw2tsPaqY5W3SZrvgid+ridWq+EUN70yz5Nrci4c11C
f4BIW2x90e7zsgIp2rzHYqHHuuASbN2Uxve2lX6Skr1JfORUfHHjmdP0eOmYLZEiArBnCFltn6WH
I+NTneQTB9t4QHfK8+VHumvJM4xeehDT/yU1vVMGQ5P31guzlpBmEM98m81qlZSPeh91VaW6WeqK
RpGsKmbRmXnzrIsw6sie29x3DpUtD9SF46/RWZmHzqZy2UPfRFJqg/BzQMeJyUxGWNt2yWajSo5a
knc/rJXHTf1LRfwENZ9nxsVlncyrmcAQoWjR8pIkMQDdBaIVyuYgVozGbbMDtTCNunMv2HYtIBAI
KTvuCTTzqRz0k3yCAOM7dAT70NTmX0nixtO5BoCXwl5I1Za5knTO+Xw9oqSnt5N80P3WaesPXU8f
663BkAdpugLAx7XN+Zk0JOd4OKDXr1hbThGJfKc4FxC1P6Xle9LrKrJ0D+no1B36kARCy6DlfBhw
wY/k+gSRumiODymkxcz53OZBkdRzwPgwDjduQnCMsGnkMx5aUIHzFc+yS2X+qiNTI9PUpkC2pZoD
keTcEHkECUMvPsmkxGWaA+fLYWXb/5/IDtcpVlanIR4BlbdZcxQBxyyuUUwBtT2aRDvsO2K/xMv3
X8uMlhHIE11ycrMUWyPMS5D0FxkRy/hcdVzthccx6YACWyrRFrmQ0cn2bb6HfGLe0y5m6iabhUOu
mgmsoCm0w7qQbVxzucg6dQOGoLAyP8SY6BtYLavWZXXB2h8T9VtASFofWGtnieYnrU7aC5zXwkXl
134et9+O/iIBUTxZ0h93r/HihltmA5xEQnbsais+nL385+wX20r2k6z8GX04VN62cUwsWppGIAfz
33TQ3M4MiC85r11SY+pJa7NXq3179z1ibtvRCzyuWc82iEU/bB9sNQtfg4OFRcdO5tII9B0Me2i9
uCJkuYVqR4dlewmzTqWrR49XC/Xkshaw+GBKdHQy4zBjJFAi/hYd0KZebr9fjfZ/4oNA8gU1sFJ6
O35ZexSQUpRC1x0Drv02PEh07BkjUZUyPawp64q1zCgaLNcrBddIpFwTzjDhiWknkyfJhSZhqerd
+mGUh1BYdvCk4rMKyF0mjwSTsjZM/cvQgNrtcrp+MldrauEntx/YmBrBuolI8N4ikDFAWC9SryKJ
yQp8Qaf2AulI2aHKo29sVRGRTWTQrwBPkT1t6PoLdFElxDHTOWrF6QSLCfxptMPDwtVnmxNgoyCF
YNF2jxHaXS1AZmbLjKXizRJDgiT195oid+aevFLaRu4fJYkVu84gOGy/RiDWNBIJ2s81P9tZ5wFJ
zz5WyixkISBvd9Cd1GvIJGdRnfU/ujlGr6wCwMFsxwddpy54jCv9+qRG2qgCQHYgZDmWasu9XFYp
Bj+LFndR/kgt+qJSn+ByeZRStmNE3H0bkWB+bt2VVbbbAtimczfZ25Q6QkZALk1YVKodfWp8OaG4
Oc1KXRe9XYHqXrc0X64B/jgM4nYm/0BBISsbGK9v7spGefWRsXL3yg012J1SlWPFxa7OiBGdKTCe
bLKaGscBgxmO2HUDUvVbdynMkP3ZNNq2P2PbCbrpIjPa9UIDK3uyBf7ESZ0Iknv8cI9dq9LcVyqf
IMdHz/7RgJFgcBfRjr4WrufAgZNvl/3FZZ6k2q5ZyFDvIr6+WafeGPq/w4zSyfj3lXL5vkbdsN52
q/Am/rvCuzM6rHgyFgIKirJVXboxbfCR7WYXJ0oqt6ZR2zDtI9jNLuRNR2ZmHiL4CTLaSL9/DeAk
sKoAM0tpnpRAhmgKS0C5cVuZjOwLicfPTnTgiKZmiE7QRa3h260a4oZViyvkXYi8rlhxnDYWxemG
v7DmRoyu7TdYWCQTGwx3VM54BWyt7jlzK5tjw8PLjySialgMv31RqFt3vNYPoE/E6Y9lIWJWFfUY
3nvYGpZPLgKxXyZoDiAhAc3VaEeYbYCYn68M84NJe88aWX2yUxBUk0NxDM9x6+SBU6oNs/5qLBNk
/M85ikeGxwFb5x3qoNliJMQ1w6elKX58sqUw6F0RtDD+6VTY9fNuZ+Oa9noC+HFWcOqBWuRGp3iC
ppZHJ3IeV6f0I5kIYS2qP6xVijfXKSIi1CS2Pd4sTvlzED2gRAzFyqwJm7EUtxXoJsS4CZU7sNj2
L7IedV+SRZGDGR01LhvrmX1K1ZLiMRDm74OTF5pL5HbmNhNgFr8JdhydP/KtdQA90/yp2ZhtLyEE
W02HG62auYgXEwUtZRscLLz1MPn3QagEecdKm6+xEJoPEoBrHjvIQw7t4OH/P9Gxix08yncvRlGU
QooElcnQiVGRJLv3YD/GyyKBu5H4fJMNyqJ9ga/N15N6AV0siq7DE1Dqn7PveNErg6Q/KhuGcQWt
xkgELTK5NoE2yB6YrYz5a62PAtPP8GW9NkjuyVvCaFK1ikqLuCjqs26j7FfcOtdz/8bWLRD1IP8C
0PT42koHM2K5lnBtbd31J+oKqco7VRZNXxlGXTDPjjYmAlAuSR9M/fJkq7hwOD9KMTIMENvJj/hg
C4ChuaoRpkrrj9APtrB0Ha0a8SctOcj6WbH+AI42pPclsnj2zpU7FvCdqrxvI0N+ZIGJtRRwqehg
xJL6Wk9F/ODI6P6EliQuVjj6iv57C8C/ZKSl24mLEyoS/5Wepm3sM66YLD82IQ3/Ya8B0YQzjngn
grUV+RT8gSCkBGru/ChuPNEug7qPXjWPz0qnhplN3fDf0YntgReHnCuydUPHihWEJcLcmZi+vFbN
RiYjhBUhWok+vpu/MWqElVHC8yXCXw+8noAO5etZ5lOwTKonwM1voqRMQW9l53p5yRSIM8g37npN
SoMEMcZ4RmX53/xh3qA/HirYuo+NE0zVdNdiEIOK/eZLhBLMus/ftjY3l1Ny5J1pGMRUOJGJuMKa
KqEa3/zn41XLkAFY5wM2xLvT0EZJo0jwovuTVxaINebz9uRpW1dM2l95cXoulwP52/8oUXrH5SVu
Rk+h9eEFoI36rujUsHt0BtPMRo1mMYc3cPjPFlL5qhEan9LG7HuRVaCdTsBNeGXYJ/wFA+UYvisi
8hVWHEGUBOXkYlo3Hchd96fLfXoLt/wTU+LfbsTuUQd7EyNSDrrPVKpsW8EbMaTzH60Iam+NM3jv
zGoZVO7qcHmATXEjXclxqaXHnyRmo/iruIxaJgL94ZgLo8YMhYIlIJcvBodsLW/wGV7NAzqu0irG
YZBycBo8HZdqeQmbm0IuykaQtcciKxrTg9y5QlkWekDZg16kTZZodKLDOEeNPpadl2Qc5WjBoU8Q
IIvL2jzJCe5wvyg9udFIAdHbGrl8l9MPAMX4RZhW/djzWXcehn8UJXxX2n8kimxtJfOffxOszDFO
sIoZ4djduzxn+AncMu0/B8yVJthWS8jwYzWIgZN5o1q32n72sjcbl3/60TO2orIJgDJ5hEctvDJC
3SNUvTDxqP7Z4Z5k3W71ObcAWltmxFUF3NILTGqc1OlMsaVRNxXwzlqF9BPuNmwAHfPCznMcLg9H
K2G7xu+x75DeTEVh+HDS7iEfrz0WpZEWbZ3tRHnAW5tr7ixrBZm8kWvAiJLjOW299Q5KoAiBICvx
zVGARfha77QYijfp7vyYXZDJ6TRJWyJfcmDe4ax0SIemqpzNNVcKgTLayMdlut7OdvL75LJFzJ0I
FPfu7sJY8gIkOKX2Ae/Ga4hudqpzwJK4NqOXcgRgu4/S4nGJ/GNThM58RGL/0UgxCYNpE0HdSPnL
NUnb0+6TbazV+6J2ppe7+O5WUai7s/AomjYUjbUON429AWjuHRZsAcLJmdcy0Q86BrOyHa8nzAkV
VqNtga0+p1s6CryBmJNMnxt5P6ZsX03NbAydGUyie6+NE99Ufouo1O6ka5ApFgBvqOqcNdcMHKjj
lGmtRc15DZedmQ8lcMUCBbS8whFLgVdXHapeJ96yZUV1yfEQ9mesNiwi+UDeNu18t/yQ0QTkFIpz
hw73xX123t65tV2NeMYMnPk/di+JMZO4GEVs00FlRptMQY4GK3TQ95XZX0EEf5GblJjgnL+edqA8
LCE6tVMrK+pBgeTQjc7mmxhRPMoXGPOJmCJ0VajbDrid8vVDTAXqdK3GWKWxoewRnD82WtsIWgyS
IkfEIBDN4LcTiYKL/Ia3T3ou78RpgSgm7yDATtFBMKFtlGFqImJRzXPlAY+PKoOxoBuaOz9eqMVy
fxqlSRVrBCGYqwfAuXj/Vkr0cUhokCnCjnBsVX6p7mogY86qpTIgCJt88ZAGok/fMcJ80S6W6A9T
8/cgn5Bhm+gIiJ+L/P7IRwHp10UySPOd/L1x6Cn/lKahn8G/3V+jwAsYUNkyxhiddrCMEsHsb5oV
U4o1IZB68TQlHYitt1CTSMpzxmMdYS93AgCC5kSP8Szb32NYI/mXFLYXVYannHj1JI0CtjkaOhld
nlZSVM6dGErZuRK6aexPbc8I9y7vllZ1C7QbBAsaIRUV/e6kQRbtWY+ICFYIthYS+zWgA0WpdGr9
UwWbbihf4pfh9j3nT4FdnxEKdKZQzs8QorJeke5TYDJ+a1FjdgcfghQXmhJ1h3G9vPopOqj8sSQ9
bTTI8Sm/VzRs/l4K2k/MlLWVYWTYW0op441/xf48dT/OFQY4Du1Czi8bqcafiRcD1MTxthudUKEi
jpUTZKTMPgtOjwQ9cPA304ftB172pvfp6NE/cxPnk21HjKb4EIeQH5gSzypPEDAGokHzOZ64E1Bt
Ku8U2SIe24Z535maf1SP6mdk47JPuS/fCyYUW0/polwvMcNRjWfmfXF0MI5mpnGgzChV68Ju+uMc
kZcTzoy7M0JF5qmKUHtq5rGuh0pKw5pAuwQ2+ibdDiPYADUWKi2NL5yubm2h+FJoZK9/4wnjTuDq
ygcyyWkw6dhX+l4zYWXbIDfj2DgykGRRS4NiJe04/0NpmVJTjKAexABTAkQmXMUwGWJ66wZZvdZV
l3mBRw4bCOuL9eqikv63Dcq7x5pxyWC1YDiJe5lqIplBPl+3oadHljzC2gFoOn82WKYWxcOFCabc
omHxZXTc61KMXAETI18U1dUmWGNL7ZUN+x1Ps6QGS3I6ohxTE3d1nYetw/TMECnTKRWGFhjDKMxi
svDcsB4hWscN8EOWBnIJOEWZrt5ZdjoveqjVg14tvAsYMcM2rm8gP5s2RAd0vPvDDj+ZK1lHC/4O
Nbm+1Ajys5Et+q7vqQzjhsqiKet2p/TRvU91btzgHgZswHqfmUDvYpegQTmdUErRO7Ii81qEblAB
vO3Ds2hizvw8TZqKVbnS0/1jQfaSXBUPebbNTj/t+oLlhf+z/f57MBR0Z6MeqcKKvK960O/wNXSE
CYkQ5ByKex5ztmRCuxkXSAWvNH8DL8Gk/5IvBR5w7YvuypTsFkzwTbeV1qJ4O13WhB9FFMo/PsZM
zWAUhz8lSfWs31U1tQcJ3Do0QinK7VtZBmDk/vBQolW+AIqaQJ/wg1RFTIUGI1gvymK94Pd9iGrF
bOOoLxt0eNCSdlOWOUd8c1NBHEsF+lWywruzFTx2/sHwKvNWaVu9B1eWBpwT67M3yH8b23lVJeVA
ZdBgC2f2OgKcSkqyGtSXN1hJKKfhLOREdYZjcdeHDAxR+zyNu4zS1RU0vxbTE5N65pvmaA63ivlP
nekf4onkF3Ebg0nuqOCGHlZnSRqk45EMm/dafKJpfRf+/LenFn10XyrcgTbDY0KZHext15FaWbhU
E8PYjRWjedM1xn97U8YMqEey4/Wor+B31y2ehJazC5vEQi4BP+Wh4+7r5XeJc2H34iNPqRAlTOaS
+pWYftFZoNWQ3wSt4h7CELzw7kSKiwPUTk1vErDSXn8vB74UAvFtYSUodO5Zagy7luzWwPAubEhZ
wSqBP0CoNgb1NhV/+JvB6dYBmLVnDzkASioPKpiMAY/jl7JrL8UgGTfoVMa5o5kW3in7TAhjkVVn
seQtFQstgU/hPbz1N3k3Th6LJ5UE49cJgzldFsxT9LVGzlvE4mxyzkEgVNFvBGi5QJ3eCcobQD7T
jSgW90qsirckAxfzI1X54OyX5tDlwN2jZ8SHwY82S5uyW8nQxxIFsBfHF7IOV91ywGAB/XfgjDbQ
uKRgXOkWb1s+0sSIvc7BXZ/Yp4AkrQzTeGQNtYF6xxsaaf4gCP0ErlJbQ4msE85g6ARuLJFJyfHS
GwwGyfasJckBOTvC6+te0TKyKMwB+l8qkdYoqK6yTKFQ5eYf/ZsMxHB3AuEBcYkkz/CvJ2c6hXqu
frPQKQLDwmNEjlRn2oosnkobx9AHeIVXfAAIGxptwzmxLmh0ATbr4fDrELE3qQw1onjii3XrAh59
xpkQEPNrbb/IC7VjHQPxF0SO30wu5EGKDGmGlLbn7KIG6FRhcEk/FfSMfHMSuApnkTllBTJ9PxdY
c2Mw+Q3UpkVngb5RTYJ4RBFKdsYG7dFsFBmZrasjv3e4h/GZwkZNS/xWtyN7hgmt9FykRZdKwSAh
tHGaOiuObHBlvSASOxnjPype6arjipZHtaRdgcc/R52n5TFSD/YroJqs7Pp1fHakhu0FD+4vSXT3
9jkttPECVIrDeQkuQaDDgPL1stcKfUK2+ulyo4dmi/RpSVgthMumf7T3YF2zBsPG44ox+qRVa1Af
LPOrEjaorp4zChzwWARAxpM8iORCZiS7RCalry/vM3EQrILc2Gak6AAc9X0sSbbfk4wOtRIeD16s
dKnq+q9Z3P/wfOmPJN7WmpQzpXGZFRCDVI+G/QkmCITaT4IQJBARZUXIg6enN6rzi3OpSAyMIr1X
9BeAsA+axx+UEH1+4T1lxWqBsYFfVRbvDL7bgBH+LHzwpe1IKTk1j0m3F1J2SzfzQ92II+j5gV+V
TzgKrY1wXrpGCdx6YbWOn8eoahj0e1iIJoeZwT+kd+a6peipMuF//zLW1oXe0bbmJpFmXuSe7aXE
eMxmLXk0bRtpoTxi2YYZZ0Ab3yPTyvIy9oE4ripsyz+CKrPRigyvTu8qXEX1LEvOGiDhaHT3TLp5
wc1ZkOnYwtvATRzIRK6G4Uu7rN1rFwGh7miyeSvuBultNY9jfOwrZC9sTGbc7PeyxahSS+joJV86
T5Eht4DAaTGnO/AaNjYDs+nFJXqnSM+RIpQa4MBYnuD2RjwDojxF3GVK86rVDRMj4O9NC58xzm3x
qyTwFvUIjvO/tnZaoeOKMNrKOrFqeFhhOXm0UPlver6qSWfKcGyzzgdS+4dymMFbqCYqOImFSKLC
h3GJs/s8V+hFCpTTEkmRU+AWl4aMBr+0RRz1QZLUXfZPznp+Stqx8ShsE1gQ/ftcOs48DQTzd79s
sBRDOH4Ld6yZSw351Y1WaLFoDMtW65miSFFUqrnFBPOvkJC0BnCQGExOlpEte+0nOIViiUKaXxzK
x3GrCl1y0rXRAj5AOnBRNiQaCTO7LSyvzsUUzQO/wdS2kOMMk8iTnKxc8w+j9AFEydYZOra7AAu0
dhmfQJALzQZqw+z4KOFez+OLgwZhPfBmchQpIDp+FvPB5FdQGNL2CM+P8SkSTgW99jZrs0KDYzOt
NmVrxkQf9KXf0HCf6oB+ReNnjMd8pvhWlr7xn4e0/poGKk0pU9zN4V/ZNvQsiDMaVe+uHpdsXssJ
0wTakwvWGZs/2F5CDfLVbamLzBVC6nvcI4a2t0bdUoYwAanmAT71ZAx/SPaUM8hPyx040tlJAu7E
0teIYzPq2KgFQNUnA5qro7Wxlr0PncWhh9s/N8mpZLjh9hY1OY7+LTv3U3DqkKiODFd3DwCAMjgk
D8wgcPI8gP2MvgKgP4M1rPtPsdbfuguizr0X8jtsGcflTpjVzl71LL/G3/0cY+RersR0Pt2kpe23
AN189jFeFRfKkCZEkFlFe7l0AUwyYVZOX9mQjlsXUzHkimXZVjLzedl6NNSk7mYNIAy1GqsMfuS/
2biq2HLbFu7AQEojNKfL+wFmk9R3ml61HArRX+Ujg+W7TTLDG1Tl7oCuKJg3HGjDQSEo6/eihlj2
F4E6jKl2vnChu1ZzeYzEuKH+dvwUgy9JTMRt6xwFe4qdf5pMvQKVf+DNF8nOr/2RAftsrzajuCKV
986RjA8qHxzKSour464zffTtUKMJr8tnGdqykmtVLinBbBcqo1W6PTEtD6eJUSDh6UJYxl/NkvkC
FZ8ka8/yEBnIQFCZuys8NEXSQ2WUi1T9RH0r9ZiiWDZDNdnV4mJePSrQS7JtXP/WJ8/A5hctfEbE
x4eI4vHO0vG+j8ph8VoO2o/Jfys2+1pI0g7OZj9IhrU3xLTG9mtpiOBjtIVst/yMqnndVpzIPPLL
XJg1oovbafx5MZltLf9oxw/OuM9iBQnnH/JGxrhYD5BH86TcWB4+7Uzss+hFbBNzrXIBXTVWRJSa
o35SgsSJWg3sY3FZyZFtricRduB3PbvNSEcO67VUz/a1+XiauM0JUkxb6p4y9ft4gtFyyWlA/Fgv
hmJBrLHoBpaWSMS3RE9kjlCU5fwQlkOzE5al6EhtBtZDrmzixxjSk51UJmPTvojZMLb8x3xb/Yt1
gaSahTHsoLOKWYNGbPwEQowCwD4tGrjn7FPGTu2WZgjjVBE74vW5UxZCfBUnZ++R4jGAnsE6yrIj
RjVsCo3LDuh/wfkzqE6JMu+PYcPJQNyH/heQqaJauK0OHz3eeIRs/hF/Jq7fYLNB391Pt9eBn7mj
OJZpQYyRcUVU1Q8X9qG+5z+xEH5Hh0q3EZGoeiv3ddds6eEWmHuDfEntgK61hfiElXykCmyI1zpe
mb2IoaAG235zytCyz7unQN/GlTey7bVjS7Rss3+jxHb8m9/rprzwiz+jToFiSN4WGkwT2feamVOW
qSjCbO78NnBeUjuQ5dCyS1SQIi55rjEBf/U+IGLdz2fKsg9A2GhTityuhRw+1KUSHqmt4wmTBL98
hLoSygYw+vlqzEuIHtcYnD8DmFKmY9ZenUm9UV6uCe8SHgCRmKAzWV1w/f3bQbHGo41xd6wRwLGB
U2T36iqOUbsVkj84niYxdNksHIXHtTnZEKU3yqGlIdQ6YovGdPXe7P04yM0AIdSc0KWfq38mcykx
2I+SztZIXJDQVYFOtY47adqpZYPLe2DLqES+E7zWSzn5xjbwraM6bcWWh9g0KsTQs6KTABAnxIs3
TcNbI3DODbJ3Kvy803RH9P0GDEVSuZl9fnQO6UY245trIYTWsZLAE56Psmdo8ZlOe5OPYIpEy0uz
aCJDIxrXsCmH2JQoIijQsgttRGGA48rFcJbcqooRjvo1AxrGjEdasp+v0MDexNcxpxSPySer/uuc
uCUMkSM2GWRob6G0sddUtlIaXzWb47jQ3s2i1jN8c2OebZWe8M7kIq/0GGCUPZHM8XhWVKehJ/u2
S2l3B3ul3yp9x/8vK9u3GfcIDpwmUZFKMZJv6tHYH/Payn9sLkB61D+4rHYx6xLAPRgMQ5n3/1WD
DNVjVnNhlK3iaLnSmFt74LuzVJ0dRGUIOIKo0vtUqhYeE1ZZm6VryEsWtW9VbF3hPPHvdWC6X+Dp
he4hnCyDI6ggMKnqIErjEYhCV/reJd+TJLJJuM/lQxTajsE5NZQX95PzRd80GIpWxz8nR72sWHcr
kkQ1PTQIA4BdH3y5rgl4z2RiaFkv8ve4nbnbgoPLNRk8ujE9igGi0hHNAXOCO4MWkndAhhW9zjzM
7ieEULdgoiB6QarYae1slia26yN3XPLFgg07QPyVeG7Y/+6bf8uqIQTOmgI2bcFKnUUSneLnxpZ0
klBE+RlECHsBXsUiw3f0nR1oJpXhXZrZcxHJ+nRRoztiOXXEk32Ua14LFO+zHaoWaNoqS8VW8LsK
iz5QbhlbnQ24JZv8azBlXNnRqoR7LhpPedeKaNuNCguYJN8k1bH2jUZfk/rLl+RHyYtr5ItAtm0t
ysG45EZJQDLjM1D4u8YC8TLiIEOUDyFfUbNssXF6khgEPrdU97gzUzPJ9fHKS3UaQV+Jh/xObfL9
uuKaC2V9jbZYHiz2RBBNv8+XZUZv0bKSuQSKVFW4HtxBiOnQQEAhsEeYWQSzqH5sk41G3fmO3Sjm
WMCI7QH8KqPSvK8oB9PwSb6W3zt+Y7Ex5OgTAGI99CZyiO8dU3sqmCC0CQR+h9HeJ8gnlcFylZhc
4QXw7VVFpWy+r/wTNwubmPJM0OKQ0VGXbDUQ5HZ9CLjAFBfQB1LFt2/WyU5JZKrks5jmhAAlQCs8
FDLEXz0VGVIAwC0Akk/i3Ci0YTsmSDU/xGRCrdT5hXX7+pEGqmJV1XqAwK3L+wx6waZRrB1kgBvG
upifBeI9UdF+vr1RCb8eHwnTb/tUf4dvzTp1tLFZWoBiWwkFfCNOOwAN0ywVng86LJ6eNfNM0grd
BTrpdmlzb2GIFNyxwEIf5dzcZsqt1tZJ7wF0t0DsIm/A1wTt3jByhs/QmhOPfoXGHe3R2JqdzliO
4360SKW51gllaPtTIpvEZ2Ev/t/bb6LWO4aofxoVIu8KenTVQl2icfCKhdfJla6v4eXd++fnvUZY
OPcevM4fgoTXNxvMwVQI7jpHy4Z+dgOBvAc28IVHpqftf34IfHkLNCStryF7uVw2KZpYyIu9Iy/3
/WmxAT0KfGzh7RH7gKXYaUoGZn0iv8/jA5rHEYuo1JSBID8XgurLfw7d4v/cYhbYLRBhHQlQH8Kf
9OlagkHwkpms1Yy4337aESWHW+1SyQ461JkfbfInhK0t7FR08zwRztgdEtwB2kEqnQSHZ+dio/sZ
fBRQPALCxOQjuuEC2YfsUuRIuM8+lPOdiwvZIYehz8uGhUBue+QXoyVh1BUxNwie9TtGbl7PD7Hd
HfeNA29nOsPgnULUCL1zcPOom0rF/OQ6tE7JxZ09RKATo1HIj5qEhZGNkM46jLq9afiJEO6u6WaQ
buALFl6RvcOeAdeyxXxCVZhK9o/Uf1pyR7Gwq1sjr5ViLGnkov4JpJLJW3e6Ctox7z9wRPfpfV4Q
FD1HpI8VOKE8EFuM72TFZHb6MFaAASA1hnavT/fA30JRaiO6Cd63OVl4d90mtn3TLHrI7ctZjhnv
xHVDxB4dbG/Sthjab9b1zPCTIKSlI7dZFHZTmlTZxxIUuCdwdxUNDXH9zv7bplQAx1fmQzX/O1q+
xb8z81eBUA0z9E79GH6HRdjDVNXcaC3dmjNAd5KFzh3ZffwaZbDkt3ZpH/Biy1CK7ausqtM/+Jhb
IG6pudcEvy8VpFsiZsgLMvdRzMlSIRQBUpgr+Kpgl9Pdn4OOzggHEd44d7FgUTrwfWDzsDkh6AaM
LNGA3aeWM+cepgcl4IvDpOcHa4k2DPtHdKUdr/JvGfQ4jI0vgoPbdK6zAfwJfjT03HI1tW7xkNYd
gWJ6rvMQJvaVRIksQ3aZtac2K/+TEoyvpXcZk7g7U7zYqV75lXRRGeOx2CcDs6aqBgnQsLq/9CZU
TJB8shlY6MRpao2puxp9QGnhGHcRAiNBA1t2ZMZzCC+8dXBIRMfr30s8qV4l5sXbUR7l1pG0Qc7+
Pki2puajF4mZpiFT1AD5KuHTY8EEcG5M0fg39v4ZxWIGF9QvRALZ9BEZvympFs+fIB8OvNP2iCWr
RKa8JPHn+lrtKWGCW7Ti2kotEE/UAl2CS1H27G5dFGVmbbSrhmz9MLrzdqFTnNreYCe1XVIve/FY
2C9pITrf2n4orn4jv8Ak8vzwgLwucLlADkznUJkvIacf5vVElZlIDhV/qJdsVj2Ij07zNtz6wMst
udJFaD5n/B7VRCn5BWToN80TJp1tUGu0yMZ9YC6OXSsPM4tMd/hPQNlzKyHexNdQ7C7bJN0A7dYM
Vy8prFWRCaaMk6gFjd0KC/03LvB9j5cuM3xX9MPrWigNCbWxkf18yQoOhasRQeWF/FrHdOQ+Uq8P
+PIg2+7Q2Ex4Zj67Yxdx67hHaYSzKau0S1jVRAn3cfwm2bkQ5pD+FfmGxvYSQuyLRCMo2j1jKR4H
ZX3p/XC0IHZQlAuDDTfcysweZFnBM1yq6xlM4dpR4ipJfOHVKGaiVLHWzr9e8GbquslM1KUpcPg3
mp+izeQKqb/XZs92ItIA0/er3Q0Q9hfJPY/ulGh0rHrVlDczaswr/CRpSiDoMGCzN004nDtadBZS
hy6x1Zj4ITO4WKwF2su+rbZ3/aLa3jjs43348sUknU/gdmiJ9j2wDcu7FXph+SL08XiJbJlgpFmF
oAM8pcx4KJNJtAap9vndLlAehxRIBmQKls4Wr1hHr1atv2DHn3Fd0EL+8svlJjmFzuJnC3gxtFML
E6Vh2EeRTQy1zq1L1dEMLJT4OYxqbYZd5qpUljSwKlR2kAziD95xy/OJtWo3fER2xeB1A3leIVyZ
TcYacYuNpPltqU//+idahHVjn740U6KPxH+9ry/VsojggQwkjOgFTooVTKvOCaKc2xj2fUyzYyzg
+5ePva9mjRhRbpXsMzHSjNjAb8itvQQkK4XbT4vBMLnlrRvxGmIamCKyQ7EFl+swq8BtNNYEZdd3
2IAVwNdZ9WuFSSGZddXtb8AD+YiFPZsKNCC71DT/UE91VMTbBRQzO6OSAe05dN56GtDHtd15kG0t
4rwRm/h76Gb4ViBMA5oPpIsmhajgLI67JTZmW2OzHGfFcTY/zQpvngI4SkBljhM8J9237E1D+lFH
0ALALlZWxYKNJrIShHzMadZ5tWL8Qy7owyN2CshIQIIhBsmukIgD4RcJ6vihHtBA0M+gMIz4QJqI
pZ0Tm7WAvZ7mYzLVyk0kBujqsmFTWZPNLEREQZQdM3YBAeg719NCyg63FpTJ/HkZjkdD48g7GpLj
RNmHMPXTfkdbpAP5dZmzOgEDli6hE8QmqbzeUgFBOQNe2OKFBXkN4JZnu1fKsBcX0I1oayvmb3iR
ZwWIXp+Nt9ZD+Ku7ujEndQIWRgsKNp0E9NmpAAApHu8pocrGCkw1oDHXF5T8ZGrRDByzPvgG5i+u
0ErtjPkHXoWxHtqeySA88GflrEGfNxgIFIFUm7B02d3lRZ1OZpq4vUCfUIF4SV13MDOnYFkPZHXt
HXc3fyzGPvxK6n7iK6UgeQfHkJ4SlQI9Wo9PT4XMAuGwdqT1dsNr9Ri+XmafJ+LCFrPTGWwAr564
8eC8Dtn0AxDCp+4ohlx+zUSKjg5fO4Fe1gYMNpArE+6+Z+A7bUmqFMAX78WJNQwcaRsNWeKLqGzF
5z+cjkpEATlL442PSDiCXAEBCYZIS03YV4jSUpAaIpWr+godMnM7fEginNpfH8SgrYTLJbVo7r2K
XcnRVkQvsNh3Dql/YcwUgNMT0ACkY03KWCVEbT7x1yOYAozSKew0BMz3lemrE0bd2OdY+tjhaVU9
ZIov+b3I5/7sODqrs5iSIdje4pkoPg9FKKMgZnXR5/Wj3D3nyu0k+QWwkAcxPIGbByHWEG4r1W2x
B/WwYVVI3W4/L4Iw1JFnsNTZ4b/bScIxJoJhn8EcABRaSYchvduJB4a/e0Adv/tRWH9ElX+ZhxQz
RSvfeF10LJpJKuAMgEykTJ7ihp8d0RpSFF0h21OGycKnRvGkhTRNmrdZBkKQOPnRH6mgIymvtcHj
pKGelcHu4FQugHEQ4zcy8ImOg3o3lkjel1E6caCz1Rfzfu6KC/D6ycZRkBdIgt7F5zPmthtMcZxG
7Lgz6xo+DrZnp9H0+Gstm7ehwJx3+pHWdN1OtlOvU0PK65brciCa6ShoaYOkx2qjQbzh1NNL67iF
ExbW29yZKY+PIm/zyT1BXioIlipY7PnJ0rtGEeO+ji5oAWpeIBH0lpHkFos9epIRM/pdu5po7gWU
RQT7H63xJhi8f5sytTCTwSC9FipyN46D0y2eWXvLmHpKgUqsqOXAguNzf8TIbs1CbotTK9RtpCHD
05cBvdHgzksZaGSyned52Jy/Benr9YZklogLAVGDMLH+J9ReAhV1tasv+x25CcInLTwKFXPVSK0d
c7WI+2Act+wsRc5wLrH3iYzB7LtQwiDWopIQzcnsiHcoHlsWZEXcEfNtPn3A4fG7pJklYKpDD0ZH
0hf2qCeLQdWOD+z0Cw8C+GWN/cNSqLM5sRxdGmNdS2boaMJjdhaeg150+Dps4//4yATtSl0x71y4
XMk5IZ6WKA34qAEAUhqQS993mH8FqXljb5QYLDJsCVXyLSrIIhbNW94xaZA6UdCNc99OXK4sdrFY
D3lv+7ZIVR6DrJFlhNli3y4ImyO67okCXNAMwwfhmaX0yAvVfPUS1BqbFm+117NJaTFjmVdF9s6o
E7BcP/+2lx0yWSJEcjU52AAQx3GkSbJJxRIGc2qmUMBvUI+AUiEJrI1mjS/FoE7vP4+Dwt4xIu9W
Kh4UyNl1JLKlpE1NlKr/i5632fJ39LQaQJDkviqwqchmLla5DpDi+bTXffDxE111r0nSJJqNgSiF
uhxhYOJVOaNhoSne1jQMWY/uXCLogmflXQc8uuqgX5WKgiaohanzc15tsXF08UZnM7qRjV9mqith
bwFFsPPkqpor26cm2LsF4PJAFx2GSXDCv8TrPqcS/5q2zJNSMxVMhMrGBucfU6OphfcoSwZ0cVyJ
OScQLabs+S0vNPsVSCDKh19wFJUfXirgIWvFE9+XhYoh6k/kIy3iuGBvZKxSoe4gCGIjfqjb6L2M
MIiU8aGbQudZr9rZQThMkZtnJyu1mDiY5HQQG/1Q9hsTGc0tgPwMkgnAdNn5r57Eh4eDTuXgruDb
oaVplCD/v8x5NbSxXvzgG6nkBXjvRgDstfGK8p5+kCZAggW0eu5RBifhOuXapEDr30hX4IVguf78
NtsOyn9kcIu8OoKsJNKlHtGU4pmtonqoOQGmQlMCtP+jqyNAXB05vQo9i/Lu/dmfr35KvEtXMZfH
1Vk1wUlTDbh7khHtQSGbj0juQSXOt2VbEns9ObdrvdL1vsuGCDUsDQYCOjNLyvFlzOEhu2WwWAtZ
ez2YLXNNtDwiKs0KcetZGaqq5nyHLYspT1jz8w2HDt2LFUdTcNTE7BbAQPUsouIcrlXKJzgckwxn
qyikZpXY/7Zl9CZ8yCoqvDcnEi7fzK68MaFayGgCcuBx8FdHZqNOoM0RADWOikFxrF6Dso/7ccon
mxK7aMrRwTFdz2W9hJeQQkofgwB0LWEoDjNOh606z3OP1Nlgo+yUFKqAY7NvxLnuueLxwQIbj757
8ij+QiRy+P7mimoMchzF3O94+7MBp7nRklAUOJgwdj3Rhu3HGQkpp7SjM93uO12RyBiz0ebc6O82
VyH9dSKS0ar5Gf4ReK07BarS+EbYL35/OCMPVm/UxXlyw68TrQyZI/e28VcvAomfD7XtOc+T38+y
0dq7NhPKWWDfUF+fyeoQzqJSYQVZzxEMJpLAKmpE1GuP9G/dTyCvep1A4MAmmPgOPPe/QxxRjLBx
f2Tt9KTvuASWJwunKh8zMj3y1CHu6XauxvctG7Oyg2gZCnAcn5rlPqVuIj53HUxMgQ/mHUwQCXOl
5ROkdSs5JBH/SrHr201g8Purof0l8ipzx+6imy6a3gVpK2Ht+ehqJSH9xIDh0IDdC+JKBjSmfCr/
9iwqWcmSggYMWFkYvHiaJ8jmvxjDMypnk/ELDUokqHFpcNifHtC+6YG8L+Q9cUXWx4gUTe6rFrbX
WKUB9usrPzD/tdPVHVTKWjWeBQelnZhmdprWaW1ic6st5jo6shPNH9fB0hgzcFlUNOuW4Sr5tbPw
uOJL2wVQKB6elKsTacga9dxzlh6FnzHMZIliuJ6FuRaxLf3DmD22IYWElc2Nv8avkgQvw+8RMTpf
FsdBZixLL9aBz7+SMT2InoLnilDm5kmBQ31BtlI9XgrWs9b0+WlxHkC+X9IWM9qjDCzoCTJVZXzS
ROKWkBjWRTruZoskDFCzLQwASpEUTxPHsRgxJasGdXtZKf8ISQZrryUkEwlgl1LHXUhfaD5+hBhY
iHkPDs7UQL4DzNhNHzF/fnrytzw49E3yzL20ePGSb9GKqbGBc5Cj4flpNsurN6qGV4+VAFBL/xit
GPok4QBfKuAHk1lKaIZKVsGNU5jUa2dn8+GrKGQayipS9MaL7s3AkntqY8BOevsQGeRyGwLm9Zef
qRkDgYiu2s0vUlKC7wO+wucbbJwjvCcMqn4gELiQMrJRNMYqTkIVR8b5z/lkRme45JhVs8mbFxk8
ZYg7Uy/ZgNwXceATy1NUnjAq0J12iLJqbN3OOI/zPYW9f6hdNPxXxhTKqw0zmpjd6GIar0djU0WD
eF5JUmkr0OpZ1MRPO/3d5p5JdF/cOv6C4I4+ukQzSNP2D8g+tcSBU3oeh33DjZ2NLfWzb1TenGAD
f2dUW1ue9ENQe9vlV/zTSEpIiBWzlWsR8SGRnPEkXf6mi96/yo9vL9O8orvkSdMAY+8fvRaF76lr
OMuhQ71xUV9loKt9ZOHWQJoHSHw+XQch0G0NilTLUMCZAZ8egrYjeGl0ecbEsPQHSalD5E5qtnKd
g+CW8DzCE+uxDWj6jqPwDkzqyq7kx6P2Zo/XuwoxDQyGGgpcvtDejz4uFpCB0epXbsWSMXDKZyhd
VVUdcdRspGw3s02YOkUbhuN16smOkWJ2Mtnkfp2KSe4QgqQ+vFjP89QP6GwDIH8foFd6W6sGeAK5
RiSv8JPrPWn4MJNzRFLqAhRNzMFeK9eL/A4VCFM4HZvd2iFWe+Qb5iWqCh+cPKSnQ43fWitaVQyS
9j400T6v8i0btmbNFwhneqfMM6U1WICgb4uoPCpjiUp2UNf2niukWZw1bc7ELaZn6RMPxEoWsPPh
bPQtQHzWwR6UIyB9lNYL8Wjzuv/OKBoYH6D75k21pX2AgfzQAayDbbt04j7ShpFCDjpSnKkUPJVN
/EqAlWRYPVNYtT4x9n6XhT3WW7+7HJFK/SIDp0iqoBp6eeOAQ84JwhTBYH5KsEJx18nFrwDH3YMO
hgz0WS2nOK3KHg9RaMtUSnsGqb5UswC8b61rHGnp5jRaZYbWDqQsRtboSFk4wTCdRMWDPHk6Q6g7
tAPpicoZkcpI1KUp2Rl4MqJFyEr+gyXTh1t0CzpSnLColZDToDcElLLKabsfHMjX/Eq/V1zN5iXT
xze2/mevvX+FCbNTDcqBp3cTwXmE7l/vcKf3AgzzuEkMdDPvWIzxR1btQUB1boWiTAMfEw1VtMtV
E7Uu14XIIA+f3oV5HvxnMZhasnH67jkYTIPoFU1AVG3KEn6/VYJ7O1RCS/J+BnH9AjTKrMnvtb3I
e32oN2aYnIBGVPolAFMIzVOUM87H8miuS+rRU3DblGA80uM4hZHOKW0GK5Bpmcfi+1EGGe0+2Qz/
U1MvspW01Qoyr5jFV+686vFtynejeknfRbgbCNC9zJ1rWQ8DhY3bG70q9bCgayK4LaUycjGiTQPq
NRn553cK8sjbtbKyoKzJjIMRgYmXN1zIUqwb61nawMngO0n7kIlatNb4++IAGX77jc4pxvbM5EAN
CpJ8u6Cqr4Uo/fzArvCytZx7q+UvwR5tAnffZm51Jz1kHCY42i/KREGd60kOFiC+f6M4kST7gPX+
vEgBC2sljV7Ye0KQTamfQ9f0SL+RF2ewnRva5rJ40FiTfhJb2Y590zI0p3kC71J81jQQ8xz2v0ca
Ra0p6TM20FvHXJp9sCJ9MO7x5b4cvUYOiN37GA+SEBdZNItaKGPHeCOCCGNbDvI5SJlNQG9HO87T
JOGOrbZAt0cxfbbMa4cvK+Juc3IPpcyQ9HHdKoxEupBWTjPV7zw9a/Y5tEts64UEC3dMp9ZUb11y
7PByEnGPK5J5Ds6gRGEZzQSTU0jLVxDQpZxIMmqSUHo/5ZA3LCfA4yGSP5zkh1VYtSk+svY/mEX3
OIIHi1iDK5zkT6OZ984ujZmNUcb3Gjba/JGopoANV3Av8QWaATjtdPkTVz7BmfPVnj3syroLhlI5
XFFmol0Y5bXkDXEj1yYQfRIDdKO/CUYD6AmHoAQ2hndSvEfzvPhmaLcgOzxfuEXtxfKrH9JGDwFN
bbF2hL9U5sRTcepruV1kC91vui9LVugsteXdp432I0TDaFoX736ZsVli3lIB03fpu/NNs//hjxTY
kNZESM/pxVbi+xRuYJ6bJhwkMrZqWEYtw14mLXVNSNo2hs1j46kzdbN0zZdxwx8qk39HMl9e4OOm
FTuCBiuAMe0deiMrszVKB4CUqhbnotgyc88fGO2otYDQfUOt7m7uQ9TOlRolzM1pas/QdKCPU8pt
J9PJ/nIBpl5utDlw2MY56enWHxA7pSMvwqSgsipLImSnv8WCnSE9T9TZRMYszqEYDMsWAo85zXnR
xVGCWMPEizSTJ65G2kVMbGxAkn0DWbG8A2Li8PfX62ESDGyL3Lmii88+DWIVNtRDdhO10QEu9M7k
QfHPj1nSvyL3/gsVOCWyo0XjuB/srOqU+LxKZ7ZEJszQ0Sxfavcb2QLMBONqGMcucHC8CxsBOoIz
aab3F9xI3r4OyQrD24cGaSQmXnNx1Rvp5UJ7aUj9Pq2ztHQyNQHCaI31RF28FKmNVUykCbED/D8q
iyCAkhm0q7MfDeFz3XH3pEMjttlUblP6T6H0G5FJxdjZFzuzIZCvLcXK2bNBSTA69P+TSZyfVATl
o+M+/xSIO+WPJLsp7tHsoPWaxiRMsIo1SfO6ziCox4ktJfudkmYmLbSYqjKkbPD6rRYE2sTHDBZB
QR7q+lTJUWt/CUO8l4ZmdhQflpLIQR97SlMRzZMWeSaLyVhCpkkULY+LI5AY7KtHjlqDcpcKqz5N
/ffWfTkXUvWRnMJB1fVWT9Mk5mZG3c/EXC5nA31jY+Z8BKoeajm7UCJyUft9r0g/Zzcr69Slc3nY
U7Pzmx1yqOCZJqvqp5ItQSwL8jnjW9xgcFpbJtZHF4+Js4ByW5oVItO4l4MYbRYfB1F8jtQPX2La
zH/l/Xq1CigMXAFR+P4VnQKjD87icSBy07Z2Wc6EozaVN2ha52uomlNy/cWE8rN22ftezyOvJhS1
6tj4LOJqCt/Qlq8rPLB8zcwiDLwTMAZsGSCOz7V1/PJk6AdwMvvD1lP0ecPHaP2nAWcJQKsZ7sj2
9Nexv5fwuWv/L3DAA7igYUlEFran4L4eZ9xnx8mtH+EQLxsOlp2YaBJp6Gv1iSsMuHoHn3TsUl/G
kDG1x1v+kejCrDvmsKblxgJbV3gs114jRozpVBlxG6qIf2IbV1M1RXl9HVwQ/9jX35LXoE52kjrs
G4AqX4BmoKaY+m2MfUXgywSgAc6ZgQcy+2o/OTDMboP6YIGsYA5+mRKon+JOhjMLIRjGoA4bNmpn
j2rr59rdgiMr35ULaP6NYvMs9mw1Nmom3XKbcFL87UPBpyS5sjHJuGVn1+oHK++3bM/VbLIOicFR
AnhxI0CE7hIddhT+PtwFAwx/MVf7U2OsvZyMH0keYWvzU/OlkBn4U//54vGAfCcUPq6wDFSNTo2k
dVuOxe0GTCSqnknKuGfKiq4JByVzT0DjXHJ6b2eF6HVUXXgD5EBUqNbYuhe+/Kj2kDNKTy7waPfJ
/n1knU0fSaYYjhwJyY9I+F6nz49Jw9twW+qTK6q0FtP9DLN6EFI8JViCuzkubFD+NGMbHKG+miLt
iGY091qKbKAKpL0oLJvN3BlCvAHCDx5bDutSUb4xMeJpaNcyLBkHeTbkaA29Ou1qpk/cScLmcicT
YotZ9RFcAF2UNnqVyjel5aTG0W5zWcPieCiYjeQNLxjqezCpUIp+NuHitm3vWb7Bew5AtuHYP9PT
bQqW5seHMQX69qYhL0CJP8pPuVGIUSHJIppyussgZFa8L+ReUWvVkO61qMKsSINgJvNGgkbujRSc
H+ZHNv4mx6XEDVbut+ii9tZIPOIaNSMHMVTIot0nREnWBMgK9csdo9fS6TlMZJaFc16FBtJ+LvLy
niBo6j6DGdB79LaJoDaOyNlD7hnY5HUvEiKD+Lyjer2m+2WUzYKqvmFjFQs8jxtJcWXO4vm9drej
mPw+xmudLEg5Mrsap0sgC7NWZ3bTJn+hL6Y8VNoB40M7wH2coxKC44uWQGsqbBFPGycivmzjQtq2
+UgacU6tJ4vMaypV9VhYuVQ9SPwXcXS7Ds5vbbjn9YT8zKemS5+BP/gq3PkpfYDvo5SpIxWJMiKs
l7TbDRu5MIvFpusMQudKG45vKsmk8obOl2QMeEtgXVvTz5vVdc9PpDIxpaKLRi3ClKrHSRHws4ZJ
utoqb+bvWkXkxgFdSD1IBwUdZ1gaJpdYioDe7OvpT3RM8BybUjGwmUGNRRfP9fFKduWJ4xop4hvJ
nO+ZUIbRwgY3zUPlCeQ9WM6KaQWSEPf261jThwI9wXmr2/D3PYu/ybmOW8nsZPLxpgflUlO95u+H
SvaNuZt1mcsYDISRYOEHwM+9Yj86R/KO63ZwMEEjpOTOEEaea6vyZsUeZhQEvMuv52guYf6iMbY6
HVsC+EM/P98+8PFRxuPpsP36nvpKOFIqDmCFV2JA1Wj62aRXXXXxVq34F0GeFdv6ZOh6T0T43tvh
RGUUb1afQONwWH6EHNpgnvPdLlTP7j+f5tqxV6emYD9XvlfDgKMU5o6FBU3UFVyCmOnqPpkbhLc6
et3R3RjnAlJ5WBbJhrj+5FqsX3MKNACdr5Y8b35TNxw73A2jsh3MH8YGbqouNHTXfpAvzxFKPhjT
gtjib/E3sfg2MyYN6PRnIDR+nmnFTVwmyGTyVYqnnfFhawyPzFmDY+RBVC1XH35zg6qIRrNN6xq0
+FfTgDjnMpbvccWSriC1A1ft/7sSsoYZPEwzVqn2JLH+zgK4oCCFvhHD2pK+aZG1+x+WK9Sc+AYs
9jTsKgJ9viVOAj2Sn+N9ME6J3X2bcOB9nuD9IZEUfRcTfXmcZm7tX9TbV+EKKQiBOmwihjn5A8le
CsHrlsPxZyMn+rQCYYGkno7jBZKv4n+95ciGm3zs0SvJyHQTGxG2wrAA2uYZn7HJnpwrL/Rq2Dsx
/Xc2sHtX4X2tg57z/OT8rpE7eq7vP0Lcb7CQup+KwGn5cKYDtIpNKMva68ZcrC2AoTslkfZ2vlBy
aiQDK2hv9w1R97IyXzNhVHT1LTP+k/yA5Mdp6mhwapWK8qZhNdCFRVPcenUk3wTJEoUXzVYikMFe
KEImGIfkCOodBvHlr941XlcDLgtPlVdP8HW7YMCVI2vD80URnKvRMDrJkTbzksr9YcN8GE+denJM
6X13vxsNaj0rB1IlyhsBszRxp9gvoCt6UdN2XfTmzAUO2DJLzatX/QcfAQ1k6YouuPEzBOekJwaw
0RuSpkGd4tQJFTLoic5qMDt23GYsCVYXEFSYY+yqfrUtUjAl0afQtIG+ACs7jpAKl5inbz8tzHUs
ZDaqMS64eGfF42qwfhDWTP6Zdk5x/BMc+ycspghwexMzZRf0fWuXjcA2+HUJ2av/PQfqW6Ddu8j9
vn6gl2mYBl0/lB0Rs1+5W198ughKFqSWsA3JYdeAKu/556t1hCLVDSW2DEJc13oOTtLabPq1MjnT
6nRz828YRWE/GGlXbU7WGl/VxJY6b68+hrKozjwlf2YgCiAy4Rt9hy9qLa5HW2cEurggviMXOrz8
guXTc1qRHH6kJ9rrrdbXShbLkTIdgTd1m1nvbwW+fZmMYfJjMomQ1EHp7Fx+b67SdR0ZZFbpWPWX
5RbzAnh7bysO9N6U3+rJV5nQpk0cprQtzl0kUnyJABArEj5TnZPNrdwxbglIwvT5WpkEG2cZK2cf
uMqOX0hENNlA+YrhSoFMItmrlA3wNea/BsSmjQRRdaoslLtnMFBsourd+UvEZ3fCsGO0ikLAYvNz
lq6ncBy0/k0wsUON1PdDTRV/8TumcQLbpJVgvTxdQIC+keRUQNCP/3GrpWp1gE7YPk3sSmgIWYW4
9bITQloOCJUV6taj5mgtjapUeQZ4aKf+u0AP70h5+48TEDIbtcsQBB7bXjE9GwTu17G0inrtrhHJ
74uXZL3RKCuB70wT8XOTc1GDjWVe9F3bCT0i9bmeDQVsMdNKtVcjAacYnk/t2nILZ9azqUqnIDkc
2L3+TGit1U5hr5VVZXouhkMC5Rs8bNR2wgW7UPX648jtSTz0+fFl0lGwynIk1VZ3hshMYSrncrVp
29WsFov94CIwpcMGGem5WjOQsc44FKw/59HkOz6AngA+SNaHD+4CVEoTjP7Z/O6XrxitbjwN4RgD
lOXkcVfRrsDFxmDciJkvAOJvpo3Gq2srGqR5FG1c5jXW6CAzEobwliQCC2FTParcrNwHRi+52S84
HS5ZC5/1Wq0byK4zfVoKRArIfKacF7nSFACunVjAVURp8vBG7iaBUXWI0ChVfOy36GUvwFP/9x0L
Xr0Q6bVhVxlF4Tro98Mr6b0h5LQqsc6BcXRouo251dlhPYyjrJMQ+lURTBYJ+y0HlmjDR68wHJui
gpIqhkEDPqadD/aWEN92AYssxg6agig7chkzGUjBE1tOpEYgECxfGnvRbPuHffCld6khnu9uAMJ6
Y4auVriXTUZkOLP89WiI5+bk9YF0hvQ/vZXZwYB9JWu2qs30zvxnri5VEal5KMDG/UgoKrzQKBoJ
OmKVhJ/ni9FLHzNOJS5J237jxd8s3WWsEy9n4dW0xkSsz7MpsQCfIgRTaDvqXAcoKhrSgIPOU58+
Yxh9jCqHmRwCegQevSCuRDgq2E15qo4kS5qqLKGvbW8w6ORKfdtBOlfEWgBwtopiDA1oM8+wUMZ3
0G/z8ayDQ/o3WBI8FCJa++obJ3S1+OoTy5x6Jr1tVKnixPA657ZIiuCQmrNStN8F5d6uMDLspaTX
zXvFiSt83aR1ofLiO79PvdgNFNUcT0qSxyJz8acp79ZVUvgrfr7MDef71ttaqoSG+7TusQ5iv1q8
PGSSLQqkka8vuQ9lEFhmIk9Gad8i31GrzCthG8cj9sBm29rM3H4q8kPAA3HSR2wB5tLODwwO8Hnh
PrITNGr0mTFQF8S2oIoPDxA8PDzT3LN4v/zhVMEndrEjdjyZh2uLbbjZubs1hbEzxjEuL0H/5YME
RmKUT1r+1FgJpkP4bZAeBnJBLU/O8ajmwmhh6icI7RyMgxBFHwZCGEpfpt3ZWaMNMIGlfhqKx2FK
2xelkdHW6FFG7IPz/gtlllBTkB5OYYXdmMvZtSV1Bout4ZcXkAARbuh6uplvkDwJP+TGGoXa+2mn
SsDFW8pSnel3Nuf4gDKZUekV+Gl2J4nD9l+dpWIMrjBCcWi5sRFXRrdOcvxvORmKhz1fQIbUxbRK
4YDmckExUhCwl5Njvh0AUOEhwY9wK8NPfrgz/kEQAcSn7L1RBAAlNvY9ZHHORo1faomN0bc1SfGK
TP4hKOUDmMPh02LDpTQX4URwXkWyeY0lBhR2jjXwslOcV+G/QeKyuXez62Ii+Ytfi9WJw/++qGMn
j6c4+VfnmIIfMXlW5zxvHQ0gX5oITGQOy6033MAef1J9xyuJKNHF/eLRgAzIkMXzU+yBTtctUaw1
RNO/Zi8/K73VoCs1Q1yjBzc7SFeEosbXkamrZWavd5FQ+LlDgN7LvtqkDujVDWBBZS3DuP0RmmHh
/nDFgXWTyKzdi1cGMoaX7OV11aZUgSTXLD+UaJYsY9JvH4zDC3Gel0MkFbbK772IJic+naGEy3JT
+tXaWX9YHcxXQ/F3Z9xjKU4YajR7ZFXMUjptaisK+C96pxIj+AKl458SrBPT+nFNDKumiI/n93Fo
aUfHR5+W8mxabZwzyWqk+vMoXrhGCVuhkwtDtoKHJgK99CqWfPod5tES8OYW5kaAw2Sz7cp9Xpa3
FSBjXy956MWvHZfw9aB+DzzOiFGVDcqaEQKEFYy1nBik0U8dhL7ZOMUtKxdoNX3W1oLxWjX7xNse
z3YQFMlEGj1BGbQ3pTciZPFElArA56bwN7NQ6XBKOLiMDuO1C8WOAT3BMBZByTo/osGHK/hkxQWG
7CW3ciW/HWtsq5amXJtn3QaE37uXLhUjpvJnqJBssOTHAxaWljinm5ejdFaRKz55MxJnZnbxpvGX
nBUoxz4IBYWUaMBmcoo0RHrDXXQY0bcczKNFEaGuGDnuHb1mBmFqDbkvjkd6aBvjCtjyam+iEkUG
RjH0+ZKrFoOzIR08ar+hCNRAW+3PZuApM9uRWbYMsGAFpEr4wUaPsbMK9q4aVq5hqkqbJJi+Vi0W
hnZS7ND2wnInYgcBYi3HuBCvwOxLgQ7EDBteoa7NHoFEytRAKjI2BzSzHzg+ScLKt6FgO+JaiZpH
9W4eeFBnVRMCj42/8qllbCc7RLHaolzmzATZD0eXsfstTo4hw0QfirMDf4lB04hpehSMn9ub6Pt4
TUNcQ7HbiJh9ZR/0YQfkOTTdfqny/aDhXi0Q7jYUQSq0JAlybJSGq6Dl4yGVYhM1j16Yc09gA8HG
ZRQVcBiu0wUXKjg0BffhocHT2nYqbDYl5QDNB/qKM8M+zozY3sU4hq4JsIciK4SSUz+00BdRPTDI
p4EMl1eveyJ+gcXBbmiOut9W/nAu7arXh2+WmlGN2HOAV6e08Fx2VhRv+08wNV2jkmowUbjI+rT4
QOmC1Pe0v+RphIgfxws+g1Ct+t6TNy4GCpo36clxuEXRgyW8tTeHOdD0qKP14N6MI5i5WrEoSQSc
omf9gCum0ydSwFdjEM3YTB0l9UubjJJSCjMxEDJga3No7tDBFdTWzK0WrRAZ0I+IwpzzJFBRz40N
r/4VYJB+iuwMJEk56Nq/CIYuq+FxXnsm9eQPkT3bZ2nXmpseyE/qoMHDxXYOPfaXRlZsS3PYvKoS
n6+CUhIT1VAk2enKhbyOfm0P4lcJpRWNUs2UbaVBXZ1mkBLaEGD78+FOl71hNsQHv1fq28ZMdPe+
yhi1oTKC6l4SsYJKN2GXQ5hdE57UagiW2Ov61LUk/+Ui7bY00kf+pdPh62dBfhxwaf7AjZYpmMOg
NRJRakHSQ7dw1DgIPps3KHJ8MCUCJnPL8H/yCwLMFX91Z6HcLntU/Eh6c8HJQ3N5u15QSFDXhyUc
RSn/PBoaxzLIXQwfiBiC8YYvPr2A7s5hhpOqefSkiDTAyGwac2SyXV2n/CO0oM2ugyafvkXcAkvS
cJ6yJRHobHwZ1ZpPJxSLjGXzrgjNkaoolhmx5FTbj8rwQUWpHYeTUxpebVINgmmdAJXMPlS8ad/n
BIrGqcYAuBTTh4RgmUvIDhTBnBKg2eh0wQCPyZsAyk4sL14Ubv0ajYtfq0gIIoE8Db+Ber7FdkkD
vpqWZdoq3rS7eD7LmH5CFk97xF5c6hB77T9Zc8krXC364GE1GpcNmUxpmuu1h5p6BsIuJZRsTxWs
9UkuvtPXpDhibjyTMSi7P61a0L1gy55UBsngDZ2KtYUExfFdBZhGJ43o6LEqVN5/wRGpZuYH/vkA
X4MkOBKyy143MzCk4BYrCcWepkb6ZL407gqOR+EKf6crYPWfmChW4XQ6KWzHAAmFYqluxzzM3PYj
Ano2L2cHCiBws252ILlUGLkjb+egUXUdLxsdAoLs2JwUiPNMlZY8jgeyD9mFxnYqgI9m6xzHzyyq
K82BOhJPZzun5vBh/8ozWGMLnZ0kVpMJOl4U5PL1y3gkbTMTgPeiVAN+nf0Fywru50fEet2zTp72
X78saYwKMV9jPH/wCHLFUsL7/jPyjqReom4wtWYwbWthdd1UE6yV3SOC6WN4v7e4ZkEAK4/i78z1
AUgAzFhFip4i+br/yu4MsUnbJf334Faa+Z7fYcaIW+MdvVwqfC0h4f3KNH1CPgPzqb8PdaB1Fqyd
uSJjBnnl37e9UtGdjf3AmAy/3OjLNeyWw0rXS95M3/e1yoQ283dKrKJPLkrusODLTLcY+vbP+MCU
iVbj9GxAwd0BmWLJYXg4RmyiB99UNB/D/IFiTs7ZI1qFlckfNW5REgZdjXZnANRObAZIiwxH8BfP
yLip88wmiit0HUk8aElYFgGGYMdpaBNYQsdYoS8qgMa+n94Ndp8q0JPhmi74zmKKWqKqCoZSm1wx
FCI+BFXwDX4HQr0HzWuR2X0d0GaH+SijbyfhR1G0AWEHBoUpPlYJaI6FY8JFc6quvVTonzhjJwi7
KZhNxrRSzmO9PgK6Uj6Q3recHiSZb3fp4E1vLGnk9npwqpMEdrOzO/1i8rXK3TWY4gPuq7RVP6C5
/OwZDm0YZC8hMpeRVTp2rGwQZiJKOGrieP4OqhGacmJscdYRFmQXP260C1oWnMBj49DlffLAzAi5
v65y4VLWi1KKak/+0kGb4LmgkivJbTMvTGyO/Y9o6IlFFvOFuPRK94k0X04dCRqyAs48XtS6HCkV
26WKOlSLQeIUt5PM5o55d9hjUKp/2Ibt/XGAzd/m8d+OupBdjuLPWtXk6SHy4N34YKwcmzm9Cmih
5LeSJeS3T1s/OdHX7Ha3znca8Deaj1z/XijoLCBcH5MV7MFxFQn9zlIXn7wCSXTQOs1FzDRHdoJg
NTTBHJlAiKdsOXz/tKjxMYiA+hGnhHfNS7t6f40oHHqFMxkMOhBUka/qxOBzFw8qbtU4ITv1y0nr
g50FTKXEuYggG2Qa6hDGo0P/BnW4HYyM8goaAkCECB/FsRbhVd+M6BsZM2MsdPL7u4yVjjg3flrX
BZOqSO2yiPAhsUViGJ92N17raRKn/fYxtgIXfcCbC7kIX0fAZZ6X4EdIbrMfVSZ9dpa/hsGLpeu9
M0HnAP4CkrA9hFHJQtjMRHt4uejNKzkUxtumZCdU9zuoYWzMsQJebKRLbH3lyC4m3cCtdLU4Y4NT
C9wbEnXtyz3EackIRjFDAmxfFCxG4jxMlT/i+00hq11DXQxGqoeoD7G0oMIql8nUhnmfP3Qdfu22
icJkL8TUGzgD5lCvi2xwJXgtU61CooKI9unj/YUjFA6oQ4Be3D2C6HFgXmiJ/lfQzKe5e4SJv9i9
s4jt9/rnCPN9vh5XOlkmtsOfuKfWKQZ+WIkpOOEt+EiXcYUXvjeSSYKfeNqlcJ4s9b8rr1M0lxHh
r9soWjgHYh+TrQBiumYzCfb+QDx1Smk7cZm97JSfEm3ROzYD9hIhJZapFpJcObdcvA0m8RdUiI3a
Dnz6pNqUIeaK4tM1ZJIpiXxMGaiYzspSBRAKGH4KCthK7eZRrd0pT61zCoNqKN/bWXXLgRHVkrCP
j1bEirN8iEClqClGsfcJyCQtM+7bra2ghY8pzs6L7vtkXFJ0CD7SpzL3jIZgg6//ATZvvLqhaW6r
2TOZ5Y96kA4udVnoMTTXe0X7hsc0Re92oQvE28iRmXfBZm4ARyzOlFkDXqggeCbId2KHXE9QbpzN
RPZtYN8Unkrve9tlQeL12FgjSloFKbaqV0vmmG9dQO98qy1777FYasu2TVqmcrA3u0f7c1PWfSTI
/e0UXBkxAQktVTGGi1h/G96pPqGwpGsRJBFcqlJBkDzkdxcsw1cDG+hbICEZew988folMb2UDzBe
zU9RuzWsIEIr6m9w98Aeuu3d/3wHiBq7h/p2LFzMv46B+u0DsvRtSyfjZzxq1tOH4XonskEidpuN
U/q/IM/ZV+8WAIf1IEuyYcxdatqxAQZXvVHtsnmAoSBXi0I7tPwplIugvWk83x3eJIAP0G+QW5b9
0XAZEo34jFbpws6ZOxi3SQTym0PAsI47GkYWfvtH4EBgAuum7pa0x83+Q9EwXdyewv/ysw3THZAv
npNa+dOv1IZiJWHYKRtzlYve6Jm5tveFijNscu4rvnWp+Q0VlNYz5I/RFCv0aWLsFI9WlZ71ab6H
uhccEbxsn2DgdWp/PXvllXGOcb+CuyCnN+TilxQs/g7D/O9izlKkWHNaSu7kQONtGP1Os8wxR2xx
T7IZFFo8OkDT6uIiFT6SBDxmpcf8KH34zjSErbZWZEk79xV1NEN5hN8UVWduq63R3nVe/nD0ORZS
mexkQzVjHBTR50EdFS2z5I4IxuyF1CO3+fvsUHhXerOfqWUSq5tw8rg+UNTDRGmAEknySDHbYBwt
bRZHDXDhxEKEUo10znmAxLbLGX4axnKr7MVVUz1xlSsrpXtM2e9af2alRXPrH4nyQU3Ws6vswG9C
UluWPw6KbZouWVgz9xKwXJlNLMjYAWzODzb64fCxgbNdqYy2Rr9uoRODI055mbqV9oLYzXrZu8VC
r5Ouoo4+gjRqbBlNeIMtqkI6bH3fqxD59Q/2WgsIy5FRjqra6PYmlu2f0Ib3uPr+NlGw4gP9SBam
vRGVg3afIltXE61Jy3pX40F29H8rrG1oGHks4X0JdQeFGJ6jeFTyevSJpYmXWNavFEwkzH2DYoUy
3Rwk7VW+tYkGxhfmM6zS73D3cYKJRrB3YyZisQM3ncOhzdLknEMYiM591bsW4tX3j9q6ZMnz8NmF
zAmtBOW9sWWDVvNAe9QmskUGSpjpeG373jMuIigKF1ek+kL8DeHy0OGGgSvA8gr2hAqRm2Nsd1ea
4ZlN9gYo7iHh40B726SqPbo+hk3GMTTGCI+p90SyvLuuLiYcSvM1Or+x6uwrI0iZZmc3qXzjmaZs
XZuHBZguNXpUDQUby0oQS+xk5RFfvjdpvQkhEwLjrRibFClK8ndNzndTfqo8Jt6awukA3mCuuYtm
LeXdCe7xrnnavIzFiGwlse2qEIBFR3uYiTIqwQnQbQXhgV6A3Wa1K5zHb7ghds/yeSAuy8cOCbp9
+A+Mr1Zc/OSrEAWAUOij/FzBdXw2XIsAoKnl9W/RyiUNPkkJZF2UwKz9mnEOamPIx9YRj/V4+AD9
NDZzMeBlPBpCQoMvELTW8JUCgogXBAYtMoqNVUz+r1GyO4R75nXM0z/QDu5ryEppmvBfFifHlrLI
T1MT9nudyaUVHdACSVaz23BCnU6KUl/CxxFkvZAIePxgKn/ySK4fRY8wcBCINslzFW2JYH+EKs2W
3fjfzgWLtzsUtfXOnMEvGd9R2J/BxVnH0CGLcZr2O0TrCiAv7PFH9YDa8TmGC2pwKy1dcLba8hjI
Ujivjt84sopw8JBZbkH0+RsYGR4RF932qcN1eTd1ck1hzi+P27mQ48R975CXaF+hCr8ikVbPFibi
wzAyvyUL0wIyrguAJ59bCa+mEb5GTGoCCe/NgH00N33ihY2+jSQJG9DkaCmEf+TTjBBGF58wkRnU
8ukpxrkbsREVXtk+IfdwOFuW0atGXWvbKaUeLi+hu9wPIRHL/khHp89svV6nWI9BzAMIzXxhRS9w
YikE4sjNE3WBWENNtf6j/QYJorCROaMh7QgVkCJv3dCp+nK/owH4UfRfaPqRlkb3gOVzaPiE/fyU
DkOaYf8v278v2zAV8x4HMwLcMBr/m10pqgCjI7KdWgxJoQCRFC/+HSE0dVTCx6hj0jHp7AlQuBxi
gkDEJLepgLuD66wCR2Q+H/lmyXInfNWQmI+F5hGQHs6dZbNOP6yYuxPpp1dxrTzJFyBOy19Ofz2n
wewz1oNlVcn+/z7jr4EVSv26zWaEh2TQLl5a1q0fjwWzxYU8zVTPA98PPLz4vCD3EQKblYh7nyo5
K5VCDJM29ZtY6zR7l5/fRDPnpJdXHFdeoVw9RON289Ewa7gSOznELnUdcQ8w6WIJz20ELvmxzgYp
td2O4FDXA13yq0nRnw0Q6D1B1sAPwcW1G5BRRUO1QHyXrdW1jTFvJoPeKlbUEJOuAYR/cRlglNoE
/v0eNzLIKeN/9txfsmwgN0zjq7msiMKpAzt4Ix6oVUIDdNivt/E588CDaIvvMe2KUDVSvw70eiXG
lWlxxVbqWnY2BJX/1TM6+XHcUAhQrH5ovOXkz4PZHkM79lGVzNIYcAnf9oJn82UYdpz+IjttqTuO
o6qNwiHQTisR8ALnO1FDlyDh9WjpVWgeX7POkGHpASlkBMevAKQb+8SzzoCqkGVt2lF6rbGaNN2G
EKA1qYnJgAXobGzFVgTPBVLbAGgEPVDRGGozmVaGDohFuBELccuvYU0vCaKpbVnCbjLQ0eyqLux7
TlCBHTQA7bwPmxkw5GzgN2DfalhhQwTkjSmK9JyDYb/cnzf4BIADsxk9TPk/EPdlu6oTvd7NJw9N
8UuyT48Kc8VBTbVtqetT5mE1y6D86+V/ob5YhqP6TX9D92ifVTvvA1qEOB3hyZqXwQuqmWs2A47d
/De8fhY7a//z2zvFeCuO1q2MP5vahnbzCdOgnA70PlRzp+sRVWRIqEs4NPCOaWVmfxgDuz0+t9jf
AVFZSVxL+4rSQgWf0zQfi3B0/wsWGlzWV/nn8qob/Rjnu+bF133MkkzrWIDhwXHLOW64rfRqQIVq
j+WF+tkN6GhoGPZ59VWpVg+IepRRWvaEJGMK7nti9BOgTckqpgir8J7VWaRM6PqA/jtgjU5iKbuF
nOWRsUsE/xZsu8QcCFXrjX/Pv0vSjeSIySxRkAvgBRi81BARxcTVxAUmgg5PLDMU1K04W/yfiJSL
tsU2+kvGdr+tGM0vAatcMsQ/v5nDsIugVq/YReZrSQZLo5CSTg/ePlN4YLNmJRjcwse2adNVqcOW
yvSb54QCl75NhFT1I374It3Wd+M8AlJzmeQPZXxYob21/n33tOq54VwIoNIzX5bD4nvbXp9PCGGx
yrZ5MgfbE/VSycvEzvyL1Fa5BD5DaQrGMsPErCJc1JUxtI5ts+SEZBt634mQNURh8j49VSF6Tedx
nCoMgwniChGUosUU23/UhigSxa9RG8t/phwigxXMeNksRRgHbCtVHoacG2X76fYJmG9+cN3ujLNH
ESIpT09+ljGuLxhQFuK8TdG62C9lGOLRFJrV4C4w22rachXU33VjWDVpt3lOc6l2+MkMf5QZbwn0
RBO3bNMC7Gkdjhix3YlKfsVil9ms9kOzg3dUUfhsHzyodtLLA5nY2Y6XMPNZmXh8icauKjO9bGnD
1YEdK/tc5mayT/IVdUwSuHn5YCZDKk167YgYONaRsjxrjYNR8OlsLnQCQBlR/8+aAZH44EnSBJ1Z
2v7x23tQCjONvwJ+8yNSv1EO4nTtciuSd+ZBJ/glzcgJn7JBrW0UCdqOkvz8d35VEHfB0vppWp4Z
dILH2f0STQaKbhM1zqedADWjtT0BYnQXRsHgzcQWznBQUhxBgQ8x/qUamV+oYnr4eJ0GGYgrNdAO
ybiyXTHSqRy/R0NuPmuBVxuz2RCQgjMh/JPxkMJXdH22AlpOf5ddpfNaXcmuLiSCayksIgUv74Ao
n19v1+8RQAi4/3rOht1Vv+twEyftQ0X2iDTrZxckBif0Y6SRCE9GdPCOe5p9VTsZ5+/p54zIF9uz
puYZpMozvPCxoM+R226AV7qqr17tiEPee21ulAdhyg6jTdMz4oEhdAfmzFOh6Z+PdSlIrWlSa8j9
yVYgQczuW9FUUnIgffIlJyMAPq/XfEy90viXZjXmAdHQD2wRjqMRwZE3Ha7KM1DtGJSCy87RE9sC
GkVDON3j+zRa3/YkqmNWk7GVPj4+KNRzYMQ5EG5J61N9YlibSVxU1Sh80c8CvQUa9eW3iTAUCy4a
BkU3G5eVNomDxw5h1Ui+zueqy6sC4v0Zy2pJP9NaiGCbVv5qqTM7pFOdzM22jUl6JAsgpYm4KIjA
MVJaxV5ZtsF7qq//AsALfyciNrRswurgI3g3FtOjIklmk6XyzHvbK/AC+7NTIYtuS6CEEBB4EEZE
SGqbqbVblDWIgCoR/6g+8epVQt+IzPf+nZ1BwpAzk7t8JW3RXcQEJrK4OdEqCeCVyJ7kpTPr8WvO
rYf82OksxeHEnjRucfMlmdE2HEs5f+R8vXY0lNj4/j9BiEWWjhR3zQafrl7BpeqB7b6k1tkBM83W
ZB9bJCoIpnp59VzAOC128gelug3UuLjq7Mp7AiaSWHUNJn651KS+wZttQn4vyaKteoqfmjHAwGlb
axoWfqYmg7xapZglRRhCGaG3Suiqskg88ziz+gmRjx03UvwOA9wIAzUzRcKWioyGACUIx1Gfdigm
FlmKD0d0S8aq6xCVvXX3sGA32CzF0Jln2mPEPN7ydzYuoU41aeJce41WoX6KyY6kMzUcPl/MNsXP
lSzq+lCWqpmTq0JT5Omz0xwOEuCR24T7n4sJPXItq3kIYL/jHlZGf5DUIXF2sokE7M6ODza07XL5
F5yPh+XVHD+VVUnWeM/q04KQnen3gn5WNtZeglMt6XhxILSkQ8+leDL9B85A/s09k7/BoamJJGit
ErzOG1gvF+k7orXoQmeuSkDrUPY+NztsmYIPnBY/iBtKzSM8uSWdneUzdLT0YEpDMWYOQpbRqfE3
3ZvnUeb5X3kJKZlkllD8S42OreVt68g9j5JYAffSytgWrXm3ABO5JsFrEnj93NnjmdvQvnCxEF8X
Syjltiq0+9IeoCtCSbcJZhzg0x0eUu0M+4PxQ/WuR0S1mG8k+wucOX6y+mL0+6slWeKckEQt85pv
TQgnWVpg8+kSIQlf+FQQmhIAqQZqK9RriTHW5W6jISnaM2RY9HoUtfSjvGWRKv19kYPyYL4vnKQt
ERC5cDY+rHPANfUZZNAWGlIBm1cwsC6RdJtxtLFR+mHGgtd6Y3JQulNrWRsxQp04S2WBs/16Y1/l
uii7wapn8ZhhKfLdLTxgONqqIhgVPMykSdEJXolhrVdyAiGlDWbrYShMRHv5Zo69LOaPsi+6coOk
FOyQthjBX0dwuviyE4T19UDOvsjAL+1mFl+WIVbo8CmbxMzsL7GlhkpPubwp/EUvgTSwETK0b5/4
xhuQXYQbwtQw5RxpGKsgm7SMZSDoefLbXzzguQGTx8+lY5oYpxdunvgT04GT8OBoUxtIHqmqnyRC
ssFdXxY20wi/rux3NHIPjbksqEWzCFDIi+RSW73mopIKI0CcCd7kx2wFmYJYoqcB9XmFaSSSxs0W
QUWu0lv0Pb1uaGvTbKPVBDbRtv4YQUR6xuhTWiBVHA1JGKn3FuRXh29xpX6GxY1ivi0UVpT7Db7x
WAmxkWsifdWNHeuxKCPHf+Nd07Tscx3TTmX0hSRfzwlucsnXM0t3OZ5M/5sPvlsBfAqrmJl+atSl
YV8/zFP+NIliaA8kd2CCJ6b1rYHsEgPzJL+lxvKm7gKqcsswBUl/y9hrqjsR6TAgho7emUAj77ns
h3uBZ8aYC2mrUIvKha6r6elW6CjusTTiJnVW/CAYHlZ/7RnX6mmsRgoImzBYi61VNHkA4hRnYIWr
F/pvlo3Mt5xqrOhzgXts4FX9R4YXl7JxgKTb0Au0E2FyFjoP6wntG0MYRTA+f++ZHxz63+2zNskk
xIdb/ioA230eC5nIPSyNOYTs7iUUDDmopXcaNfHhxLmq+2g/IbDZC/RSPZzLOfI242vmsESPZlN4
q/yLVyqHFGvGnZAsCUOuy7TDo9WG4ItUvuwaF5jzsMwZ8KQrRcL28Gt/aYMOJZ0K8LM3e6w7waKy
PXf9mZmvbAwNK1eq4OjP1G2Si2Vr9bZfByQMYOS3PXrDLdFnhrlb/fc4+p0CdS3nAw/cpZ/UIsmg
Q3QHEQnjSCdlVeY0zDOgPjRj801jhfBORJpN22QjpfRCbBJ7/1AXxa2YaLAadAyXC27mXGWG0JEU
eKQFXywROHA5RNARgekKLWjY9wVoVAK4AZXV+cQ/KsqXEjb46ZPq+1aBAr92aY0gMhXoIeRS1OYF
vL8bhbFwKxWXDtpT1cvX9u3ae0pWhvbLygcz+yUl7L648jIGPiK14wr1sZogfDA7gunYAh8Pc6bN
1DQf9RbHBE5gc84VEDoepustaYAVm9TaBv5xoek8jdW/9xUWmnXVpP2p5lTo2zKW7KRsiRP0L8jx
wsI5Qv3bFVEgs2nurZaE66SLGlxSVz9uLbxyotPewAwrodmXh1GsTm/mNLNMm/ZcBAB0ThjIlLhb
9qe8wj6PKTZrqiTyxUT6nJ4sjdW5MNDoh7ARKGY9zd3v+wgc7ficSrHEUb1Pl2AVMLsbkIfPUIaT
um7fp1sgAonOk3SOnS9uGaUqEaaahnXlwyqCBZ4nhL670oOYBBo3ad84yUbMWfSlkPwSclhcds0V
PJl+du/JzDPU5+nZnLA/qihiYMqMmeLYY78kVC/ts40563Z5rpUOaIlrV8XoBQMQNxUaftRTj9IS
7hT4K82K1Gjwqx7Rm+TjZuMEBfg1/vgEXfmjOg/j8LZGxYHOf7SdgMVkSGy/msjut+GHfNonU/GD
RWbyCFqXc5hhKcjsxgSIMSEwRYFzTqio1zy0SGPgcabbMPfmG2iTTKwVxlMPSUxM/qiqWDIiAOzZ
IXLyVaHPh9O7EHG/QIuvN7AvbIXMiROEkz1Wns7qq7P8PqN4ra9wbPq52x4+U8rr/MTJNVCzgq4u
U4FuSNHyl2yojT/NmrlE3CHeKbBLP/MOzh0kTCVxF1XNcI4rL1C7EZz1eECidCuyiM0O50/se9Jb
fceGrFJXLZVTzlTvjv3V0vBw1UdSv9hQ0PTriXql/FuJcQggVphCy5+myIluWT6qQWQJhkBMJJZh
F1FGbu+xt1anlNJh8pv6FhKQjURZ5c2z3u8lTco5HTizv4fAv61qbVrX0XqnGzB8LUmkgcwg7f5O
7lygyfiokS1vLonsJUWUzjJwIVO6aOG4l2+sVqtW0EWYw94Sw4WsB6uo7lICJl4BmwhMI7MJ+A5Q
grWPx5yCsdoZhbOvk3DNlFW9ijoS9y1bvMRNoW6zNg1SJGmWBQ7pAR7IKy+PJnyHRkOlFVJofNZ7
AS4KBp6O5WneCKgJtxh8WF5ckGqnasPZdN+mZGAkvPLo2Ch1THcEruBIagMolZfszkA+f7SWEhT8
ZHPacb0vLELpiEcK8zpI9iqk4iy8BMMYzoH+3HFrhbppcZsqjfmfomJ+k9w3PHLzeZROqRRsngUc
SVn3w6po5oQbZ5/6pDCD9sNVQgF6omQlQvK+rCXsIMLYgCh5vJpdGuy2GbgwhmyNXS2W1IFAZkj4
LrAphhmcX6C6DSVYAa9BhgjYWcGNr+62qNqcXLVjWAYfxE6bPEUUyBA8RdFgz18cbGM80vK3iSCN
4Sx/MgMBOmPVCgGoCsnLS6KoXsjYR+f5576LsmKBkAx+qK9r0ipbBiDQTqnI3giCdslW4PEVNSE2
6aaNyA0jMW6Ft/2eNX95OZ7Rmh4MsummeflVbdxNBrirxugtRNUU6HGdRotAkl3+bbKmychbhtcP
SkDtd4mMAGhRcokoF5NCSnDbog08ksjtS8m+72ziedeTn7hGEotWvSBvG0ZuKk66OqHEK4O9ehjv
SNoz4lOqXAHslyXvOUUhdUPvcYRAP1XM6Q4BpTdUYrcAvxcqfZJposQMCKBCD03WKHb8cfNNM22v
gD1HFCTpzDqo2TaWhehHSBem4kxFmqJHeJOCdVFyGPII2Fw+fcZkqmrRr6WZ1DTtkLYVGETCdmvS
N/Bp8w7A+dVfcH8Q1somtTKjekeDlfwpHdgDyqHFWnNrpOXiHbSxgMJzAgGHscjPq2OWvk1PqXps
YOeha2Q2g2REC8/WUGDMhdkwJYi79Bzdc8S2/Tc4aWtwPQgEDrCen2wGA7LiGAvz2tkZ81xf40L8
VAfzaMlCJBqu1S2KC4qt0by4RsBKCnboH+MbzIT79ddw+P+g/IQD6WGdRB/J9geA8LqFYcnWlzap
0jsjlBfHDlvgvIUyvjPckkO7mj61maqeEAYehA/yLTE7z+Hg+O8146OGLVoyI4SmdBs4SvUXU7uu
LuT1ANAEA1ao89v9swXiHpVRsiD+83TbcH5lKj4Tovyxrmr5Gm0VnHNgg0nN26rQJ1jzCr4oSF+F
JnjjrPPHI8NRDSmQSby2O7bvwZWkOdK9oelaOMRzkcOPTK7Kg9RES0xcwLZQrR0GITYfLxnx+4Tz
ij9fQPe3auDfihWTHKrqmcNJOzLV46PY4e0FTKP2/CT/sUFXvETpFxXXbsWMfcmrvcmm/KcA/FRf
1w+LX7aHpWmtwzqoGys7HeVs9yw4L1o3iKVqzsTCLxEEhjDi0G54j7OEggoKpYA/jLWIStfNm3sa
NTNS51rScYViSppEc/LC16PE6iDbW//XgGBoqOhjI2NJtap1rFTlA/qFbCslbOvs++CjpgijWK6X
EnP9nPsV0NdN5DtSj5Wok15+/gvPXPO0G3i+/Scoc+ywGBDTFJc9qa2dH569gxKlGTTRxHtI/NtP
BF9mlKadcAz2FRpXUagMKTdAZPbGBKL/5wdJQIFflytG329zfucel1IGYWm1s4fNpefG0YSW+Dff
hThBDlY2mpfdCimaxiACp1riSp5MRIoLvN5+svAgGgG9/3bSQpD3x8UMfCrlg3QcX9X0+p7/KalK
zGx63IHsZnEAtkokMwlHIQJdHl3Nx91HMoYzC6tDfSuHLw5Z4V1S/sw0C6TqzYTvvCEBA9PDvtiO
2YFbK/vc5tsqvPQkQojlhNEWmgEO2gvMn6zeFA3qX6sr7658QcoE5LwL9WAl3cxMpaRpTdz6kcXg
s8PM+EtXycL0PrhFEND2/3Vf2igCo9puZ+xJLMw9PrsbN66co6d2i7500RqjKONTovQvEmYC+XG9
6tn6L5m7RJQgCgVqt4VJPZnNPLCVN9ij65ROfjsdc3a+l+YztCKt44bgb1ob64UhC0S19PU3eeXI
gdScGWsD6hHJ0lbyADnbQvr0p0dElH+8/LKuzQAQwaoWPxY6fYWZf5wxfiYHyiMrU5MHlLCSYkwU
EfhGIrkbz75B/sJ565Yd5igFrh5jud4iCuQ1TZA1EBPar+JOBZjCNGTmVhptDhAqGGgS623sqb7k
PN+blwdSL6eCt+USAbcC7gSoaEW1x6HXTFnHw5BEP32A/JV1m2WLpe5RVulr1kc0cfIuv4p3PyuM
9qqH7X2ae/35HouyOIlKjxqU1Q/y+zR0poD1+rWhZZL1sY+YsEMk6WmcTatCdtXqBIUvDaYvpSLi
7HC2PYmdH7mRBqMnnnGkVaKIQbY0h2c9WRzOuVLbY39bfylKzzsDLIHAiO7V3oAHKWuixm3p7P7q
Y1tX6WbRcPk3/fTrKw3sp1Ns/TpGev+bxFmY1/col8cERLOrxTCZTCIx5rHuu2ogoJ9Yi9j2D0sP
ZKcvTMdsr1m8mXPA3tnzeBrt5SIEGlP4n0w8IDAxrJd4+WdNjGz01asHk5MssPQY0hk0qwo0pRHj
VPpWJjiO6QUVlKDhrOHDr2nMS0xI7hPsYPGFKQAXwqZy7jHEH/1ej7jLrfmsoOL3bP9ZynI9rrBS
AFCX/qRgRvocFhQBvWvWJHP1Hmj0GLnpKkWrEyfM9qlF5tbyr2qYWkLBIjHQmFlIc9LEA1evJQAx
v/sACsL/5wM0DZVb+CotqumsqxdawrNTRHDMWw4f0yhOrr81merLTNP03GcjfC34H6EL2SOh/JNG
yuGdmWrNySrK0Q9xNk5dMvTUCpQyXEVWQRAc1oN9j7nvxGM8ABSr+IOSVtt8kbhEW+fAC+DtjAKL
4WWmTfhnLExyMIKykAVhEa+NBwUlGGJRQ6roymfCNi7WwyGfWQutABjY9ESJqfGr30FxJh+YE0dn
VVCmWzakDQ6HhAqMF0fSDNT+MwEw2hv5r9YIj7+EKaGCPRfnf+fJWeGRvBwNraJtWSrqo5eyeu2W
HgZkII4tWzPyh7ASdxY1NfDJuX6lhUa3Q9Aor7qShS6O0Nq16zFCaALEW7Dqlz8onBRYi0Fx1D48
8xI8EHn2lwIp7A47TDhcp/Vo/bbqHlSWRkkBeBY8gmDZQ5+x8V+QhmFwXdu8Jvf22vyH1FcvYswj
3V5ajBStIVtNTIdvfG9mvCAbGfghWgqxe4KhH/C71NPCzW+4rei4PxwfDg9wpkQV7a7D3TI0nDYZ
pD+G6QrdE1BEf65IB85n4GSBO9ySXoOOB746QylM6NvXjAJ+vtHyot4APCmsxbAxpinZpnDLCrgB
mowLsm84F5w49pGJrcyo6+HFnZWd1FYjRrwK+YTSLvWp9UJBbr7wjranPkRqEkpy2qGZSBb9yOAH
WQVcBkvw7vuafa9zvT1VnQcWhziOXp6H1nxyrVtnAxoq5qVeMWEkLukcwsGSJM1enPyhIICMLtEn
y/PDoRWniDX4fuMfE5WYGzJMnCdrloJwWSakBzTK3wJPvCkLGHQtRr37g2XDnAaMrEWVNROkIntb
TR5FqzLbMzZLT98i1ypBtQxowXDPZBJvB48M3Wo42DgYNwBftLoW2sObbYilqvfw+tKOBringpRR
xV2K5xQbws7OD1M36Y9zNftay2sqz0UAwSqIcetY4v0MWM/30yO8WplpjZDjVCMeroDLS4/YQWN5
N40fGnROZTSdeUPAUNrIIY0NwQ0RFWKiNJmwwWp66p1Xm+kTzNAw60iDp4Qa7gWBLVcxvLvaeaYG
lqz3BMLnbFLEiSsDI8yIhlJwi+8ODjSojoRwLDZ5huSkj3J12fRVehmWlP4YjCun9PhCtHXaEXdp
XChZ9n1bY44dVk9EpyRMAlR624qj1R8+qOdmFPs1h0gDNu4KZ2qfKLoleSIFuaDnYoRrDXPdLXwF
UxGaLOZm9KDbJTqPP/xJh3MaWk7wSPMnp+qt7S1Dp3wst8JM9xC0ITX3ec9OxFhoxY8Q14n5FF8t
7ckljgoM1h09moQoel1qtNXrGfRnBaAUsy2+IfePSAFXUlRgF/ojBdb6HTFWecTbf7Gj4vtg48Q7
A2z/i4BlEDxhZ8EsdukEV4FyNltIOmVFvT/yR81gDGIVAOvg5wbcm3PrgU2RhRjZRWLIRB6NXWQa
OUiJJgnujRYclyysEbksKTIUPQ3QuRKMM4/jsHA/iHsjW7XCb5xsu9vDLVvdy+D7D4MGr3u5I7DT
R3TKEcOQ0hawVJXM4e2yHuQQHze8fZrk0GC/twNAQORWgr6ibZ52tqnj6/56EPEHmpysWZVnO7SK
fPjUG3+va3m7dE0s0JCxzwoVdBGFqKU+zczfNhmNutlhmwE1fLce83Dh7qbE9R4bMYIKaVTO9d9o
wHv/jDh3YbY6g9k0nqk/S07g13quRnwVsZ6cPuXz7Fr1OHc67lnd19E4mdW0fiTAekcWeYNxwpY+
Mwx3Pk9vmrmB9ARAGt7aYHGXMFKcQ94XMSvtSSIqYdzdKswMccvQTb8OZqtntOMCga9Z6h90NKli
TPqbGmOqOfU4Z01vXHOhjLTYu6aB06jLszp7Eztzli3dQCr4UFOBFkYeOZ5dTL/PJAsEcbU7f9Ef
8zIlDU2blLl90OOAQ7c3RsKqe/zmsq/4YGnHmRtZsoV2Kj7kkZ6rUggrJpFusQp7ZhHIdoPSljR5
9Ak3hE4dhfDcQKsNJ6LHs13mAJ/B5XrAxsDLwhuBJALBe+yMDU8fTFmBYrUZKcahY4aLnrrzvHZa
igA8XHRxytHtUt4h6x8avAV0uLQWtI1oZjhN3s2dr2Y6N6kvIXw/vvSdLrBNbD0spbVHVYx7TG6X
6/jhlPPHVf4djNwH7dRUO2Z6PCEHsCQmQi2V3Wb0zQFwWIWRm+HGGjOMkn5LMesT+sKfTY0tC3Zx
zO3jvbBcNjkFrG4KliQszWHXsI/nAL65sjX4FlwiI+oNDhV+BaiWlkaK+k7hWpgW76AZYpIVZQK7
dOya31SWDOtw0d0mgTDpCa5onE3FVujidc0VpuXd8SvujOfuptoaZVq1w93Q+1iCTkUupXM5yVMZ
TAk7GVqP+HYZ7Vp702YH9sZQDIHTXI/VF2q207TY7oLO8u/2im+E+yi+sUYdgscRTW5AnohXjBJ9
m0kHonZxWF4YCRq2gHkiR7JGS7VpCvgncir+2QsRQI/CqHg5eNTGWreQHrAgKOIFejU6v5V/dBG5
LTeSeNvTUq9MYYYPXoeZyRX3eNcDmZm7xcHplM6l0DPGby2QQpqRq9slhpy760lb48b/woPnEUcn
4Q8qM5Bm73rrCAwvop6NsmMorgU4ahgDHWLwL668IMCOoTjnsqYsNjxWpY5/WJy554CtJMGX30dz
DcJGts6yR1cXcNCAKty01olyUFLdU0jjxAgARYlN4y6lGz8KvAFTRom0lsp7TyMfa3oHtvTU1wBp
YH+CvyqkiHYrTJuaHVIbNzjwMsLjshDH0b6KjjfMFibEU0k2dQtkOV1BQclKZwrkkIIe8FxajuWE
+EJSBR2SMa5wglm3cM32RYewQtFMUElDNwoBWr760sR+qTE+lP9dVF12W57qLf+ErPE887ZcNYQK
ktpXasw7ZSSLEFt5v60Z/MeoPpL29EXgVLOiwSzdgrzr6DTKYK1HydDs4+j1KyQ/jLKFVt3wt7xm
Pvm06itfthSL/RBe1je1Per5Nqpez4y9f4ICKEgCRpz75jBi0ZsMn1eYB5M5DWkeDKwbHRG91Nou
b2w4zrUytToCrR6IAzoqzvRJjWtumAx02feg56hSEg4yle9kar9oC90rah6SgsK/iWR8eKLzXt3I
Gd/kY3kYF5Kqh1yVTxON9gT4ZwuYjuVBIVRqvEHrWAcH3w/qpFGo2G+nSXtAkDPvwdDUvPKsSb2I
LSTTjgvjaqEI3CjzM3agYG53pmc5AhjmU8YABnn9UwzuFzMFYehTivp28dZxHQgv+hG3r7lcUY5v
+Cr3iSAhr56k4vLOYqT6UnNdqzJrsy8b9PJTc8vcLHN59gNHxV3xhNRRoVuMHa406rAZ+SqCeOpl
SWRELa6lLR3PNdL6fWbjvCO7MhtXlkgr8mcVhjC7UIY/g36mNHINWMDRxoLtlqZfwh0Cuhq1UYBU
2L8ZPs9N0Nn+GCu81eQQ9yxcJlsifV26yhzQXx1HEuii2obYK22a/JpVl/RqNbJ9jCCLV+7SSAdf
JsL/vn2AWqcRbk7Y1h/isWK8F+5A41kBJ3W0GuFqhyeItOeEs2wqCSh5xYFGUQbJ1GhyC913FBhR
4Rc1LkbxnrsL77zAStoC/OOFQuVHpg4KI8OdxEtEHcZePERj0RUp6nGCT6fFfrNkW1kSsFF73fS2
sUGpR7PnnTUhxQ0CtbJ6CyQT2RbYAt9/e3OkfOQ89I14A2LTAY6bj0RvAygAdXfI2FtKljz7Jn93
ptJbfWwHMV5OIVeM2O6csTA2xaYvCbeh5nZJ5lDuOeLtqwWad8IfT6+FmvfMf/24cfgLUyfeeRSr
sjuSDbclUOIzNlmQHkII0M7iNr2GMe+Uy45jLqVBQg2dlZc6WVhX0OuG0YVxPcqTVy2itmSv8otG
HmuupzKxGofpJkHC8yS8COXSB8H8yrS0XXJoBux/e2E1NtW9GnC/nYHKuK5ykAkoZOV2SsATuQ5W
rYTa211z8cfyVtb8DflRhn0MswStxfpElFZdhIvb18cyuMDVXT5MRDaCVCJIT1PwchXu2tylGx5I
jnGMTgtTA+S27E3AmiUow8znTqapqCD/KYuE72BtagZiaje+0IybYpnxgq5CKS1IDEXfp+iQlSze
qf3omwi3uJEME1VVO89xiprrgDHQYnaQXbAbn1hG9hjnmK1CV3A9zUIjA2ZwuLWVPkaNlYakmmrM
fISrG5KWfdKDrZq1ZeVp2LhtCkWXDvILmB69GO1NdozJU+0sBXU3WpLU3MLobOy3ktuaIp7BwpGf
K5o9WNqw8fcJxlDDBGE1IWoEDJOvVcGwphj6yNMW1ul0APZNjPLeZcYMNbhAH5L5NO7IH3saw9RH
OKPNrlTBht49e+37vk5sPpRrfh/0/4W+qj08HnwTGkXAlC6GYMUmCm2rXOCRcRyl6sOuECE6r2kS
9+bBbS1XoAS525/pgiwvrCzPZQmMIHO+S7fFZ24I/DmPtS5KsmczuUvwqBV5yNN2CnrdpHqDH3lO
myWs6Tgtk8GrGjYeKryfxB4yaTZ31Ea0U5EHboc+mwGvLfa9js/taq2aNDKBDSnnS8AUn+os6gA/
KgfaxC70DUwEUvbCmqiToGKKygBb3igklgQfSzSnKeQvf1JSFNft41e1nk8g+2VVb3uqmpz05v21
XfoAd7HGfVvPWBCHmRdxBluKwiIeMJf0JEaT01LloiC0R7StAk6Eg5YNRD+I6WB+cYUICczH4nUj
6FmXEoxHW5iIrcPcXKfcI9NgD66SHj88QuNnFFmyl+mxW5lWvWXyhnwNC6Uqy63t48AHU3u2NExL
nvNh1Nt509Gzg2hkzh7GVG7zInm5V8dBwQOTO4lIHya0Bz/Q7YpeZqBdRtB8u7gTB715RuHum7yU
JhWLe9gTYt7E6yEuIKdw7BHbQF1GuBn7V/WMqoKl4ca8ZMYY3Wz039gKxqpqgxKWEMfPFjCE/XwY
APaufzb4x5eB2q9/GPMiRW+2+ZZ9ahN8wLx5jQFoFdXrVfWEqmLAZg2wYd7abSRmXJCwKjcQxdxb
kQ/12lUV9lW2NSdybfkFRIYvgcLOiCW2eAoqFQR5xBR+SJNbydAOk0K5jzpA2p1ZUHXFCZRGdTYH
hffLUyH1XV4MucsUJVjt41lyTFE9zX/U7qaKNuI9L/Ismzb/RigO38bAZIBVzFBBIrIu6Gy1YIua
XuHArHfk+FvQo9yTn1LdcBOyeJI+gKlJyriDeZ45tJZgeZ6MqNEmYP88qlQoxh9/AaLoH3dRpPKN
cDDLxMSmFKDYyYVnUtBEUwaFM1NtWocGhRDuBZvM0cl+RS8bexyGvMS6JjquIXUd39thqrD5DOdM
Wrt3QG1owJUjoOqu4sGCc9AD9PhXb+Jjf9g4LbfQkF98HaBOu02+ES6FrXRcn27xGB9zCExKyJ3Q
zHmdblZ/ZsVj2Bewi5n5DiOBzVB5tXX6mdCMXHR/9GvbZHn6gBm1goY42YGvHgEsHYyz20BPlq87
kZ6s5Woo/2ssG/b+Usb5Js4SSLckKl8l4aq2HjQVOmpPZuILAnef/PNWIjSMDwRgENNu49SlXErB
swuMS/kD5yC2YbCZdPVt3GUP9+h7+vjd/Ih00uJgbjFL/9+f9qeXW+IqXZQ5ndZgpQBqBykOyfGl
gqoHxbLJxsvlmxOZMi/1Li48PD/cLCmYVarAW1PUgGShEKNG/hJ1+Zvz52/+MFKv14y5X7ZdyX5/
ZRKihSGH+za00T5K9P64An7qkBG5qObqZ5dqLsfhCrhLcGoYY07Sb7tFw58zYknf/s9fOBJ0qGk4
QKczW3uHAfiuJ5ozWAYVM9n3PLyXIreIt1HjLQbD4WJJ8BYKD1M05smyzVnbzMGCTuzgo1Zb5sp6
oP6dFc+tBspraI1pqSLldcK7OiqPBKvd0nJvJKMDLOWT7PPGkiqDRDHqqyJGc2FfIdvFhnTon029
GUDaun34kUf50KYUVAJVE7wyWc5a/cOdWY2NJaoiAIxmU1cOrp4qkU4P94tRC8Pd90fRcQDYSdOx
6F0lBS/yKsU8IhV6PG02HuGw/r+vjl7VTqOnGqkoarT9pi/KAwqwBBs8DIIRITBY5Tg0QHI+5Ac1
oWkY18M1BUbpN/raKUaiIc7z6vpum2evgu0wKVF9o9Ll1Taqin0IwcUwWmtv1bCkoXMuLUJNlbl1
x6mpNHmQO7ZxgFTbEwrh7CSYHbxe18cnnFUX89wySQhPghp4e3qHWqmiZrObTqKxyLHeBR/JGD87
UJJFjXq+W/NgltB8zQXJs45svWFOdiL1lrvQjnaHwDB7gt2+YX1aAxAjCnV5Uf/roMTRvJSbHaIn
FJKawZPmlgBKsY5e0ke8DtoPTxVHIjChelSlLIhYJJOB1vuLMcxoR2rOAtqK3DeI1IEkhQAr+LHa
XAUcYMeqfuB9Ob65jK4il4loHVCFDcHdCAbRYX/x8c63v4zDgD2tqMXyj6cnu8IMqJART7vCue+R
HGM96fivLImFmcjTI9YGAVn68lowhJztD0vPdA7kZx2lYzNqFlrEfL5H4HPCXXPbjS+O6DM4jJmh
NKTLFoBesBuwd3JDT3U/9Q0SBFEPWOqZe7FIvMGv6d7DnTuS+97xMx2NwC/zL/hrLqCZyK3XASit
D+ulW4HPYD5GyZI8RYf7uVd8R+MvZ/E2wUvzjcOChLR+M9WRt2NxC8zG2bq4uxZIczaSk08as9AN
Wrfy8q8Z4AcNZXhAUpzoFUk9wfE0YLDspjp+0tHqcxDqSDttmA80VnRxzUAIph380KaXW7SHPjO+
k04abNhMay98Rg+qM0Xmk6r76/Xb3+qHVltTZisbH3xaZkfMpvx4pQLs/GsvRiHL9Ye4u1oMiXng
WP/2JtyjYbeH0GnetZnCGm2vTnVLNYDzmMZjBhoHA134Q9Q+N/1HfyXuXdlYmhwerimRf6EgTEfA
LPXoJpf6j/+/nzz2tmXHMbxxVjgsckrRhp34QSYw8J6bqvvtMG/JpBM0tLXq5QROykWM2n0T6gdL
KaSzOj6xb/oE4GVOYQAJuKN4GcUF7K4NyVTiShW6woaTxbG4gx6mSb1dYKkCchcyBIub7A9zUYdm
/YUSotFTno1w/muIOWdmr/D3UPBnwD6L+fcJGtz/25DKYTW78uuZlTXtV+KYMSrE69HuKva9tNlw
RaXuDzQZWVBb8jY4gZR7x942koGO5206xoXoORXb4i2MTfT47oNGmURMqMkeI2HrOtebC/U7FQXE
Z6w6lZYK1lBjPZeHHuyfgQ3fDU26nDfGTrhBPH9vrT5+5Y/EdfwpoRwMGvwEWP6Aq+8roh+3AROh
vuckwhu3mITMfp58pIUvFhzlkzqwx5zYbBzPzA9H8Z6UwRoaVBBvhGG8rBC+GUZe3Cu9UXO8RxV9
yxggxNoFmMO8xNZ6GPl/v+AesIj6GUBltX+VfABt5nGfVeSMNJLFng1uPTOpDm9SwWjtaMsDzjqp
/BPpvETwQ8dqPoKaiFpQZ868Y74aAbJRT0Hfo4G1gDBIwLefNshXwy8X03b8A7E7yY4S2yJa+Klt
fFcAO3bSEOqOrQiGBa0IgodkiwrhxdoZZxu5k35SyZLCybzC+EBMUy53VGDlFfb6u0QWTo/XvQnX
RkovWQsgFbheKWQuUcwi149Vl9jQtpopbtfFkZxlT6yJ7U0AgHKCFiCEBLYLO84ZfRVE1s5BiOTw
JSqpUU+70g5XfwhvpS/TIHWX4ZmARR6TmIvYIeMLVQaQ/IU3M2/p6JJYUP0l9QqzA5JTDS1HXBVG
GZmBC8aVsDJdss1hF2pUhrKvsiHUpVK5BEcR4w6UsrG2+fj//VxDV+RUiN1xX2QZpKLjFlTRR23A
93c0h6DE6YI9RMqp8mcMyXB4M1Wh33DazbYplCayS2ywLdLpiIAcJ+jFr6TGlBCqeKZzX55geLEa
ljAPbatpy9FVHEkzPMAyaGnwIjaaK9zMOVFEU2Yx+5hM0rSrTngCy0WBMNeY/pDGYRuGRXP9CzK6
tS/U4NpktsRJCbspllEzDX5750XGZWbIpWbdMl6I5+15igFpTl55Flsc+NQ2I4vRIwsfF23oQTcy
YU5PdiJ/U4tXzF2G3rHctdXmDpjJgR6Ghca/z3S/U6kQloUxjN36qANJdWl2lFZZc1KGv2cSycxD
5q1MsD4OMGL0Gbk8FvcFe1vX9T0KuBE2n8E1UfTUNS0IQOZexyflAJv5AXuxlb2PwqaGGp2zTNXe
IU0H5sswEWKguZnabXJvhPbxet1WtXDO1SZoLc4QPX3+DNTJF0xiIus1kivJEkt0ELzI0BIDxcjS
adyKQPSfds1qHYIIDCG/7jas1/WhFxY06XkgHQpZLRXhcMgZQvO1gM8R+bswosdiweJoJdtb+bqP
F/EbiTtiC/Q+WrdKy6uSucwbCUmu7MIVid/pdnZbScFdVBSwMXbttRNLk/tKkHrg9otKGL81gtdE
BtoK6cGq0Vwm36t0lgutqv7qI9sPoHggtWuvRBQbGJnP1jnCc2PR/UYkavLxlCaSKR9khnc7FiWV
ianDxzSaJ/BvMAeuntJEFm2bw6SPZNrJ5g6LXRtQON5+Iu9iGZZtPO//xFJs7OTI2/9v4MsHnLBa
LP6pnvQeTFutOs24f6jc+U6ipPEvElR75btkZ0Qwlt0yUsWsscjZb6fktv7GofopA6cOIUEL7NI3
rU0Jz4jqF2UdVpee30kJBJ4nwQztg6lhegIYwyqOSp3qmf4yaFrB9/ah2pygg0S6gjlxaL65gN4d
pvgHnRV1PAU4H9SqHcrq5MGHGs7J9WiO6t9wAHO0nWr5R9km6CH7KP6h+j+0hxgtdT/1IaP394rp
BwETxFEXgdNdj1j2pp5b3zaZPe47egbrcBtLDBHHXS0DvC1zGlXtGY98/IQhdKa2CJknI/OqP1ea
jxhnaByjNmtTLoUaS969J69K4vBOjYf+Ow+chlNkqexPXWlfoDCPrzVpXYlBxsmONIocsJkPuGmf
2Y5ds4ZRVueP3zuwX5Ey9pvA6lDn73eMkwigCeCunEAwM1xYv0rjiBBNBc6W6bEx86KNQc0gnSHB
93410uSDmfz3OXsc1/idwqydw4NkS/Wsvhqu1TzK6B5VLD9TOzLd96X8CzT+1PyaKyrtzZ1mhA/n
enmBSF205ja+DKt4ff2ebtsd04RvRqgnvCzKvF+mxmvseNtQgsytSszPKImJcR4XGWMFATV2wGRx
1e/KNBNm/vxNY7PwaTWyHhyUgW/QqVULU8/9ADSwZjIZ4eZtUgGYVfMDmRxmhqe8k7+scj0r/Ppe
q69kRq6khi+rLAkM/Y/Wt7A7Wh+PdfAFQp9KuJ5679/47mqQgBrtgpAz4kHkEL2d6a9TxjwWYSq2
XHy0OroHH+LZ4byz+034rMqL3EzhIy2KR9Kdx/qtPS3DiYhTgQgW3pHIUIlUUYo+p8CByecrIfTQ
d5122Sm/VbCA2rkBEsAMbh7tR46wVdtV9khTh/k/nm3cJ2oiGeo3K0b2vtXoiAiUT7hCR9uDBhU7
LzmHSPYm9ZwyEKFTj3ZwwVRqPfXBaJIg6oOfgvyjfIDKVoelEMBsiP2eof0WwQAPjjlBhv3n/YgX
l8tdpiI38vZvxMcZdBiEk6p07nRJOa+qyNqwafV4a7wRRNa+f+3w//2SKez4ehJtOQzHULwOwu17
pj5RYWByGSkR+rCYl+ivMLQxquWx0g1mZmaiewnmX6v7gMmJCxvX2C3D7jRn8t2JcKNFoVjZSc88
qsanMAzxg5omzmvHJrB5bf4pJx0j5vD0DOcHzKba4KXfwyIybKy0/q6pwvXUUbSMHvMTrOq5338H
feTunW8ALmqGV0rPHhNkzyTrckVXL7pzT0UdbXtwcBjsljbIpprWSXUxODoivWBqWHmWScpQ36A4
/FlHv5vD/K66fDhvYrka8d7YlKJNjsLVt0BFy6NJ3guILUsNXYpDiP8hyOMRZGR6HqMrC4jVqRJU
uT+reCsBXqghog4gb+TTH1WwddBsI2xdAGrDN/0loQ76Ic0kGem3vWBav/XY7n3XmUtldLmaC9Gq
qKz9TcHtRDD8rjEjS9LrzyRufBCMrEiFR20pJcAjpI+A+H+hyASdAGHo2g/+4mgnzk4FrlA9NhMv
WdOh3XLVLkFbBiBL57EgqfHfKLwnsV7Ftup4m5uVpshKyp7OTLc6iZOPTQ28RYpuXSKJ9ps+Ydkr
oVfhCwtJuRZvcYp88d8WGMuWE9EXojaCePuXxT0I3HsRq/daXe/xP6uRjLlE7zRFsLC657Pq8guC
rDQ2YmW1cOxbWYNkckas0w5CMGZC0UhepO+IOpjW8QkS1Q1Vtjv+KcJdiauBeyS+2bQemIHrSpAw
W/FoqHt7CQ5UL7R4QU177cqFKLIZUiV5KlvF2MNCKeaEy601njy+dohieY+NTfEuV0FsKJpCFOMO
BdBZMeoFJUP6q37ObysHcw65qLOhpfS2c5+tkLPd2IAaHQ2W5eDmPC0amIy0I3gdePeVezyaaDd6
sQ/AqtJZlIF/JF6wGhMrH0qXExkXuIl6k9GUKXGEXtueT7+539teMkdG9uqHPb33ZR/lIBCTTban
Q/CzsM/pzJohq24mOzgW4YoEVpDW1o9YN+DraiwXbQng2/MEfNDygGQDU5jQExRbLthHBZ17QuPY
cqtd2EzEN1UESlmQvFPnsHhGn2kpulPP/ctKyTty3cog8LzVLEbxVa/TkQE2ffMGipYarPoGhyxk
3YYIRRhxVrBe/CZfBe1Fssmio2SGrIN3+30yi3YBRLCfjZ+H0A3CsfFcFDlgEQhmE3IGxc7tA1S7
Ik+cb53lFBjZRDJJjhXPyQ1ohjKlfwKKyVaqnrTrUk9NmxQz+4ctPjjgN09QPB77w3Nf2cJhXPxg
4Nq3hqX/0kGHy/4mk56IY+qWZWLUG1kyTYoz7bWmEYfEOpSn818wp8HCsfi2w3ekRHTljvwTRhMn
RTehiJFd+U2DFUe0ha9CMLUEfL/pdT9HgjbM1MXVXp9aZtBwm3JtY4PmiC+fnlUBhe0XRQg139Rn
2BmMZXI8s/iPiG6Zjhyhmui6quVbu5B/U5EwHDFS+G+BuhTEJ9b+0EkhZZXYEMRIQaVBXmJwh7VU
n8xkMjcO4ymqHwetCvyKvS3kF11S9vkB68YsJcRqoktEXX2uck/60m82NerJT6PEWNyL9qvt79Rm
uwKk1h1W82v95iP5HTynfNN+xkrVh7q/cT9Ehohqs1611i5GISURqxf7xEX8/HgqQ1c38Pf+2aDM
7Q4leks3ROc9mgu3RBABq3mrqQHo1ausGW9ye7XAxV9A4etjUFymx3wy6EURDiSICBznrt0ZCyn8
LBGpp25fBgao3NGq4U64/5dhgjhGsrOAc+LaeKHiJ9AKHFARR+/1EjucgNfqHC8OWSv0ViH15sXO
whWYMrfU0woxb2Lo7oXyBO7cywWHQ5WmAcwwtlVJVjrgpTRJpGICKdLF4rljE+PJQ/mzAnyfdHCI
lEihPyrhgm5Kk0L50gw+KneEAhGrQm7/BI+NKCmxhLdG1mlSZLJusLbaXJO5q1WYXRl+i8F95HlN
F0we5IHNrF9PZS/ywwJ4p1HCfVgvjJfK+kuq8Jttg4aAQ8TcGxLSXwmpxJiB66cn4fmWXT0QOxCM
fMhR4f9eXUeBa8km2h3vD3hOucgo4ulFLPa4c56DgXkfoEzQr43FJ1R+Tq7QsuNxXiUFsRpMfhP7
KS1PyeNngoZdaO9CrYUFEYts4Pgq6MFrgekBz5+1P5CJ4x0Z17QCsTsp0itOqsZKFS12pnvlagfP
6UcnocTrclcXa2xr+uEUFlA5tWdv5E9k3sh2pUGgaX3CDOamppObeGbXmRGnvAyRn2Pmw+4OLdbR
O60lgkcqv6F2j3D+6oYvKVK4RSSnKPKgCdjwv+UMPfRCN08nGquuHvGqjZDuX5w/WmlSWI9Z+I4C
8HUa5Qi8TTbOGu69xHAzUSIaqxCXi2tJe3lKFelzP1o2FBjYpiyJwA+uuBoorxWqgNPStgEzuzt4
3NMetLJJc1hKQxUaW1Xev9B6KNVcpoys/fWdJQFFAQHR8PpaSHHAXXLXcNoDvsMO9DTW5F4bPKBy
LaQ0iWSkqa1J+b3TN3mTVbJ9SDFjbF1EPK8LjfmNh/YXFDP8r7T60R22mJCNtP6prtC6zi8cj358
umIUgMVwSEqmnjAuH1b4yKBCTL7wLig1qRWNH3ukv+9sUzHYDjYWaLB8URVOtO4t0tnAX2rsR057
NuKbjAgfqm735RUu+08RkvrtXNniegwC8wKoPVhR6t074xWr4dWMGWJKKtWqlgEIsweeXuSO6cP3
CHtCSbcTsnxwgrw04nZ8fDUZL+1/15D5avsC5DeFRMS/v+jzqEkOaMgEhwafMGE4tiXjCftUboE1
vo8g7oV9bZB4f35phpr38Mo6bh+Y2ihVoEVr92DHcxL7yrUv8IXYoC7MtVL7YdmZpoURcQ2WT8I8
cHHFunWWc0kNkkJXC7jOTQUyf+7zn8d45W8AXOgWbscUsM5e6Na2PBx9AnAR76VLif+yvR0oKBMy
R8XexWR0n9ml+5POXaGmzjzPn2XOE80JUVvTPVZfN5S2jupdgO16lrZvPI/orHevsuxpyzg+hIKE
S+tqaFIcYjAPNHOcWz/nstMY0n+VBrg/kNGB+tkl2btSRNfKYefLBRDIvB6y6f1SaCKImiKhFPC7
/kOzYaGzPlFvei7c2dWJgn3lm4bu+usUO28IOr+XtL64XgjpjQWwNxxMewgvWSYBFoK8SAvcz3vc
Gw5TjeHx4TwGjL6H6d/b7LakhDrrrqeVxQk34YDeVc/wc/G9fmzUMq2ShRd29DZjefILv4mBAtZ1
VuACPm0iu24m6K/I1YTQa6STM5fKzcUpX75IsHguJ/ekYq7xtvo7ToEf9RZLmpnj9YF4siLx1Q58
YywBd0mnnmMB9nt6ihWKYzO5rteIiNWkx45ZYaXCng2mElTSPqtXcUUsUYEyfpIO4PQjdJR+Rl6X
wn+a/ShJ9XYthx2WYa8L+/f8JvvkVo615T+xDnBjEHDDOpBtz29BJUiJkopCDO/EKGlSlN32TTKc
NM2wEPgM2rK9DBr2Yen3Omam2ka39C429KtqYAy8K05HBvA96jDfL9sqh/TK99e9bB955NUP8QLw
qLVVEya6Xok9+R9iF7a6EHi9WHVlNvcqry+kBZuhEyCn0smuKeiy0E0FA5V1BpJRDRthJsLoRA7I
oJrZzPJ0S43dh1JRkliwhwRkWCXyssWFyO0zyXvPbWcTemWbLARafAilVKVV8uWoHm9AAqVx7REG
RWu7xTce/lms55K6FJAau8y9Hk/GApD+V+K8dqHkXWu8FRgCwwjLijmJaPyfCW2pv3n9isErX2Hc
7pVYz2S3xJnb2uyaDlsBlz0xHs7vMU7OHDUcwS2FA7oJCnlufHA5sUgqTJpnsOvN7QxftVYHbwEL
5wA5WU7+kFcbrAYbcazGqqrafemFSZfTVcA/Kk5dnCxsZYf3YQZsu70FxC6D1/K4iZyJX83EZaWK
we1wRdktCryT64oiTFwx94hb9XY1IExthB+0ZJga8T4obCv9SFSe1a5teoqRN4IblONpbRpU1r/o
vztSpnLnq1Us3CjafBbFfTjqEYDUA5CTz+N4csCYYLMkn6AUMourZy8KoaHr9CvMwSza4DeKeSBD
J5u8s3BcpiFylGN+Beq0FriURFSNndmKkRyagXMHcs/YGAWarFDFgiMNPiCCpa1ypTP0xiRi+GUo
M9YpuAPgdjaV9FyqnHEaCP0C0co9yCUAX2qKXdujWiW46YQfU73eUWjNxMwVtE7pk4KfgRDONhGk
3VMk3EYR+SctRxg2DOnQdM0+DuKcagCiTTPlhWSv789wY80LWz3SktS2eWlBIz6l28dkVmEcFTsZ
BoC0+AeqH6rN0vR9Fq5YYtflfnN3zOgtAsQSU6e+7ikUCqtYTIqQMZLyCYlx4ZyMgj69KxOGKf+C
ap9+NRndFDMvxslQMG/k0cTyU8yGLHibPlBHhEzE0AZVZWHO7i+LbHWhaYyM67pnE29v/JrndbMq
43Y0k+Am82xY5neRDsEKHhLusotpVJZ8MJdm3U3Y6f4NKib0gEBY2+q98/QMq/X73MrkCkN8M1V1
V0iyCQOk3J2pGv8wKFlOPBDt+ebellsZL5eIeVKft3V+oxMxgWkQpziVRw8PnRYtcwicIFiXYNYS
3JRCpgS14cFzQWjCuAtqdXbgNhhNTLoCrZ2xVz2bGlM/MWk5rHJsX0QaXqBfRaPUbFRQsVB40sFr
DQvfGY3Zjnh0HkkqV1YZsoDDnB172OgaNu4zeERRZkIxFfjKXa078HwK1jCYOMJsJvOa4C6jfEZv
kxqEtoyeiOzk2DIWK99/89hVB6sUbGfH2lP98U0KA8wp/7GzoL7LgQRVxjMSmjl43GdIQRFrK4Ia
HOAN/PRdd4scNxqgRv/q4a9vGsjw5KDX8XOk/e+DUQ0rHR7hPx7PVlIAVRoepzq05bnL+U7oANhD
V7CDS5Ad2oW4uNBRFDe/+WRjtPyjOnzliajAT6oqvSZb8cd/pN/QJ9Gmo56rbCW1QMFfFxIE4Kir
eQw3PhF9HiO0802m3gIXiB3dYiWupyr8P1REwEnbsrUbZvc3hPNN3SI04+1lx8wcH147uqIvARcE
OuxcXlSL26Uf5rJ0P7JtvpFyY09CdKn2fZkNBCUCqDjcp42N6cTDJDNznvzbNVB6iW3yIGfy5A8r
bYnQ8e8SLH2tyGGF8KuHt7xfCtyQxKrb1MqbzLoaoelCK/P3rc3vkAbgtzV0DUe01I1BJryDN+aC
YMRHDKogshLUTTBaFyKwIWbO5GoAtzdO2V2kAQasmQ7e0Y3Av2OgX8SfbL10fqLVIfrHDrvKPhpY
eRZf8dWjndLlZpz63z5n7609ZM7/O55CxqfV/IcbFtmnsKlSvuPPzJYGB/1MDvIFjcJky7I5ch+F
dqeYpzHcU6suYZKOVnFvyuRFzjnLiXsPwjfq4E7OaLtq8gvoM8fdmRacqxTQWHLfyvJC1mlEi5uY
HcoBXSOxkzAVHPwAtAEo6JnNqB57iFb4tMoOsOwMQ5b+jD07BSzeiwpCE4+nVDtppa+IaOEevmQt
QGL08OoeJq2RM3MwNTK2FM3cQQuCKmBoRsBBbFqydi0BncTEy4cOlFXdDIuy3yaZFFcApFFUESjJ
sIK0re06sE5RaV1K86fjqa96L3T6kHv/lQercfUnNFGQoe/VgQzYvmra1UnD5aC0sCuwqkGEmwM6
pAxm8AYK2SnnMH+h1Mr9Wgu0Axfjc3xW+lDukndoJQ4aRhtYDUe6UYGfjBvR2rlzCBWUgaBAuFE3
OCMSl0fgs+VNDPSMVk6JDWFOTGtItFv1dDZVDuf8lan1X6V8hqnX5+KnQ2iIqvZglQpirUVYg2EG
0OMQu1VaEcCt4GsSozKI/NF/5sqKEZsBRqTvRjZIw8GTvLQLyuD8+2gqZ9kOwyuC0OFDnd6b2cic
6XSNKPC7Rkt8+riGFOnqO/tlQLqr2dwUSj0ZFfSEKaynwDio6RxAZtJgL4gCOU5GiyCfzJdV7MZy
Fk3j1CUUtMud/z0leiCNUFOFqJhDPFVZsDp07ZSTb/pJouqdLFMJ+uBumOSJdrlbM7ubVvuKGCDM
Y+i4EtsDPdGn0RqrAyVvgxlO29kGU1f9eFQBNm81zlFt5DWtAqPuSckqpKTXBiJkEmScS5ga2nJ/
/GzuwRS3gb2Rsr5F7cs3k+/xwnJ5KhUXTV7DpchBmjp+4K2R29UrmbH6PykDAqA6AaLMoRC/RRNA
EGJmiDAVIzUGWsSUph0HGOX7OF4qnM3KuALMwm/a6UE07DHj/HuiCmO3+eG0eEW7pprBh0Bm4vyg
VRCsKwOtUCZ/TpOusb4NOSwUNx8lXsA9X4rbbU5FHg/kZiZQE39Xq16UYEfg4FpjqBdCD5b0IGGU
m06uB2YPssoApBa250o5ZQimD0ve7xNGjMef0Bzv3R+ptjMOyuPOplUq39SX90oCllf8euwatxv/
myaqGt4Bx+uH/0du+iQ8Xx4mTdM+A0zRCGpbNyNvqxUF0TLndbOR9EaUxufacxGqpfz70U1nbB8m
ix1lbD0IWV0m3SsVCt1giey7aL9O5XAat5vpVVcRMcCEtB6Q/tEFtc5GR8ZPOHGZmT3AUHcqcSrK
9swcZ82MdTNCiDjSP98STIgRx59c8J4G4x+tpGqJuDSvlZvOM1ld9Z8imCNfaENzE8aPoMzg9Tor
le7jw3Ot+9GLbcGQqHHr0nPyBGLY+LVaaPNH82Qw92dGPlkipNP05Yx3Nh5XzKHdoC5tm1ExuGQT
GH/+AyT7IJ2s2Qo/Iu7G/oK/x7wIhDYLByO65JfYcEQ9AmXz5/xQWwQ0mffqPtsZFd4/VJTYTQqc
ReQ7VTY+4guPsekmJyPH21n3jCFc1fe0RX80LEL3b/j4yo70vqb7yFAjcEH1IWcK6OnY/TZDVLRT
00yX3xXKn0taD674WTUjWrs0U0EPZUhW9qDhhMd7qOctUn7Pz0FswXrxWelLpwIFeqxRklyXMqGW
ZkmaUY6CRlrzEbzK05DbuR0BeEYVOzzQvS6exO2pZejQO3DFTge4HbAJQPVBmKZ0KjR5Vt3Jn6h9
VsI8PZb5K1U4ICoqrOtQ+49fTUjZ9/907uv1oszLeI5Rdp6fDOgqmqXFptOAOtq+GkBLnQqU4s1r
k6rU1U42McJtZ/W83HYkyIbJBI5j+KIT0M9Tjok4wN6UctQKK9sQGEFCTH10zP7Hp72bzWwhcpGM
Se1azBBQhN5jw9F21tNo4ED7Nckd6B7enlA6dJ+kpAWDkZ3tHfmyGRfX5UWXZ/IC8FcZTWQbLt3n
zYxreDs4G0i2kuzgVJ3Uajm3jNOrFGFTwtMDZxRPYGmnNgrjxBGlrb7JHLBg15u8Cn8Zzv2Dcwjh
pFS0yTdQkAXd3yrXpyn77csvNVhr0J8FCPcRT3zQA1rNmPBx+yt+B3iY3wSkRXP4vYaa6HbuxDlL
dv6RlMknSsNRRi+77Lce2BiuXAhfHlzj+YeZyCdLjdZUSaGQC/aW+Xk2zbiruxKH+R9xcARc8c2C
Ag3jBUKfCRRblxspUxLRj3SuaNuS9rIg5HgOMnSaeArhOuNR/d9o2tIFOqsPrKY/FFfJ89lPb4gg
Mv/8fXXsNtvaMRztzSR1zHrsWgKmgpNsgcKmvw367VSZsX1Wzq4graaUwVcL/hf2GafeMQCx619a
nCd4f45nZexqiMNC70CJnt1K9ygBX4QnfZgcj1bx1Q2HQJyVuantwk3tg7TkOPnnsYdYD2CUUqKQ
bIDBl1zzDs9oAyHCB4zMWkKoC5yDPBxFxnJAWcph9MGdo0/znwojqlonvubY3vrd7XucAQy2Mt4b
zKLo05aLgNtGxkCgCLgTaas9rn5WV3swg+qkOak3WFM4s66OCiAFS4LliPWL1d+DAk4EMQye/fv7
qyzrDjQuTAYWu/LQUrJUd0Pk2oTCrdUx+z0TqH6rqdzi9yFu2IaIraC7JeA9NDSr1n2GQYz41Cli
t1xnGJoxFsvUWjl+2n6EZey8IzMi59Nsj0GHfbt0b5XrRYjq7MYe9bgQCJRWcLk5w/jMIzZcnSeR
CUYYGmEhlCQr+whBxnXzFOE1RmytHPRbANfdrtzqbXuvmULm5pjM+tPPJquW9Y+Y4T/7zaK5VpVk
7BQ28yUyvMcCGTV4sh/t04R0qpZR99OfC7TY/wU3lds3m384DWZ+TxKfYPsNeJlxogLLSKpKFJiW
hqvCAQvf/9f7fdG03S9rmkBt1JT1ZmnluTxJ+K6j+nKoYjiQOzAF2vYL44HCrk0vh4nMsXPtbnWe
gv5MgUvnAiz4J6Q27AmVtcP1Udw0kc3MMCnVMdIpaAX7oCxHUtJIfrrIGcRRZN+oYy2MbxkTbaX2
AvOXrmVr6mRpF55QlTBf0+JWEN2GWinszsckzR6a6E51qWfX2ClAE2DUILUXTdLX136EiPNoh1/N
2GTfxGGu5IEy/9njCju3Em6pMJWP17LJ8j3nUwJ54EDy95hnGC++Setl/fGIiWuGxc94qCSD8lh6
1SGibic2MileG3Vmuv0AuY3j4azn0ixHhwETETmG5IL8IalEKU3mkx+8gS/f6jsUdidm+hvVNtzH
FV3eeqYS0n+lbu3UiFw8Yqpl1KdjHychhD8+aCSNh7SvCI6wTV5yHXQkbFYqxmUZaWxNqanMw1wm
Zs4CVOaSbGA8NJoxZYIq5YS1L74IrDNbCIHArg0GnBfCEl+VKLTOJKJz+tKCMEtQVeE1FqXTgG3I
Me5M8lvoOr9wTcEpwKrXU+byw85giklm8YfsFdIZ4KEPBvMkaHUswqAAPUQCZux06aw0dpDNy5Qn
cmnmIqhFyUZ6lqV9Gt+6VyaQrUQ2At3r1B510medQhanY75G7pkB+Vwj+kdS1kl/kfHaBDSHaN7w
9+2OrZJ/ddpHY6hwDV5baTBfKC8LOx1SzKPhI20Xv5nLOe38+0DhnqQud+JOlFF1TV8NE/icQ+lm
oGVQWo9ui7fcv3GdLYsc1ST88aVd2FZGuD7+/TTRbl/31PTjh3fs4v/f61GCANesv/ezOadLhFub
5m3PQFPhKMI2R1gWg2FzMs3s7lNkM30X4HERAuCVfj39dZJ3Se0RpvJ3DTGoGiA8i6wDVYSh0HY9
Z9r1GoLr7T9ZyrheHVcCE+1dtD3f7+z3Df3rnbSv7I8RDFM5/nIcBG9Ycv/2B6owZckra2xXKXYD
A9+A3NowbyXI4NqF1ReyT5TQgx0u2pudYcY/KnLW+uopzHKfnnEtE4kV6oGqf7CJvavlRovyX4WQ
wzVacdbFGLqo9jB+uOKEbtk1QkmtF3JcLc6nnDJSNNTisEtLfcMEmXz8Pq23X7V8+yeoVf5pm5my
+DIcSQwmiLdLLTjXrxDKya1D5gF5lZhc7+KfO48rv/oOHXg5roFFdBg3Ap0xne3C62x7otu3n/H+
VDDA72WTEaNmHFPy0PH6ikeVVlY2m17i34j9jUTU++6qvyqnzFw4oPOUI5xQ6s6dnEwALufeQtZ5
CGl9ivlCeSfSFBjfkDBVmGaNG0zSE1I5tTz/CVj9oTbPEzE5mYGgRpLM/fmd9XeN2npiIHaKzTm7
IcVdlTbTnXsmo5Z49cLjvj2wzDf7Fe2Xy+8Q8SNAAZgDjvR6EJWIDR/NcvQLGQ3mwNDrvnDvjJQ8
E8a6yYNq5NruNV33S8tyQ23NBphESliIILTqt+3OOy3JqGs7uWEuqXEfK1cTNjiAIgsLgm5JlFDF
TdZ9E73IzAdK5FYf6uQ/vqpQd0L4VosqmRHF+gxXm8M3V1x1XGKdRBCU1pSoAvY7XLl77z3bhIY+
7+ZHAcZetgJtbDG4PQwsOOAJpfJEQxVUUabAf6eNQXl116JLnnPuLZVS0loXTZHMSMuNeUqBCikx
dD2o0dNO45/FElsdOaZemTy74mc+A9YAPwzjoyDrp8MocgIh5jiKV68XD8oQH3FWmWBVteEd+vJu
3+o9B2RanyEn2mb6mVCnOPzTJ7Aw5hFJHcG1QljwUoZx+ehH2i+d1351ACuosDIcr2QgPqtcwQoL
1Hi/tRaG/3a4RS0+mtzbf/+siaeWpJKqVN9N2XnUm+waqGqWnhDerRz4d+b5Xby32Euj9qc5hHt7
w1kiQl3fm2TjbhQVMBY6DNsZejrcV7ULFHYw1EfxfscF6LExME3BE7lopNZ9xdOdKI8fbSoqYTLT
6yiMV9OTMpLStRoax+LcqENlGChp5VdCRp3DpOy+0l6uuv2VUS9LL55Z2xTHguhNCTy3Pfca+XfA
T5WFzctnZlaK6/905kPnbMJRAnTUxaFrd+SuKWHZOygA+JNzzuUhhwIeqfeYv9JfZ2eqC5l2/J0M
GGpqJeNGMC7HUVRa+YYTeh4lgyvoyBQcjL+ELNBlyn/DkAfdLrMI9bDOS6VTQNQ+AtycbFGhsFzF
gJCanYq+5t2bLuNAPzR/BEhMINvAxAiDew7pxjbGCH+f1EHfhQaMFXNQR43QcMgMVS01yHSKZ7Tm
f625pNOx0skJSkZQFiIeFb0PSZUuLbR2utTFfWhlnwPSv2NBZ7WB4eAMqDVpcIp9O/MGg2aHk3jK
Nl4yrm2mye/UmPtf7QdE9LCqYvGmAFn1B1hdGPocOteASp4pEm5A7yeFqS0lDGg6SxAck9d9ITcE
54hdZMl6/9hrBRXBKdwszCbWmn81oIgD5G7o5JrzefloivqYQTzo61skKqUnh90fL7P+oPz2nLlt
U0LXyp4c7HEoeiYKGjUK2ad0hYr8TLpxN+dFnse6xKN+AzZfMVFsBSARKST4biCAfuXfzUG/9VHm
jXno0h1s1dVJt6/mS3kvXN4zWWtvmsGzIgtatMXad5VnAni2rNIM+tKaWJwqGwF+Y53i5cv/QMF9
O+6hGJz8dwRISC2Mnxb59qjcPUso0m/n9mqn5N2tWK7vbkKvLq9z428FLujPmYpF2KXC0UjyoA4A
gYtnLAFpbI7hFGhRn5dxBXjEyOEzPxUJErzpc4/bDZ32Xg0hL4uW4vV8XjkCJ+2edPbHPZU1cmB0
QQx4ngM5j9HlPpi5+H/nNYjmzAEmr3mTxAp3XySwLrsf6DTrezj+krdxUOlWNG6F32V02DFvv4C3
gTcnPh+R6fb9tYCno3ztZmmNxJK42RVjdrWtOWh/dR5wc7G61J5x7a3RwW5GLmhDixbiBbvNyEam
+J4MqvAPfRy7uItqLciJ2YyonvBiMVs0bgmwXYADTocUS5nooUj5zAVprdYnz6tYB9clytcFi/zU
14+GibOOd0PoabQLyD1QuF3NzyI1vILbtjJDZzH5iPq8NPCrhPXtv/N7XaPsqbc7bV2sbJsb5Dfd
F79rYQrJNIsV7ynH+bYRFzAScRDBBVfcnvPqYUhHFss/1yiIN2XidJc0jfFXVmeY8Mb5l5aZ29i9
zWK73UtH4HHSY1si0y7siGutDi2ZXo/5gaa1/xNwmFGWmBTGD4axzPcixXt7mRJIP7BC/1cygEt8
J/y3dDvu8iUQ15xWr3lCh59fJZK5CEe1k5yDMryIGSXf8uZqBl5X0IEN2k+hlMDK7VLJqLym0Yvo
n3nRHDNUECtiN0nO0jsoLDn4mclenXQMtEWCxtCd8QLIjNz1QER0KNCnDixRDeV16PL1SSuRhRJa
SL7FmE7Odf7FHx1/wyCH3LAaGdUIdGQONmpKL0Z2HnGmCi0j9/sMaeR3J1xUX7rY3kZRia+40rkT
znMvK4qsPCadYFF2SJOsDLA3LK7pvogZMoyo3PeTEM7J+c029uq2xG1jHzlqyeZ00gbTgEAZlm73
820QGorXphvcwHD0T/5AXmSIk9Pf2FMUI7J9SpitRvn8NPgyalyuyBHGNLCzt5AZz9gEtv9tibg3
JIoWai3fMZq2MAwaBPTnEmAF3nhb5HYsxaRG+xsqp9ViO6CreHF3a11zWeesED13I9T/h+qCaQO7
QW+A0b/Xwhx1T3dvEB2s3tYlGSyBk8eIwLLTdnL5yNptXdZItFf6mW3vXp1ME5HSyCPUSZKeJTLn
qGUYu/t8s3kr6h0uB5jFC5GBtsU9o4JywnDfR/meqa4JtuUlImlflM/7Sy5kGg9KUcmdPxoVSGWR
QQb5D3lUKxhvBoRwloTxyLIApdWgoKEOs8SBtp8JrUqJJt8iPig62zpGmWISuUJIgxd2BwrSHgiM
d+PzXVAR9VwnMbGnL1sGKLUlMXKmvXQ0Z3+f8G7AJUeWv4Vhe3ZVwV3qnBDKbL8DzTIn1YUwjw7b
yx555Sh/Mzs19CaemV8dYOFYUn9pozaVN6rxdf3Rru/+sunkufyA/iZEy9iaZM8AnTK7iVXH/qg8
Lhpie/Az1Bg9FKOZPjI6zdcmSoEvOoCsgct/tfLnAKqxTZ6yXUXumXTWpayZ3udOqaRj55F/2qG4
AONWRFVJDqj+FVqKHh6v8Mkc5cBaC11eNNJNiPcSqL8oO+WbLOWf2qg1kQ9eGPyyJzlaI390sf7n
cl2ZZuzDT+UHX85iTTe3m0hXB8SEKVZ9wFzNsrCYjjCA3v80040eX+eA6gjkdVUkR4VEcabHW90s
/Ac1OGWsUG15lBCBhPWnEvDX2mlgcl2ox52rEjwlUf+MWi3CqBN7Hjp+utGivCvM/CPepnlkpPR2
7caVW8QTP/D0ExNuc+oJNl2guhSbcRsriq1ejJaJFCtY5YW1yroXjR0xkGpZ6Q+DR0+qMqIQOSje
pshqfgiNdPE8hmLDTnIIvqHSkMPUFJidfd//dbVi1uMmDk97samhrBO8A9IMiucOHzQH2VyYh4GN
S+JNf859d9LOamD7kC2urV9JsF8DfYeYy8BqSoH3oD2e/zDPEGx/s7hgVFzoYODEPvApjICPAnBD
i7z0i/6MpEySWHuleuQp0oztjwxk5bScJYg6xZcG6r2XvtUWT1x+ORfRSFpwPAESX+hhVXCHkME5
rQI0PaODmauO0i51K2ACCpsKcppnxwMpIpabVn0kYLsfpSX9bxt3g1pneJcpzYRUy8SFb0CWMI7l
lgae3Qi98w8NyS4exuWKQRmYutVteKk0fFEp1cj4iJPEjXU3TFjJSmt8oyjnXiFC5Xi5ZZF5MUmF
u23tnJYvH32v4D8rOyKC52C8j8D8Q7Sk6VBETsI88Goc5Ch4B9WS5x5sdlev19v4Pds1sO+5Y19Y
YBqDjXOK7NVXAz8v0XwpGufkkVOCXyQe8+6WTnAW+eGosLqm12iVeZc49Y9mIx+vlZISP0bARmJO
GpK3jxnxsGDRS//oI9rYNDRlyuQbqjR51O6pW+eD5EhPmTKuiFoGiIzinsVt76CcxhZVPxgeKOHs
0aNA8IaZyRV0JzEL7jcDsItMh7uGyl1SRJbAhe+Wp3+nPh2bnpukUm3P+1PKHolyVTTrkx1a+6N5
SfviI2FQm9F3vrMmt80uslWTm8wDWclOGkifzYVrEvkCY85N0LqYmpKtxEFb28cWFaBAvXr+1GFB
XYUCDSS5Cy1Hbt53gI7s0qpOH6BAV+clYoyNh8sYR9n6gVae1sjKGxrobTZ7gmOjgHQkQHxRsm4T
oqTgVCiqi8YvWktYFTkX2mBp3hONR5JapGSor3+wFVEgQ6xRNIL+SvD0zaU0u/12o8zsJyqk5aV3
MhvGP4JT/+sjFgdxJEKq9tkZa6Dl+q8kJdqMSt4fumoyWnpuxZeOkgBV39PlQ9sAGAi/UH8rAqLn
54CKS3yrsfMw/Hiye1HHlFmylJOZVeBKAfAKPKOGw2Vq9AiPfXAEmSjwTCXdpUsBzQzc7EOB1ASE
Vpelnxo+GVG7xfSjbYjEqt9s2eBML5TluPTJUFzn7ArF8ncXD9zTi4/BplhLcF7kIPli4JHOMSUp
W/t9JJZBl6dWHLPNkAIZ44fvtENTFF2W8ittkNAY8ktykQCXiPLnIuPvy/F+ABNW5534xmG2lUE7
q+30dDKQhS/+h+mFAd3z6CtY1xY1sncXXNAsEItZLGmItXa1aV6y8T8cApG8iUXvMvY8lOcjSnx9
hz6L7Cqg2pOJZ+17wwohkMBVjYcm97o+yR6RuhHCEuBuxmvXzneUJd9tDW4Kfvq1p56LglBVBI+O
PTgnajN4T77CZyO/wBFNgFb94zoeamZvEtqI3Q+ElugEEu2tiA0OmzjZsZsTs+VG4/rGF/b2A9GL
hNgHaBUkNF1yGYXxyLRaAfzjaRYQd22fzN/iB9e1tLKfNd50ANwcTQgBzk1yw/QvU/d5coO36zd0
TRDayiFvcJ+aLSkVIYNUxINRXrrNyPDmi4p+u/jfHOkwAtAR2PYom4wBsYVWZYN/De5P1t8sz9vv
EXoPDrVh9CxEoRmAIZ6H1SG9Tkq97223cdXecdaWLxh37P4/v/Rw+Ga9CzXwLegZ4vjitleKGoPW
CFnyO5FT8y9385n8ad6LJWuwT9zEL5H4fvVGPuVkjhRWUX+B3wEa8bBDNBuRy5FRdX9qYI+loU7O
s75WGGD4hCMgNRLLT961pv2QjE6WqucADVP9ZDiAOpGYvnPM4UUcEjO1VpaeCEhqiGFplpVfatCp
BToi8BBhYtdBwx3QAlstm6fO5kSmPdNX1PuOnxu6xSD3MOsKQPN039Y5LEcn507s67sZI/G1i8H7
qMDmyeQ7W2V3aeAelFGO/d8bsmGiPyVH5NX4Jw0EqHC+KEMWF9oMaVoZ65ZuCe1m6bjPhiowRnam
mOBJ7Wug6sFdDPVYKS5zro4acWzQOzopsgI6FR+96fXI1hEfqB9H/evoL38SsunAOGHLcSIpMc5E
jg8x/gxQm65dwtznj4nfiRLRB6PfCdJ+MWzznPOiGkdpkdqhivrOPCT3XzLeneg3Ex0gcNKMk2jD
UPxBtzM9n8SA+9JhaHlIz3Y6VQvRraf/ug+WS7iw6wNak8O5PBr00SidGvrfal4nEBa3/bYo3YB5
OiPYfjS6Es/ysBWbfUExxqJUxEp8mcV9K7HtOF6gzRpMtdUyLo+R901+ueey0MCJbByq0TihivVF
6tBC/zOP7YksYJzgQCS8UA9NIMduwx8dHy19DRG8OsoGWZqb4U7hBtSkBaBTt0yrNv0H0KgBH31A
YhWWZvQ3tY7rvBgYXNHYNoIuu7GGwYAXFHPBx5h4GicH/NCfW0NDu+N/mdpg05XviqGTbaVo6INh
nfSSfEuinNOkHKKi5qNe+tY/UUooTY2iORyXXi0CTb4BRk+I7tzB+wN0BsZu7KMhDoM/Hb/u4uXp
Qtm3oUD3VQUAM/wxn4tdxW0Z7xCakovltEzPW14ujO2813Vh0CvQfepnHS+ZFm0K7m22Qkmfe2Fh
ZBu/OJIYNWX1Q3XNfzLI0Ze1b2L4+SHTu8V+G79RV6e49alx2iFWYnUA0MC4SMhcNvWHR1Vgo8a8
tp8cJz+bYSRA7JOc0M6+D8QM+5kfwxZ/mD3FPH6oNxnjOuWqjFZxAM356RfTb+xOfOEb5GR8D2Ad
T8HtF955ULDWHo3myiuUJ+0yMfcT7PketYfec6MpWydJpIPLI8Mv9C4W72rAOSlJDbULPGEa1KMk
F7ldioJH7iO4VeXVRwVCkBVPm4k+dIeTCr+boJkRFjs3o+jSXXMKfr8XoKCplO+2w2AXWEEB2ONa
N1RVHNOgkQxqgfKdpzY9nrlbSWYAJSmqZHVLSYA5bnMtHIOpztRPyPUwpBTVcTdJVhpxBrzyamkW
ee9pnQ8lMZCNRxl6pw0zWWIIbGNeaWdnOr6aiUL8J7UfrwWk9GyxpvZ9ZwL9P571xo1la2rqfUS7
xXJ+4/bDgD9H/ID/Zi0lPT9QGfPDqZIswp5kMopE7wA/oPa2+7Ut1BuPxZWbt4iZtMT4QNBpzsgK
LbQ9wN6Jv2v8bvUnLv7dvN+WlEAaYdC4o1mEIywc8MeyDe+5BH4LzJJmVNSzaLvQPS97r64HhaAm
P+Ob3Du2VIihVlKhZrb1/W/SBn0FtwGAmWV1y2wW9jltYNmD4KcjVaMxee1wDxuOhpnt3JcYutcd
rZ6ISwj7rlQsfzcP5V5+i2tZQAMkKH1YLoIO9TWKlxlvXppC5n2bIMjL1U2n+0dfojIfhjl/uBNY
z3gi0vXROQA8UL/xg8tBzcPh4ZTa35NAZK9pjexociTU+Bas/T7JoAFuoRjaFCUpC9SsAh6CMSVS
KhZjeShR1vgSaWi0bC23OXoFwvaXKgXMFkZSIVWNG0Xb9AKCTk7SlOUmHfDqvfHOCRPLItaCBKUh
kjhG/GYUBdfukPBjUX+Phtf3xA8UOqnfIH+ve6vKZLzvaWteekCTgQFPBcuNTcZH4KPl1o5WSk97
1K1ttwkdmlO5oeGD7davwCBWpxb2/XD1A0Z1il1ladviBGZYaWYOirxYz3/8T9o+sI6p/+gDczrY
KPkB994yl/2rJPKsnmjm3hsSeu4D7ixPiClsrgmqLZdCqzELy6SPT9iKKhOZQoADVQC2ijTSb8xD
p1b5jV16w5IZUPsy8KqiKDjXIpUEHcpD/UF77lCnAe7kQhEde6SVek4dGFP0XWb902SuvjD0sjBY
njgFnx8sJ9UOQyjW6l01etIFK7KvwXg2jA4AGar3ql4+TCoepusDtvQBP/yy9p63zfmvT3tPX2el
7OwN2ojst7IKN+Jz4N7gpcPhR19yv3mxxyzxeL8/W3JTqZat/wLKBGoQKfry/wYLPUM3gAWgUQOn
duk8UISo5QOXqFL7orhOVFP1k3SbeDKult2t+DZnwTv9EtMx8SJr9I9PAAQDZvlDtRQCvdfRz3XN
Z8PDQsSh+O5DAlRl80mQhMe5FXlBivRYpFoEvzUlSN1pVaU9EUfGZIzUyZe08Cq+0zXTZyDdPt3s
SEHQYyEychZ5EPapAay0g/JQvI4+1btAYuKUahunc5tvK0iQ7U42URhOCrDpyWyIW5RYOegZ4MaI
ChkjWJYMMzHBAeIyMN38bCeWwvlNL5nZYK9x7eyYbzM2ALE61Wo27AkRsFMJPLziqTr31yLb0kmG
T2FcRHabwSOOTJ61xQeqbFKIfTNn3wBrseS9LQN91QkN47sZjSmm/VHPydiTGtli89v4AXnk65N1
c9LijSWQQyH4geWwsJvODleQ0frG+VchDX4UUriewnu6xziZXPq7ORRT9IvNgpPIcZ0DjqfXcpGI
gk62gBjzmgJcYpVFna+culScIv6ViRH3dMyxFEp5YFOd3BQ3eHkJYDp8GHvvQzlLPda7OuGmnc3L
ztjtidirz2ErzADAgucJpMGyBYIndmQIlH0kZmOeZs8nY8KItGVr80t8pUNa+uE8zrQD9Robx47i
JhMNtn4dlcH4hWbXBOdAMbgYUVvaL5c0QmrGnQ/QX9MBrMcPeAZdQgymXs86+nKaJfLV5Oi8TuYi
fgKD58C6GITt+o539bf+kkTgu7/Z82IgEm+i3vkgwkNgylEEu6pflpPkYiGuaKRzl7FIh6z8BUa1
N4R6jdv8lPBiYM2chqiLwphlFu3o9198S9qSVfXKg/MoA41vHj0z7CIpc+KmRb6kigZSwcwvOjIm
lxe3uP6LW0jPk1tIVo9pyAhwbr9j8rIpA/voqjvFi3006OOFFA4v00gqdc7Zz9bRZHh0C+Yk2/o3
pubLAD5CKorDhSzD0lhZ1E8vxmeRc28YrCeTeAUUugxioOF/A9pvWMsHOIKygu0/D8flpcuhWGyg
k8kruVdCL+poV6QSfWs5dY5OLZj7c9TvOxsLObbivu9h9UufvEUd+901wZSEEKQJGeYWIbwYYj6s
pqB+QDs3AU0TH5iICs9ue522e0Gj6zZdhKv6ASSGeAHdZcNV2qZZKcijDHiPay7Y8cSwbmxKMyXy
Ykxl+rmlgvfNORyGJgQzhu7dqJNLwihXXvVpPvaBjihM0pZ3MfU57NujQXi2vZefCWGBD+y9flWH
FSKS6WGui7KE0RVoGmGYpsrnd06r0HD+dfRPybcHBG1C+/ATK+GtrR4Hnx3hzd7/SF++8Ixs3GKY
t5miIiUyfn6OoHLJ8pbZAxdjs/b3COBWFYr8hMRevbJiNxSTJuUse2Igj0iGeF1CdOBxkC6pu6tU
FYo5duxldFfRU1N0xJ/5zs/GLIJk2IsSYCp2Cp2Nk+jSbTpi8xr8R19WbC7Hg0S1G1u4RaR0fAb6
AHgrHwub+zq2NajQ7inOyXyLmPNe0wDX+Ye/ho7x7VOgEkrDsArIxfYPd8JkpR43GLfY3pjVdR4+
zmCkY6AF3R+1ysLKF6uyOo2W+3vyM+0QBoqYScTTz/I0/17zkd7x/D+rwzjOHMEFu+rTjuaxXF+B
iTl8X4Z3of9WuLMbMdXbThfnyWrUaSiPxPrY+tTo/9Og7KnwprGg1G9hZm9/vIJRwg0nEon1WHzr
ODqF64Bnm/e59rYsUlHQzLhJLbmo5zIGQPpCeHcRNeo0UyXisNtcJvbb4/3/g9Ex/DlpuZjXjlCy
qHI5Sge1+WYV2h80eNmr4kxmIvALA/RJYlJF6QHEvU52hUbFcMrWcv0f7p03jlH3QrWr73cF5e4a
jHiGc9EIvDUg9+vtOcCV5YS6E2Zf0wfmcF75wlY1PgUee51AmTAmeGPgQ1QEQtLz1UOUlpsvF4JZ
vH2PNK9vFb/UZLfjbly5HHPTv1hCerSGlxTZptSLOxxbx8Em9ZoQ2fDkXWXyDcXjyl5iJM82pE/4
gBNUhoZ2Lf+CIcmhw1u1XBuelWqS9yzJKO+8aHT8ZnaYxAP45oH6IZ85f4hen/fn1ct6fu0oq93z
PSQdlipt6SMjeVYfM9p9OlGWJ8Th9ZLQ/qfOdClHBuCvX2XKQBjO2FYTG/Ucpi2Cp+qcwZgCzOuf
N2lEkShbwSc5o5/zHVq/U3ddiyTbiBccOMcze/NaLW8ltlJOqONKGkxByRcVyvMiUtDAEvu/lIgX
Plf+X6xvG5prKvzTutSnTgLBR5Nymuhdcs0MlTgwVvP52rtS9Rb6QshcloKVzNt4JwNt1K0Plbxx
/ALRFWk0R4DHkfoVrH/VqiUm1IU/sYMFk+UDQGghB1Ny4/NLqF7BSgg/cchhctgJBfN668t+te5x
Kr7rI+ph6XlNCT6c7QSkhWq9Vt3Gyn0XzBLqrtnJxEe8lIK7H4jdEBMZxyG/OHeFnla7QZe+okUZ
cf+zhRXVJPYwzJxuPpCiKouBc2WDj2JD1s3MQoxecbOd9dmqXDa9r/SZFLkWGJyhDtNioW8f3T+L
CzUFRDQLLHoc4ocBeOyWjtEnOflBJvVZ5F3DxOz+t4e3yW5mF8QU+C/MN96dJZtLYK6V7YmH+ezA
QN8yk9IrJFsN+n/wZcF1o310tMtmeESQyHV4hdmxlhOa0lET1JUSagfDF0+hbh/27vzEdb5VrAtL
ON1IxhdIRpHSTSxXkqLAR7bjqg6xPE5Y8HoY/3UewGIwJJGqgxtLt6jB1IPTmiet6BGjMPIzWBSf
KDDdhuHj0KRMRedRTgtgV7UBcpArU0AaQlFe4L81Y+EmfVPva/s8AWM3XfsB1bZK5AuaiNesh0aN
dNPENXZ3X++6wddcS76K3OkBvgpwd0uICIHsxJ+eiEMLt45YdNdBI1s0AIQXBMi+322eNWyAGw0A
T3FM65YGEqOqT7NVf1WJFGMdRCshiNw+TbHo60q+RzDlAE0K7HFTqrJtk9mOnw+LekgXdePRUsgW
t/ziDjG3nfC15os1x1UU+G7NVryBAEMTSKBBxhwF1vKbv9S/PiVLY0swYi+ftHE/5T4GqjUccBib
tJUUAEwvuBNb9lIYXWQBsaBWN83lR9Oy8hD8wonz0u68qa7fp1nbhWacklf4e0ZeaxPR4RRzxTs3
WedHcnwmnzgYB/LoyTy/sPVzKCv5fd7JjLfE0GGHZ9ZLLk4DrKKswN8A1PSveuxSMBCMYSqxjdJr
HrGv2pmevgi5SnAgjTJ0p2sbH3rSERG+yU9h1c0fNhSki1w23V6qevrWSF7AqMjBZYI6JQylWNyg
SWRjH3BSQDVGkhBT3i+86R050IBYgTTGzwjzs7sImef7mEWkQwhXeF8uzzMJIs3KszTf3nGrUMmW
aBYicHv+VJKvOCklLKR1kmM0cD6FkbMsvQkMc37/6I7tecVJEFcya/Pw8yMx4w5XSCLgU1lFLDcG
vDmLyaZ1S8H9CaX4Wbv4K3ra20trIaZ1H/3F7xadN6QZ55PPqHQWisCdjdi3GklGwPsUJxB99gB/
vHpAGhxGUyGiYnV4Y+SlK62GTcwbcBaEfPmNxoyU6Pt1m6tLs++glbwVt5gN3q1mSwOuQgvaQhPh
UxIV/4okNvDan4pDIUta3jS+As3phi+uV9cEbt0gQSpWEUTKGpv+chtpG4NZz5gk3XSfKT8yo33W
qzv3Fe4OqSGvNIUfWdpzgcFXPOkWUMj3VWzGvLN1F4zd6MSlaIoihBtLrfNnLlAgnPYKjPceFtJf
VYSiC53D4IkqIPmLljWW7Bd5KoLI1eKgvhyFUEtF6rMfNIwHI0WTVD4qZYPoydxIZPx2hzhbA9Ft
yk88DV1y2wbCvCxssNYRjDbNDuBWcvCe+7oTaMJ41ZVQwm/Yllyp0vT2udR0sM2HkgOIj8E6aklm
4CHurhh5nq1dV2Ea1H2D8Bvhg3tW/8EN+/PoBmWy27cs+8QeRRSKrkaP7cOF6WmqCE7Z/WW65atj
4BDsPqQAwNYYtvnr7C/IzJgn30a4caRkcF2KAwQOrZEA7SXFBRRT2D4Fmk0DGK62GKmZh3P+0Agu
Qq32uGwcZ3sKkQ1iVSOe8kujLk+9dLguvA0zgg47qYfaBA7FTrsAVccsRGkCZ3pL8uy/6QPTvEVB
mU253+43QEqtDyTkbxa4VPkqKTT2k/+iiFlBVsv2fCInchNQdxr/Zg6uTdWss/4nl7SsaZT9NVWQ
kFONhaoUbcyTKG1lOdnwQnGPlddVdpznxWPs/g8sRk81dyG44uN5i9n/Plg6qzjlR1y7L4txF1Zn
ulgHWkreQs3jPqpjwtWYA9SftFbE3+umJX0bKKGrkv8o+Co+inudBfojOrJnHRA+Go9bjiecXWGY
/k6hiHvucRG4Q0AlXcfmAgm/erNZVkN291Zs/wR63HJPp1NWoBC7VazKhTdnCUGxpjfGlhvRiykx
OV/5J4cQu4ScqJJuwrCW7NGlDlQjxLFaDVb06f83IhVjtUTO9h9p6QDG3Yz3MbajyjxCGtk6AzZY
MHVKfTVZPp4L5hOY4I/6sKorPh132hHMw/G+7nDiApTsoyssA6GSV+TEl85chjkBXCn9LhvS3guS
o3YAcF8y4370izZtJb+QDO7pIIqsKf0KxMD6H6Fo4cOLLKd8176y1iBeWwpmCrkz6hobxKrO3zzf
vMq9WPywHOYfsLx9Nmr7dPqgBqoztxNLCU7W7gqUNVgPUU1Dp5UxYi/UJtUxCGUjd2hglDG5gobk
vDumcxNiHCKwnxXV3VM6v5frUwJj4uDROIWK2veAzI+mAQdG+cwVTmVPdUBK0E0CdB4B2QjUEexP
DeCqrTheL85Du2lKeqTXQXnff9QPC6HbaAB+FNm84eKRrfyvFddLbZpCbD4X/72fZyjMlj3KByPo
mDWQXpLBaHqZQfNAE3h3XaXxqiiRVRuFjwCPaBG/eZN8+EF/nIzurMuLBVxYlcNpiqLyQtVr5C8a
f7frLaBmFSiq7CXIjaCctNVS3VW5aDDCvdSmxiTYhI6lylvoDoSj8U2wMgjzXW+YeSIGqMmkkgMq
24o1wWxlZuWgKFSo41X+KATuJMoWHagwkO6mP8dR7769pXn/GKL9OKkms2/+ih6HyKWxrTqYb1F3
9jjAXXJ8n5mXL8yJv+KNiAseXVyOyRRybmU4ZOifAfV9B6ya7jshe4gzWaTDTxUppD4Z5ezf1X00
OopCNaJRcyMLPCFPorNis3gB+fgr5KZQLa5mvCzLMlGf3qcrksiJVCqQh42U49fYj8ONeiodv5Gh
kEvr2wvUK73T3sjMobY4zmc8aZu6aWjg87EBXTrOScY2R1iCLLcZt4SMZhjrYU166G9mK/MgsMZD
SInVNrVZhI6A42sL59O2txXc59wy4Zki/pbCVLxLJM1QV7cdoU1PwFOM2inFLEQDbhefaHCqhX6v
uq1ynVi0d+H4fwdnCz6pc1ULzmq3gQWoPp0s5DQEDdGIsuMdicIM9Zr/g2nJXl6MTmYMudekOy27
p66uZHvIogqr8pl6d3jRTwmALuVaeFp6jR4bHJCblJ/IRQ5b8FAhBjpk+Yk9hMdoaYnaz+kR0R01
bJ2oy7T2rCOeHZX3ZEtQ9FbYaLoTkGQk8/Ke7N/Vrsm9aowpAvgmPL3FulBoocQFuQMU0OCa2RO9
Orp3cPfDB8gDj5NwRzwmv8LD1ogxbns9GZanRwTUiAIbzhBVpbVkenFpWL8Ly1rotxVBydXiwnBM
9U3uCBp8yABHzJmXKGgv8Dd7gTc3CKAmmYdLPu+JsDVEYU/3S0jsLiQVOEljocZI0hBNhVZlfa42
+1X04v0xJnxL+lmgcOhtKjevsRUWVrJGC6BkGNeRDHBX8mmxuhVTu/xcR3eoAs6I2fJtTmL3i25H
W1t9HKBq1K7BWzNdrn0ZHBwB1HsjQnA4sdO32siF5KbCXNoAVxnWcRD3UVhlN3ayvax1iCpIvDR2
RvR/qaHoig6GLQo9QIetz8kaFGXnZxv0gZPJAc1JplGn6m92wS2O3RduEFRUHi0bdwsp49p7AguY
OWBnd5le2coY+UC7mooVPEEtwttFYVWYa4hJ+j5Pan6CgC2CCR1F8hqDK/9TC8nGB44NqDeaZbF9
BkNRRc+oWatrzJbNk9+3+HrDoNUynlrPQYcpV2DrDoznOjTJ+/iQV4fCjErLghStVHlqUEdFZlRZ
U92C6HXqNRkyVC+RV3Yax0HLMXWgMacDpjRRhfMltOy0VIU5Hoc7Ko/C8crtFKW+nG5gpooHYTrL
UXYmW8wl2HH3rTYcTG/RCDR7tjrpByzquZN/7Z8acePPj6uRN+dSio5WWWRBAPTDEpcRd/DBFnIc
MgjrcIKZqfYnjGZZk/6fJwJqObASDwl3tErsJWm1qLEX2R50EHXhz1o1DO6hQ5W6bspqmZ1k2LKY
A8lY993Mkz6Wh70p1ADSTIm7msxd7BL594mOUs47sN1G4tui9UNeM5kNkNAAoQUkue1y9K0MJrvY
0H59cmaiSR2EcmEoswOtNhQrTer3/o6DrbVsYB5u7bl+j0j87M8Mzy6WpFvgFxiTA8+1gd0pSZ+c
L8cDZXDi/CdpqYFqvCHFcbg7NMHd067SaXCIouszTTZ7c4YUyZxDyVBHaZ0Mwrl+JRlXHF5qClv+
XQ2diMYFIMA4vEMp5EILgrAIfRuru4hD8GtwYdRLB2mne7If+aQCoe7nm6TMKXyrSHut3e+dzHDf
vx9CfJu22Iygpv26+VSUvXGxTtYFnvagyZ4PisSSSa3LS+bWA3HbUyWjik0vPZjRJ1YHon2BMyuf
6BunGsnFWw+DTxoYCeS4jh6ZDrxJ5gSALiaRa9+aefCVlcwEHqJlJ+vwlFx3pn9w9ztGIB0qLRIT
u3CWA8f5eh4SvpCW4xarU8vm/JC4KTWNAbvdRM7KXU4+NMWuAvN7v3NX15JwTw27oOqaNHkIzkFk
qq+Sq2hy5kbUzlS96RUM7KprXQI85lFczQfeBH7wkY5zlhsnCVmp2Bqxks2ZITdK+W52OjlU7mjS
mute8XaLzGf4oVhI2B1voMUt9j7C+Td7t8FceIuTXuzI5IimDXANJjNdc4rurvBVJDv6Ox2I53vG
+4NgON9KefOS/di4HGhlaptdxFOWIepDR526yzI1K0xVCgwTSZtSOn47UvvzTToKT1nJkBjVlLUz
Q9OEcUYaf57kLboeWIzB7C+zGdXwDYmXWPLcLgmI5jcP9/4KXrQiEUjCJw5bxuCpFwp89kC/+YO3
jXiU5ViMWz08BIiWoi7k6ecUrKJWyPalIFUjBRX7xriSgAhKX/ttRht3u3XcXEsrvdbMfOImvECc
akRHrZ4kgX323RO/odME975AS9Ejv1F9lIJuLsSLx/xW4q/VXzG8u+G2aO8Rysa2LF0Z/uf8hgdW
yALpwiIu73rLRr4HUOGVuH+biAU0en/oPBwcmJGQgRPWTtqvOnGc9S1KMRV8TcP3ZZ7s6o1MUFgm
cvJHiYpvox4RmQiFLmj9QL0MMO1/xjclRsaj57WO4CMSURfVHyHsdSsg3fnWkQgazA4G2vty/xHC
pSN+TXWn3DQWxexdiCIRw43kw3oOKsFQLetxNe6yl3DqvuTxN+pbP6DH1i8KSBZb4ADbfsWw8y/x
ndlSCxg5sLkPMDMz3kbQSiUrBJZnUe5mUSOIvXfkxWHibBGsnDSM+S8HRadB9TzFigsirQpk6zdV
9ahTzV0ZCjnHCYQl9izchJvt7cuHBgKOA3gJSDb2Z6JRfMUrnew/5oSv0Lf4gdCMLCVtlVCqgMDm
mSkDqhyoyjp18N9WmNSOcWxjhT5wYi+pS4C+vVkV1a1Y+K9cYzd0YDzeVHxFXXJoATjbyWrDDiTE
dUK2v5y3DkCWaX0/SwxrhMfyu2eUqYT49Ur6j1FJW0yVm97GkC5bUK4n5MJLGLiHRrAeFHOJcoed
11W4UAAwC3ARPevN7beTZnh6l2mQUp/D+3xePBO3WhF0aqhUKTkvVrIYTAafGLDFyUU6uoxWWVVI
LyvXY2YM+WWTqBGjzRAM2oFnNTIYr3r5FD1ozWUGk8YD1dYHYe69FDQkh5CgMjP69RMRE/sjQQWQ
YA2qC013dE+PJa+RY2njLVaNeQ5p8Y9ZRF3pjLuy1YMttFMtcqF1Juw2pCd2yna5eKL96TjW68c0
K3ELpsLCZ1u7kM5KOMmJ78sH/4+Uh8FPd7jjh1Pdlc0XAl2R6NG1D1biiZccU1I3P6SyN7ZKM/Jv
6yRHCFDn7dVs1ELuXIeqwnEIAXUxpSS0QpU2XD+9G+wVQc0fo9WMPQzLSpOzwVR8xYEyvsoOjAr9
ZhnD9sgfGWx2mvouVtQt9ObQU5J+eaeQdwr+M0CBaZL9UCs3KC6iaEfTg2VHcy8pPPAaHZWS5rxq
pl1fFZBK83RMuOVEnMm3zGhfX14rhmOUT0OPGIGD7ReFQgti0dF2GxuxfUlVfLL1aiXLleNq47ld
6ZiYVONTtngSY5DC9QjlIdRCg1p52V2NsGpRG0a5le+bqoQ785066sM9cvQU6cJYOMq5VpdOtMxm
U4dfDfx2tD3EE8qi/lvObZB5XgeEwZlXkfAmPJtep9XvfB+HytnOiJMBlxSwtRTGCRSUcrWc+p3Z
M+fvsPFs0wwySdCymryPFj0JTqrceS85V4W34YSlmB7J6GMnTUEKpo+4HJRtdVsJGVOBXfaQ9UxR
P7hCqpWWcOmpS8aNDnecrPDfyGdzla8WIqh/pCtClRi2FHDp2kiOq1YOa1+Dtam4nd++/KZMSiS+
4Ztt5p1qTuIDKCVaouOtmy4X4+1cUiWl97Y3FDCSVJl05ckpw0hJnbA0oKdr3L1FYSOdR9geWrCM
b8nQX2g7S3M1UE+XBmq1DTCGlJhGt3f2F3koxF4FxAUX6M8zRMvTD4kj+aoK1SLp/BkCmwcYKhok
7VxFYLOPGIQCWe6OAstYpfGYu7vj9oWy6to2QNig3Mbrw/ruydl4Y9inUfB8+VhFbQhTX0x3UWNL
75y9QQaNEFnuHtKVKtt4ptP4k2aktLKdjpKQlxBQAHTvFjzcdIFQXOZySJtBrRlXFPrRIzhuY7eG
9L2Ek+95z4EDtyFQt73rd8LcrAEXUyRdguSNJRBBQEvi1U3wub/Y4fBOnOUCLb8zkw23YYSi3Taj
C88VsEj+RAqr1HC54P9xgoMgn+hDUkEMOn6MPyD4TvM9vRmKjmaHeZZNavVKkmwPfhIXnXU/OTHk
83u84Bvw5K3qWNc1/QvJEFbpFEY5UpuaY3OGAArx4CFiJcb6brQ5wZczY/Eud5oQnqxhz6RhqEWO
vnbMQBVxoDagPHGlJ5aqtsP6MOkpq5w1TprIn16Z4Ckr7fIBquOi6EKu8MLpG+5I9POS7Ti/n8QI
T6ObxwSffHDlu0/RXHSA5TuLFEP5i4/uydAnCYIACzHt3lqaDgOLGPmTZObe1rq1YMKGJBhUw6Um
bW1LRtkW5x/1JthLqs1nsa69vlNJ5BLnYIzbn/9HXQSY7SwX6eVzdFufPUAKLGI2XX+ZWTY/fb+6
/qZgxmIvchBEb++RzAWumut1miJSMhkaripD75qjYT+clhl09JiNr/emq1I1QibbIA9MCc7c+zi8
Ho0h3ISbO9aE47c9bOR6Hht8ZtuYtLYywngYAblToelNYHHejwQ0bDJfzFP60LWcAvlqfR4RVLXB
SnJwyH0Blpdp5vk1Q2h8qr4ogc+HyHn7OIZvuWPBQvtJbcLtZxvzwSljSi1mQUe+ND2Fea9sX3Xv
dYo5X3JdwpQW2fjwPZDl4PTD/c89DXPkWoqPfZg0rSzfeBHfyXvEJuO8sjil7FzGnxyNtMWHO0r+
OJklgeSbAXx2nK41tCB9FDXulCJq8AboUOO+DyNLpS8gDUyfsYHpfygn6Oa0Mwf0WMbkixGWSTNM
L0e9vUSdVcOO25IlJELTKnzQX9n9UFbMQViJkFJlcRpjQvzYN22dLcqp7ChIbFbH2a730eD4nQ6L
P2FkzI28miDiL5c9pr/KL8uCVoBX98QVE5d+OTvea5qlxo+yl0G0ZBYQCVs9AoIryhHZrBM34EKg
X3dpXBiE+LYj9D/GzDddvkdwkMhR7H0KjInxUAgoijFkwJBq2CCREaF0Zssttd9gWCYMggzEPHX4
kuogSyWqBbsvnv01QNVtI6i5Ai78q0+2ZgOf/SADTqbRpo593vTtiwZgGqRr+NKjaNdjo+WKGxpn
m8n6JPSwpjISdUgdgQD0xhO3l9vNPXhdQ4riVs0Ds9YbLP+imxTX3f5ZjqlFu8+6tgmgM0oYNqur
TdZQ5dp0TYa4w+u3ELvVl3xRzUwwmoUyBHjXQrMGM+kEpwLqOOwKKI6QEZ+wSkPbac5fmQvpe7D+
jHFKWJn1EM56HGLtzOx/8Rkn5rh7qUjlwn1YcSuljFW2T8MpVGPrdqyXtm4sGnRP+M0OLQXerACh
MUNOzl/NA6BSMS9Q2TOoFZKMf3+csM4jZE6yEc7OfcTZbBzs4UYtNWYFNFIVb0O2qLEnZcfMXFj8
YyDihye0nEzSi96NMgyvw2cqrfx2p2N4LKTJUSlGEO1Bb7wPfe2ojk7VEt/E5m8nQjxMDtOYBl2T
ST6vgeLjJVZuCqxMcMracUxTrBpYpTWD4IjkX1djvYnlzaAh+HgPJWbaHHY1nhLo36TMdg9i3SYe
82sUM1g41yTYreEhTwbx53MZ3zxD+HX6oV8LImyY1I+2DL4VktZoZ+/6/Ai7OzV5lRz9j6Bl37+Q
oFaEq9EKzgIHcT88n0QHUpJagOk9D3oArLidvNEGRfjay404+fSp7ocBxyTg5HGhW62iCT0xKVSW
vLHsBP2GX++atN2gEX9aEMqZT1jpI6G4HjT77vuM83RxC86MJij8bIDjuMIHu7z8ejla4kks00fV
Gh0PgAffmoGdzow7CnqRbFKcr4sglcCKBq2/w3XKNm2HV8iUuBhtLPyotPTXDv6Ky43ROahUcIVv
DeQot1PpIW2RuivVnb8wWKTv2vRj5zuwExdg495JxXg5u6qkum/grJRcJKUbL1iHSRvJUjy08Dh+
39XZHLNPVNR6ewv0V/98CQihwBNzuwwMqlRErgPTsZslXKli4bq6ABlEhpBQKQwZzwyaghQRKSG1
Cz+q7JR762cTOnL8GgdsyIL0pqyR1osS8WpTjX/8SymIWGUUuANcEPDuyj3WMYy7p0pLOIsLluKd
sGqzde3p/9S+B/Ug37XDKYAvq1n4WtYtB2ojP3F5Uq8N3h66xhxnVWJCziK2kw8hk7OGSi/QoHF9
661zhVEeRkAyvqn4jIkldR8lI/UslIxQEX81EXrAVEAsjZWFNzXC1b9hMjHhSvW0zJK3qSyvZdpx
gXGzTwFG3Md5Lo58w3/z00I64TtuSsUcTylO4wrWp2x0iT/Tr37KQPaHONVsoKDmnX7pTIyWhCjt
mnZ73lz2p/7nyH47jmk0IcLU/NReb1KTkAMlDOtJkCmVpXhn9E5pC4os9VKEwPpxVmZVeQPuDsgz
PNG37PPL/ByGpD1/0a9702Q2eTKnmHWY5MDdEeG/LxpxvdriKZ/ydEOwT7wjx+qJCs4dgdQJYMgP
Njf0FdpucEkyJ6OEzbgUn0tRe5xz9Pac14JkpQ4RYTdGLw6taKyaJQGcP9f/69jlZvxvRsrc3LYq
wJohoXMCvhiHPMGYc686cD8oV4WyCHwSPdPzywkb091rcxXOEu3cOag12rP0FOSTO+Q8X2igqE36
dflDD3bjECBtAbKu2Nt58MIIVeDPi2euDuEwfWnt/T3z7qMS6T2Tf4z0PKepfO0CuW42DYuk2qo2
k8XraYUnfgDjag7JjXkew+Zm29wM746GqoJXKiStsc9aY6h9HBJfirM8vfQVlnBsjW1s2pxZpxUg
GxYrIw1YwquLSf7LpwhtZnIA0Nb0KfFAVAucUBXi6wk+nljVin6GZXtWJuRhEpHkKAfjjYmxd+yr
B+8MhQnlFPWTByfcjNXZMHp6cIB/7UpXfyQzeIcUID6IIpvGOmGIvfpvibRdI6lPyP/8JUimSnUR
oYuArCUZ7Z32jxTy8b6fN9xdKLAS9iB7xx3K3BGqm3SZ7wndVts7n9QPfP10ftTkGGWXDyzwHo/R
UIAGehwqieNHl7vDeFybkWtdJtE9u1mU9WZ8FHfQYiLKn1MaoKNky2tad/HkRet64XLT9NO88ceF
f82f9AlN4/hOTY9x3c09cApwTJRqNuIIxfmD6/oNRXuD/GV3YnViZm8lwQCkCljkFqusEmXUYhL5
0AFRR3YZBXqFFIsFwds8duY8LWHUHoyXOABI2Q29J5AvsbC/j6SqnaWKjTNGupag5fg+/JxZGV45
T1PbFjbnC+Trpm35GO8roPhl24uRHOsfnYuakvzRk01JGQVN9oIdhenChIWGHO6TYSHV+uTSMUqQ
QJAmh3u2NDUFCZeP6E0/c9/eEEOPuB8CPwrxRkk6/5kImvoWXKJewWPKaGI3DSLLIHoEwAk56ZOu
WMZbJ3CJMbQZeU3Tu34/k1tOT5XbtBixO5k/KVlOCbdI4xlzxm5shM/R/KrLVsq/8WGbPiYxY7/o
x1FBOHb8SrMFsyPxzDywsrloI/wCZExCayAX15h4S9+Jsyk3SIHuvkIqm1Hjk0j42PViRU5+PZqi
FXJQfLXH0aZzT1ziaYJhCUJBWp01uluv98VtuhVWI0bUNS3XUSs780uvCgp1AdN9kWynEfq6QLfl
oJU0/vbA1f80Es8fOtc0fFBS0y68Q4Qnj8QanYLAvBUIKcDn4Y06dsj3+sOmK/qAdX6xYWJnV66B
AEUGkCQm7U2Cc8GeoF5n3e4hVDI10VfSno1tmqiL6McfDw5d1AsTUCepFQ7/fyqossWw60QoAi8F
mGHDnqHjt0VFeGzw8SeH9d+TTrmRIbsi/T+gCTvog6NPKdgVG+1ONzzi7nizydaQN+GId/CiSsRF
aHEKd7wlQFMuc0gLGf7RxOjethQfCNeK3PNrDMryTH/ppAoUrx9fmHSQlSaJBmEn5OetWHuqqM2W
Z8mYdlT6ZOfOlN9aKnKb3oBOdkA6tuPGkqwBJxtOLLjOQibH/U7QO8CJOjHO3a39jNsRhFSxsQNA
VJPrvpPeRfP9rlQFRJkhH4DgV3tlgJHMNvuHgn9yGixA0vMjS6JJOdru53rYcdKI53OPtpSr1Gr5
bNW/V9GqpA4luv0fY3RRD0D8Jr193pLGUMf/cMSNEKZNV5nSNKQsVZvLQhgaXX0WvTEuza02s7lD
GC/LvbAQn3yVPHBfZoNB5cV4Nph5+q4r2Vg2RBsNmJgjP9PdQrd3mHeNrPlTrgFlBunGHjd7m6AK
ofW7Vx0wOtSb3YFgDaoiDJdNVRqMBN2cwsdcsoSA88gV3+6R7pr3mkVlbe3QftE4ODokr9Ga/Y8J
AZSkAtqDZYivJvf9MpxbADrYFSZSJazcfJ6litLU2TgDAoLUkaUAlEEEAbyBh5zJV3kIzPprAUh6
GCLO+sbi6/WI8cNMzvEwoHdqpCLUoTQZAq2EtMZ55LOizmz13nLhBA0qwOvB/OYzRMxOSzH/kF0B
GPYxkosVwuL/+wo4zvS4Jas66CottyIRTPDuwhiZ1TWDFtozkboW/YGqFxL2r37Ut72cK8uidACG
5ub/XKsk2mx++2mmQ4+tGQMLGEz3flRNna2R5BxgYhxMB8/PpP1mrZ0Q0odrtrniJ0TtL5gxJXR6
BdfDDfNf8G/2ToOQYxlACtZ9zJgztzlFVgXCbseg5S8pvgOWKFAHhQ/OFW1CV87LyD7HDTUzVegv
fQ52dtvvl41FIjMcK5e3TePZl6KKhq0aLJilw2B+T9jgI+KatcFrXHvRAgbvmOfWzd9zeu7r8skv
1Z0siyM8FI6w3ujZtA8r6eeMWFULLDQz6L9vdKJhWMnuinTEDCiJ14SjMExfyYpKgp3iNLudw6ZQ
f/NYA1oGIP+vdS2L92yxSDaB65TFZWoiqxtgpOoj1Xe9gRZ7i81PJ25vWai5eQiRE76W6csW+6vc
bNvAaX7OVfE4B9MnrZ2y321gwYuUUz456gV5sgjgfOOsEGwu4sJv2h17lnnkt47+h0amH/Uz2H1h
xsSbIqU6jDnx+TU6VsDieRSROOYAjbYS+JXR/qKOarFs3en5+O1FxxP6HYGHxO52A2QB/MHOXkIJ
GwocdeUSgr9eJgFmh2umw6xi6kUhMgfsL9LFqkPCN7d5Ued4DL9XBc3WBKO8TL5F/oWAl1UfwtN4
0KAIT3VNlf6lyTHmr0V4sbILdzE5BkhWd+2e6KAQvyS4mJKPIAI3dKQSZYtK4ExelEC/D51n63DK
xWiK6Sw8wtvlPWQUkn2HhyCC99ZmsdN5lTOzjXyKrLUQiwrvsDkxQUR+bef/Igkd0LASxj2l7AXm
bwNQvc8xwBinuvd+Xs9VCIKMk7mPdPyfQQaDqVO1xqv5lWEFSuqCu8qxe82FA9jntIcnoN+EaaIU
wEiYemITsce+QIGsG+nrirM6hwS61R6SZ0CoS2YPknAtp8Vu7LGLuevfKvA01r4l7cre7fr8vLhh
DVe5ItlYyMUEUTsK1Wq12q+eH7BnhnBIY/4rGUDT2NNEYeL28AT/GtUfI3CpbISoKs9fie0fzvUR
hTAtL4DjtdEqx3b70PDYVI4K1K/sYQO/9vq8FnKeN/A5tPhmT8TupSAMcuPdci9SNJgxu+N+G/Nq
Djl9WUE32wgEstnLKC81/MnMiM3YlaVsAHALp/srTq/WuCZ+KxoT/m1b2nhNjboYPt0JbVPWO14C
V025wznxGyku7wJxxTQDVu++axwzDCUyAoXL6UtMfHjplIa4bNLSNvoM3AHCTYvdyELPGYOacJeK
ahfdaKwOk855EtUI/PxmcyzmYnBYsGmMtSoAnvAcU1o3LLYnwuSDccNHTUzphkSSAT8927nGAOBK
NG6gfY3yxoaxQrJZpBDzNtDlaok3zGL5QaFgaRwhKWMWPR62oDZyTZhVWwuHH7cEwRQEUISTpIql
H9lZg49x7MgaE3V6g0gCO6zi1lfMxH1sXYHHyz3SULe1UnnB20OPSxVMzicHuwCvZaItJRDp4nyX
wz7RhEAvy81fMdbssPzi5n/d7A6KOAkpM92BwKbr2WpVN9BBaClwRBx7f8PZdsgaG8TARsyvVxA1
16wO8RZ/Cp+dXsGobGooZqQVbVBSnWeS3bJysuKaEzVtlZp+hFM+itqkRRDBNg8ctF4dBPqfOyk1
77pKBLlNeH9smY/ku7FEVhHuu+d95fveJM4n75/mXUuOT6Wg8KWtLE5QwptRPY/bNybhr53YUVbK
03/S+lT4BE3vp8648dnsSyXQYiTvbsJCQCGFaIuuerAEfYdaPnjzk1CmL2MflK8IKXE1DqKV/XO+
HF8Op/H81lDINLEl/Q8JE69mVnJ2cukapVuoxLB9rA6VS1J6CKD3s1eD4lbi/mQvT9c9Z/Ht2ang
4DnhSuXmZ0ClII3K63qnOeeJ5gJas7JSUGD783+Mtya2n8WcfG3QpFcrkLJVHgyeB6OVs3vOo745
jKxQsobb5YnD72yziSuSpYd96BtDGyw/A5ev1Pybkt/zSYU/+q9qz2YelOEdwDT5pPoz5vA6G9Hv
ZzLMEfQlF3NnPv6Zl6i57mInIOUa8WYBpxM9t2BfvDNvcLaKHXp7LmjrNEHY11x/RrgYnMN+WcSs
pbwYCl/UqUO+RgyjfjibjAUd4XnxIfqq18g71XPa+tjsYqYA8fgJa7tlu0ZRql6QrQP+y2xIoJ3w
9ziAM6Hpino8phbXuCzsjlFvvzhGRBi1gEKruGYEg1PjSmrvPJvB0R6V39myIc5ZKUwoht2ebgWV
DQvsEX85x63SY3XNA1buDRDIXyXGB1HjylVET3lh6mNE1W5cIT5FLlTJy+6UwfWAt0SeP4DDAVJC
xQSZVDamxE2gfKJbRCu9Y6m1PGzPdpkrrdx06+NWPsyjSq6ScJ+BQla6oXaO03PzF20LOOXU3GLc
Ew3DTvHHjAdUiRqm3+qEIY/7oe+HdoTbKPAWTxbb5PMsX+Fo8pyl1KW8lrrMmLf0YuoZ9+sKbSKy
5hPCl/hPFHZdtz7XbCscBmeKFbQBcSTsMA8Xr8Ars+/Wirc64WHMATG9bE3yPrT7CMM8B7HbP7mZ
EdcYExXH3RUQ68zlGAklxrWInrpfWeLOXj09dv/NIc4QArtHJMu5EFaY152TlrtCz5QHBTxRzt59
OgA/F8fYsz7fnx5gcCvSAev5oeuWGcHs3GxtOnaDZirwa5xwu40yPwj5eU9/C2NIKjO4WWv/Gee7
dUs1TnVKwldmvOqMef/dgAOfkzKxkbN8EnmPrk+sOcPDA6F0EWeUlrJ0PGgujgt/l7BpCR6ri+60
W1VZsX4sRUCqaWEaiF9OpEIQFfk4vQStCwxpruDuuuSthA2zhoCb69waQHHLYfyQ7wYOhYbmvhcP
E0vcbzdqLPQe5q3R1/4s9BJOiCd60AL+dZZ9GMNf54LJXELylFd6HDCWCSE+4iwK2zpiymHeJo3m
+4O+Xj5JxPjxAt/12A0eXVqc6FVx61sH0+m0tS18v3re62S7T4ZMKbjJd0BQwPEwB6rBxahHwlMk
7i3P/xqC6jdA2D3EDYUvib2MenwQTKnY6Kdqxp6qm0v6Y0eZ76wbwQn+GK+kvscDENXCUaRJekkS
n+XP1uZ3j2i5IDlQiERVL/KMpv5QzHrvo3WH6mrkH7On+GQ/5xyPZut5m6lAgy3S+ocaV7zp1ERG
k33bq0ZPMjK14y15QIGT7j27e+wKgKiJCiBHEDPHWcqnUC2r2sxYuhs6JNy61OOXJf3THoKd070q
kU38Ib3Cnvx070XSX64N94WP7Th8SMndSWBqF07nuN6iboyu/7OyaTowa4NJKetEbXnSaqdcnl0r
zAbiAqkcyQ3Pisexux9eAUjAeQCIACt5MNy/vx4S5Byt7Xz9sbJxGjC/EeoKoDgpXEnjE0JvU1HA
QZEz5O5VK0FLGsKu8aDGWdUqHZDukp9jVLP1BPcxC8MhrcmunbXzRAcM2bVu+Lzf0LLE9WdJIJzl
HRitJjcbE7+3zN9iRdwArSW99QORP5mo1PrVAbQ2RYN+sLtwyNqpVkIYRzNT+f2gV3g+bvirHznl
mBmAhFBf6AGUGoLNKYJ1mSOEAQPK3lGZkPlnbWhPE1ln9s3Q329FSxfWP+YLj8eVtNmYBiH+PGmi
4fg/6YREpHFuctblB4ZmXu88lGmFzZL1iGZGQzqgF7/gfz3FTv26qj7CmWxfUQ1Uic/OzkPfAtrR
+RqVc97BRvesZ6X3jW/f8HFwqiD0qBIZDU1PHFnIrLsrjlp7q3hzzLdwq5DSv2tDh8CY4FryudBq
lXwniyRf2Gsc7Pzj8D50m3xiEPUxYk6EfjHM71LN8rssknmeUs40Bzkf7MrOcNJ9s+6zlt7UDYJI
PiBKvq2C4pOWuzVmR3ogHcZQp/V1e4Su7tTbtu+BCyaRtyMGrI9/YAiGoowC21o8qve7422tLo6R
sf+3JVcxVfoi5e0ba7shTxPkckBaYeamYTlxT8YQPbhTaTz9WeDbNxTgHaW1pvIP42dO02oSO6EU
loclHTuCA2m4g59u34qx4SfSyqQyWY/EeUvv90Llx4ErY8sxJTdUHSdu7alMU1NK1q15FsHNLarM
0KltrkZVhomwWGN1aMlrlsaq4KpRerC2rsrRVzhY3gECaabnYHKY9o2yeE4hPSmVTmwjSeHoHYI1
jcSoOrGqzQemMEG9Roa40l5C5/f9OBhqm0SSpjN8zPnV8UFyImT1hir8SJAtj3B2C5wov1HIZ/+I
7yLZIa6JB+wqgM5Ouw1YtwIpQ4XOYMi3Vor4LPSS+2DKmjtxzUnruKDMS3FXpSGyKo6K5XACp+5U
in+44Ie2GPqjhP3VjaiB6q/rK2A8MkWdaAWx7hjiJO5APaTQNXmr3hW93n/DN79z29hXVrK/sMSA
qtcpBULpcrpwMiHeHpefmXrbLEOtdZT3xRlZlu3pK9tOlWO0MWVktBw/a6OHLBM1le/bFVPsdQ8A
dOmFnc2jL/uJECdNiw3qQygqV1rbE0tQU2BFiiu17ofjDcgs9FaXWT6SYvpv0xPasEfrL6sIax7N
BkZDtCncrVY5oydHZ6Zm2eAZLkZKK3EPBfYoOZnKUPzb5SiQq0KVEX8PcsYZK0h1mReI2w4+7/i2
vP6U6PL5IYhwDqfbWvqqLxRqdhbczaM4hyO9wJ7NIa2dxYuLDMsNquOjB83hAlaGHYI2VDrDWrO5
thYR7nmJtWcD8umMyFbxWFvlzSLCDbURxdGRQyWgpoJKYApgMIZwAVlOzkEZ7nJMVV52FH3IEtYx
jYz5DvY+8XEjrmBB03d9pTOHSmYNBAKRkCEuX9NM/A+dkXYPMxGbiOFRcFqVQcCEfgtmYZzJHoJj
/Kev5ZiAt9o9E7XlzJyj22HtBAyo4Ux/r+F/i0snl66ljztAAcGGIY0E/1A0oiWvZbTVetJ9vI7r
nu4iFQhqH4qhoKnpreza9kxpDK8+V8hsKV6/nUY9IFUnddevTcweuHhwev47DchiILTizIDxV5ir
vagmnSOhFbGQ9Cqg3nuqlHmr1OgI+lvVvlTzeFnmpVYLPzcqNeXntP7YnmbYy8Nky5JXOtmU/THu
RqPj+gbTfFA7dBaMMpv41JuMSAq+M28qg3l79YCbnSa2gHk7I1s8IyhPNI3oz0xWjpXDPmfRfCkZ
QaaQYWDX44u3VxOMqv8uENgytlRRadXr18tqwHhH7Phgz7BOfdj0j58yyTEw1Y4XBIvWvQwFNlhj
SfJ+84T2kDfjpx3XLcgdkQg7L0s5rPjoNIf5p9b8t+VReZsmwGqkmnec1zLKn4SBc3qnM+ceP9sa
9nrUKuWGLqUJwTknNHQNa8UDQkZ8oifo/r905OUmYCQfYepV10m5rRAhDQVVdsHZhUtYUfqLULmC
xPyIE7KsGlg5Nxuu3Xde12GixLR6F8SEXCGXQci9EL2a6ZPoAlstmBlcy1q+rqkAGhMgBEK2z4qm
/CP16jQgPux6ctu6CPkHVoAN7QOidhN54Mt/zaaNWcQNpLuEf/T2GKDVDH0LjtYrnaRQESSkGabe
pXXajwEHvR9zeJt2+ik4lT7HxDOK/EoN8f3h+/MVljU1MXdOJmZPEKaNROQx2zPyX01/3HS1TaiT
eu104x2cngkF91n7tMqlGfKAYmi4Lb1NzFQdL62NFx3oXLpkh1juCuD8fyLITmc0KOZ50Fm9SOMM
MTU2h7xAVhD3uZyLsyKGCyGofz+9zHWCCzbiFds55JEfTfWedKxN0jGF15a4GtozAq0VXeB+MgOy
CLegR4sU3lvYcG4v6v3m5myqMdfzX+BQq7PIoxyQHCcVA/oIvePGrYUbNGdnPJl13oCq6n2otqVd
a/czPbKQdFRl1L2Mnh5rVT/Rikc220ivRpJuCIqNEzEjDUxCs9fqDASZ9tQmqGqXilsm1BTz6trc
Jwq1yZywrTT4C5I8apqw9sim88NEb/zVMHB8RTl94SJcwDNWMuGGasqun6qG0pvFTQ9c22svHxZq
n8VC84UockugYEjLUuCeOFyPOIA4Zf4+kIgpQk3X6Ziyrg0iOcZEErZmRc0pf2ed84sRWbvYfM+z
Kd4QhHkULAzZ+OvyQkMyfmTzNuFta1kKs0YoYYdPwSfVilfJV3PoJV7JrxbHcyolU8CPP8gAzEJR
ynB7GXMHH58S4uE8JbUpzAK4pGqdkfLXbWy4pg1La+fPJ1nX2a25HNfGjNJQ5m1Sdsu9R3DqujfL
OTdXHIt9lbZkKKa+Hq6gBUgRTGGExSq+U73PtKUCaACj8haqurFWCRUXy7np/biJYgBu7i6taNLn
d+8Mo926JzfaohFaDzFJcOyleVFJgnpuL/CRO823KDP9sa+Bi5pw/1ysm0rBrbR5pjlYQt87KZ1c
eSXDexI+RrsxN6If/sgSIODsfNh4nXkLQ1Q7DlJ1zSVlwv5J5Xs2doMPB80ba1s6/LCdZ+r3zSJk
9yDp7ODhfUUmpD5qDCKCuTyXPGqj5M44ntGMCrIE3oV8jiOxF7+FuyEtVrYq3WopKXgAILw2chqv
h+0IgM9xIi6hE25nZBBErko1BbSmapPDUA3p+zHxCcFO/THgmYmDbL3fxu3l2poaVIuGVxsvMavu
qwG7o9NXUBCVc1liFODpPSwKoFWD2S9Pw2fVy6fdlybHt4HxDa2Z4JmvjoMbOYxlZGNFBjt16P55
hZPwpDEYf3yvt3tGlxcVPLJ15+oW2X6w3RXaeQiVuQgoNBTn1nsWibBqQ2caznOQbluqRUKEx6ay
0+PIjpqNeSLD3RHoe95E9y5rMbUikkTI+lFCaYWN0duvMCsQLzxi1FWJc3ogVDNt0LisbmLQ0QYo
hQXuEm/9Fr9jdNe85XdkOSZXuavk7po2MzFogXPJwp0t7P38JYVpk2vrvqjRU7fEV1iKKsA3UzI6
dcrpq/NkBb4DUvbDt8fJSSWu8zNzbMeqzFJK2qLR7BSV7107q4kz1VYL6X2YTjE73iyo/Yp64IUr
zBis++Am8aO461uFDdoSsXZ7aFyHWgD3E72E0HX1E2+31rnmyuqZYqaFnSV7NTfdnpRkK2KSQBNE
5vuoJcc4i0vCkFtbVXXNwOLVa4LU9J6rJ0DEEErCNN0mZyhOpkXD5MWskqUkJOnddGgAU7TkIGHn
rFsDRJBLGV6k9hqK5wGYOtNhQj3BZZiueY4ehiAutxHT1ODy4LS1awfBqMtnT3w9Ju9BFz8aHdnY
VoaexfWutKIuXYnM/v+UUCLV8+OP4/fGsxzFPi1k3EJCfWsh4H9pT9EmG/PWVpZG9d0OIkCRWV+W
M/9oh21hrzLp1R3l3ntWSgVcqDClyoREYSqi1SnyS9vko7GqOpGJ88oxiey4NH0XbCbPtb/nuNbw
R4H5M8lPc3uo9b6xLClMVEKO25enKdRtRWDoV7DwS1ItHxnuBiaEArfzFLZDp9tUJwtrRCObjB3/
4gPIS8pzxzPoM2MBOb4Ib6YFwpyBpGTv61oPhCg33yFODODFmXwALxtL1/MJ2vsrvykOF5dZNAVk
fuMhXfuXL1BbT0mT3VampGob0AUq9aFNQButH/knAQNF1/PU+fBsf2RuOf5HTp8FIJafBqRU6qwC
JmJ6M06SIJNBl+yM42at8QiMtegH5yKTr//NKT7jcC6l8fOd1p8xewXCCgD6CQNikPRajNEsMBMO
szy4vctSm8slcuOxC0y1j4HbIx+dgfCuANCYOs3imvy9KM5hmnlE67gqdLjXdY7eDJcZbww4MtyY
IFQ/vozPaSMUQQh4vZntvov/1r1fVoZKgfyeSCqSmIccZ8X+ISflvEQTCiWOUcw0bVHuwGOCNBk2
HbB/cbnklfhDrOCqCQ2vBNu8kdFkkpYrXPrYn0efTQLAep36Yrz+x0oPmN3S+qtj6k7fJAEU1KSF
cLODHmNZk+eV6y0X+GOZ/LKjyPRi7uzpVDnr/TRpnSHmN8qSpLqD9DHyDYfqGz5e0VucE/VEN8dm
y2/BpvVOcDWGbhj+qbBxaoReRvzi/8RLjKIkgYjwqHaZrKfyr0mbPl/YJ4ksqRoFCol6XslT9kvr
iT+Ns9LB/RrFxvLC23vDwH+49lGFoVsYCTDR1AbLk0+VKTzEMxDlgzbjhdaNGlYXA5qykUSZYcE7
HdtudWaWqXqaBcnhKw2KOK42ZidWljxhgoK1wYby1slWnvwm2EnQCg5MCKacpaPr4Mkahqcqdz7l
aBcFfuCr9l9VVFDLsooMVMuO3m/5ERK2vHMyR5NfyYau27AmR82hcJQ1ug9hW7/Mn/tYKGjan88l
D+XNzzveWmAfEraUWF1zAHqAodCA8nlFUC+cyXwbLZQAWuEG9qoycHo8JwwMUvj7Oj4TwkxYn46/
W/Kd/Z2ne3jSTuO8bW6iDCnUIfsZhJnxn8ICgA2bJCCcDWW5I1zBJAdYH3DyA2uI4fBjZ/uTbScw
hU9oCLWiLBihnzrCb6F/RddHbYArAaE9sDSdoj578adQa+4XACGprEXILEQLf0GdL1xfA2uco9U0
7Eq9vN5oqtUeh0XtnBYAi2MtLhQWyQkv6ShNzmglYDGxSoc0Kb3G9GxYrseRQoUbt7OwG5cT3Nyv
Sv6cmYVa7Ubo9IKuhSwuv15eziLPZYplWR1wVWlF9g70yX+xna59k+zo5OxGP3b9xruDmZYsqmCV
NG8vOhuYRJnggVFGR8LkEFaudsNs13X9euoHG/trLVRCMD6VgfLE61/PMyDjXPgaEYyHe13NVC0F
n494XES+yP2vD/hQzhMX35b5aXZmEaghNiWK0+4tbxrojeB5c34VoTFYhQumWmXA1zn3VDeF6mMm
UQzpHkQmiE5//rnBvg914fLaJcYtZtJfccns08pLo5hOZTD7BidMPkZbWEl9i1UsH/Vov7cixqvg
Jv+MNpXtq7EQP4MwkldVnlrXPvv+rEMgo59+HdYO4Lk9Q2ZgUTCRHwkLQ7mrD0pR+uXMiZgN7NRc
kEewOspkYwAyyc13sWZheKtaty6/0tpwG7qkFMumvsZMV8/N36ssqULtsS+OYXgkjWbYN/zlVFzu
5ABf4XCvhqN90DKPutfVTuFaAXhSnEjYAIQk3RnBvvfFP6YWOEl2P8bY3/SPgsA5GhS0qoByOVkl
TyYVnSdRHQu4VvRebQXPlARRJQK7oyFmYKKLZngizDh2v2jKATCGkFcIyd0THfugS7TcmVzCKAhu
XSxuDonBUNHEPP8m7qToeESL+1x/8tNrYcmJurxjgqclZjU9yx8Cx303nggdg/V3fmISsEy9Zd17
U7po29nsJoE+BP39Fi9x5Vtv427o0e2QQpxhnhbQYp0SVrGS4lEAchLeSDStwdUCSSGf8H4aK/IS
jk4udxFjEUJ5utGfeCtKTSwxj3UxrttQdXt9jZtdb5lD6DXmoHy7jX+uNUfhpYALRDSDae57y7pv
4sHGOokifLhU4G3KNmqX/qkNML+t8AU8lPgQhtd8Tw54Oc3N2OsCf4SFGintjOSM6N88Z84dmF1D
gvrzFN5FzHEXrZwPVXTF3JWFyNEc/NcJNRK+HVvsWwg15WFv9TOeaFKBglPk5O522/KaqreA6Ukh
m5hb9d6nyCs/BAMGyWJVbulUH18Kn7xU70mXvGmHq0/hrQYEQNaLgD4qDWEFjud5iRASshZLqeaF
3PoDLYD0xVfDWERF3p2S1Nxx+EN8FBwkjJv7IfoGcTNwswAKvLTCs6w4VIGO3wJVQek5VzByl3i7
IfkYPf+kXDfJw3jFmF4VfeLIIBTOlmSz6/tepDYeLn+a7e9gDFP1Be3UfVWIUDq1c7+Fgq0f0xST
T9MI3ms2vNSQuHZUU+Is9iBKGoN9Tkzv6hUz8N3Gu6aJEWW+/ntG7VwdBcA4dDQ5HPEMfxs9MkT4
UQ3nEDkuXVf6FXyys1bmxerGoVguPR83/QnBnDAoVMgfhZ2RD4+Pfu+gA0YbkNFWu4FIlML9zkX1
/j+NhoOpf5VSeQw+yW0fKT0reib/n8Snjl0rdYQwL8UkNytcbxSueUK0Vhgb+wMr5Np+yOZz2n+8
dOqwx2ubqEACBX5z+SBd91AwAn1FaXxfZd70Y7CySqruvFDQzBlw3LrXIU+ZpL2fCRe8Nv0Y+sQ0
331oAmv3n+YQdtUoFJ0oab9/HMX4Ze8w/5DdfdL121iax8Pcmo7mpufqTjeUMLUYRyhudxXfmsmr
vH8Oit1Smwx7oeOa+rdTIX0QjFCEUdYoKPJEkjZ8waeNR+yxsHypRwObnEN5BpJQB4KkVxGgfGLZ
84nTUfNFK8xvRhhF92jlQ3aYWd7Hjd36YEVpA7YkIYwHPxfGxL3fZ1ourQq61SbtQf2owpCOPF7i
Tta4CLFjYjZAaaU4at7cZC3Y5nDMVecVp+LZmIoVyFwP1zMXUGsgCzXSfWHDDNomyYLPDYwzcozb
jBxc955d2vVXdMtDAuSAoJ+TM03/kniLKGqQxi+OD3SN+yOIHWq9nDSyGOELYfLjoZES6KedwSBC
2yIO8gstr3aNclLe5qwLwVZET2T8slmWtyADmUhrMwhKbZkEW/Oy0j/+4EWKwgipIZwRqIk4Vps8
0xty+ub+At13UIaikk6CAfzuM3zWWoaGW022jdx9LrfEigdbDF4ul4DaT6qkCnZxJNJTP0OlX6Tz
9EG5HV0ZlmMTDQwyJcjkQSkpwFSpUCT+3UHUehQ259ghcEZ1uisDBzmbP5APV3yYcIWMY43l6rIu
bSEMxk+LNvCCJPS9UJlP3MOsOJM6+mbLxDWsmo8OD2I3MWRUGg/EwJcILZVmKAvUzjeLfjCvQy6a
baJhMZOXA0eSItCPu8N3RlD+WWe2sOSp9R8qlk2f1RIMgdosP50gRT1XU9qhPrc7YyKHJSqgLyKC
zlXZBkMBJmJ1wKwCgXAuHNxNFG/HZoRUFQm3A9ZiYOkK7AcZBDqHOGmz1qPwqKYGnMdO8f31aoOf
oSZENUH2j1gH7OUSFPsJz/i0Z6QApyrMvZht2hgeqhx2eO3jVBBNZulUBVBEeUkyD8/CR82ds8kW
e4IR76RqAkJdXQWNy4VYoxp8JCmv3NKfqjP5C5mrNJM2uA/N5Gf25kM25x3cI1hfZr9doxegWs8K
c8gjesFGfnlFcbuxvRE/+QpeL8qC7Q/uffnQ4+KaEmVKyCW3kQ/AzdClZR+NAgUXvFRN8IM8zHBe
F7a3j4WxtvE27AVj5/li8bEZNjqVj96Ht1uOCN62vMp9isBfVvBBSa0AYCbX/lKE5oEg7JVVWx4z
oWxFCdU7LtsUxsJYggc8Ab5egIWAks5GcJodt6cVN7uZjqcXRplQoCwT91B1aR5WlK85zmrzsouO
5DwpV/YB1/oSaR+7qR/TQ+2ItCGZ30x6ECowdtaqwnaUHefWmiSr2NW5cfF4Fvfb7hk4zlC/DLHg
96kouus6wXMeX58U6v321Sx8gc/TGZPefS94GjhfT1BzAuJiomL3yvTvz205Z6OuMyYbHDlm20Kx
Zfpr/IB2QV7Jqabi6LR3eZTlcpxU2xE7d+0iFi1I9Xpv+sTbs8vHVY/vzxTcLjGGvgiK/mZDIZjX
YUP7fs5OEfKlXaREbGGvAQebEbecOEeUmER0ThGwJR0J3wX9Ev/o7wX5aFwXny9ws9qp4+LhDI1h
9lnWZ84MnHD4D6v9TFqRipnu5aKhhHN7g84fMdjqxBUjySncTr34a35MZoUmRBBiNTNTonJ365wG
zTdNvS5w022srm3rZh+KNPNh4wFvgKhSVmEjNGwMoo+nCUoiz7YaWHVJ/W1zSdJUJBGRFqQ81ZX5
c47o6f+U9f/cQG/aNhBmD/3kiTHFvHQbf3KLnbD3DmEJmSHn3l3qmQOGeltf4a9I9/HQqb25SaAd
V/1jwCFAJVTHphmsWouvNzlxTZ4v8tsbfrRPmGrPZ7rSxMmrXpSxVSspm9Td/s+xjE6Sm3MU7hdS
pY2UkhtxVWxTY1LQY+zEeaLI6TiIxyEgGC3iqQOxnb7hRYfUJt9yINWgxFNsW1GANKwQ789LCowY
cph/bfdOo2ObOddsAYDjoQr1RPYAvYoTjYLVL4oChHXXMYDuIJToPbYJjftLr2MB2mpKsdAJ8Pec
gPA/0JH9o7ibLktqqsFXzEqNzYjgjvS7L7eVBaxrl0OYLawzfiwLPWRdV5rHhAqVhULrfcfOvtnz
iBd2UhXvMSzYy+AIY1GNLwMvU6hZN0EIQzLS2XPaLTMDLUyK56gQ8JbsRwMtC4dw0aV6D1hVbQR8
sdogrxPK4kT5vfWGlClRb8k1HXeM2eWVlaQUtANfqb5dOyYfcHj+FsOD0S2kk8dnwZM1fVaI0P48
YcKEl+7rcDuWBpUN+qn8KTDK0qzCPmhCzYPq7h0+78vdrXgBVf5NgZM0PtVG069ZHsPOoUiNUDBJ
0WVtLtnTH8FOoufdMhT52Tg2atJW8+olErmPBMPQy9lAHk4uCl08/zzVgMYORsKEEOA1hJS3r6f9
YkLBHw9EolVaB+sVcQ+Nsz1B+WAGHTHsKccjttY3iSdOV70gv43xeQn8GfQ3HhnmEvpHY2nbr7xP
j/RaKV0+0rvkI/itmy4bOTV8mipMZo/LvSLRIaeTkJmD6sk2/iRE8ezQrXgfcHeI7b2DQ6Z2oUoL
v7GRzPADgldomDmRo1qCSIfetxjVo+riBgmGw/uORcb+GB11EvxjXWxerbl97WMDIRbFpTzi6gnk
MjKynOjTN2nwfG5SPKfSKcdVU/Ye5LckCEZuX5LsBP96YCYjCM72BjFbq90BUGoebjGmY6Cj4XVQ
BTZWIM42GlgvMVUzQkE2NBF6rqk5jGQVXVyiJXlZnfNIqk3Pnh5aifcsTwvCkZ+YE20SLy8B8Utf
O+wQUZ5guctLdN+hRkbdHoMVYIv3I2rDwi9WW0Viegc6gicMVZfb0FKJTv0uwE3/CIYBDzyShogN
UBSB87dnc6l1C9+0SPoKvYPRKWG1lV7ucVA3UK077zaO9jBYaKmBCA7Pd2TBJPzpgpAHZ5J3FBjy
6TRFEmro9eWuDUohwzDfmYHToLSTdq1n9QMrOLcg+zdj6/aMmfa+2vHgFSYxnjTTHFR3gHMkCrXN
mV4f/YXkLi4sbdKcCzF8s4pZjCat8LXycKO78DyIZbruziZaAHif9XYLHINjaGJIFF7lOV78Id+u
r+Vi12h1rDsweumhXrYS0g5de1IJfW7+4aGeIMfk6Xeid85WlIc1qgUpR6fQxCOunZt/DPhp59YT
b0JGEUPL9X9kAY1+GD8huUB79LrmT/SV1lCieDupvOVsjgjAfhRIyCXBrxkYcRgVn1HtVodlWOh/
yj8haQHBGRo0+jtMYtoWXY7x2zHR5jie1Lymb/hBUGvPWSFsQLLm5s2botPrvcCff1sy5fOCA/KB
mVy30998Z+nTVOcnV1RzXDmhOjfiD2ajM0dEwidVXjetsWC6r/nvkpdozIl1jP0CzrgzPGbbZn0v
plRm+6aUHA/SAGKkN4OTbaiXvGLny1Vh3ZD5sHw53+exYI8vHO8x5y7N7zOm4QVAAkiO+HSkHo09
JHf8vYzBlfXjQwSuiENcF4G5t5TOKkmcQLHcigIvUvj3R8gcv3tfCFzEoSK04tWdbflM4KZUjgBf
2rid1PSaGFiK6LzcMX+NiiWzzSN/EdTrQHNPnk2gc6a3gb+T26GZaVnYl0yO3Wa2tuE1Grs60ybD
n7kGX+LpJb/yzdjHJXFhB4dduy7nKX2QRS7JpHMHD+Z2X3UfVpFPpxQEEPDNmee2gghXQKrFpHVV
bTfNvyJkESf1TCUyJ2ujF3H9vYZIQeObEvnCFEhhdVpuEwG1n4O8FslfOIAr0BcjMXaCcAE+NBYE
xB61lG1o14EJRcWVPkJ5EC1veMVT6OFlPQgkpLA8W1VIKD8kNVLkDoNktlYA8a53utheW66nIAyw
WM4G5m9JNnNDDSdxdPpe3w2M2PSM9bsF4Ez3uTgCfZfI9d92yKnxZk+UTxFhbVe+6oRM/NnFpbcS
KxIF2eS7/G/9MwvOI5Ng+9bbtQHCLxMmYXZbh0sy2cnV/ZXyMA5E80qq5psK3eWeFE0zZyzlnOm2
MxZGufwf3VbWsNiHkglzlFqPw/KA3x4DfygLkk/cWxW0qlQdpMUnttqVUJ1oNmH2TGMTgZxCAMPq
2Yg8dq7TNOx2htkkwXySPuGrUv1XvNEE8zNzAhABJieFr3c1SmRaP+qi+TAzGPiYGVmI6kKOJMwy
VGij0QzRVKOvteSqYZ26KIhNBLKji0itR6vg2A7A5XJM25Ciszx3NmKIuj/AgancbLHkG7qxKt7O
h4u+wtiKEYn28OfFLmRRKNY84mCQaoruFvqcE7jaElqQQfJFRVulVpxBAMzX0iOXC6lElVZXeBeh
HuAChS7TmE71/bT8QFgaGyTJpXwUETe/3H6s9rvQRAf/ucKb5BBqw8UovjKx0umQW4Pn4XHfqQ5H
K5kQv0BqxHugYTTiFGx7O00gsrmUg9GNsqLOz5C02e3oG4CCX2kioxbP03w6lYx6JvEYG0gSQ9yv
xx3ENc2qeXxp1UyotpzwwbiTO5x6HbyNKDSqhFJxO2BEHpTfoIPJ3s1YURdRtqyzIakLyLozjW9d
FRjA4EnvreHfhodyV0KMmRf0rsNWrxSmN1Ihjtl1J+8czhdYf2ChYb5AKcmlQPCDYgjV+kXkIub0
JC02aKeibO1O8Mmqm94Xk02BcMrX+I3F5B3Wk51kPff7UXDebz8EiEt1cnKvDaX3/4JAjd+8QPoA
UiE4jd7CP2HBTwhW7qPRFGfaihLdvWX2Mwgxm6P+bSCkU+NQPBneYXErIU7QJGFHTnnMPbVjygAP
dTUXDf0mlt6imvwhBUTqCFB6Br8NvRrOBqmKxuZcucAEBVnPiwmpQK02Sj1fcx8cNdCgAmt4U0P3
vUK3DCqa2rmyqSZaxKodnSbEz/uahj3wBlScbsxwYrJvQjCp6yJ+WN2/2zK8k2inNA62/lfIUCrN
GdhIMM9kECSkVXA7poFnFvlIfQQwa8RRvggiX4cYpAcX4Qhdp9ZDmDS/5bi+JMNKxpCw5n/Un7lg
D+uwEf1uH5XuABIjtHqjZhi71BjRKpiXeqXoZMkyh3mwMp5QFbualVj6soc1QLnVCqbpOCQnjq4B
ilTjynMctd9CtDsY1X250MiiM5gkccvFurKDb0roEW9hDNX47fds/cb3aWQhuWUrAzpBzhFJAOQG
VRRTIZI19HqaigIGMAuYJJ29ztkCMI2nu9x04HxtTouhKHuEooVUzD4jYJT913geIbNdpEfFrRIV
9RoTwuX9pc6t+5V2BnOr9CNVLn0EdAmlQ9GCGN0vmozQfBjFk1/PEMdjQrqws0nw9T/7SS7gcOH7
uoUIM3TNxozcJSyJcu5UMPDveXH06tUQnJjMlezhtR3Td2xpRF8fbi2m04R340JZ0ELgF1mE4MCC
AHFz6cCI8gmmXGRpQwnD6RO0Z5H8Ud89RXfJrmOXHtNnzL5G8pszvJXhkMW4g42UOwzVoBtQuJgC
hCJG0UGKnQUym6mOcLp1K1ZgJ4DqiH1npwMMqoyH2D6dsh/qZJsehkjimzI52dMLxdbXVKdJas8/
S3Ucg45rB0jlZZDkYViXC6ZF4zWCgfQY5iCvijCCpWygD6YOHXDsqMfIXkBKdhe5Z1LuV4Ld/l7P
chY5bNA46lStuU4kEeDFBc4ihtAUeYTKJECGJCAwbCzQ9UaC55/DXxLCaM48+8k5eHMFXyHl0fhl
OVco3ebzRl/U5rzPwjzjU8HzAz1I++rycxQQ2nryrD5uGmufnHsjSflsaxj1u4wfs9nJoHE52E+6
WzXhO56If2KDNd4rJ29JFboxL6CZMp0saHqpM8Fk1eNjYaE8ipKhphmf9OILLngAhGBXDQcmBj31
5T14EbSf+p8Yoj7Y11NQIHLte48bCMUsVUlklf2c/VCVJ4532mgj1qerLweMsXz/vdWbnc7hZg1Y
O4bVapTPB3ZGeaGT9hQs5MgP9h6LhHEJiuQ1DB9QbuZoAZyf/Fa+t1xdf93JsKha51X9eIf7BCOr
fwIXWXw/KZ8mwKnkCDnXDAke6Tg2RpHOik527A6uB8m2o5TmQ8nUGQy9MKHyGOpCKp1LG0Jlq/Ou
8FKr6KXoutc1LVkLswYVk9P5meyJ5vETE2+of/1+h0sNpx7NfBHAANN3GkIFKi5EpiaClBsw5Vvd
+E0An5D0xJD4fd49xh7u7g6HHfxX7cZXwLb+Xsmoyehd0otWrEjIKOXogXl8H+T/hX6dh7Fnxlma
g1V11lq4lt7E8UrD3q3spE9DpI9ZbCGQ0h/rT324JWXaOgf7NhUFSRZ4okXb5o+4MclGecm5Z7uq
ZM3VG28ta/6o2HXwCEe9GQUtD6iSWQ6AigtChugKyoWH4kn4S8tMP8bN4FK3qlFq9KP6aGVykFwC
gMHgC8oJD+C419x5dbV+WZZtjPG3SNJtOjn/abd0RbsV5soh/Cb60PSNgirG7kRpK9Mgfgq6nvL0
WZQBJB57SEgni9B+b2wicBkkFWtDudjMQR46kZuQxibLB+eyaGYtks/+EfJUr2o6hyJF88mAgdYU
AHURSRHeWo4vph3G6u7Po22UAjao41wm1wvSSUjOSyxsKeeSErZfS8T0RmKMaV5/3ve79NO8pKFo
JI1+BXnNgRrCA7Hp0lSecBLLUr76jiB7RBWHtzqqpwyJHq3lkvEMT5blgUiQ83zz408NRb7lNBYl
n9pGynwLsYXSdX6T8DYabT7xvfKsTECcczoT6LlCWIe8mNzQJuOnZv15mO/hrMZlUfPt+5Unvo64
OPP2JkOAW0NXAgRPBu8pRVa+SO4xp1R9nduO+d7UTqCLoUdclxvVC2wVHEBGPXm+LCvRi1GKCEGc
Y9vm8fpvO0+RLTCMIQZvwj+22AfphsTp6yNTjPhuEGtcx2jNwbG82gywoIQ1VXEeuyU55eOk3iWL
4IkUhXxzwGc0CzNdEk0TOd1IU9g6qmcIpGurdaMIYgrtX/mL+CpbznV44n3PAB0jbWbLpm486z5H
pIgqM1T3b7TDOCX8EhgGA7KpIlHK1ISkPODjBX8FD8hG1a/WA81+kPrVU9LW+SYAqkz3dP5USKZg
ERVZwIKM2cM8zqZTRNkik5+4sVTdEYJk+sxSElOi/UtZ4OT+HQNLL2JSHa4lXR8+r2wUjEre3Y40
AWiu33l3vL3cXv4GMyZyEqvktlAyHfcLqljLdzDNzU+XVF5Y6fwPl7ypVvCdGEubOWMrjpzvnf9E
rW+VIeAD12LFuxMiaGX2C4hwysKTjATE9X34I9lIOR6QIYJuVwZ/ofLt7Rq4nGJjQ70J1Llq84oP
XckT6zUXeTMqnNJdPpdVz/BeJiEBdSIhyleA+vCTNRkNWKmy47h409Ce43i5TEOwlSudaKTHsPtq
N8tJRm1pCG9j87NVNLrxmVbR9Dy6lSaw8fhpi2k1L0GF59bxs+5aLa/bkXtN9LhNVVHnntDcqfL3
RQXiz+Wy1UjPTARSuyc/vfqyyYcw0OvSBHInXhQYpDY8TFmA03NvvFT5pgM3fB2NRS7lsQs7za/e
K0mu+ocdhV5/X8QrimbtkIcjB4iSOrfs0SHoCenUVIi3SJ3OlKWrpTkjRo+SA28SWe+bNQOvq6XU
RfGpxI8yQb3lLCzHYnAISJF1jLVeHw0e563cf68rIHpA5xHFzHUQ3nO6sA3KG5zbH/vNn+W6Rufx
Z5zlG6e4ZZqadYn3JdpP/wgDa8LGjCYcjZ23yspv6D73U8RkruWQsM4rtqepZJgQOPjJ6kfH7A8u
QlDKMzyr8GDnp/r94E4aqjh5D4mcRQBqfmG87vZzlfAs47HtsHdXX40dRuLbZODsA/J0Khw1o9VW
GEu7K6k90h7fYS5Gakeoo7B0+d2a2iZYvHATGAYZMmiIcT124m2ryLQUIkmi60Qfv+TbjTGMwwm6
BVqtSrVV/JVroIkmUDX6PmzKLzLPbTvCk6Y4apYhAi47xHer9sTYm8Buj98jvgu8KTTwc1terquX
5OkQabq5ypvHZZ3V41RQLg1ZNp40cgkLwdIPHp0hlEv2Qe8RZ4X8JOQMBuSvrK5yMUDovTIcDRRf
Bk5E+hAqen6DvXCsdnJVIwqSjo8TUWijGBRD5zDfiYn1HFQ/aJdjHzRKzNn1cj2PKTCOYPIZljNC
orVWOt4jw17WiylRANuVLr2/cvUCFxGb42uF9E2QRtFb3v13gpT5GhyQl/hLJiXO9LZr5JI9feK8
WPe7s025dHfTp1fbWNfKzwzbA6B9E7t/BESGfp81Dl/+dQ0enaf+108r+dl9ATXo5GYKzPak+8JT
fVdkXyTVO/10Slpmh1ai6Ud9IN7oVlHZ4o1s9n8onjbXMCuY7noQySO2se5Dfx89mjsbQ71tdzzQ
cxO6DKoAXm38KeBY33z1/8UNGzMzMLcehYRQFUUpBBHdn2AmQFlCAuBP54zrLKHxaGmO+e/VQ2m6
vRn7uH2kHv/hV0jQ8sy5drlhL8/FWNupmTKqf2WU9FjOGgAdOb1WNHNfzFSlsGh7tdXDlYRZ3HiH
v/poHC68POQaLyaXbxp79BZSYL/gdbv9EAQKsiW55os6ed7FSi9N1QS8TwrYcf1qSP8C1OF7pe0I
Ql6QodX3gYW8GOvVl31wx6p3qiCZTFRVOTNwCqvlLQ0xuNI3bIm9U7VLb4QFZbIjzZF9//YR+AOU
5b+caUWAp9IauUTq8SR01V3CQUFBBoyiUYUW98IQG4uULJwQF18vCZ0yuyjd2bUuOqfQMbLwrXjR
naRCd6wMtUYRNh4SrGUy/shgv7BxvA5IwYSv0DRepu3wBEWkmfQ7Qb9KAG8NKEeiCsxvzcMWZ4u4
1I5jicw7pBCPU34aZGoa/cw23So8LDpehBHaXxQSeUyZO0p/itSamdlrTIR/0FA6t1mLtMcxr304
arOJErOaWD6yQVCMaH5u8TAYYinaCeHbWqb7uVhFA2HmJtxtUhALk0XlYfnLISbH5W7n1YksU70i
9+dI67DgL4lT7gxiIP6BfIctk81iLRtxvFL5xUL86DwKAwL7cdxfADxGAB3sH6eKh6NeIVil6/Xn
CiFmVSm++xJ8j1Xp51woP7F7leBKd/FPJS6CyI07VwZTh6SW5tyKL+nNrx11r7R2G3Gu3Spf1Qq2
lwgAXtSPboQLIC8Tk+3bwwKpeJKNS1NI0zgYwZiFPtwOsH3J0YBBgGPHsZZedbT/BUVf3HH6riKL
c/5lJu8ZDZUZIwfBSJZGORjkUgh6XH4WBvSZJDaXmlXIomu6DRPRIo4v4hV/4K2BYPUyDa8TIMKP
lZ84qfg3H9Mz9xA6EAH6rs3uBCklyVAHqyFq5CydDa21xubXXwt0FqtdWSFRQTEO6HvJpesN1JDv
/mU26b++YVe+asSL2fwnXZPnirRpJtaEYYF7+jqosJQELBL3SIAGm5c5uBivw6KNX3Jb9OO2TAn9
Dw7yVaekcEmRZnKx1QiSjgrhi3MtXGDHVYF5lToiSNbSKIU18SGlviXWwhI891tX2VQ5kBIHR9AA
wFVnAebkWMfVi/v1oI8wr4It+OIGrnNW5XX+HT48MMvXCrP+6fakE3IeGwkCh+qkiPzcch63P33S
+/hNSLU61Usp/jeEohsjMAg85bior0ZfGG3jEHC0c1HQNtzxOq8Uv0+o77YO4L3V39A9zQGw6HTm
HxGEkZ0rptlPpZjQnksfkTqb5ekyENy3o0/hprrjbKPitJCIfNDR90bvjFKc/gTD214x7HYS8X40
P/I2iVCyrLq3iJggIDjRbBffneD9ieSxGzU2t41V35rDrRsA1ts7edUF58kTstI8nVVUs+usgEOq
QkYglFWSVYmUrwczhy2VYBDYC8IXXvg8jO7a9YOZlq70pFTSnvNCn4JCfEAWNUzhyGvCeGAVcYie
9vKvxI6VgUaDLqFsFaD51JUrKAq0Get8x5h73IoPFEUeSUtcR40wTrtczfhIX/q8KeWDTbRtT7bt
SNSpaVuIIkRw1El3dyxrPGCBTSZE5Dw3VzcC7fm4DePdwWaqSC+aFLvGbJTMTVycEiIsKSYRBiDX
2D1+BZMKNY+PzlimR1HwzGCgwzdaJGkBR8xXMtH7EFb1+l6+sBEMvM98X0MIqXK8e4SHepujPtHn
SFsbExQf0slk9XXOh0on0SLnoQ3GIRh9/1JWMHqJj3jPgDvencklWKlDzv/gw88BTNgE165lmsRX
frEnfDKd29ZisxRpk9lf/cVGiNz5gSWlLGkL2AU0Iys2oMCOIVvhDYt6+b2hSvKm8k5TDPVP+rMW
dYe/6DTwPNP2JCuFA5p3J7rlT03XenhMxuwQZyBsDxqPz8/VcJM0Lg00yM/yTlw4fMLncTUv5OR1
TfJvvHYcCYsWcej+DhJtbs7T0LbTDkUxJFNIwsec1INzJrDvMk5Dz0Vlobu8lxyX/wa88B4PgSgK
eVulcuaVRCMh6wKy1eoBQvkqduJD9xZp1oKhdesFy5Q9/A0QV1TXNY/2Rb8mAcjAjf+mMJcwKw4G
pKklRuFhWhwARj0PKcBtCjswPhrcSy2z4dK6qpIFoVJiNbEBlTrr1gLxMxq8NyEIBHTDHRFNTCvD
88CtIC3AFGZy93mP+v1gkxs384KDZNsYVlHfr28RmKxAdS+vrYDyknnhkBidMlbboOl7KTm9q8Px
2Mb1MCO3J7bstQHs6ESxoD9/Bj599O7xOzGrbbJFNda+kX0bWE2qf6pRU3nnCCfRPdyGYX0HZk3z
7S/oFw/690K5ht191zdhRFndPDwuO+cMxCv10q7NDtszvv3w0O2i9vLITw7yFKLGacyO5bYE8fs3
2tobslCl+P81rPFMMOWlwkpMkLJyM3UhyhcbEe1C4QlboRO9iED9bXcI1Fwi0DsEJetRTZwq5Lnf
gj3EFuxbOppOiepy35oRfoKhY/qM26RyNGkwlCqYVYI4zSt5HLgmMy84IJHadJk/xvcg6QvJ4GhS
DHUSuvJe1W3cCfymeMWVzq4KKS51xxZYoSob3e+D7ZKEU+dxozA7C7Ql0+WkhAEf9u7cMslyi3G4
Tc3lFAYeQhtkOnKWJYY9xdHk+9M1q93egkyfwJ0JqFj74fl/a70ZBSH2qUJekN17ZqP60cZcY7pJ
3szkNPaqXKoldb863wylVHlg4RZbIpgCi8iTgMcsrERfeTil8zLpzrYEkIKbDs0jTPefAu8RORt/
gwPGLCt8NPCJRf8ZZwUZ3E0qwLgPfMkds9zmU1de6dFhPSor9CIpUy4ctogjHTON/xwBxZ8013m0
pgNzliPFuWfdljKxe+OTvm7rjlnuriNsizbpw5g9htNGGtzmA8P3To47t1i5VVlc+K2nWu+dDVBN
F+j441hgAdd+y/vqZXFBPUVGC8KRci21S1I1/anv264r+RUlq6tHFfKeZZplUU8VjPoAzi59nkIf
aD6W9n7t+XRwLj2H4HA9mu8zfNxGL0t1oTYzhnuldiM7yuf7f0ne6yiRliz5k3HWLpJB4iASO9bO
JhfarhTXL0IcXuoHUFrt8LzOqSWe5EYtqTck18dVhOVNVbyekR1AWcn9WO7wPFDBUYG3jjgUzUWx
tFVf0GYjGKyybYBuNFzYpcnK3I9d0t3BPO2Ui/RujeELFTvhh73HkAQwT7naYit0xBAEZHnDaOsD
mj5UTh3GSGZy9xmHSQ0bYzGCKoF9mk9W4CTQ4kkr2PxPpB8GERepElVlOn1gBj2hdosYBBulABVl
8OYhybd7jaqs10XNH6lyLuTgDYzvPQr97R0SVvlmgQitk+c7AeNWGWN4neo43CXsTR0x+2IemRFv
SP8Y56fD2ZiAagP+azHL1xR9ISMk72C04JqvXWE0raY4gEViSCKv17ZJciPxFTUUJtHmBUmo9DS9
YHr9ZpkxFLx5/UvROBYLOd4nIN20hnEME5Aw+hWey7HIC49YpuP7JMTk8nHdrCzLfSDtjZIvZL4Q
THQAuZbQVwYaAVdWTSl7ACtgXKXMLZA4W30l3rPzeKa7FFry+ROnUKZsAtF8GCOSycX+/VIJ7M1n
zaLugClqtcTulFD/Md4DhksHqso7IhmMdVC7Cit9yLMKFPSEZSqvOeIBtGYv2Qc5wy57Wt8vEowq
4L2hVgXPfsg8+Qo6MbH5vbAt51bV6bZ6P8KtEvhJFjGD3c7I/tovfVjcc6VAFFx9PXKpvpSykqLc
NvsaIf5ZGzGB1RmyIlnGfG+e7d3fzutpWWPxr4WCS5CEkHkf37UaVa6tNst/06ah6FP8jAgaqKjB
Jg0ZGyEml85gON/yZuYFrOkGzlYImdj/6MH88/bqYriuAI5Etf9IRXSf7XSdqGpxfMVj4CvOdHR5
fomsLyt0/L2R13eEunwtqJvz5+nywI+4oG3hZ4sB9Yi8pZCWV7BULXYjD3QLf3WBVUGYE78/zD7g
5x2MLBsvzn7IXPLwYAYibdiRQJN+4JJhYtrh+QYXgmcm7GCYsz1hSF0/a8DuZ6rEUd2HD5Qgkr6u
faF0307K+WGS8AkDoOWfhRLZ16yT6k6LU+5fMW1UrPI2eC/mBnMRaFdykcoq1T7S93ToYqOH9Raw
pPkxxlamUPmXAxcQC0T5MEQ3nGUler91MJfJ1X2gO+fd8eKzUPo0gaz14Z08ox3fQkkgpL1TQIcK
j8ScpEc0LSTXo0pYGYwymXIeFQeCtwcncJC8JFZPz/z6yf69r7FBJhNal+UjAoJGrdLUh/dZRgr/
UPe1cLAwq/VsPj0YaDX21o+xQr25PTBZbYZhOKI/3N9T0bBnxzsFLU4Rx9z8JTdXUY9GvjJ//9Iq
W295JAXVtbSekaVQq4VxDNBNPJnPBDnUrS0QsiN55B48mQ+9Z2kRlLEkIAOL772w/MEnsrGAU4yL
kdxUXkkRAoLWzSXz2AAhGDvXBIBlxDsD+x1e1vXoOC0uPgn6GN6cvYyavc+hUXyoWoLFlEx/TnsG
Q7RvRMiI5w2jeHN4H5+wTg7nA4ZwclrfajZLv2F8ukDWnFMcTiThQcacpQLQcFbxCUpbAqBpiQU1
hjPnKzZxiQdzZG2Fgos7x62VRxdHEAO1ru9kl6AgVzUgTtKLVkm2XOTSJBPU2DvQrFqXelq1nuBo
sTVSoQDbDMbdW5YRRXCQdE0bNBU9C/Je5tnXLyMWg9R3sMaLtkC0NwccwF1Ig+DvFjgeoR8KkRri
bjIUND7nRnrCjUKhDqLMODatsrAchVW0Djai9myLbO+BJ+7mQkmp+Zd/lKZtfgGXZ5LayqrU5Kub
kSk6UFnWuPJoFyO1X+7+vfcmEFMNBWnpbBFzsS1tb1Aq0EZDO6WEvFWv6NK/HuTPn2FYMi4DgX+X
MVc4tyVHRRLKvjGx9e9cePS7w//SjRN9TZ7GuPFKlLIq37+ZVo8j82ds9ddub4TcvS8bW2QtfPUi
i6c11ONs6/IME4/7MqodmPnal3aS7PBHl43V4paafPY+vertvc6i6U50aZm+PscoVfIPh/1Rdbxa
fyQKH1io+Odi0utvC6+v5tuIZQtsLvqNWGb7Iqk/MANnqctLQMpIx7CczqoWWe+/QhKRxTe9x4/2
LWI7p7QrMaHr/kt+lB9v3eSYGfpkI+ddDD/eM8xuXJ2j/J7IHcsneilnoyN4gqDdfbrrXQkOa9R8
OIRn9nR4pvgNgv8VuGAsDduDGoD83zB0bEip470pi0eqE9rTOI1WGZNsuqlHxVV/DBCC1fcO2wrg
dvFvk8ojc83YmkOcZX3vDbELbLiYL5gNJuUc28ubHo4KHDhS9TesP1WNAdsJTm8h5UBQBKVsU8U0
Y2/fBKB8odhT1wiDs5ZiRlhIQ9GSiosjSywx8XX+vGYb2hUT/j6Cv3LFpd1qSr4HbqxZ8g32IfRP
aZRw8u8X672uFgcXKC/bMSx3ReKsLhH0OdtyJsEWtRQhHUtMMiMygst1VggTVttT9Cw2ShTrmpav
R3XS0hZqCczwZkLuaWlCuUzp2xGvJTkoI5jq90M5HdekwO/Ueaeg8WuFyyu03lmwyuq1rauXDpyN
CEp6uqHRFdnI3n+0ho8Zm8q5y1ZzVqXmemdTkc7tQjJhfM9LiE3nGqh0gW4tHugA2x7dh7HswSbQ
ZKWGX6ok55Zzu+peh6uTwyKlM77Z1zITT2ZNsey6hkzHb2U0rE72cKBT9d+5gdWa78HW35GappW5
QrP8584pIfP84j/AVCAgeceyTcyuC6U2AmYHkzHlJl/cVG2WhDCWfmUqsG1exOA5aUiIM8VXB/cz
8t/GwoUx+VRG3QRt5Wpf6gQ2aTq502XuDCKe8l+eEmxvDYUn+d697ufItquAl8o2VqQoHj0m+Dh+
T4f2fyo6gBx0l36+JScETMSL1vduVCmqVns5fVCVAFfn8Qmia8IfzKQIUq7/Cku7b5CPJllPE2F9
PWD4CrpzSu/nE6ey7ZBW3fC99mZJA496j7C0n4AuC0qvIzCvYn+CfkLkPm2zVH/CMTbmapgvb66x
0g66nN7Ejh1dajtWWiTlCdR36vX+rjvpM9q1R5JwpaZ4ifOjkTS0lr/E0mws6p+nQswpetAKwd+J
TNyAbOfF93XZ+zhu0eDX5JvHwQA4cRFHf1hGm6bzHiqk23Dn9WbrXQGJNCZ5xPIOUwT8HwhLPhBz
da8VOkb+4O7xE6t4AocjKNBwCvYhp/a5Igvll1iBXFb0A6GY2xeYsYp79R57pecvZyRJmHj+q5YB
7fhrlPrmNCy3NJLo6HL2wWwq0kZ0zDIZG1OFksjJE1teGZxUyFWZ/rMtCaqOPhoFBqvxv8oZU5IT
BI2GaBxvZVR1OjtX3/FXXiPhdtH/d8yeMTL8riyVPs2oRhNlI8WkDPv++L9VLtFaOuwigL420EVI
JJ73FcfPU0LHzC54y8hVK7CCMFcZ9i1BM6Ieqo5uEgM5NHwOdBi1UuVWxV0VRbtGJNAzc0nRiKxW
Q/qxKXjqTuuN6PyF5xnJ3/VtoG2ZNzqCBc56v8O1e/3S/6GsmbSRdR6bIicwD6caduFkMREI/eUA
i25Q0pIyE3rVdcx15xhxyJWoy+lrgIPTlCX3lwABMaKX4dMllQFSzVI8VTOc4hTNI2+VZqxVPOSO
9Q2VnRkVL8dNG9dMzsjka2HlPQz0UtYwrfr3lHP61LgLabXv0/VXew8zYKLOD4KTcxy1DlYM5eDq
rDRuRNgaGvyg1jzOfOXlJWFVwxhbxjscp3Ps2A1wtPG5PIWayODEyAFzC3Rykbm4Kl8YGY7ASSKJ
H9AJrFQpkBWvkmc6z9Xr0VhR8gn3Dnj/EUIYCfk2b1b7gshWBpGxW8TwNcJnqV1+QBJvXwCTJOPG
fPNPDaJKNZ7UK6+LH56e/B0dVxdh5ejj75/uwnErwLkHrI/sJob5572W5EaXTSmekPl1U5XFhJiJ
/YdoDvqBsWcln5AWkmOJWRjepDWJpcMRuCE2mbZOR+Qux274FijEBWcfL73zwdmg0+DzOgG+cVAW
l6MhAeuq2LHICRKMEql23ivMazVMcMrIuvb2OHg2Mwqfw2FrkSsv0ZRKwTVbnhsI8rbkpF9VmsxZ
LZSEJ9IpQZAVMi8YSRI7Pjlv86cghSqDsWsF5ItGry0UowUcmxQnduPQBjPYhURKKV2J0pXuAWaW
RldNS5T2W0GI1ATJosIW3n1tfqwXPg9pYMaDGMc7hysNipEr6u8/4LhYvVvWnZmE1lUxxjbW6Xtw
NkQCkR5U5O26oNYqIS3G+u8MUZF1T7cvyCYcmtHXORih2ih9THuz9iSfsckWPRD35qF4r0SbrqvW
+Ohwl8CX/UfBaa1j/qRQKrUeTy9yGV59PVR0LgFACFh5yZGB64fUXHpDZr/NLlMWlhBJma5fgaXY
um49SHv7o3/sNcLNPbmdkgLMiIQEdtlvAx42r1KcuSlL29iBglqKKdTCOWWzXtVk99CquCT//sxE
FHt+zw3Wc76QyvyqfzG4bYnHZL6x5XPqv3FKiUUzopY0d52+LWbh/NeJU3A+deOQT2LgdjLAju2/
WRF/QXiQSn0+7MQx8EbhQiT6q+a/XRisXAUDpoTE2ZHnB7oK3PBp5yWhE1vHDeO92S48NqdA77TO
qaBdogAia3HRPJvESZgq+ccJP4Yv0CwbIiPZdeqW6b5lLj23x8DBBTOI1Rccd6j6KoMX8uDScAr1
KrPIurQiFJjavEBgeHunpFr2W+eyIEEs/EMcE+SDlXivsMoZXzzxPGbr9Z4PfcfHY/XF/n9/OweZ
GgT9Ne1hFOyBdl5sxXesly+O4lyFZzqY4ts48QSMelRCMiBp88B4663youAcHjCWL8JnT9wHrioU
rlFFr4nXdvONX5SaqmORp8Oljy2xMLPAog+8kblkz62XTpTT/SDfme84EyBohk/yKhRI2bGcYVZW
rVycU+VZ/iscz3Ccgvwx+3u2HZqOFJqQb0ncbrriEu6WOAUKpZt7d4hNhxb6mjt354LKOq3yJHaa
+G/AqLrq1CeYeQxocbFLcaZBqyla78Px3SQSg7w+8qK/mmA7I6l6FNt5pXk8iZbgnmluL/F5tRio
ixw9SoIPtDhzxG/rLETLlXB9ZBFFAcdjHpfDKadbX8yTyEmz3CeCh6DAl1EOnTvtDxhKE4jMFUUO
fvUfAX3GtKbnIpvmMyIJAEQjF+T/vIsbEH27P9Rh1yxG6ET1El8mIDUKn9Ibn3wnT7fkPA1jUlcz
AIvU007h3Miw67o+upBjr94yBUHl+Nrw/CCpnLQ+Vb2seeWOjTNtcZwglhMg4KcSGSjAf2qILs3Q
pdPHHNzgW0J0MHQYEi7WU/zA9NS9pLhmA525DhSUo1Qzls6VqclOxMZL/ixI94IhGbrNvn1vO6we
z9zraAXruxUe3L1Pg+oi33vEDznEaoNCitBB5UBVnTn/+x7VqFSUlYMhR61YnqN9gHrxZU9uyiMs
7E4TuPwYYpU6xef6yLbrMb8iHvIT8/s02OHkm+QusTb5aRF71NfGDEdtexEYmVsMSxTaybKcbUe5
qzBP9LLr/+HEU86OB8vXIS4ru4gPgl0P9d8BhZaKabrrNmt6Tw/1Jzs9eyvRckN4KJC9kXd/9MNx
sulAeLwLvk1YE5e9Qw+EEOUYN+6vE6as8T/P591z1dk8GsFBqdgprSPRFQ43shQLyz7MwAlbdBXh
odTMnGaWQLNL7NKDlequX5Z5rw5bg9t+28a5ujvOhdBBohYAclcFeqEUHNU46DJXhLpZ+eYf9bFK
zO4+QKrqDM7Cl/v+HBbARnkj3Ov4LQY/BzPm8LcYe+9zFyb6vTPkQFzCTORBHkUGSRYhddsUvmX0
6rXTei5UUOWfC0hsR973CugeAOQlX0+7z1FYtbaIkGL28cf89N8iuVNvO2dUeDwNxBB4TDn0/2wv
JEXfnOB6VrM3Lkvkh1h3o9ek2PtRp4SwLew+pKey+E+9sXJSmU+iM7FeSoaWG6p2wZHhq3K1w3x2
aGoj9h5ur3bTwpOWmO/lNutix/gAxQtjCWj+hMCBBa7Rb6dRa0E/T5bIe/Vr0r2w50WCSyrr+cYZ
gn/rO87I6OIIUaBSJola4uTTZB+55Xv8deWhAxrhyDF4sA+n3p7woiAgRkVSfEed+lxn55wBfqNV
FMWI390BWdlEd+6SzMIsOFjFR62pgy+K9N4ZtegHukfIc/FF4nFg5Y+WUzDAAS4ZCQlnvF7a1A7L
tm7ksprWnu1KPhZk1SDzKWEuoESj8vhSLky9Fte1unmT0WqU+UycFpjiSrQ8oq3+nydKmSbXQJod
L2BrL49L7ACgQt8qfwh0GrSON+S5mw+vUXuuQ2F1QOUfygY+S2XdyZkRJbElNiNE9s441wN6U88Z
uhB71+wcjuvY5e2RVTFAVZlbwNqvIGrB9T/NTRS29vk44xqjmdFbR4NcJXxE7A83vRVw+2jMTv0I
Dm0J6cey+geG2sY1LNRQQOztuv3iZadMKj7VXeh9v4sHsDtaS+GullI3MN+2dLUymcIRljAed341
OnGzlbW2K1mR6kp1DGcEihU2ibjL6i31jQGh5BOII3i99q35iIKotPDL7jimX//kh4i38tYwZ4wb
fJcu28tzPK8w9bcMAdt4Na6BoTV5Y65x/QMpbjDJEcJ5GAx/RVwExZgZlzn/YitCNwMPkdLgttrw
PSjJED8lWTDgF1Qa0Ycuca3R8rdDjgk/RraRysH+EvGZTryB2tCtLxGQpruMlpKmmVqys5bChJNZ
xlCE2RYtsWaA+3DwtW3QIYajzB6uY/Y5sjX9ErPz4kuhbYhZAOzJfsjUw0CV+9UeC5iqS4WCZaL4
0cV+AYCeXAu9GeQhK9KAKSHHInotST440sLN9Uk1L2cw7HjToSSL+jScW7YEQnGSIqRElUZL+skI
3KBR2ax2Ir9D4fussnaEP/loNPIRwQZROlDSWabosnE26FKU+4NjP8H5arX++MFuDwgg73iVjYot
X1uxlbxbr75+2AZOdbGpOfnaywKwnFbvULcLPmer1/p0KJu9gl+oUE2Q1F0+2/to53xMIVRe063X
fPVbYMK7M7pYtZ6IroYygXevA2pge6seoKR+2amQpjRhg/gBNyL/t/kzBiWAmIXX0QJF9Lu71z+M
OorIbjbnSpgSTrmdzDrxHglLEenycNXNlI0MknNt1AzJcEZShEOYtVhquE2Rcdgy0U/Xhc2CYUq3
Ww7fxxNX/ZnPBIOTB3AE3/uc2lNFOKQTa6ARoJZOLP9B97/YQjrEW+1IoQwdkzSZAcLRJzepQo25
4IM/E8rIWCb4YvFfB/PEUchhVXweEJAmjsDdTjkh5JeMjO3J5rPnTrHNkkiVJZYgdoZsKgPfnJlT
451TdUHfINvqiubqeji1sVbHqFDNEir0qg8USPq/sjelXCyyCD3gOL9SD0QkAsu9PHCwHmLl0mD1
CA2Mqd6/ZI7JBp2GxMfN33CS/VRDAyYXT0z57cfcpVYetDPMUlmqy/92qb/Qpl//GQK6JUPVt3IO
jGZZwYexfRUPxodT2iFiZeYotZ2gemvBZZtB0RfFeNR9ioCCUbBIMVhZv9BzafHH2zQq0CTGwmAX
MsyGO7Za6JcQR5KZHpjtcCCTSaAAlyfOMLCkYV+kd5hx7SdMmehcxP0GhnNyU2f7F62KGi+4NTvp
Vi6M+KVaHe/CcwsmytoVaIGupRyIrFNG/bYu37Jj68pIh5qcelf1zi8sF06LIFUeVjTd1kT0Fnc7
xk6d7evMuDR9ojvMv/UiMrRroSynj0s91aUOLImMkQB0yc9bfgYr/nxAZzLhjy1vcP4aM/EKyVF3
Foq5J6fvE8VzVdsJDaRDhk3ObJRK0pZrrB4a69iz/u4p6aQrGMNKq4nTDuZK6UyYkF/EPAqeACtN
IA0h7r9VNHbIz10qtHh38Kh38f3XBtTP2MY7T5oaOcD05iK/COaLlamceU08SPTXXApGzWVaKFD/
71XwAaLU3eroIxASea0Qev3kNe0kFY+8IJBioCg/+t1DPrZm2OuN228Vwrp5myZUyZ843QopR+w0
quYWOkEfgYL5W8JnLSYcHfbLQxNtdCLlUIZr8LTp1zC5e5Ig0aqNw1ifxAzvXQ0FP90OooPko9vT
+eDYh0aRRZgoqqL+O5yNkQTRyE90qhxqFOz1RH50LCwBP2X9AtTxXmIha00OX/DIXDURf6o5YqaL
DELi607RhqVDkQ3tDIvycU4uK74s6cRohxbbhHnF2d+kqzDTrPJoEE2kMOij7VrrmGDCJqsEgYbO
D5rub6Hdv0au/XBCSxGslsg1Vo3idnp9cYSkZzn1oflHTPVmqeBgfM+VidNFSAaX8ydkFbuj90d0
qwNVFi4dwYHiVSy18nW2HAlXOKo+DeIHK77wTKggcEg8zpxO76EgW2QjQTWJdJwO3Gvac4MztYRM
2RrT7TpHA0pz2l3AHW79gGUPz5KVOErULxh431+sw8NooZMrA1ES/fbN/MidM4nw1wWR8iJmtUW+
A0TFgS8pKZP7wyI1in5sv+6s9EOEqjsfv12k5SoPEBnk0+L+DJaMTOAJNXLGMdTgP52W7jMv6lAK
IQbSvKaoAHMofxLexh0COlGncc2p4KrKaGNIFs56zu5SsXk1HPZaF0hFk09dG3LOZgajJfJJ0OK0
5O5zoGGlRWL86oRRJ8JdJHraHSy2UkOaIeg/eulLNnZ7Bx9Y/NHg93Inv+VX8KJAK/ydg1FvH/gt
gXJJS6kWyypgOUll11htTpGSGlFKA0lklN6U9D8Ghyd/8Fx0KejYJ+Ma5Rv6pNpqoBpsMV0Poqxp
bGDhrTqjG4ecKUg9LjoHe4ytRNu9T7Gm7vtIDiXFIUQ20Begw99LcnUvVcQPCKNrcuWHddOsUDja
4X8ZiCVBqpY74osPwfi5UbzetSH284OHTPVTT0tgfrTYF5BkUKKFyf+qeI/qORiAvt9StvCPmdXv
BAJxoT3iISqgMfJg9Koqti+VteRa1lD0ZEP0Cz9q1vqgh9CK1cz5EBYFH4cnfAPDa7y9tIQaaQAX
Uj6Wl5eWqrR6s8Fc3ydcPHNL8DwOrUKikNKdCmLF4mlov8hvBgFog2t7xm5lR6+MSa1YrEH0EHA3
aJKE+KHMgoCXskE3aG0/upx+gMOWkzOaIwYQGkoMBhYPkzGRj8O+6PhZv8BLnMB599GoN21JUfNC
h1sVioN/GRI35umiVnq5dscQe2FTO+ENuideW9RywKEzilZ4ASDM6xzSNh0dxl9o4PB5Rctr0ejb
S4Og570r2Tf4G69+vmjXfOcY9IJAUa332T43qjoKowRqKe/w+DVAoz5HYUie0bbBPDM88Jzny0CD
8VCqufUWu7XKIz+jMxlc1R1MvuvtoNIYULzqCRio4NhS/2wvNBn0JcGShIP8mRo/1JFB/LYpDadx
QDaBe6Ji2kMHEnCgSQCoLVzqCNeHxk9/clwdSMgr6EnldSJiL+jnnTJt6p2s+uRrlIXlfiq6WJjL
R5Sle61FWTJuQiU22+abwtdETtZl8xQXDWgiCYn4h/J99dgXqWoK38J+FNqnRQi9UONFRTwzX7IM
mFUuEHZW/LHFEnSxs3oC39UFmnJKxIcpEedSZsNNBfHqB+sG7s1o8uaVWNPWX1oN/inz/wBiMkfX
w77chSST5I8nhIfsKSLXtkTep6Vnfy3NxvVUAyCOU5SbXOYxDkOFGc5+P7rIEPGvDVK/WkdCN2h3
CqArgSxY7JPKGaEMcYd0M8c0p9HHcfjAQ05tl7CZKDolPCk5B2IoiEehj06NLs9OlweDyab3tWNa
VhjQdPDT2QTETnTV7PS2+vVJfMSox9NGqlh+FqhGCulZSHkcDq53aYemZjJEL43APh4z1gEcr8fN
F6WDJcwhK1qZ3gaFJHiT0QQggLH6IUPRBEF3dOp6fwu9lDRou4LibozdbONYGQF6NjxOAehprgYM
JcbWydHR8Oo2YWiGDKus9mkqjFKIKrcwfBX47yWAOxk4I3ISLR5tjr4LyGqL3FL39okTNkS1BUZd
a/lZDgKD7vzYjF0Qwc1zVNa3/7MnTrqHfLWb7nTy0T+MxJY2+LIHOQ5W+pomI8oAn2dIXRbZNEdN
uQ3pzFTUVS1Bl5vFhXBqCUI0aE5pCjBKN7xFYH4bEVmDJXNCtefNib6YtJtEZejI60cDdIewR9B6
dxwgdXdTnl3vDyD1vyzDTC+0aFR9snm3sD1Bpp+KV+MDf89vP+70WE3sHJLkN6ivFBCre2BdK7IU
XkeYdQV30CWNMYiexYmVG3foLuakIbuwMc9ZY9RKZoRUJmIFM28uAX3/bgciZCWiKHQvuUfBrXMa
en6Eah2IXr80ZjYhhc/T1IDGbLYJhyUd167pnsI1s/A+W8nYuZvM9wbzWmviABdu1VlFm7RaEWiq
rNNsBcul+RBe3bcCmWRz2Ylz9Ld9Q2sjDJDi61KgWUo/+dDndwAEKKkVX9ZO3XOINXz3J6BxQErJ
ey72kIAD6CgmCwLur/KMPy7gCzM5G5jkbF2a3mvNQ9UPF5gvysoCDDCK0cLqXKfHA+3CRZmREAIz
TspuYUn6cs0mRACl3OlfgPlBurJmEqdV5X3m6oQeGgqvdydaR8j12SwYSRNYdL5ul208EFmHK7EA
YUVV+HrQ7+ckhCsnUpiB65FIt+w8bKawVaLQcqKbNC4SGaNMU9/YSc0dOxYOoKGL+t7neKS3QvxE
vFXY6neMn4htpBmOfQSievuvCizUQXhJAUqRtFFu9maja9PFyhOAI9PNahSiKKPVh1NIr0lpGqqc
XBfZcLctV1u2kVgzrPKjp9C+/y8XPm6f/Gaw0oMG9dBZRYKzIi2fOFXiE2FT/6tnbNlcOq0QLSvP
mAGXoMkC16JEfvWJL7iAZvo7kVGpiv/KpbDPaIvuinQ+S+q1iv0PxUCYq/pX4NqRtnVfizJbIjqV
Kv3YLM5IJp76zKnH4/kqsj8YCEEURG29kT3L4Dn7RQ18tpOaDD3VFTGQqPHgpJSLs3OtavLcMSRC
1BnVX1YUeoaA+1WqpagiAXONm6d1HyoB9Fydtc09UA98lrvxGuZtyO6WA/GWUaTmrM5g5tPbpgWi
BYey6rL5e15pX8jhuxE24zyelOkMyl/d4qGbhrVUl8jokTI95Sd4R3W7hbnfwyPHVQ5IBbQr64my
2dRofX8B1LuOwrE8O+YObpc3S4/U46lk+vQXtvQt4Dar9OK1bHwm+QJ3/WAXGtu8FQtZKzDZx2xO
okiYdlJ9KVN8N7vANFv+r1o4AfhgnZwY9xfPgpktMCNjgGkIMIQmkm/aUSSrAFjXUbcs0AqONxBD
58aGYK0cUBqvBC6k1PqpQcby7i6tIUxuwl1WmrfIjJX/v4FmQnfOjFq/A7FjTPTTLOxuOUdlJ4Bc
chQD9KdnT9NqLqlaWktTFDhBkrEQbGqd1j1RVLyomKzRZp8/Cuv/8OAQ0NarXF11/4Bs5SN86vm3
WbBuZXydqMOsfRsuDfD3El/wsFNr5MbSq93gR6umziXn1XHdIiEaGCPvXq3jlBOTvP8tv4KG8goS
jM/B/scpj7SaGspSmNHOlBKcL+Uyf68z+/TKg1HB8iDlfYOap1X3H/KwSaoMeuS91peHKpFhdOpN
Mtypw4y/QrvAaymwtyaVVK/7qbKBiQuEIfN/P4yKumdHh7FE9F6cGO07WnUqdxpTAwPZ+qmlDBGT
CsGZNkb2MT4+6UnfKp5jsxNVvbbED4jnBPImcionslyPVxWT3oKREHpfUX+Y9wb78eBBO05Xc3c1
B3Mu5yF0/U0nOL1w676W+OxeYTZg52M0painhJVCkR1J+XeaHnfQz28kTIZZf7e9hDtPMuKckjq7
GDrjkBGgABa3hl2jQoHqQjrx5QO9Gfi3D9gaidyu+PqYkIJnC2dg1rXNzUa+PzO8nIrNnMEtBOxm
NNrNGek7+CJIV0rnjNtmtvtIQq8ha0QRgiuu1N92EWKvFQcXZSplhbbmT2k39QG44vvnaVsQoQRq
Cv4sTI/3iQYUrh1FSEa8eujF9IWWZ9k4OSSYdYpIlrIMVxx0OENbY3dlSOtnsJpjITHoVZXWYpZB
GAB7/lYfqMja8dpQIZPGzmlhFeFYW2tzPVDhbkfffvg1ik0RAkqWswKdTn+j6g9bgguuCtVpHzlC
/qDJFQnKe4chHfbKYgaQGLoIP45s+a/kyZCUk2+I8AH4yTdDfR+3zIWCZTQx3rJgiP4CYyX57tDe
JrrB7Jmov/YSoG/5bY2A8cvl0TigIrdpyEhuLH5dvvLV3JXvBVVERtdjrw4xug61J03X0wZPjKs1
P+8Ra+uZUHgTEB7oBB+AyAllxxJiAT8DpqhsI6NUzheSxbvMxpoqwvJR7kQQ3NGTvyRqgHmBiMZm
NUNOpGDzBJOxJ+FXHBRKIW9w1tQjxxU4JDICqcQptZZIFttz2exd9xnqOmnmlzxFyYfX4tDBXerK
uliMz4njf2RwyBphLFIVAK8k/lGTIbZ++SyNmTu7z7chFfhp08D7/bcIpsaQlD3NrGZwHdFWl6O0
0EPy5QgIdzXoTQ5V0avwtOtLamZ99Bhuqb0r/EIudrHLEQTlfu0GlxLXY1LCGwtROWQbW3tBSc7P
fTPH+aw3xbS45b1qk/I8eU6xiYZ81iB2MAskh6RUYThzqlNFEU8C2VOyM0KHtemL6jbHog6Bio1Q
ku9I9kE2hq5OljxdZWF29996tgT/r0vV83Q+eVMIexvxmMAH5wYnz19wNtp6VMuRT9kF9Z45IJ7V
jgWA/v68ibhHBGCzOq52caYK2Dw7GmV+pCnKyu7Au2j0np7GGAIPlf5kbHb9cxuJdbcdkQFl8kGi
AdcxsVm81eEPh+33omyizANXps9B00vRfsrATn2J1D1qCPZmqLCoPl57/F4a7Ld3FdZ7CzX9FYul
p/JlHTrYxQlU4sswBPZD5BOWhQEyzZECAj/R3cEXDMM73MXeScGhij5r+miKC7WDmANXDFc6Albk
33l/rNRhtYCkFxrriixIvM4PLq/lEE37Of4SNz3w4CydDAqQWRW5xtk6evCd8+rfmMTeXsMQi6Wf
UWV+CI92AUFa26r4/ocaLfolmHGwpSCUB6nPcA2s3iLVoJvWQ5yIdTzcRW2F7RJyp/uUJ1m29ecb
MyILoQwXVwGTA8YWVDgR4PqNPpOYFU1v7sf2u7wejX87ajnMoSE9mV8wNp5zngR+wfuSlrdHsjkF
gZKM2it4ayMjCy2hm3Z0DaKx2Vh3bP05cOeXqjZjSj4qBW0nssMrlXn68J4jMYZ2ugL2OgyjQLRE
ncUtej8MQMOrZBTQqrzyh5AHXGlZncqfSMP33RgvhXx6auoY2mL7UhItQxQS/0qmcBoKP1fg+XZS
d/YjMdv68OOP2Fsg4iaer56yfmTNeNfxwTxoevOU7s6TgyBHIz6bc13afVKCDbO3loGntWGsEU1b
r6KiC/nbg5WectYSDYFm4DUDfoAApsUjbi0FM+4IDArXOvrE2RowcKH5IwoU89db03QVvy4nqAZQ
5K4htlaB7xdjx9NiSq3pLkH/e7ua9h/ePJH866MJ6ldE8Edp+ZWe4lPlIDVMZja0tQoNnfIDiCbE
FTLncZ4ZD7WVuFqLnkvBbt0w+lb96UD+PxSxdhaZ81wfmw9rgbz9HIG/SwOy8AnmrGGI6kGrMvrc
56vgZOsgUk1syuN7mRuxsbQWeenlDlQ71wZHDA+wBFbsDt00U2Utz3Qd/gu1wfGVevBTp6nRWlAd
8SFi8juo4lnHosED6cvGPHfnSpSDDLAoup8loRDk4peLEddiSePXyxN7YDZ8OOW/yTco2KjjxcuU
s+vbF6iXb5mZLnkHligTPOH5L8TQ0ezUOOeAIioLwYf5807gFTmlC3/ijRF2D9QAwaNjU+0JuMKP
pNCc2sB43mYKs5auBu4JRmAgrdOWyYDwBDlyLlOScz26VDHW8vY7yKQt493GAOg2u5V53S2JQWe+
rQCvVkn0zV/+neChCRnog4MlB7de8+y9lWEV++NqPunsR7kz7yxTF+l4oE9ari5uX/sS2p8MxX8f
owjqBQzuPDUwRQz3HtdIsktib2YwgmnT3ldeIm2pK4WOz0OmC3s9CYnAU+YXMnBpXDcBLD6G79wO
eWIuQFXQGrI/3qNoU3ACM7V6knBcWOgtNuWz2O9oNGoKHcfpX9HRga6D71YimOYLsjJJFKcm2rFX
oBHsZ7reSm7SMrC/NtuyPLrxGkHXJrOH56tZweJfJNNHRGS/BjKx+zdsUFFcjT3DEgHzN3F3Gc4r
EQArFCbFmjclWBf4M7a91yKXKr4v+4evu2wVi3/VwKTll//YRmbypv35y2IalFc6xJU7ffcGtTXr
I7J3fmjoVhqbZVj/4mp7OaEb/JayVmBAGUPWFILMZCnOlzWV6DnE9ucACsUGXk3O5qIWAHzSH1Zo
RPwS7gTcgID0LrmJOPJ5aLq2ympGG+glA7+wxavOqtCQmTalq9Cbk9Qjvb7EoZZjo18Xet9sg+wQ
v0KpGB8NHT9nJuYqRhZFcwjXzJEC82mfgOpMZcrEa4sK4aKeFcooefbo+Dm9K6dmcneaMWv3nZ6A
yz/JUy7ePCE7+99EfGSEeEn4hiJcyXlpbf9i4o7/tQOq3meGstTgmUfmZwXd5DoKiQ56iUFauU3D
RyPGM6AKpBZfu7dVTGRUfbnp+YyCiNEfa30eOGBv32gRTLE3CavdDo1F6MWdMaqTnXClFVrPBzVB
dVUmCg76TQCupKkgXPbE88EgXF4M/I7we7gUx6U+a/SYOU133BevYu7FEe+f9GsPSK6y5n2qaC03
cDLsoAiMrmiVMVosMkaRqYfXmrPfpuakFZlu1td1KGhWGXCteXhfBReYuo/0bEPw7GY2B8sBkCFr
fx1tUZ73AL792D5ZXRaDBJg+acEPpUtNfrwRwxv+dWQiJjZzPLd4Q3P+jqHjtZ0LcMgcuzkzyIbw
Pe0fEBKdY1cEfsNlPMgTqmwEJa+OLN3qeKp2fCfafREB2Q7bm7WT09cCKPiGYJiVcyTTZD3th9t8
JwCQvqC0uXiEccWxmX9x5q+dV5yd4AwZeXMgaT7f5DLcxo+4YHoyaYFwTKk/rirnq/ozSZlAH/6Y
nKk+pSOxpgClsDjL00ZgQqmz6vu/CEPnFrSGrLRctVUcukynCKdCozd325ncR4gZoNT11JrVFvvD
BvmTLaVSGHqD3YORhXnvUh35zvDruIfNdTQauBVUoLuaVo4xco/Z70rXWKGfOQJ6olwxsSAGHTDk
zUYuqm5zD1+tIRTwHZI0yqG+AC52QtFaTeXbSIXsSuxyXGryNhGOpbebFFiNwG/bRwQzkM612S+W
Q6uXBa3A8hbK1m2xqYEx1mcCciEmBLGhptqIQNpJJhAyJlLnaPHHx+qDjRuDI+fTeJdzVItHcpBw
onRpQ2jc0nRMJGdwEAqLmHXEOhUClAzin5oBHgTsNoDnPk10VMBM/zZP6u3MhZsfQV1r+X1XnzsX
jzxZWp2pYavGV+N2CTU5lsL1XEr0DmVNpP26zZdB6N9GiiY7+WlIhs8bGqIESe5CVlEK/ci5dZQ+
2Szyi7q+r3rLbjWny7pE14NhwbqwmgZs58Nl7b3LDrppCnOMo8iUPX9g9Q+zbppyKmls2XukqTBk
PpXDGcmdtGEwJYGsJ/5D0YoCwR9vMoDt/Dgsxnqzt/UjzIn85SwLZTH6F97nEPRt5uID5g3PB1wO
dRLy6C4RCAc2P4ksWKVE7mBKxmKc4ZhBjVmB7dAkTJfUlw8d/f8OcTMiM3FaoO0WZKKqBU8bL6bC
pJ4G5XPseDZOPvA8XbQGObZ1ZXG+IdJNvlw29ghVKvsjlQRcs7Gv1akcxPqWV4cEG0bgnKixRflU
bEzOoMxpO+pAjxQfDVDNQQVdJTH6C4rfx1n4/fmUh+jcYC4+2tqupknYglDvyIXDym9ggmLq6sbx
KFgp/ueUjCad5KbrysNQm5xqYtGm8NQfVZgCwS4GEhd3zQ94SI0rfDZ4oLHRTh0HCObuZI5+5EJF
fSkmQBY4Qb1nX6utQwEMPHc5QVFNx/wteam+FfvKQ+PNh9LqxQfkptDXWdr4rUnZ06TdrSoQw4RS
TMEiKfvFTZkDW0EvWM2eeFYt1vhqtWBYeXNJVh/wU5CKzBt42pn4mFFNGE5mM7yTsDp0NQUGiI9i
YOzvGah7ggGVuFJtEW8Mdjmnrn9UqMeGg10fi7DP5oS5hlR21TFa2yC+rlEGtdqSAzZG8bs72itu
Meu+XRusPQVe9J7lfmyCuG11F1mS+JPXVeiMsXDoj9924dAnGBWeJXkfJdmd00ByyBXVtZ+gjs/j
GCaNESFoN4f6qQ2BzurcUuzH+Is0g0jA7k/VnqcuWB9ePcD2NFaxrseEUsMi4dmKWbB5p9SQp5nv
EHhZ4cljw7hjiqwWnoVgi0XYE2vO/lyq+OMqWghg3Z5mpM59xfDmYTKgUsXKddHgA1K4BdfECs40
sIwEhBt4AJJNIU3QiPJJSCHzCO6Vlh2LUdE/I6zQgjuy2JLz8KRA4uzFM8xhrfUb3BttWHJ0q22L
6GJe8+P7bDWBz/joL+biZDiDsp6tEE3T+7reND4E9/6ra8lNvIyqjqRmn71qO/HxlDniSn+3p+Wl
IP6HPZdM2NS767a5ZW8+J500WWy1Y78gdOa36HXoCIFWtBsVIQCitzKPna0QY0TiLHnrhHs6ygLz
w+kvRubq3+3095lVGE44sk2wUl7wEZm+nu9cpE0BN0zozg70wKeVtIeP5KbmVVDPENkMuGs7M1Bc
52rFSignpzfYWXXJtgtAU9EnH6xieHQ31r5tLKibPbIajU5cs/kDXcCteOehobzFIUUems9PcJYm
e/7g6NTpkzUYkpX0cW4lVxsuhyvPzHQqx5E6pHsdfO4ZdddQV03HxM1A0AVpMhhYTY9U1Ud0sblL
mPSQYleIz8qH8yIjGey9+wU7hA31doS/MyWOk0AEQhPGtbTZ+D5krZuqO85L5yJkxCTE4UjoMAVR
APuNjKpJ/xT844grbGwOOLH3AZdiHsOqd4PMAeZr/1YQiBiKxwyunU0lFEM177Ufh+ksSk/LoXl3
LjY/2XDstrupfbsrlxGT/KZbzufAHccB+v8QXcvWU5Wx5tvw6ALhBYkgZKMrEgpWCynz+16eo/ET
kngWBYmmL/tKfDHxlYh2LYjQu2Blh7D4EWDBYYRaAfwHoSiQAxYEvChOOD5Rd8Rq6wqw3YIzuJl3
nrSHZ8q3YiACFlF92GPpkHtL9dtgNtiZ23dCWhNSI04McSlnailApbcbGqLnimADVN8pzm81UAoX
djqIDU5BQyeTvYltlT82Jnjrr5etz8qlzbd32fvo4yxWRi8EsgdWVM3sa8WUIxghFXPU27GCpikz
3IeT83nJB0mGdmfgWJJb8NpTnWsrVgwgzGX2K5gTvXC2SHnNidoxPAT43ev26sywQVcxXyDZgdFD
3rs5+hyXyhkqyBtJr9aWJHqUUep/wnL8Es+o2ODye0cK7WAw7BeoTAXAGiRjSvnF28Zd0q/wqtl8
T8dl1s6+6Frg443Q74cl6QFFV34PjpF0V33VB73cdDI044PHPj1ZLeirUSHL5FmrOxFwkrrWzx33
r+AgDt7NsCdBPnTUbsdSeukct/ccz7yS/DodT0txB0m9YwAUwd7KTd5vj+sI297pszEuGCe48+dR
zgCrFqFr9KP5R1HuvC3p3WL0EADj5s7gX0jwxXMy9keJ49w6mXNswcLanLhlIilgkGbFAB4RDzY8
Sk5ma9SVTjQAuolRrj4LnveJwpBwW+LAjr3NG9NZMXyn29m9RYxPSBT4ZX2YJtvLTG/FNTeE+J/+
WUUuU1s2lrR1X3AyfUsPdoZkfhybQCfSOfLTUKa1OSeTzmsPqYyeelHx/9xuSSL4ieCOaZCDtOFV
4PCHhZvycfJdkoFsstGf7xZLhE9mys4jV2ZgQrnBiOCobIlajsk3evl5itWqyGMxfBrx4pk8a/Wf
onGzPJBE4rjMv41yD+FdCxjo4ExYeAXxKFV3FdiPn1vb/CPEsv1ItxSAs/3C75py7b8i45dlyant
QKePiiMJd7ZfIo83xqmxG3M27UVUrYAFNMmuTeZ4y5wHlSaiFzEjTDGEdy+CtXrarnrh89SDaEGn
jvl1yRnF9X0Pvupn7tf+xpga+nFXdvQc6hc0+kStxxpftNb0BsS6LNFWbv4XszSXdgPADP5eQlM6
5GKWoZXVpmOMstHwLxY5I4eI3IFA7LlNy00rWGIDN7fSVcBjsG7AyEj6G17aXgvuUyubxPq6mxiD
aZmhm6SQFlj9qkpIi4UR/5ZmOMmtbFRG41FEVP3ZDGflu8qD/tMx0nPb06WHsB1jThqX5cba43IP
3CQ974bmA15eBpGUApVbUoqdO6H8+uaQRIz1MYrOqrwkK1CfK9tRvrUgXh41F0UtaSxV0TnGOyZh
hYLSU+PieVPAHxNhY2rdpr2TNBKnCpJDHQMilQkPl6VFTG1uwTZuP6v+BHt/K/rq4C45EpxOJNIX
esx5uCJkZnLUOWN2Pw/WXmaDxzxYafUS+YaxE6i/4pBVB1zQf3NWRME1KtTK5Ei9/cSP/0A1CEeW
oz+nj6qqu9ISurGqB7hzE9+IlzaJsBLydYdo9mVWyta/IZVaENNbvqduxARwALN+A0tpV63EJb8L
i1dpVBtHFnITK3dUczr0qPdkCTghGEY/REFfvlI4utHS3pQzjepIyQSVChOGZXI58x5E/1R7vZFA
GFx8K6bnE5O6ogyfeVcbKGoHcDkgm9RA7iS7q9XhStE+crDwJqHfEDBVXrFJuvyUjMoQMDFkNVNW
g3FP9eyAj2U7idY8pAsMgPn4AeqcCeVIsv3LyhWEIX5C4uFjeWC9/A+9Qy5UUDhDEYfxVZZTJS6w
i/olS2AL0vEFVuuXhc9Us7jz5Lnn96VeGueEZPDSA+FUlD7NyZJpJw4MRxa7THa83n7SgonYAgy5
S4MT6kie68/OT1dGRxPKeRORD8VWWT9J/RNUyWMxbA/B9uFhY3Hh8OJB2GpJs9e7q/ikjLMWQgoY
leQVxVBeGrdabK+W7fkAEEmfH8rXMFkQnFCXHHUT+4GjG+8gHyoIdRettjtoPpwZ681zZ6buKGRn
DxjgCgTKJa9zwjqkwM+4V8oiEUntmpbdxBNuhKzie1bC4aJNpeMtfWLOoPvkHoh599qiWZca6byO
C+9QEefKrsA1UWpxro1Dy+Tctg+XsPJNW/Lnq1BtmsjhaQAbshxytGsdHmSI1cypFrsvvI1RIbSZ
VDJURh2J2Azk61w7Fj2Bf/NEiJqdmwo97G2Y2cP4woYFQviykJ/THtsqGutOyvb9ub61ELajDDA7
BwGLNExYbbRU0LZ9cVOaZD9s7HW5HP54nQ0haDsX2IoRponYwSMUpemGJlmAAbaLQimD1+7N9+dW
PqO/PssMmQ2OT/BOYbn19a1WaKybSPgM0jWTtWSyBe3Er6KiqVFLGDHTwPALojvK1QHZWGWiRd3T
UMUUBG6wgw9Jr97RHw+tGGmoMVuW13AJ2yM+Bi0xHKjFbyvjYVNqI4cEC2s+fXtzOdrx4lCJUp3O
b+sQfP/KKIgcmwdpdj/2UYjW+nRKALYYOWdNVgmSgbTd+oCOZ7fcZ1s8/B/W2rvFlqGxJduBFz9F
0GI0i8JMP2tJcreTpfD/oIh5HvsAIBgWaAQl5kv6/aRFXz406tWLfb/MK39LyIW71xKN1Yqw95l1
SVgGZ+YOaN4TsMQBCLxJ54L5XF9wZLfLqtnQ+4iPlgrn1g9QGUH5PZpr7FdKKG0ft9SXZ8jsxvqX
eFcaOTEhyQRBpq/z+Orn+HEXlB2d7c/GW5iAVqUaYsAFfQr6nUsGHtrgceJVSgMapz9No85e7jLJ
m47VNWeO4TRrljLMluJGiP6Z22la9bGkNDxpl4F3OpLFgIVevRwGaNaeU7Yqv7duz1026Bvrj4k0
Xu29V9RKAob9fefyCs9sCqu/+LC8GYkNTjjURiSd4GdFVkafmSW+0b5l9E8jvD1vf/AVMNAmMRaE
6zHO4ipty/oHiifmCprrCWu5MvpGDqMayi0TuLIu2GSUKd6wMYpes8X2H7OKRIX2mvgZaAnj8oeA
ga6lY6M8gta2pV+Tv3zy49zyg5bMKwYwiHyxeSPj6zXkYh8BV8HYnd1KdwMhdYPVCzeNpg7nw0Ij
OOzkXBdNCaFxN0OvDaFuuJLA4hhYefgKLFOyqr6nUeAPcxfDBAlzjQN513WFDNy/OxjB5HOvyiVL
ILfiO0ndGXpjXCLf+1h0u668ce5aDR3b/Xbz0/N9ELRZZW0cXSQCpezjLydqths4YIOtQnBUdMQC
dX2h4lk8WmYUqyHgizXVxn0iuq+6eon51Hd4hp4KW+f/nC8NuEoHe78HLMTn+SlolHUsqqAcTsTE
HagPBgnMRuYrDeyPGwC/IxKOAY8cFHlL4mOIDPiGe2BVSZUNnYWlpw0IkLCvUkUp+l7/AlIWOTWt
yL4KXKBZt1cs/MUtYqwxvBfgRn0yt+L21U4wWe2wlbdfY8MWDIdkU81Y2zSPROSZtp6ymTJwHv/4
56juKSNOzhW01sWG9ToI0B7qMKaopDPlwMaDQomOsZ2j1syAHFkVUfV4w3nlLvQYEc/+SA61msjQ
rLlXdpLa0i9eGoX99qh3RCQOweJA6T+ZZTZXgOgd8Bqw2CTxNcW/nZuEQApjctMROBeEby5x1Dl/
fYu5wwxZN/38GitW/3EP2C5bTPca23Kdr4tuNwGpGuCUoxYBKM8TkS9Y0pLzH9sw4aj8CPa52Svb
fKNl/9DR+eWU/j0hVw/TqvkFscWozrneG3ZtF5jckshhOotnqmn/iWMGsMIg8Q/339lJv5qk8pVy
NyPUq8GIRGUMa8NbwDp2QmHYNIVczhi5AYnFpEneP2IXkBx7D4KJLfAMre/Wq/zWBMet5NX2H51M
afVFJl4HxSe/RH4i7vHVpufWYjr9ZlYMDi+iV1auEq6PU9KzbDln/w0PRkTzMR27R4KrOfiIhNcp
WKM5C6LhAqiTmsQlM2G2Gj8U5teWGRLdcG+1+i5Ifdu6iwnYQsVdzNC9QzUKIo2fangc+j0SfiD0
FyLDJXDKyv3WZn8UMUbg/+jpSDQZW6DYnaHp5yPZCh/SKOvOXUMtiDyNY3YEGlvhihzZkVn+02I/
Znldbgv6AaA+hklvvAgaKIY/ClmulYwT7vHY6uyl4h4g5Z587KhLWCrnupzRP+6rKM2uvAMmEssp
5REzdH1ETSdnKRn3OQZVaaAh/iF21WvAeSKG3EjFpXglh80XTzS6dlymW60ON1NXgHGBA7Twk6Po
PX75uvCc23vjy8Xb9OsjTwcAJYYj+1t3MU9FTgLRC/xm0mCvVBLyI+Eda9L5bLYQg0LxungLCQne
HnXj5cK3inrzhLuSye4Cw67ay3EVEhEAPKbG9UbRE04H+ICW+WnvwekWLixcUltQlluQStF+NT7a
U9QvF1SnF39oJB3c2mci5mlEZvXpXYtczrm3cFVe11spK+Ii5s+URgWc7mYXz9jmByjVfg0RuYql
DjcT2QEG5c99C+z8pziszSZRVLgIYcx5OOGe3O3AA0G5+euvH4UZwmDkoML+o8cdGz7woEm8GWWB
oTk/bV/m9dX26xpW8cFJhG0g0Uu+OciSzYc9wl8ce1+6k1PmAoUeSF65j+HQ6pKt5zK6gPOEf9fa
Rhv4iAYUjOsjVYigof+vaitObRJvajZ1FL9T7M9sZaO7Sw03i3C92z57C2SVIbBdi3TX5gmd7XWH
6agotHInlRAaXxlfUd2DICgFmexgTO0kXvFUhdMq5iA6FNUPoDcYweZv4IRGt0GAVmj9WbVeKHZP
3pyty9SKgn+EudRq4w2ezw6PlHvguiUKkIPALFAjP+eXMhrDQMHCkfJz8JJhR7qQmlVeTDVa9rM1
dflG1NF8ZlURunDUl9to4Ogp+HG/wq0LbJSIGu22/6NQiK86I7agPkFJnpmxfwQ2zyHFmLcBiF5F
4w9DA2rICsyGA+D1kPBZ0cgdDD2Vn+MMZPkYBsgpjByWnBObFZxlZF+C5jCUcxY8Y/g74bcdm/vG
kj99D2479aG3jeSzppO+wikr9jv206RqPNvnPNQ/OjhioetD7BJx3JXj4M/mFJ8jx+N9oFGxg2pO
GLVW50GBUqDPuGpZsSpWuL4nx438236bniNKbMv32Cr7NRVTHR0Py4CaUkL/XIi5x52T+Ph4PQR/
UCoX2xH7rrMUY0c54BZAh+LqHQwFuHJFjnlOSI1skfgtzCnlS3/WqxIN6Bvdh4YKSBwu5nrGQE7X
GTDpaFZdzSfabMI+hAt8yZX8Fe1/jK3y2hEEIBVZnFm4Ka0uPEC0gaSIMMJ71Z7i41h2BGyUGSKs
c/zoi2BmujOwBoFjvwz6EjfTOCxmVLv3frGrEwsISTfxOKwAxFYDPzI5ZDIaZh05qElrbMhLHhgu
SZZUHc9MrrIZbvFVN85XZMVMtbJkWZOQaJ6o5tuXzRSOX0IE6kxpbZpvh77E/q4dT29pLOZDGke1
mc9aj+RUdwuzyriwhOCO3cFjSYFwjRjyEoN2nQWL8Gph9sSHapFHzjc4haurzXsWWAqKFyrB/GDa
syywvD85OsPBZP2aT0C+yta5tXNPGsAPYZUn+5+ODez21p1r6xEmx2AD35cx6cdlgMT9m5ZLZgDC
PidnuwfFkm/NNgK7/DCzHXvRFZ67ccgjXkkYPHBVfEyflcaWgocrXa8FRzfe6ZeNITOhki/lGotP
+6bwdyfSnrOsbrL0E4hFTvdgMPnc/1XiAcumliTns3AEzSa7ELZwgEIxTHqA2kAkBms8ix6Xwj+T
uwyKZPf+K3PUdIGETdTqWCbooITnXjAsZVFXYlQXEAQrbUbYM3yB1/TFEFnNG4yjZt/6xqiK1MFd
3YZ0+Kb3q7+fTPkKstSzyz3OTNGAZT1LAHkAA/MOhZnpWf6ExL3iTf5rJqUAwR5+nbW2xZ+MFfR5
WHivENhL5FNpKYSf5s+pr2vyv3c4hxyJyh4n7c4Vh8TRwN21huUozczCpkxEdqUXKAEq1Z9ki8m8
CxhXZj8J2vovBkj+zrMYjBGEv+Ne/eDKPbpeZVOssKRfBKR0nO3fJQBPdWvvY6LjRmsxSYQ90+EB
i+HuEvzfh0BbDr27NJqiEN8PvYYGZI9z/b+G1VoCfGEwVhBq1i9IFNbgrVHSt+n6b/xNAK9SU2HT
EcQTD2E7oIGRt74AEeeIjebzg5ZgZN0N/Aw7iF5r12/9OVFvZHpq4iF+pjGb3y46i40u9dJg2KIk
tBloR7AKvdOe+HZnds+9KwuqOcSjNzXba8xAxgIvvwVYZgdPQ31rWndvzWF5cSh9l1u0YA+02iVu
diH6uvrXH2hzx/rBgKHE53EE5+gGKMFsW/smbfQnsTjw4/YaOiYNhCwqJ4h+6NLiv50YtB8NhVO6
QdJ72kPchGfSQixrkwslrLYNjp0a7xO7oqIqGD7ehV3jiUKirmk3CQYZCyLWK4pznwhz4nRudqvB
ULMNg+vzA/oRDpAv4Twr7WcN1gOuGd4XphuTYTvicHig+383a1HSbMJ6fYljnzgfbj8QR8Tz0UwB
hlj/UMvlG/qY2pBdthob3QsQnBhUIzWVQE3BEiUXAfu5nv6fgpmolZ4aUXdBMeKoiC/JWuwzfDvo
p5X1qOLh1dnfGKJHvJxwO803Ap8/DMWeK9dCdyJwR2FXCmfyd1m06fViEN9lVWiILWBNii51Rkh5
W6AZbNnXJzFtkJ1zRYjqpQ5i7hWBpYSDlGcOf+iC53xoe0vcqDqlRVzELvUUFDWocKe+duROaxVG
zjEMH25gumFnRSOTuQn9pluH1JMvesHT8W3F/nExOkXhYsyEZgaVuISyHLrQw+8meQwyc4p6U7xT
qnjFv+Fpybl9AKQqTRvzBMLWtPszsgjghzpsxkxsPULFqj3BttaFD2Y4jrnGmKDl48AnFrN9aFW2
f+FzhIiI/Utbdy99lOt9rpcQqcqhU2P4kHm+gF/n/GxhPt9AkRSwyazJ5cp3pk0jSTdc+fWy+Amk
eAetIiPUnF/XYTp/+CvHgqH1AeLS/QOApS5R9JZmqvcbl/ZrsOICJaM8H/ssKYYu27GPSYpie24Y
3VgYmwcRCAyrM6LiTuJXn6Dh/vzOHYTkzWeJ0NOG695Txu6MTTbre8OK/iFLu6R4MhvlIpGS1EHl
IBJhsh00M/L7RpktcKcFA/7+xlfIVHRYe5xD4il68GKP2M7NKfcMxnZTsL3grfWEVh1bWhR4hcVH
2AKEJ80lpjg6YSt+1rfYnJt2KaRQHYyfKxpIEbMh2kkBfWfLHQhL+IrrrgRv3HSv7gSXhSFnQZQF
xxJtEl7Vu6UYY9wRB2VEHoi6qlVwVMrDLeKdbTQO/WONJfuOzjtI9wV0N6F5W42j22D/s1zR9yo/
fjaDrnRs9wYMpgJjHCiOAbhfLCCcn/yRrmj0p5Qbtvxo7/aQOb2SxHHHLwrKpnYGCjJzyJfE+r36
WWEG5pa/61PjInRQCTAoR6wGtNM/AdA2Jg6HMh5R07Tjd5xVBqVxfVxGzA90qaOvYYZjEY7NXP+D
Qia136NovXGjo+QytIcZfXcdjP5uPv68MpbknAk+YRixsUN/+nmeUdX7tpbdGfNt5p2IwA+Z/Mf6
d3Bn7sBegbi/+0k4U7rjBNFfSVLuSmPTi/DPDvdzpid5C3tmdq76lODU8nAPS4WD2Qr2/ostuqRR
WTld99Nvy+WX38hQClNc9AtK1DRRIZWaS+WcG/rc5PEn2Umj5MZ+hf+N4Yett8UvYzACS9vjoMcC
Ocj4vmv0ioXtRj9xoJ+d6bBJDilH1UzW3PHpLKJ5Icf/9BI6br8bNnpGiKPr9qqkPLALLfWKguZU
9xzZTTD77m2fj6D6MOnsL/8Tibv8JObmI9wZBNcumNzuG/rd/i/uUXqk9Q2fSvG+jSoTNjCkgRn6
Q11gFTaypEPwimAWFwSrDBV66xpXKx3W173mAOmxKhZjzU8oZZ6AcPyhaWJCUbTjxpBtvRJUxkXQ
EFkgz1SYk/ZQZJpECFsVl2/ZDP8FeQuFxxnZFQZUkjV7EKMUvnr5A8ym+mfB0I7+QgV0vFeubJc2
XTz/ZvljOhudZWRCb9VvcRE4qgqlY8aoefge/fb+XH6vfFUlWJWxLMwULdsrQCYkwRz3ucG4urBY
zFXoMn7o8PSdM0yHWVCGyquN4ZRwKAk6R1vn7jaAIoJGD41rze7NASkm52dh0yFCbAY9a+NVD+OR
YSyJRv27qXII91WgDnuPL+Z7prRQUfNfLz0G0UsnTZNYH0XGMp2in4SCPB9XL1QbAmTb8yKFxrSk
myj//j1ELXcfbXhg6bGekFP94xvMeQsVjZl71QOzw5ixmIsjCwYPTwrE8zbgdr7Pk96M/W8S21Da
1zXy4bMiPIMOkpklHXkHm4tMKCXllpgHfdFVh4z8PAz81PuL/+R6t4gbgjU1QbMHhSXJhxsF0lSE
Wsd16VxRZy6nmsUph0YIXM+jQr27VTFeS8yYxxwTccnvkOQRdpJn8bRJN21Noh6YSjBTaedL6XEz
7YWRxW40Po7Rc/AMVqUyd6jQFlC15p8uZWL3d58wCRnOIh5qHCqA30CqkcRlAxlKZQC8sBeCOjwl
Lr7FSXt95TM9aDftQIJO3geymSkBZDAm5XerOBOzH/qV5lQW//3Wbd9zY7Ma5q/l7GVEomZc2Es/
FecXVaLNsvCnvvNqxSoV+8PJIjOD0R/m9Jr4z+Umqz227/zOFYPG/As0c2Y8nCx8tG2zldIpB/aE
czeCG1WDq1Li/Tll9DLP9gjw+7n0PrHoBhkPjbtlT/PJV05wnbLzgrV46kX6qVlLpD265G3rjW34
TOy1mcfwmv3EFzygXUcQC4+NC2m0dMcXh7VAraX5Mt0VTbfj5gWtEc/FDfDhmtk6ZoC4BysrL9xv
efAfKwCpCHVFbZkbD/n6UkJxNVUWIoEyKYWmOXfp34BaVP4b36h9BsifbDl+9hsjAwrgarfw8isF
kIy9SXZ5mufuBT68pkH9LpTm18U3eg1P/cgr/w2bdCEXYpTA2yH/exNt0Dk55OPlb5cq7YJg53YU
MK9V+Btym7bDSehr6bcsZcZbPXf/DdZC8o4gNQ4aKHB5eYoG8c1uQA3GE/ZqDRg1l8GAaK93iFC5
Y+jSOwnXobaZ4ZlGACoz2ZqZfpzwCmaGzdP1Jw9NTvatXHTEWzm9UlT50EYJuF/Bq6BwwpOw3jcT
+DQpDM2bxgR14i28BtVUr+OARBnPgTwYV4mrCr6MR/SmvOF622S0RtqeR7oeC1LOz3cp+Kk0ymNY
LVYvQ6Vf9Q4ov1YPd8L6DweOAHxdrQjbJNCM79uLPbQ4J4uUN0/7Qq4QZMGWaZgV7+sSu4Rugc+0
3LaT5McoDzW207EaDHUskIB8d1706pRTvDQWlcs/JYyTclER4T6EwdWydC+PSkUBo02oozyKk/VM
qm/lALtiSj+UxNfFwd8sVdhjQ08Aj2pta0UXXSCH66eTYqRxjKLerLcS01fNtAw5MlT0tTv8Ij7b
UN8SKn3wcENMzSN2XTpeOWUKn6UDXxYFhP5pC9nKQDTbwXcv2OBbHhO4bm5FcgothBuWwgKpKbfx
ejY8Ro8HM1ciQ1nMpTzeqZOMt45EM8oXTseWmQPSK8heY7bI1f3gmDtiM1wKLNmsTh8Yydyyv6Tg
9LlQBFfXR1EI+/LtuprPx6LkanV582y9l9Sgt3yMPG8vF5gkpPL+f2EYWWtHb8nzEcsxLqHpU/4t
VrLZXeg2W+ij4lenNTrohN4hd2LfWc5j3YWvRGOvCXtxuOtD3IGe4hB9gzlwCs5VYUAzO4Vyx4UK
TXwybZQU+HySLV08wEyPBIKKjESR7b3IrTmWgACnH0kbepuaOd5CN3z85c/aV5k/qbMnaMuGigck
dU+msaqbRc762lae+iifU7KFH2yPLa6CbXnQ1XgrO+gKhKzrKogZRjqrgsXqCCzr2T61QPY5MMcl
0XiTTGFT8SggvEPKAwmBPCy0ZPvTUnxvh8b8aAHW8Z3MgdRHDTsdSaUgtOkY3D9rjUj1picIWuZB
1o5bG6ONRJf5rmAhGpIRWRKnTvN4jiICwq7aN/Tm+1edRYCJs+4k9ab372uJgh1UINkFL6qhK+DO
BMxkqjC7igomOkorFYUM9JeMlDbhoysH+vp4K//L2czrcTGCKsGj5U2rh5b1oOM0u4Yip34UP+FO
f2wNTATc2t047kWOB6cq6WwCIiIU+mHjXGiRzggcYjL5P2KzXyoU5cNGWNJWQrYTIsJQXiSPyZdn
h3fUZYUVMWXaoPMei8amJ+VyyoD1yG9YaKBZMhPuePo/7jmTek+pvCkfjnMqwx9H7+fH35T+pzKX
aMYvMpPbQtrUuBD4HxbRMy1cxxLqA8vlP7ZvXAkirrj0YzTAtQYioDZ3c53oeRUHB1YMtyMSM8h3
8eCni78PBgosC9jzU1vB19f2q5Y8hTxsMmYgJPdSApJHnbp/T7Ki1ESRfalMLm1FeqqKXEo0i2/Y
ckNNnLr1oKJStlQa4NBgTdvcIiIDfVGnXJbtf418Yojqh+fYTaL7yi7cYDlJk/YWlAFo7Fr03REL
r2u1UB0baVbqKwKFKsp8RyxJYMuUEZzT6Cf3L9mLnq3iXR4v1K7YS0q0ncVqjpozqeOjfnczyVMq
RMYttkOEOD2ubSwcWDPZ9k51Ak9jJ1Phy6ARpcXFEfCYfCF8tDw4Fmafy2EzE74q0KuGBwLd/mBL
6fB8nK202ea7cMI64P9V2SfvgJDQDqFmlSHea+1/k4ztK3gFUNbrUruxvjjZyJz4R5ssm2gKDl9k
uGvlRTrWZBDe874mXxsnabuFvZa9+PIOvmTzzJaP06sTx4IZAnpa1tboA/ewQm7I2e3F/BPipu8N
lAy2AVg4B46xMSa5DEexL56A8EHvVxXGcVKyo5vp66+SHWFOBjadD1vFV5L4W7BApJGvxPiz+lmN
qVMK+A1O7JxZvG/9GhnHhUKg0AGxswuxPaMMe7K1fMY+hhFkpAOkEfvyfMjMfEw9nVA6QJpuQXFW
+oPoDr2IHS4oe8C7DcV+/RMd26Z//uaDPBqGDZQ9MW974KaIhp0UPfjYBN6OqnuFTfqitq+PjDJe
PtFXNStkCACaMVsBw4zBjoGRqkbj5TvQC/N+xbpbfrYbBVnQSN74w+gZXvmZOthezlq1y+bn24id
aeKM5dHHKrazRAY+Se/GWHLh/CJvbL2wIvZHxWYnf30hymNOpeqhANcdKMtev9LfCOMCSDATtSs/
jMjP/gjge5k0ryVLzmnWXU9Z4RVtwqoXDcMRU4uFBjXfzjld1XqgZV9srfEDfzrY7rx9EFe5Xhjs
1QlzdNHNm+zXfFHuf6VDNAIkPynvrdOjQgyzNb9D1wMAJNGsm7QaKUFY2wda+//pYv7bORvBn42j
b3nSGX8z6Xj3X+wBk9rowYuDUSDy194EezpIu4mRbxKp7zW9xpwFK2zK9s4vbVo+oLZPPhlq1sPf
Ly8YknvJ364K4+9BN5Ndpv9UTetufPdR364jDex6deM5s9cejJjfX5hmymBYqrCxo7xb9wwnQq0X
MSSObcjVvP26i/Z4kP0xCQDLFiLaGNkcoKF2TejdpYwy3Gqj/21rhzDl83Y5vCmydDVgS7SA5y+E
cewm0hrvISVse5oBin5tAzHnpwEQyWMcBkX6GgICJHIqeRl4+/8ns+WYIXRRsGtj2oU2E5e5PsDo
8MQHbLIvpyEDXy2K1dIVNdNIsyO21l6j6g//hrIkZNPa3+xHSEZPKTl+cxz1lB+ekg+UE/DcsZhh
5nqpSo63uL0KFibBjU1FJHVgtY/U8l1HT2bVAWJAuFBPb75PWYCt6em7jdWRgt18PyMLyeeie+Un
M0K940hnIrLL7GpyEcJvy1W4mjOnb0QLLGPZQ2Xlwh3EPbIUymqLcuP68FYv/6uJjPP+GUVKV4yD
O6koyEYPuz0BJ+CtI+yhDXsw4GQzChj5KNPmQRCJkIAPI+00zuAxuMXvknEaeb+iIO2mifAIIGZ7
ukbGYjRsSJmqyVgFt8InoKkTLmUKfpfV6DxZJijZYdZuKlCN0YJ+OVYfzSVl1cXo7TA5lp2qOjLm
Ete46IcEhqlmwk4mTtLS+xBp+H/TEmhQlemxibp/7/rAI8aDQBuNcUSZyNgsYw66lRxHyYOFPbYK
GXmuxufIzkorDXuNUa8OtadnO+nUb6qa76AqZ1x/A5Cmw18mNv+P5raHbVVrGHrCK4EFr2mQ3+lx
5WFD1GTcluSDu6u9De4KTlgLFQFeicjwO8HEmCIljOi60R3Blb3uz3xIfBGsyfOJqzhF4F0SPcfm
40nrpzeAfi0s0egAzhTCLJwqRKrbjo71bFgFHjgePH418HDcFdWdxueNUSWC7JRyPBUdNQMWvWqx
sFrxolqZ8BDeMGI+qIqoAr7j5KR43EJtcHvNtYrHtUSNh27x1xmAAIhateHmi3ZwszwWLeHdCBtI
MvoG3eyVdz7X/aOgP7qY3nVFbOEMZK8w1d1NQyTWEyOHofODjLsBtYusqg9edQ22zpwtj4MoG/9p
lrURDZj7TP0JxzMqJAXr3F1QXtnY/jvEGKthTCrv3ZfoDsJcl66qmsR7jPfWK0TVpo7eXqcUfICW
fHO1TrHQJC05OKgYULN5ONcrvht01VGeHYxj3H7REDU4fvB0Zy0nLDMX+7f9m6QV8pvYd+ZE/ZAo
2NGeOu4746KNiLQ8zZ+wzI6t8b5ZuyGmmdB72PGmN8q8rntgCwJE/Hb1+RJ+c6eljjMdIWaRJaXu
tzPUgLiIowF6Y8sgLaRGqbOwolEUVUWZTXh7gRQd7YdE7NoyTYL29P4drMLLbGThRnCFJ6TJX4ir
8RgdZYeMHgkeIucLLqcFPbMeqAlPua4uIOHOc3y8rJqzxHjt28zwxGDNe9R0i1SZGhjCsUEnbzbv
HO5xMRb+Ogd5sFQXAorHI1FtXcydnsLQJ3qH0l2gpKzXRokaod3V4I8jG+62R6a1IAv9hAe0hgxM
dJNJCDtprkAXyn1V4r/V563SVSmh71U41qGUGkpqtxcZZ3qznTN5Jps0rsBK+ZExhwCIgfp8Dlls
3C0A6wzhNZcXWdToTSv8rMjWnZAy4SvF3gs1MfL0v1dHp6pMaelVbI9BZSCWej1t0aCRdrgQ3JK6
IpRFxlVi9M3/oUzDHaQaei32qf3DGfR4iS44i2EEAp7bC+Q+Y6LNcTkWGkqW9C7b7i8xVhlDUOEj
n8PT9fNcJGY7g0/kAwawqYygitlBoLECsOzGwHqRnCqbzK6sxF54axmQVvvMfUszH9oLw55wPIGz
8FlXw8WHKWgIzpStkle60SxW5eh0QK9vSjb2ntkyuWbdrMVAzjVhf3xUHV1ktsBd/4TaFfCUBB0Z
PbIPFJDMzffZL8XL/s+tzL3nAoZTS1wmzsHZ1BhmF0kwfaWvOuow38D6D104pf1XuRlJb3G/L6oI
PURnct9FQnqAAq6jLxKHNhjUyrUY1BdAKN5ZO67YmJ9auEUN5mO/hg7B+de9yIh4nzkXNRqompjn
kper0VQSQnANt05McjWOTf1OdGDReU5uo+IMzuXjpzwqyqZ/ANQMVSq/p7G2JwAEU4SLgtBzYFZ7
nXBCLwYf3h49j10zze7pukd0MK+fIFn2Xxee2u8AQlIEJNynCG1AcB//Ks6EyVm1OJ1FJQ3YcIjf
0FAZRq1t13K0ckp52qXtPbhcw4XlaZSNxDmSLkTfrwY7pyzyO1X12g9CMB5zbtGsd4kUMWGJiBJw
7HxFEqPDkaTq3ewbAAlc0ALnTrVNPT8yGGVAdGLvuYvYipJMB875hJbtA6Viy6yPm/wRZyB+0C81
+apJ62c3qxXCM/M2HqB1UcvPVlAeQA4FomBT0NUFlH5mqLHifyW5H7CQixdHymHPB8YPX8q+RQYK
/2E9aH6zS3wXLEQTBtXySN72QXtI0J+51f7Y9ATPu5Tob2U0NhRq63jPLhRv/EnaQ7nTxYQsQ9pE
1hictY8zNKgcZJI5hL7Pr9kGwvxK8Vh+xqu1izS+FRbJQgysD1EcD8kMbmR1hW5swI8gu8al8SeR
rQCRW047t2+Y63ofTlxtws0SqLgOZI77HXZ3BnjCOYiRRo5WMK6NNg8GhAWeOzHCmQLzJsbCrieS
0uw7cwAugof5+ON+6TFRNXc9RfwjlFEN/C9fKI9u458d8DpBmH/+a7oagyF7+kKgm+17jnNk+i8g
iZzMuo9HXxq4Tr9gvekQjT4dtOgnWKJPk6dInG/qnuL1LLdiINtzJTBAnQfZbaa6uCrZSVhLnemr
WmmzEFoT0KXBym7Tz37/0rd+nLJ/9fXb8JXb8V5Y/ixgLl3BTHiM6eaZ21oDzAbyivVzsgmFbPGn
W0+kKkD5osKLggDrSqMzjdXJltLt74HBDLs37h1lq9ZpB5fHFzM0/ux70Tfr8ha50w9d9sRaCn0T
+qmuUfTOfxoIaqKZLCCp3STNufQmsJKEGVLFnALwAhnn6vdqaJh9ueOCF8RyU3HeZ/yRXALRyfCF
RZ9LJlEYFO0vOIzl4UVkXAJ5inKrNIbept/kYxrfgxTRqz7X24xoJ464kfhyup7HielS3Sozk+K9
eG9UgZlQMi6+35RZptJXH/70ygXB4wJ1HngJs53n27IGWN9HG9JIFtteb87k24e4int5LR8oAWh4
sAYRS75JjJet9MYZKkI7+uJChy4zpXwVebr3LzsVRUl13sQ+BQC1qkBtbfLXO7DAtaPZ4sUqtJqt
vdTEFuLecGVI1MWf9HumVZb1g2QT+X0Dum/xgkN3GuIlvxYHaHmfPUicZ56fDy6TrQe/eMgL0fOX
6nKvXYOVAQUCXT2qx3oXKPh7/UYS2ryGmhrFpte6yhI5Mpnhs5vcVgvpYJ9q2QGiET1CQojC0iHw
5PO4+P931m70RFZgjybKq9qxZUH7t1PQFkv94IzMU9UfwhvcYVuGas88HGiLGHNrvvQAG6ZgQKt4
OCtd/JIRxySRPtPq8iGsTeWalNvIMkbgSRzcjjcqQPgUUfhpnCYNqua8XESsSUY4LChy5uNcb/dx
So3VHXpBF/yhMnT/OHUl1YU1Z/8cthBPqTCNYJ7XglCM+g1M2/CWG6fqofNP2qYlW9ZOjdYGoc6N
LDAOjeMizyJqktNtqeofCIQqqNF3WqM8JL1we19gwVcxQhVLbpU+3wPRvwhOPKEOkMDRgekQNLPx
ZEfX7pr1nB4VrTexyZSZSpqMvYa0TLvgl/gpcQ62gncNBDFp2vUcHTFyY5IuHO4fGplGBdG2Ijjj
J3ybaoYRoSFKVJjTAXuetR60Grq30TPqd/lkg/Xw8Sd0+GKsKDurC4zNn/bX0ON+N6emhCY3IHEK
64YBPgkN/N4hbqoyXC85g6C29a3XUGCvi9K97bJT1FzwvUU6RxXsxK9TCoX9g4hYFht90mpW/Ls6
14cZxpJiCt5AoVHRrJjReQ7tx4QfD9j0VtBNaTnWVMgiPwTv2IfBsIYt/DV6XbqoMVH5PDu/FQQi
Wn7z42shrmEcAZKTZKPLOmjcV8Ox2Z/8pgYo32MHHNpkfxf2pJ5xSXSp6jfyBtz8FAy2zoo9ZuNU
wKQxj8mxx076NQUv9S2Kt+7uNdVncLat0UV/FiB0FcH6i0K1o4gRJ0xo8HigGpDRV32ZWmlMNqTY
Bk53Dv8jUQ62HSV+P4JycwtqM9V3B3CEKAM1NHkC4o09vb9bhf5PXPWZkaVMSpjGfJP/Mc3aencD
KRLybp2wRuxOxU3U1cQE6wu5EbdDZ+IJxsVkhmPDkkidY8c+1McXa2MsYxFs3njHw6ZId31uQ+XF
BA8N0yPamT1e8Xs7Qfn7NEpMH3I5xM35hdPxYlPz/enHjhf2ql1akAGdjjxC2Q7LCBbCntvkZdkL
zAkTFSQf94u03+RHatQW23Te6O9JD3D0tSffBnI7OVG8Wpt4IlMBWhQobTCIx1isUZJA0PQ7L0pM
3sMmpGqXsIt9pC4omTEYHYUDpgiCLgrd6oTPHVlufy3YStANEhxvLPcgWIJBJ2c+0UV9Q1nfdLeP
us6Tb260ibLf46nHZNZbkzfWTmBt91a1npv4fSEPA+ZQN3KNYHG7lZVSVdxzxhtZ3VYP9/pymCuU
5v+A9SoxP83H67xWCMJ84BOv3MCh6qWZf81tAi/lO+22XTXz+h8B+SxIN7OQOfSiUgV19d5/TXw4
hViPACyPpiSrs1xd2zRjLSSuq0CdUOIqGh4sYLe+AE33PE0lgBJcalaJCerf89lbFwIgLd+jj/8v
6qTdJ7IGx3VadCND7d0QNCvmW12mcxFp2iW5PaDxB2jHRXvpUzIT5kxvuBCnPyPu8t/i/5j9/IYY
b3E66tEpAccxt+tR0z1pi/IzHMegZqRaqqf0waH25MmQ+VGx1Mgni45h9eRHcFGgKjNPzSsSveoN
iZ9pbS9Ypw98Ip6LJMx4ysa8poIoi+S1fHbYQU4djV5sJtykVRe+z1QLeloHgc6BtcLXh2Gb4k/X
0BRkZjKHvCLfNcfCO/0a9lSFPhWNMmjqU94jpTT3tgJXq/20ZsHBhxmC0FBPSVMwGpXaaJrz31Fh
OkZFbJFFLL20kuDV5OX2y12HNUqVmIFpWyoC2IzxYjakafjl9n9usWxb2SbMvjA88+Dphi4UDSKN
qQIPgG/wqM8TD7nqYlVXbatyGQwJVtOJWEkF7sdQe9WJ8o4X8CwKg2WcD7v6ZTzYW6+joALhMrH5
GvPP7NtGrangIje7uZd3RrAZRG8wQVesW3py7A/uI+z8iLjUePzcTw2KfvCSoMjA2iw/+SUTCSIN
ZV5VGUbbBf5Fl824GxK4jIgNQWuCiElg/XRHMyR76iLZgrNQSvlQsBz4uUHdSEnsV+cv8vR8N09V
VcAIDMxCf/Df/wbk6YLxiK+EyPTmqvz2qgOCnpPXE251Guizaoiqr/n+eI7z8v5LrXwUL3tbVlO2
1hh7vvigoclEXSnd6cCp7qHvdfqSE18x4qUo6fqhc2uvvKzzZJ4ZP0y9QCDDhirke8dLgZh5ohb+
mwftubzaZ79iksYSmEWORu98JfkbC2ea+UnEW9Qo5LjgPrZNV5feyhJLfCKcuMa4CsEF6X2sAK4D
V0H8mw7qcYO94+qWYntKzlkSTRcNQKr9aCImKoA8bYH0vJlZ5569Y/nsuoGMIgj4e+8c66CAPvrm
HGPNrhTnlCT4JJ0Oh29Hy64HIzC9JD4e+DL1TE8Vtm8t2FzDVl1sOq8do5xXn0S1eYCE0v8TslJB
rw5mN6g4OKLqf1FFw4Pj0pMsIjIJERaUsLiGvsuu6HnPcLBhZT/xhZkLg1fIfSntGsLMBvP92w5I
u/mLE4HekiYsmXBd5tw//yJ8OgggJ4de92nxhHl6Ib1WTWHho5eZA5nsbHHRyzsgkf8mJ0WrGvxh
OvWZk21sBqCH4l4jup2UW6laVc4JDPV55Q42Wx55/LzE9Eo4ov45QHv8S4cjSqlpY+BF1C5YBvqn
Keti6OLLhYgRtPggRU1QFTjPRDdIpsjk/pStwNxwLOQcPZ8+lO99eQQPLADWGhp0kH4WEWt4ACfk
ut7Ui4BlPeGgAGi5lNc/9hY0rLkLTZ/GUzJvU8Ad2tFsQ9QhDkFExUESbyh0dVH5AtH9cdBEKMsJ
Wa2dIZde9Kf+cjWXxEYyy4oHRO4GTJ80C52uMn8ksLGKWaj2kP1tBar5VYGJjsIt7WkvEzAbn5cf
TwKYrCoLZG+6C9Z4QyS1PFiansdfo9EyAGyO1pszfdAPuPCNgQ9+Oix7OY2eLMHOAT4Vi+7hr2go
yYcOebDIcSInN3VgcniSZL65WfG5YE/0Aj/WGzezOzwnUicFdFgfT1ix3yRIv9N8Ddv62Jng4kq1
Bo/vOA6eIkmAJGH2LiTX6aBGdHeuTGiGsHedgD2iU6ZkMuiAmk9WlTRsNjGL95iggHDfq8XajVYe
Yi7IUeGU7BeLnI+Ay9fqF1jUEaGSkE5F+iXs6jhDXe+eZ9oXkcOZ5esQf+7De4cmlFzLaXwMYb7z
O+njFbR3gQyFyzbmzQEdOU3fXMI6ydYcHUnYHEU7ozaEGXgC5ZTezqEwRpYZAevua5dPypMIS82v
9EyO0A4bIo3C2Pay2hNlebmX3idJYYKcNdnj0PpzVnSDX4bcjh1y3vW6XmrI5D2zFa5MESXJ/HXb
Lmei/URIG7sXJGeQ8p8boDdr05nnGbaR6jUVANW5rvAHbng4fSvg8tH4CwauBLU3uEhPQ3UFA2Kr
VdfYNBTVgns7haplguO4lHW8+ce2AUzGivzljeCgiV+rLfmYqiUVWgaWs3BU1+2xw7iU5y8pXQpM
GGwd9SjfKUso/jq5oBHD8Lekw10LFKHCBJJmsVlYQLfOs3LvIT/eZVABiwK43hsUUxrtWCjJv9As
JRb3Xi1VPJZD+fJb+AcsXOgqMKhFg40cUkxag8eXLfSQoGWKv2RTarqxsFD+Tbeuf7S+j2kaoS1v
CBfPFaoI58tkc6Bcuh+hve5pDWE9suwk4v/CoItopeexFynCEkWBh6g+aJD43US9YeXNbetNAVkf
g7la9a5fCVMuJHxkAfQ87hssLhJ7i4tE6uH3rcUFEnKUn45rNw+bCaAnnXGYbTrEp6Ushpj6/9/0
FmguYvyFzxR2A2x63fax9H9NIp0UEw0HY66VuCdQNsGhrmKxU1mJ2Z6O69Kh1b/1KhNdq79uatF3
TrMq+PQHwTuKLVe4+tQBA7v5A8KRq4mjZ4jV6jbMUcsXWsQ8NjxccyDep8rurPOAYo57UuJ1kgm8
N7iqB94q+2ptuZ1MnHcCzLtwwGHXuowk6yCUFTZYiexZ8bu/GKFZzdCy+fjLBKWBgpLCmJ8bk3Uh
emGb4F46TyqenHHsIfyicJHQbciJI4pGAwo+7CARYUICaH+htFDhldp69gD8uyBthoGmoCp1OefK
LQmF5TucUzBkKlIrtjHuQPRQ9LAu8+DaIn5lsQ3359VrThjcJjbXCP4mZQkDxeFDKGozICcvqrUh
PbBfGdVfDHTUZZzpsjRcoJE358rz4rDVcqLL2mD6JL5ggK0bBufmtrNv7l+qH6SgPaC5nUC4fkS0
0WY7fDSP53bjAutL8JO/Y2ircdvfwynRMTN2klUto4uFID04+50qTZTEfWA1mwiQOnSHnxuwCZ/A
DfbZLCveDTMiUKFppvRaNHVDjy3F5fjzir3eXUnEEoJySvXQJ83BzSC0uhP1ym9QY01Yg/wG4oBR
E1AAZHjt/aQbJ1cu9UxuBRSq73QvVHKrl9W/dd0Sj+vqJwDGCEMQZ4LJaLnDalNUaTw6Clb11X/E
NzTQle7Bp91XbryZSOzoz/cJICRCVyv18ZdtA574zDkLw+O7BbD7c4SKOUtB3zsZeq/PjLzV44Dl
aZY7yYvoCQpDIF2ZVBiGohilsmeHGKCjTrYTnKloZU1GsKXL8sprzY1EiyulXadwDneFRBPJQnuI
jxQreAtf3qdoVvt0SY9rskbsyM9GSBO8pzzEmTkLjBKkczvBc4eiYb0gTf1VLSSc196oxXA9BG4O
SH6GUe4J3/wJ4ADDAolb/PFYC86JltsTvmiTg4KZ8amboyB6Lddp2BVsHt3J0R3Gln8VyLZysliB
siLUZ14raz7wyn75KFaHHsSyaW8r6hGCTqgM3krvecOpC+p2csLDhjXro72MYL2AvbtPOkL9ZBBs
93tGqPdniHkn8Xaq6H8ZGDrfbi89sZMRlQQNxxWhs13cUhAD9kblE+UcRq5uLFwWXSfUPuWh8vN6
TJN4z+TNObyAuYL0hBGbjfwbTWv6wqskWkidmslWPwnuXmuEsmPC9X8Tm+aYQrh07V09pmr2x6bM
pJRfUGcbiN5I6hplOtR5k9VU/eJLrcxbV1VG5l4ADou6PQGIKYlOIhON18JhoJ5X17RkEJoNPnSj
Y1b+uEPUcWvio8ekxpsrzxscK32uFAcj1VhwKf7gDoep05ebzKrxb0P4oS8m+Z+p9W+R6Wj06z8B
HlhPfI+3KW256q0g8hDSZtA4FhHtlRoFtkjUF4ohewVfT1ak0TDUvpNYmzMUzbhTr71KUzUZY1MF
+NVwPtfNf0On27hqEKs8G0/1r7nhiBGWdkZFwjCY3cTfDpBj/NOPtt8cGC1XtU4aag9NGzh0VH7C
ndIbkUZ06LZkcs/JNGnndSET+i4qOpzBtMvsZ4spfqBzld6CGVIVO8GFSEhiRwjkrDUxWDZpE1+y
TxCdCtCPpvONil1ejNzDswriuGrkCASS4Ewtxkt+rLR3In5G4HfZY4ksXNFmb6sK7a13dM/kehV6
FoXXHL/GVDhXR0Y2r9wV+Z8v7g0iDn3u/SDjpREozAVZp6NWOgsykJckBirYW+2Ymz64tMCHM/eV
icTUY2Mjmd4whZB36Z6DgDmkXy8cbK8KmUc552siLG/2X711gFRaC96SGHJjkGV8nHlUaNptHrBS
cRqmC8LBIBkm8n51OL5ohYMj74OPnnGH0lWrI10mlejn4eRV06v8+1Rmaa2DqFFgcQuYq7zBgomU
hEeM6v/dByvs6kgRz7oExaCZTrEw/aGhBJIMq3xP/IxSAaGmdPduWQfeCfMlnYrkyCFZNTrfao18
0h4gwT8cel2tbyAd1paA6KWQu+aRx4rK0VjLFi0i/sEQa/lYFk5DriEonJSOFxPH7AB20U+TFkEY
EFtBXs7bpRukoq5w8vWasV1M/mTOJuzTojhTyMu1VZEhGlWYoly46/wR1fNqR8FVWXQeiptRyz5N
hatTeKtVnc4PdCEZU/1fHY05j+O5Ux2hqhA9Lqf7FWefVHKo+yjqdyuc5GE0NNv63KDEQFO0hNJz
e2rnrPj+1e9sT7VEYpkl9wyRBnN5nSzkhEMipgARMGZR9mduiOIAd8cLfIXrwfnI5PZeqvISt0Fx
pJumuzKZtxYzeq0t/41pgB2q17gcsSky4A4YC3MquMc5aqNollDE4F7B+RWhCldHW9s+PGAxEm2u
gyADFJMHy52rEVLcdkVrvDd+hxJH4RvilUUigb5sFjXy8CDnhKXBZ1X8cYyIMaD5N7qeCRrFc7W5
/tcRygndHjtAPx0A9xUIC+0nUHhJywqxfN9j6HgTWUep78D/xcLJe9kSDcJxQYgyIKo9QzvKs9J6
BV49LykDFUCP3+v4XXiHip+aCAkDrZZaplB630UbVinWimejUCfaAMOuN+/ehnST6HeDj7MuTJys
ovvrjLUC2b0jsKrSqBnbsshgzHR1gE7UYPDveQEqee+e+2laCYofVuPRnSmEX/2yCgHf17TyyBiE
gXc39oSi0NzhChwSF07grlSpmxfLmBAycWhHbP3J45nqkwxa6Y1b1LJpYk6jgadX+T8cczNMWLEo
XlXNS3JaWZjNaRjcdjJkNZ689a23dbm5Way4G3m4BOgSe+a7qDSWDipkUYlfbtLMCSrnW342GNPL
zll9MgyqQdV08qrr6KemWYQmDxjRbD2stO6bv8v4/9Y/VhnjTdVZASOJ5qrestHTGpBgvteP3BLX
zjttfhGTX1wjCdiGytm1wga7qlsy2sMIUExWDeCl5qzDju8l2eMIHdG3w4vl0jVJ/egPLS6UXMEo
fcrAy5Qz37Cw1CXan9CoqJN/eUu6Wl8k6I8IC8VDABexSE71HP8CXC86rB3mbh5ecwUwic4sH3PY
pVnOnbYD/sLciyXL1ci/eriBlDJfaaPb0/jqld/SyazzL1ZikCq7wcaGfSADANdMtLSzThqa0x3W
y9VKOd0bKlLBGRJgJJet2J4t5pyt9vpuQ5lrLdu3RDDnmqmnuK763YLISv448SL3j8j42sEWgSS0
sYIsXypng3SrlHnMn/n4eD7BxpCtRE9wKSUDslGNt9trJeEhqkdMyYNDxmf/Ss0nGjf/yb/mEj78
eoIbz7PPX7/xhYKmxB+34nOUZg8f2knUMIQy7C3qHL3sz5iaO3aWAXq9K/e/jH7jRguDNyewF/a7
fXdfQ1TcQSZeV3yVujA0kcOmvolAa7UGCQXEcLPBQhjUs6BpkGIzS1tewmP8Mg9Mo+DOrVhRCDB5
MJZ+gkSAkdJMgbr68SEUe0kQnfvXhGOHnonCexsqCpbm/SrB/yjI7SKUT0xdv1gBWGDw2Ldct0W6
8V2vN2oMuaJ98tvYrVzPi7uGMFqi3iJCYk8uA41hjSXLpWIsUW6eq2JgOUYkHn7r/DmaE6DudFIt
DL4VJV8qIM7Ar+684m27EL5ENy/sMir5iuLOQ4mUdOl6pTqZuuV/hTwzvo8kR9ar7k6UXB/sGT1e
0kf0LX7HYtlH/hJhftgwHsBbbVu+UECEcpi5TJ2aTNUkEYd6hIa6PNf8ig4gX0bYiygfnWDyRAdo
BBLP4IaQSYtk6d0XdQtU/NdxplQQyV4PDPLtICM6+ydPaztC8fISOfqdpkFfq7LIGV7AZGP+GqMm
++pnT3ZzzPT/9n42/JVZFKiTLgZ9zah/G506f5V1ofg9sH0A7DiSgQg1Vz97dnnXhyDTkHaxNqX5
dDhga0GRhxPmiQWhb+DI+vDvxk9l8vDNvp3b5Gt56AijoCLGfgHR6M2ca3DKp/Qf11A0ZZgFOXQq
YWiTnUIyn7uHZeaW3aoN7AjrttSh1CkTQsRXwuBdfpEkZpxQ4qUqh46DByPTIwJFbDfraw2X4Zc0
r81FUcU/lRx24S3D51t16DIN6tpDWyJjr4on4qStf2fruZjoCpFNLqP09UPpkhkUfg4MdDjrQPN4
LL5dOtlR+pcU7x1eF1LfY+zVGlKc5woMRuBRlChFUeEfZk65VJzLB9F9StiUk5VL0xjqJ/6oxo5t
r2IkfFoT1rX8ifsXZZiiF8TToBuV2WBwuS0JtIL5LkSM6Ki0O/9OKwbJXpKiE/34G5uIBS1HF+KC
CxQvVUUYs20x1hlopXZ9EU4/aCTWC3s0jU6yviQeWFn/3LJ2dYP76qKFiwcSjDdRNFELiCYMvxa4
6Nmr7u58+cVvdROvfeBucULPsX/Ffqi2YkXutkjJd1C4grm1kU6BGGNQzqbEneXgfc/0YWXRE2M2
Q73oGUGM9gLVZW2fatuVOZxe5Qd8x1z0PEVQwqb9T8nhap8uyDrHyYYJj94f2RUphQ67U9kgs7pf
F/GvCyMUIAL/NfpOqiI/Ia3KaWadAsLSrLh17j1KNrZpEArPVgsPfodcVE2hURYuJDntQIUoJ1qk
1UnEFSrYDHylxNcB0wqEpk0eCH+nb4oRKzcYgoCG88P9BIAtkckm7hmTv1FY5DzxFTfM1Jxz62LL
rEZlpqA8hW4OelXvbzOZ7A0oMkU4/4VAyHwXpQjoycDFfyLWVAkWHAEzDpe9klVA1Pls6UJmUkaW
pYywZfHy7zeccwPhw5qiEihRBdtyVXHCHbWpgA5x+FegQIHzdxsmSJbCFbcT1iNOnUh4LpfouxZc
hz14gloDWjFJUeDigzDSK1UeEdDm6WLbhIXqNvEI81MKY54QT3cRTpnLlGuPaBJNVNk65E39efEz
ZGdyJHuCbDtJx7wh0qm/08TziR7r85sPBLpj8UFDZz4ZUOv2oLkk112TVqUWBMWCxG+uwIZWRrqI
WkWPM5TOiDrx8VXT26ZaKlOQbrtulkYRtwafdYRYzBxsx1XyyIW7zumlI0cA7/eTcmCTrtIgtl9R
zjtOEzYLQoCfonIhnPViS7Udbz23xyQqPL/Za5WHDmLaonY0ltmUekdwJT65SYqZ92wwM0rlG8HO
kTZDkpAhtgCc3TqGz0JbioMWIwWaEfXCrMqkUdl7aN4iaaE1T3TuoUjOKykcIJW6/S9nG8Rgt2CE
ERBYirXbpj6uE/0wVQjV7vGUZRP0Umj2gHNBR6Mn0ZOrqY6FAFTRaulHcHAU87n9zkA952Aoc724
CvVqzmv3jGj5u+Pnd/EFEBov2fxOg3tUnlcBpIF/1dIAJ0rNx+HU+2S/UulKFjzd6W4QDNrkJKir
g0PjW8z0Sf63ZxeQ53a5D33SyGGqXm5WvmOCDiCWT9U7JiuEO789N6jKajiauZIj0Nrcvnyc7M5Q
6rujYcRrWEEU2qyBxkn0x2qj9UcoiLtbxdrLI9nOD9MYD13BAnV6vtHTxJVej08JfblnkJ7F6j2n
8HcIOS26D37VOEZT4UROn63wBdOXwGbxb243MnkI++GSiOkQ4+JMOZ6laC0QAawdeG3SBmdhP15o
+xa48KSZ/eXlMthDn1DeK855Fpkxee/DoEiY9yoHvc5tv0uUkiWlcBSO0L4U3zgqOFlnn5SZ1f7L
9eciFwr6VxXdGCpeDQyf8cxkLkFYgkdNgDcRwJw+N+Qpm0lhGU8KO8JlrArPoIGEtQl9AhCVo0ZC
sAD4liGpXZdTiOr9Sh7MvUZEp9+8B3KdG8PZd68Emw0IgFHdGd/lAUMCyq/Lz+I6C4OdAkUmqnG0
EZeQ5eRx8MpyPdd/j1tpJ+xm/kAIJVq76cSqqv/ZEvYmsU192HpQ4YV3+DsVyd/VViHmDI4ojn2k
XN4dqUzC87PzzHjh8OY9/pP5cmwuicT5UpndFpQwFtY0/BiQX+oY3i8gQCRv21oWbyj68dAEzOcq
5KV+Ll6Lnln+6DU22TlLVPx69N2MIEndA73DnzuGq4+CKNFVaxgkJQu0toRVAW6c6zcVO++4jntm
bKSiHzTfPbblZXn27bNJbceMXdpBRlc2dpsugGBDIH/SEGVrna78HeIFI+mdDYlRj/wUfArv5so4
cnljod8MKf7nnS8a9DTSoK/QPp3MWTUsgrs0xG//55Q1B0aRii2mJA7ZsdN/Etgwg8J8SL/Z6qtl
tKzrcpJ4GACAVBjgQ4V3EPVqN/95iJIl5HeBjKBWhLnrjFGoRxZZCOe2KIcEKKE5TvZac9u0KhVR
Xj5Kn05xDVvLdl3k2uvOrA3kVQ+rCoqQiqLswSkZXnPB8RlGKxyUwhtdYJOOayO9ZTvLX/qLbdQ9
MkWA/d8SuJbNz5pNWmMW9Kf+PAfowL5B8pVcIQz4U7A0O7YOQyQT1py8cNAThbdiqhP+qaKSCJDH
UbPJqFCON+Cm94OWtFdkdvQJDc5sFQEZw0UsadqEhMrkjSr3R+97IpmTTUSq14+7E94x4yqFc84J
4YuuKv72zns+poBSVQjYzw6gNGH7ry5aPsUHNqM1fnY9QO6N1weWmiGzxxOv8Dptm0P7QdRxS1MT
OeK1KroWsIb0RXIG1vmXHp7INCD41RkZDiv1JcwWu+B06tEFWdcc2K54eVWxmrmY8TrTvkM/qJB1
nVTHLg+Caxqk/dmaFPzqKxgLLu7s4DlJt4fqXA8xEfINXT47/3eLNgrjHkGl+gLU9OVEc1o/raFx
XTc6UKRWGKkbyLdHKmrUs0Um9pDz5LWKbvvF0zQiVMh0UkBvoUPdd2NnWCNH4tSqn5lDbprRbT/9
JGn+vAdo4/WHW+mO+4I3B8CKJPE9WaHwXn57clZdNDbOomvUaV66UR/TLOcwY3/MSdsVrVuu+1Mb
XQi/6kN06YQY2LXXLYfSc4/Iz/zxB/j5yAdqnsNmPNbXNbyfbUv2Jbs5+TwJdbCtJsvgklkoOaHo
bFIPfJcR3a857hBLVzPyMvhZXsRS7TQD/lj3n4Ihm18BOsd9duMkM/aDcwEG1OfR630N6H8tEMwf
ET9ZJu3Aow61jMfqZODnx+ZG7bEt3EVYdhmOLKJhMVBgUe1krbLUZSrfS3I1Z3muP919aD8XFc99
62/m3xmLqObJZ0NjyfZUyVXzW4w98vAfU/x9gCQ7KopOGJa3SsVeNjwqHdg975GQvigpvXs+JaYp
tn++vbsR3+2kG19mkPVPnx3kVuc81KrBSrMM0HfVWmDKeuKIKS6HNW4QEQzcrqDKTdWijresO0UI
8NVSHvQO/C7yE6oR6Z4sLpfgsf+rTx1pLq5FmEd9+NcroyxIaEMpi6M45CGwBixC/UCkM4p4G+Ct
v/FBSf+pDncNQABYIrpaWkBgX5pBAZ0qA2lRxO1v3ZERWFu74Zy+NWkdel6ImJJzP8k0FlSsa32l
l25LifBmhFcanBlVDnGB03f+Fzd+z5/xcieHbV4kP65ZtpB8IP3AFvscK++Q0ynRVP7l2n6HMSND
64YsgcBqc5/ie7p2EnWjXr8NhA6zoxf/w63NELP6PH21++txfiKYh3I3tEVywcCl9CmozJYRZS47
T+z5nBvrgIeJ5vsnEl0GLr0m/xmaLOzx2cDq9zQ5/pLq2PlxUr8zaifxLclY6M6lHZYTUeXoTZz7
Af7BlM7g/0rcRG3PVs5IHOLDIOvu3puZbjKij3l/EYnlled7yW6zqK8bvxv1zxc9K4fjnYNJ8pci
OJ1xNjePyTzwBWLYeKgZ/hi96lzs8gr7eGwXSYn7Ydz3Vls1gpB6pUDeXWv6fwzvPgNPNSgRIlyw
IXkQToGtXuqW3D1utYtXo7b3IKOpYaxPtYpP6F5McjXMAcWeH39uMoDRKJjZYb6Foj54c6iC1JQP
NVE7in3aysRzos68RF1NK13AkyiCFGTEKBLNnbgWyR6lPe3MKuqyb5+OnSgnwdjxobBcOBSfNyjU
LIASPRXUUPZU3eOJ47k7lpq+yD7hmrZcYAL4Vg2b4Dm1QVEVP4oiNf2XGRFC3pL/64NwmfJCuI1+
RJAiEhfvHitfklntaTkZR8xrBUAVOloM6I1ouPnpUargu+Uc4XUAm7hILdAC7EJd3ZmDT3WcB02F
WOTgLB5nvsL73CblZohfvkZSy7F7BePrkKTNkFQUOztXuK75xZZ/CRhhLbFB9LmITsxkT6/wpa3T
9Fkp0q/HqLDo0AXau8fquze7ne7H0UiREtb8nYJ9fvEY/yzMQdzvaRpz5EqJnqm9jIHZy+X+NiOF
tCRgp2Imwm8USY02BC7T4T+fjFgPuOIf5DyOEiRCEfh07PzQbF1xMZUXyc4Q8yBolQuIVKrhMgly
+ZMCvV9zxbwxZxsUBwu+6dc3Vg7KYc5PS6euL8ncf5TeXbKwiXYNi8WIvTJzeCxE8w0MKkiiU+4h
XkcY6DQzVmKRVyaG8oAfI8kZHTJHamQQ1dJvMLmLM/j+L2Iulg9V7sVyhr4W6sO3UAKfgLownFE6
JCzewd9CJTwg5sCiPVhitkwZ7G5ZWdu3BwkBd1KV8YpHOG8po2ok16w1net0qrSPeDXsjqXqwKdh
3tZasfKBtGjzwIhfxtSMvrb4f4YzMKH1NhJpqsiA8jS8HzNDNC3dUlRzgvQUIk7br+pVixIX97cE
vkiLARK4EZZC0wMfb1+vntcSF1WlOEz4xt65BZRYoczLpI9QJ4Hjg5WxS9SYdKZpFu93i6rjLiJ5
AVVm+DqJByNpLKijpBch7zJGzVbq4QuXjTJB7sm7aMVBuRAD2uSdGRWy1FJho3Q8Nerauzs+xoSf
aZ7TvEfTZccgufkvg4A0Iivo82y1db1Jn91aOJfM3k9laAyegCxJXtxzRbCUVFzLkZxxCn8E6Jmy
c4aw5tIDH1wf1XcAQtpshm/jXsSzpPDklkNLZaoFwEg4inDf0ykl7tOQCB/heSRzt7JgLvR06N5k
slsfDrYtZ1bDsUtFAYWrWUcDIr4QWbxYaKuiWuRFR0wSStlmMVX4a0aNAUrwf75TJrielE+HpzQv
w08Dszn+ggIQ7Zv/aPGqGyRI2G2Cp7/EUQ5Y0cYizYjKuUIN1cxzZpU0yPx8c/5UezmQdQItgOgr
k5bUE5rMgjwGiKhTdd1T/301UjIYoI3P7KmR5he3jOih3A4iwn0Aha4yYzTc+pm2Nr4MR77SaqZI
fixR+zEBxMb0EWZJUgiSNhrzdG3vDskaavthao0meRzEdi2pvl6sKv0qViKnEFJOJ2VIAqGhqtO1
MkfuPbUav6hn0n6kGFdUE4rYdZmsfLA7h8MIYJMQ/6oZmTdGYC8b6mjGb89jTebJ5g8PoHJTT1kl
YAGdA8PUcz91fwD7lixEG6kmoSUAsOaV336WkQuls3z3J0k1KnhfN7rZ+usUM0o2v0RG1YBvXOY/
PrzYrctKuE2RNgxpQpaFMY9CQ0U9uzLTE5PPoXowmdrPhfe1JU1VZbQdSD4NW+mKXE80o1yXSy+4
jrorFgundcDh8VmToDG0dGxeIS+R3DdDlYqPW7PYhXqjw2RFHRqR/sSxdenTwfIeuKwlHpEwrmuK
ART3bMub/z3OwErb5P7nhwEjtInE0Qlvo2bEuqaqEoSWdKZw5VKy30VSGJyiI4xh5QB5jwJSCKoz
xnZQPNe5pvFmxNoKrctqyhxSC7kKWy4c18DKHpcpSL1XDv8vab19Q+z6e6wVNwST9nIWE8ycOLh+
D1ybq/o3rZ9IpYKp+KlSW9SjB9nISLEl1ABmlVuKbYBFVmVSH9uizTtnMLADMpthz743xHJV6EW7
/B72rztHftWx9T+zWLJ4bhMoQjqTITygzxiyzwlpZkCWwfAXMlZBdP9H9aH/TKWoLO8+snuJU7PE
zy2TzF35chiEELvcCiCsBkmM/F74RJeOnI02qzSULl76DE4HkV4uWW+R46XRN2Ym7PlXxTAPXLD9
4OqVB/ZbzgZ0Eeqz7wv0uoLqgILzjAEe0UGeu8+uDDBokxHxYPIs4F8nyx1GMnNwWtrUOGMw4Uxo
p+Nl8rG880iy3VoObPI76o0D86c7BOy3x0GNBt4RNtXy9VUW4g0N5+WL13yvwxirwdJEni0qhSsP
Qg10R7T0xzTySyNZil+W/euev8YLpIgpSPqHCvUpaJfc5gbjRt5W5Kei/IBSgtYcCs9tUZdJrLOk
TYplXZwtjThRQaNp1PL0EA+OXwdpzh+q0GT+niObaQqOhEXHyyJB6uP0Vy/GTyYosIidpSye9nC8
X6l+6hx+b9Za2Eebj5EAgRkKL8XosyAFEajThPHz/Az27rx1WgXSF7znbGRodMoH6P/6kqFqXwWQ
OFJSyB5rlhIskZA0bN2xbUNfSVmJYFtHNHjLfHyMkGmYyriHhCmiuF+waNC05gbx+IWEFenpcZYP
R/X8Uh/EydcVcQAR67Eb9krsYe8ZTu+YXVZG+VcoYNcgn63O7MomJ32vfADXQ3pYon4/9hNWfOLr
+IdqOA+ZDoO5e28GJJMcmx6xAwDInjIRxPx73EGXcfr0qr/lcCRuv+pYGO5LdSYSS6nx8VDS/2wB
iiwd6z6slYhF/FU1dOQkBxe4yI5NOgXcsKC3J8VhDyBaW+inVhhxyip1Wo8FxrVFrZE7sDcWvu6M
zuaQ0mhvVT/btfJwIhv02WbNH0RCgRbsRXE+8ajWLHLsjMj7fE2iBS/yVNba1h3hVXU5y+htBDYS
GA9jK2e2wubbW83Qlly6OGGwlwFDmWU0HLCh32ysFNtZQwdexE80fxbc4q+uV81rteP+G59Qqxxq
rrKXZiCa+BPXQYw3BvkLDQrUybf+UbU9Yo/C9kevCUdual+EAjTt9RroK5v4E+CsHXwNEdkwvmZI
MMwuQcCvBE4DpjJYpDlSWs7GxQFXx1khLZ5oxi8WD2Epfkq5FdLZjjAI4Acy4BwD4RTJVJPCp+BD
YzsA6HQ8b+8Qsrqe752Gj0C2+buyDeI1UMsJ0fT/GTxYWNnRErVw0Ud4ZxBnYS3Ju6tDD39eWcec
U+zAUFDo9K3hAkljcWsLD0nqf/TrVl3UCObZTok5UQm7TVSNjvlWechRZjAiI3f29BKZVfeAvBBC
3NPM8l6Ilx0Mcs9LbG1yk3f9tRoVJNSPskcX1o6Ga4zNi9wJOxJgk6T9sjM4NFjdkbiqVcbke6MQ
/xw0WBVBSntXgaFVT04E8tAPhR4nP8XEb7Lpp3Sm3bml2LW6vRwn+g2XOp4EgI554rIHQpi++U5G
xRNv0LkM2Zc7/pSeXt3QBXHVJ/+FJ3ffrr67GVVUSFYXMSvFy4xqj5ZTH2BYGgSe41GeYFhqdZ/s
EQT2a3JYYIeSVWLwZgCqT+goDHf1pj2Qgmd2e6FhrfdSvXSScNFtKz10kR/uneGvd+9tGPwNJME4
p5QI2fNSwCMDcvahU6GoECjsC7aIrXlXtPS8S/vb0pJmuaxJbTYP+vsyOc7wepsgohYWNQtuxEQL
2cvhm43d7jNMbFQrW6qBQZuQZWg25klARQuMR0fkgLGGhvuCd+7GmocaDKIW3c0mNspw6k4FfVtg
go1sZn2qe+OtMvMfYhXr+82/gFNzqVcxzdbdniSqZSh/rVm7z1NCfVrvCT1ZMx+y1ktJYyFo3OR5
u+u0ri9o6gW6bdCXbAy5goKUZTNT1QTNHbiJJKDJZcZj9n1R0lmkPM9UPuVM7hrWdjsPerjHy10f
nT2G8DfFlA+sJAL4aDo77XX26iDclSsWz6QD9zUNGdd0m25PfOW1Ys1zPUeLFhs/v8iQUVxvMKac
8cybu2TQ6Yi/CQgbGYkkTbEdJPHCWju7LSNs47C0I1hepGkQ3xNZF0gwpQKIdu8abvUZ/anyZ3V6
FAjMet+VH+ul7CEKGArNz1N0+UF0l4fjR6y4/x69KsihKXDH79saEdGGF4SbW9brVQzMEeztGI/4
RjNcTZPYvB0EfJOTzp1dNFjDXAwmWTDQiA7q8XmXMCZ34ww2HNEr8Ztswf7M03iMzY/QySVu/UvB
nJS2WJPGxO0FuS/xdzwusxcxG0Tc+CnbNE2fehddygynwv0TGKqQlNfG6n8XCiq4iz966roc69mP
K9RoMaYG8t8ebevBjtd0U1thMXhPNmUo3f/PL5mhbXhsAsQ54TH3Lq8PfgB+u5HBza+NfMgX+D/2
anzJGGTk47fygcYQ+5/yqTdOtV7otwR7/ZnXDIWNv9mFVrjgAhcVdgdE0mTGUFhs0k9YsZUKy9L5
vBHY8KH4H1Jz1t1Q9UOHyuAWkQF/lalSrRoP1Xv1mYrCZXBmApB27UxQym3xYmVC0lc0kTVllhLS
yZiI8jDmcfUA27yMvyn9ElOYRfGEaHj2VBb/TMUS1cfcc9S8wtKeOZlt2d6nf51bkqDOMmg1ZY2/
jPwCHzCiKU3e7IS5m5WXczUGvhD5qtLIXKhbyH1fi7r/jY9KBzcsgXFOOijvpVsQlHmgoxZRIhW5
Y1WuEwtzId7aFMV/36FxPl8II3G74pDS2DRyQ1+Ntgxp/IorNTiW0LGHFIbISEsuwZo1bOW0ZvRD
pjBII+doJoms3hWHpTmlmtjERvOU4fzjQsqKunetOiYicpv5WOgIFHWaOuSwwaevHbjIfpijZ1Rx
6YsePzMzjMI6zPpa9Sw6Wwf3dqjhX5D3qcJD+fmy55+szvB5TIuBS9EBTkIRtd1fuaxtgCkNWezc
CjQext2Lw3N6jVJj0qRAnWkEKkDCdSEh7z7FFeEnAjpG2emYSvz/VMgUjeCDEm3jybHCnJqGv1S5
F6x5gxddl5LRD/7T4CbquATJdmyvsv3S5MtjuwTPlMKPgu1px6DpAgUjV7+JcH8131XBgob5VmWv
4YL7c55pHUKpyXCzXsdukfGWYYi13ShFcV3sWKhR5Nu0aSMqj2c15qrYoyKt3pau0lKZxlcmdSsj
TtO2LA4BqSSlRzHTZ7fvcBtD8Z21DoFgKkijy2D48p8v2WXMn5NCt2mYqW6Xv/lyaqmC3zo+o6Yr
4G3VgcFZaKWCbKMom2L9zpBhH68KsYrx2XMtOfJIzZCD7s0V+nsqW7W6dwo4f8QEtwPQjsaGP7VU
PzFULF3aHYZJ3WX9n1QoAMOVMRFQFUBFkeLbLh+wZynQWSXUrL5mZjK55f1IPl/72klDoj5d7smN
VM+yzSHU3FgTWPfle50kNBlyBPkWOqvSaA/4A5DKaKRS25hdLoJMvqtGPXfO8Tk2/D4R6qu19LQq
pLnGdM5jVU1hjGRgW8Rb52IRK43nzmW1oWv2E6ol6XTIFbmRA0rcXMOQpsOVjgiI+FS2R2iE6JVp
9Lad4YvyE+E2BeXkqrGeHrFJJ9/5KcNubxcGW1BAeOgPDuDk5JOcjuaVUE+JgBZEGJAWlvIOWTZj
CWdDp9JWr5pShMowQrTpBF9U78felvVPg4Q8ERzZcYKmPsdTexAhdg6QXX7Bn+cySMqeOh1uP3ja
pWGNMH/iHiD146N3NyEoKFeMi152YTeiZFF8dg68Uf6k6f1BrytlEVOuY37xjcDSC50Tu5q9/Sd/
nnAM405pkOW3Mo5CRweK5fmgWzts8TG05qfIu9g09Egq2G5pkHyoxVWaCbfLft1YjYhbMlh3TG9z
YkV2nSAJDWGKpN4fGtgtzj1/SZiKeGb43s3OtNHuy9LY7DJ1ZxR8LmSL9QbBauMg9IKs8g+JR/TD
hyIkdMnPQZ7a2+KrhcyfurkaPYsJwpQIOhEaf901UNXfjfynsgrBIkeTF8gaUgovBhuLrD6zEMYu
dxFMIEm89bvTDRhv2nZQyxlCSZHpcCWDYPy7xy8mqN1pNPVHf9KHMrwg+jfjWj0qtDPEeFK46kx3
Ks7g3hFFkicJQze9AfXHZcrLEDq+ogK/v+DYe2MMDqcSk+DaDJ6HcPNd2iXRMwoW2o/IGV3oTqPc
38FgPePz9GVnYn8AksMKVPcdW/CZje6Bj6502wwWPSV5YylX4stsueHkM6ctMOmatQ2cPvmCmgx5
wJRJ76OFqmIK11x5z/agipkMGfGl9Bo9iFfno/V1Be9QuGBxjJcGkV+51Luop94afLqUEjQYCdWc
NyLGInQIa/nfDshj/qyn3dQ5wPAeqZSHgvv61jOe4CPzuxuUQwj+Ikyxlx+tAA2yWxhwYP6Oniow
tYGdlGgemLX02//jfQ4f4Y44cYBJSvzyNz9LyZRUSu02+VKFQt8kAAsWSd6pt5eYkW72TV8zs2fg
PFu6FMmtgYYGTM6KrceIfXT6sK4blXuSv3otZ151Vjg7/716AV9me7cYBUo3g/uQg1hWMZVCZ80L
UKVimjRco5dmViwuwmS8/lphoJj1aGeydaNNb7wpd6BHBqL14WaBC+0E/rbMM0m7uGRvoGLNXIhQ
yTU96C/e3hYyUD7bQXFiLMF2FePVgvxPCEDClbI/AlaB6J84yJP+yhesmKCYq9mNaJGwnSIZJt/K
j20PRAcu1xevAhRwhg6ef1XX+JqLhrsfCaYGBRljD3r4+RjWTMJNBlPEsBMW++NxVuZBh7FbkpGl
Jrh1bJTQ9jHgxfocG+7Mt6X5SCmRFNl0cJOoGQPAkxUopsTOrAUM47AZaZDGsmijncJ2NoaYxPKr
tZWi+9bis9gWdlneo8MHHmsehQVlKOnxfqc96+BOLO84Qqmd8hPXNTOmwK6NliYHz98++YSaEvXy
crUFTo2pcoBhnlCKd+BkSeBu3ylxd7xzVceg7ad4CjBaD5I/+ei8+6CKF9tTqf81dV4iac0UWhlE
Eo13MxgpizTHWC2ZuvrGKrC+t1rZga98/lrok5CAxSJK4Y02Y6CAgze/jPV1SM5N4UOe+7ip3WzQ
PzZWOU5FeWaO6PF3bxJtuN24SKzoXPHpLUkRapeNsk8XFElbfHqK4fvreO+8if5s3N8zDQhDsUUm
I0fTtcjWIARGDGkmyN2k9tetQR4c1VV+1jVXvleQPfL08Kg5BGsSVciMe+hrbx7OXV4DjLqdM1Rs
oBmrLVKb9uDxRmyWZ7GnMXa2zS/yIQW9WeEC7qBjPzQbvvJ6mmII+KhLDmtO6xttUbupod/IqsI6
t6RbIWoRNHqVz3kVc5fj4c13+5pyVid6KcB54PHQVevFk1jOihmrTDG7Fq7Ug7JJwdzRc6CmmpCI
9bBpzpHfsQx18pPPUujx1IaKio44l6pGRfBg1UY4iIxtDcxsx9g3Cuc1TH/ENIgkgURmSMYIIR+S
760d0F0T7Ah9xXdmZRx5sgrev+1c4wVJRgcuboYPa+zs1qB4WSJe1/cONAgJctaEZe9BnAfsT1eV
Q8VLCyBmJWentuqsPYbkcZ4Dq6WrP1hJTfpaRma9O9PgoySXYeNNp8UDWJXH5vK3++IUSJe3rNFo
vXUGHzeV6MWXcMCEnaqd3GAgJdouozZQzrto9EOLsZgldqAWbGXmrQa7/sa1timin/S6BDHq5bHm
+jHDoSgY8Sydwo47Dl9hYNr1JJtZ3EWWCCobkzqddlvKbVcHbMdDF/xPmL+MJo0A75NUQFtt8QmQ
1VRnsn/3R9x85ATm7CQL+uqShcMp97ZmxpEydekmktY7XVvo9aLA49okorgmF7SsM6cvCxm+mF3L
k/xUNZkrZqtaGGbGX13DL5qSEgO3eSpVxXjcZxDs/43Tb0gC0t1zcrWAf5xMOrTctaLPDlSMEtSu
bRX+VTToE3QstQ3nCeogiVBc0fptZ60h2Lyuv5IAKmqSAgP5wJwnIglD3ybqTqxHOGlYjTd6TvSG
wiovBq1NyIyEr1xSHI4P/mEKzRZayvq5s2rgE1IBuq2gWSC/CYQvbCFCVWJ4N3ObVfoUvzTS7PtQ
Ngh3N/eBAxGcWYpYBp/6xrynK+AjycODDq3rEKYMT/SyTVk+0GzBpjvtkx8pKJDvkyURtCZdEfgF
7byZ0Q2dZgQsmA8HW99y7sIc1++6MBgI6d2sZTZaO4WNvRUgA+WW6ZWyDv3TU29T3q896iAkvz8K
J3kizgnNRk1FKr30LItNZAgPUu1m8ybCGuk1jadF4X0RAXGDUaKVm/hbUBD/6f8OxpgUp+ms/TK9
OGAaNN22ZEeJmC1zQWeiDE5/7PdTH7yJSXSHGi1bEoQQTAHxCMH83VnTUI+x7QblzSRSmj7E8K4o
CNq5hNNLT8SHqt0hG52+SKgZPQEBL6aTHQqx6IaOzPApLgMpE96GS9EIkNlUshNRwUuspbOeCMvJ
4DpEAEDgY/IqWykiKwSYGB8biobBPx9lgBWuNpcYmFbrHYcgrLyHg7xfXnPlFU6KSbtT+s9h8L4K
WWBaOiIzX867hKUqWC7BjFqYUp1AqGgrU59B7RsAPH63Q2D2J07iwqI3xeVLZdbaR8p+pNKQ8y7E
5+JvUf0kVVzdE1IezYIM50Gfzn8nJafPU15TEuUXxznchn8aAT4QlczXMep+OPLaIt3l2TjBBxtI
hd2WIh97RgEEOVL9tzhw2JCWjcNwfyjZwF25VzZo8lho3Lw6ZG5EQ3dZrFxi/o8M6UeIS5zBEwU4
qu+loGO1Y3K+mDc4RbxEvNI8FuRPSveoZ0uY5vHnIT8QPEhP8GXAbO8i0d6dMvxTL+OieSNQ4jnm
8LSIN5F+hz7nwvZh8Xf2v8ZFG8rbqxPFmvSvnlyO6iX7CedoFyxnXysrEPWRMexQFsxZ8/v8y5l7
F00B95BtjYLiOfGNXBB1sdpvUN7Q9mktrJIU/J6PrA+s39oFC41M3p46phsbXjFIasF4MAjfK9ic
LTxjMgr677VC3pxnvOucD03Hm+BLWyHbmsg4m29PMmNptvtxEdIj8qPGhKKTErcpRziP77fLg/FV
5KJvNIHQLAVivE8fMg8q9vutcHGEoMyk0V+EwEYgOfUY5+0SE20PPKrXhpxN0mIHWm2aFkJuA4ND
7BdjZscJrO6hqeR2C8fdgDRZADMQaqI0cvj/Ie+WhvmXxjQyRNETxhFx7scIh2/uwTE4KTxAGf1q
jNrnzNe+kAk1sq8w73Q8AYqnPRUqXdiGyX6axQENKqCOj7m21Ptv3YhvTP2u6aDkJPhnS9k9tdd7
DSFVeCbAlDCmsOjTcz7zLkyj/o20wiu+62zpXrM9WbVkqXDOUhvuQii3cgB/KWk9u3q2GjnORHRH
CKsQ/ttMK070tx+wZ0lk4wkeEHOtYrdbYGjIvRPmPU0+QIJ5+HOCUyz+DVxUFIWM2ODZtKf/E2cH
Ys3NRCJ9inDRkmDHkCx6xnv27g3i9rQZReKZpp2wk2iOTjnm6XJDYa5Je2syyIb+qycgAUhwT2VO
kq34r7UqIW/1FOGkDMqAfwAQyfBDEh3CFPrXrBOBrD0m4UgN8A280PYs//uoVGsd9kahpjD4CiUi
ZhLkNxP5pwALqGqRmMCKriRTU8bims9UZtfJZAcPX6ptYzOepahEpmQOZou390YWkQ+0JETGcjNL
iA2GjQtxg8fLS5Z8LoT+DlvEFyZKEJ4XcyiIxHMyDqE+Hd9qsisX2Q5VGljFkk6ncZL1gncAqwxL
WJin0k0bACyLzOrzXz7QMdn86WLKnRaceU2w8dU/3aRPuVEAKMqYVmCAuilzuE8uiOaJ4Rg0NuCc
KltT9+AUk7rFWjrmb7mBk4rUUoIjLQ+wSY2eWb4LPqoOrVhoaic8nwId24Qh3JEwxBf9PAhL5RJN
CVJoadlgP2KFRMnuuO2QsUJEAQ0KYCrMj6DGMAtxsfgwDgrqsI96yEStPtugleLhBJAjGfcM5nAM
XFYiW/cts+4aUgRFwpqRRM/x2zIWVve3nf6vV6UeTtjTrOxFd8mJfXltnuvJ3WUAg+ANcAoH2kcA
36pyz4vejBgXA+5fHcLKzSbeu+rrmVj52gELmbtTgEHPF0W+oNHNdc5sDEZGXAi5Fq7d2ysRqxVr
oyy6Y4pN/dgiDpXRmK5e88Tbhn/ELIWMbSnJ/7eXHkLspki9gUMkLIjrQPU5gBY2zIt2n1hWl461
lztWvH1/RPZlaWFe5TlfXOHpFXfLfOmCpEIIVgKqiPlqSA8kO3SJLOjJjnt6Nr86Ap8BNlwwB6r4
MJtjQlMGvo+ZyfRs6NN8gKtYMmzxUFl8LDxgCc2/IFHPvbt5hmLXM0CVTdry0LLRbs+VqwX/1QL4
QNZVHB2YWoyC0XggWhxJNfcNwHRXQpir2yggbn61iz0Qn6KgsZc7MostA49RaeWns0WEmfItlKsF
20Pm9y2Y6EiBNjgYx84uVWQC4/wqtT9OsMOehg0rH2QIKdDxMeRVENgDsDs0Lu3WRj8XRhW1Olj2
dsyTTkavKIE88sfaVbONSL00IQIJn4kFWuQ4b10yz3158uJm5Xcs5Nuk3YNxEUb9AgQF8d3SOVyw
Pk8UY2kljuSuoeamWYyX8saATrT2CD51W/T2csHrVAJ0qTFPYD3En77KJgIiVI8IUJzl097MgWsy
lXVuQ99zWIWNgcxa/LFgEbTo1mdtl9sqIKqUYkKt7NHF6Rm3LD86a3DEzIRZ4e2nV3jxFcVm+DyV
8cynEMmd8x7hIa5UPaOLoESKeG5s+ybQk14d1YEPVYg4BiSAeKz+aySFCcAmdGBdOY9ImVfN25kD
LOANkE99JGNbxtWWqjYTCe5mrs+b5b6Su46+unfBNLjTCE+D9QqloDP1yELw3+/8XNURYezLdf5b
/FtVzphFJKTZe7t5JTSJvdfLPDtXrQ2I3qy51DbnLztwV+jqUSoYJsU6U1ApwI+pweWmwR7IFVma
NjBt4Y0CyCcWuyJLTx1V12WPU9/umvq2oIlOOiSr7FiiSmRFswiRGP2pe9LKA+G/WeMB9R1BwU0B
Ph/oIHbl6fv4D7WwF/8az1RKwuMJ1OTWVKW+Nta0dW9LoFD4+KWWIGQH/L26qWxOclmPegITma7i
pPJxiCkdR+yW9rc+TdySIyhiCO9jcja9bGLM9MlPwmFLqhllUCQ5G9+UdqJvLkNtRgJyqm5xaOpT
sCjhmRYUt6zQSqzcOCXjwJkVbS90tjnipTqxeiNTpt5jhJbj5nAAgA/lv6SSZ+QUe4ZNxOu4+X5u
sg9CD4UGOXeoNG8q+q/l8v/jQrAhntpzVAr9Ifi+JEuX50AnidTOEweQ5RP5ZgQi0Dweohcint4n
tN0dJv09ehKUO0Cn73AHtbGH/aGlfpiE1Llcbw79GBorgr14N/MZYZKk+u85QNSGV0wDq/XiLE+T
nSywz5MXeAY02j7ETEauBlREQXPK8PdQpm8KAWjfI6MpiE+WH3aVYWxXRO12/EFxOihYPaRTt9yB
B/HQUXTLQ3slh6VVYEnn9xYDSS/Q+WsYGHnn7p4kzh/GMkpk3tCDTbe5i30eSVeXHLV6xZZH7a+n
qEQYXsCB1aXYg+yckT29Rtsv6S6W+kaMRX6WpNRFbvbvzDHU7+8NtY5mlfKXsv7aaMb+pi4+lzUK
eFAWVPtdgMP6CUrjxgyKOElxeKnKSrnzKArFqYhkQ16e+qZVrUntYXXjZoVMvNPadySSQAetrWcX
OWcXNGb8OCRg9944ufvkw8FKRq//ZptElxRWl312DZBysLhkjHidGOGlsQA+9dNkN3n1D1PhETXi
UVPxc7AF4igFGkZMzrII/YogLxvJhTDszcJ8sW/pf5txdSe9HaTdd/8j5r/1273Lv86aILZBOdJ0
XG9619jmSZvUnr7IlFZ+kZc/d8WRDnFJbsWAMCDIV7FmNN8SCcrCDYAKsUbhYxblScN7Zt/8/9hl
sUmisSqnXtkWqFxqrI+UCXhIp+tTQ24rJYYouk1CKa5yhaXA0sjq5h0zdsdorOBJ8kwkHdeq1oa7
EePCHWZ0zdImh1oIRs/Uwviae3oK2i+ND4gaHnhmAIdlwZihw9SXesuKW89ugQpnv20M7wXLolj3
fhUPmQwlNEpFxzTR4c+PX0KsUv9b50+9nWxZGqHRtYa4dkYCBcpDNwoKL3lwkQCExzhfOuGUmiSV
5hrKek0s3bRIU17PlFlnHoglCoEDyqcLjk2k65dLw1Z2NTm0QrI6P2p1k4E2SjtUaZ9hH+Tm8EVh
g26vTYtvHA87CN9G1LGCMVeTAteWXa1IlDEQL8gPtULLnT0ab/Aubcx1JDcHlZYbxh6L2oZqAaFm
KuRVvn+/Es6Z6/tONRi+2s3RMRcox/CFesSDF0rlXfQRvNdYOzvE6JMUzcD1AhPVM9LgBJnFgvvI
EPCJGkWfvrHD4R3AhNf1xysrKOhOyxw10m4DwAAN6xjBVSdAoDhtRdLnqsxdcSoSgcqZq78epoV+
fgFpqa2KsrnvN7//21z7XAOIm+5nth7WJSLWm1C8DX8iDuK70houAzvqGFxG3fH7aREfcTX5Vbec
whcZUT26q1n6QTQ3Qsta0HBef/rBNgvn7RxXvMEtONZvu5sAy8iRQ+2LCd2UeV33u9/a9TYZO5km
WhF0YB4+3mXxpo5BpZsLjlMJ4adm6EiUqZCGd8coNggfTq8vSrCmhphzNWT/yKd9CVN2OJUY7xiS
9j9tmLOALZdCrN6cx0d5lanSyxEfFMJGzU9Ei9AEGe8ER2mzcs2t9P9JM2Wb8CudK9SUkB4Q5Bzt
RJKY0+l2uNwDyYeYw9mWC8On+1PmgU6PtkSqCRxyUOzw46FXmRTYJjr6+13Lq7LRlbeIqLxl5qJx
qIMALh1f4ImokTXP8etOw9d3/A7XGRGzHbtVKdhaA5332YJMLkxZkpMOzGiEAgNqBC17so5UAuDi
od3mZ66T9aJqanUKnLkRZykt6hP5o7OLB96QxyUStW9Fy8/c+xLoLqHDUBs7BIAZ94ctuzRYgtNN
CuyxeAIQfoH41+CD8sHMJmD+L45zRgZq43oTn0Q2HL0N6aafB/Llykr9Q5haeBwE4Oy7QxNSJaza
SEoxgaWQsXz0gqyWKkjsS0eQnsg9uyzyM7hZYyGZPrV4VKHgyDNgWm5/zoIDjry/FJV+UoKXdOnG
3wZbyrU+xq+3SDhm9VuE+5zFgqfviUowf+orq1BcUiOD+2SYmg0Q/zehwOVkzi8vd3Td8oXLv2p8
YWF5x8CAuRtgoD3wVd5O3OlumFcm0wNBPUeiVn8E1+PegI1UjHCiTX5Jd0QyYF+o8X1BHcnKJEfJ
xrBcTQkvVnka2Va68uOV/006jLRwkv3muWS1a3O/l/9mDFdqtsUioC6c+mFKsk7BAMABtZrkrSZM
+ZR9pTtxephn7TwfoRx2S72UOno3a5nnFP8VdK5FPwnPR0JSWBlPC+waRrwei7Mm0UdfE5ePRDzO
WXfllK+OivcBjjpzV9VmNOgNCoaS0MF4J/qVqShPKzqpO9Al4/Kvx39kncnHURkX9dtNmpY6EuJi
ejHvxngw1lD21B1j+raXg3/hiUMtVjINuMRBp0EphH7AqRIdWL5tfchmag/AFCXs3DqTIEM/wDSz
pBaJEnwAQ06HQDzXpHsD7zPRhj9VGadIUaiMwMPV+ce030CDYeHwSxI4SPZcZI9yWZmBWF0ru25p
VScxuyS5WK98GDdgJ707uDkv5Tyg/QJdaYh38k0kmXrztGKhXy0uJ6QFrKtTLW6rML2I61+Plp7g
OvEXNvHdgZsye2NFvd6pcb+PD1D3NS1ddQZzJiNAXG5HIV3xeJXpMsfaWu0qnnz7wHrlFdKhKY6m
JE5zbjTftCWCkvACHJe4er03eUUZHZ2wVsNobPDcqEfrM6ZbkOrx8sQX/YMcpNYf3a6cvKBgIhdW
1mLyuMa44r4u9BAQayRrvJnjA4pfHdS/7eoHzFxiOQ2QdfNyFm34frfJKInxAs7cwOmvLY9sLhkX
fIr0rrMTZ32VR5nvD4pcCi+GUbegw4n3B1SWeE7ZKlp1j5xLeWgblhUquT6KkH80F+yJ+NMFOgPI
sGjV77C0tBIkJdhXhMh7QDpPxlNmJCfvJB6c4POmghQoTkfa9rYUIcrYgGqN+StTjCTtYYJV8RL2
O1ATyIQHoj+K7unc5hoH33Mq4XrI93eAiGUqFGTyj5YkOISM4HvEl90Ac++aervvmQZUIlfCAHoz
XqUW/TNW2d8TD5SKSSAYNSWsmV3qrgSRHAQZyCEmw292Z/uwcgnfkSXLSksrykFcYcoJnGAY2Pvc
7DCrW8/IOPiSckjJyMvNP2vb6bAq6bqvODDFs539yYIEweeVs7Ojxu7ZFCTkAZeNWC+3EZ7vqOZR
VMbjTvdvg9VIJAqvBmcb1IDB3OD9nXyYyFjWqQhBu68whvM+QiM2IP+UDVkxX52alP4dwVPfidWW
MIiiQuH8XouG3A3CwXYAFlPpzhQ/SQWFFcpM857745XHNh5/MSTElgrk7bZec/tyWdsk+XQEigkO
5V5YbEGUTYiJsS59L7fKMycXfDRXF4mWXu4s8J4Sdtfg9JoGJ3hik+gTDVIGwD7115Pj6LNz+sa7
fXysKimDP6ESPYl2AtGrtiChVh5gbEF9ea0B5FtQ7B9MruPhAngamvksLjflvE1Rdi+i3FoSDrZ+
UMSVtZwWadZJtvJO2t6u8kk4iC8aIS9BexSjSveuzG1WG+dP/EPw3lnY/dhmd48rRwrYto7lM1I6
zBjOpWZ0rjYXH5OUiwfPfZLVsxZjL9tZVrrbfvBGnqZHdKCMuzojwd0jff8VK0F7//2PmwlC+m3/
moyaVPU0DIpn6D210PXV+OisIMcAPua8GMYbylWaFVH7oV6kgXqCcxAZvL9zGUOQdL49hmtidaru
EQOlZBrh0Mskb7xSHANUMpBVAl6cKYpnDZp7NHFOrjvNVZ8iiW1Fd1zznYxIdo8wpwNKJzmL9UXD
GTwQuCYlSyE72IkFl8RTfpud0qxWeAiejRJZZfhDnW+kNatSlI9LTG3WTrHMiOkYnHD69e1BfHi0
w5BKYhXAxK/m6uQoKSyRlgDGe94uytd/objtZ0QacmWTjXLS8ekca9yrotd3y56twisAOPY9YVHp
aWwQx8oSL6Al9TBID3KKFsQ2nitil2tmoKwbCyc7ehfCNKazUF1+mvXFlP2TAlGacy+0xHaFkuMq
yZDK/+viNBONWPGBo4KhcAE5kjGlGz+Z4dRUxNcJ3c1h+Ltr4//ggUxgfNHN11aGuMLsurReY3uW
Uafjmnun/ODIJiMNRmIgE5P3pNqwpOwvST3oPmCPIDPK8xaKXpnj4yAogEJIYaxdHf0gsCyarfKK
DXPFe8Xg10Xr0tOY0+bpzkQ04oEXofAhbk6o7EgDhakow0wXsNrg2rs5osm2lZXwVg6tWFiyM0lg
TFLyV4IxCh1ZiuaH6zVcnTte+j1SwM/MY+a4L1s2n3OSybhF7T/9tnbStrjPV/h5P9aTTS+g5WEc
p1UoHkQhqfxtCc1SdobzpPqUo7WmQcKlZp9rRryNVxm/BWLVh5rXme0Fb/kYrFukp5xf2gf+DVi3
GhjKe3/H6qWVBEFK9gZxQetpRjSC3Fk9fRi1vIP+bJdb9afPzDTPEk+85pj8EdnW2y3/R+EpvVZn
5sN6IP2vYeAulU4G9CNjFLsqBdUzAjvkx69RaaHWPpj/DwRIOol0CR+25koGoZvjuyliGBxgm/st
EThoLvlYoQi5x6Z4c8c7VSmUNB7GKXDxZnpBhe64+VsCBprjVmxJBNvTi9lHEeCqlOcL8lZLZZV5
qyUJnhr/h+VbYhJ7rNqn1gA7xaT402gWDqOBoxGDfCsR38zn5U+or3pQLgRClvUs/Trn95/fePSP
TlKecRf02FrYeSct0wruVp+qGb7oKMuiuKLtenzYqH3V2nBl8FEc6uk8k8cL2K/6MzL94i0j4lKV
BAnn3uurVVTuWHjJvzfDxFh15elGptEsQnMhS5tJZs+HtCv73Tl8HStyWYoV8+b08Sy9ecEMC/vs
PaoXuJAiV7yJv9cnJA++DIk6buPCjvSzAVMVCCewmMYgZMlQjT5Eb+muZSzq5ya8Nkqn436YDXvM
20uDXbTuaDxaVKEQSuYrZFO5jzot9RqfwbDS7DHpBPCvZni7DxIjGux7hg8Vp9r3V5M7YQZEE2LL
TcrTkmb7GI0VgVy6cRrXTIiD5IZtRfCUbSFg4fipodPbah/38NLyAMHIJFaJnQzmj8ibtmLnh5ok
vk8qHJh/IQOqkcXV3fjEVPLC5CXDs808SXzsov5GmQXyla6Rv0IUJOBM/F+vUkje0yzwymn2nPPF
gQZZ4qIjfruFQ7LpACRKt/h4jJoV3tLi96mETebQxxeybQ5iprZv5hzwVgW5T+IycsJ+O/gYjx6S
3xApzKBfM0XAAYF30H3nASrsraC0OmWH5iivO7PB5mstGkpkmr3h8rdzdHLHJbvXS17ZFFh9JqBh
VBDwW5ZcicHMJVTIucibVp2XwEAaQ6Bq0B1x1oT9xz4MUTHAkNzpFVweeXlVoaeTq9/NVNLtfMgD
w3/qOv75PYnw+sr0f6RdBKMIdZA4HTyDUfuC7DHklWLcDrBaigDivGcIRMU8P+lx4DEXa2nqvxq8
sGDGve4Hwc6WCEbIb3W3JJuvJUQUd1bWZJ1B2ebeBHgXqovrD8uG/SEsRgCpHwY0cyZAc7U988Pl
1OMO2Sh/GD4icYFZp6PpQEIJ1JsQ3DtW5yDCaroJnEu0174sVtbE72uecpnuBr1WWae6RO0M7vDs
o/Gg72w3lbn4nQ5qkPditShDnkh4EDdx1d6aYoaeS1Hq/jM5cMw7m5LXAnZMMYukcb3ffsja8pZ3
p1fAHWHHPanIEqGt4jXqRDFphowQVEIYw9IciZEvA917vAcFeyHaUpFGGMtz5aatZyj69gU3z/ZM
NbDjduQH23xImP+3SWwdi2GzszAtYAeK2+Seev1b6Rc7pRnZCgbTjPHirEBWkKimBp1u5apMSmRv
VSSEaIhSEQbfSxP3TJXNnp7zmucupmoNj3mONw0R/osaA+4kNleZOjSrkgnPVrCt93EpOU231al1
pS99j/bEKL1WP1UuzNffE3k942ZevRqLJJWMRP4px87ZQiAKNXNRePgnL5bN49nqtmUQWwlLFc1/
vjXE6oJECSIHDOn/CF10NNBAMpe7uRqpALdDBOUHXFHH1iNvao3agMznnuNsdtdrlYhcuw7G22Lf
U36D9z6uo8XlbYhZXZbWn1Vh/R8bi1wjzNKUuVeF+2Zr8j2f/1wpEmK1TZQqLDRZa6uRlX9IziX5
UNjkQFj45MFRcqN7vbx6+Jd3kMKJ4JIdqU3PZVAepWMu4uuWbphLHGc42HVVNhPTzr2JXLTTAB/k
oYb7fE0fNmBMtM3+QtGCGhKizUhduXH0df4/huftcZ++L+SZbPaw/RhhmHrHkrql4Akj/QFp/mnW
nCHxPHxVNIuYRx11Nmn2rR5XZHAwsa+XUVES61ambrILGSqXCBQvpHBG26/D27nb1kfv7ei9rTGj
UAgy54sLUSuQYgR7JXVhRlIy1j0UZcK4SQhV6Tg69WdL/bj1jhgFmFFGw5bipiJz7MgH2w64y9dl
bkSpE0wZb8ppK8zrgLBeVzpRt6DsjbxuqzM2S79b1HYdmDpGdjvGvNpw1ZcAPvr/hUlUNkTlqkC3
ysOGuQWfTq8MPcWnIrdgxM/dTTVmGNzVQp/ledgxLTOdwjGP8lN2S/o4e0+zEgPPFvsZL+tNF4SW
xP75r14eFR2DYDiESXtUAmQ9lgXsgtmEuQjLdiq8QcsWhNWg9X08M3x7ttOU17ERfdCXI1VTO8QE
aXJx2aS+6YftTeN0+ibuSabiHuNbNSA2US7bSAL/eCrZiOpWGZofggZArgokLeD1jLesnw6Mr3Zb
MNPG8Dq4wHx7Qj6Njzgoo4oRUxSsNVddOONfKuYQ8Vbu6qvW3DgcVNtzdIKw6uqnzC7TpfPfWvYv
y6jZHO8IXafX63z8hJhNdmEoDQoQ4Fjr4E6tOBRm3gMaT78CCBIzn9HeXa05dLfq1vKFa53zIo+q
65JlVP3S7H0hzKiMVAKfmmWiUP/PTZ/TzhBmqHez5K8eAhsm5dNBxyFmnPZQVfD84YSg1EQK7/Bz
XR4MI/zBEfHgh3E+iwgTPkGNM8DbCMdm3biNXrOBrvSfoO8L1oX/cLCf6pHb1lWVKI4H+WoNOI7O
JEvDOEoJIEkWHEeeHyP5nk0V/JAbvfHfjc7EfKYoGofxsTuBHJ5p0SnJtlF39h5zL1y+h33aFqO7
AmH5VzKi5Tp/DtJipYrS07rqHZKpKAvd73m1V3QWrGpZlVFSvKGcoph86PolJMluWNnDewY43Umq
Lebquh/j7XKAQq3CZ3YDNGIe7/vjgk6LNhSsBEjqsewrlgCzxl1tZnJFOO7awV6n76awwl32aVdU
JkAWxdcSPrjx9oRAjJZ3z1fKmbpupd1kkDUnfdqhNTElEtz/pm6mAiK0AQ7EfeCItUjnlXqXZNli
sFIbUMKrNYGZatgw65z7T2WFSGWZHbNniL4gc4/qbMOTQRsDEF1v8PECZbVEPIf5bssAC4gu78on
bJ2vHsr496b/urzTpbXVb619eJF5wUAVS3+Ypu4coVQAFKiNlc/pCCzDFoZBa0WCut7zSN9b1mN8
xOiAeap3BctjkTwoNtH2NNDnrEm5QbIUcXQiMieKvr17RjpP5QnaOPhy7ZKuryTnp335JcDiqDPB
ggxIG2DYdLfL8+bgHUb06sgyTK1DqQUuSgZebdNS4O8DO0BjQbm3T+phiJhfnV2rCQZVwKxm1Sps
uez2tIEBSxm7Lc9y2u+OduJLqcPMfTqYw3b5GHY7dIsbTKQdDJPcwae5dx8HyIvO81VswZi0l4E6
WDAKsttSzJOnYUXcg4MOb7NUGvdAQu7moeQ4MD7KQkKBdj5mF6AmcU+UrMNCv3wGH+lipKeRZCS9
CYYLz4ZLA5BK1Fwc0RKDX+V1eu/DDyapn82jd5imTzdhZnpd2HDyrVRrGkwhHf0OomzEfTFjZrmo
AYQMwmwE7Q68lpmD3OmAarLrdcgdTZCIfNp6rE2BbGyBVtIYPG308gRcyIodJul7ZMfqEHiUPQZ9
QPaPFm+r2m9di+HTLneIlaSJrG0CsKpWmEaSVUNOA+4Z9yzJfRjWID4ZdKoLdfNUoqBGJdd84Fec
6EN1F/anCe8hJrpW4iskJMOJQFMe2nehZfSz1OnEKygAPSKyVIajTm2BqqbQ8sRjedmHFdyn19Uh
tjKZUnJJctEum/qZCMqMla3A8mU6BMln+/TYZYLqjry5nkKW4QDv1sEyWc6StERBB0YMRfxXJLFa
p+oQD6i5m5ljI1Hn+Z90Nh/pB7IDpbNfK1zYpfZZJA2d7n7cwV9iAzGNcp57CgLzPMB/+RjfuTA1
NWzUsUW8+vDmVBCgVnkfGmoGm+qqQ099HyPqjI+O0bCQvro3gKpOlTQnpp925MQf999vXDXUSs46
b+bXDJ2aL9q2JPrWJDFecjd0F4EE7RJELiN1wIhIJqYo5HCmH3QmVEnArGZLlkNB4PqCg+i3/N1c
VYdy+hHW64ldE8U6/pTlvhOUsqGZT96prk38qSejrJ/EAAWEWqSz0GNGY3jwvpVWsdNQ0ktgXDkw
lEq91IUOCPM2ZSOKqbpU+4Gsdd5Le06I2twLFZb8qDcCGEl/2X5prPp0gShxNCQ6Cvtx/bvCHZ9D
ZUlcrQF0RumYFTnCnwejISV38WMd8z0KaAtHUYU7tY54vnVv3pjGSxnfEC+B0zD54vIYD7Z4esCX
ndzhey9CWS72Mg+KHP9fUQe0Eb5LQX8LHZuIZmHgnf1FtPcAeW2x6DMpWYkcDZn4/ccQXbmsw+9h
9cFGde/8R5kZUPnPGaWs6eH2+mkckaLHFJSm1pfJn0DmAgQL0sKfx6ERCcOunkBH7Fomjnk9mCdh
8t/lJuQdWWLTQrQpOJj2k7GH4XZP8Txb5VRT+eawniifV9HAeTopYIU9MKlXkMOpfZ+0Y0LRGBlh
SBXLvGQNQWnjmTGbcByutx0MVbkLPfew7fB3hieNP/ec5z2vJeMgfo1Fcgshg7DBqjP8WxGAQSBV
puqe5qJDGYfWi1mqtCCTY4mCRyKAaMGPfWd8cMa+kWwIFOQ+jNhP68XH4ivVSmO+BnJhLq3i58x/
Re2AxERANcsvyXB+8CGWDtKhVjc+dGj5zexpXs5UdJwe4mBScX+A5bnN+VN12NxZna7IDItWyfki
OYI7MnLkfZL5LBWIPgP9jkWpUuMcTW69Lb8+y6lkyNt1UsBbIiNiLPZGkW2Y/WFE2zqLWwF6ADeE
U4LfexQTWbmC9kPk1z3Ca5Csrap4d7DZiTcwLWd0jjLVolmL6dg7abFyA/WO+3aBvLvvzYdIA2I5
h8Dxq9FDugI62IJXlKYZaHUKa4RyCqXY3823bi+8FeIP1T9yJkcJMy11o6NP43jjFJEA3TDukm1r
fbnUV1bkHNRoxplu+ExIO7n9UP6AqZSxBW5OLSx7nF63yFnYSKRKtlsefbjwzHU+ynktRzhJWuQ2
mUIeFpHZEjT4x8R5WgvrTKfqg5eD/eZuztywCyx/kG+3XtsXuuEUZ5slczWtpJEiWx7ISnrv0JGI
ZptoDqBOxtoYh16LKMlQWkgfvz1av2BxuFXr2emOry0wPs/qfmw+ItIkVBqEsHbcIfK6NkkfSmNw
sdRFMbl0zwUyq+67Z3uDm7gAFRE5WTOfgTwMFsRLg12D/JfxEuqTvSIUGEofN4sjd888d/FLvvaN
nWf5/2gOrc1l/tz+fLgEI22Ug2ehdMe6DMMdhS4B69RRp//NHOyn3RG0mO6skUegNUJA18vhdhcw
Vboe4m7mzrPwhvODxQ5h5i0XExmH6KCvGSSRf7Wc8+uw4c1PRbnkQUBAxbQR6bLeUytRLWDL11ae
RkEQKINoPZBoQXiJVzoyQSWn3wmuk8NUD03Xe/bzFntm1ErF+dou20QCbFS4S76SntvyRiGQq79v
Ngjg2HfpmNZaUiSiRYEjpjzy15kCujSy+zQoWw84HC8Eyg2l2ODtS51lp+fF/j7/O+JSKwCrHOYt
54hPPve+r/88DqjVjTHiEI3b0ibNk7XHzVlUfEUk5U60rOn/82ucO7TIMLTC++lFOBGx1zb/QGsB
Z+u4F2rP5YPz0cLzGytd+xOYRV6Z6JpbffS9QrKzEx7HhcGS/48V1rJFXFu8KRLahWqXXmKv71Xz
xKVbw1PYyp2NyS+UPPLe0LSYscm+1ziHe65KnBQdH85S7+iQp0QKi742lWM+K4I+Uo8KlJRv4Jpf
w291Tmt2Ijsv6CrnYdUanNe9Lvn6VO7k7yEny+TW7MGE7rSnpyh5URMrYKzBOlHo+fFquAMyQVX6
+GS/3j7w8sTO8KY/8nodOpqZoASIlgvbQbouwzjExHYNNYaG3AXxoJVH1xwPwLiSPRtC2fRvCgjc
tZh2sX/vUWxH9merL7x12tMjOGYjjAkoZx78kXiAdkxEmoH26e3VNkZxNRqnXvSnZUv466BYaha8
ZUrdyTfY2FqUZz9vf49cWu/AHk8D++LCNwrF2wGHa1UHAZDtsoXfRztlePqivhekrY8nwUTV9xDp
xJeDpJzXJpl8faD5B3YpJT8kQf8k0MQep/hfoQjpKbEq3qTOqg3SJIK1ONmYXj19RiTEl5yvFkty
4CRJmN20Gn79+9bRhpIAgFccVJ7vRgsZlAfQgo6qmi7vo1eNBN/fCZLihc/XJlgxzx7E+AWZdSVO
uxjbIB9AsrjtOnB/yYdOjtIyaQsjYs24XDHqzgQ0iUOLDhWQix3ZWGW+NDKUFXYy7qsA44/xarZL
e0BwDb/VlHmV0dfd72uHIXO5eb9jtJ90WT6So1v/HEDjnUuG/noRYEnc752CFIcSEbszpkMDm5sp
kfra17BrGATOj52JcR1LL1/Z5YVOteh0i5WWzoztDwyLdGE3KCS6uxKOkYRZOnntXlGUefHi0fna
pHS5R5ysqFIBs78ybOfiBlKlb3mANzQqN9RDT6WAMM3O0JAIX8+AMFx3O8HjhxaGxgmC1ijDg0Bq
bKRZxdEaEewQr/s3s+Qabws2xmRNxf00c/tmcwbVkPttczCulhpmBaD2f/fFnzNMcaFpBeQTQblZ
j9re+DHVZKMOw4Vds0Y1gLLWUhu8QAw9Dvnb2apOX6Psde+RUgeQCnooj8WBBDOEHVe3FkyCWnQR
uMdYIZHrTnGzFzIyjetBGgJ8dRNtWoo4+LFoFXyBVGkHyXWFEwrNq2gJiq86yKs8KmVUPKWeTYeo
5Z+rbQslFyNLjGatPBeAKCjmkQor+f4b/iy1KjVE6TZDCS2c2aUQaElWeQOu6tOP8FpK7QphiKxU
zT1suuu0cH5RsXWJXMMFblGpAhwCEj9V1hVpNTl7T4Dg3/lnDI1c6VqS9D5X635UaqgPjXa1Lr1x
hSj5UzD84h/YscZhtSCfq7bTjUOQ6mw6tBl8RwGj1KKelFtgd1NU+8ahzntJrvgXdSHakFst/GrW
3t0U5ugM99x8LdQ0uWInxGVrBE8Eo+OoxQXLOSKdmiam4kZOKxEUlS9OZr2dZ18geqv8xAVqh6BZ
OLGQsGpVFDAVR5/KctQJg+a9GoWMndRvlLfWtoR13EZ80NmOHg2FNKF2oROGJIi3nfMlgLYHWIyr
CbyUaurAvVYlFLkznd8FNOtgSQXeWxJAZkdYIzQsHv029zLBeeoIyrL9mG8v0jSlIPw25FFrRo+E
Hv7ihDTK+qNNj5rH2RPCKbw9n5TGlb2eVGUpn/7e368tvYOxC1CkdXDoeKP3hcL1tBFVzOsxXSMi
FL29ntDeK43l1jWksefMspG0Twpv9h2pk8I++UvLi8Wa98hFJFv4rY6Z1dKX2Y8vZkaIUyRUBVfp
UGskTlCYGGGJZ3/k16N+hd8z3M7xPIGgEE6EYmhSICTOFU0kHAQgtHZTuQSlnDJAIBHV/N2j3j55
RGWJkyNx8bmlvzrZ0e+4rolwRltABYEyRjR+zuMbeb2Am8qdvVg4HQiHL3U9qAoUo3ozv4EiE4KG
03ovr0bU1lgEnuwIX72A4iDzGe/HpbuaXBstoEaKbQTrnlyGKG3FeEc0gFsivMcU+ZWx3LAo1tK7
uepBd6JRo3nNxb7NeYLfE9AmdYDXompV7CVraXcMkpkjWWlEIiaTnJphgs36qbC8E4ij7rSUDuKz
n9RbnWMDFWRq01SIzEdDi9M9TBT9OTqFry43eCcMJsenZf4i4pN12RzxRR2tXDyU97yxAEdFkdrH
ap5wyufnLDSSXU0A5d0++ER8rcPWXYhHp0YpN6cEXyIKSLINCpM1R/jjz1b/WRaGA8O3bpXqzcB2
DIUbWwlaIdsZJn5YvWixZGjmwB8q+LCzDIFE/+sJa1abhT7hYlTiW41Choyk6qeQe8UFrvYNrAzM
xph2wOM+EuTIatbIVdQlJxitpvxaKCg25CIAqTSpsZnjjMO5diVgzM1d3xx6r50FV02qpjH3shZe
7J4Nroksprz8xLiFxFnMPBi5lgAAbfEBRIJOV8HV+iSDT5AUCmsUk3oWMnq5mf/MZ51SssDNGLvF
hjhvGtXOzqA8v84NQ5Ab1yZZwUoy4Ilvm6ffii9gKGZLineuqYA3175F+7RJ0UYrYKVQP6OSnJKQ
/FK/7KI5QbMjGebUoCsgoY9KX3SmaWpMOet/lOfSXvjOw5Nb6+rt1vbnYzfBn43m5L+POn4v3WSp
czJaxYe5tspL5elgHD4pK6+xpcgRXercdtoV2Xym5nFgtWwxc56hDiBDPtIC5PDkJZ3+x4YRF93+
94emyfEvWPSAhhG/0ly6DQIZ948o1zj6XixX4pma1VzTvoWjrfbMVinoJeVWslc5UO8FYTHk4Zre
GfG2TrlbN1R1Upyt2VMYbM2hWwqaaptZqUn8PvruTET7j2+i9j+ej+JEMYTyNTbQhevKhDUp29uE
tdGTB97TObFa9IjuBlK8CSvpCg1VPXyKs6Ry7FNaCRUDLXh8QDtQNYVcludhidMrV+KNwhIwk9ED
ysxG8gtLD7gaKRczZH5eAbih1tbSmDDvkBiordpJNVfuH4ajMkZXvvlHsYL4Wvb/Ha7wBN5mxffP
4yDbj8fRzEWswdXIOcMcEFeQO/oHUr29H5gy8d1Xqg+7yAjgOh85nNYOhlalA91L73yUuhvIRGqw
udYcXicmuXKAD8DnGFUVUx1N4dtE9cnAv/wr/XeezgihAd1edcEb1S24JU1Cu3D/y3dxsAm5Z70K
ZMkHW7TourKKYZ90LXbfi6EuXNjz7TSBBTYWIkai3pcx361IW8NkXSZ+BtPKzrrZ1d0Sm6WVVH1L
pxbjPlQVuLg3j2PBvGRRGUEOpDS18uaDBVh1OTGwJmX2pRe871imqQCv4Vv9sMRhScvvzA9aUG4f
xXRfAvhMtqIHKs5PAQBb+QExAvVIvLyTgaQffNIOPWRa7ptJbU/WY8CwGzvlEkK5caNou5ZFyLsI
WVNc+qd1an7CevVJgci9fNcbK2nAZtPvsVjzir0Rw728i9IVvViiXx6eyR5ze0YrkZjqlAfWtnWX
b/OfQoU75Jv0M3FJWm/7axNmiW6/0medhVERvWGNLmAlWUNmCbnTRyjshg6ekxVUD37Wh+o9VAh9
OzXDeSX2BW4EJ0UT/bsTK1wUf8M2+YPWOntxBJzIfn4va4yangNK5MJ5cCvpSx6dCF9tjCTWDUuW
Rc9OMSxHSl5CWmAovJMHlv3zvTZR+rlOHt8DI1alXXB/xjOk0JADsszHaaGmLtr8ejP5F19djMQX
naHuaj0BDrW5yErCH/OveFHUrhKch/rg39IqsYNQsHjR1+WLI3f9vTMbnTZw0qLRS0gd/Wh+99W6
X1NkFj89+6ig8vgU7tVhIblYA7Jp/80MD32QuxXNzasyVw/mnB7P0z1YsOo5KWgcE3KkshLyCVPN
NTTI0qsg2herczDcwq9sX+nxfLqeeVw8dGejXneg+9mORaXcAgOfQqIZlIpour89qHjMOBNFaYH5
KoXAGLGiAbcJF5VwQNgksf38sWVfhRYv2MAn7i+o8MHLjXZbmW9tL6EiFVLGFHwYx7BhnNE2reAN
SNfNWkybRIDO0Otody4F2pZJ18e+Xi9eoPcIQx0IhLoJSJW2M8ulPceQMVlohsFMS5FewwS7eaHH
qCb39nlWt/STMZgg2MwKsbeHGkRlQoDcIWQIh1kfgGSg5X/u7MHqnog3ZtAoPcTFGvXdP/1Kp+Ol
R7wvkUOzHRINCUU8NeVwxrHoZC75qUlAxKnWAKp/WChvNOG1RhYiBQopXtgRI2lYiMZ+z5x+Wsh8
kINWy1P0P/BGEsOHKiXPQSSxlODKRNslJlyjVy3ClqEXWDBXFcMH7P/2Nxiq1pACUoMeNPqIAUuG
6NfjvCIt5idFluyAmE0sU6vIoceSHITBp+HgEgoqo7jWZJRPABgqaQr+/xMLbuD4elEiuk67G+7b
/xaeWZCBSIqUgxw22sRU/xPjsF2fBUUDHwpG39yrVh1J4UPXCZbIDho+UFkxgCbbcMIDUTVz/Zgv
c//SFbyihUuvU550Tl4OAvkVVmqVR3ghCoP3VAP5gI/V7lgOBoy18gSMOYwl4fftiHmZQmkdloCI
HoU454SQwJ7Q2D1kGcjZGYh9T4E6AzEHUZHB2UZ/Khp7gc2BTr2v3uQBWrKdmCpyKE0u+ZI6+zCW
9+ZpQFYb0m9W0Lsl+xLlXyMpsXkk3RNrfoYjz0dexbOF2+KOB3SPnImfB4FZCXqtcsL1m3oTLIDX
BXRR/YibruqMmuHeumS1VNpUcSBiC4kfVkH7tC97pUSZ/WMmmqB3QBgJRnVv6rQONlKd2KP4Dyti
eK9k8T076BrTxMQTDfkhiKA47KKXVWEZWmg/ow33r9fi1JbV3rWI9SQ53iQEDYI1qyUFIWFv4MKk
I/Y0wVDghyEvKCTPlfo3YXNtQKkRLemZ5gzACZKp+kWrLyTK2DXw4agrjMen+Q20yQGGVf1RlX2I
KKf9w/tGh0TALE6ZBEFStXussJKSzgGr4Pukq5bBXcLlC5cJItJbqH58s9oP0hpIp5qOjH9tf3ho
bj0FDplp4m2VZU3ikeMBOL344zHo1GgR6U2Mwus+GvD18v5VgCKNlw5ntkFm85Wzwye7+cvPjBkg
Ighw1klALKIu7UMgdhYvxNzsOizARGEEbuhdGW490Ck1Xeoejm7UrtmMh8ARYS+qLuLyYS/DF2Q8
CcIy+iHd+wNOWQ/QA/8mB4nVCQNvHy3uJnZRps7MsRnzB1Njfl6fS1wzPRb8WGPSYbKTEFP+DVpG
4oKgtYM27vRkqVM3Mqb+JwQu/PCfAD85Rv1EASdtM/z5iC0VwO/RH2+NZxhoKIP2H7CwI/y0vjUg
xwhFT8TKttscoDqqpHeaTkavEmArtz6euEi0Th/uCj7uzOsy5gAzTAH3RYYR20VEGR5/QiGg3Z2u
zBmfY/oEmJIlJyFboOobHv/TTu6bwdyi68HubUPiKx5amZfvivbmESgp7zZlM0c5oJEDsKnEH4mo
fkBtF0fVv3mlwnXpOhKsCdLbu1l1UMNShy6csS+RMpQA2qOL2fC/B9l02jGomOCIqoDX0xm2iVs8
pcd1oQaPUqRKtEZ9lhzbL7EK9zoyPeU2u9LfS7MhAGHyGpm0VfQ2oKDv7FC6f9NOLhwd1JIh2P3N
Gq8vuOuUCrzFC6N3qfchMkrXFcpILlIPcERlWvR1YvdVK9R5SnHZD9gUBS5O2aKvjzF4JRBudfTt
2lLujqdjIoI1sEYVlyqHxonUUa8ca1FmQybGbY+qFiEDp5jwfRaTh3F177FDz5iVc7tuzGpH6UCX
P2JqexFDbfLqHd6NL639P7+NQRjB9hi5qTiEIv3chxjzIu2UWURmPuqrbE6Y6Za/RhwHeTe55fw3
+WGLN+KobiPgUqh25jqXw9qd1Tpd2DYBxZ3blEz7HYCH7kdyQoKSUqo37/2uVKxCcrfD5li0pNiN
tIMq/6HTAdgcMZEI8CUJxNGQFtKAqosV4+2lUkl67BA=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity fpDiv is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  data_a :  in std_logic_vector(31 downto 0);
  data_b :  in std_logic_vector(31 downto 0);
  result :  out std_logic_vector(31 downto 0));
end fpDiv;
architecture beh of fpDiv is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \(FP_Div)/(fpDiv)\
port(
  clk: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  rstn: in std_logic;
  data_a : in std_logic_vector(31 downto 0);
  data_b : in std_logic_vector(31 downto 0);
  result : out std_logic_vector(31 downto 0));
end component;
begin
GND_s51: GND
port map (
  G => GND_0);
VCC_s50: VCC
port map (
  V => VCC_0);
GSR_96: GSR
port map (
  GSRI => VCC_0);
FP_Div_inst: \(FP_Div)/(fpDiv)\
port map(
  clk => clk,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  rstn => rstn,
  data_a(31 downto 0) => data_a(31 downto 0),
  data_b(31 downto 0) => data_b(31 downto 0),
  result(31 downto 0) => result(31 downto 0));
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Sat Feb 17 22:16:05 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_HS/data/fifo_hs.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_HS/data/fifo_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
FQW+m7qV6K8Sf35CP0+Pii0pNDbWNo49VzSEu0DhgDLMhOg4ikDtAjx7viGKMCB82oIaTpkHhCC3
BQarD5SGL+ZgwbvBgHZE4TBOLKMsLoYRcuNlBpbGm4o4Op2Yn2UHd1N6RTgsc5nyC9fXAXNyOg5v
oKRdzWHhjR/TJ/iFiib0lsF0JFveaHV9bGLk0syGo4B9dleAqb0n3B4N7eSUBTOrBmcbBjcXIK/X
C4pza2VgZ2TZEprFKsAicQRQypUkg5enD2CINOrAXukpCEHF7jLRgcQJW6Py0hWmHUW5Uhuy43Lz
ucPvVlGvrLXOxF1Tuj2B3PzwndkJyRaChjlB1w==

`protect encoding=(enctype="base64", line_length=76, bytes=804960)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
+w5VaxZCa1UXQ5eFqWPyg36Smk+9VDX8BNYrpiFeL+9ViSmg92TGGvYA7IPmpRLB8B8Jv3Ldk7Dg
Gv2LeoXFdZWeDPIMYc49+QD7v6Gtjc7HlhOkIl/t2UKs/0ixT4/pxWoRg6wE9zf2JjFsszfsPa+5
KqDmS+B6QP0/DSRfGZy7A6um9RRqhm2Kg5xlBluXFhW6BOMydUA/QFUsE+5Gv8++mvT1/6L6vNgA
hxR4A3bHRAZZ1pHIKEsCr2+mr+ryf2f411tSQIQQj5TS0oId42G0CXQg5qE7ZisgHQ3xczP1X3vW
+g+I+dnyBoxNjL6yklkn6qDnqO1VZanh44v9yy7nETKQTMVNRyyfmtfaRoTxbxhvRsdHKGGFjVXi
C8fyHlistHsi/Aq4WilqCyA7ITAPiuIdp16ZU90KDYsIbOydyME5ghSibrLXylKDltcEx3mkN8vI
Wfd6OyHmwhW5cMhcRuUqn0wBTAKPqJXZUvrG/Nlj3NYwbqSIF3d3oG8ufOxD8FdyK+uGNNjhhbC0
qnI0BMct34LkG0woij1EjEKrK1h1pNdH9A99zsi+Fn2fpC14/LSwhm+lJsYHrMmeFACWk9b8sVpt
ZFQM1h49UKua7e3z21EseG1iwSTyb/EmOCes891+BRZZUR7PpFuIAaScksbmv/Xjsl+6xiEBSMMQ
P6iMbJbnJS2IkbmWvEydFq8HuRb9FKgBl7t1S7mGN/nLhRUw7Hg1p7s9707O/Mteee4SWT07PAKw
FqFwX6yFyuPzY53F/+rXPEMjwJYdNIzMD8nmTNnNyjgkoVB4Y3GCM77Uq9ddWGqntKVLW+nhjlVD
a88Hz2mmkyuIRTeuUF68ZhiDl7bNYq6payUbCGz1s8dzTOvS/vuq91JX7QZodtveRBA8WsAyhlM/
fvLNnxYtn9Qitw6Eg5T+63CsjOthrMeO50vEsnp6pvKZLnaGIIhwpHbylQvHygROBGmOKUiNegSV
3TDGpD3z1RSjMZMxuCJvXDgQlhJGGj3BTExzAM9xFnYhRESo9HMroCpKrlzFb+stkWZi6ij6UvWR
8xdUtzjTkleT4TKs4iNyM18UXuwBaLRsZ3knENi1s4fwLVEIn9xXughvkgGB7x/rh2cSYcuBSrrp
mMb6U9sXMsbQoLkZpZMyo4oq8MxVt5+dg8yM8jhmc47Mzjmy7L4r66IFa5Zc/lANhb17dcFq0vVz
F0YuAfTTTspueOxIwIwyPtfrwwDWuLVp2XqsEnN883BE1SInLcFAK5thc7mC1J/92RwttiGHfrn/
lC2V8vYYJ476IC4AzlLPgLNVau2CBxN/ubl1YgQwBQ+xf5hDd+e+ZuDJiqsSljjz7vdFwdSKnYbc
SHPIT9i8r/rsn0yulj080izMU7P5h3AEGttbHVSEv55b+GV8SdT1R+F8cLrIotaTiKEqxEYJPijz
Y0xDIr6WDMCw/KUeqm+CS404LespcQ7L7gex/AkcVUPFG2wmvs6beiwWQkSk8dCO1BEuDucjY36o
sPJLr/EcIskJMfajKd9Z8erH3/kRaILax8ac/y8GILOu0+zIsOuA2k6qMNOTULYwNGT6hR4wwzkV
FlpzK1dh21QHPFuMjDM2BD+W12ZZ0QY+Uwe6eknByAorqKsaGgLLkaGZKocN9Kf21ArP4o9XNGxM
sce6D033FW9xRBFty5aYLHVuEFlrWZmmuqckm1BOYEyQyS0QQCB7oSDvygaXAHOI8j2IpR/px6Ts
D+73nySGGIDw6WkYQxATvY6BICX99E2od/SFOLQ0daGD/DAG4omJorWlqT4g3P4D1sx9SemvvVgB
JafyoASZXQ6WkUoOGvQ3zgRVthhBffGCDQ25pzOkRshht6FdnZOTbDoOTcR2vtCtuhXolwffOQSw
m1gDA/piL8lOYG4KTUd+MtoUa8xLkDovcKYTsKd/i8v/0pe1Vs4pCBD2YkKo8yFGk4hZC752Y3k4
QWwZEbXgBGuGp/Nqva5bWiWeqHN6EGH9PE0rsLDhpDHUxEOqilK/r9oC/ettLQ7yWtXHEx0D9QLq
iyKZUU7rUjAlMeHtwCi8HFLqDE2z9BE2CxzmdbpFE+ZLjyjtcoNLSkQZGADZTY4JecLVL7NicRDT
YnZv2UFb9ZK3S5uxv4u+iqvIOzK9F7F8J/JejLzSOV4YiomFwecfWy+8MmJqg4addel/HNH4ntvH
8ismhhXLfI0zkdREgr9JWijkHGJr+PjZ48N4ItS26z70+5+NB3iaRSO5+FZI+KS2xSk3rwHSJcQU
0l5DytoNk311ZF/SQfD+C01xdz4di4a2KXCPqQaTmI4t3fwK+6A7Yik67WSQTB0E87FZuMff3VHz
+sbDFO3z9/vVRAzh8eMXTAtbkpJm141u3H/1TbA5d5gLIYB26bMAmlKgNumO+DbpabkFHraDeunD
Cox4pWVPhPnug1YaDI2nglXmoPYfq7QgYiYl8i3w6yI6w0lUFC4hHutxo8eAB53Pc49lQrBR3OOV
E8tt1map6xLBBqwb92X7RajwIis8QK6R2ofVKCA19hXD9Zp4qbfoa72d5uSYAVnJRN2luLDsSxqp
YqQA3iVRCnaBVrQKNwrhr02dIVAvzQjTrwEeJsLW4jUlfVdF6v97kJP1LjPTruaUaVrDfDeODT4N
Zak6HyOZFbifGEdLN/zd19fJK40kjm4IOMsLe3QL5QtHG7K221AjY+Srue6YM5JQIJA9+HMPml61
ZJSBOR3vOQFtpZp+J3MnjXpTlKaZ/cAuhFTBSNrRTjNFpjlboKUko+qIwKF2a7GeBJ35LSt+teeD
Bmfkij7XTUYrYT3wDPcOPt8q6WXwFxFK6xVwVwEe/pISb9AW1vKxXY/DS+Z2IuCbF/nZ/Fo39Jl4
5OdTl9A6viyHcatEu7LyB0S43HqNF/NVs28FWZsV3xRzsCF26lEtch8pQs+6rc56MROcpztVuqRS
l9l8StJD8DaolMdHt+rYrDUUZAOX3hHKZleACoYNIAnfgRaIaEOPH2BV3yDbwnJv9F4fr9KxciZC
59j/AayTIhPTmqlGuq9BumKpVTTokkQXu08G/I0/FvZ8ahz5IIOPRuIoaby+tzoZbDlxrTCPSCGF
un66ShLdfgQzwdM6muRQlP0P82vVQSVHpPoJAH30ZHp1a4kVDo0Y5+PWKe0/M8/ok7P5+Ia6z1W0
/hnDfykj3dhCQC7G70VhRWAP3qC4pM2UVfSdbsc40aUD5DrjjDo4ut3klIvi5AWacOFFJuGscJUW
drBI8mr07pkXAhtShmCs+UI3R1K+iaU7eV0CfaJIcDNfcwCIBXk+Osk9Q5EeMKaVrrK+DTgy5WYN
OMHIHKid6GazZoQ+1y22n/QHUFWQUFR6S4C/EPf63/w3eCGF3zAgj+U+RedPeBoOLHZaBPL4+QTc
gR8xVtb/LeP9k+jcbLdUkmKwTeJeywZQmso0IuBBq0tqP24uE2GC99cm7LFNxyC/bOg22sbVAfXI
4QWXz5KDK/OOkatd8JHgkKYf7X6DLyuD9U3830GuW145sdzlZ46oGrLsicybTht2+7dofqeosOwa
40C8ncJUi+RyIVTB2Ngo+SiKo7NnmmPWkHyKAgNb47ZDaW9aAaFyPJ4JJh6ZEpcGBQyzX8DY0ikQ
Xrh7OEXYYNRAemv8Xg5codm5MQ3at03e2TvNJ7cC0RwtdD0LZ8QmDX0xMhLaWv/UI/xStRPjhgmv
yhw/C+J066hTUsTyyXR/bffgRb3TR8YPaf2yHKQIirnIUIeMNdn17QyrDsqfG+K14/3o5P1Esuf5
sckL8c63kKurDiggPCmohLscCitJt6Xsbh0mKTuxdVoOsvwt70hMVTZkWydKZRXB75FJDFaYgycw
SDbbh9OPkinJoDbWx/XfrYIYG793ypnLWYXtsG9mC0AEIJzTyZqqSv4WXl5z96Yf11GcpaLUBB8G
7QWeu6choQ+rxMkeLFtRO+hwWVUtjik6seQ5XVhCIUr3wrhMLVDSArhqcYH5lTNjyXcmA+k/jiDW
lEbJ0dXy4n1IpRwW1+Ak7KbYicW8fzV8XgaynihNiNY/HhXDqvGmVe2HYWx4WmtULxz6oaPPyhTK
UoKixM34XGWZ39UHstUQ9MR6DTwKWGzt5Si82oWIWyiq/9nGUvw1ffYhFewI92RU9NxSRI+tu/JF
tI5aZ5a7GsTlQ0/konoF6SGdW3kGymmrHXD5DCkUcnk9aDaqSjZRsKzo4iLu5sENuk0gGzr2/qLk
//eDNQV7jWeLzqI1oEgrPBKSVNko96JewVj1zqlDyFMjJrWxLn2kb3XQVm+apgzjE5RVpUr+1n0h
+Dh2lUhKfqKspFYzTr78dWd203WtyZ8jRpOILJtTqCSWUwwI/svYRmUM5Rt0CSskPHd8NcDamAF1
Yqa8ItZyqJYaSEmJEM6pNHd/ahfbCg/Fy2J9Zqxp3MzK62t7Y5mRHX4XYKRIJJQsvnIxvhuScD/t
hb+BeXF/46DD2rC1PnjM27KGqofxRdP1KRZpu0CZ8ohUiqEemGzzQO+bfrY9lIF1SaRccOrKSUef
6iVnCklPykNjGvjQXnsZPH0183tJys64icc+YHNkufTadhPPIe2wmAFWVL8AOMB2007mMZkDP3cS
EBCQKxGG6DqUqlpJgpYDhQCqPLbDDMZJYt9YUSj1E4pMhhiT/UaIM0J6wV2CEOWTDT/XdvVDoKZ8
4ctcY7zqe4klqO/AJ3iZx0eHzaOjPYVOta6BfEcIrxbDucKuqgW6jFa4t89RH+Kc8W0jG6UL2o3n
2sUqxTtMuP8m96XYFO78aKFxKnqBI3x6N0teS9k+BIuU2Al4kXNLuQyKBoYQwu617I3GqvnnBf+P
X7zHNyvkPeeCN5inR+O+E9/I2sPqInc9ahs8mpg6bb9BkgLJDJH4F3qjvxDK4aHQp8A5kCP8rJWo
qkdpI600jj/dHEFHWlodR0Ycty6cOm0kq9jaEooRoP/uYN94dmap6oFQAr26Hv4lnFKfN9xaFASF
V8xnRs/k1Wjk1AMr5JQeJQlA1zFbmEnv+Wn4tvYFYGiKm60cqRwmnc0rG2YVu+kVw8AxXm+VxvH9
S2ctlA0034ml0zX7iLLBH9pdqmzyp6CClarSuEGV7WIr51qZb0Zm19rXP3eX3qLTNAJnmsGAjdzv
Fe0xAAOLn82Wz6Xy7LxSF66gGeCM8Ud4N6qpKV0x9X/fwyVH3QpIm7Y6B5sEr8Wwnp4Roys8zr9T
PN7Y+w/JoFXgdMVmhhpMK2AiOkq1jiYCQeOxbPNva3K1A/Gm1i0UtHfuxq5yE3RKlLObC0RLmaWZ
hu2nuTvuavmmjHoxME6HaDcJUqHJgYShc0u+r46J8W+kWP7VdhYviCuXIhTS79e+ajajIc2bbxQb
okwgTGFETFStHCv6MvRtwNYtaVdNMidlxLU5gKxWaImofGxWUXRPs5an7gVXUjygFjGsethAeyEc
vndOGIF+ybHWpWMRXNd9ZuLCw4iVy67QYu5fg4KgyJnWL8RmUBNN2SgYeOKUUevwykJFkFgzPHxb
DYyQGW24WHrbkP4kq+Bt5hkzLMXqRK2u34zhgr6mX+vVofKRjmqa4JOj8/G/USrpgIILbKRPoCzi
NS4j4cPRNfv+uytLNcnvmghV43X1cTx0rKrTex/VL6JKFaIdBD68MCmjZScP9s2lZw5VzjPNsnfq
dH9g7VL4GOWUpx/bCamqTLjEvLRI9xWqTI5Hpg/SVsn9kRBNqBtmoho/ci6KAYwY9RJ9uo0uFCGy
RYsh/yD3COOCvWgw4YyUokWcgo6/3UfKm77knkhrBHH2iwsfohZjRpxmObpc3X0y5IoCsGhCIeNj
34fMJrY/2qEvYC8Z3PlHDTvfx37TMYeOYwq2gxsXFJmbZPRt+M0wJ6Y47NAjW+fjMkg0cNeq/Rlu
oMyX+D2lfL1xsOLuDmiBAkrt4vSTmDlXC2lqhDxPUrQDgeyrR18Y7QpBA861hnQetyEuE4Oyl+Qu
mtwJa+V0F9Tb4dokycRGyzn8A4xc7qvz+PJvPfRAlQoZkoKxKHCPBcgVdNx8h6xJCCEJcphrn0WX
po5SzwTQj3WHOWARSbLgudpRjnnZOKrPVV1iQSXa6lrG4PDLwwKFlGWN6Hokvw2XvhKeBLHYf3wr
8eN0ysceX+y2TzgvELkOcZo0avBvFo29X29O+5ITVC1It54YH5Xk+wfpchiB2f+NnP3v+EPqI0oB
6AdTP23RTeBJAvfKXfrZuNi0YhSiIv3NhEMZQd1PUxAMS4rChNw2QqCg6OLOUBy0FA9hRfHDf9qI
EfPZqP+O5b2u0dTkBmPO8mPl9HwhymOQArtJ0Kw2jqP4d8pEXeYX2qwA+shDmTqD2ghPR7EVRoLR
rn98t4ilb+JGzz4wDrBTxNTAsXBZ7+RzNtF3BET3vgJXtaZg4Vz3AO+TVc9AwWJxW5PcE1rqIWuU
B0VQuBL7enXptTjth0BMV4w0qt6mVnO5xwFDTj4kQzItRUAjxY3ijqbsBj5cKI+weHsE8DP2kZXx
NjcjFCJ2/+bS54eJsgGZKQ0zQzKdtFm6SD5+ZfAKABlKssBXonXsb4Wgc16PKlao3d0f8px60DzX
aaxgiiOS0rLYybHDsBcPHIPX/TpRwv1w+HBMFmrR6ujtklMAYi4QsfydyAMyqPRpcQboGfu4CsrQ
adFWglTzZhb99831FmwW4C5S8XG8WDyf0vMNQ2nb46Cs4vFBfwjzB+fWAcwFrZvHtcix0DqHG430
mgjexNSVIasJesnDKnACCbYk2+iVFowrLsW25H0YJMcE8uHXVnZWiH1HzmTGB1CELBqogV+HokvC
bL90sRaFq7C3RQqx7obYOXnt1awFGnRnFygzjbRyW+PRu2Izsw9El5Hp5zKJtJjxHlJNFw5V6c0q
yCytMZUYtOnlS6YfTGV4+EYHY8WGW0kbGZWC4mDSgA5R2hx9+rSzwhcO3+9ACOjUlVNFwuaDhIqB
8ngy6+O9Tdx6p4aHULvagMRHeOY08oB0axuUyOm9a8CPfYiit/tOG4+MkKivB5wbW792mccwtbTL
3HseN5aot1eYNfC7E+2IbFeWhOAU+cjanRaOo5hfTpkEMyw6P3WPdDiTwHOJtktWlja/kX8vbdmY
QvOqqfmg8VqFuVrY9e6cZA9pNRnUc4bntyCRYDb2eX8H9qlUMTavJBtyvCZfyeChHEhLZamNiHfc
+XlEunNN+C/gg/cxyjUYCzbedP4qGIn//q9fAy4HEXudFa76rGsDrOZjQhC3eUQcGlGBxJSF6BMM
b43LqRte54WHZUdMbXvTVf7gTSf8gQGq85xNIi8zy4Sq43DGm/Spd6c3oYD1YOVX/yB+GThXnHuH
Q13an732hLB4D7z1WWzbBx2d+belcL2Hdq3Tjsn9YcshcCl3sxSSi47gKfBUXaO7B+m+vxWQucRP
rPRnILlS2Bk7QpptOPyl+cuRiyflC1xt7r/2vy8g3uFnRBI7zGyf3AQPQ3lvJjCex8flckoijs+/
wrNQl9Qf/GCTnGcVWVBYsjUzSH123J327IgP88AziQszptbvGtrQHApuw+vftjptMQrTMsmyXnEc
QolbimZho5trLB6FQU8uUW7WWRNcUILN8x2STKtMamk0lHFMhBJjAO+YZvFq8oK9ORPuGFwrGGRX
7KPy4f3FlnxnvQtBxu+v0CtpbPhTSqIxq2saEifdNMCqb55IZ0g7AvR/voz6mYDJPkYpf3iWIDCa
mhabCdqXcDnfU8Z8gouTOECskUe51vYvbz9kSFKiOJxaqqX0KiiiCcaFTomZ++vCQWdL1w+I6FLw
s9sqS+Rz5d+OTjctelSQ9F/dfEMZ6SpscUDSE2EPm8lg+hOY/4f9tcR+u6N7ZTfWLVBlNEgFpbaH
xodW4e1FNcBifXrEZ/UzrJVyDcJnOezzyWu19ZyxE86qesSNxnfa16BWPFhCefPpuE+6YLILz6Yn
EmKjgolRa3k51UErrbfWFWmxGFACJnu5BKoyLunVitDBVkCsrBF+878bPAfmNzVE3Q6v3D1nltmH
LUhbXDa6V60cTJnqIRbA2GWrelIpMhXReb3vkhxVP/VdEuzfpn0IxbbUnfDiCm/fDvw7qrT2Q1pi
/GPb+H5k7n2y4Cx+dGLU+yVksJU2Di6uojka/yqRZOCJZPKfLfUuN2FAMupMK6Hu0pJkvaEUZxbr
DWtVUDGpqoLqdw+cr4JskrW4bsuOk4zUyIGIEW0BYIW6V8zMhuNZPnX+NbRdNrEVipS7iGw+LnMy
68rf6GRlKjA9gJ2TUtyIKULGMOXtxaB+nzboiYdR293HwVP8sWuH7aRRxZlbR0zZ6HpPKTtoXMsk
rh2OWzD+f/fB6Og16EoiNwqWqh4e2AC166UPjfB8LByl6WMtmFmfsJQ1t9pCEjiDQgu+8kfAe4bD
8/LG+NB5Nn2C1bJw8ohAybE6arvZqxnnZiYdBp3IpBPvajhf5jZtUmgODxUVp0j2B+igw7CB0aYn
zlpXZPxkGhpNXji8lPFsV6w8TUwC/nxZsm64uYXzWLqblESbJU279vtqx/sP+ygUfOWsOUH1Qq64
Teun58e7IW7QrMaNZz/JxI1sWPB4Pk2eHlNr5vA4UW3FPbsCdh9tQQKnP4mKEf/UhsJoiuaX4TGc
SgrfkPcKvvaJHb8OR59J+vGeFo8EyXJYjT3cp7KjmftonDHH/ISy/gSbXxIRBlDKddwbt4TraQnN
+HyeaY78ck5qxMht7Qeb6lGr1+QLQP3xKAWLIFkiZbddrqqPNEF2ux0wsMPw6ENYrPr030UE2ANf
WQjbST/zWs2J+eyp71EGTGrMRD9U26PW7eFK8sfe/rCcru0lCqzHkO6JLS2LS76g1EMo8tilcsD1
RyJRteFg3uvUsaWQF2on1m3vJo/pZokFthxwXVQCD9kGMUw02cWkrroyTOh1cs+lXG/7sLQiUZw2
omBGAaYDda1CRPXS7Kp6TQ6z7Gcnii1LnhuGJOHoDI2PujfennOqWcJP/+BVbDmRell2Vf+hsvhZ
XFOLVBprVzKTqjBmIq5PwIs7dS/6Xd+jgW9vTQYuu1FAloF078Iy27IG0Fl2ymSeyrioigl+Bgqg
12Wv8awTV1p0TjZ8VK6xiy3IX6uI6gKeC9puG3QeDdyzqwGq5uFBQQHF/hjLv2L/A3bd8v+XzVFP
XWZLkKWZnaT2zM3xN/YREzLzAUsGaqx9t5mGRcY1O+YMYUW8Upmw0UIwPQLVmZMMZ9rpxVigMNID
ppZs9tfRtlo6wuE3Kmo0ODK+nvip409yl6X23ETNotCN7/SAgM1fYTKh6HIHgoDZn3KskeFAp9Oj
ukbtrrhhTaS8V2atFFAXPKmBMxcnxVpN/EuuQZfCuVWKfGri7YIgEqvd5PN+mtEtjzbFBS4F3u5E
LAre7u5vLH0BL2j3J4RCrV1EjwKKILbgQDLtPFKoGbJeBEwayXpOk+CTftmd5moWETzLKL5Pwsfr
b6MOFrQ2mOsoJJDf+/04SS0GkQJolYmS5cgKvNs9P7xTR7c9yZjYJhLRKM+8+hYo4Iw932yUzulU
LDnZ98ooxMZNvqXUkaDijZdCOOVqNt2hgaDavhoPdK0CIrAUWjHMglNfiy9EgVVmGGpiPOjXCZfA
kuFKk2X5zxuoycVt2Oow24/BKyZpcOJui5gk+I6LGNoJvnbc2e0m95k+i3xGfjTYHf9TX8DDmpvo
MkSN4VJvn/utYYDHWHVChUn21si0eoHrmWpe5jdIIeqM5hQyXe40e7QwnDtEC4Iizn2c8Hos6G/y
bcjb1Nz3W4oHRwCzum3MVOPPRq0DA5ui/HgjtHsdfavINpdy+jR4XnbdcIPn5F9GeoGWzt8feqY6
2TQHPaTQOcY1PKStQQZ+vdxlE525RE+zQc+bE3yswwZjF/IFlyay4mLaAkX8ltp8MjXattYbvvd6
0zx77M/vDHqJG+f7Iq9LmrEd9Ta8EqlAlLf3zeQHfJaMjQ38RpmZjYfopaTIa5OYoWBHoHBWKGhD
0xfy2bWG55ozcRRCRjFT3vgPZrhYryec7TCoZRtzoeWPS0wzsU9K92ddfgeIoG009lbIcmD/VmT9
qmNNzLCI4UF3wtCTTlvVfvxTImE2X4jLTQZVOXyuMBO1ajQ6Ju6ebxVGsOWbWgCnG4XMo0fwXNnD
ZhJ7lf6ij+l8/qZaA9DisrnNcERKg4caMEkbehw8EnKfDz/+3in6+lQQ+tmIEGuEWPiLX72eXZep
7neiAr1VKl7NjPFrbO74PqhgXELUgYTHlYGVNzlezydD8j6sQk+MLqKSZM0xOe6DB1ke4FNz6CPL
nzcGoHjaGajTp/aR5cPdZQh3ue9LxbDLrr8G0Oi71DrV/2L6VfUgnHA1PlZN6+BOdQvGsbRf4ycN
q/73A/h1WcaPGfDbyP7PYxMFCvwA3o3KWyFHs9QWuKnkHP0aibu9L2cXOI1vxpK1EmLo79a8hLbx
yell77hoHp3qvETgSaOksY97Ghv41Gzf2seXdc5BMm2iRD5MwD1R0JTYOfc+dUfnPolVi+cn2dgd
YRXRQNviNpJkaMU3tdtUO+npKwtO1Frgtv23ykgDA2yUZdetQ8vVqUBmTH2KqEZsYcXpqyb4AQ1x
IAWKS6Bu3Shhofr1i78shPyPlnZuEPGyzN3K1ClNyaKynma6IpwTfdl2r5f2Z00Bw/DQ3AGQJRpo
tvS/9y3EdaV0KtBdoKHs8CNIN+PK4Vc9vleblB0MKQ0och2EEuWAqXJnPmSr86pi/fDGMGP9f5sm
d0pmXRjncyI/gteDGHnwDwtZGWe8OUPScgflJ7EUMackB870bS+KNoLgl6iab/YRPt46uPAtKGHK
Z9EyZI8RrbTIXYR8Ir08hdUOrqhaJ7kIJOE826lHqjR+LkkD9oRyyUt17cI1r/Cj4q2d5hyVTHvB
K06nGOaPtXZhzz4X9+dVKmqKuqt70Ue5dIAME2aoI5jjlNCvmSIpg4S6sry3+1WTm9z/5p4Bc7dq
wxVm+pt18lWZh/PYmcdxZhgt6fN1XcaAgHVvXpjoNXyW2B1TbeLXv+gx6DmXxvQJZNf0bkwzO/JD
0gcxuvIBl7m26zgkYHX6ZnadmH5OiNP6KVZOswzf4UeUMhuTh4o+bNh1lwD6NJKmJVDNwdq//wWq
vh2GMXHdYej9X70AGPXj224IGKnv1AhljLy7i47710mS2fROQEFBkJs38byaeqigyaBROPkwnI+X
Kntafcrvb71Gww/XJFw1BW128AfOLIdu7aYFjXRodyymEN6IWf4re2diJyqzw/wl0Wv1pPXCdx/i
5R037pQQKHH1pgSkVWxwi7wHBonaYsNr8W9VnzdYBrlFXpLstlY//rTJ8ka/NosOU+XsOenFS/t/
W2b8OIb5wu7ExzcTYNUfeAIAprMDuGikmAb9hBdJ8bg5S1vcapjUhb3xKlv9xxFux5wElS6tgQMq
rZn8wUaeWU3KfbXv5g/NBLUEt3llYbFV7K/jzdFNxO3j5b82EelnH9+HvC2X5rmUdu2IKowC5fQp
ork6wC3OA56Xu3PA+573/o5hb4CuO8lbC8ZB0wlJqHsYtPg2oRCIob8jTUi8jNwX6A1/VUr3Y/o9
340mNRHBO0aTh2gDf8Ca33yA3ibSCiaj7vEdfdU9oE7F7sB1bPQrdbTN+Rvu4a5q6xT4+Z3NTLJ2
j4eazho+aaltvVB4y4DGcpzxzm5gY71X9b1ouEyD4RVYH+XYIQ9U6T9/sSruH65tr2RMl/E5LHrB
UhxLQIUlDDizSz4FgcwW0L9cT01DrBavuqmdLQOI8QNx9BaUDL0lktdXZp7FUN/QwSulq4IAowzr
38C1Xnba2u5CxadVtIno3Ee1N0//kJ9JTYszIAHEI3+bVFqjOUktb8oq/jTLwxRUQnB5A8+EieQX
uJUzETPetU8hjF2mxBDr/lppjJgxiT7rdhTW/RU3JPPmMqDEaMj3F2IBD8x9ZWMLCUUFRd/qkPNc
LpQrcpzrcdMZyAZxd3k8lE/dPA6N4abh8V9VAibPqCACYG6HTVLTtx+GbAFM+5jmVQ6ddMNfmx1+
VLMWy3AS56mudDrOO2AAEUPVSFBJYa5T+3+UoTNJq5ZkNf63vn+fnrdFzDMTns7VqzNpPWx5cpOm
U/XhiShtoxA3GLBaU5GcIPAhkqTxRXWhXfHFs9BGm0a03jTTsSbsmdBIVOe0ipwbLKN1BMBFIqKE
AkKZhHNoyhw+Pv7cbF213F6ESerKXc/wWU4U0VEuturhbSbsuXGNAzfut1dYRIgYFyjv/duMVGma
TOxYCU0MK+muM/gkRTl4VlwgWFUbxZJPIJVRI6O+fFEtXcaMTq5WIICMxKPevesqTBZmJg7doZJM
Oiy0SGlzVH2FeWjIAh6OPzuMJIWBnedBUPhocZcpgb57w2KQU65FZBYkpq28qbmGcTtauqFqIAt3
whZRVwB3ugSt8p7/Zz4xF/dYw+/8RHQpWyj47MaETdMezBJLaR3P0ghJpRiilzmFEEPZkYEpjeNZ
Yb3iWihOxoJvzSld1EoMZcW26m1QO6fCxG15XG6lV4TiLbEwR0l1vPd7o1slehkXaCc5kNwEB4hT
hIK9vmBTVPKayU/txDTMJEVw1bHzWGZ7ZH7DUVK916zxXOABBGvZD/nLieDdpCUXNwh1E8/9/R47
6fEBf7OzBtiK0CVhgYRY2W5YA/itGJnbgK7T4YzTjDvjpHFPpfxh48n3pYF/SeCH9BKOwf6ttMb4
1W+MBm43HvRbGg5jajW4bPOYXqblp3WauqKPy3CO8yk76eOPcULO6GF//CS3IV/vJeDJxhL7U73A
QVqhTSV8TEJMPCSU0+SQ5Fz+z47NAOgUVPcckH1E00JVrFc9PGO80iSe5cKiQiUiKI9iNWbyTWTd
D4t3ubvxt98JSZi6XE1WC3fWeWew+1Ny6iJ4Biy76tkke8zzAJSMB8fFjFEQNxjZxtIv8idJxxbK
MFgWsyb2Mm9OsvtUADxyCDkFZ7+SM38x+cmbXbXMa2cVnrsH5wEOU9HajrskmOFHkBeRXfA2Hvnm
+mU3lVK1oe7t8PBm9tUaMJepug35tasXIECC+S4GC/LbFF6w1ZKYZE/6/8sGRZIMxXWtddJ+rZo8
5LuVXUTeCClzFdWjphq0LlD6i6KBrYTqy+tO61dLeewJrLjfJ3AYrrwJS3z8Cr3G3oQRK9tGKBYj
o85xLKiHeeS6uSXfKiR3KuXGjs9G4uWziJbxkKYQIdaVS79KCsxxpENTekgRsI3zR1hv5Hx+0tzX
cTg6SnpjedFWgnv1hpdyADBGrHtjlka8Kt08aTM/TvsodvEgzAXsOqyNoPeuTnBmeRHxC5RbEmJ4
UKZbHwT4Zmt7HD4JmnmpzuoPXzq5T0VeWYIea6bbjZTyCLRA82q17CIVZfj/qjuBmmsTXRbPbzbq
SXAPMRQiN9k9wPEPX8DdF4WDvKKlS2WWo4hXUo818C9uvAPvJa5f9j05sTeUzzC+DH4NDSlOWRrT
lIUNUh6ybZlbnQteVx4AZfi3PZMmYzAF7P3wAq9F+9RzjpkI5tmnjn76ICXVzI92x6uzxRMuXaxy
l9EySb+HMN7qkQxTQJB8jIbG9KbJX8tThOVXOv3pwnIgdYkHQwiX9u1p2pMQgDezvwuqP5VA+Ddt
HDlGANJHVlXsm+LPIX9X5I3aWVXK0YuflaxMPDiViRcI63G01oag4B96+hLcTXXr2pBEgm6FPONq
Mp8O5+1QBJUoDQ5g0Oq2+YXHXW/XrQOhPMzTFVXFjHtCyl3hmr9OvMVVB3yg7Ilht65GGEFrzdKS
Rp4qVCU2BrjvPX58qzsRY2FkT1Gg+C2BiKeuVFw2JOyScNZ+P2YL4Dv30/UzQYFYgoib76SKnHa9
xGB4Aaz23ypabCKEM4tS9pCZMbh8DUqFtIXKpxahOery9AX4umSTLwy8km1xp1afNtiR6MIA+eNJ
EKGRKAq4+d9gEoGqWTV7rqY0Ry+ZRPkvvDKqoZgJy+cXWrPkzKkEXi/C4FDQFv1NbTICLfk1ggks
gX9PGqO77keGQL5BNrEhZnuv4+iCoow1wnqmDtHRxZUfp9ItWcJz3TpXG5s4cnHlsmnwmua8lhF9
soderph97lkeV63gj4QIS5J3eus9fJNMviZ0omG52sjQU3l+Uv2+KiD/5eouM1ydW31eSC2OIO61
lpqQHUoWR+UaPcJ4kykWL3s4uuqWdtvRwgT2Xu9MSSl19szeDAdIr2hrgau0rAfumEh3PhZ/bxxQ
34HbNMpT/H8XFro/pNMvnqHCwqK7tuv37UBBWFW5D/anj8TxO1aH6fgPMQwSaf1Pg/rcnA2I/UQN
s9SoBR+2hrIqYwH0dq0u4cEY2Zp9y8DySCKjZUO9WAf4xLLTafI4Fv1nYLs34urVO2Kdq5bwbkrV
DX0b9/XOVUadDNqTht7HHs7DkL3XfAw+0uTsomSIzslCssw+nNav83L5vRdvM7fAxrTi2QKaOkqY
sIsbHpiaLjIPSDnRpuOFflEBzJ23wacUUq3lRPiaXrRXugtFmYdEaUnk7CVytBr4zuB1Td2Zx+uM
rmAc2PX2R6A/prZNpD9+kuzjCMHCOjHXYTozp215u1FHDnc8hIqVZACZX5ZCKgVMBUkqc9I4lige
4bQ+8sj8Tae+R/NphxvJuJ3O1xmG63mptiBVBdhhJZK1QubBiCwFhfLpUWeE24gdmw6Q8X0HS/nI
HvlAi8gX8AQeOWNONLuN5IoBucpBbyv0f92d148ctZcPm2TpgpkoEFKaLxbSCM3GmNIdOPeoJAvr
RdNqS1xH/qEj2iHDVE8zjJhvQn965xI4WOmuwHJullrA6Kf+y+XEXLN29pklupvvMtgifZ2UNPCg
mcKl7hfjn1RR2LtR73zMSf70cez2B435I+id1bhFcK63fYg85BO/7b9PV6kXNHAHyH3ak6JZZa2v
Y0uQ1UuWc+J7QofIBgRgo60X2vWBjYLw0pC/xz6O8i+2xWd24BSdVJK8MTv0MFOg3YGRcf9h/r0w
bgTYJSvmS5Rbutf78w+r2cmRBca6VEElMq/WyPfiohi6Wjqhf+XBGFjF4eCkwzhuRJwtUn/Ut5Ds
/ZVl1teG2EAiqxRAZtiWRiXFX4O23IQl9pzt9/CUz7PF3bRZqmMizuKJA6xIsndJhhUsp3vDWpaP
ULl3F1+1KKZLYquKIJkdQWUDdWJn9bqLLHmjH1G9YW6M6/87Keff6ujJCCcvOpvzTCUoeiPhyQOt
QNuFSisKlhpxJ9NspxkhoXhhnjSAuXz0bgPr8g3YuBkNoR4upibvBh4pEyzYza8AVMzdCCGzkJgS
4E+ICq5BePAB38T/tLo8DsE+QxSfDrpKcx6dnoVZWEfUDiGQY7ZFw+jIHniaoUNrktLCNwvVXXOL
nJ2F018Mm6IY847EjlA6F7jtIRAmHV/EgW0kkDG9W9rNNeSNDZJTfiJ52UYDj22iyHQ/RteVpKDk
U9t3C7xWj7aaBfNn3Nj4ffOU7TnTvDRd/mHRh25x/HjitOeE1SG93PaYSlkUgXMEmbsNWZlTRYCq
Rrn3z+dWBZZZgKBiSpdT5n4iQ2BtWmTX1cYxZEvq153TjiaNw5GC1chzKdH3D748S4aFeoKYzyeD
k1nfRm+sGMPpG0H73ZIXtCYTBP+lxi3SA43v7IZ0ZbmFOpMTiqyWYfk41ll1ELFlk0uWiqEy+vON
GT3oS9Swr+Af1W8Oe/oq0nav78aaEcWrMwDeAf0vMQiWwpdV19Sd5R7Be8RkGL/dJ7aMrJlm6EIl
hGhxEoh9Jx2EbFMpO7ARVV3boDKRucOzUUYdcL+FvJ7QgR5mD9dt0OkjUb7AoU2yXvMArZWECjFv
kMUu4JWUmm9iqCr2k4c9cjaneDfnsBEmy8DHSmFfgHA23gL4P8LODiXCAexTiwr1EzW0i1ygmIlL
tYPUoJ4p++1q7KOgzLQvvqf1MZAE6lvTG7DLn1iHiaNJ4LZE07vDMf3zLA02DnFLjC6j8L3ssGIP
84q1PhYU8Lw4Btny5Y0mNqNtv9cMFkKYxW3u/WiFvqGJhNX1YHirBXdVFuNHNr4dtMsjePVSmoHk
bKghEWHXnWchn5AfJLtkozYLZQ+Lk/htqr5ipLlnPlIxJvMb2puT83rgON+eqBJUcBn1qWSdBZS5
f4GRPljLwnDyNpvJ2OIYB6mJ9VwDF+8rmF/87cBxbPWSc0r0FPP9gQ4+S0ACP7ZbWhL5JqeUBUpa
7NdiXjKPrYZ50uAF1+C80wiZ8eYc+Unc4L6O57HnAheocyssPfDt0DwCQWxolMMyjtZ5lEpDh0aE
/sZHQC7Y3plVUh1ephwBFLhyxx6ILIaSSfzhFFkJnU4YCPKi2CNnyxLU4/Ye6BWvxP+Fot+nQJTL
+SZd99v0tHabQCW+nHQjjMqDnktGXx46Mp2J+9saT8a+X6eNjJH+K/VdSY3UTXlhDaLh0hMQzNru
vHmH02QoDEifJ29hSZ9fqHF6bKFMK6uumLJPaVPYCbmDWd7+c5WOpXQubmgm5gbpPkVhbw/M9x1M
BMUnn73kh7JS5CfPvInFq8RUsAeP2IvQD6YHumUQtkpb25YqVMkdCqhHHn2fwl7FP6UUhOWp8FXI
Ep4o0cw+ir8plGA0ELEhOdk2uzA6vrt3mIOoi7AuDs6EFrhIc90TPg2Sih2ccwJdaP3v6AFlu6t8
vDrlJTzG5o8xHNI/nD0tLI139ORuqBR3dwW5s2mneDfuaeQf0MIzjEyhZm8oqDvkITE5aF3aMZjg
iNEGHA1fWH39Ez5L35Ek6r/mBCsk0eMbofDe7HtVVvuXA0PDD5u3eKqmsr0gt+o/IMs1kLucE4pw
iJ+RHaBU1UJLy8kgIWwK0fVjMFydsDH3k+3GeRftGP6ywOHPngaLkARcJO2Y5hkQQnZx4hs6uz++
RICmn8oFvmp9yhHKoDM7+JkW6+Jihj0YbL7IHWVzj0Dh55a8e1kkH4qysKF/r+/uIxgRCWcDj9ul
EfYMfyiFOgvCbHQZJHhxR36AK7iQa6PlFpro9lLTSeMOiBSEGPCdI2jVOnLKteYkJHmLv0iwJ6oR
9zYGiWO+MnQB/Kx13QdgiaG2z/a15UY51pmxX4VI2mjwI1gT9K6vTadvcyfeibZhJTdgLiQoUA6y
K04q1nYsHWIcFHFh8dxxGDEfX8SyIFzxD71yvLldSxDIiWsSiLrPwUqlhUG8wC8mY6uIhlZgihNj
OdtOZJe8ngtT7tHVnBwRbIwf6k8RVo+pY85ldAjgZ80TUl+IDU8k9b2JGbf4T99l84gXlRZTHR+o
9XV1sw2gxeyeyZBxOTB9ikeL8fimz0BoFDlrCsQ0Rx8yjlatdlMD/E7kvHn9OowvC/AqnzPQqcp4
D+p0Ddo7m1171T2ySp0U15DNlmemAT0wwDDZgJFAPEK75KHWJtazky53HWvlcFiI7PoS0Q+8ZdWU
Tc6WvASidMwlHS091t6QMeqHOyp1k+fOm7nWSjglXSxIb3RBe9Ov2vUZzouI8bD9nhug+eKSfiMU
cjNe4OcbWGr88B2PrJqFWeX8on5aZ++mXvpIZYvU9ZgVlHD4fY81H+dD04G6OfRhvOEWugjWy9d0
hyFMgV8mF1KjZKw8m3aSsZI+K0U3QsqakaEJ4DcizON+XcLj0tMOS9Sc47Bc74nQtVr3pAApjf6T
zi0EtAOORLid+PfqYj8pfLheeVRDDNVRSQnsi2mroe1XHzJClFF6g5oqes+rAz+SPli9i8QjANIj
wLqhMd04CPO/Jea42SVC4rca4exoUBHLOb1iXKVK6yRXzeK2pWABl0yTsM6aVravXgz7je3byaAN
/YEPqy5PwJGNeTYy5WJXyE5FhAcj0YZMf/Szxx/AwD5REwyNjqXtXb+FqOjYI5wI3AjXxuTB1SU/
LTf3uQdCo+rIvqG34TMQZ1apMz/JvMUcKZo2Zd2kgfqoPlUOKxnzl9FZoiADunrMyC75Wow1SvNH
7ZDm7o+hI4gZdprhDxcYsnmJR5GmtnwXXOKfmyqJfjxwENSYHAzc6MUORk6h+yn2GifQmpOaK9VV
EsE738ejnGRew7eFpVOTSm2nrPiTUvywo63HMSzMbjgiYJLFuEaX9GwUiPqkE283eX8GZ/pcoSMK
QeOfJrlAx/oYBNm+Dl/eK41GHM6EucIJZ78YYpnNALf1eHjxIFHVprzrnOVRsmk9toP0ZALMxEtK
KvaZ0eQZ05+kUXL+RXvqkpin/Iapt6DQ4TvudbDJ34nzk/nUyDsEu5nd9411qVRvhWskzuVbOI1r
L+4nTL5FnCYDjCRP+SFVu63espVQ0sLXspq3smratBpIYP0BoEW3uuRcCPLa8frlAISh3VvIWkdQ
zJWrMDNV9EpXczt+5XZCgvMkoJVHCwyMp/Oxvi0cuVhZRqrA2AHanyrRf0j+yJJHJXdpi5Vwxo3q
5wXqWNS1dZqqB83m/DT4TmGEZ2k1gUlHCW6Y7nmlTyrw+a7mNT/WVU0I4urQA0qF5vNTY4xC0KJC
Wj6xps20ITixeQzIOQuSoSwF/mFH4docCIZEowefLMAASZD6kIgnOjEjzuJwHC7MTm9VLbPXiXoP
hqRSQMek5kIhvQcau2SWovd8bz7qvrHEYFLNLbPG6i0Wtow0a1/qbWhtNgnIX6Zr7mI/NXTvthJY
Kbxmabo3yIB9Q85X2Bgy+TGhnThHELkYVXS2ORdvPAzWl7nnGCzKujoSS7G5K4BwN26E9rM6lwtb
TDgwcVhhWyR8nSXreRMZnOqlgRV/m8m2iuBDHCAMCahAiroh41UnwzAjcFtylASBhUffhWDNW/Ka
tTaEoe4HEYGwfoXq8GOO/2ONAugtiZrH2r+SaThoHqHVn33DtX5W4SKz5nuawdQuADskeyB3pc4X
3oRiS9NgH0xPTNgbwqrwFsWq0xh/9HlwFBQ1LqHPN+doydA8TuNcgsvG8g7WrgA0lw9rMi823ApE
IQl6gYFRmB+yY85sFf3gw2X5jIvGju+ynOBbpEPv5V37F0+L/aPQ+OKrkskwkamUKB5EkGG0k2oI
d3PIKIQBN+aGNQ04DUCA3rFotNm1un0NPzmJwpYi3qA1znKlQhTLcR164b15/eWFv3wmtxAZwtzG
hbji8DPNq5jW1bmc9DqE5Y4ePa57rs3rwWEK1MjkhRISCo6STMbOyos7xjBuM2P5IhctzhkhjXOz
Zp+SGKSUUBzUBd22vR2AJgSq0BkFpNO1hsHLB7L981QxEu7omNft4URQoxRmj87zq2z1/x9OqAZB
nh3eV2lLC6LzAPw2+VFeAIjqYaBn0BRh/K34lzGzOqr7G2ers0irmF9Yho/wd6w2NuCDC/EJeX9P
0s6Pn8q/axtlUd5dqEBLxVzm9FNl3AK/jZDKU98zgbxYMYLXzLp/pOC7ejmR8Q+3GAkGnBcsdyIg
YleRvMlThnTgKVt4NhZOdB4uotk4ewTrU4u9nMx2z5Uafeo5FWPSlymrngx5s9jvBGjj3ehsRBlS
LfII2sSn1zH2/DUhKYbSdVkKC2XPdGuyNHnJifYMM8xa7KoCIlg4cF26BI3R2hML5zVtAilXBhlK
GIEkT6l2rFch1/XGdFst0dSPqEfi5dj76/cpNG25fGfTEauewdAJl0qJLRCK20DzaH2J4zDw1DJx
+RlMu6Fqg1nyH+TlRXwfc+6Q+UTxbxFedMKg5GDFCry65Byxx+rUZ43+4jWg0leWNrtrEm6cHYKU
cpXfcSMZ89tUotxSNpmtXQYpYci2JGNmRCiy6SJaCvFO0oXPckr2MEwh3BVnozEzsAotfUx9dIVi
oaRN9cjS1gV6znFxOWsMqZ2JMFI4o7r1YJTJem1qFgB7WFU30n6lzt4D1cur3eiDDcbxYr9LEshQ
fYkPN+WBb59s7M+q+02oC3/3DHKuwWsbI/ZsBcwEOo4hFAnPikZYwsLNtsNXq9SWoYGJD/BSVsVn
MvkhXWGkbhNk4Eh1ghMRCRCd8rsiXvXVAsLpFifujPM3+swTLhka2dlYoeLAEqutGMq/jZr3l6dG
TuKiYUC5VyKlIki7evyMT7vUrPiviPwpjxfOm3DEBUt1q3n6p/haxfWfaUJdVd/ecrct8yIBFy0Q
oxp7LUG7gvGBbZ8Juett1L00ij9L/AIGdT/I2/vfxs7mOUGMJzrsHHKXORLq/Idq3b3fA5DWwin+
+GP+EwXomU8xkI7cwHr9ZrQRlNWxKHZ6KdGBhBe0It81NYNr9OakdZEB8jm1+5DKiwcVn5pl7UQp
j3DF9UEHqvAh8+vofz1PkoXSskE2b6OGD0h2qKDSp15NYtq0EOeaoSJLH56s2lbF37tOX9QC3lTd
GucDGSurMN6LklD28uOG5lbhm9rF67MDrGjI5sG97XOgiA5llzHRnfWIlZzwb6/iDx/DRDtmA5/T
zp35mm5qS0R9FTQgm2yWKizbtwxPA/rY71KxvK2WpvhBKT69Sx7RrJwaEqc8WpsTsVdmYiYrL4Hu
pfbdVcRo8MMXAyx18dvjy2Q3bK/m7UEIkzCULhQJtosOGHjl1etc1xi73CcIKIv+4ji7MpJRZ73j
zFB5eFlQI+fzB1uVQ/MKH/B7O5NqPtLpjtrv6SN9/deZNzOR1QpvfYaDoBzx3WGDpdm8DTRMxQ9P
XNCjS4CEdt3BEtYS6pzNbGyrbnvdUiQBq8fss3lFxdBqOU+i4Z6QE3uDEC51ztvCXVGnaYJ2kDyw
186X4gUH3jAG36svwwGeOBefiC87HmeHjr5ynmahM2iehWG6nilP/qrKpV+C07tWSoMKP5ZlM+P+
JcHkSznK8xdcSp29UkxX7+SOWNXwTmnkouBoI6o1LlVeaCnBGU1gZpwNV+YRvwUZIq2G9/VrISKY
UVqFYKknA8V285JQH7s3vh1Eihhv9oBp2EtY+PtnHTJfbVI1bmsRXLC9vCdVcAmoDcW0D3JOOy2O
4zUw4hXkFmYUNPWN6ywt5ZpFTtEP4/v9AqJyPfBUsbAOe8XfYpSD9qWwBH775it/+glqLCQN7HDU
cPHNvTf7EejCDcHouKPXgMjD+s+AUODnsnE+zcYcB/MdLTYKNUGaSJuljRERGUblCOcOpm+I758k
TJBk6MmbTiBN0jU3FZ57vwyPtBz4zRjBjPtoDJnCFt2auqSEkv86+fiHhL+kEy2yhcOTH5cGcLy4
FxrsWRAaiGq4BLtvJU6MQF1CxhpBCo/yogD4BvV/qYme1MVZ0iFmJ/MXnn9ulcgcbv9vI+SX2bBr
tx8PnYkrN29Iq/SWHBNLihW5Hqeq/QxhsO7uipSxNVK0yREdCDfaZZADFj/ODwZ9MyLt7/IY+n3z
buPl1e5UWkOGcpwvO/C/Dt8H+ZV2Ds2H8TInd+6ppdIXYsJvWj0UKSPLVNdrmwVlDmxyuNE8ORkS
AjuxS39Um+ZBxCMAmGsE0gP+DzajDcYEv3fIQIRxkkAIKSHiDKAI6nkfSe7MfkCWi19Otu+jG8BH
hG1cHCw62n470abRbWXS2JhDWfGoOGkQiJgw/iLvDfjK/se1rXY6ZgL8PhN/roP9Ek7z1+0i58W8
i+OspDWd/r1YO9Ftktk6l4Fl8o7jBfQPPRXMTqlsTfKXdLwiTTRlCWryajOEMUfgPJQiWymWfEk0
aepUQd7PgWME14XbQn11wuEW8RTZP2oyLy6JVLqNJISAVOZym1CRau7sQd5Td6ypY8DXl8Oop534
jKvKr+BunVx6Kvo+Sbu/DY68boWNFP77ulRL6GM7UinfUxGG65iB5dIn/gJkmx0YWVnAqKUibDEL
fBXjh4N4zAGL2ElbxINcL34OwoEUpDqDdwtNjsP0btZm+KoGaJdZbDT4J/INmBCfmSZEU8L8dOXz
+wE0mQp7zCrsEufGB5o1Xzxk1MJNTAhdIBioG2S0PyaXbXWDXRfhzliQHvs2DCh2asCzt24eolXh
sBGykQH9HL3njtaUb7D49ay5SnwES9yAgkKsn3Q7TksL8aDtJsIjhwBxSihT+NAA6iRrcQ8vdYp/
kiRBaBFSEqFt48TV6xKjB9NhmYh0//4FcMLswU94WcsuTUduRBqVUKhOFMfT7E3LAeubrIVcSEiz
PI0OQnLb1tu7z0o11EYq02hmK6cnz4I24g43WCS+9aCT258ZVe51q+pWoPWqnJwbah7L0dZ/R/ee
nynjX7nadx3p1NiYf2uI1ijQ1SLrFYTnh2/EaK9KrgAS9oBq8wmrOzJ85sRLm3nlgdQ5NhIH3xXc
mFpiWLy40dZ5FPD75ry0cwuh804V7A6d1iydtC6yzueRtz8lUtvupU9zrfRgwBKl3vH9rtFSvf2T
0AfCFjeMoNEtWA34sRgeWiz8Ciqj+hQ6QTTC9hQ215b2T1xz5A19XfTwayfJNCSv9yBcM+mDlixG
VpgcSC4CJzmCQr/AbXcduE0D3/siWrnnAljsZ9FDvixgFsdbPdxI73Bf6zlbwQ3qjFmqGSgw4Kni
/XbhOXzujF9Nzo4zJbPJMttMPJ945bQSjR3v8NXsZkFl5BJGkCmh9H1Gdof3YECB2DBnz12djzkR
9neFCyChbqTw5pvxYI9m7Y0yIHnB55eg+dty9ukIpbzICS8XIOYq47R+tmLhvg6EgsLyDZt38qxs
F7bLWf/K+9wMY/J+XetV8lfZ60mckXqg0bf0Tg4X1zxvRZA77oU37JRpvIlplRJJrDNaZ6fry6Ck
o+jvTns5lJLFmPShUp8st+G0G3BpaYRiD2L3bkmKAkoS1X8quAvKz2bYceV8iTk7f5vuLGa0FSsJ
h3KiWFPgsJ2N/iAVKTMG0URkK/Q2QMPY0Geg2W58hxOYgR8CM80GBbtNRTrI+IL2tJ+eoQZ4bwXq
j8vAm+/XSED+0g7deW7gaBg1cEACfgSMzoHDrpZg4hIaTZlokJtSycW8TzIkywgHM7ffqQJKcvBE
hZqX1JD4eNYKNf1SZKaeFFjM8l9d9jZrx9+Je2lYM+QslCOMOpY6tSMj546jGBVX5wA1Gb+PeK5H
vwKwPnS60ivmWCjRsivpBjRdw7pblZeYJvL5lQ42Hvi8cbQYEDIReSENpdUVxh4c+QUxohgYwh7O
4h6GCgu6zwr7U+z8woQ8Dk1+7tazwu2d3TdezsnXM8FHeKr/2gMlCT3AwcSe25iHn7lJ2FxVAHD5
GjAA7psZ36kr8qCOjNKPbdoSztduFYodXeZ4HQOFqiNZkTCIlLDmMl5ROQKTc4GJQQbXLD+5my1j
U9aQ43PYWh5UcT+LWz0JY20msHejpQJEnNvObvIettTPoznMEp6Rrpjyu6K2W28+0TypQUg3udH3
frPuBNQDpeyEmXu3CFDqqOoAshf8MLrQmpt3W1lHRU0Fn8bAe+/pmVvA7g+uCILxEyhY0zeY66YP
qnxx/ATStwEMh/5kQ1UIZjCFgh7t80WnxlzydZ1+VpVxi73PzsiTpsp7WfBQqamWw2bowZbOGObw
Ys5w0xE88oViPbK7K5Px4hdj41RxHl3HeskgC9gvrCsztcIdPJaCX1Uw+qtjjorNlNTuaqmu5Vqk
UlLKmJ3jafwJX60YAQ4r3jrF25Qg+pXeLpAdiS8djd3cCpXT8XMvcjVUm3EZ/kxcouTR5eyJD+aV
XBnoYgzk7G4WpHCNdxVkvPdY8hzKtdCPKVTv5JrO/KIt2Tu3YStCSWR09mvuLlbWj+YktAVNTf8u
qrIFjY8o8AfwaF0FgRAT5/4Ynh0wXNFTqucNi73y5PzYvXKUgVQ/GpnQRhkXrnI7kKPeECDY8GNw
r5CGxGvdeLEQsr/3TpWPnCCZztjfkhXSbRdnobsA07tDawu8+Cm0gDD16iaxvKcQbpv37Yp4ed0Q
TmRspVs0cayKGhjzyHNG/aiKJetakZZtYAlGxP21ZmhQfsKsBlp2RFERt6gChjVD1HCbGahOdt8g
Tky7X3IvpSNbqrDUHP0isgz8YSNFfYmBdYmKYQMosnrAaYjn+uygnL6XwYqUPDfV3rRahW9tmdmf
DAD1GrZAxiggNkrSPMNZYAMxl6It8zj8tonBzoVBvWmt/hkortCB1ctR2e63KgmOGiFLe5xKtx2S
AN4YmfovkORBUTETYmPRaF8T/P7ws8YW0Ufr52N8B6LSPiNp6Vj/I/I9+GxBYniVBjzdUH3ZMsaL
IMdd3Fzvcma1W9p2EEwm8tH8aLW+7KfDTUjKg9G8JidYTH/ABS9AFDVfTm4ZMWmqKFxEwBHIK8tu
pzuGIXqhELLFTQ5vTkktFzhhJjMYDIuiyK8PUa3Ap7T4fCT4iLuSGMVu0z57M2tiO1tryzOD/JaL
1ImTOmEXTZG9EHbsLA0axx0Qb1F1Zz3gFgPzQ/fiHRJ49RTl+6tEugsOINfD/BF8LMryvYD5ryAJ
t9rH2yjAaFPBr1Vf3Q5hBhSjme6SsPL6pYSjLCdAf+Qpyra/SRjG6fAL5fW6FU7EUKwghpjvPVp8
7iwJkuHbOS0aq5rDL4ZzuJXRv556+wLbkxOB8Xz3TL3E8j1nzx+56dYsyAxXC+k8KjSYsQ1+vmUa
3qlUI/uwrRNgolZsKK+ptwmskb4/SToKXWxkrha/IWIKxC3IOXAIuxIysdnhGdaJIP/p1h/PGZ1D
7mZ/9HsQOwjNOlJwIRJPNBiNtNudAw84RsyrG32BZn3aOuA1JucHpaq+Xk6Mue1eQn5emsH6FsVH
SrBJBsuIKayYPSEXJEpaKFKcnSL8Bw9HWjnvXxciZjP9Bdim/JfINeaHJEz2A+RF+ekR8IhWA/NO
ifZtY3GdFGh8NR2uWb7BpD8KQ3BJdqh6CHRTWHD9uO8FSV+tV0D3IWb2+oqYwf20OFHKks4tJg1R
w58cKeZ0NCwsurZbYbB0iYXQNGU/xZYh/xlwoQnxATujBHYO5VIZnt6Wc+IiCQa9RXtVz///1NrZ
QdX5okmZkUn1fB6iSCMWG/e8TBtSc73WgVkrlrM2cU2bYv2o5L1s4Wej+N+RWAQqGZb9xH0AU6SQ
M61OnbgOtnycmeZxJe0+ny2f62n0OmlrfZo8l1n3zLtQIFkE9XJFk+iCHGsNd6QGwLKSyGlovXP2
fhDaMXc+3XBDRixA3UUTrlOHkbtPu64S3J50JmDVo8tsPmikqk6HbtvCM7Ca6B/yxZxXXloYtJkh
HIBC8vbGX1ABSLSwHK7Nz/7AfEzfTupGoRA0NbQysjQ4IeTkeNgjtYzRERoXC3oeTZMRQO7ckp+n
K4rsD+6ViV8Z95IISLjIthPTova6Xybg5RkAToUDG7OD//0SjOcUStoY2kV3aCHOSLaVtLelf/fX
ZP4PwmBoBpKmmpxH9TRy0D+FwiswQ3IiTccbQosOHFd6XO5/OYR8Es2vGmhEi0j6v2gFV5tykmk0
RFJm8qzD4ItTJ1dD8WkqwQlMCgD41tFukN8fN/UFUuCrKtK1OQEjhQB//tT8lrgf/8ZZ3RPn6mBY
dMueO4TJ80ejT299npV2gZyVIy52AO9fYb0gRLBOs+GcTlsGerRaQ4EWDOAHNPpTlElHoKx8JXcM
OFo4AQd8MqMd4UN+NQlAFLq9bmG6MQHjtGItzvGAdX6fnb0Q6US+bOldrS5pqeuvcD/ZpqDdRbzn
V4ICx5v95gn4Jp4B+7gwyCNNZZkLOv7aJTCv0fmkiS3zHcoxOtit8pV+wekTUGCW5HabCKZnMuSy
7ZNsbKo6HnNJrtVDb3ZTgfHURcXU1pn7fj263pxtJZd/ino6ugaDidxZrGDyTnqgYsZncNTzSC67
h3SmbxErQStrV8xQWMQ+9/LvUJSfKEh8UGybEfNgNqP6eXLQtZ7TS3mwHZVMVWSXtWElH71OnS5r
9/lqNmKJmmiFpw21WIKduQMHtKbH80+YOQyPfBqnXyMdVvEMMyOWY+jakVgFISW1hna3/poFfGb2
4j1NYIsyBVSJkZXU9kqh352JAwa+OqLZJDtXASYpz9cCF/C/+iXHCPNoz1SIhve1SrpUlVLYy9P3
NjEGYGhur1dLL9B43yl2a8t3toeJ9djH2zHtoyjsscWC9gWCbKa6nz0ZRCyChz3KV5UCUv5sO4yh
CmEhPZYIDG9BfOjOXe4ATqEw96GQ2jUtuVRswEULgdThewhHhn/yKYG3RqrXGOqZsGSsHuPoPR8F
6FoWHAxUoHBmPAm+F89wocawKtIyHXDud40kvZ3QwPdYn+nDaopJ+PIho36nj/qULdB3PswCCerS
W9vKZY+bm2nw0yJ3c0o5NLoSOuy2ccKvAw/qK39lz/jcdXzfWggb1sQYDR0FNQWw3USSwzfyzRNm
5OsK1K/7elaac9Gdkef/70kTRYxEemHIIjxBmCrnoARfZW5YFdCbQwoTjXpaweDUU3IOLryl4rr3
Hrlz7o7WUXJJLJ77FYRu0xQze0qoAwyFnVQDadPHt2oy9TaJLznFdx12esTu6GAh1DOLWQGissMc
rykUAgreCZ7RRMpjvwaYDXSD0S5BVPiVUTcWyHdUsskx8vcqOajL5NMOUEgoGAAMV5MTgUoD5CuB
xiRBOap1zdgoQ81/onKHLIAfMXPP/o2UiGqE2ZAlKY9VlTrqX8E6Fqwd2YPp3XX0uUg5B0t+lTgk
NoxJiNddnj7cyowDegsZuHlBxsVx7Dzo+a8o5rsJuvvFyhN5VHVbnkGehrp8ZjK1A6Ji7xKxNxMB
6ghJOj23goo8EUxc9YbXq3Sx7Ve8CAdZ1rb+JgzpvBv/pB+gMk0DAEfWTD4BnodvmTvoI5JZXMB7
wDVVQhURSEFB3Zcu4LgaZAEn8W3lX9HsNNv69J4lJx210/cT+EP9aMN07rNW20fi/QA+XyIhV7Vo
KN1Dfn0dM+LOLq+lqS4Gj4oALwyNycnqKwPip60gOEoZPrGKflSC7Kdl/4Q8jLSvGxPV6/8xzHlZ
4pLKLrxcW+jf389HZQKOltym3gF5pYbQPGj/4BhnwxMJOlUCdAMMK2RTDB6i164kjmrfLK4ciXvj
lrFHQ/98RB6cfO3N2muEePtdbZ/Kn8c3iX0UvHzO/xFmazXAIjZqCptMw0Z5HLPUKuYAF/jd/trs
h1/AWejboKP8DaxjKjHOcPm9JcgNQvW5POObbWqvh0br04+zQEzPUN7HiZlfPXw9BCen45WWP+PZ
AQzYLI+Bhn2PUTaO5e1CnoUaITkAszOC0x3iiccwmooUJnELQfEGfp7foF0o2HcugLjM5KtA196M
4/g5M64zRsRZVzx+d9bBBuFUvFz9Q+dUnlaDgelSGK7YtSyW6UyCUNeFNYyPkq050b7AfMXPfjG6
Vkrd2X5k5ps1G3h8tCquKmcd0AL4A4hEcZZxEYwVlr0LIUVSeTfvooX90ZVKtNGvPYEw3rt3Wgxb
Nv+XGXkYxOYDmLzK4TCgKd0gTUz2g05jxrHbflhnyceWToFx9WkJrFc/vDmH9aZFGaG6c86qhqTr
c6wxZpb36Z35rTcOwstK9+KHO5iw3ots/047gGJNLLIxDHmULXzRgWTInqQyno3DFlIq3A80eWa7
uYxZuOLmwAGprzyJ7SJKG4OeSl9SEMMjb6R6wU+3bRvn37y8zqKCMk5jq95NLG+xDuBSYSXKlc2N
r0PQv4bAMmfDXRbxepUgGW5E1udemyy6XI5rkOUFu0H1KP5jyG/EqJorTe49Dg1VujqmoeOl93Nm
kdaniFjvpyZps/fm4qn19XfT0MYhpF2QWbranWcyXKX1sX/ilRwuzfgvDy421bnwIVftOJAz6MFb
2GOMM6aQpg8HcJJrP5BBXnvaI8zaHy4qrhX9Mo5anZztxT0zGZ8n/cn2lhg9AeHo9nopLny9bLg5
2q1fb4yzZF66EPop9U/hNG2/D1Rvo2WWj0lEzPlbjlH36IXSmihkMn3fOooNcOMgiXfSg1thlFbH
glXeh6ZUNVAS+TrVEpF15pEmtAlMC7MR5TjA2og+AFgfSEyLhs8NLJGNNIM8HbO6h/iyKlLnnk7b
gYBFYUmYzI/F9pJtQPC/MMWCAYVpXBJ++1qgAywH7BlSoz/0/Ok0m65H5JYX921DG+ELrQzwmzci
FotP8GkAccot1gP8A1ROSRI3mIIN3fLBtbZHeA0WzC5hzeky8yA6eeCT+ifLiUakbPeiOo5pZl2J
GKDyvLuEr3CXDaea0faOye/mAZeuTsXCemlok0tPR7C1Mzne2ZwPbfnxqs08PpIJFftZWuznk5xy
fLlLzK59oxiU/MA6uYTByydn6kMbfFOhCYDLy3nxNPEisCMaETH4h2WwG1+PduxXfoVWHBg2frKE
ZYIYA9h+O8+XWTZ+LjOQ8VrQfR6/m/nfbSSvh0PtCv5SmhNk0Ujrh/EMv8+lurWBRg0ePfKTGAyj
/YMqLSGCwWJCDCy4oy0nl8VXtrXyKvDRgwjwU2L+FFSrAtZFXoOV7gpdsUuvCzy2vB7WwT9Sj0wu
8kCUrqyAoB1bghE9Qs5bQwToTbGvGVs2RuaeUmh5DNEzo47mHzqfeRTELjQgtoXxL58C9QBX1fU2
4NzmU8u39lH5dcEylyv1FStNr0mu+s5xIgc6pvd84jT3gpzgcC5n2RLBfaBMOX4Cd97UI+icDROf
2b4T5G/3utBUtw4rQQyTOiu5qDcMRx83F6tl0z9KD1/3BDRDbXqJszTtOauSS9ua8hhhQ+T3vunU
FZ8N/xhLZJECRJsaXZtgedqe3oEM+qkMql3SMlcWDWWI1yCBUDemffeG0fc61VnMGMn+9xdcE6gz
I0jHqc2PBcU5i90ROkr9h9rmURZxG3Vjcsh5l3Rljxutjmqt+Nn1spBnKY5Ik6eRg1feAyYth87T
7j1yC8386fSzcV/VkxjvdoOJBigQYQF4uU02kK9N0we6tO+5//FeSM6VOFUBnYy+ZYyrqk1EEdv4
d6PwTr1nQgM4BqHNl39TGdHfZ5hKch2X3NmO+zA3/ogBSDCetdyuOHQeEDtvn7hZ3Ma375FZ2Svz
X+tG2ESr5/U3nfaFETjnb56PJ6E5vbtJe2iOEisrgEk3dntpbuWsMhdoXoszVmjHBBr/gFUxIMTh
it/7jmLyilC+0crPSuXOOewzU8dsjC5N0KU/Z2TdZiGFUJLpRkuJryijs0SOGI4tQODvbWwdpSqZ
ED7/pftEeLCM6cE+zFhDue8uD8SNUVIxu+clSp9t6HrGEfqUXa7Rj6kurz5DTgU28f0RHFPlPZzo
kMbNCIX62r0/fsqyj0FglWTxZ2UwoY6Hmls576SMz+h7CTJb0Anxe4+qQ97hCrz48ae6wP05Brn5
D8Ezmhl2fa1e+Dl9QLEM0nrzHuks/1KbBqigG5QJ7CJa4DO1zMxJwuvDR4JawV1+hPWQFIhQ3wwa
NIxVTieSZ7WrrEbgzsuVlhC49PPtgfu8Cif/48vMVc2sj/rvWEGZw2i0cZehaBlomfH1NMzL5d7K
rsev/ccnj/+7SWBi3fq20hUBXB19HJHUtZR7jfbR7HE/2Rxti9HEcablT1s82Wk6t0t2l1UGGtz0
sLVQXfxAJge+OaqYEyd9YmKeI7EBrRlonKtNa7pK28vo0sW8WVs+a2dm0/wacqAyy31KOfP705nG
A2FK+k3yGbi102Wi0WbsoygzsJq+PIuu7Ij8yey6WESepFg78GNS3PiDSJotjvccreQx/5+sArku
Y6/hNXac3mE3/AIqOcC4vl3dLivS9TQeSmMkXGex55bA+w5uzd1TM8vCEMB5pLxfnkO02w3utABa
2WTOUPtnph1krA2K3qeSW0kJr0lmqQ5JN1bgi4f55AQExTqqT4HIDabNeFF8zPWZikYrRK1rlk50
gsSWUEuQTPKaanGr6LdfFbPcIVw6aKCF6WbLHh+S9fyp9v8UcryJrtTGQ0rXvqukOZS4V9Clp94t
eI2AUP4bpYXjbhD9jMmAENMAWxbvryr3oyZ8jPkq/GZyEbT6DoMIY0ndCSS4igql75tdLjoTTb/k
JJP0fzmf4AKMOacBDyc3I6qd5q1t3gWHB5HxyWQQ6f0ibpU+PeRkljCfknvPBPqI4LMG3mTbo4fn
xiWSYeJ8KH4oJVea3PR2RGgUI23iBrf3EteBq+kbq0X3z6zbqTN/rmX+jJII5da4pKlupJY2EkQR
jjadZcUPdEPVui0wNLhGcQLBHMVbos28F8PNjipQvW3K6Ykxp2WfNG6ln8BcWdXOBHYLqQX2wJ3j
NCJ/qwHJvaJqsGCfTa+XCSN23X5p7BZt6hwIuv0i7x44y5j/erb3wA9DIDn11Ei9IqLkosvcs/ON
TVaq7c00/SJpU0ZUN41lwdhaGVMc7oQnZuB7+qw0sKuwbZtsBFPQvc8dLUvVQ5l8f/UnRMreX7t+
p0AF90SirTI9mC0JKoq1Ab3Wzoh/DN5y2hIjY7Z5/QGoOGlHOdmlIYIVfAIy0J//Ux7MVtzeYV9r
PoNDyv7ypTVKwhHPv67Nbqw8hdCU84ceLM6g2rJV+ZRFm0ko2Gh8OvlDpk2Z/u7CZw13hiIzXUwJ
/5R56tZzPaM1NFhBVoYtAJZZWYtEt1VkIqiIw08pFdoWBM5hTqMZV0nau7z8oOPOR6uuetdQlsML
3O2j8V2Hg7BQ9wDs4EC3xaETxPxBPBtiYfyRHGiX795JjXXsQZBag2GnrEJGVbBPlTxNGynCnhDO
Ff+tA8MGaqkaF8MgekKEwftaK7DPZhpYq0uM/MCaEtsR4DLGQ8RuXkKzuek7Mx8EY8A9+SOc032R
gXdNyGW5tjPlQH1pdqU1LyIcRoKxwzFk2czISoReru1J+AKoD+DV0pDI6WF1rO8YV2pxfOu5Fi3r
fcyM1brMxbJmI0ti9b6xCkJfgUPEb8MsXylqDOOJVW4CXiVCPr991l3XlVZRYJuMw1kpv9mWOFrF
LIlKZaJr3LBX0fgQGYv41YbnZr246fg2scVgZhu8WLjjYPGheOjU2ANYFLw9iOqZY/QLFY9joRA9
VjGdxEfjsnnWnqrUMCQNFunC+Ic5/iRwAKRO7FcIejtJHllAO4GimfimjXbzxrydANnNjc5DySNO
1n0qXS5Lxqfm751H1H6H1h7/ESR6ln4qebZz8SvwqAfa63gBr8Oz4DEdOiMslVmneNzBY9yFFopA
ItW/pk5MUeDmkaeJuk4cnHLMxoN2paCiDVF5yB6bADb9n3xtb1drtc12KdHhtOlBD1R7mrYDtPfo
m6DA5tEIDNrjGjq7PFK3NnAbna0xgCJz4JP2QIus5oNaE3tQNBmSWn3YlVMpKkVgk4j8rvJlAcmN
clDjyeR9D7+KO6IzheqCVT955iPXDbnPxoXu7GA5BSWVkdlxllv0EQWe2y5BKqr/PvLwbH+dfBB0
mJyrMLeXeMhciDNXU8gM1qyy5QVmoUtz3Ntu/S4gbzFiZb2exSGtvGU1GWVLiOiOBRvkS+3Amgsb
nDTOe1VTG8gXIRMnBh6vZ2Zx9Jw1Wsa0F5Q5nniVSWETx8N3EmZvU9LyqvFgweXszSxjfU3VsGqR
lDnKRzmLL/ESsVo+GMDkH1bmi+deEyUZvXm00oPlnXeJmPzYTxkzoXTt7anpQXiVPCcQbvKZbBqk
3PDG2CwTXL58VEn5SALRFLRq24p7xPJNOqPl0GzMcNhNO5spE0wxqbTlsZzrVaam+hWe8RmaVWCF
UjAnwt/oo8pwQVN7gxKzjHolrH0XdggsSD0Gi954e1wiI4+HB6WuuN/nHPGVhB8dTmrw+HwjEUX9
LO/CEZDJAp1Dnod/q5BplM2vUZqGC+RSZicgpSQ7+vNgrPV0Gh2M06zhH7pYW3o5M6FcMPoID9E+
uT1Q6/EPSXf9CO1OqsoH1WLrHEdECLH7HjTpFJPjCFqjlJ9zuRJZmjCTpXH6bplOZuZgYPZfQ1+c
qzJS9pWH1JfSvnrDbA/YSdoFD3JjeYqcZbTm+7C0eK/vAHYlNvCc+uNJAtnBr8BrK0LQYCCVbCXM
LCHp2w01elkhn5xeEE2wMDHjRXiH9eVSrN+uEH7hOs84rCcVNV/VZsTewDPpvfVSij9daH6CyKU0
t1WODUpHrtqOOzFD23fEA+5HqqyIt5XiSRj4fkBmWTD43LTq9TYIHmY5eZHIWz0ok7KTIaYClTdI
Tu06HSh4OaF2fuaYqv0ysv3SUCjIWO5xa2TOEclUNZxBjQnT2EuUnfSRncAllggrVaSroICdpoTR
OX2GHicqKl4iJwBT6jtXeEqfr39rNLruL0BDG4t7JQz0hkURFbSp5HeZ5mOJg2VfUReMCtiCY3DS
C67bMmX3Gzc6pGSXmlO25C7qVaglB5QuNuFCfBDvccFk5+hlqQbh74juJGIv267H3xpH7jhZkJHk
9dkxLW0WB0V1SSEouGWmsiMHqe+fg5hbMGFN3vzjkQmhOc8RSPncDGn6ntOhJT3CgHeEj6jvgFOG
3fhnqV8J9sHY15UkDEKHjERbPjOABmPFf40X7xNpdjwYUg/KMBhO2yNFDz0pRvmmtfaQ585pRxXm
2Q83XN4Lt8ISrxjrDGrwZk/IRSYKwDOE0IkJa30ygBR5dgSx0KZTOVEmnGdi68k7AktO4d6Dk4Ri
7mFArteU9P5ftPhm+6agVNi8E5nqemRtOOmdpWF/Ki+DyhfcN027X/eadeq2Qd+xlKN57f545+Y1
bcbZ9QuBbxDSRc7G5Wnvq/Tm3uyODMN3ROoOAzQXqwDVASeZdsUZ2MjeiSzRPzfaT6E9tHjSg7Nh
T+53fbnX1L7ZG3DkzxWt0Z5VD/p2IKTcvjT7goNGoyB81JxCQAzHah25oZMbTByPD6Z+z77ZU8g5
QHcCr4ZLhGP3K/vOIhpccG4Xu8ZCqplgMMEW+1tbcFyCMKNGBhAZY9kSRfo9Wm1/OnQh3Y/Oea1h
hypJs4ClL6FqbbTruEnJZ1wVTwSBM8Pc8lW35iuqlfZbKU3WHU9IAdewibhG49AUvPefiARoB3nj
3nxmzFTeKFpK4Kwd1eBZTGgbs1c0PhKqy5j84lCbFffGDkMomTG5yqFWiF/VEWkliuIO6JRLo7u3
huvtXL07OQgtYOpae5f5WtIMMwBO6VlX9gIWQ/9TJdHF5+E9Ziyorn5JFSOY2+VQur+otpEjLkLY
RE+HAT42l1JLz4NhPbYQ+jEcU9c38+Z4PrPz4yJMK3qwpwo9psM4RCaWza/R6Hm8ObC6rQHI+PUp
oTmd+7YB19O6mUvoizCZkHEONASK7TgFPQ9bUI6hmBvyotjco5DnpOZ66kbCo7K8tDuX0Oh6BqCs
Olfmiz7SdN2BYkZ/euvoOFFcmJHGSPZ3fE5feKY9ZVYQK99hPZDHUogO6Z00omjKaqEii8b9SNtq
0wmlfXirIqzAphideH7JbtuZMeB/SYi9sw8eIlNW/qcn8k2zB0/TTrEAxVVcOH3/HCYQf0YQkwx4
4nmKrgvZl0+0OgErJTsmjOCHuzUg5VJcvkIZsNGxyz/MYQ5PNdWGcETMj0PNa7LBeM4SNJD5cYb4
fmWiH113liIx97IjBrMaDKPOsVd1ctZBESkHgeRUS2a+T+hifg4uvombZ/wZD6eo0RPuUMGLu7wv
Hs+S+P3QsTgzexdepxlcz5RD6gxjmHjRffDdq8yJdHlB2wpcmU/FqjTZnVFpxB2OiVXrvqOXmRnM
8gC3KP6YhENX4hPzPlKhMEnKlW5LJXCwQN5w2l52iY6CtDJgZHsrB1L5Zg96ZTPT1783tK5JBNkb
0ZLJJ1U1p1493VsPEVoYq/bywwHe9iQCDxoYhIugxzs7m5sOxz9joKYWwzqrVI5O7Iz9qKnNKqRe
BGatd76WZ+tZ0ZSJSIJ3dxxETS1QASAiYGVQ4Uc/Qns5dOBgK8If3s8N8kl/rAsyYQF3Rt3zgFjs
mcg3ancR1cofgXDejSYVAFDe7f28bqVDavpgtTlrB/t4GUITygRQxWc74i/DhQrjhKUox/vOIR4/
oEsLKaV0y8F0hQ5PBQId5p9iB+mkInQhIt28k6wSnOgtFc5O0jMRxhqioBVX0FYNA+IjQWWYc8HP
wuyHgcOT5pZk3GKxkZ1MuP6wwmBvU+U2sCtnNVNIpmhj/pt+WE2KT8LRODllRXy4dCAaCDOriY9x
Jt6UEUFQazhrdSYKcbRnOBy9Bx1EIgMbx31kiSpOrp6MpGxg6f6uokDOItPGjYBAqcBOQPmoAN/s
ZkQ1M0y8g2sidvjjx5uQR0jjPKNrT26uP+gDIekFTOGFfFZ8KYYkGCpYPCGLzW16TkscFlP835Yq
gCJA7NgkFGmDm9ZEQUIVfm8eNPPfICuMsvTp3lt5tOlZbu+J1l53QG8Jk10lYBLco2ivjWJFiHi+
0LuTLK6DAlh4G9MYfiLDTdoibDXUnL9Hthoniy4SFfAJZD4ePX0qFFOr7TdJj5jywDFfgD9tKQEU
zO6GCkZ3R836v9XZ+I1qVHbJpQF+d25ETIMcMtRKlHL7k2pV/dxoutp55YbSKtipIErp0shf8jx3
SBxFO5XBH/bmcMhJtbNB53xCiM4uO4D4TaJs6E/aRv5nfu5JAZtIZJQUo74n3MVvOZq4NEi0MBID
Ls7K2fma+VUyHu1sx3vZUqWoDWgkAyih9bsYDKVCEvz1CIb6jAZWvJ4E1HOafZzPENZLytSYcol5
A9ffAebQu9+Q1TdVeQbd+LJLHoilqUbsahxHshgsSXz425XZqOmhhByu6ox3SKzcyCXjRockQ1zW
u3TxBrb37xMkC/GqvYGU0BOt8cpf1Q8vD1ORV6FNuvTRf9Pn4i6ou7JaI0NSo3MQ2dm/H5IPQEFI
/suZOrg2QbLt8Tx/vlGBorWo1Y09BoDJ8G0OBaju3r9DLvxDexCW/mInCgmWUiwf6/9WgTC8VUMH
NXsePGnXYkLoHjmUSYNbL9bgQkbpBhVk/YGlP4sdhEGJC9rvGGjF17RVVtR1obtGsXBP0AcZjO4x
gV7lod60oPzppGOZ/qSMOGW1Uv7SsGkkrUq0W9+Ra9Cdnm7Rc5gM1cHvd76tIvxEncZx78RDkxXu
TeODbp8h0IKUtKQEB4YKwHGu4DdcPk7wlTHNM/RWYr+z2GVMcDf8Sm/iFCVtZo/+UyTUekxL4rtt
oVS0KJvpxKbFLz7BecO27iO+id/NK1fMEozIt3ChWA13Ik+wXcRl9KnzirqoDUgZmo72HwQFuiuc
46dBzcXyaKmR539Cbr5da/2q0kzLz0ThQ7rOqEas+O3WcRVZUEAU+LnN/+Ty91nortk2/PtUf2iw
tWM6WyzANqHQo93IxvjHy+7cRwGSrq97atQC0dVIqf2qCSfa+LZdu0fj8WOAqE0Sb8IPmQySYOQg
CvgBXdiCkxTQWK2/onXW9ztqHMTPv1w1mpD30Aojash8/efWp91uoR3Fxq7/RJMBEq2yYSXNEaUo
cCpF6tEbWPd1cjVBTvr0aYgKACy9W2W0En+byERnhT6Eh43kdctZoHdA5UNFDMNmfT3iQkDu9EY8
Vo9urjwbn17wkbkEtdFdjmGyvuo0o21RENKFCnjGviP6g/CCxS+dbditZyOpuRUOhP8pM1UU+VZH
oBp+XHcEgd4MmfiYcR+vsWIq74bA7XveJuC1auwjPdXP18nD0wKZg2d1JjLmI3VvFceNBOPgbxZH
NISLERleJVt0SLslnlEzaISwKyy3CxBG/meMWC/jepZnAHvooaONQ3dmU7FOhATNMvwcfFaiytWU
3UXmQe0ELfLNTW2ZaItsVkjrj0OMyDRB9zZZhRwWIwxIHdd8RQN7AmHwqWVBeP9EcYUjx0LJZ5VO
EpTzqDfNKZKe7KJ6eFgCWHk2l2H5oGTJEfq31S+AKW3wbs0q8zVjPt6u/Tg4A02d1gWdImPSYWg3
ytj+D0a2acSoSH169G2dPOL61/c2Q5bcDkm1E8AlvNhZVsmLUzPqKogOMOSn/9t5Y6xj1HJcigev
rV0fqr2sFrzjI9GZMtKgiufe20o40ioANv2A/7YNF1H6gJPfyTK6GkvsGIglcur9o54J/fs51nTK
04QWlGIwDHtSE48E5iMJD25cFVuHbJ1BnqjOro/O4DKBU5L82l+/2MiPpP2wlSUOoF2FR1e8r/Im
zLei40PUul+yBGYRiIxaHYPQz3pNtfQfcsm3sP1DbDOguDiPSbVvq5yaUI43vQqf6itnCG4faHmH
5JP5rvCNcF76IXW7kTVN0lbqtPGkZV3xdHbCH5DaT4qnbPZs5O1qSQQzu6WhL6rB9oIWnelYs+Qv
PGXuw4sHq3f6rf6kSyaPk51hFjppJQo7XijIDvKaijjRGdxZHtNIxJO6SoD9NsH37kNSVl/hbc4Z
f5c8/txx/799YvA0AgWWLPO3BR+3G87i6QtG7x4KbfOJvuUE7C09dE3G/+Npx9qAwsh/fEOMyAsS
CDdJ7MY3Ojmq4xdTpTrhURddaw3QDVdxLPagzacNue4W65LfWHk3kKSbKat2BFh3J8RNqsO6MbYP
b7zQNui7sV9R55Yn9/4OK8Ii2xrMHUZ7XzHUiSF12Vw2ID2HuLe2moNDB51yMOZjZYXhkrNpsY6M
QsqYxp42v5gfdkniJpQuavUiYSMc1klCEqN/I1OMB/yopGKw6kw00QQlO1gxM78YZlBgA7bA37kb
d7cqrnK4ZlKVLfF0c60rv2Ma5eCrwBt3OOPE5V3XXZC6o/H4WH2RzYaPP4DtSW2NHxgirJZxYROE
Gba7tkWAnARduO/dPwxTUAjyP/Tn4/i1PlpbciEZd5Nj66r3S46E7EihIPWMzBmUkkMDMOA31hJe
eEOo8kwKfnOUT3Cpxgngc33m9aNYuRzbVhOh+62awpQYpkE2qOx8eKD7h1/rqK1NO16yYiahlvga
/QHtF4AmaZ1bQEPBOEVz0Kr+DBvdBQXHwVRhNvDzBSbvKTkg+PRaKzFksSsr9XBcK/t1hoffP9I2
KOK2JNARuhTyVrROFICS4ZGyI23Q7tZ50FbVLAkLVVmGNj0gBn9S4m+loa0oIXVMTRMsJegnFRNz
0a8uMfZIvCEGQFqE0WVRYQmtjKQRzb1IcEy3uAVMkeBXoCAE2mBzIoMxbq0UdktrBCLAKthNc2aH
K0ke2ytrrQ7uN1RtQ3yJplvUI0IG5HIYYynHZq8NsoycVVqOgL+7/2y/DZxNYSMqn8ZiPhozlYvl
riBbACQr3Oihog+LJXxWczXIPNgMj8m4nFemTyipzNkw2Xp+JsUzti+sbFvLji8O/6t0Oz6/FXLm
0Y9mqCtAGph+nGZMRiiY8yUEqMxzDNeNryd/+4idjMNM8O9/+18Rl5RcyalU1RqLs0/aSJFXlGGE
AD1KLC+suQptE35k5F/sGC80RH6ixgvuc5kAWIV0RLvF18R2Ywe9da4xrFIqQgjVbMvv+lOzM3O1
AyvAGAmt9tQhIJvETs5gjlw8auhsvvryqdX3W9GdFeFRd3jDjwepYD9xBaPb+dFn7SNbPGk+saJp
o8i4Q7lIaXJ2VhMMqkVzCQClslusqq+n9PU0OIrW3hbhWy4KfgOcJrvfRT9B1GrbQPy3vdSFM38M
Lc0Np0yMapsckLecCehoe2V1IGYuvTwuDZZLuvDfPeD1Qhs3EFy+FVTj1YKYqVpmg8sGPma0Sipg
KK+MPbTGQ3+YK0vS+kdOQO/5BJeFt9jDSB6E7yU0YoBNMDwfiWXZnrI3E7/D5uJlY1SX8Ntn6jVE
cImIWYR4eoABjtng/m0Uo/0GZR7LvlrSD2mG1EnsBEuP/T9yHLLwcPcjf4nkQ6GRltIEISwHdHSj
Zv6QIBw3kOiyJSGySpobjQiemvty6oJ0rZChanFZdJvKN5ZKk2pgcNlDr0XWJIWnL5L4aKOm5EFR
0//S2DaQChESpyvAGmgBwwmzeg5XrsmOHq8zhSaRuBsee7xcrdgAX5RXBrEIIs+k33FCczh9MZod
xDu/jXciMtbJiZjVZeq0Tju6El/Xus/UQ/UEDlfsMpHQtTz09oWCJ0/1QYcOzgUUDtDh/oMLmPHw
hOBjXYT1u5XQhQGaiNU/xK/b1aSM66jF006Do2VRxR0eyRHuKlAT1kS4S4Gzs1x80hQXZccRJcbb
9ycMz0VahW7CPy1+OFLTCw8YMDvgty/c4/Zlbz8nsBah9JPWNlEFB/B4F4fEDKgbAZQvM7AUj/Hw
X85Lb8/uNdedNVr5mYp4t5/o1tdHSMbXEzGhOf4KtGSEcKMKU2vJDGiYsFqH+x1/kwjKzQ3wPoCs
nui/fluPdxoHWH5FmBUG/QTOEGhnk67I7y1sWfl5VjTQK22wEORvRlvLkyEeXEUZntcYq/+B4ev9
aMBYRSdAIKVhHh3KoC4Aqyu0qeJFpsof3cFWMqgTdBXcpBq2Y198JSoRj2ioknOTfbWZ3M+bzd4/
XRrMzwYUTY5ubcjCIG/SQpj2MJct2j6pCw1cjbZ0ltYrJWByCq65rs3ZQfiunaouzotdFDRud/pQ
CWdSq56sIR708FnYKIT+r3KU425AyL+SXCn/4oi15sPlDG8xYZ7UfpkydRcStwH9QQ3RCbAs/Qfw
Z5tMc3hPZ0LWiky1k/3eicCdzICmsPnyjiJufYehVvxxahHtd/+I15ix+9L6gKwC+MZIi08dHs+i
nYuTgmvw3uoz3dOyCtrbAsc+v1lYg4Qn9qyQ0IhwJvn1Hu/u7+Dypq/IdnRoe0ibsfjsBvT7Qhm6
AXpUyzen1ORvSAmSS6yRnSTgb14SBMqJ+TSeLw+rIDcuNomrr9DbRy9TL/we3/L5p4alg5TnBTkx
9X/oqUUeR+8wmXo67JtlVP0Dt6UFrquuw+8sNEe7M+653Ax3/afTwXYAni35x4SvCeuklHS5QUN7
rUbfJ3Z/FfZ4fDFL1TKMl480BmlQq1+ZKnT8u454eSgMV5BbSjp6mm6O7wN4LQiyDGw6Z/MLfxLn
TymO5BeeKzTUjSg0zV/Pz9U6U4Wk7v6pc3NcVI0dlnNCoQu3nfCAS0CVq4aEl58s552byLv7JGE2
ncFLI4VetHszl29ar3mf9S25D5aptplPBg2E6sixOziaSvlYKjebb/RuI+UKQfembBlHmdAx+HsM
qwwD75p+UpuQ6PdLr4BSSyZJfymWbBNXfvSSTFRdNL7DwjRHno5toNW0gwA5TSAipiRh+ZsuIPxq
6MT0oML051ArAXHVenGGlTbGoP9Rd7bnAJ6eNerVHSOOc4hdU0ngUJ3s0UDeYTQPHbd87dFYai9J
84eqJuOyyyzkicktkSYanxOBxowzr5It1uLqmj9C2FmaV8M8u4+IJMiQBSs2VUyqok1GmUIMXmLw
u+PYTfXRcLbIPkZ1D8Mveyj0qQevD+OFA8WQWqXWkp9dB8G0PKnaufqCncL9VNHNtmFUs8G7FDYr
VzEtrYXDxHERhgEX4FoO2A0YX304vs4ULGe1BzWHxMvHH/CuLuEhdt2jMgE0tBvNIbTXX9Gt6Hh9
xBKV7te7dHb8WJXlitbpBaYAfx6Kc5QwVDYkUuJoa9pSnPO+Mgxc622wETe3pSKqyW+0GrvNhmSG
CCJ6APfUADnREtG5/SBlKaXvBYkJdOg1ztcUyeU9USC2z1BO2FRfxRjMoBkdw4V1CcRrFMu9lxjj
MNUqY5zxUwjP+fVrzJdJBYnyiPhS5Y7XWV3aO83ub57lYY1r1isfvjyWymqaO3A+qHbDOMhLZdNg
1eeVBElIRlM1GsavX9MYRrg89QT19YQhvAUdPcJ4mpve2IWyslRMDH0eoJ7lYKIRKZEEb5gC/5po
ylh1jmT6keyzZn00p3hPO+qW4vizA8uy83WqW2xKb41v2RRe0c1vbX42+Lae+MRhaCy6JolG1hz5
Im1tOQmE8BdGzGg3P2erVzsT+Naux2XXwFaU8pf//gH7l/i73NWdUWV/7MLLZYqQlfnzWRYIm40A
nePiQASSgUYL+7PSNuQ3jio32xkDjK1znsb7Qwhu9oeeT8o9seBj15dXHt3I9XTe7h+050cru66f
l/obqXrqxhwHmUf3AZZ03y31X+CGSTCckJeKOsHfK85KFkoo1k5buJQqbukzFhu0izXi/UK7AzKP
TnZCOq+VdFQZCz+cQAtyqB3BlXC8UOGzoyTwAo7pjr7T95VSH1G+HgWsBBNiYYTLEMrKon91ivHW
ZHfOFsZSlMjeUV+NsI0JfjHG6CBKFJH/l3f59cWnMurkMWvdKV/geT3x5klbygs3kvdEehHz1682
C7j9fpfcubF8yX8zVB/YEFRLplrZzLo4+t4EBJaAMJK93+oWYMmnDJj4CnHhlsa8Ef/lFQ6GRoSu
LGtz3MWRK0JrP95eNVx8uMXR1MpFs/mnFsUJELmXoWsTu4whRRGVTEJq3BhAavt9aJ0KLoMQ6Q47
D+ZqfdHxl2NAmB+qmQdAg5w55tNVLiHl0iB4C5x5+ffClS8lotreEsQi+B/eX/iECB2zrYU2tZW6
v6lj9JyJuQQ/1UYtARXpg2Uo4xNhuOcPjmTW8GY9LqSTD56dj0DhD3/6WzTnpsMUBfZ84rA8KEMk
ZbabkD8G9q2MISe88JCZultAAomXch26P23+MhSjcpklRljOH3bemjFUwoGSEQ1DOcy/56pCUH2D
tBxVuW3BiudUQFYm0+g4axSQG1RuX73hPzLr5vf2/BCLupw+lJflD+qVMXZFx6or6+OXOko6dHwV
aE7aVtNR1gkIvKb0PZLuPl0dUHgNsKVXqwA24zx+EHPeSQLem6y1vfBwfAWFWO7GXqo5lm89h5Qw
RIi5xggyG0U+K1wSQUTkkYnxJwv2dfTDhRszkKJmIAo0At/MFOqWvS0yT63ylQ8v+A4EXsNPGASB
Y8OY371Qjiv6HCKEItbgYbIDh+WwLYyQnGdtM3qLExmUpO+4gYH4hzEOVegq3R9PRWQCnM0YaZqC
MePENga26zcHjwxLWD/auaog31041C2pBK0t3wN7viWgcJJK2Cpi2siLfy1WiIdZu0pso5ypexKo
mNwxsNJXBIVveZhwpc94hAWITojTlVzQu4GI2uz1/A8l9nHcpmsQMpmE4ELNArQdG+zdy4Mob5G6
nWp1uw8/HUgvQl96ABxs6Ibbz6E904xFajNuOwRWSU933uYwu96B2K5sl0pWCTJSAWhmyl1kMC3m
eEKDEcyyQ6is42QUH1Eejl8CscqErrJT+kaZMVN1mnz++nQutX1jWdN2jB8qADbSRyNoR4+O+v6b
CZ6QB4RKj+dRRXpmKx7bW2LZp1y/1WkuWoddOyZx02WpVJgipduTudBNZWdZZ9rG+eERsJC8R2lZ
qkRE4be7qyl2HCGcm/yIQ/ui/RG2usV+Sh9hI/LaFV5chsC6FOc72bOwizzu0O7X2ChF4+jVwEWk
VxXmzBrSNo8kaAiKcx4CPMv2v4Pwgf7YraqDgtaDaPVuwRub25w5UegNCMAL+ZRV5BemrWtGLIX8
pHfRN0RoPtwbcJOSn5Xafi5y4w93BU04Y8nKRXCBGYAgwZeoF6AM/3q86wpKUidPxP7C4NNGLeTK
MvmKJQLUReqU+qemmvzYJZwdOyyon3poyO66lblFmTdGwHkU+99CSNP7JvsDqYLfNj0KarwgsZ/n
zQfmA+ohF/qVc4dtewwgRfxV68Gc+ymCu99o2eO23JCMZGhcle1hBC8epbc50Lgk7pNCyxC/s9gf
1XJ27jA6Y5VtEswGDtMFh4xwLBj8B4Mu4jCkMcVQP85HRRkyx00m5tvxIl3EPtJ9vMHTYyraSdM1
GKXoMT1MVwnYjBGwf97B/+sBMLwqj+Qc7yKNTpSggk1BsjwpPOOJSBEFP25a+0Nz1fHkluR+Ij9D
fYkccg7L+HqsHl8GBqn99A4tSXFvfl3DWMxkxaYceXhatzcsyMQEoutQkj0jnfh6OXR6SYOoj/Xr
8Uy/GiPASWcSpqCzjA1oNnbT2HFXUuPaT3fLpZbbV/d7RC/mcEgFw+YWI1yZmvsoFPHGxd8f0SyV
EZnkiZoAZLmYgJgAukW1O93tTP2SQMePOssjIr7LXx6hZthzx7KIHs6n/IMhcmEr0B4EdAGHdOfa
IAvb7LPMSZMFmYjbI3tl5G3ttJRJDDP3cxCNKv0wQPR1DIXE1UgR9LT1g1RCYpmci71JArNEgEop
CIKIikGx2rtn+U4xavNtlZc6PPtGK9afb+3xUNFukHjJ05FpIzolJNprvJh0ZLTzWICxVKPlzSvu
KKWK06vmkBHG1niujxsmlZwrqXq6p78ni4vgbuYaOaZE6cscl38bNjeCqdtmgkaesBOGpPEko1xP
1v359ao1pOI+5N5u/r0Xk/hNab+9dYihVSDqIdTCF5WmFWR7vk2Vvx/ph80JlbBJqojWU6d5Ac6L
k0YNW0CGSM0XMDIWV4YvVwDRNb3udFi5+EQbQ1LyH83c4/xwjFVKGgMVZB08mXVCE9hjD0i88DLv
qBQ5888fojRzlqVgOBvPD466emlYanojTFyXPRyBogdcyOCTnK+CwZlzsbc6umKjrbX08zjQ9q7O
NU02da9++FPAVKbaRtEtl9+b6+qz9LlWb329Nd71bte7TBiDzHtxVLkkpLy/m5ElOOv81xVjNksn
ZjTNbytMHmfWYQv60kgBmLTGKEYDVO0M40ZrmYC4EyQ3AbfnGIh7W2dQxIZ0TJmLNW8qqn6Xet2P
JBxNyCSZCIfcaw1x4SwUzB3+pT4Rn6vZFm+lkx2quD7YTBXUNLXEsyw1N+O1UtB+gYX4xAzyEioe
FCgUZHLWecSNvVfF/VR02JeFidaQ5rBzBtkFIAx8xuCIAnC+mjAeOqmoAaGLLTzo8bxyrQutBG8w
vumculXSgmPkIQXnylP68IYeWNcGbXkLPIkzA3Muo4gm8BQVWlomC3e1Y2zBGv5MqbtRqrRN2ZdY
b38DWiM1IqtVgRJnWaFWVP09A62o+IdPgiv+ARuNUs8HJxnD2N/bN/ErpOz5RyaEK2+YJkdg5xjR
Trig6YVXEhmm3U9qgnxI7Y2vkI64SPmb4bN8RrSepVfdUR4SB5Ejqi52X7Xmfgf3cvTKJOfHA7hj
M2y7hdlyFRxLZbRaqfQ1ydxYLX3of+doy3oX/KsywCwslgUYmE6gaVwchL7FkzdnJX96kngvuLFc
u0Fv3LQIqT3IDNQB9E5XXkyliN4U84lxwGD+ks1j/zi9JqEvU+80yjj8Nl+Ckqco5JwgG5gm1LuQ
WLJ8JufVjx2FB1AtS8VBoKqeu2NrB+A5ngWLE/su0vtbGyzCSZBjgCulH9eCSRUgrDQJchry58bQ
wwquvF7L5NY138MSGXSMThgkKPmMA3wcyZdscuJafmbujxldC7KLWvbm/A/VyYa8l/L3xGJyDVDX
KBRSt6uwsw+yjgY3/Xkpn16y00B7E1cnHBTv+/hnScW6hoK4rcnrPgVzkB1da25cU6RpOVvSjb+M
8xa4b2A4D6JzfQ0Bmg/NF116jdhbdgEUNuJj+MEvEpdYaUdKr3nf4GiUd0ph2IWMutviI6DOYvYT
cGV5zdLiYnWLRduFgeyLlJGzxy/sumXXaACEUnSuQcH8VkziqFo3Q/VSp6EmcZQz+fiOJO6h39/A
nlbVf7MBXurgrC+qgdutLZciuFrurqhENuONBp6USULXWydlRqCd8vwNNXqK5RGdJlWOSOGmhuXH
8GcOKkXM4eS8wnqifu8pz/Y5UXXe0V5nFRhPKUJ3ROPOXnZT6RfFt4iFWk4hSRqyd/flLXJRJbXs
5h+Hg9s0R5xSpygfY/HjtAz/4R16uqR+2MiJhV09aVoMaJ8IaZWCfFGEJd2cmknVlTGdf538ZutV
moAFdd2uoix5lYEJwqAyXNXNl0L+GEHdUWDbpavKEh/GB+7jhNdnWwk3mri+QB/iPZSjlp402b7O
g5o8u0tptrqnL0L3dDDcWGDt14eKHF2KdwNx9NxlcI/jXnKeRwY1VF64ZyASiupHCZEnQPyaiLfV
s45yW5LB/+e7VLq60ACgA7fN3QGrpEUAHt0NolN9d+Bj0bqu0Tv0csW5q/x8TwQ3d+Zk9W93qdPD
6G8VIY+uF3E3zw5YtbcTbeD5bbv4bIAcRkPruH9Mr9j7zmiPtXy4t5nUiR0wrjAuaZPeLy0FyvQt
SxEV+Vy6Cw8NgT7aMfs8N2H4yMm3hGsKhI5IpajjuVdfomC1wyFLP6nrMIg5ZmKnucSqNhkO+9RD
c55P0P31VKIv0/W/4kx9Ybhgmey1AK6YyV6noNd6sCfxYksRGV2tliM7KI7EzmisU2KygtWwaLHB
LM6udcZbQC94OJdFdgU9ksZ9czDQzF39yIk3P+ZYy36VLTtOn7gNTd0sDsIMahp3cyD5qRQjLurY
jqBbHcgVDQ80s7aaTH+Y3O4zdSBbopXpB5JD6B6Z4Q9Wmbr++9EbAPUSlSeUlVB0rGC/KRsqXWIE
h3RTe6ecOK6KhPtRreSBcJUk6ohGG+IFKkgVzoJICywAnZkAHIyrr9xduKWl4CDcgr3oDBBblCs3
O6yLU9vIKX2j9+bTbXAV6mf6siyQi+Yv/LClHM7A2TNRI+qNeikFbXyXzMeoWYC8v9fT5/IovQuj
CEH1HPsj8vL3C92eONwCvEqbQPR6aQkDFn/nunK94TQH6wK1YFDLa/YJwGghP6O1b4hHRJcFWjqf
PXehu8t2kZuBcpYZ8sJLFPRP0OSwHdrcA4QNOzP2X56R8V1sU+TOndfuk3yJBAF2dpOxb3yCG88q
mVz8Vuj5hAQ6tpcC0aLSLpbDChWSt74JbJEt8e5W8HhrB17iE4hAgoPNPMQ7DcwAVqAvBm/Xc/W7
0SnUZXZGq8CeFXI3d2yVb9yNJio1tvBcopOvAgo6BwkjfFgXxbe6YPv0/B8Ed4gH1HQBhjYKf5q1
gFoo1OwYMu90Uf8SoTS/3RnxuqAyLg+fWvzBnOmA4Gv7DQ2C5xpMmTUlVRsozVekPO0JAMtxQ+yf
8O2jxxBwyQjHxicPx6jW50RcPe66Fe/6X8kI8Y/ADU6CuUWIubtXfs0izaW0YPGGV0w7vN5CED/P
MVglpUPhGB53ubM45EzA7/VzPnlxABvyGKMcbcDwL9tahpYnBSGMVpzI80ZSrOJFInE51Wvt6YnM
oeX/+D7Mv0qZtA6jQNa33icuviA4ZujZ3LoP3HBSM6jgMGBu78ui2AVmI8atsAFYyhsli09qvYvB
ZKyAB4RBqaNkD37ggshdVS3689e9+6L8pvoHGiyYHXzv+lsrD4v6Xrtf3q3tprBHaCJlJSMnFvST
MYnP+WGLvK1C5XQ0kQqtdeDVvgjhqnpUYGsNq+eOAX3ZAp2lVBYbuV3A1J79oLKsYxfDxi59H914
Ing4yQjvJumLDZhpwPvpV1KcWR9itiP+tJf89waTFVfgpdyb8ky98rXodLy6GzlFKwX8cyTokPsn
Vq+B9zxjW1PCd4VPutKlwpoIEtdDrzSVklz0V4o+s9ZWky4t14kkGK5pD1BwY7X4llBeZ7strvO3
NTuTJLlfi0uy/tJaxGYWKpDMKEvOyTy87J9OltZIvxkkxUa6PrigLQ8HusTEkA5sSGtVKgDfPz/C
LL9JIoDVXkObtPavkpGAiMgofciRRYfnNkkwTdVKFlUT4+YBxYZR9j75vv1eryv6q5KUyafwnvO9
L8nHb/E1Ho7QQnVa9LHDsuTftouLHVxQnjdRxGfZt6LFiqTnA/fakOAFlfQrYJMoWb+XxnhUduOp
GLe6rzULZuZOYQDJCYQTqoRiY1WDegUbAusCADWG/p+R3xdEprM3+6SyK0RJ47XMUGug/vY/i6ku
b2Qu6zvALdJGEJqOqzyGcjGP4ylfs70XRCF7Mui7IShn6001uTZKI/ivb00CdmvF3ZdRRoTZuHIe
eE8DtV9dh0H9uten8T6OFJawCVNwJRUxR6IhJimkK63Z7THKgmb4eKvN/vmnJbvjWg91NotF7vG4
2OnKxlHjCakulqeJEiD3a3dzaO41Qa9il9ueV4xRDfhGVOT3LwvRB6vXPy4M0aGO1r80ZfKCPvGA
No0WA4tl2IzthTrjvgJ/RSJDVnTAdlm0cpv+rc6E6OdMVuPCTyKC7CqCgejbE7w1nU5p/qJ+uJlB
BPVf07CdNtv2u5433jV43mH7WBHUce8uhaH6qJnCjQEiZZqlhbs30BiBzhgcxe3vz9U4pePkaq+q
MNZm4gBwZ6e03WJZlk3V3nfaPZQsbgleanX0P9RccwhAdXgWn62GFQF91ZnDEZ/TI04FGzMzgsAE
BKrtjLTaBOxhE+PxVENNpS2k5pn0g+XYzaJpIXK+Z3A8lCfzQ5hsDD5utxo432XAp8NAzpaHthrX
M5vV2xvlYwbScNQPx1eqvJylkOMZU/7P7QQ6Z/rV1kREUaAohZMJuHGvVh9VcsjlcI5nFFM4OWOo
d//S48Rpp5uLZFymzVnfQk+suIV7ajZepvHCB7rtTy10eS570JdFrd7vCjxPCOrw1MAB96+vAzoB
KoGHW1+SO27vNgKfYFVrGPZHhfFpX2mIcpg1WcKGrqz8+D6jLHZ8uS/nbhGIdpeycaLkmsJkVKon
VBnlizuNPA2nWMiw+uO9HUbS8HRIwmaXpCZIhwtewAGxk1r/218s8qUYvdOnF5lGsLmhOOeRkmdY
9LWJkor8A6qwNX8Ck9CygPBE1jzhY2jBhrryP69q4J/WzWDaMzilvvOsJhOCvwFCL/n9A0CJaDm+
tntSktHN/M3hau0vQVbjlvAoZIv1qQ+FP7J6ZKtIwtEiM/NRunngHJxWbr72zpb33mOgyv+gpo6E
5kCyEk8Oru30ERklhvpuwHr9FVVysCJrawKFqvTyH8zK+e32njE+3IbwF3IHPHa6ypKmP/kXPbX3
1gVNFC7p4z829+mOMb5buPA0R1HH3V2+WEbgL65J1BKi1MgU4DIQ824JJNTYgG1pztqGq4RoqwKE
yBTDJa+z1je5wVxyAEcPsot9QF9pwB5BnhTanGnRS1unA2ZfF2NQEeY+IX7b00iOLBGraxCewtvK
Jm88Ixv8midqkiGskuiVS4ucJOTfIYQHnaXvonRLtKyTS3CLDTGG/TfGiBiuvbDsyhKxOt8x2Hx+
df/Cgw6JXb+pjRoh3qAXN7gXg6Hy2eY6MjfrIwU3EAyRe2yGGtebaPFvVGSJE8MyEu+ViZUOmDMz
qu98AvW1X3FajzjyK/FPXe7D+CmaycX0dXGSVzQIuVHejvxgvd7NoQ53edUaIHxi2BkqPqyFANUr
LiAYmpWIotZr9rJlCeFnut1GeQWtv4mdZ8fpIUiQft4Wt1ycH9Xpdt7gmB90w34NsqCVHbIzcgXR
/nvq71rNdmJ88dRg29SHakLhoc5Uv4MAUpV4chTlrfXEM7KCEZMIxhcEA5Xu6Ko8KAUN/ILaTn3Y
hoxBrg11H05fPO4k7Cz+m9QzkV/uV7W4jnNmWmFWZoi5OQKYHxlJXMmKea66q4kVtWwwXWzM8myq
LIvaZoDF1b35JL05IlsxrkCHA3bmCCgSRzmxjJHGV41L6f1qYrvNvJXD0W5jKPD9s2uo+oY36PIi
BWt2QXFWKDNzjSCOP/8qw86B989wjmUu2vTiqpQRxgRYv3uavB6t/xwx4Ex1tZbT0jIXn37TgV2b
E7O7zQDTXf8fogMWx+eK1Fxq0egdd6l5sS6K1VS/fRclkZAvx9s8jB3bGxmOJ9nEBmLrgMxVW2Fj
2B8UT8UP4jX8s7dyea93dCdJ0ZfNCFwqfOYgxgeHtEJu750yk5K8Ydaz9ClNgn19qAbMeiT26RUg
FqyKJS+yusmYImuzeIr0V5GI+QIkn+SYCGvi1iGVVGlkYZUigAePmmIToM13iLhu+R/quEit+ujD
F87feyduca6bUzCJuyVd/0hqCnamKQ0jnDUkDaq76gb2iVtkNWBou2xQjF0utvJbKDUAjNVmCCJQ
2oQUg6tduVBuHZUUoSTmpHiDJdne6Q2Qx/LHLjZTjID/7BuCH122p40yRSs561Zr+RaoAc5IQmhw
SaBTplS1RC8mkHFfUbfAXL5qmBGoYA1Qci/2Uq+PAXsbUAOPLR0HzrkDFotDNhsGGC82wAG5xvZ0
ERp2xtXIp9nxNbrYKwtaM7f/x1K23YdMqK3vXB6FPSzNNjkdhB1OKrmjeAujLq9gpaNBMzJ7+yze
6mPbZuOVaZNvycAxiACH76LIo4MpoDj+6V37zGmXAGLPTjZUfRYJjsatAgASacqI18z9v5AB7Ya1
RACO3LM+4hYSt2wtHIkekSW2xARM9HIVRw5uPKBAsUEeI32BT5KSpkV6c2UZn3uunw7G+GqkY/Jl
aUsk2fmPhZ/mYX3d9yj6OJ6fzkojvWcw9rpRBmYsOnuePJmym19/OYDWoZjrLnJv07xVLpA8KnY4
01Fok97B+JIN0U3UCCwMuz4HVjj+iidMhzsSP426ql2jDSR0tMSu/LzwP2jPyIqDUcQZ5IKTHLnQ
pP383o/6WlIsrktyrV6nFR7F5G3zeyrpbaHhR0BH1rbg0EnK9BQ2KTetWhpJbGYrxtkc3Xej0laO
03JlUpJqUFULr2HqkH3nm+lpVrCzYLSGBwXIwDKK6/I2o5E0XKJQUBBsas21SQtCUp6H+coQQenf
yitEujBs8SHIYWx6C5pbK8Zw0bJ43Un0usfQ23gfCQW7EWX6+M+Nuek4jXajlsCMOTL1XRsTmpuW
ksQuFa+QrItETW1rPSEzCcgnRw6ZATj403rogfOjQCKkuGLHCV8bqBmF6WH3HO9JStwRcH47cbYH
qTXmUm7TtnNht5jX1rxn7wvev5Dh6oU+/lLlduhDwbghIGCk6ExMnRA8R3wlPNsOPIeGxmobEKom
6LaexQqhHX4r/WxyCFSg92rV0/e2OlO7uJ8UiydJmKZJBH8nu1622sHOibjBZA+drfOrLDwWoJwq
o5OeAy7oE7HdVKMDuDfPklOAk52n3QdiUz85xSHL/9paSYWN487vWa2+mj6nhXcfMfyj9dDsNKIW
C9BFCqU5CHLDnFhdxG7eBXHvfJqiLu3XalkoSfngnu/kBjWCKrvoE/qzFT7C3OQzY6rXe7p21bGW
wlS0PUC8Q2GyomX0zKmRI8i1m++cv+6up1yl8ifjU2ly2IuL9eDVr20U4U8QWsxyWLtksSdjPsj5
O2KZqV8pVuAPVruVEiozec95NGSYq++YaaCyDUcWgGCfGts4ZQHqi5O1W3qAljT+FiGUYA9eUWgO
aurhQtTwe6Rr1YrTO49BhngsH6a49FVMKVeX6GoNGURdtftmqNVxK70HDid1OmJwZcWD3+vOzOaI
+IypSWH/j/udISwiyw7R13F5ZTBSL8vkqqbG6Hf1B75cACFE617jfgHsBRL4MFEopogBiTAblPN/
43YBazdVLO6D7u92WP4Jwaq2316Fw2upAiRHY4V+mfp4m9W40CQKYwkhMdENt4iN/985Vu3M41AR
slc3Napx0L3BcrCIDpGWPWsk4kgNhSZMxUdU+NsoGxDFxJS1JStATFOmXL94sZwz/INd9BB3C7h1
gzTVxEPglvg4D/T/+Sw6itOycvp+RjSB4JnyukRKEorYUSMvn3FCT5WAFmxYwt7k8yFUsDDGQ/cc
fCqHnGloLC51fJjs7wEhlEVce+rytJ3YUbAEu9MZAzEkFbDqiGJGjvRLnyaJy9Cor6VI2BT8xfvq
csYrvipG/h205+shhBFftcTDnliKQdos02dAL2ZYQiWw8pcK/P1HIll75i30U9Wr0krp7i/Ze8G9
4eSro/hw3s5bGOZ+wg1NxOEapHS/Agim+KxBagw4/Upm9zd6vUg2H5s8VQmMFAtwnrhXRthmvo2o
tfIwFS9ugA/kd004EnD+sKM2hIc+nXaCiSM2B3p9LvuAde5pRrjdb+DqEt+nS1Yc0gbwgf4KYddb
GL/Rm0yX8JTfWAPJeziIyHrU5Xmq2feisdutdZhKTF9VqQkZbDwS13KzIXBdwOMFmG3Is4GBs9e3
QnvZJtH2e2+f8B6VHn9KAWHhPuiAE6lH38ZfS7BMJvvMzm+5BJP/G3p3aqJvEFqCFSc5Lc64l3UO
Aba//ocni/evGfGsU6ZV0l0emiCqJRkjUNM7d3nMwTWLSZAMaBcNylFCfZqnhGJRnQDAL25cDE2C
sLdAAQk+LvUvbK/uFbkNkEFUHu3A1GkTH2pLaPJIxSgvOL1jg3iZhVXJJoDHh7loSuQuWzZ4w+15
tWBwW2nNTAqfPekC12Xt9Dj9pfciFerCRH5ivpvcDF9lfQ+nlYg9goWLiB4JkKvNtgYvytFvgCXY
AOThQh/mawbpZNhe9ZWMJrxNdP8TpzWalfBnrhFNgStLeUfzLhVvuBhLsudl+4/t53Affvn7Ejvt
Xz3jCLuZn1+TRgJ+F985pyhJXHJn57AVPaxH99CYCKQt7fqCuCDYHcOuRNifFhgWIMNaUxf0pzem
lGhRZc7zPWcPKanzuPuk8DERHyD2EwR8YYlfuAoqLgCBkNGu5KYyujlAdiZCqID3M8avIom4V/06
PweIisQ9vxp14rsSrtuT16PcmwmFWUg8PKSK7A+jCJ+UW7Sad/BkgsPOjeqPy7OADV1tuwRerw0A
A2ELFMcVrleYut7QY1kbsqL1IxXt8sVVp93G2cGfaL6WA4m1Cm4ceBu0m9rsySujoiBsZ/vtM5TQ
VF7beIqGYtzV4y7msUzfTiWTsIIS57XZfxC8ZvYmhIvmmutnm/lhUWIboh2aPKF1KWYdd1iA7gxo
BO8RhwvZkDSIqNjD62H1LyeHMzNtbf46qzd15BLsAh0qU+3Ji12PzYnbsuLA+HfB1ez9ajjh6h3F
tT2DYzDo3qW8S7QJ5XCsZZ4NQCMDnhHGoOpTay5q60lXHACzNaSw+KiAir26sHQVX1X+RunopoB4
j9b1yU/q3UKRkPyGNBD8Ql93t27qkeO28KL276D2vj6zklwTNM7qhZka7kfgpwH2H/NkkLlveKTL
didepayYlaHYYkvaYBqcc+7jKA57FMA2HLVaOkN6XZm91m9t2tyzs+DHE3fZWo2SoAfoB2L6zhAE
BblAcsOX/XOO1L4CgF9/CBiZw/HAU2ruNUMqwShOKKz5CFnHvkhF1uL5Kdfcb3MlSzHkKct8g8sQ
er09ztJoet7Y3AJnRWyB8Rv3oxLnuoU7HMBL+CNrOJAr8DCxhV1nstPlGv8TM6f+eOKMLYURUAq6
trr8rqtPNxGCoO/hj0sZJ3gvF0Zgb+cRXBIL9aAvOaffJJid0Vcl85/e4VsPHC2x/V/XDBfVmk8r
LC0uO15SXljEtxFLCymA4OXl5e7GarwNvqV7EyrvYQOl0E/8tfr7ofX1sfdUmBf+J46laKR6BXXu
9LmhrHUmGYFnoYIfKWVZO8QjcK0jRnXt3TJ866w+L7FsW+6NbedZIgOQHF4s1PhlRd0eL+QMohQ3
8CG6/qCeVDrKLNJuAdAjXSRHl9S5Ny9gUFntwkiFDrV3drAfJflGBTlrUu+Wicaczn+z8gFMrNot
A1CL1GW0vBvll0oU9YWKFb5OsNgH+I6m4FefyixKX+1PZf7QX+Osxx5vemK8SmXPrq//AzzAEhGZ
nfLEwnWv6YB2apZ2LacsOln4u34GDG2VYB8AbFeW8Y0sRgdo1q4ZYWfkm+CVm5bq/UIeuoRMmAKI
0Ua7is93j2M7DxUhjVkSBOkgPb+E6ZXXaYtXiWYckGdwND/YwwCE0p1rvryWCWDT7sqkE9kjQY2a
RjA1+gIYsVfulzoB6phbwXKSVM/+if7mIXaXsP3boo1LyGfiojS5ifnMnWF/yrSpuSmVNqzr3vko
HY7N17SOJTDToqwLuZt9e3ES32xEE1zMdOXvAeLuKrHZhx/6Y6WxoDRxZYHIts7DvBQpJCzrD7Nr
e3zEUDhBt8eBjKz/t22r2AZq5fRzxDUij7AU9A0mFe07a0eVnJ6y2DbgybX8OIrmd6rEN4P/NoqL
ZVcCGm1F1ldWpKCKXK1fBWCKn80dQkxPIZfFBoYPv+H/bgIitYWzF0kTrRYIP2Z6DoYZIXnxQrFZ
q+Y3U3W9BBiNmaK7pW9lHiMMgcvVm8DSYGGYJ4zvwdq0MnBL7XzWAOgUpt4iBWBOgi8Wrgye14RM
8N/IL7bhiDaEZJnJ7qQjS7GYFe2GjhV32PjMzXByZCHCjl0/4CzVr9THtWOW08W1mOE7EVrluWJ5
fisNxTAa1o8kG+JAr6k6/1uDd92qXqspbvZ0sbfuZY+w20Bu5zXC9Fm6L2dwbIz7sp2dPm0Ti50L
wM7bErLp3hs043thCy6KLenVnwetIwosQyr8F+Y0zWgX6n1fW8x7izoFfbRlrTJ/UFJVJKpOtYBN
Zmt5eoPeYs3UMjKoNpglo35yUDGJcAaTUf/OYHqhWB52hRqPjvIP9l6fN3L4Dc5oxXc5X8epAJvp
x3v1Z6+ig9OhqxaCMxSonImHJ35Aa3Hb/zJ7b6nlxnez0UoYz660B9cAFvTpCmK6AIQ2WUVEZABp
YUH2FuXnbcixqgn3Kvg8bu0qiJX2zTWuUDcf+ZbIfhpoEo3F3fXKng73jSp5KuVuF4UbDtLNkmLl
kWNlvgmwIGNO/tvsQTeB9HqMzLAlAW39ewqIY7zA9+xmeoYrvJT5oSV+b4d7236Pmx8dALbmmEoW
guC+dCJtpc7r41hQrzRxMayUCXVJFjKtn/U2wiJqF7OA0uAIfgLRj+oqYpbuHRza9iDkFrafHJ6w
V3/WFwlhZZbA+3o9aWreDOmTOW/sxQ2lY4CGhDx69ZD5VDp5BTlDNGyLJJYki/CN7iZqmldwVll5
LXf27ADs3XSiJ26XEha4FM7r9GV4xjKHjmeaMjDjkzKjObqt2XhWaw/Pslp1qFscGrona1sBM77H
WlzFsM60dGycYf5FWJuVpa5V8qZPL7YIsgZptODMUJ2gNdlMBEnDCQB+eSjS/n5AW7bruvhqBrfh
IadxM4/dsABnH4qFe0zn/KyK7reFIzEw/z933LSq3Uy+lnMWeILl1bJQ1ypHw9zuqOlzNdvPyAft
X9ITSF2a+PQwawc3tkAAcTr+qkQRWZR3M9oh/uHkomZloOwt7b0FTfRCJ7U0e8+jEGHrtaaMOrWo
PJKU9ESPl59hwqE4DyPQqrYaOvHoRzStJ1u5kOattHRZB26yM1cZSX/C+czTGgWLp+dNcRKBfppf
SO7N1jRnwqOfl2MFfzCQxJAop5FZ9PYRLZOagYdPaGHX/j84Dl+8UJX152nl6zieRSiacyPitm6M
wh/8rzxILMXaIR7YUeFf7FTiBxZ2Al1lbo2X11j3d5ltVihkDVS4fSCp7ff4ZettlL/IB2Zjq/65
PNopFrbs4IZ2YTGZ5shsO6xNGyCcxTIdAUH8uEYQ2OdXVj86nFsxAj+UxV+0tQW8JDuDDwUllhAg
gukZdj4zivSpLddl1V7ZU91+e3s+8U2CrO9SaevI3Eq4UmP2S1SS2eT9KJvgGVhDa15SbVWcqXr4
EdT4QJS/U4k/8dkH7jq9VDwbreXpxbUWlgZGz/h5u2eVUREQ2T+AJiREc/M9kLlPQT7MRHNL6QDW
CfGmVhz0FJquj4i9RO/Cny7F80hUstsQ/JuOfdR+ggYyatapncMwBOJ7M+P/QIu0A6mo+UW3M6CA
lUdD/T9j55RJx1KWNubXmNP7nMboIL/enJmVgxOV9iLqKbLIb48Cj/AGhnj/30DwbvtZAqPUuXzu
pCmrl9G7YUjDCkHXFCgcoiNHDpNdajrcVrHtKSOTpDH13ThQfl3zq04zbayhUg5M+50W17BKVdMm
UXw88KI2rTNKVb5TK3rPqtbqHBb+NoAsCysKRI5tCxPZaGkqUJpJA9WrgNm2l/2Lp8X8xrRzMKz/
ysxX5cEbpgBLMoNnfuakpeMaiHqvy1jkYM1FImfZW79cj2GZz+fKGa0AWWYiWa56jPOYC4zxvReP
Fu3kVsJmzN2BqGc2wEGFEjwYd7B3qEtIv6LsqOmyLcWrAZZ/cyC54G9Od4EjmXasRnJqHqPJoFgI
SWvN27lY2S6FyJtPjatWsrzWQLqcFEv8dBT2RXk7o+jWo47iFgkh2z2AOA+xom+2ED0lylIj+1p5
pYZiA1itu2rZX5qIT/j/aqIvnHCMfHNm4hHMGeFrDrglNJgLQDpCxq8PQkKU1cyV+sh2z5gRF9T0
GxsYWD+RiKiUQHOJ5gg+3jfeEim2GkCJUwTOGjGnaw8zpouUjPKbHclNwvCByRY6FeJlAbnjNIYf
DdCWFeTUdqMlxK+HKrkbf/gv9EtpWTEqZC0SpYluiN3oiHh0FP5ZrVUD/IG4/XTFih5LfqWui1th
G55DuAOp5mY1H/RnlIYXul3PS8iztLGX8UUvxEaoDPyTUes82jdt06IfLZiMMsIbm87l1xjJh4jh
bjgElWxgfFPMXiIRhVYJgNVvvJc9B9aNVjhSpkvp6lX5DPQ/o9F+JO/2J8mxfzjubm5LsG90NG8J
eGZOgu4Qdvf23X74ShX4xFBWl/UUeQI8Yb49G6OSq6LXAZmN6RYeYHQ+L6PVE5XD0BImSarjq0gM
tFR0D3nudDplMEfBeSlUTiHej2uo9ZCurgpjPIGQK7SThsZk3l8/j6QTVKVP59hMfuROUP0auQiN
9EHtze0w/qFkmrJuNq9bGDHWpUsZGI2RdzsLnS5YUSA+aU4ZrBEmIszAUCuKcvv+BnCwNky/3mfo
BXzBtHCF+On0NcN0I41j+OE91kHHL5rMndvc40LqBNVUPIJXfxJZ/2Ne+LYDDh0YVWHxrJ1kWdnP
EXwH689NIaWjOLqXkaxi+XeaYhkhKOJik5yVYf3qWxKDudRPccDazfU6UiRIye9KQy8iNqIE6r0V
rlW6A9P4E2+RTZXt49iEiAWmqwugt60ShzsIVef0Q2EpYJsp6awT7AwqSIu3QpUUXerW1/S/oN3V
gUNyAZyJZA9PPgcJ8E4b7K6exwJsoNdv44IbOmuvuPmyHaOZbrNE2VrV6VfrnpgZHSuBWTtJY23v
Ydy/YSwKpU1e5tayxCewE7NzMy5DSizpPnl3QODp1lT8lYh6S4jDtLTL7eivx8ZnHRhGv7eMh5p3
T2IkisCZ2xAA670q102b4h4j8cPI1jmc5m96iZ4PL8S7H6iBF7EJXHh3uewkbtwQGbWfLVn7xv7o
jLTVHvz4y4Z2Xp/bkICKPoY0jvrddIN8/jEk+z7IECG2AyySwAFZP/pz0/xsKFekfdVnk+SXsuk9
V2CNn9ZSieXAF2sFuiXYWv1wicDO516yKuKXp52ZeUIsQxMnHnpn+NDeks81NDhA56xWGn0rkaYp
5yaLFOu71rJr13F8kjz14121l6+Q4sqv3NOUip6YmU+XnoX8qGxd5qeBXx+rFAYIC4JrxxZKoqif
cjtp/qZCqi2gqBF8iGUmO0z0x60N5VAq2H1+Oo8bE3JQ0hExIHm3KIXPS5LAXZlGwzBKLxpT1TPT
xw7ilgXm7AN2jlB+7y26+O23oGja5zjnBWKwWdTN2QamOSVAltJdGo/nDytsj4ifPHMR06GxpfhK
9GezsF4mCIqC6/02MkBkZODGx4RMFmGBSBb3BwdIcauSuQ7wC9DDjWCQZ9kug2py22Yxz8W8hAUi
TPQOG08I9jTLt4h6poNfEkSuh110byfeRkvz0Bj+rHMfEPQh6CTebmWH0hcG5XBG5ustWumJUn1f
njrU8TNxnMKEjo9QujDJwKkvAzOY7fRGMrzXaXxmWFO8l+GwSxmHTcjTHLhFbOqlbKezf7ifgwd5
QUlhoyLWku5XAehiQDIHgnwiCia0MGYngWG2aeuga3cVKd2k/DNS9jpsYCziMNd5bdIfehmYl+eo
Wee8nXyUZGS3TKH+poxoIjUDoECyxBQ9JlU1NUHf8+Q7uBmOpIUBsVprpvhLtbxPPgnGc1ueWQeh
nY5ukW9b6WkrzXsheXzSb1az+NJdh7JNGtD/vrPWAR7Os2TfQByewOK5zV4iBbZhpLL+Uxyw7snv
ZBZ0ztCEulwSPzvLFqpy+kipaQcWBCOhrnbK/W8K4oXdRYlB15I/gmRGV9PZaUY5fMj7hG2WMzZG
Fbl2p7ZtzDXIYX7ByzUOOBZZnnLkcRMMmwBCHi5wNSyidaQe1Qdz8KgEPcesdWDWwC1VGYSdUTbU
r/84KpoSooUbxFcIIdNlLBBYopjp2MJ2d87PMMRBYRj/OOETFWxhItMUB48qtF49KjrFuUqTjRvH
u9zFfsk1ZKZHnAMMyVmj3b2lSfQaxeIlj7dbSMnOwcKKRH3VP1YsPcC8eXtBI0bqe69xBUIsDVkP
dOltiaRFsKvZYHqXPjPNdGaOrOvgKpKNiuNu4ouAqsQreoSETu9iKI/LtTUEBsp6x8A7thAkiyTV
yPCZ6AGxr1bn4csyUYXpG22tJCF4qWJgqyy64GSCAeOTqjyssMpGU1yu3l2JSv9dTNk8LxZBd7Dm
uEQKnM/a+5Sh+oBaBdzrf7s6lZV4VUNnfOcEzTcGQF/ihAZ+mDyE9xpi6+0ZqXgherNWjM8HGkLl
oqE6KJsE5mwWrBBaUtWpx2VGOBH1SRcLXvR2Dj3QHk5CvNMhtawaW4SbHeoH8FtCvxmtV9PTAGLz
p7MXohoJWREtBZA24HEnr+MOXW4gfkuv0ZGrJ1kllGx/l0Cjp/OTJ/PD2mFVYvpMqyOhaLm8DUVT
WB2VGLs1P9FP8J0d/+bueecwbILdtWQmN56kYYHfDzsRUZ5GJ1jPFhCZSHwAYDIik+j/kpWlX0gY
C1wsa1+zWh9Us/OnUmPKZPiOfSclwLMF5mURyLBSQzbjnOpqjcIlubrYz3PzpeaOy05MtdGzP7Ge
osq4WEC6juUIlHKSfIJWqv/B3WX4A4vwdg5BlHpSX5ZGsnZX0lPqgTkMOS4g0Oq1WRSAQTGYZSOY
JOCFIBBziRYPXPAxS01/3qcPiepNwJ/w8NCC2wkjO981n+c7Dzy2/ppmi7+vA8UX0RzRtKcABZc0
pyZxtHROYEgcCmUVDzVV/mG37voct0iiupcqoIfNm09bR9d4/YHzaXMjrxjLLRCa4oBuU2VrsKue
uoIWF+QgmSZj19zYlWpSt6vd/9D2CjzT4jsc1LOuRbGmiT0bfCqtcMfgqkhp6M2LwWdXdap4cbkq
Mrl4pxFnFhuM5vF0v3eis6ombjJvpoG9hgIHa6SzCNJwP6I3MubVNk0C/kfdI/LJDmpUgDGztQq5
Jp6GLJZu7gF6p2O/FMPIy06XfqvnmsFva5vWekq0HBAP3W1rdtGbT9mdBLVmPECIFtevtkrjKL9k
yCInIdLpMSV+OXX8fEM596wU155OacdQUAzdsA6ZvJEnousYBf1wIsKCRCcFf3mZv4qYTlnX6cfN
z4kT8KzMq+MyuFsg9ylpmLgLnJjGILfWqV2COne9Zq0cOtI/VjAQZWadItkoxPX+rjCTwJfsOHD3
whd6MhwiQXzAXwJTHFsHMM1XJyUFQXLXWM2h9JdAoGNyDSfqC5fK+YXi4I4hM7VYlUIBV9OKmYpI
jz13BVRNoyuzE7jMwffsexNRgDgWgYwJu/ebH6sDnvlTDiqjNZzwZnqbG2NVxhUoh6s+DrAZwr4c
TxGFE/WmriWML7hpT0Tt+PJ6j8b48KL+UzHuJ7ClSF90t1Lq4Cy6TMvGmWPrXlihTY68infH1xxW
o/OEFEyZiU1nx+AmjS+T3F+Fgrcc1Ggeh1Her1g/RfryiX4Q/vx5+Ant1TDme2By5w4ozV12fmYl
DxNVTqxlKpWVJoMY2YRV1G4T4TeFpFGRdJs701n3g41kkRFMsLn3JJ71hht/wDp5pzE+jriy5Vcs
dHeGVsNAsMYhlJ1nWLWXQkZWq03FFNOLbcdvUycRzD9I7JgeQAWXt85EZ+lnQrOtSiD6Wbt5eTQK
+HVn8OCmG7oqETyWD/NvWqlW96x0qgjpNeoD2oIX8vgMf4oTuNJJVhF1rA9DTXrmOIBdUbAQk98O
Fz1lmZT+x49jPBDHjl1CJLDit7tC6xa3LBON/dc1bnYR7WXVQqnumbX02iA2uGQt3c8fJ2n5R7F1
LMrm4dBV8NRVL4FsnLdY6FwZmK96tIdv0YSYGpNnJyl7PghJr53JC97AOtUSD0q6LQdfSrShQyMl
ynB5znYJCdfsW/EDEwWU+jr3bnRE2GYGsrfMHRjkpGm8V1M6SIKFHOqe8x/XSeU+M+FQuTEOCboh
dY1WSE5GHm8IF+tBzoMj+S7ff8H9NXpNX+cz2iHBn8cM4HZss9/+Y58bwVJGfZiEi05N7LRaTe3N
UVbyCTgpY4DhAYTY84PLF3a1M1v0kdnIofcg7R54sOVJPyxQ3tWd3qk7XIJ8cKhlC4TdpAQryzFL
vBHiGEjD39pu8p6O2tVxvce45T6MSp29qgPwjVSP5vnahrj+5ayjiCE0VNWTo/Ny/z+z5dJE3ftb
vsq2N1i66jJ2DBP2sKvMaHOl7DSqcl169cpyGbN9NxMeG54WJoWTmgC05B1+laVGNOk8Fu9TTSXT
mUPrAinYGZyCNXdIeX2kZRb/62K070GuvhKsDUKm8ZJy6/eY96Kj2B+UWbnVWabLk29fYKQn58U7
MNk8t+AsNMd+oPiezgnuzZMIhxJvpasujKY8xvGSVw7sF3Eo32EtJrpNlVLOH3VvqbKxqb8ccRJH
u+Rb112V6JCA7vM13+CbJfUxzI0gAjlrgPvIeUPVj97MzIptkjI0lCDrIiNoAbfLZSLNdm6CdAy9
UwQa3h/otL6DCx3Ouz4TNj339fAPtY2AdxLM8ms8h3bmGVsSXsYZcszduGLnLzU/wO4k/NaK0cqn
CRy7pkJzcYTJuGHZvkMOHAA2lhEnMviH9d6c6b8IKNYs9nb72I1L5vtiI57bHqxGHeQg4zgm2gm9
gO69854znlX304kYgyL0JaFuFvjAnVNDGeyPgwqd2krvTK6+q1M6j/Ur0p7TebhoLCz4odZM6DaB
DnGHD6ld8k7edntKub8PaRbRQxvezZbQumjUgJAef2NrGQYlN8/ZwNQOmVDFIFWTVSjl6DAoOr11
ZY1qFh+ihvLiIc3PqSA3Ey8EvDdfTYXBBchMKhNfKWhVM1G06XdOB3NlkmrHvhBRAIvSZLQj2330
EhPMtdOfdMzR2NJSIlKkZvE9ZktQ3JpPewYFV3L2UIPfjwdd0vfZWv71SKl6SoJqdn6/JQBjbQUi
F6T21FG+4SuSEf2wHzThNbHMh373Gr2GxKw9fzka2GGhOxRtJzd5HyTQBdvDVHTsZb3XEkrL64Gz
IRAMUeE5ijcWgf3jVDeMuAstDwX3bufZmfWOP+tj7CXIIMqeRTSbr83jo7DhRlqvffL77E7K1bXW
rTUXx9MjWgJrf0ntAdQv2FF32+YojVuuSPEIPuYGcB6KRs1du1luTr8afHdYQnsC9MUNHvpPeHf8
Mmgx4ZXQIAwwni3MZUKiurwWtRl0JUn+0AlqwnQLb71ioTGfd4FhlEmd4oghvDTieKqkB/4sD3mV
pOG+OR4H8PkHaSXBX6II4EJyuxtOIQrWWSLY4pvAsS1BzoiRf3QkQmhJ//Z9DkZ8kGUgXpkem1Q/
PGYJvfRnz22Z7pCD3m5M1v4+0GLjQWRWQEPDJxN1dPpXeWHE5Y2Elv6pIigdoXYvdJKyVYaTwn38
hIyM6t2zaorakzOMKsq0z31eqIpRLPVFosYFGt4gFCfoTH6IPUVwHPbVIt7PLtWgzCGTpXuFWlWf
pk26yxqI9/8ffWM4BAlYQqOjNr9f1sdrOp2GCHZZ1xgnMsYzCJX0WUzwTJgxxCLsZa5zLaDMhmZ0
OOHaPIpENfK+ClTicTYpxPMjUEsp/e/AyVJLqcK0iLdybMgvfyygzCqztrQEBb1DnNbgbz4xNh0Z
fFuhTlVGuVfhu9kJjtXdQAufj4l/geksRsP8G9xd9bjLfrqb6Hx+yePoYAhmOaMcfYJgQgZSNTRz
z7H2y4NjQ68GA7EsJzeKLMiysONYlKYAtmT02rLuqseUeEtjlGZpsQE6eMRzSeqlkDIu5OkpaJW1
FxEEicQ0/TwchueYNCfI/DA/TNk6pyS+2REX/+DLHZixGUH3L25M6c26q4P1bE2OkNQdRGN9+jg0
Yf5q8kqjqsshATJ9U6aPakCZpd56h80tQg+x1ehzq+kegFxJAXBNUSi7AHvWmz2Gr9FV2xDde/j5
8v1et2RVaaA0xzY5N9YzNsq2vlLsZbEkpPtAB94ywmMdnpK44XtXcApMwuDCke8o4XElU6hNgjRg
eFM58fwE1y4c4N931E65K3oUDVxknW+6RCDDGklDvT8jp/y0PWNYkpbcDAGG0ZaHw6GNRA9to2Lh
6AQh3S0GfkMcWhzybfQANBFa0sgaaAR/Luu6T1nfptNMnclhkwePpRtGfkOoJLW2WH4RRmqlrMQ5
kWNni3FWUpLMFy1n0qnPkI8vwMxHabG1B0j+oo3ORaeh6qNLHboV20E1BLANMn7+3foExRpwX14Z
vZ/DoXd0LvUu9Gck+k6T2cVFv69aPDxmsFaaGbV0xA38M+uUHP0QjH1DtnZaLMalV1sMvjoxPlCJ
UFOX6Fk6uviacy+iQQeLaTv9N002pQZ5Lna/qamEmrhynxQiAi4+q6u5nmL3dM77f0XvRyGzKD9J
hMniSQgRtxoDtpr/LNG7QBUY3sOVem5Z5RNk1mmsuYeRXlUjHkZabHSMd5LOooJitvbpwrtOQOhW
LCUoA1mZjIjiFOq/fcGPTl+qsZR9vdfnu+zRrByw2GNSR8I6fq1WTqKlgQSFIWZiQWeWWrxdaZjl
s0F/htE3RgB/EccCS8A2mgdBb+vbAPwUDm4nPffUgWgxrJ8KQiG3t4v9YBbbgIPyswgyGJ9BAPnb
BcNtzCaMDSbiro58+lPAAQr9nvLoLc8rNgvriu68P4Gx+PlLG+nb7i+vo6KAByKwM9q1e0jn0A/B
HVvTBveE7x8EhonnNv70D71Ikf3B6bdBOLjt4vzVCS9d7CUDNGDQ1gl7a650ABvfjwGAUwjxDWjl
ABp4zKtAJUevKmhD74eYPHSpxW3rQDsNfrX0EUOWIkZUaIsGqGLtbBTAZ4gISaCIPPOOXfiDsZr3
KMkUAuRA0wPhCBo0dLk1Bz7CKlqivwdafTsiND7iejf4uD6vRJP/0CGhBPf2xI7yNiWkka4O46ZS
GpG1fszR7ZH7rkbqjz00rM4qmrUm+tfqCB2QMa/9SJDlzeyECjEiMfNZnr7J2Zzrv4FUDnt96DZT
Thu8g1RnOoNh3gvyJiTDiPfQb/0DPBDhupmhntpK+SDZDp8KPi/3jbWFbCKcNc2cOm53CMiYv/mP
AyNLCcoLguIAphyRWzFEjCXpDiCqjqhTB0mo46RMJVdr4nSkHHgcICtR8vawdNRsW89eBOEe2ANu
HwE0RidOx0yYLGpKckQrqAMhQMlpxL2tTYb3rOSkQQ3Uxdws+B3t8X79nTkjKgAvlcGRjANNHwuE
boCCuvm6ueaZdp1DphwPeV15DgiLzUatqB/OyOkm0VhpU8yQ4dasekvU6HJ1RzGyvXgdwKcHRF4+
NmzBOJQdQ3Z0QGEluhSWVxpL5u91al2aIdlX6wpMZTj0g8FDODdB57a9o+QMY7XF7frs2Vz4wwdU
deEDTw7rhMhho37yfz1rn5+k67tLUqmY4NUWv1DyRi79/6AaJO0GQNx3igWaLHykLVa7ecBksYuP
YeGOqhgu6Xla/SyX7VXJRqWQOlZxk6o/it8A9cgsKDtT3/pocGGVF3MosO0LkVkaoeCFtMwPfPDn
huT5SqZXmwGhokUOSAgJgxNtlvFI12PrKGZnnrVPZTGN7uKMD74Zp4WqEfNE7OWsfRAbC56aqCuL
Jcbr1zsTWrN3kNItHuyJfwRr/Dqstz0ZGD/WZ1Q6lbCUbRnQvv0t81Re7e2u9PTSMc536cWZu4FH
6XVL9iw3OWVsrbgnU+T2D+nLvWorRyEhF5Qhjrln76+ydaMNY1YbP5ByncEwdufnSW6p1DdckUQL
X+xxBkIQlhYjcM416NGXiNVDrkfFxBZ1A90ZsQu6mYbyh17SbBXIuaau0FOi32PSAelFiYeFiU6x
XqqFnMqB32Ho+ivEiqq49Lk6dCPtgKmtRXhIVoL4bUUW+CzKahNQX0KeuSNIPgNUobNmnHAnEzp3
n7SVE2U75xgrF05VY33L6eI933rhZfBLYbPJSwjxDuds0yKvw465iffMOrCXyvOXBN10iYYcRqdt
MuyH+e3WaMwSALQ/CniySVqvcp2cQzPeuuRpMmEGZvR+tLk/ElAaJ2aO3Yn8QQgAGJ724J7yh9Qi
bmKtvsS7KW3grGRal6Mf/ALkKpFDgT92DmJ8UeTRD+iMS5aen9IFJZcyZIWW+GIjcntJTDtxp06s
lv/1epNNzHPKwqUXQcfMgop5//q2nh9Ef8EdJxITEXaTgEW3MIBeJ7PfzAZPhF/w4VKWvF0gnKxM
u6Feoto2YYQ13jqtwtxez6adsMJyeqtnoHzInUs25p1uEn3CQ1E7kvUige+YN1/hnqPcEwVEBeRt
AcJhBVQKWSmGSOpaVupQ0pbqadwEbRx/3SHtwKP+ytlcDvUTCO/nU7J5WdbeFFjXVLMDpTXoxHBg
u8E/3ZqxLIdmkw6ZCYuXJnyvgxD2uFbroVgMzeRoU3+oyq6X+L3FBBgFZ4oBQlcWAHJcgpx7gTJX
7/FiN5i02GG7mpjRWub/TmhdD4r9YL49BfMu8zax6fuL3uGsgFtHh1KMamgKvT+y4xvl+S762slF
BhG+Aohz3tA06uqdIfrfNqajbK284N3xlMr+0hc49z9Yval+KxpGICAgteitz9ui9h+cZ1djv23u
Ll+5uXH3JkxL2/NrkIvArPEM60SGUixrGaSUhbI6aAUlodL9tPm501g7MK0uUCUF9JdVAUcIggIN
r2nLUdfgX5dB4yqr7OlOjAmtkNvSiaO5aN+m7SSL+a8If3mmOlaaq902gBDkg8fBsmIJjkELHfmh
jwV405ERm4Jqmk+b4LBB0CidPm0YIzJuFeHBDRo9C7DTjP3PSe6X47S49F8W6jLONwt1kLvlYzJM
FcESCXt1WdabyVWE+0Hbmab/YTz/JJ0tabUsJijvimkCzDSy6mNmPcU/m/1Ekez4V+sEkEgTsq2K
rhAT9LVCpyynslo1bIbm4mve3LascRHrWcvhPiqkJ4PwwfbTKQIyGpJSRx4YaTEQXNHzV9RVZWL8
+Tgo9fVeyC2OBpywEPwxK2yiLooELvT1BXapdeRoms0iGmH6+YvzS6aESKMQ/ZMn3XtGgJTwDxNd
DApfI3zFPKRoCv4odUSBKKHLUvo/7fEOspdrw6PmO5sEGC+2zssVqJDguIm/h5w5VKT+t1wkfnhm
ST62gog4bzgRyKQOH63Sx0wTXSG0FLJ3vuTHfo2AQBC7S0tLaOW2k8+GFel07cosndfB7TxYh9bm
jknWURKO6hQ5Iyyes0Vpf269576it9Nw8VTr6EwFj/sHKu8N12Z9yAqnzoWSKIB1IUFyuj47GTMc
mZmazzoR3MyF1RRXR/KeGhnamhZL3QtiPUxQM6klngetSrQbOcfLdawQih9/4I8ZnN1UQcBMGOdP
ESSY8/LkAZpE8wi4s90qjlzq2u9SQZXGBmlPdp2NmPbIsiOaq2XW1qEthp3jJ/bx5zskad9sYwD8
69Sml6PQYOyjUhLEbYUx0q3HpOSQWj15SMKuGC1+LnLw7BuMtPYUqBqRNGh/yJ2Czn0IK5ImaKpW
2IZ6+N5j9mVcruhBvnnoH9TTaQbN5Mnx/kp+9mQ8UH0pY5W033v/MYwS6q0psaAFz3kOqvw8G04R
p39P3DvB9so3FzY/U2SfjMwyekVs/x+6HhLPvurzSaMDlMUj1i6jpvIpzuQqYBtJyDkqAOfuFKu/
xxFRmAI3yf4EPqCNzOqQfJsctdxnxmmeIqBkz6BO4UYD23q673RvATqkwpprgcJnamKvEOqs6LvH
jzaUrcv0TtXcFUqbqCp2bomEey79nen/Nl5L5HHRWd9EZ+V3RTDzE+fHCuQsbj5glJEaRu+y1wqw
rTL4jFF+UelKSAECxDM0zeM2ZsOTD5X0oh/0avCGnovXGxeDlFiKbJ4pZ8a9+/ppeJ9ovhIuVffD
Do+F0BAH8XFT3IuZvKV44+3OoMYOnQDqoSsASG8a94V28h9jlv+g1jymMQkgAeFV1yALpXKn7Ypy
2WsUsOQsUWeS+ng9h0w+JPWekT8IyXgeVBIUU9xxBz/H2JZcZNUtx2BOEyy7JTJRE77VYoOIc1oe
75pXg2M7RSfaJxLMYGIonxwRmxMCSOiUFtLA2DBTE6f766QI3ddfhZiBwX4s6wqs4RJfdR8nb5TG
i5CoQ9P1fXRGVmI1+dMAXbemXt2eznJhQkQ/JUfsjl9ZpH8dcM1b3LRz+j219E2LNNe4stcuCYIk
1YNuKm3Ng6WdtQ/nzSowIOmIVU934D62WP31JtGq6d/rg5ZPMNb2Ve9T2AenhkV0/7DwWTGWKWvy
giVamMMVtrnpWyyw9mhITTQteoGNjCQXSIxbJj1lMWo1zIzhFkxSf6JTo0gVdLzaamPsTV6KSHvR
FfiGYPBNNVKpH2jsxmooaceW+EnvH48QViuaMS/QBiGWGci9D74y70/b4qApbY3hv/JVGrCE3YsL
+yj3PTDwzRFtFfKdHLeGfT8Ovlg49CDSTGl4d+JEIo6FazuDl0e50bUoEOorbQ88EOc5el+Vybn3
oi9Dng6AmB+e64cPs2dGeAehT+fcPClgWgjFDg/XJ6oC2EBnpYpY+KG4nN6MnCsYzyOFFD5hbu77
FuGgyUxqcRxx9qFUlBlldSmqy8Fqm6PZscIXTHIKy2+ERezr9UwWZWKhW4Lrx4EpYFB3DQnOjvKP
Zw6HE1Z47RPzp+42aF9XfFiore+2gktc/XFuKgqp1ECz9CJV/kuehvSid6oQboyrXSCFXoggiOU+
3HrgDIyy92FLF0AwmslzWUk898X5VD0Aya4bozlQ36oPSC/2aBkXzsVv2CA1BnNzxz8PRWKJBPBv
lE14S7Og4JfDARPwwJBfx6K6lQqAvqVsBMZfslfmP5sk6GmVfLmPNzkusxBMQM6/Ufyahu0yZYQm
DN+mMsVcfkt5ICpspziMc7U7fGAaY9nSz08FQvG+4ATvEysEspeEzZQvm/ycN/ev8mWq9EKVl1to
8UG44cY235WFxdRNPymyor0q6M1WDfqmiZsaIHgMHpdhbFAMCmbfI5De5fR/6EBu+429QnpAHD6P
cutNgpXoaIulq9YEz4sI2ZmzHbiMUWala9ATNBYNSL+xjZtdGa3OOyuSskrwuJiBSHy44ogiahpG
M4fu+LNAZGS+h/gTvHyCzMantwNT9xnp2oIrdfukytRcMjGC9gPc92YUXJJs3uCCwE/OX1PGDG8E
Mojoyyv4Q2wFcgtAAkY/GffGOabx/G4DjfaxVupe9Q+GCUZ2j9eBZi8fqJOQWzr31vAPaytkIdCp
QCIUC2XBTbpDHU/rO1WtRckq03Y2XOed1SZ25jx2Y8E7qDdyOJok8vmxvAWAYb+0D9IAJLjUN2UO
ZrcB425C4483t3T47zgnKZwIm4U+zm/kxn8U/tX37rTeAQgspXNc6z9DRDNg/ulh4FRKYjYv34ym
HkelBeudbHPhJ56RGu1FTqlLas6MsQrD7M/OR/2G4MFq01dI+n0b9uNgqWB/XZNv2pYuY4dILX9V
7ad6SurGkoPIXqCna2WL+iFy/rUVgF0KG2MeuYH+cNpFZhokgs4bwHW7KcA8w1V3trIWMcCBBgQj
A+yNA478jX5xnGJ9qoWeE5YAkCnScZc+OUiD5+D6aQrZu+18hxfFikTc+718B5NMRVQRTm4IJV5M
YlwrJftO1SvsFfGLMCWzutAhY5qWoIqU3eS+vmU2tffubhi2JqGjpJwtj/dtGScg7UiW70Q90Uz8
COdHbp7LXWiS07IAnafLQRazOQWYRCW2KfQ4QtmhzZlWb9uHbpHq7XYtR1ZzPxDWytLgRetEdCQt
MqN6ej+8YQMNPG2Y/XCbILn5d/fP3HeQDTkv76JNBbvv6RiNtSUKF91CHfmGoUVU/twcFrzwbnIk
GqOTflhJOrvxJg41RWPyaeygoaHdQpxJiWvIvTvGinsf0MKP8zTWpNsE3swvEKCqNIyXtf8Tp+VD
UpNyxd5ZTS1N+3MaPAIf65mG8vGyJfjcZ7YkfFQbbCyFoogETgcvyyKKd3aC+d6i4pDZpYnYDWbD
XfTPtKN0uAbLhcirCMPcMf9+EMVJVVNeUwgVR2G07ADX722B/6Fe6UEMLZOaC51FOfv72GiXhjqM
k/VeC1NlfXuPGBIJ8r8YfX3yQJwkDkC9khIj0lzYuUtaZ+A6a2AMGG/vXmsWjtE23JKxMvNwSVEy
DvS2CBeLyuWmnuW0ZjvesvxdNmZgbvlrXxgIlGNmo8boSYZLnDV3fTTKsxBAzhOZb7VozyehSHb0
cUR4AooY1zwqJtwsuTshvKRZD7Lc7/ztAKHiv0oj4Jdzho/ip12vy5Mz7WBl4ko3vvjt3DiNTZYW
2tNpbLmcOsH0TMvDj9JeoX0g9L4NXI4hyzVaDF3YuHHu0aquRKWgjePEJGmYB9H0bG1x02oWd4ts
xugKLCsyKLNe2j9LJVIgkSxFQKjzB5NIuxxXpdHNxzWbe1byl1ZpCXMl4hSo3U6FuW88WWV4Gbxm
zE5fHDrEXM4i/lhiGExirQHtboqgE3wgMHWzdAVV9XFeZZIb7j5p1ulpTgZFj4Xti7VeInMXr4Mx
gI0afm/K/4mJaqdqimz92FFqFTjuOMBpFA5YeURs208rXLGAQca87cX9jpAGDGqYoWvUHtPPEG7K
tdzdVwLa+rIx+fTXBHuSS4JnK3v1Zb/w3UkMCD4fSBZUdUUKSxUQKvyQ0WaxvHVplMozuzX96hgc
1FH4+QaE8f9knkh2hXxBX8FrvDZe3rJwiBTavsB43dg4JWsYCwxohpODBAXdZNB8njcZSZk99lR4
oDCWYalCjXHbrlbbgfwb4VdZlcsvJ7Y/veF+uoVdBgnc8UZ2ENxGuIuOX7By2ptHT0FFSq41Vhss
ZAXD1xxB/lRRmCpPgtzdKHcIlwZDjdXLDHy5bUSuTdPBjaXILZKySlC2/mN45l2KXYvU8XmNEpfp
1aZX+/yYbCWt+wpziEbqjrv+msiqz0CXRTEpHfxV5jUBHiu7G2divjIp1a0LYd8Jqn2CsmcrNGqd
9g/+FmcbjBJgX8LnkIh/r6Obcdw/FzgHncvKQ5HA1LHBgqdtKMblaUO6W8pGixN3GHUtSPKsSQUK
sFiyQ7BVlEQ2UUDNJcY7SYVgqeLDqxw0eWpxxyJdnKKReMiUT5MK4xOB9HbAwaz9NRB3BibrLCYd
ecHOxmjJCRp3fLHIkWTxgavkhUjREtwRgHwMsuG/5pqIi/x41Vaqyu84K64m7Fi7aKcauw+jI9K0
4VAhNoA0JIHRCTA6LUr54qUDsvm5IhFZ/qAVfkGp9rXsTirvmicnImCu0usbbxIIwInP5/EDlJmI
lwO47ZAOHwGQKNDmwLtMVGOSsTwVGGLFAGESy78zm76o+9RUJyiudV6Jn84G+kOg+knM++XuQQXp
g9HbH1ut2B3K6rJU0o1OPPvusORIrAD6CSWqeDggiR8vd+dvTCNzjuEO7dqVOiHTgS4B2+liz66f
rTkRMXNmFYB9/MgUtjpL5IMjXef/URm86NLep/5qq/T0Ar0EmQPqgl13QJDhbGJlhAm6s5BGlC+6
0rRoG6jl7w9b44/2126pgj6F/PMY+a3LiJoH8isfcSH+TX3GcRqTg75EKfvS/v2JHoFY8+Z5ynNs
AqOisEA9u14hvt1nGVxWXQyONev/ZJrnRjMDDK+cJQ42UGSSz9brqI1wFS2GhKLK+txEL2WoY0ZE
bPUPkb2hW75FfRoGi1VMjEIs0kWSBWSUtJw9LwXk9sjA8AVlIlIImSyshWE8LOvdnzVdI9CyIKnw
HRsSnfy9U3dC57Bu5q4sfdM+Q3yUtIe+fs+RM4mbChnUl26xqFIUXKzQvlhwfD3MWgi1kscRpYM+
NLmVC3X5zjtiKB1vSS79aF0aJpl847R7gqxHHjFwWqLDXpAd9EX3FWEOx3bfj0GzquRdSl01wlmM
ugEjjWuhv61QA8tzQAr+lsijWMnrqPMtS2hfmDFF2YgFk6XGCkAv3RwFeBCTCvsccecURXw5FgBL
wfB+7N2J6nfiOqMM8s1eATbhTsC2xRUG7gvR13Glw3/WTmXzWYccULj/Gvufl7HvErV/DeyKZPvE
GV10qcZeT8mWrUJTteQTW+QVZGJXgqHuytkAmNCegv2k0XihL0BpO6WHfWMt3m8ajBpJNqn3Ru2Y
iCDUrh2PY5ANwYBtOphtv1ATAVsbHJlrfPMquMTVW0dr93aXpJFpLGQqe1SLuUva7+OfW0gia4Z8
qlnOo/PshlQlFX8MoqG4r5oSa4Q6dFSY21MRa24Yn2J+ya6PCERIVAXJbiY0FM/7SLgHdRQKrUVL
RiQwjWw3iK3G+KmQGmZUXMqvXUlDlT6oNsuehQw7PmPCH3OAfsbYGkiTxHTTvF1R5BZpIMJNFqbE
OMRQUMDQFhVFyVsENszKX4S+cWY6Acty4Kl377BZB7OCCJvGoalRdUIe8SUNFSwQMQo5Y33kDylh
prS7c36wXV+uibNHD4aRwGNyHMBbe6pHp1j0MnXaSU1xphfjbfO+JjxyR/O2Yq5wFT8Eq1hCu66u
bUuuwrq+q8nBQE4tYpKQNeqcH5P1TMMBZUmKSuyIoM3XTr5aciRGMgsZzNrPWW4GYPDONUgJQ6WO
h7q1c7oJF8Oyl/it4TXU5r4exvhC1cPo6DfJZv7N0tJk65/9WSDM0xNj2HKT0q7raWVBpSHOgi60
2fAEUZL74pWM30gi4yxyN7Ubg8EevYFZW2C2BCJgYhS8QU4hG4zbE0UU0M8jpNW1YYbomaSlQjAZ
5kuhZ8mz6JifpoOZT5dyRcPtTZeH0M8AydQE/8ZbZQbL26RTwX367fhiwQyaMasF+T7Aos49WBmL
Xw+us80MWF+fV/Vpd/ZNMUmEqHPRHtbBrOMOrNERCocRjnvHiInd3XnWMNFbrKfK51RF2Dw0Zf3d
vOXY4fCY/u4SbVGJZ3slYPaCVh7B+mIQzrtp7FE1EpTvWN3wN28PExrMq2tq0wDqLU4jLvtCPozJ
dLhyLmYeEsRRTqZ7LuBxiitKr7J/SyOovHcgjYO6fxfDIMDfKpkKGy01pJnDMqB4kkEWhy24LX7U
bM8RpoNlt2ACyM/Urs3I96W20SmWPTpjRfEzngr9Yb3j1wkbdns/Au3KaE3KYTYX6iaNl9KL0J6W
F2HrLuvtWNougIgDSyAFdXylWhlEOVnb5ktwArCdEoMe3Fyz/CxNp1VvuOoZ4+/CazFNrwJCsOtP
9Y/fkRogPENZ/HyNksZVhYNh8n5etJJSvm2F8xyjbMkU1ShTC9GN7N3Iio5u50pXBiLWJxA45PEc
kJttEY8QjMntCY7oDSpQJ6mybiiWPu7Bz0Dt+dAIMj8Isl7ZZBmML8N/ffDIBFOpKsTmH1Q0N0eD
6zZvpCVRzIEzQoSjIklQ7B37v0VfCIfx4KFUHmVu5rRpZWzHveq4//ThksORiG1CJ2uiXlGWh5N2
5RRDHY+/3VE2hsnTvVIJNUxOG/2bVoepgyKbi4cv5OqwHE47vh+CtNCKpOfqogaxiXvczmjuPmXV
/RBFXSkD+CfFrZ1VJlxnpi+YxhPEgGPXIixur3Ey4rS/yrqENdscW27gBWsI6YUZhxZm5PcO2ykt
KnlQTDs8Z1N3AygGh4uzFYf/FlElOAuZcL7ulW/VOxz8QTa6ILhK4jt1FJKLMu8W/ZEFdWGJpQAE
nzoxUZ25l/B/UPHlNszIhFbZEZMNc2FdZ6ewAf9ASIAiVMCGjE2ryeICzWGakOrfAbBF81u4pfS4
nQKHFpRadWLSll8Zu2edhSszVQQlPWj5Uymaz6ZdzfSh31Wimgt5mUmFDCf95kKmnvWQD2DHSHYG
gVoebq1ghSiDnorDdUm2th9QQLsi1hIR8vpKgqmiVk78+jLdCxxYw5xh4EAfKSY7ffnj3HhDHUgv
bJLuRuRaz0RvOubvB/f9JpQQBfCMROUhsDJIeqII3JX08h6gYVhFMeqwyHaUk+UygHf3NABYxMUE
QbcGnpciNodzRKpq4a+atPUtYNitZaMDXEUkQP40RS8cdnkA+xUhK4xQuCy7MhSHbmLT/XUfvVP0
/Dv0vWm7L37R9JaKJDfGkGs7sAGH4gkIp4EqDEby25aOVvCMtLGpBc20+bzE78nKmNCEYHtHJyVO
dZLrqd5rb5GLqZpSNXu9ntCOWV1L2Vcwj/o1WP1OO3uCNGRv+sEAHAp4ugNFhvmIIPeSjcdEY/IH
cttn+Jv2VEA+dAQ+JsM4n5V838yQi494aGaStggP2BTp0DEBRuK94FVMY8ZMsdTotN+w0p8TIrsn
6EdLOV1dyrDtCfb7phQJRrIj6yKaEPZ6HbuU/jI2DimU9Q/WXLYEpk4Wz3bgmS8ItSvMECgAKrci
7pn9/tgirTo+4zmxph/jrL3WSWRxrFIl52p2VBMUGVCOY1GjQ2GN5ljbtbtbFd3fJIFcDyn/9qKu
Qw+d2MKDMIgZhg1gUv9wnrKRpVF8fzhDt0kYbK+TvA/LuoxlquXQZYjMNWaLQGcXcQkGqvJ1/o73
VAlwnUAajdzy7pVWUQrmlWEbYpGHp+7vbVQfobud3s+gtiTRXZDLTCa7P9D6xaWZRA2SVJBmGvBp
iyaviueMrVX5jqSyAT0E1zt6AfAEZ0PaWSvVBLgOx7YsVOeaWsH21t7tDDjxlehnd9PPfhipEuNd
ON5GzM6J8hamiQ3TW7yX+Vrp90bDYdT/4qpGkGoCmjNsKHVkLyXTwCh4FeigPCO0LmWJEV7lHQPU
AcXdV0Hp7tfsbGiMvfDdCZkDx1p+PrtZtIKoLWaYpbswlG8BDztFHUbnvERafh9iAnUFJ9Yq7was
BBbUvi+GMLqIugJEwIL+M4zrb2PipD+PcSFaO4DUJlnraTrT2EmiYywSveGsYN7iEAkYNEvJjPsn
fzoN/mfSXNOJU9Wz/62kuigaAwt7EQkfUuFA05nBuqcvYBWkQasujZ2JpII07B+st/e2WtSh9ZJP
yPNq3RXQCPJF6anDW2f4n5DrmAu22PAek0l+Dggwhv4PU386ickrDeqmbJc50LxtHfjb/BrbESFI
h75+vgIQE6c6WxMSlbHb8STsz2SoTciCxZoVnSgQQwBOtdQkIEA6IY6whi94XZdewamQ1eW/YDX4
T4CAAdvw/tpc4oWQMyJK4PYB/mFx/AHxfdzkSWWYM7SpV+s3Nt5UyFu5NnpN5kyPQ9ZedwRZck1X
4efcnATpEq5eCqcKQxZhOMiNBGPSVXARj87wyKW7AexQOs+fRPUwNmjry3vUFj+csMiocxQvZ7/X
LmXLOtj84swN490VEXbk17jxxI38NW5Urgbk1NJ3FLLO3BLl51sJV/8X9grJ5m9Xs9gL8IopNWM0
fZwr4blGLQ9orcjfNaFg6lCiK4ZmDFrFCblzx/59TdbvN0T64A16j4ipJ1FJzQ1rCcoUHV3Ij2AX
FelQ4GhEsGcAfkh++syuCImd/iPYm6C1TyuAwzgUzQ6g1DyWMymq7pNSE2vGu0M7dZSH1DVqfTn+
wmKoePV+kEIauOHWCEvgWvt+siPr8zoFSMnuGGlTdFbm6Lpo13uFgToBl8x+byI/3YrruSXoKpDc
kPE7a4q0kj9mY5MsfdbQqfMLqBuoZhCOm+SAEa8gKzwzGgg45guuQbHTgwdrnBOy0J9Y4sT4MpHn
dRo2oXP4AaxspuNVy2wvFEn3K0g8jBL7xAAUXF4L+MFdvjDn6tQ114X9o1k7NEQH8EuBLbKMcHYj
lsleoxtfMkRnSlNeIBr6WesKs3QDX8jN4/dwtUnUl2TDaemWvVDQJkIlQDSrNgdeLucRSF9ypay7
alLahJL2J17b9dBg7cAKnIUp/iQYLXWbPFCYf/ZV7g/v9fmrSuC2EbqbuUVUFeS9/8Aby04QvX7Q
tKsDQxhZNg+ZXH1R0Eh8/6QYpKgWhai44YPxyOHLcRShjnt9zdNR/AOlJebprSUvbfUHNiE6C3XX
yUnO/oKQrTEekABNCFcBKwoeiVgGQ/hiW/FGekvAqCUo8SYg4pSlCCZpqcuqbmiaCmV43U5GnzQ/
SyDHhVPgcaqdcu3pmbIrEAOzMvtLhLqMmBfRbvWrldSvZ1Gk0oHfdnyXV1Uyik1c+mpxEsT9Fvtt
Znm5GsJ64Dbkl4MyCIzKcC/GB//qOvFuxs5qiRwjF9vMhpVwWbwtUcsWUqNNzrF05Yu9sShVVYPN
pKHzHA7aXGrwzRvN5kpHw8ZHyJb/h6GLa0yKaA1y+eMYW/bme+UFFmbv8k887CH6i+YK33TxjCX7
SrR3ZQuyWyqai4fB4fMe6FWmWFnIjqErDuuE4Dx0MoJQbqC4DyckO5RBUWhWXrBDN4lZrMklHLdF
LQdLm5czUlCRSueTiuDvtJF2Agulor+s50oCyY7JjTRJdM3Mq3Qt23VP4mjL9j4Kka/wQ3plAl8k
e4fCmXddJvjUSbUxQ44EpJZa0my8zaj+0lvQy23KGNqQUv9Fg5YQSePI0bFufGeRAemkNJtbaoLf
sw+sos8p/dRuacblvfyB24ZWvsY1JPGv84O2kV3XhHa8pJbgGkjwkJzS3/3yMPvxc0VVDXbAu/Ru
0J/LtcAIe/2XnDCgC5cwGPf5uvh0RYjwyNo/UV/7FB7iO2maJvsJP9tEMatIkwngUbi1NhWXNj91
SDnbumNC9Fz2x/601dTSmS2OkSMUBiCvtwm3Nae+FlBUrLgvR0Cmz66RwQTWDuWVsWE5yuHW33m9
m+kfsJi6K4KqRC11yliB7H0egSBDTmLQOBVbqHwO8li8jzCFdQkG4AveQQu+U8JgwCHmR1c4ufzF
O1cOPM6gaIFgymGhNQcpS19AAcoX/8fdkQD0iK10x3nJE7NUdyuZvapfQ9fKIpTgFXTk0M7zMh+W
ZLXT3q7QmFpjdPpG49PiHcxB5UeY04cSidkLcOk/tlovy0xkWlXsZSSwEL7p0X6rcwO1cgQKGMHK
hPDWOKjT3SOR4A/mWsSh/QF5QyYXXxwyNHitT18FQdNIVMKa5Ly+doRC5CR+WtWXT3v24N69Haqs
bBGhFFUMZ/zFoOoIbHFBG9u+HkT0s308R8KBjplk6lOQR03yPpt00coxA3mBGLHpeMk+o1hnp6k1
eGt4RN+0IRb+watx6hotyhIbp1kNIBkYLOHawzCkhM0XhCUYnx8zTFXkGk2ZczkxLP3UdflSvHSC
CL5R/lcfMjoGhJyrhGDbMndvYzGdbuLOOK1BXrygBoSWpEDI2ufQuF7AFr1ZBr12H+IKMstoAnMb
siH1m3EPgTGedvReFJBBCtam9ulqKjD1LlPoMb86DMkOfHZYmTnRq41lKdUlVWkyH5bG7qd7RNX0
hwaVqoWBDTLycaZGDoBSaOhPgUVMjTMZBDlLHhe1BwOu1luKqa3Sz8332DnG2tQptIibGG0vYUtb
l6gOYtzXdIcQLejwaqyqK5PwVP2K3sSj+3kezpGs3ExFlrXwvkCRD3QWBq7bwaeDEWVmA/6yc8PI
WmVwkUsd5BtK6kOKHtj3s0YxIofbCZhXH6+w2BvUknhkXBtajeXucACUm/abe2Uo8SrDXKZt4j0l
9IGdKg2tk/tuoxUxiRj6GWXX363wjxG9B/6jASkCQTfVF66KHD41CeSB0wX7yqeCsL++pa/Tf39I
MEe3W34Tjgi5TyRM29lgTM340S6otKkgnJbZnf622Y55JrrbRFPpADkBmesm8UkconIj326XH2P6
shctrcDoHloGQKB/Oc0H7GJeYmI4HCKOw+Yeci2zp2Gzi8HJPycAgtVS0mHY7+DoyKZvI9YVsjzO
YW1oveqojoRpCQRikdVlOSg3/tV+0QLO8cHonggQQhyQpT/5WD0D4okTzhHMYygFQx/Ns9YOuCq4
4dx8tifpcUDut2Dj+Olk1gBOQ6YG8UHjU2bA1g1PESNXyNSFrtiIgs1IpPpj1wN18jOb8qHyqRsx
T+FMpmhYeJK8uXYU6AHG65e8xvqgi8UNsBdmfKaELDih0gg1jV+e68eSKNXn7XyD+h/8Ma4Z8/Cq
cLBECZACv0eLU6co8wFI7bEJW/sW6zByELRnDe1Kqhw68adlDeoKctgmk2J8tUflWEqWanbYy5dc
hqTX3mXEF3C+f9YNd4ah5Dfzq9oiF9Ea2/KEfwpA1dX71UZTrKRvkJH1vwaC8SjjgrunV53IGDe0
7gs7SovesoI5vuO7ZASABoP/pKITn9T0aRycrbOjudodr6fubcEqI27A56CrS8/gwnNdFKr0DvLM
Kav4i5l6TgTpRbCx+YhCU5bsfuNPucbyuHUdbtyPjhGgeYzCzvCDuLZf9R0TZGrSlbmU9yWlklQb
r/KMGaEai/kG6Sb4vJx2DlQEEGy4Zb2/5pcgoelz6QF8AkbOlCh7dMrajQYc6juV8yZbbCQAzv/1
kx4a/zEj6l+8iCSci033PIHz6JjnQ0JAwgp167Lcb6RE2QrRgLGvxUYTOgJ58zPih5EQs0bljXb5
8mgyVhNdt9VWwmclBLLHOs2bV0Fx6prYc4yCb5LZ30VTDCYa73k5EEIVedQX3rbBh0wXp7ktUKm/
bAtNFFrKvDdCHFbVANB75PXgnIqEhIWON1LHNQoNI4tC9Vz5NTtoUkRQSkHTupZFBEg8VOuuP41f
pgPhNxJ5ojT9i2aYFQ/mWRXqHcOUIi4euLnVuAP+z+H0nYTnlzt9mJxDejL0vcaDSPJVGDqnbMyZ
pgY/KS3TxTd5HSPAgQXfCLb/psViy1W+kEKuI+PviCeULhGzSpzwg4KPwm5+Ppj+pRMaiOwbF3wU
EGt4Jcuhqssi0qk0Hcm8BslCpaC5Rp/szfjxmqrayZQVNIO7XlNbx5kts2UT8o0oP30+uOoL0aoH
9HTS05ootu9hd6bnexeNg/RAB3qgyZuTAa61+Vgf2TsnVJKeCsVP0mTZKlvMI/v0gKmWgv4yfTTI
gkaOUW/EqmIpdg4Jy54wBZi+Qnj9X5r9hMzyrgT0BRijJIrLl2LJFIXelaqr+T9ojYW1U5VRRgOo
+TwJqHLe3lk4RY06wlygSye/pgTTCX4u5O0qGr9Bbzf1eyTgc6ujgqiy7rSoBiZNbum/fP5cIVWD
SKhPXtyhvAMsDgIldhJ9L5kF8Yp/R/p5HFzFSoSE3ALYMTez2Zq10ElY9Vgi7A4r40EXUsiEQzPz
w0rdOQCHsKUIxKYn6sLZfPkv2FLlDqkQoIm6SRkwWp/IeRGhBmTtjXyDIGvRIdeE+bGfKOkpAfh4
3IUMD0MtE00NR8qQK3HcYgHetyQqxSPnjj5il9IMax5+6kP6kBd6Br3hIT8WUf/IGcpAWgg7A3Ch
mhbOcKd5vuq4I0y+0OjaPta1HR8ROp1JPGAF5VDFJgnoGCmb2KFg0s9iwaU0XeG/ZMk6Tmvjix28
jGlKgur7kmOV12erGkvbFInhPXX3B0Ql7DDDRv37W5tlRgwJLElW2Wu0Qu3GXmT+xRPn0xtoIADL
4luPsI+xbL96bOZe6XeZgJyWj/drusuzgteWoJgFWUnKcruBZleg07ZsxwG8Gk+cmMWO7SpBNfno
gqFwopDCdh8Sv3IzC9P+ZdeyE8kqhDNFn9PsUjoaY5DOJDJkg/82DHYCR8IKvYArxjqumKvTdAjA
+mGNc53SiCpccJ5dhfcW2zzRD0GM6JIQt+CWzG7ZReFPP093n8Mt75DkyIhSmB1bEa6AcR66mBOP
zgrAu2WsJ6wYgWeDlH2src6jW+VTLjMFoG2Uf6wanvhhl097YGABUDbV7JzWLmKQbwyAJIu9qoQ0
oDOVZ+XidlKBOqgVqlsS9e1FqctNf2TO8tzlz9vInzSdbx+54Wn+l5UzwtlW+7lvXE2eSdAlj1xC
9uYhwxdkX4sdRNOQ8wCsSzQ3+22wWd/mhpsV2Ot3PjRypfSI2CPl9Se/hZ3uDNfH/wdfqi4YkVbm
fonT9xzGb9iQb+7xbpD37gdmv6zfAk3YIOxkbNVHPc1MeJpVvO4G/pUpuAhQ4STXRwD2MJaJMhM+
KJNnz6UNdYPRsTsoiRLarW/zqwrwQMWbUgQX0UIyYU/j00Gc9svLX8zGqH3t1xSLRHFe0vZtKrVf
+2PzzUUN3aWLtGq95ZHgU2kkA2MUclEDH6E794hskdSOO0Zi2nTjqnIF+RMgXOBti+ku1CWRXH0F
WIZIDqqAkXL7+Ff6e8eGmUmW0NCLV0/2ZMeo05oz8IpVXWX6PqJONd7lrxwU9eftOLpcONbuTRy1
YbZq52jdir7gH9Iy7eJhiqiapSG28fEsMqyFluYwOj70gtopxNlXZ/QkwfA/Msuz0yPgetdp+cLT
OQ1xS3cEClB8Ude2xR27Gffc3t1xB+m8Bq2WGUkHlypX9l6gZQ0BHH5HGL93K2N2qiHrA2Ri3U+L
wHhMpc8JD7BHXmjJyB49nNPlKOTk7es6OUOQnRHbeyqyoKM/cynhHZf9P2fR77nk7rNAqdVRyrTA
UaMFwIbUN/BjALaFGi0RAe2iEyWrbReiXE3sLEELiwz+PrPTfUnp55Gsm690zGpuc6nhsgX4XQHX
2/eKg1XmVgprImos2wVhXxpK0MWhvBcKXM/4wfrDn0yk0Q8YobO6Ack8PKnfGmHPfLiIKbskpbIT
QcY6Aq3Z/HNhCGiKFwaWPZF8nKiPhawTdDAge8MWzXeCRdt8puEe7BxFaHm32QpJ0Qxb0htO/aJ0
gaXqKX5FzF4OiWh5g+R1ChEvnBUnOR2S5apkzW+KUHtLv7CnLUbAnHI9VsuqiY0v8LDpkzcnBKiY
MSxh271/gCIHMZS2EAevXdA3q3UrjrqX8U+9x6Akwv/wWBRbpYIlnPZyAd3Q5r183wioEtiWyNda
jBdD5+Tcaa8NxlkhbUy7zQS4keFQhHIODjV3ltK3cbm+0aHa/J2xo9FEetXW1M27I7bYrODdbU8D
sN/b4A76nI5PHegv4DPp3Qttobh4Ha/Wve8X+l3iYjQrC5P2ST/6lJlCFf99eBVf4ZCRg3amNnCS
kRoFnvyR6KsTP2Ufj80LZPlE5aC1BXSvPdkwdgJ7JYGb+PcbCcHSyXymFIFMbNkrlXEzHsBxXpon
KQU3yd1GWY6tA3enpdN4mI42d5qhdTXjwjwl3zr9lfJIJhx5AMfChc2+r9fdvqKCdU7keWGW1Bl0
1UE7sPHxKd/3jkVX75LwdVwR3ArE3l4k8Y1QumVi3V82fK6Ub8Nmf+LWBvIg95jx0EHxoj+2CKqd
qbU9j6AVfODovUR5ANCWKsKR5YIzzspJbPB5mFyXCf2xvNYd2yPyDJQPzoEgBn9ZWDaXYk/STjs+
ZPnhsWL8uNKad5AmSsMlTsctxQWb4tlj4GI7YLIhXEeVXjGXwbcZvBSjXKxpd0w9dWI00z0jvqsZ
pyGgQeCGleCQKagdpUekw4W0OHHVuI+qmckfQGaW2yJKYlYnDZqlhcts+fQIsR753ziD5WP2+9C6
FzZuzvzJd8GgsUO4IB2kiIjNM0v5v1IfVYd/E83ppBeWx4WcqK44/5NsEG96yr7BkB3cusa1e583
D7ZmiSJFoIcC1iXbiamjj0tF1yzSngUS+EWifannUhxX7gy6kAYE8bi5jtYtRgcIbZ8mD7TUEy07
2MbFbvmHfH+8kyPTmvl4B7im/VwdGryljRsBBcvLLwntGzCP+stFPpohvPne8QlGnjajWKn3+dUr
Y90ayxuvS/RaLskRelnsKI8PTTPcCm7LHbR8RqCuZbL09U10yXdFfLSEds9Jh/fF4p8emslQTZF2
YJ9R/vFfxzr08MTVRRBpdBthAJncWfamsjnhcnHlDGcyOH+K1oYrctgxxipENvGSncsGSjN1IAqo
WBV7h3yLS8+8kGP8os18DcRaKpUXlWtm9SQfxuhnTnYp9PXHLAXjGhToonhFC34hoppo3kPB0orG
AZ5m33NMyObaejCKEyf0E380XI1Fp94nPGWdyrmzW70ujm5tvpfEVPM3ELYRdo7LUUAzdkp4AwEy
kwQ35e6pnQ3wGqpO7HqfwG+AIbshGZ8Jfg2sOqpDVE32cRPiZPrVTfVtHrQZzEEEPdKoZc0BeJi8
096JmtakcdaWJ+26CHLE36zy+FZeONqVOllzB4n7vIesN3cxnrYWkvf8qPYc7SAcwVNzk3//3HjK
Hk8Z2GkjgaeMyXD9nCHdqKgNas4dgb9+fS3d+/UJWXeKGaKuYB21jWoNbLJzYIReX00pLl+dQUvG
GyjsMQMOb3qePMNRDeeGclQY8TFvAsa8Ps8THAsZg8edYw/r64/FlmJZLvKZZyiCx+HBnR+bfyzB
0EH54j+D65OqxJB2eY+lKCLFAlEacHkJh9qXPcUhr7NWfqJ6OVjDVEpRPY3GYLWvAGlSrlnJxNQO
U1zjqGXZIvjxVHlb71QBzb64PulLHENW5BsZhoLGju/qYgQbDH7Tcjv18RaNxDh3j1ZfmzqoLARR
7wgPEDR1K2tQqRSPDud4KE8R5MZibILogoRSx1gTcdhnP5ZyoZrDY/z/lK/+hzm+5R1BnbgNuN+2
y3BZZEAB3m3ZyXcoMvGu5xoVAti21bvY5vTO17LMtMbySxOn66T1WIZ9s44U8QGVreww9HMDakRH
iUF5HqRHAOZfzRvmkwH3LBr2Pftxd2y6GPCP20MLhbTtGTYQ0as0cQejNEEqNDHJSQAQPJz+iTX2
WntLe9SOv2xPyTDCCrKxvQKZVyVC9DEd93edtTmTPh7aiRHp7XQXa1WtAn+S6lde/ASCxYEbMKPR
DS887y1DXfDVh7EKi34EVH2RgL0HxpEp1gHB+5pb7hrI+kcGnRUeCxczPmqvZOtAoxRotB52ry9s
Z/ZeUwDWr/q1M5Zsc5hpRVHTKLkoJWu9R79mvDIuRgSZ2OiAMEn96ME3MN7v5f8v0KEQsKcvtEHP
eQhum9YFSNPooExWSq12pLI2INgOfDUJCdgyIZKHFiRudtOd6bCJeu4NgWYvzMzNcI5Eg8VHOBKz
Bb9iTRfc/mvgyjCLTGqBfW3pv4LAZFrZrLvxPoziI0JUEZvvJzkjyhyKRMEUTnh8XUnoPtIPG1ZG
NiP8Gf6bavDU/PdMDP40uP37ceIoumGqWTeKOh1kZakKKMe3tbPyCdH6DNLNyYDwBbdAZCh4DfKR
dGG4OQx3BRqe/fJhi6wYBrhbTK2QHJpAU+ChnRzEF+XM1R6s4IHRHnWENpR6SjKi9c2tLKkI0Ldf
jxoRJdPFzQFkjtDv7Y6aVpQ8l3e2BS32M4BZrPCUP6TlzBuhCzCgaZzka0qyq2Z9ePxP+ztR+gvd
SvBlYJavxLDawxEbiXZA0uQ1REqbgnFUiT6131Smr2Bsmm5W4Fpcud4OtzUB9O5zLIVHbjXfB1N/
+6tdJYJ07RDJrND/1IEE1tQsIQPcuqq8V+vmwBW+nPze5Kkvj1ZIfBYho769TmulJ3MUHkizSEO8
m0ntPmvS1krnO/I2jirL5TgYFuQTgmK3x3xipXkQXbpsYR14l81QFl++P2JibGBs/4QoSBTgk0Mr
5rhusIJS5v8bQvXM/hkXVuw8ou2zre86ZaYrAWrd7EkBLslJEC8i5HT53WXS3FVdz41qPWLlXrgk
l0w4cwPFaYkVZmOVqLddSFEu5jhQFqxvnuL+wDvNA1b+1pJpvNXWnDaqpaHyltC3PWIozSe2xODE
znvjbYWvKdFB5LFxnB8bJamKXtyVczirW2YJ/YtS4PBIj21WiXf5dwWKdQgB04IITHjwQUaRoJJy
yRNOhG9hoBB6QJdr5MUQ6eRoBeFFGQz88Cr9WaQar3e72XFrWwAmIF0k+lluREE9xtR9WZNMbIEj
+Vk/kFqKlahwmyVbO/G3MuRB44aO537HZysIMbTWCIDi4aEyCGhGFwkEv6nK8q3GoHhkxUdkkgYE
SYzrhAtTBGM7ZJIWnyJLmB6UankyU0Z+ajBQ6K1oDpzcrlgxmjxOBsiRNkESkYHL2/sKogrKgBZe
gpEq8zHsVYB93m2MGTTYHSpwpN+G2KMVmx1YFg4TbpKKML6uqX2lwcBYm5n7ZVDvcJqJMAzM27ae
mmPOSQw9KDQbPI6N1CjhF4VT42fnot4068d/3GQG2f2/XJqI//Ht0llFMHv3NSTxAdOVon5DaT0N
eSviNieKq++er6Af1dLkIWe2GpgYJb+7tx/xIXSxFWsMt7YcvECGKJIN2fJ/WE+k8jbAtTY6aHIX
NOow1k/WEpPPSR4C+owISIH/EQJoD3qI+ciDKCvouE2erouGYnyhOaAHpppTPkjFzKYUvN7Xc12X
GGCJzFfG6LcpjItb3t3py0R7V35sjjx4p1XaSrBbr0nAQsXk+dtCqEy35jf6Jcf50K4Hyp+pWW4P
QzJOc8jqjXg7u4vYaScHqm6oILItsT8bBzCoMFKNrvI2wdABj/19WIQZjo8GHNjBEBVFOhvjf/ki
+uwblq7R/RwVP0WXPqByaIATyt6bcareYRgcjl0qFEHn0H6ih1DsrGuH8bq11IkjVMhZyP1oeai2
BXp2c63QlR2PNSF9XEDEPtS0EOruF5SOFIB+jWC5MutMITae9naAaHaetPLrOU+fJkJR8RLqJ2lW
fLanhRvd8kgmqoJIh8W1JSyVCKj55PrpC3IjoAggLO1M11+j3pySQXwN7RCXGxnGf2EPZx/ntBmD
lcTcghk8Gm/R3XpOJYUcTx47f+o8Ewxyd4fU1+u2atS369DZ/oFcu6BXZ3+R3WUmjR4e9HE9nHL/
t+9v7kYHvzCpRGeEvz30GfBoxXj1TfPqpfW0G9teBqcx522WqSYv7Cv2CQGwiu5mX1c5Jw1QM3sc
eVAr3CH43kmAmqJsOYRbri38rqZpiqvDfzksMYqrcfc70UKYETGS/d9JPon80S4FZYWSsfkqcXI2
vUvoBhvMsAOqhmYItbfrAqwP7+AraQh+a1o3GncRWdjpGHfJQZeGxsY+szL76PBQ8pQTWWR7nZIU
Nr9Ko6lgpEyDD3l7w9bOuFZz4hQ1/dDvQx/HXIxXpPVzdMSowmPMLpkVf0GAJWVrbjy5ehpaQURM
JSIDNm2S10mLEPecTYFWj/FSY9c2+B4ffo+cDnxpbbdNYO7rmJVuGezWym+52hq6Ab7gNWghgQ9g
H+EASiBp07NKDPj9e4iQ6zAHlwsGy4YxYv/p1uJR0uxty4C9/zXrkYKR1ONAApMgDdcxfldz1/Yp
GbjDZe2Pg9tX8RzeWiujd4+5UTubLVnUYN1VrguLG89QhqphMvIDU30Cxo5gSaTOk40+Sr2n4w2C
v9Mk2JrGyVmZVsq6Pytde76nl+e7M0XlEroaIfOiEswlUPqbfWBgFslaH1CZWy5L5CMsrFCRlfL/
HeIsrFAJt0R8GcAuvWh+EdzY/6fnK4Ap7wZp11KZl908Yd26C5kNTz0i9KNwLSovzHE9bnpP5TrL
PMv2FgDYdRYPpM56+Y8jLygoTgvCp/tHvZBjx25gFOBYlN+HW0BrafBhbcWX2xWfX1qDenY24Sju
KTqxDgR8RfckNWMz2vgkUZh9V0CkHFZmQS/762kVXiNaMdsO1TbzPueRRF2hDV3J1B5bQq+wHk2Z
1gFpp318PV0DX90JMnN1+xPIcYwcFdg9vdbEcrqd6rMI7CoaSNOy078VwxRz1h43FXyeIK5xzacD
AD0JfHncvb0NCsAhvn0a5nj54mXhAXutsQd36MpuCi61C/xQGLJ7UKkoX197x3v6wQQ9No8EgHhD
J5QW2Zb6DjMIM1Y1yo0p3JN92AVW0VMaW6HtqlJRF+9GSxMW+MhSt2VU6uCVUhRg7ljPDIROmf6r
qbHeGgASeJDD4SufIOfgdrr73l97XHFSQLh7KBmVIRVT1Ms7KPWoDGlRrdpmIPshx5rqpMw9zZPk
fDBXxsVzu2esepUpqTDh6jy7h5uMdJGE2CJ191jtuNY9XG3ft6ssADiFuBmvmJeqSOkBhFuVgtKQ
2XugJ+fEhxp3zq936JL5sJwHY0YK3mHa5SGggzbmxUlNBNMZSOjCHtdgcTryE9TF5ATgv231aisc
k+wltbcRxNU6Fnm54DE+7dr9at9ocs3l1CXFpyE6WAgw0fKQ4+iku1R3gJm7+rwsB7BtcsmND7mV
FZPwwpSFmwUJ/HgASqTJNLZnSbk5l5IMTQ5vU6vbaEt9/p2N+VJKWsnO61V0/uKhz27fG4yORQBF
cFRZnqWDadDZWU6QgY4o1Jaq/vwmtIhhDsq8dWsjz+AZOQHzg9wwItQJVp9dK3BUp5HC00BKT3iv
Zv3kNJUoeSj4MGZvCgOn93hK6dloSct3VLuOqHVgWj3TqCwsLMqGrYLT0aOw+McasI+IGNRkPOc+
JgBiihDixlusJq7FVMfectWvjJXcbopicGQE0KgZ4Hdr4FhDF5I3OfbMa7mPSfwGS7/dxbTDjbDg
dHUPnpJT8Y18f2HRF/JG6vqfz4uQufMtlyBmOmz8dEWHQl2BffluKTcU63D1DaqKMUIFrI+5/0tT
AC+0oX4ZBJKGyUN5E4c2XJIPUVTBbWUgxbuafAoW48nznKSj4SnDsv3habvpsdlCeW1QK4njKt+O
C8qfmaa8NLmcH09Q17lr6HIMAkINWasU8xIrOtR6c6zTDqqTYtH2WtFpTyAZtm7520h/2Xufqfpk
yluDhqKYhduYfiPPDrMdNzCZ7kycPmfG6msd8Hfh0R7vLm9l5j7uSmCOPC5liFT398v9f1iw3hGV
3bv1U8t2UF8bxzn9eWxg3kf1f404dgVgy45WOrNsk88ZVy+Uy7h3NrTv8PEw3PYbWiPHzxKH+KcB
vhcR84Pyd712qbEht8GECloqxlFHXFPNU/57D6Z9L2x5aMLZ2SA5DfpDzInRn423zuLpB04QWivC
EtX5PUYsXibxyeMnvsabOhAP8ejUnGoqU4fZUf5XU33tHDPiz5RufICJY81OWjXyGngdOmr9QXCL
Uxx1myjqSuAQHyFu8cUhdGzRRi62YJmplEb8+AxfPQ31vV2ODVP9ih29n6vmQy4TSumRCsVWPUgE
cRTb8T4nbekw5mcCz0OOWEpWfm216OZIz3hBXSS0LRnlZ8BwyrS9aUIssI2VB4kwyjM9VGvaGeZ8
V2wPbtbgJ+FiVC5WS9l97tlwUBWClnku0CyM2PD4DA45ABpaqGbcmWmlEhwh7Ql86R3+vHe2xYok
BoxqMPrGttPX2zQDUfwYQmNFsWYQ4G+Zc5DPe7XRBBhR7fEe7lv1DfVmGuhbVa3cOkBzfGQ2BR4Z
Ybgt2kVm5Sl6oTPF9fR1grqdBZiB3ipYgZH6R8o9/xw2LLM9fLYcrowZ3exnrOs1P4egPi+R6xbj
6UiyYYDkK+UvbpIEqAQqX+Xl8ElyeOHa70ozv0sEANKDuIW2BGCDwRB6LvXS2dVEV5vme+zSGU06
EcR2zXFqMatp+STXdNnMiL/bU8NkRRy/N241l58XXnVYlw6qZZdptdJarfgnC4bqi8Kk0RggB8N2
TraRnTs+a/AHv9YxVwrLSYP3VIvOkJwsm/H028JMTrXZ0ikIA7FzURIqVOQadJywJkk0edfLMaDg
hl8evucvohA9zhN7kIV9R5PIOOmZHI9ZRiXOIHxsabmZfqY6jSn5S+z6k4nJOXgLLcL6A4BJxSYx
dkR7ixfKkmciml94oLAwaxOIXTvmKhJbRtYw0InZ/YkPOyUeZCmHJiBz7RwfxZGeXuY2OoJs4+f2
Kt3LgVPiQ1OcCW6l7XyPSyE6IqSQqYGRxG/1SC5EbJoWLEoyMPGulYr8eY5oePBCLripXx4fN/RA
u8wEtHS3RLcF7eFgcwiWugqLxhTZ82G115MGEmpIxE8H0zcVt8b8Tr5+IL4BKIfIUvMt3zt67i0Q
UJpS5W31I/2pgqdLFbP3qj+Dz9sJJKPSrWWh1ynYoFptJvWizhb8f/O6NEzMrciyJCV53IIKqOkR
mrO2RYHokE7C3gtkyy3ULcalr2+7tH4M5SvLIBIgZLonKdtPPjtsFTlY70c+eyHM/kDM/2u33Hcg
clNzpzAyonCuKHk1DSEU43Sz9SmvWcfTecjyTxuW8aeVxJIxe+xbIp61bugBmlUJtZJ7dPNW9cdk
eGKKOW5JynOS2PdOIHveryR7HKDN1PNidpRE7kPSI3SwlVg4Ye5fbQExyh30eRxdrBcS2vQU9cVt
EMcKI9X8gk37Qaz8513z4gv3QVG5/sBjHTFe2pWVUM2CEtNJ91sPdcTGUGRXTeRPTkD+KirTalJG
Bf0e/57Ni6s291vMLCpc4E8TsCz1rJRnMJzPQ95GA1IiVSdAJzR19eGe7fgo4yeaqbChTCn01OME
4SG3r5Hba2gfGKvHsggLendiIRffG7kndOG+zG+qtoqkFKjR6YVXvdeh97pZbTH5L7pNYRn6wMYp
AZ0K/4WrjHocpmz4MlrDip/7iSu1/cl1qjcizb93BrEZoIGAlY5x6SHqb1M8VVwkTLU67JlJLc4j
gSVjmWTRYHxXzY7R5+u4FB7P6Omq3TADyEIvvilBZCkdp0bXxUCi3ho9e90dmU1psVPrUcLJpZKc
i1tQSf3I/wsEbPgPVwgwooxzhXeqipAwvhG9V6/XyfXPlHdK139GIgV7NWaaOAWUPOPKlK5u3EYS
Ys0SXlOHzWUZP5IGrGNvwzlilWNNfnfl/Jz4HyiPaC1YaInFiI1jvhyPN+bS6r9vDYPQRMk9Vfjs
TmqerITmeTfvXScTJD1YZq9pw+zCR7OMQZWJ0sEs6zB+3MyKFQn0fy4q3BM8yLbYYInXJgJsPYgH
fh+b3JT+D3ERllGJ30Hh4B4cZtMh5uIST7PaY1YaBpF9OcBDmKmV/bih0LGEA9OPy5QIybT29eW+
U7DraMl5jg0k76akyggUk8LOeS8PJ3snTYtw0prVe8ipmUbV3bNPl4fSMfwhD6SuRQS2soioEgO+
k9qabe/y4vF6N2qhkYkP4meI/vaFODv4ufFm9DkbNP8lR3n40nncy+sx6GjFbihsIzPWewbvWK1B
fm8PHUFzcW++/wcu0JxcnoI8EfNSr5oufLMIy54Ggj54HoIC4+WZr7gDt6y2XCyZXmh3go4Lxqv4
jy9D+Rgx0ab+iGb7gGzltIlONeA+4u5k6yN9rKJMh7nGX2dRXn5g2fMG0HDL1uz+1iuiXZ6C9Vh+
JslJtv5+5oNJhncRr1IBdKHgRrjY8GqL1/gm01CU5odEfK1Lyyg+68NgJtPaaI4UOAvX2SaOYbh4
DHfoG5Cbsu7YM2kP294PPZ4gtQMi+Gg0dCh8Jty0gD5BicGd/oYk11hSRZz+Q99F1kO/KhcuIZJ/
IBM8x4BvWjVyOlW2FWUzCZfxTQg2nwxxcv1g0ySD51zherpZaZL4TdkZsvdkNUplEbnva6nAbs9T
KFZslZNPJgpA1kzwlmVH8j/qTahVXSbq9wkM52vMiQPKdbVahfLihfWxEbSa0HuiKtTlrzUkxOLQ
AddIW/xGbv3bwFD53fsGK+qiYbzzVB888FxX/nPROmCWNqrbCWpVv8FZagZzg5n2oidonlGgF7I/
alxPKbJrlbPa83kL9/t97Rh1xNbZx1rdkqfqDTu6HC4c+Sk+p/WkS5A+m2PYRUOGYmD1CO39y3gt
FMBwowmbI5IWLsfMznw6VPmwxZCJ4DEplBUIdu6OYMY3d8YS37yMB8tUtxRP7twES+aLu6V7HVuY
cXNHb+kYhqiVt9P7peR5Bbo9j5rkgZrMtlEa5dUdYWYe8U6tii69kxnukpPbnWHZf0XI3oeUtBE5
Dv1/LGDn21jDCzqrkOKpT2UZVXHfekFIYOIQNtOgfKQM/N3qJ0pGy7FXF7w0TQP3R5JADmRKlWQ/
0bs6dHYKOOhvUzVc1OwVq/dAxtWVn7hTP98v91RE00gsqbAOmE7fHukxnGvY457yzu5mdtzEsmMS
qXS3pMsHATkwfSyfszcldfNtRTyKpfnhSzHjRtUoQp+JIackC3g9oFU52HpevkUerDd9JPP16vXD
IF+O3MDVCuDvPdJsEIAPn6sZDZgLpgDyE8SlGLXon8Ksdx+Bso/1VzLeBOr4scmenufnw7k3aGxM
+v1DsnYJ9LPh6T/n7rUuQNZ2QZWN4u9YvNQ5KfY67ZYBL4c7HFcqFkALQjr1QaDhBaeumjVi9ne9
4muT2zGKbsasTbVpaEcUOmrVKy8LKrTjhbi8JMCOAJBBAD/LuaZeLox0UMuJW6UDcThzF2iTY/nr
e/xHpTGrjmk+hUQ6I1exC4lTgI5fiMzbb03UWlWO6/MaRfebv1nT8vOGil6oOiFeIUyGSdbE/bKl
eYeMSkTAXnQYyF6v1MaiCi4qORnHLJHFOhRz/K4MXBucixTbMWU2VpAknRM0yHEnaLanhRo3gd01
i8kjFqqpTEhlBrah7WaY+IbXXgpJG0s3q05lv9hBkLX8yGs7OBC6JjWmpDEd/N+3myaj9IPswSLM
y9UZaj9d+yb3MS5ejlTwYqflVe6EgOagQtRybYV9c4cLwcfkviYVZAq5Q++T1vMNoM10bE4EPE4w
9EDrnBNrJ1dYZEb4IN3IlAjBOJRg9S8LTtU2RrFU5/BYnQpvejfyMDRt0TDvnGr96PVvYhxU5y8K
2oHYU0CQlX3a56WHBXxIJUi1lJJYDcnSNBQrbQO013a9VX7c8NfO+41sr3tTv4anzPKtfPQvY9FP
XppEpImPN48anZ3YXYHfRcl4brSXZT9Hj54tdXxXJxiPWcd9HKZRbIReEkZ7VuAB9u0yercHdWqe
V5xnp0hGKcAe3R+enJqoBRK8bB0Q5y+uE44C5HaiSL2HQtuy9etCb51qdjZArTn6cjdAbgq10gsU
Twkh8a9/OQw24x2g7O9WXBXPiGfFd+9xRA+5KrlCb/L4mu/wmp7VW3ZgDsrdNFDlEv9sQfjPajkn
H2lsi7hErJgxRSZn1OXu+n8sTORoknsCVFOgXJIYkg2OSkJUltGaNOpu5C+r1a3SGvd/sU2p5Tp1
1BJ2i3fJRDKW0mTaPuwuHiZE9hbAcrU0bfQl1nLYqvZ4WDzIPYibOA7DvM2kAvaQJLvYbZSzW6wj
R4ssZRDWtu1fN/TQ/qnVPkEBrSdcgNI8yeTnHEs1pIa8IuQmgRRP4aoEreMmSTg1yYka8x5TE+LZ
q+Z6JBW10eIzQuyrfSHA1dg8XyDbvaNNaCdb5EyYcoy9oHIOfGgs5uCyrvTDDHhV3gDu618YeCrM
FB1Nb6v+XQLBLUzyT9abQfC39WtubLaAecTj0wbl+gmrPM21YXzOP2Ah3ckqnwynp4uUFYr+EbKK
+43ZPhiVZStMxENA+zf6gR1mcoYjNahLWXIDabb+C+B518NHCosym8ORolo+zyvAhkjx96OLlnxZ
9CilGftZCdBpEenTGWGgj5MXJ+ZL0d2WlwA6QLnTfmOTtQAJi7I98p4HRHfgrf74JCWFXhgEW/u/
ImCxo9Yp4PIbqE/x7rNyPQtkZknZki35uUyAOfRxc1HLNG5kvUEPvtKfdL9XxB9Iq0iFU2Vj1jBr
Om0mRjxhTB2xklLpM7keqrSTHMe8nYA1Ucwy/ER5Qo39GWQ34UcC/ehFkb4CKQc1OdsVyTzkA4F8
jYXBKxLMiLZnr2rOkNeTjK0BvASUUlqCKY6zree715YasLl9gD6qCu3jpwsl5ty/FPTvTF2sFS2B
qVv+jHgEw4CeKdprr8rsc7aFTQWNWnfXioBVtnX+bdSvUn3E9QPO0wMHwhU7NNcqeGPX5d/p+sBF
4B0JGPyIFTBrHbioLTKzZwuLvySh9IbKw+G7aY6Ywie5WD2k6iKYfjcSl8KDkWsg/8opzHlD8aiJ
T74ZRS5L7W+OY3nxvtvOhO9G6rTnr222GQ5LqLGXFjXXRXahFRsGY0t2scWx/gCHhgGUxju7IT+O
hl+A7dsTeN4ONWt5cT0UOSNfz9s3pAYM6kV3mJKbY88xViiFy1FVNInA9g4S8pBtc+uLPxN5frPk
0Ws/cnCvOr+gC+qGw8ZF2ppiSGMilxe8H/vqhyVfcsK0ln6TjD6pbjwmr76hvYEFJOepsQCbCJXZ
hzUMbPIVEUX9jrqDy172rrH1A5aQzhZIRcZBE09EBobrIyr23w0dKyftNH/Nd4nHDTFisbAPQeBG
zn+EBS6McwukLN+plPBvJsTwKjqmDTi3nQd42XrcDLeH+qY6Nrl/RRVY2/SnrXJVZpxms5eJXNtY
oZZb5szS/bmLeaNEPAkE7QyWN081uuCHn/ajpv1c6+gcd2kVerB7iqgx8J/xfbtISafcfYBgqAYs
EXKxwBZls4NUh85RoTCFbquZfLDUV5j3PtDnGrS78eXigcFa7Jfw3qfIgA6R+obeJE6u87Jb0yto
EaqfXnZJXLOUduYmpxB0utc13qr6tDeev7Ewv1NUTt8UcNnpOvBRYXzX/KcadBR63PrkwMvzQzGK
w3H0hYrgKK7+HQtJU8exNdEy+UBfxpcZuhqbiPRGp1VEWRfYH8Hnr8nAUeCcg6I5Lr2al2FWe+Nc
WnNVXpfEZN6p/Esh85ASi2ojbcO5xZC/1crGqLlZIvwJig92ZxJChZkCTm4U07NWaDpCtpje/tWq
WEFjH0grD9MBsHSAhraEBR9L0RNxGhedkaiku+aObE2RFey97qG1GczmeCIlbGRkOS1yRXtQ7sz8
D6URZGCEWXSE/oa2ifqLZJ4GLX/ryFU5KJDjlRLVkQj8aTMpai55/LZwQUakDcm1BmhJEbCIS0R4
zJRYj4ADoB5xy9PDweuiCqbYDb5NYjGmWKK5x9n1v0fc3FCaWhFVG+g+zOfYOJsROPpk+uCtAsBH
9gDvxK+d7S0fiL8TdMBwqhDSRhYqP+gjCMWrFpIXHoX261YscKiCgCZmXfmFuc6mDGV6zWPwAmzv
MD99H+Q9hzD5hdemkyeJ/kC36zwLfvEvsDrTUVL94uMp7E0RNLM2MEQtW7pQBuRVcKWg00Tsrj+5
yneO2HmJ4hg1JlV1JTTkUaqswLVS903QPIpsM7ysvY0THNJJWZAfAEOgY5qJjU6deOoKhSsL0xoF
tRebw8dlnTinu2LBEbF6B0G0hXnblT6/GRGWUPV54qvYY+oa2eYTfXDMaP0/scqovhXyyVkU8cyb
2hlnpxrS0z74g03zJHSOmeLMoBzmGFM7ezS+D4hQPfRQFJjEKhe+mQCEMvx18qCYxMKEB28WDjyt
8nBdo6fNc/vuyD6C6yzNhIEg45pYNAhSvxRhr9Gto/sSDjp0V8sAu+raAzTLxTjwJmACExlqfGfL
PhecbB3ql2/ifZL5uQAqcAHflz5czSlI38bvLDRr/e7zDZtHvhqkrM1Y+BE97gr1+5YshzRqUi1+
9eeyCrFrQohFjaA1O0ZQwPxYHGEz74YvbsXW1L6tdWUagObhRMAtWCuKLsmH+lgRJH5N6xM9kZln
tPcLlPbsuMHD8EC52nsNCu4k5hk+f7QE/VhGvd8vi+isKG0lUxXlcbNk3uj3/fuFHwkphMnXs5wo
413Tt1oiIhdXoVWNLeHXVvtzc9IHidOYbqKqWDH86GTi1M9qXn7GU7c4LTI9lmpeMBSOKZZnyj4C
kp7DW0wOCOUfnscZWYHyb3988NVclfKarr7zILe+72LlhU5IMO3HJALuDpLegLQRydKFtd92Zr8N
tz/ihq5kEDscy88cjuZ1EX0YiXNl2cEYLHVfb+zla/+qrqpR51VbLKA3S7//60Btvmndcx1NvdnQ
mx1+kMaBhVxLl8YqqhLyIeVG1vOCe3kPKp01WVaiMtDdoLIWlQCKWhhnkuyKEJ6+IGEcN1wJC9zc
rPEa175eoays70QQxzbuJ9DikbwgH50xuk5f1rUNDh/ajqZGepz0I0NUBhcNXr5U33T6UW07Ixuc
nCqJR7T9MySB3Hv8sltGkHRgm9XJ9Dg7vvSa6IICp9qi7vN3c2XQ/YFFyfUEnLHwCq8pzptlhPcD
5v4H0APHZAJsib4/0sV5aZGI6dY/9FUGrqTj8n/Kaf9Li0FEYqrN0tj4cwljdFSuLivNFmu292+N
f9oDXTVuWraG7Ka5C67+pmjv6P23wXQ84d77jzidrnwGFEzgz0ODWUeIHcR5p916AMlfTBq1Edvf
/I1Jm0eXqjYzaw7Ijg/vOhh/ettLD3Zv8dhyB7oWhNgeRWxEzTy2QstffUcl3vSejy7Tj50poQ75
8kNIO9u75q8m7Gfvi3bzuEFlAWKjn2zVMlOwmlhqxO7oUbaWMWRgeIbH8u9KBnMlLVDKkxN2QM+O
2GPH/ZfJVoxX8SufeD0i3pStKxi09Z5JncO5BdXNx+UVOHU8XQdnFkWZByuA8yJhRZcGvx9KyQBo
OdFauh6rx4+oXxbDYE3Yt6GjuwjT3ozeJ4V4A2KKX/JXvc2+VTzhuGGn1aFEHcgtKx8v85D56b7i
ukh6lyBMPQhJ9qOn5sFdOHci+TSoASilc5ocunwkLxVY5Sb2wKY9GYQco5trvQSPiw1A+xfDXubT
yi3BcSVGCtEqYXIDr9dos7Sly44Ki2lqsntxNu3P1uUzO22ftu541lIOhkQ0wO248zYqAnLJQVi0
+wy/WCk2BpXJtUxzww6gUbLoY2EnhhMHO7fKrj0Bg/afVFFjWMWEG/A8nBbw4pbksfNmnts2FHHD
/LWwu76KUEyWSIKTGycv73UracNQSg3uf/PLGRZyL44wEj08IUfLc1/4LJDu7Eq0lZZsnKCn++pm
BvHkqtGihI1Qy/2msb8NaUgqgcr0CRi+RgviutKhBPjPQzdgeaEw4ozCdWYATql6Db2jIUT4wu40
HUWF7YsNpVRYCIYixMYxbbfbDscGXm502AzlRyxvcv4iNaMPEqzfUgDkSC7iw7ia48hLPkb9mSns
3yGe1yxBhMYr+O+1Dh2NLTqtroyw4IJK4LJ51ss9Zaiu0cA5Rq6z30zwLMvHxzP6Mnr45/gPaTmZ
9Aql+JCVc5yBrB0BEi1pvJ0bUMvqqOGPbhpAJbzj/4PciYcHn3b+XYeWQBVVQ2ZwEN4195CfHCQ1
GzkvUEPRsoqFlllkFZZj4l70kXJC3m+w7wZ8krup5w2hKHfKJ+EwtZuOxMunhjL9oF6Cc3g0wk7F
FJOCCNecSrO46AQKbdlC9kSADKpD5AfXDgGE1amwoIz8+TJXfBWCIDw5lzNyNPqq9/+veLH7Ucfa
hjjojOULyqR96cPTZLh34PdZB+HSrHhS+5rh0TNCHb2xMr44t5svy8YHAleDB0jgU6W+U2XvA5W0
MfEUOuaesfffP8zbZTetWWUyNZw4ErBvcf4au6s+nuN/+fQ0Z/eHGjlun9bJdz6nVtU9pzCVLMMO
K0xBUTlDC1OyyDzzi/jZ+H9BuB6XP3vusPz7/8UoWYNPerPdAb7hMHinp1KMbJ8NF+RZQfD8SvvH
5tZ8Kc0K4nqNhrXQf9e1bTmBbTP9oAjhsUWCzSL1qPfpzPehaktQF2rock+Q0k1dfrFOsRRlqbjP
K3I6jectAtVeLi3RaySs8VlmjM41XYQ/qJi7EvlBFBzQOSr/bRaO83pk3PnDdwxmUDzEpnxfSJjV
R9Dm6mG7KFE4fk61rRhLDnG4bGw9CmNl/3lyTTKl22RcgAUKG64F5DSmP9kxrelClkmExOFa1f8o
pVYmsZtyuOmGrN43MS/wAJHbcln3IepJ6+9s0dSdf4Z4xIaCez6djBrx/7Zys/4xyeFZVgnwYCPz
/T7+o1tzuTYhmjImm4WsOomYNiT39aJBt3XGkKlJ9zQqIc3D1zpHpWXCcaOqQM4YSJ2ijuvdlsK9
B4k3tZSUd6jgn6GQKl1XOELpOYRcmPs1Pf3RWUQ3QxaeoN1a6X/kRX1WAl3icSVqiufb9pl47HS3
2jKONuhcsC0+DBQdB4nOeasFpGKKSWv8l+9NHezSrAwAzzeyOG+zIZHfPeAevOHOIHwb21bKns01
QOlZh5BLEnVtAbLQu9RhyQn4LrGD54gj5CK39JXHjhMA2Jy1DIle4R8Gi6EiUcpLwQFl9NhqupsS
Ll2VjkVAsdmP5h7D9MByCbtGQ9oTGdbeJJNRpG/qyMiK+20upPBxCzrmf4n7QxTRaDqTMi3i1+dW
2vttmqEJ1hUJXtIXXY8SafoH2iT9RDLxyXAieCvzXSxFWsz8XD0faLRpoWCC2dJ1fLWj4R+LtIFg
ACauCSNxk3UMpEsa1KhFMV8YKcXuM5ri5dGDboC7vwJZmSd1BwwilpwQtQLRbU2LacCXztWLznWk
jr3w4TAh7WfgAiozvm8omlETpHydP4Qmd7Z9Hd44Jyh9yqkkcqf4UKa8wI5wabsUWWgiblOjLca4
pqm9r/cULMWnOaWrkPLLguysU81Ep6UTXY3qNPxReMpUyLmEWp2O9KsL10O1jBm5FfXhYkiR8AHb
DC91ehWio6ie5Ac82TLsGViAFaCt38GBAldSzfFotDu7G0jpa7y45wec0Oa4I6XupkWU6rN21a0G
tl8dS0GjzvZYv0cOcC4Vurx83YVNXmR5OY5/AYPkt7q/7DLZqR4smwO3ts3mcS80zp9Dz9kDUtFF
NOi4z8kKXZf6/Y+Fg8J1igKF2sLarSv07eO64d8ydEyJEFy5pOL6nK14CRK3xHJQnX9QCZwisEHZ
q00EqZk/OJcIVqVRKlUJ9B5P2nM3I9vZO9hHYuOPl+Qc9gTw3kxepwDBsyuPhm6BnISrnxtNZ9hI
etu+xYR8l0BVDsZ/QkLmDRQ7kxS/YCeCof/PmIczv/5DDS4aO83gfgJhg5vfZtTPKaj3U2gE4uCL
RPptQZ71X6ir7sx8U4R9PEQu2rjks1XLuph/Ieid6W+bX9R0orhEbmyyOYE71+RNlyBT23764sS5
ehrXLQHx1WbsC3PuhQLJ5sQAbU3UMcDamHBqNFda4sRKy1Dd+dgIn3xemx+jWQX0s626M1YlC5sC
+n1HidqciO/07XUuLC6Bc0TM0uZukeS/My8MST6n2NRWvN5aYkG1WyMmZskF82PHB9WTCZOxacNg
U+2FljrcspCaqReSj/ERzYz62dpDbTIJsFa6CcVsxbEN/REyRA92VvY4o0mZ2zOg0JMPROoMX812
/eSnFWVah1xxdQdqonBaluE5cjSXqx+b7PDGrQu+h79bHZAbA8HHaOilE5UO2RdzqHRqKpjJSbY3
yPWcvobv9DZtpLllNhCCuZ5a8qSHHwbfyQZzpqYatEzFbQze9fJEATF3K0+JHA0CO+CFPnUJ3BGv
2bAJ90w9Ph1YfePFI78cnZKF3CxDBF2br2h4QFcpG6rJp9rijkgPfu+3LSGuc4wEiA1VyRUgMuDS
YgX8SRZ2WRFoUlrKxkUE0WrgNLRRVOX4IgAPP+l4dv5/E65RgD2AUpxooSPZQ7OGazG5NZ1mUGjl
d5TQuQtpQfukUTzddppbjAr6jlSMsNouRUwUj5WQWcJsPAru0Dd4kByxQUqb+YJ/kA+ZxEFbL/11
2/FzoZeVZjixgSaMesoHBVmXq3JvGnmnBoI1SIkhmpX9GfQsfUIhpcZ4NiT+Uem9JpxmDy5gES4o
pxpBHJ4r2Qu0Ky8Lh2UerMIeBLk9lNmM4s+a9mf8Lb6N2OUkNnHMmzzdBR5yTV+0wYpJGwS/so8l
IW7kyiMLNm1IlhgT7ME5VZerE9+MVhPB5RuXq2IZbPFFYRAic/wDWdoNy7bzMYOlUHrb+ZmM7sOZ
5UKnwGg4QQuM8e3IXYSvsVZWRgV1nrBMTyKLwvkmpR3p2QhFKp09nft0rBAxDXJBdp/Jsp2e2hjJ
IjcPc5iYNsl7zx9LgUPXEe5hG3CHBPlgRJCE4HxYVOoY0reR4NkHDc5KyV2dpTObPRx4R3fZ1SwC
DsjL1jLV//FlrH3ji2Wz7jWzzFMEa945XgfV8ALKo9wKq6omfKOU1cpQ6G+H6lg7h9R0e/7yTHcP
oquUa2URK/JAaaijVSg3TLTzEKRMCyc55A5A0qAlCU0ki8DePDZ9U9Vp+8NxZeCpNWZIcddTEzFE
W3iY97UUeSpqppUbr9mHWb5BsrqUtFAv4pTfMp3/erIHA6ReBoDGNYjTQWI7rW/X5fINRVJbhKzH
9KXLRsKjSLzqJOvw8qLi88q4zJfBmYj5T93lCqDEX4rSO8uzFSXLvnjOlodNz4Xau3m94Or6FIsf
LV+BJj1Kxxh814SbKaZspX6knW+qbo5PZOApEnjzqD9OQ+tk6jqQZzakCIQsBuGGu5sTcohGLNUc
5bcHlqJL7sSwQMr2jsXJIqRgJp4P41nGmJxRGj9YjJQ9u+hv6OJ9/vCUOES//goPTObGlOFKkaKy
kGD8Ugb0VobRqk6WkljaySFMD/hVNuDPdxjR2aIttygK/2g19sSN+oQFqNiv6ke/wRM73Pa5VtvY
WrnG+0LVFeqVDfFSauqUIDbMNG1RupGsExaxNfW1N7aaxG3NinYyD/CQmVSzAxxZTsmve7sWfwQ4
ifKdngmJq6wpF8BOAlLxcllVeY5RDABO1sOkEyP1Kq/uiu6glka33WDknWX3L+i7XxwhyZwXmg28
Gg/zk9tkvmXPllpGrzwNY4lALdyL7j/wId1vEYldSrODvezjM/By5Gb148CkAGerOVZ03DLD2sGc
CkDTke7OxPN39o9e9pcbMT2mgXCJwFwRGzEv6b9AYETgkMwDfMzOdmFSpPTck2nIP3PeTg/9FB0K
ZM06RYchlkuYLyaoEGqKRv+1/Kfn8CZUZDCz1aXy2VcJMdkQidWtOA5kF+hAswGme6Vmum7WZXrD
KZXQYyqVDVK/ck4MZN2RfvPE5SLrhIkRhpLFd/8KHl9LpIMm1nS/XAH3T2zUcVscTluc6wQ2jRbt
cUxUjkis7LUG9Mpd5GXNCwTPNzFfrdf1SaiUKsmf5AFDNGJXVpwpEtXqodHMBDSXqLgKM7Pu1KDR
KoJCvKxQgywrAzNdKKn4VRpHFuZNT3jaNS96iiph6LLecU2rPTwEAEKZQtBFPmQCuIkPNNKzS2xq
8GvLSRRgeRN3BZ1aExmMNQc5rY/RGyBIHBDSTohq+aHXuuXCfpTnwKoA4DdD8KxRxez9+f4JS8KM
1D8uox1mIs/agjqHMw21p0Fu+dvt55s9sDDezIsUxPXEGTfE2jxcSwR+PZ6R8YOBY15EeO37io+f
F2ZqG0LcSZSvAen+9ZfU4chtdDsHXqvqOIhAGhQOKIHY2A7nTO7kzD5BqJH+Du3n6YtkH7dVAFLk
TY8py6OA9TZAKtOqcLQUbVNp/dSFih6TfFW/fZosQqrj4WQJMy5O4CqBb5h4BarafPzfDDXnGkjB
+VdJc2iL4F87+eKS0xbjRBEtn1UrBfrmnQDDoT4VFQuZZaXroHyXqAVCRnn2hor4/b57cuPLeA1L
Uweb2D54TW8jYXD6Z2FtVBZZHndbEI5A+TspUjk3u9PBeUIP66ON6+t4WTgtFmJ5+CpFq6Dzsaoa
pCNBfth2buJ9S/aVu9nRKizWTJfPPg5JrO4/fnqZQrbGq7v+nVxsujJEufJ1B19xcPXkgDG8o13p
EhZvg3vJH27hGjX3l3WDlcl//8euRc1kwRr+L4f7NL5f5gFf1BS+PNMlCg8AULkDqYCDzECWP49A
/CH1r5F0A3ENuw3ssCAPgPuAujAWK5Ze2ndusOXlP65dedeqZ2aM54ALiR5Nhl1ZnyCo0qOtXFFt
pL0uugUHFrzetVKCB7LPLK9HPZbNz3RqY85p9S9N1612yO/jOYJiZF0vMisjdEE6TEa/wV72LCqb
v/WB80dAeCut6cFMu9oEshnDaFIRqK3d4XySnKBqSD0K1SSOwAwva0NtitQZAgyR5dOnE6hrrNks
3tcwna6WZeZM3wjonXGH0OVfxmV+48+8LNUB6uPD4MTnUFBm8BGJQIZ3MnLydpgaRShjdzE+gudK
D0rWbBopsUCc6r3h82joFa9yCJeUyUpDA7X4vVn6yI9rlbYuHjyL/tUa4E9PqAn9q2+CtB9bkRRI
04jcKsO2ZnIzJ7Ggj2iSxBFcpwe7/0WwHFul0F6p3uYAwhgV2Lx0e/UKT3Gcdsm+/mCe3NibMBRJ
Pp8VeRCwmVtP8jrdbveHbjOUiyb4bJlNnc4YSaoZkwF5IZ5nNmrpoHXEGgS5w/+yqenI64TXWgtI
QkVcu0GqrKItL/LsMpT0fcJEfIykd3hiKXSMkMAbJuOkS3RBd2CbJbE3ogzpkPtVSBEvJ4IdtziV
/XAt/2Y98O8RUGXgygxv79k9+4hF5rsmY59Vmg75AOBIfO5ytZaH1wHqblJkCutxpXOQ53O7bdr+
cqw93fXRN7X1leIsq/LflKVlhSjIcutcTXQ2uVBbfyfw1107vNTGyw/PKpNAPJ6UQ2T3H9Tq1Y81
jeya+KJQDGrX/DOD9aLDgKgtVdFRV8adivAPoidAaX0WPKTUgjkhoB/f6zUU1eWGtB9dYWkN4ire
rpaUVIOAOQugHKcCluwsu2ZEzUQoxmOgksFllhWOe0LwtFR2eSkMjuoPHKaYrsfe/UmBEftKmOPW
QNOTebRK/j1J81Sl9Wnl8XiUZUIJeYdYOYxAFqxQ/sgHG+dRqKHQHX64x80EMC2MD9q4po4AUQBb
LiIOn/u73fbMVsT9DoqTaoGJwpZHlSsLypiWj1zohKS71lk/BXvgJeXNeAIVXpgtYE+UQxO1cW/0
/W9zYqcAKvOnaqwhPnEw8yio83Q7/0E3ZnVhvmvEDVaXBQJKa5QLdbjlHHVxGIiEOvmSFgrZ5ns1
Og4Bid2Xs0Ldfv94fHC30bIQiEZS42sbW12VbFkoYUQrL+Y9QK0I3C2VqYCIFGQvJAfOqiuAoSsU
V7fZwPbzPyRi9xMTkZ0z8B01Z+tX4ZdFx2pVeN6hqwy5n3Cnrd9B3UiLQ8ueLib/utW2pC3ORKCp
Cf5uymqF5ldx+TidzfD0BYrALXq3CsELHk5ntRfrhYN1YOPkV6/m7J8ncHbUFiDLVOSbXnG3Dg4o
MOfj3sZTLJFUfAY5dyxNlu6Iu6dBE/HGByt5ExHtsyWMNH1bbAW0r9UkO+8L4JA/zcc23RGTgsEn
bBm/O3aE4ER7sNE3vv2R9UEraVG34LEfJyeB/4+FZ1ttc5M47CnTI7oOQGMOBfjUudKU7mCmNFIo
JF6QvxBXNCnzHRCNHqz6X3zXpmC0hx0IcXFmZ2+2XzZzk1GnyL9xUibwrlar9MPb5UFfelpDPkb/
jdokMEwWRWuox+v+KdXUQg0OPcQJcxUy1C/OXRmp5SEe9zQ81ZE+iufRheHcPsHl5kMtM54WVjB9
2kMcSn2eJA3CgEkFLqhKzz0ObkhTWQLAQ9NzLcRu20mrbqK2T6YxCONRRpxEdvBJype+U0jHHKzo
r7vB6y9JkxTtYgiceG2mkpnChaxubgFzKXQqMMptRGZkn0ZqXheYOwqdwjvIb+0dhhFfkp62fSL7
t5mTiLpMd5R2OXwAc7WCEOF+lXlKc9gvG/eg453RUdiqza485o005LsOmqdQ+PeXDMBvvyLR5CeK
K2Y7X+B77QhjD17d5G+EHT+GcB7oQN4vNAQTYiGdl338L8DndUpkbWfOQxiKzIVcHF56ZvHRMErE
HWQjkD/8qpee5uzagRfgv6fxWaCZWorYFdjL4HzjyxVsk5oJZQu8OlOwqa63WPwEB3x9g98ukFp2
f8gQrxVzlNnr4AEAfn+2Gr0clzDKoJzjNpmhNBXU/5vDXkKhj1pXr15lXeAroOdtLwYjQ6DfQW22
+AAhfVVu1EL6202mhgnwG+kHSvusR6sD5C+/FO9Rfj2bqpEArBlYoODjvCrIZwQgK6jrsqbTX9fe
lntonjE1FkUNXQWLPq7jsjlOE/4LLTdvMYXjwwkZWlwdcJr2CazCTR6nXmzh32xhMtt7GNnRjzWx
VHgV5pYife28mh7jBar/WoXvfpKiJnKcAtNoueDylC+G47AQf7ZmCSBQkGozNSTDe9rXZcOqROlL
mqcZ6Z+igDfrVVNFcqeH62fHWEODX4YWsWZRvpCU7/pW/fNWybEx5h+FoQ9CJ5MxO66mk4sKOK2/
m5lZgD8czQ0mAA9xPLEZspOLaqyVvGNMkE0s8fvKEO7ROR8qou6+Ozh2VLoxW8WQqtPC5lf8WuDm
twwdUFff7ron8XO2iWCScNJDhukJVGeUIfuGPF7uvZe6FiNfagPA2jyUbiD0y3wlE5Q1TrBCRNRs
emV7kZfQCzD7uyxyDW9m0mNSsM9sIHBfywxwwp6D0+EvvYOh7/olXq+5b8FCSNUvxmGCvsE/jnEq
jPwJHEESJqQIfgogntUNgs6QHiDyYif8neoGcaw2A+aSPDJdc9vWD+vNO8GEcilDMjz2+5C51XGI
rWtcp5420RmgHZl3yWVjdYk0uhnTk4EIhwYpifdbL004HxL1gAtAJXyDWJh5UfMT2/+NShnXwkHd
v1WlRGYXkZBm4St3ENcNQUa0jmdv+AYAxkwkDpl1YS7rIgP6dKNxibm2QHUdXzY7yBqOAhm2WcJs
+tm3keFXljVgdkGCxcZtxVhd3NRtbXn69Pws2Zxdg6wuEo3Uhqgg4UpVHq3kpm8lsLyFQYR48uzn
5KMYdtmW5S7f956gpNo7k/Zlcs2k+j/DY71lrxkksiCnTP/AzcShQnhWbGQPkuOXcxAaP5NW+8U/
3JTO9GHd8qI0ffks91D40vVlLByhu4Jc44uARAXRTlCiBu0P6RIe2GXWLxxAJoPsHLaBHo2wG6se
9/RkBFy+A2LBMiPSxBtSX4ZFRq9348yt3Ltre3TJeOCrxWyh1J9ObXRdX9Rn7J9uUKi3ETArL+UY
ToOTpsUtC6EUODkiREYaO/wjujv7wC6KcZmOQ9hpmQuc981hnHjQzM4uIO4qYqosARfEdklgx+su
80Qdw46TK0wkgnCeP2L5az7t1E3MzwWfZ+MIxDjABSAyoz3WlThDEmyJrBYGNBW7N0XTiKd+879m
FdlX0OZs+A6R5zgerh08nB9BLyLYLuYHO/86dIhiqfOW3k9Y1sWCJz7BqJIdYq/QLxfkM4+cr7Vq
vPm/z+AfnTDEF//X0RmJIzBdGgRKfu3dGEGMqa8JeXaX5unIX5TUHKpBupVAG4LcP8fn+j3Gxo9J
Ot2YDNHsY1msfPZOuGq6/4xZ6iIqJgNHbjAwkFATg4yczKq8Lz816bj90OT1QZ7i4xlbaUb87zGG
Z17O206cGKDFzVQT0RB2FNp5mFYUoUMqZ/jcchxhL3IdpPPH92naTD0WnCPWVqe2Kiikkiq9RqJy
W/Fb2n7OV7Tdabm2juNmjyf7pND7gJe8OwXD7A2FVNR5ONPEj3xtwg/SoENGkPAecONWLdowoCg2
uUC2mTqRbF/izLgEdSoQiU4//d5nQxkuf1PTbYSbVtPsFEQbBEVR0prGgV4fxGn5jsN17267xXqF
8Gdplo4zzSiNhImy2eSAWGB+RnyJRh0V2wNFicM08vCMGHFeH7zxgm8H6QPxhrcciXPxq3cTieuC
dd62JPoteQSG6cM1SHfrpOI0YBO/5WiqqW482ptyZS1xFwzdd7Gt8KbtfgWOIP5OErmskVO6gG2J
MEZJHkEISl0HFhp+5xOR50dI4wpWaYSpBMv2apZzDdoqsTre1om1yAWuNMMUY+52crp7VjNGl8eA
VtZSgUNESob7c7NjxG8haxs1lv0yEMYdCBi3UkY7g7QJQL7LzzU83/INOv8/kEHyXf95RymFQOJ1
INUzrgv0xHXTe+LrXHLBOhAzRyhCJeejnF5CM+tDaneYGgiiKxmv3nxHmlZbVGzuKc4XizE/txvS
wa5V/IebDlnZLO5pNmPN7jE34buWy0OVDQOyKS+G+WgNpEEy7au2umcZqA7c7X1U6JOic6XrqDZB
Ar0q+dn2nyEhcr9QRGDgf9qTBcNxqfXb6pncoa9zBqXT9CexycJAQetaOus1oyBBQw/J7eyiUrQP
HEt77UyU370vbQhNzNBERe/tUK+7NdRY6687JMFK88oHuyFPs6jigAb1lYe0/cuRc7+elCRA37UX
xlFoFaGjd6x34g8C8bpOopZ4MmucBlnTU37hXK1f56vYXxfZQqH1QYLnVUA0xhDBRNtHHVnqjOIy
Iw+6GJopnVdGX02PiVT6gVXpKQZ/W/fZB9G76YJkSo/zkgyn17SMk3lzhbAe7zkhrSM+9c0i4xbj
ozjVtxV6UFSva5johLn62/LOP/b7tTwDsxAF2KASQhV/2h6ACOufAOpCkoIoNWikdLt5tBafg5Ls
Fr19CPO7PAnnlrNugNImuTRhgMe5e4GvJ+iOL8ZaznqK5kuSb/WST0s63V+Bzu8VMrD4vN6qmIn0
hkrXMELZUIOpZc8VtK55MFNd0kMiSMgYke64FYdYYN8b1PnGrPxzp9SSO51yPOOedUta+xz7sGur
gn0//wOdG2Yk2kSdnV6UfClXp24iA27/y/EvAScGvSqrjbALEFsQ0ELz8twB6W7qWGY5tqCNvBmT
uUiSbGCRTdncTgxaAWkgKcxzel/MwqJI2gH3k/tJP7WqUqwBo7kTgEqNG2kim35u80DtW/cq3q8i
1ckuxijYiRxKTYMuzCB1uIotImNhbwGKudo+Dsz6OELAFWmKW8+knH4q4j8Afqtz+2icuUKDAThH
9IdxhGpE9fRORZUbH5/44R8O15JZSFQXEUQCRNl2HeiaMK0IEkz7XAKoBYuretqu3h+02xNasQNy
23XTUzU45WZtffs5tFvQU77Ru809kI5L80R+G1vSs8jmla9kN76OSa1OdOB81RJOctgW7fc8wV5v
+r3cbPAO0ZmURzZzfrfvCwnnGcWGckxOagtmLqxpUX0BYZITLfVyKHdnEYd/LGkA65qdZmU7Ag0n
Q7gneQWyfOcWeq7/swtScbckQIzSvkid06nuOB3JZbRYnpC4E10ucBri/yViCP5A/mMSCloEYWJA
MxSCYep5tzgbu2jeKwKpeNHG6UE5wW3Qa0RMThzYKfzrjhUSiVmarVtU8uB13uHv5YigkLfkzQY0
6F62XseHrsNIfffV7qa9pC4mUG1COOw57HMixXQiEbYSm6DkTHTX6/IwB3pAaIMTLxHHyAOMvY6t
YeJZzL1YlL1rtj5kBaL8kTyYbu0jzFuzsxIviwGOcsTxB/XfGGjXNwktPtFPyZ/osFoOZFOjk4hs
BB4+s4p0ImErYIY/YJT3M2qzruIZk0Ie7aQkrRjVWHwuLoibbQp8b7Tyv6sdU1IGs6I2/Dz7TgVR
s+7YFmaNMTRnb6QElmryOINuGg5eiONpB5edD1dzAAZ8CQnSVgwf9bLpESObNNrC/+TBBf2KY46w
gWTVQopiRUQEgqERPaIMXcT2/MkR8R9OfJJ/MAnGzKK41l5MpamLE69Ewi4hKXpBD5ZE8wYUEiaY
xVS0IQ5rtqGj6a6ewhTVJEHP7RJIcVX/2fBQPL5jlPp07Zf0KHjuywc+g5N4aIZEtVcV/ZflPPlc
yKwyU1gh1UqAj6Y8TCgTa61pP+sb6eUXzTwSrBejBPNs+bTUjuFx88V0PwwLoZohqcoiUk/IHxuc
yMWp4bVfZNYv0uG7rxe7de6hNV0qjJm3sOPnUbNf25SJvoTs2qRlnhW8da4njmqWLAN31sve2962
7H/hTVFLIyO/NSvFnHoolx+icZPOkohOVGhZSg2StA4eG1tHxce5PhgQpQWNirx9UHvV/CzQqVAB
Uy6e5s83kNVyYv8hAAT7yMNy5bCDwdAy2jkXIE07XMWD3G5kAxyKkyjUbHl80HXeBRQ+pzvRTi+j
ny6Ss8nPBpfeIJu4zu+AE6KWLsPn5B0JyKF2AD1x4J0X254fZ0WKTFyZAHS8W1w1rm27amyPcgPn
2r9Zc/VH168yVGHZj21k8OEdcRlGKt3EgHa22/rfFCpTmieOttV+/ESFu4IHvMAWUl3vxo67oHGV
Oq8FmUn9AmYutlp2aqELhrlYUwu/yyvE0W1QSw7yaHEEbIESE3QaDO+AbFYxhkMTxAB2BgyhPnj5
GkE/ItMOEPEyIR23t/WMGF5cSeFiyCY0iWNB1uXAAYkRhZc29EVbfFnUVsaWGx8oqqwgKmrTbZ3M
99rh3jm8wns0a6t1ikosGKeLmEDJcjhng2SsbsLzd+LwDlWBlUDtlpg322alsy65Xf7X0hBNm9VS
HX01K0dRk/SiAMYI7rppGZMSrsOAhojgX7CYYXsv0MHWJERHBFDT4HFDVUz4afnxA41NLY7Wm3hw
+jL+SpFUcgb5pmd6RdZIg8+JJi7HYzKnkCGqmlrsBJ+stoBLO7lHABpEkTSgSumpnRzctHhtkdjC
0VI0hb/W97IxVgtE03YJ2YuUyWVD9WdGy//NiN3yMG7s0lCSp8X0vwvZkmLJL8MixVsOzmMN86kx
lkBFLxe5LK5jzAso7PNrwVA8w2Em+r4+BszZV4gIar73dc91KbuBnhLJa8U6HE+DZNskk/Rr98Ke
TGTKVHVP6T5cofDbnHRwgtqh7iGEXc/3eZwinysxWIHKc7k8MVLcFEmtvvNgrS2K9lqxaatgkZa2
cklT0VqHgB9wz1Akbm+5GSMQTUYCN+KrE5/rJ2H/hxljIVrrfQ4nnNJh+1MU/lFf78kATK6Eq/7B
wXoSloEat84oa/jjhj5rqhnw4kUAIbKgpwbMu4u2dte8duVSK7AFCBNtFCXXrDsqH1Yji9PmXOQs
r+uMHWz7TvSdiiUVAtXS3ZVSszoNb4XvRWoOXeBj37s2pr6BMCzUCl8w7h4AW0xbiT7h2IKvxWMO
lWPpmkNEnxb/xyJXWgDhKuEv1wIHc2szX01tsvXKAVe0eGBcW5f3DSvbl/vAvzAqrUASAmstMK7V
SQRywQOWf1Kgb9zSGozpEVBDu32WSHOL9hUKP6qE9w1aUb/K/Eg+R/nR0q/f8oDArbksRFjfrna8
APFaoa6ydY9Y09Mz/6Qur/eJffHcIjYn6wxDFA0vg/dgI/8XdShJXEVKiZgUXLuTgqsZ9g5mnUP6
3Hd178ENse/hoXGtC6ae/J2SE7WyuQ+JSBFoAkz3Buo5HC+Rq5tQVwsSadKSPdqrEk+jyf3KAeAK
px0kImZOcxYYK8C15+XPJnwvblCGq3dp399Fd7iQ+3X6ebq5qRYfXgt77Egs20bby8+eM5MxJsA4
5fnJN0vom31SjODvkYSfkYCT/RWDEAueFadsrXd3Sgg+W3CVgtcCwyrGCbBAeryA+VE1qeyOuJez
6ygeDYrctITmnDdr32e4Lg90FyTR5jzfDtQsbe23a1SpagPfoZDy5phMnt6UyKZtqD2zK+Rh/Xs8
o8IhGE/+o60ewfiZcFLgMahGkYwf0gIt94Dnirx2NDpySa75Nz3rUV35K8QRBRFgAKrJwfbSLitC
ZxRosI8GYqC2bnR29sEmtAmtkOm9yG1vZQr/OjDKmjeZvheSDDtZnVCgjTUnb6e7WXt67na320/v
MPxCFZ2NNNGsFlb4T8Jd/9tqHgjGzLryLcI/AEU0DJCskmuVnVfKPyEcAWRdFCwi05ActW/yLIjG
bjgzZRbGZ+fOS1+GDWdsUD7rvVdJ0pjjMYyLTqa73KBrzuoXgP2sC/qklBfvA5d67PKx3NkQjXWK
k1SN1vBxq2X71wkRsbliWTSxbwvvbEVCyY9X7N5ChuQsxyNLHAsB00dLa6T+R2IrSENOWIJtuV9Q
XqpBttcUur5k+9OA01+wlOkFjWEBDGNQcOzuJiB2QhRWRjpI5cmuorI0t3P8sf/u+6I52+aTiu/S
T7Z3MsK16fDtI+v1uk6qtH+ubJUpExWVyanOeytu2iaYM4FsrIXceGXRTPglAbVt40ropBFngIKs
jsWmOjgyBIN4L+MTT5YFT8q98wWvqvt9zE/usMg90Nw3kZPqDuTkoew05UhOUYC5vLOuUBur9QUX
H2YMsfG93KEFxf7K0EK3aJJq5tPxc2QRAW6zmv4CvJ2b7AIw8+pioBNrpBrZDC/K66y7wksyY16x
Ok3MstkuLYPCwDw7xq9KSblId7Vip2RM0wgozZd5RgdDAsx1Fc0Ze6cvFuClyTJsGKAAFjenVzWZ
9S7WCRVeY4oJJXMGfdZW0m+jbgSOGEAx6kqCbntmm00qgIeFFnLtVSdIw5MYzbtohPHvZS7J31RQ
d8JHksMlrh3Bd0VefHCokm+0WVUlwYZqSJYr9dlx/bsRoxW4PAWhpEmv85uYH8MemlssEGJniMjZ
o6pZ5ABRpDjdYT4r6mfmExiYf/Hx7cUbvV1wRUdUzOd13tKTmVLz5VdGhDJobr+dUwqfU3QzBsWl
JxXOxUClC0z7ZA4Lx5EVsbJO1EnFN6DjmKrRwfhBV8WTVwIVhuTK0kWYEeadHf7LuHbWbg+xQG1h
V3vls9M2vAYb3K4RkDyAv1P851+eZ74EOux3rwL5avte/qCgNt5fSWDGzjKUV2pvZxAW8J1FCirN
HODKjyWuaJ/L3LMRBkp7oz386glKbFygKcDSuL1R2ThHj/WpZoASV3NxN8droeh8BYsX8pCByuLi
t/H5JpOJ17KVFzriE2CgnhgdxfyYRWVrz312fr2oe5ZcsNTU7EsDY7AMc3BQEPCO+hNenY+mwoUb
ddMSJwQS2knWJA0egEj3VS3U8EIMuZomVONBTzEijngjACG3eMvEdWycFbAOWG47gp+rH7xRX6t3
JiGdwU5eWhl+Djrr9+rG+5KbJ2EzH/8qwWChl87ResRWAqdmQao2NTyG7bxM509kfaYNky2Dtv7/
GI2jAnxsCblR5196vjVqOPKupaXpRWHkZIFrgmjuHBHCNNmFrdRSZOtmWG2W+h3Z98gZKOGWlt0j
ee42mPe4xHgrwGuOYOtXDDl0caYvjgw9ReKX99frO6GqAYxE/iUYdpXwCty8p2q6rA/6jfiym6Qq
RB77FAwtTzKZRtqefBU3q2LKYnIu0x9iLq4MIrUcHQE91hK7sW1cUkK2W6xm7U+09BNCGNgiSu9E
otk4pKAk5YHS6cPn8zb6DaDMb2N5kE+csP7TAskIa9Ja2Y4z6HLhTvr1zDC0P3VG+kS2ZMtnkuAW
O76P5c31MLwWbSbv7JW63ZEywAiaViTKi05Q5ryEOkKnjSJTM0Eh3/C2E+xOGXG0vrxlEtWvFJ7u
5/iwnl9+40eL9O2QzPVhAAY2BUUPcPOH8Wg0yBilhszXZ6431QkdNwIsuy9Svcc02HhQz0DngGJV
c8O/wtzALPLoXDNF6CBAy89P+pybWsdIq5+67CNWfYmjJXyDAWP3qweZrV1gynx/CSAxHYlgdNwn
avANR2mUPrYGltVAEXpBm5SGUcjS3mnxPHKhxIG3t0RrKR3WTuuzLIa4F4h10CD48AskMrY69qam
GDMIShRrKnxvCcz/XrZDq9uoClRRlW8oqGbMKeQJ4qy7Lvn6uSW2hAK6YyE0ujlsBiZqGOsjoVLA
4kS+RZ1YIg98vKqvH3nsCpDybm0UXjEJK4tfxbQTFmnJcj1T/XUE6b6Hh13Sm3NIdyaUL8kugaAr
oGJlT9PdPp7IdIGMt+JW4yx/01aXOpbvD5lsufWr0AZ/Sg6iW4VrpGQzkKIJW0CuYMYr8Z9J36ub
9IYMxDJNX3jJErqPU5sXyXvNdSTwrWSnYcT5gDLeTTeRAqhoxaSnYTQ4fPl6Rz1b6qmpF+PR1wf6
hghdPAUaARgZlFePX1rMKYvjjKkAuHcX1kiDqAvXKl7HkS5RMlUm5XBIKMaa0CA7WYSSnQDpyZ8t
xDY1gWd+2W7+zYAPKZvg7DPWuSNSjdkwbyUzjNVsNrQhJPgn1Rxcxt5vVy/MXQwV/sLOHh/YfldB
liwkpO6p3V2DWhi5dKth+1hSqqiiUVNmTnynqmrE8IXUyi88WZzQ4PVRE32akx60h0mv7FMEjRpD
LU+VMF4dXE7RRjxrMnbOOub85pZ1oSEl+58nlRo2cHerVlJC1csbgoAWTKdctRnE/F6epBSSSpPZ
RbkbTN+G8rmJbt4zkh9Rnl8deFWNFhVnK9x8p0yycZDRlpFW5Q3wEb6hD78q+g6V4WkQwOT84h/4
AJfn1Fj9YkyDLuvdsrd7lz0wnDx8Vn1d5e0djHALoYeHZPlw/VDieLIQp68s81rKYueLTjCt2t9n
5oFMRG3hi9H5VjM7kM3x+Sdg3tZ53ijjHW8IgHrlJbPpC+tY4aG9xxtZh2FW9CCsHFd05AdT2uGt
7btn86jl1TwtcfXeRaBwiNuEgyiMDEC2cbrAsddlVjNYx5uOaQvv28XsT20BA47jTwesARLdc0bG
4tW2CQ6CJMrJGYzBonbMOP0ADXS5Su80HU157w56KZwpJ0sE3RRO00HpB3RhYkMQdM3GoSFgILbM
rwt1Qq0cZeYFdRoFH7H4Zx15YV//Hsxw2D/VTqFKYjWbkJSv9miNKPYrmL6OCqgso6ygf1/3xRw6
nvRAzluN2X/hxOeUY0r6rDFFPeuvc8ERmvitPBOJ2YlXNgmP09pZer7fvpGBjJ6CdwGMP87LXj/u
oJ/Y7tF/n64nfuAQRuzob02U9SIAb0+0TY/HztEFPs3xD1RR49TJpREgzKDuBS7+UxNSNJXzIA8l
OPL4bLJVOxWMgIRIiKAAbNNfuz3Uet1Yt+fPd3fQ5AypKqQGdIug38MK6hn4x6PRjW60YeCAoyDd
9jRyeK2zA/eBrhN2zw9iNN7XSuTkolo07aSBp5riCwGK7QjpxFd/BSDMvRTFFvhfOkhSwYYRYn3r
XLI8cf3ORw1sDwnfBF+1Mvp4AR58eTTodouUnWiEvEu4pBubBh/uPLe63MCz5WdwRzFXIVprXdNR
Pxow6p9jrw+6OvKE7FIkQ7R9GG/ryT8+h+PuFS1ECGx7qvzgEJlI+Od44Ne3f/GnSq+SaFcIQpXf
8DHLlt+zGX4bXA04o/SvP6Cy4OPl22bO9bC4IOOy5IKAQMyRc3MtGDJikQdZHkl7ZZZT+DRwoRsf
WWsj7/E8+6KJCjX8+woxFw37rNaclDRnDhPibpxj9omtEBIea760TkKaVPyr7IJAWe1IIDwwXVN0
XENOxapt8veW2nAczjCPd2GwIXRo4HNCDB87t16I0EhHpG4XGlqJSdozQyNgbxxBEpkzGzWOzB/A
1rDmg/3CwTUflVOM3uNpp09zuIczLnACJCNWdr6MBDsICpSLbKef1ofKjcaEZelEwDM4zL9OPwtr
FEuVUaVII1k6Gs0acpRhWr5MpnVE0NfadBzQ8dVvX1hkw3nMnHO5z55pgtggRe17YqeZv07ufonu
1/P/pQtErQAZLM8zlduDT/xp/0CuSYMilPo9fJCGdLx9WCOaAFiicq53LZgC6XbG0m8qx8TYdqqP
URVllI3ykzc/JLV3Ba5EqWZu5RxGBXyvVyd5uTvbx9YlML40RxpC5t6sxd2fk+M22uVjOhFx0LEO
0yjAhlSCPd/YGMsrgtFTUA47KwXt8TqA1wZgsFJ8vCl0WQltKRoM8KEjgn1VaGGr66hH/yiVHyrS
+SA3UxTKLJGW9AhGmpIx8e+i8UZ4XOMF1yionA1UyksJTK8ac6IBdxaXrXdWbXp+yWyIJhmLxMmg
O4hTxf6LVZqpq8dRIrfebS0qwkzGvyMhxi+5wCD3lnsGL3vi6fzeoz4rsr+3/9Y9SAwfuwtEHDnr
FYI3O4E+YAUX+ayxN1cpcBXc5utvUL2Xas15PJDn5L3YzJdb+N7zX6llz/xdpWvEv+RaUfSaP/8l
kOYxbylJyRsqyC80pbVeJ2CgVpzFlRUZQGrHUeh723schx0r7i9rTHeqO5DCDRVlrUV2n7VvCarR
ADxb6djX6yHzD/jYJCeFE9LioAKrCztwhEH/v6vILCEtZ3qAk8jpoBnpbov1pB3VqGmCjMpITQo2
6IaUJPoGHRyh3Lechw6Nc76KibVuaA1EXn9Tla4pKHtLk4BHhq165GJhV/74O36DzIaMNrakOAOI
Vo0ND09nQaUpg15MRR8YL1m7GqxcNRIlxAXKdRF8gq3OXJFjK2al6piYeGqZeXqof2LFZEJxhwFz
NG+UoyO4ZFLg26XyY5DOIVJu0gJZ1JRU34tedr/dOKcL+vm2ioqY1yGV9Q8GWmubVJVdCRz9BYHG
XFBuawqXeqdqmoU5HUq2vequGESx7Wgg89EMzQAMbiZhuczpNVBdifw9zs64D0sa43Ho9TPiEJge
e/l8JeqMmUO6LbnZmGoWByFqyY+YeCkExHGeHgHQoD5/fTAGhZA4sWbQ41PyP5+ElofMDbi3xzgh
u4i/O/GWQS6ekuIkRMB/JRZIFtI71nMSCQcm/S7IWNSCRvaDFBs3FB875QWGMztTK37Yiprjj+Te
5XIE+IXSI6opZvA2faFV4LwnsK3t9qKSOdCLKxLZUdVY7bsfQIpNQydOVq/TfqLY1I6OFz5ESBZN
E+R60FJxxD4a35uNuBIIpl7p29NmUjmVhDqY4940gb84UmOI2TxcOWFenhho+mzEjXbNDX9Efoot
28j3r/WK1NTva7Z+bX128djmhdL4QjKbO2d8X14ieG3qgd85jNpp905VyKLv0A7iLn388v1yI1fO
lLkSnxP744q+z88lRLrbV6+ZpPMX0C3hRgpdlwdRl0VX8ZRaGUQMuDv8sADa2ECVjb8Xj54A8cVt
7jjtkchkzTjOyhBU6AZ1pl8f7jhZLhLQMhE+stAkhBmlCLcsS98p57D8CTZLTZg3ljuZJy6T0YCS
5QteHa2kv1aWwJHB2ymFar1iioiQrSB9TSCA98XV/eHeY0jKloK+2v81s1nQFv7kOnHxTFNXOMfu
YJpsURLIkik0XgMFv/a70Q/TxJwEWwTvL0tU/PuZNwB/d+ZK61RflgdfcIj5V7HkHl8YHvCZhcbz
J8D+JUYEZ8xAts0hCoccVtlF5ZMq6zLlYvZc971tynQ6ZvabYzMpHV0eioQLy9l3nTZXkTF/vRFG
O2fNy6vGiwfouzYoCAYn79qTPSdtvku1b/5fWrT6nJ6w2EpO+55oH9Zkniebk2PbTuxB8lV5iVMq
kC43pEjK37fENOqINEYpA4MB7syUvUoAwrj8UQ7oF5A6sEP/3J0rmT1stwFn0kvePABklDDczHs+
kU5J7ZRfhOZZdZi3QJPYaSeoAzUgERgpx3DMI4Hv16CGD0EC4xu6cQkQOf2iFdYuYtVP96Qx9FQB
hQoROVy3QLipOvlj4t/zttBRHT/jQ+Auy5EtaSIrCKpFS0jAmSDWY58svH6ITKRfGyCWOnkvWFuE
FOexeqSw6GbCqdv02UPsADjfJoEAVPxZqY8gWP4tZ/ElvyBBpgRLXp+cc2qXXdzJQdlr6gDyIa+L
GKMI+DrOhq/WujAt56Sg99tfGwQ1H0mBL/m1NQv8x4hGfLdBR5G6PU3odSVvBC2J2paSolIfFyZ6
e0Z5ZoHCZjEBJK+gX4amBGaI3JsFQVfpAHO9+ZE0nSPMkUN8aeVYOJ82O76jwxInsr7ByK0fGkFs
RoAEKsAjunGf/GWjZ7myUqeB9Vms95+FAP9Ydv4pXWVf3mIt4dHd+DIcbEAZjpPOiSYBO0j1Erg9
WeFvcxi0vRqFWYCRQzZfVShw1j4K2l9NJqjYuiazp33uOk+FLP7KV83SxZmCl0OywXxugu6tQ3ap
hF/ADJ2Tv5S7DZZ7u5oqmuihxJ8GHAeiMzCJFn0aFYcNrJ54/Pg2pIbR0Pf0ptb+NPSg/NpX+t4S
etkdcNubtpYm8mZ+5TQm7N0qnaKvF35wNfE0LVuDrFxenF3Z/e3gwIoX37MCeXU4mnnsKJ5A00Ex
F0jHa0SdZyFFXL+ybtOVRHZAFM12+Xerj0EDSFnX3qYQdN2ukprxTtZJ6ry7oyyWskPUB92DhmAG
x3sMwk3GScexXzBrlz4RFYFjq0RubDs2A0+tKqf381vwmSJdcY1ZuFhJhd5yMwUZWAriFhvKqtN1
iOffFyi767I9VzbPsK3Z/u+QHhmcCv0A9olUNc/Q6Eyv1+Hf6Kla6Fn1p6a1w0PDoL4J0AihZV96
Ztd3Vo8gvzViNxT/noahJaMLYfKMHpNw/2bjhlMszj2cxn3Nu9PjZhF3arqeYfRHgxwPKz3EDokg
JbAti0+Wuq3wawQpHJfYB2/ciPHULajqAgosHh+rNz5gPgBudTy8d73cSJFmeahiKxSfotDdimwE
iKTm1ZKBXO3mc6PToSq+fUeANNOTh4BpHa9RATozuRCvmzqlg8JUsaHAr4f3tapOoacTWYP/IgAs
GJw+KKFqFT+JjmeU1XsvkALEexCC3vva/84z9998neFtm17sxjd12s+Gs1umGuounvZW8LxzcVS/
zttqfyDjDsJx9D/lIuqeBFbMqkwRJI4npRQyj4m//x7sEobPxJgFvjdHc4EhyuwYTCmniH2QLCxD
kyXO3Am6ejcxq7U8T11EfNsp1rGLRfePaMxJqrI+V+WkHoEywEq9/zesyyhsy4oLFVKcc4p0xoFr
E6NQFh+KI+HUdqqKpAY4AQzhLgKdHXEtaz8EeA9+kqKMbD9LTZla+iRZS+51TCKWa8zkY59AH8hr
EfbhsA3ZRx8dUZqzYAVYiYKVYHcCSKRddscBGjZ7Jrz1prz9SYO9m6Ki9lw7YELdhhlZDN84Xmyf
A58mndnBBMeDPoTcbQwetb0NAPOekqut/SKVlDqTEE2WT7MID+OBnzwHh1w6eN5Mr2B/umRR3y5s
tUvi6sxoJnX9mFyIa6chHetk09I7ZvJcjkYVamLix4CFPaPPgZ1NrYPQfvqSJdwuYMqRsh3eNxHv
lpyLAv0y3Ewnti4p79ydq1yKKhNVdb4OYsolZL4zNQVdb4hjbHpWNumFRfG4MGiAd8GWvScIz71U
GM4ONvtP9f14dZtTAhH4fM/R9m9KJuHDn/3UK7qNbgHlunlVXhvE6zXtnL7TsaXjzGO9zl+IpvJZ
U6AOtQ35LICWoTuSbaAY/UNFnhpW0Nzfv8NGRQRZT1yQdLoO65Hlm6GmOPkmT3zu0hNAjumBo3sF
5FJdWsny2ehaxdRhhnpW+Ei44ijuR//NvVYlRJSQ65BJhJ/GHVBkjAO++TgVKCOHpZ13h8pkU7rZ
gBzFahrQOoNEPRxLxmg2beT2FRYbQZO7ycI5vIbPvJi2JtixdHdMKm5lHA+R6ngswAgYXbLbZShw
xQ9w+kWLefLkE7lcjWyZ4VUgJnONu7ENz5ZGDKh9RI2eF6yDwaGw57BI/f0nhS9nAFKbn1t/47Jg
yH9VlTnlXMuMqKEU48iKgGc6MLt207/n4cEqXpa56LffNLh1IqOUOSTBp3co6pQESLL0E5bOU2es
3JQHt0EXMWdouLX0/Zet5M8Z91MkbNjlWybXjQZNgW8jNU3KXJ70PttUW8y/eIINiKVoSqJWF+46
DepRgDa6KG+uz2jxIrINGcHN5sdUXHoIrhFthydRnwGbEnyhNEN4LRCwGeTE+ouArllGfah6k/d8
01R/lYG6uEMHDYvkRFJJGD4/2wvGm0wU7wC3Q4OOvAkjYDW3rUsNEZGVyZmApw/f/Sez/98ooRb4
mBj49jT0csEBssY6ubgjoCLZIX+5PjOa3FFylRvFGJh6JUiyqupCVJ64IC1kwNMShx/HQ4sH0Y17
3xI8KdclVrGnH3h8CYp03U++ZVBYWyjOeBHP0YIRhjCbmdpWp7HqJyncguPT3QkXJEvNuxIL5oAW
TFPCJtAeazCRhotjRBM1aIf4LQhj0mmB9cBFQLEiO9xPPtH1+7L1EqAnmavJjG9HVNNNI9Ma3uZU
zGjAP2QaMfZglGEOp1lSJpQC0uNlulzhZb/CDUQjthc7DAtU3GDxaQFsCaL5KCmR1t0SMdlgGHdf
OS3tS372YbJzs0A/SVeZJOeQsOqLrojn7qZQuY4YdJqgCQqxUOLV4wXnLFTGURxf47KQ2jPhUktZ
4zlh01P581QAKn0yi1JuGzBHifU0TDCrr/JCQ/su8Be6c82fEGDMIX0WQhWkewmvbGexQALcoEYW
KiBnDjLn4F+r0NB3CkSV9IHsuQyZupaO5lveVidnIbnv6jfSfEj2CLxXsRZw/iW2kF6Z8JVFb8wC
q2f+dFCC6DjukGH2fdKVHwKBBNl1jbYJhjhQQHG/tOfyZGc7/Dkfq3qIGeyg6vCeScHIRVJ5ztE0
cpNDZ5PtEVqceCBtHPb6G6Lk0o5c7HGF5U2QpgU3s/GXux+nbC5bqdTAdYDd0XZYmp8f/jATsJUl
RVOaricYs+HnlF7tf7av3/O2okDjSEfyw8LBhdnf7W9uxR72Ut+ZFGhb1eaLbsarW7qbHHajtulS
1eTnvKtMAHI6hWrNbs/y+dBT462hprIwrP5fsOcRxP53jRA1v+EykH2BSnSbqdjGBflLHqHzN6tI
lRDpik6AiuvuRJsPuI4cXar3BNueZWLJF+S9tD4SHc7vhq/b32Ti5Cnma7r1yR6GgnDNxY2g4U1j
HSm+mnuC0hfwHSi2XKFBaa3JdjamoSMwHhuusn9jIBa+FFRHirBRx0qNRNA5JdlVi/KFHkLw7EGA
eNcqEkkjHS/aKFldQrWlNtvijWSU7wCcXLEXLI2ILZfMpZtshh/bV1m3Hzd0uYzuLJ2cYFeksR/T
IQ6fa/BTNSs2G06QecZJYp2OlNWm/9gMc5t3vKsKzrXHQ4WyY4HxKlKLYK4+CBhOWA/3kgWgB+/x
GyDP+q0hZF8S6cV4b08X7JuKHEMv5lKcD1KJU2AQnmjupf5TSNSLII0hR9BRAHHhEUu/uYfRTZ1G
X0dhCjezynDBJy7odlX59nN7+39+P3d11hAF/wzOtGvSXrI99di2nBJ+hjSRLD+JXAXH5x1HVLv+
RQxNq7SNuvUBjh7+E/IRWuaWGtNxrLphuKA3KCBUXYs+Y6+uXpH3MHglbCUXaThrvcbBWsnMOh3f
1DpR5tG53VYsB0E4RNKIv/hKLaP3zLNV7S7zNWsiiZF0Y9i7gJy3mj97Kr4LIPZYltw8YXWU5vwh
pQwgBbTgdWfvabLjfMsUVdXgdjcDShvyDUh8vfMyY0CtxnqNzMZjDyyTGuclCphleN2DRfW7NEc1
16mzHbM7GQ6/yS2rSaxSrLSy38jHjU/4ZuA9bI8Y6dUsI6VaMjkkoi0nhDorEvK2vtKJO2bU1+Ju
OjNb3wlsmBVp4GpHB26iB3cfm4X2qx5GVRNM6CpmpSfycUmXfSPeINHK3kDmBKEp4as1garfyTsx
r/fGsLALJ6Ygq3HBSdqT8UDJ1ips49vD2yj9/XfUhrCXIMw4twlny+GaSPKfVdiBhOL+NFE6/znB
6Tuys3wa+VbuKLwd2p+Xn68kU3ijz451so08KE0bIS9KzKqrPbqOmwQiRFjJsNXCUxPDmUKE4Z76
vwCQ1Znq7dsLcFFqd8qhcsRDD9ooChkbvBXqLcQXFlt2C3CQdb8YT3dLBfwI1mYkcRHOs48isoSZ
yQ4Q4xmsPJM4JfKJugn1oBfKF3vkcZkSt2qIDOCeXpQKEbXcbj52lEP0lBd0RrhUxqBCdtlqePiu
OSo8ERVPgkgcV680grYvMyDc+4TIaYb1Oe4TuUeYMqqx5CTbsnyKBv+uThKu6uSqgsSCUQ/Q+r+X
IlqB95NtBpi5KFJX+7tIIYLTGVGNqUckSNfHd5TmOc5IyQLSbSrrT6J6J/RvwaPje+Cz1zVqL/Uf
xtQN4/IGy/fgIcPjK4cu4cNNZl6sKQwxU6hEt26u0F/rQ2Cs3PXguDEU8fcyZd4chGf7HNZJ4+t3
wUKBLKEFsFsQ0uJCJycgzBUr89CrBZe/cfoG9e1Pu/bs4jOovmahFSKlthvFzXha31XYzQcbHrtx
LJcAwsie4MmnssxAzJdv6BuJzHekVtU9yiKuKFvX5PJwe6NAqgzpLtlmPz1RzhDsCc+OaaTp7XFu
LV7vpigRFacjwFyicgn/rlGniENEYRxobB0Df9CrlH5VQlL+ZPwkR2EdM222jPmWolORa77Us9Ee
+QhkO1J1b9n6rPPbqzkM7fqTeMAtjkS624GvHlcxmsZNJJbzI/th5eP9JM83EFuWYtPKDTFyuEjA
65VPek0y4qaeqn67ML/fItm0dWrK6nDebE09lMtOxDLmDIsvkV7fpSVwy/TC/Eb0LU/yDSUa/CIm
j6erLFJrl/iQdzKt80wOANPfhnv8YMKAwo/QHNxZoShaaewPE3PLgdP7mN6DqjdbSnWe25XjATTg
/+BqnJ1TWEwx7qiM8zlzEIfZyUObAucZMSBXV7XqU3/qxT8zBSMpdxQRVX9vx2mxsj/Jli8hcU9r
nLDz/YZwN71qncIB9KvuXeK7QMuWnkrCjtTXWXRhOQukV04Mei2LRgvRzqshwP1ZvedzWPWwpwb3
thF1wN0qz4ZffxcgDYEY4IeiAA0hE2Dtyn70J5pWU9LqgS16qQNfpL/TyyLo2Fcz70gCZF27FmRp
EtRve5oS9nZsTuzrWF5hQZ42JK8iyWpLYqLJ/GWZ8udzbgLitExo7v8cWJvzeuBiGYofY+yHYGVh
JyCgqGJiTrkytUIgBGPBe+BktHLjp1rdhcPYkIiMpA1uB8hidi4OkACxrkfAbZXqpHXuRKlEpCUJ
CJwwSg2Iq3wNM3JIcs9hKceBPFruCXvkAzO/nPE7Y9DfOW4Y/VZy8frCeQVZ07yEi+tlF/T6ke4s
GzTqyCDMy17ONrC0G419Dahsq8mD/77E9GgZZzOUFaIUdwGr6CZz4EMN5JgfC/JTbNtHSRJt7vA+
gtJn6jgHNLqesvWYsCG6bM1sQS94Pr+AE3vxOj+aw59MMUuSkhRzzggexf8IWMoXWqv9nHaFS/Jl
Cb6fgurZlhpxMhGim52FrzwRZlAkQ7Px5tWBhUoh6fP8ShPWW3IGTTjCveGid3EXNJwWVF3x2vtK
zg+c5cawcWCrURMsjLufanMWJaslamfTTJLNzI6A9s225Ku8u1+xszXDk3e1pexDsSFwUPzuiv09
AfIx+cdZTqa6Zp+c5Jy/7Q+tWIy70x96vSxGxnKx9QyvuXBT2zKvHUE3p76OSnNH1dNhWzVBgMLp
1JdTp2q1bs8Q/PKF6Y3whk72++lYkCj0Yu0JgulmtB7eRB7LnU4ltMMCdgqFMYFf+lkMGv9MEErY
E6Fn62TJATrXaEh7NwaOMy45BTxNMKlO3ZA35L917G7qqCUY5tqx8z5An8HjLEp88dReYQImG8fN
3J01s5190qLIn9Z0RaR7ndGrAh1khlz2/teYN3rGiuWQnNNvqwsvDJRRk+x3KHwFEArWMYvDhjhs
xF92kAnTaWut0Brk37syluUdiaogHPypUa25Ds43fqQPyfXTBr8jDlSMjUf5lOqnHDl+k1qci2Ll
kwJZNvKCDUHJLZ5vzF6q+n2BPvP0ieTRIx0oKP6p5jJUvORftpMTu18NO//9SjS7dOBviYuP3EOu
6My1WAG4/wfDxEQnBxU7NMo7yBEX17ZygCQLkyZo8QdQsHWl4qECnhyAKYmVDzS2jjc8ycZhga4k
MxNCqx/xc34Vs/eJ1WPEVzpANkcJQe1l/0xzyy8TbXUJ4zla2V32NYVN3hdewXrMIo0p/gS/0sG3
f9ujXlpxBp6aWJwLdcyKTnmRjiXlK4qldNM3Iwa8o7/R35I/oAxWB9XsFI0nM0vlvqGM5oIvGOfx
XTL40v5qimZDPQvsuoHnpPfJuW2qoIh9RxURr7VrxSNHMkAbyulHdXvzZfPPTYZ12M19sj7xuBmb
P0xA8sMO+nHG+165YrjwqBU5C6/++jNvs4GIsnySwkzcBjCNIMXaXGbGupM1qq3nCBw3O89XytMY
g+zKcRMo0jceZ2ct6LZ4jUgCBexqzBYa45zC9HETz0HiZB1cyHYyNDpt4atv4TT2WaawkePiNJis
bTJYyG3B7aU5A2+oQ5BFGYRTiIFo+kPQEd6089aaNrkvqwjuSsu0jZJ0SfpDouveatF+Xvj0QZ44
ZBrk85MWl6CHmuVmJCxNtvYLvuMzjbS/4S1MRRBlGsj2pXHgF1B2cVNt2zEbBVJ06fZmI+OI0/wg
qqhFbsE+fuCMIFL8SfTV+x4V4ZxvkWQg7MzT5Z9AITthcFSGjZc0sUvVmECcC2O4VyYeYN3t+53z
FLJxhk5265jUGv/3BzmQbvqpg7voAdXVcykUoo4GIwcrWDIV16/J5m6l0AzmaG0ocIRdXREFuvNQ
D+IjmNtacdx8086aOS/GvAQXwbjiu4KpZTaYOsdyf7wtoDvfH02P+mG7duYNcKgwRbKrhfHvEcRo
J0M/rC4OEouSD2jeWgMU6IC0leBqxRejEKUo7+s1UruZIm/3vz7b/nEmKTKfGbIFVVuKvS72tmJI
bArdJttFoDJhBRfsUywDr2IvabIcr3HpDsun6aT+4FcnO4fNa8MByC7yo0+vBBFDLVUMyyUScAWv
fVT0W2wGyGbzTz4rGQJvQBQQgHJKYZRsz3nNEs7deMlceMXr+0RSCbuKvTyKOJIywA4npsN04Y6T
yobu9o7zlA/RJx9+QTjW3P+HYIZEt/ieIpSbg2RfmS6nxLaHKNRCEdIUevkCaSrWKUq00tNlealF
R1yWoX9mgVDejD8fP9vf85cOPXpibWC0GDsy6c9ml7N7w998MwoAsKx6kXNSKlUmKpNprih1l7c1
79VMJKwkempkMXrtbcwuUfLky2NIK2XqERiovUpViBvKT9T4wOJFg4PuaIAgoX40dJk3hsV+n4Qh
T3JOzJTdFUb1PyOa/uXoOKX398cl+umkcNP+/G1IxDoD+G2wg6/F3t4qswCHwXoEI0rbovDPQU1Q
PovlO4urKwro6ivrsYIyj7EouWT29CpHXBbgs8UQ0yjudWNT3xD3yzIupb2CZjOBiqFo/9iZQuN0
Wt27obwL+8u7yAu2cIu9Je5JWLDItbAY3F4d5amA3C+ScwuXGqXXtRoOCb0KubTeH++e4ITp/Hhl
ECjD7aI+X5apE5d1AAEiRL4WMJYWDfSBasGJkeTzCki3Btgu0moVJi4uKTk6sRupdWe6KetGN7ml
tn2/Rghji9FCq1j5PD1puJ0upMccKJzIXVl2/2Fppz16BfoYoGLLzlxEwB4W2jv+A+mZA980Sk/S
GbxQeYIN3p8oWgTOUJiENYAwdpRnV3FCKgqZPfwPBi4JEAewsL1YP8sR04JTMa1tsihDOw52EkTd
slvmTQ7lM0z01C1aa6fEy9U1r8z731t9IDwSraa7nKRBIn6jXbc3DvsLbdYXYFuOgqv0xRA2vcd8
BERWfsnJ2g4fkdPXc3a+QUJGl/CnSCFJc0ZE6y6bdc7Ho9om4MG8sJhWo47Ii+ZZGW103LtUpghr
65kRC4x6lWnChkkv78KCkd8BWmIaQTJfCjNLwYmNTBNwenEw6lH93WvLdliHpOePmzKVx0xRAkm4
QkoIKJXLKEBPoiaa7576j0fKixpUPBiritpUKBTZWQJ10W1iyFHmJ4pX0OtE1Cnz/zxlIjQ/PoFa
klw83mGi65geE7UNqmW9K26JUsMXwwJJmP5NcyqXvJ5MrJ8/r+qh2outdCALAmVJTBnQrnlwBxFO
qednmf0H/QyFOLRGcj5m3kgXQ9BLVbhCv5dzeP2vCiGnzRkLCgAMTfi7uBDFLvAvz2gEhapPw3az
d0JASdc1zUTzBM1Pshmyp1sBnxidJAi7WtWtjW0FZ0aGmyXnsbiL6sbUAEtjM03GL0bidRi5m/Zk
k61r0mpoyeoRz1RUX+if9eRxqFvenQQMhzZ339b31LRGe05FIqHMAvrCdDNdqnE7QOri8vYEKZp9
Wkb64zcVkfGrF8Bnr+zZcMrwRKhApgczeSJcnI24d85U/8lu9yZm0YWoYoV7jxgB5M8R0qayQmnG
DNlP8lTttCFeeSh9Zf/MmES7xA6XIVwnnZ2+Tqv0SeAYBIZuBC8eMAnat8uh87UI17hoEb9Ee76M
E3lX293ISOVnTqZTZH2sUqWQWtkXf25rw5a4lmjkK5sqxGgqFpQZgXN4zd9185NaS4HoO69lYQsb
ClSoJt3BbksNjH0FnQUX+WZPQqn1PfYGNHLEPTGTntKvi2yfa66/JfbuJFFyKUBj8dCbdbYoi+o7
eQo3920Gi1zHmQRfVqc2ifcyX5foTPOL8B4SoTXu2WCg6O4F3M4Vh/KvhJuSRTOTVde6JRhrNZdK
4u1JvbjLdYt9eaDCYy+5L7Ij1MIGpWOeTgb0c57N25D7TJKFieD43I3FBHXFSTP5HAbfvI8Ds/LP
OFwMiyUB6xcfAvJ5L5mrZjcGZ4vVGpdNDB/m0LnRO+8U7NtyY13yZ7ffYD9ZAVNQMi+xi7wfabuK
0jLuwf+kYE1GgEjT7vHi2VA7MgDLc6LopX9gKhLH6jvnJtbuVpKnj4eUC2aSHe4dd9S+1OmDpV1e
N4PT5bkKIV9Rvv9aThdzaHRvRkF+m2tMtW2NK55UiaIX0K7L72bxxEtkgcQFuQOAW5tA4z9j2LYf
TqnrJeW3Qkx/mZGVxsJ3yzZnuBgm+cNNobcY91OCnMjC1QjUrM55NNm/DgI1fbaXXf+4GuUyYMwT
i4k/Z2aApthhDbqXfhRXyEZ5Y527xxkWLZc8tpYs+6i8yuhrXTZQy4eqjzLF57a+nhFNa1Q/+7S0
Qg5B3X/LANQ3reMSGg1H5Thl5WTPvDchD9y0cU8J7UnyarcRBCv5XVT0ii0RSN/BDBFZXYKrv5wb
oFSNQqqeecHQWxQ+9cJ7e2qUNiNg5tCpiVukzSi+SBGuyFofnU+lCKKgCBlVz3f43WRoGUjtXXa9
097POVf/6tWWh4JSnN833kLxUZk3ELD3w48zhIza9d36cTEnroSj0UCKKSJ1X1aAbX6fNIA+H9eR
2hZRn+q2XRkOxcF5sDoLZwiDR88HxlYd+GQJr9sENW7U6f6ERvpapBFdE5lZP7VkjvWgluTvKjZb
L6zRVBBSWfH8Kmf1vgYVHluGO16I6E5UxPeZmIuvWzzV1IRl89fI5JeSBKsKIS20YokS+sTkIXPT
QKftPnEC2YdrjKuaad6RQEMKPxysXnjcuWxraBC4uGKaLWvCnMiDCQ79CfFQAHzHyiCqBoXOcyhE
6ZFz4XttHwzN7Q9V4AWSa1h1tp2yR4wFx0Mx+RZdWEdgIVyzIS0YqF+uP2kJotszw7erOiVm0UKD
xC4iLx7bvV4kMuOR4O1XWy0d9azI9ofl3GfUpl9hLjIHr0z6Yx4YrE4vi08uNTNGs0DQJIfR3TwX
xFTWcSwkOD7HHlN+IYYon4JFBWsaA/E4Ao6rGZbQzvwy5wdtCFKhR4Nz7NEFkcB2jM0Y/ZMsIHVa
7Cs6H9IAWymK7oRTSJVV6BzRw00qm7X2/Oeq96SBk7NTbfdLaQ8RMgP82i7Krhjef7TGp1Luyqze
BLKiBTryOFu0Lee/H+DX04htMNBroIf1MHNUTK6DSNDoWR7a82Kljl3xkAdyBKoUaTDKfOElFhhL
ujg/dm7HDHXS2YlZm3/MHjbEKdg21dhQ6TfNw9SUjV+6ouBe8uwA0QhSuk9bzhLFiurArEjB/dlg
jtGPQ2hS/mTPeYGlE+ekAKg/fE13DooNgBo6p7lsB2k/CR0Zgfl52zmUXG2GdtKa6Nhhm7XNSU0o
edEdSczjRR3XPI/qR7oqMvc+3cfJUfIQfx5yAuuXu6tAW/VZj2bjQI9iV6eJ9vW00pcCGVwvJWu3
1LIwL4uwHeH37orn0WclEIN766t3tscoa5Ex0tVuKLTyFLMQTptD+EMHqY7/Tx1zo9oGsAEhe6eL
1mQE3Dmh5lt4tRRo1giCDGYnpkbdsaY9LiI6d5F2QmEWk99BEvaa4YUjiDu+hUW8EeIJ7RYB373O
wP02DBLxMJ4l1JiKTK9LcjDbxpEponkNuCxbj8O+waLHuzkcYCmN5e/9l+NZYu9NSbWd98axwj1Y
i8IYliradP6SxGaoC9vmX0dOO7QV5Atln+GyS/OH9g/bF22Rg8rw27Xk1hO9tHW2l5pAmMeaR5qX
fciNnztGfO1hDGJiy0o3HEqlqxCCMC69GDKdkRnxP046cJTrA69dz06cbz8HSQiLTmvt+fRJnrmj
LYuw+yUMalPCOLU/DT4nrHBuoOrjDP3ARNCmH1vj9JiA/JeAKkELkUYB8lXJmQCCYDOeGp9k38f5
0FfjzRVp5vIV+q8GN9hpp4aWssI2qSYeYd9PvrDw//G90Ei7hZEcjioHxXf9oeZmD+jiBmLGQI9g
+wCSmkvp8/vZ0rUptnnjxLa/nBWjJSLFE4c45EWaP4GlqjJI++zE2ZSkAIuy7Q6G4HhR0MpJ2B0j
hRL0fjO9g1pGJKyvu7XgQ587HwygJ2Msj+zGab5sxGn2fDyT2QRzr+z1CGxC6DRUQwSwlIsBytUi
9ySDGr3liYPUyiZKbJFNi0Dhdclje/ZL+4hpi4P3JrG0cyCHFHgv7ZhKhIJ0C2a3/MyMcXJqlZBR
uUILh96CfXUNoTGibHXaYomPT+1S6c/a+2pb03pkmMDTUDmCUgbIf9pDS87qNkDWsP2d5ponU6bi
UHt+ci6J9OEar2gmgZxAFX+5fF7RF8nrS5dOBAt72rP1wZlJZzu2sItrZPkeLCLlQPhN+UmcDh9M
77NZ3tcigLnK45ktd8m9/mysk4A8/TkJkLTeBNZ4bzE/aWvDi+hhkwATZ9HYlcXVklXM2u+95SWp
OhSEuI5gyQa42vsUoo13zOHQBuVDmmeETjxMiWdKD9vZCn0bzms3WQrbHbjXK3kBTu/vUnUleNlo
k6dxAQHeHfIgszPGUfzLlSs6qqG/+ZUVp9LPSU+at2saY5aO+mOMMBiGftt+YgUz8zlcrXs4tFDo
z3Km9C2KTDQuqyu9VnyTc5qdOFOUCaqSIhV/cQfTDjSqagrvZWi7utL8/iRFLwrTA4olp+T5aw0+
QIiW7stkA1tOoGPXHvwr53bcq1qfZItwm1F/X+PWae2Vtj2Ts4poXKrYQ4QKu30iqgkChRdU0qy8
/l8oea98H5z8hq6UbnZJfcSnncoRZYpgUB8RH+tdHHsDXAbYHso8kJZmlDSvEXTaR6Uo146Jbl08
QiW6QjYQsRONBp1goYynZ97RMm5ffQA+1rUnvIl5jOOfAxupX4xQI6O/M9caYZ9KSpusANoxQg1G
5XQq9030cDxfYaOowl+uO674HdOxuA0dkkRdMdiqGUd9SDg4T47Lv5QwxOHhjSzuykcxNOKOBfrO
zs2HhNgVd5DWbckbKl8sXsDoEh6hefnQeNlJti2PwmRrqm1AEMgjyiPoZVJ30NE8Ycnclh1pbPJw
UXmi5G0kgvDnqfAeZADzIP28vFM/6KpSSde6x0wyniiW0kW1Hii1T6agNZfFuDyGgBHnIO49rvnA
pd/yAZkNIhU9aWDSBl/sdaTTIiq9iULt0RyihxJ/vjlpS96P46L3kByHOB60f1eXn9Y4rNICTNzV
CDxIHSpJVJyWq5ZrWdLdttLJH3nV9ibr1Ov8nbp8p2NMuD0lVP1TVxq+nfxG8IgsZ0L8k5lJjmdi
1JO2g6G2EuxvaLIJGxKzX0jH//7njtBMGyf40aBZBzmiiBI8YvjlkRCWoasHdSmmq01rzDDbo0tn
zcTjpelsMJeahOmikZ0MJbuil2/CWL37QufAwSB1rwsdLPNFYjZbabxRzJwBUsg13voZKJ0cj9uR
qic9qCKYNJp3EmeFVifhfsrPLfX8JvdFfkFzHtmcC+n0okyzdqZWQ2hbHA9rcFYskem0v9F/hSCS
/+qd4vxWj5ZBnmZbo1hZif/Sryb2xygB8VwP6jJv4btZuR+4UsivslbM1kzIRViS5ux3nrFlJ40o
MApubVfaHXLVJqg+/xymKw4g8CyY4Fv/zDENAXOObjDLsdTbcjv+PmjFHA+hLhSr8hxJ7lLtJEAb
l5yNuEPw+qPhZwL1A0pCr4iHJP+kVDgjzwmAr1IVGtgdXivyyWhVbaz/+3e6qudL2BKzI+KE0nYd
mNvBm5HoMvG8xa4t0C3Hmkax9qIG0eNUvZYrfxaEljnfvGLLZYF2aEFVy0hj4aA+jVG0sbDg7W1h
fYU5b409KW5QBkAeujHhcdHhLMYpCikLr6kS0EUzrpu1KeKIXePE6WTDJ3E2HJq/TXhRFlcLC9Yb
LpbrEptrj43k77lrHxCkfq4nfE+E468BSQgdQM39yIZzZvCYPcIaS6dhfIVaiEhqBpFzI7266s1B
vGZ0om8wNSR7dMrrdTrvmKcSTJlv2QLj7qx5bNppVy2eB63R8eJ9bAo4QlpHi841ghYWjTZjT3w9
w0aN2AHj3CCq7fKs5PKzmGuogSdrId2UaFjkPBdmjxPt+FwBmVhdLYAZcflX6y9sd/qdu9UtOQAw
wVS+2k0Bn3mSG5vhANNwwED56gmAgH3mmL8Tt6BWQTITxm5H7hgiIp+aCYcBGjynou23QXULYAM/
j7da04Bf5QzJLJo/Mpyc9swfKDWjSzachmo63/uBNzsJGUX7iQTQll+KZwQ/yNG+0knvabh9635Z
dbB0YtZvllrfwICLSJmahmz+FJ9K7lZKvLTl2PIhpNvkavx9N7vKyzazY3otMWtcRl5A8YCdJ3Uq
YfpjyCa5sgSBwyIRuXB6I0pl20MwDlXjz7nsGPlSfq/CSKt4y7vL4lwdlVfXKvPVvRmocczwkCr5
NS0iOvRA7FTKWvglEn8f37S2a3+a36EXNxS5l1j2UrzpDYZDvMgmFTChcCbAsO8eGvtJdhV7QGq8
Wnl/jtVYNgzJxrTfIcnQ76pXS16Pv5KGVWQswz761Dw+5mLaj+u8CrpT+BPkzjwG4t//V53ncCVS
Y0pOh8IjE4ihTSx/I8fSzwTp2TGYDccGgC/2RH8xR6lVjMlexK55Ga7gx4/8GUyDFUc7tsnAvmJY
J0d5sIZFnp4rtagbD2L7PNh68d920mOWAL/WGyJaLL7u0eUvL9qrVi7ha+CXyrmayOKItg8FXPpY
m632FhHcmECC6YfAgcOJPaTLJSqDOccNGBw7eJe40DwPkl3UT3Z/Y/hWxMHXMHqFBMNGrTSw5i5e
uTSIbCDEinmBcMvo2nM0/BbIDaCS/+n2cFQ4xvnAzY+71TyhK0858rhlG+nE/8AiLsKwYP893iii
S+985cRiAvneUyVhvtyqEMQiR7is3lI3Y9V2puMP9nJeaHDgX0iMWhLJJL2v72UMWQxVD4KNA07C
5EegfuefeB/gW2D1o6M0lRGkevca/Xyiwllgh3s0LRxdVKNGI8op02/tqQUWAas8B3st8d30tCQP
BMS03xBdAQ/EmJyKHCwCKtfXjIbp8s8Rq6AASPVNhzUyahdcinnfEUwO1yTsINWvSyu0kin6fpXl
Bw9eHDE5VJa3sp0uY/R3mrSsUm5Bvj0f0JNHvQqzrG78GHYMOG2cBHANOQiLY9SFmVbe3SqTpu/m
mSIs/SXyUizjURjjR7XY2wzbGz7IyRWcNDWwoMK8ZxaloAMO4t7rHo/6uCkCq2CsmG2s/bCCmDaH
QwWHEnWumHx4/NaBwgZ83/yT37/7jMXUU76FDEgCeJS5tyPK4UoNtPxXt+D9q1TY1xc5RX7SzZT1
PtgWdhht6caR8VJbzcEDG/Poi+OPf5dZBQi9G0eoJDpGIEm1w1IxMcEyOYOLoifwn6JfnX8yhcm0
Fl8JBaJ2RV+Skx35udIbfKHE4HQXHS2Md5KbSWl6B+ahPAAfi9kaFNj5WRr9q35saXb2ttYZeziO
Bu6En2q3ucVTJQdmOzDmQFcQnzgnhA3MEQ8v6m6TyQl6A6V+AZTxgoBDSBENhrbNOXWe0LLGuPVY
d/51Gze/oYLOHpD0JyezbBJetsMm1WdO2b77iLAPzh4Pz94Mp0z7BNhN+LjFwvfbyYkDG6FZh3U6
e0iw6+NWhx1Rp5DHzeL0Zmfhb+WMrJYO7z3dsYgdI3F/LhBDoPvaOgWGtaoFQRUXXMeFUJn7Q1SE
fHz+NnWZi/Pc3wAnwbeGJXcRmp4nI/ouAL6C6ibzgWXmuB5ggnrSeUhHTxh+lMiCvx0DS9nfxuW6
7lj9ff/ZerxSDDLR6Qto49q3z6cFNrepYaxmcZwxDmS/d7Td1LOlDKERMtNvYuWKdo/lR+azFmll
v62Ejie0gu1KUtkmgCqEhTZ8b9vk1elqxaTb3NRmyY+Jxf45PofbUZZX9n8hPsAxRbSGtQTcuaAD
/6jeaYddPd4PAm2aWsbVnWErR3IgoAh6w0Q+xiPOtN28094YeKMcKbIww0Sqtf7BaI0rJJU3Cxl7
KUQwLPg6tpi0yqla0dWpgvFepXwaJQ+i4Em5giSqJl3Tv/rzZu6VYugznQ1PRCmh0DU+Ba2yFVYF
ece89pDQi+Y5CYgygfaHevJ819x8FxaBftqfDDUYm1k2GgR0MD6YfQYuNp6M9jTQ+c8siuYowzwa
jHjuPljREAiWefBxq8esbivxz/uocaDdeKgGVYdYDbHrsb9MuSzVOPHGlztLc+uLqEH4bOc11Q6X
wem2zsHKcIDduQHpiWeh44TjPWPTxZvysW9Qph/yu43sMD6HuL8HM6Rbou/A5WmCGy/swmPNA/1Y
d0pypW5aJkG/jX1bbhofXPz45zycTWSAaMe3K7iJlBhiVckCpByVaIh5kEoKB5hNDYmcfos3zOvH
stqgA0Oj0NloRnjX5n3x9hqIOv5y6pey7+ulBsq+btN4qVWSCcnNp2q+6X9PqfCJF6Cd7Axi+DeS
T2LuG1fQY6reTqTK4AXaKFtweLc+iiiLQ810U5BE4ae5fkNOpNNruwgAm72YnG1xmTc43t1De26B
6/JMCsfE6LH1bmkmXquttnC0vtWyGu8P/fmO9AHeRQ98/9pjkcUuHXSixK/6r4R0+w0GKGmvcuoQ
ae308kF6uVD+RW0shOUv0HFIjdqXn+XpF2sKp6Br1zusvnoMiSpsHaqPesCGkzi2p3/kBU/ib60e
kNvXfAljU8DD+TJeMxtQhnTkpNgiUuOIKFZfjRjJakg1d815Jua+DX6LsSQV9eo/GA/Ea9ArFrfr
sn+0l9fSEjc27rLUco0IVY1y9PW2Fuh8nza9/G0Y/mm2bjmZK/QagAGpG9gG5Xza9qcYcpeLty/D
iC6PJ4u3Ruod1koWyr9Ofe6ST9mQVo3xBcZ1CAVzmJLQPGroIr/PyZfxKDnY49VzoKa2sCExKkRr
pFTwiZEnsiDn+oatOvaPKkZg700O7aJOFuZi9wla3JUKlJURhEPsVewyde+CIX1g7plfIDKAj6pl
vDWRypnKmPb6/7dJhzhY1fldwE6fUr7U1Zx2x6EayaJipoDkCErdAaC48OYuDFGWfWfr9r4N2url
Dt2b5ETgLfDLPKU7P8Xy2QxA++jHaVt9D5Ys/Y5k8eGgCPlffKpAzKzewQ//43MM8/fK4kgNr5Fm
3VDP3lgpqkJ/hDNSUOo9Nosu4uKtEof1IeXfDx9QYxqexhmqIqoPYZZ82bQLTOC1wFJ8OTdt3fOi
ZuL9AphlzBMM0gQI+8qpTNydoDcZmKxzKpJldTtNQNjM/aJFUITxiIbgy7bGK53kMhg0y1aU2Oei
egp3/Tp0kaoFE83eX+Bq18a8Du5kVfpBGRWIlgz/d0TXBJqG+JHqk62Jf5vKbeEAW9hfsJoUCSdK
h6qXGf72oCG87CatkslccpxVzFcHCNLjTvp/Zujs4+T9D9OJEOKkBwVds8bhDrVRjHGsDGJv1Uyl
2fCDfEyCLvzZRZMN0LtJm70UqFOVM0iJQldPZVAo6Giup4prC/4ZqxRzP2R3dUhAZE2qpNdUILPp
H2T/KsISP1bDICuF6RHYANpRKiMU+nezyR0nYcNOfL06+uxJOcRdK61KezOe9goeUHso2DQ4hZAY
/4K2M2H+pR5AnwXJOtSxV28ZrXcze35FLSEIAgt2fCQ9FzHS84mNQCUBTasf2lbxyKqfH/o4F0wz
dfkd1wlFb/xc7nVrNXzP5pfe2Lu3pPTNnMarhd8bkglLb5RkPRm5JftcNqekLIJRxygrWWEn2I9v
0ZMPV2ECMf/r2tRKcmIrvUNLieo+pzczI3sLUV2Cs//ylWcKl+gXky51RhTgT7jgNPlhOb7WNeDq
KNBSvIU2T8PWMhGBhe3NG6z+1Ek1VmIxmBWzbfatukZ+iRw1VZQD3rQN2rTBBn+g2rrh3dq8zY36
jFF7Qejk3+OtYLAGqraWNz51hAesmaFA36Y/bvu0VN7LDmSHAUq13gX/3qHalFkNp2O3ytGQew0a
tJ5FA22GScXCKMCzlBSSWfcb++UPMScCdShYsuPC2gY4mnCzd5ut0qJE9PAX680qxnMbUhkaTwPw
pDwOjdazRv6kjVC7K4xBkO+YnbpAt5pddhaEQJ5wYuKRIxUWnzLbww3+nckPBL9TEGTeOm36b2EC
MCwGbFzsvqDYQdi/kd/FZGDAFkRo94IcROCB972bisda7aSx3i1daHBewLX/8pCgC50BAt5Did8a
OV4CegoqQiLzlSK0//XwbkZ1I8SnpkrqaSWpsJnYpIAUkNr8byUISBek7Wb3xW4vn+oTnt9tdZMg
s+4NUc8oDZyN+NrWVNiH8gUxmMOozvar3EmkqTeNADZy0iaIqdi7zUO70dBG+gLkFlNDjlGcGfme
PN2kFSS191SGIrkwJcWt+Tmr+2mW0EITP6F8glxrrWadcH+f9tS1KvStHvqJzIX5VGDI61zepoZ5
pmdIuEKgMhIq19sFZYYhrqojBnsIkrQNKIUkP3vfOX5yhNjhfsdg5BkOjUWca9H0frx6CIbuz1JS
aEqEa2nlN5AsV04FsE2H/KNM/g4NzD4xOJEbKiHOQCbkSpn4p015cktyyAS/2ork0qfWnJQTWQvL
yfD+SchwrnQ5BTs09ZMC5Gd8t97JTJBN48ivWf5hbOXSmGYb+NFouXpuO/YApiwGQkF51TuHKFHj
9zblNSmQTIDqi0RNbQH4kLltMMAjUK0Mu4UtsN70UrY7c5tlEipnCTDY234UC6U6/OfKhWUqsKp1
8duN2Xc3pGkdss9XLrqaG/yfd4mX4kSHUFCoAiZZxNVX5SbRM7YGS72+Tgu012R8Fnra+IaQG6yo
2nAQp+mO2jrhvkPsKf6g7aYtS9WcEFg5UfXkW/F5M0MDlSGLG5+g0rUkQ1Fwpw3sdg+AVOnmXOHr
+RH9ds8ZbHzJu+elPkxSmA1q+fuN1Lu6gCEs48lkyY3ZKkbc/rpXrGCVFRbE1eUwJPAw3P/B5wCb
dLPF6zJGcMxNNnZ2FoKNco4BFQhDOKKKq5jrFACmUYv1aDegU7AWcjWFuzjQokMbNPsz1ihomUsk
63PrM5A2+wbjh8IBUuPMZYcFfha2tBxmyVVfKrDyoykQ0MQnmkbPyTMV+Tf1ev6ApagzvanmThCM
3y3uOpMmFD6FxVxU+QKrVSKXv3OZjRoCGbZW1SAKjoXRTn1cfCWZpCed6tb5/ESQWu8pj7hpE3M2
7+wWtJ7Ud5Vicb3X4SKTUgjTfp5e1g53R6kBy2IH1BwQUs+UIHq04aaNKiLCFkCdmILiebkQc2yR
sxJ2fj7Q0lymLcALQxW9fX/zq5Qy5A3XEEP/XZcPHpX/zs4oyN3JTUfbGEdFjXWqo7aHB+Tkitp/
1UWefWyBQblU20YHfDyWt0D79OjIpKKMgCBVOx3Y285Dw4QOyvTnMHmTtlFWy+osugNFob7rdMBV
GDtFlC+d7ldcv3mw0PoXmioy2uUTNfZjIzr89xBFVV6Nw2X5EbeRYWGV3PMO3b837kWrmDKgrDcz
KOsWVxabV6W3T74S7V3OkQ7Kt4VpkCY+D0oPf3GoA+g27emJsCiQrte/sfTVTJAlaxaaKKrgDF4S
bw6oJGmmpgtUE6BZbhUu5Hrz5gVC8gzbmkNpkuijNyGG3/uYGi0Bg/hRJ/ZJ2vDrPUoQZ8he4gBi
wPCnV8FvcARkuDveF/bdU0PoaAAp3GD3Z0uL2reUhIRdGPzPeFzDaYa1ecV/ZswoPO0nyeI9gxJ0
njmQMDC7CCieWSP3DtMv5q6oWglTOt7cB5xjFhvTfcfoC/92OrGt7GDUvHzaBUrG2jnsGQiYnAbt
NgOhOkpLBJ7sXGLM9eGWqTXxziyFXS8CVlepolIPSvtrrcny0FEzvEnobkB4vNHnJlI6RVC+ZoGy
jMM3pquYg3GngjnXyiTKJh1jnqp/fDg5qkXyqbzidQNqW3IHnaX2tV2FPNRp+nS03Y/xe6fOvTix
Kdzgxpq8Iuel8ZtGHfXbpCCwZktlK3lFi3At1sWQfTLz2G7h7z/esyG6dpcwSnUKRjohWr7RDBEs
M6bvRzprGqchf/cBahTR324QgSg1uEXW8CovHbMCm0lRFA70GsfDhkDHVN33OzFK6DM0D3pmyBQY
QTUY2zDixz6gUKJRKxph4STEMKjQOOp+s6pkio6dYGmiaALRxnsf2ViOIJirVBdU0xiqeHGQx7t/
pJThBijIRmk8KNs3A02Rqy+33uwzGm9t8CMwBxviN207IvpAN6SMHba3vx8RG51oV6CedQ5zbvlZ
skCqwtNNFj9Bcd0rCreqzFrLEtqy9AgBPcFu5kyxSPDBTPgxAlcaMAoEQAlfUcw8a426btnhGqXm
9XwuailW7xV8UN4yKZfSteTDoa3avKjjDbZ1xVPK+N3NkLwU/8rT0rCRBUxuvjEZU+9qmujB8+LG
UhS4pcz3CYFV1ZOgBxsd+eTy3aseZ1CGc7OqCIblw7J8IVGnag/dQf2vz0hfZiFm2VxgEg7o1bbu
VALgafmqG24lglIWHOxqEzzLjHfCQtKYqX0DjmGwD0AQXaEyAX7C4XfXn3v4uvxyzGi2U8Ke6p0t
DU9MrXTvJXZMrm0Zz5yBj73mpvlzUJfmA3AS5dm4C1BRNgzg5R3MQFok3UhFTgzXzKVZMOKa7zS2
7heEkgPB8K61/BQI0CrVdwX0RpyA5irny3rlt5NeBL1RVD0Ga0s2kFCA0t+WdBqbA8G3sbUGjOKZ
DIoykDzsWsd2GOlLrB6Hm0K8/JbccsjVMv4Jhpo0IUd9aQ3uu9OMQJ8XcdoTs9yH8xy45+dKrebQ
8fsn3Siy5aXEzyZFuLnsIJYsKwXZWPGEg5lKNfJc95+lNFJUfzAITR33oyzdnNgNW2VihNPvc2ri
I3Rrc3x+8bscmTUZKKy+7qynojWA7zTAdkdW0dlmbtmlWqMpzCS+538taT16D2eeOo6FGiPd3rYO
hrrg344e3TxwZ1xoxkMkPwbX0k3NLskAuuP0VXmTP7hkx2rzgPqgcJxbKjxFEqVOFvSQkO4K3atl
yUwir8OPrBLASs37oiJnfvnFazPG0kcID81Dbrm59foptU8rbDQx6PtFTHukyWeR7cqPfovybYvF
z6z5bwyVa+tWy/jHG6SjHnAWnuBi4cif3ZYf+fc1ufjiAU3Fk4J+c9v+esqg6n6AcpTzgTkdvu09
CMKbMMCLdzVOEygwGvKHr4BKREnJfp45PCg5vsu2ns+tUBY/K/7qfzlyhrc2bHhEpXMEfL9Bx2QV
GhOkUivjCuhEaGyQM3HT6uE88Kw8qdkXvhvLsztsvPaofPEHK6AGEjWOX6Iex098xsj/MbesPfO8
VfeLgDpV2VyjnwMYWfR35Hv16zP1NU1NzzOqlMvnMOBK19KSnTsXaVHIPoY9wGYbb4r4AAErLNyg
N2jkyM+HeL7MyBK/NSjkZITf6elwyXOU0ojgRmwUONLKbBMbOYvKOq5peIrvN57eTQqo2SLCfCXQ
B3jo+gvWuPKNjMpVPoWlQicO+aBo+REYEbgmGSSxo+WgJld+VLr3ikwbAYu6NfrYi1E9gCZL2AEF
wit0H7a7JkzosAW9SPdnNUvZuFgQPSRrlXo8buGv7Vlzw7bf7pNFQ1lDYCf/+9AG7VV2htFj+ZyY
VnUaBTRnDWmF6HVMIb5w3npqIdWj/LwpJM7m2S0643rfqJ9ELzrul5M0eKt/u+Oj3F+tWIpAKMIV
mH8ql2AMd1f3oqeL7fwUyW6tjHNqPdwu6PwO8MpH11nGEawyiVx7lkEwkP8mGsAxMb9kofktuAto
IJoNjoMY/LsaO5hC+gXVILVjxbr0frAbWUQPJN170KGkfAAfmCBMg1iHjbM8+7ZoTm6n4HLMe9BA
e3b87Pw2xq0m6KlFXYDx4FLxehDPtuRhjBkeSrgUKoiWa8f4IkVoLYpkgcPGzjVqbGioTvoHrye9
BjIffaxMNbzuMIY4lumpxsPwS89+QeY4uVL+2YAoBHcsbGajYRM9i/H0yKNVQ1Y3Ko6q/vWSBomp
aDTwFSz4zbwCZ42n2NtqtzmUh8XR5xv8/JZJPV6o+kQKDtkGfc8b1tygzqseMdEFFSo4AW6m8Rgv
JbgbN+5JoBNAtaGsyoPwaVuOX0UbEQYw2pnSTbaRzEJDx+8qM9MplN5JNte+7Qrr8Fb/x3+iynFG
gDkpq2Mt8PoRFDdxCJqNpgNQK/ouDwQTgLw4zkuS2GUrOi9s9rqMQZ84u53RoPrwrmreO2QbMelE
GyIVdntIpQOsGZMk2zvE4EIke/lkTQll/ZePNfU6sLj2hori/sAeaP9NKJl8Iek6Jys8tDuFTrBs
83SqMh0nMZnrEDSgm03yLRxwPbX0f943HO6Y5yixA5qWzNyV5ssO/asroT0LOt5hRUnJEF69t1QV
ZuSlztGV1Ao7V6yt3iCRsMAiAYEwtdAr+Wg4SOh4rfn56vZJ97lM2+6Az2M+pkuyyl0BXwbyJ8Yu
M82IGeRlFF8aAHYOK0fFWoGmjBq83GXR63vcFNd1ZQ/jXoFzg1zXUk9s8dYLN6CTPlt69W+/1iZo
HtxxV9tiW2u2FtqoD3rouGP4XsBMEbVG/i2roCE5Dwv4Gmp+JOrTrQGOi5zprm7Mm1ZqIhsZQ9AF
HcP13pHrk+/Hef4omUDKypKV8n/cW00Ok3yFtsndsnZpT0PeiRuElkGFrRp5CLXrolmAv7YX/C/u
1iSwPXr8qgUsosVgvUb2cbeU33OjleMyN3qXq60xNGu61prJ2MT0wd/gDt/RnE7OKmMDftQbfl2Z
UIZMFkhLEU0AlHIn7Tth5Y7co7EuRX7nyDNV7vtGMjjSwZTibvTZzfu74MB5Kri1mhKKPIHDIPtk
SapIEcEtukwhXwW7DS7pWbZ7tkfMqS1ztWWchkKwS6gpCmuCtZL6FeDw29whD220+s8n3NJE6OSV
71yT/Y2i2Sjd1im2V5uTKEdQJGILCltAFXw3p++I4dCzq4mp+su3LUjR+OMOIStGW2I0azpP0/+m
vDAZn8xvmOV1fvxXJU1w62iAvqA2EVVgoFBszKehcWRS83cogKeleAzfjQptouU55Ta2iG2rb3nS
JX9QRPFTDKeAnB8Q0f4n/CJCqljJzS9S7hoWIDqN/S07r20x5nGBwx3TJjwEESIBtf7me7NtNPPQ
INqNn1MuD613aeLyPThbXt9MP/T3lQMo14xn7+QAu+mBpGn8JbhcAJu0TTraYmmPSj2liMpvif+7
rcK9r4URpUKlaH/13Upyf9brY84ILLg+zzr9LHTepgiM8WKUJ09dQs/FJ2uXNyVvOSgkBP0ZXt/s
9Z+MHnBOGpRil/KPRbDk5hy705IQoMchLzbxagKLMHfE7WGEFvZrsLMM2XVrpJceYKXDQnpmop3t
SwP0y2f29xg0CBqdfd7XiH2JvWOYRqdBgG0oUf3mB8jDD19ahWh5LTuVveRfjlrQ4Wf7ZVelEgr6
Sp9bNG8plcTRDg5cnf9Vb1+2Zhs9FPh/v1M/4/y4i2ZgSsJXPWUrZrnthjB2Co+41a+ZDQ6RzZA8
GWFCSGgLSWXVdxDRoEcz8sq8XAMHCTER5EtAyzVobEv8xvkrjQjK7iNbcjVy4RNa4FksbcXUjaT/
3rLS83RpFG9CDJQMIiHq90xpjO4RKfhivZb7keUJotsC9CwI63QupBqaYIKn3wxqGtew9kMlTOSH
vKc5xYAU8p3wBGjKCTo18t1Z2a0MZ+D8LqglBE/NRa47rAF2QOt2MX7LGRKwr09UA5IeAG2E0vs3
dMAS5UAW3dgZPIeWLP60LuSl9fGjmuH0ENjEZhU7JEbYseori9+8ByIjcJj7WfLdtM9j8JpnkJZG
RNRp4Qa+wdVUgorVIm8i20RK1LNMJM2LsqC5PV66wsShjsK/Rb5cd7tThgna1rYMnGDoIrbIj4Ok
6QWpR2Jote6AoQQNY+9ezafUIC9FT+4OPxieCTxuwNZNlO5ng8t2No0QIC0Fi0SUFOnFR5M3tEBn
bc2B1ondtQg/h+ru0NQbAlJOyd41bQcuYEtnSJIpv1DjZk3nW9In+ZfAyKDOhS63+EwHxjkEWbsu
VDIs3aFypcJjjzOC0+CqsD8OWOBjmx8xgNNOVmf2sWYCjh4OzN5aRmIvLZ4bUqJXlrvBiRjevz6G
RIFZzmW3GfratBrrWa3toscxO3ITAoaBjisgD5rpA1S68m7sKehC3MXbw37xXLlrjHQiCiUqE2vN
+fpkVjki2rIiveZjxH2JQJChtcDx60JxL87IBjzYFZBlWWF4B0dqWe4XppymBL+0hyhV2I8XToR/
b3U0Gm1o16GpR5pWvF4KTp53SVW9BPoonrrqTH1425SYckNsYTQ+WnlOm/Ja04l3XYjHZYpQoL2l
29ZIi1LERufhz0iqtxnHabC7fuvCgh6EzcrOeK5heOoKF9k9OPDoROY3fAOMa2ZLdusr9VnJaXGm
56JJ9FHGzB7Pu6ZC4j+w5RTZQkNfV4T0l1ykZD7NRjguRA+nYBUukH0GSfKy+/9B4VxFPfU3Fg4U
sKAt2lWbq307ateDf1gRHigbcIRxLBfPrMEj6sOHnEsBHdsXZskrwYKW+jP9gxkCOEVtdczXsmdL
l0f+3zCUXCkhQxav5UoQu7Rcu7uCgGTO5vWQ38HpMvWObdSHO8uq1lZPCoE7opuIx+Ke0VYaTkli
p4c9QPcy3zynVihEGz9j8B7fEudNZEK5hkKzgLPkztE5iLGKS602/N8NQsts8eA4vRZu6IKkfgzB
fRJlMjXodOAJKmQgQtHzFp/XuLsVo6E/w30a6YOjds3GCvgUhIBqSn/iVLFK/MRqAnVgcyIsjkK+
xXVZnicctQtmESpcdPuE5YWcvnRnL+P957tlrEhV3Svng/U9RdFBzVgN5ZnW4zB1cBpkwbJzKNf+
EG2jWsK7uIZusoY2O54rIaFLZJzm3qi71WF8CpBD5GtzCg9atUe0i87Mq6CkDcW2g3CrgHoSSlMN
DX0qFO/2z3PGCWUWqEaiGDYTFgRcFFGkfEikL5F/oYtqzlnh0Jks4EY+VKM8TlkIN7QDEzhZAcp/
JIqRgTKOCHzj3WaY7YwdVMNJLjaURfMawGvayeNFWp6NnokwVF85/2XNDd3JDaj0pQGY+xzLoUOI
GDKoBdxlFHjukrKcMj5qyPvBTZktdXmIpM7ranR9dduBNDj/Ci2ep/f4K0/+b89+/8zK/lNEJrYK
imK8k66RsiImy0NBWg9yznGFKhNAJGm5jxQxiLgQLbQWyJEVKxM4/hgmpOyRJCKu6063um751qVL
ukc9raIyHrMgeVxRS069frOmumSMYJJGFiVsKvSDY3jb9V3IhGH2isqM2TXGXv4ooNCxmWNs5D9M
5SY2sCggKN+BZTmzSfR4RCqyBJrcOE7RTqlgf9ME+0o1crXqEM/SCWTl8SK4KPCW6Q+gs/HwhmIR
3nxbI7LJKNJzLwDdriKEzhExDOkKZK7IGiAxoJNN2uCj0cXlMFhkqxAaT6Il5D/COkQ5rDaVK97x
msBr85xkkjsGzO/9S6BBZX0Bq1ru1MJIpwPPhdmVRpaV0vmhiL3lvriYlBVaXILBU04UZbtIZrfc
TZbp4xTT6/C3xKsuakyowhhHjwjTyr4RGNmSBxx6/Y1RmYPtELY6jYwt1pxj0I/3Ex3utsfKRgKV
igQmfelNArtzPFH4/fUqMRQk+eBp68hXDdWlQuwUhAwUiROtBrdP3H2BpUetBF189WBjV3eazqW5
LMeTMXnAvEHsTpqc5V27zXXFR/ftE0RBV3nh5m6u/1xlwQJomTWgsp3YtPtb7uvgAS40fUlaymtP
KqDYrlsJMGErh934RDk1mp/vKZmUG7+fRyg6o6e+sHP+X7VbrrRzbQs6hltTZmxjyRjZFNtR1caD
fJ5zptOHpGiIuNr8bBjpxxNSCRHJoOm4fYGGVqnv7ibFSInVStvXEZ2Q5VzpHOCzCwvbV2FeUEXF
o+dE2HxzJoiM7+LgFGr1nZ5BtOp2rPSsK1yXDAjjaob3F3AptD5INrQtZNmsmyWH3nCNEWwoAZx8
WgZPMw3kU+FPFsS8zAlz6L45SW/++Nb2wORvtf9Ynj0wwVZL48cvRWsUN0Dqg2hXWxRqd8RTam1B
t2gYJ+zpBeB+OXzfrUqqmMJlTVJQ+NoKYxnzjDwsJkwuoj9FQMFUhhALHJ3pdBEHVRBnvIUJQ60a
NPUFGiY8xEveyHFdqRgFx+tjYAPs6yO0w9wFxyBD0WXRJx9UO7KvHDx9OgejKMle2je9sxR7BCxq
74/3McJ9JmOkDQ73Rs4VfhKCjTW25GKqFCaAzf+l4HCghdn1SXl9MOebeaxJ0U5laBtBWUDxx/50
EJwaoJqQoMW1xdDo3yufxemfixAqNj9Y/7IMEweJsyEvCsQ435WvPRn8AKV06JOfRJDojhtQz5nO
2ceDXIBY2TdjWMfbsYIlLnJ90JicZpjYYGbn9cyqRKa/Mr41Q9y4r00rU14/fFfU8FavavHpHqZ4
xVF9+3kbCdVQT83wb9HZ6NufOKKcl66dRrFR4bl27TJE4Cd525kUTZgcVhLZqzadPn45Lf/aEUvB
fQILxjLVojSP3Nyf2lQpHsxqMj8OIXW4/zDcYdOxkpmTNQ4rh+wObBUPWI0GGIS2+Dfnb/M+WHbP
Vc0TERBh71UG0O/1HrJB3yvOmJBS8ojg6NCxilT8gPZLXLZmMd57CaBV6m3TrvKzE/JhqP+CL59z
kVXzmlkP5doKRqVCp+9AWLqXNBiP295yJcNOV6ruhM0Knkg+cD97sgNBDSDc4fqVJ6Ws88d+jhYI
0e0gypKOz/2SgHvRX9H/ZrLj8JZ94KUxkMe5gMo7LFmQyFFLUcM82/ezT83B6iTz9fsg5LwFMDgn
mhgh8DLbgdP1pn6ZBE4z+ACxGVgKN4jydU4pHjPCnoUetEKIcDHf6oVVRnEg39l9MV43CQ2cqlji
AnDD5zDlaFsFp+QAIVlvGiVE8miuwZ0RmyHdh3nSNs+Hba8fk78O6lgpHPVW39QQAwy/kGAf4Hsk
kZfq9mTcbeuaPrap0sOe/iNOqQjQr9iSh51MplDH9TuoAn2orybewllMIK3P61DzvFKPLx4Oggud
a8q7iE7S0DLMJa1Ua/JK/11SU5E5KGFIZ3lEJwAtwWZU51co5/rBHokAbQ6Jb52A2Mp1X4zYU11e
BIAtjofthfvtgEy4cQGj5eKiysf6S4GLdKrs/FEvXXC/NsjF7/7Xg+NZVsyemMXR/5CW2u+Maax0
XpzXOOmh1jOoYH3B4/AZ0jlGl6BIcuvX/A18JAzJtmE/U2xahkNGsLUGkWBxvlD39OOPl18KLRBN
wByPM/i4GDjmHdkdz4PS6Budffh6BtMKH/KFDIz0xtvKyvgfnfX2plCDcifk0sfz/Q+iQtlbAVx0
pXPiSMQBLkgFB2GC5fur+PtoSrGkYE6KxWaOXNZORwgVtJBvnTm+YxTQk8rOI91EpM606Z0q74oT
eQE/Dbyo/PMLPr+5sNGlPYyDVYjMSOwNtnL1mcL/DpkWMFl+NVmyA+IGYet+ruUsa8Q80Ghw8xRF
30bDMn+QJ9cL47LNhAy6/LAeqbfLl+MdHWYK72eKGKXTFLbkHVsORmcN9/tIMvA3LhpMvV+T6FYZ
PFOKQMJM4sqZA/+n5ula9zCCK0bdpCySln3GOMQZblsDfu40aT6FFmCXWuiL1mFXONDzQJAOnoU0
mxAO8bXjEUMrczFdQS07QPK3atPMtiIvXmjepD5HuuI6oSZWAsiKfJ8y+7DJmDJ6U4dghM328gqj
jptPwoieEnsPZFxQstNuoHKfIKgW+fmSm8fVMYbbneMsl7CEKvDS/9kUZ5cNZJwK3USgMlWKpHvc
28HY2IrtcQC9SHc6CZ5iggL9tAQ3fFel1wes3O48vyWTrv+23MraxcwuQIciWq4zHeadz8TEoWVh
eZH4LMKfvBdh1gxspVQZJXRREr+VSld7DcJl0lc0Rri+5i6PZkS60IomMMHl0tmi57/IC1nPp9PQ
RsHhsNKD55tn4izbwEryRZqYzWKy7hgaob8Fcp892LgqZ50SgW9GTEbvpHBOXXcDF+POko1ekt7V
8jP0AcA8H22VqFfrol6FQuRiKtGMK20QmWUIQtgCRabL25IsjJQBiC1cFuhTJ/u3IGGv93ZhRePq
FGgPyXG6U9qLhz0fWo+XfUBr2+SLvrnqm2YXV4Yv98pmJGoeILM+QSvnB6/2b8PXRMhysIQQ38mZ
k5T2cyIkE1sH9aMtY2dj83fA4NsQjbxO8VGn6Y2U+Kzt/zJ66ixdi5VBv07XJMWwex0sjmoDi3IO
SsbDyw7KXTm6iAlxHFlsuskECFNLL0I/TTKX8ZKkea8V0St3UsRCl8rTvumSp0lBH1gVK+uey8U1
PPiK10EkQ4eOULrbL4oP0bG5PloOPCPSLojEcXJwRaWNYDYdKLvggXzvl8PWFrQJgCYnjnsgHOMx
rggkzU1VTQVi0I5JXm4Atskpyah2kK4mpMKKb3FLdj+zey/EPaVpNwNkh0g/OCPjKRT8vWDIEORI
HDZXBRjDgyN4hyHW2z2Xmzq8op38X5rQBqTw25L/iGM94TMfR2jyfCwqLLIibGTW/umwpoxsXKGs
c2gIYOOpyi2KgOjzemOmVMNB+bPHaS2VQZDo4bILV/RRQ6gOIg4MHSuEllclbuJCIwrbzidXIP5Y
IM5h0UM6/bqaHXaglzZptL+A8LIEjlD4YtoEfviqPsX/ivMMHbkGZTBJBWgGCE95ubypMQ6T+z0c
/H6Voy2o8ai8n2482hTz8+9ceE6M8PoNtGBD6iFSlt6TTapEvM13KLd/AnwCUvtP75N+ODlVvxFm
kYxphvaOO734CTLC036CKEqUFg3piiZdo1A70magz3Vr527u9EHzAMSjiiqXXDE9CxT1J64sYoNH
20OL1U0TNgx06DHR1vGlKNO8oWARf6SUDysWzNwcKT8+JWEdDR4W2napytTexeqorwszhN1cxja4
4LFrwrM3QbW+wZLcFKL7eV8dnEYMHtz/D8SMJ7LybXVAdlxHDZgNLQBjN2R3W6mOrr3j78ZS5n3A
aqV9lesVpPB01Jb/3hMK8AwSPTw/4VovIpaswwv7IHhE3XORRf1O7AgQVuC7y7T/k+OCXpk2Vi4E
35r2HjSNFoa15dY+gnjOjFyRbxY6y+AQH1ri2xwGumeI3IEUNS+iiLvowZwcnLFDH+g23sKy/8i9
mN1bXqtVuOzoV+aVx+WT+7hZZwEf9vFIqwgAClHMQabiqSRH8hdgE6Y+sM6VD7Fc+hRTW95ylXd4
gPQxWkX/tiL0xZkVusoMwerqeOejz02DAt9xvXAfGoZFRNfB8Rc/clLY1++CRnGde2D3fO5XAoDx
JAJHIDNPox+Dlnk449eG5fmxF53Ll6Tv8a+FP+WgrynO2AI8Mp8teuyBAoyG4a2MFFg0N45ySsuH
OCcpC5fdgtavE9b6+p89bqLkfjWNkhjeQsfAvgy5O8NxbkPTKIZbmqIsm0o3rP9gPD94Gs38YEw6
h0PwPPnxSvBChL/CnKU4j1LnvebIU1sr5E1twYUpWNYT2aOWpN5DtKYtWc+2CQSwSe2HGOpD/VjT
Nw5Q8/6odg4+Ry4pUAb2C85R7G5150+5iXbvIlwTYrYZbu/Zcsd4kvoklJfXjZ7UFY+OwLi//o0m
dC/2eDDoleZbSP/dUIq+hrBi9YUf6ns07aLdSrGC806i1oWsy6gdrfN+xCwwGz8Ni2bfXgiSo6Z1
2wI7gWT/XwYNHzoWo96iS0reU9x5GfkQJixCshfEUI2MOQMEeG3SxEraBzTq7Nc268xWW3PnwxeM
zqnq96eZFFR1+agLv6AJSxS/A9YKd4sJBieRwBxFmJ75ozsVpQjldRRUjl8xh9nX3TvyQTo2sS7K
VppxRGFG5S/zmuIFIhuxdputsNTWRsUma9/c4m9whoygF/ULpVKYSr3AtJGYZoNQfeJndHIe0SgX
RyK755jVpeKIZROZwo7h4r1v0X4QXerE+R7zmXgleSWORSNUyHcAolU93TSerMxt8Hp3qRqxvdbt
wnz8Vq95uOFAS5B2kTSyU6wpRdMn/N+mc6PIgXjnb0jfjZE0t4f9Z1wO7qREiI0Uag0dRbScr+Y6
7kgmVRjTBn9breoZWA1Av4zNmzVMMDVPhb6IetiIY1LOKlY24A2rkG+a3MoNWR3C1SS894hkBNzz
E6KunctUGijCl79Ff5uXp7H10PcjeIFHPxBFzzsu0t6dML24NJFxbE75ljtr3CwnVt/fOcsr8exc
INUV1empOsaoxEUfW+Uf6Xv09/Z6QPZ9DUQJxbJF8etVbz6izHU2PKyiB55I5NQTGWibUX0hEiy6
o0LoTlkXuaaP6qPdj4Tj2xXtMYJ+iKlxbsdyZ/YRgTSO54OUlDneXGJiXaE7IKqkB04vr906qhMb
MmrOh1VP+u7BF5i4p/wZlPputiq5xEWgWlc5gOsi36iJRPMoifNjLQzBWfb98Z7onchMibohfSBG
7NQIiy0AF+btyUOrFrsO6FELiphJMm4tkcAYa/1kbtaQGGilFCgSZdxF7aBTBpNBPmH6Ijqc491z
Vn4URwCNs2gFHruQgSIh4ZqieCTSvV6gl/W6/wlbkW0pzmXiG+jDsrS3FbzF8YMMq2d7C1pCeIV5
CbuTGHQmdGVEIa8HWcpzR+sAsRtBwGqfs5FAZWT4dhIVeauUBnhO+VQ/q8RFzELjjhBoqAI/uRfA
tuEitCtgPN9QJ59iyUtQeCFCwotmSmtO0whOZMXuc36GX7pWTPSpGCFPN3/9+WDA/C+vjGpm7wo/
zGcq/58Dr4rA553hQvYdq2AWgP7Kna+CV0IX0ZNTxjJTsa7dAW984vxNLltYnN3aZfN1SBFB235A
cfFeMd8mjIsLxpq4rjw0vceGthaE0hr8/A7hcByvxRfsw+FqRMhWbvlOz+umcodgmiOXv6EOIRam
T99dFIetzzdJzrewsewKAvk2p24oVDmt2O0evY+ahHqOMJVaLYyrdEsU6pZNgKsFzpptzX+fdhcN
aWzwxx22UvlyHRZQtg6vT1K1OF2Tx5lVaMUpyyO/wUyHvLmmOc4QWjBLJyzHDAI49g1jn7LgF9mZ
kCUJxvxsZ25d4lQSmQVKS2EJ72X/V/0jKpLo9wgydv63GDNsf9EbxEO2gdXvYlSwc2UnPWVovZ66
b/Nan5UOqS19WjTVk9+dy0eLWU0R8Ecn9DfqLFt4CoLRyh065V1Yd1YE548UJ9rn8uYVEGgT0DhI
ndkWI4BnwHr8KNfJ+nKUkPcWl3L/UpPESF9PCLK9fmqua79XFm3Uj2cE4R30UYoLewgx1Qs753ub
NSI1Cmyi56NPFjT/J0sIEYijc1B3O2P1WR/7kRSHr7Hy+MlUvkthFXcojyy3Bndw4luHCQKKBU7Y
h53modEXqxGN/E/OqQ7DJyu9XbV/7uaH/FtJ/n92mG0YooSg3Wp8KQqGOC4OwC3WVxlaoH+Wq7ES
jhwUcjqfiYJXIsq7y77JyVxFc9UUdX+sr9W/vnB+wkTm802hRIshWxqB0uD8gl0zuJ4fIHSP3GQN
t6X5urPZXQEBmeREjd0st1/dcr38AU8YslVpgSo3+sdWbbwJD4Pe48eTzHqued5II6n8ACMRgqnJ
re9EtvNrUXHWJxMPA0jOTgwb1Ds2Q3e0WUDBV6UjhrYe7H7fNLOEAz+3IJyoenehAa9sx9X320q0
6fholBLRktGno3cWYnAsfiPSy/jFVQf5QdZehXMfq+iaMBIpSPWgWSlv7IA/o7ynInzGAfvXG/Bs
qnSoEQgxwG2xQF2x3UHYf1jdfOSV1F0c7BLE0/cDYI4jfA9bo55MpVajWI10hXTZ1vS/CzuaPCpj
g8zoUwN/jjvE7k6BJPYmzNQt6+0HD24Lkdv4uYh+x9jBg9hZucZLSLQbHVMIA0/LqIS2hbXgnNmK
BJIMTACbF3dgmajXr77LP1rMC2HgKGipclGpbXso/MQaxnjtDqrz+oj3+LK2tjBp1ZlqgCjRkYZ7
LcpR8MjpjULyS6zkMNsQGUaP0RDzp81shD+CNCd1gVghEGYyQboLS382WrbPG8lgnLdgLjjWA3lx
3cePBXE7pKQaRDxIuRLPLfD5XkXWrniOQQrbsQ9YXSuVvRyIUAFPJUMniWwTnhJxcOQnIXS6x63c
HV1qOlRc0uBInAPTBF+4Z889/xG0hnhd33DXXDFUIEEhZyH9HLmgjOAREY+mWq2Ru5lSvJydH2zW
GiBGeeOgTqJkUd44dp+OBGguR6OQpxsVMB5YvmQKklmGI32gW312LY7lU/PF2XOuaoH4iy3Rsn0e
5TchmDo2ll2svqRKkRm1tXIB0NziesrAM5POfoU6sj1q2swIY8lQ2ZbUAiSxJ84qePpE6wpQTiuz
8mNfyo8+LIEAVc9hSLkeNFKImeEDh95AE2Jdajk9jTrqjrgv8DryslGZFonuHSFUTQoBsQDra11B
vEYFNuc4y9BJiF9v7MF5jf91LA5ZVPw2RVp5rToyrtkd+4gA1lUkjggaoml62rfQQEZ2m5hH0aLY
l3tAJCKyFVz65eIGn6AVN2QgfF9R3OwpVijVAD/ZLG3CxtkNe48JnDgHMM8hVgQIp8ho2+DGZ/ZW
6bgiMHIZaeNeSwdn8Bl/pBGWnbj43qU0ebkGhIA8IcQxjfk3w0PCU7HkxLMh5q+Ipzt1qI3W//gk
ilPIkKQPxpq4Z23OeHDYEEwjiwDLH46A6x+FJ4NkyIysxfg65nFVepAEOWAqqkGKoUen2rEocNMP
mzaiOnDYj0un93Cmsxlp67jY47E8X+KXIM10+vv/Qi4Pl42u+w9t4HEr6R9nW8M44haXS8TUSECG
S9dwT3yPd+8JWwIvG1ukl3TsosCJQ10IwL16QC5Gc2dUcL89CaTA6lX7Pq4nom1l+ejhEaVFU00c
o/zobbzY01FsaEVm87c5TGgLx7qCj8fesNZ5W+87I6M48kXaHFRW3WvYF3rMZuBeNbm8NU4DZOXb
wtpfhp4E28ao8p+s8aMvV1aiCY7p9WLnLa3qG2xadKyBDF0AbJv04cK2V3W/Y92t8269rTr9RI7T
Tlx6M10fmT2pEJ3wW4tG5/50lTgluX4BRG5HgzTUG9cf1QGyvFq3PXndEDi6gZhqco67/UNhdcBl
cclw1uVjVVq5efzgUivjWKpl5P+wGNHmSFGgk4l2nivLfK1ah24wi8mI/bg8sX145mW5e0b8aQSe
WmDjoq1WtUo+05A5aFTemv8GyuO4MuvbuMCicRxtCGwOcpqarEuPhZYdPjSuZatGYxGgGszsdawo
JaUmp0oTMxyxnSD1A6fZRpsF/9LnRUKEoHF+Px2yxdmX+Pi9TMqATalR3Es5mRES1/t2dQb2OAvH
o00gDF3BfXUFQ4HC7NrV0nieqLAfJeKt5XenYjyD43vryxa1I5688QWAX9Hh0V8DlKGsvvE9uI1Q
GNBSixpLq7QJHvS3Nl442teaGrgMLwSTp+Eje3Mg5mWKGh/tT7ScO5sUXH43t1ya6Hc0UYjyBGWx
HKpodElCCCRFgLMoDx3j0sy3yU/1f1HE/zHaBTVMuhvO6/U+Qkjwj7SVgTAFh+VxxeQ92GbSxJBo
eQMDbCQKdFb1fpH64ushor2ajqqf9ixD/gkAO93mqO4VELjUb1Jkj6ymhTSvEjN2qWVW19if3MJz
MWPuE0R7zZhWhaDRvXlqdPH303Q8gobFTDPThOrKkW2XNgsi0Lm6UlrFZA+gFJtO4htiAKUBFXH9
PJUd7Rbhg3RkkI0F8IVLR15iF3wyV4b1ts6YvwXHeWZXWWo1hfPhAjzWfKFkmlbvC3C+CzlLQSjl
xzSRo8XCahOMcBkD+YRbAyaQDix01XV7n2pb4lNt+EcAsqFFvwWyknnEwD0M8N+l5+Ffo6sxAZj1
CchGPtXvrW04f3496/sCw8HSlcukDrACuhZhmIX9Ti0E4N1MGkQvFMWt97pbNL4Mp+zfTfaZBN/R
YF3zT27wdYhv0ZA63wOXNx7oVPFI7T+WwNAChIZ3Az6eYyg3+rRICOEgRXx1YGxqeGrD2URtmjT+
2opZ+zYtX6jIueWcJ9W3vMzq7/krv7XEBanWvuRwq5VE4FnbTkotoNsxyGWkhIbh9N9EsqXC2/zy
oukI5FUCFRCUQXrhDGci8033gw4MZKss4OQ4z5JMm3052oDcax3kCiA7zPkn5hnXWhCWGdkrDM1d
dCV6ymNZnfFvXr1JHR9rlvg0d8MqTEptlxEXl98FQ/D11eyRaBTWyQ4GkWnCu389pYuewwcy2PR/
CZOuX2SENBtU3WQKfA18nh7b4J3VSpWP2T0TSyLd3NY2Bt44+TGlpREwabzX/kiNJBzn3/Qn4teV
xhKN5sA3aTwPU73RshVHY36D/IOjsMEqjHjrJ6HSV/ji5DsB3xEUcVvHtkXvJW5MpIBpUvaBSLpL
Sd1Z56jintLHCs2B376k3M+qyJ8qIy1LKREvyNAfl60vyVUXGyalIUXTfURUQ9iGj8/EFFqpUMlF
1sUyMuHZBHU3w2FWqE6kdtUQpj5p6iBwqqBaZ5x11Ky44BvDORB86K4ZSC0P0VS0vijT92cdc831
gwJ8nttkEFTUbHsgfsqFGQR7GafLbjhh79y3r/oUVqwPEEVfMsScdOHZOcGAnow2BuVliqDwjq+Y
eLCR0li6PNIfRTgAgsqyl/AiZCFSY9HeqwoLMi0slXRxNsOzhOMWj2ikJKIkAzpBC5oB9zmKodf1
Hxu+uqPvouYdYXopNA6P+jOQicKPpkD0ki2dB7Wo+ApWV2CgDmqi7V7xQgasbVaXgYAIP3HW6Br8
S/6qyXIXDBERo7GMka6Ok1jO6OGJDI0pyaDsxtOF2ECEfUWDd+NKlJZ/hSjymWMXjBAryUy0iLEg
eo0znUexlfNy685Z28XZshIkipI9/4UPpxMNczsZ7LeqDE86kY+gABLDTw4xMBY/6wvYejz93ivB
d8zldMUYE5gy2Sj7LMVVvtb/JfkoK5EtX31xRV1SSomJpett+7bYa21VC/b9yE3VK7S0qgnk+E5n
oEzIQ8gG8cRxWWPSS/pTxBqaJySnvXfIyJSRoAWsMKLqucTQNFnsss1USNiyq9o8a/LdqC7oJL94
Rh5E8LuouqJkitaUcyf/CCTmzHLi+2SVx573xv35AxlLSSLnO/aDPD8LMCpVoidH7dOigLo83kVr
jU47D9iUCa3s2g1oEIO8BmhjtExM02tYE36YtT0lO5hLwGI9VCBb3KQq/WW/3F//kmAf7NUn21+C
HQ7PJh5lcGK3UmZRJ/3aZAoippaylU5YX9TAcxhjvsL6DzdGJqjVVesXH37IkN4WyJKOlFkoCMDb
PHJZdsGcH7O3vdN0h4nHzBKtA0yf9Hza2bx0fJ9W6oh7HK/8LVcYBrnXniOuqhVuUUDJ5JLO7b+h
KNygO0ZSpYGc2XObo4mAf/p/MYzdNuYJl7eXHf9+r1B36epk7op9rCENaMeOtguyXEWJcidv4BKl
aBKHv5neV/TLfE+LW+/VcaVvH4TjQNHrzeaP88rfJguKU/jvXj41PdTKlovKe+9mf3joo/DRbyfk
iQtAaqojqZ9wtiqnfXpO9CXwM3OJv4Fm6RkeRminT8Ff5LiT3lctmWp8RD4bhgp5l8MeJ+jBA6sg
4wbPVmK6RLHSeqkgZyhtnCHcpz/KkeEh7/gjV07lOaOoKkzyKpEyQbLAuj1o4qVANf77bITjgZc/
tvnewjufhXvoxHTNHQM4OiRTvW7MDR/RVIMFhQtd4W89+F6FjcNMY/rm/Jk95vglQwgTR8eMF2lq
tOz6vqovZn5RuZF6UUHUSMzZdNfHtkHluMmMhDRp8TEmDDKfQn3+meEMhMGD0w+Tf++ppwOSLFWH
cNrMClN8Z9PM9guqPWGyl0BWTnkdsC9S5o0AnSrCsG7LQQ4d82Vx+K6MptrHSLuihrb+sxI5iXKb
w/Gxu/zWpA7C6X+DZRE//r6x9AO1kl2OSh+QzgjuXVznbOn8ns8F2oEVNHBY2uxypxKpPbulWX+V
2x2uSozUSfZnZkYoIZ7WdpLxttvm944ziVTe7VTn41XNccCJRlNkDqumetvQbPZatcMNZmAbX19C
37wEjAE/e1RTiiWR3zYgwzDxY3hzP5kVMSaKNyrKZtFZWginagPpY5MMk1jZ/0xo4WS/WZ8aoBSy
8Kac1elBoyELl89Mn7DhT/XaQ/KcqDzkmkPCpAyKCXiMi4p2rlVkUq71cgwKgIBNAoiuYcUO3BRy
tkg7C5CQZNZ3VdynJIO+wiw9pt3F4GJSBDrwL1hrN+XTJMlllHcwlcta3nbXrD4D5m4DzNBthM63
IFfgaJBSB0rRd2m9aKCnbBlItExq0uZkjLOClmBcgev/9uZO2I3wiJGlEJs4cPHAzbQL92qHtAmh
PJjjhdKmocSs4/b6r1MAA1ujOjlK7Io3UsqXDHAjAcr83cY1XqPSSi+75VA53S1ttHHyOgO1Y6C6
1vLsOX5ZeFg/LS/ei+9Nj45b247QktP2Igoe/k0sP15H8easFZzjmlff1KLXszsFgJFdf+9GYXa0
hwwnwGoR7yJcCqT35tZurFet0E/lr/gGFV+fB/uVv3wpbC32o95WXvqPKSXjOcgFgVKlpaPlG4mj
O6rK37mFKtrs+AiGS7nBQ2851ACNnIqyxfkqH3x85KvR9FYU0nkwOaigKhGpReGPMLeZlhQXr13D
3TjBPgm8iNivhiQUHJ7A2TRD6VSbh7gxEageIdY1NO0tMEP6++sjdJaxZJcPP0R82PRordM0P+wG
iECbtBpECsU9uSU5mG+RvHFOMwBD+UU1kW+fB/SnqSc6s+tldaMeYiFPKEsvbWx94YELSdQlo0kd
+dami10lGxN7vnWO8zXps0IWbpvg4HggNrRAsnCrpOmAQtpPpP83yOJkF+QO7/fbJ34pSoGOlmgN
fxjG2ltKPVoC6MtamvDVeX4+7gkh1WJbfg5toHDOsqsqqoOvUQQU63qmQqOejHeES+QYYWxAp7li
S1Je4SmuR5ALG4GL+l2D11HGbRyh5WIpI8HcW0b3Kv6jiNcGwFKwSKbnVrQ2VycUIWmE2UQUew7q
p0HBXbHEwmCkmQzYVqpe813/OgWHmGVcYBG0Jdn9u0XsFYJDdOa2Jx6R6JX2sGOprufubemWS8Hf
pfSHOp7rcznY4n8d8XIp/eAJgTB+rYQv4mLLaiWCfqKhEp/9MDTlvC+0d4eCi0u61JQzLeXJeZK/
UONWIMAHv9W0dUfsPYbtsb0A4Pl4ygG4y0loGvfDnVemcwb+SAxkJ80bf4o9ZfIR+E/gtxjUK33U
PD1oBSf3ssbyGKcX5JA6YkRvzxfPrmipa/uxuqSwma40EjSnYg2KpOQU61bD4/KtJg3/V9i5B3HL
hYRpg8Nd3cyCiTXK/7RZaxtmJAqZzs9yJ86cPibFLj7j+ea6bvcwXZk2UUj0HEZyUggjMqJt0ruU
Y3yikr/bArxSwSAcksb0e3dvlm+DqptLLk8e2MQeNEBKafduR7nJ1FcEHNoTcewlnIZ4ip+nz3dd
J2XDyk7xnlxbroHeDES+zk4y4kFTaetRt/jHgvFEM//1kx6NFfPMnwRK5DHIaVNJs1ih/dwgKZnS
vx+lFW07ITFYu476/eYlENrJI51d/rRsbwpFfqrjM7WjUbezulfllNysW5tcSf8hf5gljLKF9dGL
h1mFNjzHX+IpHuqZQdtxeK5Vsm7n6UOAQ8AxR3Ct3ckapuF4hTuMt56yATqj/rbq7qfVEKzY22xN
dng7Li9e7p2fItSFiPNzlyg1ccoJRvkueVkXAsL71htiWG6JItPEW94TMP+0dI0Lm3fDNNkxB3Px
TKWiH4quMnTO+gHjNYDyq+fb1WivtiFtLb7XN+yENPpgTg4wgEhxG5bElQ0aCfcKsFZFgcsW1YoL
1etbsbWrU8atu0whcS87bqnvPrT1f0O30FyK2y01J45TC6biQWPN3tVWQDneYeGppL9sYPPKcEDE
W51dq4Pn/j82/n2WWBZ29oOPFfKaL/5ma8WM28TnUDAqg7ALjkJQaBgcpIKSdUaOfKOCkQ7mGfEM
sW7KJK8u9TCGiNUY7HLxEZGtpXN7gu2qjJ0LTJbTUL4jzrC0JJwjKOROULWTkw7BpQ0MRtdgkzZR
w5wogK8Ja4jz+dy+hvkyMPoX6zpkeeH4Llt2Vdm1kATZaY7VE2sygd5jO5ZAojGBUHFvdO+D5iCh
NOzwGUIbmlRqoxgLTu2FBjfqarxXgpjEQ7aPwBvTFs+M7+hdE4wpzWNJ2xifKS38xgGejVgUEJVE
1nIRhyEKoVYzcsawLFjstWDNEIY5W1UMAWOxjeHZO7NQ8q8RRc6SKr0loYH0xIOnwdOBwBdOkSOh
qBIiX0b5MfYTsmeGFts9+LG5gK5nHvDM+IGkf7g3ssO3B/WeHwy3XBGWBo2yHzE44cn0RwTlFmOq
Ksoelg7t8HJbPPGjj71UPRpQcJGiGg9EVgsoVTnlQ3vaNqXgh+R83byolMruiRGVpZ0Tr6bUh2B6
DML/zVMs9sD0nBZgGRiiSgmAlwsHwPJbCjkJp9qDG2+hRwZ6gTSGb9WAbCA5qch//M9yVGMob36/
iXwS1ySEuxugbQLCwpfhltR1vwMnpmgNzKoJLebORf1EpVGjLcBDx6Buz706vG4Wz9O2SQtmDu7J
G6NGnZG7Q+xautF3QF54cnmhgs2qcYkpseseo/VDpZSlXEGnEBemv5coTZCJjrAtamLp7th0yb2K
KdNZT7w+YlmR3Ppbi3U1yc+RkQd5UAqqvm+Lf1WxNtOq737g/6jaRWu418BNYgHmvWDueEioS/YQ
2eb3nTCbrn1h9wXg4urHjcvEssq66j08z80Oten4fCSXjv/VBVauJUMc7NwjAuwnfiP2sJjQtXZO
BObh14LSY3vcyGJGeOaNp8p5iOQN+tkrNVKG2ChIhw90LQqumQZJ0TlaovPHYkR7JmdWO0DmmXH5
RC5yKhbVVtuhFIrNkkv59vtoIq8ylYeU7r+KhtPQXugkLJMm8ksi1dLcntaj97O06zlYnx+bRsnv
d5pOKkDomn9OJ5c+0nCrS41hQHJFJ1/GEoTHmXXFgAakaoONXUhIHri00EB4d+N57z4au+6+AQmi
hDYUV3Cy1TuQfSGGkaW+SU3k9RvCpk/gcIhkP1fh4ErDXGkvxnMW56QsIdPQ4w8jONrAlY+hRDpv
vUYSVGCDD9wEjQM8uLmXFRZqhXkSd1I7lePVp35OT7RHkGgRal4UFKboysp2hCj+7/qmphYCr6Zc
wVCvqw9xLI4PtUetTdw2jl15bCwT7oIoIOaIbeGBsq2ZPhgVgj30sOf4g5nNy8pUsmZrr4dqN74F
eOXQ+yN8ubbNpPeAzMsSSITPvE6Bi3cwUXYnwQGhvI7wsWzXofvVDWzWuGCKayNJ6iDyAiETIY6e
1mY8lsDVPIvgyX+Ym0/9Mkx/v55bniifQqO+eFddVSAFbgC5cqCzcUINV1KIoexRAYkHtnxbYpW6
LdOgzXuadu/9wXXkdy90RwEssu++x2pP71/Nfg/A/+v6b7o9nJrY36dKQSsgFzjJlMhmvmkKc754
vMKAfZJr7HpJGaRCCQpjE6icFhLr4D2aclN4kEql0/Fl1BDlvNqGk+2A5ptV5qoUmFIkQJQmoGaF
srmRguLmHptmeQQq67DtGZHEYx8Jdw6i/U/4K8Hit8+CfSNCnWlBT8F0G8/EEwn1oVFXCqesEPSb
Zhv1zpuE0SOfelQxy/AmIgKPYzGsTnzUGQqAaEylxl1wBYAFsbaDCaE4mjUlK9lAnUaDIgCsGQUs
LgdfQkfrnNdH+0z3H5HbBIHjrflTbNVuSL0anarx/4Ka8mXrobDRVA/P7GuHiRvT0tZTjdjzP9SC
lJ8gHjX28qiZiZGZvhqTpr3AxLtzzUzNPF1C9TI1LlRrPsXOaIG/UBsiY4HThX1wQtUMTALh066A
F3yE0LNAHVFjaIfTJJgjAmphvzBJudbK+3vndiONhaZ1z8cxEnocmf5nZubUVwRy0bNHibuBUP2s
r+XwGubhdmiIRgli1aCxDBEj7UPOB+/u8SppUUStZgQGQ1rwnJ5AsKpMbZ81/GCZli3E8eZGI6PY
LIHLq0SOLNFfhJiE1ytvKNRMIleRvAm3g/99FwKPP64gVTfGsixs8mArIshzxjjyJA14Va1/wShT
vtSUFl4YpBvPoCvP5JL0BNYGVNp3zg6T/Tbr5TEj3hACX2rIph0yp4dj/9/+QImcEM6aXzAhFMnk
Mb4c7NK6cd1bozYlzpfycv94BxwPseIO7CWZUQ9e81ZYkIE6G531JN70BvknlJwNVG4R6HqPNFr/
eHD6TNqK7si8/ehDFXqHv5mKud73Sra4BDoNmTCMzQg7TXkeIv+UZTN9SN6AhGBjNxwBwVnxOJGf
nX1caQ1zqkl3POIHgcNSxh3TkF/a3VrvRvWaIxo6u6xeM3r1a6KFNanNAOS+6WOpmpuA8q0b5AmN
AWi3qZgTxzPdvMjLPPacrClrWTB8h99XtFNSWXRYjvsjB6KB7CNoWizolPZHntzEWUer3kcdIOVd
qIcsKTqWT/KrnfiOuJj3Oyt7F5r9S5E7q7pCpCEcQAz7cRLp1Dncdel4ikqS9yZPi1ENN73b1rJ0
8iI0VTCI9Y0WL28/iIKCVZ/wP2/PN2lxmBt3nzPMglNskW5SYvLV0AISCi2Ayne+6nWwKHEvDRCl
NUWcs4FTagoF6lWGOfyjbw7URCerfuhyxy8mPV9MvuASIqvBpyRrtVeOVjMoUAMopEOLWZJJD8bG
tq3C+ZyqqHe5sZKXBYb3dIfvsx/mChmogmnCfwEPx2kWsqnSaWJTlBiyx2Q8YY5eO+ffrOBvCyy4
pc2kAsai/lUQZdaPLjo0/0m/5ZfyB0qrXKGJsZWDOxD4QN8/kDIEyk4DmPnDpOdnT1QIH9XfbkV8
cFYzT71IUCmiv6v+TzPCIIhR//s0CxIoO0e0d+mNAI2ZtWTa5Lyk7CD60dguUSy5YQ49grh7G+2v
jIOhvZAnaf36cv+xN/jYmnHqV35hWwCU0dj+2v/B10hbNDQ1P/gHRk2kizpSby9n7YCOeIgkJcmi
WSxEyRrChTJoODdRYVP6RdDK4Ry3eayx8aSPGueGX0sJxqRaG5Jm+IlojG5eQy3ysuFmb9vAupvX
r9e3DWZI5yjuECIYi0W+FdHHCkQhEutjhmVzbgVkMhnBROGvjeVT+AjGIWdSgEAFr5/WBkjC4pmp
zhQFaqxFbr9bZojBSf7w9G4bavf/Vbq0qx4XCzJHP6FTdBjgB8k16c49SbZL3Hf5UceC6IPTGrKc
uGDLuj5QQ0YuWYsSR1JyLpAsSSCH3UcAuvAZVErfUA/sb+TFWNOfybutUcmwCd2iipH7ud6EYhMh
CjHatyDo2Re3B1WTnaq34JOte41sCcJMdr6gMOfZV/zByApx7hTylFdrwR2crZzot9CjxIs9De9m
bhxHIK1K0ab+rAESuMRVfNjloU96VNp/OT1qhUUkLM52520eDWO13anaScVPC8zGqmnNW3yU8JHi
V0i/YqZlfFbIn4R+CY+G4t3hcPUzZlp9OoOO7MsjicPRfzfMM58vbBzsalcfodEAcBc6QWEB9s5A
ZU3O6IEaTTA11wp950qjS4XcJxuKFd0iMKi5bKw9MC76kMnr/bfT2IDP0zqUOwUTXCGsNNRrRcqr
5hRXsM/LgD5KG7FjgejtOGmpKAEDtvl+2gtvyfF4P1opGM5iUUeTEo9N6aEXfEDybSXaVa80E3Pg
lWiD9AlYZk8HGlFrl4Ea6YwaZuV/oV1CtRjtnxdIbP4GY2a5fxEsqSSWopkKtys4ZMBzk153nvGB
uE+dwBRLXox8D+ZMBX6eVhPv7ZXXFOXWq+e55My3Yw7gw0j3d/q3nkmWjKCt/9CgwYsFkATfP6my
jcmVDSxxBbJiIoPlspcbA2/7pYlnfbl4Ras7GfdAq+PiJgvhb9tiwDWehpqyThQYHaAsbzLYHJQ3
APwhMPt6S1ctxgqX3KoiUskiYXsBJAlYCB88jj1TV54BmTFyVFKAOGqtWqGlfB9qxJiA3rqSeYLW
ZUSo+XqLvfGqmSBrEoZqnF627odQQp4yjICW6TFiyJNBtKIo517t91tOlx8WJtabNCu3TQhKDs+4
9J62D/7jGcX9tq2ro97aOAq3p58228vbYXLRMfSvPUjhbU28SEtlvO19NLSAOuRrpsU3PO3jIGnj
jj+7nzwH9xepA9o61xpFfnmvHOGGqVJ798bY0pT6jmusRu9nqj/0cLzbsdQ1Vc9A0qQfzsv9EVnR
v4FtzVHxeJFTRruBk3Tw8Ff52Fj+eahoxRwDpv93jmtBhGLK6UHsj3bKCtk6qJ48DNGWMFbhEEGY
Prrvl5urxQm+ik4gU8hJYfDIGaQbqR33/ntrZdY4i+A+tyCH+eZ3N3NbVNY4P2pBVy7ySsHWAAKB
YSoR00utTiKseaZ3Ws2gCBnLWB+47+4RJTLcV488F4/+aAyiKuWrlU3yUBp60h5mRp0J+8083147
rUDJiT/GzIAdLPlMeqO4PePDsXHcXn8gdFmAhYT2jQV9PgwW4nVIAGA2vAvSGdWmyw5ffuLZqZFy
A96oj7q2rvo+DeSpUObMKKjN9Eawx0HeRylxpS/rJV5aPS/oUOhR1fvLskQ8wThVJ5tmIB4t3/4z
qmKbrhhtowqjHrzXVyHDYK+CELQOPh1rJpOcNrKuSX6RCyyJYZ1Yg3lxd23bVs6G37RiSAPpjrgs
gTFEheq834m9NrpZK0fiDhE8DnlF7o+t8q3v46biVR2fbgOAomCfwAyOXv3ivtnJEBiaSYFs05CH
hv9J8qHEQtpKzVKiyKlQnpYMg1DIWnE6XOkGnncKMBYcksXylvuOZTb9dgRGHC5TQxkoZF5FSpJF
8DptFjeBvotjLZavr2+Wy1XcgVa/jHOwozgJOlVDrx0otgi1aznVJyHzKUMyRp9WKyU/T8LDVgIn
6zh29xbG9QbffW/RO4ctY6DJGhQH9/0MYhzusqD95hkq37/ddn1stnk3Uc5gbQqF6zSvvGSSGlMt
80uh40kd+LHND8s4hF9SJgfjGnMPZJlv1HzU3ckbmE8Ee9vaX236/8Rt2QXJs06oSiEjw8twP8Ei
PARX2+yz28zK7+vNYyI/j+QhGicDHrdB49HHlN+UVko0nmgfZAQftrpnr341S8zSOBdUZi3C21uc
hCWJC7lPZ/clKuDFUyNwjfzHsjvKDpCG7mKnI+TZ/U7haVABS7NnTopcqzvOwd10vYhkgMYrYjB7
YWV8RKUoupqAsnBWBkYIP45UWdpJBThni1RnlKCVfesez1ZB6lBH/uDGhBIbHyXtXLCP1gv+zJGU
FHIsX5AtWMFbq72pcDpmgH9B3nxRm1SjQATeTTo522uPFO1DXsDwXe7V6UqfAeDpZ3z2Z1WnRk/F
SuSi+nmSEeLu3b14N64D02V+3mP4RGoHuLHCjypuv0vVnVSweWDC0QYx1X94jhD2EnCJM1WXrrsf
7eQd8baQx2gFyFNKl7IAKBWMss67qqRkrnLiFxjn4KcKGZOfkaAZ+QKPn1xTlydJ226VdbMjqUun
HhH2Hl3CWUA/njujwv7sqLjHB5XRZMPZcKmIRgzRJ5SyVf0BNBR0+CysWJgf7OLYwt4btS6Wp7nn
ywj1Hqy3qKerlg6+g4lpT3HVA21zIvTfxhbSKnhW3nI2mqvHw3AmNS2dwdOgc9MDgMogiNDL1qZV
/bfedy6yKYdBz7SlcXU+uW00cN9ldNYT5Fd/n1cs1HWspUjm4zrf5Kh+0PiJs5R5oZNqTnyW7EFZ
1dSxNifJcuDihJa6bP38dQ1RPuhmp8AAiW/A7YoE/sA4CfQQfM306XRPs7Ei5h9gQLhsGn87Cz15
8Nlxxq9Xd0iiTh27ZoouYGVD5Bio3IVJ+k93V6YG8GlCxS/INF8E0CqgccJRk9lJS7BrTh6BDRPH
VPyRcYrDx0xSQ0Ae2Ubvc3BMSgxztvt0OqLpFvsdZfURw2aB7VOXIOSrB5rR4teyXzm97HGylLpB
/31/g/crR0jaXXn516Lvd7bCkQkcvIgQIYYZrq1TMzTwS0eO2fxs9NqUMjGNcTc1avDNqJIyXSFI
znUPZvKXjIeA8OaeSXRAaVwjPW/AjY2ZUp7hfCgjKs6JImoSgzi9ruOCw4EZpIddBGZOSVXW3SqD
yY4Pzu32E2Wk2JjnC4MAewIOH1SwJK+UE3LY9wtbwCeYkTPsqM1b+tpGDwmZ2lnypoBE9ZGcbuuN
PMrp7AR2AFpIV+Bw/Jh29SnJ46FdHt96Dr1pZl/vankC7AJlawb74S8zrSKOrHrAXfrwwYyc5lef
PaRTEye657fLker9BoR9aEeuyi/oskG6Urz3t9vtMlmIDvqx4qYb1tf0faqtHWjOOTYAgwqKy5CK
cLE9pbfkizHByCTK0rCybia17hlr+aHebtg/38yVsLL06qiQrmNTaPvhdwKTCjZmbxHmNelVfWyo
u44fdhYf7fw5oYtD7HVN05N40/vi6j3hDoRgxR4DIbGOI4XkBFHUM14ntSqnbwWzBrTzGGiv9f8K
mdccl1sg3NLGHSaLHnEpI1v90rGXI/kK9tZw/+5TvDmRWNFvWFigFgpUB1CVBGWTlXKCG/TYcXaw
PjD92ZrjZ4pmVi7h4a1VcSRNvmzmqDep28+bY00XgIKg12PUlj6bppUhHA5OCJumcwRfYR9oGz2F
9NwWCM8h2amYP78w7ysWeCGVsy3aEFnUWuL57sUxvenF2/v7iRfHhZBDiOlaHs7cjFVoqwFfYn5U
umAW+Pu/I0PgKlsQq2w2rRfxWqMj5jzyNRMeqVMZsmWoam6i8TNK4zNB8OmvE6MRexiABcqPB6Z6
/zXqyOv+voT2GlgvPRKytivyMWtN7LlWNNXOeSviLpGHi9y6ga311uaWqb+0TbWzDnNE0zJKhO0H
Qlgf4ewxBM3y0MslPTx4LcoLanY4BRwEqusDOeJLZR2x9UD64aBVk8YqUJpz/rl/4iGAHq1EUTqI
VA99tNi6j3TMSfZvTZfFI6VlR7gbhvjjbYZEO821dYgQQYY6Mnm6ugJPa8hIGnhF2t50pa4ArSJY
+JSA4b6m5n/o9rjAfHochCpYb13E3QbZqqUiR6YyEDM1BQnVOWgy1XqzCZ+kQVDIQrSmYLdlB0dq
G50C+iy6LZV5+cjC31T3WIjYfolkQOQnWbLzSB5/rCxbUm/2Iac9xiC8SCysemfA5iNy+GxHeqai
FxvDkZowFpkJiiTMUKt+i73fapWRJ0vWiY8RN9aWNdUFwxILMIMNjCy0hwUzlW0gNoESBraRpdMf
vpxWPgefRuS9ezhNoKHo52GMbmMuzmj52EvpBbVLrtxGd5sUrokw/LvbcaCVLxrxRTnbi917B9BO
5UQxG4E7CWqI/EAsdtM+qwJRkRlbLoOLHK+f9epRnhTgpeYXeX63a/jH9Fh6rX9GhCYpTn6Q1LAv
CsPenPyk8vu1m9p4YTANJREMBYJpFpZG36Y6kbTCrab+Id49upzIno5XCFu1q8QRL7XEoK18hcDk
h2fJEXmcsnJZD0J37+CSQM4R8JXrdmAxAtl89oLYXs7K/wqOzybahro7XjmcRbPH7saT9aeqHlN5
7zGDXpOh8HwbYCMSgOQ/t/GWF/q8p2qhA6+hcL168qSibCGR0UDLTKQ8TufqlhzQzuzbhjLEO8/Q
oOMaQSHF3S9jATQi2PqBkXXsyzvdonSHhyHvN0ts9YKzXRj6mRkDhhCDtTxBZAHw2km8rsBnfAi0
VKs16aFooOzELqm7p53kcFdoLJ1Jg+sUZ48yvu5uX0V6xOtaxduXAaKO5X7XdULaWKwmvzO0ISFV
nmRO11g0jsyoR8SBC0trT/kkSvRd4UbDA94KrTp8fAtq+jt+amala+YW3DHLbwBptDhPNb5YdhyM
4XSWJdS3We0s7kQfsZ/HWEo+OGR8kAeZh5IEVppe9WgzWNjHIWlYTO28YA4GxEanN+JY1hoy2W6N
JRYddepDbLwxxxgXo/DCA7j9idD0sfgndwoVQu2St/Jv5RxKCgfy8zpZuJfsV/C0i+2Qczxha66w
bJjuAOHcSk0mzIuEdXGswBQ/LoTBSP/1DyrsWhDQNAxC0FHqSXyV+COoCkFKYuYe9/ZbRAYu1h2v
v+BRUa+xHHh8x2f2iT/PbZdBFAki03K6YFniVQ2AKeJ6M+jnDxOC5kamSsSocYzZEsmCWbO0yJvj
m5KKnkP1+YkmSN7BXTq3xVL0hm9ZqiLqxa6U+CCkxRL7NbADCH7STIe1Ak+alIbFJrn/4qVPfHGV
uUno/hMS2DNat0oXgfi2zG6JEP242Q0+9kTOnsHLUDkbBkbHBUDzd54hvsVPLyHQ9GpmAJ/crkFj
PZFM/cS2KCnNwP9zNKJZpYOvrHCgtfheouDU8a9eEibW0OWcsdKNfDneXpo+8wCjY9V0ORAZ1Fm8
gBth0wVnuSOeySNh8H/+hp4edSqr3LsvZEh2/KhRDyMLNP2YHZ6rUsgrYxSMmYqXuj5MuvTHVUrr
KjOaoBCtuJqGHGYGT666OyQdDdDXp4JwImZN0CkFi4g/L9xw9746Yd4UmjP3N5verNvnx9uatZon
5h5kapKDqqSasUpw76BbZpNTLcq94+wkMz6/uFs9yXb0KwtCpNZuJSUPwFzzUILPBnV++YnkhorW
lMPzlWZUfw+/BJp7pVFqtPxfzTLDKOqrTceLPE/NZafkkQbCY+RC8tx+Q2qBvOhXSrM/2dYeLfMO
iiROsKTmWEp8cOPUDaaZ+J9z1BNrAV/sQzrKCYbFiQKmCs+8ysGu0f9GkArPSddeGuY1VFA1TEvf
9+LPIMywQg++tTIUp1sGet7A7MRieaEkZnkR7U/N1I8AmdC+J5XXE6n3O4kR0aVi1AGuFNuAp4E7
ihOIRS+7+tWvPVM2t9gRDGd3C0HqF5eUIkpMGz7MAQ6pOGzik4SJH2Nr0OxFoaEk9LjyZ5TnCAyD
st0/fUENx/y2ifZMs3V5nqGZlPVtysPLOHx3KV+N0VZvrzTsICMhpllo1EKgPDIwkkA4F6Gk1AfP
v3cqfWZaQAOrQdCLBZz+WE4rdYv+qDJivNbq16YR7S2cP82TI6fdCulEt7wuO0mx+Vj9AJQSOxQw
i9SoSIvm30Pvqcx8Q7h4ySlmlRehqC5IHCG9Je3WYtEPgAP3smeokq/4OoKD1yDTDbhNFhSFeXhI
rhQh6l0rhNVHRMzMZeT/AcVqXUoRoPS87fimn/EAOQt9W24VsQvdOI4+xbsvbEV7AwiwXeH/IOiv
Kxx6ubh9lOwihmnFu69INwUnKfhTLCLZiATZx+oYB35DMi0HMrreBjMEdVrRltDXZb0b916JpkD0
YDUKJpx98slNA5HoIkKoZa5qvAx+xj7vuG1rq80ZjC7/1BpneXnG3P9vL4m4zKSzW4HtF/shcomx
H1spZ5rxzdwmnzF4A3fdJRbgnrO5s7t/Omk2X1GgzegrBt5QMFfNH+eMyclI6tuauSIdTh8ZuQ1h
kPeLYY8CVdBLXLwbtO+VdiDKS+raDD4+m7mSfGE2EndqX7VieFhoHiox2NNueT/OwAIoMh1NI+Ze
t/qyC9g35acwSsFAfqkj5hHFIz4Bjff0vXgmj6oH+LuMJXw2anuzFWLwLpEVgwGWztE3TJWzKbhr
eh6qLNIp+56OTOZddjEJ8KlLMbrRJlV2BoL7hNIUqVloT4IOPODDdqa77z7Nyhh1oMTykJM/SEYi
il3FDiA1ph7iG+f2TMLeJafHWnK0qKUPCobssfcnAhNuJVJMtgEFt+PliIGvhPBVJoH871fHc25/
egQuGM5jdiBLezJEXIGih+MCSFgou5/g7wXf0nVnk4iXa/NvGVGX7R3ZaWN0UXLw9BUlhkA43YeU
m+o0vsz5p+lWQ1moINfbUkyp+LNNzyPOgnB2EIk9SODelDjhDa/EiV6dQLKge1E2YdVXJwvrg/b7
IpdPVRKfpsSYuWXlwLh5AeGjW+PhVxZwWDl9jxYufZrQ1axqz8pVviu4uSpXrUI3jLTXAEIedxFD
0+p6TozqjEv66SQhHK4ZOMmL9BMjSi4ZfyRXLEEa+4sgP5xl8S0vMnK3J7xDxNZI7PWdoOsXHYbm
cdTwDEHFzzuoh1y6h1FVzBjpq0lDToBx0CmP8VbIy1WCahmapjcqYOo+zd8AohPlNfUhQD2Rz3f3
xAmZRkQHrOdWqPcmXlcEf6RZXGWlK01rl13xywDPyDi7srAeqGoozX2mld+GGSuga+NKxHINjL11
LdyX/BTdGAMvjnM+GqHKUzoj4HSlVYDUe1ZQgrYO/zSZ8IB1/NNK2dZSLkqnpEKZuY4AP7jb02cc
lJtYGkGT4rLi+zOyE6kSi2y1Qce9BglHXZcLm8i1USQqydXTO1MbezKfJQWAnZ0C8MlIoufK1LRU
cNzewnxyzZT4FFrzplpSQTlB0aPvxElpaovYMWLFmS46C/GtX+q6RO/JuMKhOZTuzrAuW1dJGHXl
ay2JGdR0bV8Ov7FyjfQNWIcu1TV4V/4tEaA7oDDmrIuqxBsidgtuT4Sve6v7FftRRNTgeeDp0R2/
fLdtWMFpd40vVV2P2GIB9h4pvLyO6zrP0UR6jrm9llOf/MJg03F/efRRay2PtWvGvIIbZlgMXPjE
X2l9V72NicD/BH0UoJnZOoEcg4w4dXw9ETRP3bq8QQvIfLs1XxDBgp4VAgqvlr090tx4E6JjJGUl
e+9S/V/gh32vM/0O+0B3ibFwVa/PYk++nghwiL/uPjAZp1bdoFHBIK/btcfbc+lGJEbP25Fk6LCG
SvteQPy4J19QaBHWpHUba/2rE9LVb8iRRC9d0WHn6wARGqbobhsBpQimWkQcozTzu+MrDOOtw3+v
cnAunho3XzhZafp8Ap+YKnyaIIqMsDvHzbGLzcHJ/f1iOzE7aRqyYSrEK1g5F9QWB5ZZV/ZNnke7
tmHmvrb5rO1NtobGKJFFt7xpQpR0Cb1EZqRf70g9Hfz0mUTEW4SuAdhYZ7nHu1GbRQcTJOO4cSTS
FeJD418J25tqbCMaTu4krSOetT5AJ7xdv4RVQ6dR0rC69FRr/1abfq077bUA3IlPCN4yfjzDcr9l
Vyt7bGn0m5AqX2gaoo9YtIhALu2S6I/eR+bmwvyYvLSyMhs7Z8EiD0KpDF/bZicoXHKeqjAe2ZU6
mbDt61wiBCCwqWJ3BvC8b7PdgFUVoChhyB1N4AaLaHTuJsxrn9zWc9ia+2JMeVIpZTmd05U5t1rI
f/HG4E3lKRp23WRRq6gFJkeRpwN4EOWMP4ekYALFN0fMiCUiXLZhxZC4Q7ki5qCtg3TuSiIrqjTf
1Y3UmGuvEs3Nx8AH9vfR5zNcy+tkHgEXOXUc0uA7BZT+0gjcA3CcyoxmYWwnihzezaxG2GPsU2CX
yS3CELm5sh+igHnaeTElfy1HybnutM4jTbfBuSj7HJF8nQKLh68oz8VuXToD5b2gPW9ReASKf3xW
z9RZoKSM7h6IXEtJuapZ9LJoFNlHwEi5r8n/guVcbJUOqRbx2GdWvqFiHzLCzDWPScMa9xiiNV3N
SpiwWJLP1hwBYvOyos6KohfvocEDpI6LHxyZ5LZ6iHUAGFD47urcdU1Xtw1Ae6sRNoTt0UJ5nLVE
F4UEZcHwnIvjzdhoykQHYpSorl0OEyjrwFDaTUkh1NfX8DvntMRikFapmZ6LUaYKkvZxiEbTlcwU
oSHYhNW9uAfBMGIsi0veE0AwFPZsYObG7P9sYDhXMfe7pizASgNbWcjFoCBUyNB4yv3ypQZVoerJ
/eVH2CKcOguQIZSDGj217MOIoMJbwYVEwy8Yz7dCamkX4fPIr27Hel2PgIho0m0pVqr1uylAiRd+
GGMTxoEe7HxFzEI3JeS9cZz3y+8iDYpuYA/AsyFpudvhMtptqy/U8eoMZOm3dDK7jZFO+xvGlhti
zt4cExGiLyMplk9lXQUsVPS9QCZzzBe6DzUgUdZtA7yXE2awaEL1kjbfLF+Fkhv2liz1P0eDUUHF
MzYkS3O/gZsWjP0py25Fh5IwL8IMJRjnjJwQQJ6UD3ee+roG9Kwjghzi4mnMafNzAvx0lvM1qKCy
lWQIHO3+YyEhRnyi818VllOkZ47blj/uNlDFrHQFR2VIe+M2BU3VMnnv5rDYkeBJh5qEOpm6+fPB
u2iRevfL28tSpHRciNGIiKuGy+6o6FVcWVqtjZe4c5L2qfNnniHSTOiMMweN4HS0sPaHP/nwrRvg
kLj35vtAgLZdfsYm5UZ6FYkF2XLR+MnVhZ0Ux6A0X/EZq+8tcXAIstzBSTEDdokExjoNXqZ7KNJn
8jBNXcH21xpMHm9O1WFLa25c453BhHE5OQtI8++c1T4L0qv7yx0+xRG/oNzt+B2jOAkYsYWWj/Hr
4i7szpeYmydlYdDuwWvSOObBOyVRP3URPFtHmp7Ro2i8xEZiSQTmVQ1N7II9wt11y4BRo+oWwopt
+ElSYiqhumO6u+RYGV3ZDvrQkC1GjR3zzcJz2jb5MJfYeWer5yiY0AqPhrtZYnZfNFDYNA2aee/z
HjwvNpEqRHz7YaCms+2Wnwq+A0RopeUKXOp0MFB0ogco72+s4OEP1nXS+QvPUAH2THntu+SzmzWp
w7tS4MLR73NeB6l8Z+6PDZAG8jGuCiG+Ct/iwq6Mb5iOga5Rx70TWCBJmoPlZmKVO8/hwqNj+IeK
4LyFpk5M5AcO27A9mIgn9HDgSB4/tuulDGRrSSnuxDuqsIKHY1+VnwHMFDNZY+Jgw65ocrpCuwPY
qAPn+4UXEdwaoGklMYL/1BXGS4Ea+KMSNGmDgjvezI37v4M52Tj+UY06yvbO65YFHEa2Dy8rYDe2
leiciD/34+b2oovBkFewog7rn19ORsOYNutvcKxwDItxyYDcWB8F9vuZ6v3M0yNf7VRVajsepdgL
j8dZwGS9k0HBWG3ZDdS/xmfofeM0RzwQDh3o1JiaPJMf/RLCG1Z79UpiQw3KbR5/ignzZu4HVw7r
5cSLRI1o3NqfBpPxUQxw+Of0DdseecBaB4hAJ/IUMvT3BsAShjUH7FG8Ixr8EDb6MUqX4RIf2cZc
8WtRDUXJbMo04QSfAm5bsV/HYfrSZdTAO7kJlUk3KJndjX+Ibnp7n1CpzrohIFHIa8Q4ekKJC+Vh
7Z7XoI9X3WVnFeP8f8SOubsV/BnaivYMA3h2ezhI7p7oVUbXgSrVbuZF/5WrQKKlmC3ct4W8ISkH
oS5CT9o9uR6mY76AqcxzTW9dllfWPL1Brl0K11gWoUsA4Jj7JjtDIQTuGK54SHZ/2RBDujkmYw1w
fX3U3bn5lH4bBDjfyn/Ki6rjEdSJWv6JIoBgWf4bAfebOaheOO+sYfCi7k12unrqod0EOUwtxWWw
xHmi6jJzMIvi6FWHbYVpoFg9cvtgNnOuzs58aFShx7+d0RL3dOHyyzOrOBNg4WoU4CTclBcZNLbp
8zis+ntAWHl/Gq9tyauTVloDq7n86sfv5AfbQ8cSjPzvgl8Zo73MlHSOwl20AgAAT8n4nwOrpwwZ
9LirxJIvHh9SfSf+9IHKzYwBWVF8nSS9K7nQbLRrK5MSLdrHNj8wNRfddIaE1V7Mri5RMUsI9d0W
l10p3eswsQBX9Xe+WQhlZx+UZPbjxwdyjd8X1zT0+nVHzQytDgF9AMfBe2j+st6zMZSaJLwANjuI
uKWwHjT61uyFhLdZh7c8J+pBbvoP+Pow7aHOXS9Y2FxXXjhh8fJkSVybr9ffJn1OResShnRGhUMz
5cVR0jRmzQVnE16x17o3WjuY04GYFjIO6QwDpEH1ETu890ncB8TcFG+viuGyVv+FqGUn5/HGvrAt
Z9f6Qwgs5PCiMacLn84G+YVSPmNtSMtnhCgGZHAcF6pnFObCypmAz4Vl/lIljYQtZnhYwYRqjxjk
1G4X3jCMasdQ99diRrG0jjNv2mhGLxFOZx+hr5jmQ3C1Z2EQPJlLFyO9m6rkuRZ8xWkWeZA2/dFb
SFa1R/h1vnU7Kl3PscD/N0L0YU4iw6QyBq2XZL3DzNGHs0WQsuDPi5e8XGr5y6LIlknOwfeGOBGB
VYcVoPEzHtqVE0OWvhZYgnhEGoAAFOT0WCPjUPGtIO9Z3pZTew1IlbNg/4hTpCk0KrkAg68NYXgo
hCak/Y0Y5VFc3zgDh24gYoiUug7389oLgCU+gyLu+tr3ltzfXb48SS4U/bfrjPHLlrIeNN6daFYb
4/WOodw5a4PwZmr8cM5lahBEBTuCGs+zFHYVRqjBuDx0M1C18rtIYp6aQ6BHh2UkyDfQduYlzhBB
4tqMmrwaZzcg3g7eipPJjQBGPmEQuOqK5qhYezaVKumimJqPOkPeXgr8TBCHo3awd04C5ADaDf0X
aeBxuh9+8bSKcqkGNysHneOk+Y1BPztvyGZLuOSBYQUmQ+n2BQwV/sUmKVDMean3szy0sEmE0etI
QE7H4snRb3iBAEiiOnT8QTNARiH+s+4rdO9m8XMeC2zd2f4PF3J2vH6a9oey3OZnmM16hElsx8YI
QW/zm44HlCRJHNpB98f1qXBC5MlGbBhiw/Q+1/xk6mE0VyJ/MhBMM4u0tfoOreRZK5k+2Dm5ixCn
ndCAZXwZOKKCVZT9ET1EyNyt8+LD1dvCfyMRiduEAUt8pqn0h/yAFaLi/TZkZTLUVWyc0s6Z8z9k
jVJPf7h5u7KTfABGezI9LI7QsL70tFhzrbV0aWA/gh8Ji/x61Cybut2axGedEONGR1+npA7xGqlg
cCQsJs5OrkYSBN6cEQ8J/ZJrAk5etZebevnjOxOdkTaJkH6rNOo+xEEW0clqYoszP8rGbfPxkCU+
44lTBXO9yB+KmDBzysUiH/aHCeDP4/5DlF6UTEGVYM9K/eu1ATkYaOPo5w7UwqHFlMv54Nom8mUb
3W/ct8pw49FtA2F6b/SrKm5RCX/IDWVzrfTtBEloXykEdqXrU1VHesiSmzyvoronH6VeMonO2by9
pVFmxhfsW7zT5oHA0G5vmsvte0XPKcFKQvOSaRrQxR8qVZHbxtBohq8FlZfBJhKjEHfy2bYd2n8T
KKtILZUBPrDmv8Xbpc9qiXdLfJ8gC3EBiDZ6JLdoC4jb0rr/e4SUGqPwrFynnXd6/XShszI0jCbH
Fo6GM4WZZ6x2vN5HPAYof2B2dxWDhYAVfHyjl0341RTdZd3XnrxiL1v6uBTBkNGfUJlSFZ9nqDcs
k2+Umu4c8ukzfpd0ppAm6UL4tclHkXDDlQSguETmL22ITGa+huRxigc/ei4tKH6ebF1s+jYoQ+oM
ubnvHoIfagVU6fSygn5ocE8TiZZS6SaPgLt0OTeTtOyJKK4ZQSPOEyjArwiz4UPesSQshyPJ7KZd
f8uSHJfzb2HBipJCMGGRjVMelHyIb8c6uJeAfrn6Q441GQYTOPbRJay4NNNmFvnPuWjSDUbKXovd
Ak++YGUVGTzDIhNSTaKcpLLClxT14uZYrra6uQlTLrvfPNMt7bF4XGk3/u4CvYhGJDcWoGHptQ7/
QK2FQjNojTvfmMJa2EkOIWkLx/SsjJ8bvLv65zHdo/Sq+4fUVPJWsM2ioio/6BPOqC2I5pItxGcR
+tvzpSoi+lhgD2CtKLFyrrayXHX9sUUnStyYTpXDAeKYYY2jNUpDSqLyClMm9T4vqY9rYbrQGXEa
IMIe0l567X7sPjKijO59rfikvwnuLmbyUKnQbpoqngE/ZDop0YVYC+Af3KQThYmTKTURqwmnDzPI
mcwJv3DmI3FDEZgCpKToikPidyONX+rTDj4SibMGHDNYx3EsFITYYd6K5AAd8J/H1W+LnwrNCshe
UpHr+EqtlrM4R6T7tt07/s9vJOVbHA1Mqf7xuYEUfjXmmoDgZOeo6jQRhcmsugpiHyebI87oPYLJ
cnbq3I68JC+2s8ee+x8Asr0+AneAu5d7HSi5XfLnSAuyPM5gNC4JAmiJ433y35G8ZMIZbJ8aKq5m
YWYF6X+rK6Xvm90/niasrfzsKsQYb+j9MClu+1liCzGa3dDk62BSckX7VrOy46rj4XsOmD0XCjlK
765jYLcG4/jx9GsuhlMw7Je5BrB9vnNHwl/9FBYRnCYgbHMOe5FbSVQnPzGcTGd4PhVl1iRLcWFm
bg7h1pNDbh0uQtG2Cg1xtzJ9Z6UE63/bfZ/bVOtAtrUwiEv4YBrZLXK08+uGAuO3SmUcve2gFmO/
j7iJx5M6sz1Uar2+MBjhXygyO8qkAqfaxLoNLggyUDOU+LVbUrXIdndY0+ALgLBpeFeQeID+Q8re
61m7aTmIjMQxhqfIdR0/Gpu3A1yHtUfErI1yuFCHw7Bg6PBlk/0LU35tGHsNOtOJ4khRtHULHBPU
maRtnTRvyty/BIoeQnQ0te/W7l7oaYcifwGuGwjC82bKyh3Xxqvyvnxtzkc4VzlbAAMEUEGEFM51
KPS33F5OD/3tJi/LzNj7M3ss20uJq/aWEhBpeKGBTkjHPN8Vd0BXOdvoi7POdqyWy8wY/zYz4ZVq
oAZJUt+vJqY2dqkPnnZaKe0RHxm44HpJ2lpN62TjOBBL2YgqQEcia5j7k0zUJxeMyW0upM142wC0
35VpwsyOKCY2+EhxVG4ZwqGqZuqIgtFWNayAbd6q9+wTtM/5QK30RBAiqdN6v6LS8gNIMK90w8ME
xNOFoTlv0gihPo0XFjVAEhdCy+kxW1yaXfcpXb+stQ9BN/diJGPCfSWE5AFegbTCQ/Dv5u+XK3pQ
QcKV8x/fjCHfzvJ1C2uOfvOJQeA263q9YhUPbUB5FUqYJ5EsbcxZBqUKcbA/viX2qO4KQE0OnXaR
dLgVoqiptaBVR85BNRNXYAV2OVFu8Q1ivD2IFPIwFagEpJgzSfRWmOzZ9+c4UlzaGbvIgio8sd6P
kX8x0kqWgnaHLItlb6Z6nzCFK2odrYJfmWhZDYAklCzSUZXC74Pnmns5QEO83iitVC/JQXDMC2mL
g0NR3Sr4KgDp94xtRWwlIXONKSnYfKy6m6c+rl/2GD/VfUWen1ZUJp3vMVlW/WZemGmekyci8rMf
IurvdmKQXyzl7hV4h82zeJ7NjxUm6+4j/3VYyGCfrOc2VI6wMtU7MQOpKC9/diLo327JZxRbWaez
1RAWLT5zH/edO8Kl4Ncup7H5jnG9U2oYfKBD9MvVB7OCQgzYvOWK/4DW1N73RQr2QU+G77poAcXa
SMeJNaOIy+rnnhHjOL8OrXbqHl3nNd2IKig0ySFRdhkjMClq79ji9i4CnU5FTMLrfpXwiaBBimdS
CQsAlMVt/JpbpZ+sIoQPObxoJX/YjkQGgvCiLa0T+6ehKGuTlGaBYcbMvSUivBPJSJrfkW3rdOG8
VUJhO6zbzMclBEBDUcX/ScdOcWP9TdmyRyYDdKJmXP3ikLNPr+/SeLOe/94BXXpP7rfPP9D4R/cL
Yl4wU/lXydw3Z1Ga9Mrha946USKuNRcE6Jvf2hXKjjz5d88goh9A96WcZGCt0RrzmQDlLK/Auf12
c7iwPlFXEmRCR9fb5OX4KkY2QPDhDb9LIUpyNpg1IctWq2n4Mm6c42lZKGlGZkWBnZlvPqadLlcB
ECj6xoQ5kXvq7UmBcEv0YAE97uVrIHUlL4dn7wYEIssRID/WaWXoJtM2tFer31tXdWtdpdLsdr0c
Ut9GvUpGuqxlSFSdfMJQ04m5iN+jfA5sFtlutZVuQELnCVJnsq5pugJGoS+ht2k6LfaQKoQFRo5s
2d1YSxSP6wgYmHYlb/h6mkZ66tkyD6OvM1tuWr1TtazQjObR5OoWpxzAeBdchV0Q2BSS4B6EbShF
hWeflEkN9z2zNLZlp8mRExV5EXupJptzcUew0StSf08xBBRCSDinucvTwYRCvy/zV95wNB0EuQag
0LeVPMKaoaOLGeWKTcguu5JKwJ9VYQz2zDF3ukjO3ciWKGjjChmfB5PmVmmHi2578CEN4GAQisSU
A/EQPJMVLAiw4mPq/l4AEeBQW6PCM8mwnJwZX1NzgzhrATSIItIa5ad8jDsckenC4ef6EQSXfRiQ
2j7k64LzfTEltUDkmyOe9EVdLSTQU8zqTfxfXZUaPx+Ly3Yct0tm3IEpZOAyA82eArS5j0CsdkEJ
yzeBEM4oqmzcKFkFzE7BQhpsA842nC1Li/KA08ZyfDg7slYUWULqxieQ5oqKJZgpvuzEJsatZ11A
dJ1IoouIQfGLOy3fhAY5enurtA6aFDGVK351PQHt/f1OiFo9M1ou8UTM64CGLQuvHGn07Ys2FFfH
uqFlAWVrfnpJ7rrH7NqukzF+Alv4s5JY2WxdD+z8ROr0ndUIJwt7KmKhUnMK0GSuYuuOlXkT3PKh
oGNh9GwIO9PRqQ2BI6PeJiDK7yjrJXBZU1W/rsvVL/jc9CqpGypdMyKkUnEXH5y89V3LRXGGkOU4
QEbIptk38K8Xn/ZkorIDpOwTnbXHJifReBRhAjjFEq+VlsLOBFb9nT2rA/MjYLvS3417xDnGzck4
GhNsG0slEnJptfb3BkYj/+/PvBvZO4nrE2WTH4/tO1iUQSC5NhCEJQusT3zv9feqcJYxJWc9ojvB
HqKULkrs+IM0I/w5gTDnwnDFjLlgynh9c62Qkj5230zSpcQeqHG2OhTkmuvMrv+L7j5zlBrQI8AQ
4/pgwYnJQShJsr67lLSV0E/sxIdvYWm+Y6KSVCeYiAmbvz4mq9Y4G/7SownuCwei4gcAae8+9CAD
fXFco4vwYXXWv4MaUxgRLBG8S+LN4bDzquT5w5A+EeXN6l/hG0dMzsLP9dCTB+XCOkBFR25A/iIX
Vh24QpsZTB+Jw+fPShOGl0U5O7xCKrwVzPmZpy3l3w2k661nlC3igI0bHFKEk76p02Q33j2Rcubp
WDTOUa3NwloLnsPHOmYxppb35Mzq/jYiBN73zr2A4nFc/NG5AcUpVO8DgKzme7HcOC/8A6zto+zR
FHsRU4kHgUigeP2G3RWo5czNcQmdh+EQNSceSsIfgNs+U/FCycgKxojPaf53LvKcZrL5ub2TnQTB
cpIDsFqoto4ElSACJnfshGj6j4lugp62JeLw44Z7s2OCfUjms5o1nodK/2u8IuAaARhUHs2iVUU4
/IHZfY7esgH8sHQBzVSl93hoJES2yuzAxclfNW8BFWybEYQr45HXiU0fq3ctsHjXmaHBmm03LAQj
Lhv1cJUJG5LuSLVIUlFHmtEqpQUiOUBTg+pcsCK1iAb1tg+tP07ea1D5NDx4CHlGSTvoyc42LqiT
HFlcVtX70jxwefBFiE1a3uxpgaBT9/g1GaDutMJ7dP0hNgGC4RZnbFIkAi0YJUdG8JEtK/Vb5S8w
twDW3/TqBQPcPA9s7RrWYU1qwVEUQnRoP+aF0GIs7KzpKeL+cKFJkx+FFt/GXYQS/X29cFaIw0BU
Ogbmk6t0XJe4hazsIGvvQVoYKNY0GxYjpMW9RRqjtVaSGpEw9GXbJ/+5oa9gKOm3TuidMbwzpb5P
6mRFKW+xLE41Abp2SqTYpUAsZIh1z4k7j2i8K6IqjwNRZScuia6Yo5PIg6h6dvv5csaST+3rWWxx
nCsdd0i8Eevp0iVQUp6lPflLHe8je0jJekx1lPn4ZiMHBrNM59p7AxDiY3fxIGOkkyAKhqkHIKQV
M5sLEgi2B+4rOClXgnQz9aQ9Rs84oC/g85wtBOZiH1CpGMmtevYoUlWVYc3Mf7KRN6cCBSI4gqJv
DQSGlzCMp3RbSXWuQrCwz09gcBVMpkj0M/aFGlG8jdF/7T/rkxlAOHe7fyp/PqS7ao1r/yBm5moI
i2UR3c2lwN/WVc1y5WxiZ0wxmejREjAJRuS8yIUh7J8rBBvZs7vk8SEKEq81ysnztZajYJGmstTB
/wqqOtWGMvIAIIsYNS4ZciCy9N4v9T/+6D3Kbgmppp8mnXXXym1R1Cw3xbW5gVYnrUsRLKdLA/kY
NbfL/jzOLjjJ2iWR7rQzAzDT2uB18aZotvsoB8bOqGGf0sichC7r55u+tjCnihfubjo4xyLLjPfA
hH4LO18KlvEpH2e2p8i7/56RXq1uRIA7eRH1QNBOZiTf+90wSXqfm7Kd81XjGZ88GtnmOEXQNNTa
bRry9Dnkw9L+w2+BKbYh2HiI1gLQJetRhEi3rAzS9RFx4GBFZ9ekPN42QdLmNLu8nlWVohaxuTay
sPUaBBqxsL9cjG3G/bY3mTRi7Wc/E6MHOlT/ansE4RHgfLNk05zDuoRf/log+DNaITkVxwAdSivG
/1Lll8/pp91vuIZV9ULbEM04nKS7v5+6zvpNv+4dj9NuIBUkinrOlPsxbgqzMeUz14hMtTrMgXqS
69XERlZMip2mRDexyVrSxeKl3VoKG1nQ4u4Gy0kyvmELUM57bRcznA93kr7MH97rHYHD6udJrLyY
U4dB7OCC5SaqgportrxDbaHAaFyvYkn/tVxXT+nqidKBIFK8KpzOA/5jHAehKXDkMij6ZBdwGD8g
sqXwsli72OjuSuwvrXK2ZbRfE+Yny1WWvLU3fntnRLcdicLeJYdYWT0ucEJf+W5lF7aiEV7B1MMk
xqM1RAlhSlRGkTJsRO3hwmtauyH9v0OVH1CrS7SCMw4wRCFBSxYx2FqVp7CoY7mEmBeT0iKxyWEZ
9SgsIIBCR1iUPWruVyHJ67yi78jcu9yiwYUytY/gUVqjrflLlAK5gfARuggNEZCSqOGz2bN8cTF4
pWrghHafZwzz0VXzhD5sz2Xw69mcxZGyqCBoKV6muXY4xR5KCsRBkPrHrxTYNJe5VFFib1cMBLm2
8fT8a62Ia+c2KLPy6b8yJuuJfl2195T0sB0n30PgfZSbm/1O/jcfwI/zVvHweTIYZCJRhH/W0VUA
T7bc9G2xKn6N6Cb+VfnH4Px+eEg60utkez7FnwbVZOP//7Ss6EZFFXTgFj8205+sNoQ2GjQISLKH
+LNFRY6ARtj+GWrIQ9CU9Ja5iRz5vkDUX0n8dUkI/ns4sfTtYGO5XYnYTauhtEZ2zUqE5AdjH1Lc
qVlK9okpsR8QY9ZR2oxRPfTm1wDEQzO58s7SDyHeDPnpYg45aPz0HJnyOTemwJPEd+/hxtYjPHkl
zLCFX8Lzht063VJA6sxae/IM/Ql52lCVEPoxfEEj1WhLC6wk/TOkdsDBX9S3gSyAGXfHfDO2d7iY
J0TgprlY3SM9aKkxmLo3YijW1olibNytjGX7hNs6k9TS4k+dJ4TR4A432+3aGknyuXUt4Xzke7bl
4n+eetjKTz9qdlTjRTc2QXmwLszc8Z6QFATO2oWFT2S+cKK+v+zGIb45/fnA1UJnHUNMpIDRpiGJ
P5EemVid+SpttEdKrByr80S9/0V6RYH/UI5amCfvgpTVKx961UBNxsOEGGSjCmbl8qmRfRyDfXNr
I1i9B6wb3jkxdDxpClG09iZtfsurOgFNG5F/FbISH+GxaQj2Kr7zRe3el21UW9L34HY3Ztruj4Kh
qiYSLYord2ghbHhJrC+r7jjtaqJ6vpjxnxXPHKsl/LGjvvHBEPkTt0HXukvbFymG+JuFXYzAafyI
CvKh9c4Hb8FhvFag+tXeXKDHFVV6p/Dw3M/jtJB51ryBwnJvT8Tzj4qI/iD5F7oyaMgI0AMq6IR8
VNp/ZSsiLe/CBXcsCVfPJUuTYGT54gKQWQgw3ELFV5XjL9wzHsdtYRpA+Q/vZdAx80MvAtQCwn0o
k4ly7B/PzKXghbgUGvKNeHPL6aLiDf6Lu6uN9EQNTHu/RE9nrjs0RuAVmwaj2udGxPYt10dMwOm3
bA1XKvm09Er/44FFjGwMJ3oqIEcyMNV7SG+RiOFTv04FyKN8uM7zjVdugSKUdG7hTKjzQzEHK6/M
t9s8hsgnCi2PA3nDRMuh3obX0AhZBL2xvbc6vwhI/mlpXAt1Nrjihg5LVPIbp7mxvw+XEcthnFHb
A8k8AAkcXXTfF1ucOF3DYao+GMYhPc0Z7Lp5OHGMIRM36e6/4Y0NV2aiIPQdi6tEw7wx3phsZiDb
Jp/l4jbgmnTFsjREGkxSShxk4WD3ZhzU06ys4HZ9S2a5TyEWEeMX8sQNLLRbnniXf1UcPN4YRu39
W2jVNwA2X+I7dOj4qedMuoIUn3Kz0vgV/XOXTgZz8DSDGT2OcQS12UbPXkBnIKZuqqPUtlHgD6TJ
ITalvH9s80lrRR6+SP3psQ8jD+ZjyborRRbt7U0zgXcmrqs9Z3lOeGOg4C/FuhT75uwfSiraUCVx
oQzgaoVg5WYW4SNcboHKpdhEG7snplKBV5Az+1t4AYeExVGpzmgmk0WhYqid1cIQIw0yyKKbPJo5
vR1fCSBYa1K/EkeCkejUzG/+LtBgi+833H2apLeR/mG8ZyaG0zFpoPAKZrhMiyIdcSuGZhG2QhP2
6ImMgbcB0dxQDqasywUHmAzLturERaVUnfifG2LFuqseiRRTHYsXT6ddF4X9nMWPI5pFRGi1ZAYD
Vaj0Uhx0xkyaDe6pesN6RoAEldjv9QEsDafGuok+UvDBgBidwF9ZejgDURovJ/lsFp+Dd/MBO7Ay
2NasjgMLPupHevAncZ+N47jWSJgbH/2rEHY48Z1ctXckEwJhHzzjNyyfWPW6t4y73w2+G+TxsbEH
4Vh4er1EeQkXavjDly0hcs8Nlz/VuYVk7cIh+L4zNZc3us+y9vGkolxHlkaSGqmLvQbZYCGlnyII
TA0On7lJVUJk8ZuDATv+X3Jt2ULCO8MxR8V54UqrL23ji3v/UQc/e3G/gwkg3aqlXcs1uSkqoXgm
hOCQT3AVR/lb7D+fYD+l/KZUmDXrFu8ZIfTEBVnolJhuvmZxdkdz0NhjoU/b0/NrgE3/PkI7HF8M
bbEG6is7B+P84PX1r3Bz2W1Ix9rA++q6TRqEo0/GrMf5+yE1MPEFMQTDnlyks3DmE/hrqJJPl2BE
yg+oms8zlnjkPZeYenUtSCsmwkBVODLB3bksQB7adi6RuITBFhaVXGKCMpOPDzF9khd4PC9VOm9u
5DptoiK9AoyjN2fAkc6r+mv/XhdOiX2HlsLJAdGqKTTJD54ogXhRI4cbhCMYNoLMlAANQTZoUl9g
m97pWXXUQnvHS0zoBK6k73dF3odIoE1AbPB+PME0toEs2T4Pjx38pTJUDgyvigHd+s+c6QDqOwv7
D243Pp43zIz8CTZNfZH4/Li3CS6JAbCyw5HnIgGrffIPyST1iXC8QYwbx+aLORQj0XxOlK6nUcxY
2UZH4jwQBHyOFSuTQ3MVIr0fYXEJMK7s0NYygYN0jngp3F/w5/RY5Il+rn+d1EZO9BkR27rtvQKT
Nn+9jIj5Gku/4pFmuF22tKBgyrudBDLZtsnXevePR/x5a8d9hFRWio2OP0F8Vbmb3NdcDh9/g7uJ
zrr0nS8h7PSh/0fYVW4ZrZon9pU0shgCa3xVJFMQoq1LonMcXCylIsecuWrK82F7Na/4guFVBAAO
bqrbfoswF52oLsQY3aX8yLlTJCfhLEznf0azPxRP7c4FQI1Pu4kKed+gIrWxgXhWOlRJu1hdDdIl
JejmE+sYJWcVhbnZQXfMuWpvveLcw5XFnkLe7eIa6hPGvSIHqm3A87ORAGoWV2+wQ/3T76UpCIYc
Ad+23TZoStWCZPGTdzlfp2hK6+eTOQkZ4m7D4LMOEE2kAU4eM3MhYGnGedrl5rO/zB5xiprCJOF0
HhOG0Vb22A8VLGlg9VKJ/Iufc6e1xxsjMLrbAGvkmlYcvtye/nFDj69Cxd+1/MxTTh5J43zbHCHv
DZX+ci4R85ylm1+HlpPWgP/vzIe+e3max8oY7UPxxoy0VHFqxC9iJQPxXqwpSJFtAchp25JW92zi
67tUdgNVPjAw66pWx61lN4wGLKdaGSyE3rATif/5Jgc2iw74htS03aCCHyUsMLCaYXTg40zx9mNs
cm2DclEzml2jdLPqfeN5dHlhE06eVuRp1e5WkybKhjSmhuug2UpOwR7DN6a0etYSCSrBT4gdYKwG
83WQq7R+WW9KJrVwwk04RoRH2M2UbhHl/jTrhu8y1qVUJV28xBUCkOwX6AWZCGI8PlDJGSsbOra9
SLJrbI4cJSObOSrN/PI91et14lt6rgevFpM3ZsMFBV9eEdZU40bkDfeTJOcAXN5j8va353axgWPo
5r6mwVzupvEtAkn3Y/r6/niLvHzy9Bv97ylQTQbviiK4kuZjDGRaXBzgJq2R6XjAcp5t3TVaWIfz
AsA4AVAP8LEe7GqDLRsuVCZ0O5Jnaedvz+cV1y9fArI6ExpzTeOEnTAjCMlh9c0KGse6UnA5xFH1
R2266Bjl6nVQUgdzfB9NGodNzDipXTH6slufHXfKEUfWwQAmvMrx0LYsJnhTkI6LhxC2gJhyqn5y
X9iSJNyGdboSot3bVjfJzhFMUSxH2sSDVZNW8fs1KCi1hoB5/k0GWZt3+DRNAbflwz2Xocq7TJRh
Fi2sfwWf19evoNpdqM+EtMFroA1gXMvh9PqSTkIiaIfZ8DFMbWlXHzNiAT/R2ZogKldAUZ9S8Lna
i4jUJOHzkLeUTsZVwV3CxrCUEoyRA8Ck97VW9RlS5eW0/CqUmU+842jftM85lUCJBRJ4Do9sKVBs
e7iQToSfo/G7Fls0hwGaTYS4cwvlNFsLoZUatSbqyTFjFoXkXaa2ctpRQFqYLvRk5qpfVAzoDDK1
m0vW90dWDQa8mpicVVkfAfIbSwBixRcWFhwmgljVqMJBQ05upCBhCPuLrKcKTDBE0xGl15ib46Qj
0dcG2Y/xKRyNQWm8F4aX+TA2heZhLHAF2rdgcI0w8L/RJBMr4ZYKTLeCSibTkcfsgKgq3VPgHTnJ
BiibulssKxEt3V2lq/KV6XsPl51aOV17cyZvYVNvusvAU7P+mUY9ByTPImxoh3z1NKi37X0uP887
LcM7q1G8UoO8N9+a3XtIDgDuuQr3/ZCsmTfqQl1969pUd6F6ideBizz7dKzEWhXmJ969KjJh8bvY
3945/AHWllViOlSJq5wnvu6UCyobjMQNPVsW9I9PXEHV5Ps7y35XcwC2eVuYHWHL7eqSit+S+uX0
VbtQzh5FDJLN/aUjLjVO65hMM+7nxLsGYcqjQ+Mkb7dNZ/zGGOtdpsWVYtIYogc9wUuW9I59IjMe
USzp6bxmwv653qWYEtN2FsflZLmdp9nVHPM6R/nYyMAHhyX3284CjD8rjZaSVMRD2SLQ3BnGtK8L
576OIOXiB/dv1SXqbvKCYgw8bu6KggJira462aRFx4fjRCtREwJacAjtm/dHv/bPnKUrrvXbLaJ0
3q4Z66/Py2FVIGIWaE4WxSyV+HicFjLkqjAEvjwNEnvd7UgJmHjKp64nIlDUO/9fAZqotilmg1u2
jIopR+hu3s3hd7yIrSqb5C57jR1nvr7VwrdTBQ/FTCJIoKs3QOgP+ujfWfJRmOcXOYtFJeOdLgRt
yIPZlG8dCIvFr9B0AEZqo86c6764JAEO+p9efRZp1wJ5OLCgkVCVjW0ZdjVHF4u+cef8sbE2lkB2
07aZqUCRAspp+i5xVv10SiQ68OP87xSBCn4RYdjKIR01POJKm6Zr/R8mnUA4uIKkkACTDbl70GgI
qTiEWV6F+ocJXY8DlK/bRpqsITiifxBLxaOUxUAEiM8wzvF5s28jczPsqeMH4yksNiQk2mhJnU84
OMQlLMBTXKJ3T2OzRp1OFL7VbWFviT+MCJ8yNE+KFpzH86PblicGmn7xAxCMxTrfaBcQ0zOljvC1
YA5dbtPBTgUC6RF6kWEJHua2/FkFxs6I6aGnoZ9GjxNQlwZ0WUGE+CZB+8h7SxDP5NIoyGc6FVSm
cYjBnQI8C05tsTvqKnenYH4ZGkKml57hrFihIb25Clu+C+O9cHBWAziDZcoW2vpdwJ3YKVY7KMIu
A2YYOIC/y8UA1aEqmeqwGnQdVClvbwc9cU0+LGgbEyCLIMzAN+L+pEtxb6GJkRXBIryCYdCD4wjk
X33cyFIGD4vcjLBnY1SeUKEnDfam3+X81D/rijR07uUnijWag3yrnWsTmt2PwQXV/ffJhB60H79s
7vFlia+uIVdajZRTuqv+mgmj+spP0IZ+KLmmW6odcv0Rv17t8Idi6AQyn4oeWyA6/nTXrRhnNocc
rnK31yi+UdT8i20tdP8WF8HKPyDpZxHd7ZbKCfrYHjkeXJpgSqjCFfS76Zf7EQuQR778fRGzptdj
nNQmOboYVk4BcdHjfs6mkrPwx5eVf8+qfnTcfnanFPi52BF75ZLXCLxIXBJZcv//LQcDIYhUcxdR
Og6e2Mand6VI06efgvl1EyciWB02BSsw0kmnzErMdxe3vmC67Itwl7cHZ0Gi2N+Czd3HoDnwi8a2
tNnUwlbZwZezwIHad84d4onN5XzsFiGF0ZqrZFxCMC+QGfA4/zdVBvtffkcjTwDFpAGJvvZIhLlH
7z6r2zYio5UlxqXRWMuMtalZVIwKLVzIuG0X1WaiUPBXW/YHOCHkBdViJNjHZ9C/gHK6MhU59e9q
3KbYD5S5XCuI5VTtKHS548hq5/TbPnCExcpaPYHllywG5Ay14Xi+itwS8Fys/mnemd+L1AB697+u
3H/RnMfYVtxM5mB5/9kS/ut2qASTmqjcE+RAbVGoT0346+1YeMbKmEezW2CPuYs6Aw8Y1XO6XMHv
ZUjGc7tedMMbx/Pdar8kn+bbCCLuNRHw6/koBcK0ueXrV2koT/axNGFhl5dTRl+Td54m5AZnLOI5
96JXjBfDpQ4blPdQp1EBZ50qKws2huEIgNuJx/OjbJj8j5+OxCZmj9Max0YdcgomT9iPki2g+HPa
puOIS3ZB3IA2kV14/CXudmFGHgsagr18xk2YqxqO6PHbWoMgHF5mnu0pSVBxUwZM8pNp9lkTt4vJ
V/VfySBWHj4XhPSDbvCN9bNkPJ0pRmvzpiSqp63L0LE3/JzchGIgVKjWVSIh/S/GRw3fMa+wo4S9
baULDQzibVojVuqm2I1HH1EqRtI0fCjCsIoWl/UHOgPlQ6TC1HAz9s6a28CnBA2pIb/puBT2MuUJ
ecR+U8x5E9gvlbvHMX2kP/vtYC+g9ewfmr+6FXYaknjfBrfhoGHoq20ks0FPrP5NgBZRQ3z74SkN
IihBoIgxSMIzvarOz37hT7eDoDMPsqKi1LtM5uvSXLrUPqTSkPGdtJSbcbn1b5X8YBAlqrAL3A13
1W0wzwxqRfqBeDIFHaUPpQRsTWc20pQFE2ymbwUTQ/lkMCMhQudjmXOOKDIME2gZnEzzT/SIWapk
7rUhpDQDSrsAgXsoJqv9BdZO4CxfzA1/5XGxMn/3DnYimlHNavkNfxcEbpU29srmw5t2gH2QdBSg
U7e5x8ZOH+Y88/bDFOBSZ8b119QKbZVzNsoAcHoJP8bPXZLCZkpMizcBb5ynuwY1IsmI8EJlEybS
ZuQixBJgfWXs6lFszJqBmT4qknY3HUq1nfNx0Cyzof9tHGYu+vbXz3aTli314thKqfH3RM7ACHgE
Ez1N1nmtta/SRdzuPuh/P8LIAUPt1saji0uVRiUPHz0gQmBK8FP4x+lhWGRDhQbE6kYzJBCR1JGw
b/wKkadVYtkKPWy7LS5Pj2zdygpOfaW+mxhCy3w2vHVbEO10d7+V58COZNrwz0JqhO/zzfEOj7EJ
EcCJa9kyK2Hl0B2cgOlFc9blt+RqOs27vgHuugr7nC14bavSyMWPcev3giFsBdVJeZtbYCDmnhnt
Kw1RvQvydStJ7mDBQQYB1NucmCUVcB4FLx+P6/sjGkw3xnDVfuPakAzZ0oYst0D8xPm1OW89Dsje
EnryrOExRGf4llIXxfBGmZcSZn8+zQ2vBJgJndyYOjCD7ugO9AgGAjtWpqfoVm+3mu8E3ylAhfag
35HZ0PAQ/S5Jb18ArGZf4QW54+ljUDIrJ+lQZqZC7iveUZsUB/a9pzmWa2ZoJ3wAUgDL/zjMmyz+
ZvT6IXYmitkuCO6l24W6sN4YkMMbHXcCF8mRIa2okuE15lDXhWvJDCnJupw35FD0jrVAooh40m0K
0llup5Q0lpPkSzssxCxHn5eyyVG9zbO/RnZp/OK+hHmSiLkipC42rMfrbBGYFcpc1vL+CGexJ+j7
DVo40sp4ZMDYUZyusMCFhR6Et3KWQ9TeIZu24xoXHoYbeU+X118cJde/yphERixFR9hMwNKYvJXM
u/xXdiA5IAPuGw2wne07P/9kFsxB6VK5XiXJ1tTupZ06GZPPJ0w97urYtsEXx9Px5XfMaTcH8Z8x
Yk5vhMhGdxx6DRQN70pS4e6vlq7fM5yQzM41DHUjUUSpi1/i2d6+5jMsmvrDCGNRJP2nc7g8emVf
cHVsZDqo976hD0ZQeAz88y9PvwbS2/NBQpJGPkFr//WhO73B+8+HDKxiJc36KBgoNUjBuzRfQBDP
a6nPHl86tQXPk6uAyiDR4DdvPRKy0MmqJ05+C2w8Ul9s4hE/0tEi0wg0FuNjgYULVXcsR1GTN/sI
LufR5wD3HYs6vLAoRF/sO6DJAhT6p+xfeHxV+XG3mavt/hU8/rl6uOz8FKd4XCykckX8YIPZTASH
qoLI9jJTrI0xhBzyxWZQlY96nINI5hvsYEA4u1Wmd32ARkvQB6s8d7nJ1XzwbuzRfql7bFVYJCi7
JjZXqtRVWHdVPmItepae7/+WlZ9LVpxWx6Bi1WXkpEsXHdRsrIpaOHNGwh6K3cL5ll99Ii1WR/9v
U4AOZx1oIGn2PotVHSlI5qaxFRRbd9pa0HOX6j4oufGx7RJhG0lAedOsemrIsBOcU4pPatsItAax
4eJqlEJDBA1r7yPdrtIv0VvIxvhWZ6Ba/HSI72cT2h8ixay6P6wHUieWK4gtEzb/8VvQ/40tB3Hd
8CLLakNl7uHqli42vjM5DCJ3rnQ9DOU8ETpB/+D2ohvtvbZQ+GDRP5Kx8Cw07m7hSmSHpNzohRl7
RbHpfJ1AjMzCENoDwFzH8y+0WQZ66wud56tzC3Hx3oky7x6WSYkeUtq8stmK4WeOUu2fznymIpMg
mCFpH2+WV8cfgh5DN5VFmDV7kByhQoBNKD3gp72ROJ69CGnqLZVSZiEtNdTqhhj1O0N0zSp9SGIh
BY3SiB/30M0GysFjq0JficBpfVeeMi9COiey6/Y4+yqkJmBhUui0KlXMhkVHfc12fhmTMmHa42Qn
BPK0EdFWIyx3kMrFJJjputI9Lfsn23sXDK1Z9wutjTXRhoHUPNRfH4MtODPJasIQ7znjBaKRDyXf
9XNVz6vlUyCGV46tfs40HsflbwOmoCwqnPZW5JLqh+4NzTwWtaKk9U/HajEqdgMmRKvdwBjJcUS1
+wpLVoLSA3nZWplCKZtPJTwpGn7BcnK5z3LNIHS4gK0NloC/105RwSkZWI1kGGl27QYBOO8fxvW8
jf1K2Y12lNVrgUeHjtR6dPr13KTrXTJgfxh05YB8fTrEIGQnQx6ldYAPptfe37nyWkgPbDMEo4K1
5NLKCAQ2muP/dzuT8HSPJD7dzFZDJq3kA72qET3wJsdQ+HlvWlIrzZiocVwR2ZFOy3rpwuX00z77
s3DtMaaETi/9UMnL9D9phrforhIYO8falECoHkI1WNRNCpp4jlmxbpQGWjhopFunD/tojZ+/ntDG
29K4HYFdllklKDFh0GahIi83EsWVOY8l79xH/hP02gk63Vayc+ecxg7SoL6HCHLACwo9FJii4fom
mD9nyQDYYc7PBdjWGOqoZFErFUhuZzvgKqWOzomhHk2lIViZO7Na3cwhhK8lLvi92aOTHeBOWOC6
5fuWLbrBWhxicnuVDBKuU/45u3vEV+cdKccIEUqIAGGgd5gnM+if7tbspGHzQwkMe5WlcZtAt5WG
gPGd19iPQNl6Fo7uaRaD65NztqSBhMcL/TKqRjz+JOG8R8OXREmjpVz7OewGMwQ5sRx2YUYSwodk
YTLi1tR6KRuu8/3q4kBib4EB31SIcRXAxDGkE3v5VJl1UGoYmsJZVmfdQnwJrJO2ulz4hnjic1aY
WYkYSZ2BdPhELMxsvBJTwATGsQwuiiygL1gAGXsA3ii8Qk6KDCypF5hohaQWTu6kiUzUg34ccJE4
E80qojSmpV5e66csdvw165RRsW0kiX1TGcwYTzVW+CJt8ANdb7JjAPf3wE71kQZ4e/LPNSHBYvg6
xnuBa9pgL7d08GyTQY2SfNXJ7a5fOJPGUnfpPHhuhiby7p2Lqfx3N75GAAUPXxYqlArzx1i+31O5
CfxrONJIAWpK+tPAanZj99c/Dy17H5iqUfGf5rYnO11U18c3COhwlNgzO6+FvdZb3u0r8dmC9+sA
PpmsZDqZ2xfZaQ0Ay2UHzMh/Unk7L8sFHYOjeSkJRtuim2QHVseo92G35PsdUn14tEOWk7w6ZcTK
yP1wVNWSdpuZkCHlWBvu1hCWfPDhM7atR4F7dbqnPhhDghT1bAuOtKP1XJQjkUzuI0NxqNo2j20p
nFnyWf70thYMbYVKDt/oWg5LoY4jDniQ7TuxDaPWqz/sK3QbgF/oQrY2bN3elYVzpy3YTlYxVjqa
+vlbkhdT+K+Ei5aRGhnCGVMUg/DiiXXapUTljWlMqoXwStlZOMnVhV+gu58NvVHx0wnU9iX4/aub
VXGJWA9R+H1rPD4Cha6mJuQDvXh+rjlFRb+ohTu8MvHq4siLJxDeJDuvez1aiHIfdAxtXOPKLRSl
sX4X81t2zMErzatAPd+0/GQNzpMgdKDAlNybv6EithAFsBwmLZEHnRCSsdpmdibTp/NwxzJVyqZn
6yV9RTxcXvNexThRjaxemDO8Imb3vuNxzjsCGfG2VuZhOU8R4hjiAyjVq7uoy64SUp4u/6thXh9V
qox+QnAO/vckbhaqbDT1XTQDOoP/olO4/aZOAyZI0U2bqdmXz3+R5RoWLXAvzy0632sObI4XzHM+
ZOpcG7+aFZHb4Rk4nw2K+FwcYgdGqyYNPFyoGzHCT0QlaNyxgOzKE4AOPBf0A7fMsxG+1tQgqgSO
xb2jYmqZORHhJ0K3YbDqOATceuZUUfvJUOA5HTQ9aYHvXc/7FxDVNrJOTOWIV7AaRbdkqRKgh5cv
Sh1YYV6VGKFFEUy2OP1pGka5J5fKaFxQf8PX8XSGdDF/vEJjfSaFDvDy/U8tMRq1nknq3lm6mkSi
FFVxfr711W6KSjcdQpK240pHylwEUWDAU16ubxcobC5G8jhWZ+KYPxXQR3sDSu8P4dCXU4vvo0wA
yZYVsEneGq+6vQWigDeE3quzOBzVASAWm5iJxWJdXSTMZJQ4jEFcX43ez+69e1LKDtXqSMCpl7Fq
WCXwnh72JX0WmtONci3asTiV/3pZqQwfM4CNksPdGURbryI/PHG06kCfxqUlLtiBL4L5H1ZBxGJG
GdjIlUDyTxNGlpBRQd6qRDh/vLmF8TFsr3D9hfvnCPRBem9ewqg58hijRNYS3WQxjRri40731JDZ
usEg1el8dsQMGtBfMPWKJuH/2FuJPvkcjNsvG97m6aZGcaTNKUFpAkRf3PRrGFfrtxVgFLN7M5V+
gKJk11j8RsYIvSej0zykJgGWYZRvkHPKQle3qwHqeuQqwzLeHFUno2va4BoYBLLwAX4BDLcJFWhI
lzQcEaEu1b98TXMC75o/TE8SIekD8ZMfY/ylUKLNWTVglgB3rjGetCPhDE3katB2hGZ30Ax0GsYq
4hxXYioDxR3TMU54mh/7a6T1BxDvrJNafWcZofHMR5XcejAziSnuHAsnNPj/TRYAslhNqMioJXHp
XkDW/9Whsq3wJ7GAdpqQnstlSi2QT2jwjpjvOrecw6K/Ln50doqK92fm8CSkWTTdJbC4cLdPb7TN
jf3u/z4MXxiNW52O1AeW4sVucPoiyR7MHwyXCWwzkcUa/lnFtL2myZN6147NlObjZ7Rn6Fh+LakP
CnkgUny2sCXRLhrHOYJcLJ2QPkb3ZPQqwOlaBQvj/FYvYE4edVESSyqGuNt7ka0t0SFy1vJ1nTkf
FE9XbY6iIV76u+qypnooXjn7BmolEM6Axvz/asMmcJGyWLqq+KE9tygA4jrb9tyx92LiF+l7STt1
4RUD6ynjDNrVIgdIpO9qC2IUZZ4X0Utl8T8UIJbvJ1XCkyYMn5ev6AjDmzvCJ+OW0kZuPHgD383J
xfofjgBCDQFgwWDa5YP+JMhIWhJ+UC4n9C5vHnleyZHgqDy4ES+9QBW2wxPTNGXuOWlB7jTFui1w
4RW3lrnwVaHZeaohP5GYlTaKZaLlyiq6gSgqja8i8AOXWdTYcMHWRWRY6oY7kViNAygFSwY40+R+
glfNyHXXSFy4LZi5PhvuLN3Ovt1PfCa5f8pLXFo0yWw7r4fg2yRwJELcgnGdO42fmqIvJFihZVv5
1sRKxtSnl8Z0ma2vTkzBWYSK707tHCAnwCaIR5cK366ou6NjNc1vv6q/nLb2qv2WFkKnWiWxsY4/
97Zu/C0LgOwx1iCq/eY4szlWgQ8jnjIHX0BXxh8cNY7EtYZ+ss6jWnycCDNmaEp4bCDpgimIc0Zm
wkSJ2tekCV+W1yNZ0AgPBVafgK4tEEnmbpqWDyRqRJg/c8SuydWodVjesFVa9ZpJXOizMPW252c3
BGmL5Nir7j0GqU1Llr6e2gDH1lX98+l3NJRkSefaLzZf4PPqwerJu+XSarib44HxpmgGEZECpF4k
2KBXjY86zIRfdu0AYM54xrQ9rPpgv4K3vS7ODEAAG1UDDSeRAmMG2IarW30qkirMjBcKQGViwaqq
j9YVr6P3MV8ExWLIFTsI+hHYBI0Qz6+hqvexQ7s0zq9lyqngnf29D/SwtBJFJ2Skm+DsMnK3WEUM
w/4hLsDFfs06+MUqvZBXMl44ZxL3ssyW1DEJgXj8/3XbO/Rk9xbK5FuezwVP8mfMvMZuEmxyVMgm
57HgM7n3z57x+5liceE//guGszKAXfJZmqMxILnF6+o8dRFfqJ08BIfHeyXlt222/0RDXI11XZ9A
ha2nGRP4fW0dKzIJWs5zulNPaXZXvYHUfLQu/dvpIyIw7frOEUFxUKhkORN6sFZHW9K3wwez+hL7
3Gz+wkVS+Haiyd1A49WDXdab4ytInfnYMaiQMH6SneWXyginm5++6U6jHbA15bv/SjfMhuIKs/Fc
sgI1SvWVgOFANFUaxWDvLLRCYDNOH9lZsWRD5FlMPiUGBi4aVZPybe0rxu5qbRIob+cLHp8j47O+
/LKNfoDSRQtjBjhAZ857oB78VFl9NVpOByMWsjCTxqKvysXSTkEwVrjLwd6ZBc4ARn2PmcEX/W7D
v7SK2HetVQ+58QmUM4BIqZDBANc4hzNSWPfDg8ufpYjw84jZReMNYJTysdXrJm3jzPyuZmDld11E
6ngnPJG+wDi6b4J9NspnkeAwig4COWXj6rk5ybLjB4qsMMNYvM/fbBpdnOdJaSNXkKQ++wdRA5JJ
16QY1d5FhUFIsczVT1Z+uZ2SBLDwzjkzIKVVDFb6krbb6HT6ogOueI3fYT3+xO4BNEZqt60lETPl
UeJBlQ+4mJ742L+nExH7kgXyMQsPQTcnr0mwtsURUimXMvIYdJWnYyWCQSVVrJlqEZ5mkrT2rlv1
lMV5t8HsbFG7QxbdRZkRzM72lLn8DLYLfZ9xm9okHqAI4XhChsvD/Ei8/CI3xwsD1LVwUjkTEn3r
NWJM1iOfnCwG7zySlHbbYbmLPutXvjHyHgvOxa2tiMfdvjdoeCERf0FMkdxHnMgC5BSljlVEPfKX
dumdme4a/C8XX9BgM4hF2G4eRWvE8fFz/dIMwK65TwoEQy0RvMzBqCL8wVfEQVG+sxVuybvqaESN
XAgQVEqx0pBGFU0k/5WvTWBnbUGHcaxsHmwU8sNy1R9QmfRsZJHGfxgfLJMOY0G8Uo1OTTaQ9TTm
hsWfkeU5Nkly7DkQv+5tmDGVhQXSTM+O0xOlND0d2YaP7SIr/yjCf8yHoAcIJMNIwhtx95QST7kn
Y371cKHIo1TGlaoSKJY6dxDnAVBKmoWggS6drI3JzKQ8v6a/GTPwH/VpV7XRDgfaw/RUqfekxdOK
iB7sigc2Bxb5o+EyVtpuWhIhmDZfq7NAaoxPv35o1GxRSG+KweaFunB4lvcRP4rWVhDalK3Jbf0M
1r94r+16NwwOA/ToxWLC4/1CdPOR9noN2wqao0LST9XTmcMxoV4d4G57Fw54VgQftgUVadndHtf0
rhiAuYr7rFFJQL4Sn5ixKfBR/i1dHpHFVIfOjtc3KXh7oqw1m0MOGI1cE8g/n06ytz3vj+aPX0vl
ORmdFoLKO9aXW45ldmuQ7oVesRfbp5q/YH4Klw6jx3lzFYkP3xQVycWjJbEwb9cCEgs+9gE21aYr
tFHj+HgroG8qN1alvM5dMJKN3U95VlbEtxYgNy+NST2ZPTTqaLYIUuLdnF+c8gFU0bo9dh6YsDyg
B8pVh8e4gvyOjoZFVS7Jd26T2ql5UQgP4trDjlyjwTXisJWA0zeMgVzJNLduBpmrcbZYSqs/C306
+yb/PdaNA7BcZ75B8bbvKpcYSy/bdlXk03di5fAieaV85LtP8ZNZ1GLUaQrqTEZfGeOfk8qHG1/s
IYpf8/hpJ7HaN8ZwlWalWnY/5tKKVrdAvTYsgwi0sGh7pwHmJV37qoT7sjHBQqedGE9QgvwQ2OoI
ulgUa6U1FbX5ZY1Hp38Ao3eV4I4/pQ7sTdPUgMKpG9e+j1rJV0Dr7gphaOBd+PxlyffHH+gRql2W
6Uaj9yelkGAkF5KW3UKxthHJvKw/52QyrBCMgsBrkyb7pKlvYmzCeTk5DSA+lUJMbnEc/lmqdKYG
6n2EslhrNzPqF+QRAr4S3jwy88dNfFzjj8IP9pQqdhdR4DU78IgJNHU8rqZ7N/rRzbsixCSRvWEx
wZmc23RxhByK3J5JV47wHpaeXPttyotfNrueE+4JKEJddv4UCsHsc+zEB6jEJ1hFIN0FyZwv2MTt
R6mgyXTZ9ouThrY+mOELfLzbmg6sItbPtGcRWNwCwWnP+eoO6L5CbVKmTot+ll8tPetFh26or0tE
RtjN5j9EnQcru4rdInvPlayrJr3txlDbS73pGJ+qjXHBYQCME4rDPOOfmTkPzOxLmbj7y6Awg6fE
jlxVHJvMkZDD+D4fuOEtfij/7Ukh2gk2/F8dFoc8uRwmEx/PIiemMhJvqwNjatBbPmfeRwnQ9PNM
hjBvGql0ehN06iTFsB7DAAdKyOLXJDwDUi5rOcBrI/HNKaPdU/G6tcwphxW3JR77pnhMv/zavqRf
c6OEffp5gm7iJUFFkw+waS7bv7x+1aPfL9ht5x0Gv5uAvFVRD8OBODdWmjhzqMoO67MvWqkYWr98
1FC48bPa65UVV2WP57NM2bl/EX+PwRdzagPMoAhIHdYOkeXk9e1yOsflMGgLscCjB48nO9DVrDST
XhP6xj5pzu+d+EryQIin4uSpM+68s4OIdZicruJynEoWgxeQZRvAySZLPn7RQCL68sk5skjRSAXX
U39tOj8UrqNp8979BkJ9EyXOOK2gLNUW/vCMTMZbLPcyWRYgWXujU+6oX2QxkoyQAsC7IC5wjnGh
HeatmJ/+z508rvaSscHo82GtsjBRLDGglVR+NOJ6JC/Fk9njfLVv12ltcNly1KV6t0NtGR1N+leT
Rkjgz2WMF+1donguLDrDWPqeS7b+eHwIjwkviPyylpxRXz8HPSMM729xNZZxtQiixV3+G0fNSGm6
qnxkVNn+9cTe5exSUBOy3EPkd96tc/F522xHzKVGy1RqQlyFKF4sPk/XkMS5UHllD3g58/+Cmtda
cuo0TbuseX54taqnFU5T3/qgJ6L2On29xf7Qx4ykop3McDbUD+7F/QJY+zntadFpIgDeb4sOGeZ3
6Yoj5gkRnrxqINGbP0OFMGDCYHN2iBWLkpE3cJgc/ZpKc8mvQ9JQgKuS7mC8tCwi+Rz75LYlG9SG
tAcS5vPjyOxgVsw2I9oYHT6O9LBPYLWl9hkyxEqFYahjk+fURW5nbK0DBwawaWb143iZis1VWkRU
ipqJtBKcxWjroBNePpjKtIkWR76ohpLiD6qISaw49JU9eZq3ORPQQW+0sZzJwDfX1y+rrTTYATWB
+WZBSQY5XSYEHOazbDzTMtHEAaB3VfnNDODeWDq6IpFiJYg0TtWeq/W7BoQgswa8rf002EwTY1OG
OBZeK06DkLyI01l6gZi1TsVn45swTwKUISWxF1dlGOZoFi/XsbJEeRpt1jZiFVBwc9OpBXWl8Qu2
Tvs6ASeWf0yajky8HyTvDGANVJPj7flHfm+jYWxWHDxEDHUdNRWehln0tSBB2pblveqoI8NPqhNA
5s/lmuZxoZh5EAWQSS2dT8gTQn0Z5pE+EHg+4hhOqro3m3130wQE1HMOKrrZtWLjABpfCAvyR042
PJepf/DpuHqdMhD3PDAbcSo20cEkb27UiiH2l4xEfMVxqDgCZ+8DVc0jETXaEmKHa8UY46F+0HTO
QWPpWHpgieFunJehlpMoosgFLrlgeEwk+Tfj3Mn0wQDcDkQhzwh2TZjC8WvWuGzVAMLFamAc+ELr
y2o6d6CFp3NDL8aJPxSCVsqMHcKeyXhX2DWYLVqHauxNqQlJ0IVdKWn3Ik5/zI5BhkuZPaSinQu7
Pft4UwjXVniLuO4K1GJS4/DltXBHpPYenQgJR54n+kPjotMPB4Jm0U5sPrEIp4/aC/nwNaBu4vXL
Aj2xd9JXlrcO3Wm3f6KxHEqZOgoAAn+BBdKg4SKVDQ/HaDYiIqwiHPUEhTyK4h7m2CIcusMbvwQY
MwCE5ISHcNJvSS7QSegFh9nq/oAIOhIIhzaeWdMpvpJhcXNUAFGE4iwUDZqPD1ePAER3ae2cc+0r
YoWy/tlvvc+ff0+7rgpBYN2tOHASD62ZwgHAFzZBnuIlfSPPQGDFpd4V35T57BLqFnw8rU6vD0Uq
rH6fOpvF/Psh2+yJasZ2rWII8udX68ZnwLSG7cVl1VnhPYgx4P+q7Dut/gFraBm23cpAaqBqmPfv
Fb5VwcqX38D3NzVV2cLk/qYa6vu9bO6SJ0IBcCGOqpXIwf3dYPQG0egPHdWIF3N5/BvuDFtH3z98
u3WCuk3iTMrzYh7BCpz8YRy/LyAuVoA52gnHmffI3FujqLsJqNpwmLxgVkkN18SC5KGwiP7alDWB
osx7pgYe8bxuyAS/tnsxnALdmvWFL03YAgWanHBlpXpKFipMzLWWHVs1tjZv54YJfNWp61JwvCeH
QMlL5YOdE/MzhPLp/5YaBZJhz9kAbd2wyVqOQt1V7ZOitBLrkFoq8mzQ6omlX5IbabuFVuKO+Est
lBsKWXI5VBTmeDClWTey3HxG6BmPVVDCamH8LbjxAueJc4qYGSmRdCsuvWTUcPwsvGi9XoexB7S0
HYtdGoPTItkJnghKnKNzi98O+CWPzuF2HIqL0eMwcBSDOklEON1cSjn73c3HFmKsrcEUXTiN+gjA
MtNq1XJZB9sOt34VazMchN7qpY7uEnaak7+vWjJyIC57De3flU7CZgmW2hIPRm9uDgsgd4JIx9JO
VJxK+zb4b0DvukOsjc7zv+QAqRV6RsconkSQLe3tCLpyzOHq214nAP46oQZLWhH175ZO4fiSXGHI
eGlkrdyPSmwZoDSIcfn/cK0z1PEF9Nu3+UU9quiUPK3JWS10det8s+Zup8iZU14O2Z2eo+yGh2FI
Kmjy2/rpgXLclRfaZ3hTfvHuPTCwYTnRh67Od16kYHW7NbTTIMA0jOQLFmXZXyHjKeT+IZcMc+Zz
cCuTKMZEMdSQsElJM1WsWG5uJz5Bee7bC5vQal/Tae9pv5mYBBg983Th1IWJMevKemLNN9LjsDN8
/u3QAXuUg6pBzd3s/BOpE0YO4CdesMOAvSAj6m4O4jQ/LAgocQlhN3Y9247JxP3VUtEc354eJ/lh
nBJ+oXsMvGIijR/dzOYHuQaKJK9uF1ydSkFJfmwaLz+NFYzQqoZLm/cAkkxbu5WW5tAFDO+pNBLR
C18DVSFHXEg5CLjBqpVCl/6HVNQY2yU4gSrn8649VFAmMmDLQiPZiFplwFYXG0djwJMd09oNgFR8
E5dvl2q5GUUHIKC7OR70aWrdBuNMhkuyir/tobAjHZ5xxsKPQWUo649zgbKYD1ejOEjTVD0lVW45
CtpEkKfaYXAsCHDd1X/JvDsIzfWLeIR9nlIWVNXiY0kOkRxrX+nnqhKILPSFd5YxyuFMG5Yea6Ey
Vharwrf6anCLg1HmmykdwItEDXhrWDCiVe4WJeLAiXnNJqJ4/gby3KyvBXqdlpyXik4QXGxWbq4z
Z7x2cI6SuWYHaqwIslyzbMNRJbe/aDf2TPXV3/D+k71IFkDeFHz8gxUSwjbuLO+E/Xi9RI+oeogK
rnZN5LC7HIMHH3p6zpm2sZ2C7/ivQ6+q7WIp0DRTEPdk2ef0JWumHcaFJWKGvQb/xIlqujhPYiBo
Sh+ktRz3GbeLc2Al3nR+ye13Ch9wFusrqwzVTpsj5qTuyKCe/6T69z+cWksPx1kG6VAmvvMG5muX
He0vYs/MXr+BWZzrC5B8FmTUDkqgty3MZEQORC5iId4EooierIaWH+JNic2f9z8Xn9lL4/DSBhbp
+uR26rtjpBJp3BOceWjmhHdOiRhh3L5QeOV2059NSgXL1aytRFhCffqKXxBlpfZJrqJG8fFm2TEM
t4VuGck3kisrAEQ584DxE5G7uYfi5nPJvmyA+HdVqnATGOdrSS3AdMmaqGgdN/mfS1VgBUfasrXs
+xM7aSKE4jBwXyK7pNSG1fV83+rsP19/h8gIlJmPCaxZVWa7JBlLzaQ9rTsaap/Ijwe1PWKm/Dom
GOpM5u/gIzXVALatUnzwQ/EYP8GOEkpYjw4PIvICgzD8HA+dwsSRjgWqfiKVmDscqBC2qUkFVVSQ
Vt+4PauoI3uPXWaNo4+hW6rq3NwxN04qfu/BbkyFGweHLmnV53nir0afYK/YVHn+EoW9MILSMbEH
hnuqhI8CjKpU6LmNemokbZOX6pz4gbt0NzQumASd9/SZ//E7J/Cli5hIm32JsRJj7Tztc4Mlg15t
BzGY+JKIlvwHxt2tSx6xqjtuVdGGbOFOG1D78yXnPX4AOyW3QASgGTgaWuWvpQtwO/tqGHiHMhow
YZlncjQ2dtX2H/O/ywqLE8+8xVj93sFArlMuwXGoTltEsG/P0xfODzavi69iVHhwLiNezxzlq6ON
mj8/T6a8lUW4Fq9tvceIv0xhBkP7Rx7U6VhLuvkd1Gf7gZ+k+yrlb3ugHLHSKek45Ks+Asl/2bwq
EwcjBurzTwf05NR6jhRAm/Bm1fDlpgK9z8EujqwZh9V81ok4hqEEL+Wv0c47kF031TETPAAs1B2g
e+1hJMuKRCOSEX+wySHyhp7ysY7kK4moUJ69PNKkur9xC/oylf/O0sfFEZCIsmgN+bXNsquAH/rF
aotZlYWaiuIt96qPChUCXqooOENTyo74FdNpaJ9qG+xIhh6VcqDPb17nLQNEQXNalR3+IYZgqXUc
jRkliy0fTFsk6bHiC2XpcFTq9QtuPQFJ8om3TDmRyRERVKSWyFYqN+CBZAS2o1850ITfzkqYxmX0
tWHh/yh7YBdoPZXLp2KkHg6+87A/PMeVTTx4t+CNQzEI400eTjvjt6eqNtlUNKhOs/PXsz6f1WgQ
razp8kkktwQDE+1roSLgBWYoyJ4oKUBCa87vCXJ31lU5QxVR9fUzch7CG7uh2nLBvvBrUuELFWa3
e9syyp/dQ/j9tIP41FPNsX1NSoUSe9Iglx2KHSSPCHT3OLdue3mHJIsNCyXonuV2zYcSXtXuLj57
immVn/nz4Kfy0Zp1xBMpvbE1YQAY5L9GTY2MZKNzVKUJw5/PuNVTKK5d3l/j5SAHj3gNXDQegae+
Z40pMVBNbbnPerN+D8s77T2xBW+yr2KhqVAimQYy82DNLFm2ELHL+48BxS1vXgtj5h5secnENUE3
icziAGhNMSrgh0gHcXFt9VJz3vj6YCNOrm25UIClbMRnuo6MjwPBxqL3jt53RVDvpfcUp8QY77+p
ayoyq/C3pikh4BKV8k30UAKG04/FAOZgmSeYSOoGDWkyKjiQkL/lfBotWnOtSrmxR8kmgzAoEVV9
o0jASo9+UyYTIsjByunDZ9YqVmV5xdcEhVN1lc6OW21meDMvmBH802XDj8zZU9XaZCzXwbpwPWC/
0hdijsP4ylJd6iveWfLh8SnLWJt+LTQHroncXilnyXbC45ISLWxZcH3SKBvZHMtqSWCmrWwIVjCH
tpVYYp4OzFcanoUGfDmAAEub1ijRpKtzo5PRsBmX6Djb12BOM04HItYNJF5mMkNmT1op879E6UpZ
ke0VXVR10CXLe05EpBjxJAtvxl4Z+7qPb3GnemqldnREADtY2JFt+ms2vzyNHGOr4k35b4dw33AB
hiTfndhaU/PHcBhzFMP83/9mvYWl98VeOig5VGNQEKi2KGnP3cvzOpOMggsK5+Ffi1MZCjqKOtba
HEG5twvQlinl9g9oGyaQAwkDx6OGer4JwrG0Xgqv2l18+AMtG4RQnxmqvuGj9H34GCqDXRU0aadK
xhxg4iKWYBJFk8LfvFYCXMWKarCpyn/ES8Mu/F8YlDu4H3Lqpv4PAYdPs+DHpYVwEWxA4ghkqXXg
rD3zXY3uSRDzPpWO/U8zvD/RBCIStavtgjJEsS+NYtjeEEbobIXQXBUpIVR8stpqCWQTdKhPH2Em
dtxsmloHqT5Qe+T584qxD6IDigkIeXF8aRu6huX++c1w3Szn6OdN4NvF8O1TVHvgpcKBF27cjXto
xzddtwSVFqItXZd96D6V0u+bb0O4QqgnQfSAYnjSI5UzY2OLgk85T/ywOB7Gj61FXnwoLC1b6XRT
ybLvNuwdRMe+a66agOsR1kqQncDkIGYABhXtfwUr8cMG/DBd33l71/LulkFQ9KGPEMV6+CD3iD4x
bOdDgXb5NDHyIY9zMc/utmX/pfjbY2+a9DPPA9BiWRzIex4Cb9+T1rdEjYtGEW4AfzQeFchNey1R
iMyqFdfHYMyp5qCP9P7DbGyvWFEkoY/u4y5VWnMnRnaJqggck2Jp32XEGNY9esBT2/2HSyrdY0g3
TCH95p5N9m9h5sY8rl2t8qpK+COqkuVeOmktMV6HR0dTq1UwaeMCAxmSoM1F8Q5ayN4Rx6nZXrzc
iHMQmDeEw6pyj+Kdxbu7szNZAzSTRx5I0H6A5ulBnMhSr8UlLzN7OIFzdAQjWp5yzZBrF3se7wfq
7xSGfwz/e8pT98RZOfB9pS9+APNO+4EqIaANvF9PM+VRN/9tE1fOhhO7iN/eQgwvfMAACX2I2T03
vWqVo+5pFB/D61w5yDvCm1/w6EGMlT/B0JldIJmr4K0NuvG/bIzhRed8r/USwFSfd9s9WNO1xYRT
3pC6gFpOCPcEqfVFqZnK6kp8/MtDvEjmLtv8kozaTsslxds213OadO/dcyPdVmc6YAoda5FsA9CR
qpX7VR0jD6pFtsseGKfj7ERjIELKGtW6zvh5YNhxRohG3aVpb/CaWwvIBIVqoh31NcvVT0hfuoZO
k6A301lGT6iz/sGIZECAkLpfMnBQI0ig1jUPfFYhQ5k5fDw8Va868hxvmv+1pojZJiM1ZVp7GqEC
c3SLOc8WGUB+ifISiSJwEuw6STk432/KCup1/9GmpXTamZHpBv9W46g6WW9B0u1cg6nSiLFT+RY5
gXE72N/hkVswSt4QtPF+qMR8KRIxe/B82b6HI5ittJdaa9OIBvSezCIcaz9XxWDdbO0n1i/N03ad
joc/5QCskcdaJR4y/Wt1ilVDIx4TIy4/lfxfp30RtK6qt8Gzactl9hvSd3v4NLUWZw4sfbtQ0mJH
7R390hfepy8GHVWjQOSGucnMFInHIkj/zgTO243nDAkCW1WJ0p5MBa/apEYGbfRoS57fno1Eb9ut
JRJMb510A3CJYph1qv+yyNO0d59H9W0w6flXvXM6i5aCP01IPPzTlpdqFFQENLzCjfs0EK+wDSyK
Slp/seCskzOosLqGqu4agEmca84ZUljmPeP682G6/4N4jvIoBiTiW8uuFH3tvTVBcfj5jH+WHRot
FdHSuiDTmmpyExol9mxUuPo7K704x849feucr8rz+FAjTy7hN7ZsLT5UPuoZq4cGg8v4bymAt4ZT
D5tROvD+kQENh216IqYDvDD7G4uxMzUfK8plYG52rZt18oGfw8xiF4RJwbLS5a19JkD7kWo6KRuV
wE6qo6Ev1uYCbGBDbjF+Kz8h+RjYC1rCFsA/EeYRcYyO/rzMI0ZSrfeb7p1dPhGSp/+umiR+RZj6
YEZjUH4wX4A6xr5LcmR+skncAn00rnH4yJjZllaDQ6leeH0/ZB/IzxoNecUfxp9BoYCoUnB913xn
l2GL8Ciu/HUTQOkBdx0lJ668dHMGobgV6etqx2+WXmr4IZLjLlqgVG1dAM9z6LCsCv/L0kdDHOMF
P7s05pwLrI4vxuv1nFiT97vdNO4Rt2taKxjd+m46LPwUvJJUv1i6GMFM+ui1tTxMGmvAathwUl8w
WQqEf1qHN7RcGxc+0hzgSzUvOb2h5XwtPcObNOfpEAFYn9U3PNS3tuqHo5mBSHYcvOpZ/kGDZFp8
EKzWdTyDtaZuwAmpk/kOU9cf7Jt83DUtmvHe9eL7lLt8GM0V/WkEATUkkwes1DDNVef29oeuNSTM
bFOoW+WlZrVw++0GFi5EFYb40eI7ZmjvbsgaY9Mg2lMOClHoVo6BhbXtGM4oIz3Q9zUiovoRDA0b
oxP8K4MmpF1oAMY0oIdJDAjFMWMyzKp7gwrA7ajNR/yCorycgD9rVDf8dvn3uIQu9iV/l/nRdz1a
9qNO8yIxLfiA+BJwVARKehDpzoPR7KXKzLVUDegCHt+52OBUhenBXMWYceqep9MEKxKCFeC5uvD9
zxakxv1+fPz4f/BVjJorCoHdlZPvtyswexC6hJ/2dQzRCaxyDhHumP3KoQkzalLd5id5SmHLWVMs
u4QWe02O8FgsAYg5SUslUP+8uZ6yo3ICcB8e6P4Vz6Z2hULm1slOyPzYNntbVfTMnlNJbPVr6zJA
Bng99R5kVjCub0II67dGKVWbHS0brUWmdjeN5+vtGxBRRrDRvogueLXQ16Qoo1GHxkWu5rb8AIQk
G69D/yzYJpjE7uu7MDG4P/rzd5umEmjHA7lbJRFOMBViwOeiBkK2eyL/jCHMX+TCF8qisMillvZL
X14nYhfQSSjgoMzFWg6So208AseUM5Q9EXWg/SUtSyvpEZMcDNfWIPMGS7QUY5LxtNBMo9HRKuet
7KPK7WIenH5qMvD1UjAgF1MpTISvvH4DB9NmAfBk6msZKAdATRqUQn245sn7/O6bQNJg/Yi/Uoo7
oK/t3KzfWuGYKUPMcyjxLe1qlOXO+Toi8ZTR0pjacsgAuC9M2NwTo3Yw+TZtBjyhbmUwbwgoCWVg
aON5paLI6zTMCgbVkV0RPxviPAfwmKh4wOArJwK61TK4suIBlUz+Dj++MvdEzFYmSQkxR7u5Ak6E
7FfhA1vunD6lTkgkF7JoMeQxmCyIywZs8ji5FgM4hZmIQXtkgxHEwtVVBnfE9wQv3gpgsuK0mMp7
BZTYVWese9vqTyi1RjmABu9Yrtr58mgun/Q9QuD+8n9a6aI1DPNvmIv6pOgvvr6ErxfW0bUoZD30
mH0lV8fRH5UxRJRmGiAhgXIuJLaVubkJS6afn2bHX60ubCidIpYPcFYdsn31ojwtks5AAHQzLnrU
eSlW7kR8cvTs08bBw1nH6Ieydyo35VYLdJ0Qi8qZdIzpxVc8jvIC8FcPVhbZt2Qls31nCduhbY/c
ztpAiaEJ3q7UhMWb40Tps47zKZ8rVuiZd++5LqSij4eOdmiCjNHoYEkb5euImvITDY0obplr8z2g
ZF8Gb6hIg/eFrS5TUj6A0+P2mvbIA9HnNBCL7WMBaWuZ9pfPhwS8fwtI3H9+Ywd1acXOTpNCidcn
nGf2wL7gxnDX81PgT7STuNRRXuu6l/wbbBO1tOA/YaOObL9VY/YRIY2qJqphwgBtu4paXhb1e5tc
hOqnjoN4beoW8iQlp86v25u6qBaVfTdSLTUaA1nYbOCzIdKmAMDX0pVI2RMLYbSoMkECh790raI8
H2/aykSmCtHZx234S/ZHfDxIehe8vfxNjE0+eQBGuQZJ+xMeGjHrH6Ce0l3U2RMebwncul+2SlQX
P6f9YdyA/aI7++yiOeuxLSkJlh1T+OQ1eK1tgfqwWP7dbigIPg1Hkzf57+ZOnmpGUM3GW0LKtmuV
hZuSnTrbWq3Y9GUuyNi8aq812vYCdK+s5IDDBhYN7Cp4LQxRu+R8WhDYD4Yn98SaN13nZbmA6asa
0XW6Id1P0AHDdYDX1XFGwss+fKNRKfnCjzM47IxbUU9vVAJsLEAo9UTvZBYLthpce2azRysbcUB/
TWVTqkRV92FJlGEHrzQuUBoKgP9IgTfiqBP8bBikgcXyuyXoHvx5I5pk4VGkbu1YgWnVD1SQfUmD
6klZ7qXJSfplis9TZGm8XhHZFW93ZhljPeF8ptIAmn5EfS9dxLw0QCmQBBewLAFcmibp6zobjYQo
LHcZqeMUJE4bl6+t2/U9n6VVLuGgBMYByLpTTsYxv/euSiECMh92wtg9ofqLlClSRQd0GuReblPJ
hGQGSJ/Aebur1SmyA9bOmSZY72SbEEh8VPP0pGbYgqtk8TBcdevUs2I0fVkwisnrlfVb6xBf3CJT
+K42I0XjnEOVoB9yYeSGrE7lNhh20aCvUkzq5cXN5TbRD265WYno9jwAgcju/Fmky/8AEHZXLhLa
k7q51QsmHqTXdy1r6yZQnKGfy8J4Mufq80Pbj2tlh+JpaK5tEVTxmV6/kAREeHApdxdpHEsnTYW/
PkjEIUtdqOX4HNGYL8C51oeQQXJKfo3PYTzplacyughqHgSNswS+OOJGmN0mS2l6yiP+my6ESklR
vl0vCULLqVuu+idcRqJkS4aK2bX1jX9EIydzhWK6ON0c57tjRGsTclK/ADhRJ0+Xg9OikkNbSXUO
8aoWcf7U4LmemVZBbd+QHRYRvi7oJ/jP4QRIUYSiSF5L106gXHmeR6OKgXHBpHdlJDY+oB/JI3qT
rL2ZlyhtVbDoW+m8g+C1DuxghJ1iRNhkrFdt72ItZoNRqD7fo4PiZnNcN1pgmdF8o0koiHQ9AfMT
9o7IyUik4GDDIyKBxpbseWmQ4FOLgsu+BKDO6/03he3r4WgSnwuRlID3JBeghWDfectfI9VqKKde
YpynH9UfaiVgzNeVQhYIYUALkbgrdbTM44l16JsUmG6eiBCGHAlprK3I5+DC384cwRDurYKDdY3Y
iCEbf0ZqWBQ33rEVxLnPXe3dAjegD98QDwab0g/1X1EL4aVN1JG0SGvil/hp+XkFUWKU0XhHaazN
2doe2CECjrVO79TGjpaWXQja8rsVcHsa5MHUb9fm8u1dGtEbrB2xuZBMTz5bewfXRQKorwT6g/5z
vH8n7694sbYb7nVFlQ4Ag3aDdrDoOQ53yKs8vAmuOcMWq/a6Ux8Wj9s3Yj29juldeyclWDfj+BBV
KixTpkyo0Y4BO/95sLNYJyTGJDfZ4Srjf85NIxPyZsCtzdkynyxUUS9WNSWkk6Vjw6plrHtGOxQo
gGV9LzkGqdeOtFwMriazGy3mcZ2umaRy5p0B9JWSpKyECoQxUiqvupym5CB9wMsmTiYh4Zxz/X9e
T6Z4kPB34/GZZgGhI3mR6Nu9CcriAsDGcMz7WgoQCY/J+/A/w4YpuCq09KE/MmpaEZVHXNy0S4S/
Ga5whDceJLhZZ3kf1i35azXwmFrqSzo8aeo2zQ0wpeEGtnn2g8rmtejCRI0144zruLxOcyyfXPjv
jDwzhKZNcMwdfJYkX8yn8RBPRaVJKrK/XiV9SFbIvB72OEEij7WZV812i3Tkfm3gH26Dl5xEr2IZ
05dpc3NWTNSe9QHpEygIZr9IyBTu11E63NOYlFb5IaHRzjZm9mxZneLyiMU91n4zcmTLOJ4oIgY4
G4AfxnpvoAnqXU501fOfV9ISJD3U28TVUP6IGddvej3Au8wDIgLfJnmtjrQxmYswrjYKz7sosGo+
JZ0rrWMCgqfA+KJo0XNMv0zBysC5uIj9bKH3BSSgqza7RPRny+GJDofKGTO9/DSKy8ZI79Y/ofw2
VO9nrLisdk92M0nF2BVu+VhAqkRSUxc7biyDXfK7oXx7omWNwKuAWp1b+bLab+PsgtR1dbCGF/UQ
dXwE2CZM8zsU94aFc2eyCCNgczcQjppc89CPpRrH1AmI74QfKOGqDd5JVjyCUbiaV5LO2oyL/03G
O5GeNYVOLyxoO6LaVLzLVGSuU0LVOLthBSwuj6eKM27k5Tsw8yNd0elWyW8oGnhGS3/zbUs8c3Gj
iCpLYYNMDwJ/KDVYWKJOFv5cK2HcYjO11Iw18aWbuHOpAYnLL6gopg5XpDizWfdx8iOqN/Qx91ug
/+idZh38Ztla34inmcmLTgVGGwq/21BWn4MBMLWeH+XOFdXBrPL+KDk7rb8xfELiwZQO0VRRGmFm
uhUja7jRzhKoBTnWn6HHlWEZ/aAzNMlRTJByfeDb/4C07B/GBDRwTRIrKV86Lplc47iqVd3wt4dz
5XtE1eBxiAzYlcF8hnMdGoxUKuOSSfd8dJgHCFnIK2lEpR9yZWa4NLZGGP4Af6vYkTpTT8x4KhdP
WzvMGBGUlW1YMr1Qz0dozQXHqC0Kksq0fMG4+LXpMxBOFrIAEjZ6x+zCQ3bMIjz7TkgL15G2Lzok
Mg9vtGj7ehQt9sFcO73fBEOjECVIqvT6lq/6BOHisZRzY7XM3dZLQ7VBDb5prpuDNnMMWDl2RzDs
1hJduKayhBhBT0vPa93G84qdTpbCUm5UlugbQjFK/4fM4mQTALVlLk4ku3B30DcYHy7Zaht/bcBU
qtDb5AbKbtPkbJFUOURCNVyC6EwNkDrmu2zxen/Wy50ZjLC5Wfg1RFx1f0CkHK+epM762F9f47cm
nq+gmXt9PiWWtDMQXQSoHpi2aSHfYIJ8GNdmi+x8L5jNuJCgWgYTFeAF320Gok9HGh4RBOzvnq9U
H9b/yTc2YzeYYwKcC92Tjl9vfiSp6kwKnoK0yzdYzi4zwLAI1+JmlnCamNEjrUEYBk26ptV0O7PD
lj9geOOOeA5uXU8ljK8aBAWQ78DSvCQLVifKh9dqBERU1pWGOiAOPU3FJQAf7dQgPBmVg5QpfOZ0
x7Wjw2wKgjFejm0N1qymoa4HpJWFXswka9IBuTJPEM5LQQU7W2z9Z1auP7t2QOhqtDkdLd7Z8+uw
S8cJnhbaf+qhSoztJcmJ2EgR5vZ0BOhsHLTtk4ABg8LQ3MifrIfDRVrMaf/VCIQ8D7+IX230TMia
AvjCwBzjqAK/a1GKPoyX0/m+NHEBy/N0Grs+5D7GVbY+U4T8hRswoe2woh6A8eFwJ25gDnK79ccz
HYgHs6jmPi4mbAymyYoFNKbTMNbD4NE8fisdRrkC7+hEWLw7Q/yhV425a0dcc/vgO7a3aK7omGtg
cABZKIME+I3XnX2tk8ukUFEmF9djBVu0cXVJG7MUagTw+F54NSmDPAyBj60DcW6ajmn+BI6ZH1bz
cY271ClsygGws0XT0hrp7McN8IbrMvtCoZxPTDXD2zFDFYW20KysUtsEPHAYtgRM7EwGLDkGsdgc
JlkWJql/WgFdQAB7UVsEBPffC7ek9Ov3n/jq8PW91oDJlmA8sdqm0Yp5LDgDKUJd4HxzPJrgdFux
NjEwCn2Z7lYhlL+cdpqGiOHng6tpxQntiX48W1ZCfuUH1URNNgYh6jLGTCGMA9rkjNEWcmTvMIhi
R3ePK21GDpQhvQk4qOiOJpwyznL4l6XcLxpxHO2BT+RmbWJkWc8V8m0p6Ka9sRAqsYuEhYnZa/hM
8btwy/kUAEHLxsXDUscJ9CV9m0PoD9PMgD6VYlv6jdqHOqZaNQT3/uHasFwSRkg6rveroNswz7a5
OiX3NMCbgCsSbbQR8ZrCSSegOjPy8InNpMGkHjmQMN1XYW1dWfK8598g7KD/D9MRHT0BHzBAZlvw
0LuEsORRzFxdtUlaKn6SvjIGVgt/4zLtXCZN/OUiWvz7RjvqtGINjqsJxQqsF2tl6vCB8xVmC4qQ
HOip5koJvAU3MSMMKGEwyO30aXyC5OW5Ox6qmi6Zg9NGXT5nCeN2LGs0njGJ2R2/wchtb2znW93w
RW7wVEigz+rx0GojGfDqu2U5CKIH6lvpruIhY+Eyjl7GP0sKz/AaiC/gMuuRv1ESaDM4WvByHSzs
Lg+EKyCF0moWyE6RcTU90SAqJfIN1pgka2LQKz7hzIPd+TvIzRAUQMJ4hYS6eI7c47JIFGIMRLuY
m8qGLwBtYtFDS8Ljd1HKQAPJwdZ53NHpTl8uVU1TQLnHrh2YJQRVmuos+UWR7tpTDm1XeG07fHUD
3oD2OsRy5JGD2tMo7e/WYnvxEPSUqEPks+ZJGy+GZGtqgUgAeEddwX3mgTXKJVvJXCXlAbaMMB2v
8rYpQsQYkwC1W6qNYlgFp6sMu+7lCz7zPvxxHPaMbIEZPuBrAkt5Z2KHmvAV66oUUbZvLdxtsbqj
6gOAVXtO7xWDJ/i41qpf9quyIPlnyaAbanZFo5EUQ84TH2BrJGvZQcMtqRmHvVP920wjYCDWr8bH
xIKaKkrbIueZYKNYVWHFsjeuMG3m8hB8K8fnuE3bOR3MTSys1TB7w8Q5JmgS+CSjzBPXKsTptuL5
H8jR7RpMjtfqN7WskzRrn8He6utWWCS1CvBTPBGem85gS+FxQOa3h6c69UqSnJuxDV9rnG483Sdo
hLK1fMhXuSftmt6Q58+HQQN4B7f+cDPAH0OLY3H4+L9RN8/rUQk8IRtnBGeSX88ZmyS5k1r3jO+a
R0ae3N+x4IDWob5F1+Q0h6/UwKxVd0h2WL5vxQisFQC1FL6LcCCjaEPujYrblNddqT/YQmEFV2Q0
HGH1sv6l3sZ1d8eTZPfOxcKwT5GVlI3Axbj/gpZV5yvCXqTju2QceR3ZQjSeHXF/AcMAPWE6Tn6o
JiniwfSk7oaksgqDtnaJgcdxaNmHfC4MtvttpAwgD5Gs6Rs7dGDJQpid6JzbiCpCaOpb7OjA2NjG
T3DBuvhL1z5vI/AUqPxPy4alenZi6AlKspW40jkA4UAn2B3aB4x/j1Ffq8YUYL8cUdbRdG4q7U14
p4waW880tpsW/FTJHrcQgAgeT6BMdCO1Lwdab+dTFxZUB3RJij+jNs8xdLRKYx79D+6YB0UlPI+W
Hnkq+a5rna0bpVLQPZ+OpZMsIRX3gz8eC4f0+YF2cMdiH40rRt9r/o0XYqpuPlPm6NnauBpz8pVK
IN2iFT5ddImqkT+8xFfAXBVx6w8e5bw9bkEx/rx+eF/YioUrXIeIlFR8DiDDTwTxIt3l5w1OUvLy
scqCy37jMlou0Wfu96kkKgIMqQb/wERK1FURmk3VBbL/wFuiQbb39a1XLzWYUDjOV1eYRcyeEw3i
rA2yNnvnBP16U4O7Tj9dY+H+dow6GDWQkJU/bVlf/mvGmqYcJtLX9Kw3pGTOeuTX/sWf5Bzr7nw6
k2L6AP8+u03c4dvlkZhE3mXycW2GWyGVuVel/jAd8xEzGix8n4DJgwO1JYbApHfrdIscLYO8gNUY
j0LUXuknmUisLXXtT2TMaHKwXOrAt9+fQrlhaAQiaJKxIlIvmTM32zG8kEOR+OZAwDabQfk/Fhb3
Sxo2cEYNiObg+EwOH9/NnUsm7+aG7dZoLROYSOcnwK0OiZw10WEFqr6S+w5rR7oeleCJLhFk/VPH
7cQcoBkRj8MZEV9c/bzuKv2dADJ3O6tkl7Y1uCNGyPafhsc7eDrfxX8EPTuvna1wQmAgXZC8dCfG
GEetCvg6vxtcUrOjsw8b8W24OHkY+3+XKoZFEB9TlXwsFZJUOfgyFbFFkk7XDV9moiHiRRi4FPo6
ZLRTmhkNpIKnPWlaRPVy4QJokP/0gktNm+bfngdfQ5dWdVjv5wOG8zLMMxlo78SsdThktHXTu9nZ
y3DvTprywJcZI+4V2AALIQZLlTdFuQ3g+ozXUG9rCAPC7EVL9F7dCJd0K4Y6ovYYkqzukzIyJ2sU
zGe45bCcsZBdOREiyuiIBuEjROM+0N4bv6pAhMSBgCSiI9VQL0krY0yaG1Eet9oO91IZcgZVWeyd
dYNOiwSXHb+74jOcgbYUn+u41ukVqk4el37C6pVyIa6VdmQudRhaY8stoSB0C5zlkwZrslkOf1LF
bI2tpRrEvQ8FJsbJkNI4UzQQl3WCuWdTtaoNuBswfMb/B7zEApCv55yF3gGr+2VOJNH0/RnbttnE
62bpKUBg7w1ulQPSOb5V4oSb7mFAXUvFVPLgJOWQFpNnyxUCnp8QLICiP38vMuUeQwdi6m5Kd7VL
gkhaEw4Z5DB/3Be+IqkDDD+Z+USdSciD56u5m2Z0I7qXhDJOBwOgfd40OiNh3kfRNnB4AWZ2cWLH
oTctAcoBcBaogn1FDpM11LyFgyFtqV3N5LtFqxIPFUMtz9RyLF4xaAPmHxDWWFQi4DM4F9SuLcud
oD8CxZ8c/cPD9E0MonAIRojAa+z3kQc5mbKtqN8khEPf+CtX4PGfAg2wjfVxMJrUMrOchvJs7+cd
x9Lyywlu62bG6I/e1/JgaCAnnNiDN1fpxDLR+xGm3Pxiv5df1pHV8m2r+YckWWUFS1r6U4p6B7Zx
BBh0TzZG3oNADmqPihcpZKhzMLZbNeyZ13egTbwCwC3rB9wERc9VEdtAL/w1OqyZwTzF/QHaVPy1
IdI8YZmDVYKtSoowOJrWEKp4Dk6T6Fx5dKOjpu+aJq/mH01OP9/lz5O4+qfLDIXEqXMTskdjVfIy
LB6BzV2ypEhUJYghTKNji639fr06mZi4N/NSps71emGgaq+0l9diQxlAly18OMmcB8gLM/qT+I1t
b/2myMuNs6ECD/c4SDzWq4BNYqQ3paBng7tAAS9F5T9+AjS7I7jEyC03r0C3OQbn6n2gvXF1+nem
OMfvRIDCT3CcylOy6LNLcWiOx+1EIQH0LiHcjyoRiGqCUGTrqTyeNpipN7k89qbKPjAQWq8fo03h
e6cpsdpR5X58UxVoi+Kf16vywuOZK+MnzXqpdOsINAHB3uypZrDMc5FIWwyMa5A8R2Oo8DnrDOvQ
7D7P4FgNyMHw2H3loWHIGpn95683ploGoZUFoVypMC7KI7TO3SRrkHSy6dL8R5AZHkEBfM/0Vx2g
+xF6M/5LCliSSjmVmPEebwAf79AWzbjYpJ3vck8b5AGDNAbfFRdy22kd1llQJyLJzyqPUqjnzYKu
SgsBI6CCv+57CMRVzPzhDtQSKtAzNVedf/cqCZRLilhXe6VBdEtSgfjl+vncRs1kS4GPkSLliBmT
LUWo+I0lTg4i4H1PzzbY+74Un0hrnEeJWYpywtzkK9dcIv4oOExk/FUm4Vkg6PVPMqq1OiTTDnEK
HcQfIKQRfdNPu4mcqp4OqeMtikii+kidFjd2sNEnV1UiLFp8HrWmbWWAv+i8otsfP+AEZ3VuJK+W
9kLyOD6/r57IDYf5GDdGytN9J/FuiujqJ5Fv1SVSLZLRo22+6/jozHrbm7mrzkF9Hq5WjYf9bgzv
MYj+GD/TrWLU+zXTbBmcH+tWgdSk5R7ZAXmV1Hvt0EXv5NAVFs2Ozic66z3gJa+srhqKhktML6Ju
oY+8qlye6yCxByD5xS7HFs+9X1zsCkXrjZr8N1pl84Oo6+G3NsfbDDQRdZf6cTzppkZv6j5EF6Q+
b/3RkFgImuRFlEtitUGLJBF3/e7WDSDsNrZA6CM+ej+zTB82lb2y0vDT0lOBjbCP1mDXGp5euE1v
xSk6ZvM0GW2QJCNM+7jHUm6lmXeOmiGyFLF5opmIhmA7fJ9/ZXFVt96++70TIakMJq9crjRhVLsY
AIMafTS/J84XrPlf2qoL2JxhLgrBA/aFhRmW+QDDJNKYN+5+ta1lDUuZkO9m8hIYiQ1XhFYm3ASV
Hyjrh69LN3xbA0lbjSprUVJdak1KvragHFNMMIyICG8tPA5KeEp/BD4BjJtlw20R7tcdUs+vWaGL
z3EtRTcFQboPlSAzfhW1wdzLcyHfwLspLUKEoA3a+Ih8gj41WWG7g3EV4YbaJ+TTtMIu95T8hh1D
AkLXoBqdmswO5OdoI4GMCBAbo18uMWbC5yw9w/ea9L3UFsTxeqa8iLPQne8zt+7GKz6j1nguoLEK
Y9wEzS6XdzpPT7d019hr7Z97Y40rfKXweMEeYIbxKHWDQ4nQuugnol++kdciGgXri1mCC0ZsJMa3
oJBSJQzixm/CyR/nYicG8PDAJeGBG+yDeCD0UgSFts2HPt/Gp0MDr6Ql2LO6+mwWjHqk/62M4fUE
AA+xKamijkySc7A8U6rfUb7Hu94b4mx5bXUowWzAtVA+mq1hVK1Ef9Qkc3xCeYh+w1+Iff3Zt8zQ
hn1jXDJaxCH1BddteK0rEJRKlPZWfQAGo0Zi16ACx7lUbCEJtzVri9y8V9E3OrD6Ng0RJJNH7mog
8TqyYdv0jFWW8aXRRGyC0t3QnFHnJ2ESj4iiZCI9vmnmDX7jDDUX3/ybRjCE/W9NfwHbIfHjLPSc
rYphK1peHWprtC6DRGIx7ly0UhLBJowjTq8DGrovQnCJymUKMejIYDWAkB2DQ/OQRQTJY17JIcaL
/eG3wbjHA5NVwy1JdzVfbsDHHBQWiXVoYQQOvRfumC9sgprrqMPgGbh2SCXJok5q6XT7OQFHSqHT
Mkwu0WLehfSdwawqeTvQiZnk9XrJqG2eU7woFF6NtY7Eq/GqjU5rGs5dds9Aey781rPVx87BnWZd
UOtHqz7zmERfvl/hy2iN87c+CgE8cxCZLIkz45VOVb2AogNDOx6smM4oYhnuaw8gsEN3hpqMEIqc
rk26O0uLiOaCGeZwiW0FLDaBhNx2FhknCuRXEhLWoVCjc1hi78N0VYujDxzzAEqrlZvWB0GmywaD
4dS8jxMuYaQpSEMBg8qIfJpgVnXyUb37o80F85Zc5tRvtQJEaXCJdG2OUGqjWzXm1PBsS3OrKpFt
JjDTazv9J15E19zMr36GZ/Jgli9inpWZvIcy1OagGmAdCsYTOYiQiOdSjQuGfR/5YzSzopjXIvHP
YLnZijGQ6cbkbhYVPa0FITmuprDAtmFz9yPQq3zVlK/ZcXelPuNnQSCeKJNlEBheog5E0uq80s39
sP93KiWRblLIt6aBt7XcZFvMbfrkbRkUWLZfhLEVLN2Fta/UHlw0aKkEhpJlGjKWFAYqX0r11OyV
WC8EVwe5H4DZZKnsh4pnzQbFRm3PAVqlrar/RFtzH7W3OILFLIOyanUQyjZUTyeki6M56iY1BgXg
MI3H9071ineNqXFEfb1F6IhUMfw2xra209rbWTnn6R6uOfdEp8Rs+BiT02BqHg5CaQbO+wuco4Ga
oOfzTG6QduPDgCc/ufOv2ngHRGbnCMRS2dSQJp2mYyyo9Sk5bwHlPba3k9pNve0z0qVZjju7+q+b
HAc2ADBeX55KGCQq9RwrrJD+lqZ9HaQPyZ17NzMQrVtIoNHmGlkJDSeMXmVmS0qmLxvbWzBrMSzq
ueOCBY6ubmTjyan0ypF831DBqjnKQYn935VqwBgRdUL3PqswyOsCCPvo69JpJFuyZIhymXjgGRPZ
uZFifWpVQ9ZikGh4OxJpczbo6+sZEpyibM1SRPNfBZrxBmVG1+t4YjyJgj/S41Uwxxy21FdvAVzQ
1lPD7uPJ7TNT8WCCW3NbsH7ujpkw4DTl+AX/Ft4k7rfHGEFelaXIK0/NlxjhIWuNNQGFoYp6SzLQ
Lb9WjTRDlwvq169PdgDnEQIuYcSFEZ0zg8kSzdBw5bb1c3ebr9lV8Qo+WZNnKk5vh9izynbH5D5l
0na+cMRs/pYMZrPGNmlsP9o2gUH1FIJIKPQ5gbCONaiKVadZdd0C4SqOgWwqxbdMDdZdB6za33st
4NDmrx/bCQ3CVJ909zLTu3uRA58HBUwcm+gsyLaP7fxnEnND0reeSis72yPMl1get2tO3ek4yfIS
YcBsu7byvxgg3b/o2NYOkXXC1M3EEzrno3k/TVOTCzXvfeliFxeE8br8lxGBiYE5NiBbIQ29AgDJ
tSDpQQFKedG7XKaWfDMftyum9C81u/3WpbND9TAjr0Kal18+tXXFhJLiiX7xzVFSdPDn5WsGvB8E
eD2O2xBSIbnRf3UC5xSdqusqFEQiDOCY8tiMxqubl8yqkBPMHxHQveBZEiNpr70cHk18djAp4L4Q
PKw7Oy6BRThXSDLOU+LiQYAFjkt8A0i42vfvThK5lDVyOOS5YGwbvkFTSPb0JH8QjwUJwAJFjaJq
ah5lPujG7hKe9DJZHhzXZF1FRsLGEhOkwUtBDto8hUHAnDd83wsAMyBXrsYSqp3V9p2q2crM/iq4
ELvFcQJhgd/tIrGhem4V5CLUGyys/bKmsstPnsjhAeftIr6Vj0T9tbIZPFMFmapFLmxNIZx50FP5
xYqu10Q4PidgmNankKvbI16k8/vLm1ZVB/tNNZ4weqiEhE4nR5BaZBmyGpBP9J2LlhCWPYRJkrgy
6sAoo8VYxOqe6okHaKdtrLNo7/rKS4plAt+hPgIOXGE4po7URZ55WY7gaMNwak3oRU1j8wAg2+U/
k/T0jgKoEQGxrbGH+w6aVx1kMrIWChbC+ksJVWgoZ3jf534mA4F08Kr3UokrRN8E7DrzHjEBQXCO
h5l8TV8fcZaRZUJ4u+r7VDGMr/3bSA5QT4PtDMO2NCZQjrzjRy19eklZ1PHVEiam5kKrywRbdwyA
H9wcthI1XKGKUs00VGzpF+UUNvdt/154+UBk11Rj1BMx6yTWbA14Y3U16PywSDdGxAi81XAGpo0M
7dZm8MY4fZR7pI7ujmdsLlbaNoCNmXE6fOmDx+Q2wsiwz8KTSrYiHWTJLKk5Odo0jGYVC6GLY2+t
3KgYl53y0mjWwxEwWjv4pSJA5rFQ0ZUmYNpIHMxDFTDtuK1TyF4rIcWR0lSNDdXQ8eSQLqMnE4hP
vCao5m8Sg3aUcRexBc3LnKFTdXNIgri3crdU2CajCF7l6nWx/eXgaaLrljwJSqUGE0oc2SQSRRRh
F8tFSFToSKaKGS9FX+QkpVpffW25pUzyAbj8ri1qEIKTJknUqF7uQah5omTDw2PFWJX/5ycfKSgY
sl+laVQUkJJ0oisBys2BhFzI4LNTlMql9s7V2mdJzWNV+p8t5QO6j+2YB4OTjQTj50HEo40qHMie
ljj5vzSoloktMeeN9obyn/BcrmLJZJ1CHYKxoo1IOSunizEPZrC8zlC7ThonwywRaJAvI7DhTxz9
5zqB86pOLOO/7EmYAECq676q5mYguhPxPYD7kKmc93kn3ZGqfHcQ6oadK/T/JTwvx/kANRxmCGmV
FA0elb5MVdmj3GCEugQWQK2RQUF7y91O7ZWlcQjpwJnlUiFUk0eNG2Z60185YhT8yyi91jxqL+vI
ggQmw2DKXWVfgn3MW72nTCwlcpA/WKDrbCdrhdgsGNu3SAShId35ZH6QPXx1ptGTwgaVz1uOjkS9
UY/b3bRFF1hGxjp2nOAeOWGuqUO9moFEa52GRmg4q2dvso7cMAxRe/eLU1QcZfsaVIk5HSeqOnn/
ciJZsdL4es6AJPTAgG1NK9vMvMiSSRCiBbzd3wornWwZ1kge/bCX2kUGYMm3k+cgBcU6xUf7Cd2+
sNc2xehcMAePgIRUKYMXxJpKFKb8zYoLC4+Vw4oudSyFZda+sdOHHNzxbnHkcWXZ4vB2Xo9wo7Sg
boflZayxESIS5YPWsm4R70cbSnVogP9LgCpMQ6a0s7X3wcBO+QKERJBU8h52SD5u2FAl45K0V2Ij
hVUG8fYYEvRykJ7TFubWm4zdlyz9l4RmJV4DUy++JIUuBtnNwVQh/GjrBVxD9bi0lorMnKgkz1xC
5sNJyWywbqO17p9rzQt64w/6wLdoVhLFJf4bXsvi6Uh+oegUwj9jQgzBrMtj3g0NQ5/OyY3xv6GR
pu1obU7KsjzaIe4YiY5+KyRAid2mc48TqLsee14bnzt+k1cgKEMQPgTjK7j7zVmb0BgwUShUPzdD
G7V6+xKvDfRZg5p1jvHlR3FgaoJahSXYfZY6h0gUJxax85qSWF50sHzfdf1SntKcPlQsfZrlw+tc
r8tZEPgynByKaEEAOsnOiplju5bua09w4uhnmeDn7Y9qE46gpepx8i9MWvicBeYpuhn8w8vC6Ihi
GKUUsV2tb7X8l06R1pMJyT3jN8+8jnT+walX4F/gMp8GZw5EOJeaKboEpJ2kWtneeRSPUiYT67ex
Gw19y6A4dgtIZwUVfoeRiL5WfQY44W/boAS82Fu8zZCPwE0KKOdKcCSPMeTzyOELCuWb2Rc0x8L7
hm6GYQEhj2dhBcyPeaIwDZK4zzq/eDrDV64cVF9VAW+MF+WaTxSEX32BSNp+9dSPOzE2ZYxFEkEX
FxP/dfrng7SjaUN83QMdkU80FUoyBzI2GCnOuBHDUEnR1Fmq+KArq9sDH2PPpUVNqPHPKL3FjBeJ
OefqIKDxcHfSY7ANa5hF06vL5EmSI0m8tS+sHOjjVlh5FRmoY4q9+l22fwc51+/Lh+2OLK3UtVRs
/W8oCwJlroKlvQeGyUYWlqRJT5rAkc9XjXxMWIpp80sE07vbLRvW3RC2MHdWSbFSbyBjoHhZSOfk
2n3+yRIzPcxAOIZqVSyQ4lUySXgCn+JasMyzp+VNniJTukb6shuqxChaxSIu+fYkIx1dEYknesAU
iK0O6WbyKooCiEogHkHxcUm96/iKeJGqomyw0Ym2FIgIquwe2Am8qjf25CzQ1I3XeJUpbgCzhsTb
rPxcGWeiPgEzshq9XB1+aeDT1vsyNV04yrraoY+5YBbiEsAtuCfPAlDTubRFXoerGcIdMSSSSkwd
QwAI+glhvSS50Km6zrva5XuYLUHmhuZpT3ejZo6IEEncSXfSSYaAe0LBURvAbbiJks0UFx38CJeV
neYgs/70gpgJkqReBvj2PutCpbKQPPRyVAbKcHgKQ3vjT0+LaoTqyNL8iSON3s8T836JYRiC44Y+
uJjhkoUdGQrYtVM9w2lpr7VMwqd88Cw8J4I21T01b+zk2qDxQbT2yOSPFp3yGzFNnYZkz1grKYpL
TIadFhcJJz59ASMI9EjvmrIgtwfXfR+ySDE7oh9Y5+ZrAjZ9b3YqHDWJiQAIGfES9CU/iLfHckfy
lv8/sP1uwh/2M4XGAvAW6RnlekYwWOXju8dPneorMzesPPAAshFxyGp1+l6/Uox1RZby7XP48h17
StBoAD7Sfn7hmoMtqoGe1MEavcdJdlB97VU5Gmv8zu1jTTNd2aliZMaaHD0WS7pjUWGiE7KTENtB
s0vr9nk07TdjQfYTwErca9P6mU5e3xnGX60azL2mxe6JMXyefS/p/6kak4rl9Jh1YIl6G1/Mmjmn
ap+7O/xMSzRYE6uluucoUuQ/5xvsIlHZdQM0GfkDxSlcaard4yLh0maKa684mwl6HqMsAnUKZ2t6
X8DhQP8V6OKyexCvvA5jRpLTTpS/XxYOg8fQFp4GkPuaYNGjEJ7mIVnEQJCJBarWhp1jixNt14XD
2pBRhSSdwVY9AIj4Nn4zfTAEPfxlUj9N1OuNR7OcOhBEmyTeDuym8Aiq9UW/Cgiv/+UoIk7DBZDB
QcDLrOVBwLEzi+7yTvet9YjDw1X+idATAJEsbWUp5Xa0L+7yWgIFQgcaUqVPtDQbZAmz01YAaIWD
PbGumYCsBC04qRCVcnfU+tq+goX2R/REi8xlnXp+H7XGIL9lNHHdbh0Eh52/etfufUXHxUO4YMHn
rB7T/iOqk41k1blqht30EXPrOGhrSzMHf4rMbjB1RUeiLVyXvCUdbLYeb+tuFA6Yw/9ZrHTQwQJJ
zvRbIhgRHSkSGRAkMus3Xl37qa6OnmaKHL1oBE1i0C7jVLbIDr0FH0LQFophRufItkYZX0BwT3FO
oI5wB52MZHM+p5wy1qMp4wxE0JU7diLQeH4RC4Ii6IbkhfiEyjJo8Fy8JN+mhni2vuXwEkPgZZBR
jbXPZvUEDxBTRAW+OmX6rvQfW2vD3mMBmuRm27SB3biszkj2n190IjBYrDZmEMhbMmEpnk3aMqhc
6iyRiSWUfQlUOQwI/yvLFIdEdAJbQrIqaKp7yedLEnRpmRPY8jaid357I619K8sC7UtB8iMlzBdL
shewDVsciULL4Ey+wQmhmzig2mFMMoRVw9DkklWHYO6pCyYePsbX8TMgGgFrseRbHqTc0gJjuK10
JtHrhhhsU7Hac50uFe8k9WpQb/3ra8Ahyd7uY3nfTiVP5HPjAFBbI2qtxOpvckiBG+qNyRiy3FHV
dzq5ev4TPdtvfxHehAsthbPf4UMZRKRcqXkYCfiykDYkipXG3i+jX7I9eqL4m1YVBQmRw4Q/svf6
+1jhP+9p+QhH27eOC2eFM7EXq8NYGr35ej/DgBIc8KRAaHZzXP1wkZr6XVqMumRjk0PbN1HNuo8w
+aLwXy5R4OJpuw1bTmJvAw0U69Qc+uUkJs4mdwNBEtxg91N27YvTAd4cO4yHOTmNnKiXNrJ1XMMJ
kSkbrh7Y/kEig+cVyfkobSKOXNd7VaQAvrL8OMcGSVnsJL94hpWrMvYG6w7zxFnhRSV4YDnEdeSF
G4atMtUX+16ZenzK3D+9n6yW1jWGCr1unPv/AHKcVcGpZ9jAyW4qpjfCSC87Jox0zP3yvZ/7eI/6
jxCh9dZ4xtsi2+QnpawgxX2tqk0zluzGKijHKrsx72E81hETQhfquIcRtKrInmJ0VZekYYiV9NJ5
1//T+I/BancmZzhHloyvaX4ErWNMcrO+07WIWQy08WDYxlrc2VLWJlRNYi0iKaOH1m499GGzAPKs
95y/KxMrg/tgs1nZaILPmpUpu9T/trCCMhwf3FDu5/yF9YPsbeKCiGCx1z4zKYy+r8JyE9r9wWq1
on8cwcvuLSfYj1u87vluIY30gdoeiyUE7ITb9dZli0zo4qjqm3kKjiVWuxIwHPfmL6L9Bwo9BTJ4
URp3GwZGGKcRnp4bkr/koirWQT1U/+h3xiHMnIfF9A5f1TcXetv9lfe62DGPdLpCwTWX1MnNgOOe
Iuy9MZtix9r0fDC4u58VyrOHEpk29Ayu5Dp/XSIL6zdPns4xyrI6rLSwW/JDb0By4v/JFT79RaHJ
jRw8GXuCWnO0ptYJlIxnpU15lxXChyNbGtuRI4N0jNOI2w+9+gCqNcDr1PqVvfMlnucu8geLOisu
+Tssl5n2w8r1R2fMRGpLt1I3L5E84VaRh1+ZRK9tuEW1w7xegYtEduVY1LJ+BFFatoIsvWaC09A4
vDsKUsL+Ue97THA+Wmx4c6wBO0ShtgPYsDebklGhDXIa+lYUXtKn4AJY/UGMI+NgnLC2j1rnOcT6
dR/1ChKVG71X0W8CxgfSmLbWcEcMYUjuER0pNEA3XbI+RXc4vho4+k/6qjOlasMDAaCkURKxmi1u
BeLMLTcPuLcOktpHB1TWeZiyZJEA7WAZD5OGX95+MS8dJqixeiDz2va204gpEr9GleqR64ZLzwZW
mjIkI671AMAeSBqjjHFjRdCwDeZ/CTFrF4Ll2s5+pF85fDQcQ4kI78rHFwYltXymVFmAE6SEiOb/
x9czg3VTRYB64mITXkVBq3kPi4Lm5M83iAcP4zUEZ8mux6zCuZIM35vV+U0qBfh8LbONbDyesRNG
Mb7adh86b97iuIvazmWbDlavLS0HTsSIZalzD/98Ea8i35EykueGI5etoLyiCfg8o8VekR7G0sr5
nPkHyyWiHPzEQbdtvIhGHxSaZ93CHlowkmtRUrLKrVY1F8u7KhR3bYqiwSCmZkeOwUDo8fLNCtqm
CadkSraJdx7YZcXwgpi4FKLJQcbiVz6olxoAZlnZFZorH8LSklBl6Y7JH0tuYiGS4busNmV/WEYI
CkXveHlYtoxpIrFfcD8x3kjsGSMg4f+wW0y/jH961kuXTAst+znuDTf8Z85Z4D+gr/u+EBIGjzyA
5t8bby7m56xnJDCoEBYNHj9EZxdk48aglb7S6f0BgH0WKbU7VpzZwUx+g9mAv8x0h+YjTpr2XPIR
wcpW9q4d4kmIcQBFndp8+PTBeD1fY1FNvtgh9SvexhDQbg5cRB4Dy7Sklj+tBszBH9Y8jW1nPido
7SVNzi8GhRIi4n6Yesct2HrnOQgyZoIXH+CV8yzjZNyd7xld6gs0AnCg2mLB9vq7YZIdBou7KJJk
ssZZ/LUo6F8VJGalx2+u6zykL+lzAXU4IDIU5devfx2b4ippz5AUeM1F1R3Ef6poMWoqAly29JiX
TeI1+sOCKhpVZTHgnl9HPmGUXtpZdDVphVNnDTX2bkwLN64Av4gld2Yc7uzO4TtR/70TQgQPKLI2
5YhEPZMdUsxReIqWbJRjUXxb3AxwHDa0WGYgqU+MeE6HmVF6wjTgiZdv+xaxINanHGTeCs3KUXll
ZfkgTf9xZTnDTiMdL4vfiR49KyOIZkPYnGtxsu5jRc6oJx037HvVo21MSdXdy2smw/RqfKa5JIXY
C5WvxLBvLz7LdKESdCfEOXbp50VDXRdd9lV08fK1nrKReAhpxknY3aB1H2Nn9QAtVPd+2oesO98M
d5x81GiMPjsFiusnEHz6O+8JIpUle4hG0r5sTcyGfIqm95z/fgNhkVcaPdavvmQgHarz/Ay4NFj1
/eXRtAbmYVVc+5s77FmDfbJTCvUXV/pKEWI0ABnLLOfvWOZXvAzeVLpsW+bPP2Pk+ie9H3YLdO7P
P10Bm+qIoAs9M+5JlyJ7S8VAKHSe8RJxHbnrJjuWTrIdprPeN5zPKZL1+Jgmu6M9VIZqd77MU3+4
63jyDfvSYKuMvc8/SJIAfxPs8o8Pa1PmSXRZv76I/zst/ha4ALykXGiaxs/+ONW0hm8gg1IhIAOs
d+SyvfdaLlx5XRBcNaYMYDN736VSVitZov1RDM69YuNtKTogZcJvnA/KwhTL6N0uDo0eQdJvzrFz
YRTEEWYAv8Rr0qxNk9ut5r4r5XHxY4ggS+kJXlob+3TlRWT0/aLvhoHvDszt743TfTqOiECiuo6C
OTyHp5hZwj3RfpxHc0BtEzl1rWEGJw5ZPAybw0eem/aW4n6CAy/Fg4kQN3/Walr5MnIuYer/ytga
QUSSqFa/GdeFvjiQvbg1tVMwk4d6vU+zzmOY8CJ6GexrK/Z8YgapUUCrJ/8Sl7y4KIsagtqqHg6k
iPgVwIIN361WQAnYkwXeOxAmJDNCSkXr+YAK0emYuzc8MrnvrzvQOkXlhwHx+A4Jyl1FLOZl89/B
mUGS/C2iBafSY52CBL2HDznU0d3360sjQs43wa+lDin3dkn9o1erDxsOX94MQzKgRFCas2/pvV6L
la+UG8BI6AIkwfIU1WvJU2uYe0y0tnKF9itedGlNbqfNJveqAdHVkcUmnJI84F8qm9yVAnWTbBxA
kxLzE9kDz/cSBlvbigKEnRp72iaUCgLhA0HnmKGHb8MpMrxT6cwFzX6oB+kWHdee2M9U7OkC3PpK
Zos3KtecaoH44VxLuSukRsxSesw9/T+ONJe7XkO8SNb/qGlwiPgYZxvuwBDq+Wclq2a0aASv+tJI
Dxw+l3p25s2foUwpUdn7ZjPKXBScxL5wNjmM78VFBq6HLumvf9HtZZEv9L3MKzlUnhAZvxKLm0Gk
/ESOEplsT4WrqpI5EY2HZTPaD/kh1hZiLr0/H6E66gGQaUep4GNDFMyKveucmonyX+3b5ldKnYjT
rqnd2bma3udZU5b8iLn9S42IxFS6EvTzESWnD8EG65hsuULAtz78gLrRgdSu7CjjctHbag3sm0hE
xWNPXmMDl2AhEzBnWviSd/Fen8onEKntW3mgXKNslsdRFkANGuRZcGWg0gXfB8/X7aeDcYYwD02c
OMTwxEQOPT4FTrA9vlZkfx1EXLMQ/JauaRnhAhN90mLZ7RrVT50wczHY4Ti5sKJ3pxubNDXuR4qJ
H9rlp51FoXgQgIvk3vUE1soojsLMPJZWh4klCu/qBWbEVwBKtzood3MGlx/wKaGO8/8BCyy3GruQ
GhKWNjNCUGebHQew5jI+OAuWHWVPdjz+dcgsSWSU3eTjZY0OFCXkVFVDObk1b2WJEZFbymeRTyEq
f8ZefK+yDyEDvjuOhVlnyhA4luTd5EV7mMKKiMGKKIViXfjYarY6EWCtWW7AoPBN0Z23dOrbLCZB
zLaSsItkidnlQiDCIFIEe5uVbJrw9MkB87KYWhwPfBhTp6rO9ePX3q1tMP0Kt9lmP9EG3+Zi6t2P
X7KU6v4l+AcvarBv3tif3/Bh3KgHdhxWYCxpNfaTwlUkmUSFn0Bkq3POgph+kMbMwrSfArjmFCKU
Ad4pNCpMqart87mxk44OfRks5RNrEyD99N926EiXnmTov95tu/2LhiYhXAim9MT3tENhTXLK8ZTY
o/yLAL/2JI7ZUPaK9Z29d8a4hM0l7kj5sg8dBFRlLw2jwublx9FYckACAgjWnf134RiJ9Zn9zHnL
YJwXj0kv6KF1+5JWrzWFaJyS48slcXF0fCqLzq5wbvzPk95VaRFvhAu7yk4XJB32MVS4w/2ZbGOO
XM2CM8uY7PoYDAAwElk8Q55SGWV2sMyV0EO0rRo/zxLuhUbVl6BOMpyL68Q6IXP0W2mBqQryqkV/
I3FL0Eul8Aa7CHGjFfVIZEzWMountaQ6eIrtIjEcTaxwsyP9kvUtLL94mwGBqwe2012d4OveLabS
78pcjzlc6kajg3C+1NyPPIoZgfO9uhHCKy/B21zP+Wxs7vZrmHBZVBd1gMx6/7RWSPHmI2wExdcs
H9Y9kxXQF+ECFfzsvks7nj82xRJ2eHeoTo7PV0fFvpqJyl+y8ukKmkiVddosUfTSb9NQT++lQv/g
yRw5vIY2pkEPDIrwmRkva4oY8s+MlIpCFiYMamtI2YhkIn6N/IBDRnsmXlfP51gmvaFO6WIR3QT5
p/2o8vkPOQgSo5Vj/n5ObuEKMz6KG5TJGSyvauRak22bNQrJAmqoRw4RwpEc2/ShcTGKJwPzexCw
SdVFK4SW7BTQ56MwQo6dhCRth92i7FeHXMzCSwIZ1igWdZ1eHox9NpfejSuzBO+HXm+BbxWCMHQE
6apUed+WnjqWNYCg78LxBTeOT+jS7K4OkO9OAD5N1RprEAm1Z5RrEhyjfOzeR/6/YFrP6mJSW/N+
d0jK44Sz8FME1vOmP6biCuKeNRMF/LaTgzMst893HZzE+Szd7+m9ia/0+wOlkw2uNhqCZmJv1YgH
kU/mQ/A3xwb6meyyr9/rZSYtonbVGX+/jPvAzo15WjxaqKB2KMzg9aqJ5gk+3jCu0g0hIMAjYMeC
XCly5XWNVN8FNLTVQoRAunihTRA4Tun7ejM6uDXvDDta/7M4OeeVPOrOQ5L+vsbiGTAXiztdACQz
0kg08Lt8u177nsJgGj1VQBk2nRhmNIrSJPz0oAyQjAeC6YX19fCM44BIyDRDjU9UUUYjHp7BwVQr
3alsuvaRz6m3+uGoryJr3m5tRYPzwZTVpehDT2QAs9ekvuVSpuGMDNWsx+VcDb6Pe2fOECTy1Hgr
9G8XiNnfaGnsg5h5t1nhfpeKjJncVgDXl9LSIk1QpDT2goYc0CSzZ0wGOEEmlMnp6BFIbIuzeY6X
RmNBRjKQq8xpVjov9Ms93HB0iWZUMYWd7yYdJ16X+eLgADKNb5+lZGv2LXy6kYRwdw6V9i01svOt
G5ZeFyMktfngiBvdknF1nddCXa5f42nHByzkS0tb7P+5hwoNAt93GYAvSRfjRuWzzIP2jwUnlBvr
hVYWwdlJRSV3gNijJbcCcPXJjQ38mF0o7DLDFwZSjZ9a2ZF1xhC0XH8x1FbDd0awxy2BDmR2ISRI
rBEsSKKcSQcbGJmDPjZtm+hI4m5yj613S4VBfj/3wmpnHJkRDIUdY0xbvbSlDb0s1Mcbq9fGcFGo
EbncV5BSAZHw4iXA8bcCMgIrW5C56RioaVOZEV1uBYQbkfVXOXQUrxzrOoucnpbL8qk6/Ot4jEOx
Oew//EsTqOX/obrCaKqQCB1TXHKgPef5DtTp172I7KsCvVG0v5JzafaHBdtdeGdwDs39pWQGwVwM
Dp4kbFYKFQslyBXgUhF7gb23Jw5lj9yioAfPD+FsHDPL8WOhcbnwIlYEzGPT+SR8s+NhcgoGJBCt
ha2IHJTqlil9cOvBhRy8gtqSi9T2wLEKYt13e+c/kNBFN5kYBn8b77ek+ld8sSg3YZI1MRFKeR2Q
VFkqyW1XbI7UUiPhr+/qgqaAkIS6bTrob2u2ZlDslLOB1fgKw5hx2gDuXyFuSoW8dZ5WA8h5ajX4
GEwezJ9IDzagXCJbfkV0li3JjV+1BxJGBKHtQNe2EtUylVeQnGydjao223rsJk0L/NX9TKHXeBMF
nkAnzpWINLQmySgAqoVG0MKzKDIb3RTWdKwdX9L5/uPuX6H83x8d28CJpLZZMfdp53NZkxHADm/I
SSCy9KREdyW3zfYFflX53pb56PcmnCGa6xLPWSGXtdVi+S6QEZKo2nBSpVeQc0UFOkV6lmkoHgCL
4zbaniUTfjSjJKWgBTWGuD3NrqyjgfQ/pstGICFD3Iz5dIRTlzCPgNxTuDeT4xSsDLAZrZx86QQs
l2eJ57hr/v3Otrr47P+WnOx+vis8xmVgLSBJUyGl8x99QGKFd/mVtmco88WFzEiiCD/7pTY6asLf
WiA2So2NGnP8zsDl90a3VSZMQ8RW48jhRsPidZ8Kocfu1WmuhJfrBNDmLKo046JklU54dfdrlTaH
3ENGcTWI6hnvvaPjEnDTVg/z+SqDGc2lPfRaJ+xJj5YN/s3izPQ3iRQA9V7noYDtmJcpfrF1V0j1
sbxfi7K3jn/Pn0POmBBstVRgDWqoAlbPaZ1f031gLQD81YkQz2oUve18ukfiaSzOkn9haiUKcszf
YP/iQ7CfG0ojrif4rcmc1rjJpqfaPDf4+IwbLOmqxglHr5XfkYI8NM3XL31PKgqjHz1nk2CTl10D
iL7hK0+TWKssYvTJC2p4FFMfzyL3NeNlJAzrkx0zlqPfEMLJmhGGk9yGOqMsJnNAtY4J3AjdXH3T
yozWZE7dGPYPte/mIhh2MbEQxDhKx7G/FJ41kmUFlZuNOdlEqCvV9oetZe1OU8DNVjiaLkm70Tt1
W9ajeYb9opNcH4CEw4i+hrqpVFSYDHd5HPGceZ40m1rXD/YVbre1GW8D+t+ZOnV+btjDv9LHUpjR
KR9EevlnLdCOK5trK4/sjTeLWQzErU/2BInfTa15rBhhWfPQ94vuhXpGiIv841LWRaqDbizzURro
Idg5EpzxqZCaSUNRbLWBxcRP8cKorwTpuu6nTnD2oLhs5trOzcn0oh7y+bXcY7R6edYtEUwv82Sv
mNr+25Q3B+bWMAVCLGzrn5f1UZHrOqsujXZ0lKwq65Je2LG2oH1MCe7f3t8Cd5xuwVeLV7OtC5Lp
uxA45ZO2ZAo9Riy5gi01anblzRMqRhPpIAwPhgEvgBQZkT4PeZb3Zc1TeLSrMupWQ3HOagpJHN/C
PsyMZ4GZTT2JOSZIxJmV+EMLwS7XuU/hz5vGUduRyZ6munMlH986+ruUya77hQfJgvGlkFNdj6W6
r3cyvcK3C1/4ebc9JU1MlLWTr7Bjsqpsa1MEgiob6mTgO1Zpi5jqMPD2nR3X57YA0JPVMdP4aWYY
giSxq+I7Zia2TaWbLeMOpWsqVPUDMx9erJymGvrvPBY8fkqSvEENcj3Jhq9+J3vdkNIifyza//aY
t/gB87xQpnOKl2SRvVDteTfwj4sX4k9EsYkxlDfVecgcmpy7PTJ10v/Odj2vfG4FyCPr749wXNvQ
5UiXeBYQPbCBNOWwNcqVnOJEgpp063GM1K371RMPLwWnn9+TFoFDuJWO/nKbK6jthn6S1N37UYh1
ngjygjrIBol2wEM/J/7e5z+7xfgvyZs854Y1tcF1xzXiLJnJ31bu2U+9khj0+BwGdU5Fquv8THY9
mgE5H9L4CBAs9r2zNZbly3T363WVyezs7gy9ha4JoQw6ovQ6RdItvgLSWjYXwzM8YKiEWS1cupI7
zD+HHtBLvaZCUwJY393l+RsQft7m2vdXIfk32/WLOf4wYvj0x03z3Rnz94AD3/60kKa9Ym2Hs0Tt
/uGLznoYo7eq6pb7hqbQDBt6DEvUxLzW5sul5FV/nS/Um7qxt9XtHV0CS0n+LPBJ3QeLOy147Nno
peVnNdcqWCuRCMOGRRcAqqWOCeIUqaCdeiqgIzBfVfvgfdaaYYBjcrdvxolR7y9m0RvxxybxWtII
QPIq9rHxHiye9ldMupwt0Xvg+Yu4LjXQ6SSwh1a0xteZwo0nJSYiAtmMSMMcA+6zMIgfCe7U4/k/
Py+JqqXG0E2SGPm5FKP6Ui6xKUdUo00nPE8WQaJX7DqsV9YD83JuKtSRCQye1xxQtW9CQwaLQD93
dOzQjbEQ2+C8V/LvASJ9UUh1zHAIgxSvRdUoGpzpzT0GcnlWH6mX6vxzDnaheaYlo7KBiaNsNtpw
/bNcfHQM6X9xmhLivJerCJ9A2ThvixV5+kK9UqhL5FPBfBh7CrDjwd2l7gHxpolQ68iSBXYSTr9N
3wLyptlCQf3FQjirvqk8hXPclP4sgb60XUDlBzDoSsEE0ODZ/IAU9DvhIv1xf1abJHKnOFGYZ2P/
s4KQw9oAgo05zY4tO82A+bgY0+EA2I4t5kDHTpvGUDlJ9b9gwQcYdewqrJuIBBqo4nlf/WyqfWkP
Zg3FxDrKANocr49jaUMz1caWc5F16jbq4i7FCQERoQZ/MYtVD5AR7vXkELlNAxhhpTRCrk0zxU6d
kO+46darIbL5CREnfRI/r0PeRbgwkHzrnEYaEmoB3coFb2pK/45nwa8kefwz0Kifp40imV+ztLdL
3/iY/NiBAv7hdfVq6ttsMT3e7wtPNx5Vms0lcjqYE5YwkFYbYy3J708N9VuwG2DpZhWOSnKK37px
QL8+GJcgFHwmzopuP7CeA9uj3H+XLixL2g/4XVS77T8069ZdPptV41cSs/7rt+zwYWoRhtj1hrQO
osKc6wyOWklD3V203nIKF7LfDjZutuLibjqlhDYqN9YYCJZ13EoHtaZKazjQIWoMuKWw39cRdsS8
c2rlsPU/RmFhJc89aKkEHTU8IXYzTJK3v7l2UQq4ai/5LRPj3nosFI30F2aodNh8TmK8Kg6vduGY
7xIbIs+WxtRzIgh9sPz03mY3OGBSl/CoJkUd3YnCCbrfj38Sxm87kisKfTj1AEVLyf3a/V3GhAHX
l/kVR7JAOpKigNZF0rXbemSnj167EoXboehbC/admwxtmlYousqeMRrh3cmUHwgGTEnDy+/Rw9Zh
OGJeDv+4ZIThV8UA/MRzNmOwrhHjgmdn/T3EmoQz+LfQ1x+C439D8UGTERc4DEaIxKGB88HQvK78
5JkratFcW7aa53lFDJUDV3UXjmmEN6xNDdrfAE/AVjUXk+wqjNAjq2jHd2hrK+U7iAXRzwmPypU1
49/RMlxl4knuuR2oXuhlfcv9IYkJjRjOf0hT+OZt5Wv6fifvbtNyzKb/141V0wo/f54ohhp/aSxy
vkCjV32fpQPbl8qB8g1FUmTeV/DKc3wDWUtpbRFFhb1Q+IZEYvpb5j5OZQc1UfBMyGX2/QtFI/TH
YQH3e8oNRQ/1efZK+0ps6UJvcHXbzNInbtRMold+5kLfnbkavmnBFKc5ncOSRdGkWZpbCadRxstP
r1g5hM4Zl2qxjW1oSxY4YLa+dJXTLwAdqpEYFILuMsL4ZweEthYF36kqoWWxy/N+F0vCG/3R4s/m
mAKJGzMX82bIZdwC0xzdLhM/Zt5bWryE/49AHtjxyooG9GgTK49/LHfyHuxUaeMOXNdZkRdSrNcw
xslhpWOx2g5jFpz14mbxYg2tBRZAS9n9ncccVQ6Cr/QqLk0TLsuk/s4S7dL3OKfWWaCuC4ndTQz/
cr5ZcgVLD+4VRXAcZktazkDaCBqg07zMe2F1/LIPXZ6LDw4j58xePGgF9V3MtHxPjvSma1CVyPt7
BH8gZPmSPkw0Po2Jzrmd5uAENHdvX2LUk9l3MZ3e8PMxMExHbKku/aYWQWhsH3wxN82hS95zzEeC
pyr209Pa08RJtINmVTRxeMUTBsAsmoprc+4NgLtB6Mf3wzLlGN1Fv4hT2Ro5e5xFD45ILuRVSKoI
0E2K8stV5PAcC4Yt+L8XJOBhh6ih11wE7bQfWrF9UBZc1bD3eB/pTbvs7gRrGzwk06u1fuvSSauj
f45Px+S8xemrjlRi7+gkHxsPp68huqLD+9emabKL49i/cR6KKgS5yPqZf3d8OYaPyHhRFhMC4Z3t
IerdVk+1F04dKT6/KO1VGE0wlDXnFkJUEYV8wu4Vf6gAyICG6eOIbiww0YLyhbFLg1dXC4iuU8dG
8Bj6XSZhCFGh0Q1Ccv2u4hr8dnbNtJMQAltsTn0Hdc32UVYnah1aPBHiCpExCqGm3Jj9/L3pDcug
w33Ep32xxxraBvh6Oxgya3wkhm5nduLnxuqOvoUnJ6BKWZaxbHwE8ARYMGZ7eUuR5n+SPMO0mSlf
MfFtmKrpCNBJIsrzHaa9MmezWm61+8I6mUyuOvb5wrD8DJCE+bZWwRYxmS3OA1NotK8bOapLS+kk
rzw+ccLeTuu0aUmrP6hqWfxW3wnupheQYsy80BHHRzDibJkPPrnZybvvznRqxRcHc4dcwmKT0QUF
2S/s+8Dv4iqB5ubYhNhIxbayoJPf++rukaXYR007UNdcIbl7ULxsTJdNv4n11+Zlg2o6iASLLud8
qKB6nFZtIZGgow0WklsVz7K5mf5AL5aJKKMrARLmyhEAza5kyle8zfChpneeEzlftOoa3ePT0rt1
EORrI7j/uM0Zt+9hmmkNFb2Kfmi7BEngFBBAWmVNLUOj8rte7ERkR81NrJo3TKy3rUosN9bpNTv7
ohyTZAHu+uuh5uuqnNK4OSAijPO9TBgJt7IV1ciTm3Z6M++/azOIH2Qq+rV1ZyhNs7juYO49cqNH
VtGEmDHownj5tt0DQaW898tku1cnFF2LgxSJ6HSwcMclFWXiJrVHqm4gFLpdU4Bl6Kfqpo8A/Kca
xAGmNJxL+V5gQZ+yLC767f6GRhyl0u5J9JfyShYqXt89PwPRXTzvMu/W5MUxfL7rS032p5wQNA6E
W28pLEEnJsguMTn/X2DpN2skTzQC5WUF9a53AuLz54ktIjsCX0esGMFaqBGNA6LNMGk1F9exOU1v
DAkf1B9EGYMlu98MU2kw1Qz+anzmI7Dkz6KMdt6DnVjJ7we1LNsSqMwbyetWz31F6pfz3/hSLJuz
1mQNzUFplbkLCoPgASVszOal1PLuP4meJz7nYmgQUAdDiKPvzozfqTqCj4QqbWQCIYnvbI10Y0Q5
NYuO2ozTxbnZIZkntNGBX0QBIC2pE/vyg3AaZZMtGn8UuOidy+f5aOjJrQnUk+zu+TaK1H6y4LTy
5NQum4Wf73xOig0ogOLQbpPOhaVVPzOcm2yCdVSHm0t6yOLm7m+OUPRrz/B4RQpfwl5xBSs5C0jl
IuoJbO5fJnX0+G4GeYyl0QlIPAWLi49yW/pvAH0hQLEh1NVY5QWyLZ9WU1/qp1kTLMYTECg3nc0Z
Yq07KpI3KuJM9clwRCNph+MmnvFXGX4lHPeLDF4hvXF5jnmyt99NSpN9FzSwS05qaao+qI8o5dOX
qwAfHnAR69WI1Oa7lQ3d6BOXH8YDqGJUXeDbgCoUVwIdnQvR1PXBMGjHh2tUWOWr9beE3lvOJ/+a
/g64aTs/39/JqLzISUEyvciI/hdmEszQdFH+F0WcT5c/FZB14a6W8FSlmMOB7O9tLfBUB9JA5US0
HNw8M3tdZJApqms2AzhnKwwXoYf1rLQhCo7bRmYfczybgpin4ZxuYvOpJBzQICZlodTEEJ0vX4UU
TzI6woSKtMqy3RxMb/9blIHtx2duEv3NBi2Wld7tQwnre4IDhSMUKe1tkKR/AYte3VLmga1jdnRh
yqqrcGVwDGjvnXX22XPaMZfzYG53XghN5lFixA2do8C9KMg2/VsbaPC0lrOOhxRYMNSh3V6aORj1
P+XUltE6KvEZYZroJ7quR+RdtMlwo/9TsHOB+A/i+Upc4rRP6er6NBusVJgdmNRUUzqRphT0JdJ2
E2m0v02DwIUGaYMQjQWXMQXreoI7r4kPAJfNO6nIqh38DSz397A8FKWJs2hPHsxag8jaXhhElZ/U
QIH4GSaQswpyAAk+LmLRzIbPRx2cohhakAeuXQ5nOLsSDSZncecyC72PiWpO3AIzELhCIS4yWR7Q
TfXDspeLGLEybKAHG5ZqDPb+MZIFgpV9N8CdCti/HW/nSt3FHhhpfaKjZaBp8Bx5Naie0fSGULdG
RT9O1pOrcC2rSOu/G+H80FsfKdZWH9V+ys6p5eP7MH/wlFAnj8vDt6Y7nC5GCAiZo56iYr2jeG2z
bQwh0PLFs1c1zy3oE5xOKbQ0SeuRIURzasiJsSJzYBi3varjoy8Ud6gIjrq0zYucM0+2MCUK1YAH
yjnYkJ3um8U4Esq/2M+EbDpuKqXfNN5ivx90qdcJBLF+aNr8vCXd3Z5U3PH6nTRTbVKRvN9WSL3X
qBQwulfXp4FdMRsynPW68jAgaatE69w0fz20Q9HK8H79h+HNSCeggMyl8hkNJYylgX3PUyzjbwyK
41zK9ND6mBh79ui3N2EmgcdIn06QcVHj/3ZqnWry6xlfBhGh+FVjrESHGLpshGE2H7ebMIJAITLG
FRch0MSlHtfacFJtwWS54ppY8WZ+YD5b0wVwV4ywbQILEEDFt3khQmyImdCOc8qxmAanll7uGFNk
KUxQatMSW2F7i+qY7jNrEHkAYCIm6THPqPWRtjBSretdGld4mm/Kr+Ki1Y2E3yYII6jMcd3u5OOE
2Fl9jhTIvb5LPhoF3FhhW9xvy04oQRYuclhZs9mVGjAhCCP4lD1ggSKWQqttJ317MBvTaB3aH5xS
B4+4wbVjVg6Ep9QLYOk90k3q8NFZXhIPlyq32iZ+Rp7mijdfSKpDs2Bt8/BRWG60q37ptrZCpP9F
WOGfKnm+ArsO1mLOcArCUp1DYLVVl53ea7/qz33fXvvPOktkX55AuKS/mkc2Q+Hi9ft88bZG4n1z
RpTI+JZmycDfoFbGkL31rkboD0vlBiz0YIWHAcr75SDEFxugLFRXhi1oVx8ME8v2ZMCkxJJE4A6H
U52x5tIEGZ0VTvvAlciifcUxGTEKJ8BMJWSd5wD8Fu6+tkUq0dHxOUmpnaNZ5aAQV6iDn/Ud37T8
VW3Qp4o8s2hTPO2yEDiyXtUAcNgsIWPjHFrWIJfELh2JqO7rYR9iWwLsWwJYDKHpHQc8vRrG3EHs
34OFsNRMJCGg22cD7uxYSfBbIwGMTXm1EOlQ9Ce21NTlcd4F+C1rk/Hhc9UMzUQ6qO0TMIEnJqC/
7owL3TfhvUExQJqCigGWAnt2zGxDbBtDrEBIacyk4wcpfnGqBIQz5xZoJ5iKYXgH8K7sC+QvEaJO
8TWF0b5G7v3QzVzKG4DRvp0cvaWQj6TqZvBh8E3E3t0n/Kl8jivILA0tNuULeod+KK3oMp3usfn+
ocIKZTxBAsIqSCkU57ydHDgTV0HzdD6GG5mLM7xPzZkuQ2sXk9iSWYd15nYvlvaGoZoEdIAmXNWq
NQi0/HBmUh0lVdZMK4E6XZJL965GeXeWuOQHsI6LbuQhTekwvkGhFwAc6c7RyRTzG01A4HSxW0Ij
mgTYTOElhFdUmR7KuLjvIZCbZ7YxTPyWBoGnr3LZLl4XsXyyCQq9SAg3/PfRckxinXvVeyWd6UjN
PMj+NNw8QMHXcpyF//+5rqUeeFPkJ3cOVxNHoqwyrMog5t2qyEWbRZ/HHN8bGUC+KX/ABBOKNpKu
BTq+R5K7zfjQQUcFUVvcYEZJLQc7k96h3kj2voHDTvD0lV7sy0Z83qww96t4AEdCpCRjNxgpem9Y
qRU/azN7QSLBPneSG7fc6+DcHjrs9988KeecYhLK35x4FYqkxo40DmOybSzP+upJouTsAk+uNd26
BvJwUQ7ET13HJ9/dsvRTHejCRKenms682l1Jwk4XTRI9MmWkyGDqPUtp/ATEoB6LbouQn6ZL4DpQ
0Ks5F+JeSRMJnBxuL3ja7LkNjpwBRWasSlOtw4K5jS/IzPzqfCNlrhfq3iHpmb9pBacP0HNVwg5n
mZ1BBz0UvBCrwIaoj7ljyqr9uXO73GUkpTQ7/uQyrZoNVg/k++zNr7g23/RvQiJdgXhQq8a1Wr/S
t4IBxZ4ccXy/Qw4PrRgKuuyDfkdRdnppsebQl6nYFyXalo7lCcr8zogp/+ZJDpMkAyZ5IQaxS9j8
75pQgnZae7p/rLYrz0o/mN2VrU4zVyfMUkXnAB8F85+mJbA+wUQNvV0kWBIsAghdgwWTuuQR9aT4
8OE24mN4XCPd1QgAp57H5JXLGXkLlTkKSsaxqSf+dsJPl9gcQRedJsKBaig5m2+59DoSu50amWXh
bQUu97gShUgTuMVLU/SlAKa0hHJn0zSEPINHKYj+JInnC1UDZsshqp/RO5rlo/kpsfBaHiFOuOi3
B1tPeQkkLk3e5ITeIOw9lEPG2w2ra3DSIa8xbezwY8T9nR2dgycrWmYap/l4LSJ9JZ0f4nIaz5+7
p/Y1J4juTg8QgTtwsVxU56VwKuXwEPpF8lACqCRnLCywlrD1DsoPjUQkHx3UZgo6EPNdkIJNPg1p
SdZEpKjLvWuBVw4QmEkClUcDMtl5a74hgxwzcHt+MMBZWe4A3bcuAF+x9jHGGqhtrUeTEj/IyCvX
R5CyF79E2VrE6GVcD4xH01DwIRAC41xysHmBX006wCaOuRctDLcap+PDXW6Fwcfg8DgfKk8ljRna
bfik8CiU55hQKsu6shHidLfeTTBsbgJtd+RM37kOdTaNxhn+cQmhdT9+kIPN4xaf/C63O64iQiLO
t6I/NxXZDRS69COFOTgOuhpA9gNRU22cu4tUU8VfweVjKQyueFf06awjm6K0GrcRI9+bRQOyjPBj
rzaA9vxQGIGLujBvtU/VJQGWpW2Jp/QchInrMAtIzIcbjv5WQWSp2oRcoe+WA6ghCXxg5R8ZGCZ3
Zm2sJK2h1lOPr8XoQ+MYWRZUK97v3yMDMiYRqpaxPAz1SejeQGCKEwWKmXHHhhFfmbugrzCk+FkX
JHniZw4iQ4rfcLvsxVLkS2JVMASE5dyrIoudJAKL4dzSOI5RPR0KATp07KV0nvN0syEWXIB3KtUl
JuZixhUKOmubPOr3KdzOPEfUO5DyXxt0C21Yb9ePrxNARzkBwdDXNsZO4TVAT6Wi1odaGz/Bcg+w
4IKILcn/3AF/XFgPzXA8XHvm6dFTnwLkK9qCxYEwSPcy8r5N8yji/SG+u+oZr19W5vy4PK4VkzGj
T8b0zyif4Eg5nOskK5xMMUZvMrEzyFOvhXyICYFrH9G5pUJypO90X67z5acksJ8k2nvfuW7lDRyi
iR7hEgnehk4pdIzwm/7LvRuTj/nXMXo4WCW6buZv4Xfa0/dnrdQ8ry4QCswhe40oM65+GSt3raYM
PflNmX///Qs7u77B7CntkSilcxGZjG9sKRiBvmX2SuOFLAEeTNKs+GSzFmUAXiuds7RJuHNuEMcx
h/FpB0rCo3RrwSNZ14sUiYqCyJesaLM4R5bs+S8LmZ5RHZInlc0PDoY9v44j8wgAdkpQ13bWKtY+
zvDu7LkS6QZnkxxgt1X6DFV7ZuCGcX5jfgPmvZvClyuU1fQejEv4Z851xhB00K4J2tsSDY35FL41
dLzN1IxtdKFsJw+WKtoBUogJxOIkbCpFw97cv0hcprdhXEscT4FLi9X7Uuw5DmrAcdxPKBlgVvji
NC/tcvVpISfG9f1CxI3S+eG9uO+ePLEeBJefHyFjWcYCaq6oEePu/RoeB/3BpYOy5T9e9pEDGAsW
26b8aYMz4uxnxXemmoqr61fsCmlbCQ0RWJ9mKFvCBQ6d74PAAwMswVnwcrJFcCkK3ueEI2s9AZFt
3ZEcuA3xQpl9+1/PI4Wmb/3SL0uWbNEF1xQ34h21zaZFjOLfxf//Rmsu28iD7u/OUWM1qms/PTps
fhIJuhL/k1pLGG461jPknNpaxBHWJc0YXYiR7yz0lwVUbA5Oq7e92UDgn/OT4ZMIpPn/MN4fPVjt
1KgiCzmNxEd1oISpem9Al1VgfZhfQ4g+Z5caKOTa7A9QiNt0aOsUp4gv+MJrn79++BXRLKlynMnQ
Qizn0yiLtF6iUKqOA/AMfJcCe1GRihVzEdrWy5HIMo/VJN1f2dx+kzqo1+cKe0gggIViBWUkxJ/Z
4fgqQKhYLM9QumrCO/cDGCFwhNp8wiHgtF4NR5E7rlKgZd6K0r0Z/TZDcDFCBnYSCLV+2EeOUTNh
7mbjMtmNnOCY+ZlTBZZzOHgVAfuCoakhv0EwqTI+gKQ958E8OoXj9psId9gtSfcq7AiuYHH31ttp
aY0Efb54LTtXX+air+z2M7AzNePqcb0OUHNCATSgysf8fhrLo62UxxLAPOAudDelRc6JBncND2KT
ycRK2mp30VAsbwGtKL6y+C1SdA/v3cFOxG5QX4rOzLm8bSA1o1OenUvOjL47qIlX1uwm2U/jgZ+K
6BQZPfg9d3G3q9s4LsyOvoEvR1MeGyZxQipe856NhKjVCTRTE0HSRbOMJUh2Bo+L9vDQShRlc/KA
rQckb6KyzNLNmkFr7kYn+GMVTAtlQbvIPCB0zmnzqXeC78FRSayw+bFRWd7pFA4L5KASTFupa/sA
2tsZNt5FxUh0+KPVNint8kLtlh2h2Qyfy+uqkCoNmLTbyylUhtTrS6ybJq+wwCBDuYuuedVic2rj
Ys3B7+rQ6AhmLPobPVHWdIWbLonD9crMXZsRy39YKM6DgQ1AhZ2jilorbgsPyaPgeEBWucxuttww
/Hm4cKBiaQ7AhvZhhg9RxguAcsjD46xtJmFwwWsxshNzONXlif+HqwT+rQ9kaOPq0VWCZb0CkUTX
ZR6GpIs3zG3FaBMEh4wCxkTobz6VmHsALQyLsfJ0TGgezK8NnHAhABTZIc+RXhcguAFw6u8V4tMS
S2YtQxtP/sEsnyK6/P+dOgqCKTg59JhbC9iqtWgYvRCY0ZaAkS9jgLScyEyCl8wcgv+WlJhSDqXY
EM/bdWlvIZ0vA9nwbPwSdLIT6uYqAa2p8e5KhyGJpGVQeNfRbcYNpJOTXAjIna/63rhWqf7jGzqP
zGExmoTdxXl7H0q2T4pDBHYUQTI2duaYHkJAZPhVuFrURFPe8vjkx9VwZls2wZY3CTC+ra0t/1Vl
QWkJn1FGvFnfymdR9d1eexCK+TAQ/CbIoeXWz6ojS+EW4KIk3lUquYYM46HnhmKBFiHsTXQ3Mwcu
thOSorTqvgp+hKLVxC81nvtpobAnWu9SDwCYcuNcPQAQJieqPdVK8HgXBg11mcUpis83f1kUfvyy
vCgjNPjxFVVeq5Jq2+mwM2WD3nh39lTdrPlQNo7Lkb0fAdiE7f8hnPo+DpCW7RQ50DJkL4/6ZqnF
H3RyHL195ihIfE2ItY5LyfwrNB79TjBI3Cpc1aMkcIro+HA109yaI0ijlCxQtHqoioORt+MW4gAp
jzMw87ZQU9HMLfhciuRwDsfSZbf7Xw26/Ds/VneStiIUGbP5Dt9dARUtoR+CWsRJT78OU4RXilyF
KNuxfSVkdHWGzrV3k/LvyHBtICYABEn657zT/TSMPo0Rhd1dNpQkYF9P6bQKx4HZZQm/TI2YZgdo
85oE93UbT9IYvGXuvj96rEzcWagYAnenIFQ22/8LIgF82a1ZF0AHsrduGogypVqPXujVl/xdr7gZ
iD3gQ5jq7L1bh/0puf8Sb2vCnOFbb08+eqZn6PQQp3oX+Cc8ZOr6oHMt3vKp24A+a6GMqtsTPk3H
6t6cw2l8a1EaxSgcCwDOFOnTQftlVGjK/p4FYXS2Fs5bBmaEidUSS+fQ3UuGq7PkdZe7Y3cUtdR0
NepnpWFH6iDcTcUQtliTNhpxHo7QESbRVN2+7Q3iCBGws4WZtoNMM9bOJ5ZCYqgE0E5UvxRgicPT
mKPl+peTZkWFp9foCCNRYkV7F8zWRdmVsAtpOvdO9ijWZgNEleV9OJCvIKMtG3DDTrzWs73rLwlu
aHAFtCxOK++PeHsYTv7cA6mcx5X53evN/LtLHNIWGfw9ijnoIYS8I6T/EWgBCcM3+HD+mDCrmHyG
KxNRq0UP0QcxiJ8nwyZsfC5Y/nQLNElJqCoUFLcfh5pVPsukkpUzWUF/DpGNQsCmUbeXDQYpMN+M
hveXilWoAXD/KhGrPMZrtsAcuKHE9cL1FbEUFYUeTRL8kRvcbo5IjpFkEdXfPLaQqwGhpP454+k1
kjG7bGUiTn8fIcg3SP2NtWPNPf2f8L9AFvYyIA2FUHqebxfZBdqBQwi1fs4BHbtzdjsSr/qFUEnx
Bhfzu2YEsbms/tvw2aR+slYRcWBVnkKL6QKUZ+oCe/5NzpJv6q9Mxi/7T4mE6esH+qteP7NR4ePL
WpEaMXEMzaZ15rG8tJjYYlYEqX9nHxr3VMPeHz6Sx+StDx/fJ7B23qdHNEGJpi7C4/T+HQN3C9rF
XNGjeeJ9ff2Gz28YCl/3ftfkwju9KhC84LQa+YcE8t2gqyUhq9ZbCEMGQQdGd2au55Oa6NoA9gUu
ODtthXgmSC1UouuyPeXEbAUUFBNeUNgMVKODYMwKMwD9BiLkx8gcplr4WJ+G5mZ8bY8wKpS/QPai
08sPxKdC7PnSQJHV/OJhm8Rgzm9OcPqzf/gg6GWNsQVMXinsquFJMOvKyPEYZSSQ29YkXF/nqKMd
UnSftfv9VPHFeLozw4UYqQcECNMCHSiATx4DXf/4GyA9vDPlaLBuuRCFJFPjNlvea0g1G0hvHk5H
pYiQQZTLYsFLvuNBZaT0lvOFRqpryabTQ4kD5y0hYfjF9qAt9HvhbCUDTVJnN0t+tiLSZIasFOUi
/VpaNMuoGzOhL/tAi0bgerLlx+Fu39sebH+w+KwOMYP9l2v/1FOFXTWOAs8CZIuDBeYe2W5lJch0
jS1W32Z30Uk1hhFsew87I3W4Vi+6/lCdcYgfv4XWZYJm1hwKQgCJnLkoUzoTZMAXxZzx5spZkdUI
a7BKQIMnkshxM56xzbz2HDuhZpC+0UXDoEHjOMy4ojwoXp/53wxXflepz7LRFqvCh7aQajRviHud
8Rd6sWfSjgkYUPYyHUTwW60FJBiAWDayvFRtIWif5BqsqRQqN8i+yylG4ThPCHFjM0Jlwdwv2qSL
WT3UTdlRietrtagtECKTNk4QOEHHFQm2lwoxDwXcrUHWxsb8TKnJSxIEQyqj7Zlk+zyNKJyjfzIf
3Tizrdo2cRsZowiB6W0jzotBqNutamLlAkTMiJHqK27pUWetZP4VW48Qz/s7qBm22kMbdDpTIoC7
RWeB26pJgrIaHUAqpY0pD1nxKFv7RbSx+VXubWUHsBJ6MMJzn3lWTw9rGo6ty89TROphICgQLyft
VS6R+Pket1SqEq2cq+3nRV36wNapLxTezv+fmAa/WXTFOCx3l9NvlkcVG2Qsx3WwoPcw/qHsWa0V
momZoeE/rESwZjqW19qqbPj8M/z6w1ayVmIKivIytnUuQ+n3K1TQfXYBYwdxpACRORWfky4AczZx
FzjmplKI3l301iUws8m5QONaL7XY6NaOol6BUTm9GCtxotctq3MPg+3a4w4zm/2ODN8lZ9eXexTG
qVKs1uRuCoulkUmSdkEbtiS3kRt2BEC/twUMci7ZFqNWPLMh7Gaz7IdKTBYAtL2UdWcGVgkRCIUH
tBzEx8ir90tzzEW4Iq5MAApgJNWCDA0ew3DDrPpKgVfS0MLWAE+Y8FWdKAgRO0Gt44S3Wi49u8/h
Hep/e8fJl34tLg9qGzUHDuYYnOJhZm8NtwkesXAR3LXG99bvppz3UvuBh8IBrSsm20YD+vuXJJRG
ocf1md0hC/TzArC2TxxdYXYKV5j/KArnz93atGsYpDtOnjnGsJY6jbnP5QylMikr4Burx4+fP9tZ
YLw3sFOvKjWssmVsAh/A77QKojeJ7ZKM1MTyFEBglrtbAl6GeXlneEYjFxxO15J19bDYNjn7O65K
JgAOkSEcWjjtKCCM/BbqNdDvnjonkaCFa7ULOc5lrY9hjUAmVUuxxZaERZaqARGRDrH4oV4EEs+b
vEEiXID7CftKaGIG2oqfIxhLVPlebEvKsnQxVZx4dGJSRNzhEq6aYZA428jJLm6LnM/sMCVq8VHj
o8warT7Q0l74SiVT9JCsuc9g+KlMxFg73xERwZYP/9MzIrlXydjvqvvaoYfC1xCeiW1bVYsKxf0m
w0n1LeXQC+QpzGuVmMFkrHXyJCuqagxEEeuNgq7LPNFJFilz0bAdtBgBHMD55JGBsXDXdHjU08Pq
4mx50UNfVY05/woa/0NTq5eTlcLauIugpeOY6ZHr+vg2CZDxlTnTrbGcGmmdp+IAqNx1WoF4UBTl
0Jx+D5vgMJzhmvyxzvDizXAg0C9Lybv+DA58lpAGoAjdWwMFmXG5ZifJDpc8bhBlPkl96n7SEqqe
K6ow+gObud28zIfJspaUmtZYFAy6Hu6it09JSBy4lycPYN6jn3RvigOvujHDjRrpGqJeKRwa7wkC
1aB5GqIrotqx1PIZvVD4fkz9yqrHWCuNxu7rzM6mte7VAOGv8l2iGfmFnV/DuYO4kV8lgAbvFEFQ
RY0HJ2A8i4HHJ6NOeHLoMu3FV5ibokMlBXEaoMa0oy8OGg3yYXgp78YZZWWobzfi9dFoyFNj0anR
DLh8qnvTcFtWgqIR0uTFIGcVyFBd6JNvxdWJTDG3b5m13OlIvsGJzRsLw44VTZ2NgXU36hY1o0Ug
u8jkLjh5tmapTG+42X7wMJIlv5ytwdWP+Xo75XVTl2Ay9UCKslIEbEklsnMA/nAgzJ68nR+JILwO
bok73KnMj0JnBPPN8w59GjhCvtdX70geLRlrEZUPT/fCGzlF4v/0FGqZRWVQTd1l2pYX7i9B1HQo
pFVEU1iFgvuwyy6xWeYIzgIyRu6JqpOGHEt919Z5C3NGtGmWrWMDpDVWrXad2QVVxjEHVdpl9RRj
oHt2nz6jTjUzYwV9yccWwmyE9LY4brboQdb6pu93DZHlFIYUa1Wp7DWkwhDjSrBJMBQHyDTns+XK
qqykn98EF/rPgTq7L5NfN7WbOKoUhcdc5in9hmoVlmwvdmfp0YWnwMOr5Y5rf2ToKTadFIm739Wv
1xa8O5gW+1bguv82DWNcAszXNWGushxNL/EYCus3bNtDe2XMHY+nRaplW3n4IOHlzjXs5Gqx8a4j
6S1f+HWdgSUspSbdvoa+QzDWdYxbQ1Rj+zPEbNfPLE++EfNP2BJcDSOuhrWCSNRUbhrYQAUR0Cce
Xj41GTlbQL50Jh54i/wDDJLdZi+BF69F9GCiRk3MMOa2fTMWuUzsLue5F8bUahZEscFvZAVxewEN
oS4jiTCyHFWnXuPDAV8cGu9eGIN6AQpoEX7wCGiEULtXaqSpsxuRRblKrmXD3lSYGwFFA+PRhOJy
6FKSorGqFKz9P+LRxPcebyXk4HRPqUQUf4ncX438IgBZTL+zPTBYXkIepGxayemQO5R6Q6nBDoKV
AOlQERuP+qUdw/PJOeTjGiotpqb98Ldtv+J9NynGOBfvTysEFgL74HsjG61TLApwFqYHuJAmnzzo
uHKziJLyyvgx+DWaEkzwy1IlKehN4GO5YP7BFanETEQAjCeiaZLXYskT2QpSfy/toF7i/UEyMsLo
FllgWz+3CJPOM13ww70B+JO3DwewCmr25TDu3K4QylpvGfQA3z/4jF4LSXApZRkNyYTRSEv1Wlm4
0ltnhOcl2Fsu3FmgaAyLSbWJnOI36gc/zqJS54DljZYG9WJMjdKEYyUGuCpbhUWaqynsBwGgGVrG
tMbk08DQvieyoISxv/wWQPUsNiwOq92RTf7r0qc3c00tspVdw+92oyxutIeMCXMwOl+0SRxnbjBT
jrHLiiN1SYdMkB4e61hWV3hFPr1KR5ipNzecz7SOczeAiHRr/0X0S0BgINxohwf1i5SCCUDvXBzp
fCrRtr68aHckAejmWo0TpPqS62UpfTMEAnAipU5VfCacQrcfRHB78RZW1uLSYIxmIAkDLuybdetL
epPLFO7TkgGVKe7E2oixb3SomAG6Z9zhu3PNgHuYsOnrXITnRrM1JcL+LEJGa4gxQx86hJPFSj/T
DmJuKiqMknaNaYp8rRLM7IPpoQhg88ysp5oBdCL81eLveUJxBzni9AJCkhpktjAEsNL6nUDAO3GA
OYqHUnI7HC5QYxLrArMAoDmsH+b1bKO+SiOeRedvoBjXZZc3qRDtwclCqAvj5NOAQFsTM7r2jqfc
z8pcMyTBIpHlZT8qNpIuh4dDlxsMFyjwF3kh8X/dxARLwl5zrVPi70BUchQ5NAHL4sjiOVcz/HQy
7JVHgyv581OYv3CZqhrNgQc2cPYk+iuwFyYRiqEeJoCdtGxrrGWHRolONtGIRzADWZT7t3FF7mge
yYI/j5HZt0hTE9N/Y8SfGnbh8QVkc8THzzbeEng7UtIXJp1lFOuO27FdNAF/15d3VWzPlwgvvHVy
E1FRI6OaWFhhiMMxCgwmqLgbh/PcZOcOFy1dnwJTbis1ML6+iAOdRtruHbnjC/jDRMVQ1YAa0Qnb
MWdoTf97EawJ23vHWdIOmov92uX/dH3/I4wqd+Dpkt/jj7ENpXLYExoBCiLdv9XZZeiF8Wu5yzw5
4tXi6ZWqC0i1B4Zs4yL55Zj+VwDeJhiSmNmFdopI0qnH8YPpJYygONeqMwtL9Q1IuBZcBahVegfJ
lJ3gukz+mWyHR6DfhlWk/Q3uQU5xaCkNd6scaqTBQfhAuBaADbrdskhnzqcjC5UNhxzo0EXardvN
VhnjNlKW4Etxn9J+mV66SYgp2lHxhJgYmUR8q3d/eUnt9XIBq0fQxlZpX3bu741JUNDX2+YJjBD4
wnbLYmPi10RkQfo1rD4o9wa2vdrurEYWvRmEdCaYhq9pA1lbItqANXDdw5CPYzwP/kKOBakVXnhX
VA7WNIRR09xr34/oc7GHGy3gjSGcpJnq996NOTLA173ulZqKBObbiVW8M9LYZVspCnmeVj89HJLf
6lAHZfT4UXqiFwBqX8Lu/K+eQmK+9y8rCjDn4JqOdJwhxUNg8jZ5VpupTZ4ql8lduwoxVz34+Bvi
0pd/XPfTiJV3HmpwQFNxdi7NfSRJF/7FWkZ4M/RUlswlkUq4N0jhaCOKeYq8RrPXAvkaR2AfipN8
4w99fwqXPxAjqqJuSJ0gyxCUplBfJAGgMKLzNMhskUOx2kkxxsmhNgWiDW3roDiz4fbevQGFK/nk
NZ9Wyujta5q2wJNtZllYnMjIggSQJxOwyFy62vYOI1+E/0R1JSL/eFk3XqlxO27zpNGHxgQQjI0Z
255+ZFrpLiLbtXlqlMCsOPNhsO2guuID2+YgnTH0hAYMTIMW7k60b99GwIj4iCGCSXO0Vayz0vHt
ioMtm/xpg9OsS2D6kJLcUB+1RzTgxUoNH2lNheUSDgJ4WfzOxYLzagfuXSqPGUUHOAXUpFTobCgL
K58qi5N4XUvRTT9ZD3mYW4xSjkMWAEmt62Hao8WOtQT5vmsichQQb5GM47Hn9ExnC5hJ6nlUxwau
s5w3vFXxvOKtEsIk/v2sb7wzg5qi+lcufkiFaE1Ty2w2o9MtTMLVMb+Za+/Nab6u838ygApRdFmq
IZB1HL7oH7Z6jNmjwC5hmsVMA97dArfLA72VB7vW6sRvpRkxeZmPkLl0V9BU1/rXcyVHZRuPpSTv
a0vqzLbjnRbAsHPRQEu+g4atiPn6TwO8wHjo6Pu60qsVuChRZvdOg7HP/bkbmB6CYYNLlBphxmAU
SZQ9NsQh4QvBQwxYbHzn3JuE+Os2RbUq4LSOXoR+IuhQwECH2L6OpsKECj02QeE+rQgUtqymKdeW
c+DjwlbxH2cZYRMMW8HXUAsDlhISNXnJMhOCJjR4d2dhav1Rx48qjNSvKKRPTVGmxbbgM7+P/L7X
q2fuexn1BPEGh8EPx+lj9ceICZTRCxg07HnrYx6+SDRkw1NtVnNTITzd+cgDPemOSqU2nALMm12y
eHSMbem23TQkt/fIlwWGmnONm4PWfdtrX8G7gQtfI/nubs6iTPNjPdbOrGNg/y8jepchpuNuR0vu
eSCnO+GD1v/wre4SP3SdgrCy1tOrFkwbnnafs8RBBe2iFvihAN+GdcIQQEhtEU0WHr+HSQt8DuGJ
SA+aZzhO3oWjawYmV6V9DDXEjU4RSFdvQ+rzxQ2kqKdflVhuzjkucjWk0SDRDS8tQNEPpDQ9Gt5U
IcPZOfxnF7rQmBXG1ua41vIqptodAszbq5jDPUqez1bbPO+WWlLE1UzmcInqwf5chYltlSIh81nb
pGrqNXQiLqvHg9Jj4OH9IhY/kHCkeiv0lwn0zd/r7FAoQ4pjgpYCZt6CsvZOdJH908kojLTQ/9M+
BYyhS/ZwPQsEXxW2LV46I+jbubGcQijToy4FOw0JcXy0Z60gELDcV39K9A3lns1rCr05Ms3ZlTIQ
B8LppPfDl77HnVHPXzVR3tSDk1DuH0ec3Ry38p0/qOPTF8YdZjdpvqmteqIF7HADfXbyrOTpBfI6
d54f58fMV8IrM0mWygGsRzpYyofUSoZPdKtAPBDtDly1gGBU18wp+QZO742v050uuO32mlRK6hFa
BFiJlMIBhxBQ1vXFMo2+Z+XX7agl3eQwq7boT7MI3Dnvvq+BykCydIY9oJaD5qSrxvSZKtqGJr5b
SX0D4VOs0my911Gk4yhScyQYBch9tUE04YNF1KIhIIik+aBlqrnYcCS/Ml16gKl/rWnG68sl6dkj
OmiHn+SCO+PAc25in9mopguRRlhBt4dkqGQbZT2IPtc9q4VxyN4ye+vNLfA6rFUfCaCE1KISqJHS
mlRgqB69gFAJOyXZpcQASCZ3n6Ox+kB5TdQ78JuCco1xjuBqpqsGRK5ucs4UcoHhOcky8p/q72Wr
XIDyMmd0zAWnrxdczaeWt/R0Lo5FzSLfxJedKjyLKDrnzFBlP6RMPqWIKlISY7GBm3goh4kW5mZI
614tkpmQlYdjOIy7405SXrX2MYiIilfWBMeJC/FL0bpiuh09mhqP7ROBBolawC+RsF1RexfIkrPR
h8aHWfxa75tXbU03ZZf4mZZCsXx6exG++ISL2i/xPC18BoWl/CfZ4/8huxyln4qCCtu1rvqmDZNA
phruRtDqQNkpuKKmLmeloHDZmpWztziCX+ZhRuif7cQG6ag2OLAVNVyQjRWX/wLPfohx6cn2jvmY
LMNQW2rVeSQFrvNK5cHiGxzw/mqrzrLTwwuDB0/wLTx6rE9bi5kynvEid0sICjy1VKLOfArdIqR/
NjbR8kW3LP/gE9kvRff9rP+RcyN5RGpt9hT13FmwBtbjfWJZWHyLO9PrYhptfsEexlVTU9wyGHam
4//eNN/D/NnF+dMaGvgKBUgDLZJ3FKoeRFPJHZSTjT9vTOV0c8d0GRNAcypHh8mWRksJU0YJNokx
zULLPkMGbeqTDH/Fvg3jttkX1Yy4HhO9N2q+dX+gazpn+F4RG66l7z6rimmTdV2YeR3w9Y1Z4kqx
Ij1s+9LfZrXzssU9YQ7++EX3cMAbPphXw08NqYjQb2zqpdS4B3GyYfwzU//hmX9Zo/aSepkWzpge
d6oBAcxsKGTfUEYePJfpoYpV7D/DURTp4vCofS7Y2gqB5FrvE89uDVRhH+O/aeJCF6N+yyfVJXlz
rGK8zvmqUEYapWLxsJ/4lrib1BbpjA9+RTwgCRvMDUwfzMoB7p7uHPaEt/smT3dS9M4AYuZ0Vc+S
W9bO/6HpKL8JQoTEAreb5lI5NDtTMdNJTypRZ1AL+MaZ9lPl4eAUfgs6cTwkgXy6OyLeWB5kLWB7
anwcwIJcJZYtnIgU1haht1Gsb1LC8Z60vqoIlXOkgtCuBGkXlONWUWn0vFVbr7xAvwb6mVN2YV1+
0JBD6TAIyOMKW0jL94sZ9GTg1s4CsyKMk36Ny4gFna55YTj+xlMtzvA80J4xfNG68UraUm6RHhzM
dbPeyQ5cSEOYTTAoE9kxsi9k3Px2ln3cVaFDR2iV+iJWt613bWKbVkaV+1YrKFvfJCBJAnjJ8sWT
Y5SGp8kdBGPYrKSWg1ucyATl7dxhZ22/0/nD7vIom5GO23+QJLlKgG9YZOf8EOhCjsv/9Q6WEMqx
dbVhLoNUQj8zyLLZTq/bhPWiGC8ilWCUy31saYKEzpdDRnYf4liKEwofVYSpepKL0tnidd8xI+c+
k4ojiFRKLXkHe5FaSj9ExG/8bDdB55dudEPrQ0AyMDBDxdUNQOBnao2UlN//a/cKLEJ9NwbVPrK5
YT3Asz4bppyTRxvFM0bzA5UijF+FTP9YeLpm057I9LZPxH51kkbp+f/BhJ8leOAE1Ei75NNeAjDI
nXaxuDP4u+dRxilhyu1JnYBsKpwLoAICZjQNtqJzeVGQ8YkRSDCLVENNC5GE0dgt6JUeTdlhllpC
JQGQouMDUsMw+LhtJVDSpRgT89/yj/+A+92uCbwOFXqGPfPASyF/MDdV9G0ZmZjjdivJj7lf475U
XN7pKYdv1XJxEHsDn5JlWOSnp6cje6gLZn1c41NivWfUayIaPvv2O6kOiOZQTSbWPhWfbMCVwq8k
yJvka5/WcXzUYxUX0aJNk0d887PdVnE1mH7/x29FtVyaRkbJX7uDMBlcNO0UB5F67V+sqRXFgO6t
X26okwX1ZCZk9m8DFMPhdXuq1SEO3du96wJ58BL4SomWrPpgzbBKU821SIjkxg9CIC9kb3UNI+n8
bxh/geQWCga5JswMpUN/ZUMOpSJuBuqZ+Qsl7vmuWnOQOA9essUTnutNJzrF9O4IWics1FBvinCb
ncxu/6b2EzkTb/+anKbfx/jsw5xZw5F/CDouu2dEzzLKZtcf7JwWN3IfUn2xK+oVpkgVfc+T5Zlw
rxEEG3o4EsVcEhfqVnJfL03nazexfgxstco781xvv4rpcymNwG6UwnCd/1Vjx01EeDPkKm7NpzzB
Clwb6f/oFCjFcQP2pDhwfw0rgaBtnosUDl+U78PTvAfCkTyUvaRyPwKKqnS3d8Tv+8fqs9U5zyDd
WUSHhyqt9wYfjI03JHK3G0jQRxADQRVjqPSLkJCF+IBxutmu1E2ULjg6qVHDFfOfKfiNE1tD3owj
CDCrrL83l5vEvv8jiB8LS4ZcCFrA/s6It6EhKdku6RCvTP1oizgE+KJXD/n7WfwPiBGKMUS23QvK
L2a1fpDeyePelAvJsS6gAVOISvx1crsSIiC2PJQ60mkyzZtUjxB69V1w6Os/wW/IOX6URGLGY+g1
Rv651B1Zk5mZzvWFSF3spFYjeM+GwhWFDJW3IvgCxyu9NojJnO64ikwegEE3pN+7razWvSEVaJWt
7HMHV4IHWOp6CIQFFP5tXoSVBpji/5DybP8ImoCXoeRjvGV5zTmaiahDjUupTVvj/ruUDhcqp1b6
4uYImwNHqxpn4wRuddcA33inPNv7LrX+rTHKdUmZtM5wcKy2XhKxiEMV0Ej9ASefXg4X31Ek1kJx
sZuU5ORMrk0aV151RhFYdKPR7bH7YyiOObW31konJJ31z5uenFaIzOS6Pi4TdpMAeEpI7FDTlgxh
R93CGoXny1ts7rbPggQ1Q8LCpeyLW8ZHa437sBfx3nKpOgIfvJnsdll0d9wZSCMTl0eL5LZYiCbH
f9KegkAdb5MRS+FQTvX6GyhAVuVbLxYwCr9ihodYMuJ4FJMSSya4r2mZqeCzgrQzy88RdxkmwyvQ
3d+ERR9YJZfQ0PadwrI++9QnSVPNbPwREFKgBrmEMJ4Oiw4gwuVLinkjaolLYZKkriWXqmMHrLuZ
67sJScO5F8jsVbwsd3DqyxA4gMAk0Nv/jZ+WrTkn93W2g4HWm7btQd/NgrmWtMGS1ZsZDozjXyGM
YZ3LtUzdQVE7XpjWCXxPAKuEx2IY2Jqlo/W5EXVUbaNFQRHWajy3BvBZhgZsSuec9UvhKahd/BOC
KRIAW3hWntdlCeaO0/TYdSxCVjNcjms9aNHFzAYhAEPFQPievKuRrybtyCE3+w1R0Yw+4+VLqH9R
/Tmy/ATYzc0lB6Bt9ztegRLA1dzxr90NCqeHbVjocXozh/aQuVTHmdQ5Re5YK6/NKJl/04IpTnPa
grlAQVHQ7pWGgrDrBapOYsW8u1V33ypWK2uSOVeChIbS+MCBf6mwwOGq2UPYj286YPry5/gc9WWV
5ODvnOMeR0v2JSTsh/E9G8rDk4sGY/+sFR1qqm/6JLKzVl7ZhmJT7Hy1IYP7z8SW8EjSuSgdWKBN
kkzSXzP8uE1cxQ2HuuPqPdkiZj1cBM5Ti4PcMf0m42VxDOcULiXDWiE+no9BtBe05dpQnzkCb6ZU
RMlsA7nFI9pEPud8nj8BEUxqbtStt+yDpMimWqrzmzag+dtXFIxFYa4wZIO+DHZ5oEQrzRV55zjx
6hBiAiY/r0QjFftoC0oFAwIuHh7rbc6cAm9ouXMwAzBIjDg81VWthimzT/pgqsdfJ2ndsLtNmIch
dCUT31emtYP5/4iE7Af7n/UoCG/9fOl7ZfcJipR4YX5WoUW3iuB+F4I3kzT/Tebedgy1jTIco0Az
SypcSfS+/yZ/kpfzh+zZ3N1xF2iWH96RDFLuKdEWGa9djLUZ0L5Ra/VFFRBBEuRSZ9ZrISjJJlYT
XSILMJnLjjhL7ewBXY3s6e/RURvGwou9nO8EhRLylNB+d+hoatl5pVu5+NFs4CQcIchRAt/z103P
h5JTvZjv8MMV42ywkzM0Unh51h/ozd8x7gcc1sjpXDjPDslvI9xijBui6mviAzsezpIw4+e0yuVa
zXZjX21eRv6czLHQs7Hniwf7FBYzs0qivAWTY0t0+ffu4CZv3QKubK46glCM9pDXLmw9eccJ9WY8
TkRXJtCpf6ktMUiSSRVtHMENJFxCF41a3M+PXCKz+2aLcWDCCUnNNHr9KlUL2dk2QgujSCyQEUXW
cED+IrNtIzAnjvBdBxMHGHJUWM0tUQoR1eCNQFa4Cd8KpwK3f3RENGT1KLKV+jIoCLnQCEt3Y14L
ML5SwJRaHK1wo2yXxgCP//lcInX2uncdwsMHUskjVSfXKHMtvBiHV1gaqlCWW7/T1bmbKUEI7Ngf
fvjO6eduU4liU6cVyzMvTuip8Uh8pKxX0zzeGOYep2Z2MhI9+Nu/i3uuVZuDoHFXIGSjgZkvzbXC
MenV0/0PHOfG3ktWoqtxsS1DChF0EjTv6/lqkVh98IB+tatscCMG1JhDF5TFsWMQx4eaRgY6iX1c
7nkaJ7ZCCklZo+Ne6xM/2+P6I3L702dFq+nTsDD0IHP12/hjm8f9rhf1erG/bL54FJbHLDg4rXw2
bHFA02WfEtDBjVkDhcYtGbZWLOXDXkPC6u9lMvg4cyvxSR+JXUDFVnX5Cm6mS0PxGok2nmcZTsEL
otHmSaS2O2KsXRhlsqG7LAc/z2w0yhds8pH3cSTIy7sFMrScfzithnlgHJ8CVMvLEw/idtZwjdvx
uezpv3w9XK0F1K++Pc0O0vbtpWLj0EwpyS7d/e9uC7+GP7GBWrt5EStipVi1wewLw+n96GPLR2bb
ciOARNntfoU9z4u+qy+NUJQsphuFWn1OsjVrv3kHVZgqvZnwnQdmSUn9grJiApqdiBBu20as1MkO
5qSFSnhO3VclnxPeDG6hgddKWqkHB3Bg0DIL5gY/siIGnXdd6MYrQpFM10KXCYIuwaZP2sAgl+25
4Q16+HViXIqmC1MBtqojo3GPRYARJy/voREoqDk3rhZlam/Mnh6jqyao3scfcLKcGq4V53HsqPzS
tuXFcJH4s4w7Ufv0Ngt/qU/OC7h6JzqPDl59d9GfFvJa89NVpfWopvJ95X469sUkbv1k50l9uNoy
xpHaO9vt5MD2V1+EVOFnyZOvmIdhw+FPlPjI2mhYXDgUMZJ9/dDDvqkr6hHDwAhus4jJIuGw/wev
Q2I1pMEpaMlzxssagfc8ndpBrElqFgxWhn+45OaYreiCcXdl09cVMQfeBC44MCFGhS6WEihkSjo+
8Kn7nBYpoP0j/ejsQTBe2RWock7XMGf+4gupsZ/ifu2sVgG2l/k8RpUTqSBdQ5Q6U2uw3S7WS7+e
sr3Ez+3G8AoPrsu9y9BewoFcD0Jtiz8Po/RwGe2smiLFvpnroiqri8p+WlgtO+XCns/pjU5Cw9Kh
7f1sG1Hd9d7YcFfBgUlOD6FCWeCbTtA9nh55D58XLz8xJHrErPG/nrSZZlI0f8WhQW3MbtspWarH
a2hqsKjqdIF7F8e1bChiQvkFAxqD7BgIKjLOhGAqAbxZkVuRqtO97ghU0hAF9JFaoqFy9ZVa4RtS
+d0+NbWs+r8a+kJY8rl4N3kDlIPm3jzAb2UANoD5H6Q5NsjTxWZjoJ0JpgC497tXcE0+lbnwJOkn
ca8CYkCUsJbp7yeIQ84q4FnOyzcoRoqa2OXyWAF92/KJipBCkJdCFHeg8OwhAVPKfgU02MA8PKKV
z0rNDcG8LJH5Y8jHFfYJ4t5eY4hJI+AAGiyGEBp6//5Xcq9XCm5HM5zMxttFc8o+mLmFQD5YPh7A
vW+IgIHr8Udf9iAEG9EcBipqWHoHRy+mP4CUVbxdMguQK7qZmdPqWIoEo0nEfii7pU17lR/5A0u2
sv5q1KwQ+6iNVqlFmX0Cjc2BZmQW0UfizzMiUVpMdWUTYQ+OhSQHItU2yHQakA+MFrbEK9jdsrx+
nyvlV+0I/8hQtvYWpj3G73V+ckLJaYWZjdXcHDHQgSIDJY2MWqRAaQ61lQTj+4+oj7rF9GCoy84P
N+Wrasq/pSFs3LEVCt3khVldjhgmyiPdk7kPY4bZLS2OmGQoHnjCVirQZvrXzIMUNKnAO3oYcfqA
S1uyuVusAWnajukORPCJW6xsS9vaPUK5LXA3f4WeU4xXlMbEEttgARnHkj1WOcM33h/wgkAigx+E
TwO9afK3iusFtuIr6Tdqc+4FbD4jD1yOCDA78nOjfz9TcKufGGVn1PD2QEXSbNIhU/cK1eCwrzmL
7VIwEkaXcvoW0Cl8QhKaguQih6kkZyl7C6q1LvPYeD71OBHWw6hl9fN8CS71y/pp5uOBxgKq0r4F
fq+p4JKW9cdl8q0Rj6NP3k6bSM6QiopFmKy7ddXjwEbBoG/RO8Y2Cq2SIKsN0aB1o/bjhDewPs1a
X18fVOW1Z+4WdOQ2FkVp0uQwqseuP0g8rpjwRaY1irAYf0wI3+Gek4pVBHIOO00R409Uf4N9Y8Lz
4u8xtCCPS5GHvbQe16uPzoWm0NZcOjqtLRolM84fElhchdQa6aaPf7hxn5dS+1vvuY1Aomt3xjQ2
x9OHRF92R5mVF6hploqLSC6po36A3KIc/s4nWYD705WXTIzI7dz7d4NF58d/Ov6zhYKWZk4Umde9
42ZFrq1ntML0IwsAe07u4yXQIsaTsPURgyjIw0l8Ma4/fQq3/rsOWbHv0z1W16mZyMu/xP5qW9Qy
IbPuRVoDzE2bFisEJD9PXeiRq5jVlYv799HfRb8HSkgfA39qQen6hhQ1vkhWwI7Q2sn7pzpTumdi
HiFUVmeDzeZ1eFBBGZwUOvQD+GoT2Een2QEZaYhyRA8AFpaTQhKW89QxiHhY74l94CZHoNrybtEo
rGfIctnl7vEmvrfpJu6Kx/sZ/YdgOygPZOlAbKEb/HiLwmzUjjiC5G47nmdZTRdgoGcTlZcD6RnP
RSOtnzj2nitvG9sWmgZmT7ySNN0GNCEk+Bm4g9avGsz2ver2U6x5M5Pcm7QsTkg+I6OEBsz1mD7b
BLCKnSC7ZYyooP4YMWloCjYHR4DplLj4x4Ij/Wnqw7EgxREHHOidijykVmzL9HbDJP3m4c1Ki13q
Vk2NVb/01rehioFXbCb0kPlM9j/NzjRUltR0DQWafzzDjrgcoi+XiExxd8sPN6PQ3yZjyAIKp1Bj
mqhlfGPrYWghGsV0YoFywbcqh+/lYwpKRy8xYuakAPhhVvxbuB75UYIKtLhR0yuB+Tw75a8TRbZc
MtxjY5pc38XMdEE71WBkiflUKnZJmm7+MWuvU4QFKgR2IIzmfOaY+DpnyaC8RW7+EI17hdPnHphz
V8wAvSFW0DwMg3XYcscLY9gkHouSwrvSWnDcQVIjCcHfy//5NJFYb/a4e5qio+ArfYmo7a6iI0Yo
CpYOkWQdw1dNxl/Pb3RAYLui/25arB5g1FDwP9Nd4nTtI46iSsNuiAtnWExfvTTmuNviXuiLrNUZ
7Y/f7POvRDlSwYuBSMiBF9ROFt9ANLTl7yQRf2JDTtlM+fj7VGbpC4Fv7IY4iaYrckjApZ8rtA0E
HH+3nPJf8KMP6RqpePDmA8AkYb2bKMedPK7UDSLrDM7OGttPc0sRGLNxkUhxE/tEsO/MYK5WdI13
3j60J44dcH+RTkLln3qboOHLFkGjHJ2HBSwu3uhuq9afFjMNqERtsYfWAyu6CVu0tspmB2Dr+biv
ALj5acJ9Sj7wTmGgTaRG2iHeKfVUhzpdg0qiZXBe9HrxZH4XLZGZ9JsZbk/ngKpHeQQt+gkWz0KR
vKrTOy1V/ANCOl969NO5jktjcigvsWfqXh8oKepKWUqtIu9KqdXPxVBSswnPvblg/6K/uX1t/aIU
n4OjutRGWl+IvpY6SlZCIJB/Fe/p70WKrZxJSqP/HAlPV5s86cyckpBdh/MA6sRS4ClhPKkuXgDp
B0xHGAtIQKYQ6ZtvwPo+nPe4yFdJt+phyQPUbjbGt1+KaN8KUi8Q4AgUM7HB9H9mm5SBf4bZui9L
HYlbcCs/fZLFvyvDCrGtEOsxjKJGutwoAsWM9Ol5+vQn2MCQv6Y7kPpzDBDNCaoAiY7ECzY7h87L
gORYsRpj+DwvYQNun8B1UZbJWPVKixaKxZIKkYs/WeQrikPvK5EDhk5Wi7ANhAZs+cLcAN7UtE90
gwTd0R0okq2VMiJaWL9FxeMDM1bcOwTVemUZrnPll9FzHomStwSOyYdXEm7vZbOUpHKS47VjKSGi
hg9ef4ud6nldfnKUMcUlBC3T7jx3+OeJjR/qzbBAB8kd1xSwhDgYz9ovLfDDdFpc80+DXDTPdXE/
sRV1ZKtnyiWRnKGQNUhldcpgB9Zbtf+q3m0DhkBxkzpPatK5pL6P6JcfvydGBNJK5IpBccV24Xss
vA+JBOenGAwk5320F0L7tQbLtd0W+aJgqeVPwkF1xmIascBQ4xKRNVc7s6EFnb1olGQA2bkI7Lwx
O+gUoHmRJZMr4WTA0LnbqRTFty6v1ahmQXQCL6/aM8APWcdpdSlhSa7q+6G7yDKxoTLNXLhdDXQ2
A8aAd6cVp418KohIWHOCFOAd3KVSTdbKX1DqK2BzURBWjAOHqbDl9QwSJutoKEiPZ8LV1FkN4GXt
wtxifGjOKbHmm+Q1mBWyNAQjFaH600QfMre2yHdCL7I7fBKL9pNFN7dk7OaMn7Yf6f7FAFXeS+8m
J+QLBBnMnZYekHlPuiIQbAwhwdczcmuqWDt7FWo+27FKi8ANKWQZ7JeLQEjdHv+6T0+fjB2RV+0A
gQTKb/xrJqhoAegrHIwrnQgfxqPcCiHIrP66WN/D3hLyFwwKK7nVtYlo4cY2y1+7olN9aVHMNuVL
9J3+YW/M/PgF05yrUR71zNf4G9JQmdJqhjFE0mZUfZ9gmXqBH7vshK9MsPz29XvUq7NJTVXtdD2R
N9r+WBZbNPMab5qg0HaLRsbwHY987wl/d/+3Oh7u/dtyCzYRbiYVRZs2+1pTFF4zVQXSG/mCrzbR
S06V32VQ+JqK2435FS+6sHXWKDWNYqV/nAciYd48El+bzDl6vr2tivBY/RfAqcExtxsIsHKsESSv
SSoNqemmKexUwWPZihJTLHdZFh5PoXLm9hunJHRec/lcMm1GrklP1rbWHBiSGsnXVvdtqLA9Smrd
gydhpLlUh2cfQMBrRWVdWnUPWbNsIq0bU0h123hZ81tjhscJhlWE6SqNd6BmzuffZBmb/qT3sKO6
/16E0n611bHcNYuV91c8n4FU9t1tCBSB1W2I6zD4VA/AYjP3iQOKqYOgt19n53Ji81ej24N6Zt0n
rp7a11cVkdAjoTAZEzWS01gfDroWAirkFGio/UsEbdFlkRZc/QJLNgoi0AhK6ZjWUEJ3i/jDYJ8Q
q3VMWXDZ1kEu4rMSiNFuK7LM6387zDyKnJVIgfKzQ5T6hIE0VySARumNyHNaHPIK5Ep+19MK5ry4
UVk7kPpMBKx/yHo5kCrLnJSYtMARcHMvv0YggZ7ZpOCtvJyWICE0ttVKqW6IhbJXiazZeXbthqUf
Y3qN1YTIuVkDYgv6aKcDxafLzkucvsHtiM6Ra/zeHx+uaEfNoBSlu9/DZCs1DzOjkrFSqIRgk0f1
S6jc57ffw3vWkMeA7ks9KvlakCDVa+Hjj5feRg24pgzeJKfXboUH6l3sEU1KvJwXW2yMHX681szz
vFb335M2UYjSckAYl3lK5paQB7hMP8uioSB7AgcAckAIhTy5ACsOYvgNoFEWcW6HXukNvqa5tpJW
/kEeF3cV1pHlPk4u1AJuLB41/JgsNJoF1dXqxHu8wHDvkHSqxtujCpiabAEm2/PfHg8XFg7JSN9O
XFNu9sVnzgdJZjme+m2G4Ndl1LouM1IqELXPMPCuyXZYN8T4I+uC8bwXMBS2Rk4S+L58JKufQASJ
t0TetSFeICYUENyRD8ibavGQAgiDbBfxQnKyZ2O6XJP84bXKw2PoGAyjuhDheiTt5YxpBAnc64Xm
OTbXnHmN/rCA0xQQIZGf0B8G3K8ATGNNlse8yikdAlHAKezaMwF3x85X3erfRZ7VNWtHpl6MRHNz
6x8mUFN17ba1DbV6oyehypNE5TvZhuiOlP9kzPTxaBQAdzScHtoAXFAIqAIG90AzYzS6rUnbLmei
/BgMMm1qA4OLH8p1R++8SCwiUYzQ928TmVoz78Pgj2qqBU5QWl+OKj8g2ygqIX2l2S9wVirn83ac
vfEUO32eVBD/+qG8V6phtd2nK8nLz/hiQlxTFcjcslqhUXi4rffLdP5TkNVDwEHP2JTkjyRikO4k
rvatTqH5Y+DKFIHG9BuMLpRfB7JVrM572scyDRT3NNlcfTnxpGwlDx/15NOQUZ9NM7/+We19AUTF
3VpbNuxZ67D7s3acY2PMUvvI5HUw1s0dy+sWtlfOb7lnxC/vAcRPtlDs1QhpRoMBO/+xazTkTWhP
KT8NBtQDMorfdjoXQ1CHeWrhkM9FGNxKN9FZ5Z5JkJe5NTHNH2bxxgLnLmYrOCY2QqID2/B9vAC0
PKVZoIOcdOllvnc7U7zetmgQGumk+0rwe114NANFdigmnv8rbmv6rjYeQ/FvcU3Z1uRgAGmmrPh0
A+bpIa6H94HZ45m2vyzwt1xrQXd1HC9p5st1H8bUqSyyiG6y79vjy4glgnDXRn/Xgwm0/QzhuCDc
v2Yb0N1x/QHynkMe1+P2UtI5vBc2CYRg5SgCa/JxeYDt0h4mNaKZwsFFndfnRLzb05AHU0HoJRb7
gxu3NE2XXTewOnoLe8gpsXBoMLqUI5Pkezk72OXEizNCqaH5EPJV6/czHX7BbGfJmIOZ0bUwqIsu
uZMbXVPtcjKuAdcdSK0BdOCFHOLU/eHIc2rEQTU4i1AMcWMcDq89VPGNNP0+Ou3/NTl7zAaMOyN+
hILL9SJZbWUdgm7lCTIpU/juTkRnHxMN9ARjulCJsrww+51uBEvVqolOc0/TPffN+8SogiVAdqK5
yGYaAMsdSnsbgDTQJFw6+HMMyGq2XkSNGToJLjBwLwJ0zdv/XK/iqvK6OYoYIgtDtmrDrCj+lIme
6iNwcb0ncRh+xvMBYwnW96XNyJJEstmazZDumKVQRmaYTxTiP61NxZ2E77UPTL2ELBvT69Lo6SWe
6OEEYcnxcLHAO/OgSmDbM2uyrFjEKmKvhDOUe2EsvhKOU+KxTDZ2hKRc+ysfX0cpXJDyBg5rfJi4
FoMyYZSBk49BP8xfn9cgqahm8CBhLCkkUA61zhUB2yfe/nXY5v+UfuXJAxX/ZHNGY0M9+0/9wXNd
eL5Ledoo9qAHw+T0PjoTN6t0j2GNK0EluJxRU5DsnWyf4iX6vXhzuzSGpoQZa6SmL4TU5QnB8y9Z
xsahTgTKrTMOWdfNKb1R39SpdoEcboTwb3yn4gPWTF75wUVBoxF/4HUAgIRrkmMQ6k1nOMu196bu
ck1phRrl3yVhqQFNl7PtkrCV5HbgY1PNdtRtm0KJk7xS64OdnBlF5y0gZYy8nVp3lrHtLu5qYSGT
aZ4T7t2tAEIXVmfhqhZgRx5Z5I3Ypq800XQ22Ot9xygeDGnwhIHwYS5P2ZnxeIBdfdhxYdAo3Ca5
GHNz3XS2D9lthjJlsy5PeL8IfouHg3HLswb4I5mRhjwatbHJ3TTvG+IM3K3FosZWoKernLhQSG4t
58zN9bPXi1AayLZwXICDN5N4BfB7zT9gBRknj7fcrWvfX015u4StDKYICeOCc4c1vyZ1ksUgIL13
v2hGHbZCbOFdCBdv12rf7PETGnrPCrUgCVtxs6e0yCHVEg5L/qyIIXT8dkYxR+JWd1T3ztzmIIp9
i92xdaVauco5g0vmx6hKUBU4fCoUDk/TQvcc8if9OkcSqlvPucGHVrvkW/0rxUBzet4Abd6eshxA
y2rAwaFohoWFBMygclueyt53A9D2w0VdEHzbhS3UqnoOWfeYx4Fm53yFaUar7uIv4VC6DVWb5+XL
AbY29d9CideZt0ysdGX6YZRE0B/UUcpw2wjs8dx6GTQO+NPETnQe+xzPtbUHdQKkFAF9KlgrQ/0z
Q/IkSyGDDPedrOnix8R/YgjScSPrphZskgtetUT2KxN8CbVTUnv3FW4j5FsS0mewLtcd9iK75o+7
GGKUlnHQ5Xowhm4TiaoG6WrOYO5mkGyvmQm+y0kJpxiAzam9Pewr47HXy2I2ypZpZdBU6rAe5kEG
Mt52BBN+xQYa2nRcNW1qw1Y2h6pD3hO36FaFlpeuY22M5CcouooHoh5fb289Cvz7T9cz/RL/EHA/
216kzf6sPe0v6Uo9nJjXUrpADRk6SKkbEUTb96Sk948ug9ilB8MD8WaBOdWwRoVnB7R2zY1Fozw8
qaxOG42WefypglJEUpPMXjSrVGMZ3vwQM/xMVB9BXWVfaFVv8ZLv/xfQk4MbxEJFyi0hz2r5LJET
sXY3a4W3AAcGuhEm/3byXI09b/+euDvfVBeJ0AOuoZKy85kfVoRMbwbamKa51DukpHH2kIQTgI/q
xqkI34w9M30ODFurzDvKLPsNAUVrXrlTu8KAPRksiiSSf12s0JXDu2OZccxKW1mWlwHoXLJ57mC6
SW31VR1SMATi6z7x8rVoYeYLzo9WRSG9bOjRWZy3C+WG9FFmjkTBUCt31hr0mrwknGG/HSE9v+fr
GcZ+4oCqFZOyuCWDpeTUHlgmO1AFgI6vxW3HVzNN1T5tRWydVbHIJlSw47s7gLz/Cp5XvcrHqs8Z
Z5KU3COtIYv4/H6/7u54SIJ2nRiT1TgeHuKufT+xHv1jaUOU1M0pelBsYl6JrNSe+4ymL7R7546i
KGMUzgN5l6H7b4HPeYHIc4bsxT2mH3PpE6+gt+Jcv/iWJ+HD5BUWEzKcrfSX8MxQ0yLaHYsUdTSR
xo7WGm/QDZjGHWpf573++sfQ/ryNAa9T35kg42P+Wd8jYifhk4/o3IPLeSiHZo6OpxxaJfBWl2Fw
6sDApuUsPFBgqDXssgAgmJ2OuIm7Y1vKcVGePWSye6Oz0yg2jr1793RUkjs+AjUtOQiymXZC5Pkt
3/BReW4XJiLY481Boja0SVIClIkS1y19klRCGPkN0nrIQvFFa5inVfGdW43ANElDHb2s33K1ybmA
KuyNM0a1JsUxi5M+0+P83LYQztOhaAyVCprCCUQOV4O9on1GlhXeYUtMsVfkvo1kaeAzMX95CyUq
4sSwwBjr4x8Ns1tRYcq9PJ4HdKba7xSgry62MQq5MmswMjUq55bD7Rb14r1/95SroPZ02ge4Eh88
y3p7o2hjYyRtcZYan31UAiwO7zUsbrMbp6jDHGbIoGn2Q7xNcRWy/kdeDLdSLFD8cLiRxo1gNEQd
pTwvhPqDLJweQA9W9V5xXFt5xh5x93iQok3BwXdbdUJzKmbg6dz404lYwKO5YNjkImKaOsXSHEUw
GMYCuolOCP/ZDEv73441YotCKm6n0zwxGzfvKxDsPjeoBQnqN7BLRYk8toVEEH20cIYYBor6US1V
2D/38/UPWaKk2FkjS6JzBTF+dZ1PKoJeXEFODE+W4CXeRlXlve3Xnttp+uEozbte1n+Vu7s4y6sK
KGufbt06JRmjJUiujW1snzImbl2wxPhuujGZAV5L/qfqBasavJZEByMv8c5HLGhciKSYnnUc21pm
6M4htTyCZTD5VC4ZNrAlSecYZK3DWL5v0SAuzjdiZA41md8O3oxUEqqhAWRsx0Wxwvl0C/KLfsLE
DWDZXJfmzKfX+Q3aEw2HjfL5lhLEFFJxFT0V9vyOTH4qQgLEvreld+QYA71enYckiA6tZOfac+p0
6xVeCsau/SBsA5vWsSrXdpZbZQgd+lcefqqm0x32lNRrvlzlI3GUzofgwrV73q/pk2UK4JUDA09I
oVWQjnUd6dfz79RMCAd1Bp+844qhs6QfjHY1xhoCW8yP1FsrKrjVzaEnbjCOa6KkoqPD5e55+eew
ytPgFEqtcy7TedUCgB8zN+8sk8k5MZUEYZnhqjlh6hzO5X1DCLKQfYeB9o4LpJ3JpWTgqycC41aW
OLVR3u7ADIyzh8Ip6dtC7VLLeOT+TT/y5xY0gQbEd5/yQMNgCAYomnEVekDsyFI6ucVbbwNo1Jfa
aUdZlfMg3Z7LaG3471KmlR6H86otDDCUHqguT3n5pg9ZDfR4GZOGLydUwg/7kqFhtF2UysG6/mu5
9tc7e8hTynAFATRLeMX9w2gBsihSoM743kDwlW3gmeH0BOjvmizm1UEw2jXpnh3Os3vunVDosueC
014ZsM75ONtjhzuhULfgd1+GShEvpGt/3dy3cXVVqxTh1jLtt6L3rARCDFQsdNOxSja+tpl6+ojW
DJAjF87cMl68nOcH7g2sMAkKW5GzUCJC6gMQN73W3KxkGrOVl4PX03UY4qXiJV/vFEf7nrhlCDLt
h7xDbrSej9Nrk8DnZKl34kpTECOBBd7qgH1OK2SMJrEChtIixfX4Rg+N4hvuOJODlmqpSc9ldzth
9+MAn6j2ienotO4kpJaBDYzGCk/40YV2zUSpfmYf1xCOTkBwFFEByViPDuHVAU4B2iF2JdkJjK0c
l4hyMde97PRnMkN6V4iB0u4+teriFKJhNZj7AHc2v94NhkIB6G8dZyNMwJEjETw/OMktCM/0jwAq
5LX9dIi/A4HchVlL74iwd7khGX2q3NI9XnEcLnsehH3OjVZUb2OEIrGJiHj0WF3Mse6eE+0UVxTd
wSIyfS9ujYV8ijri/bME9Mfx1aNzio7+wywCPVIJwtil90ohJkF/mxifY2TyGbwsLE4VI0WQAhsC
VWkgKSH8J6sejeupW3f5Wt3iCcr9kBkyg73YM5Ojq+WnrILdLhy7k/C4liBFZsOAKZtsG0dV4pAX
d55dFOHKZLRSMP136p4qpo9YT5sYunn4uOorx/hz+D9g5+bSOqTAd8gazqf563Zgv1rHcw4XjjOy
5M0+xLNoZ4weOOBiQCkbMAJMCXf3pzuf92jBTCtQUg1h1TT4KDkGPO986bsrI2Z8PVE5cIygButk
8foBSa0vumwxHCARfWzzFW4jN83ZznM6GrWuEfSVrQ58uJh1V8F5T9X/IfoFOGssuEfIOqLHBzqD
SbeBfhPcYRgqFkeOQF1hlrWzdXFINI/G6gZ5lCXm6dUQ4YeX4j79kdHRnhF7nUv1jmCYQdI/DVRK
E2nrTFDOA2bbF9d28MCNpQpl6vfh1S1rhAKCN4g6/23nqui/qJpw4t7BXbxjhpMb/NnYIlmF6TaS
BY8zquH0ynFsvDhFK7tl84eag0ShJKqIyr6+Dggwp3i3Ok78wfkVEoTTC4GY6cM1I/T15SAMlJVE
+xRvAk9bpQ2YVbihoFx68Ive9MhoCCYbePO9p7+DyW8fwSb0KcRGEuN4FDHd/7cNJcjzEYbYg9iw
rJC8K1z24swyYgWjVFzYnNam1+TfQxzvyJhrOuRW/npyrprnm9erIxPzI+TXRQyxl/xnZUM9ECSa
F45LYSCvUqqI3UUYu6r5YDDjQYWCV9JP0qwB1hI9AVfdFwpgVki8nG9Bm9G0MuVzs0lUF9d4wYbf
XpS8TpMi9/q0rXW35KZZJ3z45d/zKK6FqLrvivWtAc6RA5DrhGSIT1jgbt6FVZfEjcWnZJ5xCWlv
G3lCbAV5plm6EasrplfmdnFg651ovoPji9BpFpokr2QnvujPNTPkVYRBL3PjmZH/InFkEB0caMcD
IsACYhDXD0brgE806uhLya0gJVEU9xAkphN5yzVZli2/KtUfYXLruBLt27Ogod3kv2NSrZa4NI7F
TbkrAPfCE5mZ5fo9HCIkN87EV/F1L0kL5eOqaVyWZeu2dk3lCB3iu2i7mb440JP8eMfPPWpPXoJa
RG3yIOLuMNc3A9uGICrHPQi3a9ZNRXSWusfq/nz6inveV5fbxLtqmnfWO0QCq/IVt8wCWjr4PN2G
ZXsc3X03Ir/ZFv4bITxp8zS4vcK574XEM2i1ciJyLGE754j/KJ+liOr4Y2xjTGxrkS/kVmzh1ipS
/gWHCUQoBpzuBvVjPtCcocEhwSq2RhnP8lWOFwCa3K4EDujvk/cUzN/+GzI2920XROf/1cjEOd2d
0zjpdZhfX5/otwzSH47YDXMj7Fs8De2DasuuQji9E6GwWStz0VFFvmu+yomUGJRp5gxozyS9jPLU
Al7a40rhlP1NfhUoLRJP5cKwdEi1BY64R1wNObrUPXzQinHsUzB98/TQI3uEpv5gdI1hdc8cQo85
tEw34F1LXRsaWE9SPkBjcS66yt35FJFR6/ZM1sQ+i6VhyIcRDoCgc1sMC5tX2tSL3yY2UkXENtLa
6FjqpIvAnBgY7JZ34/rf520ZQsWqIigkb7VA1cI0AH1o2Z9tdbY+/CSKfGjbicdTTTJ+to806DgE
Js6VIiTf3tmXYSo4OnRz5gJSZLtCag1Z1FBfH3jiRrM721sJ/zudOcy/wpiOwsi7Zvrgp2MQ1Zri
qx8eNp/50bvaqAp3M5bO7BJcnY1k03mbqBawy662SfPMjsdKBiMDeWS28G6eHCss0XB48bVYww4v
cNqJPtrV9tr2BIoKotl5Wj5oZl9+5QszM+e5d5Afo4l1mYmI6kDWYabHrFb34IAWCa+Xtzh/WSuh
KOQmJpo2q15G3vXeOrlJWw1jCuYCZ76qyyR5ne/Jhbpr6GPTiTgUl3f8ANFYEkUoZuCWIcSDXp8v
V3JFiXxH4RuNg9yBR2tNo/ZXhxjeDdr+owEXzU8cwmMYNCn7zRDgwIbIF18ohyRYrnRitaKfHKsM
kdCVpvUAHp4rLctc7DHvLEfXErM/u+QV7pNWq+ouYjxE3xSaR7yq8vhr1Fas43LyIpQtoRBJ2yG7
CM5zJVABk2bfrZ0O1VH0Lzu39eE+np0bJGkbgFrgi3lZovdXFjKij0XkfTRh8BRcE9lBxpY3Qtkd
eE9HYCXkJ8keZ1FJGCcbzHLPA7u2PP7bLYOCX4IkF4Ha1eTbZ6uwuOsSsEv/DpBpNW628Mj5sStj
QVKLuDSRVocgjo96UMjCGNpn9k2UVXvJgHuCmzsyXe0UmP4Vf1BTXfMS4tyuHyn8HpmVya1+Z3G/
jf5i3x+jOw/Iv5qyh4XVFqlhvw1kf3vJrFPP1r+mQnWEuA4pAaUc8mNo8qXp4r52m2A+rPnSiECY
rhs9cek5L5T7h73J88umn3GF1tBxMVdYk+Y6pCEGHJJzmCBF1MS3Q5sNugcPxJChHROSrzH9OlrX
dVmCWlc0cr7N88FHhK+M9Wq99UAuOPk7IlpmcY7BsHqbE8sxFLklxIhXn0ieSfVn9gFjELuwPeMx
85DuIJxn2ojOU7TLIq2HZudUcz+8RoDDWxZgwhsfwXwZcVskCRQJb0lPecAHsybW0r/YT4/0J3Dn
lHPrWcomWGiKLdU7mxAfsjJvQGX0ODFxiqvU8hOBTibGxMjGUPexps5++oT4rYgecTaj4yS9pR38
nIYBzLYvHHUs0jaGbDcfa/nB3EdOXedwG+Ayk0577I5UPTTmbmrjK3G3AajImeYml4z+vDuiHIOF
5AyEPec4BWYfA0F5KGTnVtCEKXzJYQk+aofl4x9nvXoJY9YXjHcpoJ5xF32e3hOQ82cl5iI/fOpY
xiLGabOAvNfORf0GftT2JE8nNlcddlYyRk7T1v4bEWR8U/uFJCs3gqHJvP7Dqwma9Uwxu2D51aMs
7FnnZWH76+W1gwWXeSFfzpxo2k6RKwC1aRHvNIYLKZ3AnqN+Zpdye3KUYoL6N7sEb8xW+Kczw0Vn
PW5RMExeMj9NWuGCKGZIjuw/4eK77r/SgP+2KuZG8+qyHVfmYCq00I1f0EwWnFN3AkXw4iKqFfPH
yQvubLxbR8K8n4Dyyz4FadzmE2Xgw3DzLzRBZg4Sw2fewX/YrWY+wk9TP3wKpznWu6L1XmltuQbN
QUg703lylcKb9WML2RjoqfHs5vuLzZIFT7HuyBX1L26DjgN7uoAwKVlXttcru22fbFSqftiKWqH0
1SIVM3u+7RBRUyzDf+L9GWchnJYUvn8525TF0/EUpJxQedoOhLk72p9B9S4jR+KyxEOkt3r2cHmg
DS1nVwtaJTxYmEIJ/N4BxKnrIW4MdtG/zSdZ1S7cpIjNDUmiW8RH8rf2srAmnx/AtIuDQWCAQnZV
SDgMkVpIgetLwyRmg+NDK/hPnd70Wpt+R9bgWSDZ8NqT7R0IQTk5r610/SXtWYEEmgI/gFvL5j57
lYDiGzJxfynvmGLonvVvrhfq7fpeECKmbqV5G9TnEBB2UvKkgTXIP6mvrqkgpYDMlfob6ZlsmXv1
cXbXk5riqzSHvezEhh/BOHUY/qjyREEB77QBRslPCAA1easipQHulldz6gePOdm5qncyFWXVcihU
G3UmJ3iVOa8naIr1/R7e66jNr1+6Vz64xsXIO2tXeuqEBzToVGS25ZYeC2Xl1qMUbvv6tZ1l5MG3
/R5esjt78XyZrjpkgLwPm3hgBzGWfizB2jd6ECuWJhobpwOaZtzVQIRXxc+LPiz8WolwNlTzIA0j
Zn+WdXFgxVhnp8sKUCzW/0Llyofq6pMySjrBP0eJ+ujKu4AqI/Rb+X8S5EVSeGtPhvd8uDBAedX6
rwi0dACSnUaq7IulvALuvIj4He2MGF3bbR4NLrSOY0Rhb4n3Gor+y1ptxNvMQj1equxJTfFzterQ
GwlEwh/a6C5KJ/44VklULxArqoCtco1fJv9xnQJFd3Id5ogClCMnvRg/wdihZ8/mh6XZ2PVqv68t
v9rrbW0fT1kEPFGdYmMFrHlm6rAZ9PbMcQb4cTfsCXy/E49QxwrkRrGnhjav0XOEoqdYPsqF7Oe5
c2E6ZjJtXtjo2uEPMsGPTW9UEG8S9bfU78aZbUPtmy1h9p/jyvoYP6885QpGAG/Ii4ZPsVaPDBDc
vEzPt01dA1ewUG/YcvTL9taeYnZnRJZ4N++du81ZFHVADHrZkw1G8q+/P0oyP6AdxuPNtNPHAvLi
E7C9baRCDBEUDCeoHUYZRSIFEjbY5msmSKSs4WTboAE/yVLdzIw/BOWeMfH6QXMSWiJlN76bmJJ4
6fke84YaC54eFQPEhIQ8KJ3MCVV8kXmf0mjhoOoLvVRrfjN44R/AOorbezIvRFbKhT1mE0OyiHb/
8SVwNkcGCWzIg8TA0m2JeVMbjBnfygU+XaoibufAQFbvIfqVHZDReBeBaGXcJhNGKMW0HD0VfD8z
U6EFFQSo5O41Df8hvXQgqIguVuvHBuN4mjgZsxs2gRee2G/WKHXZcMn66MqGTeAhaLUj2vNLltdP
JpEtlBwzUWMFvmQ+Sb9ctsuskPMNn8ZYCsnHhrG3uicHPJNw4bfKomDZwNIWEwLzdEdRs2YnOcLZ
WZ1wTU37JHpLH9Iv/DCCoIbKUhpOvtesbJP9L+ObDih97TzwgtS2mZMOsW8hVEUqkKKYUIrPkz0M
xdKXtR6uAjN+RmFivFNrDM0CA68GYdhysdQTYjyXCqDOMcrNruT+33PuGJC0ZSUL0pXceualEk9p
vTjvU91BRuYNqXRQEeTVvYSvp0TWNTG3ne2h2rRw2OEHB9hRPIyV9DrsZD6f7nGMF4hAHt4S3y0e
5nzX7euekzwyYKXkqhRO8z22rsmtVxEdgtYd7S4rvYz6nGf0uMzJWFtyW9V/v61TawkDtVcwf/QU
KWM9zeESNeNy0cirK+EcVT7winZyXCUg35WG09TJwumEMMaJn4D1BUByUEseC9StjC1LdE6W1Ypx
BlLB5U9Kv6kthevoRx2BH7Ge20kJqyAMTXtY4SjNg+OQiphdQxVuWanUOrBMp8681hHwNzVoJp3F
AHoC1qW0DCMoyHUwYz/1KbFxnzGgJbUbf/Pj30XEH7RN9TQjQ7wTV6KstQHteE7sMe7s/HC5jZ7J
vGyneZV5FgvBQsMXJdteV4FzzLm122o9IxxQHsQgitORitHFIe9JF/Rm1P8ymx3QetqnaWmS4Jl1
cPbe/+K+ljhzIOcxiNGy6FXmaDnhElDbcLK6dDmfgRestCqyrmt3n2P7uHc2Uc4Otk8M79W9IVxT
HW/BOvXTxdCWPH7TnsCZVCpbeKjAq3PQSnT0It0Qokn7NaKXldTemLU0joTeuUFOIDfT4qhytw7n
7RbYvMOuv5hToh3H4UgxyGRZbczXlt/3QD24A1ua0i/fzZ3v4x26QSTjhfY4Hs+imc+dNF2l/WJ+
3ehOPP5akTp1zblvIz/3LPH4J5o4WyTjsuQWZ7XBfeiyCet6S5OPGbhY2TO4IE9uZ/XTPqnqLWsf
fWSsOaU3G63XpwzlNIKCe60KtHq9mj/5ocjoX5V7G9mppSuDoXvGyGHfD9XTTJHRwKbRsUfbwwkF
OyCG+njuXVAy0lLIb6xtBklKrmc10P/mfZK0VOa29FUgA91ckqcyduSh4ByvhEwXt7oA7SU8PTXM
FRDjp/M+bDtjwdRXgmXfo8fNxrdkhpywSkplP8A8Oy/j2MujphkPpM9mYo2lJ0ewoCq1koEsvnVO
WTwyBZEnG39FxDNQUYTGTdztcVM8PQ+oDCfb5MPyX3F09ZMofb8RhPRw109CUO3TNng3N3u8uAz2
iPL1Pdme5Rxs8759Xzn839sbQ1EN3FZ3Te0C9ZKy/kPwXPwXCG0pxsficy7QnbRCy3yFz1HL6OkN
pFPFgBlbanYlJNjfG/dJATdwnCDuSaRHhbdTm8junujMBxSe06ChwpSCVDCZBozCb9BgRktmozV1
K90iT/+U31GAWGpumS2Cp6jQ/5cUBYuznjDCvL5NavOeKuLoj46jaFLQ2MTNOtHFJzuX6FnR0Y03
aextjj4x5Z0J8UI67whRClzJfHQKHYsowvieMRXWC7WrWMnBtlB/ExsZ3OGKt67LfMFZ0CsOJgXb
iEojFejUBNqb+MNESKBJhu1UPMVV3DNBs2nU0dJgIkD1yKPPPpA+Uc2d/Ja762hJE7ilOApxo+XS
+BVFRdtz9cn4m8QQcPCxFNZA/eM6zVXBIoovINRJFKR+IYawf3kFOXiXQOj5hKv/Fht4v4ub4KLk
6Ygvy2Q8mkSg6Mig/uM6j/qqSXX1h+hHzurKivIGMrmwIHtDc4auti7YlJ8R1mZNvoTnm3WSGKKb
oJT3VbHWsuqBjCvZyQEr8c8dh1o0iELP+Fxr5jRZzAwF4VSj5oby0aPFEdax6Iol5Jetwgdaj1oI
c4A6Dv9PmdaY/Fm+xKqFHjEZViy5tprj/NKIEjaf3DhRUvxHHF+OULFEbRT/YAtYJw2+pZM997tu
KV1+qWUUEqkBOkf8zLrtgAx+czqkP+bvLeQGThTsTaZ1GHyfc2vuTpi87pI55eNsc3fL+bClTLGn
IbGE0wcqT4C6oFumD4VkvxchswZSSayO3uAWGbP1BkNpzefJhR8KvY0/dE9kclIRMVJFVSmViX0G
fojrZVtQZzNf4XRCdhLMvD+h1SblgnzV0ZPKYrK4Vpl9VEad1EK3Ird4VgeR6LNhaSAybZfdDKb/
G+fRd70GP+BadWhb89CZWOGT0tATGqHCPuy1gv33XMuZeDDIAoEnEjFXfqLg8t2ag76yZsjlsdf6
qS7GA3p4Sd5sG47Vg/M/ivKVEmDQXI/XP6SIa52nwEzBH2tAtKRpTkJdyXgE9YMpqvzCvz2kJ+5g
ihiaJEljQv3ntL/1IAyIIJeTvfiCJ1ku93rn3YmGShzrzjw0MvcfT4WOzI4877cFaMJSY7WjZij9
8lbJLgLjyr7Wu3AMts2/RTj0TMukLD/wGG6ElMkNMi4PmaO6UdD6pk46/ujiqHtRKUUa3AOONBTm
8eZ7L22S1YmMFzxV1yBizeSyRxVgFq4KgUIR6izAc9knP/66IdsMjExm2Lrdj1ZwmzliCxyNkLtG
vXofHx16+y6a+YWXA02nCE0sQ+O/XbVUNGljxiutI++ba1F/NBLC+p2CEk8EinwnY0BF17hm5/on
++tkTeKwv6v0wIemfy1m+wbKMzf6MbcOx7wF0EhGTsWxbnil2PaTwSsjrIr268VjYzcsrs1lK5uG
CpBDc2SN6bO9NfyPkYcMCuWhihL/V6VhBUAuAxiI3CeX0d2Un5sta2GXJr5WMoYvzm/BtcosKSBf
K8XpJIm+TBtT5tuGVNSKc2ZiTkV/yAaUrxjh4+enlEv1lDhMkhRXL4JqCZBxF4wauJETyJrAL+6p
ATjanVR3w32JMscskx//uSGTzQsxebKx3HDm0Wuowc6h/feMlxrg7SAhi/FgIjG6xm14OkxswWUS
eeGsMHaOUk/AIE727jK2rIcQ0Sua2bN8ayx4B4VfChF+Pry5sixOMgH5A/pj4BxUqP2J6lBF1IUq
rKTrZuwd5nZZO8cx9ajocQfcork5IT+Qokzb7n4bB22V/zubHOcbDWf/yum82iaa93hsFH3Bv9yS
pgNzsfHOcqbgBegeMVFJb9HR45Ox7GCInZuBZDgx4UWFFKriiLqWS+mwU9XGkhsd+do7nUK7xWBQ
e4XvAN0BpfevJ4g2Y0ckO1mHafx5gpXUysRumwwDVbuuG7TS//NEiFQ/dzIUxRWEB2HAkBfIXEai
7a4EFmUDhmGHQV2kw6MY2Fh7OQUIcjwQhfafXe7rv34N0OTPgj+yusMRcIj89/rVTGCbpT3YCWhl
vvunyOkpdbsgTVsVYfEZf0k6r6/fqfUNpIiJSzVr2VlnWiHqO6i3ldEPXieGwYF0VVtT+S5Je2N7
1DBoSkVlpmDKBEiDJnVtmVqRdgSS8SYe9O4NKrffFAvWcdTj1JT197hfW3QUGShy+EhSil+S2x6F
hWHdBnoAM3dJRF758cX9mawd3v4MIZbJ4ME6hyqjlMxOnA/jO/StRXy6a4CiLmmYRzO0AowhcIoq
mXEXfqi6BVHSZ6tEIyolZ9nRGg8daZ6Mo3/5a8SDR9CbXuICZsDZRe1MwFHjodDjPeOOdKO1RaKj
SriCPY5Hpc6T1uE+zh5rRWD7Gy5sMaWKxRs/DVZvaGV1BXsqRqFjTUJicpjiww8qlADaS5A48FF0
bm3DR7G41SvctxuiTsLTYKReHvWtkAyRSVTnqxmNl88gYZHeE/sBaWCTx+9fMJgnQz3XTaTffVQB
obK4W+IhOnmKkqw9mvTZyAaPfBhZkhSUWdsWPjusn122D7lUQfHVG4QvTNaLPDToziYjiTVFSywS
pE5EJuTa+N764dzylnKYzbDocy6xMCU9CFoHMaaYvZySwCL+5ywLhBG98MlmrIPkYqiVeqPktNOr
ydSE3kQmT1323kBVglno2Z6pXr6IxbLtNTTWbCBEdbv6VgZ2n8SH2hxB1IX1ziyyMsY0PcMB/VMm
giVudBaXFeXDn/bU+8PSBkh+EszLznToddToGJXAclZqwXtBZO4ox9svQbnykVLjZ5erSq1kFKmu
c2qHGHwfyo5KDQgKl6C4JO2X34lTVVZLViGn2ZO7DsnWflHX7PswMEacsDRsxeCqnA95k9ccwYOD
7Ma1ArxY8CkrClrh51w7B8Geu95Iayy61HLm7OOaA43eemlB2yyN08xUtFtXGfg2p269wbxlo5Hw
KaslEt0bQc2bJZDraAYNuRkWNsr8gq8+QlmqvZXqfxFwUmFFAc8BSxpwcYx2st1XOxzKzwSciBlF
j5Rzx3XBGDQbNdXbsXi+9R7+OFcRPAGJlVesY0pleIgum+Bv0j7CPaVzMAOXAVaP3o3RhbfzWOwX
pEj6tWyMj9oZHTGWI0oHvuvnVwUZ8WQ0Spd7GCC3UidSLzWqCGXqUR1akMholnKQpiINZ8ul+2mL
K0IWbKal79Sn69XIfhUvRwUObPXSJIQOo3lceRJ0OQiBnmaNXTZHklIADFueipp08EdfRinc/Ora
eptN3+KQ2xks1friKdlyS6JuNmtrvsiNPYbd27onlLssSKdedvoUV1ucsp1/2t7YA7fyq61vZtY4
TU6DS5W4IeoOFDrsjXnIA5B/V/r/gpjLOj7GFWCcSnDpx392G6HZrx7vWC2RXcmnz3za68iOYvFs
OD5pPiUx0rpodU2mFG7K79cs4qd5cH6F0D3UObODTM/dK7D21aRvZAjsHDVEU6rQpklDkoHm3bDD
sVvmBMTQYTBufup9liK/4mqsTougDAZjIWCdUDyCrMGv/8YNLxF6OvEQxwzl3ICZd1TPqmIxk7xG
+O7AvCfsMGwsIO8UtK80aC7lYNmyOGe0BGGL8ikhVS/4aQrNTo6XgnpdoRA0Q+rU0kZ6x45wkIlQ
mD1MwI13MVPMGQx0qOuT2uB33UKrRN7MlY5dj4dZuU5XePyDZRCQxXr5mjKbglD+eUs+/cIGye+m
IG6V5mfAGkbAoI+ZxvQWABKAbesC/5uNU1OF5VOAZLJneY8+7aK/IrU6Nr6TtobqYhl2MOFbvIyD
ysNyix5bzcd3eitDgSGum8Fsc5gkLYOZaPhKirYmRG7Tgzffgasp5h4ZN1DYnKD2sW2Tuf48+97K
zGMaAjgtSecELGCGbZ3PEldOLWfARQeRdhpfmcXMKco8cFO/GWnoMziwqRra/+nP7Ue2aMYsvCtX
BPgXPi96MzTHXbpYs68mAVqdOhmnwjf8RuowZrHT0ArKp7d0edSzKNA8kejhf5WPwSNJDycYecJl
9zuHJLv21DQdEJ+uJgpHmuWlsi2uc3+qsTC/vcxDKl+qMUHNC1IlwK66E4dqdyLfDZv3Tz4VZFuW
8DGfHPYZL9gHTSNn3C5iufsqdLJUtF1PecvuISaeSw1jN5Qs54U6fJiIAAQI3bFjfvwDOSLvD2TU
1OHZnTxfKZzQ44jl1IFcIHC+kQ0BgfxA8qYZgVHbUsJ+ZHfsDf75Rp/21+1nD+H/lXpLCfgqpppW
ViFmmRf1lnZONizW6i12KwKrs158loy7qCXCJQYAvMgTM1bYLOI0QG8a7KFgOqaIf9vyClo36Pzz
jdyOhdtDZjCTa5s7Uc1JxudAhKed21hWjLgpOGGPXUil36ua7T6DdBmVdTIUM5rxnv5hO5m7DlKf
Hyup7RvTOHC+Ub5bynAGpOeL4b73LEAe7tOyawgCqeRcsbfDujpqA3OqHMBCRc3gHbJddUlkmHjq
wBYA5a5/eXDaHWLrDAcmATpKqzZxz8V5Vdmvl1YEe8JycvTvRY2Y9RLHSuv7kBkFhPxWou/Nh36S
b31DjZSNSaB5x6LNiRki4lph9Nj+ud9UY1y4yQWevQ4WjxHVdFKzcv1m/2fvwHLUbV67USHBjohR
H4gtbp32dzWjjPuTT+yqOi0NH/u2p6/HubQ/fFrS9PJ/aVH18+mptd5jDQMKDy2Fo6TGPOmXpj5L
9w3L61lmPgN/xRbWASLHsHd8ZGQ9UF42YRomnak5X+EqM9NLKKIfpl/bgh77XBtc+toGm/AYjaj+
K1zp+rXMJ87dwbQkkFOrss6u5YWigpzDB2zaIlLC5fvIQ2z05lephsbwldtTRSYL9K5imdKKCF5i
bNz82JWYBoSp8k0SJlSdxa5Ojh3eliCxoxsKZrbWuOae0gva9touyMGv8+2Bm22PfA/XsTLZg5s8
VTy/Bd27fMNEayG1WVXzLPT4qaQvkDU9i/Al/UjWrO6zG0p5E/tF8gw4TnuhEUi54QKxxK9AT/Br
JxiOZQ4585IRLjvxYGlBr7QMUVy2+YbqF7Gx+mA4QyQjcegVJv6VhKuA2gi3mUdT4s2VWmpHO7GB
1zQ2g/XzyIOKCIhMRmUPrTF5hWnhLt5dxQZhiNvAdKxprSk0CHOLhvFrnxhMSKml+bTR95oMagAU
g+wEG0zDlSDkwTwxqNwXHTPXl3RnzIqQpfQBAtcZudk4Yqm7ALOJcLUdNOjG+o7/0wt8XxHhdsQQ
9cT8JkQkVfCudAgDdJ6GYmk61/kuTPyQA1oTfKbr9yrY1OnjdB/DiRQoiYYMPBzzugiFlRqHoqL7
q3oiJ/5lgf7sK24W6UOm2wHfqaYxXqwoaeDuEjNgtlbqmkOFbnkljngOnlS/34isjmuLbsmG64A2
OIC3241Km25LDYOoISj3lhZV1JmjgfM2P7RIe6eyFKqoRTt4eRP51JQl2FOWZbv/lDuzM68Q0wW9
tfvitF32XaLvtr1g0FVekY34gnyKXbX9kfTydz+hSreYrlx4yxtCP0iHdMgJcp5S48aFrI03rnl7
LFMGez/jCBCtcRsZhlTCKMkqRL0QSoRQ16DOnwTTGp1suQrTmCSq/nl/4rp6ne3M9Mav5CJcRdMi
xR3+6OAaKUmGs866jcdC+Z5gOVvO37g40gwxb0kUf7R/m9ORwjFtvRaiEfrHXvIz8Vma+lRkZuIF
P0xfZZgRlTQE45Roi84d59rd/ljYz2br+M786UjjAy67seDz7SmqvpOU0nN7HfaWx4v/DaP1c0cy
jubc2Np51df0P8LSHnkspJVoqfYIIVVQUir+WwMd7TogsS5baiQCQ5gOrIdjIRTCqcEi6lxVmRHN
OPKOiozkd02GB7tjhT7BRZQB7+nI7qqcGwAqOcJ3vYirGNHAgetxjjZbmliva0QXTMr3V60KkB6Q
jewkzVaFjXzrH8fhtYjpP4uksB4IFUX62H9+Xd4aDEj1JJfaF3TXBlnxr3KJ0Su6JoShHRBpdP1N
QkL1GIliGVhQqD1zm9wtvQdavzkpzb3Y6eLgYPf1C5rE6xKFnecEeuCDsNPmSZtyxnD6aOgM9819
A8EaiKI5/oEteP8/ffs1YEQ9F/7c+f3WREXOOX3HX8Gv+p5uW1Cdg8VWZ/BKwGw79khjBldMMScO
kWwfj6vUi4QgcaKguC6VgdZOJqIahbOzTqc7YSRpvp6EEaiIgbFc8tD14BaBJBEgtW9CNte1j4S3
Z/zucLQVrviEiCo58sdd05wLrrVeSAebEVA0kapP+XBu224qYUHtn93L4xSPc2rLOa6QX2dVRU+9
ZiDVHNVHIwoJ1ewm425V6caVvFhYkab8kJJCI1uLll8SSqEEE4kSiHA1CMCGk3A0HfrEbKSa/e7+
3XIG0r5k1huwOdQmlJevnVe9xAQDKJj8Z169LPsk9BUBJPNGJGAgOo92Cu+zZmXnx484u6+z8IND
UvICfgqiaIDoYVnI/MFW0vTmmWLk/ZpNQRPObonGcQ9hWokS4k/x9EeDoeWHQRD9AVEONIrtc0XB
3BFJPrNl/7oKpAoeWKj15IBnkNJIsKYpy0b89JVaeRmJskqjc4/4UX6mYthgLCOAWoWY1KxrnNKF
aSTFliIOIF0oJh/E3kJqGmBcqCGfkCZdtBE1eYMlZcjWupR2Kw5/TbpP3utRHpmqrG3L6ws5IYMk
js++cBj1CaQEElizADdBvkjwJjGaLtUZF/uMojHYvt1zF58qTAmoLcoJr1hvtDJ0GWcFmR2a+RhW
WI4XLSE7/rlYk1kZ08UxIzUh7nwC5Ke6ZjeZ7CB18z7XwAbhNrzwvm1wU6t8YVln7x29BmVDjpmZ
MUIjq9cnA8fwse5svCddxIARdcrG3hmd93HTEb0oRNLT6PjWbvze3JhS3wCSUwA40NS4wv+qzvtH
YlFE1jTFXjQnWB0ZWSnWz4HNnW2uN9TSzkz/267nROZPIey28nymN1/qdlyL7Tu0J6LFI95LvYB8
6xBtcNPz657elXyhcqSkMBFD4W/sZ1jXMOlL4xq4MwPl0mqkMlrBptI0PE2rfdBom3zngK5e1qFB
IyhqdLIaOGVc5sEecM02yLwvW6N4YPqUlNNHfl3vyTlRlX1etMzETMJE4RhnQOkdc6+xKvm+3Gcx
/yJ0iaL8tUuPrCpim7TPPWMqSqQJCbk/lkjRQbFID5XThMBe2TqbGy3Q1833Y5Jor3YzoOifPF6D
rnMbUsRiV2mK6M7daaD92uhOaexTYk7A0L/U8S85dNr6Ap8/vPjqPoPBuSHDcaYjVeereEkW77gw
4Y1l6F4tt0XelcnQloNzrO4SrsOtHbib5rYvHny+AhIdSvG629SdrtY67s37Z4LBwRH5Uv+fpCRg
BEkUZsXfsu/wXFkvZoc7bgrvxINCeUvCevzxCSlq1qbkzLPQGU/wAN39DnSfu76QeaEBiWqRynnA
PWAD5qeloEu/AyNOb5AGFk4+SHkJ710ulV+Ott8hlkPMdp+Au2+vhPVDXEc5wvd+hxeZUvTEBTbe
O4fSN2iSeBDJHVpvM4mBxVcKCY9eoowPmu8o08lXi0QmF/9WcpHO+yXuHFX9GMVYRasARm/cmDXp
DOoxxTuNLsVNy4WgTaNUhWNZI1NRha0I7qsLeo+1YWv+4o/kyIf4Eh1RwdfDmMVBZUfoJqx2wrMq
M6vBRqDbKI5EKOBltTu/oddlJIutbg5RZE+Pqb4u+YMlBcss540xshUMpv7aY5mW7suNLtgnNG7m
DboBqTuWa00xoGLhy5UBjq/SJcklwpr2DHCH+4tzworNQuwsvHcJMqE0zGNPHJ78cCkpoGy9Zw6o
9jVAH19l2Y4CVtaaJRM2xnD323ikOZQdVwHajF41lMj/tpB25AnMXKuIwvF7NyUaJBbrLD5F90W3
l4Ga/RYNfzLg/5/Vew+j/V4+X2H9GSXBB9kSgxtRFGIUwM1diMdhtVxi6dqp0StBJ18RNCUmdBLq
mFqo7VLLnq8tIHSty8Ek7avQcGkiK8zZ1NkIi9okPt4H9Epu7ZJPWBRjBrdKDAwam8vn4mIWxOoH
d8u//xB3WAzOYeydyZhZghykrY65K4tSM9zPtHmDE+kRgqpIG89rNLEAWfAkMRHsCyHmHANZLglB
zuEkLIgJBfH9RAMjEunbA94hgLOqo7Udzq9zBl15IOHS6oqoEH+B6EADQN3w41ouH/HWJpBIE4+w
q5nM52+uDMlMUW/n7E7Kkrr57hcgZvqIQ0MaL3JN98cOKrC8Dga3KmFu0PvC56Nv00byF78+fq7f
nfuWSi4BwFtxpBm9TIkrBZfTHkG1D3YBE0pFWXEHmtnxs6Lgal9WxpxCeTeTP+jxRpdWodOPvWOh
uD6FmuzGFuoRBGuWv/Oz3yUZ9S8pvZfP6pKrSYX1mThmdMDitv7rSoEZRRDgQjvNkluG3g2OpVLF
HzNKJOhvk0sU2rqF7tOHd2+E/WU8zBUmgO4a0ceq1I7hUdP8Y7ryzwrgJKHg4ETlcjh33/OPY3qN
pWEci5R6cGYQwwcbJGZ9AyumM7bgmUl/+suPH4tmXN3SZUipCeZWrUJG6kT2HCXvV7FQAqn7gJCK
E7Z2I0l6qzW1t8b7wflqvwOJsnaPenm1Prvtv/kPsCx3Cuo1pkAnsdiD03Pt7pLJfvzyjEgyNczU
RwVLavFoLEFoPIGsdZAbVJL2u0sm/CBsfIgZJqPYwDsDl28S8wiOLZlHtE6N0mzQ1qSeUCzV7Rj8
ZJEryYh1qR0IWg/u9MKGgTE4RqQPZpiL85SZJeBC6RQ9bKa6/lPYrOVSxQrAyzqQRKq5dI8qQ4gb
Mbyqy+U2WSEZQ7uXwZYJjvuAi6Ydx5ZWVQcFpLGGg77BXXHO7oVeClufru6bJ0beWtLC03MyzIyt
badAmW+8O4bAH6IYZX6mjkL+kc/0xwyUO6dpniz952V2QpLQvkPTdJ07ij36fHjBxibXos7q+L86
I92oeSoHeSgspWsowrY+uQ5iwK1I/yTNXwNQU/QlcpsifJwLNaaixoHnHAMQwpE2r/yOt5chHUSl
ho5WV9EANQzZW36hFZVwz1ucKiq5IGIXj/BH7aKlVKQUvYDC7ycDEOG+WQmtFBb3OsuU4FZWFpL3
z7aHPOraaZp6f9/R5Hlh5wGrJNjGGnWIs2wtMGO3LDCJn3bSPC3+yUYWsODqcDy5ELOiLP3/1yGq
YgAFoUEDZUCfzE3iB38ZNxYV7/qDWbx24zXhhze/Gz5PXrs5OG98nbAYqwkUVjXMJiJbvMyL4kg0
VdjqyEhHGVu5E1oomDFo3xDBiBrJprkKqhcEty2Xk4hupLIqAH4JrIc1seOFkRXX/WyYyYLs7wHP
zN9RrOFkOPMw4rdkksP/qvQL6Gr+7EeZdI4cioW0a8DrRtFWrZOXyu3fjMMYvojYlZjzpwoUTT9k
sUjxwQxUVbDg1vGBk1laYh3PESSvxHU6yr+XuUMf7PgN1NBg/h5yQYgJm2PNFupsqgmMPxow9mHz
3R/+0C8y2HE687laDTO84+AQrQ6CnB1SSMqsUgoH7GvJFMmVjiqgy2W6Q3z/950kg+w/r/aQxQLs
d2I9k2yeEcaYBBP+9G4qOuYa7MVFZxc6/KY76O/jJy+T4NTZz+CA0h+NCFhvFKhGzJkB/QN4UMri
4m6eIBb8l3w9h7Vsflj6LnMA3n8l1KkwfjYSPnLrrdhnOUXYIbcdYf1FoZQDYSykRlxFv+2YssQn
S4kOJUr+Kzh/vdHRFYRypox/oy/EyD2AhF9g9BgnNnO/6mCxsaSDYcc6C+txgkXEIRaq9bpk884f
ml7l1rdfzmxPpeqRC1G1LjDAD08jgwvSxh51qXpLmYr8uMn85m91FvJxJOJKSgy/7B4NqOrHAnTD
G/pZIa8i2PhMiPN42T4syVC5IeH4hs7lay3DvXSe1u3W71e2iBHPnAEfFAf/JSMFuNUO/P1v7dQk
Bb+R57zfi2VQdVEqanSN41qth16MGpWdT5WW3k6PqgElFhmMOSt1GD54jcipGXWrnWrbhm6kFaWA
fFKeS7SbNMJPt+KAWmkUp18BtNefAi4TmitpEQycrIrAVjm4C+CpJAlFtFnT1f0AbSY21FWPI8R1
SW5s+ts4iUxrxL3uhegkA25JWcFk43/LdEiYbNY4XSoAje/37kX1l/7q7qP2mRz69GzhlN5LLLHa
jimAt9wcconzbIt/RDIpYn29wSovjceua7gq+EYRY4rqcW6BnRc/ABqALmPEv3u78TvuMEA7i6Mj
lokRLrvOPrnSZ+Vl3wZDmBoKwHd/V/DmUZ284FeN653JKAFQAAbSt9kSVyjqMmLP1BwhSygCXOAH
8geVrdXgA2vi2EztPrNwyiYKh8xN+1kgSxXN08F8wwSfNpbwZJclq7brZsBwaciato5kdomtK0k5
2T9HyQZngoxLIez4jegYiNLwaGjgS47OUhcu1YH0RpKLax4xuMMg62vlnfzIOzMpimcq+eeEM2wE
e+weyMNDA/dVBzwbbStjC4uSUeMHBS1mH+q+i14PeZ7bw4bIeAyK1+kp9K3w6XDomFvBnBsgVdGa
HOYuR2EpDsE2qvsdc7T+seBhpu87snvzuuvcNSk/d+vs+DvLWX/dMYgaSnqghmEHrPvi6x+nsXb3
pj3A2uXISw8H6TTwGgZT8/lkd6nnYZzmVIgzyrCHIGSWMFUBPFabAHZntnWndWhLUWpKIJj2Upnm
wvohiSWAB5SWCG8DSti11grXuA8ZrbzIiAgVMNqsTyB31IqItjzRGxe5wZqqDCuxI+s/RDooWYve
lbdIQovBmVLSimOFHcIgwll2fVe9dl4F/UiGV43y+n08yLjPemCktGdM9Wsm1uKkdxmBTM2bCmRT
PuCHVPitu9CmQlamzJguhTDXsTe+cFXTC0icvGXoYusO5LSJF8oIXbXttmyY4Jb0qO+zTeqV5us1
CYaHQ5tyZBaPMmJNP1/OseI17HxVsnQaD1+alHdrzjcAxLjftq93bJHeMnWIbJhSA2H9WXUNBBlL
f+pvi8BhsdytuiE/NkoIdoGqgMswdfGd43/I1MQ5KmkcWwoHgreKep8sNu22rQxxsMJZUnJrps1N
OAnrt/Dc2DmCZWTYzsjN6/h0LZJEQrMtt1cNS7n4jbV22jEy0UFv4AFpy+3rs3Q7n78puTxEgVCo
bMK96P/Ki+WFp9papIYnUesMd0bORZfqkEC/1BULYR4kFwbg4LAc0rRUZYXtw8hHs8lQDfKVIkpQ
LFbulEfGZdi0n6kBIJSLQk/ESJ4ON9XmXBa90zpuu0NAm6JL+fz6oVNI4gOE70+bhusQe0z1haQD
m8QAqYAaIsGRqck8t56Sd1wf/eSHUyoJr6g6pZrzCxH6GTLIap+YHpXeWWBzK7FfAtnVY/sXhR+W
XFojeAkKnSNGEm0sNBc6+IJfeJFJSVhtRDJMhqWv25osOBlhP+49uTmxmiVaFbEUzwnzbLGjCjRz
IaIDd7067CTuixA32H8x2GaPuXINE0BfQt9TCjh/fBfpNoYFU3mM7pMS1WFlOYyKUnATsuefpvgx
sdIBQNp2pUWlRc12AKEDU95LiscO0498WdYSmn6HXeiETSat9kQHncYQVrTgfSbvBWfpPPLzXxrv
yW0kpV5qdJ3sXMJ3fJlvG3e2oawztSlM4ijOPzZS609PGr8HGiyt2nq28q2WNU1i1bF1YgYsJ/ml
XYNErG0ffQB19nkLiiwkZ+spMvJxrdbEWmAFgkyWbB/AJKErQq6UQn47Zzo+dSSH8TYFph6CeuJl
KPrU2+BS33KE5pYI/d2DBSf4kDEonn0fIXjbjjY/PAk6XstzH0QqexoK3ZSsBXG3T4Ndpnw0Zcr4
wWGPr/849JchjdERDUu1Pki1TJhGo3+9DaKfQS/F+/ovQ/xbhgESIxCrF1z3QXh9ZdFnD+Y0YwHP
5EedpL/dibAM2TyfeBx21qNCtsmyJiDzn3+MWFL2HZRqts13/yvmSm4Qu7AilSQrahMmh3NswBkT
2fDH9MItCDkpOYkiF8CL1K8CeilBvxixkygkhTROzSYjzwa62mhfHvgLs5n7yXQ+x7TRv81esNj+
xDb11M4hrIBUZnx+dLVuYMgBmP0+WL5dHqfBofLd+bzVZfMVjeDPxHlMIBQLm8fPTxf4qStZggoV
PMMfhT1gUFjcjDfRCPFP2mWIr6eKkrjePs6AxaKLE1rSxdNqY0GqbHUUqQKk5tuplUI9RE6M7aQW
Mc6ogzAKjSUu1I9hFD7hbWCOsLI1iLbhlu1eSDoLum0pwvIvZ3Js67A2RB9/fRBN6bEAc0Pja2ra
Kwm/gi9kRWDCzDuT2i74SYRHLOdddUEU+GXUtmKBjNv3ATveo8dZbXLNpR8+6b2V/yyi9mzYQCgx
D5AEhBqRE9AsTv3dorRMvZsxCSltZVtoBGWsqNV0w84ql+LInVoWUp3kbgejGGXYXF5QER7CdPC5
OL4YGX5ww130xtukfd0auNhxqSwbiwvwKIdsSXlgoDN+bR17OBctptpp3t5liSzBfJZjxLsBsr/M
jxdoyKhb/B7IXkdKNy/JauCLDCE2NWDu3xJWqpiAaWttL1p0+i5jyTuCecj5wNvygCiQ1CABc+qi
qM9HPSdXkRnEfRyzLvb/dj17t6Qp0vkf2yD6qp84BquGK38BbSOxHJtDjGVMc84wF03dY+PzD90F
SoyMalpl1z7YfSIYD3ktDKkzWvh9bCSbQ1+CEDIOM8hIlbxZ94XFkuOhTISHBjokKmDlbR/12z2r
JM4gr56CrTW3NfT6vf+fKehnVtJ+DyRS3qKbXlmvLiJOFCanEZZ3e6lDRWS/exAhF1Vcb43hMroe
Hw41v5R6o8epmibQR51FI5OaeZcHoLIqMWWLBYs2c489zzCNyRO7lUKmYUADCWyKGbceR/EjItU+
QZjlQKwuPUhxaE8hLzKuQa48pFOPwxxqJnb/B2rIlRYUxMj65Orld+/itTBf6w2Oc2fHjVnOmoUg
wr8ntoJGnPoRmxp18dMCRcwqZrsUIFRVeT6hVbDpXyBNLg90mGu13CzYYTpuYFXCY7dJSjl094wN
W7ODSZkyTEvGIZyiFvxki15R6kLqJ7FISTdMCKI7Qt2mrbcQlEW3hQmFfClurTfiD4QfpAzPY4V2
NezuZv3IS6gOgRjb88bvYXR/ctXmacEZrWsEbt65ZX+r72vohpz5tGaZ9tQEuADBcLUMKXqBW1F/
zgm3iUVnPgGOmUJOiKQH0W1vXBmAbcoqZLqOmHqN1nlyM36kDo47z/Ufv+DCmIvO9e3S7k+BTcys
TxlVaSDks7z2V2dSTR54b6CJzXAq0XjHp4khRDFEP+d6NtwYTPWfsfBLSzO5hNbtSdagujKoAbrX
eoPdaEds6lukAdePsNWGf4+NNnfCHMPesWdfhcUQBtpkuxsQrRBxAaCq+O2xz9zz3vF3vT0THjBU
sI5vy1XOzIbIwF8XwuMunAs+ZzRfy3Zd1OFUkXUphIrciTRIAVtPc593HIFovFVa5WtUetQooG6C
0RNnyoaYCMhcknd1K5O31sPUlD50BtmQOZEgur4p9klOz4qXc2aokdMmpjR2gfKaS98EFBFlPTjg
Q5mLdldShlU4FvSXMfSE0klHH9ttt5Y2KBhPxjreHMlwYwePQV+G9NlNT7S9KHd9XJsthZv9J9ty
f3jUgU3OZu2VVFBBRs8JYFqekphg8yaMa+cbKInZqh4arcfecsYLPSWvQj/qxFEqhRP0ofBO2LN4
1BYeyQg94h/qc4+YkACENLrYHvASB52dtVJ3Hj7xIwVJvJZTjh4b9mPhLodPZOBnaDxwM1MrY8RW
NXQaln8+y+s4WXXCpm8rEjXUrepiEyNOUnyQgvllWILjms0T4oJjes8P0gPeQQ0uJx+hAf3THtW0
Z+bxKjQKm3rDYAB4asfjuqzoQ13ul4R0S7wj4LfFcHY2W37LfAxyBJB1q6yAfdVygBYpcZ3ByTNR
nT5xux66+IJ/q9vrOaMjrmyUIcPllftBu2xlEgJ9oFEzdiib7ckuSDehRtY5L4noftOpMdMM8lUH
W++G0DjMqzA8ZFT48qtbwD2RU/oOyPbPY6f6c+vrYocbKZSQgxTWJWSHzOxrtcQ58f6Br2H9GVkb
ENwQXBlGIlMjoH7UcczfYQVR+2Hqb181vERUk0xhPE41jZzJmMxcHfIWBEf3kV9QhMw6AIFWkCD4
9etrTqlE7qTTB+9yAS8wokoKTwGcQ74zZchWVg43QHqwWwP3/uP4RXq/D4LB6ojp5yzvI0t0pfjQ
mOrS5x/hp9U6xVJHkaCI3OZBg6wnw63eCH//EElkK6vxEQb1+wCZvaXnP8SJj1um0TTHBdigpPmU
9WPUuQGzGP4rBoD8jw9d3tQ4Myn2dYAQJqUxMvkuCqegLsFppNX7IjYD89TK8I8/LBrCAXV4jogA
B70rGIfZfrAW9qERnIrZ2ckMHQIBi3GVDOBUn4wt1GhHU0kGqMYMVj8YDWKsJDZ/mmt1UbUuiO9h
iwQc0WYQLviIDK0gwcWsCpFEYuI5u65MGaQEj/ENGODSO9OXwZPmVLvZPYi98BST2+mD66+0SDQh
1gWL4lGkxN56vW1CyasDnb8XnIVqVa/41vIq8+ROW7nNIpZVpZ6auZ5aNOJkt9WYeN0tESozMVH+
bCVqtjmZVLLpjYB8z8JFCQyk5uglVdTcTeD3z3k/xUcZKlQ9ejD/RsmgDMmIWP9qZCM9HgYefBI1
/o/7vyqC9ycSbAiCRzRZNvFfHovzshwSFjMhf5XtD7tjWLRWRjlbUEocJftTiylQcrYNQU0LM9Ru
7EtxKoMbtX1XHfOQ/2s/LW038RFDr5RXzrd/F/k+jcmRmO9vc/7y7dOxLy0V0zZAdAn8yfyggJ6Q
/HIkBZrhQND1Ubw49O6GJWOjeJcNjgVwqBeOVH0zbLJQowj9mfFvr208Ls2+T3ui4+C3dUtLE1mr
wAdr3RTO35DWhX5auIPzztrovnfyJ423jg1z+B0wzfR3ppeKsz4KIom0ZSjJZ5KOFCZDIctwIZCh
Ln+0OmzQaEx/kDhYkhwCHpPtXs1c59+XD8wSJpzLfpKiaANDR7dCAjKEv+/UbmgRAgNtMH/5OgoD
2uHn+BXFMjZT9z8ThRbSBO4RFAEFLNXkUbeKcojMaUBHYAmQzd23ZqR7tmtsZUznYQeFTG4ZOcee
d/b0/22NlIoMmEtggJNug4veq6dmQWpEPad4NNf5JUZU13I/8VLp7LigTXqvvca9C14tqRFv/SEc
IC3RH27vYczIP1r2eY44QFjok+7AsAYOGwyqob+nvarPlkvIfBu7uf5kBt0+xfzLEt2BJ9fUrZ5B
7S10ZSctlp4AGDFDn0IbIuKNSBJU5iEQ0+YHW6TggLK26UkO4Q7xqZs4gWeHNDZ3JBDVIL6rRZuk
n709LxFi6pebCH70G/et6PC1YJorA7RqztaCqmtMcaIhr3R2wU20EhBqMupaIAmZ5SRdnfGMR63W
x50tZK7AB1LHsQ2rAIPwz9hUenaooqJ3QW2/UAvCqJqVtsF+zUMYbbbNIYU7oRiILvu72kj4U1Vv
utIR5OjvU9LuUTsFxjLKQ3U05KMCjU9M+J80YBbtNv9A5H1Twqy4KJapiTfR4PKPMeABjXZIBdJ5
YKhBPf0xgyhwc8FRW+ll045CKY0uk7Bsjae3rCcyTiPwB2ZZuTZDttMCGVBbVLeMwt6mLfLZEhz2
HuvWzXy1FPdp3YdoN8OMpzcqHDayku6MOdjGi7naHnv/lvgWnMNTzv+i0xK6eAPXmvArAaTsV1uZ
+liwIdLqK0/e5gPpQRzluoaHyXy0/khGjz9S1pmi3y/owvHFzU/62/5pbXsHAP2ts4lv4H0gkF2M
VNC2gioxXCBKiGCoC2uvJBMphuMMdokebqXtGMT2eulc/rj/Ut3qYwTPC9KRsPWHvyjYAD39ada0
GFBy1/PiB8DGWJ0BB02QyFqNxky82e8v4G/L/yrn9KboUG7K/DKuVvUKOx6aq+hsjNfcaFxvkOal
S264TGo+Z7cfr1dXc0FIEQbEsNyJfHIEVJTpPy8m/93KAN/xdjrAj+AXkM216+cr1fyU/1txBZ+r
Ga86i2EEP+exI/4oHF5WNjJyR7ZyzTzI29Jz4/YCNjwsfrVYsTJak/vWYscP6XigvGNZkmvQDRUJ
3O5yPeTtrk6B7G+xavCWxqw5+qwusXPivSAY8pId4UFJVy1y0sYECL7CyYK6WqDgfi19Z11JsJE1
xKv8ivo4tfDKx+fN6d74Nk7Kq2GTMR3qy9Qg2xoPsma4uug3qcPNUefdho6pHy+n4shNqyETsbVh
i2XxWFy2ZoJ/aAKoLord8HNWk98d6aKCm65C3ESOYHkfhD7QDTl01b8NPCCrkOoZYIb/VlQdSklq
wt+tMpgx5Icxr8B9AZOZfCFN3BgXQsOPQXL+BGe7IsVNPOtHij22Jw5i4WfdZ4ej9o3M//Eax1z0
F27z/+8g8Dfoh1PkZI3ZSdVTby0jCfMeHHrdnbZMfD9Llod/qlAa27Zq/UCGjl6ZBiio1yOOREMm
ZZiuUZ/FRIR7RL7mILyQHzQ+r30OU4Yt/AUY5Feg7aYwhQ2kxE6zc3Btg/FrL3bSJIMCf8KaKyw6
6vt36YRYdQSpfNyQm8EERIFww6YrYRsMr8lHcgVViCRVwixNDAVl2rgy69T1439Lr2GFYFBv7ROx
CSSvk86Gg3YWLflJLDiKs/nLEI3oUdRXXm+Zjv4ZaNoV6Urg1Q6d+G5GODX7V/l3L/NnqHr6L03p
Fb9qJTCGEGtb4NIwXKDpHxKg1c70/MJ0A0dm511vJat/gnA01g5abGFkT9VMchQiYjZHwYpwQsQ/
1LjqMAph6SSejYXhiIhHGtnSl/HbAmGABcHH43g9HvWXmMseLo77ZfKVlNdtA5nMxL4eIvxZb6AG
D1BVZdNHoYwRUr6v6fLRA5skggPyh8MVnKlYm1GjyczFVYKK5Pi0ZiIpLr3258TLNl2yzqBez5CT
MBehpKFvz96fOVMy+3zBMqW0ulMPU8/odjzgCMQn6IGKLqWm6PQB/odEXtfFJ4D6P31jzAeQLhnB
6MmirOEz/g0Iu5bt0SIRI2yg4Pgt8gGUzTqSXyE1WRu/Dw+GMb6WTnxYOFwWgbAy/jnS3BMi4hVi
kD5Jo+YDjb2IZnCLbsPEjLwr5mALTJBMrPqDnxGRsg/zJzP9zW4TCnsUkA5u2NhDcTzeczWkPvok
b5DNBuvzCGMkohMEpfah73qrLmqr5B+06qtKGuXn1iQCrUJ4t9kHoAVTMKqpISGGvwA4QgQaPYbv
R4Wqeh5XdyJmiCAzSUb5EvwjNrIu0Uye4CZVT+PPiPgrzTgyO7Z8tD4+NuB/GWiSY1Ji5MclhbZW
Yu5fKYpB5SKjS0L4fPMBDhiNOTPR60ociG6NSEOxQEYI5I+RrYObnT1hEW1d9cpUedaxxsr9OnGE
A7wG4N8LFxamArnEtirQbDgHm5ZyF/DqlQsxwPvm5jF4JGBpDVM1oZTs8I1JU4JsVQf+UOYJfbCA
Age9ef0lobn7oTvzPbvqkCtKXTyq6SgxzgyQb1jRxsMzgU1niwWvaTqrUV3ZGwFhTgG2WqEiDMXW
EeIfmx4u9dEFGgVgug7MIHaoosy6ehgOAeudVEQijie6QkbHq58Q4JuSa8ZXbHI0FCwgHrFqa/Gt
T51E/wZ8HBFDzge/2XH8U0pElAmyD0MrZk+6j/zZld9NjuckdogQEWy91NdgY12SzgxX8hqeYikp
ibLxCbad7YFmm1eKriC0ORxhzP0p2PfcJ+vDcXs5jp/m4bltwLcPOy0sHjhnfBG/5c9tOR2IbyKt
37cvRVihinoPvavi3unWNYuTelngyKpNQrgQSj26nleOtL9sK+ft700GJemLhF1MryFiBn5D15Bg
r8lFM08pP+tSAVwBNI3/e608gHsX4l6Xt76ixSklcKzxLM47ULy36lpYpgRrae26fJPj/Ylil2u0
2pr8ibRWqu8ohMnqsMT+1WAqclYUj0IlYTbyG4Kt7Z+lc7ez5g7io4Md1EHBVrYcq7kVjLtn/brC
EnWqlp06UZZ07uVUJmXDqx7xMoerNGXK4eKPAoQ/8kP+Hqy7jB8easrndUtJdCdKIIjePEy8uqTM
EsPrszuw3tli+2p79kuzsjd2nXTKh1lbKDaC9O8X+RDS+XGArI6tusU0EdOz0MMn3AYcWKdEHUui
787vvU8vtL2KEJTz/JEmGRK7ARZhW6WiagMDZoNbRU5QXK7UCVcjIFc9ZU4OyrFxTEW4sbZXncpn
3a2quNwtio01ZZZLjLBh9xg/o6Zw0SjUOv02pMCRIsd6U1XVBsu5NIeIxPMZfkJk7/Y5D1o1qR9h
6kCVs9ZF3YfYcxk6Nhq8VlFzp63EdTqCrluOBJpLKA07KeO+naRUj7mR/tKNtbOTC93Zh1UcoXYp
m+gqSCXfm8Y2syA+hp9j3qKtIIkfS0AuEAN5JmbwazpkeQEXdTuweUHaI8lx0uXzK+g9q3X5lWrk
uLjE8w7/nFtjAyf7L6Zrlgbm85PeQ3/9eK6NQZ29q9QEdvI5pR1iXCIwHyZN6wNJSeD7pC9Cla6+
MkKGIBDv8SAm9HI0lm6KeXLxGp5xaX2wcpFUcCM4igsQZLOSrZYJ4NzKz2PwtjRwKmILZlyAt6a8
RZY6A8aP0GSoU+yz5MCams457D7KU//gfHQvMzsPXHuQMD5t96QyMYTangWYJ4COKk8u6gq5J9pD
lzpm72B4qsuenTW40HpLSeY+LhlwOerKijgnqhpvQ0uJfndgkqDhxP7Gc9r/o3MyXbmdlKj3msmH
jkC8Teh+T2A/SdPM3+ncNf1hC3NcjqR53wZu+tTaszJQPafKQlb8UoltmlZ4GhzPi31jxnpdnSbl
XQgErRLZoxmsylEm/9sRCh3dXhV6kIXbrgm97uWL9b0iV8fGg/j03NTvl3oQFCVa4UpRVcCvn36Q
coSb58bqfO//z3JxE6MhcL58fb4GmawW/Og1/EeEASqV+Y8zhKh2e0EWdFF9hO3f9gwnKn77H2ds
CHgwsthqYCjPB0BioWC9G1k7HRjFWlf9tMYcY/9L6QR/knKDU+EZCMmrG6ZftPEYm+XEOzDEPgf9
3Mq0IHuPIGQmlYoJXuwzmfanbiNoHupkkiHVw1tC1rT60SRcjwF4bB7WixbgAR0Nv5Pq7wOJngfc
Ppk221Em4MP9QQG/U2IkyIMJjFlN5p9OjEmZgMyTm1JXtNt2clb7V1luTEVVtRa6ImFCU3jhow4E
feCGaK1OHJGjILOYVO7uPYBzCk3js0QlwdCkvFyf0M/HwnZLMgP9gBMwhrYxlLhpZU/u23adSDHj
MWCtC5KL9sa/qbewRWlJLUMmehq0M5kWnd+tP8EHe5Yhh5g7q9Oduq+w/rKG5ALPM7l+r0ssOTGN
ugYADFlBs91CHwZPuvD6tiNAiMN0uBTrbWUS6RrEC+JrNBIuDwxVcYsKdXJD7FRGdOPknfml/KW+
ic4A5sKJrW98tHRccP58UWXXbqTHP+rZ6eSM0QQlnO/48Krpg4f++l+yd4S6yoGSDf+d90keqMRv
AWPWbwnn+qZIXfZEi10bZvoS6UZIkNGfaRRIAxAoWzfw2SvncafpmneBL11TE1nx8+pkyslgEgKF
MqzjLGgCzo5SvjGfmE7EppWWlQSAi5O951jAUwQmjtr7G/zOhXKxo5Hll2Dawb9kPMcnVyG06LPQ
ydf7bX5fKmWcN2fUEOihLtQMPtWKIygaAaVRSRP9yDiPEVCpwpLQ07hcqADJRCDbE92Fe7+OF6CR
Ik5EFyBqjwaEYU+1dgwSV1jXt7Z4TqVJKmzUgwazcPFTZ6DsTFitwXLcCwzguxhoOM31i2PmcRWz
hazo6mBl/cCZYrT+zasp/Z9JDhHZQxb9twVlDilXdsydX4hT4LuQoVA0g3nG7fbcZCUffTs4kXga
lQewO57xOAnSXAsFMGM57VvmgE9En6vIJtFGfyUpcw2sxlSBY+xq5kgVpjfPqOjU7687F1aMvDvc
ZkfVYrrI/qZPqV77n0Zj0ERV/aSvOwRlL+dlhFY+P2BeqFGFg7DaQaHQBAmj0eQmGS8NE1ZljttP
ercZJQJxBnmLPuNI9McjtOb0k3ZbShqqTw48bSwyX348TWZ0jFxqEViTwNj8dfhnbNOlnCtiCYq8
JFMvYQ0zgdVoskTCwBlBXxNm0cjW65nwZ4pnEhOKhACqMezpdP6Fvo1xLB03UUvgHAZ6u2+o/zCo
w6ADsr84j96Oheaas47xo8H/VwmrXFlz8lSOjczOrn9ZG1iz5rbfpRNekpNsvBeuI4jfkZvr468Q
PoSu7ZXJbAlL8J946EJ0QutSbqNBSpni/9YhDBxb4jZrHK/5BWBl39BxPxgzQBiO+R6TpP+x/xsE
bZOwNOzSVWK/iCIps2lax4rkAfO20/pyLhSPX6qO093sEl9sMs75HbLV47wRTZ7p6iFUNigKtsQy
43XNcevI7UMSXT7+bLdsvcM0eGxZVhB0iuVR0sfDegF5yj27V4BTeXHbKo9G2nh1L/Zn6MhpCG30
y6RaXcnaJGFisFALAp3Ax+Y16CF1kgHotb90q2p10mfMspYMkTxLq55d0BNK2PCvVx1oqaOPHX5o
QRQUI9SU61zZd0pRtPAGTcjYDzfeBg0Kdh60DF5eohj0dizpU96z6a8MSmrxLagNFr9jp69QHEvZ
wMeakStz74IEdyLR6WOMYxE076CgR2rfFfmor3/D18uMkU5CYc6bnvwpOTbPGUJAv9TU57wBc/FQ
VQhgkdqqNvQYxQ1EnniFkTYtgO9eJaHY8CVB3Xi1//IUGYXM2GUyIEe38U+JQWW2z5jp3/jr/KIX
4zQNRntcXffOQprmuA7maZIVgcSOQSXINXK70TY8+YAqS/ikepyxikv0aI4a+iOcd8c5tZFZSYoM
MFNiYgUxlktXyTzlgKLOHcTkEzVNKL0UgUczrL+fy+zhxBt7tn3GuvB4YIfyTmb4IGrzQP0JPEz3
uBiZy5iRtWj/h5/awqvUtNLCK6t0pZOGn4/3sZ1mxVUdGSPT4Ln1YJQ0fyfNV5Ovz8F3hKQMVKi7
P88fNNl/LIWH/sOqXPifLTRl7siWNRDWXkXUr86CyNTf8YkXXIEsCTFscobVqWBxNrzlPPiF7k5x
qbKRVKMMOcc46NXfkk3TVlV7FwxNiX7lSr8Ii0H3pqoCTFzy6Dknk1NcloMBemR76KgEWHEmIGa7
3z34wQ0G+2PBY8FH65ZJdmIeeBsH1T06GcxU47ViNEWCYgSJANIFHS16gjNMMQrRIBYZN+m22OmO
aOgpp7gJFTw2tPcF2DxukQzhwUAEVoXesNVRWWzK/tTkzlZZip4ozotwtkG5rjxyMnZU52oVe/lm
HNu2YLv3JJ25dBIIzA/YYrD2ASEx+jxTOlONIN86IDmBrOH5YT3FFJml15CGhthTYuEeyBGcZWuZ
yGV8nF1r3miD7RD3hIWVulCaHoNiWQ/DN4+JoWRB4+b/nbyM4zOcrxN9xN/OVd6uUh0+7f84y+It
D/vH0X/Jzq6XPx76NIIBFFAkBVFeQ3w54IBaVqS6E57VUV+4/NzwXc3kRvTu5hBpB16HB/Yx2Cfn
A6Zo+vCTH/Ea74r3tBmKkaSuBLA7ku1Nrd+PJQwFDbQAd1P4+rBUtOwXJc7i1mnp5VsYD4Pm7B/b
ucYFa7lzeBCLY2u4WC7JsXaStJv2lj2mlik3ZEyaMq2Z6u6cbkU2U7BCjPLP5paA7iILPPZQncuC
Y5XqnlNoDyo7uWgcdSjTKxQqn/jDvK5uh9r+9BTJWC2BAYAxU/ubY7J2oqpOLreYZVnzkKyKFi5t
GNnh+FVYHGnYsvxT2/agQ/BR3ZdJJrBLBCbYAGs5DgSesiZ2WTPybFiaKwOpnUppH2mXLbU7eQYo
qNE/OUteNO7+VoaPlPSdsIurWd4oN4xiCzhGJ0WTj3rvznJcSONVLIX8mxhanLZ64C0TWAw3vlvD
Zke3QTGOoi3wnYorgrQxEA198QShZTnFeg8GWTg5luuy945zJsoTdCncFnu3FtKbz9EpU9vcJmyS
X3Dk/d4Ve9ZxXgQe5vfUMdGNKI9p8t5kTVoFo+9LH6fsUtXJBs8n0h1nFBm0VxvHNY3KnfkCEkx8
HLngvwnbaWZ0NLooEsMVkbP9C+s5mKXQYtI4aIsqCH8gNZA/4VHIwI65UX02wMlGgP67Bezg4kPB
adu6YwSiHfimasWCaz3y+VBXdI4dWdTejKjJS8JjFMs6qiw+fEEOrfvKHy90Bm5GCVvsFb3XX4r0
TGpfFlkK54OumkKwYBsyI8rkHIoaHVDgEEAbZyNi5ufO93qrhKN653qiM2BCh7gWXV2BN1OFfEfD
X1PQRitB4LXxOiiyX0rvDYjyHkGlBWgGPfTYvuR3ML8tTGvfH41CgCe+oAQqx32s5jW/g9jEhclo
2NexbDNhGJIXyu9+fX5AwCTkOHs+CDAGZYkCZFjCg7tfkrPXLVzFqi9tmY6rhwfg72RaNpHHplvs
qOnQbhurklnMItdCKApbc4P58oiTOp83c8KR1skWkkSNBwoRfxDS4nYsFDz4ojxAyd9VHvaDNRkf
4wQknF9JiNS+4djeAQQuFQjvHjk23SgKIXbF7IZ6mrprRmn7GiKfWE+Dq+NGXkGmFbB2atRGvPq4
6s2bH10VbdvTwUV4Uf0ma8Wv5CwAfdQj6mNak7HDwiWhHpJI7KwMUcWWFD7bssFrQ8phVTBblAll
T6tVrHWUhsvB5isKGRep6K3Wod60sVIq79AbwN2R/UdYDPPpng5zTu27j80qqGj9Id+AOhY0QZMC
VRoGRqe6a+TzO1bvHX1vYkBMfPZICVdEibXTTQ0niFrM9lx8sgOWt+nEelvStdfbHFsOpwgcnhV5
qxVTQrWX28/2fIzelTlMQa4/BeBqUT+55Ym1wxYifg4JLRNqK/V3lAtWjIXgGlbwEPdPk1+ASdbQ
oeupk5T3c/SCoPyFYvu1fvPt1M0RWytfeqb8NHeNl4YWneFo3EmEwRADyjxd8O+wasgOXr7tbAua
s7M4w3f93sslRIv2nZVl5O/E/73pxgC52NZ0RGps/sIi2TUtKGMdONEPIKI/ledIw3GDmDLwga70
lVupYfGP5G+mCCXkUqikKOgGUSUhdMZ7AMQbWulY5va2e4OUXXrj8kjc4anWAZoDkBbvkxUoFvPr
TxeMMV92WoSDoS+LEQzQMdB0F2xHRxJ3WTHv6npOiWGvPW6UI9wkUb8zRL5nOhkC5nIVT9qr8/td
ee4Snk0DDjuBB8jkFO62RVogeWuNNdQYK0zO50jZ8+JRx19z0uxSPSqJsi8yHXshO7kPBJH9c9jp
eJqb/ld0+tyttQ9uM5MxvJIhvdjgm7eOu+p4G57pzqL/H8bwME5R8difjqZE2yeCK6tTuCChd0Qe
cTwRyS9Yn0GGLxVMeAoJMvcTdK6p+2HoGwRGth7teJvB+E3Ph+Ql2TFZFvEjMQOYPJYVZIoJRWnh
6JvZkgM0RZrycgSoWZifP7X2+1pc+1zl76luQ9ds3Uiq7c82USIpl85iE27iHzSHjgUFGTTMsFhN
MtzMSob92lHXE0sUptMmmW1+0twDGRvCYT/sTqqXYKgDCW9y1p1PTIe83iLZZY2YU8vVJ1UMhpb2
V/BUHCR1yJdXO2+u5SbXlrw/SoAmrMy/ZjC7bfNe0AguubnK+O9/O476AL5/fGWxJwH4YocDmqNU
vLkdmOj9KbCGxPWFeILBC9aCxEdPqQSQUqbOrPDZca+OXsQ6Kapl3W4LFGjxuu+WCfxDjTlmio05
kK3gBc4AZWLZFUmM/MOJ39QUm4ErhV7Fs+1BzU6RfDCpyN5s+TcEo7/FeZuHml6MBH/uwJhFbd+0
u3OcXEZHu+68fPKYdlqBWFkDxe6SVn3UefpoVEkSuimwl17lPs3f8lSXK13GTJ77gYxw/XfjA14E
KkA/btBklBPOcBn67QGLTLhLgYJ+eSrxEvPvAMWHB9oVTmlFUDb04GN//c+H6Jj3FAxSShbr+jdI
zrZnR+qhVRLQw6n9HcRX3rw11Hf8JCpwsNnavYvVUvng+9lZe2+XXBBakBy3idbapT3wqD5VY6yf
kXW2mM8PmGHN/rgOZZgDtZmBVLC6yJF2lbVwX4KdfmuurOEI7moOMu4aZ7WL7NmO61Vb8fl9s4xW
hFZ8QjEZrTr6vi2+4iBK8w92MeqU4CFna7ac1X0e/RjNLoU7+tZ+/OWGkUmoBDEoLwfN3BexFfUF
Iogq0I4U3Ydz9iTCpLCkY0Pw1wztfi1EUxg6ksHnEztkF+rlUQvkauN5Pdo64SscGpeEIoF3nOu2
tiNyib5j82XhCXG4OXBTbVY7trE49AJ2yxQv3RhGkQ5srgHIGUHWWmyARD2WARinsh3WqZ4DOWbz
9t0K3nib4p7CTS8kgq08vTMc3z52FbF1DMeEyRSrg4/ZO/A1BFefTxVrjbME7JsKztbb1CRXP9GS
F+nqWe8uWUXdNZbGMSCwviRLOvDYJC+OV+CzNIpTk12VLuTl8Vj91sz2sEXzbG9YE4C8OzU7J5mY
x2nvBD/jxyCQdFP4su43ECZOU+FVwX8TuWHy5Y+TINMS+ybfhEIzQERB+81NotVw3qaPNj1HgT+6
vs7I5r3FoaCwHH4TppTdtN+NMpl0h+6YSMKHPqqrJDIkutJfuVAvmfyoAp1EKkoPN8ybhFeZLh3H
FhvQaR8nOO7CDH/GHAV3ij/lfqOzfyziEzRXzNesE19f3sruQCggxBe4AHHl6pv4UXxu+zqQ6tJz
DrN+mt3ftXE45KfHHCDPf+brAlewsUlu4WhANf9pzqJXayRIVFWAAhKlOXXBE9F1MB32zUwTON2a
IijouBD4qHCJuf4RqwKqc86RS4YW9p1SrZEjvyPJlM9UZG3MFNpVg+io1KeqPM3inum9mJHIX56X
IHkEWu7s/9uUnv97kCJBaw67U8zLZmDKIgu0tEfbCCzimXGVU0XjCZWYKPX/zo83cd4gl0ughsZt
XbHJR2ONC8AVRvSkqMhMXlA+LGCaTLIvII9pAsg+ZAr4W1nAP/2sRR/QRrZ+IKuRg25i7h6nOs42
7TbVlUXkJ4f3Bn411YuVTjP++pY/jlzHvjA8RhNN8z6sim8Zj9nkQBr1K7YXBCrqdvhM+oFEqK57
iT4L92XRpwNg98VI0No1wj8aeidiENP1n800k7yDBXBNoelLsuJujGDsTQG6HAH5+XHyYp9o1ZKM
UFMqmmjbr4hk9Mib3+RXnf7DB03QTIrqcxNM4g6fdt1lAJX7rmgzbcxvnOOUiOv0k+whrss6b31P
disQHM3PiO7r5ViXLobIvvfh40IKQg+IEe3yBb8/fpMS1YcThrMrOBaYTT50qByrCDFtXxQ6Ll4o
5gTLKVKKEVoa9w2c031HWb7VJ0Vzy15tyNJzhcQzCyUoSD0jKxUzQKFksGihIRK/PZQE/Gs3b2lV
ZFA9nGNq5UDlj5hkm4moT18aghtve5HuLBrtO5cSAN3qiRpABPHuppX9lS+TM4d+exjGcabMtull
r+8P7T3mOam1O4V8itt1+y/b84S6eJM8DCnueJK4H72oQilvQgxhupvSO7yAysfCfAJmG1YI/23Y
Do9ipFgA9+oe7ZrVzcutcLINQd4m9MYIf+6XZReD4qw/liJ0BCaV8K0dviriKtEG5DsCnG49OEi2
Lzur1Tb/utbcw5+hYEC+3DNxJGlEyGbSpwUB+icHq6ReFA27UgsDJ76w/5tpa+Ozsno2GVNVgiiK
9lPV3Bhk/ORVcgO5ko2uaAfTMZQaHLncZCQyAF8GoyRRJIaLa4+X1IYCc6Zj4NlMytLdNq/AU1gS
iPhfbOxpaVW9ODwLlvnL0mngGSMu2rXLRwEus+z4F+5rL7PYUpS5p0SkmYuPQ0jQFOZrAkPcHP4R
UGrxCtXfeGTsx4qAq88739rcaglDaVkpoVySOj3GHAWFZWvG7Bg2B8PErldluPsauQ/hqjfR/se8
w4FhiqtuXwpYzb1zCAiEa1L4XVyC8hXdaSi0eTZOYmp56VFXXr4PPkwtpLeMGCiqyN9xWQ53DOeR
DgRAuPZmGRcYIGC7hIde19LShMvmUtV7ABMRp0e/jrFv7xaS8FGXSM+tIzj+FWE6Hi2FTlhvw7I4
MumH52ddA9+NfBfS/ZYxS6GrLhHCrBlYA+hqQfeX9DLXF+a/juHfWhCy2EPUEJNA34ZkX8Q9YmNb
iyiN2+tAathgrehf3s0IaLj/bzVudmLN+d3dSer2IQq3suPvTbwTITAKS0AL+zBGB/wuQ1sFJMZ0
y2T//spsNhQ5i2/HGLzk8ysQ8VyufURT12UZywFl6IWIr4Yw6Ggt1Qi2slmZs6k+AoSdTT5Tg8eE
hlOE6+yn5Z62+YDYGwpeszsIiZTUk20zB9OOAT1V6lSTxmexukej/btRzlmZmGcrj5ojt9boRUGy
KfTOt28Cs+RIjAX/WSs13dX3/R609Nf/3h6LG5NUoiLdo6KL2oB/4kWHmSToyX3K+NHL2nKvKAbU
s7O3eTnndxpG6gDSq9mJ6O0C2IPHuHTNGAu/whd3DndFPgEuwvfpHMZx5QyipTZKTgaRrre9Wh7Z
PzHwjNEioP37p4I3f9LN2ECh9lzxJBXcm76eu745hcMqRcCZyEZzwreHPVX3zR6nB2+/1PLV+GrP
/qIu1psmbkLeBuH1C1Xy7b2HmUNuvXvMJmaQnwlxBBkdSfSQLrKpFEVmgnngk/js/8YT73UAn5OK
0BFD9pFYZUBLQJYcdxSyKd9PfrkicWj8bPGAD6IxzjaHYPalAuBwZxIQzDVQ7boBIJ+xAVx9WuGt
m+AQgayShEF5Y9duy5LYmexYiKWhH3WVdnqpEYBVMtPgA5hjdNazOzuczRzXUQkM5LTBipY7hpZ7
FnFZ8lJKfb3rVyhqZgJwe+jpr9AT1Fyr+dFzbaN73OL0jcUir9LHtsJxNYQQlPdQ9epxg0r1aBKj
jiJTsrAJTOrKJ5HxAhna3aoR+qW9iC/bB56/2FAvxUoA+SSv249JmihuInd25HcDivDMGLTomcbT
fc4rI3n0gaAiV7Pi6DUIjURdxoVbE0F0rgIHvSEq7/wWo7MpAfMn/e7/u55cH2RaUYrdpMDVO5N8
T8/bGEKOech2l4J4SW/a0Oj439z4h9iLwJBxQPHke+Xnmarp01SNyLUbgG2Dq+sp3ilzj+8SJfnq
BaoIejyLoa5BvXlUlT6l7h0RdWSgQRegZsHYjncgETCC6LIPrP7//8a5C+1WtTkfFCgLnTI8ZTGA
sziTDsFU3YtYNWZcM+Y9QNuv8ZCbMFZCq1M3HLeMBRIQopuMT+DTiP0GhCT63MEHvLW9VbGaOd/0
ku7leSqLXzNmEpi5l1pthLPUMAZZ1BUd26SdkzTzlEdAnHzz0TiGCePDE1jH5C829Fn9oDXKrDtE
JFt+hLpcU1FQVySbR8RTyLccRkTbeerISe47HSWAv3jatcdhL5ICqR7/cXdq0pWalXUBEBWB805S
Av00CDW963uxmcf/fZTjaRbh5eImOSMgjbDou2sdDPyEK7NJmEVZQ8n38EqG+ff0Rxepy/J55Uzx
YXmPvis+B3o2y9CnIhiCs7fk40mDlxV1lJ6S+udc6QOUeJdJB2MuWil/XD9AOT0DyOgDxDZibfEF
SElzhVNOksB1JDhuoHRxTVV4G72Kly4dxkX+6j6pAIogE+dV6GK7OCPk0cKS+OEs2vX3A4N035Xa
oZB9ZCjaoO/HWPHlD4uwck1gm8C8j2qjXDzdyRewjLKthieb0HdDYMNNi2htDlxzQtOYdVWrIHhK
UgOuUp4X8G2gCX5Y3FR3pIXigbKxG9nl/dp0zJa/JB2XJCLYZOYD+Fnfyzfu9MAaNR6YVtUp8JrK
ixzp3BkEHni00N5sGfziQoc7252HKT0GniLzK6oMuCoGb3es2ollyeuEoD37vgDDtbb8vG1zJG3X
LT79aOFJlD1lKzQp/Hh9rKjgXiyn6KsHIqJhOVTzjgTdh7LS0AVGgF0SytL6dHZx/IPKmbwE99eY
5Xkhq2XlGzI4H4fTCgQlKdLTf0V6eueOl9IIEoNOIU17E0rjnivz6Frq8ez4GM6x+u54XJi+/8ah
8zQA0tgCfG7l1/Fd0QTPmdvQJpHgsw1YNhzNqDBekxzJze5lBDohtWKsD01K5TIYXQO2pVTCrv0z
Eu2BqFLbmeapspJyu7mktBkUzq8vp8obhlWYV8Vw49KecM9RRoIsO7b0rBVO6Rx59bHlps4qElkF
x/+ENNC9Dr9QW8olP7iFKI6fD03YDHj4G2HbYy18jc8xfVZfOwdK5N7xL4DkfOBbssxn3NrFtsFL
rs+eUi3E7wmAar5HPKzYDcSGYZaboJHADsJPkZymK1AqRmwxBqXoiedV5gHpTmSHvUbqxHfRo5ZD
OB8YA/O7P8GYm7mkCBiI8yf/tIUKSequm+CoElW60xNg5QcQmerOcbZN23LsHdNoY3A9GmKAt2YH
z6SgYi8VIqstTfkTxeja0iYo7aHJBWyonvC3hdjizcHCuhQaOEsH4VcQJX1Gc1hRUB1lFG5V4VO3
q/lrCl55a6ngOfUIFZ8hLnBsdP+WEQwOTet04HkjFw+VPkhWTS9F1Y4J7oUf4XzzBMUUQJkjrLoF
RO5jSaMSuJ4h8+ER3c+Aqe4X4Z6ul++V5TYD0lYvI5cssaTntnXcHpRdbPHZIh8FNS0KdQVshYLU
ejMAHO5Ah2aCCwODkT+4UMl6+3/PV76RL13bVyCEL717YevxUnaqSQ4JjC+TFowmKDytBt4ixdRL
N7CDV6KFhhRfDP7+sAERyPjW/snosWtr01CaUdxpujnsspijmpcHe8HmH2HhacICvzBX6Exiv6Ch
G7I3tDsTIFCU6KL4P/qIcV23p8OZAqQ2ryUZww+AB9XSaVUPBF0XisVqGMl38iGZ99H5sHQNnYQa
N1+qtt6FSVMMz95xwtkM4JXqMp5E0d+k1YGOZfQmMoXM4YCvPN2nx/7UwGx1PO6Wjr9qdlUxUf2w
VIm0ZbLifokxmTQGAqClqwnQQgdaqoaU7XE/n6+o30wfyi+p+f5LLov086+fC6LpnVt7oSqFX5Z9
id1Zgq/XivPfkDi/aqx56WyzQdbIBRjdnLwbhgOtkLZr7Of4jAxBfbqhNR9E4qlD0nvRyt/98516
hdgh+PQDQx5AM9hTq6dmUdavPBJRKLxxwVr5A8MWEJPcjJ90GuhQGX+F33052Hzf1Rd3zBXE/Kts
1gem4FoTw0ZzUNztVs32b+iyzxI/2Yc+hclH5mZmRe75brlIiYvII02dCMZsjqYlbv0QGypaja3b
oKjkwNyTbApbbmsJJMYQmoEHU34Y4aUxwRNi4NkpLIVLfufasFGtH5piqqFMX2rW+TkczgriS2bi
dFN3ojf0EGaM303cYiBqF484fCZI/33JItoaM1SaRzy5aOs5K92zhtihNK1ggAHhiT69aAdD9Z9l
upGJtoolDMzIWCmBAjGA9W2CEU3lAnjalSa6rkEerUuOuZyb6NvhmCM1fdEidpi381qc46RVYutW
2JHW2TczMfXXE0YVRaxr1BWN8YtMa2v+O3q9lF9a0kPOwlYay8/iA7O73d1tABchlzLl+zBbAQWz
lYVL+YWeKnLo4uMXCBkHg+ZHLkNEM0X0LIjR1CJtmx/PBm/5pEw/4pdXSHDxqIvanvkvzEI0x0YN
i2y+47hGcMLM8f5/jkn70wGjH9sMxZdGUEhBz+wyzQxjjaalSqqPpJpMaPVFh55SJerN/U/D395d
UwixcM1Ti8mvP3ith3Hb0cGicinZIysQSil19QDPjSvEvwcS5hSpvdr4E/drE7kpM4J2RHXeCXdh
F6Nnr8AFX2XBMo4YQubK94A+442BKQWEL1J6bg+fqQvE4YLlTjhgXsio2lCjT1F3p4sCOX4q+Yz5
OdQJBBGRfDMPcemSJLmcbHQ9oEQaB7TwOOyyYW3m6D5lrSvfegSH3lQ/NlMZ4I/lyKz0sFEt7hJ3
UGeBfGHSolcNHTG2WE3yQJQWUsHELvjybx+YaXR1xcJcuDfONqlfkovz8wqgpEucIMw5IhBvde5C
S/Cdr+rP0hBlWr/bV7Qh5YxyuGAHypFxJHiiXZeyw3JadRViPlN88r2eZa0g6lQsd++HooQ6KHA+
5gQ8xuPE1Rt18JptMd2Wyd2rVsof/f2QcQQKsNPpGkWum+Q9MXrd3QgqKNj+gndF+1zk1gyPB2XC
3FDMxr/khpbTp0Z74kIUTYv6e63baH1QGN9whSKcCm0Pu4oFHQ1rElqYOo3u5mL2GemhH5h4cdlC
4+8kuJwMTfnOxdQ6mt8hGpnnfbvHRtoNcrBvXv9vAlAa6s6Uc1o8+AgNSa+UTpmm9tboi0SuqfV9
WtzUwjMfh5FvBnJMI4AM8y5YMaLBpHvJs/8+toIhMT/PwE8HhFe7yrGZ9857ge4eH+1LRs1FuC7f
Ip/fXv72Y24jB1AuiGdtR/xHziinrKBEIVnnUCa3g8ZmDDkmpP/7ANbkXHbg7LB3evqpd11gwuds
3fGT/lOIaT2AHGVNIghXBNTOWFraBlpBzZxnpVmyrL6V4qzZj6pOrIPhzhxbYj3FKCWKJXj9sC6K
HTG9UdKnr3IGTZE8GkeDAXhwGJmJS8Ki0k/jCWjptIghkeNKcHquXbrugZTxn13YOqHv60ntHB2d
KVKOWd0Brxx6E0y44n5QuUc/Py6X/yTdz304ZyQlW0CreorWjcpcr/Fs7IJHB9FpGqT0SeBETaYR
jrHQ57LeHM4wSaqwbKHhbcH3wyeGpjVDCLD03U0TxxRyfRNFlTG/3mwAhoanmIeTd8v8kUn/RDTy
/CnOdH+ggXlz7U6P6aWB7gru1A6cxb+jonEmvQZIDCHyUBpWdI33ibsg1mA7TiFXWxl/5XE369Ra
/qnWoLGog3JUXNVstP2ug3jyMh2WGqPocbnukyc+bngDR0hibvDHHmN+Op1SUTmEqqyzdCD2fO6D
VJjcF7ozGsO3TjcpY94IrC8La8M8SClT25QSI3+5DdL8QR14taaqrrz/2WH6JbbuvENeuO6aeDCR
rtIPhzUrwX+kKMndkcyM9OTdYURWWCiK3CrQC372i8IDzk4gVqGlacBys9+ezwbQT2dCDLzmZ3ug
6jofPlMt39Qk2XeFZl/WLT0TYZkdrUgXwYGzWF5jWUWIakYQpuo1cCPNeHJe5KV6XWyKni32ncoe
2pbrDIHmZwDIMqVBvys3kb6KcFrha4GFclIiuaO+/ctvai6d4rhEDCU4emr568OMQhZdVQaa764r
EH9QVslFOyrNfDYp17UodXJDYwNQko8g2QMAmsgQAyorL5eSAVG8GaF0gWwSgUG8BspbJC1laT+B
3WD/Dmkgz7mvI7k7KS8Q9h6V5RHIpBV5qCVsjzviShGd4GBeroA/ODD2BR41gYUCg+GUOVdAPPwu
cg4WBWXafZLRtyKcrRaLwUgULX0MuLJUBYiHwlhn8TJHzC6gusWHD7DlmYaWqQYE3tE9jZitXIhf
o8lxe6flWzXtntDwLN+c8RvFy1Pl0M85QIkY5XdSCwdXpuBUNenQLq7dsgrR+AouBe5YzIpzPmiI
F9eioo7VL/Rg+4MYlS+U3p94znHZ1rkE8sZ7Yhm6aEbztWfX6xjujh9W5/DsXhluR5/iYEsQiyVR
53cQECDC71JgSNuh1ad16+7ozTrHdpizIl+yDBO2hE4jDhfvtkiLSezzreIm2yVDpmihSyWrQ3eN
4rWgUbp1FT+srxnRCtqTkKxswgRf+DbLgrb+3qG9hL6FpvdiBoQ7FxXhHX2kxQ4E+AYuHmwuIfAw
o0XjKFTIXMKZSLuKLcIftacqsim52HPyOWNdYLLBPYWrLt4FQdHbNOonRpjgLpJc+vziohO2NnNK
eZ3wVi3ZFxI3E26a3K0AF7yIOGnnimqTLzjjBjc3+QMj9vGtSFZJ4iLr4oKC+ggIQi9yKEZmFRJu
xwtku6ce+b7o+s/UxshRiq4CBr4ble6gNQFXBVnaeokED0k3cXMggbAzczEDa/amSLvmBhr1xiHO
fc9b8ZQGz0MsBJ0UujCkXe/8pMvQsRXzAarQbvxhg8KDn9pD9ruEPYs8lTVV9WiTGsq7+Y4is0OY
yuWpUnE7Qeaw0USMlL75JjHeqWbLFByjdFhR7Ze9ZrpNQpiLxhekukaTu6tmjpwHpkiPKRrW6tX2
IS7JZXUjNgyNuFqSVSglcQ6ZylJ50V9LAysu2LklVrsIGxaYQKWtyR/DizLOjJmFRWHxeaxQMo8F
AYt1r11ZLvx2cdDPMqnLsN8CV3W7j/ocVbIZQKiAMAEm411Wmd13UF8SSv64MHO7Iv89FVM/SHQo
bjM3QF2Hk18x6koViKsuqdeRX49pebGy9WH1RXDm4Gnt4Z08kOEbSsHQJaDto5I4VGfmvEyg5D63
PYsIjb7szLRHlfK2Ws5h4BJPNod000ak2y46j6HoyTcva95aGOzjsjepZg8jPZ8pIodkjTQvHacE
B1Sl/LDDz2CapEYHeonKViT7j1bvbRUTOnHm9h5G8WyoEfEqv4IkvSWxeBc4rxCZGNZ/moVyoxoI
dx86PKWzHmXhLRDp5gjTMjAJcSIsb06IX0W69rV/0Rsul33n1UKzGXqlZ/wtBK9gmE0+tcnnd+3I
U+YSlDxNlVGBKORsu9f276JDy3Go2nf04CPlrfpSzYYEM+bkCRbF4DvxB0wfyqr84xs0W4R2GnYo
OCYFfZsFEDv6+7jVmppXzF88kI7hI/5Huai6W6GnQW8aZGcZQN4D1vDZGcQmrkNwygpPwc/PH2qh
QOKI+FdTPZUuJhS3srEF9xFn8njlRI5+U6MlCHgWUqB2GQLiM9C2rr5lA4uyW7YaQHHzCepkuFFg
mO26W5MuOD0P62CNwtE9R1vY2FELQsw3jqkOW9oU+qKwL000Qkg25zxqv9+fbgex9PfzRGoeAxqk
G4otvK29EGupcKm2+xv2gj+4jL8dYL6jvTDh1qysnmUnHRPbpa3XBBn37rMk9cxB+eFaXs6Ib6IL
Mm2fBa0x9ysq7ouYwvE7a8zWweMRW6ySFA3Y84FwBL53Ez1ZyfpjiaLJpCy4AOTh4gnTzPCKuNGA
q0PWBScvYPbRG/XlB+DIjJY0JadaWcWO5glmOj848uhHKR53RERW7NNr6QitmqvcPqaTckxOkAxT
5HGbZ95I3gpyHYGtz/kZfQcnhv2blel6TYN4BbRvOVdRT/uFKnPPbP2CSDfHIKg4/+SZQjQuy8vQ
zwmQix0gyEGaeANYWXrsTt8jjDsy9JGe9k/ybffprQTJNAclzqfbA32QlUcgjN/iS6VVSS9e4JMN
ryBFFdlSreflbkNZSz2ga9VwrChHenSCkM5HiaYBVH/biLSQ6zw/7QOsNdoPlKfvEkV/FtbBfzO8
GRR9Wr7M7j7aOJDhlu8EHz/ZLTOb30OWtDMhhYKfHNQdkyh1WYY34UPOgQ8sWZQIYGMFXzf8Mi5+
2oxAQ2NJEAjkweeJtMdRFa7E0HjYKBpof80jmOK2IVfN/2mMwXAH8hWL0EwxKuaAJ3BRZXEKPydy
pg77b149Ijbs2Kcj44tcoEFRT/XSLtDpMApBCNucqH7KIE/nAXe09Yji/lx+AQYJ1NyJz69N77wH
/2U+cAwLhobcE5jb7vRF7HpkfbHOlKtNWQKBkzKW1ZGK8RhIqiFtvqzkhwupd9dhaVb0qpj4Zw0l
QAKABCxeEF2m1BQ2CSgaQI4LMhyGYCeAX6B4/qLtWVo+O0TUJ/aeG/W5wajmQjSEquZYIWxbSa12
TqzQX+Oz8efVHbtsaqP/9JdsPtQ7f8AE/+EVBYrBuaMKf5lVOGtmitQPJcsKUMpz43yuoJefnSJd
M5K7dJZKX7Cvao4JbrAn6EjTUjFnW1vHmJIhZowkAV9j/rk++hH2x1JVfZYlbW7S3rI2eETuepyQ
/kmM2J5GZsP3H8qj/WAANQ4cx6yHGvL76rRVtRl1Etf6rqTHAAKMFb/ME/lXaoSQSfmu2bbN+ZMA
IkTvRfb92DddRiQi2e/KDqisRHSf/ggU+tDji59U2qgP8t4AOtmKTxNv5th0Gfwvm55aDgXyLOMs
sQFmRRJnf6w87GjI/IU3QF5GfWyXt+vqlnfDfuetIG0ou5CCxX6dgofGjdjkvz8wxMu0hcw0sqT2
vHCF+mvgPDSmpK/kV6BszGTKfqpSpe32eeNL7dbkb8v9K8r2+1Tycor5Uc2XOFHetYgVdbibciyr
recA+YVn3T9avPQTduaX4RumRiQaWn/2lWdb7Vg8SlF9NDDdjUvOWrK/grxcptnv7IgxhM0E1LoX
7Ofw/xN0J096G/wAuH8PMjkLkhEWRJL3Q42pfPCdY7Fh6laSgUD8vULHfKfXg5GAgEnci5Nzk0oK
N8U5tfXKqi0xZ5iQXx4MZwNY0R4yveCwHRiQbBnqrIkiVqGDmZPkGlSMJ/GfCtKt08lJNl/BNBnd
EjoWvowMl4bVmnTrvezUFdkXEt+ikDFYjOi7dw3nN+pgJTOkr9WnrzRVX1VwO0V+/1dEV0LPtna6
pY6HyFuU7nr/+yz4EDvGolC18n7Tog6rqmyieIz3paWM8PNOhsAEIr+xC87s0ThXAA0bw33llKZk
3/rF38aYIEqO9WROE7VULq5ErEyXJo/8VaXI6F25QHXDOZZxTkXcjVtKqmFnnscz6A6uIzZiqg8K
yPdf2xUxFdcFhpJwpT7Ghg3V3ydboIlqzkecuH9M0xFObj7EpsnxXkSKBfj6+MYmfiCPudQdv4/E
gcRCFLRRhX9G9esoN3uAGtjfgYMaDCdE4rJuU65lxR5NrQLBESAkcj7/o/dtGUh/ILgY1MLZWMv3
XzUE3GM6aIDV0BiJ5bJ7dBS+th2/kR4DYM2bI10h//T5Do83jZpIX7TvScElbDZZGS/xci8c4fNg
7Z8FBC9JctMZ+tSIPzlksu8wNmJKKtr/b6DFTiTQsDdibLg9HhWCIJfDOvSH5nIF1ADUNjeXBdj2
4qBfVO/EHO11+RmJP4EYjIxsmZeixdUArq07hJSJ+xf/neS7Fwsctj+HtFbH2inPAadYmXtUy+Fh
v3cl/eSOodpHGWy6L1PoSvYgXHiNiEawg9oPNqzGR62ERin4RabA5/OcDRRFojtFZa+04rUguD1F
ULYxPg/jiNA3IbPVnZHKJOWJZVARoYpFE8JwX6sImTW4sUa3IadZOhPaUhsd//k/p6moXASs+8qo
c0g/251+9niwVWpYYmBQbF7fU3zdzRdBYLFNryqALBZFgmucdY5NPg8R+o5+6zotEW5KHwUKUQAd
nd7ku/NO48PQbhguOPzPiS6FNWT4oaTbNNvMiQO4CsmWFLzklL7TUrdftaA77a+1nnxTQY7RsBql
m0PUChVDSUKK4Kjp8bLx7TT6l0mPFGbL+KRBRm8Gv/tcrRIb51XWk3LNMI6mZdo4vWgN5S+2UKbD
rhwwDrC7+ot2KRTXFg1KCEUBcSvzTa2edJkc2jBAk5sLF2tviHCf5m2ijhG/zLVIc9o6qVtN4yt+
T2bdpMX4gR4QaqXNZn8VvhQLsAGl6vj8ixl9weau0Lxl913SIJpLiETie+HC8X1sW5+YXQN0Tz6S
NuWkKyMVSISW+y3rRZW6J2asO0GO06q4J4Bvy1J33nReWgqQG3U42e2vw6cgUETL2IBnR0NInM87
TLycFNGzqPr0cWt+b7xfsG3QWj4No857T6Y0FAhUzq0CLdom7ZDSWT7VouFDNxGKCoky7dDnq/sr
h8pxe8o9D9C5ra5P367SNPDKgXHPMZFHQqtf1XX8VdreJmDy6stf+gxP0iJkt984Yj/4DUfjyC3X
8TjwKDESAVPL6l3ALZW+jXBLN/RChZ7i5dZL870ItJ6Atms+1PQHBixoCfe6J9r+q2q1imlRBNxZ
oKj6IUsr2Fz2u1+3ri0e3WdaH1pwp1z0yc2Kmrc7EijLv9Fk07LuQSTGWgD19bDpmGW6qpqs5gxL
qpmqozxR5j+XuQSvXWVfj/lZds2+Wllz3ged9tj60IGKeNFPOtv8ogAkgkhXWYFRRMo8Lw4NbjQz
2nGU51pl3fPeNiz03+5Nj/3qZle5yLgsN40j1Oeuy5Bd9rjXWQVHxtk9iA4ia23TVjQZ7IbShjbG
e7eFFGJyGwEkkVNfM7tX2xnKE+2WQP7e3LUNfYGI9c8VwyoESgGbubtr1ajzAM87VzRCAH2kRBv3
uHsFff89GCUfhV34lOeU0tnKsjVOqsoM+w8mjHBzw4atH6iF4Y3jZ0AdQAP2bfGCBBNeHR/364Mz
IgnFM/jJduI0ciy6F+5ensIpdHSgDqluuyV1Pg1+00er6C4u9N95+ZbB5XoiPyO2oYyhEk1bJoWr
UnsTcmngEODKWnH68bUF0beIQuc+QjwOM4FilCFdtVrtkF6TpQ5dC8iuukzR+YF7iLKUTfejhoo6
/xZOB75w2960wY5bz4shAFkozOL8+5tkrO77SZIBHoMdWKpExftTkcRIdobeFnW3PczJBSNj2Wzz
lc2M7S0RxTMKP1z+fotMiZCoKzvxlYTJn0GgDitR5fbNjDm4a5dVr1yN1RMX7L3e2CgZ+Coyl0KN
sBfp0vhV0BNLbdBrYFSN2vJX5328NqLtnY/5OJW8vpW8LX+2Fb/t3E95ff/E3npueP3hcHpEZM5c
ZImD4We0EDUxkz6teOtNjxgVJSJmdF6F6uYcaPHwWrRXKL7F5ND3J5LQgk0DKrYEaHotyh/sMhEN
B5QbJtVRd6jpCoSFvyE9P+oHUAmyPzDGYyI4wOfT7PYJEHI5mhx7lZ3w7U+TZh+GJu6ydI4o6DUA
YCUyF/d3VrqhVwZMi5ifmKUUGy9YuUxPQ1wpbLL8bCowV5pjzIt1uIF2eZpEVygkcbipg7uIPQxe
3oQdnaXLDkN/AFZMVUTg/GHszrqiOgie1aFt9IzEs4YSYGjVJM8nVpcCyK/DhAsgScLs5Jbeyftz
A7jNsK2WAET3pnOuEU7gWWxho6W0r9jFrNtWpZ3c4JRdS0UmyMmc/L6hzYL+4SrCpbZqpGvwgCWP
9gJpFaMFfo5tl5q5HyKPfYwtFWnGZ5CAdxwn0GDQeMiHrR4qfwOgna71b63MDFpFGbCdWKLL8Bv6
LSEEkx5+ze9Cy1EdTAGgCUKSUp9sCNEjmkoVhlva5b/5as6YmCMIsdJADRtxWGd7maIGSfpS0s9q
Kdzu1kQbm1jjVx1UbXnWDuWJISNSaY2wuUdl9RoMrvpqQCKQJC89X5/UbzpfIJj9K7f1MwUR9O3K
EUfa46MBVmjDzcFfyUwcueguYQ8+NsKwyzo7iginUYmg3Om5cqY5IyGdUgFqdaET9YHnl5Yr9ezP
aLZeIBY8rrJEC8P7lv435rP+LoqB/LPYmGVfoM7jfeIVdWPsKIxcmGRAs5g2WTX02k9C/GBDS699
nXW2Xcd6k5h9GMeTdEStU14eCMzKTulIvI9PUpdzUGysWH6Ewh6IRYN2Jeja2tCCtFJsZngfvdsS
4y0z9O9cZEPLNTURNVmT2sHsJ/F2CSn1owwOzh55tAzthovI1ZzO7aObnyUyxUtwmbSddbTYq1RR
Ugh0tvenpi7CrUDdZimChihGlekEhT6g59CF95V8mnk3+qF1p8M8QR1/VJUWHe6KBGnIrPVrlA6Y
1rAQs1Nrt00xAVzzxAeA9Zp2NuBLrSuAeALcI+EcZ6YLJT/2GjfTRgITazMalE0FtHMyZA1o62Bi
+pQwC+ISlTwBZQ+i60u20CDFysFvqvCS4eIv2/QgtHYgQYnMAJedmRwodRIXL8ZvrcrcSQUYn3Hn
u3WeNi/4QHvSEl+mp14aweciQk40yUN7wzbNO6Q6YcQQ2awAIinUgPo5gi+C6VQ/Whor4nXzNlY4
thA9qHxKUC9A1Zyqjxjb29V/DJIsGvxjGI1D2DT01BUYQrqCgWTWTmOvgXjHHMiezxb2BeAo52xk
d6/FLkE1EBefBfeTHw1TmAMcy57y+XCJvt9WTvpv7PKMLvUr57HR5jDuiOOdR4f0AlLo4J7+X85y
/4ovMA4KFuUeFBY8Xd33hIBTpsMGmGAAGCzGUhAMaMCtFJh++4rqRFSsaEtJuS6n4GSN4JKp+N0z
pGqFbPU08zUWmf2mKu7OoA8pn0i+WJFCkIl9amZrgK9Vh12YRuekrA4GECBmD1pu0bh9uJM7B2x1
jq8eP1XfWv6rcIYSQ9CKx3FJ4H42RyHxwnEUmvl86Ttuf6aeXKPu1AspMZCkolBLUtvUSLfKVdia
k81s/ck1wD+Mqq67K+D9GGShnzimY/7II+ymsG/C7MziHQfvxIL4gIsG69fdPzZrDNbIMmvIEFZy
q+FP4uCT84LvrACbdr+lxOrHHxgAGtlClFXJ2imDxXXZuLksy4HpI6MPCUiQo4hdcOCFRAFUyhZu
xM3igsFEUQl0K28IkxC7RUhZwLRUbSc2++Tdfjg9YQ5TChmQGZQR3BUg6HD23GZ7WmzH/Y5vg2pU
dP6yrhWY71/1kUBsHaq48OtlBDcoIp1mq9Qov/CiHEA9JdB66z1Ka2fFzzf6ySrSTiuVTzCcWFcL
FUU0mwScamnzrWEgttNDcrwdfhAXyQN3X5jSlG8Al8XZygXRaAWYJQPCFNe78W188yCzW9KtlGff
7Oj1niaEtREdlwsnOZLAVSxggd1ry5rQZBL6uMLqYH30uxQRVEFaPGtEzW1+1vpBhtACER6XLIzZ
KzFG6BAHXMu0stw6SkTJOh6/5N/3INhaEn5XcTA1C/f2eZZu/4ut7kqdu4qqnvwJVY2mGO7LTIJ+
Y3og6a/LU+YlVqZFSL3kLBHBejR0WM/1hdx/hyo+6Vyv/Sy6jxRMxuX6W1/nBxzoeauoEfaZEjbo
Puxos+qsS+AFooJ3ymU+R+aEAmI8FhUBi/WCvzlWAKsEEhjluW+FTwbgurHcZO7zWHQ5GhLCCYdV
2BJxZ/wwXPmXeTgEnKJav5BD3JS8rm+mLH8CxlcO21FWLzdADRCfL6i6RslWiIKW08dMtMPhOE/j
MZfRxLMAvykC08O4ddDDcipAINqRscIRJK1x04AFyRapDMGQWUHdKMdEesY2E9qA6a8MIxelmG2+
Btlvw4pcWpnYiy5vERA5nqpc18t2EJoOfK8O1ByE4R07sk54JTtfWQ3xOSjieTtZgiF9Jn8kb1Ms
ZGNguQYqQDUIWqNnIW69DmEefkx8kKI9QlNoKywweIBSY/lkkV1GW3fNClh0Hh/nRajNcUswv3UH
jWCDqjb+jd/Y+5cc1jlVhgB+BQum4Vcxx58vJxWGnv372wPsb8IB0nr8zK5HWVzkn59bXQ9oDQXw
3ImgjsCQj9VBeCoz0JBTJensHMRnrCyzOFjRdYm+eyfyAJS43GDKL7JL61pfpq0kMgtJBQg1SNbZ
WHv7GyPHuLRaaU382k7vhfUHUu3fyyDb77R8shB02WWLrpCv5XVhEkFSNvFwBmAYCDRXZHQWtCKL
ttGBZ+JYFE8b6LxzXV4fT7I6m+g4EMu65L/Bf6LSAL9JVV/ABTrBQHzxx98edA25fOf48kbJAi6b
4gbvoLRvWVg53LyAHtHHCzCAhP7UJbTmFJAspPPCuj0BuJZ2yCtB3GOeohX25xT6lMfu0OE0biCN
W4CnquKvlL9xcXcTa17SmUzUJf5njqNupLrBmJBbCENBR0ldZWQDYHsQuFL7Gz1TNV/o2c8OifFk
WRq66pmdIa1P+t6ULrl54ILHyBt57vQ66SHwJPSGrwLlA1/WvH4eFtIVcScZapn6TA3tZWEGmGfx
XSUm/H7F6YAzjrKS+7YcuiYwB3uf8dDDKJisQ5q9zuRzxRgRekK4St8+J2aPg2QwkI7cP5e+wFo+
1VE9GKV7TbuPl2/W9D5FG/+lmV4u+muREz/U9JZKC+lwRFUtrw3kRHDrXFmS2C2iUvAdLpwXQeSW
b2lPxxEBD3wevKaaQFclOpsz3oJylYnKaVclUlIzSVHHzLHkdapupQTwkyzlhhJ1p6vh7KSVOo8J
yN7VdCzhbw1P83DIcYUSdfOLAZV4axOYwc1GQO9bDCB5lbnMpATW8OJuR+EIBhuT6N/fbCR08VtM
6ohDfk4r4EbbJv4g7Geu8+r3CtHlSxNpyhgf+BQVGaDrfT4MPRrdZD8doj4PUepEuEuTw/S3Pl2w
dlMYtC0PynVxi5udL7RDhheBd59Begzjlz2I7ZCLZ1OiPe0Vy6ljuAEZ8WrmmNycfbfHfHniS0Gi
fsYEhQxcIaQ6+SVXqcJ3598NGR0CBXTlq5zOCHdPlTVMD7CGP+ANowmLfp1BLUmXyjrMx84Lm4DJ
HrrJvZ6WiRlcXeUv1itFU+YXjzgHgbkVUWF7W9vt81PnT6h4M92wfl/9qQdFM35VuRlUG6ML8p7g
Kpwpop09SoifUOWs57QmIISrVKbT0faacGijEgCy9Iakkd6hocOr9n3lDRgnBo8lbZAU0GgTymNM
DKbwIEfUbakyEA5ZRAubJnXwqkSSn2v6OKnYAHkJvbFlRkHvLOgfiSASrtEk59t66PV43nJEmK9y
3NnSyZ7qCFJEsON9hQi0rgavcC9tW3LOFYAm6/OySV9iJVYVVQV18JgepBWXAmNdGCU0hpHpGqyl
ev/qOOiUYOt7SSrmv7Qe+3OASLtgxQcHCTKGajEJY/7jid49oZaia/JTOQSkKVBR5eaBPPMCUlNv
7nbw9ZxUfFfZWgUX2sa8CS4sAS1+AlIpbrlAaSd1mgKkmOSvd6LsdF6iGQXSljtA4HtS21WBcHJD
Paqp1S3zjGQ6iS3AHYLwzbaCwqBAm5ODJD/z5UbLfOkBGbJt7Kduc4tqDQjfrqk01gQ3ZgFFKaMF
wmunSVTmaUG45cbvg+qm3mDDA4OW0tHzo+WtC3fXwRx+o/70/bJJBu9YugBAp4eIfHCcmVR0q8UM
kHhGpExi+EwDFanGlPPxToSVLkXcl70rYNggT67F3rPkT9B3iR3AgKt32gsx9otmtTJmONQPOETf
yg+rUGOq0PkZnx/WoStC/VER8l0jTZ+U02PtuaBNUChlBA/xKB0Sm2exuqcHGQQmODtm/dV6LDhQ
Usnkz/zIYHC81eCAT3pa1IlyVk0GE2ukfGiAjDt+otTBufbWql8T6VcvwMR65fQ4bDNfVry3mKI3
M+GMPrII8Gojr0c3kfGVifq+wKbl0bwPu5LCJj4rXXJVWrZBzsFmRVarF21RlqzGok2qTWqYGzwI
TiAtanwtq+SiG4SHTsaRd5CKSbbFVctxc9wMT5HL4ji5dGpu6QcV/N66YTK2Yb42rXBiCWLKkUZN
Cu+197nuoP2lZ8Y5aEzfwLooxioXp1OfIqQr4J7BZfgryplDl0TmrvwOKXMQr9fow6CeFLw2jJRZ
rYGeqyvlhLDeYOSdpvP08cKFoxsEVPbK3dRXIBGBb1FVtMxWiVasu0E11BeHXsuGXC7yb28TIJV5
yxqTZzWbA5sQXk6sCxHEusJ0eBQ3erDfKmXJaNx+xUHckkAiTSm0jh/vgoitpHVGO4Oufan2+HNG
hKDEVmCHcscdDk/pMMVN6NrukivWTxD/oMS1UNu6nRwhUsCmvMxXecEu9OUTe+HEpZUKAVagiPjQ
8RqSfyT7KzwnZ0vZkU4LLePAZdsPaPAddrgKEzITBiwXTcUROlaCya+dROW6VQAeTxgaJoyiBMGF
rx3+/IiS/M5KPo1IMt83yB++tfTOM/fK5Dl7Wwuv+o752+AwQoD7L3/ep6JDDQw69rwH5NK0dpy3
snQff5Kh3S0rN12n+FHv72avPCJa5iNPf1zh6dXPh0tyqNnOcPvr/smi471MCnwor6hJvQQl7ZlJ
ws7vmWVA73W6T2tiKTtWXEg7Sa9n90zKoDuoyCZMfSc7A4nyfDGI2paqiHpwR/Nz7dKjqg0RIgEY
LoJKJsbn1qJaP0UElrM3qBbt7FGFZFnU4PiPcPcWeLhdT7Vqk2TsYnYL3mlXRN8XHz+aZoAzdiVl
hi3P22R4jlT4Ch1rTmc6PW9aUVe1nLMWFBsw9b+75R1l6T35uIivHujuaCzOMHMBv8AdW7My94tj
pVOLz5r782ZSYg+HojAv/oLSj1QanArW738O1NZBEAbK4iFYNmwPnzQWGb6xvZJguYEa3A82NOiN
G+R7bKZasLGNAbUPb+AGURufu4CUjlLj6Io9ysx4hOr49XZpW5xXuSxbkshbRQx/ecEgOaLn6KoK
FMbbJ2dRetcAhL5/xeUty9zSEj7OsgTpnYpVB3U2DczebuMG3K2MvHk3cjaDg22U4oT6N/25kSai
ohUFg5Rc8YB6Pgdi97o/4AORNtUrDvFM1YaVsPIuc8Eyp9jGGsJqWAoV2hpmHzdnw40czSzYjM3C
2VOO+iIMkUs9Q44xyO/qpHw62j2Gmm+i2B+cqggPPv+SW2s6xv/X2Otxw60d3FqiOPjaVsquxjGW
AV0hiXgAe4zTiKUw0bsHuS9WZmaxUT2VcRX4igWpu477+HYcJpggNwYUKTbMWm6Kb5dWFtFwFz4+
T8FLnRFHQclFMDdQDuCDUr9RP3nPAtcRwFDvrG7hmSlidszsM9CSokfeReZMAf/xcxqbd8jjXS97
ReUhXS6WqgXqsI1VlVButacIzNtzb6Zy/AuFUDye5YZ15jOZInuvc7+k05zz17Uth8ZOlHWiUM0k
pkxk5cupar3+BbzE9I/wsd1LevvNJKtISu8dIOaeQPPosbUby/meelcq2JYacj9p0g55Yh8epllS
tWjkFcVIhUa4jI8fGOjuILxPwdSMVfgN4oi1Oa1aCnaZxMvKsZkWUMpRE514AtAW11bCStq8ES7C
TXN31qgIXIVQTOKshPAk21Bub6GV8LXRY/4Vg/+NDvatfaER34PenmLhKSU1XEc5EHxsdyOu6H7b
Xo78qSrzgezD8Mfw9gwfz/W3EH0GUlLSdnMLYSJbujb6AMLOgYto3sorSJblAehdIv9fG2nAiZ43
ALs5n5zsVhkRlQHG6FoJi3kYomzzfeHSM1wzsW7k6lkvXmlrxtaEscOrbKaJzpDiYA/68nuiIu7O
oRaYkDhY/2P0nlwU8Zf6u/EXr9jMco7GNgvVqnXWF6bV4guzR6sNU1zZ9mF2PDdz+nCRQ6E5//gI
9ozeIuT21VnyW6ZgLhRxWQ2/N62t87ouTZ0J1nkl9o+IT88s+fp30+gGXRxjAq8TmGr0Zzlk/ELq
3WKdvTuHembdw+cndxesD8ttVoVSf3s/rLXGWK5qWlZMwxaIFwjRrzEwEjwPSIkvLV+EWBwpUnyS
Dn5y/D6PrJ+5CG6JMgxa6XErtZWrfQ5UKCVM5E2L4Td2s98UdMcMDXPqQuJf63wmqTJWzZzk1I8J
Rv1LgqYstCVSg9RdCMw9at4qGWu7UCz+4lMTC3xS2/5PaZJoXlv/p9r8ZjNOVYm8Qqny9hN/XdpJ
UelzRi2ReG8R4H4vc5xUqIQEYPuebblLH73DNpZ/hwSF5hRRiNv7cN2S7aUE+N3+a6MfghoahM3Q
FBbKSXih9XMF8KFuVG0qDBr2wLe06I+G4ezDWPuBq17VVEqda0MbzNEplLz4hR74lM7pCu6lEUcP
0QeerHoDNz4s90Y2KFFhqbkbNBXMqCYznu9yLd1Cy9V0vDZtnpqFKqKfLlCgrrEDOrDIFFNUsUWj
HhW4ni5aHY7Bw+E593NBbpKvNRlJV7p4WhlEs2uz28I876D01TccetGwGBpmAJMuwG8bcPckMCTa
2tI+YqSAMHMOtvh/qX/4HwDkxmPE9M9mbHj2tqi7Ge5YU2QCk0N8cFQEyxT9JEnnC0riGiIyf1OO
RBEqtRE3980M3Ytd8ZF6GvKpVfjBG3GeOcLI+jaMoNiP6sYjktGzpA9ufBhkbrk+8bW6JKvBgV2Y
MwDX60H6YhNlc7i23jW+cnl79FAdxCnG56HkH/XUMmfwrMaYJJTh/38ZXkLWClVIBxu7gHU6THb8
7fPdNws3BHBdMndF1JO7Ft20x18rj5mNt0h51IxQLpCgie9qoaLjmkxvwi1GeT5t9KXBdBoVVeds
hdMGMA736ihJ6zWB6bNnxGySB/JnN/H1dXFeoogiVXYlnDyXnsBYeWRwSeGtu2b1h7jZGSSLIU6/
R7s0CHc2DMEqxKBhGUITtNEUbc5wahtrPSuBZZAzp+yjyo/iYs2zY+SgORywKw1I8LwM7EJioGOu
rW6sCyR/WRFPfQMVroqY3Omz2g8QBWqetweQzbDZo7W+YDu7Y9oJEQiCsX1gHaTxHhrAb1Px/v9c
++XtoL0ltQbiqleni843yNOSdnadB2I00infShjPoP0o3n3UvzJ0FCTkcBy5zpI1K/s+XBjpm5yh
2rWksGTTTF/ZW7+8x+52gJtwJt7Gbz0yivJTzxzWaFIROKnXcjwAOnRs4LIc9sbvCq4SAlQNpFwd
I3wJBYfz+cYQB89IkEJlLoqS5Vm8YWVDEgR+X9CbuRXxMVg1+w9YKlKwEY4MTxTAm7O5PmT9fInl
GpwvAXBiyHi50qKTLq21Il75IeOaECr6YAzvnLKHsR7Gtay1VZdiXV7D+BfjPVQUQYFl+vqiY/nM
YYAFLAwQOy0UdVI7kz3y3PPFtZdNpPURAqbD9Gm6NvAjom5yuyXr79NVUOZOUyxIG2gU5wiEjUEi
AllCMi8BSlWy6+D8pMdPWKOdK9gKrrjEg2pmghCwDkvcsD+Gyc+pQvdZDlVBajuLQzH5Ag31WHcL
ldw0aenr8oKelh1xh0Nh2dql7PRub/bEEdZM5L7KlTftRNrHP6/yZYSvrhjY+Rv7Ma6Itn2EKpQf
4OGS9mkoowp3SNtIpwmmewJfat5xbqiImv55rtbbU0X6PaTQUOrR664P5ouDMEdShDuToTvWIW5I
jhZVXtWe0mEDLjqXotJHwX70/JSt0az39ilItOzaC7zOS1eDTdUxQ6/RP7Jfid3xYe8ahDL+S4bU
oJ0invMuDp9Fc/YTh+qAEf1GjTANaSWJFTCVkGR01FdTpSTz0i2gqJgiZA+q7Qc/R7Mg3fnQ9dpW
RxiqEp+BxLABEjY71FUBfONwPJOmcCLDsEZFqa1HxUAJi8XGj6PVswWQHN2fXOGfCdJwpBQ8CHLt
AZEdVtnDEDtY+HE2o9O0XrrXgmKkn0bGfXF1g5o2uRXMLJMwzsZN07zGP2YPRsniimm3AMH81tQ8
xTpV/tgpku7VvBp5DJboBwFRlDgHQeiIwFZKbFXxQmIofG+JYbeoN2lW4dUie+UHs0D68dgzVyuE
iAocf9iy5tFZAI4cZoyCMKMZzFa4UkhQt6QjXQuhD1gKRPumbvSaZU3UBXs11dRT8hUCT+d+Q03M
Bllg98rVXpuO/wuMtC6r3DXNCQECYR65Lt7jzehg3ThKd+VaEiJxgkGb2NGqQvaJc3uPZDsfHHtm
N+csiY5ug1Zst/zi5Vc8y5Q2B/PSuGq6Uo+5A1PnXl/IZ4ZzDOvCgAymtufUfenCODCVkzpb5ULw
20DRyL6kNbVpC2vf84skwrfdSYGTiXxvm4OSLQXEZegAFO1iDnuh8InmEx2089zqdZpE5BIFin9c
6TJDFCGXHIBw0nqJfY/2bEEjvHJeioA5mwDhcR6BujMD/BeWOQKvYc+YRK9VRaLKJjS+Sv+hYpIa
/SZpzAv6boJEyDwRBpT3W4opFaf627lxO0+89ADPV9iUQ/ClyYgWQgW3RYkRh/rK04vngq03O4Mt
K+6jNRR2VoFJelHTYlx+0+w3BFjeOss/hUwpgvzuR0fCfIA9Fh3PUAnu5jpQY4Otip2wc8sJGIOz
6pBoTb7tDMG8mh9xBaI7vM/eUoR2tcSjefd2rjZ426kfE/zfnXzHt73iXDs7S/iwr7xm7eRGJ+wm
TSrBUGWjefca1y/aO17PWNcbbShLunajxP/7VZUhoOfMrxaAPNAY7nCI1MjdDJj79WaDWyq6gich
2pIAOR4H7OaWyKYJ+MdDqRIIqCLqpqcR9GxcKgWUnDn58Yt4CLDAg84FBoHpv6ine8lebStNuc9o
A9i/a6YPSCLhpWJ7HFXkZV83oQwbaTpZwSdCSZfQXERSzQl2WJEu4bCo+EU451s7lTCXzc3yuv8W
Nug5UZ0AIzdRGFQTPz7cQipuTqgFiYhnKyc2iVwRsDj0hyFPKYb5++eyeNGA7plcstiD8NC7jqKS
HTuuenrhfgqJPPDboFCqs7g7fl5XVHmmjdoZTJxxY5tAfpz19cBxBU+G8/DsKpomLWCuevVfnWCv
EJ5Ss1HYeUOg9ps2otyB8AkuV7FcoRMN0f/XadiSAZwq648swu8b319TTvcKdCB/UBc+0gWe/3Gd
zwzQ6M6l1U2cOgwb01AeloVJI4wrJAjm01KLz0s+97BfSP+ar49b7WrPhFrF4EHHu+w6sekZ16nv
0/noop7zVDy+Hv9W+Mm9cp4/F09eJuf+zTD9W3zwq7cDH8i+5MbGO1jTtjcquEZ5J5x/yWReT0Mh
KXDKyf91d7OlWssGCWMF1rk3f6LTjEaCZyP5a0yHcri2yRY0bAvHVUk0PzD4ljxWI3gDCyf+njeX
mrNZ3iMyrxiwlZ4FnpNJTMIwTbm6Zl0CUzgHkoXjOdFsuaXTk8azIdFIB57p19cHgFCaXlgRg1w/
lE2FTMH1yfNyxkiF45/NVNEsZCnuPqdo8P/Ia5UPcpxHj8r1zh1S3NK8AaP9JRev4K8JSkCZj8sU
Y4VILzZoYi7yUxJWm6WwLmnKuu81q5RSpg7JXp+nWGaiy+SirQ3qwZ8N4ckfqp6w0xG6WXLt4zHD
JyyBvNhIXY/goDj1Aa1zg/cpEeneaPdus24mWh7qpDYC5AHgesZRADz0eOhCcE3wzm1cKz6CZjoS
5ta5JyMxIsa51ntB9HwjhjKV6bD6rvVloYd8i+cQyw9u51Y/PvMUH/fO6Mcd0FoHjF4KHBEePXXX
grbYTi2055D1G1XTEtA4RXM3DwTKrxvuVwbKGC1BhdWa9zCKuTIxn2sf/nOttgkD2I7dXHZTcKUo
H+B1HJoT+ylx6uOcCrhprKdUXKO09k7tsZYldNlKW0+RdAaoTU5VH7fBPCKi3dmmzqFMy9fVQToh
5llZpvh/ZlyZxCYfgqxR8HUP+HZUW9kO353apTjn9VxR/HhxoOECixmPRRmHsXJKzv48xPbYdKuD
6h75EaIRXiHafMeFfLoWpg9LbH3e64z8VwzBJWfhxBKAs5ZPtqIMSgFyaUPckN1VDVZls9ffchuU
BXS38tzksjq+yCUIQPgMltC1K2i/kwHAXckTSpTBHGyblxjgRRJChKCaR0qY/CblXXEs86Jb+xSI
r80TbblWoO1KklWc/m0eWrGKtbzXDNVV3XKjbQO9A3T5Gl6aXo8/9BH8DatBY2xOGGibFjcTUMzT
lnLekMDqUamf8BGIkzDOIVes2Teno50Wl04oXR8ydt5s1PilZIrFIxT+wG2XKA1VhXL3ZlsGMjrz
MRXts0iU3udpDuZWmrAKQ3exHd474BKJUgp1h5rSJYtV9M9PFAVtw+v5m4DWiOrUYLW1Pa8ZiriA
gIS0K7mx1XYwppcv5e54ZYeotSCJ54ILQK/VVrlfAD4ah54om+mSObklCTj6DzX9qs+nPEPsRXPV
RD6nOW+bq/EYMNK4OtVYP+bmU3jowj8N9XaUROCoh0faO9bI02gXfsSdVSL2if6Xlxv040n7Dnrn
d8ZklFTtBZYikSfzCmVBoV9A648x7SijvmfC8KRi7D5tYlY2tQj9+Bmn6d7nR5mXLPjMTJaqSzy3
ZOfNbqjbt8R9XFGSaNiJ5SSS6k8+vUACz+5kEgDLIDMt4lC8gdXZu783Nb07Q+yNOuIp318UTgKA
jv12qhIoIMMhQqd+QoIBaMiFM4atlSFdSG0WR+Za/JVeIyfPYelCvJI3CXwhtLKqx7jzyHR5/cVJ
danzswFi0pvIZ8q1p7x3eDGOOAAWaCpc2/CMbuKbQBh27019/T9mduKFpVd6HO3AZFzunOeTT8AP
Cocg6bUg4959ulW4cMwiy2AWf8dFplQ8DZfhZXZusc8xUHurMu85XcPa85m1s7hXNvNBHl7Shmyd
uOdiIKEUUFEOFpB1Zaqx/py08OOjl7wnZcUf0QsEAcaMOYCF7yVaiXJz25dZ9XE8r+cl7E7C+Z0o
edhCztWgSiyuRnT0wQjurIZ3JLJkZMHqqkdigpr0dnKc3UQybMn+BaeOoEZDGmSXt1l+TNxh0O9v
fvlECKz3pRn2e4k2c1pDkwIGJ7xpDDRG4qJO4rYXILQkEZ0PYwPqR0TWxui7IVGzwytDmV9SO8Z/
c3rvwx0v2U9CakbTVxH+TrBIsvODMjc+h/d1luAIHBkgc7m+AzwwSO412C1lLi+xOh/6syf/o+3e
J15v9vA2Oap+BPPWsg8p9k4STINP66jRgcGnLrjUHDhbwADUihjzubEjRHImtDu+v0gXIcWvJ6ev
3d4it5m+gfh1IPmMy9JTxxiuK7bCGMq/LWAiiuUYYlX0lDnqSvaJs2F/kfLPmugOoGGU+w0scev5
MJa4GlFyu8VUev+TrJK2YhW/JfpzzetOuTp/650U0hCNvhjxKIeuDlF64eESG7jahbjlGvTAi4vI
vuz0GEvoAwC+aDoA5OiJDmf0w2+DWHKVPJEr8NXgU5gHM5vVN7TCkrQ8/N4eyZY4gEpX7Cyq73Ol
sxseZ2dFP2m2XDm4khGP3LXL8u2XGOmmUmCocft/l68vkaPUJLp3z9xJvwiv5nolzWlykviMeSDo
N/z34WeaJh1k6AcmaRJ57GWsrxCVu2OXXckHr+na/4FNcpE2PDPAI27bCvH2xA7EnTtMvGdex7fJ
UGMwhBnJ9uzHmgdn/slUD8G/uYL9FuHPNoaR4hYuUVYXK2oVRJA/m2OGKMOrdKY26/WLVUw6fQpd
fZcZYD5zWpih99cuhmuby82HmodHExqWTn0sX3v7Fa8B3dhk7tEQ1/DPqWlJpskPFzVn8jrqohUm
FLtLs/Fk0jbyYnAFGMtXE/GEUgAoHtB4y68sk4ZSt1HyjhFMiguTrd8N8gAP2jd1MmQ1vsGDNaQV
Po3eVOj/X9HF34ujQ0aWIS215Eq6A9u2eJhptA3YqYKH551cnPcsa7M4NuC2ixfbFJGv3MLDTyJU
wB9NvB7tD0httV2QoNwUs07TOh3ZMVIqa+5BFgpX7w3pCJQDsgZNJicGQg3h+6yOjJb9sDVBvW8Y
RZcU4XEf+RN67xscz4TOncBVp68yk1NNg0JC3RZlfLFTEh6LmJqw2jxnKvwok1pfIGonboiYp+bk
WVSJxOPWbR3Y3ExeC6MKXVVnPY38pI/rYkDIzpf8rnsjyaf3Z0w4SIHzTpfaNWKdlVuJnwjMAdmS
Q8/rXiIqPeRu73tW+vS/e4/DOAk6VbFWHcadBmQDxv+OM3Fi5W1HavEdnoKo3uI/xx6kDkJyTbgx
c+AulCGLTzry8moG3BG1oBJulJiWKC5neA9fWQcf2cqnH9qaqElJF88gD/MRE9haE0lD/5bdHG6e
watO9uNKm+deGF4YJAFkSSjhi28g7a80CJ3zF5tEpBxogJJhStbF87pTKj8fVQNavZmgnaMx89mZ
GI9Ir9TZ5pbFZbX3D61+3U7SHcbuA3+iB34ItfZxjtAFkKlaAfISyuvGAfSWoA571fTBgpbWcgB3
J3qqFnE0rXV844CAmqTUCigyEFIL+Nln/GNm/h/DFCTiPy93Rr0sZDXlP9TYNnGmXotwmDqHRrcn
W19BIW9UjhbBFSIXDsQIF2OMazhRl/0LjsIqUFfke7EdbgEDvkpkAegYeJsRJh+IVINf9VbFjhY8
oCSWxcc2lUyHPCgZa3L2tfIeJmBeYvzBBn4TkjNWW0h2kS/fwzqyjbi53SkMyLm7yyF/BEb5kqk4
pSUpBc/H1NOXYTR2GmGGHFzu3dOStbdIjJ38FHOvEFX6bfEVL5/bwfrubu+npQCW2evFoJOXQJ83
8fxRdQVyj5ND1H6Ldq9ASVgAa+CZc+WtMYBwghy2o6Zmw7FLY89ek2F+rfhyjSGvd4U7+niiITMs
uqjFtqwMWOGjzeKYqqwkSkDMtRwnq8S1x3VjOwJp5KOmemkz64DKY9RG8byedelbZafUES1XKyZI
kUK2AoybkmuOWiL3rxZ9Tff6ulLIpQd694p87+nUqWbOCXdeytf9NdwgXGqMqZ4VB6cpZqMIe/tI
2GjbvR+1ac7UqRqKOWRKdi7T2ZpuPD/xTwKtxku9HbAf9DvoTa4NB2rC8+qKSMaQeOAHCR8GGnkm
Z3OvF0U8Ef8sSNjFILTr7kUuZgMHPU3Z8ENmDFd4G/GmSn2kAs22b7HfCt4SNwFNMlDAO/oqa6NQ
0f4iF5A25NA1GpWkSoIAR05ISWjmyCkavr/TTy4Zf4d/DuSBQX5B+67uuhdCaBLM3J0qa6vcmVWB
9F0b55wJYJZLIBNAr3oBB+2o2R1rou9u/UqeMtBk7JZo6tyZsSsA/thcAvYrFj3C3sUe5aoEDqh4
XQs0zyi07cO1JmvDRy4JP0DORo8W7SjGuhrPxb6SH6H/Lcq7iSE4NL9IqkWGIH3WY2BR9V+aq6uV
bQGoXZ3hNVSpRhnKVRgv7p+lEl5zeYUsmrBZbniMlsly8gs2ynu5b6sRfuaRNXKPsGiRQLVwCji6
K2RxWUSrqRozZfhmbx2Y+Ya7kAgx9ExyESdqvcZt58EksU40ovum7ypDP0KqwLkJcoVO1Xleogvb
2rKH65A9tJCYafqA0EntKb3aKnIUkuE8sW2rujw4BFarlY4Fm5Mt8jdZkQSJfTeHscXEKO3pn4rD
Tcsg/H464GqUhqzaf/uBUdcsz2F/echhEko6A7f6YZt13K2Nc/dxt+KHyVndOd/Ic82+KJJ0DEvJ
2yvPfpHZvyL8ZVQQs6LPXlKH9GjSUAYAbw73EQB78+qU2OrDIgXWrp+92+Qef+PDyPjtg21NIcXN
zFnRb+a3tNKdjKG7rYZW6dMVS6o6X3YNdsh8omKC6oLn7rOrjmRp3HJxRyyTeBZgG/CDhgZGP2Fo
8ygKKbdvrhqnYna7Ir4rySi9AnB1njmuIJtK/1r/up6ho6Z0jsjT1Ha3BKAmJFIzkgVNJ1MvPdBO
NtN732X+UKah67F9HczwNHNhBt9l2/7/bf7xFQGQNUlyaNj4lkcvJio4F4V6EyHjhBgV8Lue1IYS
GK/nTDX/WjW0yQOBbO26lhbdWjfwQ/HrpDKUn5Luwew2d6FJ0s3dymDOQERpyKxUELalX152ShjW
7bNsKoDjDcUU2gqGF/VZznS1bn5WQ3JtAT5t7aDR1aJmbvTMX3qfb0Mw+2RtDThpVBUYeEgJ5y9G
nq8GrojOL3++9ClASmcd1DyfX7oqSX3S86ieaaPLSIkyl3/oB5vzRh/MnC4rxNDtrwsOl8QyNWtw
cGfAkcBp6XxAIf92F5/JuvLbo8Fb6UukL1PJRX5qIlBwoVvhCM35JpqkB7Af4GNRRMVDCFWL57/v
k9MGySpvocYksy29k5lKrlygULkZOICTolU4uzQlDI4dyCc74vaP1TT0rZsl8ivUvGLpeAsW1jsb
ihwOXgVy3Xneabjo/j43slozulkwY+WxLcUTz1wexn0igod5Y5cYkc4P5d2N1O8kcN3Wj7Z8LPjH
4ac91exIeFnPIfcWXKmareVDoWWTkB7xlPNhNo/jMjsob+EqI8yOdh3Fj141auhn3q70Mx0PTzyU
ar8r4P/Q8mrpAek/svLqL2a6E0lNM993EcXwyMucXJFrkDz9Kc89eynEj4GXC0iBTIpVurdAcz8x
nlvteMY2h81D0o622CHa1kkHH7L9zhDP5IDL4As5JlpI+nG7XhS5Y5BMgwqfK814CIrOiLdj5eZY
fFRXuBSVWD7nsWWnH7XXAYKLZQXfgsG2QeFgjoiLoGWfkMqIv2eladRejgixDGRnttTOwNNtCnNS
Av6qjyFwuNfTEvMzxy1+ozXXjb0Y/Und2kVzXSwL052du819kgDCVDqIurQ/UApjxPc6yhgJk/JL
aZhFWi78iAVskmX9IWJDEEGWk1ccF7cTxggKJWJcZSjTVLysidV/1sq5FM6JDnritNxMyY3XqovB
EGBIGlcoIY4CTuX594rw+qludih95I09poSu4IHQkWarF0T3LMtZDMXc9kF6wGrY43Akv4Cjw2Vz
kjxZIi6AzulT0HyV75/li5WcJeFmd3NaS6jTwGriyXxtRZBJb8nsqAdzd5WDW4Tfg3dp/JdkdgBd
i4ufDuJuhNdpB9M9gnRrO2P0m4hRA5Jw9bzSjXSp0rKqTjsbbPizktz89kmL3YbvJYqPH7ZVCr4n
3odF+GWvtBJ0vs1E9D4pOl3rrGTJVEVSRaxszSY2ybFhIvnJ8jcjVqZU2/eixpAGekiAekPOYZoL
yYk1tNYcK6k/9ByMxWZN7djG1gNQbmv2rmgwqJ/oqXvD+7DGXsnB7dlvAt6VAdHj+e8nAzzG+Gn+
qpP9Uq3giBSbwBz33h363DBwQ6HmufodFtPakHLDhThKZbDvJWVwLT1fuXurjJ0oAbE4oRg6B5gI
o+TFV+euOfLnDkywcdbHeiahlIuFZftU1XuvgPmCzfyhzRQUkDGLqZf9xIDF/3em0MfT/SVEEqC+
3y4q/E0Ihk4iIr8Q/AoTvd87u5wl2ZvlgU913BXBA1h/ld47ZjqkPC1fsX16MjhPNfrYIb9Cp4Vn
GW0b7Z1VM25F9B+a+P/SQmLtlF01RdbKWvubaA0Yh66KsoK4gqyCpAQIVqNd1VXUOvAp3xEo6LuW
6zumVmMMiA91ARGGdJUjZb2tbya0KxTH7L8ore2l+2dqBUOo107+tDXsTB+dMtJGOJCGPTfNTFyK
fd8ADiCqNN1I0JXBF+14LRXjvaf+WzsCL2hO5hpOM1mxwDAjpew/t6iovbN+JmjSWuZkhA+/gEEQ
2uM1fViSQIFvhPUo3pp0yCMB92b/TlsWOj1grnyE3VJs20H+j6pF6SYQbFxS3/EaXpqpCqO8CXZC
lwne7B+uiWvZAryx73uyXV9W+tOISakubYkl1c3IgC6rIROwbrXBiWbzsQ9RXcjZN3w+G3TbE67L
sodH2Kdqm/eQoWcSwuaJl5eiMxFO7YVL7ztpzjMYa0YgFTdU9/F7gTU6NPSRzzDqtuEsZjkS4WrZ
HdoppZoCCn/clNubIV6V38616vTrU8u2R4jYx485F0LxwKOdC9r3V2hCWHscskx1E5+CHUJZJ1EN
V7CnfKzJUUUopz3kcoHp0EbInFJEWd0NMnpyYjiiC2j+/yV27z3IEkMSaAXl/XJm/mE35B0LpJs8
LGt9yX/udXc6tsks2mE1zvb6UK6UfrjaL13jERtlwqHOccTUeEQfoGIRiC3vfpmtuVj9A3+IsSin
q+7+lRrgLvUxSRkYHsfB96+kMuHbKZaq2tmGR3/7G27pJt3dxbT4ksc06F/a8LZjVdfF3iXmLlhl
aeHACaGH5vX9gw/d56pXYUruIA+QxrPYCXilP3VkBejn3nY/sMohJcEabdO4Myq0qHiwHqYwndCT
x5sFKTAAsP0Y4h2loVrCKLYaYMRgq04Qt1MhQsC74oKWpLf1hZAsBR5vptdo3T8VOySWhAL+esu0
VdfQPB+ohNtHBNLgcQF7jjQvCOlcDSWvoptV4oNXbaDpQa+zcEvR3KOjboxMfYjLelifZfXnzLml
bHUEx9CS5GpM9CfiwqDNDzFZGaU3tzcEGXjG90IW/X9NvlZzSMnVeEyjGxIhRZr3V0TBhrnOlnWl
eUbvAjRk1uK3+QK15dlpwbPpiMeun4KnTE0Jr+yhLwDuU2iVg/pg6Fgo4TF5f1sVvXTpV0AIx6CH
F4O+TOmBAKGfWaF6tE/LZbofdGyXSHpti6mbViS8lgt8PtWvgNZ0+jbrf9nUCPzYVIzJu+ENvZQ+
BUwxSwU9axbJvK4seVHdHzm/dlWJPxzzq1RCHzUQh0RpPauLBV8W0VvK2mhOKGsYsSZGmjhijZNt
pnXCi4kQA6/olVaVUt6qHQpZ6M7tZwwS+paYQssavf0QFKOL6o0F8/ZqcrRzd+mXNqWvu9KZ1qhk
nwinOyiI2/cuDA1neHOUjv9slviG5Hrmqxbg6Z4tJhXgB6Ms7zR4sUfDPonem00UqIdGEe0ItTfE
4T1Gb8EwVHDHjJ7MvznbKLjuET5MptUT3SPp3tgIOUDJHuswLQNztHCN5UPWQdinSbl25oYevwzH
FqPU3d6loQ//dXq/Gl6r0nPGo8FNZ6x3txkfj+nkWhR/2m/+GG2QK5jquBbG/Fo+dRpAL5123Z65
j3oNDSmhuFK3SWm/d5D0IlZlYoCwzUyk+GXh1uyawOm7YkUYbMoO+rESHRFv8AURKIqXcFysyK9j
zU51GkRj7MmLEHE2+tiLHgZWByGC+oAJVxlkbfBq+jaePviBSR8Bxbl41eTs7JoKe0C2Cl5M3na0
G1QuoG4JJbsRjC6pngULB+h576GPZtjojnigIX9UNd+HXvoZiUOsNPnCnPKUHsMVfw8eLpq2rKrS
QL/JtlMzEhqICuovY/Njd+QMPcd2l8vY6BMTbBpt1aOGxQh+LxVi2UQvGGaEc6caGQUy+bBpTDog
1tIkC9J6ALQ/IW9rpUErNKLK3sYQVKk2mdixqjGN37T/FtflNGDC9jAacFTKXYIxtAYXeTZOOPRE
Fdxx9fxpNKaY9QLdZsCFZFXoN2eWVeqvKhq7vMAuIeeuxQvvl8UbpbNJyXKDRqEfD5V9EcnFSqNH
qY7/tPNvyfu9E8RA/I7T0k7MG+pW9dNjai0zd5TD/yk1EM7G/XDbcvynAbhS3YnWMQzVezj18Jf2
mzghhHAbSCfENRTjlg/Gk+S61jOqn4zmt5s/C4Zgeeiqk9rtywI23c0+E42mCqandkeHY4cxEDIJ
zlHXp+lyzBpFyozGmJ9zZ9+QSF9iqFLRJ8+HrmShUdZu13XIsonsh2t0v6wPAXc6oJ9wh04w9AX1
rb2Zz57yjm9YFAyDGD49kHGKXZ0aA6+OA652JcXbEprCzpICfWJ4/u5M23/cRh2yip9Ni9w3j8Qw
NOMdBMIWO43XFk+lvCJy8wFqudMsLx0IM56MPl8QVZD3IKqBlJxQ+YLCNLBjZJAHckXTg1uyq78D
8u1k0ty5jZmhMdRzUTMvERVZXnQWO9Lp1JWKGAe+O5uFd1nepznT6RshVoDpLtazTzNeBj+mejSj
Rcoq9/lVmSgOr05jF5/IbT3/kMKYDlYKqE3xQ9LnAh0qIHE0zfMggSPhkMw+wbz+WHC0+JNmejMT
up0NEJ4L+A7WyBEw1sJRqm2XYciQXttXm8Bvqnea4/07YcLuYv5uqoG3d/WUTHH99+p47qE0KIpY
6ZHtxQl6xhUZs652w3AqzQR1rIFftegBSnAozcESP3TvUCXqvfzkIBLWZwWclGSWx+do8zR0IIto
B0dP/1Ej6sRQ1WjTLY0HEnsftF3I6MZvMGRSrC3NATgVPex7telbqPpAHQJt+885diaWvq50TUXh
csdHu0qaqRCeR0Cvsybn3g9NxK61UF1abVlEjzWm7LE71fGWJOuQaS1bfpf8G02qxAjlPRDDhatm
bAgrNAH94jP+YN1NkKbVnFk2viI89Q74PvjjUDDXWlznEZCs3j37OOAjAw4qRa7IvPOsXBoXAh2J
6QjkRdsbaVUumnFmSzlLCwD6EqNPx3hJLfcm5oFZbqxGAlk8bcNk8A8hKaSzvRYhMoffGU7/SATn
akJkHVHPYpIBgJ97zYSc9kWCRdS40IOPlOtX+93KxpesinG3iL6LnbZRsCuaF2CcpQCQvXOTgwAI
1WtNMIJ/SqO3xkAwKSdeOqURyIXwYiWKq6lua10KA5q6lTRb84CBz5VQs/HJdLc3NHDvrX2i+Zwv
RWOm41XBezI4tvZRRBBCKfifHC/HjxS019a7J4BjGNYY9HZ8AO5NmAZyau0Nu8zWg1Yq5nPHaoCD
AEc8j0YbLLfwcWEcKCCH8X4hJYlAAyTVrjO0FhG3zUInFsOwdekxQoyWiorwZa24pZwaB/bYtSGs
e/ingpQG7+4a5UhgSvv0hmGdX+luD7mzMH1aeUABb0O4K9O+jpM3yrspc7bS8xHVLlo+OIbAd7mM
Qgwe5iSOKXeOJ4NP91CqC3uFx4VR2S7USYW5/GCLPgd/mhxm5iG4LX5vIng59C4wIaUW5SmlBs/6
2hPlouJ3c82nH3cnFvQzg7VNu0fE7SG+LrkMRPWDM3Eza0RPaAXWd2KiHplQTl+kWtD1mGHJAr49
WZzMA54T9gqNoVV05qco/yCskPqCDI5Qv8tl655Zzs5s9ueLTjzrZaIdxv2p8w8htdrk7BeijXPE
BOH2eEVmmcrb5ATVX5aiMBS9DUI3T6IqclN3g2TnHAjjRXvEK4hr+w/44Wd/pFDwgmS1Mp4+xPck
a3+diHz40QwLbFMJoephsBtMZyAMQrf5WEq7HY7vzRkRn2wzaHwQQrYuIi1uGLJzCBI/1hhUrBVd
esiYLjO2YHb8yO4HMJN2OHOj5J9H3RZj5Xsb9pD7UrlFzRpb7yt9tSpyNgs2nzdh4zUQJJynJ1Yl
FyJnfWAAm9kslBXZ9pO9KLh8hmCaCnOUqtFFFhcAV0fTyxUAl5e183gDWB7l8jyh71QGcdzfRSTn
A33fA9SAJ95I5cn1j8Z01tPlw6pThhoZURNHyTfw/ECCFDdzfKn0bXuXo0P4KMHvlphuFBGlnFtA
7mEYlSZ2p8XS/SFS9dVN+MDakddyZvbjyRo6Pm4vRgp9u0cSNwzVO5tOf9L6uQaRnWyw4n1EenMM
q4r8QA6iLEAlaO2DJl6ocGIpRoeXslz303w6bvvKVKbXyMJXtuiBhrWa6scYzzkQkrd8tFsoh9zP
9lP54lgCeSSEslh2anyfjS0OC3ka/ouj/2GaGnuUn3p30x/UXFiDicGG1gcjB0vNZuurM02m0PrF
9LCFBkojgK/c67C01exp3d+pxVEfScVuOE1QCeCRPDSpX1d/UnatNOy/0U0G5nH0hy8j94IUoMnw
fCaggZRSK6VvOnwWbrnt2GcJqGrCtb6NKEFF04kbIIvwZXPpUDx1TU6bQJfNmtTVN0DbHaV7GPLo
eUhyJMnNFddBo0ctR4KRnawApOp9k/shEUed966DvgJqgU2LC8iaKeeTUhSwNy76MBma5uUq4LoT
lSm5TBkCHOSIjfsi6dlILJ1oQlLyBRms0aQdonFClR80Uqev0n0YAsN3NwQLmKkQUzoIDRbPL3cZ
CVWp/xW4zHDwoUjQyfBhANsx0Y0A51dcfdpm0jv8ckbWILJPN7U34KWxyXsZHFtMDoJCd3lszgfn
kcDqrNZa9WtufskdovNXqU20WtPn3nNGIl8A6LBhC8uabIj6diGSMV3NuybqgTFsVI7Dgq+0zmaQ
og0FlYM0udt7QvFiqmx8VPCBOs+zPm+bbeN68ZMd14LJEGRTOsExlRmXOMYsEv7n8m31N4kAnEIP
qRzg2+eNXnLCs61jAlZrS66eJiNN2RaMZpLTEFg4OTPqECAsNSPqTfwQRN5FzcbbpkYLqs3nPR+F
sxNkFJUnwsefUL5EVa66DIMSBWr3Al6p2Nt0VjKOd7HC7j4sKIu9VW5GEi8C0LKMTKbjfaNUHFg5
fvV8Yw6uTjZHhq3SX9mD9/+eVQuD/kCZpT+f0gcSzAC0vwA1MWfs76EGhadf9QMmes22jmEiawFc
6vMEudhMRsLSrFi91FWiTDBDQAs/UMeiVjl4laAVXS9IfqMG5YszKnTU+JbOLE0vmlGPBfKt/SpQ
EuNx1/Fr56GnuH4QpwhHIjli7kVqEKZl1wKg1cdehAopm6wtN8oxjSC9p5SCm/9q3PCT40otA+y4
02DLMPegZ8I4NJc2om7mp9J0xczIq/6Zgrvyr6Me9LtkDoorv2fyLqlqzBNVHYLQXJdGqDorz6zw
7wDTM+c87XQOlvcrbBjI8HHCKjpUhfKOEtuM4OTrPEZefLAo5flQk//1kBaN6Z0CxfsDCgeJyb67
xb7/puNladn/yUz8RR9L4KpwuNj24PifPGubQ+RLlft9GtP29hhw93nIZOETyu6sKELCpQTDZ5dS
hSaPQ4jaJf30+TeVtQsGgvpKtNw0lkzTEFAqVXgqg7k8LGdEUtxIO57MPqn3miRvicU7ZEViF6DP
cF1WX9dbHbz3SBIn69TRVk14dcUYLqzKNaF0DQIMsYHYjtGQW5p61OSC31OsYgxlcvHeQHNt5cUm
JKda3kc02R0ECE/vnw1mBUX0xQEaWuVRLKUKGQECB6euYglimN4+P7m6WH/yE7dE/UR+l55/GWVo
HUuSQ6koSzK15Bsoliyf70W8ce5y8GycUbjxOpp7igiJrbC7ialU5TDNJTi3bJGYaV5Arx/AVTfv
EUMAHKTWK5hbukPgUDAlOh2283/6J5sqZg/mKnxUQDcVCCzG8FvP37XJ1zyfSg53eKfYyiJBIfHl
DE/u+qjhP0BWN7DJQ5PILoIAtpnWOvKu88ENCcGwdN80+avqG7I1gxJ/nOUAK0fYomB0rjj2KPT4
MTw+ktiMzvtOL7N2SvUmrOPd83Nqr/LSL53xgTN81lFXjrGR3E4RWb00WfY0wq3Xn34lexUEQ07B
BiIa4Bz/Eau4qIBC/PVk1t9VZEDLfY2nJvGD+Z0uLVLcWkoMZhHuOjwI+rgD9GORHRCo9rWqYd9F
XCzMF8eKmejfs5fDtPp8kS5jxK4MIF4cDNueW8+e38p3eEf7J0K0EqH3hJaTRY8VPj4vY4m/FV4p
1jblKxsTramrsRTQL2tCLUT8jOTs/K6lItIw0tIF53uxOh0BqmZQhIj5Vw7e24X+jC9uyY8wwCSb
XpuF6mDelqPU++nkv0eov9ibHxJ9Ib2rdJlSd4ivmJjuPMpeWXfQfpZ1g1eD4CY44Qgjdots8DPg
rEhi6YduF8Wxy8xqIt4hBuCRr1pVpfC6YSMcPPagBJL6tmSBAYFaLicps7980o5BQcrPPVEi+MrW
X2rnUA/4WPdElBJLuSD7f7/p5sOppIRv9NaNWYwPyGs1uEY0+tyYtQAXja7lawrK02gExGFJ0XZt
mpAcirs3ZqLyx+gpU5aE8GV+nMkhe/iZsFnywY+NM89Gpws8z9MqpyNw9LuKBhKj2ZujAn7y6EGF
odaARfbXSXXWqaqxjKMljRCWOQ9C6CBupRU+bHMTB7zrWWyuLUThdFZkZbgVlHFmi5mRPB4zgC5N
lh8SjWK2g+q2gJw/T1h9SFpManIq3L60SYjBbEqKi36eAjNyHarH+hiHVKCm/yH0Z/wpdK95QzVp
X3rBJGAc2NelXxll4NgEiRTuYKaWKgqNRBynD9kJf1K5ATGGIeAQggmHoGrFuhVMHEGzMcI5kHu9
XRMyd7pgEaA9zI6oSopjlkgawN/huEDxnKxg5XDdd6GXkXh1cqii78RYakGZfpKvTii96SXYWcWG
q/9GEP7Jz0unEzjTikaI4g0D2su2gSt8vQuNRFuU9ft1f1cFrZz/hD2zSnQmcN4DVOO3FQFCVp3d
mgRvKaxC0gKaiTq9pMBCx6OUR61T1yfzM9Zdp7+C2Sz+bDCH0YIaFUaAAckDeZTbiRoLVx5d4342
XWxwYmdt+zfkqZiYOC9/Y7EFhA+RCrhC61KZCF4ttLw6oBju3B9otmVam5BR1vy9kcuSz6Em9J07
gjSfxKFxiMqsE/Oo3605kdGJZiKP5cxO1LwZ7M1cAB4wa5Q7qw7NmMb2UFTu1hhpUpSg/w7OtzfM
5/gsoB56TAOYBHWlsEj2/lf0MAa//KZwoIqs33QiRBqbJdYIdu/wWzKTv9/6gN9zCkflgrKzjJDw
zuV9Fg6Q9f89vBf3fbQJZTYIlcZKKMmdJ+rznqfuWvn+wZ6ANG4o3R53U/u3l8fRNhz2WyDsG+6G
pVf3d/klKwgZTT/lNQhtsK9fzJD08buGSyptpfcnpRCC2CNvCY5B2SxoHHo9JnUAiobxMXNQKHCc
3US/zY9ES6QxIvCm3TLc7q7fQL8Lm2n0VNL0OsdpyYQyHbE0RFXbLOIVbWeW2HfNHkwBgKLUfr7o
94Me5CA9KnKXKAlR4oH2nuuubkqK9/3YYz0NFuutvW2rzcnk/4t9N5It+hLaQHV4EJRGp0+7RKUg
5XEVZR53Ob8Vs/DicojGq/u4M5OijdgOIRE6zjJEQbwMd/NBaUEkV0C39jopbby1PQHTQFi7Z1HJ
sH6gCRkvZnFYIuFz998ERX4rIm8d1WzZh6G2g5r8TCKb04H4CMv8R2Ed+aAmz2dh/Pvmkrnf7Wch
qVDiU1xYXbiBvfsGNpbychLr4DzUDRHxO3TklkMNzU/SJaMR3xHNRuv00xRgI+bhpJWsjY1swcQV
m1aeZv/aogNCrttuB1fkMvYr8ehe1im8tgjgBz/0utq+ihhs2kTwNcPQ9LTdovbV8Q6KhtU0l82W
W9S+qMyNHaTDFPO+fwzRViCjz+5GP6WW+OH5MU4eSFMY1jIGKBEeChcv/Y4mvrM0ZEHJj2vTYZxR
GbV6fWnEywmpLV2oBTldbQ9wLcu+o8j0UBfme+QFI+N8pMmgHXq1UZKZhgoo46hqtS8QvGIjMD1M
BxjWdjHnPFnr3B5Eszi9WKeDH3WCRMZJha3USyes1dpXHSd1iqtRr+p2jEtVRlP64k9EbDjT5lNd
2+yx3DSVaibNeQSWLCQdKtd0jJmftO8FiQWWzHhgK8rD4F4jUXAvzilHpuuqx7BW2zbxfiRFkGc0
qnMNc44bPe5KZRSFVRZm6Rl2kSoaTYAxCGBeY7vHN5pr8IuPbn/Ny8pQ44xM93AmwhRrOc5BeZxv
eMR2ggR23k1UYuAtdF7xwQU+1ArPHV/FBRq86GY/Yi/7cAIG/ZhcxFldGmkLm6zx1JZpNUaGMzmX
zIwlWCfMRxB/RAGk4mlcVDpT76ASec/c7dOSQG2vjJDl4z691iW7VrP+kIj4A58ULBJsS+bjUf7S
xlbh2gbLnuA+/5owfpNZPkMKM1ki7lQeiGIp61IgpAQT6dXA6CrCTgvSsFA/nfAa6vvjUrYY+2Pz
eIf9/OYoCuJJfHvvpmmajgYLoaAsX65Kj+BgzGyTCcMeeIILhcCANkaghEXKXSTHsRI3WPidYCuy
8QcnphroyJw5GCJRF+9AZAo2RPbf4+sOXxMbmOWhHui7dKoFquTMeovniaaN92Mlc9l1dA/dceez
HloTFVzM1QXjwgl6RC6mRGjsNhx5hO0qJHgycIk7NF84cI3MKyCKQy7Ya1lkuhLlxxOLDKFZdSx1
ej2ofyzHLgf8bbTKFod1ihYqomc38/UpjeHeyNAc58qj12JprLbFUBQQjk3W56abjN0A6NG2wyUg
b7k4b23M3PiqY8d3gpTMCuv6zs0fq0uu+kW38dBvtER6zW7b/eRYfriwe0+qVJ3KFsAQBzDRQaFs
Dq5YwT84TqWUZiDjBMqMktpJ0pG6L1crRDqU+Za+LiuheOBn78kRDkRIVSoZHzAALlMTD4wqf88w
KpW6w5C5U1vMpqWaFrOAaYz33inVCumH7r+bcpJSXcBIxN4TFpEGe8hBUO5c+yTDwRx4+HVj5yyo
MTLdgpgb6m3zT92+VZbTEo4QLMIdJCY311r0tzj1f8j5DJBWFli2cjuxkkXRBWB2c9x10SyijNmC
sQrMczFJQX4Ox0pMrqYtzrco6JHL06oAeCeU9RAhxzeBIxiJzZq2gR+YqhfkEWfHzKJregr8YTxs
W1ZCkYg1tF1bFO6x5bYPjZhL+krp/sHudAcY81kpqPbg4maMeCpRdVBsadrNC03eCkeH0UEqB3RU
vJCs2rerD53eMCryYuREZ/UUHocvDYOh/+juy73LMr2Y+rRz+DyaKSsAShU231Fs229YJTO+d/1J
HNglMWcA2Dr1s2KF7U1TbTMJeLWz57Sqfg9tak3Hyyloj9dTbnoWuidRN4ZyX0QuYAi2YwcRKh8y
z0MJcYcaygxtXAy3Tvu75StZnnrIsBFIG/GwY8+vT7EFIbKEJGt2YtanTJvEmLPnYwVx1Hqt8NMG
+kLYLkCdjqnhCooQrwSE7U9VSCrYSQBlj625B59rV1pvukXGIZ3jWv/YKQEi7nYb4Z1Xk9Fnfv80
jrsTp7BHYBMgMhTNleDZjale9EyzImiKL6rc1L47lTsRcGLoOmd51mQcVOlZr53+zJMJN5haS7kf
teUB67Hx9wC26BkWiA4cDkBM8XW2nQly5WrEfqaIbpemr5qAkvBXIlFJUwgbNHGdib80TYOCzLtX
7mSQEVZjmptHwbxoYxd8OrwNO/rr630mYdjsvIlcuHdugGpiljcQBBvv3vxuuIPC0zvx4kk1jfKE
q09THa3nM8Czu5Rj/By4V2M4hwFILppXaCJQg3yxeSswe52GsyjGRNB1tfabP2hVqPSnwNdFVsSR
jZQC4IMEJEfreL/QuG+SEFYBLAScdIOxd7qzA0IhhvlP3Vmfvbxt5otUk+fccvwmfAC0wsbjoMJs
hJYR37jnF2xrgJIQvZmq56hhxUS7ABbKRDhnt6Srk+zuMffAnjAZQ5J+YWK3jIRpvlemwVqP6H98
79D6G2yyyXrDuJSpZpr2JWEkh+EhxvqxiW84E8A8A4FsdKqUFqX2vQjIZAcv61KvNpHVwGhKQx10
sWVoc67E1nkHb4wzC1bwvL3GRl6ax4qOtOVCaMv3OhkQurPXWELqyokhvR6jROX4FiLkhttf1uZv
6KIXlUBFu74LuNShbVrQ5FkJZZB45j8EjFc95xv8mQ8XLr2NKq77px8Z4/McFvq4llXCGCPDHo1o
R8kntVduJWeAgK8pTBZ/tQaotC22H0e9BhDxQLGDBL7XylTZu3c2bcl8MiKOO17B+yYIqWZW/PvE
7xwix/7yDoKjIpi+YFme6rq+ti5V1mTlC3FIQHRVmBLbx6h/eXCS+vErLop1rHwlCdukqGGjpy/S
bzmCMno5XGZZsPO74Z/I+NeFPptk7frEBciGRMspTJ5Bg+reP+mC78YIKHPeEfbo70DPEAXt8jPL
Uozwc3IGvjMDso3srBB/zo2RTHOajAneYx+fe+4+uCdImUdcoQv5BS+GnV/w2LLGtO/kuM2ioih+
ShScIdTCk4Bsu8x2BV554op3R3Bgtlc84dEofTG5MBUwHLvCbtNJq9fMrMX3exmrE5e3Cn/kxBlu
EyyrlI9tisAfO4JKbBY4K6dCdy8tAvP81ZA4raiSlG+gP1woDGN0utN8AoN6o9fKtqPg5xVmVT3m
pjT9pBm16x7y2WzvPIU1rZGhjalrbtoPSnSKIR1JbgprC8Dy2cLESJrSJNXgA/VxndiE4Vfu3nUj
dhbe3hwYbpT6Gh/S7DanGyF5vLuAlrkyWA4hqlkKkATMERaf9OywNyXBPDoVV+BPlBkA+6XuGjCo
rZOb4NRNFYR8xidLkPmGgQI6U/TVrTGb3k36hYdRrga/YIgUiLcPED4gcIJ8rkdzvBJXkzoW+Oqb
gcYaKTAXY6j5fF98q8z2+EbFESGDRAZNOqfoQfR+vYytnmXfXAqOY8WDGPwHOmHefonB6rTp+z7i
BtWJcutZ1XfQ04mYM95Ex+pbNAgKulX6WVNcjkPWQBOSDzCHD5pXCa0Q7iCCmn0pU5hE1mMoN8tw
llkET79MMHPdmiNXrmdNxOZ9GWEX6qrWVCHIwPKjXai8IzDkKKdZ2/emXQc5Br4zzinLOoKW3vYy
K5pWL0BN/wkzSIlTipBjUOFShHU5HdZCk9QmvL5TMhWgMoeQ7SDLRD4x3ctgfqsLKNvw/i2gUOE0
6tr+dMyVpR8fnDPl625xmx3c9vl/J9Glke2vEzMpB/5zNNF3TqnIq6C0pt8gvZaSixGbdiUlhJ/p
GBZoFP8Oa8FEt7klIckc7c6/2nLRHhp1tTE5WxwXx+yNgrPJF0P3Gqc/BRB8U6sDStDfzBubV9qI
tESS4x+s7e6tjKLxZpivR38/KPDMErIVtVKyZfARfZgI4mWYGU7hTk9eHY7797xbMfKmNS4npfpt
uAKB0/uKCWl1xlQue5lFsFxhsuFv9UgigeN8LMhE4lZiLiGO+xdlyT/VgzN/Jk0NJhDZTNwNszV4
qI7/R6DLrEu0fIUru/abw0CWVllyBkrn/Ur6zOLVR+IanCQXs6VoWfNc2HoESxf59XY1O+qgwhQ0
JcCsOe2nNwl5dueB9IN1MXrMclMjXYliy3Mu+/38oR+5hPNfBiiMntQi6KWvbhA++gLTYrUtCPMg
UApQvGBgC2lQjv7dtjfzfsqCeJneG36ZZzSheaLV18hrhvKKk233vWt6143s9BpH3LzlQPYfuth9
NH7NjMllAZdZxkYCCs4/7KAQPLdZmg0+Ylhfc7FBv/9nu3sHW62xVZpFPeETydsEdvoMbJu1Zsfc
yoBJDHhvsIJiapwR7w+kbpOCJWKH6Cb9ykBJka3ozC+t3Fp+sTk78ESM5kjXaU50ze61n/OoibJj
XYKcHuBltecTKW12HJn9yB7/1tbBQ4Xa9WdVYjVHF9rNro/TMITwbpmqSpEHk3hbRBwf9RyAENLH
ccR7LN4Zdu0sUabvfwuyBjqGCaDQQA9sshPbpFJHBWFutVHpeeinlmRNxO/dASeKuAA9yRiB91vq
znRQC2Y0nu0dQQgAYTd/eEqORs+XtJg5AJfizVE2UzunZlw9TtbqQU/Had3fV+zzJdz9vS0Xw4Dm
iaDnXbCDbSK7WWTq9XML2Yw6dfVH1FygVh/nQG8q+5alfC5GhoAfm8ck7bvcC2SDoDnfW5UGkrjq
s4VZBaRMVBBUBuYsliGAgDqzy8kUcRdadgdAnV57D/1QwChHulXTZynzsqXWPhCGhxx2RKtxxZve
crU+nLsbIN5ngSYuCUFKRqn0qzYX3G45fR7G4zCWFHtYHXyc2HOVPghPl1Oo0WLxJE2biV0J13V6
E4DpuJn35kNtiAdyb9FqUeZurfevKLpIgwlqHxKQJsBb5PS0NAdDp2lZqimCRlN3xig+RPpUWIGw
yNqm3O9XpVomyER8/Blggw+4R1StwyPyT/yI9EImsE7jNT0JyUJoby21luBd3JmSdWfstWFoqVM5
3T5jmEtsgLew9he8vofIKff1Z3cKssuYrmSrrT9WB8cOAF6UloE8RohCVuxHfBv+qW3UkYFWZRxE
MGihPuozQLdKLiagwvcLqbLN+PC4PAKnASsnJD/Cz/mU5bbfXu467ozg7RKcT6WOxuAfg+1iLw0y
dD1cKqgkrTo0cm1pzUFqJ7R71tWLwXTaMJEbmSa+qpSjH+/2IJB6q1OPFyWdBUv7wI6ThI7poRiS
GLObYbw5032CYUwL3zTSMmOtZtwqiM4hTuj9x6dFAW4ExmUMR8Ig72bc1yXEmhJhk83wdrCyKTlL
PRSRJaRZBlbG61C1r2AbolxQWKoXDsEC6D5kkQGGNCuUlX9CJ34hy654ZGrp5ZKUTVK+yzHPz7ML
BWqSir5WD8UY99XqBaRQ7x8TavJgv3GnGyjRBOUcsr/I/FZvWD0PqbqD6hk1VbTUXCyQ1DfDNUuV
92tvQAeO2u2SeOX3MpTmi6k3tqBHzVMpYN7O82prunljq4aWIxe1o7/WV9EiK4QRkwJ397bzGNeG
i3fs2B7nTlepUrYF0LFZucD/2GfIlw6u7DJHZGiB6yTN/1NKUr5booiNecJUJHlWnFqrxawrFnoM
5yPD4jPPP+GLSJpzH83pJkXehaoE7KnEmF+ea2eIKfvu3zSsfcLd9lfFdoQA1TGz5xlqkn5RGnTW
o2UViReqli7EC+uA/i1RslETdvVEnyVTdUiIvbh6yBRr2Q6c7Nag7FFbp5oPrktqXWeKZpD19Exs
SjfBVTA+fZKUGyBALM4aANSNuTUFMXc7pnUi96wvwWl/w/Ag9bz5cVpQpS0AzfPqw/WYNOZ3C+QR
sDpWKlgXTRTTaUw5RDnr6x9oRHQo+zP36H1FFBMK3saTEN9OpIrDiyaj2Fx2GuRd3V/qvAQWUaND
/YNbN/cfGy1QB+PKmBi3kFEmeKHkWXOeU9z8rxeg1dkEjVn4WUBEEXJDL62Ml759DcJ2lS3F46g0
VZKNVdOsBkP5joDZDIa0uifKf6557xZifTdS0JWVneuXB4JgcVUEKw5+32tEDba9lhnT53i/3D9g
pF2HOTdYIFqcvRJBEulDz8wiUQA+65QlDDdLD5DQ9p5VJd2vHPC55txb1iWA6cZQvO0ewVpzIxG9
xuhe9rSkJavXWTUun/anhzeH5lswiQhsOMqoH2RYPMPtyV63Czdj6BewhmYe27sud35mW9gyFEII
cOUr3ZALGAr7mTEC/GeuULkZnaIk8O3tu2X0008aTnp0BzXp55TAVfLF42V49YhVLYcaTNraI1Bk
HADbefi4uFufLwwdPtcsJ19j9BZx58QM2mg4iGbPHVSMICjsE7HRnYnN0Yz2Ih5/N9Ti3P4t2vBN
hYLnyMLT8HxvxHdWckmaUiJRoe+5d5dJ/jDPZ41BmfbKA99Guf2XCuOLZSiqwFdVb1Vfc3MjhFBH
+K0gC7/jkyOE9DBnVoIYoLyif164a9C4T2AvKcAYHW6//MSwj/0MvKY6rhc4YeyTAwYC9QQPtzfa
fEK746id4c0nUI4oeIuXWfbEzm45wCN1AxZ8sOXK/Go4dEDMQsA/8LTqt/WJ4x/BUVeU9aDuqfN0
VD78fzaESJLp95IdoF0MRC/KlQddzTtPtRPOH6hOej+xk8tQQiIRr47Vi64Fw4M8SrvKnsXgIU0x
HtgB4i6X2q49cG3vJ7Y7ZB9DPILGIkB0+xs/wGFJCuF4GbINb9D8Rr/GqeO5ccPSzQi05BBDy/pv
JxIjaOIgDGfKTJAj4x/Aagn61SlOoZ48mIVbFct6WWnUR3PhOEOWkE39hMO1x39x0oV65m0Z5v6r
n2zfKvoaTgG5D8w3B+QUWL/dZzQqjf6qgd2NYVi1Po86RYr3eAHDnN66UUlJAw2AansAKXm94DTB
arfpPXz2ekL0kg+N1c3LxZkhJxe864zgCQhj8h2wWfeJjIebyJIiQWj+o17CarTrd3BelvreLkTU
u8vhThFAm1/X2aebhYai4/VHP0r0CbO3fuxm273SoGawIgWJvQV61EWSZbzwoK1976Zo5QwFLq7s
wxoUJvzzaY+VEeJNOGt5j1WfjG6tstXAsxWEiE9oMChO8X4OOtLMxYYyUxIoIc4F9bjA2HLp31t6
s/n3PRhyh5L0ooHxDtOs9yofAjilowAuwLk4njutMhaFg6I346E+rw9rYKqJDZu3m7ZPhAJLJa4A
tLm6esOA3sDgpdmubyY/9C81udCv3+XU03QBo6EdMlOAv8AQRwwnpSyOcHEIA1Dro7ab2qnjLYpa
Be0IYlZdEGFLvJ/qIe1T89/fOwQX0CoT1BoRVBJ9sld8iNH6yf5lFba1ZofGa3sonFg4YWvTJYiP
Cg+X2m+1qS+iizKii0W7PyevkoArnElu6DXMaSmY+I1jSjLAc0Qu9ltcPOdBZvqDUD2DkXvdWy4G
fBt4HsHWJULHR32g81zG1CHddLhcfQZL7pfIdQFewPxc30FN3QiALfksOJdtktN2vwSJ3GLCCTu7
MkpAZVoPPGXmpwBp2geI32f44Fc+KRSMkTnTGMP224RzoeC1J95jNdeESOZsHsZijrE/z1PDg0IO
NOef1OeONW4jgPkpn8Atfe+AQ/Hw/qD0SylLTHdRbihG1GNQ7MgxzGRQRfqoDDyZ5ylHCBzE7bFu
8crH/1fAvFfSLjWb8KFf/fjiWaYPzC4fM1GU5cNZ6XXi/2qHwMYkAI+aR8Cb/DgQzqtkS1I4S9Ho
Kka+K3zwznAbYS8ljM7dw74fzNUfPJfO5jKLG1CZsJNSB36pNmfLIY5Pvp6yl0iBwePibKojHMyv
o0f1cZUJDcjg1+E/eP5Yf5yOGQjLvEavntrzt7zSL33PTmpjxhWutwn1RB8Ockvx17kufmdgZ9yB
FnaBwzqYKltf7acSm1Al4gfSRAfxxxIW4FNQEi2GXYjkhoZScd70lU+JbqYQ3+xR1Fx4Nm8g7dFS
hvEgba6oCwFyNomgMwEXmyQFSAcj2CyrpBAJJeT0sUZBHoRV+HjvhXR1ag/BGQj2SEkHcRMqURaB
cYxsVWi31XdHsCERNjjym0ksUPcVsKcLC2YxjrJtBJASB5xRfETkmV9wQ55MQH33iqmTcYewvgLv
3BpIV6OdLRqBxtTZKzAUWEqjUPt2Z3ygPi6QvgoqAY/xYrSWAo4ESPVC93WG0oUqHv27qULQqb/a
CLiJn5bW8X14YGcz6TIiGQfzZADrpv50z8cOP7odiqN3qjZizQOMDW+++6VYXb9h+5GC67yWWPsu
RAN6wMh74qVrvh4mmRUWMz0/tOCRQCIXHIo2QkQMyMCyVOc2XvvAsVMkCqZR5d/usS8e7Kjk9017
MjHl5nzFCXJ6vZp/2gNgrPX1UTtQpv+pq1zr1kUplGdvCWGUHMwHfm8KdWYuHmTaFJ6LvLKRtoGK
y43TgvFtThAVVKe52BVawLKoTLJivEdWM9QlCuK5Vzt8HF5LEjy2Xqw3z63hFr8OChpv85g0FM8g
yTSZf6r+44JJ9oze73SF1wavIXUXfPAAgJMV6AjEUlIzMRKdzkbm9D/tG6o1OuCmENm8dZCgM+19
B8b9Eb4JzDKknGfvnwbhzJlwn5eqJGSRQDlFY0IF1hqdRvOkLFlkW13VvEc2+VFqrJvCoeuaRMlw
hXGzW6GdYwjMd0nwtthH3cBrolhtHCGXHdhfSLDYJi7WPjj2P6uVIRl5TLmkYjNl+oRs3qYyWkZ/
s78ZqZ5ARf0KN/LYSgqVUnDMT/kZsCIGrYyMQpu3ZU/VIhLfpIZNpON9zSIj0jAULsy5741ZyTZL
i8F7paV1P5Ka0fwVUwQ779jJkmmI65zmh8ZMVN0uYVIJ3U1aE08aFAbK+pwHyh5ekWn1xL2dTwCd
zlrMM4qaUs4IVBfTEtVByjTX2QJY7cCcoAZbOVUeUcol0StfhvRPnMds1Z8gC4TtzYzIhi7k+lVt
4b613LJiUDmlWPmjEJCMwCs3IFmwrF9A7i2HWzR7Oa0TrwxoHlApZhUlRxvKrRGTj/F+S4I0hH1Q
uBTd1lEfRqLdWggLfejL672AENZ8GZ73IO6Tyh0jv5O3CxKIQ4r6NUUCw3W94/bg4qB+HO+aluQU
XMzIXMKR0vch1Sz5FtyFAllRjkKQj1oCQiKXTPds9ioL1X+nH0CS76tGKbK5bl2PCvN7JNWIo7ab
hz3t9xU7PmyTC7BYfcRlyKTmrEUNgnGS3MmdvFs9MAG+CSeptTJ1XFISDuOrPqzrmPVYRBF2rSgb
WqLF6iwCg2ONxW2Kf0cKldAeji4NnBlDvtzoQP8cCaGgwba4ARdQtgDJXXijAkuOc2eU1AqJVy2a
QALaOdjrL/WJezdRawOS40e1rn+w5kUNM0CofNsdBeJxDubdeNJHvcgEii5ea1xKk3e98vNfMVNU
FM+S0npEFQpjXBDeNT8XnsJUvDljdQlbXAKyVPDVW1OBcyZIeFVE5l+c1LrPLW1mwhSMIwp17cxl
EkKsz4ZtrikAZLPYa/gPhKFBKD/41MK7VQjTWxji17lLAWTsORyALLDD4HQvobiXcDkMvbpApXyf
jhJlrCL5Zv6XPsyHo0KbZSSJHn0utD5xJkbaUnh5t5yA5UwRXbQoEMW6WWIEXFJhBN+OMNjUxo9M
DXpra8mJu4/W+aqBw8R5OrK1Q0I44wELCMmbCXh7lzJFmmqGLGpK1Pdd5LOED9+GsZ+kvVWHXJYf
Niqewznb68vUUm3+hwjLz60Ur6/dYuqjrxWGneAZwBdcnFQgg59/NFMt+g4P/kODhRdCXW9qR698
E3tXsnQrfO4JOEQeoPp5W1vnucnp/KG935MD96xYHFg+SGB5FPpRJCRhm87LAkN6fCN9Vp9j1bmM
ODtRi/OYbWXTfE7akUXlCSDYb7z8P38GU0umXYEO0BdgDuXwodBb7u5X20YDs43d+dvOVz2PacwE
4SpiMrr2VS++zLc51wbU903xktNAnLFPX8PcytZHL/Yv3FlodWWFZDuj4YsE0bwFCQhlKI1AhvMn
yZDrm51NPciI5+8PTDw1jDWQ/HSPB4l54ME2Tuzn17y2RrunmBaAFzJ3km8e9J3wojRC2zgY5JUa
GMZ8GEhPsyeXEeeAc+GTkoW63J+UY5JGworJ1lviByBgDAlWXvK6ytfyiHXFxQYitJYIJmV/ttuh
J6E4zdur9mgFScq+W8OXSByyP8ydA7cJvhZyCdBKj982lzrHoFYmplvoVvMOcvbryg2iWFiqWWrL
StsYC/Wx3GdfLJEFnQ1zNIGVZqmUsUu0ZFQECftMs1fLM56N9YjK98gMK6zNgql81deZFxK7p7s6
v7qGsBKIBDO471F9PhqmAgaqEjw7W+PM90g8en3TdyOPGFFuEr7tQvY+2YTxZ+qg0S6VICbmI7bT
PusCYdJ2WdiBWHXQp8lO9MngBySPWmGIdVcZdu8IIpzP/i4d/WVzBWbP0F7U3sJKEDiF0iWsf7PM
W1yfoMaRQg9zQWnV2FD9+A85R35a7RvAwga5lE18o5r6TZU/ratmvpsstlx1Dx8PqpVqmvPSu7HA
Jmf+ND3sGn5plT8ljyACK24ly4/L3uKrKCwrak5agtg0Jx+dOytltuZGZkv7ZHJnpOs2caEt/8qp
1HWqUtMa2L4xFbTFXdoz0dR2fWClhEQSNLddUn+vPBB78uv757pA0oceiPV/A7N9nUmUeydnGUrD
1XbTiRnFi4s0zQCZ0q32NA/YGkwIiM/VWSyNE1jIdGNwiTRzsncaqpZoRuEN29AjkgReO9IUYpJG
DOUM3wta0m8VhQcHTkFtYwe9G4laQeLRUNTJQi4wWMaME1BgM/55nN+/aFj0qguJtWGEA5ouXXZ+
1uFOiZKdH72p1CrcfI4n6vGL1u2ZAjkiAHS2yOTxNnkZ+9bXAqvB23MTQZyP2h23coItANPwOWjW
3kmEZZblA+KMfo51DYue4RSOIQG7NuCnzpsuLplgma2JEqSJOyho6XRbrUyv2RD3nDnsWFcvhV23
hylgdIwAV4SQ7lkH43VjgyFfQZR58HaxykEQ4oX49OdjyGlsLPhbuf9/etz29+CqZfJZ+eA/35fe
0riapl3/n+/D5P/caqlvNZDwdONv9I7/wOAdzctipsITmHKfEwI2pgkiaf/fLKsLahI8RkGvu5c6
xqRIbvwd4LIuSEJB7Q7IPDO/a0jIejeMyJ0/NxKXyUw2kYWGpUPwcktHGW1hP841qsodk3qjF484
V3a0lMeTOgdiuumpWJuPrqaq9EFXEpQAyKIRWDi90NgcY0lLPolgtCxA77UQ7iXBTLFrIaMsnrvB
ZEeumyYWQm4b7UtcwbSf/BUWk3jF6EZEgwH3U/4hu4SL0b9Hm9rA2HFETr51ed17Ji9FqV/m1tof
xHUd8vZoVgZuLcuu4SlblyzbPOCpAYJJyE9pmnGmpYyWlhbVf7SlkOGayNq4sqZ+jBoST1LA/yV9
WjNuTjjnmZ4W4rG1KWXVFydwTaygw+epO4JssHTQJyZng/x79Jtv0GcPSW15V0JiFdEd4yQ/0wfn
wm+RG3bAOCTK7Eht887VlxLTWgGE9pyLOfy0BxKbO3d/UtzIsa2rBzOOtVLC4m2PVdcl9tRPVgYe
3DGLkHrVDH6ewdw4g5e3cqLSOw5lXVkjH+8qbMLAnYXZt3MGXvag7Yirlmepn1+udB9xteD/AqWY
qyNzhZbCZMsJJ8BjHHJBa9uW02KVY4pM7/PP5qnQP2eVN9Ytc+iNQVSxVi62Kfa4CN/ZhHM32C1b
xs1iWlQ9SvAPaGEiuHDCoFLRPzLlRhIRTtXqqrft1eqCNPLem/3+rEEDP1C/EI6x5s79b7L6tojX
aAYTnADK5PmYqHZEbGgyy/iB1JxKgbfhCBcF+tTeyn+z0ylXk/z3YV0iiyMo9hXtkQCvJ5mWwV5+
FwvUWpBrZR59VYvkfrm8swF7We4U6RvnTYKGFiq9QwL7eHHStu2COa18HbBO1A1jK9DWf9twrCBy
MTi5o27WCRiJzt8+HEprIWFrdvyjV/euLKbMkD8Mg1YQ2UHwaH8yqOh0J+ZJhWO3SNWe8w448mNZ
diuLGPuCFkQWLWxqWfIAQGhmjK7q39M7EBL6mKaXbrqT5J5P0zCo8ISPYKH6LlpVjIdmubuenw54
BSdTwTVcYQdrMAM6SigBE05yjy2/ldYN7Vd6OEApaevZQ+Ev2wMoOpqZFQvcCWzaWkHXggX/7Yqp
XplX26zDsIADLkHgaWxxpZozp+v+bsPM2cilcfJbwrh26ASIicMa8Zyvrp1DWAVIcWv/wzTof3Z4
RyWbaqLwrxKJ3mEV6EQZYgoaC1YEFwvu33DktKFgPDCxkS1r0QUIYhYj6/Bg/vtNB3gxlj+DiMYY
Mjp78j89GSGtu8uGKDQ1ASQNZj5QafRo3izhRmW5p/91VfvwGar3cJcuWWYa1OdoUiPQ7CRlodym
EfZ55GQqoXeXLTOo9+LiAY6vN53VTO46a5ihwRtssf+15OzAPi9DKNg8ucUZqcNfMy3ZxA6rRsLQ
A4nR1qpEOMxXduuo5y4YyHZtNTD5D7+DzpsQiSjSMAI+oHyjvVsr0gEzzJLkoeRG3r8k21BcI5/n
YbJVYyxGKphHLWuoerhQo/d6tpYga4Zhv+4c5C19rkYLYEp/rPnqYH7v7eYCWnxh/HCKYYPqcQDt
W8nThVPlegiJChmtdD9ktYEi5L5mLAvYGgVa++8bhPy1UuzO2EQ3oLz0yuUlLVG9eAn6vh4Mg+3I
1RypxdACNrg64Z8FSislr3bXVu3U4SV3sc4dNrRZszXiB0BTHJVPaUNgqRUhlOKNKoOEUuOKs8zg
5OddP3JTksBewcCI6jD9UEneiwNcudNAHMxMciL1ZaJUrKpgDVr/R9bzUzhYLHDGbFYc0hDLscNB
/BdV0//pplrMJRYTnnw1Gj5JoZA/vUyz1YIn4NQmgTMH8tnR4cA7Zu7Z4qDvB6640jeDFpHpLmbw
brGFnSMvvFjacdJqwjiafoxk246UctVHwujWmD2yMtjjaC8Oaq5xdSw4BBt6k+S2VGVhFP0gavD1
7k6GJD3hdvFwD0CIGuz2ddExSia1oUI9hfMGjqEP5YvSlkNfqICum7U345wAwZJr7rqObwWiCN9h
S/N+gdRLXEgb3jjPC5T6nowc6bcn3Q1wizWXbzNOWScxSsSE2JaKaJra7gxNTL44/HMRmtBquV0o
XFVb4a7l3w2wU6mFLFR7nqBBcjG8K3VI9Sm29l+C4ul7GbUlRjg6RzsxUPw5JO14n7ARZEoo6pXG
R1iXe5VeTESt2zhJjX3n4YUBPnXurZ/+VRducpTJ2vCHVYrDLXswaouH8lNQmkjnp/o9+wmduAy3
5fbD+9XUF2xEny+HD1nyT+nEFd/cNtEAuHxZMW+KJ8KUnjhqv0WV4vX8UscfzAMEfoP45URwkdcv
NYemK8dI4RSq9Nhjibu016SXlQKVV/8bgd0EVOyPhu9yXhylihX7/ivR7j4Zj9KbRkQzJ3MBoxIH
TlmgcxxdR2P9S3AIRo4R4hmm/KPn1fErS5mK7EWypqoj1Vbr1j//MaBPu84hTsJm25kLN5OpayHy
wicrZwPh4ijVZh/lG0ZSebAs3ODBPODP25LjWB5X3G8uKH8ok+xcpII5+Mdxec47pblxq0n1mBfM
mzp6K9cwz4M/FAEKYSymNZQiiJYa+V64UCigOifvfu+3Qedu9U2XGNcGLQObhe1NYZmd8T6UTJCj
i4M86C3CWS5zLXIffeNJ0dMorP8AWnhTiKIDhonAigVoQt0iBizDg+Xm45Ip7+DnZvlLBlPWTmTH
YkAnR0IfscZkvOvm581xy72gAuuaexsk5rsxSQZK3gkmmeAjo+6wBBPTiCm/dT1qgMidgnlqeq6Y
3qy1Eqihkq+/hskmU3eKvUDkwS30aZfQZkQgrcei/s87XemqYhX1jqMJgEE3ss+QW+5kB9pS4+i2
rtunouY8PilAuixj1NSXs5z0yHxcDkui2esINA9Kdi0MhdKKOABs/YKXAp7tRn8vRvYz+TLRl0x3
RC+7MTpE0pW4v12sd1z78AvGiRPC8iMAjZgh+rvRf9tyjgtcymLAJnlWu505RI7AwcoSijzx0uvr
zBFzZKmgfHX5HLnawD0VuU6bTGRdCYduP1IMgODKYcjUqMSFQgINncoO9s0DXZgAiP8FvKtUtmQb
5lYGZCmTJOPvhLGzD7yZpuyy0XNIKwuFB6W3fn+uqtZzPxkkTXby0ITo+IcWRAhz/L7goHv/OHVZ
Av2Js6oHkn+xLWsCFIUX5Iv2+O9Dj/Tj/lL5eMpYBwWnweFooMFAfryxAkpbv+KagWNcVdngTq8Q
hlX14BzjRzKFmz1FvIUluFNJXaIIipjngM4KHEg3WaNvpz1Ph0ZHFSVZ9yPMAeue0Vq+mawjj1jQ
+5zKt8U3lCBa/NzgrgDk4Sokru9iQ+igDeKUXyoX7jIS/D9y4sH1HyQmml9B1NtUmDT6Rgwf/Sez
hXRZ3R7SaPMM2dvVoHtpbuJN5lLnh4zcTPrrW2kXs2BpqGJ6Vlf3/FqCtuNz/hl539FC6574sZXA
fen9cZHvOWzuDQH80b8dCkyAb4IoixO7hGNeJRswuEU2AEecoRHZy/OyPrZ3iRiqPR6fMz/UfOli
3gY+1dLcCGUzFPd3+rndSM64v8BjQPW3kt2xZjUzFldcoFTVq2iyLWuSXkCcLen9Hq8Q4f08MiA7
8StknMZ6K3LTnHpQLXLswjX0aZJqqeG/VWQSfQ7ULnTskCqRhP6LjSYAPGIEIOxy5qYGaBzJ+O/z
KYW4cGJ1VsEiMtF6gxpk+mp5QsiqHoqDZkkrE9pf0hBUwcWlxEjza/XHogj7wItaeBWncu+wgf+u
eiJU+j/oUvW48CpJctUpm/1Vs5W3ieX0zmUButgJGFeIzpAbsL3p++yCaVdecL5dxLU+5CWoFfVT
W1MgeaeBgg7tcPL8FtLcc/soBxr30Jz4ukSGlzfJ5qbka4BRHWKDLddf25UBofc8YUnr0uzoY4up
bnhLVE35kfSpxuXfKU837OnLcufmvi0PLSVQfTLi9Y9KH6inQs7b0oeWsUbQAEwUGEZva0UxbLw6
PPrpcKertjVT2h6CxhORSdsgEa1aEbpfOrt4gWpoFAgJflwAUVOfFRio4AFzr+fsFe/pdnbHSJEN
oIuepfqjUXqeLjWDwexCUpwfdMauv3xHxqiB0I7YPlFKOr7QzLuQ/d9Vit+KXXdlIw0BfaUbt7X4
sog43XxlMY3+cRb/vHU5rUSGvnamWxsLh1XCPvnEH6gv0P2RVC4zokJh1Tw2sXNIeaE1IQ7Tt2ou
9kMLQ6I0/6JAOOjHru+u/CBflcWku2pygzmAotXS+6ri+tEEunPf6KoaLzWzz71rlR4LnWf0+r/S
t8QrbSYodhDpr4ukyrwiLVrufHPdI2XJvu9vsvKZhMIksL+zAILaZji8ibTD865qKOSwft5FYAbb
OGu8w6CKEPmJgr4UUW9eoK91b0uu73E9R5XGNb7nMM+7KD2UN4ZolhOjDQkg7nZksK+9+cm6F8S7
XMfdPznyaw3k+/MGxoe6NOsZCn3pE2LHyOwF/jk9EN/wE+6myGffGXxeWSylOI4+dS7lI6g0n+iP
mZgswk+Wv1boM1IiQefo+A3S7Vn6dRUGvgna21VXpKLDfU15UHQjp3wq/8kHb3CC4jdboxTx9Q30
13mQJUV3WzmV0Ogenm9ajkZTYIT2gteljM9v05QBawhDjSahlXlGHrAwFM/UAVqfh/E3FBK6oAGz
VQARe+cEc1TW/jdkb1DIS87236pBYDlhdbotMcj52Ro/q/RKmrRysa4e8Bn38/27KozRFoHmX9gy
ZGE28djcwu0boGhv+UVyOhq6noEiYI9K/8F5G/vdO/siYK0sMCaCmgdd6YLGiSqRAN60JlhCGJgH
C8GqI189ERW4SJi3hApRYFG8eMu/qwYuuxSZ3lzHa2LvuVEcLPWUPW0Te01uaUcPtQhYeY7pLAhj
MZKaQdW9+ty+oUme90FfHcSVks78U3dMHrA/Q1uzgP+ChTCgGHIeT8YHXpMkBX8Re/MTc0I9rFRH
vzN2WJNNX9yQfe8DpL0GRsUA9bSzNL4R7nTgx1gWMUilqpZ/DlrilesoDmBhH8k8tGBSUemAQFla
ewuC7yyl/cDuEO0+jIMam3ByOzYALxgAxUH8cAYvR0kn6Kj/zrbHeqo/GglNZloHjx3TFedz4MFN
sA+CdktsF+mpGG8FKweJ2UsIU/9MTyTbUjSYEWmvT875+bSuejMyAp4cqy5+jGzMCDXBV6kTA35C
uEzT6jFQb8ZmzFW2nVxbMbtOOssXpXqo/QJRpbuEMp51ZzGKQllyaMHwkbDk8rck5GYMzqKRi/A8
475GdOEDbFzfkKxWS6Yb7Hkmh/dxguzZEi2tERbhGzJz0CGiNlVxXL658zfdif7/9Z10g/wGDyS6
Do8YNYfWoqguCSTxyPeXERhyACqS4SkU4R/x/mNsrg6ey1Y7QMbcYIJni18lxuOq0itxWYIKxuPK
TbHIR9rgHwWdNSOxxKLWMo3BWQlyPRtXpV2DB/xnBLnmtx5bTr7y9V5EO4Hp+toe7h2dAVOGdiHR
CZH3zsYdNya/tC1yuHbZenL3leFJRuwgxNB3RVTNJY3kZvNwNYaxK12RtR4s1EOATHBM4PlGuYr6
BEuW8cCch9DI0tueGX2U2pwDTzGiNh7vq0RkEEz5a1AZwvWl2Vy8QQTgbXIYCUc7T61G4dE73NHw
FTamwyhYSq7TAGjRj74TVKx2V4fpLMWWq9wPIb+fYVcQYpAgQ4XUSmvlCpFJw+LIvzstasUmiuaQ
/2CN9ZuAdM3d3zKFBT4mouMfuOzpCn3y8AyzarW91IAa2ODF2/UdUIhbjRcIPtq3Z7OolcbH49+Z
1LcVuU6bNGhQSegfjuA/FesRhrab0MXOQ6ZnAdwnFwJGv4h9Vv0eIy0fjIKlY9WGEQ0863ukaafB
sjk9pAcGmwOCIAtlKLAeWxb3PQQQMbRG1uOflpYPyR736mAA3JT5WL0D6LcxlQE2UrzZFSbflExr
b84JjDP0j9HZtm4svwyRLAD4cHAOLDEunaPB674270dNOgdRC4qcnnWLK8u6N4lhxdSTq2oFB8Al
9zie6F5ky1Ttn+p7i0kfV99CQDhvHv0eOFuLhPK7DeJe8sQpX67b9ZXz1+dsqpkE5lg13CAF+w4s
nTvCjOAu0PFxTyilYvltTQ0xRyB1kcHx65tpChmIKtPsxz/UDbF5TOn9G6fIhxR+6BW6l9IFfema
CgaQIfOnRR+P3yjEHrFR8UsFAMpT6A7EwiUguCI3JSoUGag2OBB4sKJXOzldB3B2JgwmuHDWMkYY
xs4XWKQvpNsBrxhRyuuF+NVwyupo33mt3cX/+fq9Slsi6H0NywkcwOxkyLcnXjSVN5ZOeiKAJ9Cx
TX0jNJsmvgL9TxDBFeguTrt0TrZS6t1lk+fqwZqDL3PRH19iqK69TN4g4GuYue47A36JyD21aoYq
jaOkg2CjfepaDg+qaIU4p3Vf/0x+yKNSQB1Xg9SRYwmnVA8Itmr9AIt55dwFr7VM2HLNy3eeSZZq
XgPASVUn4zF1M1EQKDUEETTIBiH+ReSirWhzaudvggA00YUWKdfU2v6he7Ru2ok9jTFvr6Zr/O/c
4NQHnBgWXgoFxZjYHzZkkpkG4ZB5kn6G+DbtojRD+cSJX/ddPrrF3Q8jwo7eoXBAq4PjlzAhjLf9
klcLSf0VTCBAKOVoTTNWHqp+DUxNpZ67M4PrdIzLpJDbha4v+dUmC9T3sT+euBM70XbS2+zB7Trs
ObQtM8dxSqlYx8K2QtObnjHovuYEfujG1e+D55lnBCIR9mqXY6ZHJLt5Z2fjCJHcV42nCE5BdZTQ
ouGlkxiTsJAbCtutgBpG6eMpYVmy8oIc0M8gSS1D+rrDq4oDFGx3bBbUM6+h7zkbcRPTyKKR+u4q
oPrQz3mTxhfD3oRK2FAPnmvlVbSvxwb3xbWB/03EHE3q7dvAK6sdTbwbBKa2X4vch5128ntiFQtg
dpzOrUMVv/NYTyajK+ANWSjUJ56xbs1TLT1bzeTVNDuFm7owd+eibGKuUa+qAet0cYe3XNCqDS+n
DD4eycue1oXQ2fb4xlLnh6XsV7R/cKuxkIGUXBiEp5jYGViAmuoflbl2Uk1f5gBNnlL302MeSY/r
85pk2A3u/IJoIrBVguL0T1h7PHbO7kvC6w/QTX9PHISK8WgjcTM2CosoCtbQ/X54tFquyAUOU+qj
uDpzEf/H6RnUmsbsZoVWM448xDimKlDKsDIGxLEkdp9zgnrlqbAVWb0qFEFUlyRaS+yg7AOG12Yc
PjhSS08ZFkQv2NR89sBka7zoeSPkVJvV1y0YR62Tyl5PQKbU45gjOpi69yhN+35dm92FvPqiNyvC
IAwZKMk4JvQnyjrIUGTwXmicQcybLwd16XhLu/LxkNEzO3bKLOUY0sTqKYXkaylDrZqXKmsknwLI
tWANwL86jY+KrjfodoLWC+PUux2E8xEFuno5V1F5qfRdBJfAjjdsWGJY76hgw58IsMWt0SNUPVGc
NLqkutzB8PK8AT68xz9bC/56ggqgA1nh0oZ3sQsruNv1RUGXcUSp3jSKWMv87HjZnTGRXqFcgPtq
NvQX0rJ1Qnbx6K2a7D2F9fOIYqxv2DnVRkVftAdFc5VdocNSwOKRc48BKr8PSpC2hfdgE9GiSp+A
UX8UrJUMPGeveHWAiw+6sUHH4hsTL1GpN6UEHIdPMlv0g7IMU0D3CMyhYaew3e2QRfZ7rhzTEm2f
Uv1Ncdd38YxJM4oSO55nzw1r3TBYsbDy8Kf8rT6IeX6SGeAxleqasqRDu1GypsxIwACYDeVdNBxD
8A0qtZcpCfRAnWstg6ao78cewath2m1ultJC+GRAMYSy/TCfNy+VDP2kg+JX2l5V0JB+RhvYY/U+
KvSk+Bc8trX1h8SN/KgqqdI6bx1f2Mlw0eZmdi3S/p1XN3pMhSKQvqvuSqUS/N9Vgpb35Q1AoyhY
0SShcELIPCNjnatX4i1lVnHHaWll5nuc8HyphrDDNqP7KCjUFPP0j+TPpe3cgGqM+RAwfGUNJpuX
0Ed1IxOLuYEbbdgBUBSTRrRMRaJcXw+Z8VvygAlcb+AOAvQLQvhpDYk3bNToBrCKRlJBX/1IzLsN
yfBnV4D5pAvUyt6sAr/QcqaYHYSvtgL0Q8bfBWiHuUzMr7X3uEyq9rHCreJR4OnsRTBBBiJtV/us
3IfYXMfP+mwj+gM6YAX/pWx+DhFyrLXqNFP9styMEQbmB8ZvZY6RXfiPiqGC2j7TGPgmirTIdxX0
jdGUx+3fJezhSRkFsioxqE24ldHOwQBipNLOdUDAJbSv5Dqe5s7ub5nPf+7KpVfP/Y5zeeZZnitE
QEVoMnVCmb95MBMajSCVXXEXj1486uBE+gzVxItOefF1GL+eP3ZMKNbbpxkVpsR9UGORguPa6hLL
NIWYncZdi8vT2OFO2wtKLbjOwMvYnwo2a2d0Cxl31BWd/Y1HXgDh64IYxKw3arm/8zbmoNiSm6lB
OZFWO5yjy+NNaqGZHYXson2Xf+8Mk1az5G733WO/VWeppztDFu359UPhn/siNs7HK2DhsQ83Sxvh
chN5kyPqhyqsSHQN4q9TtY0kyvAlqxVyeagwJWAz1eVcq+R5KFfYjlTDbaheLILxg3taU0kctTbF
flL37xEWO6ajuG4rl5FYBrAWWK5kPCkpH3JgYFoRdSlfNksdNiE2ecO3PS9GGFjyHkYmgrLn4InI
XYR1U75J6459CvCLyDc5t7JuZNvjZVMxPNnc8XNhuvHTisTkN/QS7AqMN8TytBr2o5dFZihw0LxB
dqe/BiMdv8kMjSO8zB0h3vdS2F04t5Ri8fabnUftTMAg8QZDt2F8xW1f0fQeEi7JOLMrIIUlB05Y
9h9QzdmHCg8Fo2OCuThdRdmZlNHsRGpeEJPwGSzne4ISvVTObJvhGrBoqirtV9Em668zrQfJHDdy
ZgiWKULrb2a88yDb1wtRk/BfDkHQxRIakt9d2v5VX96YikH5jVvcoyzlJIIr8tIEUmP0Uqd4YKjT
y+b49SwO7IJbl+k5+ZnzlqMKrTRgY31aqyVYhMqSIth4c94raGNlUyKaPYpmZB7w3AS7ZioOBRSc
B67BIRrhoiwRCsnN+nf7x565MrWlR16bmx+vVaN4HiA1huUFCM2DQgoQHsNXl3Sa553TcHN8pEuR
nYebfb2JGqek7h7+plwpfMwb4FPxECG7H1iE6qHLENSuWcQ537e+9ZZH7R+XH7DIpBOf2ruhdl7O
NN0VLw7qr+PbcWsUt4iTVozI3lG9yXlUAkf5W3DTwTGTodYw/sh9cXrFUc7XXSjvQINqdBYyYFhn
ubmUWu749PyoePVUC9LE5fhVtUFyQWAUGgbQRkLkyGO87P3DroExBJzBvUGJ+snOQAhqQnGZMGyW
Qm2ma1VCyI/WyEAdUFDcBIi8Ar8f7M0X0l4V3v2bTXk0pVOzhxHV/htFwFBZAZWVPQ54CXa+xlNe
YXbZSNt6WsFoUDkJK2Zrj1++9xQfxJ2DanprsBwm87Eg+xB3CB3knWKMn3e1xEOZfwZK3VPZyNQ/
ki6s7nVf3dxDOG5EKJ7R2m/QTqhYm5XzYYf9+ciOtr9qYa1bwmeX+2C6U4Xo7+hR5RiacfDQgR3u
pGrQG6L2h8bEj8BIYGTDmermmv+nBbPKlsPbC9cx4czRxky1WD5sPc409o8qJRbEJRhFH3BBdn2I
rpPD9WQFwdxPBr27DyRzkywN9bvYc98Y8VckpLc8i8KLzhYSHMPUvlQA+oURGfuuU6Hw/7Cv1eaZ
NUUYzHl0aairGtELMSHkJ+pFpuimZDP/7C6wx7Id7d05yEWLGKN9Ez8FeMf7MH6tl0s8ziZtPydU
RZMURKL65P35JHdm+HyGlmydazegXkNu3jbQpguffCG/j53Pv+NZSykPomi5+rCPWZUtw4KhL0Or
NIv6bu3W7hJqjwSo7cIJzS9DWNqpLCGdaZzvPrrzlrVu8WpEvMC8hurZSh9BhxNzzLFBOTZhbL7K
D1KShXj9xEN/QWzhKOTDWtp9v/e4PndWbuB3w7YLNGXRkk4nxl0G2mGv9pQQrnGtqNDGHTLdGnNw
p+STatqUw/G0kkKUIjUxHRJx3+/KWCu1keOk738+KT4SWo5IJFjQLJ/m3pXgw5PWucAOEwqdsdkI
8A/kTzxq7ASR2raKvO3T/8CY2Nr4LTpO191jzsO1IqTTvkDYErH9HUHqHWdXPwigWUolG+unxcgb
uOeAngmzMw9y8TGuiX+yfSLY5sDkgh0/d6AJLvXMgZKJ67S2IELXdz088ztv/MfnZMvOUGYokEqU
A/2WakIGc+Ff1mNlFnNswrpOZ437WxPdBhtAaflwtcw5WWrKeDcdf/CM8GWdXSg4N5FwxnBGun7L
JqiIL7fCtXiqsc5AgKW4GEb3LR2dYl5QXZ3vTZJGGzFaHlYDusTrTRE5UStqG6Ne8TcO4+X8Cc3C
jtj9eIf+wjIM1t8Z8d+RZZE3bYOis1yxh3QpYwLf/orx97E3CpbjqdN3Wnvuuh4cmykL1uO61z1b
Rt+OvF4gBly+3t8EGUlNbfTAXyGlDxWHDz4V+dakQqz6QcVFS5TXNJ+aGmUr7yn5adHI8gqMIspa
rVmSR3KXujNAxsR7TtFn8sJYTkToTiKHS47eBisEU6XMKzih4GT/8tOIDCnYZxdAVwuhOtchWaqy
9DT1xLIe5wrtELv5KgZiRzYYMmfBDmJRb0rhYcaSYpzRCBsGAUZvArMpmqVLjIwh7rvxdhni0x/A
fFsStLuz23LWl9YhSD5Er8XugDIOFd2jEn0+xHoLxDVO7Xguwg939bW57CM27sSXPdRSGvUfhSER
Dk4fSmmTQIzPZmj8ReHlGjNz5P6wcJM8PHpHy2MRIpKQyZEPWD5pxyHkHTtyNYbFvEmnKMKNrD0x
kX0xS95GgiSQJT8nd3a8kQKTpCUEPSRKlcAi+9qHwfGUPAyzJl15KDPDaLJ6WLeFZwwNuqiF6tba
MS8+JqTNaC+pSPVGoqWHzdcWjexG2E1VBdQ5lzs/nTGnE48vYazbJk1sk1+N0Q//6M0t1n4XocAG
4MP0/o8xyZGqiNkBviixciEilRd7OsMKG3/jTbEnp6YFwT1GoSJPbMZmMawB29mryJa5Icy595X3
0LJadKwtdJjMMnO8L1VAEELFSXfzLOWNK7nn6aHXBQH2JOowejvTgpYkEqSDXjff5SYWWTsvvfG0
xc7ndx0QT30AX1LBUCfl4zrjXkntQdMYW+8586klGUtgmO0cC7QdtJFCb/Rgw96l40xczN8EFqHU
9S155wMVUP/PY/4grGD8e5n8cUADzbR0DkmTPRTvB0T7boJOL0/OLKGvNzLtWT7jC2720C2uTETj
hg+6H7zHBdxHbFMZbK0bVBq7CL6nerz0/Kb/aODKmC2G45+NkmIzwplqxaGXg4DeMU4ptQYTnJsR
DnW/vWImIbZBY6QZqGm745YBe1p1m9Gd02L/xFqXQM2rfviitM7oVxkcnOv55uh03CH65Ew7SNf0
jx0GYZSVtACQT4uSo4AomKTUWtzmnA0lgyCeYm5orObm933JwwG30Dhm0eXbP4vWnltVLwv+OmVN
we9K9RVvwRt+WO6VaKW+FEhh/FlGyN0XSw8Qwu3vTV+U7zkxekm7a+TZrxVooIfcLeupThNKX4hI
s4aGhHxBHTt1BoN1mYaFzOZLyg3RNzGWG0pT+KHs+tx4TOzFmWBALMmLGMVtveuOrIrxL80B0qyq
ANl0BtB3BG2Tuk/LIijjWphKuR+JZHp5sYPaJrDfqJh9uz3PGnAgcc1CtVMZ/mH5UUGkqzxjlsYq
i+qdAanxtPzWGuTQsVeaRfDrHF5k15gJxnUXBCc+h3IitMviiQxGmrKOJxke9Bspgwk4tJfGZekk
RrDtpeVlYU7kr5lDItMh+HCs0ys4VjD6VFfGB8fBx26c32Vexm6/s4C0tmaKRacaNDPj0bQoD1uw
TWIxsyx3Sdu0IA3ecZJzWAAu56RweIWy5qCq5PNYCGzi23x4gUxF5CWsJwYVsZopupdMDJFk+2TL
xNz/UtnjdATBASB+hjeWnCjx2gTk8bl6il7cTL/j48Lnj1QI4nDlLrI3BUT7Ld+EdXILTjewLDkk
Rq8VBj0gSwajWc/6inDxc254+kI+B8I+BGnLh97jRwNiLlYWUMzmkupyVgoTUfi85OA8L/oru5NA
jfxBJgNTW8Vo8WdIvpIkuapkVcZC2PHJcsQicrZJmhhcBz8/xqDGvAp3AzVbEZ+q4B6Ck3hXMs7+
GTieeQBtQ5vUx9GxBtN5fFL/zf9RP1XlokWCWvj2riSMPWFdsPbEhglQSP921de7l/ZO68Np5FVD
FPVcZKWUL3dCFD/KU5SUCMApvBFETiZAfJmFIC9pyK55dIB9i2GOhHzH81YqemWKyHIihJpFAa7m
RieD25aNNFnL9vQhNOzOO2iql5633jVkJf6kzgLivB2timibxxFGvvtX/BHTNYvbllp2D4+/3qVz
zWvhgsw95DCIMOlW+S1+CMCcoAGs6xIzoHEpSUi5b30FpWtiX46ms9FMSkXQSpd/3Imf3/+4xBGa
5GHTY0/QG0RVgVZZKzYl5vDqs+VGhootYt0K3mZIi0Cf6O8BjtuCaJGGTgiD4dGQiYT1OzgTCseJ
DcG0rkfzojWHYah8HOFyK6wmEMX6bA5+ilTlmt96V8ldHFYGTmdXPr7JYNi8Mx09TP1UK/rGSanr
8cANQdSc6aWN0wZ4hZ3Vul/Zh8PeGI2aucoT78PRbQome6JICwzOlykOMf/Q5fDq2V65Gw01Ogqo
p5XiJLZllXqb0Fbg4RWTKOVQId4bqWP2W3B2zNteVtZEnE5x9eq54/c6o9H+SjWowy1j3oF8W+xB
p/owS6ytvJXlwc9Rd2PgLydbUJkQoVthDYNMvvLwFEM+SR0C4/tbJoF+mDYijVTShsjhocIhXUBp
dK35IA2bysp2guSOLEZacC7WO53NHRk1/xmC7ylku4NztFQ/CE3ErmjnitXoD+ft0dvsKNE9Z9uR
K9JnOI1E+Wun7dADF8Pieqv/rJmz5cPoRq8T14xx7Dlm3FvW91FJieaKWTYYjEO9GPaEFBpE/7ra
31bObeq34qzI/WyeMwCMZHlH2zIxLfbOheUi3lFPQqa9BD/D/cgHqDJwA4r/2SIF2+aaDaiShyTw
M0n5BnxoaTB4qTQ5SoHDhimXqgO0jDEBZL7U5k0Gl9sZrHv58qeadPnycdcRaFA47k7rcnXAJRhO
+KT1zCzh2Bfq8ZqEoRPm179SC09ep1P8SbJ029KAC6TmUPzTJvVScuilm8OLfZ3rxuoXyHmENOR5
hmxE8yBXpFekNKL4Zwsyxu4SYUfqbWLeB5Ik2G14R1ZZwGraucLmpbBWu0rgS028Ijl3lMvUBIvt
DII+y4kiSH8PqJNtBiNXBNj9wkrMw/seXIAYZvhQkXuHtm983KMgfrpgNEjhkIcC4RG2fLHbUXTs
EXBeEegw0jcfDC5Fz2f5FEIvMYOOJE7iQPbHt/bYHbi91/i4EARztR14ufzu1ht/VInoWVAeMXPT
BTsVc4X7Kgs+vwJDXPFbnZx5zfm29wTeSp+tQgzkVrx0QHYnZ5ZtwWF3DoFEnlY5waw7Q22Ppunh
3K6QXLlRSGeIClcymKOKseBUEsHQi1vyBq3HcrFU7H/nylR2w0TAeCJslHkL1E0f4MRUFllt2tQo
VhrD1opGVb4rTzZEm3egMWgEfv+iwJfiG+dNCTbEqpIChU5uOg1ayKZwo52h+8oEcfGf99cujBPT
VMmjiWe/789Adr6tdIX5sDuofm0m19n7DcGGgDg6z+uk1NxdtefCb0Waiq9kow1SdvCMTYRAzGJJ
BOVSB6RlTwhsVR84a0FkvapVCXQUPinwQoA5gD0rA36EMEu8qLBDDGJ5pmdDgjuxG5b7S3FO8F0Q
Bn2VPWN5eHaOAVLdx1vOIuAbXkFAgc22s0fvGQRMXC5DLWBcLnSzIDVq51SWLypRLcm1v95cK+yt
YNb3luiyWJwud8bej4PcGM1Q8ziuQlXwtbM5vOuNHgUTlkbE/QsbTXXaEDm+IvTXMmr6cSkNJHfu
jTc0zMilkeouHUQRx07NY0fgYOczSx4PXkKJ1IxIQoyl0/Ld2w8M+SVWdV0X4JYh6m2AY2ze8bHO
H//RjUEJiBr0G+gT+s1tinrX0DAfKyJWH6aJC860mJooLJxYttVpJj2jHetAhqDOormJrbL0a47l
2oWNbnY9ZkvdniZJjSXBM/ZtJzRFY0LeLgrnP3j1MtYwFXqAlOWBRPN4SBt0zjbFV1qhiT2Mg5Ai
XdYMUUCcjZWaYR+3joxieUy0MqPmyuKzPFr9c0a6n6H3qyr2RFvap1ejz9jIU/ooGJy7O3k8ju9k
es/qccv5WH98gkLJyQxppTBhG3iI/Vi2dB9ZexJ3fVGgkdrKf284J68mfqtkNgllpo51T5UO8Q8H
IYBQCEKuJQTnXIz6b55bInP0OwEb+z7WP3pLnRly5yapugv9KkxgtLOg7N/2bx7dlrscAJQoZf9o
q88xtiYPr6yFzlrOZwWVd2HMhn2rU/1+N6nMUpG+e9BOjHGLq8R8h8HnztNQ+YeJma9RloHgGNVa
LnTJ308xfjCMuuhFWdOARYVRB8iQecQwNC7OACGGlFAFhn3Xn65qfiMx5fPzZg/oU8tcye+Ox7/x
7OTaGkfEGXzjhixLGmGbQTBSzbOg+dhoOT7L63zyw1+00G9lbLkXBXtIK87Sjyu6PHdyOShhAs3/
69cMogypCkcWZTLAMtBw2MMY8WsuXWH5jFOCnR1gfOWTGOL4ehIt95EcoUkHKyLkde0Rnhi1aWQI
5fadxowHsFU9S8qIP4zKHEsD+67TD6p7PjsYkFohxYU2teXc9zW5Y+7yK63WZXc6cVyzNgbWyE3h
YIH3M290qROrmCcll5x9FMn3ij1G80NUc2/B5ffz4KlqGWaMslZVFI4HWd0Y/4K8vc9p3sZPZ55u
it7qVsyld2/wBP5u/Vld9qdY5xpBBiaOHUBVRqrR868uzuGsoU2yajs3X0ZI6AP7P4CyYEvDiW0x
+BgnPPyCLwOvVIhWdVVbBtvLKXCy1eOOWsHQNTeK5MWr2l1QKxtQs5/kBfWp+NOWzHOG3yp6vmyv
fF4vFNMBmTAd882mpKS7ZVxtUICxiorn0GFZvlTDHzpu7jFGKDO1MZxP3KjEY40WDsVDFSi42s07
cPeO6MBgRRTEztUlLiL+iNapVOJMn5UIoVGTm3+RKimCJ8lQFPSgmsEP+yvAUVC867H8CrDd/vf/
S1RNpk5eJC3Di6l3ngaDYUHFm//4XShJITXGRT9erGr7a8mmcPKPRvCP30OsVMena9VsEw4ZkiSK
RHe9jvv8RQ5ra/29Xqn8AaunnsVUnqQJlQVTQTIzabCJPSYB16QE8udLD9Mh9JYw9ekD9y2Q+KXw
BPqXxylpgiYhDpuVTsSR3J/acHlqzbyZiYBRGOCuSzCCixfXyVFxZaGkUf7V8bHw200oqlHLARcS
nJ8Jmf/yd2Acl4+f/Uk/q943RUmzI8hRE/jqknGzqDsnB4yiLh7CHw/ap8/wLNYKBRzeydMWpque
zgHmwZ6N7yW3I0avRfp290g8hDLTyTytGAnx1VMkxyYvmgboWgvuBfUSU1E8lvv9q4+0gqLs7rNq
FURu6TPJHqA7PxwR0hzXL6XHyG7O9GtvN92w/u4p//1kdKWh7GU0v9T3ThXUG3XSMv/9OuigHXAy
9NuB6Nbgl815B1vke0n86+Kl2o843Cxs8tLDen2hhx9tdBiAbxgGTmtDdR9O7fAmTCrNuJhxjxWb
+2S4rBbX5G5T2FIr8cgkF0Lqof1z3CG+Quj+5j/RhL0N374HeO/aJelomGTQKDhLYwTXp9LmkObU
iDR2Zx5TGfCZUvlsWOaXDHeJ2E9AIgrGx5Ob/8lrdC+cmK9IXcsjhP6BQCzTjSkvn1xebKZ3YitX
rwhEmgn4k8Wffd8fMBcDyqbAMliD5Gkg1Mz1wMuLeQACKHxoFSIU68Ie3wlwFlyvgub2J1AZ4rMS
LBWm2GN7XnfWP5+WqNFV0MpjhXGfa0epU0U1UCY8SzDz101rpV4jiKKEJACMI5YXfc2jqym48vz/
qoYt+XVSojp6xvFPayjtIpctR+0hYu/kB69yoltvdiYgN0moYGH2e5KcaW8uyjzJDJwYykYDGKzA
CxEWzSvyEauDF2wQpZ4X2t7lqsJsuGnnT8HxxXu1OyPCFp74Az9AtdnzjMsJw+WWoOpLKLsWLMMr
4sx2t4Fk+xw+2oTaAtk030+zy3YFLBzbUgYq1t/QDTd1br/ZpLsxwPOAQz/xseazCkBHiYhAwIX+
D9YpaMhkQinSsW2ENuZ0V46n625DzUQ3DqJrexT7RN5kAB2w/R/udv7gXovdIasqXxgTIqaeeQhX
GCTdG5wqLZOZeJfgAGuTvKvrG7RJFtB+l+GSsb2Lxa1FJdgxHP54mtYYEENx+JtG9mZNxxHwnOgy
l55NrypYhLb0UPuggE0zYtnmQuBdKaPNv3m3UBKFPjdwefWSi8TbUBGOZz+OexGjOyJqQkdRmy47
eNobPlzfpwoR2sSyqh/woEcuxBZkqHmrsw/gXgLz6XCxdasKKuz25ndnFA38CUEvzRa177BAUj30
C/ziSsMESspJFoWUj+36R5Vp+D6u5VFySMrLvv+HfhI+NP06GGCnamygul2g3YE5+oRhiMg6F5wj
YwjU2o0zCJWRoJ/pmiZhBfBATkzZSH4uZt+DmglWZ4yzh/VhkuwsJZwr8FWlp619rsbGW/583Qa0
2ac4tUVwSD7lUxKxEtuPiffodGZW4Vcy6lLddl8TsFdE+kpgRSH/HfhWJ4BlyoqgATIonAVFy7ZR
nO4H7R6ztjjwbt3uQyaZ7k2tm1hMpibpKifAuw/dw9AjnA8VSi71BngNRSycnz7/q3E3GPrXOBbM
ybJURwjpi2pGypi/7g3mspYIIYzp3bvL1BBhAMekhbYKwUgDyV8Wt+VIF1pNQW+7nDOYrmXFz9Zv
L37OvSKlazuzjuYwdSbDX8TESjUXHa3JFaBrBuAY4WiyUnYVtRRKHTEIEzk7PUvVbdAeDONVoOPg
y1WcV7nbO8zLsyapssBSquIMJ37cDYzloSCe3+jJAbQ/m2vKrePH7XaE1yjGUXQb9sNQkHuXGpnV
Bu8bJOMSvC7SFFCfCd9174c22Y9zjcbRBZ4mTjdlffa4OpegsIeBIwG1d+p64/xNx7wXwyHmGdh5
cBSVY3yv6SXjJh12j1eklsh2FHgr+yTBhtH1dc4obJ8hYlxboXyKmU7+Zk6lsbPceZJyvh3WhleZ
UxYYyJUU0koLigiuETJh9WoRmKtSU+BXmlrTOVIjAUIM7kLVWJho3w/nsVa1W1EWtcoXuZQ9hhQw
9OKD2p0fH8okZSlS/Lgh3wubaDQd61/f26e1Qqx6nYCoadMHYu1O5hixSOhvzuT/YSN9j3mRNLdV
MVG17txMzRBvcbSo/BHAyEv3f525IOHycNkO/ybhUc0UF2bHIPyq15zsVfLblv3XdNhjKNDkuZDV
OZISuj3lK04Qd1vQuRE/UgXr8dmGyckUkBb488xZaH6YxxQjqYJ+esjda3X39ApnKUwNiqr3RU9r
33Nvh6xaxHD16JYcwzeIWwYF9ck7TTr6F1vXfRJDT7CvAmVEsFHeK+tnZA+fAifYXG0eCLzHHs8D
vnQTSbAmP8+AUol45FC8++3MvKTgvwS1aojKo0JkJP8akqRUFud2hXE0lH8wnHArhCu5WMx7SLDj
03lbAVktM2dlnVvTSGhwFZDFsfgXL9djN1Hf1tC+VqCjWkIyqcFYGphvN7u1cQ62NNZ5hq01lUAm
fESe7iM46JhQnkJxdF1WVCXX95KeSyuRrL96EWh4ZdozsSuVqr7bEl/v3eBJz9afa+zTVNjbnoqx
WKgXHi/IcaKosqo7I+kFKPNVZcViGpWPBznTfN0+UJrg3+WeT9EjUWsVPX0xClcR5WXLReo5Cxtn
/lWhXJF7jvWjT7pOJv1SgrMUEZ4Z7aCEfH8WN5hk3DjBLiswR61QHgIU7pKcdLbjlAzQTbW+lvKh
3jOmnQ94kjl2juYDka3GYnOC5OVUCVmbF3NN2hFtfw8xqFZa+m+c35vA9E97DexIKNuMJa+G/q1R
KBoz1lwQQZGuvNsyFKQv/sHUQEe5SReKTLvxG95j9rInJgfsDXFWMC4GdGreRjyKDZ/9Ydvjlt6f
sSgYfcT9GIscbindDwjw+bmGHwsH+EUMZ4nsqoBKiegITl9y2sMMlIPm9uJdP2yblB02jsFcAuct
DS9e2hmXbdUtFrYY9m07rm/Tw1tbJQgqgAGuAHDrzcbj4EFN9HU3/iaNAm3gacmzn4ED+mAWg1pd
KoB7eYSWYRdF0MziMWYD0ImTI3g6n4MCv9ytHbFQihOA1F8x40JjcQ/MFnyJNB7g1bXVpYf17on2
oVaSG7PQAcdSH5snPvEkhJuyAXGVtHrne+njOoGe2eb18Ofi5J4VhR+cfA5+ikAoDktxghgumU96
OdNZIgKbHAHRGNfWZkwOVAj8xbmcPCCrJxxj49hhhKdEqOmh1+1DmgwPrBknXRnsZDW7CoETgL+M
+PFdaOIquFtkymTygckijA8nH2wpql5v6CuGsJgEhHrwh1ezkD4n/24x0R9f/W7X/vGo7I6o7Urh
ML+Kvub1qhebh4+N0o4YKHvIiRR7C90t4Radny2lGSLk6EQ//kKhD/FrIs433IfcjPGCz1x4Pm1O
vGfhC0D9dSiCJHU074UqhMIWKVGAX9ui/YOXxzUjsQns6ixvMHQ9r0sFafmFJc2Q+09LA41fcrT7
sB6z6JqQmxUD/iEk8KtN4h2NNYfhwkW6s5pTDBnOAe5Oi8b+a0yeD2QsvrzT6WbMPR/1dVCP3Udy
y8o941Q0CZhO2Mrd3mwYnwq7YL2uBM1Q4ruDAI1IEfP/FMJhJdlJbgLSAedCaFDVGO2ga6WYCUrG
3G+FgEqD2KPK2f1lZvk/IPG0B2FMoUXMC1k06FfLL6nJ6FrdrK/YIQ/8p0bcV6lc/sFoHiWS6End
7DKhf9yteaDtIYayHp9IuM6oe9yZte423b1zcG398AJHcy9Uj8aYWg9LN42Rh0jq55eGvxbon/Su
fxsLI2fbldv2eTIyo7ZValjLLxwDsBjmIxAXWXhSfIxzrQwHomiZzOtYxtmTMz70UVN7O3+aK8aL
wrlKIrwFg4PRyyi0xse/sx6OUhuGbkPtY5tCvEyzgxerTgwmdT1aT2sSG8IV+RK4NM8x+84+yb34
64cVsYtzeQeBYsurdzHf8B/G8PDkZAfgBixjYt36y/qjxZ/UeYQhqUASWuLHczTNfBY34tdDm5K3
E9rQ9HfovOmeNb622y3K4J2JLC2+LjQicjL5H43npTFbGeNFOWITV18098hyuqta68nlUznDAD2z
ZuD0iu532BOF1UWw8CM2I4pVOtxhljMcauDwob5gUgSpyS8sqIhyNV8lmqPYKYz/FzpSd6MO62Ku
C9TX7QBAYimWCRQ1SMa81y5sTHgoPnzDRVH86m563B8GhN0IIvn9M90ENqCk3bOyyH+ePiqgJXcb
KxFe4VzachYJrYXKsJHIaRDVQE1mSIHOap59KB6XrOshueNMWSzA7gvILJcgqOgL6Fq6G+bhfKKT
FFt1wihX+bPmC82tXeMz8URiHP0kvXurp3qgCOYB7Ett7rBqXS0OCcMkGUfP7oMawlwC0TFPP4Vz
FOh863YIFhXSynACOx4jGWoDcXvsj7kaPSVj7jDZHYNvOuVYW7hUeFMhCiLKCzusGQZiFuRgg9+d
ww1XWDiaw7fPOWeYJ4VL5QEVGZlNnyUEXdcGoX2G7MSgiTO5OcD0w5wcTIcns1K1sLvdceM2jFco
zEBHtLrF1QnPHaM9TuAkzme/VIEW6c49bIlwQvjdCnfp90hfvNXNQjDSwM/tk2eyt+P2Y03Us6D1
xU8qJh1XFc/Dw0dkc+hpk63r0P5nYZLOkCSNdHNFbhQWXAglywpEN8wRSY43IgcvZlNVanK7bPQo
FdbbC4GdaZgoIKF45pZ9Qm6UCZFynT4zLT8zl4BD0+GYyckYRnWrT8+eoem02kv7/k0w4SIZyZbx
0WD/oDR4/XuJhYj/RVBoChFE37xBx6A0HA/efhe3xCriggup8g5y8f3IPh/vBOFtaCypv7qJW3vD
+lY22aLRuwOn6zcfRtXq99fhYafZvJqZ1idkesW0H8q79tpzcEUbGFdyqXHPsWNUq3Qs0NxY1kFh
dXB1l8AIcd0DvdsO6TlWY7Ggq991O9GZp8rYDjkBHTCYFvt/A0+yXh7ljL9XWdeaGyAg3yzQwyxP
BCdFN/DdwH2RUCcHxLIMjpB9Jxl4U2IIFZkJnoDwI+RZRJwosmXTUBKLqFV0KZAK76e++IM4Vwob
FC+7VVL0NVYFRzdJzDVfJjlGRudAUS8ZKdy5wHr4JKiKomn53xEYRz697fhjK9c7236JXTse8XNW
XCT8ll50GokjqSvBSFKXCsg2dZrfIljTKOx8Lr3PbGPbULc2fQpaw8wa3oNqOUu43BL3eVn3xbGe
WhNmHROqeEcO6zNBtFS8ZQoTWwqfrmn6QGEgLRUAm8s/Cx9ezfjo5S1746lqTQV8jbaf9+NnI/Rb
6gAsem1mdJtSjsMK5n1vDd1zuhI/YApGxul27H3+0BPozy8td01SXL4yFwlcJYHbRqAC0Ue4XY/S
djul8d4FFScubRMAV9wb3ReYC9ApdQhDMrtXutKNpPqb9CwKQm90x2ubOB6SKG97UO/XuUB5fx+9
QwEmcxi0ZPYgvsv8CIw11w3kA2aqRU9m9Yl8DRURCjFbOKFGtLkSGMAbu+KGH/Ztt1FeHxg4Gk/k
+2/uAfwbF5RyUvSQr01rYbVfUSdwM1X/FeEh2saxSdE57281Cg3BvGuDx+dRpl94tBMxxXtCwzxZ
PrxxqibdCgckCp2DXwUwYQ23HWZRgFkDih9qeqTyGIKWDRD4kOFaoC8AeysYROtSbZLv3dCW7hMc
WgPmeCffR48nk0+UfZDSUfFFBMebmNpPFDr7UCKVVkv3jzj8c4yDTZn6J6DWlJr1lLcHvZ19B6aI
WERQC/eCRZEtXbTUiCZmSqqCE8BbMeBbeMhcygXpllq8SiU7Uw1F/m1AMBhnjK80Q8FAe62KisKc
rV+Dwjh7Vg53J0/G2wp8SkS5qY/TvF16/Y5ionBU+vgdZdZTgVAnfetIKredC0rMOj178D5QmuAK
8xLM6eF5SxmJ79qS303ozJoXPwCSIXCTtAnlvn51cKiGZxoTwldFsXz3KqymPB2S2WP3OPJP7FoY
Pp2UGCxguQ4OcON+7f56Yvd564DeiVx2nE6pdONv86nj0bsW6fH/rsjfgXvD+FMF0tzj9ytHhyzP
AQOt1KMfcIcTKDCLI2cnj+EY0tIiKiMJlttjHqkYh+BJfhE/20Dh4o2+XSHzjFoxb7qkF6Np/SSe
a5b5cokkRYKvFH/VQKI9MwJ5qvr0US5UgSK5gzszy8aYuhJv2HwSA9qrjQ1hSUge5TvUe/8gBwOV
p2QukuEyfQO7NjOmMsOmL3Ss4ncg+fUwuxSIS9ELu7knVlGiA8wOQ4wMm6h5l3fuQ7ppTsf8rH2A
+UqkDG9VtTOOeT37oNLMYOcP0XWqgfOqxb1Ev3c0kpANv7Xyua1Hu4c2uB8HlSfr+ggdAShCUTeG
y5UjttcLTxbGtTP2e4s3c1BBTY4ImSelhFmS1sSJlz7pERXEokB6Lt1eLx9WL3suDj8e8kMxRsBs
nR2YADF8YiUKw9YS15A3jpx2plKWw5chTooRS4bjaAYWxPrhMaDZmWdZVFV3iMjvS3m4duJFwnWC
T6dQ4qbrTWF3sdOxjtqdbnJZqhr5qaD+5ssT903KMCgP4gVUF/J/D+wUMlUkQSLu5TU7X6+CDNwC
uo4dRHHJBkN6RZ+dy4Ov0XHb7uzTXiAXP5l9HQ0PbkUjeQbu7Q2gMZpnGrHGElPEaEJh1fGgdF0Q
7pBw1V7R9fI3x/xLH9wG+juK2z1+suwLa7RN6kaGQPP3HyXRLDjscum6nLVP4lTXflKR2rSkHWH1
iVGvE1wvHliB9EN3ZjCpbtYhnMQ7RWMyOjRwH5ogjs6CXV45xDMghDNBOo4DCDKyvjYjS7jnzLe7
E4K9MGxMwnUCklj3c7LAi0vllOJyPENJOvLhrpuKHsoy1CmtjT4vNI5VCK4Bn6aRY6YQQ/0bCblA
m86J2l3SHaSpYyExU1A//Q895G8Hp9WARDqqkaacpZScOPjmoF50X+zxhRhavZYwndS1RP2AZPWN
ezdlF4hENda7PKOplO2+7ur/8V4ez7MG2lYE0FqxXYkCYrtBsI4O/+WruQR364dUPnsYd2XezXzV
Cf08yPiwDSXibYGA6ugxP8IJl49xDk5q8yksGVe2WofP64eBSQmJhRFhNUPEOS/W7Iz0MeGBEPqy
uw6g1K8q0ySy8ooJP6iBA+h3kezXoZlwuUj5E8g5FVX6ZsZGIIVGkmgGOjf37x+0pEvtQA5BdG/c
pkq/EREkWAk/uEQBqK3xA//WEp4QuFP3NQa9V3MmtYcNToT6KOHWA0FQ16r1gznxaLR1JHsrnad+
qfzm0/iBL///AaXUqKrzLQy7FVqpSRDlFP5HhFn5d/5z6lC6PUgDvgPDmmUViW+CZfEdGKG1sVvl
40BExd69nUst0EkmvclgoHYWTq9jkbITDpd5r95UvI4LJRdP+BTS4s7cHLcKPNaF7OohhaypxUI9
GoBrIxGVVus0cFgcuN3bhuXkkVxIxPKObrGWv/JZ50qlS/jkLy0m4sQ624rFg8taWsVJudTBRmNI
ZVMqedlMDh3rgRpSLQo2e/gGUVmmYE35LpsXlgh89khYgPzq5f5ekpC/WSX6czcvdBv8EeDDGcw6
iIQ4jfE3YV181yF49G2nQQBakiEqeQZUMUgDLu7Oq39tLWEnzTaXnAzOqWpMxVkevEQ7ofpy5t8M
Ku/UozBroKq5mPSQkEOeXYODVOafjeWE2f1mldCHe3rdUFuHWTIfkFkURCjy9bdVKeHC6oD/Ym1v
3OBF+7HoEnk8CYz5m5FSMqg2RhoJazGqrrL+dzHFDYv6ceuYuNusXnX1d/BRVzAlJz1n9pHZnhF/
XqxJ6BPtz3zmNCdLp62TbDaeOXCFnz7E9AWhnUndx0y8Mi0iIk4lh3t4fmPwkVa0EUkM2SsMbGv7
jg1hpxfExmlz11wMc3LxP4/yFcg+3LJKBOU8ucnU/bmbvE/8yK7LXC+2/4nH5OEgo3VVZc1r5vYr
3py2Ji0Qo+xmKF3iwKsdQ4PfSgqC2FX4DRSvVySWomF6VouKAYz/vvyKElO+kufy6vKjE6zg7gYA
/k/e3JCTKWzd2o3cUuoHeAvJ4YoVuzxlfZH/9/MpzNTQ0krvzD2W1Cxr6uq1eAGwAG+dU5pix6Ox
98LuqG2qf5YDoLkAOmV0N9H0HVxE8APG3ymDPfWfelmm6wRmTpOQEx6PgVdxwWvWfT8wOokxdRPK
N9XhuLAF+MGoIzT0j1k7+Is4stk2VaP8ufbhCK9cxAzP6jILd/DzBeJMRltU/Qjj/8KPJASAgZzm
YfXpuTcVZx8adlBV9GpTldzJy6/+Sh+H+AcLl1TCyU5fwqDYJopCzaoE5x/2wfMReANr6fympcmN
UEaM+a7cS+qQh3LqOhax5vC26lw7K0Hqp4qZlJT9a6tQ7RMH+/YNo37TG+LRrEipcWQvFGMvo500
V5xAGblALJus3XnB0DXKDy0lrfdHhlCkYc9npHLVqxWFCIa9V8zBXfzI6x/7bvuvkBCS7rpKTWS1
vey2kM76DE3vZuRPqd1GqS5+IqkJaLtw9EnZDKDK3slPY+OgZYZbJ83F1dR0kUmmvBwNMxghHk6B
ziBa6et+UBnZE/fisWzJlzD2+hSF/Tht1H7d+honEQ3x5V1cQvtyB060h2hmAGFgg/nTEyBkzMT2
EkgVz2qdVVilxWY1BX+uZjcxftTd7invRQaalrhUV2/Ty+GH2l1bSIYY8kLVFo3yN3it/xBKJfYy
T9iUp9svAxhtLgae8wYcVXLSnfow2eeiXSRjr5HIWpFh051ZmKxjnFyEVjomCfRh3cjHLA3r+0Qh
Ov5IIi2nmAmqMVfcLz8YboocyPZsl5y9WlS6LsxCFk+CWPUZ/NsW83yhqlHDJQ2m+8Id6dGXSZIp
DntwkOGzcQanBgzmtzxyKEEJUYL/Yjsog8VfTXU4v0Fld+EciQqo/1kAEabdc0ADvO5DjCxoGy1n
h51BoL8SAVeVYOmhkf+V/3GbB4EMMHMneLlFqGGaM1yecos7bXd9Rgxw3hRIvBO89H0iKOY4Nh1R
3UVDbuvemjTxO1rffMTWsXlIkJyi8GobKshD+uBE72skaN1gd/wx//ZOWNwITxwoDrc/oBCYFWEO
TIwYvKBpHvOE7gOO54OaYQ5w8xMpKsbxBZa4qEcKtPpDCjIwq5UI9VTNDpWUViX/hCaKcImDM3VK
bgJkXpqRI3+8eET1zPJJfFbyRpswyU4K8u0YkdB+4ZqZSbifJYIKq7oLxLDYD21w/1/vo+bF1Ide
Az/HnSeKHVFgvkNsM27O7bUf6A3Fw5EZySWkiLb8403EC6Qoi0lrhqR3FSTQTCBnTWv76UAZfJai
9OVJlkMFhWmb4Xz3hRyFUgn/hHlTln0vab8bpKpROMSnA7XvkiKdaWyJSY5KPrGMRtIIA6Q/xRJ3
b1gMaFCc56VDHk1RQWGtD+07+FQBjR4G5qZ81VfRUTVRqyOMVjDrr5+o+h0tz3XUR8HhnUQdUybj
WoS6yF415nAeQIR+T/zGT5JmaeQ+o0HGhDy307bnA5AF/QWKt131Kw67LcaCHgQAx6K6bY05CQdf
0jSChWxQ0I49+6jn1zf49Ut2kA14gqXXub2Vs655I+ErtJTz04uie4BlRcOq6dPkY7IwqXvA48ws
rKcg/20ElqCSzzN92whAaiB4zbJdqP9vuhHzsbAtsh8s0YezTU1dOA1vQ8WBHH5UYHXp53jitu17
fqkxflBpZunehl7zOXbgjVgmM/lpAwEjzy0Zkri3r8gGJ3mCS7CqrGfE/05P3W1uK+uE9kYHBfjJ
pTLFNgzAQC8RkMD7bEEB9uu2kjgvqlnoy6BhmV7h3n48m0CVnjd9mCf9a0OOJ1pGiWIVqHE5y5lu
bu29yU9+vzvq0C0UsxYQknUhE2D3ZYO2SAXr3bBlClNblrhYs5W6KypRjZ2ZRi+LpZMszV9Ndf29
u489fyySnb0dX6e/XXTMPxSy1RbaKCdVqXq7TfMHt5rNGa+urYM0xRusA5smeA5YKA5683ZcC4nl
Fgx73FKcJU0izf/lzYGAQ6Am782OT9bvhK78h5bGG+jmAxH1OADJui3217p/JUOiH2QRM0MKC5Vl
zbfzH+DuC0dJY2JRHU/1r9E5EVLUqBxgOrXoglplgDwTb42yoHbA7wN/H7aQ9SCU2QwTpVq6RQvN
/ryM6xQ9g3rLOjVE4UfKG7Mmtcetmu2eHOHtpH7PjPNKzOLA1IRMEP42P7E1EPpOelf9SeiY26B0
bblPFoJxULVYjQbSZb7+0zNi0xoa46p0uud+gly7q28qlOAL3WyaqGK//u+rtzcFdDyhhUBz/I9n
WjZ/uXwd19ThgZFn++S+cADUR/tXgUJ6piUeLuc4tPczivq62fN/DPjhnMoKylfY96tJfXopqv5J
Kpjkp/GomWAD0O3gql6RMNLfXBAURqBJohy6a3F19NVTM+ye3c6hIzhsq/W0Xhb1KmhNVPuUV57m
INCCaKPpCrCfsXmeDFYoKzeGzMzw23sTjVJPthBTlRK2x2lADMyBEnDxej+UvXobAj5NtkHBAm3D
IaaJd8TrYzfRAk33/XK/Lc5MC8spxVdo11Tv4LSzxXrznGF3tTzrZz2ubK8EM/TDzoCZ8BOSctls
QTtfZMOwslMBKMQVGfsIMzpxbwutX4qOPpCki8VjPiw7bdCyFBxldXIwe43yXrDN8eHWyXmqF9ew
7bidyas8qFAyCz4rq5zE5Rj01a1dQmZkS1G5QEZUn2TIcR7+eG5QdGw9fJIvNptlFTcHYWonkcUc
AVSp+qKWqDNkXL9XZnLpecHFauItMrsoIC71Shl82MN8TYFyUMKEoqNq1lhDp+61/FozfXOji0kO
oSHASOWYd/57gImy/0xsfFb+8MqYHjqhzq2kLugyaAR/TYtLqfefIVnP50+qvdTbS8mPrEgAsc+x
qq5w8yML/+ocDYiLjljSs/RPuML8qH7Gc7Xt8QEgJrHXaL0O2j+Ahf8a9BpcusFo4SuWXbnZZK+a
Mpsls50wYUxBqormg2574AmrvSVMjx5E1RRTjbe7VLyDal8J7dJpit7TB5su/0Wbu2mSkDdsgk3X
TfG114BDwlDr/xfHJzgTUo0g32gd3oNxFhq+8MSueoCgwu/STLNmibk7lBsl53ooMsuM+3Uqi3eq
OOkacFoN4bVQK+UTuSzH1N1QhSJNOT6QXCkgRMoVmQYhGO+hUivh4+rLPNfSbb+jknTFv/QP2eP5
MNbJyCVKy3NaRhAkhodyPUtRFSdaKzhKaWF+kG31VrCuM+tQ1PloeAZCXqy6VOv8DPHyLvcHFUjG
btAvU6R8fyv/9OQFxTXN3y0f9ixgBr+Nh5tMgpcWOJCwQI4hf2IFS/S11yqhd5W2ACf2D53mxOJ+
IAHYRMexniNg791hB+E72PJfGuu8qKFtdQwtMxnZ7MgkUD2lYR/82deYJnZY6pmCJ3sx52+EYKZo
omYlBHd+o3DvoyyZfSnBz47J+mVODxQXlrPoz4dXAJ/SWa1A0CnsNQ2Zqo9AM/zjZJ5WQiUzBvDG
RDT1fw63SXgPOVIlrVUHhnX1sRhyqoLuKF3SC4Af6qqwb3ED3lP+FFS5As6QrmKPv9/ZwezJMQmg
eUgt/+cqtNr9bgYS+C83ONUw5/3YAfPaUvgDAUnXSLJF41Y2ZAZvKyFJKjjm0iA4PPuVbXI/nDcN
gpB5J/laNMOo9PuKGjBER/n39ZmR+5dwSe6YMj35YKQIjC3nQWpP945Rd+R+GS8BP9tLuF3Y9xo0
Bh8YDnCCazhOpaWmY5SR488zq68qmSM6LtQq5DRpIJz/8iL6QInu2t36eRL0Ku98Yy5pyvgGvW8M
MHnzmDU7fUDEUhlSdSda0txjZPmblsXg1aMBcd49fYxdReO9yt29tFLNo0VfzVt+u/nk7gXhTkmy
IJBCWDTNP0CPFViEzGfFW2CYYt+IxIMbkL3jSxaquRYD+/M2+1P+pMxwKco2b9vsgH7P2jo5UvjO
n6vaceTGINHfDCiE0ji90TTnYk6EfA+RSbHfKxLsYS/otf7rVC77wFvPItQoeVPtuyfTA1/x2dR/
iXnSsOC3rsSJ+cHZf0/tvzPgIdLstifn+I/536k9CEH5NDlxQWrVMAm3x14f7tfMbL/8TKrmuBYK
hGCU+hZcmqj4XX7RzCyTvqFxYuCg3LUcBl2pgRs7NCah/cu4vMsLN5ZwjcHsKJu4RKMB1/2oLC2j
LlcGCsO1oXMgSOSOHIEJE0+gd0Jr2FyTGv5u605qQVVB6VklwtsNlUX2GPdsdardnPuP37Xy6b3f
oaEdJfatc8kmAEXeDOClIwLUH59k2rDKYXkdR6NRIOW7qZw+kr18rvxePahi6q87n5zd1IChOtWu
FmRUQdphViaoVlwN8921wBA8WZcws8ZGxNOWxK51tFQ/mlGbPWndPx/Ma0KmX/EsxOFzZ3bTC2QY
rw4LiNppTYXLIAtPchty1QH4oRt+YOs38OVhFv/GFUwss+ZTcTUbMaOXmtYSKoFIyPTOno+DyDxF
N3fclOjrm3GWb0Y5nE5jnliQa4d3pGX7hKjCI8rYdSI7Yfk9wV8T5E34ycjSV4kFidUOeLAbEh8I
Nvn+UiewxQkxXrBiytaBSkF1bJMnbHxzRx81JUo2EOPaKP25jTigLtLdgnM0cVEvAV92hp3z7K4Z
LBpQ14XZMkbYvlWduaedw2/wbF+QinJvzcVek8nrdAPezWId9TWEWcBy9Zvb3UbJdSa9zJ411/a3
zQ6bQtGYIV85b6ySIB8GbkNZsa49npeGhaJxTz9h8yvjoPC1SABNOni3xhUwBx/kJjJTKUR8126a
AFlQxEejC2drpmswzbw63g8LNjiJMaNkGcXT3zpgNbMkxAytrAp5+YlyAIsJEiwTUA+R0M9TbrHR
ZuvG4eLmywHaC+pEdZMR+FDyLFueHlD7ZMsY14EQu6VOGb5seTuXBpqjxzcHo1ZhYO4Eww/WGW/P
KM7U16xnP7xwd0kMt6jnSR4vYqLF8EkpENIhgEN5w5OeUc0Q8DpGM5+UhowN/cATPwf7jrQOew6O
WS+ruQu0VIaC1Js2acnKnfFyAF4IxRM4Kb3fbF+wNTT4suIuNlsVxVjis+hZrki+X7Vqe7hMZ9Hf
UCi27h6kyvy5WSjACEuwUv1Y4huJuRsLVwgpyPMBmROiuF3jcCoDouqgjaABgbbfWlQ6d52HdrF6
dl4CBBZHe/pkd2ArIgNaByPr1qaLPU6Nl115p4mGDICkNbvHt6A4kEUan5eBkrF/fV5TCnt4K6d9
eRiD/orJzffk0cAko6qIR+5F4EoQ8CzE9nPmK8GO8lStsuNvCWuvfvDRLcqdYH0wW1mmYj69n/2M
S4DzjrAyUHwi8yIo7qwv/Yo/TcazwXKGOFb/W6slzqLFWcuCrDRPncQykXb9o5zQ7VteiH9K9rHl
7/MIdMnoOCMs/fRTr8hdvSuO5beaq218WUmDI6vXjFbEVVT+DKJyL7VLBtmP7nz6tfAInmkjD5C1
oG0guXM6CuQ33QcnJutmrrAixd2uB1432NrVENkyHNNeNMftQe7xsXPbvmYD4rF0+bvqKeGM0LXr
ttx9hBEW13Dv9R2TjhCa+zmb5xpJ3FISiA3xf1PQii/GtsPlmFFzrhn9sngNgEl7GVAU4vqGvN9v
aZewoZbQPZg2O8mEnfTWaSSthKDHkbooSTDwdEDcCVc2Mv/ReCNNzJUIZz3fqhhy76JYULOsKiAx
f5+8pJcDiPEjDwSQ3mTxeBXRvIDhimdF49vOBolDEzmfVFrPBAq0gJSTQh4/2/Xr6MqKEIVdy+zr
1MfO5frADtoGyxv0KdzvH842p9ndT87Br2m3fyNVC2kyKVCCZSCO69XsUgW6hWCwsnjOeNgEYKZA
eT0ictyE/gjSRT4kbRzYeFCRV0Un6oSH+ZxikmkQyo30p56w3IfTEtBeQmKUAuqA1CqBdS/Y1a6X
w9nTvAb+p3ER8JzEMowIeWiz3AcKxzqvGQiTUi1oOmy3jV/swG9rTbNoVTHDibUpxm1iUZeO9yOf
sCTWks8/kbkBI9ZCCiqIWwjKefGXJBldCkEZINOjrYY9EVRdTTNabPKxEHI4DslbZFTOZT9PMTEq
0VA4itjLfRTr2HiSXuMKBrrQrydPKmxXl/JhN/npyF2zvnGcEicC8nnGnemVsde5WVGMYjQnAktA
CKV0OmB0R4MVlD0QFjvrXr5VljEUnCQGUksP3noHWWFDFhvO75iCHWEgUUQCfKe2DHrUH5Sx1Fw4
krFXINh3R7OueDKNtTrIm5Y3/2VljOr0FtYO/MjJvKSnerzFDdD0sPc1VHgbjopmQqYTXdo9HSqG
+xmsXUCdo6yurNCkIFZMMpSVzOqQ+dIv8mP8Enmm3fSFlDRjgwwJp3Wx9uN3FH8TW4bziS1bnK71
eU8JqFXKksm5KvJy1/6BOsJg7FQKYJ3BWs3eBVmMMgFAsayZAvn7XGnH7xJZkX5cufKAZiyqmc6b
mXjpPMrk+crHfjcnm4e9SPVEkRaNwZqhvqU783mK0XiImgvJRElQRaXMRuL99c5cAVuN08C/lEed
4g6HwW+hIQCABQIRRlN+xBYvSVST0neNTppzX45IbL5gDg4RUc4S97Wlzw/wDYVDGlrLHiVIpKwb
EE5/KMU+yNA/wYUSBJNnrkA/NdDNZX/jagwCSl3rm20HoaSIpOQ8woD4qt5+5exd6sbTBa58jUew
eDMmXwGAfH0d/dBJLx+zGOycHIGgUOf9JYzzWoxUomsfG0vg+bxWRFZgHSwu6XbjA31qli+m6f8k
6fpsiAbZ/EQ1Avr+G2gyrAk0efVzl/2AzUZYJGQYZpqPkBRy9Jmb70Uoz3n4RMphcxgCTmOloBjS
TCWxTYlyjk06pe61P2flI/iUBUwWAMQnholaU4Cj0oHGs5E7PSmFEC8UnFVSeoVakv2b9bSZV9dp
fHokFqM4wHKEmOx7CF3zuH5NRJTNe3rNvIyQ/WGlmsT9wiZUdd+0uHhOlmSh0vQxxgRVyVCWxu7E
TuZmlHP9EkGgeTXxtasj+n4HgMrcZJm6W/qQ/GrEbn5p518UdnNiJiv8yq9TBDUX2jXQDABEoF1B
2SJcK8CwE8dyi0zr7oNjG7LIrcfa7FljMtlBMCM9h2A42F77tVEgOyLwStAQPM4obOC32ktT7QEf
EtPKrx2xTsf+IUwSu5itakNmgDrrOjMPHok59vczyT6K3GhjssiwrsiJF/vW1ys5BLooxOa2wo9j
z2Xb5p4ygrx+frasoRggoneKizRvemqJxcnmQCLWS7lZNnBx4Z1xfzy2NLWW9LFRNUoeBjKfgBd5
5cHnrpOBxUYH0Dg/vHg0mFp70ImCtV/kCRZY6Owh4dgu+dzY0WVrZPsv+T3vYkEC7P1ViqPPL8bp
qwpHaLUlVKZ7Dcl58gW+XILkLs1H/35FpMBPWr0JJm+thykBdPkygYFduR3/mZAWALOzIfv5VRoo
ifiKHWhW+Su+8hA7LzOvbw0A9bMuk+KMjbr9nnkQ9OmNAdrvdU4t1DcArtwt0hTM2+yuOnG6jcDF
6qSTZxy3sObwv4aPJmjz+i+I7AXuRx2X69b5m6Y/QhognsvorYctgkVktotbhdD33lfKaA5l7qJe
hq+GOxRs1O9tiQidUDTU0cB4M8NYjDuWROzP8v/Z+/CdlH5nvbaFKjT3H60PA7nEDj/5gid+UXnS
D5KZn/JYDXmhJCY8azBX70ooQHRvQ/IJXQP5BjjryObIly1P1zmqJspeHQyRJyn15+162BRc0Gaq
Zs+ilbeSSAXqwfW9p4dOmR1Vnd5qbbFtBV00Ln5qHyxDE9+ccxQaMMw0mDzQQuRE8WzW/GwZI3X6
6uJgeicfJTDvzvDXLyTiiwadnodNUbS/P0ljxLpEs7T2gCeUtd5+458xrGCrBjJixXWLlA+PJgo6
59j61B23N3LLdxONQ1lB5ZVlDwqpTmbBgHIcITOF+Q1dT94Z7cu1mmJZsOPhKMSKuudOZSz0gdZJ
TP0/x/PVU+HRJknWnSgTYzHNq8oEB27Hc7viQjg5Pbs/5aQc0OiNZlkeej9wNPBnAqhRsG5aeYFT
GeXYJPaaWTbGYzrs/TUv9LKXopcU41eSouuyuTeHEr0qjjczxR9tjJUmkdZZEaLI5qgZrwmO9Wf+
6V6Tok+aa3CjM0nrZgmqGjtEtgqOM1PAKLNCSV07A1ixu8OlhycnYihaOwt20JSCT5c9ivYPMH+b
Pj7VwLOmveX+Wlg93s8B3QVFPbYxDamoZutEnv1hshtFvzVAnidlMsjVQiK8BRdNVrbj6icLYrcL
e/9hYwa7cMGaZRfmB6ohadqmWEVE3vSU0pOfu9W/5gCAQVC9aHamxTh84mdvWCkGDUFSoIAx8un4
u5DlPTktR4omENBNGzJvoSUpbH3L9YZQaCCJ2+NqrYIm1iXx5vGqtzaoJyYWTU1PXyXC7PAaEW5f
LHAyoMRExHbyN+wuxkFvsYifgb43yMhyO7W3v8OBcg1MinxlO9/kMzTC9LvRGjoLNp50/9g3IMxU
+CAMAwZU5I2/2kNNtaTCJJ2OKKnjbw7u3NdOeIc2uC+gZBA0osTs52Au4jhM8AP0D8AuQVC3HDmi
mzsrOY+V448+yhRWiwApNSB+3IcW6uLqL66zBuv3AuhkjOQlUutHF+qS7kmjeo2vMRtEZpEZhRrE
ArsJKucSxCWitz9wa7jxwkkRciALqSkIFjM46y431zpwo03Q5KyXTy/+5yoC/2wwjIU703HhqCfl
9IwrxyrXnm8MrJZuIUQa+nWUrMHHsGIX5MmmRTjoqG0piPX/2a4FS9Sv5JUdf+uBCHjdZrJ+Mibk
VTntfgDkUZbuQTBIXgTmbvAmMklRFV4sK+eCjjK3cqdUma9dk2MW6CmJWlgemNMrRV17a6kkNYJU
m9kgslfrrJ72zKdiPGSk7aQewfCx1/LC7Q4sxKpUtyDhLhrb4RvBhJhB5ymYrfE2wgCplp/U2PVV
oyS4OOHjQ5U7ZILyOc9TP4tAFHrAYGiUZgls2ixnAWaho3ul1t3BW7FFB2fuVodQkM612qAb0jyw
BPGHi8MSsgbURdR46GdC0KhZU7yKPHiszoshEpNDYRviFLUagUAEahX3AjFrKFfFs2gSVGrPh/jV
I5a54ZTsmIk0F4RGPved9x85wtcvdQTx5KnY5+RJNbd8C8IRq7uiZIQPv+a1RF9sbRTh2MI48LSA
hwhlbR67rymU48NQxoraZIyQDfp5sawP/GMFyEl4WCsAYbL66mbBAPKTfy/dj+Mibg1+3KwDn53u
nmb0El9R6M2EDEROesh1ABArY6S8POje5xR0JSAlQgrezhtKqr40KDnPICtHiQOKZBZXgrf/Xyok
qoiusXHKA2721BJ/5+zdtm1ZHnN4iwJh90cwIUXDvaEWSNobKK4di8th8lNq6Tw/XFIlzBObCspD
c/bQ2uH8+AxsnTZw3ku+Fwgfywa74x4d1eiMQHhPNbvfwE302JxIXrfa4hr7RGXHatI84qpendS8
S/5BvAIfiuGJq7ZBiFEcl7u5lSk0wQ041n3oFmdnWf6CAriBFmJpD4lHz2s4ynQFeBPHOBcyZEj1
ecyrfo5bhfmhj+nxhGEC9yHs0ELskf46YWbWUEVNXAKBKGK/XKyjGuAVEe2zD+VwMJwPwL4mOWvR
bm8FGdRWHWkrt83ke17tv3Z8YrIRtwA2cVGs0FhfK7YsZUL43uYyNl78Y3uigXM4KoOhaIuHv0yI
AyNMhPUkklyjgdrlHz/1TPu+ET3M+YqdCQr2CtvtlybrTJzA3Rpems5h0RzLhkmfc8zj1E8cWeCK
DoRZMIW502q1BjtK4MRonlNWbzfhoHyd+Pw1Btv55W/+mlDo9tQNgVJdSFzh4zrBkzzGpxQbfQx0
L0JkjUC+dJtkSTqYw8o3Gbagdk7dtuGWhEiB+cjzX/KTUgtVUuLmyUrw9KbN891cQ/OogF1bX+MI
uIx8/cL7PyAWTtXxebLPm8kDKZmNKLon+n59gx06RlO4AaF20fVqAMiPkE4DiJLo8lhndy8MhF3D
6Cx/A9VrJ9oC6X3bT5bk8FMd3RNYYtwqvNqTBwOjaCplCOusa1EFpT4PJLaauds/0iNs4CD8dHGM
5xXkULSLLcS15SwnofM1Ax/ydJqjssHs+ftqDFykjed+eY8wmJIn7DKGqwsBZeKnRBVkYNo0rt/i
XTCTlksynQyUK1TwMk2rV6j7vz5N5bteriF7GgUlWkm8h1om8vlAwPs3dU2ZmQUbP3iyr70TC7vh
rx8cHFvO/7uIaLHyNaKB72q7TsVMLgenctP1iWubmZ4VJViEOBM9chGzkkFNnlqYEN2aM+ONuSt3
b4ypwpowz5MFMS8QslZC/uGBoKEde2Ty4oPL+V/mjtdYcKgmgAM6iwBeMTbgwsDHyQmmylxW+2Ag
Hw2wdrh01GBXnrw+qLmTLCHbqlbfpPlEujj7o2/nDDNH6wIy1nkqKHsMKXeMEk1yxegIZNS6SrZc
hqI3E0Vv+6I8E/uEBjNiI7Ons/UvNdqBTJ2/GiYRjLhbaDW76v9rqGoi7Sq27jUf7U+STxBVwB7I
4RRzG8kQcERmuHEYODF7LEL/TNzJ1COnIozOPbX7rr/Z5npFAwXNrevlBRYA7OLegrK7nCm9C3I0
62lbFat8aAOOgfDjsH69Rld5PqC1JuD4bOHFIy8FIhUMsWLCLyGvLLPaA0EAGTZAKUjy7g5w3c9l
CRxkvIT1Hy6WqrpsPjF7+DGB93B5hikzAP1z92+YCnFJhcUUhPzrnWxUug6AEGrjjr+D9fTFv2DE
GQck3xc6ONUsX0mbdvWxJCrxB4ew5OsFoHAF08xpzM8UJIFwC4R+/C3Gy8lxieigkhl9nv699ZG2
JXmyoLjuTnJoOHhJ9sMxydYRH+hGPTQWyDAyEFz6ajrSVVbvS/2rsH0ZqNfyV7VZsplJUpFZKqWc
k+k7RNXt7zqRJWV2f91tznTmNuD3MYWYoc+FFIdJ8UGex0G9Qrl35J+rAYaw25cxnamwneXb5Hc4
iF2bKoiCaK4IrsoOP/4EXqEreJscxBsTvpUI5KuRID3fsMJMdjIChE1kRQXWG+DH81L/dRqgLYR3
wDxPSt9sglGxBDKvntMUBTRWLhlfHM55diVQ1kNHYN3jVRgRmfyWP5qJx81/ug1pZ51NntzhOqCq
GAuhophWWr8U6kfRsnv9/TUEBP/BPV3/MXcWWIR4AcvciLWN8VDenqV1MVmg+337o3NWv2ih0fsA
Z/0Okcr7DcP2RgSGqJht1Nb7m+fm0RSzfOZVu+uQ8L1V+fTXHnNNP3kY/NLmbcLpdr9RQ8uIGG0l
srsr/LP2UgucTZrMagTkJyzfZ5+X3SU9JE+MI7gyLVpuTz6t1gIGwYyLk6LR3Sqkje9U+L50vb4G
W5QC18fQ74mFqGwWRLiiYq/aEXtkrLH6Z4kkFEmj9kk+Y3q+jPp0K+xjUpz6LCmru4YlDoY3AB5C
ehpue1GstC1hOrCg7T9jcqgT4zk3Ux9/gez8IkMl4W6XWETY2IZ0nyFUy+y7u19svUrMxkR2pvVl
45VBQyXiumEGemNzhfenBEeKitk8//kN+W9rCfJ0JxVCHVOM67dEjuNNohinzz7pIIwGMXL1lLaq
+Nhz96dnP6ci2qhCZ0ijk1r1b4oYQ1tNcb4i5celw4gfXJMO6lXxG7NMwiL4pj6ZUTWvMEOKQg7R
ODWj2RppcrikzAKTOY96V0Jeu9PMbPyqh0i2o6LjapYrSklGGZq6K8qpd0vBsfkAsCRoEeVSDeHt
ksaAth67gldNLn4b9rd98HLVM5qPkMsFiZtEpQgpL3ekYCfVJzu3zDicVWcwA919+WuD64YFkQ4J
CvZ9+bZWLhVMfv96KwKUKYj7IFUtMFOjKP0MS06hPMEwEFF5bsSQHmrqBld/FFwyWvHaZ3/h23Tx
7dKJETAZiboSvFOLq3mFtAu5TZxXGEov3p6WlfjzrkFv/5rftUyvBdLrBA7nPtvwF5+JDK8IfB8w
SlisNv4/rSFKt93xQfliAonnxp8+NS6y/AcKNo1iCw9YiwqSXTbx43RYVjgLlCTR1hhEblHhWLHL
p9WUccJ4J7XPIgoTrdyDCXhCkfwIbVBAj4ZBP/1yLAsz37CveldKmpWI5fP0ebfmhIuUV5Yj3dKQ
r2xD80OLXnMTT8GZ61RjhDpvFW8L3hyVLKcROeVRDSAVW7+sZk6I5LEL29T0wHae3QNh8oo0cxsk
TU76WK5Nm1Wfsj8FHOg1qAjbrP7m8xFONooXQ+tc9KlRXfBTmuAPqBD5KvQgCyUwd1ZOAvi3brsY
9yJUBR+nsStc/ZpHF6QNipgRokNOGwRCAal75MTCVbeTtMr88k4WC6y6Z/ISaaVCOYolq48dQmbK
zKfLAQT00iXoF36M3CEXl20r7PwSRWbMsLqx+sTv9fWbfVGMICCiswEE73wAwyUoXoSKiTffXimB
Q/rLpp8e1Lvw1exr0PYT+u0sbjqVzmkOYzvOFhGQaCh2ZfL7UdEQpn9JvCKmUWIQDqklbXEBjegl
UTewhMIPIJYE8ki4hj4NLpW/3HJYcI+cSP5JVnGKdSbebqDxJcQI71yGM/ByiUBNPP1RakBCMph0
iJoE+EBT64KsP2ZQSv8SDkanxiELGDTGrtVpsQNc9KPPHbU7LSwHj5RyfOtWEdcKSyp9mgRzJhV+
cIgPds3A8dVPmFslJfC/YSAnB8X4wEWqxeitbZzU1CN98kQtwIJN4q+Kze+Q5YzxBkMQ9TK9HCG+
9fs+Oz7KhY7eNreMQ1A5oX5durxMKBwr+Y3adDezT2IJe6/1V5S3SCI3jBJ4lfQnpfArFb0wc7nI
EOKJnjBAv94Q4DzYNTUK4MNZ810FmjWT7fi12nXd/ENa/zOki7H2Fwkt7OfhAQAcZBM5GiyIreQU
GCeulr45lnX+4Om1JMM+QNhCahHpQST5X06gNYVD3eI5RyTjYIIkB4EVyEFcVmtXIPkwsg8jVlWL
XGjYcp3nQf/F629Xhfut+ULqbsfZo4K+Cq7mMI0oKvWetvCrnzUqfvHfrtLsMSkuajTd1buzdq6s
4eLPe1LReAo5XWl4UXFDc43AjA6eVFqeYmoHZoLUy+ErbSZQU3qXENCQlRLnltGKEiPddgEclfZj
sjoj95AO/MQAUR26NIyZe8IYuQy7Us/5M0o2ul7Ur/jB6nS4ZLxbmgZItYjPwy6LFZS2xP4HsDcJ
rlwb5GyiAymC+C/fVzqGu2OXOlpmKOd495iZarD1PKx4YZE5MYTZBuSwFTQi6NrMyXQbJuNixrGD
j5VjM0rtCUg3xKANU9sgiI5Ec4XSHoQ+797wCX6a8NoUcyuxkTR7/QKpFFfhPFm8bLyrlx5QhlG9
SCZh/oNMuDw9CygrwTRsQMTmRbmk9Sc43Atl3RaS00trY+rBQquOGtikbKJL1/BXCu0eErvZyk+E
3mXMth1W26OPlR7vJjiMZ5Aaxbyi5Pm3Gcg+64cIkKZSsXu9BecdUe29EopGai/AXwqWRFeVxb+3
GHGbkrNJBp1uDYdHhFPRBHiKVHoGnPuJpKy41/V46kt7a6L0g5VD/oKoCfIA7el/AL8WiEN/wCNC
/T+e7e+OJKAe+7fhHL2Zcp2mTP1zzTxQoJKC7zoRNbuHe9GZBb5C85tBo/Bfx86nbfJA1xFmd1t2
rMXL0QJQQQIoJlGg53yKf3kqO6kVVa4kcVUr0Wa/WazxnhmBNkex5FHFbMRPGIZb39/9allKgiW6
sKZnnGDgHX9oNpwUrrUY+sjIKUxO+4jc+inkUHbErbFkfCcONNf5W1a6ZQrPYKnIVXNbMxR20l2H
9qZ2hpLpL89dcOyVhO/I2GJnAasSDjgV6wrs05zbAJytdfIZgvvN4BYmxybHcos4YAQ9P38bIUMc
JpdvCOPJhw3QeDdDd+fBWPOcWE4pSx3NOpa8G2PrY0mgupFYNxZdyqj30qLubrC5G56RPC6zbChi
Oi04KpaZQaxjyZ6YFAlOHLa8yR4TKlIXjqSMpPxBmGSHh/uABC1ZdqbCpAHAkbe2u7I/2KuYE5m0
oP6Q6XKXMwDutKu0mka3Fw0e9sasyuUFwx51MavSi1lqZPkC990IWY/+AO++ugyBw0tPtWEI4XiB
Dxma17VuvayoCIczSMEtpCOssy3VgRsiQ6Hc29DcbXkAzS5IXvfbpYb7TWmaoQP7OAmAbVw88TgN
1sVd0aV01vJxQs/KfHQHbu7bgQS4SUIFJUQ8KVu85rhT8Z6wC3iE45SCKV0vwY9gApjo5YLdzQH0
8eu4jeVdScTgL7hRQmzGx7d8neO09lBbYE//Xu5+GWlsfaxuokgyWOcJZ02M8Rtoag5s9ghBhxnf
Hv1RVzASgju3R+/AEaRQjU3WcpeqrBVXrZE+IM32mB8F9Fv0+RDeYz1tFWRdKgmj+L7+8jsF1fTI
+7kU88+qYTaCdbDjVYECGTwGim5UqFFua06u97MpsWvhQgj54WmUugXDg/6+RgojHq9+hCGka940
3MR8WjLkYsXxkoXUXhgrITTSjB0TRAuP7nwV3yr13OlmoMcm8pLeoHLp0FbT1Nwyf3ycDaJXDrfm
fhaEBTcClRH1yAC+ZbFSe5xgslqP8Jw+/YlNsvXxhcP9oJJBF26YykfWfIVqxLFcXbAv0UCuErt8
PGQ+s9wIZal7+tXcYG9DsOwsQx1NAMl1168W4MvlsKpx0yUULODQU9QZ4sOuBGxMcma5EWgY8jW1
138rFAXN2pUBHpYW1ao5/pJs0Zp85F2OSnBoRhNGmWQ71C2MGHOY5jYbg3Wg0VwOdeHVcpmPU9+h
3ovQPrdmRRqksa26wSBPPW48eoU2WPSOcKfXJiQZt/3ndQbqUrlIZ1dQLS5mMHRNPmdax3FsWq6z
3xROp76jqRak6xzL2sJPQ5RQ5enMGwXZwF4m8NXW9UvC0cx/hS3b/c3kaoxBEM5NGxG1QSytyGzb
jj+c7OqLgoFGQs+72MUSyp/9mHD8evGdREJxGC0zajphEtM1jI23LLVkr0coT2bAib11IL34nCsQ
3JVT/ahgcCvXakW1jXNNLmxbCG08JDitFjJrI8uPtOkWcewdC5mLDzQX+bvA/r24nYHGYbleM38q
xQGZlsXmbo80UHubCANhu+jkFSI057FriVTGnuSR46hq4As4rb7LajCu5NqYPIpvne6/71OZ9/Hv
6fuSM0VPYEWkBhhr/US3/Y/pXDnK2cZXZxRrzc+7GR4bDVZ01YjXUWCvbQtmJD76Ahn1wnjvHbpA
wusVb2n2xZTOVV4waZGio6SbaRH29uOzo2V44MJ/ws7W4PMBDssAvsk6IyLKwwRaiQjXsOs996CX
v89njGZ3GlQUB18/z6CxBJKElPxtdcolg0fAnYfdIWKltzkbGSYsp4ALlMIqhWNQ1TkcArd+ZV0m
sAX2OIhYa+cX4eJV+ShJziwCXGV/fEhkcslACRnel8oo31NqpnizuC5mQiQuqRCRFVzKV6dVIH7k
HpZ2wJiVFSQCCmQ55gVkXgsz7eGUB8A8Lpiocl8nm0NvcH7vHrMWt/K8PzhEKb63c1WAv04QQR9z
sv6EMd+lft/IHwotZhQ2sB8cPUvPvrOCrmv2vaT3RDsh8GYXBKhfkXk7a2UIfS9gAu7Gy8ThV1QL
nBplZ1OGz9CA9SNIrM+kBTcwh+DGLFozM0hVq2PAQ0Uj9TFBI0a5vkbWmjkUGE6nRZAfbf+pYH3Y
WFSTGM0bD5M32xXtpEm4mDovwq9tH73EBIQMYZi6GEE/P//Y/KELjQg+1XibJAxxkTt3p5OcvVwW
kWciNVMmFOMm+j0VU3Xk2xE/vA2oE7af/ZvfFHnwJyEPVMeczBptqkiHEkYWTt3d5GctBe6dk2FN
9O72oHCs/IowTzzY8uWMxCeBdzZn+zFXMiVQZA7gq958A0HAglgZGJ6Rg2xTlnV54bQmlUVII3zz
Aty9YityzT74r0ISP7wVYGqrKATitvJp3RCakK+9ON9dOt2WACg297DO5tIgZB1Vhxmc56W+MmGi
T4ktTnT67ahjm3YDsQyC1KrP3mybHe3DEocl9zWYd+3IakC6FkHmBU2O5LwjjgnsR46sNVhFMzsd
G/uXl7JZvfBCq0W5p2nO21rZO4NmN48yGr+j0pZC58VIhAgc7SiaOTlnQV3+3f87x8vCK41o7/Be
BJBI8YhQKdJCSBkiHdDu0SSZIc1jEeCCkAjDyEHRNsc4QLqNBgJOXLoY+mzul3jDKT6pHMhcZJbL
TRKYkbXl4aptIrKCRQNtFDI65ww7OBEcO6RwMv0plaWGq08nFimSGi+zQVJ1QYzSPBRmFbJUBO3I
s2V2NTsgxUNS07cULPyTdvs7o350KyU83LSc35eJN9UitDvpnXLCA99TTopjih2kDzYabzYpX1HJ
I+4f70USSHFvdKhCIfWwlp7cyS6W7Y/edvA4KEW96BicuwQc2QVlQqLbKHxruSTK5g9/NFjZiHfX
eVTAK0Aay3oVI0KyTlN0t94zSF9pviMPpKQkCLY7NpuVaElkiSDLlIRXS4JrWZNX5wWGFOdgD6x/
C78ZK8spLZWrvP0vkIyx8qSQnJqvQ67yLBczXhVNDTM98kPgqGFJAHknQ+bm1pwHveqJz3xh6eMG
rMU80yxSfuqXHfn72Lc2321Evf1lJnIX2a6Bc1SYYPFZcnHd93f36mz+I4n3R/DuCwfezHZeB5A1
CcNdiDykW2WAXxBPHu3MqMYQvYgCKqWn0ieWPMpXm0kfhfrD1pxXEaSZbDa7FuPvoMbaYvdH66rx
ozI9vcUHLbGIKhc8YyN0lOZXiXMDvSLfS/iAg1txax3gtk/0JoHhIr4uEvSAaEaz8kPPkKtC9tei
VoVyPH6724EDdOTSvxikgGegyXdGHAYiNZaiRhh7BRsi0YmZkhoIZgXusL8dPy8acr2VZvc3RThz
9sQz83rE9wu/r90BHSjAnP+yLlBoICw8jhJcddrzJpAsqHeRLcTsIXo4ylXD0T3ZtihUf2bxuGY0
+0r+Zah49hTTP+pP26Ky1Tlc9rlAQSoBSV1cbuHW9VkHuQhTnfVOUfmRHO79CQBLWhYqn8EChKhQ
2Ne9aId37tJ9sytquWMVjNjT3pjdi5W1wzkVG8xdRKXMaKbFoJoTD+0Nj5kDMnmf/x1Y+C9TpnWP
+M0AviBXTC1waZ4IITXIPCZPaMYGEYsOo9z9ShqdkQ84+1XsR1FQ09RXcPsYy2iIpNtRjs0t2LgV
1OOr9rDsrvr0o5Ff39sFRLRDJY/m1JggtqpJKtHtfZvy0YiHNYDFX01bSG5AUfEdKH3lPFxgSCek
B/ClkuWzrS3Iamn1OA8w+oWpwVjVmQnittM72hyGvH+SM60v/uvMVV6P8bmcy5C5oFXnEEZy901o
UEx8My/TVjDTtQpqtd7bdg+HW9Y33HltaxbT87FrWeYH1JNrRVGoUD2oyP4mO4+JuyT8BJOWUeGx
5Dc1pnCPH6jS8bkt3SjhrrsTEXS3uX0sLKIqb4HPQhxlthXcvetBEWk6u/N9TDQ0m7ap6GSYh7XU
t4DSOWoqdWCa2nYwpiU0aNcuCA8lqHWTLmOw3jZQii/BI2Y5Z10c1imA6sMGc/Kh3Xm/Y2qGvIJo
Rg7uoq4txDNJQHDdL9KQsM40WgC63gCoEyr0LRUAaf6gqo1T33I68aIKxaYZ5705HCeo1hu4nfHO
WqNM2GU8cbgOb+83k3/TwojNYAqm0F+wC4Pfs6d6kUPZkOGsBgyUCl3dAzzZLhPcjpLuDk8gObaY
wTLEOkZnhMjV/S2bqCB0oibAYM19yO612857VrC/1ah+COj6e85L6pzs1ALJqy+vKl+l2l6rqirL
3xlkaFnZ1TwlFSIHbKTVv1ea4TwzsS6vVHh/D42M0Zj0WH9eO93NmPEHhhsTbY2n6cG6Ae4chIaf
NOwApvxsSyK8CBbgKtQJAz4ZPNKsGQAQ306cR63H4UaLYM3+BrOxP6KyeiOrAj0bcJBC5rmFq2nu
+hO7okHioP4h/XXnXY3zFSUXxrM4l2rr8YS7Wa7W+G2mJ20xhgN+hprRmJzUc2kMhwseZqQxaymt
8gTw4PK0rtOZKimYzTDJOhMEpWxfCO0HRg3dG+/IVayQLIFLDX4IroPVqNRpVTx8ggi0/x43Q3ay
xiqM5E3UJ5NwPvx/d+GEH+h2Tyh3Wpu3dxjoYoDFpgJfCUxV9Wb+8uXLlSv42GHfHUuFP3uv4gz/
VOgk/Cs61c5FYuVXxIwhqCSYabGbEUM3Ex5BlTz9Nkgu8MAVgtAPZcNBSeKY1gwxx6hKReQt9UiC
m0wDg659JcAMla/qoJEm5hdhZ1PYBjBSuogc5qqXRyxuhk3C99t8YdBOVib8Z97uryK2L38Xbpk0
q3YprtthXDb2dhN8btHMbw5HMAniwIplTf7NP/Zp6Lg+o8vtOlzED4j6v0n6jcU96g7b6RSNEhhL
yvKhmpU/5NwJj3EsDYHTj6732DMDG9bHZnkDi1jzmflM1cBOxhqbTtZTYfxUQ5RDDAMDIV2Xthk+
wC78O5e5OjsHt0JZ4S5koymGmScDsnv3Rq82IBOwUJ3fl/Ae/MnsGbHHISc83xE+42rz2IqXlXke
L6QATmc3KMUUIpSpsydJLuIp0DYdX4iEweR9hhmM7YPFmQDUbFmmKs61rP31j5EAubRvN4sx2xGd
0gCSYy/JamYKsYbWAnU5pzk/wXxJkOdGLq+L9jIxCKxynltMDEFE9Sk7kiM7Ct3iUirbZ+g5UaaD
Xd8gY/1YSTwkJOwW26ybvVfGudmrYWF2qRefabB9qRIyp2584iRptL+hGXWlEhsiikMnlwnOasRt
L8QkZd9gX2j2ScZU4W821DzkUplR/y5KzXt3amkjWVdprwsuMGkRD5kGFf6AfLL2RaPjY5bcarDv
cDQfBqU/I73jgTqJMMhMj+EwhiUIBZrIbrDlg5FKS+eAXN5CasvwfkoGmOvaCwODxHOr+s2x+ZFi
mG4glR2fzge5E4uz7kD0hzi/F6yTIpL97o3uuR9OkpIHKYjozMyRSvzPTH2PBTJjDvlA5REyOyXA
iH+ALe6URz5CzD2OIYe/RGyU0fPkjgSLHFqUBTmynM34Tfx98uFgl5FpS8EFi4MEHt5Gfq5ZnODw
G1qTq6QWcEzQiJqfdzfHnwWoShl0FSFHh8bfpSfc61MgGFGduKUwEQzhrgyRqWfMTWfGPdijq2EA
ptDaXIpNFeYknKdBp1njQZlDBQUL74jCmIDfMEG02QXWAvT95kuP1ZWUlEYtXyx26sYFb3o5IUep
R+NHFf/npuyGD+uRQAzkISuMuTq1EqyZXLe8cb7yXcDuF1YmoG7saWOtaXNkLSaflbM3pAlxEsrx
HpofUz/ZBYSPdXdyz5sEpvBo1zLPXKNynKjU2x9TEpL7qDnLa6kyR7Io8Lo3l2aUGNuUM/crMJ7e
dxmKt/HvO2US6+qOvqEUHm4kQioaa7e0Lk5pj8th1ISk8AZEs92ogiuJyb8uNBSKplWElNhrzD7Y
ErBjzPppjGEwMb0zdeEOL+zL1goUF6HJ0GnJvWz89flcP8btHOoz2qIy3wxk3elIbLACfIjnYj9m
6Ewv13HfcaZSECmVGqJLs4whAk4NMcQZvqP513ti53eoxZr308DRDI36S2NpklPWot727c3mnAvD
UqaHcrrW7vC6AfYjK8987wFjtlLZiXGhSqS9PkouRiCMN80EHIOHhPcJbkitfiPIUGI+lW0Fofgm
L8DQt9qYrOkTOSrY7EUE56VaEOxZPxtFNHhDZL1FnHQ6xA8ACjjpaic1tEWL621vWdCNV4daAgjC
JIzkOKSxZVCQMQ1cCfOEPnD4GuyGaL7Yp7K/3rVwk/JazFefXVOD67vnO0IVs1bg7TDxwxYcddzZ
QAm1BlmEaH/mI3NB2Fu1hGAYByMPhYNDb4DweLm1LvSrp7zEhhC6cf1EYr7nK7BGTTn5ucOEQAID
OGY3UHqxiGRon/TCP0qU89vq6qXUv6DMHrb+ptksIOZl50GAvUoGUrBtswCUxfeGw/oYC8RpI5mq
zsmvRYmNZArxHHBqKgpZWM7L9tmJ91dfDOE7sDN80AJFfVYM3bAz99ePwks79dYZFku0IyLCjSbl
tSkWwM9ORxDTzh9OVUo5smggFuvMK1ayXg3MucoOsqhjMFLZgmKakbhhsvFeFPrw3n9JDTBBjyY8
zAWEhzHEQnPLSiUHZ87MZokpYnp1ZcqKYEAkcABtfME/Jo1NUatpAMsM46aljgolNb+qVIlLx07Q
TC5UJdB5ZhmgF9QPc/JY+oh6L+bYsGra7gJF9tt2+Ujt8k8wownCwFGIaArOLliEsZetsSxyWVzd
0OhwnAei9EsedIRHvPEwTe6SQGNNoOUqjXwdNeECNpk3z6pxBUJI4++HJYcMVQ2Z1lD/bo5H37ku
VE4ZKfxYOmCiIOCntnlyiged2ZVdhXTsnRVk7f+QT499/+KRQwxsLYpS9zPbwrjtTCYYSQVa0tsU
bjdTqFIexil40SEspQnQCMouuUrn2sIWVn0noqY5sepfmZL2IveCzUD0pKdFhe+ldLGdDD/an9bh
DsCtUjRBFzWuYwspCQeFanCZMNI/ZeGcgcSIvKCxP5pRRPGI8bxWnoSN7DKI1ZCpIO+rtD82r0p3
gqfKblXWJvhOYOFSPhW7CsgeX9Az5Ve4ZjpR/VqZvPR34V81nLEaRlmoLVT0XVEJEXTdJU0tM4fi
yKst84YeDGoXf6odVmg8+AyjDqlENXF5teKxcK/08vD+jd6d03rmA6XXxrGxA9/Dy2j6m8ITmxd9
nWXsEb1wQBM+cYmo54JGPw+SVq24e02AZkgiQ0Du3gmoVR7OgufU+7NkOgYvxQOwTVFwmk0DOfXw
dbrG+scqDcp1XV2RVZ4QqJFCQyMuuIinC65ByYLFkUfovklf2dZcEo956q1hJRTXk36cC4haRV90
O0sz8ahBQHtSIE7rrnlQyBfL9h4o6GiB18gIBy7j60lPqorPCt10CzM6U+OmqWM/0wox7l3pvUys
NbubrMLNkNzOOHFAG/b9XQKv5bkRjKpSp7HXVE1UFcP4L7/vXgEoIHaG5XCq3nRARvLb4A0+Uvz6
++INOdW0laLYQj61xnciMd1UuMnZonyuL/Xq8mTJUI7xRUU9y/8rWS6xWTxCBPWv1cDlIFz52gvo
1j9U1m4ZpeDra1uN0id47intPpbycGJOlPYh28ZcQlmi5p5oW6TzBLII3MklZL59jOp+M0lOX3JJ
l0rDC7sZ8OrLFLBKnF8sFpuFmp9FC6uZvuilQwJ+Tbqu/7eBQjB3q6OK4h6a2Po6KTwYzTQbzU/Q
QgUSRICd6BaQ3I4dShG7nwrnoBZCXNzEEl7Im/vQe/88YnlqMTKszA8C47RpZgmQuVyY37bSQpb5
e1aa9x3tBYCIsSrWom36fJixBciC/Masp74t/wlYIIUoMqukRI12jFIocwHAyzwCVmhkCw7XPFfR
4vhXW1gYCmCLlb9LrWVapHWeb+6PYruBSsUlh2VQAeEcqe8coX8GCRrpYKq8eIiS/beHIfhpCKd7
bk3lHtaN3A/KxkM1rXGEMc/sDYIjYE0HQS+J1IyAS9mZK4rjyMoEaYWwITT8ox1bYhnhGkgnPH8R
0HncgClLFipom4XfIz0bFHUk8MBwJayvQtuKahOlvJmDfsMtoQ4ELMbYo2kSb8q+jBpXcIlgO3m8
xg9ffaczWwEP+BLFE/zy0JL6Ke5kPdHcSqfsTD10hLnfRjRvNpYMt9R5TOIAw4tbP90SfmAaB/Pq
0wDVhzzD7LgupriHLJc9mf7R/xYgk55h9cZxcYA7kMmlrxNFRsjvSjIv8lknPPaDSeUaRJUfocl7
oB2r36Zlz4MuDshJX4uhOJ+S7lYANXAGsoWGd+f/04hOFBy/80hpnv2zBhso8ldPOg5znNUrfWvO
I3WopG7dDBtVypMlaYQuehxwwej6euOhOagv6er2yynmjQfh4CCWgcGI+h1WYWY4OAnfxAer6Ryh
ILD1kPfcxEft58FtpH7bAUCecI5Ts8KofKlADsJq2bgSbUtIJ8Wof2edNrmWL5xaNq31+o7Qk8Hh
E3jy2VEJimsn/s5m5RjJwE5OxqXuZ0aFYmt108VDdtFzoNVKjd+Dv0CtmirrUGh2P2fWRvZVo989
4/DTKhurKxIkVrEGhxqUZ/iZbpIyjkZiTQYztFscdcmmmmV5eNa2sbTF153QesBdxTqL2cg+r3eo
h9kXrAo4UNfiBSxy0BRk7oZEsloB97usTDQbLHzDU3g2uVqxeE0I+QtELJlyaMw0jbBARYWajCXZ
NLQa7f6pqmyRVwgBeJ3V0kCX0hvQQSLlTzW29Jb64t5mxKjY8I23QuvjfgewiRfUUhpakvy0Szbd
8CV8br74kJ8PTx1TBTnTG9SF3QeoRZ3I6nc68BOcU2AywE7kE41koRbOGFo5p2Tcr2Sxg88oVqdT
78RmDtCzvpBMVHxpaAxyQvYr+v64JoMRSVSwh8YBAnAMLTysoK5ReI+xY6RMic2z/kAOQ8jl1d+n
yGCMEPcnb6V1iuMJ/cmuS7wf5HWWHeICuzfd77iLJD0qqYK/0tQN2rOUMzLDITE+twv5nTCHs9HW
8m6DI8x1gWzzfZoA5NPVmjbQC+GcVJA2qdGfEqyLc5+quwBLO9ZJGk0LasvDIjbZVcGu/NP+2lkN
yAkawNmPTbpU+mYLQ5cPSL0XYjAyBM7M71ntBoRpkjuGjENxRkHdJ5DsgbULwwxUbxalNufke9rl
OUF3x3RfMPgPwg0DeOGg+elKAt7WmfFmZcv4H5Ut83B7fpPvF9JyNLrznAMI3w/qhHBHggk2XHxC
kGzSvxQJTkzhWXx5eNls3HRXkoZXAAbGViROVj8qPBGM6CoIMPJ331AO0lZeUfN4sRmttkB/DgBO
eizv8gnDUc2ILqqDsOOBhuL9UiRXZVrS/Enf1KufwQAjXQggmNo0AJCSJezRK8sTBUhNd1rhvA/W
RYIAqTQRYGoMW2P9yTSkf7US1K6OlGGjqHy7jpV7Xu1tv8uUuqUf/OWb5cEYnSD6QrawRu5psem9
j822EXdPsD3Lej4s4YX476ZwBUQC+KI1LYvv943sa3uZRxoY18ufHABprz+TKQzzGthFDYmSTjQK
UMdza3uCVm4K3hWJHlR5w5mDHvLdSqTlvGOrE67r9vWKK6hSC+fY1iuG3S9FCjN0adCJMyK5P338
a2j4+3PMcK5/BeUACA+Jr49jvFL83euP8Qmc5zWEFXwKOGFyk/WI2sw5GGo00ulDR1dxYflE/RGS
IsqLpnmrqj8e5iRsvJw42qqscq5fytP1KYf2WNX3S5B8IljrMWc/M7i8gfDvKFaIaM0RbOyT+Iw6
FqSHSmYEgYYWVy3j2v+cv6M0WQXWpHqiIW8Fy5u1756drJfvcnVslaJeQIuvV1a/BxT/5aHSN5j6
EUz8FWEb5HvgR4m5hkqpBbAZbW4DmYKKg3go7hRcU/kACSjaGaWcBkvEtIU5bkKQXG46p62nAxe6
CarhJRIFNM+r1CvyFnvlsigusoK3VO9q+TIkwxU7QGbRcPrhtfyI78SpvkwP5R6ABj89Tj+5EBjj
oWzwXi+iVpnZw9WPKZhu5jlh2j/+0Zi2PLfN5yu7fNoHzx3FtdT/BVvhFrcI0nYxqgOs+a/F+wZq
gG94I+Xg6I3exXjSEEzXvg3j7vffn2ffidR6Jmh35Jlk4X+z+shMeHZuQhHwyvyk/Bm+XqpK7Cuj
rv+Xu3yiEwJGBNnhnsWFyLrubhK856tiy2SB69dKSp6uUwaCtT703QEdFhacVND2ixUj8Lwg5MEq
EfjyoJaCrrpXPyn8WcqgDNsL2RglXOlF47pZ3DQaErpwCCKFwzKvb5xtlsq/Jo9VyC6jbECFVvg9
u+incA5XCYADjO3aZw1F/XNaMEm7Mt/xCujyavf3uzQZ8nRLK/1cxz6k9UHVtNIIOoYXcvCOanEB
7NJDnTlyW2CTX+gVSpwudOpjJw1gO6LuKZbmp8UCRAjAb4v944bnmAQmgOfkz7smnEU8wOWukS21
7nQaaQgqQrJbC1cbBMJWJKYXiYOXeS1FMq158tqCQjSUuys9kT5LYEVkb1zu4nFGxYO7qFLKCuaB
uyrzhr7rVg4b4KCwSHRSk04Q9FDZ23BmtjIjxf5Dq/dZF7I8NH30seAp3KVL22+ly7O0WpLDipcC
xosqQ7zKYbD37Q+ChuqnlWAUbFXG/gJFAY5G7jyH1L8JOzdmvolFVOBeTFyzruERwLvE0tsVu+in
7rnoa+DKCsxJAv2Sfy3BLLgP3r/0YrI8BqWQCT4YCp5pyn81AOxI/PvTcp97BOm6qUWSldx8jHoB
CN7m6zXEP8abmDcoGgI4x8C/U9Gx98CYiocX/ENyMMIiulWwAS1cJ8+KCq+pB8tOrIaZtFyUjTTU
JzWeh2ZFgL/OPHDYmoJ5zb5QiJuPyhQk4zUeQOq4CwJ08RHY8eiitbuxbV+9uMbDfePbAE7Y4ZAW
9s+UKeRhcvupZYNwQKIIJxLGlOiFBP+9C1qrJ5F/NYbJdTCsVjMu+XvULszyGjB0SPZXm/EnrNGm
XcZ3jzB9/h/qhBDPDDdXHLpPXvdvy6MvvgiqYoYxtkh/bqNZQsH6L9EIR9aBykn2+jE++PUh8EnN
Hjs0EFyJdBRd7qniJpwwqu/KCfQlcqXCRUm/w7RswBma+P3Qjpe5qlObNShUfds+aGVq8WW3JnJB
FD0Q2l/tVyZMhlqXcdvmG55mtCiUpqh4X2zAwiKv66fLCzua0Wl6IHPCGXUHCtoqOYveimWtQ1ab
WHnvlg0tRch0CewPL3QtHR8BEiZfq8KqHO+QFXl6KbYz/01Fjwn++4nqi1P6lmncWDClO346nfrI
/dgA7EnmLnG1lj8k5cMiK3VoYAh36eXqDUL9gpQPGyfo7xHhQqLtwY54bvSjS9IQZZ9Y0f4pY471
44rHVMBPCXGVE7Uq8oL5/wVPFmnZihpWCNDiy+41RFw/6r8C+Svl1PB1gZ728Rc+HeIxKYKrtryE
7H7XAvvAcezz1hU7iFkfK+aYiTg32djyj7X5rwdKtp/xa2tII9sf/yEY1GFtk+CZvgv0DhnyhmP5
GbgPL1tT5ZJPae6JBdyLS7myU+ogU5W1Ie9uINgFqgf4vdZ7IlGzkq6j6Gd+4FaLEsz5BCJ8bSqv
GMdRE+BSul/D5W7ugeYp9jP3/Tv/UL+qhyCYfuPd4vt6plK/9IVQyimht2ulbJwgxXbRRjb61Zev
qMyPMMhGc3s/+BvNuSmtDTGM47QOrnnAB8yNYdbzxXPKtax37jPNOUQz36cJ1wAyx7N5VFfmKGZ6
9oBeINkqVkPT+hD3l6+wzGG1S50Q4abkcFbDpaXpc9DBDA+wWByuRd1/AG8FnndIj7LaHwGHhZ9S
u24UT18Znu/giC/PZLq5TsH6DbtHqnSRIP/8WlLnUApDqI//jE+SPK5maBClL/0Te9KJ67wPxXNC
xuRrrC35HHhJ26aE2UUE94eCRqvHp8UGPW+EGSR+UZBQO61pGl0Gcl0XuDpnN9ErStf4YeWZN+cL
EK3Xbp4TTOyIUuT38VvqLA1f6o0/NGjDr5nY+PitoudutqoXPYM0oO3fEk8fu6SxjGZK4BI7s4Sz
OXc9tYklZHHkGlDHIW9UXjPQNtffSOydax8JJZKeh4N/9J/cJnrUeBi1kjdM1HdFRyhmHOjdsm5z
jTKM8f5rHfdG2wDsuJmczWYlolyqpHGFeHm2b2t93cFzoXkfBm3QhWnzd9Ev4B7s5dV6pzahQvlU
D+L1CyYbaEUlK077AStNp2pUNl3Lkd/XIgzDXQ+zy27gSV17W7fn86xPmiYUSA3Kcy5/bSEsGnJb
zCrnDJEGvqifMKYGtbTmIbE8Qfnb6sXQ48XvRNVT8xba8oIHhstimHLfQS0SlKMJ23jyMfYQtFSu
MWMwkIvxAikdeIDgwFdmMeGbIAKA2CLhOnzwiJ7p0goRVjTybsoL7j0WXF+PDDIV+SThnHLnVQiu
0OfvTBFSSWu8WxezyjaCGdK+TSkke3J3kaDCrsIXHTyVi8YBmvHV3ym49arc66qYXZZCGKRUjiky
qOyNyAq4R3/CZG17rAnOjQ+PxKEsh2aGdmEkUsIHHpUNmofsI9deUQi9FlytNxkVTPtEJTf1GSx7
BIw9c1ciw2or3ALxL5OhLJ9wxgTeL680PT7rJkBciTyBHO7ZxaA6eKmVT4TQM+f8rtK6eJrqUFwC
e2AFE22qinDN3KFEITkMw6fbq1ojgWDFd8CgSqZgr6+6kZOs0/rd7kS/HnRxikJmx0wd3of2QSgC
E2voqy6XLEmND0iBUfnmKIgVn31V803eCs0Oc5JtQ58Mn8weSt4xHCdBRfKWaOCp3jvzneA8Tt9y
O8ml6qgcYhGf9uTJxcDpbMQS+dCvBMsf4BkZDf1qlNCPj/rXAMwT/fA46/nBPdxTSEOoYzXI3mlL
aILAwL2dOQaDXZbRFx+OfXkKGERiYeKjBNONEEv7ks06ptQy/Gs/hxREMmeThMqGf8Vx7h9TsM82
/f4/VVkbsQ2w/dCHj79+PuLD2HvnuTQV1Pbm4mmV3bY0ZySnqNEph/UbJTNv5sHQnMwgpoj50rpI
VWYIc+EybCIsXdY5ajDkXQ1b0SoZnc7pVd7AwCabUCB5TS3Mw0dLRznpue80HcfUfU2ZkIpUAeId
oDWprd1i+AH0p5r8L+RB3ROdJMhIPYNpR0bD1Q6/le2UwR+Q4VrRb9kAiCZYQyNfSv0vvkyYnPkx
vXcb4YufuBwAyIFGsk8w1JxRyMi8QBD2mTpe0wtBQ6Wm8OcycmGSwZIqsKXR5RYEhkv6H0Jf+7jH
/cqiLD8cwKWnil3t6yLnDII1Db9wViJVtxzJhOEp4/mMsFthZQw3O58TFfbAqum9xNoY1A6yhKv6
JRz5QYMY43B0tLKK+dwWAyed3m2LiPGgtBlCj4NqaenjmfT61dxJgI1ZfC8MMmErNTrBE7CMtGLC
VfmF4L19b/XmU933YPxeGUsQjnV2pBADtevYnKDfw3p2pIPWgnsu2F+dhfDgH89mvhUP4Mk3mZKg
ebyFOzXNl07o2yV8tH1E2T46RCiVykBJoEB1xNZq1foHQWCbAbO0imNJwJZaiIg6tdnwBx7Vv1kO
EyISWT93DMNJeyWLDfSyQKOsNKN3maR6CZ1eTiKg9Vrd1ZDpNTj935oE1Z4fF7IwocWytHO+YMLx
xBOE7YCB996L2bFKyAkcKkAIk5o6hjb/KGYUsJroCkwVytDubz+IatI2/QS5tKE1uQBmNvs7gNhB
qircIpaHXD3oRZKtxNXULRPoTskFDT4MTjwNOO2AZUOe+Q6tCditWMvg3j2YVD3AQMv5H8HPw8KP
ENwHGjAmmLK5gobzARR39Iz68jD2h1MyPjLRYjxnQAjuhLEuuGcGB9Qx/PCYcJHsmUkxeltZjsOs
Br9R9LTyhlX570qoBX17Vmy67fXGl17uQ9D6eorJ2e9NamWiNjsXMn6Dv9Gof3d6f0C9mCe23rdz
SmqyzPbvQPc8lnavKRq8KvQLXC/m+3tOwvdScuMXd0iEX76xxKJK1undCpqSu1WgXWakgbyUjLRg
5aLMeKWYkW17c+bNcN5TaBGhO9OO+UgxqkBSnELgAHm83XYY+Uc+y33RvyEOUumMYCzy5lKl8AT2
WJ3GuE7mPBTzT8IYPrU/AWA9kbewmTeNX3XLRyJ0BRkP7kcUXrvLp21Hit4NnzukOoLmGv+GOxzy
dyOdsZ1xX1NvmSiuEoaru2JIkCUgVC+XHM1xN6w5WfsTOdpO3qeDIQxTHJw+7OC0m6YKxduuvseh
h2X+Qnp7iy+s5KNMCAjlgGaXXY1RZcDRMUePdwnJyHcB+b0YSbEhP9eV6xxbQsY8yAgj/mAUEgHk
kE6u9owCtfu2+uUixIncnggmMULhgDznizbnZA0cSKmUpch9aXnzGBofkwDl3pP+Hmlp0gzvA8PA
vUaC+EAtIjg+CApWPzpQZFFb6lpwABsoK73KddvzgKdHwd0wFPcesZruHqKc3t/Vgk8C6/oIWAj7
x3HI8gReH9+9dtDS7XnfRLOBz/JDLfuQ3X6mHorgc8NkAYrJW76JcAi+Fxdo/TRXsfWabGRwIwFS
1T2XTXW6KvGxsqa1CqDqjp9du6QEv62bvq8crYn5DTpF11bHdnRKQCs7n0CaoyIV/VyT9wpwsGmY
eGyB1LqXYznilFmpTRTV+rqWWfC19kFAVGvIxBRCk+buWo17R9GVj+igBpmN4Y2U5oK8IKlhwuL3
WPJA3NA7xU5DWe+uCPrkME1WJSBsXd26UfwMzFgf6YZLnhSiwww3uGW7l2r7tE0QixXYphwO4Cmo
RlMPtqiWuwiuN7/2PqysHvKnSrQIt8/GrgNj6miAueDeBGJ2SbnneTuvZscNv5ulJRjK60ZCtM1w
shKtfOuPBcL69T93x2FmamGCIElop3Jv6Wq06D4RlZJyXjKd5Y8URbnGzVh5J+d8hrHxjVYl7H30
gxGGymD2WOCnbs2C2/xipCJySEQDZNTlKkHHXfPNoNA354KCm7wrhzf88fYxWHG3ldoHKTWVZb72
YN6inPxGDsrsSmPNuFai9OMcuNcisxyFGZUGdc83UWPlKgw3J1OLX0iGhs76gE+R1y1TlfCUU/c0
K5gZk/oG8QItnXPrA4M97LpAgg3VpoyERW0gsq2OvSNYIWahc9aD9tkvYfNBUEwgRDZVsFYFtW1J
qy1+U0yAkwTQECFUitT9RE7fTpikGBBW+55vNRJhHGF3UhGNPvD7NiXxVTuklMdlr2+YDEL2NEyL
yAyF/9O7QkOA61wHi3a6cjxvuSzHwrmGW752SOn8JgCKYsiRoZH1Rr4zumaYXF6NDxo7FOedpElJ
WwwfdkKaAk4fFtw95pVMe1prU4TZjX+tt9A6uNZrCscRbQhD2HXfSjcYcnKFaSa5pUhdE4x8+oZZ
6MDCieL9TLxAVSRL5Y7P64zELz2HEPOD2ZnxTwPPcxIG/T16vNFckQwlqTTifYGbTKH5CCiarkwr
S+cNUnHSjiKaw5UJ9xHix4RXUdT2xkICq7N/Ad8EbiwxmvQ75UaRNOmOWHIBe4aEAUyIyRsZ1GqA
7mZbyYBubOw5+R9DfqJUZsw3WVQdHRqCNMo7fJKB/EQFuHNlfTEe55Ea+8UDI06jHpHRnrj60UYp
BEyDAF85ERZqRVTlann4BCslMNrpQZNMJf+nGzUw7wpjPhkc6AfG3p8oSI3Yr6qjRk+Y0bDzGiOu
pYqYoejgx74EYh0ny14FFMiIpTlzqCGFTRatkxjYoHVMScRH9NXbk9EdaD8O2K2nsaD+oHitETi4
OUiNnAPlSTvLjJcvBkOf0dCIDs36lGX4MZmUOQR9eomfpvyfWnQrdjZrWlpxX7kGBx+PsWVdZ+Fe
OsozHKNR8s4m1dTVW0jTQTBrGQ6Rj8y8d6GFCKf8EsOP4Q1vpf+wqITURSGsryTceo7nzOvL7pXj
VGtBKgQP3sxVtuzbrsuLTa9rlNS+E5KzzatnBldnzeU/RcvRBWbVYGg9drBYb9QCzgZQoc5Dc2ms
ICJaS8AN5hUlB+CanQQEAvU7ZATsKjxaOGAorUl6AFKzimKZ1CEIvG4SIdtdoM5lauiNzmv0f9tj
whfOaR55E+k6cxQDAOiCELDw5BeCRp5f/l05ubcfQiJRPsYgwuSYkq4hTTOxzvUKAYJdlNWY/gua
swxymDuV/Mz9EDY5MMCLzWIpBG32anlXE6myESVO9f/OIckYJIEYL6e0BwVkcZllnx8eiDZ54vMX
8rwj9waoMkXE6mcYSCzlc3tS1hPl6ive6UXvqScZTerCJv/29/D6K6smeyGzl2ZtvqNvJUCfaCL1
5TQvAvUmfaaktQLY3Rf0m3Rz8KrXX5jRFUJ704QsLU51o94iAsaiwZ01JcqUjiQT1+Afr4ADH43L
q5c2mP6VkXTxjz8SeAQj/vu2aRp+Qdoca2XIXBxGDZVXIPNnGRsw2z9nb/mEou7hl9xd+sperSBO
/vxw9Xod0YtmU4lItIigqKWRaEUekCkwYNZ5fGXXSrVN0+eGvgbdwj7h0iD0J13o18bFIYsPfmY9
eFhz2kA6MLeyMLJreEC82fxSopsKhEt0Wp1orMI7f87jRVNIeSyaLQwpRPvM25LEYeczH0pn9QeR
E7BgElOEfP1vEZ8h0ubdNX0VCPF4HvyRshLM93j85tG5I0TDkx3GsXzpqV+fISBVC6IHj5yI5htl
qup9vbFDRoLFfXItcDhPgDILitJcGEKk7xPXyg7I97MFZX2vr6baEHiFOE0RGeGidQX6szUJVDpM
/qN1qXNTwUb4My9MudFvAMwy5C9mXDjhrWrvhNeHtztUDMYoDq+BdQj4ek4XE6WP25qLCZvHNVNb
MMeOyRzt6XEC8ZrW5DaNNtjtYqibT8aEZ+3j9aYmGWWfTmVnJPwJ6pRS5uEI2X0zUlfPBxgJ4KvP
kEWWanpQ15gq38Uk7xFoof4BPg8XlEDTt6EwA5RHTO/vT44oCkvm7pd2fHAvonQEu0DS93ix3ngS
W7VRwXXDlZnVQSjx9nA7NWkk0xvvrP3Fj1KSae1nAxKDd29mw8iokMz/jKf7opwpDWtw2VYmHikr
h3FIfDz4pxzT76tl5EqqaOmXwf6fUFYxXpSKY9D6tk9LtrmSR8KnKy9GsruA4oZENzRBWxEIiQ+O
OgqQp0dnscWE4Nqnj2RbCMLa/Di6OAz1lxWbHEoZbfOnptaO8cVFZu/kC5R0K51/gdMxcYQTTcvA
IthDQPfCutIeAOL2ElJU+TEPsx2Ok0qogSwJpFtsYQWbCA7IQMm0fP/j9PsBHSRth/+YkTvk1Ms6
7HZtbUM7nfo3yHTBXnbzBV6+wx/Wz+eKdj50ikD9WXdGYJzlYHCClns/3Pahgk6f8SK1pArspz9k
ZxbHJka/l5Z6+8zlHvaeV+i4JEAgCo6zEylK5nA8Hv3eULeJX7/Jf5o3W/L/6WO1sQ7pkMG3bZN+
1YxWT9ELG6VikQPldL2TRYx1TLhxPAVhV1z1Iq/BUduDDFhCi6o2o8HvgNqCBG+kZCUhPPBfQeWe
GTmdhMbiCEfeKnc1bBZZdZgp+DW/ICxX+ML27D2oCCHfl1cHudeNuI47RgXdKL29dbnXX8CjhjIH
u383ufsBnAv4m4bZms0NK9l/f4Di8JFdRc0o/z7ee6xusvMGlGQ4P/zxixHNCs571SBMvYMiBhgR
p/tY3VUfjIpD99yhsYBXtZbALkvB4Rr7PsmES+3xl0tFLu8kAe7TPmkqKDhbDGQXxRmupO/+WWxj
Dm7GA7bi9HqrFCACNDH1hvX3VTDaCLP4orPWbZRrJcpq+F2nsYdMfuZFq0/lg6P9iOd76k2COxlg
dHdATqml7n24jYBiZwPCohkQtkaVpDkgN59MmjKe/uGprA/ZmCAuRMzkTWdF8vOw1SkxCnEkuwwm
6sRtcOs4oX/Y0VLdOjThsIoYXLCMciE80uyU7HiL9XMIEbNi+mGjwlEUe75DhRUvXiQZ4DwtewKO
zCfBEDPm5ODAN9qz/8MZKr691qhUrVU2aLPtvC894LQphQcAVrNSQPNHGrhjDZM48IiWoRMiQGu4
IRnQ6nNZipOcKgoRDoAaYz4FKcFd6uBnCwqxClt2nRyEqRgjHYyKV3AwMXchWoAq4XhoETAjf59X
44LhWssaCX4SahVlt6U1AOXYXlP5uEwzEJ71UPDkRcXR1OU06wnIqO6ui1TGXN5S8huHPv/pHMFA
tKMpOefuQBTIEVr/xGY103qjg7HB+1zBF3l5umbRSw1gvU6YOOprFk3bbr4nWoynfV83kW7KFIsl
0EcD9UnWX7KF3/QTq6iEsJCDyEpDYg23qxFpZMIHyliO/U2sLBmzJr0MxD4x4ZdFWVTcCqsFZ76z
BttyN0Rwir0T1N6IjEbzZIDdPdAvGqaK3Vo0p/5w+6sczX4X4OpPsNNq4jqfYtWma1fYrVoost1O
YL0xyH/4kbwusIa3eBDAB6onoqqROOG+GI0dDvLsaEhiPhPNRutiNYzP451S+tOaIHpTqWhaUMuW
BRC9ZMjNh2U/QacP1ZoF39BAFEWQ26iLkG7FEss/l03gcI6JcYjNrQFjm6NPKSJRNTS4BORcKMrK
aGA4bZrXxPde9nNqcd6VMdkV77O8fmv9zZEk4VfHBI6KK7drWP1kiy+nUtcC+BXGxGCj+2cYvJyx
eNrE+5u5lN39NR5rObswKeWxk9bR+erVD5Emy36Fp34oVbS/IMbd2FQhkx0BwXFh7NM0szmEKmb/
zXTyYAJe7VvIW9yPltDNHdHua66GpaTVa9EbTC7aH67L5FVlCLr6Da32UH7l4i4l9KBQjtip0S7b
bRqYT3IUkYQYwMtJ//plFSWifxNDJyo5ysqWq4k7KN9JzlTk9Ur2fZUWKD472T3wZyOxURHRc6c1
TSZ+OG6tRixqCyAGKMEsqWxIVo0Lagug4SIFeuuJ0oyD/eg2gxxr/EUa2huVaQ4N8X8/YTASis8e
0aCNZg0sLRlf1PfaZXMxP14h6n+WgR6LMXqe/ZCnuEc5iAz9r0K2OCsTexmKKFijpS8mw3KWHLpg
gql/yfCOrLS/Stp2KCxs7T8z4jffNHYb8x90LWKo7GDqIfde0LbPPP9MfPEnuVdTraFdJKZpmj5J
ljB9BXwWqfibw1T4TnfELB+IKFBM1w0IS5VcCekTCS+bUzV7rxkHeJvVeuiCuO8C1+GUzE6JtSge
vuzEbPTNRYhQy8MImMbd1/GPAD2DnXKkRNk4naSMPPcQnZBgJgZjepwCrujPnrKo/GQiSNPTP3ug
KzYIT3vcbF3opSsHt6jaeiV2BljSpwEr+ivZRid6OJeSTFzN7dnGKiRzSGe+Zqsq3xKxCCxnQYtV
zSm1N8fSmNsUVS4hewxYUrMSe8nmCQ37ecrDSytQ9lFjVSiV2cuGpijxr7y8Z3sq6uvPaOCSjgY6
O8qBhUC8jQKA6EKZ4kUtRPljMBAT7OMdak4kzP8zNx3yC0LwIXTErEe0hDKXdTv9hFpmVYyRnhFl
azt3cqIFgX8LRZ/+4uxXVfzcxiGU8mwjUeh/BuOOghBE5YiAIjw/WWj7KmspfY06v4j2zeXTM9x+
UOJ1Z6jkhQntTtXy9XIPLh2ruQMAkoO4G56+orvq52mSMZlxnQmZ1fUvSTKzus/WHdTOD8oANlVB
/cyUs5xtERuUHWMele2lWweHSZuDJyIQo1HK50s2pcxvHSwb3ElowbtQnXIYG+6U2YThPhLGRsWI
hBCa16bKa8e8wBruGbPGv5Tb9cgcqQxv05iB3lpp7yPfX+LyYW1Ud81dT9zW1Q3kwePmiTUVTIbO
MUmNNAGrHcjpyMy1ROouWWPqWoQRRStX5rb1DxPEh0zyuu1FYW1LM/5yBm6r+Y5zNpyUsuFF62Bc
bKD3gizFKQeHUApZh9AGdlT3SvksMGwA6bVu5ChnoUYWbSzJRbFPbmBYu6nn9Uy4uXRdq2SkvUEC
7L5ulsmZ8tHYo+1Yk5nvZNUqAD00NQOnS1LSnVO7aqXp0PSeGdRERUrBY/sR6eJykV1kApYaKSLZ
8cmvY9msR4AzeOWel2mUqceEFRC/QyuA+1yEdnsoqOoHsxRwYzKibxP3lj+5aIKhXuvSc9NP9TXN
XqHz52vY3f/SSeMVXDQc5NJxzy+VUxMAnrZtruFRvG2TFlfZe9K9tb/H5526mnvUxiOKEk+uvYI9
4ggEHvdPCoFSD7dic3kwI54KAoH7IK9mN8xoqAbIquQpKeRsW0Qg8NSiOWmKDMsjsdurR3vaP3uL
O5cLbm6yGnF6LFOvboofbq4A00115EZDx68RtCTuGCjhWFPf3uxYB3702gykZ6SaESGb7MI7g2lK
NMnXbkFQbYOSEDG+cb7ywNaar600O4adPI7aRMwCIrOGzIrkbvPu8ZRRC8sSU7+7Dj+5tgHGRa7K
kuPgD/1uP05QZIUzdMP2WxK8QQEMyTaitP6hYFDLFh0e3KeOgK49kK3ZE4qJrGgx0kZXl53EmhyL
XKm8ff0lwNfIj+gL2kzSai9G4IDs4ohDpXGwzv9wpn+73Fm9JaRztp4qjWu++8h0XNFmQZgWn7eI
9qik6LHAtRd5NDyr0yqdnV2BY80f/+dGGgWJne6YPB/GeP+/tTPLOXgMwm83zfhWamW2eJd0C78J
gzojO4g7qC92UUMBvctTPnmQ8a+phjBPys0DSXVM93OfzRVGhEAbVDZbe3QiXpALlDXGPd/JNKNT
QX+jSKQIOyQ0hVKVpB138UuylhfV79SyQyDuG5kXFlTP4lzvdfY+e9FpSSxXk8Q+9QpNMn1MebX/
vJsN/1mX1MXp8lOuNWovrjeZMU3XsCN+Ei1or/kDNhbdfubJ1JymVq9EhllLXDdpbYQO9FwawtXi
aRoRY64bZ4zLdlLxHCvvfgWtrwCX9kIT6czgAnLZy4+16HGesnKd81RvSxs154EgSiAoT3B7ecON
GMhXUfEETARX1Qcolvae/VDeYXhkbYpzz7Ckx9K+A6b1EV7uDnjwmL+r0h5p17P1XR3ktoshzXBD
d0UeOGVRnQ+quLCKm29s78IY4gF/Rc2zdrOiil0LnPSu1XSUwwm2Jp97GJDL9DOtb4wBtQxFaaUT
Q3nLLYXJKSuUf5lzm9CdFHchUaVViKNBxU66z1dFlZKrMOY2fVJ+gllcXIsp6254pPX9bH9NkVNy
t6yXMnFDO2+pkSDZnL5TrenOO72KV1X4r5hl3FYybZHA0IcA86Zp+qDLY2ow3e38LdVCEhZ0/0TP
3KzelPwAbZyoPlO61EIXxyaqoaRJjfbxHMpNBiUp4ikxWphnxJd8lUcl8ugGbBDpiVsxXkiFgu/7
f9QF+qermbqFlahlgofhGY57XHEJFcPTKJufkZjhvEmRhanjUDS2sQwFIo8S7BODCN8ooJvV8j/v
1+QckkuaZRvCrOv5oFa2tMmeFaruvBro2thYqwpIVgSEPADbqlLMJa76xBfc6t3ooH3Wr9EHMYFJ
8MC7CShXLIgRtdp6qUnsGtRI7HSdY9zwToZaz+/zZruieWsIF5MW9OavNuZJn0ka69NIlUvZJsFg
GLr2mgbmSZnBpwVYNAB1NlLkJtW05XB8FveuO8WQl87oWo0b2a0WSk3agdCZ6KDJXs4YUr4/tSvP
4yJy3UWMZ/UL26/MDDkf3k4MfZ0LU88aqGx/XQqv1E9Cqp6UgzOpDDjb+cCUNtApJ0NoZaJqLDOt
HNlfTvu7tZxovJFSHkp/I2Bi6uAmSb2i/p80267Jn7oCo8HIdmGGgHJq3DC0k+aV2/3LjZ8DklpA
kswM1C7fAPoSpobkXqEzOpsnPTZMJ5lAmOmuIH1VM0u9XocSizCJCaGFes92Q6TR2+CrprjKNunI
tRX7GTwWg4cV7rlBHNIAYR734xMCdan940fj+6A268WXS/OZKuRBy8n7Cbl7gNohFyVyEWnCRDo5
rOQwu+zflIeSuc4WI121/iQCgAyPUC4Llico2MIglSvvgJDuLlYvQmKr7yLS8W7cGEs2m7DVn9ud
aevNBZA5AsZq7fa1J37dZo5FC1jMPjpr+b+j9R45cZEfAOz3hh+BwigY2r58PZ7t5LPm9XxurjpX
etD7gN+cgYa8DwhgNjUFcOCiRCB6jRnGF1l1hnsBf95LLfUV/KecvpSSwKOlU3K1rv6mAJ2j6uWv
GpvUg5POp3tJMrM8V1fwZAMn/8ZQHTQfUjgDFWp4VsL5SGlL3DgK4M/d/xLNbl4ICmP/H8Pe7DH8
Vr7QKC3aogwUrCp4FAMM+HM8t2QlLMj73bFpIR+xUG6Hkjj7joGDc83oWcsVjLqMfU/Xq9UH658D
NuCfcxm/mE8cpqQppHp3tPu2D3hlcd8Yp09HlIIjAspM5J13C2p/QGy9uKW4+aHLSaYjL2W81ahw
1ilKSJRWpsFb/66vD5MjHapeyQL4f5KOGYPuudKN4mGXYFapeT6GO1IDzFcF+K+zv+kshaGuuu/c
AGjJtfnHUh4CV6AhY9iy5WrBrBL7fs7uUq+dCrb9ZugDv84g2loLv8yV6vnq+Ln3za6Hs3yKdGcX
bMV4e0k+pL9frmuEKRngwnM5Iyaui+BS/7c5smVSE18RkQzE+ueqYIwDrnKO1gUho67JjQWrFDeL
rjIAofMlzHvS3MND/5si3KkZq4E8rZSkjMefHkzmgUxlKyplSB/JIWFcEo7VVD0U1ud1V+bdRiT0
gWuNbfHme7WbIrWwLGhJ+5K5x6dfJmGhbhzVoe1VqhHNzKZho3YlJUTRwj0k66/NrULOaRkvHn+L
rdhqZsAHielRQCUgmcQX6bbNYHunOvICz3gkEEwmYJy45+BhUmeEj8oRaA8/zo4HFHUQZUzKqfoe
ca88cV78zceptLac9punRFH4RblU1o0Zoby5MuKBaQ6sZ5rVMIKox66p5pmDdxHNmijacLjWSFhx
oG+lpltXC3pf+nTkit/VBE0g8rFyjsO2kj+G5E7Ee3T8Ptkqxw0Q9i/hr7Sv8Vq38RjJYJtKK5ZF
+ExUjn7d7Qpqa47tcq5MbNiKPWJlBMRyHXtEi0m0tuXtmiIlzPN2ETFQN42QBDCFoiEozi/dL7vC
iHD+nq3FdxVRf0BtbxEkns0orIqyGtEa6QVqEzrtOREutLn/i7uafIYMc0uPTcAwfIH/a+vHqw2G
t1337tAcne4KcasN6541WBD9LdeREOiz7IVYfFxRcWlSGCwDcrPWhWCGSs/tfr+0wv8fDLU28WrQ
8GB+yQw7lSv/Z7fpcPUapDqPepjNwQtHnmu5QnjCum4x0A84XhlBCeax6U4Xq8oZc626dfM25uF3
GxgPRAaYIhZBSkNipzOy9Ql6mteZuR2wmtekFKIh7bAsB4hML3Qidb49a6hsCdqfQgOXGryZeZaM
hLcuaCoNSTmjCLdSU4i1EfGVBVFCBdqKyqXdhys0WWgtB3gTOVlO07iJEaoojIfhaAx22foafqc0
7rfn5rdsP/zIb+Ze3frjAlEQ5tAPcTABul6jXgWS7vwR2CqO4nBSaZiqpKrOT6XUEa027rLHHRna
vv69GfY0BF1paNXpANJcUaezeG1tYoGOQbgUCPn8HJ3FxHCqj4oFbx7uSn4MfYS7gkC65lmcFVyO
sVmUa0bpaPmrkGAzKsmmqwk9CP1IHR1CdSQUO9HGumq8b9DcDqMUb7gEJHO8HuJbDLys0FG2HG7J
f9mVsR6AHSq6emZ2NnNCSGb8TX0PRk3vDgAwo1Vz6qTW4tcAV3za7vD+78UxZ9vZrMycZ/87TKSf
HnMo8oBkDRoUCP/UaCrUff95uzDW657xiW+uCmZ3dcvsVVIS5i9Uh6WutUiU91IpMOsGlP3sIeTa
jIIaFuwHZBoCwiFbJqjcEQxDmZjAiA2J1t4WwhZKmLNEZTWzquQaS97z9taMqdqVZRX34osztZ5d
9VKL9oYYvbctx/9y/6tr/Cbvwy1JZ4irgz7O+n/zPLNO4pfwq4klTXMcxS9QWYotGv3pk9XZKA2V
+8ZqIqpewPsCLUnQe9ffJiXujcVYHMlJQuLJOLO0o3HR+sTVkwIwBLi8Pc7z982lCIt9uL7Pp+SG
7oqXCtJ7dMykA7xbqJK3AZ2W165lD/pCguKdFa+scJCb0n1x9q2MaVu7NCepgNSXiJrGllDNxeyu
vdfXDOkUOVUmDbk3SUuoaxpdNe7YfB/THifq4PGcFSQC2spX3I/RggLZwQXz9GI3XeRyfYCeENHV
lBI/YqqD7j5P5BPIWs3rdAvYqlj5AUzg6cZKYM84sFbG9w36TOGo7ZHDHzSmEgQm6EMYth7f0COr
lgoasKYzmBJUxQwaPq/HVImQbhJJS5O6xWV3QIdQoAUmyw2PEQrUM17v49nyBypHi6ceWTdyp3o5
qafuBLBG2kE9H+9SKKZ981TSl2oX0ARG8c+BI8n/lmQGmQhvse10TCLIzccAdSGnEgx7R02MM8j2
1P6WXqqNewQ67yjl3laoeTJNXuEFdBaWKRx0nrRqi6QL60hj3mb/jNXzZZwIB8ZVsCKVNZFQQtuS
kEe0wQIxBNBI/tgKj0uRLBYFz9NAJNjT8piqucw5s35DG4xLOlXQNpTMSmvQtwKluvaf1H6TndrT
oEe4xJOruUXGOlkI+OzqYpbVmXn1bc8zWFbHAbY25T5xB7lLoe3WMJTwGsp9gnVK5Qaou+qJlyGF
hY2gcHLEnJYn+Mit7NRNZuxo5uNrwNjfuc01HX/wASNJKPSnjueq6AGFgbyYIrmq6UdUK0ta8x7W
JMPZtv321l2hhoi5iV1PLICKBnk1uEcuqbuWj530I42nKRni/+qFmqiuH9HYNMPtmPT0+ielBw3r
OzHJWWLZ5+HdsOj20DfQ2coNUM2RD1PXRtnX8LbbzHqcJCHJeyAqATWGi2W7f9oN3FwJrZ9nlnnn
ixu8t6DHSxnzHV7rm/AtHvVf2yqAkn2y/r/vYEK3mkvXb5Xob8e2yVGxZlQD/AD+uf6iKmqrWWXr
iJLFrzI8G3X7qNw4G/MF/c0bxSt1tw/tfFAUVWOInHWJsqPyNiQv6+CIc0sA9RJGJTJgFrXvfvFW
TZNsJZlRMbu2ITBOC7NkVCXMr3qDUmjQuaHPwR4kriRNu2WO0GAY7qJtEtekDvIcp4J7zdDhmsVk
cnc2myYpQ0zSIVULWzhSP1qYuY/aLXECIQOhOhZzKoQs71iq558oqKJSw9X8qZyFSeo2zyhS4K7X
qFXvKZFF79SqeQKJdkP+S0eZgsVXMjaJOmoqCtvk0Lx/c5wcIc2H/xq6rooQq9l5ZUWfO/5aFC1t
JiHOLERU8X207tgbWJNxT29xaLJVV/wTmiBrKenS9yLZpToPI3hBx6Q2EussbruP8lFe4MhAt5Fa
6yVEDxhwVnWEWvDimNhjvvQdiess37UwLOEqTCmNw8nHRCz8bMdFjaBtKfhbrlxdBEaULiFsY21o
nQAWlknZEsKaMNQHEZ9R5v2pWEM1kET++LIlKmM5yOdmNyVH604oPHm1foTGcPi16CwAbaiPkeVP
CrdKGrqY+9LiCdd5LgRCrmU21rRSCc47tLZqEdWfzh2YWUdCGJkc7A1QBIyo2quHBfMOZL1rJ4pW
eU+KplC3VDvXTQFBFEpaCcLtL5vZ1p62GI9gsFNd6EW0dHJItVWGUkT989vE2LqI9QjrGmo9bgnY
hoerN9MXrYPKFS5SNwzwJvAXphFzSImLZYVzP1nzTXJRaOml5bjHd6eN6sFFDGda0DrA/jXUTEs2
q27Vw5x1luBCXzoYt3XgeMnsgB3IgG76/J2drTu8HxqvlPlEWP1LWbxRT6SeKUI5qEzLgqvhQvCo
/UAwfrG+3okbnj7KzSw89GC/7kjVem4lidbWPrddY+de/gHE5QdmgtYKpMtgXBMuA4/rRnWy01vs
vE5XJ1aynU8NWqkGTr/vu/R/q2FDkAJV+9vzvifg+UcnqKA8B8EqpQ6yUzJXG0f06c6ZKAL227Nr
RGNIBSSO6wvnJlJWWLW7gQ3BnoPOk/8kZpif8a3vR1EjvPycVJwUusm9VN799ECv2chqhUm9TXSt
gc4KMmPnrNCBJIe0FMXAYyVmS32FZlKbwAX11oExbHaeg3LVSO9ljY+ie6rEifTpfJci6NVNweDS
kP04ec41jKflx1kXWTT53uWMFRK010ro/Q2bSOpMl50esQ12iigU2c4G8vewuTBLHFQXFBWkzpFA
h7wrpz430pZNh5HWjA1bZc1Km9VMvivNcSigcfPortbAk4u3ivcJdRK9O6ECcRS+R850YJkws6Nr
09HK8C0ZQ5iUk3iGt+/wI1hPUnZuJwt3Af83Ukgg+oNMWd+PcWIRzgRb43ohJ/gmMs/luM7yXBsi
GR/RRlXfpsVRTGmFFX0r8ZresXWsIpq2/Pax2e8nuCJ6buS6dINbj1TgXoyoPkP5i+Trv/iS9Sil
sf3pbOwJJ92UFG8hZCfwiR2s/TkxYpBb/rDFVo85b93aFPBga6tAU885F4ev1J3TIt1FX8NUP7IU
VjhXq5Sn3NKhK0SPM2s0vmcLFN6gN2e9+4UL2Xg69Ql3RigQCM0kczwfNcWTmWX9gjpheOnY6MfL
01m0nyN/RGI0tHV2uz3UgBfx+nUi1nVek99Sh7dNU560qsTiSafNgvdhMx6HCzbU9jsphTCzr2gH
YoMM1K3eQ3VgxEvGvgu0uBusqfPJ7jhskGu9EFoN1j/XoklvDlYk+uB9/XTTIueDUSk2JAl05jGj
nBX4H4O6h8AUFBRaKb5OmwxH2DkwbxOrd+m6MlCEImTWLvXgY8V+qUVqGmNlyqgOJ5bfjg7psILc
hYJ+ZMSnFv3cZOiTyG2zmv/Elssw0Ic1khF8hseyMpVmfxyzePMTvwTAolWN+7rSBCV5mj/vWmUm
eArpsZFJuEOslfLeTmQSBWuLphig0WXMWPdXZyXr/sDyOU3UaEILeaqrFZustxQ32aYEndkx/ySs
qhDXVtOijXHRqL1f09YK1feu8Ft/cZSa1WSGGfldFKGFrytYEjRw87H9RhiWRcEKxH+amsGz1lYj
AxPH5DzllAsndez4Zia16fZjTy1DdRju8wGMoV1ROiKqBvgnYknsAg6DaEg3EDQriUXsP/fAQ9Bd
H9twYnrBhCeST9elgPtKlkJgTZB4KIKrJO7N3rxgTGDPWs9pGMK/719+nUQnx1DhD2GQFwDg7LaF
vohOMePtwxTzkqpRqZWnk0aKS4UZwbd5GOpF4UzYPaunOSIU+Q/SSl1lkzMSwrHEsb6GDQ8zj1S+
4XIApc56pgR9pVVab8eIGAj9CTGhDIhggVtMDlVyzMhaG70a3+rMKXxEwhamW12roebVciNJAq5+
h+ey2r7CbWEKVCI5l0tDi3qfEFOPDof4gtg+5oMY5WS/zRIPmhwaPIblnZVXsZAjtaBawoHfGDF5
Rc4gf6yU0MsTgzcP2940xRGQVgDjaSOy/RpVNcaoNBrQ83/63SoggUGqCM8aWn4iEF4+UjB7/0lr
2LHaa3diZcL1vsTai0rbsHGNAGn/PMMRYX6w63BR+Mfm+uHE+aihBcz7gFUirOanLNzWvP9lvA9A
kq7uS8T8mhQuQUUsEAakKFbWyAB0+JGX4xImBDVCZypoY/2X5BGA9dL4t6pjg+rxC8eg7s6dVaL0
W1rLsO5F9xqzU2IhsFgHVFZNIAgaPy6djXdhgTZQxlYtvFuvDmGfODzunGco3Gcf1ngsYq7GgAKe
FThWZJHlPLZNE5ytntgiM0pjZDuytXlKDojRXDx/XK7W935amatHYqKRwDTKFvA1de6mL0QopjU0
1IJaeLbnmP/uJuKsEQ48CXNHjLMShw8DAEN8fcJdoS57OQp8vIkQ9vu0lqm9FpbvfhvS9G0L74tk
BaGJqQX4pvM0OuVYrAvVY/4ANe3GcRrYlfGwm/sMUNhoz1EvYDTg/JuHJHLfMtLhjZGIXiZ61G/M
GsxUQB29N9FMdTosxYdzk/KKCNSlwQuOYdDawK8SfiqekKhazRd89BToD/sXUfMloxXbg3d3DoqU
ki8AMau1Yv2v84LywEP3ig6/CvUYZ/58UyHv6XK29dlpUkV+shnEq3iNIqbmiS3Hgq3/gVfLScnM
UYe10x2O/m5bDLLU1pus/FoyUUu+BJ3DQ3dKh5SXECzA+6qLgLZQm3rspP4UZRDV6l2StTBhoqot
uxO7J4TtiJXEOs5ZbrzTNik8GL2jdwooA5qGkDV1SLiS6ap9xGKT96UB9hun/j7MgNW381ppoukT
XjQDJtADs9fWAExWwvpmMWD/KIuUgr3qvm36M3ouVXw4qWtJ40Kb5PlJCixvugBAAgvNF+CpeD7H
sbpCCp77pWYDxEup2WzAZhJ/HnBBWv+ILyyM8+bhYhAlKniqaUqIj+pji8bC+xCYKHPfs56v84Jj
EfdHxpTNRfEOXsxFCMKlRd9H0M6tZN6PaW4vpz8K4sTEVhRBCEQ+FaUO+wrYZUzTPUMSUpuv8MZv
suLmHJ2hqGn1+leJiFnN9trUnqUSINJ+TcGsmNn46MH5tfvbQyF1QPioJDFK4PL8q5h10BwhXbis
SpvZTUzdZrrTMtZ+AiHbrxM1RMsr4VrMh+fblhFu6pB9RxAIql8rvbT8AejEWU+kiTf66oTVuYmS
T6GhlQn367W3lXwIPZNVFUTaubxijGxluNki42UI3+2bdDDNUFnbPIepbsxTuhzCsXRm3jL1W0mU
yv+9hQLR+s3BsCmStcDWtYYEoi1V5ED40R+DaUCZcxUS+iV8iqeF82x3mGueaweyACiMOn+ZOX8j
UN9TNXIcXSvuVJtxpr5g/r6Gxz2BstnAnujdFoTFFz095/8vMugviBuZ/O1JkwqATm5phi1fukqV
bs0LBbb1l8G7Kia4cPJI+A453SfIbGPEcflU06HxllW/cfITMJdifKePJA49AP8gmgGh3UXUiq+R
aQjhDDqc7dtozw3IkGVz4k8SQdiD0AteEoxtfTIr1IGZUbh+N2QZogjRJgBU8YLbdeWqEsbRWnWP
0UCQES4drDb7tXlT+efZNh38/fZG3LOK5OOr3zIFq+upfx8tGXmULB+70aNATJjfsM7Tom92mHBY
NOrg3kFHCeIy7z+HLZPso2Xfcj2u7sLgwd21Wpdoy4/ops46fGib4aBEhxyIUwM39kHLsQq8kMdv
6YQ62ZluC4UcqDVNXzqlic7gjyrSEP8tcBmObFaV6aD7/219rH5bAuuGdBkNTlHrMzK/cu0qCcBL
KoQzt5oh+8+GL8SJmOmsd757LGGkztYScUFbrydbdOkFIa1igbYdxg1D2uJCeBlSCdM6dtVoV8WD
oQHTSiTw44ht2l1drwETUqr9ckOVxg75fMHevlMiUw620V3dXCeK7+TXqrwQbR1ZHUW8iKF8gKm0
2Bfd/yEAIhGS+cAXRrCdc3SKboZFerjxu6n62IYhjBT2z2NF2V/JR/M+O2Y+buXTTs4Fp4hCX08k
qKYN2WRtwaoW14LGYX1/CxgyysZ63BkhMdK64L6c4E6HwIVXjUSEwuvSzkZFYY8KflZOqwHcTRow
AvhfIZ4Zkc/Zj6L/wxKy1K7pi0UnA5hwEuul6im57WqIvvTLC61qy+Hx9a7SME98GY+zUfJZBE2E
7P1EMBfBFSvVhGbSLNrMlEWQ1xFAKF4jrSH5+K5A0t+cbU0DWSs2nzh6X1U1xuZP+1JPZC+In92a
dgPjG3zBBZ538J3M/TSxnXKSvM/dC8OLkpa7qW1DvGxtlUkqLyKUvCyanIYSSorwEilkrUOCtE35
52uL8KBMzlrvzZCtkqQ/9F1Qa3L94QSrp09HsOblMFdvdFA9pJHMq+fjjFVv74NPmLDJPIyfB5+I
pbTm1HUSnx7w2qmBJ7v+14ir0gutvkRNTqg7+x3a0zTL30McUHgbXAH9PPBieiozVPAn2wtmivc0
X+1zRsNgj5CUvm+M2bVBPkNerRL16+oSZEXL+vfRjeC9W3uvldPCu5CLzaHpH7YabyzmnBeg6Afi
LS1y63CLnEdHgMD4Xov5IH2cCFqe/6+FFDEAnyVX0aVDBS4A9Qwjs7K2gRVHeMTDuiyS7stdOTx5
TOvpoO5CDD7c0nZA8AfYmpN1ldHpO6KK7AfGh73l00HMzcJYZVhXFdoNHwhWHL+bztBQJSN3B07i
bJRxBU0fyM1OE2WxDmZOQtfj3r8wMmSOp3nNFhpOQf4jX9US0ablixJ5as6oiWcGSQk84QdSzoj4
EEc2GxnY3dktYqjw/dLl6foDoA7GEDOloCmvtdufNjJf0nnfCWsxXDqxt4OOmLkfXgcNO85BYBq5
djk6m5KA05CDP+4cUHBiglUyT1YJqGgzlWy6FyNCcxFt6e7yWMdR9flkVuL9jI4qr9ZPmHlqezEz
S86Qitp5LphhtIiL8sAM1Ps8eCUvUnUUjxfVKLfDudY9zGoffw9QOWhLuUNjUg9SSYkskOwmZLTJ
RztcMEz11oAhtvpB2tEjhtWDlAjfnYdSJW/S2zAz8RGlI+jWTLUdtCIrn+G2YW2LQ1Kxe4YVuTfX
zqA19DHlK8AtEvK/gaMp+lIxpMNCmN/lb9MjK1tDNeiWGlNaWTwiwZZZdyPjfTMDnsHCBwThJW9f
CU7dALMRol3O0YoFBgQrixezWe0Hwjldf37Jnj+17zbMMpL+GTq/Tz8ZyEsz2WFTaVAxsekCn7rB
gLFuo+Xh4YtnZk6etr9qHwfG/tDQ7nsgUxV7YbYMeCPQYHpnbG+C1cmxGbumq95ugoD5AIBxuPSy
/FPrsfZnCPP77muoVl8JS7y7ifnuZIXROzq7MwppBiekA0vLtUWefLaaGfTgH3u9wAciOxk5Ml4I
ojSuVH8mX0SBUrtNBMSTJhd1kYGCPOCLIWtl4IVgAjz6E93b7ao7vnXeQGR/UcLSJQDCMYrt9vV0
JY1jW24elTk4DD1gbZM7OcGUV4lbfq4G/oIZhZRk4JS7ckThoy/9pUiQjAZDejggAVtmJpnOzUuW
vE4QTWnktQCly+HaGwB1fAyMO6taBc/y9MyZ/UEdOxlCgyv7XfHzlzGS0PEB7wDDrZwLP8f74JVS
+lvh5smp9JgY3DX407lkNiKbAlNYq56vY2IAlaf6Pdf75NviN2KG2JBCJQbu/eW1EyNP4PWXEzFO
XRRJZ6eVYGKuS7mgJhBHaPxOfnWdbTc8gpzJdlhO32Ub72G3hcRVf9Ad8SRDZNsy1dxrY3emy4Z+
oMBRRxEfmj+Kzl9OpM8k/XSt6DOXn/GPGweqX5xwnqtV1fcgBpXX5CW6m4oi5DL/EPInPrNI+lk7
v1w9yo7NwrGPfY3j6GRNsI4WuEdl6CLmz0hvmCsGO12D41bbTVPmwzx70X7zEqpLJNtbv4EkUWxX
lw9PwL2QantdubYVt2vf8slPmQ2c7qax6cB9Cpa9Uq4KzeKmfp0xdgHjET2dWTi88DMEo4+8SXMi
HDLv6GD+4nDMICQ6uUuvhYqR06m9F1H8LrHt3d0/s6rTrb55QySXkBDdYq2iSmZZq+ELvm0R9ln2
P9oLfLmL/PAghUOqfbDaIWgOXfdg+3v7ZBlfjxd9StHedndQSzzopsnITR2DBuZQfOe+emAYt29g
9aHqrbqhJhCBlrFw3miS8Y/KgZuPPVOebWlowFsUNTeWUZgEw7zcBU1mdPY5h1foax79/A0+w+jQ
iyF1KjDQtXLa2xVX48CTcbXbFUfwq67Zv+pNkLZc358yWoIO0l8Y5omO6sP6Kj8Uc0QkbUoA5n0c
nZ7j3uUfR0yXhHLZwarODJHQkft12afuyULo98pCQiL51aLfJcWr4shIe1WFwjYQvY39x6nYGDxq
gp+1luwEKlC1Fe72nP1u7AVJT55Gt92Wm7kWKca2brvXv40izWcsNCB/PDMx+dUvhrk/zWc15Yl3
rBgGm+E6zGXcIy0tw8RfRqWthQxDEigLu01iGFyMQyL09T+rtBna/iQV94RBHNBSx71KgPwt0DXf
ZFzvigpyAOu+in0IM+5MTSEGbmJVDlJtZjclQtgfq6sZC7/u6oGtjRkch6CkS+5XFj4osAc6q175
c3wgAIsP2apWZCjNCoDVcipao+TzJ6lgN40d1hbj8lFe1PhJxdctSQwDFrSrrb1XYadVXdA1tsG4
E/zq0VWRtJgzvbhzPfkdRpJrQhW2Tx8lHEi5vTAxNYJrdZcsChg1iSNGWIOZ9X5Zjq9dekVW5W/A
ORejU25I8r/ihJF0wHU9rlPgNV7m/+MRhPQ9v7TUwkRVJ0S4Um5Y3ynxXmbnHDo6EecFdhzCEi39
BLEP4oUw8CoXBjRahGKtt8P9f6Xx3eMLBLSmJhLTMPyYGaY24Pvs9Gxna11tceoqnLitzP/MFdd1
ZwaSYMdlUa8MI1zCEgHYM8NLmFLw1v0VAY65E6pnslkEZWL0MSfPtyNgzTAe5Hg3No10642CXhdE
HpbtgyQuz2y1Rwx1hoHWUQFCAfFPZvqyhLnx6mkrzc4DtS7CXVGbah4mxNr6MjEffrLPfUwfL/yL
kG8A4QGjG4RWC4teeNtu+9xCm5laqJZTJQNI6U8zc73qdiPgZ9DBBMs80crwrxNuYsO0GGCf34bG
1YDJHMxIHNniKiF65A4NPNEyPrEnw9nQqQ3mHgwuKsW9kwzIpJMqV1kHi9aNsXGwY+ecOziUKNLg
DVvnj08Z18+xF9ntGQvP9iIsJgMFWFm/Yczf6K9TbYanunIuUFnr7bQE5GZNzrgRGWhE/1Z+0x/+
DvlZQB8cPot6lwSv1+WEncMZFLUispWn+h0zjjwhxt9qeF1CNUwBHzUUEGXBTrlEnBXJmt2ptvIt
5u89Ez9K+eGtS++Wlp88gqTvr8Rs9pxvDTYw94xexXFJva+SIWlCcd3v8N7Aza0yeyX9hCIy2vXC
p72LJ+u5GGqxWxIj06n8m1Ickx+XgwAAmAPTHQt9oTkd2GsIcw0+vbrN/q33RG62mCZY70fDF37f
EgjltRinXNhQ0ZVUNihJ2WAJfIh4UcuVox7Ik5ZyHsjZx7VKxK4D983rbu24txObuDSUYbY5dVPj
P0n99ck50izm4ERLXW1Yg/xD6Jr5UlyUJLpkVj9vdiFJFteGPx/l4iMelwFpVy5ThA9a9KjzfjvP
sEfszBEAlNZ0SVP0pFTEAtuK2NkuFHkHDW3IqLI7IXT5rcIH0x4hVTFO4zju2/uYbyfu2RCcf2De
fhhWo9CizlGYCXb83+6fRZYuhSFViX2v7AW3WtCG4K/eCgULiLsPz+UGaaPpezSfeRKeRDjSbex+
kRw+UqOhkiJxgJ+DlvBnJT2dW6kA7gkz13nLIVBJWSLHkRfLqCWqZFsGEYLOZjrsAEQeMgzE/hNx
PMeNe1mXM6GUB2++dFopyxnf8Lixn8UD2eOzn72igYRbq9Fr8BFNSoE8Yjhkys87k9C5VswyT48T
1m2CUsjRVFsDkUIPrmUlwGrNPiJLNedTSMN7HR6blM4vuByMokLH7bRqK1wvZnfjlLNTBAjlY2h6
gFe4lyG1914ow54gAjs+eEOrIeyR7ImezsX/Hket4UbjVG8Uw1anjQjgznGaQeOfkb6USnIMOp0+
Nm6ij7ITrng/WQ47LIDS/TLLyBHPKcCV0G/12JcLV/LQQSdmjezWy4G7DpKN38567GEkhF4uTtuo
MvqE+IdS8fSIZSLPTFiYD/+KajW2M0b3daObN3BOQF/jmy2wGvbpUxML2qMgD0SsRySjBU986CcA
90nFS1iNTDgbHdTrT+lXIVAKZR0Tdt0H781azi3AOjm+/ic1zWzaY4iR/U+byoTvDNtzrQlODelZ
u3LWfPxdRcC1fQ9n994nPTqjj19anbI1WQB5evqAWrF2XRBPyKsghOgDFthP9q0uBT4IuqpkRTAj
COnlVj0tPE7JqS8/X36xtmyQYmd8zNs+2KHdU2fFQB36WX4uxq8hvginzO/7rpMsJQoKcPPLgQ/z
NOyXLr2InMbX88U1vmtIxifRm1OCQH5UX5EHnyq+Kl1PKIAm7xJyfiXIBMCZDATvcwhqlEkKRMtj
2yTIwSU6dvupYHQNeHd3Az5vh/VKmdoNKyO/FW9uEu+IDEJNyUUfod5q/q6dJLr3nkH8oIPJInAZ
iP0m99rq//rByLqfjkwpAZgfzu5IGUKl+AHn5xT0ghpQ/vuwcZs7m5naIMTahpMDBiEXg29ShYz3
KVIDR3YBZQ80aX0jOZU4YuiFPtthUy9triJ3vfD1H0RpqG+D7Nxw20YIxVqiqMtZbzLWzpxGSE8s
8XpUrLbg/MFTEIj7J4TAL2To/jmY/8WmGBKOof3cFK90sgYOt4O4IMV7Q+V76Wl6hs0bFdNHEHFG
PhTgI/tRyuIYRdEfsin3oD2pWyieKo83spE1ue63XR1Xw9l8OGAolP+/ecCdQEl5GbBYr0VRkMWI
Yz9MD6840txgP1bocTJqrHaHgPKM98uTk2X41mJLz4sRoDbsrxbQeLPMHnPSxj4spYCyoIBRmLjm
fYBkzOrTENjYWRUIHksQzF7V5hkWVgPicrexg1JOJ++FgK/YjLtfOvYtri/jJiTElhv9HN5SeVch
Nc8ZSH2Xa2hclDdM9rNKlRufCjUK6uAwOrSE8dJfbbko3ZXsR700Cr33XD1rfOtate6KgrgoACJz
eTBG1pMHR3NUKNHXimTPOvbDByUpReaxP6WlF0y/RJPqDR7i7ADSSBs8U6fuk0+N6lkmH4S8QFII
LQZnyHal7+OapEvUkf9hBS45uAaS7Aou+yOrqcMYpjBRAH7755v98VxCDAUpdOiZkxmt1u5JS6hU
15QlKbdk3XXWPGUl1Yfdbqsush8+WlVtzvt412JGod6XdmNfprl6XtUPWN7V482AELEE5Ul0iRWc
G+dzS0Ry0HrmBqRL2lYNEkvUmqZxvCTANVZxRks6EXmN8RMrz7+q/E4XQ65fcCdRbYAnLkFGRt2X
rw7jUPNfr9V+LKlozYGo82qnrCFZekS3dnzY/FcYX7YTQgORJURlLjdXXHAN8zeQANQkClTZoWTC
EX67le/SuXWzL3a02JxAJ8pkcKGukw0jyEhmysUZIOI49bUDM6ZRsEhE9ltHFTR+0LSGkzUDMrlD
m2LLdjE1EyTkuNn5dd++AnpwcX8vviC0rUaZRdYuBvTAeM3w7fjnnYngSrS9zvjmiytW5HKHoN48
HmIoMEdwzvJxadddqk/uF2oIF54LCorRbl+DFm2deSjGEgr71+sSr54+j1T9mlT/FkSPf94Hyz6q
AbtuGZKFmR3WbVAefBLBQ5YpXBn0SFUlXFgwZisNZXNgVJZw+PXPyMexCs3YFOtQ2kWtF4QPaPGx
cqsT2fAgu5ZQWPgzR/+pRuKlGkWxZ+vKKRyo01z6AWwDwVtQ0ClYMoBS7lRum1Aa8MhWLoZYFQsy
r8hYID5YOpqJEV+iOV6IB1q+hvNd4bonC5k+yJu0gloYLv+DZgPKrnXSChJrLr4y/gO+SZ3BJcLT
KwprzOaaidTN41JOQZDy/MKxsOs4mANqD+J17nKAZhyl4JLNzLCzPsA1OYnGYSXjuGCmr6uNVg2p
Lp00TYtxtj81FwQOospifSA4G13ydxNK7Ll65jHBHW2IrUF8Hg4I+kgbBBgrzGEHxPxMdow0CkR2
xZvQyvYyxI6aQOKOPwEibMkvrYS4LD2LG1FrslnkHSrbbCNUj8N5f7pRVqEA7JWzpn0it/dtrVWi
pLarwFc137ODC9wn37264O8S/9SgnGq/r/9noJXeXwNO4SEr8+ZZp1Czu9HCqWXmNF9xgY1CutxM
eEmOsEKosEKWpdDqRfJLyLtvUTLVbIWs2HuBPyiX7K5930ewvGwE/v/7vvU6sTab/imDSP4hSSEv
PQnFz41pFheOpqDNz4QBhuUlONOt20AzNJrDL3n/BuDrVffOWmAGoFr7r7FmiX0yZHkanqK3dPy2
tayV5RwN0gVAaHO6xlN//VNEZBtew+rEctWsgkZ4UR3x7/ZpgNExfssQ9cQkDQpHhMYGcXdB9Vht
WY11m/tFIJ+z9W50DYv/4JjHueIaitBXDpx5K7geD8XbSm2Qz61se/8eT6CIN26JhOQjyZChCR5F
W+klCt88cZQJXahleMrQpt0i9oDXXOK4sS0WvQK//hqAxBtuYUHa9VBcs3AH0SCxqTlKYyf0cPwG
hkPm9YEq8liAlOJ3efix9G22x45LWGyXVBUlIY+4/bD8M9hkoTPy7Yrky8jH5PqkwZeS8mqFt+2N
DBFZgrRr1pCj8mby4xGLp3SA3gqNAaialIoqWdm740wCzdg5w9T/9sEZLW00C0Qo9mCWpMzUEnCS
dIW8Hq2pmqMo455qDguW6DwEZtsj3EJF/sZtwphlTUHzLB2KUUe1/guFGlBF7x13SXXloJ1gjGqw
D/fezNrdm6bkAqlW4c6Zx7sCqeyHA8vCNn+g5actKt9kRTF4BKH7W7DhcLpgffWgxhJsTnlto9g4
3ZpgHkcljA1hCX9EYycUtohNv+bsX4OiXl/HFNDn9NE5QnrgnwKQTSp+RGm72ZhHH8q/ljJJfe2n
5et1A7hR7POmh41d8mLmyOeF0VoKzBROWeVvHYJLj2HY/8SoUyL54YarIR7tpNeSZZAYSmCsjQou
nv8Ky6V7Rl7LljPfvepRSERDrgYB1BIsHQmFMx3KKOKzOwO6/jy5niN3121pyaNf/Tl0IDdf+mvY
lp8nyY0ESaGe1W/a+AFY9OQY7ZVBrX5kDs58997ym3oxJ5YeIBH1hH1ghvix7daiW+DVHaMnJvf0
/daFzcLuXLsx5SsDpK5O1EpWMav6UcPW5nEWVZN1co7YLY/G5Q/8U2Y8cpNvfU1sXMnbWuhVtzfM
CXUKPsHHeeO6uGwonviZM+WJKVeA3IOw1rxjTBBBfrSWcODBGRvvz1SkYDG9tH3YGr+igSXNQbpv
8+Jj+LqPnMyl6PSuAyDfkb5bpzgGvXGfGoj0POUC87mCmW+dowHxEbcxZsDQB37+l4GceihegrFa
903PtmjwmJkdMkeLOc9tZVgsPsNInFh0uucRrBQtcNQaKstIn3VqW18g7ojgmQAMLcTITouRNwzh
/5W8iI09pj0taiLTh10D5l+VNqSzQQvlSdwTr+n/wMejssA9QPUggQ4zXrnA+Iw8cVxhg0ao2yDt
4N58PJTQ+u7K2VpHocvy0jTedI5Fr88MA7fIBRz0dwHeWQzSJIE+jy0K3FWza7Pyq3g3gPG/3qxZ
BbUmdAeIOV0h0Z8evSo53+Gjo1nSd4RsH2X571h1Kp60zp8kG1uJHkXc3hmfNjKhHElw9vRJzyv/
ugyndS9GOUYik29erKRWqRsy5CxffYDPYIGPZi1h2lWSucsOXisCHskxAeFaFIL8nlVwgANKy5Lv
SVOW58VSsyFh3779Hx0LkN4KEYllnJ19uh7f8+CXZMx6rPXlwmJox8renDAkLEOPJoj8uNulC/mF
Uk/N58gQBijovHaWHcrz0j5uXKzfQ9OpTDgafxkJTCDZZjBJ2ONLCRO7usYiaAj++MzYYYG1/V7U
6YAVFjrSmbxJv8aK4wROTX6acBSZH47AiQgYW8M2ZcK62AkA0Uw6FLq5Bi8mrjPX8IZ19yXqoE/Z
5R3gDdmZkI6Jqfj8JEkFl4ZubeT2cGNRxEpi3pV/lZ08PHpmTPJ0+X+mbwC8R3W/tAQuMYRfKrts
4C0BxaIlkA+Cl7tBB8INJsg8Km3gtSf5Mp11PzD62IUjpCu0ZgjojCS5o+vuEpy/lLWJ10hsLDL7
3LzhHT56QgBh54lbyZZOMA91csBBqOyDgRZff6cXe7Nh9ebYF2SUD/KMbZ79eFsxm8Zp0RI24VID
g8I3uaF5DikUkweQBkvZXRZXVK2pcgv6rBFl3ZAVPa8UFREvoAVKLgxPD3vwaEPToxAPnUBPps8F
I/ox09+3KLlTQcXE0Bl+2/ojW2PyIxE7gSy909fZh+XKKknAKd/J4dbhl7rdsia6/Y2tMh0d0dS9
9o3Q81+QCfTZGKtu92c6HZnWVjAaZg0hERSfDOT0l/bAjEpJbXz1iLcjA8wDWeLgMf2F3R0DPClY
M7/+10Wc06RRxxxvtcBSu94mNUxh+bgwVc7+uddY6erHCZtLLZ6xkMYdI8EIiNbUCCdRwkxFsWfu
63iQHE1f2gd9VKmHUOgez7MmQ6KkwtxmbMIEkERlhg5HCSWKSRCy1i9J++makT4qJyIyvJZ+XD9L
5gj8PdYQkBHSO9Joy+P0uLqxubYP8LsOpnGv+C+bb7C6Z6xKvcOV7fl59I7A34+S1Q7Tno3qSZxp
EBpx4wM/tpgZESxgN5NeEVl/L/3gFZM0+CwuvKJYt0SZchEluuB1SOb5i1zftxqj5h5eTuSNs29f
sQJy/RFMDwBGRuwOItGzQxvrM1jBBZD8ldnyHHWP0qYSO/foTsbPxMpDemVwcXye9mDrEIO/Hg5X
tZpgl5HL0A4NSFauakCIVz6ffxoaCFbz8R3NMX6ouJJ3ox/96zt8tFou7ySsiCrYyYLhz2GoXl2h
EV0+BOoN81kEo4QmP24LbSCGXcLb5/PqqlUrXod43a0wSmPsHaHVnM9sUq+bfNPX3ttymu6GhPHe
eyJTrzDIjmBY9duvfkB6vVEzKLAR+EDI+i6eyjn/t1Gz4IZDjj7o0zQWNCCUhPxzYoZJ16frmi3C
8ceBOBaFkzLv1cxoYqoYPeSQRBZK9+Zl7JdwMpDfy1X2iH0GCqozOSZMgOVZ2piyG2yTNA+pXPbE
AnZFC5ZZy/9zat0PYmxOARmkAavPWynyO/XW/+3JVsn7dCoHF0WRipTNfVMr/1KDBef0fTbxhqAm
dMnHcDkjc9Jac2gk8nhRGjD4EHfj6Cfud6i5DmVd1T2Ct0QlC4cLY/uTVzSy2SZXq+UNrUMd9tbw
URZTIiOJFhYXqreboPbfkwPPmc8t9MFFEHOct4ezI9yFWANX4vI8mcfiYdCsaMDX3ZCZIaNTENBi
Q7Pkh/ab43M3D+2vH3zj4qdySub1dvvNRaQnemp7FZozMlIugCbztX7l8jMwotHDumvXUABmseUz
PXN+PbZUGQgYT4Zwa+zwncTKa1HpSoZesPzE1rB9xjh7HGbMLZEywphlUw7T6HpwGgEbJGO9TZUe
X53yK0y4RvoRiG5ZUAh87msC9n75HNcRKB2/TgA6LZtLh7LFdaTf1oUA6WKCDATGhiiSZD4XGYQu
aFfUDq7DnV0fxeCgcg/49L3KR7NMBHaQQ2khHoyCyKMzjAvDn7I9DjpxDfJE5mTQcsGKxbWVSeXE
DTdeeSbl2RYqJzANvwyAj+3Wsu9CCPNuXx6tFph6WbLGgM/z81RkXnN5KwvAdXPOpGktTsGBIypr
DmcFeUqBcWVL7lZ1lYpS8vYI797/bfqMbiUAVSW2Qe28iKLStxWiyBUs2z9qwL66/tX0ThLl0ar4
ktl/LzVPeWgRgOnjuYq1zhVxW4scS8ApMe/g9FCXgX2imvX43NRFpYq+MlqFJdnPSyLGc33Eei87
O/9T/839vsKIZ5m1LEot2BcCjItuQGdVAQnFl4FjNgr4yM9VKKsfYG+7Gl9m42PX3wL3LT3/JFLD
zJaLMyH/WAZthDsvDpTjpUIv3bQAySyouzYrz3uNDl9AMfrSoST8r0B5vSbK+GVjY7D3jYCiChFm
d5WzSuGGPTGMcb4mEsFpArfB2h7GDN2aov7SYvaj9pdwHMcgqPg44O9yeGJSTDf2QHzjLKCwEpW4
4qrHpq9zByE3nN+PxqROxqOkbG4SD+CRwtxtSB3J+Iltg9tEoXoT52MdYCGQD8kjvC1QmJKGAXVe
APlmyg/JufnjsA8hky60/qkEWak6+AlT5UpNUWlpABPyJXDZgmAv3F8i3cjlA5cC9jZhWzB9VDcB
fS31pxp6LwvAl+eMv5e2OtcLOrodcJKbJXIKz6F5H0Ip5Yj9qcnGETSuHIkB8CJGAh1V5yhTgIfm
w0fT2VqcWTIDnsfYSQyEek07fz34GU1HjVamIPTSNvQ0ebH6KXyv+GedS/AkZKgW0JGDrGwU6gCm
QMZXrwrE6ef36EoxWdEVHqChVDlWEbRRJd5C2sQKBGE+O8ytQGWGA+Fq79DvYjE/kpFja5/YYvvO
mvDEnI6yuZdPEGG4NT1GLdYPotXQcW3ppcPhXHhF3AWX3KO+VAHVWVeaRRIy4ZAy19by0W1Y/e30
yg84Omhw3aOg3F2elRVgW9x4n9MQ37Ijvl8KyUAXm4GJ/7gNIRuaz2URtW31yB0vBqtgoXAztdPW
fBzdrmoFViFwkssKJznG/oT7/EVqfFRrCCQ2qSrYzSVL8vYMkgBWVsWrJF508071ya5QZFng4gl0
Q4zHS9dSTSbf00rnCB3krByqlxG/nVfi5R3SacXtRLZWMIfSSA2jwCIUWmYxsSc+QkpNL9hOwe7Y
wnOwkKbim58v1/goIWNF5UMONpLchUWclFyqoAcLwfTv/ekRWYPFNN6CKFEO4B1mVcosiX4i9eBR
PQoOTYl3FA0Y2+VU97m46P2T+gmfueTsQCJcCpSCHyyWcC1HXVzwEyLJ/lJmtQNwFoOo6CqqBhDd
CgXv3L35495fcojguuv+ATo5oUKoJvVN1NoOaDQc/NOoP5IOS3wNkXlqVAFIbntms4ap357PEVaw
+EPpK2gXMcVH7mDWSe2qI0tiImCNFoaA/BEKjXMfzQMX2vDkKHCbjYmeGtJvYEdammdKq1L8s42A
0gEUrbMiHSnubockvmnd8uc4nvJYSbnHs0394sczf3bLBvxsd/MzSGqJlMWVZAqo9cFGgbq6HHCQ
SV4r5snvrQ70ppAIUQR+OmO8bDO8lNcbHYmCkczziw8xGJg87TeYP55cRyNB5745JGOwWOTlnE6A
XmKiN2nC9j+KtT3tBHpxSZAgl5y0OaNVvtWfYoGrVEM+uOb2i3MYnc93CviQO0Kk9eEgFvQORWNp
dlE4KCg4ARsSjZ+guUdhdIvGtnb+Y3iLIewHPc6QL54EE4Uv7Cy6Y5ejlTbJZ/fu1SuJJnnG0S2/
TOddeUlW18+bDEBVUaphUBVf6KiVgzdXczUDQeSUrA8OVR2E3JCbIIy2QLiP4d9qWo+S+jDxKI5E
PNKFPMA/gMPU8c6LsCw0/7luRVpH6/k8EAPuoMXdBOrCOZDJuNTwCOC2GrVlezjWK/eSEqPu3J/k
vIIfRPeP5IlefNr8olTf2uNiw9IwHFXwFZvbUx89Td2kVazhvd7S2DQyWbn9AG9QtwP85pRpx8oW
egOnJQN+dbXmhoukSqC9giHASidEL6rbr1EYH1Mym8LJOMbHYdbTj/cAqDOICPXUhtsNHiKYDpAy
FGSXv8nu1M8nWVhuDel1Ifdx3iDHhnBDw3Fz73rXYP9Yt7ygyTABplPb4bMMoFY56Whm8hHPLaBN
hZZ+8AEy6zTo50cf9gwW2RSMF0AIYET0Bb7/l3fYiALNjPBJCLSmjgflvbxTywrg5NS1MMj4zUW9
8w+HrMV9sPPFflBSAC0qgzbmdpq2hDgmmiKxP2BQHylMxxM3+tCB35vXCDA8oXoOgq/o5UQlcypu
Mklb0vLG0f0W8SBnd3kj4zCecCWT31pTwv/7dCMSF+FU/m/uTYWhm+2rmW2+X1ggoGtFBA+ZcN1x
xitgu4eMw8hUmlhieyHSD702xbFEIkShlfYt26iI1iOOQS4n7iZKtDj6wwu13rPLcUEFyQWm/xII
qAlNL+Yde3igvcvJ/+neeWTVa6nyFdgkg/i832KD5YwFp4bE9WsXDjJl3LAVIco4XcChfkIpuBSM
wubTU222ZF3VAN7LGRmOhd4xXWBvHAB/dHHkCktt8qDRZVEzjcUun52Ws0DsyKotGlfQBeyFAzIz
OR6EqNuwl541merIIPMThfTIxE+u3mZQeg9MAKNGLkmQDE+p7LILDIlExPgIe0uDTpVtt3N6UtGf
76ZOOf2/c4ZeWX2tFWsD3qd381AMxqVqmu7x3TBb76K/0AF2wbeFJqdAvyOm9B1WNPZuok1BELLu
F6Dkp+4JRpiA/WzWXpuIEATBZZ9gbuSqW7ZfU54p/aLOmSUhyZIph48XMfN+balcbcfVcOV1W3s7
hNUj6xUzXTYaYJktimKtrQX9+udwYwIiKi7btFMmby/JTj+x/LbCTFMF43gFpxHOUdxMXDH1/jHq
nH6FBiQgFay+vueWVgvBbfU793W4xi5VuvCz/r7RHE3MRctBBCPAZUmjl+qpQhRCJxpf9EH3BTxB
jnSuGKTRNo4OsxUL8C3PRu8JPENQVKzXR1z9o6tAOuBb9iPBqSX51ppsW5JN27l9c0cinuhh59qe
efR34I4kH18M1+fXx6aQEJdvNKFAOBieI4WrkGRyEt/XnXV9kfSmhldZnJTwHwWUmNvCM0bWwqsY
uhftjnQ2DrdFGIaZ7QJQvqIQj0UhdCyUUt9fRasX/IVHLRj1HndmO+E8nRi6RVhNNPQs8A5bT+jN
CXSVFnKOkSecyarGyCYMAdN/ZyZ9CngTG1vINwYDdXJFsJpyggxnyXe05wAP1lvwAlxjgFZOV5NP
dJCMJ44XO2X9obtTscpxn3Mr/NiBTE0xFXGBUaRtAozfjHJog8y68zsUjTt2z/f3d8lJaXYNIrU1
mKhoqEpEmCJft8BorGEnZyJ4gsbN2tnKtfeJLyQ4F/N4jL38rO14RToW6RXRb1ydHUIvXgB60c7F
wbqtXIApYtzw67vVLEg093cjmbkaFEBCjM1DIEngo7zXFE0P26kgSPKZeZKZmTQIS1NahlvYxS+r
QLc1tV2ZjqkS9X/iiNm1tls+/MXHIhfbz5nZqmFoQ+amn0XDtcQigJ051LS6OFJCQr1pIfxCDelE
OJBEDuEwIwEgex5N0migHipV3c9x8wGIMOZWNLe2zSeGkiF5+n8Hz4CjGBREW/EsC2qmzS41u0yu
Yp85LS+jHO7dtMQ0IQ6fVOQ5h72/6FO8wTOqSwm1IvXkl/EPOHahlnlp7HsPDRxzogds+37hVuCm
J+zy6w79GLC7fiafEAiYK6L7pHj6wCgOCxjIDXdt45wEy5pBo0zf9Vk4hJYd/OVRrRt/eWt60Ddb
GLfDwgXSujP/YU+E4EbK2O0NjwHUC+WKvypkZbc+Sw6q75wykTnNz1BiM32QAYQQEKWlQ0DRLdVh
YHANyvnoPar/iSiIPYTVHIDvOgG9LdCqJQ+mf0bldryeCXp5eLXHkTaECbM1Xw8VuccG5ahyysMT
8okx/CXNspBzl72mt/YlpzQRGSNr041LEU99mN6yYdvO6fMWunkMRU7LCiQ26AioKV3ikJ0hEku2
K7lckJ8MubEA5xWiHtk9Jq3OhThoFjnc0UQiV1M5w4GcR3VJMN8O9l/J7AHOGZepAL+G0BLBYes3
XrTlSAzJvH2J+PnaxlaJOHIhK/MKJhtxYOa0CNUdNkYprFb0pfHv1zlHsuyVSkBm6ESmH+5yp8mt
fHKccmzuwiKYCImeKJ/4EddqL+YwsnVmhtm32nKTxri/3VTgDCPMloMF2RoyvaKvrWJio4dFNWhq
w+MsRcRuZqGW8gsxFbzUMA2tYFWyCtgqL8h7DRJMLcXPq2+S7UlTZ3nDCN5fn0wHoitK8VzUg9Bq
QwRUmGopNCT7zu/YJQs027ffQhucEM/p6A7aQpAbVcCdQpbuzCryvNb5ml3i3j82hYnBCc3ngGXp
VN+4o5OU/xkzcm3ViG4c2MLSUw3w9GVbfNhDcj7j5RruSwhgW99s093B9KNb9J4Mcdz6hj98IKxV
0Skdj4LlCD/9nYjkHiDWPEd1D99oq7tj+S3QUlN8NsA4fcGCAA+JtpjtL4C/VIPBTATlO0FIDSEI
yqY8AF4LybMIe5xEy0iDlktE089vFQ4dWm45W8I3w9bdc1iqiAKAbIvFjdcj9po84RPUZE7P7vJM
VDUqrm/cnpc+QcAdGQqbwQtbF0vtZQ1e4IzVYL67CZ5W1+WZMrwSSZp+PK4tthomVLBs55YFm+eN
5VtVJtBbgyLLMKAuHCxsFj6RWPns4YM8nF/X5ROp/8/tr+5wm0S+B6lndrIQPJK41CvpF2oA7MPP
1mHII2kOtKp6BIWeFhWusFJ0XVFfd5EQTTk7bUnwn3BPJX6Ve064Ra+HEgfCSvdNGn3KyQBTdeP+
RcY6YMzGc3V1tZrRAxWnnFJ4jho7/PncREPalvjEM1bZOZDWBUM4tWwNitUFGRrVMggm029zx7oD
5HTGR5nukucI/fyX1DvbJnq3W7zaavHrFCRpDMbsaVhdfvHknTJGyA09x+Jl2w58l1EASffAnJ/X
ZDkhEY8Wgiazt2LwhV9sIHJRN/r0oJ31FvnLMNSsubDuKrfMLMNtibggRJLTwumIqAzRnTCl6Kc0
JYsK30WBvAAk+/XWLiMx2MjAuxy6r0igjQDQX3KixO/2OYcHgSfmLKmzm16CP7iynCJqbP+0og68
qScdtR/GaQAUemo/hlaSJpQxscYaY7l18gsGCJ4U3of2Gytt6EZjHCzxJ0gtqgnqK78jNLngLVQA
OxZGWCJ3LV6V0ubd0OQ28ZnMqWHT13p6cvUS1UDQHRZd7+NXze+dSkMh+Sa97kpAczesImYJkUiz
Mmx2eD9QaSnAQn9RpWvUkHBZDS0N0J4f8rbnK916nEtldJKgaXb+3xh5eGagRTZ90Wt6E27YtmH3
ICJOzlBXAWs6m7+0l4arc/LGvEL8U38U2s6Wx9mCYvHXY7JAhm6XzsFgbooJnfLF0ZEtyD6tv2SV
m4Bt51QKYLF9Yq/KDiGMnejhmN+/xM7RbOBXfqpYjwNM9MZ1tA3PoyLWfbH7bd6Bwj0RIwxPrh2K
uL6LpHC7COL9/w9BQMxty5OgOROjfTuvem9A/zWImuAQgUP41Pr5Vu3xeCTIRmL/d6GpQ2YBBy/N
cX5yP33V4A1mFtmZw+HYAm2LVL/PF+OGrx4SkEWoOa24g4rdj/HPA5x9CR0HLl1+P3GfADLq46nA
amO1gVOjaESN1+jUutMUWfnHX9Ok/fm6VIqoRBfDsRQ6eCeNA22VebZVURnODEzEDdOliMWBA1K7
6xH3mlfCN+iULJYMDzEIfbWWecZsERP0TI35sj4gpn8otJjypMIXZysEVoCavCNmjxzhOyEn6dwp
+O7II/sYl/ZN4sj5Kdvqh6vzXGd/3he6K0JOe3Iqi66jxAAq7P4HV53ad2MX3dC0vknV2A85VCpT
ufOUGChzOYzBO9j9YgxyqvEt7D3yCbnLLDgMjW88pf0RNcDJGV/3BW0DBxlZHbJfVzuhqWPjy7NW
xWNA4CHEjY7hNsUvAsdD524oAh84+o90G/0n3NWMkJFaB2pw5WaW3Ya9I2wPuRx1eXfLYDKNCP86
OFMPN2dyjnPqW/IzFVvYIrdSj9VAGE4vOTmbk3UCQUSOJsa6HCGX0LWFzu3LthHtC8z+UWTHzMGd
6Ylgxl0hIhI9iPssalEUm/4JMhEOXc34ZA5skhKWS5NE5X0M9V7fYnzR7Vvf/sG5+nGpkLPSJ2dR
d6zZ8x/QwEEBXRF2b1QM9BoEH6uOlA0yVq+1kKfxUM7frHHb2PeDtG1waw/Q49AvWS0uX74cA4qF
ETr3BS/vsdJ+BvWShu43vvvon2QS7QNZTUR8vvPpOilz90tb2VKs2j6dG+0NxtaWqdApYLUzpTe+
IARzWeTJa7W5ZE3QPr9ZYe/ygDjdEbZklIr+MhsTW5xEkKJ5MsHtVaB6GIwGjxFktuxvZEOIOC2f
s49kmRcfmqE4SnTEzzvIyB4BuiFhUowJooKJoi02IIMa8YV8Z5IvuzyrLHjZ/vhQRu8SYZYzL0Gi
bgeJspH4OdPslwKY+jG+hdkhIt9th51QQvSz+dIPNlMNwjexecoKwjSLy84rLlIp+O6OeXatLcmO
k9LGOIR1zNj1qiP25i9QjDEDkGJwApTLM+m4NZMQqT9uvnKnNmRfwfP8Oi1RGrVzuZI0vcLFdpMU
znsE8hsfL+qCgBQlsKaNCc+pEr5PYynSybOjYh7zkkFm4Am1ikSRIJeDUmVAfxqq4E4+W7In5IMb
Bg6gisEAOoTOuIIZy7l1EY2dvMHgIx7CEHc4a5GFjYRgmqgAUisN4RuOExN/jxaCGUJF4B6ZTO+/
KbHLkyg0Nor4FlzRHakuh3FabpOtSdI/o7GnH1tW7hOmIr3pPk+g6lgQ4Gcu+hgV9Wqkb0PQdEFu
1ywctS5h/wfYzVmc6drLXCS8SkE3MGmaZU2uvKlz/DunbbPIvuNoXszZxs96ZC5Gu+p1tOW1wNNY
e727hFpppWIzK0o+9QH5eJcdOpMCmSlaU4hDQTg3o0zA+DK5kYlobpROsE6Pl2IeeLLtUNHRyLwH
yHdsDX3x9u1841EXe4aLEQNd6qh7ql8Y+7HAVcoFQVH2bcHbPc1/e2DTI/xukicLmI4p8fzpCNJn
bkhJ+75s/3zLvshMwWrXUNikTtc7bXnoM9exs7sOJvdkxUI2RNZO3T9CSBo6OT6hhfIWaAz6bnTH
+bm5bnw36ZLWgilI2lZ+lY7/T0iuzL4ud/XERdD5lSym1FzcryrxVP+iWcXc02fPiHN4d038vSLs
PexrjcxFJPQtnI2xAlWWm1W/s08LNjdEc/AcnugZ5Cshdl8SYxpw8LxyfGQACSYXzEWHQRC/SRRE
vsp3M3F/oT2swI8ccy7vxglR/ldy1Oi7by8syPuMlbyVzMyRCE8JuZFPNixK0k9ojgoCzTzMck3p
X5tQVTCffYpVEa8jz5AS0bpcSlqbzCddE0gVBrRRyYqF70XQMyWjfOmPeTMeg1QXQfuMS5oLn0q3
ZTVVJ+gBxm1rQifaB9dHsQYfR0VvQKhhXr+IKOZlGm1hBqFOU+MUHnbgq+09lFGUjP1zaNEy5uPG
CBHPCSvX/oOBR/66qJFnNco6hk90bK5rH8R+6PEYBlzrr+GRACK/Wa0oV5e5s5wkU+cGSxXZvxtH
ML12UhS+gQhbrEvmM92a14YnQI8fgAtp5qcsgk2EpxnxsEbLIrs7BK+Uy9JoB8dj/kTVNjEgMjn0
CcmtgOtkQIiZdxgRvgwAfXpFSY1jd/XCEazAzLDhqualn5b0ocvOCICpMChUpC0V2B+NTTAN6OQW
+LK+NpYrj6ariVHixdixm0VFOf2ltl6KApm/qC9BDdChexjuJ+ZPVjQVSELHJd2w+NRhTWcuoS/e
FcOTo7F8UXvt2+JPGV6qOK2InPcGjvGjXGD+Ms4z67FM3SthobzKZektPTE3jhsFoGcRgtK/jzyv
OUXVp0xnFa1MIQfq2VLY+HWn/95tvlRVzM45YEu5W7EdmDJ6DniJQienMcCYeUBPjTGEuOLPkd8q
uznTdgrdcI6YaSPblpIDja/0iWTPvL9szGRi+Smxx6rX80Gr7d9UHQ5GiU4wCSPPCY8MoUrHVgjF
+u1qGGNld4MThNUHT5e3se3JlH/cwTPnr/sc7x4Pb9bL0WNCMEtbOMYT3+n0Bw2mnrY7jmUbL2ip
J376S78CapvSCJ6VuxnWqdN1xluGUQsoBr3igUDCRjOl54zXCyjTAp6pquBzpn+wk6EGu36wpDep
205w+X/j5BrTGSRhnaVDs/ET3gc9iC1JEoiw08mflzFUFu59Uf8KmvuqH6c6De7WPJbH/lHQ74NH
+nEc/K9prHPtzqQhs6cWeSYHQX5uabn/L3HCSj6OYEG4YXFgHqrUnbvxrUqogGHoOt0QnlP/fLe4
p3cs2pL7ugUyCOdJcbWmpGufVR5zVkiFsIb0FJChCKl8kcvBzMCAdkfI6kmneRFoDoScHHhn7Ori
tH4YoKj4ze1Q7E/K5lEBGmNEDZF0lGc1ejY5YyMhfjYHaHIFdUa1A5weHeP6O+WZ3m7MVC0g4Ymk
7l/3otRDwkEy8ASePm9TdcyYx54pjPPpunzi83ltOIc5MneCNOk5diSKVN+PYCdtAKTd59laeZAo
h/iy025KI8kF0cpZzf0XPQ5huCIUCT600viz4pVo8gS56rm0Il3r87FCA41H9DMPlUGGT0nD2ZK4
99VWeZ8RWyUsBWjZNzI8oK8qBbxTsnQ8GJ/REo2Go6fG+I4btkItCNgKRlNTTBC2UEwjiSVlmgTV
HxGzyCH6g9xrQtNncpfadtdynXm4+eHfUWnSW7feB+PoF/b4VOyAEw0yscbJX1EF3z6+06wYjX3T
E1txDTZvLZAhYI4ZArecill4y8XmVmwQsaG146wnCJMs3bXPctD3jIJ5ekQswxRAzf6nY5nW2JcJ
6kcrKRfJPITtYDvIZBSaa7yjWVFWLg4KSWFLw/Io5MOc/R/KCG4qJaumwEedM+UHQUNsNxkjy1Ai
6W9Cf+c65FNO8N1sCAACo3Ry2h4FnwlMyDGUoopNcqD81WGc24ayBlMC5YxToCZqWeyUDRTFNWX4
weR3byHvJZl0AWsZcWkmnB3UoXSGZDP6XE4Rqdn1Jcl9StqbQN6mxO1BrtNqmJmWGS/4QgjAZ1np
6rv1946ZYw/4clpQof2gdTodyp1oEfE2bUGn7O1z3erLYggeIB4H8LtlB4QROpqU3IfXLgcZy012
E4+aSg6iy61oXChxSGrtgTDX3cHH4Q/cZ6Nbun7JKaYscUabutcQiJ1MFEjXvpqvidwlikHvjGJz
7R8UVChMeJIQA7Rgzozc7ucbmR+vGDoNl38NpcPRSnAI9Y67L0zSqVrMaKB0DlO12i/BD9eb0zNv
Kmawy397Hf2x5daPNyXELdMl2XE4RgVfeiFXL1WANVWwRg6mnXRc3EH4XTryRcXlS2MAymTvcqqr
M9QOI6nEigHwYud+zonDLmAG6zZcOrW9CPPHTgYcg+WHXIonC1Z32CmeIVT6o5lvulb9krf9wKV4
P2HrfYO9Dx2AtyGhnPMdakVZJ7lOWRrQPnJMaFtd5SSioEPOZvyCdcGRY/MocxKmTfth+JvmApxW
Bt3NUCL7SprGhxhkmJHgqUmxSNNMsIYVi6hPugKwxW4xIvgmRpoOV/j4f1T7sLk/EWdw0NivyzA+
fIHXZuzjWd7fbRc80cOQ54f/i+Q37iMX31PENWh81CYolSVoaoYMpton6SdKUIRDDdYX9i209nzm
xTH8Q5iQiofhG9AHuSkJBis5/dgixGG5aEjZW6qkOHpC91+tSuYeYER70p0ccMGFEoAo/P/hQUeL
29LrsdMYVGArE4W9cu48SuwbEZN0EFmwzwZCAXiu9vZdlAezVN5WsjViTNaOOvKJXOJl2QGFqouy
A8mbQ3M1aYNdIRkRk5NR6LO42aFkGOH91Ax4JnxAAvBWDDmbm9AL8DKzMYiARzbnplMqYJNriCy6
r7u/Y6QmpCSjT4GUMADP/Gq2wfSv7X7pwNBkq88MUufR5QgqfU7ygkoryK6EtJH3rN6dgFAPUkpF
EWlOczs97y8X82nivNtnQaF/P78UBNAJfTC/3blvXa25EFPtPMx9ja3KVML41C7/psFW/zwx35UV
sz4w22D3Kk7ROiWxPPdpkIF9f5diTlnKDWFkGaXTRmP8nvww3Lm9fjUXh1I1LmZVHSKx5gYUROpS
WumI/MyNJipnUP8+mw3UV0nz5kqIzPBnlrrhxUEB4FJV3m3xBKlS9iO1nH5w4MtEsYP/joVFVXMn
h0rxMcQX+SwagZTKYFrlwVaHeKA44bVAZ+pXg287akiYzbOteQdtM2Eyr3vl29aPI7M5blrDtLvC
okOO+uqu/mfiRtY0Zj/R1zlo+KQkKl+oVvzRD2r8wT3NdUonFk5JdkZqeXUYxJ87Cb40vtz+QJcr
s5KMZKZrXs2sk21nrpe2g9g6LqqbQ6yrb/04U+PW217EJMMg6kk58qlX6njFQpN5WuaUHIjfPgCm
Y11UaB088BT6zrqW94gpZ+HPJ6we8bmfKfh1xvoF07OcqpMJTJByTddksfguv21ORY8bzafDuC/U
n7+vMX4pkoUSJNQHmT3pGm2UemCmnvMS4MT8DalOkJxLjjXqhTgT45GqOnEclOd3stOnUkuoI8md
R7A+h+HfDDKj/knHqPPTQNz6FaXZFWkyszDbVHZbsjRzZONxmDcQ6+Wop/kp96Cy68RlU/BPWqa8
/IqytKs2LB2fsx/l16Mp9tKCXRl6sFq5kz6Q3DsmrDeQFhIIpqC6PQPjYWHzquZxAcshnO86c9XH
CwQ2qEoziRxYrCXZVNpM4/5hRNwQsggGoXaEvk5+t9qW/K6NiYPDThxq1nn2djHepU/UEukyn38z
yG/WpRM7fnj8HO16BOMNCMp2qqqql7/1grfF8sXNfkQrm1/RIy6fLzb07zqJLIWGhCOnCtbmwq6p
BU0KFdCTMjR2bZ8jN/gD2ihvzlsOnIwthLs83CEI1jNvXPTqC6WbWT/DWfMaH5t2xkAf861XXmYp
QNykA29LCMfDSZQI64cQdaxfH9IrIjSSIpSxkkls4S9VNUTgvHWjn8oPQlbOqFBxkar6jjFHOF/+
83NXv+6Hpgq1dj2SyQGmvQbqyj343QfdPAk2Wl4mVdzAM2CADf7krwPZghBvvQDTU5EgfTgB1AK7
MQScHoFfTpuUCQkgQehhR2/Bhkwx3HDW/VNF3/tSqo2DTsjcmqpAFr69huyXG9KuLFUq4j5fmgDT
7rOSb7wHCXueiFxVvKq7fsv+/VLK8zoCTeFnIWZRyQZQm28sdOOrBfRC0l7sRT9PfVPyDPEjU7mJ
KA6YRo6S8f4WygZB5l/jrmCTB5sJZXO6yB9XBAcEsW2xCR5/7HwBlBKZwdEU+DxpBrCvCGReSxLK
Di4uKeNazn/bgtrfPt6RybI/WmYVtGYlA8tAcJmGjdyzSOw8VMB/IZulA/qvjvUkgim0Y5WZ/m7P
WGSNTGTQpewIesnGB7okR6uqIRzhsSkh7K0D429AaUpW8T0YmSh+L8VDSPYh5IU0u5WSx0fHc+Yb
uxEyNRQXHqBZgjyS+LKCxf2HawvkwcxPqWtvN+Ouv1cTyKA9NFwR5mrJDh1/caIbH1aVmBGx9x6W
thjwmzEqhlIsUsDOK/1Fk8nSTL4aFJ+OPWXkNLCgMC5JdFL792DdyDtawNNxvxUl0qn24vyuM8kX
MGp6BH02jhk5RnbvsI/HSB0YcYMfgYEEyxE/I3vxMh4k1yXGumN+/CUFNmsZ5ZqlA6hYcYJl9uiw
cCm3lwGm14eRLVSXz8Gm/Q4LG8YLSHthWcEfLh5tcL5knGcvSxuXsF9e8Bd8EZ4YmNYk25WzFjPT
RsXrSzujdTOPM/msMkwep2LQYHZUR1qJKH2uXp32AIn0ZNDnsG75WbbVuT7AYMsD32Y8DTsPPe3E
lGp0XBqms2BDKIwNLNObFb+quFkIxMVsk8WZgTBlDbKwDp4iqJPxJxleF3MSPruH8z5XxgyUOamT
9HBwHtDsPLQ5nzINryp9nEBFhFGRPCEVu8LvLkJI9/W+cYBp2aShg6yKruxhqtuqBzxrgp1AGgIE
k64jWU2CSutdWBxJKypmT62RLRXzrrWPdrb7ZYooBFkxvffluvbBqlcHTPBdV+0mbRDCmOHDW+44
t93Ha10NJpg/nAtKlN3h+8Gy/vIfk60GzDSYvW1/bs9XRPLca+oyHgOpWmBqAKgLHbPvlMMfK76q
TCZqdk2VNEIHcJ16O7CPN5i9SmUiF53LsrnrnSyGdP7AxmptGeiWhbM6NNjPpiSb+pNx8RRpKJF8
/c+ybZT1+B8PnTMCpjvMz66Ta7xxdePLphsUFHxu3thSyc/b8zc2Cz1pr1u8VzK/CXZ9Q0SaDVmP
SGE+7XHmM/2jpq43lKAWkzsV0jfXELM7Mn778AYBrX7t2Y2Md9fqduJHRnB5XwJWFJ8G+0R67cB0
zzJo8XvlxNU/w1OtB6W7TDmN6cKSHcWVS9q2w21Wue0/Kv0Y0itvILWESzQqDNGgwjrwwMe3FYUO
rmP9lVd3b/7fx5IXrU6ypgqWDmL8JFuKHeh4aGOwD35/7QQG75LPGd03+lYgUC9QsK7konDbn5ce
C1oBIy71waFSrCBfAZu4P8Pq1t7TTjc1/B8NycsTDYNZD2SvKLychXHkH1/WohmG8BAkTiOg0zTb
F44+qU8/POon7d5z4f2VWpUt2Zi7ZRP6pDzIiI57R50SukbElG+hWejYTqvyeCbDfrs3fzohxOVs
37gdxOs0zE8mPkgX171Qg6PX4UThyCn5setALIjVOampP3OCq32YX5qrXl5NQzuZ3oP3xAHfQ42a
xzJPHNUscf8T1wXSG6xKhHKIgaSYPJOprdL4utaPjcTQXCYm/+vuo1ltdRJQAY+xbzXOrIJ+h8LK
xT4C7E8nz/x0gu6CnInAuoX4ZnFPc4CwJUCuUWKRbW8B33rwZGp1eQMKlzERD52ZsrMWa3zXVHZQ
vQXgxMHaa4122ivzB7UVt2SP+fdC7JUyP+RSz0bHQcrHg06mjGSVtFivyWZnm8qR9CkNcFb+oXPC
Iya2+ZOU6uGL2X0vcViZeVeWHCQLvK8MTM1rSsTVnsehM9SjVz4dkToUkzGtNtz/59iYyzi2bjgl
oBpVzH3N/3Va0BZho9KK6xopqhmRPeU5ChsHPknIbEXwa5RhXt0jyH6GTJZsDxehtOnELSVF/8bo
y1hRtw4Fvhp2D/yV6MXieA+DfUyjj0dCvNxMsSNJeSpkm963iqwJEatkr+wm5xtOfAZegg6SqCf7
/k5+muUIpn1PVNGGhWusp0sTAUsQkPKTlDAt+m6FeE7yVjW22S9QI50A2dTeo3Icp2krHm9cSr7j
vpLEmt2P8/vOa6KrHegsV7fw30QRl4ax/QnPDl+N9ppnHnwXreAoi16StkJ51NRgnEs/25VH530o
P9X8csqNEsnlBfvbhl02XIJglHMofENtSRD3CL8I/i69ae6VRDGfHJKXtAt7hMzbLtdmfF4Rf04j
6zHJXs8ta520uz9iwRUqt/o5qibmFxh1ahv6dSxF3N9+IkKGa94XIfdvb+8wrIp+HotzKzwCIPpw
26PEeufSUN0Yj3FLyvYuqxk5GpKyx6oWiDM2advbXqVD1roQLrDYr6r4o913JC6ImS724tnDfWmq
eKVKd6f6BO/stZOfLGGJMv1WzNfUPFY6XKsnXTi2H3yYg+9W3a8ybalDxXgKYfL+JtWjU2owpR0k
04r9C3OZPq4MC9JcrNL0Lb0Bj210IBB2Id3z4rcWqAsnuLm9TcEwIeCi9lO9PHq9MpeKxEwNR2BA
wNhjYuqrtV4DqECdFnJTSo7g8xfKNeILVcrgHMBmVDBv5HgND9i0beMwgynDDFXNVAvd3v6C3DIS
Th/27NnGFU2yjY7v36/noIkNMypRTRmWCe/0vcQyvB3BQQEjfbNxAguVB2laNH/hO2q09UaJ9MLa
XbqrcS8bqYv8HKyTOyg78SmGSve6jfDg1cw/4jcDGiKPR+jtvUfbMZf8KXKWtDDh4pFmIOogNJk6
gARog2BTfI9sLud8dyH/SIhJ2yJaBR0YmLoow0GBAnhBbokO9rh0vj2SDRLMMr0b1TRv0rfSIpdy
5QAN+qdtXhgNp/35JU59HL0NvZYUpeODosj/65o3FF+qmNdUoZge2eILr4UERMFRrsDLfbgMNH5z
aROCZ3lRke+k0Gf7uB5DxYAzRj9MXO5WmyNEFoZEcnBGYPgE+who4wGrbuB/x+yXoTzOS81sqReZ
RqPHmCJd+K6fUItvo8K1PSzt//FG+KDFGQ5hXASEsjdDawnSbit0cyVM0x9kOo0dOtTwR3a3p6kz
R3LKapz0/nCOcuAoKyOAygmbJFuwWuYrAn2QzzuA1U+g1OHOCmfv9DUCQXb48Bn0ZAbjf01PtLgE
oEmFCgUWxWtaCMvWyvWwU5Yz0d8SYqLtEUmrGSuJWX2Nb5iBF/u7KveSC+7IxLtI9C8BLgd1IKqE
9iPWHmPJOsvoK54a01UL6+AhLm0WwhX5SWSbL9wpw/FLbCZEh/6IJ6NkBARk/otnr429niHgknTh
BeANfDEqvZECl36T2qDJWNkIvLOoNdvXkq3rXJVMzhj5Yc3zMj9tJ3M78nJH2hP+CqBgzCRrWIig
X2xfdZ7Va1c6Yfvw3788Z2R3hEJUdDV8FTlBbMkswU/jMHfkA/K7rpj6Vxxxp+t7yMFTXiYHIRKH
tgtFnYoqp9FFcmuI1dgfB79phug/5F42q36Q3AnObsxYWiiIVnCCjBAeAsK3+KQ/jbTDx0fLmMH4
twczqAfKtSEo3bIF0tam3nWuku0T5YZmuRrBRgjc2YZ8f40rHCw2+IWemxzmKXiJteTsfEyEIwRN
lmrNNLC7bQW2pevzUlUFXJL7wGueh+PFl2gZI2WavOHznuh1rSP1mavOkIPShlDnVoACfi8iHbbB
IxmNnkuGZDJGtAKCiRcUCjhd8E5m3F/CYAFYMtM6M3c1vCMVixHF8ghodN6ih5b6NAAzUB+o6JWR
/mOu2sDx3Flj1mW9ROMH7V7bi3GQ3fjZm2U8Dh7ov8z3XK8IE8JyoVqJDCqQRBGq7NJbHXvKLlYM
dfmq5DJTYR3/dffqHd6C4rlYeL5I45aDA05icxgR6heKzINyslf1hPWIgBYenv8B4MP/M+HBqfyt
9UESuxq9yHgUW2KQYJP4O/J3lhN1V4g0i7o1VdljXR1jHCiXTEQG3g4D7BRh6kg2OPHjjNptOHXE
Mg5VGLVQnVtnkxE6tVhm32ce6zAc7h0avi2bWRwQkQO/73gCx5nLDqo/MhCuJ2oizCP7/651Vav7
QXnOJgm4eF43lSCyIMW5jnQ4/Nigu7bAu6JBqwa3FjO4YrjXPt0p2Uak5yFQphQw/80LEJZw/8Yz
vcW9qWeL05Zm/grCss7O6Z1CNCcTtSb3jw3RdJC0Q2Je9kcmfIyAbADqKbHYeWvVd+SU+dEKdJZS
6ei1bjVG2vXJYQbRzcXrUe9eYsHbvD1oK2+EdjHD4ctUCv1W1W0/q/GXIQ4v5KOe+PPxe8vL8u3i
VLNr0KPUU7ZV/bx9EFp9iHRUg6RK2Vl5Xcc6Dz9YCAHybYlnxyMOyqKRZ981F/fOgsY7hilLj5Su
XKXpVyvIRNgwsz74ZRnYJES5C7Raa5NyrA2hfQp3AdP3bMJMRmVnYGYz8w6yynY+5PAZMMRoFzo6
O77nXVYFrC97AHZnaetHXQ4VbzWa9lMOnu45Q//vFSMvL6t0eD3McLt/TCxEC8GMAbS8Al4kLQ0x
wr8twPo1lGuYXH/2jTIm1LWdYaVk8YmDLJSM6YLk5uP3BYK39LlKkTjvaXyC23nOowPQHUvsdy2c
XuzeyCWDOBwzfPb5Dx2lgPlC2rA9bBsq483pqpgdPyxc0B5k4Qh8+a0PTElOifUGYhnkRXq0+rxd
4a7KS+IMU1F0CwXxZehUdwODWMhIwUtKYjyH8kwrK46x+gjsrQOmnnsekcydfARJ7IZRyNqEyC2T
N9oIoj+xhfzeUfC1PCHfA/T9t4hTKuMYKKwQyk0ZqNA5EiJ9yNC8aiXdWFj6O0cWu158GFKy62Xf
ygV+SGQarnMwxPpyDBuoUT515sw30TsBCRZPYNr14SQB1jaIyKwz5RHmajbXwtHm0oW56SzOOgB1
NOUoLnf1kNw23R2qGnNO7khEQRjnP+mkjcT4wqM4gUIWcQAmIoj5Klq2rkRnPjrvIot3moRs9XLR
e4kQlZuM7z2n3Vqh6KrVRJO+Fkfo4klnFKPf7Hvxy3RDxWuI1cB9bU1kuaUPVLao6vpfNa3jaXcY
ICh3FGaYgTA5cJjIB6Xbn2EWN/r2hDRhbefc0GE1axfrmsQnevVsB0x4Y0eZOFxca5IA6z0gZ8cS
G+hjfbfcTPHFb07H7ONe/RSSU40ANeC/z4aE3iY7klG3RzKRcxSa4mkmCZ2BqK+OeXdtZWRzUsJd
87u+vUsPCOikCPbQsEk3dSbBJJa0jfyV1UKCK4PjnW1trOp1auo7gAt4+z800pwF1BMc9ZxFUVvN
vQGfkJGa0uxi+70SKKP5odHnoY0ldj7MvVPzWoxbgaIJvIX6TfmTDcIbo0uXnVE2EMndqx64zJYv
IqY4ELTxwLmr/oi2LINaAWqSrtAnq2EypEUXIEmoP9djnpwZzqUdmFaITNttnS1PvGGIfZ1tBHmq
9FTqggQVsErBrXVE7I3GmGrj+WhX60yz32wWSAEkT21swC8hz5jIaYLrYTyuWkOmNe45g4myLmAb
32OgBbRSQa/ls+ZrM3v0eyqpJ0eKSS78GDCFtiyRcoiOTu6jD3R2Q/Gm8eeb6QnpD7TE2qhOIYIe
GTijLVndwl8tz7mE4QV8LzqUR/1MN4iqiGGn5ndQSsglqu9olcA+ZJLW+7LsB3wCzPgwXxRgnx2l
u6+UCv7aoroRI43FfVFQ02eOtQr02/DOqrbvPLYd6/+YfyAT4Ohld11IVZrFfFG6lzy4UmPsuddY
mJEZIBF62pibP5esPutgaPww0Cyc/+F9HyqMNkBfxwI+g4LO2JsPhmKyUAiORQx8tLqCD5zBcbrL
iWavN4eihetP33h6mxdUxUD7Ai0spS1GXrPZ9ebYo3vivOL3cvDTgCuV1uJNY0IBQJKXhDBLAiPI
hmnxun/blHYdz7yVO3l67kpUFiGjj76WejnTXLwmCBRTWbr0sRs7swvVzIqBg+ox7USPhFktu84s
9RBovkiEbgfTKrjOmNPXVYUDJq0YOXPNl64VWrsYRZo0AvgaDzIklJTfPWPgajeNbC45SEHhP6ps
/46VD5BVw/8XOddvHShxRWWLuf7LaMV7cYg5XFdP0pb2LqE8bMPR82K1T599uqRk1jg8KaLyB9jE
zqInWYgkMWozlwYh1XxLQvtrAgRJ3TpQbxaFS739zLBW79H0QAfFA1sJyGiYYAT65rEfyADROWac
eDtAkE0hAJDYFemOS07G+ZxS10SNEgIyZDBpz1BhKShRZo+NJSxn4bOnrVIELQoXLjL546JJ5Mx6
mIDeQ0kmiNPFavUInSRxsabZCPXvkluuR+l1gnENsviHDI5WTRQYjSC9w2JWpovngLje2mk3SIUW
Hbq3j1RViHtoqLol7rGXCzOexwPzuMkWLmh1B/j9rOUefKMJquLfCI78fjZfA8waxdjL1CyJmuvg
Zwd+7qfdaV9s04lXxXLh7XMv3pyhTVopbK8owwOr1jvvB8LPl9P2lPik1mWLCG8iDdGRjJGc+8N8
MaYuH6z1Y6zfpXTpTEtdkezSs3xGzfGHThcE97J1J9ojfXyuQfdveXK5FD5yzfhjZ1GNOQrE9dr1
ZbHneD28IRzvUthyE2xckh0S0uMEQAtK3QsaTeTrbGuIr2EGreTsOimNDSe+jYnwFiOHLdeE063P
0dy0D8WszyM7i9S6HdnS4dGQxGAqRwkRP+Ls7itEp4B9rqKLrtcDG2BPWwDWjKI+jipW/lzbQzsZ
+DqZYGA0OMb07odvtphlUfP/lWhayOeEcKYfzosBI5rKccGggUxhzvum29XfNvDh1VaWU/Qt9fDi
Lr1fH7vYDL9eZfbdEOFoIXFXrZ84GmdGk/if1bNkVjLbGUOg8ZAqDPbvUCUAPC6Oo6/pbu1bOvcy
REjnw1CXY1sZjC3+YgXzElUJX8MyboZQR6x2nvBq5ZIxR489JD7PDpUhLJrn5jST2qeAp/MOna9G
N1eiy1XMjwR31mSqWI3x0O0O1WDJ9nW8q7ttVCZSIjtE611DW9PLetc6L3VFNkbIKy/Z6tS0HV+o
WHhGHs3lisyGuAx3AvrTFCNSJ/vm99kccj8qig5y6dQuDM/1tLoA3RgTmbZ/q8BCVKN3dw7/pVJ+
tavP+moYvE/yZjGYYvcQYQ8WYr2L0jTO3PhGf5Ashq8RgRSjdU/kPblJZLd75MlwmF4QpPF4YdUt
bfLdPRryzDxOphNTligfUKfch2tme+KE5975IVj+bPuWCml+S7UQGdpP9IjmRqCdGYJk/lKwEXD+
jtlRjUF8pdgHyMY5ei/wkuJ0OjSMp3bL3PNC0lC1ZwtkIBc7EMNZSXPp2IEtcBV+wgAkrv1r9RfX
edWUw8KhqYte/atBhJP1lMOMqnDeY88jko/ymng900dnomAmcpQVhWEkvWoK8R9p7FAnV3emIzOT
4hB8oxaRSkRkg1/VgMR5ZaLCgs3NnBTRfPCQpjaQiCGSHX6PQ6PA2oxurpz5KsR3PHYdCwbshUJJ
9WhwlSFxwU38JFzvrVS33u37TJRUmm5ahOoTdCp4vwDUXUqaq/FZ6wMtPWS62NeNmLtiuAMiJLp3
jigrJy+6CM0DNkK2geuLHhOW0Cnznsvd5DE3BlFYrJSyespUlAchreM7cezjmDxqU57Gs+aJXT61
5ZkEz8pbw1EdCoUWEA50oB+wTJHliNw7jvcMxZdLUOZB/rIJVzitSMXgPEkHJaT1P5HwbMvQQSL0
LdGuRFyN7CsfzK29Ixmzr0+wkP7lj1QDpyiIQ+XSU74tEBtv17aQZxYk07/HE/mM+MVmbzVNAshu
+a0ArsBP6kFD2i7ASkCCLzZLZtZ4PNaLWtbz/mgTe3ySJk34Y5OMny0Q7Zh9Yifft35hAdeOgtvl
LO6FGA3M3bm/ACq7eyJVp2Ool/bza60zEvO7FOVFYWpzqv29ti3lw8wWKQis+JGMmu6AqlfU9Oxe
y+kznN3TbDzHNaUg9DiQ8m/hUg0wd7GJ7B3SR9IbVQMS47yd+30qHy6aV4/AorBcbRbNob3Ld5Nb
k8CgzNWvv+3I7w+p7Z30UjqMs7emFMyymISOcRkdx5mjb/+ehXk+7NyQgPcBre6+VgVy8pGWZJqw
Tgxn/6BPCQt87387GdxkRKNUuF+JlVXoVijh5aIB1it4nY3vi2+MgMnTREHMuC9qHLgR5bvrV+J/
jGcgMUfTzAzPnonQEADnpQgk/Hq6RTBVrLhLt6M5nwzmb8IKu6stqEVwWIZ2B4MQeggaRWVZ6LHu
GoGOhR6VSNwV5Jr4bhyEOCS8AhmabvkxK+4olFTTWKd/06nkkcZhrXW7rH4l0JI6/bIfRQwACEzz
CHTe4F769ES1lfGfu9aJL+Np+m/hsXFSx/YK6fPEhXz+kdlK8Ljw3os1Gsb+sEFQOVU/o3zeTmVf
qh/F8IJmmfAJP4/uykMakmal4Rx/l2LCH/85zpU0Ll+0wBSfxt4PmuOKLHROcJRukgLwoNAA4ZC4
cOQyoTzbcxtQbB1dmLt7SRH8AxxYX0Sk8pg2PsngGx4SSaf7KHZUEl9ZVR20x6/PeRZCnED7fFT3
ELQg+9kMuql/X39JkarBplkGYFyEB5FJq9umuxC8yZN7Ecp7ZW39i29oczOIpxibtTSaaD/m+YlY
WUJgq/ODud6GeoJbxFU/vTEZtvfFiHnSWxewkMUM4W0qTBP8554RMA3Uvo6jrJhEJTWezH5smI+K
oFDOFZbNz8Dm7cw0Jv/CEgPpevAgu6Rn3KpiW3ytJmg8wJIB1Istcby4jPLzo8+Ub/uwc5/xhlgk
qdK7Pg8tvc1ToavwqzGXB2dRW8pKgqg3NUowFxZFjVfK7VeE+NmG1yJE9M7F/SlWqHYsleyPL3Qd
3TLzH59aRkSlG6M/25eeeKYRGID8T9ZZDG+ckeTBtuBCKG2eU4AUxe/uk/SYQPkyXsvZ6NsWzxaN
5GCzVFtj/5m0O5emY0WYbrm9C9lvsM6OzxsqCtIUOUQ6yUs2LcTV5TdQLmATjKyCMJcIAOhjtqkx
BMCEihfHkslUdCYKofrN/MHq7CTXsLNbuDFuiFRs+lMVIBLdIHV0J6y67MmoRu+a6e9n7f1jzKVA
RFHsfHj7Y7yseOvt59PSGDfAsspPhH43MaK5nW/RWWBwQMsgcCKFs39tLW+VohKyE48WLtsI4k4n
k/N/AKzKbZlN3PQJ7m0EUeTjxmyIyQpiGX5C0Yf2NETZXhuu+56Sa7/x5J9isDfdmvBjxEDmcDl1
XOCchGMAaqKzThDNLrzv/yQh++/0Jgp6WuITw4Eq+Meo1wHxx2U/b0NrUEZRiFK9kUDs2AL5FCIT
Q3ffqhtsK1OhCmn+liL44HCp7TBloGueNwL/WSkzAG0aMu25BGo/HcdoOnNa6rCLSLHUfuEyORV7
5U8ZRnC0l7bh/nBHCxA7rWvhdns++u4pLxi34ty/bKf059fw7SoCU+JaoXFLyYPFL/JPgKqjd89F
LWe6rbI6dzgkPEPIbK+sKoCbjnM/fbRqZHWkP/bPDF9LTOsMZYGRE5OBqLLXh3bfvqIJOcQ27OSZ
XYKi17128jum1IxjwcykNyvAeSh7GTR3R/cwlt9g+1SbU2MgeTsmtnGPIX1IfFg6YKDzJ7DEc1JO
mKsNEKbrCAeTZ4NWGrFnCbGh7gSy18ZRzQ+E9QwhLHEI8rjlQoocYWjIZ5ptzWYfQI41kLYztKNU
jnoVVeFYwZ8WOaWPA7C/B76CGIis4g302td6WLDiTvXb5V+VtzmZ7jIfEAKRgn+dn4nD+2TfarhV
lez+PkRDbn9HbCtngMAfOGzSTOJ2Ympu8VlC6DD3RG2NWQa0f5Udv+yXKE9so3p57S5loi509bmC
TYt2iA18TCyCueSxG0fUm5MQH4U1ELtt9WqIAVezryUDsHMCHu4hJIYURpyMOGPeh4rly5aWAkza
iwDVuns7gerlbTzlRryw1L0qW2EXXqK04Qn/ofzVYLcGplDDS+GTZvwTsWEP9VvyJK/KNN6RVmhz
+MkpePDCiH82E4WtafA6JRNk0D5ozpaB3gU8E8sfIUGBBZc6QoR9xbvO55XPbiIE+X9CQtPMB4Dn
pLcNt4x2QdnjmjO1AHJ7kzenWVFmhNHHrjH4dGH30C5isH/236eP7xMDHboiti69q7N4U+4q+D9K
MtBx4+zueKhGfcN73gyTgVNaOi6h9SxOMnXjwbkbj81IeKKarzEkUkNUX1liScHfHwoGQfZPRfk/
sFEYx9mPK5Wr0g7mzBq0EXyIvF0gZNg95fhyQpGeJ95uFwVtadXDUR43/pEZ1Q8lvfDGWP08r31z
sibaUNdiUxQYv/534N81cUUOxpRCX0M4168JWlP1Cj5kvAnKoBhlIkQom/of+jzeNfq4lKOmw8KL
ACEW/TzmXRd20zRkbB1kR7ty8CPTeUsYv45/MiPclfClGVm6gdmxvbVTVy+Fkp+7WlTFX9g/cZCb
Dfj78HLbekBUvHfD8cq7uN6hL5orqrwQZ9kruCZzmhslsIj6iY9WfMEnyoNfUJPeM3iKTfan4zaL
gcefxmZ+gbcXhkdcFfvt7ukLJlPe/5kW9Xuc8FEUtNOt/R5Jm0TNyuvq0zHBFQDGAh0BcSYImRrq
QXoZSKI31JpkH9apNHHXVUD/QViNBOfe54IGvWzs6/bNHCIXO/68DULJtXjbUWxaY/sbvVx+/C69
0m/fooPd1n42jiQyQubAQuas8CjK4pYiHv6033ZM4MiSjhYARnDsVYOBW4zpGoEFwACzqYzh1UiR
Zg5OA1a543WSwPyRjme5TDEAOvE8ZwSmRPOiIfEw49bi0H2T7HLkKMakHJYRHI6uUIMSnF80vgrt
YQLEUUtpG6N5VDbXpPZmz1XARC4HWQz4CIcmxeASX/d/cFf4VC/BJlOUEfimvvRKiDkG8sRFJpSh
pXoLVrrg5URqvLb+x+J5OsQaB2TW78bm6o4DleXHUpR3nQ3vsmD2OAVni/JyryGJtw0drGQtjX5J
BABsYue2/xd/N+RHIRyvMG9FF/gaIAtXyfsabxdqV2ZOMIoRyAmL0IxNHoCsPOLHXokMW5015Rm9
KEmDUp0PBViBuFFF3nArQsL/KJgnwpAmmzlwmKeKdvY0by/iG+FS8gRppRtC+8mDvdx+JldLIa68
9QiBLT6EZy78RYrl6be2WvttYBbTHkWhwx3mB4U9qh9+lU/i3noImRFl5ImMouWYiRgvP1F1DZ1X
mmJY2wgAVvuiIUwdKlGPHl1fCLq6XNjDQQiCbWxH52jCwqTrB4/FchP68kVucvODInuA6btSalQM
DOE7Jbx281S9c33q8LhcvZWAtmt4p+kPI03/ETlxnB8UwyIQvJbcbrEt2g7lnFgg40+gWYQEhLSN
7p35yLwseZVroJg3s7skTEMEarywXGzoHC/LwbtG7awit2HsFZRxuwRw8I+di+OI9oQ9hpXVEIKx
wLGpeQqLPud9R9cM3XMJXZi5Fj8e2Yq6E33UhzlG9ScTtY4WZmN+QOm0Sr0Zz90JRCkWQcUXkcWN
e+5ad3m3uEhXo7a3vRHgzXa1ubFj/m6YwqcS5as7jQK8iG1WOpS2rV1GE+BXKx/tW00OtRHt2PTM
TIx2R3woaGDjJqPo7trKSJJUUaN/55PITwjuh/kfFY4WwB1GBB26Y8P3uEl5/1bvdpE1ZzcT3Tiz
+Nw9pmJPv5hROoEAjkRjIQzBvA5HOP9IQcb8ILAMoa7JjoG/bRMKiL1ddB6Tii5eaGs7eEZPf66a
VlehX0BA7pn34RsFD3AFdb4nAvASJY0SDfzgeRontdAaWj5OzxXY0KflPNeknmBukc62b4sVZbP1
sonKfxKSRaXBV7l+ca0yhso/zsSp11SOM9itjK6US0/fOgj3PfAtcvVyxcBuC4lSqX23jHajfnd+
C5Ekg3nfHx2Z4On3TMf+c3JjVGiOGbR8SNm5oYENky3eRVf2wNkkd49C9ZSRKcEHDzHjqL/UaTKM
P2N06MXbecqEz4qRwdWuXAf1s7h7U5PtoRKI3mWRcPAlnPnvinr801nzr1F2Eg70icH8UcSgIXtV
6/1/24DCx6uVP4Cps55hMBnp5K6i5nmQLPq0GdMhv9+aB+vnJlaVB242mobkv9Q32gLEE2SP+GfS
QnDK69ryV0xhrsTIomLlLZ663b9Q63CdH/1DE5QCXv5kvx1mKy4Xe4Atfod1Ul93ZvCuGylsoK1t
G/2dGVY1vrB1FTJkS8hiaqhMickn0CNvUaDafKrjGs9pDVEMvd70CYUkXwGksjGusKKMSV0dFLDu
iBBjG8xZU6u8AtHG5TmNnFEDLbaPYOr24vnOp8cXjhzWQS7oe859b4QMeIjAMPm49+uHiUMcRQap
6u39swMiK2H15YuhjkBCa/rQ7tvGZwMnM3Hccj7pberYni6DVeikMZtYrc8BdpKsuw4GDXsKQv0X
nJfvsvgSMJ/j5R09xj1WtpLhtMiQG2/WF7kZ0eoFubkLMPUma4PUmibdkuYLmB93MmHl564Y+mMl
wl1tRkoCDvtBJGSN+EvsuX4nQDF4YraTC78h72WREzPBWYvCBvaPYfS1Mbw3Xq/eXEKQ2K6DBb79
kNcuyqeORyIDAC86Tb55doa3r8ukwOADsHvFvdnzqQ6pFAkdX/r7cgv+SKC5UYnEgKxNEg2mnL4B
ekoz9S97Lu4wv5mycEOxq0aqEtR9UbliGS1A7VuGSDYdVorvuK6QAMRVV9Tg9gLs5Tcm8rtTsN7W
QjdKYbm0KC2NdGKEAZlsdUMyQxc1YGDy8Nq6M4tUaBjjgyla0Y6UnXBIN2FXnluyvt3H2688UFbH
nXRlDQAtt7Gfiwo1yrqrpu6ED74pewUSSGeqNqZOm1dqov9AasYSHc6FooO06GKVMBoLDzN8Odw+
cD2YJyVxum5U0A2o0c69vbwuNjvQwA25mOPiRs1exqD8HVxzxSQ+xrbU8teCqkVTm4F1ddTIgWSg
DrfhkqyvyUc+sFn/nnrk0t4OlCCeX/qQ/3r+ey81QLRDoRmtJo5U+Cdj08XJn/kGkQZKLWsOjjVL
w6tqYKcnXcMjDkwrmfx4eHlRzizSQejovGBw6xMqnEfckKhiMZFQVcpuACXsLS3wR53VSniUxxIi
pVYBpQvtGlt5Vzk3kzT4H96kS1rc+uVpLo7tLrX8OneQXOriNC08b4UnRd/8Uet1him00xGcWPko
d1evhPfqzvJM5sEFnGah9VNN5xqUshK0Z7hqlLNoaW69in6Do3Fj0xNEIm0JxwTlwVg/izUou/KN
2JwKjO2IHsJJk+dBxELOiW+k1Zzji6mRQN0PwOLeOAxQjn11+s1PWGVGjdRfPldHMR+k75aMIfIA
sI1K5LFNVqXziHGpqBoy/qAA9PObli84ZVDtwfj5UOMywUcEIFWTqXSq/98yY9H66giIy1T4/PIR
+ob/w3K+u4rkFxEI8pNYJEXfn9KJwK5+WXyOdBpUFmLsGqIH4KODCFj57DZuqbiCnUeLLi/OYmB9
KL1nUqoOTGsEIwO3LjecBaoG2g2Akb/Nw1I1BDLNCEQbg35y8SJKYjI2CS6zLu+iIPq8u2ppiduX
Azsu7k/6q8nKf/k2iP8QhvRFprAtTArwQvA/EE5Bfw4cch0rPLAkMBBLdBst3V1Joqxi82qofxcP
A7nvEJvn06NVi0aSP+wM+lHT/XfL3XB0WPkEOysNQNRIv1sT4Wpkl9U6h2waMzDEKuyNXXGLqNI4
4E/2K3kizxAAFN+JRhBl8Bi0D4S+ocAhkXwAhQcsKm+hd9/fVNQDnA+OZ5nWrF05LQ/hkDQ7cM5o
oZ1mTTjvmxhVxKsEWQC6PmgdAN5Fs/rHLm2hWMO6HhEytVYdxIelRiCw51G7QESdLJVQxzttZ+hY
Y65icUaHy6s/i7c5BZ3YR6WnZUvrZ7blHHNMcuqjlRtX6Tm+W/qpCexMiBFjwQkGnMwz0Cb6RzXE
+mGVY/NrTrpL6/VF2r+KltiXfXRTiitJl70uIELVLm1QHPt7ZKWXeZ1DKKH10MYHdvlH1HxSp8oo
Kw+XBuZTKtsXXW9JJ4wofBQo01gkAu+C156Sg6S9lAZRqAh62CW3AOCm/IMpW+1+1Ev2nB9vNCu1
iUtdQgFZjua0/X6Dq/aCmsZdZ/GVuIqXi9YeasI5/dv7jq4Gzsi+6/FNjQ0oXieIpBuOibimfpZX
ro0OPeJShyQA+PDoVRCQRRksPgWvJeSKsCnmEfo/F3jNXP39tBt2m9zkmfjbCAjqnFDe0aAyBWFy
iuuoZBMSQ8CkgLzz0kExIXlGp3MAaz2fHPpaKLuol8bEa4HD3ZYTobXeufKmC8jZgpwlq9DpPOYB
80JJOnnjcqzIOSuLSSZlk46PFcfcupmbvwcsjk4smNbEPkFQ/GpD38tOnOXHEWtZQUuShrkjGvCO
F5WEDYlCS1oBU3kEJls3ZkfeiM7UJoNGy6jnbXbdkC6J3yMH2/3JYBijM0eI+yEFzyz7Wa9VptxR
nCV6gJ++/ljgEb59ShzWvwdeYxmUvj3CAXyircP3aFtEsvEY/X/Zdw3bogeOR5cVR6xbRLMZa7tg
iMVlarEDDlFjGDT0Pf2G1iUvLdkxwVzoE/PKqMF9NJKJ73sCw/SxGj5re0ragHBfT6blDuCiOCd2
6xt3Qzm6BI+KZqbk5X4bkjXPZ5SDak5XlEDT+2neuF96wbcjwuKdSpza7mM6otIXnqpY+ODxlOcl
VdwMyx56Yt0JyLMIpZKXwkfzYuwTjG1ApiPslAo0AeMrGqPt+weBvdguSPwBz9QWls7WtlG0Ugil
6RGdoB7K/zsAeiZK5t5XSn0JrLO/18sxi0SAmOxs0RiNVjqPHnQBoaWd4kU7BvuJt1Z573KfWgQS
7AYmoAb9eLU+31C907r2+49YOIxggi7VWHeS3VY21Sgjl6h/XC1JNQUPfF/g1aLrn858XpaWb7T9
YyHBWU9FOxEOSMGk4tdhvKlFwwL6xoiCIi1+SwUNFgU3QQSL9+ygW/eHJoiubUCjrmeyPeeAKvS/
UrWOpaA92uEmlgRp42UFjuT1PNnMQqACwbIEArK75CqgUw5TJ+lffPuxVM03sVQ2V9vY2gJZSNTy
jeAnJ+F7J2OEfkD370PwT9SnRTK8E0WURyWQoCOYCiULiiO13jMVRFYv/pYTPE9pjzS1kVkKeStB
ObtyYlSUqaSPowmzLZq3RuAlDj1weD0MusrFDxQkC2SdmNTQ/IDdxEn0jhx0U6nELIA9vLNzD+b0
j7Ja/xBNrCWr0htQo4rVg0DX0IRDUjhEVzQnQzepSXgdrprXoU3BsvAziVS551IKAx12F4lcoEwf
CMWbxs7EFO5iG6RNr3PUMqd3Xm6fXs8kh++PdyvZNGrjsk8o0LTFt2RuLTxVymh2lAboqMgbbsVv
eY+zCWA6Unzn63K818vp24zUllIygc3sqhMfj1vYEb9T76CmH4zlHRG7O29jh+mTT5qK3KIhWN9P
PcUFUouAZverV9lNTi8zdndRdkzubJRmjUsqwmRaNqu/g4n2xXkK8fK6upZQAKTYHyvCSlODKrzj
5lEMfIVHK0jJDST5ZJAfgFyB+V1oXRiZ6U7hLX00yYc5ORqACtoiAhD4OXtvZmtg6WzZ+y4+/G79
zgB0RsHEbRPFJvoKajS2nC2x7UNYWLWm3VfTrSTTokb8keZFkPYDrhplQ0qkXedKmZGaF4FathgJ
gtOvXEfiG/l+JzC1A1AyV5iZDBHgamI8Om5K0b/R/ZcKM1sZaUjEb6/xNyOgXcYls2Lls1h5hWTN
0KGmq0OwDPR6pShHj0Qdeo5alj8kHT7hJUSA4y3xQpbfeTmS/J0tz+cuS36D+86Ih1KwWkFCxSMW
LfBPl8xJj9s65fc4bqj9Oq1Stu3VZRAikF425qkDWqqkAqETtx2Zb+Hhwa+ssOE6xhp6N/L34w4R
SIygrH/XtMsC28GI1r1/BhXDN19fGJgiA8nS9fKB955ake1wyoFVOCzslyETfWckhENo1b67DCH0
mRyF4BkWp900ZTxvlFOVuQrK6RDs8t4VCx+Kbd4fHAs1UiPv7GdTB1+qiIdIFt+x7AS0pNKEBDwm
SbD+3m5L5R9TYA6afGpe6VZrkHVj+26xCYQPzzVmlwB4shtCcDRpwV40IOM6tg1fjoJyZ40xaMj2
+S0M3WzVTmZXT8qxSB0Hzu7a1c9sDIjFloEXEWPALJpNH9BnXOHc5l1pHphQx97HMpCf/DiIuoLl
QFSPZ1U690EQTDbB7LYc6JngCrIA0dIPLjYh+J1ZDOmd89L/8tEIv3Z41FefAR6NsvBhq1L9P0TF
OLPMWenvcFdai/9L6qJzKrPqprB52T5oG/pq48kRdmw0m91SdtGAUpGPvKZxa6huY6C8+7F+Lphf
Cm02oZGn2qExDGTMjAB0WzwZ5nm4ZxB8qSUbtkjQgGkrqjkMKZe7CQLeq9qLNdzXHzxOq589Vr6m
ZRh5NtYsfrmrkDjaQiFPangJLYny2Uh4fLKNqU+mCJNwiqt9ryOde5YoAO9UaEzrhbIdcj007isF
iU9TBRpngZZV/usGtE/K/jM0UtgWpX7IyXyS7Cv0E6dcMRiMf5LfiTcp0zCCxpJ1Fe2iIPoyQwP9
sifasvRqAA8e+osKEHnuMxBGfUxH8kAHEf1a2Q6S2qyS80ThOis31g9u4LiBE76RBsCupZJo8jPg
wc9PXwjBtj0LnQ03u+9yMg47AsKR3W2DQiRu78nYia+k1P6vorrNqXHjA22gUPsOmBIVH+jimUzC
ZpsRL+xGm4eX3G6P5yHy/CVnyaJ9AOxtQNRHJVAorSvK0BvSd9bJp6krkbGPEwgXehgW3VUXvs3S
7xxoR1bxug1omn90DTypZYcXdkVi56kAALJ1pdf7vV3vnKnRcibCF10J81MY773z4l135mTZLecz
1gUu1QtrHPyMkjRpibcC7JoHUSxSrmV90p0jJratCEEDbC0lNOEI2StGfJ8CeBXYjqsZjr2wKlik
N4LLT+LySkLUYhQCtJRJ4addoQL9hCaAP+dbg6S+alanVgxjR/vj/JmY2NwmRGl8zMi1mMaUSfad
hcE4bqmFHJvY/E1SS8iG3kuuxnv50GLgD7gbQjze+nPDzx0QrBoP5RgJPPfLNNXYtN5Ok4tpaicY
TyBof/xbYkCPp8pxeUga34QxZSLFGfGRiSeWMLGc5BH0PwdIRnhk4a+qmBVa0I/56lTpBvzHl1Ws
YqKeulqVuL5xS4UxpqKI+n0S6sPrwSkBMyJtn+PfxjuoDiimtuLatQFWqY5X49NQ5q3zn6bin4WT
WT+Klaq5ulxbGFkm2pcpzSVmZhZ2b06pC7S4gp4hmmX1y3y/20Jy+kNUv984zAL7UAVWFAhuGFX2
blS4gNppi9W1TRPDhmKtHOl5ARQGCfQDdDRGMTMfEHTHsIEZBw8CeAP7TUxii1n3m2rDTK2ae2ew
LJhc+1zHff2PaXDecEij7ScxNuIsdwQ2UIN/FvBvRfR1PT8MeuY6R/J3xcR8sp3s32+zUZlkYZl4
mE//aj2wkvpePGyt5rHSacPmWMTnSE2ire79CS2hbRmP5B7wkxjrhURx71nJ6P758OZG1vW3iUwy
Sk8vDBqzUJlVzkOkgcwt6G6mezqSZOB5JpLw2jOjkVqnT3OjvtyhdHcpHs16CVSYD/mps1rzxmev
aljS+ePz5WyUAMkFwh05TZIWbuCxWR7Vi5zHYr8uhDL2s0IQBIY1BZmuWmQVm/g5ho+OQR4uTmN5
SWGg8qu3XIKJNrPC0vcx4Ry4zHFv4PM1tRKp6/qEOp7tpAofRAP5hiWW3Oc3R8mNBPJYF7O4I369
9EDcLWZpqKitSBvEOSeNxWQk35LIqusHj+618ciiznsbGbvBrwhHXWDZLMTKorP/VjKA46TpTpty
ZBN0yG/iRlsv9DmjCaMv2U6HcYegJ529Y8hGACE2eDTKi1kf8Te0Ll2E8/slGi5v13TKjMIt5zYj
nsVcQQNNgOInIoKgYsu4OYh/EE4E0vEJsLu0utK5v06Mrp4F8JNTXTe+6MJYKkNKqIk+BbBaMD9j
MBFlIZr6sT33WgjqW5EvETUzrGGnTYHka6XsfZzIfH1jFs3oJuuwm+TaE109GL5OTUYGY0HtRW2n
AKJeRX0mGC+lQN0tiz2ciQTSR0ErhjEkUrpvhCAMFwlusmeB4AZ5LDQfw9yPnRMdVYNI+Yh3bSPj
vvO4nIkHO6gt92A9Ahn8qceUI9iNqT22GppR2Z6hYxA+DV8Q7ct4w+CNtmej6GkgFrper7WX+eYd
JEyrOZaLJS804FMKRLZHOKndJVVbJcboCruQ/gU1mJWyWGiWMzcwGHIbw34zm8Oqa9z8XzCcdOSb
gJ/XZZA5NJf/wVe4ge+xywhx8xjVudyM104LRDIrJ+tf9Qbr6epRztdglrgkJLxDStu+fQwVyv5L
9JxHt61wA11sxiVnmnEDesev5jpaEHVEbniIIhcbneZF5XiuOJP6jx95wMEMjD9kJZhU+k+h6uNg
pVm6wRGhZdC05PG9gYpepJAZ23dbfDTmOtk/Z006W9WLW9s78bNnL8YiEdBmKNweVLSXHerSzXtU
vi5io2cwsfZ+GUcLTMlF1lLLAW8goQ165dhV4wHSMcdvMTs6563IG5Khh2/pXYt4LkZtuxSQLYsX
NNYc4aN2x45PT/mB9SGHmPiFJdwbbpQxRHWFW64b5EYExvf115zipqCMbOj7aZau6UqUfo/Thth1
f8f5FGFgETUesF14GwX8NL4hHVHwnX3LpeUpmy+KYSH6ljrtq5pNqGeQgtBXWV5WjwTin2cZln6y
V8oivzNIlK+OIoybI4j449zGDakE6ob2zd+UckCzYrhxuvCtxtG1RT6sfRh1wm5yW8wcGCpk5LUz
01sXPjAf3RXQfi1jR/RoK+1oMFtaT3DWVqhI8rjtc1vP93dF/xEYLCZQs9qxRLlv1n4arPDWN+aD
LEJx53QcMdSttHK1s1KFX2nH4pHLZDIs62t7/MkzvIGpuEU9rc12d6uV6XbER83/Mmy4XsRcC/76
YldcNiO5ecDUfscxQxkt0ILpLolKQzgLagwYq38GcI8+E7L5AeYGrkULJqx3QfuX0ArUm1qbJicq
yCpiF1KnMPtuXM07ICpcgk14VgbH4oIQftPLONreJSWPqpNg1fLK6BBrq6LDWTpoXwX7HWlYdFjY
ujMkl11/BVA58bgivwxE2QGlAy8sfFocBRJdFvYk1AcOYIhb1U6cloFTmwxvTV4Lm7Gg9tg62IfW
yMBBtLJfJDGKpztPjzFKC/ZGRCQ7mAWLqlT+aCxr+f6p2SxRWrCokJo3woDiwgqWqFfoGPn3Cd7m
YDJwzfE5Oy5cAT3Q3GxMWUp/Hvl0QwgaVdWXn97pd1e+mdGSCVCr2Oh5nbrV9zoFzvX0WOCgELt4
bexQTwkNUeVdlH3UxyCdwc+AOmHHnDFDl1AFGmD/F+6JETxxbSSb2/8onQnCZMzcOXYDNE9RxHbU
85EUOioDVvGarQm5I9G1Er1qaWIx8AvTEsUvww55dG2NXgYGjuJ7axIdaBt1dn2tPogkTYB5W9LM
t9crZ5hvivz4rFxxFpyvkdps4kRS0e31TqSJOAq9amKgnlKLTWbyQ+5OeRBq/P8wccWNEwNn3U/Q
oCKa2Dbq8pPINUYP1QdyQK2owT2MkrcL6BxWnJmDcdeHYqwSBvdmAE/hye2wrSOeJBYeKTIT8y8I
pb94jx1pVibIZSwoQc1GQ55MLXAKHpYyVPtfyRkoAPZY61ccCKKpc3OaEkoQaLqkanzOEuu6R8Zs
LjcizE5bVO9m/GikLWFvVK3GqkFeRNj08HQxAP5lF+rMC02gMwvm85OJFlG4mSlN4mcP9ml7pUM7
IX64DqwHpsJ639qBXsVFj2LyYPIXTmIyAqk5qPxebvsrj2wMWqcWBdjaCOEv44j7s1aEwgbQfR1Z
MIX+7JL1YiXShMoJozUxXITNmZ6m8rBi/tEDyIaIRLneQJ2WcEeoppygu9UJgYq2Nbf/khKvdkOR
fwVq+ztU8Ly2Msb7P6S/xBTDowSI9px4DDWF1HrgB/lCtl3BwcYBtiWgT6ce0tnBMFhglYgPqOEQ
l4O8lv2sd+tpuQswG05QsB9AHgKu8PwPOGupWiKmTMe+qg5GWn6y/UpYebMT0cAhN+keE1IKxJQN
bihwkKKBInWuzILfCYJhLzkDlf4Lvt5ZJAin5KbrQxK5NdP3mGa4N77sxcFuKyPYbVPHRrjNVbTx
m4Vga3YyytMOoneQ4pnpB5E9JkQ+rSsY64abgHQlWJxhLSpS81yH2kVi/Vsa/DGx2kRB6QBelBDA
x1TPwBkySB1I2+NW1BcHgGxYcKJMwMvW/cRwVzWqdGHr4UvVYHVTjH/CRXb5JjdEsl5dRMYDU0rS
JL7dHb6Z6Mq/zou+6mJ6whjqL3cyPMH8apLlc/4u4WtT0dyCvjdjLgadrJySUPRBAyy1dme0DYmF
NasJBXD47ZXO4mPZhedl7Ziyouhl05rg1iZh6HsNRjmHk9NylaVRUfMRTyN5DYQNUx+Sp9OmTbM4
7Qte2cyNTPQB7b5OefrT+haFcfmG++HOTgtFxO+tRzipc7e7wo4fkjFX0sDaKsiFJXZXgu7HTo5A
k7OGeGWkVab2S/CADilNniEEsq51SncmcGozymdalSWhk2kNld9sy6HzF1CCs/v2a0HkBiOhMB0O
iZ5FDMYi0Fa6fkjkcavoM4MtW0GcpxfPWk7Q+PHC6BQ76E/U4EK20Eb/s0t0lrI9MMFulhx2D/KD
rGSn6qTVw4KRGoTbtjGiHtEkQ8d7nI3/sahec+TR7EHYhjf4J6uvtjIkU4EH3DGTPtpItLAVbCg4
+qOCSDvVg6WfkWEzamgKtS7ZEuJichF1Yz5gybkVG7GMmNVv6gLnSnb1T7shtllgmHvq4YqvW0Nf
3ox8e+35kP3uhGAOUcHyGHQYAITAC0C4es9ge4ODMl+FFkT0iZvmwm7zQg+9Uuckb7fhA7WhO84M
2bIUQ7u028PnEn8CIT3EWfs/ogPeHeXZ/2vDk/N7/zk+d+rrLJ4RBZl2/dmzM2w5Lu8HwGZNAC1R
T24rR1lV/Pppk5kDILT0Hi6MqJGdou7IBVi1dSQdO9Vku2DFjY67ItWKPAoM8tHoHk/MNX6qFby1
Nx49+aZenOhBLaVDtxmG2htPRLJQOoM8I1YkRUkjfu8YjVJhp7I5RIfjl5Meny0LK5PT16WtDN4e
jKNPs3Yx+gmvkfeeOGzkC9VH86f89cNOzyCq9mDBfeEXVYKx+ixdYBc4piVexZgbtUKKSSW/kICZ
GI5hyZ9iIEUTgYjPVugQJdkkPnCvT3lD82dDNnU0wv8HbMC2sl+TC12B3eTmRT8Mydff2n6i6jyA
0RNfaSwIo6iloGMmTyAS4ck4NTGZUQ8rrMDjfYh9AM5BctRQtPltaVM2Wh+fA0HGlJc5eChIi/z7
L5ajyf8ITBrJpZU/sYCDSBTNXx4dxSyEYEZsSSiFUpI2/I3XvRtbvwjTKDl9HDbaOVHwhWx0WCdJ
xLEnRDXZboJARKxQC5G5Ppw+xG+cFG6Vt29xksqq22istiaGJ+OB4oqbYxXepGh1J9GJr3w8CKAI
5Bpmd2E/TsanPsoRpmxifvH2uXB6n4nCpt4Cxa51F5h1tJv6FciISioYG9wTZlWbM8HsVldZeVL3
xzEy0Q8V4OBLMeLFYuy8IfNmzJ7GWGBjvPJhyzoCFvsu9IH7r8FmXXYlq/IBIp0ofr2VyULRmO4G
42HzK8ZylCiweSO14YsynSRW8tcWaKbLicmlxMEGaT2N95S/hPlIg84jORfEk3dlrr5p3JM09Yvr
NPzerrnVfLsD4ObE1GzyaAqfmC06aiBkl4CCF3tEqOT5Rrn8SuDFPC8BiB0S9THEmryhBreMcrNP
vrOBp/udG7fm8TUipkQJUIzJ1KsTlWTp7+WXRCLrz+Sq8+N9aoYiVVBjDHuPoj9Kh9UHT/EaZ0GQ
RiNQfJ27pAS80VE6hFO2qLFuOnYK2j2jSaXahmcripz14N3cwHAUwt/IoRX5F6hifx8f9fyv25XZ
O7eeRrtw3btSvtIpyX3DFBlldszfYvq+Jc2xrY5EgBnMLRAwah5ovGRiEGBKE80WppNv4zc7hSRb
04hDHyD0SpY1gi18nvLP6yxWHWFmzGv6Q0232qZioEHdp/hc2hVTLwRTAoKCXegBeAIOW/TAg4AL
aU+djF1FUHjPPRp55fBQ9doDhYilFVcE9ZZ3oI+TyYtVxhzn/QEv1hgDr0MmPzr4nazexGQvl7FC
SUtlpOIBEjaYrhUnPYIslv5CBN/GU7RZZAHhbsTYZp+0hG5l1B/gEIepf+qlmJqc9FgRxDMQDUlt
hQJScJG7D9ocvgxR3rwHZUQQ8Z6Md/A9hZFU8AiTZoFO5m99Hwc6QM3HqWg9f8MDH8pJdkpKuY3P
TYvBYI2GDTqj4sTGDDGY8JL04uayEs8dKjqehYEsoY7kqkpjrnhkY/6yfhnCAdA4FvN5VSN2ndWr
O/pCuu5nbgxzEbLIhiwydoNSnTt968mF3FlYIWGY1u+Fx6fLPvIPrACZOtV76pizR+6qzA1uZ0B4
8dg0cYl/ca9H+iZrmmLffqU7i8V0bGowmxAzN49dEHUWXU8zNoPs2xesTpk9ucEcWN/K5zIt7Gsr
1t0TJDQBsUTrANn1SCxEovEyyCPYkDv3XFZcU5HqynkkcoaUMGXlBLFJaJYjf2JEQOF7beW3ml7D
tud5YPOPIv6122ed/OglFhFHXzNb3DQ1SGuDSw79RkW6N0Ql3wrnyDk80G7nnlD+5UyY8/pbeSBJ
SpTxbJpFS2LiWJKZ+SGASnS9Q3SCTEGaiaPcnrAV3C9IDAn8dcAb4X/21UBSC59Rcoltva/MOum/
siCGHKm6pImIhcmHc8CItDOtxUEcLNJzSu7AlRmTAEtbd0wzxzKYy6QKEvLUAoOzg1uo83xfGl37
QOmTSMA3gjoh/C9h9Y1sOptNH7M5kLoGnfkRrCw2qaDE/zf/5vlegygX/kE6gnetoDBwiYQJ3FqR
9n19kY9We1LToVruO2V0Vq+qCUUvWytd9h6BR4gIjN4HJRShDq6upT4OV65nBLSMy8+KxlEbxs8g
k7GxDaNdoHAitMgdrPlsP/fcrs9fmVYpRiMFQhQpHvPi7k+r1R2BeqeCZqOfXf8CfmKJPEInrKHi
z/bMa56ZPbLaNhZhAoNlck5paU+ja2x9wuhL9XrN2Ngj8FdNPxAqgZEFvkGhB5aiBivo8lmasTO7
C82D43FmHEKeY6CTnUWaxargz4p8w8rnj4NlyYMI2JgFJkFGUiYdxTBNVODz/mBIOofDobNb50Ue
oVI6EDOD+kl21naHYkQ9l05GBxu8b3Fr3YvZxeIkF2Cut3qZudq/4Fshwdvtzg8KxFi5qFlLKe1G
mR4fzW3VW+gpD+We0MQ3rToQvLMLvw++vygtpqbm8F7rvvkoDRZvv29y+51qAvIoPg/kklSOR2US
bj3kMli2OFH2c+ralDV4CsjkanFJzO+rh/splgNd+yQ/przzFi7Y2K2jN0gWme25+KPo5uE1vfY2
+gQqUucTybIeE+Gv5n8rUgmSi7ZjTDb63QknvB4HJVa0s+dxQHr0zY/AmwSbNLJ/nTu00AFjPnRP
LcgIIWjF1l1bBH+9DgCMFBTbUwmeHo6mEufbP52lT/RTj5lK8PfjCEWWtuBCSdpeKeqPNH8nHOFV
7KPPwzgFa5k71Ljz07+M+dM5n4AKPbwiu6UvDhmeR3YjS3rcZ/BENK0iMFWe+TdOHToiTKGHRmj2
0zv+peeitmJ+bPW4cr32hsg4ET8suVpfthcG44IgpTU9rk7aosPd0WfDMbWLvy426QdWwDc52Mc5
WIqQeF6yV0QLkSCVZ6DW+G0WDpjuUQ/TrFJzeFCmTZDqGvQk/pr3VDSoAtTPqw7enO4VfFNfEvR1
J4fceQXuCpDmX6K4FmO9BVOgcjiwt289Q6fWIur5U61Tv+9vnBMHi5fAp51DkTo455Nvo/77A46S
Fpa3/+9NP4HM5+PMQ7IUoDvy3G9sGsvDY9AWExsfc4lZIF7GvqBBV6K771wHasc9Pr66LaDCVfc1
8pFvQ05PmYDjbJbEYt34n5SOB5KiBuKlvl6P4g1uUbfHCpezPzHyNzSjevOoPGB3agOwKq6BlF1y
mgHptVwlU0M5g3N1OaYgrZ8j0oJmEz9QpgZqxNht2xyG2HAdqr0K/KY6IFreIO8NnoDt74gXkFFd
l93jP9rh8Uk6ovBfFTpbuRWzYwWv8QLIrbOpE+qAZp26wYdMe/Kn736ylmqpCgxGZBGFiW6iVLL1
A5xWb1ORxGhlMgFfE2VByaNONShOOgQxgjHg7/5WWM2F1E/bidDlqpIA9igMXeCMMmNxFRNxx1Wz
K/lyGD3JdwehFZ58xxafqvNgDFQ9Pzh+4soDoKFERO5b3aPHswAzTzGL9FdvjRw07oZXo+b3tI9W
s9F1dnOxF4+nQROXRKkXgFfMjfLAcaJzRU4mtBNcAJjaM619QY4nwRQqNF8pxf8GNFRjMEbzy5Tm
/FAdCvSvEkX2FubI1S0Y9mrL2yBqDAvGs/Z7C62FO45rr2RY5kLd1jQSr6Z7S2e0ZvOtAgsjSGh1
1z4LSh4azzhP7UccoIZzyG0CB0fBDzf7mEX90XddeGvpN0xlazE4DjbuiODspBKZZ1fAYEUEj5nW
rWORGfTgl9wBsD8G83odUczqAiu9cnbdnSeCdICULIEURfJ8/95WfwgGhbOZFkPhdMEei2pyiKR6
qL9mSnyGx0z72b7iXVdaehIyjpjp82yeKTVumXrjw/I/ej112MAKXM2mAYQCzzlApQr/rUwnG8SU
/oIU5KCMIDpZgomXUkOJOdnUK2EdADeYTHWcFzmxvbywB0q3DYZHOzsD6iBYlUnLxoF+TVOFH0cw
qrvETDtS3HxQvmLNHLNrTcROgMnMvC7mc6ExjxqTfE5wM4sYey5BKB3d+Gih7b6NnhrZLFOUTbJO
B/5rGL35O4EuCd8EAtS28RMnJqWXb3Tqnz2m2oF3AyaQfohYBiOWvCfNs6Mf0QZtYlAJujWLdvj8
D7yXSLsQrEWdoqcKh/zOQkc9niDCIQgm0zZh4gTe3vxz8uG7FNCixrDQgJKjXNjXFhshX6gCsnJ3
IN1bUkPS8LovN1brCy2Gcv4dEwe0/ICFXkH8zK3MOi4W+0W7YcYFfXyK+QyEeIEOitptVXZK/Cko
5WslLxFpPlXkLY8JkOQaKx/KVzFVCFA8hY16+FmCfVfNEUKTr2gVd6UzvNO36fA43j+JqSV45DEl
pE8pNGyqf3a4sNXPS4k6gkxu1KHvjuUqZGO0dGIONpLqrj89ehXKHGJLNh/QtlSkD4rBP57R6U9O
NdpoctnM9rzgQS0GgtOCOoR8E9m//SmQKEUXF2GzZ4hTiGcqnv0o8J9Wvk7tfxiJZhdifwsVOP4T
QLPdpMxUM3DZ3QZ4lNELsnEJ/X4CjeSham0MuAL8wrvPbbDEPJhedBx0LdfSU3yOwi2HDCJISjJs
JSjtruWjspDTemDsU1lUsp+Qxnp4rVEd2T6zyKuHER9/hrY8Agg84FVOIQCTIJkwkj1iRIzhp67U
rgjz9hAy4jJtseI93bPuOG+WN1kGlf3NObuJR4L09yRteID+N70hDO0oAixkYBebQiwVuK5fS1Ah
6B6rEgktOu58WZ+vA7JRa94VUQL36ohwXWPHafCEKA3qWoWb6p3ia8oSrY93DfBfa2lV4KbpsYpI
JjkQNFTY9W2aJYv3D2//q7XMJ7FOLNY4oamYZstJwUJyZBCxZ+eLEw+UojVM93xa0IiZPsva7hsy
2pWQ9vUIs4kwaI2OxVOVviZTLzDEXpDjuWQ5bbZXHWUCohz44aBBB95/u9Gowi4saj9TOHFTyN45
+gzex83zWgP1JkpKGtZMytIE+4/IdQu1xplLjSSzT4/bJm9FOoHpf92frkhbhWQW6ZDFHGFHm4dI
86wuth+Bbd/mfIJRtXAiRiad1pdasdM1orKmDnUqfkBsfIXkh++pAVseWzBV9ymgnNRfET0vUpAW
s9wvtljlwyBhCCkXeL4qsG4p/iEogR7Gnz/m0jf5ryqrMLGR6Jzq+BjhEJM3zCeyooedixPaIFbB
kkxoeVgCf8mklmVkkV/Z5TSsErKr/uObIoO+kV7BMpvL9OGZTFH1GNv+BX1QvbpSj+vp23cSHtsH
pRcta7cvygc4KxtvX9IFLPiHF4MDu1hAuw0MfiufyQ2Dn5atDqgEhmtRbLpGbpZvPbjQ+n0CfdfS
mLjhdnmuzZv5E/AMzcEn8WOSf4t+rkWG9byiqGfZ7MI61sKhQz00bchy706AwvAH9t01nxkbon9s
wtOAkwYsk/eF/43/LgFAlXQlP3Sf7ceBAU2v/Jsn88vrIEYHRTFDQ4jMPRei2+ktr7ykBooxRKnK
Up+hckaIXYrqrLr6iYoQx+BOMmB5ZBJbS26lk54xEb3ZVNDOPdZNI/by87KzM6MNufR5wvIqxmWx
lzSnZoTiPqe0OkFXZo5yR3kFqY8jVdvgF6ogOvTpbLybCy+ahpSQC6osOBTgNl9mKmdyW6uZIy+e
SQFdJpcKrutc1LVbDG1uhdhoTmGgEiKGClx6hj28XmOapTfHSa0I7uLwjw1vvM1TYjBc35zFZuMb
mQIw3fhzo1WxLzxpHXd9vR8yehg6Azk7LcYmHwLLOBJOEhZpJx13jiOg1wOVWB5+kJ04P6ZCTVfE
dm56aEh+n3KII5Q5uIvOKugIfXaQxrY/qf3WnFOxCaLKF+OTEXzg2Mr8EaUzOJJd9gY4upG8xzMS
j5uBsbPWGhxih/i4QfqxmL4Y3PwJgZ/vBpq9MTXhYNTtg9pSFrvXEBfzcgPzc+WW9auiGNkwhGNJ
UivtZYJiQp3KjoiBCrf+NkmcA3iwSq395fGpzn5N6Hlp7ZhXv3WOj6MUHdJHzIzjSJebLyUgPbO/
gc5LvdelPHoKoHYi8GFJRPfC62LwxChnO1KIZD/fwSRpJgEWAXKGyfeRPwH1jYOqTYuwau0NNvOB
bHhcD7xIQWnL50iDRSn/PyS6+boMzy5RFCf4djC0h54hffZWfd4KpSdOlgFEgAUbj66duhbWCJC8
3wVQ5G470A+5DVpn04DdwKL/WFchlBBgEHib+JPa4V8vhV7kteh5sArghq0zUTMFCn9wHuaXCRTq
tpSsqDefTnn8d0szaKp+s9AW9qEuZ4I27DzK0Dw7Z2eLsW+1q6/qwGsYYTD1ZpDEiAm6BwuG7dZd
JcY6oD4qFMMYZ6qcUlmKoOFNtO51v2Vplx7mS73K+gZCyeVTccdHmQ3dZXQDmSLUunvWxvs/FTMZ
U4UOrB8TIOPK6XO/HCkUhSjWwgtDNdapPYXyyrCeY/YiA91gsBgiYoxR6VJYQ6/nPWSWAFBnUjAb
apKOHc4QaAQYdnFDaVIUNgbCSrHUqO2pdkOGx0fnfVbUwcf1jA3Vc7UTVBSjgpgR60Of+Py+q5DZ
Xt6J1k4d7SbGtZUmChgyAwIZjttMMXdKsO+t6+KJtAzwLK7imNZ/tNwX3wkIaZQ/4WQRZMi4/060
bvel3icpyrGp5+BBPfpoY/Tsa5Sc6OOI9PJao8aQHln2sHoc7XrjU8RdF5O2ChaxQVmSlUUubKCR
vNDHwX8EzoUL+uTAIhAZiCnm3kByAk8uh63jY4gSKLnEH2Ip/9lD/KSbnaiVItaxG9QCRv7h4vPu
MfE0SW6QLZ0W2U7jBAYGfowqjgyjSv6/jy3xg8iWUbV722FBdFE+V2da3aNMLXgaaQ81QUPopwGK
NrCGvFEgArqtaDT7UuPe+hDM8gWX7DKB6+o/eGBpuSBAkej2NSO+ns2JBGWZ/dwLeI1hIDWvJB3R
ljBSjzt3BLy+VxPz2A4VasQMO0DCNMljnx6VuKSx0jb82aucJcALZAzZ5/PAjeG0QfEEWoAPBt87
ksmEQfdJMie8IB6F5CPSE3oD+Ohc1OlFj2i/XbX8083uCTa9v4pa45Pft7sHQmENDVydfGaW+Mh3
nqBNH2L/0jPwd78qQUOdyHgc+86xnI0forVv5QynSDkzAf+/kmOGpKjqs9+YCaG7yVA/Q7k4rDXy
XncCW2d+BUD987xGNUiIOtgQOPs8cjqxJ708LigYHb0QscyRrlSzyrDp6U623pQN3gc4tFiaXiqE
emk7zwzScxlqXvTLDGbGKvjZ4aTUY2YZqyzvIoyJmsyLWYaT2LwHuh1ztj+rARZCprqo30k3Dm35
MRg3KSmW4HJE/WTaeE7tydz8VY0BLACBAI/3Dw0fT1IPe10iAKQ7rX8IH6mhxoNip0XS5bJyKqXf
bRL9Q4RoPMU7YVrKJcJZYXgoHOT122adieOwtAqIcaaAoYFFArOvsi6Qq8VDleTjyGras3UKQAY/
6yiaouDFhRz9XVCHBDg3Irp6YRb1k47UREi8N0+SNQLjo2d4q32fZpqpX42NCIz7VL7Zxcx9NQ1U
pV8dK+qsFefGU7UKTG6JFTCw7GWleuyDvLqhpERgm7xGHIA7BfReb/wQYDJZaCF5O9v9S8UrfmFm
NS5zcl4oERFQzvVU6Ryr6KmZrGPoX+xJfa5Phyu9qTE15+Hm0wh1zYGPFoKkkDVi9AVRdLYuEZT3
y5JFef25FwWMCKLrOP6v5ZeEh5PLKVwBL0FETjWS7QL23y/AbfjCfoHSTieOSYS+wOagTQYd1qjW
yoS5o6bG684WTKm4y4VTymzSQw7y8poNMgdfe6IePViLCRfLE3225z1Hv8rioeZcwWChdODRw5sb
ZERCntOFuXODOF/KkTE4axlBDqUq/dty4M+kYHocYel3G4VDg/JXsxuXOTHycHIjLFVVMu7EFcwq
SLFDcUVUF6/NAwYAJBmTo9oYc9oFWZwl2f6xy4xg9I1KHJaFoQfBYXDaYXqq+0w4AmXhY0rXsajq
ix3bW0jVOh/ruypp/Ygqf8dL51naRn+pPcdLtMYJZznIDFVrOmpyvrkctK2+J3YUba9kdnnkPLdd
TazMlzsToyLGIV9RgYHJi/glItVSq9Tf9iKaPVwFrKklZzUf7N+ZxMYVgJ8ceyxYFexxeSxXxOu6
1Gg/3heqzpl4Gw5QRqptzKuSLQOi6HXrHmIZ3smYxccpnryME/IeqVjQMY185lYZCekaTxq90Fwd
G1qtok2qzODIfcJkUDLUNb25ukaGFj9XBrcppnVHWvoUf6g6Uy6vdqIr8Bc+U96+5EEAB0ZgXDhY
uNvgIJWQ20MvFNKWlwVOcsYpDDz9LR7i1pfTI7RGslSigNqEP/rBHHWI4ZfcZi3kb1YWqETRyzt+
cqEia2rXPQ1mlPIbPtdXPToF41SDL9x5WkNMMShD55p8z7Ye7ZXUkM5wnobsepDU+kNh4w2kcDkQ
/WtSwsrl4KRIw1gQMKCVZnvK3ttL1tylrNEyt/cGsmzGcDVPile4ZwDNPPZK7EPDUzHHqnpvxRPm
4KbMUMqRrcF8XKMpVmO9DNnv3faNhYn5bsxDASJur9noMFh4zwF1TowkqZPyWunQ5UBbb9LAx+Rk
MpgJQVo+7yQ/p0UqZAROwSir5wccvK9ISOR3NJiEJlWYXlUtAoa4eRAfKf17qbpZ78Q7v89PvDET
udUI5snSMfdj24q1bUX5f5/VtEOoM5i3ojxRsU4gTlYXWanAru6bo6XAMpt1eTfty8RNvdxpR7Y1
23RQw7TvhHU/Y2gwM56vNgFuA5n+kAggf6j1TZljOfWNdhQfCACoZfGYt53DetuT2tnbDndzWpDG
Fu4i7b7177zxp06gzY7dGji+Y37mV4bbOcsXHIItrxnxnWtDOWPSbCihkSOun5wPaWpiut0M0fax
zo8KLzGesV0vP5wSmB/u4LUr+0DpJ99jbNUApQgFCAMZA6OUBA/DFb6R/forrYVJAsqxbZuo8R8U
IRvOsW2DLFxbQ9w3N96SdR43/xCTMRcRgJxTMZlqQvyzIJayJ8pHtqs8WozKtjCC+cKqz7TCsrEI
D8lriATGLxvPgTCEiPKKD8VB3DWzp3OrNBNbaAn497ZgKjpkW3O9QmkdEZckqIfAh5KdX8ulBreS
gNWqlpGYjV6tqgeVCK7gvh9vpg0pCqzjYoeaUt0llFPXjm+qMfhX+JNKUmbwd6CgOO/Xq/rUpbGB
YJEVWFlrK7RVE75ulDGC676WMJK2uNapwkReBYc7ZQYqpHfxnPcrGXR4Q8yCtBFS4xg42uH/hp3V
pjttXnH3ii2fhlpgi4cLk9aBoATjft7OtLlyFAGtV/9RrLgejE56WQnfdaTe42x1KCGHxpjL94fx
ZHkaf/G14eh2Fy+T+FFtHkVGMNWWMRagWXuLyu3tGpu2rMPt3G/iX6gfOnoCjSsFbmYSJk0KZs6+
ziQ5S7nwougm79VOOK8j+UQYQrfvORNs2OuwuANZnmmDUUx2GerqNboS/MsvOLo897SgPRQxp1Bi
lkW81UNIkVlX8so31TMqpLRBPfisKydVhtxkwp58VxyRC39CxpO6xLqABPvohwfCakO9YOXu/71B
AQp3An2HAyCBaK642LGfjvVk6AO1CVHgea+jBHrdMkyvpgr1+hja6BBd7icPGUResHXKFSBtqCTW
2Y2qcMlqo7IEmnMmCXar0yQZmqOAlowPoOwcq+i+gOhFkVzjIE4jQqkge3497qFhCq1CwjMSjjV7
oyowc4k772QENLktU/OwGr6ifDMuwLHSuI/ZAvy8b/WapWS7KAik8D33AD6Lbqquukq5x57Y/0cs
5aHudU9gGdwRBSFIn/wAX5x0azfUE3w49xyLbjWJzO8ilGI/10ae0nH+Fe6YHxKfKWCTxQTmYe7D
gsIyTV5VCZyZH42YhPWvdTlhclZe9FZnRwilfgLS0bhzrIYpFC352V2K2IBOpP25ubGtzc2PZe2x
J/USdCZsUPakebvPVBQvfoWvC1Mvgpi1nMMZXat4WzGy/7PZy/6c+koRZPtdzL+7q77+lYy3b1GQ
NP9LjD3DJaeG0yKzLHf1ebd2Sp9s8uPvGq2SfKxotUQFDrDISzSEKYYqrWgs/vgsKyvsbFn5J6fu
KEPfA1tFZxPlHvHUJcbUtYYSeEKUaY/kqWVqtfey9zjTNeA0uy4t68YTUKYqFIGZbwqbJ9ob+4H7
RGkDZIM164jNs19f5HNzZg8SH+zzXy4KWcGMrJLabB+oj3+HHicMu6XQk+7vwLxURWwnEHRe6tux
mCVZHBpj+F7MKIzDmtUhuUPhGM8xsXzeQDihkDizxpYe18XdAzjTEbskRuiGjFF2/dD5GGNsaoOs
KFyXk/HWyrbKi3SYH/e7H4qOuhRksPyKWlLayzbKyEKtaY5eIQ8rEzf9A+tivDkuhZDnj38Il47x
NwEF8Pe+Pb0ffFORM68FsWhO4CKTogQKVZ47HV8/C1c0rPwhHbM+GHc9IVk4aHBWF2evWqiUHUU4
w6aAUnxSvswFbPxJ+Ra0PGuASBOj08exuIjMrVh3duPEQfHUdn9ApicWy90v4wnny+NJumwgX6i8
OU3/V/J1VRAzPUoHPB8JPjeSoB34Cbc81ShbRdMEX9NQY8IiT02t0aeqvSer6DsoZePe5vUH+isz
bPDGhnOrhdruDYKxsYMuNN0v3S9U2KokS6U1YbgAdwMTB70+4lJdeiXM5yuCfasK9ISr7gqxCu+e
7oj8fKNq7/JFO0gHokASWPTn2tvm6vkAkQJdPMKC9rViS+2o/o9+YbSS0UZW0Sqs4x0bLaAPLInR
Tx/AhTCbK237IZRHFRsD7TUlF1ZAjXJr7Nkg1uefpl5BMxFs/YtBuPQjAgf8sV4JpLuaarCQ9j+u
7xwz7f4TuocvHE3ls2oni9QMO895TvjrRUOdguEs2XlCf/ci/O4SO5gLB0EL3wWgSc7Fkh3cknzh
jFZ+PkrnSznOKWEBJfEdXtQjv8nck+M+R04ZO5t5bWKCegFJxEwvTE0QxPhns8LLvOJuoOvc8Zig
FZkqit51/DFReJNM8W7eFn1W2GlPA30hRAMNyuNotSosRy2Lym2hWXWTnvH6rBxfSF78J8weWi1q
Yk8b1Xy/ukPFGmlRt/kDqL9hY5qyWzD+gzV02qp0MGhOBYF1A0cTjbjkc0NU9KkYbaPgO19fDof2
ecQq17lhLhgKeIV1Wz9OjgsOr117fWxdhoDhSUrB/EeCnbzwb08iFhTQ4GkcJiUvGODaACczTjY7
2QjgyZcmKYUB4+e+fjcCdUFyDFNasfTwMuo/1aMsQlxvBdaDoq/Uuz9jnONyQStQyArk9w9Da+hs
kKTDtKjq4Ih9+CJfur7N2o3tW0eXNOTF20NoV1IEf3zPlGgibreIo8h1RAxgtFBg7J4EM4ISSIGl
SyWy7jeKocGdtd8x6PqfIlhqyqRYkUatJ6RrYyWYUJBGwkcZas4vEIpudblizMPpMIC78QnIUiRK
lFb1jPksXMgR7DvIlT9IheUNFxrt4lkCBFj6rPFeM4iaxraJ+tMOFvhCdWTiKl9AGp5MCJ6vcP0g
aEAk9dPlnHgkYDG9W2Di8ZOh6zNHJzGhXqfYiNsbWlma3hOOiZ1P3saUCAQzG6iFs7ceRbvh/00d
d3imv0xbRnA9lm4CDUzL5TNhhOhW+hPULBaHkEhK8+nxe4dqeLnO7BB6xza/Pg76J31QVbzBHDzM
uwyoSnu8pa+AyYu7w1c/duUhV0cGgNFQdSz0OgDwj5WTwebUnLONf2hjY6aYnbAdrt6SXQ8BjYaK
09hcifJ8vCkjbbmGT94stxpLCTBU2tcWdhRWfR0l7uL/TqujXKKW4I5YOTHUfDIvLoWov9ieLCf9
zTAFCwHHMaVRQzGz4ufecuCsHPAJjnWgnGsvdbOIl2dE4+GIX5IHTrbw0sMcQYnS/pKX3tKbsQNV
uRlxPMznoAwwX9jc/o+YOIda92/7PXgzx9TyxZPuYTgbrnioXe20lkUYJ/fpW7pqU7nsPWlMrMgw
PwEur6fEKKOZZJRIS3VJmVmNb69VQAt9wa3LHMsoxYM5FgOfXiyUEAzAPOeren1q4zGVgM/G5B71
6f30BPmXi/JZf6i/zqCrMf5XL1iYa/rZ+yZYuFizJ0fo+ewc1gpAKgPS1AJGkMIP9ZbOMCAVP2mt
qeKRdK293t6fX5x+Koa5JECdO95/6dm2X8z3F8G0NwR7LxlmUeTszVM3NBj27BLe8lxtaC5Re0Ep
89yqjLBRhNarAQMYSk5B8uzMh4FdvNVri87xN16Xw+q1eyt3gX9Io0V1kBrmM82ddvjNzR0YVnFe
zVdgqSguo3K2Cs5JCzmO9liYMdKT0XCc+Jffy/YEuFuoKoD8uyYk/E7WOUvs+iUgxPCop+jjAVas
dAiSBMtiAB8sqTITgrthp0qu6cIEDhKAkyDQmcB5FsNEL9kYMkl8KMzF3+fkFdgx1ObqaxesYYdf
Kh8nc4Su+TOOye9nOQnzh5hPQ9dxxMdh0BWelk2CnMWkHUVMJQRgbDrSGKSLYqbI9yvEGotBOJnz
Ln/B2DVP/nr49B5XTIe5sjBeC/Rah6h1DexWbF3tfmNjRm44snnY/Yhe3uanTVRRvqp/VCDAKbDx
Qpr4xviS5DDLUSeyqEiMCUUWyruyTs8zkFLXkkOAlT1jBzKH49AL5EfUvOvC7p6gWLF9rdaWzYXq
c9dRHtmljhieKrAQzbnotgr65PasToLjQcQz/ZQA6InpvKkFmhdc+mPQECQKo/kML1V/j7rHbjaq
F8W0eNrl5Xig3W1c/kkjvIbt6yMfNnQFgEibYWM4yvm0g19Enu612dQFC5lGXj9htHNrp0IYGwlK
qEXAsk4DqTTu25s30YS91bN+S/ynnz1t5Ue7kjJPuF5AUBjcsa+YT2noR8Q/j4XzStLxH+gsNA6v
yTVpc46Z0l7odCowyOcMoMdVS3RfL1oricdXCKpf8MWOqSeP5QDPEemiNg8KfMCAqTf6LXLAloHt
kXHtQFXu3R6iSbs7fUvrpVbj2I/1gWSsYUNrQHNrkcQEFR3TXyEpibw7nB5nXl1Hi4cwu9eeLFtO
o6wfHc75ge3OG+XhICcSBYWA/jliLpCwDjv0N9q1OMu5sVVyvX3nfus1nG0zgo37/BOKPIg+u6nd
se67zawSFmw1jgVAtQW+wKvDZdi0fvMKGE6kHYOqpoOim369+OIVzt06swaVy9amspCxDbwwLvj4
9JTRPIDet6tMfwiJfhX9rajSYDJWZA+CFbWZ6HA3zlNg8EMYYZu2GgEgbPbLHIl9T3hWixmfc2ht
s/hh1Hx0whaDIzkAuR20An/HpkVydYvXAKvyr4ur5X7SGKvtZcdvft6gs2mKbKb5EtN+kbM0q0sN
+oAwuO4fG2phv+rCSu3XX+PoxIKAFDcC5rHZvlBmHYwsQHNR0eVaBBq8VLclnXOsX3VpibuAcPRx
eBX0sSso7xhi6/1D+rN6iiKQBnI1XItd0s6ol52/wlaW89mUYSIk2iNVHmrHQ0qJ8BVrD35PpJWr
3laqF7JznnSTBqQDyLHJy0zj9OHR3xSOyPr9LBJoKFki+pD8OI7/NGUSjtUuOl1+gCHl7lFqpIsS
k3/RNmpDTg/Va+zZb7DbDEc8junE+IpLtzZdybZzYxw4o46lipBwOMCMvnb9WlBBqCHSXUAnhn0r
GPUSsNVlwZFQtVpEL9xlI2GsCCUaO/qUcBzfaFruY+PZ5wJeX7RJ0DRGENLMoD1mEx2WL9LUG82R
h5RJvRNGe1z47F5nlw4ua5KJkCkENO3k7+nM/Q+AWs+nCegN6TAv/fT2//M2UyAmPTDeCHshIqvb
C3xD6bjwCDwVaoHQJmO0tsUz+a5DdYJX3xifF9tLNNiC+OM/Jwu0NugpHTN3MoFNnnhy4sQC/wul
5fSrTdUCryx13XTXmYz3b37/QfCYc9/LSFEUBFp1eiSMDDxb9cJhEsfLK8Au1a6L8XM+3rDgX7xz
VRglyWfg7OnscTOrkqcPMMbz/G4zmi3w9RjVop7UwVJGPBmnP2IAaokqVh5jJkAHCkVL00WG1fdZ
406USVCaXYj/uWI/tKiH6pkw/oRdk64r4UOEcMsoISx4ljG7G+9HZGbwWrTk6t+kqs47yA2Fp6z+
vJSIG6ZWRdlj1ltAozCXlAGmu5kilKckbix05JY98RKHSuczBrWRe2YlSCioVkEwz1RSm6GEKkc0
gyFBlK/RK6uzhU68Z1+5uLyuzzC9i8cfd4a7/0g9ntxuVN14TPSkuAjsc2Utb13wpz+vbWD58ygC
13/SpyHVwQhkf1j9zddv98MBLKwveBDVGe0wrzfRfg4JZcFLsm5gQoq/QivYruk9DSl2rbP5YomU
afjUL4s96qqOYRDlC53g01iL3e88QSZOrIEMkbk6CP8KoVVHZ/sFATlwS12AB51sFMXbQIuJZsGl
01pKGV7IcyTD3Agm2/4LGXB+Q9gPLZj8qGoqpyADGatIPxNlVJ5wd3O9LbVniEMNdomPocu8MzdA
XJyiRkWNby5u3R5s3czcX0JUIAksoJExnhJ8tp2IUi+8+MRkIEuhIfThJb+5hNXXGYtvg+3S5oy5
PP3Q/U5DTLl9nzjKI0PBtMYrRrvUcMjt4YClitdTT/nyq+rks3Bk63ct/IwKcGdFn8xl+4V2zudl
elQmbX6pjAhKiSbPzaEXyQh7o7+1UtzBWIVGk8Ku++gvtPx2vwXYDZAMy6N7ABNWL70Mn7UvMhyy
8xhpFigA6i7HtABBg4uHkcpWw6GlHLNjIdIZdgvr4MSY/AWN4vp04NANpjJvkV0iYSqyGaWeQ0jr
5lZG5kvk+J4iugC2avZx4prGpbGznF8OXWmKWvNRg4gefgY0Q1fvdRrSuMZBgm6NG5mRznd6CsPq
lzk2DHdPS47XspJdzlSWGEkeYbVT2HiB49XctXzdHxxFojlDPBT9Khgzi1OO1/g/VXnGZXSlnx3b
JQ0P0RlRACTiFATXI+hcFzvY+DJR5ywfeB/+cnVhipEV5/H39eLVyj8NWvMTeCqxwPsORqQBLzpX
t7C1Xfhwa4qJTjrS/Z/o8xeqLN+QkUEWlJogLtlH+1deUFIU7QJmkjW66FSXzFv9K8GaOZ1ehDf4
lxqkXxFyOGHAbbvT8om6//LQtEfuzzAPHXRYuteKHlU32lMc9llj47THTGXSRJo0TXepVNpS2stC
w4oJQKpDAYwSsId8AB6aWrmGV4fPMmQ1CHwcCN8p+1XkrLfb+X3y1aAFkCYEivukb10qtavqYklP
85YP1k2LpYqFjF6h0s9L/Hc7SGVpzHdoVO3BxIRCJz+HHH7iZQN5SVoZZN++4kakaF+WqZ5KS+Nj
MsJ670X9BYmWxbf1HGbDBUVNulgdXRGW7F61wbPzEuLovF/C/5OzdEWYTFfQmdwMtluYpxHHCuI4
P7TVXWjb6/ZlGy2Zeh6uIJiR9RJ26c82bjIIYiHQRgVq2hosAErzVjGXHHXQMgyz7GWHtLpUxb6H
UM0tztVuYTs1yzQonXjNEvPITBV/+MYkTGxWIlbesATJD8si+OtCjD5jLCoxt9X/8NwhqCMB9Y3J
HRqV+FKB3eGv1CMD/vG9am75Eoy6EHJnEvVHE8awJTAZyHHboyM+q9iqBLsC1OW3J5NoL8hZGChU
/4kl01TqbLSS8+E9ctiF0dBYinXylDaf4vTM0/M5S/1upa66NHEUaNer2bmWRCGL+4pthMKgeKGk
ys9/B0ILYPvIdk3vIXsEBw/YUDTN6m3AEDMBDYV+1SXnWy7wdz1Z1Qrkyn8TEk4+E0pfmokMld7H
ClegVoWh8Md+DThzLP1AIxvLvy2nDMF0VDHzGRfdM1YaYQV229uccXwTDFozQkI/y8yZLzaPJn6Z
Muop1c0MEjdWojvBYrS1ORpNNBcXrCPlxYN6XivE3JoAFQUz7Gxs9y3V/VFuV4KQfwxGifkOXJpU
qTosflhQQZGnaFtNm9GDY+LbvbdZpuav66cCQGha9w7gx1khpb1d/Ke1+eLACnT5/m8ZFtibInq/
6qG7nwneTGBYC2isoJ/XIw6fxbE6QunWLzsnsnefJ9C0g26BDMlC2QYWFm5kqtZpKdlkZDac920f
SnachEIBrz6pmtT+raAwnNNAieYqbw+DzNMFRRASohhKuCrl6jSVj5oekcsMjmFUauWPqwhsXXVl
0JYjfm3ZSawhwZZCuJm7lkX4uhpmQ2NVCPyOPo8VLw2q+kmTGjjdqv52pXzys2wECpFQLmnNzCEj
kJpPN3/GPfyanz1UzxF0lbFMGXzeMShiirCZlS1disa7E+hURoXhO/22wCwzhUkmHyEjb/oER90B
cAks49jJdI8ByZls4jQJL7LIwAe+OV4HOytPTJigQh+podCbl0K/GfQu8S/a8VAMTe4g/GDpvzav
yiB1wc2sbx+slwdt0NMf47Xx5dWdLzieIthbTZiaxFxG/OEycicZf1gZTxk0++CvNTiFDZCKZtnG
VNzqVUaJ6DRUWNnNvMUjhVpYXSPkcNT3/M4/Y+2h4FAg05b40ES6HRTT1C0lJFu7tg2fJe6eMyWX
uWqIEImdIjO3zUDAfWHlOVGyAOgx+Bz33Vcx1XY1U/IvVIB4g64rnlRA3lTzpueBRanObzdBjaAP
z7YdeAU2P3RfBylBIDgxe1XxozjOLXFiqEpX794OF+QMnXvBHJHG4NQBypJoM3M8qZCf+369soST
QAJ4vpaA+wrFKY9YN1BePpjzsY8czJzNHnYfgPte6WqwN6oLDcKvaKxRSpHDlQh02WAIDCcrHAxb
PL9eBjroCg5FFx3g2QmdOdznqyP2ExqjpQWBttwJL5eK0GVkH/Pr4dZHHwbpF6LUpLV2/oZnBoES
dB2/jZvwc3WXSUyRjERGIyfed8Z0XbWPcm2TBIISYpPa3ciSQWXnOCrvBQoWV3EDEKNFwNTEJCJw
u8lSacCjGyJPYp62kzqBfqdEKR5UQPMODXVQd57Gg2eBT5X5MWnJZTrFIkyRKgi5Dw2s0THX9cUN
wavzxYNecFfXwKrUa2KvjE2t+W5OxsI3Qo5w7Ej5ZZXCu2kcHR0OzVspvDUY2jG6GPDIfOuR/cA/
lWCdpOnoqW7YmCcEPESPZzO8fLJnvoj+afGi1IyevGMApvsdCj/5IY0TOgN3qY0MoXcxFIZknsHD
1Rr/oK1go7TanDuWQtWfEvUH5Go4zP6YQqycSX/dk9MUO4Aq1X4joA2D4Qne+Q4SoUaFKYi9hFMq
FqSlMaSVBoY8msMFIOpfe0j41FLtBKohsMjI5MLvtQfNXF1/BPdLVJWH+WxkBZ1g3kgzr8/j+lRc
FAWpuJHduCVJc/5l5C3xgHpgcvbG2x9hQPzTEKRBY+8cYKaQC+nwgni+K0ir4VgMdPdU9nvVpAgo
tM2JGL/M7TqCSWxC1upPBGo31QCCkipZS2UO1+VmbQbvbg6Z780p2fhmnb0tBturXJyGzN7hc5HB
J3+ucRI6cDyHVROBVJHRpLQdEjQqDzpNODuVUfPMLipWF5XGAFOTXeo/d6b6exIcAEA+DmGM+Wvt
OiKH5ixrw+0qlbaiZCEQefxNTHxskKiyfzPYgNxDiKcDhHSN9Rd7Of29UkKnv673/h857BbhRSrS
gK8p1nohmsvFbjuOh6ZnWqKYoTPPsM7A2PMz7lhANjNJN5rRzeZcfCQY/L4yzTeruiN3BAWJeXIu
AXK6Uev5vDcHQfcOAynXxO4XYrLLsivIe5i5IcOo13dzpbN9We0UXsCp0RSnpceirB3mPnXQHR6B
Kt6cS187H3tG/IC3zQ29hAxBNN3PByd+hPQs76onw2HABVCALy55Axv+dVd3qmaj/SBqLdqRDquE
w5eJu4ARdZIyJRnGs1ElDkB6sunLx26GTGUswO3WWxYm/74LIxYyU5MwaV7ljzaUK7M/SwAqmUtY
w9EWz9Cze2UwZsAj62peIVmoOnjaKQ5R/gzrCpe5OoQYZyQV/CF9H/8AZdcYRsAxWH4rEKoQyLAU
OPPn2AX+fbhi3dnHYlqIkNm4dmNl7gMNVvot9Hb//Iw4Pe1TcWRvNRRAIOVEe4TpVahOUlLqdg+Y
8gcINJIQLZ6XUY7XqN/IEbM0qiP2prEIoFQDhWuCIDEVXOMqToq/G48wY+n+lMsVDuPgLmYjnNo2
ao+mWpWiw9dgwz1aF6nGI+emcARQtFZS173HmfEcC8XpYR9swSU3quUg9mqpo5V4zhTloB/vOZQm
Ai2434e3oj8xHZ00SwzU7nDjMpvcvks88TYYKb0B5O73eaNxjGhm2SBXmOAhBw/FBKDka7Vc888J
exuIVmtNExTLmRIPIqUv+J4JsXuadLuAgFaobOkSyJQepmiKi+VXAkWNAdJA/jOiS4k+INWLrDG7
Ipc8o4C+YY/7S8BtP0pBZsNNsvBO1Bni+XI+aLGGfY39rbrIqneoQ/8Au18o1sljE8Txfxa9g15k
VN8+OhqkReAbz8gdjixSx66bGJ7UQjcLPFxW9SBajGfw2G9Nb0hIRg+FKvusJZLASWHZ5TCaRvhQ
R5l6eaeT3lULQNSd3U2plELMwOJyUl6++3s/I1ai5KPKMOCSbsddimBu3MDF5OClf7jA8iXYeWrp
917YIZLy5g7Z5rlvQhEySPEQstU/g3lvBCSoh8RXq3sKnFUZ1W1VAxgZsK8FTQ1O1G2gByv0XtOs
c3XNhaARowl6wB32rOHnd7makZB6gFb5Lxup2bphVWXOos9kYHG7Iudk2K8HZfu0kxl4r5NYRkAO
oRfpB/PLQemFRGrU+3ox4sgGY4sXh3vzj+UwScY4T8B4gK7XKr/9GlD+OE7kWr7cEv8QYRNYGjdV
W7nlUaWabwwC69jpy+fD2Dq+LsWKxiL5qUcU621Zq1sd+Pph0+biuotzGdH/TNA2jB5kEPDGnBtj
JGD59+nxQa7+zRtmr0xHrQqs0I8nufoKGYlCT2dJjiORAx3tt6ajMNCbSR9eu2PhL+eWliRZgnV+
jn+kHXrXYjHGdRs/MejnjRDTEgAuJ2uQv8eujY7cbWmSUm2qHHn6xLpG/nwo9T8ZzRLQVMpF0WtR
XMiv5ES8hur0dv3e2UYsthRz2iWQipQBgVs0aRsfB+rkXqtvFAk0IcDTKw7KLZyNVrAYutUgkLFD
Vm68kUzqTioVwMh999Ci7IL+H8WvsnSUlkbt6IZ9CL2Dk2l6pcVud9V3Qx7/xr3BLd5SS/Dxey8I
Mxp19ViIL7vbgCBftTTClVc4kv3jMuIhPn+gUTN8TwQYiLzBDzjYXFKcfZHqQD9PALHn0dkIFARY
svkH3RBAhyk1hdsFjMQRK6gW2dzp55ye4aZkq7QHs7AJPwyNgoEaRrYx5cbz+8hoZtrFR9jcL8N9
Ba/oOgzittmCDCKr+Z6us47CNVqKDJcHk6jH0mdgyRMTiGcGUbJXZmYLOTFNyeVi0blkSo82aS5E
HV5q+SOEVXf64qiqHSsLJawZj38sJmjFybq+Fm2+tmrnLZ9oL755QmblC5uR+R320jBZZsxHWFq1
nSBleO6aaN7tcpIsKazM69DdEc10LxertBLBxeMTxBsstg6vindLgr3tim3nxWbxT/hd2Wut90Vf
YVSjnMSfk6HIeMjoWYjF8TaNrR0Eur2ZnUClKJEHLMrZrWRD4HscOkjZEKQqV3FhjX2OOARSkoGP
CDBh4SpBuzYJ+W081inOH61rl1bCpYslB/p6/lLn22VRGX/l6U2sWA3fW27e1smhxFLqMqHDKF1r
7bPQ+g6p6Y5kvhnO9qEynvKgE5RSSx7ReXz4WYBzKyQwG/CjiaP+yXTBifYBKmXdjeqWzGQ7raKM
z3UmLNY77dSJRwMO0IZOb/vjSnC+1Ba/j8WcJ30f1oK4PkcuSFRDWLvwn9TN9UaU2v1qdfr9g3Oc
TmOpFnVBJ8sNMyxb5cR3jABN4duerU90Z3Vwco3GePPL66baipavJAU3EBcDZSOFX7gAptmrV5Zq
oqGtPPb0VcwsvZkd3ZloUTAjBLaNDjPM9sxI659yzxVT0yYySjQTfkWMCmcbd3GmrvKNSccCCSUp
YEBjyQonIv95zGmAnCM0My2GDrQ4GOSvyU3URveNDDsqcD3eCod1b9H5JxE62Tse34RcuCeoJM90
2IGEh7W6i9S//K7GkkcyOqi/4+EVfvUXXZxJCe6iaOGgzxyg7iD/ozw+Monfk4Vd4nOztwWFVEhq
tz2pBn9lpS1JnQcD0OVKN/QPDwDEbWwFJnd9d/vx2x0E2PzrMe6qCpsZG7oC8y8P8CgDWxqqkwYa
ZMOuw2gD2ffDm6vSTLRE5OkimLT88eUu6ehuhIzCyqAbCmraRZXwxNmu/bwrZwGuFtlbEx2mob6A
ZZegw8+6QPos7QqjzZVsagaeGndsu0BO0MB+T755PnpSeWcTh7XW4yl5snHAhSZHUqcIwQhd13ab
Mrn9L0RZRkfGtPad714D4m5E9K6czYDXGpoOoxra0zy0Ec8P2gcaSbyI8hOye1PqF6CkVf+uHElx
lptMZA2fUoP7TWyOtjk1IvF0AClvd8/U2Ali7kp5Vdgo53l73KteyDlRKBoVv/l2IW12PoehqD6L
YyIW13VBVl38HsZsSEueRvEle0Uw1rEKMhcTDBg+F9sh5p4al4tv1t2DR8PEDHx46Q+Sm2SEwxG/
MEV1Se/uiSaqTvHGrYAT+R5zDsyhApz8CC5Xtl/DaxHb1fm9Doazxz2uMPTDJh0Ulqi6fz9M1HAw
PJqS8rkXOSqmF+2c8BsEbEunr83ZeAsLZHbJokx5PhxXUPp3Vf+NoZ86c6efZbueZjZfkVwR9Rh3
V9QpNTkm0dK1FPTTnLoLB3jSauWgFDee96ziHQ9AH38ljO+0WFk526NIYOBJLk8AfAvesbuIX1gW
sLILUlIVq33aE3jUvK2dllyBGGhJPIOxOY8FH/IJ1j8pfWNtCeSCsC+38jZLirmjGOA3X8BuWNDK
neLjvEYFcDbV1jYzPctgRycJDqcng6H9oWaWutvxjCjl7py2EIJUhj1+iC5Aj79ZmxbKROSB65jQ
bUGI8n5tnUTAOytn1i4o+P1RgkEqZ27sIMoIu8BCJYPnS9MYNsw5Gao4GMhtiHQVoAKvUt4jvLZS
HRKPfYCiZarSQP349tO23uz/Fh6l39/ab7Ni2isNe4hxwkyNFxfO0rKLAWsqNtB7ivLAJ9baEcSy
itiNhZxPDCKFn8sGM6CyudLrIIGtM+J8n8YVDHK0CaXSWsmawlHqMsz2okKmgxslq7yR4ne6qvIW
4t5mpIkwsiCW4LCCUqfB4u/nK5qqlyIl/6/IFGjZQcC/QhW1N273kbN3AGDv+DqGe+v4ydug8CTL
cWaegjTMe2A0LMOB464k37cJlnIgU9clKb0JXKybHOQOFADzC6QvRcU4QtO0v6EY5zMZbdW8PtdA
ohdGVUgf+bIwKxDeccgqzbvFWK8SnrEg0ivG7FNPZJJtINVE4CoCrMWunlvXSBQZVFxnq9M1T/Ja
XUsVRVZf4VGZ4UCti9k5WbtcuzpifNTA9wGaWJlNm7k3FqQiVa0Zg+lgmtzsyeq9QDwaNYGysgiP
M1AF3YVAxVqnJQuxLL5Ch9TEuvN4IK+2CjnkjPln8nKQZsIQGgX04zb5F/ZMFLBzYMRJHoQSC6p0
0oXwASF3x4gBA/UhTu2C/8vQicG0kn1fmSgQ323XzR6RYGWNw/S9BasvPUjtQaQ/CRjQ0h5Vv+nA
X8GgXpJl6b2oFj6+ujMY1rt3QeruVaGISHsNAIbj6ZvG/dAzXJKBVTty+8LM0vN53AuSePx+ZrCz
56QqTx19KxIFvV18BtEGnJHtcgB0KT0uSqYxgD3Gzd7N4iKMv2fuOpdxwmOEcb/eAiX5W/z4pS80
AS6lkfMd0o5R9xJ3oc0W1jGDbPofLxySctsXx6o4dKwX410grFhB9xP/DVlXf4hEcR5B0OZY+j/v
mK9RLqy6868TZ3omJewQmgwY89KwjVJWdYRNQL0ECviXp3vhQ2kG5qGsJNURApxbcHN55Y3+WgpP
CZVoMwew4g0LDt7WLkhBe9BOCCv/uUi5FyypWjz/5tVYbIH+9Fo7cT+fUNYClvq/bWQWuZWReSj6
m1lxt3D3snj6i3aKLgHobzCAfAZV5pEDADp2+98cFK0FBgK+mGTixn2fJkp/iuFprguyw3KAK+pf
FnTFV9ez/BRGHd3UYAkgVqP361obydPOQN1t/FlPqHlRKICl+cjTI+71UuaG8Mnzrfg1B+8Ov9mV
w+/vz7x1cvbuO+K1pizFX6Gq7tIg2xJo1fuRYl5Ij85i5t8K+4TuuKd0ok6wsQzECz0Fn5OA4js5
+QjOZMFH/htEMMASYw4KG3bC8YfDCVxUDwavVvIiO30SCG8B8vbwMuyIgnEd1AQT7Vu9HH8/pAPm
tPs/rYcifJ8u2uTJr65jS4wYH59vWfqC/DSJMBIWPXJUGRc2OIXb7DvbJCyjzZyW3HHpQ/auLCzv
ZYT+21wyY6XoEb1DQVx78KsNgleo5GEF1r47ZVF9QHIMOUuOCGo/aUi1XFXJWNqhmcRsQ2EFHU7k
g0QjFZt2JcAOLICgQF5/A86kkSsfY6Dp3zWNSa+/Kqxb5A8Nz4GdHN/EcE5wGFKVjiM5PKTZeWgf
Mo6HDhIrh/T78QDZ67Cwv3uVUI32tS72RMNq/iOHW/VzMdjhN+8kDz8dliZZVRilVWbwjHpUw2vJ
79m4czdQkKumdGEb+yYSBt40/0occ7LwHJWL37xCGhrOncOWjDZKuEEIGb6r/8sW95koasHBgQiv
2WyZJTHASr9mopWv2Jo4WoyJd80ktCU32bgUuQ404iD1OOQCn+MezyS3/0b0Iqu5iKJNpdL2ptKg
viHZ39IpRRKjKHEqwrSfaJsLJba0Q+2cyf+o1uvnlEif3EQ+3qBmFv409e89+a5QqZoh6bj8+8I7
ahLhSWe3mWkaSvEOufqJuPAtpq5VdCp2APPLt9tT2LGG+5kUPJ/IFJEMwvH+KgAvIV61R2nZjKsJ
dbKjUZMKeZeseMt7h+QrR3SWsr8FDAMY/Oli0OfBUBj9ICP5ObiXIS8EdkAiVfALYBVgiD0+aeRJ
t3v+hhQCmUVF26/fBAPGMRoXVShKqyY2Prrb0NWSERj/5EzhLkRQwlJScafEppuo72DWxyc9B1fJ
+kEqBTH2KlPvHEzg1Bts5V257smwAAJ7hJ21LJTUp3Kub9Teov8+uuOUS5hyRF5UBT/scCmBAo4T
iFhbtVwU43kdIx9MFkQtFqSj8VuFRz0xYLkTH/ICPwNjTqKT2+We0Pch9vgo8eEKRNeesw//UWq6
rTLAhABeHBm1srsn4tmuJTTsSKZlGkjryZgKj9X1xiS0Y+pr3Co8BxbP7cE4xdbaCKgDnxRR7JU8
szAQni137SCSmPVjM8Ks8pWNS+cnniQ23CVRwYsVwuI1YG9WXi3aY84w2+6JFC/gece95Zibrbzf
hyykhfI4JfP84+2vGmKarxo2w04sYXpG5CsxMAT3vfnf9po4dLqibuDOf/WKTxTl0XgmadgAD0yl
z08QvOOD1GPw8CIOin6Iwg1LHVXqKfY8WOy3r3eOrMFHwUgmydCooJHQHRbxODzPWJlUD+XjYaD4
45VvpCcBKHit8nscCGlrFa9UkhzUum1vS29LYGNdpdGttlZhGEqdUSSp0UdQwWpYw6M/o6k2sumq
DRPheIXoIN2kl+BQmaPUvBlw9Fjbycat1MXl/VlT4JIDCwMqWSZdQWf2RNpFcWqTSVNLZ3jZRz2L
Q4yC+5OmGDvKtqJPXKlPRXvO0+5d1BEayq0WstxCjOu3St4sRue4EFv7VtLGXzVNsSKHI6pNrg7e
tDJC1JX/l8w7UKp+GCVyudpfBvO8/g7OMNjjysxu3xfyu3krXGFOvkRifyPE8g4me//cNA4aRkBa
tTi5UB3OOW+a35ublvDrovVb+y4XjiE0aIa39hpATLXovOfXVRKpTZpcTy0NrigHhOzsdJ0z3tQJ
RmyWDlkDJ5nVOrZQL+SSW5stbh3SujVQDkdujrt8zCKPW9JtidSKrnAcxS5pRO01NWMkVhGhLcxj
e2Gh+AQiA/cxB685xcLoMW/giLVTvNlKUc285hDhQn/HzGJtHAzk+7vv0RfxwGFpGfjqx8ELzaKL
MyCq7YkK3FEfVlpAVoZJvJgc+H16GHhNB7MZOmUIvBNZWAf/GIaIR+kzZMRDOgen0bZDTxULffT/
n4PuRli/rvQB+9Z5qjewMuAGGedJQ7GkB4/WZEk0rxbYsMojKxPnnCFi5C3dCEo+WZAXotoHauLQ
lFhMWbT1oSe7K3eyG5fknu3JXfQJLefbwzcxpAA1DGJzlJ1RYcfouJW5cS4jaBXEZ9R3e6ayPMqn
g2KK4UEQea7aK60rp+mCB3oV1s0Fov0rLwB6CftYqXlfALrE6mNKyygldeyW8bGNbzughubZ2rvv
VlgOk3B4UN/fcsHGaCsmDeTZpuiVE3NvclIC1Efumop6NsX0MPwkQMwX67tAJxD8ItLaTaLfaK/s
Xczz6HmDY9L6B7fxMeTP2U/De+Hp3RQUhdv/3ZqJV3G5/QSR45dkkEeBdsikSsBlX8xsULOyRica
XYjJsi+mXA5YcIpPmAezcU4irIE1W1GNTNVIZBl9G9QxaowvLkGmQnr09dGA/XfY1hcHnydzQ3r2
DqVeQysA2Gxc6lwYiR3HvZbU7n6b/MS3auEnjocyHD8Zz78zqIvXQ2hiLjDwKiqLSxJ2bQqgMi2p
bRi94mKwG8VGN0zY9aig307ZSLKRsnKgJTWQktsj1sujXQQ/hUrek8XCphrE1jSuW78rTeM5uvi6
VW/I1yrbyTBJtrgvUFodkL/oRjZmTQbX0ER+Dw+dLyTaogshuMRMzv/ebwB9Xzk3iBVKeHqKWGlC
bQT2Tk6HQakSzq6JV0rgcK6XbdD3V98aSI9q+T/02/u3mRW6/Xbcs8+1yOskQnjlKVmcvE0tdBJK
fRizR6azbs3r0EuhDfMapBw21kIDJ2A1AAFoVTbsjk/hatbrX1oMb7YWQbyzl4eX1MdgtubA5zHh
z/dd0UKwtSlU9QCirZ/zHhkDM8c7ClVGnvYEHZfZwTKVDZeewcznZWiBT6QhHxpYcNPSE3Q3v9KA
meuyngGwQPGxlHJF1N3ecUU5o0OU2twRgDEuqxQNVBkEoQMkiBvcl9L+6pLLQl795H5qAktgtNrp
T+JvgNshJ1lkh+yNzg3/nTkQfGJfL5lx3/BkQFDNoFfdWR4LOHjnI8RvvxQdpW8q97cZwlTaKoVm
VSuECUZHP8KvkmmopXD65I+DrxNxQONpvfxhvMhoqu7rS9D/SU+d2qlUto+eyq14xxjeXMuRgZqe
QNn0zn8vXiVUFTqgkCLtILwv929wgEzXEyrld00A7fqN8Roon/iFHh1c58rlg6VvSWh3RQbOZoCB
0xOzZxUDTADZIhrTtUgKECqVUPmcwLdbG1BlUNcXHdlDtWRxv1Wk77pUKeFbdzPF8XbILMLngWSA
rbAZKUlpg/az+OzQsirOFoOXRwd4h+3xJF51qk3SqJ30Ds/yv9XsXL9HksMJ+p+8MFOPUrtmRu/k
bXhSflSeez1JLMT3WAH49pde5yM3wThxiQRsj1ZTVKmWOaDFVw/blWAekmQwUxZnfxTEUB4c66qI
b+HlZrNKWDBBOJnSy486hI1OiD6tE+Te71xRQCoXZt12dw79Lhx4zgCsY+qN0Rltf/rRcxXueXwm
9ALdD65F+9IcrQgYOEEq41KZP1KZ2i6ABBYyPIzkeqA5KfNcr23vAGPVt93B/MWRNrju+EnDhlMd
I6PCgi3/+dM1xAg1WljUbcd2tLkYFx742k76/fXGXLTrpIORSHAAyGG2p3zBfMxQVkIWbahmEhgk
Se+Cyo/hJVUpA7q4mWYPhFrB/7+CHsKEHpYEFlk1PJo5w3HdftacBIbtJaUkpj7YL+mVCl5OB7JR
q+vqAlYiqs/95e1v+gXE+5Rz8L9mqPiqG4LcPAyTZwFIktkft07wBayZiJLET+pQRhvYH1OsZr28
HG1L3UP/SElPbt1+8jNCdseOnvcYsK7ZibpHd4+G1yT+VOtHND9djohaWUJcgWsHoKDnxLVcJ8Ar
nb2Yjnv0hk1iDSeENvCQDq8fYpKChFRc3YU6zXsckqnHEb6G7zA6IB6sswZZS1uB8PG/dMuAJ6rk
dg4jaZMkvwGriQe2Lcho3rSyUYDOleYVtPKuJ8oDrOuTqwraagjYCpVZxHBfWENCV0VTb0EdHp4T
8vVH1h/wn59TP3cde34oYRZs+Z3wnHQ1gKKECifcm1FhM3u2PBknlpX7TuVtjTYosptrT451idTb
CLFw2lJ8TXD3N+JFl8oOdn5T+k5ShWoPHz/NF9KGmWifnyoy2GGfDynkQ6jzlsqcQ6XvS7UP3Z18
RFRg2b1a5HNCwhtwfY7whs7fYesQPwT/44ZCChv81coC91aXnEBdd6r3Q7VNVmRDJKG3lhUx44C2
fWzdclImbL8ovvnSqHbRBZYIueUJUC5DouY6jkhhWEynGuGFQ/KG91MeSaatFucp7DNM9Ttl5T7m
VyWkS/aA6dK1/mI5zT58S8uIoSaU+nuWraqrlv8klYAkNbEC2EGiC5EMvYT4pDF1X0f2JehWGtfe
34ooqJUvSlT9tF/OTEmElsD2cljUXmE8Iw5Qw5HNmJCGcrqoFYn6YrjHZ91cqBsRysdvVVgYdT71
7c5YaevetIrf3XpG0fh3f+p3S93KfODptRB6CXCO8p+7iw9GgjhLmzZ6WHtZrxO/xg1icLKF+Fuy
T/8vgMfEi6a+bt+p4z7fPi+dwDKM3AzCkhd0y9dUW6fV7+AGj8RGHpmG2GpSie8MPpU/qw+ZJt3o
n/6Ff5RJETjF2rU557QetZR9wp5qhbGLSCQesmabFLLU8cekvLRJN52RSpe/GXRZt/2o8vMwrvjX
A9bua+kIE3oOtrxE4v1K1yiisc9sUjcum3I3WzMqGD9VkhJSYiPaBes4iwHm3HI5cJhGSzNAKKSs
KxbNyE9mtI7dIPS6TeMISPRFxtbnvacGqLWCdQMg/a5kf7vOiFYNag4OiNi+KHxpZflLtOYQg75L
KiuvowjSyoc36mJTcUqYJpqghPWc0LSsUocZXtHlCyHGkeO2TvbdrpXFCS6Gk/X8vzEvOsJA5/5m
TDi2CphViywhXaEou59s2Y9+dO5XhMa9mkuF/NHyE+TkL0U4mBe/xyjyGwwR1nrwJfycv74Js6t1
XmVW3hKMu7wcuahSqe7pRrufkL+S6wGA0IwOhYPw4B3DS0bkZIgFrV6n2nw+cdzi273VfvDAmuk1
dNkWcPuAa+71kXi1ne0+aO+Txb9h3xYR2Zh7qoyADyZrz3dt+Y49NrB5+T5AE8uY0xFcENnWbrYH
OmO1hPIhHJC3kxpKP8p+XzIWPMiZNp9HLu6ceZonw+lPMVLWK2uZD9Bf0nh5hZ9bjXN8HivU5I5F
o9GuPUBgFiCGtPW+zke+m7W84u/1vhhqd2LwG1Ym2PgPsWMWY9C7TYL2AcFSMvdR+XB2uvld8QUE
vU/c0qJXDE+pt/nQKtAJEalK6//w77vyUroRRhWAEyJ7fJv/JWYVxexba064Dg6W4Kd1LacJXIOT
eyuK+NujeJKwdJNk3BCoWaUXpR6V8hnigWz8nzBzNGnJewGZfBh/dAkaviY8Nh4sPTXa6toJvSih
Dsv/eDqhCMVec4Gh0Xp0uP/k3rcNz1zG+rlX13IeQ+Fyd/C2QTEheLsyRAD629+hJ86HmawGwqHq
vxTva8NIswhyspx5NIm41wReSVgG2FO1jM3E+XwV2VgdNhvL3BPVq0UbovVnKi0AYRNeudkBccLt
srgPdjkDIxmktovwTgnJNBglIZw/u5GOB6xjWPaREnug4erpgnEvV1sCaLv0AqQjMV+zISG61pG1
c8Tqod21UbQT53FfMUT2sBF6EDJjwEkUR1yWbvp9jzpiewzI7ttwKRhiEfCeL4Ev2ZZ0YkStYiNh
xmvXhSjYLIWPDfHd/hM1NfQm/eQlIYTYyW+YHAHy9mlJFZ+g9B120BAmCQclC45dHsa8t3hvWEh1
VE9+JOAbffLAEo9Zp47lfA64Uv5XCKTJ3BEHKcMc6A+Zjwm94zLV2ijWNoypfxiwgfVOhDxUzvdX
BM3kmRT/zDG3CnbUhmR8uBhL8yxYAZNcUlBwiAD9XbSk4KmBr/sAynWrY92x8e/k1ej9yl4FkJoc
im8zppD1NXxIflPku4zmGqXOjRiC2eOZJIE7SHDNtJrC1dnGTN6zp9EdrSOcCCifCao3eR6hdGkh
YML430fPxkrcwD9P+xPF2I35Xf1UpxuByQ86jCXxQ5AlNzEz2q3oBNsnQ4xJ3hi0fDLHFg93+UhA
2DJF4sGaOW2KTZgdQbNcpMlpJwDRJDGizgmdd/25DhUNmqSxqa8f/2sfTbnGGCrt7DBBJBwjaZ+l
CqoH9OvZHJG/Q+6xU8+AxkDmijF0sXtKHVHFJwt62FkrDW5j13PDdzU77oh2WHWOO3hQIXd7HXEZ
sy+NLZgi+1D05qxdCiu2qwev+2vuYL7EDpqqHg4uyO+i/NKFD3Zv4gYEvPGsOpIitSk54gzFmbDu
NEiCKqx4RJYbIO+/NV1P63enutyytCpcWDWpMSETfHbnfk729BazB+xNJdZ+PN/5ET6PNHcAFVBM
AAUyFvzx02FIaOYzgy8o88N3rMTQult9ri7Ms2676JQB7kLA/v0fiW/LTPXH9wp5AKaULW3tJy1A
RwdXlkWCbD1c6YulZD7X2VhL3LFPAltd7c21xtQ5TLlaFIB/CqiGzNaAKsCc0kxSAkB9qDKVZIUv
/7rA/+A7PgXNzDPP8qqFa92mD95IlEEW4Hr5dl0CPCGtzw7Gi9HmvL3aw2TvuF8U2VPOzRjGyAkn
vQ20uACyEQkX/7mFOd95GzW9bhTgpIXLBUEtOAeoAXWHniuvw5IFtPtiX3PYexKSL0vWdjkUj9JP
CYSjTW17+bIOjoE+3zngLtsiBJ0vVOLaB/gRnkmCjgjhNK/xJJ0gfYx/GR+cqyzGdSPn3vLZvPHv
8ibWk+rrs6rsT1aPQG15I1Ts/hCR5p+mM/yDqohW046aNrvrqx9cwvJxvGro2GE+9Q087tJHnXuE
Ra1AB/esO74Ykh7gDpZapuV4EzGk0tnkAvCbxroOFC9YfmOZVTOGZ7UoQXduZpNP4ZKdp7GDTF+O
gDKHP8O9G3Pw3FkLcKc+AVHETkQky9YUYM8WVwrnE/PGZM32OPD5fM6saNu77xXm9PyCbr6mXLqT
Wdr4CD9YUC1XdVETXycclK+Hmr548GYMdcztiCTZnvGI9cjTKrbqPjThuB8aIc67qM5jMj1vkTft
CaI8RFWYr6BCdETPeah8t9rrKHKimtNux5bu5qL3PypHQ66gEa5cJkJZbLyzPyKVL+nALSI1JFXL
7gyRy7MqEGW87i2Dc94olXONJk3+9e4M/QT7DnQVhvhbq849nnkLI4JA6QbZJGxwM1/Wq6U4sLGN
ZYnOdQj1Mszl7EnyKPM3kD6q2Fn6zITrsuEhInRIMunaFgRfGR5SqOeoW20QIJhSGexgc2hTF29R
FP9uKWf6nrxPjxG+0+nztNOycnQOXIGJidlUdUkUulqKpMVXOXPj+GTQBzxNCzbkjxztjXwf0PuA
TR6LGG9XYxfd1BxgcngiU3zGH5Kx0xOa4SdJiaYeRlVPKLLtoOS+KshO4UkZrCqnfwxwmSMD71Zx
MrS1vmY/xiyG/5pMgWiYGMVsF2Df54c3EDFnSrdXeNW+HYWwCDWb6awquqg4RGty53U/HnErAbqY
nXsEeDKpzALU/DhbQloCQzD5ZnCmYoy4Q/e240bn2xV0wimMW8kUEPO8EpiXvzYV1zL+ISyT39Zc
j+4L51kKkq7ahh5e8mZwuN2uJw+ls3ZZhHwaE9+7qyPT8X/cpH+QhRHn4l4AcdCthux05Bi/dciE
WFaxZV87jym1fe5PILMbPlR/vyTwfJRaB9cTSwcRfWQUspKjs1uoqNOjg8fKxI5nqH97zmihAaT/
Olu+GwrE9vtXUp+2YQ/qU9FA0sTVULdZBwD9BXpRnyfsHiq4VT7FmhOe5wjFA5y8QWf3kVDwfkp9
FCd49hkwB7DIBPZlDUxJVLo+YgeqnjYt+DvGAB/WioAPDnbt0tSGI8LxOfZvHSzGULQNAiGmd/gg
ns884JPqu4amJXcl0OqK1Cm8DqRsUQMU7AfVuDPJtmtR612Bb8rFleEUdVXJaY3GdTfh9sjHpWNo
aMyIF/3Eq9AM0+4fk0JLSQcuXRgRtAWj82Bl/VpboWqNY63/07zpMqrrdfaqH5tgs1947kbEB1ZA
xSkpF+FM4BdkhhJo523azbHVxoS0LCP4RsZ9tg4EhoEAjHzy/OrnJN98h02DFd7K+8uIV/Frgr8N
T7mNHXY6lQgp6uXzJSLTRjCI+WPxnmSjjNBZhYQWxU5eoU6fdEmyCN76Aba4BL38cCVSt1fV8Yki
z8QEQdPRgV04GVBszlfN+O6gUbASifybDK9XCyAYBy4UxxL01LkbBQYBCBBBTHuwAQdoW4FMXKA5
lJHwbev1GTjb5/nd9npXISO/fS7WufEoNYh+X1r5rXsfLuQIosR0l6Lr6vfHA4R+iNHIYXbGo9RY
6MQ3hT3rfyKCT2Of86t+eY2HsUh79uxoT/pr2z+NsL80T5bobzujrt3gNR1xgZOQ+EwxuCpqAt8o
jdYRgBm+/pQYRImAnAwcVVQLUpKNvwkTjePk67CzPoU5+XfOuc91b7Z/6z22/XDLY6GuEi37zfsn
Vd2+E+tEA3n3pl7+927AwfB3w76J6icQm/lN1GgUPbN8zw6eMwkaZfK8+9BO1bOO4IGb7kbUCotM
he2gUgd8vRTkzKqiN1ieuVzu+TPPXe06iU0fcIgiBcqp5bCEHHeZZ+wtxG2G9jSP4xlL+suRh1q+
HfK/uLvX/3GIHASRgHdGCQ1+tmf+mzD2gB/+rTN25/8mWIvR9MzmlnCTaebaPrhnBGxu950fjido
yOKfB2ngP7x8BlUBx6bXfvYjyB0kNk2nJWHh3dsmjpVKkykXDbxopsQzmNfdnfrIbMep2FfX5Evv
apv9YI1GinpUpGXbpHBvROXjwBcYAfMVUumoE4HXzSFcmk9TPHIylz78YKKTMjFTdAdxsO9v/Sht
93s+74LeEcLUxYjkJWp/D5ZlfAHlIns+VSZmMsslRgehJi56j05XaSQ8HrH9/TEgFgJ163XNX9NP
lyt3UfwssW5iZeHm1Zk96NhgQuYZbETwG80VpmjC9rYxg0pBdSvuoz4ChNafz4s9tisplJH7G9+w
dO0n6Bj9CqFSPJIx1Htwqrah6ozN4ymLJJ76zzRtFhFVPjQsNAnRnrAafNY5wK8yj2QJzhEavNbG
2h52pHOYhxjExKtkS9kUT31JptjozLqn0x9AxXNsmLKH6t5btrRnYg1oGmlKQDDtr7v8T8kdmXFO
5jSMGsxZY93ZNOIcaGL9QlurrdUclz6qcWZdMlkETtBm0h4QwN0vVI3S6855iPnFZQvulGWOzUzz
1SBAwYtgNsuAdydw+bPb5F6RT9xw7Ub1GfxAPQsCwjwsyPtm+Fq7jQz/upE6tBIbevCxf8MAxFJO
Le14JLawmVpAWVoB8mJioM9fO61KkpHWn32fJ381Nk71kDdhxMGfbSDTNTDmNHiV+K7I+F9TVlaP
TYyGrr5MyMR4HkR/1PyXU/aqoe44keQJospu+6TtQar762/Hsxz4T6lLFiJ2Z/E+2JjOt+SZjmKP
UKUYuMaq/2ismU9mGklV2yhpf/fXNG6MOwjbc+uvQ0QuDXbOdlOFoLmi6k86SLWFkMKXCAPtEAMS
hdodgM/QOgMQD1juJcQwMhSk+/PI/R2WXBMC+PrMxyF+MaufYBYf/izEof78BbImBNa5XAfMdr6+
jPHJmEIqhBOW0uIUca2qLkoHOofzhNF6/pXcVdf0mlitfIM5GhxGtB/dh8H5P29B01sTqWVz3nge
JDeTNT30MQlh9wXc4HA+CTs1wOL3RMMgODnjKN+blAHn351RD97U0WSctJTeQ/6Wua2ml3uIosby
x1TERM+cgn3WqrPT9QjjQ5M/oZTH6KwFT4oNCFfu8orB8O/ZUi5jVGdJy/vVxhuTMRby2sc+xpyp
6JFqdcRya8mX6EbXn6VKV6gkxHB/iHGwNfORNxp+uJuaPZfjFdNmeeP+QxQeIe2jw7xVijnIJlU2
5MpDknYxG0eux1r9nojy1dGmvcBM2uxjvoFrVRMXliFTZZUvizOc+Jes91s9cwuBAZUplg91FrHu
CsfNFQ5JSqzSzpEOBil/aTIhfrz0oxvGw6eymPyMPSoyPV1WJdSj3VFn+kFcqEGtQ81SQfNU5BYv
rbeZI5pSr2frqGJJBOKsn7ao91COXzI80M+k2lYSCP9gzIALkhVWUd4bSvVoM6E/a72rFTcbqeUm
xHh6WpXhumz75IFSL37WySiYYd6aDqQfR8K5sJVw38bYRPt2VYcl9vQ4V+AxgtZOZ6qGqL7NcFk3
jEo30vdij1wgGiizRuFPcg99dDC5LG/VyEh7k9NA24QwiMX0Xm+Ek58DcvmIm1NN7BQUP/MSXd8A
pg8OSI1JwoToqwruw9h7xWPM/8ft70cdliYRiFBrsaLM8CcpaVZZ9+Z0LsdbZVkdE0v2T8C6bmVm
+ONN93vE0EbDOxew/lOpb5+xaONhPu6ahFe/J2E7ytz1RTCHvaZpCpGrnlj2N/9Xw0DzBsM4JJg7
NFzEsU9Vfczq2WtdMkQECLb5TIzebHCL4ZzFF9za6BOqmzDS/DI4FEqXgPuAc2fJM+nO5mbnIA8V
wkJ8eEZg1l24kl/wdqkoNeaRgVfKdxmJfZS6iMy0Y7202Vv0qbTCXfLSyrbGrFd4DUuPYVQealcQ
S29NnEHY+ueLs5YjFJUOJGOT1UASOvKFPLjpi3Kn3FI3RWPcyg1TqZxhKXJ0F7jFwPSMnpvxPEuB
zuqj9Vw32daZ9Mpxh8Jg8YPFTsXgPdl1VQ5ZF52fh9CteMoHCLbDnhY5Aa5qrDhH7VMSV3ntro8H
r8WZP6Yqxd19/8il1hBjS+pQirolvCa0CxkNWejtTK6cGYHePyr5n/EdQgPljIw4sxrAxngK7gmC
eGl+THRPb+NHKXrfr5C/GvD00snSGP7WQJL4rx+pfes7LI3oNgl/pqayKw5jzcEy6hTdHNFzhB2Q
51x85wW0fWAqTj01/fSaiTtmZ5nPcK98GvflXLe7DjAjnWq89DKhkAA7Mya22gecWmRtuMHTVPs7
5zesL6/zs1m+tgTgxS6IbasUijzy69qGzE1d55/vj/CaNtFJwho1HllZm6kQbOYfJQAJyr1VXdjj
YZZZ3ItCpAoEkpwBBbWVIXMkgt5N6LMPj3jFj6TFVsWdln0cf+EdtjpNfGqzIjzNNwqOZytMFF0B
QLASw8EgsiZapGmR6L1AwcTM5K9G+Ax5jQOTpNGMjnmUhNQXKqIefu4KFXm3HbczhIlQPAa9bauK
vG/jkVGs0thU+eY2Pz8c4c1CHdgoH4EfpCb8p5e/JMBq58P6Xhwve4nWWblFHTIyu5zdOAS2MtxD
wNsPrIN8DAh9FeMTfF7IGijyZOtu7p4v13Ykn9tfZ2IOsxXpFH4g9w1oSxanNGiNO+YHEq8cI7tc
juoXhaGSmf0BlUrFz2AutE1iQHhJbX/KCum3wKcQvSXkCf6hmjBUw0uGvh7lJl4tge6cpx4uFS/4
a+VsbrULk8pTR/vomc6PUo6xk8kPZc2IQU2XgxbU8aVUlG+bGWl+FLpzbRc3NSzQuPaqdOgIuBMl
oD0Qf8sWBkTN9AHZm5JUIewazcfysJfALE418AURs2RiyN3+k9SE/p1gc/XviviCF4DhNRC3PZLb
ecf+qAReiSXBgTaQ3Yal2mJBVY9LRdAcMGMFDiGonLLihDEFf8oJ0LejdG1TCO3YV0d70ANWkcGe
SOom2/vzb5QDx5KblhQkdqU+aWDW9EYGGaD4lSGM43U/vejhVAJYkcXLkjXB/9FFD2+xjWiYLb9E
5oO5i4zs2GlvR6sD5VT9ycqBg1gL4cPoluQ34A7qKzvYAxZRV21Fz6eJKXjFhSqsQExDe9XYbg+3
QOXOMv6qob3OAJT8yKpNWagCFfwndetUHtFbVIFVtxZ8EtlQa3UfmdO9gb2jLttXFZQxkq0UgLnh
CGT3veSnnHm5b9+4iYNnVD24Iz5H+UsMZryfpvmvKj/rKWZLlWz07k4AgXjJ9K1eY6Q8n/g1uSa6
tBu11Xsdrafo0Kv+sT5Md32yMM62Ar7e3TTtgRN9igVWHN383jLh0fCdeTf24DEnVn/iLIMf1Uc7
Z7EjCurcVSVMDTs8FUSbi37msW9vQVc1CGTk6G785Ggkf1QfeHTOkrB3Xi6UujM3QANmyNSzZphT
iTQ0mn5jwJ7htxVbyskXoxmeThsyKGsNgxTbCsELPa8kD3rkVi1/7vZ5OVaqlyt7JGrc/N+Pl/C8
Nit5huM6ZEIuQEdS/76tZLqy6a0gjd6UOAYpbG/gjCdgsC7m8gqUoBpTluQTh8JbFcBHLIGG+vSw
O/NHspisHBRPFeqr8EspoAwmIa+Mwc1e5ZRw/1zHf26B8JdF83Wy4AXQSQgl9ZqmIdn1OmDyMgSQ
AnnPQmJjEn6mo8YnAEkcc3h4L5xAX/jVujOMKU1VWl9rCBagQyTI+CjxxgJCups37iA5hoV9R7TL
YLpb0ae1KQFwoJ0eTCToFdE0iCLurLznXcgLSpqOEeBqyGYABN/YKBxoHhEoCrqeVqbiznu/Arjo
xMXQotxXhXE/ZwBk2YWDJCWov1LMckpV3KJMON3FG7vU8VlGaYUQ7d/Ap7p1NwbjKUep0IJf79dg
VNnek0qG3WPp/cSkYaBjCK0qWAp8z+myLSxv5WPJdnpu4go0PxZEaPTBAIczOiDUnfACTLwY9OJ9
XU9rL47HRxp2hWQayl34UDA/g79f+yQ1pudDGgrFNDz2B86ys4ttdkRAPTd/bj6be3H7Toe8OSKh
r73jmGtwyJACtBJBeV0Bnof9KfogKkI+o8DC6mqzcLwzRYPO3WpxqeCD43ITvoQa7EBDiNu29DJ5
pb1rdOQ0EIGzx9nk6WNIJJJ7Z8xa7dYOQp2Ratul1++uFm+/SBXeJdJdlEiEy62o1HjV56YTZP/Z
hDz83v5OtXMXKcs8AUbowyKzMgU55daBbCHnveMqrQ5UXZyKO+tHrfm8q8fTjLxGuCioCZzjFaIT
8iQOpEd7al98z2nNHb4JvQXSKpxlHuPqpaeJ3eLGxifQTaPR5TDIw6s/AyyqBO6HqMYjDMvnm3q+
yRTTYS+Wwm3PCa+obJuly7fyMAaQyzUSkC3hqX4blPcZydC0CZZLkw98U9x6BXuqHPcmcnMNuFVS
MWH+gdduIcIo1YzZNpMudIJ+Agk9a6SKWAaygyVsyDo3OFz9Z7zad+MuN/0a/kkzg8gRs5A68+dw
mJ1xGSS7COjmuRtw9Ft0htXeOjLhQkudnIOiXK7765dyXW3lQafDU0DvemvrNJ33YLjiVlh2hG+H
Kt5vlw/IWfeD/054RnsoIz7GC2GaYW+45U/s9LWDR67wXIVibbHwI+Nl2Qzbfd9rGICIXRezLaYY
8rU1MjZLClVOJFSgM2BO2a2X2nt2yHs9fJuI9FVbTpwCQf5jN3wXBMAuTHModagxM9jrR9/OdlGr
Dzq/ZaWbrQ9WSwfYrCrclMqt942662iA1J6ZLvLLip6ODGqD9hlb/QshfBMlyuRuJUYbDHj4nULq
YdG5vrE+fEGucJljsKUvw+bZmXMGGmDBmJXul0M7Fy7AN9Fzt5Bd+xJNBahVigBBF2N2xtXjRQIP
kl5sUMDdrTcIBGmLa2xrxidNP9fELix684F+Dzheoin7u21ZNZRb5RBP6Ne2n0N4r7xAvB/gAb4Q
H0grzDe5GvFHQeoBk6fMILu2HaKjluXUYA58w0ZJPCgeFpP7sMBGsFtWkNyR1sKgpepiTXCd1rpr
80yak0luTYPYGdzoQVRYF9M5aPzudoAxX0Lc9AKMiVjDwIy5ocKB5soNB6LAQomd6/sS1FpHLWt1
PT9FUA3D5rCvrdE4UZYlWHuBG0v4ZgkxZN/oziT9jTX3kRFf9h3aW/PAK5HtrT+RBk1u5Kudzm4C
tTtHhloFBL4vkF2jya6EgmktMcBVkJRqYb1l4Gb1eXKsYzjQZ86+EVAe3IhbEwcRUlIBUX8w65Tl
p27pL7ARdmhZoQlNkVixwLgPCQ8jyhA7DwAi3P4252h775ad863fxL2iDyPeiw3tUwoqhFdxX9xo
GDsjp8NexsBPOyds23fQnb5ZtVYwvuscQuu8UUINY4NnqOCNw8bMu5GrpOGn2oALU7Ce9DyUU6Wh
/R9ah8qFvqytl9+sbZjxHpizUJ87fAppH5aLwv1O0favsjei48XTG6UdLK+TClDs7IsjYE73POB0
Az0lYKQ7azo8y8pmgSb8kQP04PS8FAuDI1ByNgaFO+WvkdFIstzNwG5kwTGQA2iuWyslSFw5S8Mo
Vk8zDUk6apc/xy+oE36Cj98KQdYPcUK6Y5EYXZJrZ/6y7ADEkA1GuQXT69sRmpCK1rjsEANj1+gY
9LU6cLvSGAVBUrceBtpujjV0QUcJakMRQj2K7KGurRzwyb//ERWo6738T87vpCGlpCz0lUVdfiTs
B6KggtakiByr3luAAb+KvxUXkmRMNvrUe58B3HHJ9EcLx2JzAWr4ZtpR/jndmYVboZW0iG6VqHTV
Ej6c6BTK2Jo+qXgmxdX1MsQeL9W25ptAVlNVnKyxP6kE/etPLKhjH0oGkN1DvJTEHgAPX8D0q9td
WNFV4dqOFtd4OzpE6+R5m+Hg3PcCtonQYuYodmc70W0DAHYARck6yM5c3SYq/AAp4qzRKod4WxtI
K92X7Yw9y8UORzFz2C/3GIUxOAQLULjHFwgQjzNH4nmox4+tM28DHf+T7em7d6QUNbtD8OeSCdQa
AvgL5RA+Hs7iL9GTVenNoM6CELwUu3r3EpcaRmg45SWIIl6cx/PAsAS6G7uorzGZsJ5bDSyjQZYf
MIFPIwcgZ641xtIGqzLkstnMzlJiCdWZ4sf3kaJh6KzVftYphEYZdHONpOoqyzDg65Xh+dg6z3kv
zeOx0COsMFELyqd5R/yxOEsm3/j9k9qOy9G3J8SC+F17yWZD004XsFcochiUpcllBcL/SubOB8mG
IYWziwoylRgY3Y77x29fh64K8946LWSBRxRFuHAJMq8TQkHD9avfswJULP4DOA1IHq/td0i7Ykbw
akOxbXzsRSJyzDbphi9Y9uUO6UzyXBTJ8j7sPbYvbrGu2kJEXoWSMPZX1reUbEVLmziXtwEf7Z6C
Wv2fe2uf1C+U+pvPDR++k2ZkJAKoRSsPHgjANyWZhNwkiEPe5eW5ZJzcx2yeJ/UHMY+64UpzDZZM
OnJMjPDmDaWD/WyBNSNcya5FZjoGIz6Ck6/mbBnQtbUlulMqxlxTG5Or/1hqInGp2jOIKh2mFfx/
Q7o78nhsgs2dY5JsbqK1EDgLLlBKJCdsKl1rZfq3t1qI+r4LyeIYyVjElIFeL9EKiIdehT2sGXD3
nkhQKnq7iWmRxKKOtUTMdD0g6WLNPvFRbTiKvtra5Lc5YONU53JIUPnt34j9mQG8OC0fRUvP8oQK
zcaCY2hp/hJL7jt77bruGMvxj1ocYGdDN2zfjhsbZSP010Sf49fazPurKFMQ2QIe825cofMjRqSG
qhyCGrMTJMfInAU+GZilHj6r2HOSdpP9lUpZ08RJElV05JinNfPG1WQAOL6FaQK8JWLTIqnQU7d8
zyll/nh7Xp2cve/gAW7KofEc7ZJu7o1AoNZqUg4k9/sluRmmqPrUrhtVbmZMNp4HkSLAHopyPI57
/suRIxi7qSNq6b509/za6UgM4Ia4pZhIF53O7veqTnTyWMdemmOvHAi1rHa+MJ56SHcLrDu0oqma
oW9gi1nCtVZCuuhGiE5W5ltRwGF9X19OQ8Nguuv+TAdcU6nUzOqR0k9ChNFYANOTxu9CaXn2KjQg
PtZLwHdjSTbnRK1DKXAAabPG7LR2QZs87sjTE+w53UR55EnWWykDTlcFfvPTjXITmo4v2TbPhwvR
FQf2zJQjnKoEbnfhDUHZRzLt6QQBxVaZLJaLA2UzK0Pvf/ipbQ3p+mfrI2DFRJoG/DZ6+PN+hjKA
zBQfuBvUKDRzTLv+rLbYxpSBfPOlrnFSHVeSxx9YGBrAEonUHwh5UDij3zH3iXoNMS2E7RTBZXLt
wqsij/2784rT2mA4W/lLa1srtQ4YVGS2xnu9Wd5SqJn3BP9sGwzjkuCQHhOkYXWcYIlasqTrKGy/
K1g+xCk75Br0OMDU/ReL/DTk5SZGFSIOjI7/cyGw2ip3lhdEOzp4Sogn5T8YE3XWxkwz2P2ikIWe
/KHOBxRufg9pXKYYaIoUA3PaunFsQ3gr5h3MHrkbaIN4h2MQe3fDMh8da+xmCFKjgqEc9wzizlOr
gnMvsUecbDXgrT9kJYTsYQOhnbKn5rtiXXgrMBFAQ8/q4QX3Uemy+8vU3MSYpvM/5bfdfRdODec1
75ceYLLrPBOv8piXRZL/FwijoSUupY5zDK7XFyk2aJ4MqAGFw/cdx9iezzjxRgY/5R9xqlxT2wVt
B7utEMuT2zJiZAUmHKbYWYeIWyoY+RrCrrJ32H/ZApCUahS3cpvoyIWulkBWNxV+V/n9b7C8rMS0
yzYLCvXU5dZf54tw8YoUn/xLkVCcLO836i/j6t/Bwc2PNiOzj0oADV2TdQStpTgfFIrNhZQFNVcc
/pBAfV1wZ6xggtgBZujHYr67lO28QaKchA4Lxu8c4JsRtnVWYrA2QgAR9gh8GLPDsHn7Zx7oPD+A
/l7Dx5w0bZ6A08vmBW8ldMpFk5s0Lk1vtvAaZcvAURnwAlP3WNxlLC57RY4UZHtVbxlCfCnuyf0X
IsBoFLPRGCOeAvhrxeQr3JbiieWyGmg5h3pdbtlkYPhUukzXdzTpv044hWTMc9JPqg2ym+5S683F
X6apsCNH5gsOmd++l5mKTQmCSj0lONPChUezYQc5asoiOpN2Lt2fi+GXcVxhDNkczBhzKsnQxseh
UNHwqd990bBOn1CGYuKI3aM/a1UbfVsw36stV4AeSSrt8MKAGcUHbE+KMC9U+XezbZ/70mw0WJbZ
vjZtYiuzLqu+/AyLJsARdFvSUUks0AkLjQbY2jaSq75+JroYhD2IkB+ohGBfss6tA6LBeChMeKag
N3H5ITohYr/U5+tZiyv6CFA5D8LQ9uhY/gM22/JSaOd77Tlf2Ocyy5daS0852hury44pAJ0C+kJI
3KYmnD6kbEpTpoxkPDJUDOy9b5HqQCvQ8S5Oy5GKQ9uGJu6sj6szKelpit2n0wprgHt7fKI9fyYL
gzxtjsJCt5mXVrxGQ3kZVSzyfEgGNx6PPVUaKIVCkY8ZyIxFFD23LtAaBtW168JEUDCD6DHHGVT1
qu5yTya4MGzBgUyfPSMizdSblET0Abw3K3TeikEyguuovuZ+Ix+MGXk4L0nSvLusEw67uaeq9Xrk
jnERWg9BkjbX5HBJUVks6mk456cEAXoBHrzWSg3BMn+LUIscYB9G69dj/bBP81/V0zC26RwBunPC
Zf74rNVPUJ3lqUr7SODMvyQ/y16EGQNHKvvXx4K6ZdZ+lDz3N+USdlBkRQZHDqyowkV2L/pilCWG
O2IpEJ5DyJaCj2jZMrp8ooHZ1GM5LMTNjbWsRqLcoheoxPbM1JryTzNUFcM5ZAaoRj/ws1Qc9oHm
yLfUeduseoJHogDk8LLK9NYo0t2OTG3XTHtBWYJYdLzOG6KsNWt2y3yGjJfudZOhjRYEHGRUSA0Z
GiBspwlOlnHy1taRRUIyT8sRQkOprJtt8iXGKqhpxYXXYezZj7K6irRIWQWqLwQJ+AM84bXvC4cZ
Y8hzOLZxFZovpMmmNtzgn/ut9zLQ9oyMMktRTZdwFXDjXy1F5nb7rfgniCw2pzGFuqK3f4G64X52
6LTbz6e2MJV/620KptYI/zbeiuhXjQecAGsgHQgLHLbYUx6DvBqrUqfLBuxRI5T3cKF5pNxyCwcN
gIrdM4cPj/0fP3qOPtMippr5LM7jmoub27+7NdeqVd5TiUF26kQF0EH/LWxtdyiCtOZFIExVwHc5
be4dQbLreuRX6AX/pWm4BdkMExCTe+YyeRwfByQJkoJ2PGzQLZKJor0jTg2tpGBdCHnOIP0ERSzG
+RRc0ow1dzqNIoNLNlSYvj7WuRI5PS027dAAroaCu+N/5eTRnuKvAw/NIU77gukVt/A4aluaH1iD
NjE5vsN0I82CX+UEzIrw3sADgCvFviQ2eM7/oPjbwzbF1k7myjf4HioqlZ/lkKffSx4la1fXkovL
OTHwPKjZO2lUEqkXNIh2Zq+bGSMFsazWk8V1qBXUepzb27FAAw1g5I+a5AjVSc2fboLt189UF1ub
Ro8Dp/fK0uk/WIHgWDeWWm3fuBKtqXNguW3i+tCNqizw78A9ZAe5pyJy8oW18O1bFhiR+qO6OHPQ
1GIuuUvw1JfgaOQ3xOJ54IeKrNWiyv8oROxl2Dne0vnbcWeoCqD6AvvPLR0zFKTpTg9JJk0oJMoK
tI27ujgpDEBs1XxosIYNBMzm0SEmFw2/XmaRNhKyzdzGuSJv/dDb4+wHQ+IFrpyFP5DKgBoQS7EG
VjEdB7sBUDxCeXgBhishwHTubsifr+U/nfw3Gyy063/yZ0IZHgWHF0Ba9D3ueaHUFUwthuaTDci3
UGJUue+oiF9IPchvSd2Ge7VyN0hMlViqIlzLf6XtjTT3JsMQDEZqIxs+Qd1ekzlaUt01K7uRPsM6
Idjg/L2SBQ9QO/T4M+j/kjbU1eo+YkfkCzQFWYuXeBrQ0kRYuH56yAcaRDhBoSARuW96KESmH6b/
vCVolJbPAB6uqaJZSQ0DMZTGvTAQhWv6Blva5nIzF42AfviKNnF6zqM0htx++FJYPzEfgt7MpGeA
TCApVILYJEhLuft1Rawq+mc524gmjQ9UKABL0ZUbLHZAWCPEJ1fEJsdAxmP9UmtqGsyX/4sL+krN
r/drt76283eNh4CBLT/FhXnoLV+6Tr52TizXU+qzxNSUrTu/OsPC9s9UjDXW0SJL/EFkIBAgPm9o
uB0VJaDH/Ck9oK4qSRnoUaHaZVIqrigH6OdY+NxNxD1K+0XnM93SBD8EsxyAd2FzLbovhE9XVTCz
u2O/Xyej/+CCCsQyN1t+gmgyP2ZKJwO7iLG0LcrOnHzTVi1u+umKyKncOUjlTeQzB7umDkX1Rik9
YzmMQvuDEaQsY2afWW5aXighaTrm9BmE/oMIRGl6pmxucJ0DkSCG+V1uNcpHET8VLRoe5gp3nkXv
WTwhp5bBheqrajzjPCFpMZp/GZaL/J4WCbWHyfusbTVBdsOoOO4y3hnuRZgy+s4U+4yxGY0MvIsG
eflRTsoyKPPpWzIQCAfpblc9v5HQC4azMeCvRfvqSd0B6lqE34cQNl26ewLyYGO4na8sJ/puvtpk
f6zCzEM7FCbReyodI6MyxRPtcSBnC+/O+VZQTo1yZfdwNWEulMtxOZ7dVi2OskiG4zmBTAvuc/9z
L5OzEDA/36vKTc/cnkD9ZmUotCaCAMqYHpuxIxkNjgswRGw9QOOXGIcO3z3KDBY+/fFdX4p8YArK
1FyD4wsvfhpz2o7qJDH8/tPrvubSstHrn8U4t4nBYkU+xrdIg+kLRzq0BPQa42TgAGhxLy4unEho
XkVe8KeUY2kEkqCyQeJhsNB5So1x5iZ5fWATSMTVZyA5tzA8+908iIuQ8lreItxq+ozDDmIiMLpm
2sZglmqUHZaNmY6H2sl1cJzOVYS597Gr8F03eAkOCITTJH7WwoKMEc8Hl9teoi2SFLfq2eEjXi1O
J8W0dzMr3t1oCQN0iwk4I9I/VkGdI1NPd/uOyHIwbUAfjlstg1AhHkE4Q5U4Rq3scbwjaHvb33FO
vB3QoW0ZhHKfJDcGKEF5SspHvIwjH1Y0JALGYHNDQ0mBvz8xJA08QXWVenR5aPG/W2rwFSmEq1I9
1vLvGGN+0WMQpyYqEfF7RlLwG0FXEe5AjvdiJIGTlW6bEi7DLW+yUyx0h8MQw27yE630t2hA4p7o
WMotkdKXWID1pdGuk9WAX8lNrVTSMxR/UshW1zpxFwyaKtKaY8cdPBP1LHXgYloYKg1Cft0RKGSf
K+YCNizmkQF6A4fPpwUM5KuIIpEV/lBeR4pEhB0jij+ICsdRdgCecxGnS3xR8wpLqR8svNuQ4nkM
lkXoAbg70Ai0/5gVc+VmWe4eIZaeLMS20fRAMrKcngTw0JDyl55sdvwFHcuJ3vhnHwKYRAP2Mleg
tTfeetjOiGqzrtpST4hJMsRaxlf/54c6knuIOJxzR+wFZc/nX5mAvJNGXRe8SVng6FveFTkCzzpi
arotvYbdZo62iyegREXCfXSUjudnxszWPyvMLbX+ctpqTl9qoS7RFq6+0W/5BvP58nOtIIUYUq+P
V7SfxBrA1YEcyWG5FzJ8YBppAIL21Jv+ntIQKT0PKhqxDzyY77taY1wdkLw9xfS0INS62ohUq2ck
uoDOQkk6vLbOqM36jiL5WbpGetJtGAOLMFbHwkLQW8A9DcGuiuQ0UKNQkOwbbK5/q5A5YvvhYL5C
EW30XZ6nHX7XU3H7b9kM1m9pNyzLZSPSX7x3y3JQaX4xmG6KgTK2Wyy6AY/DR3ZcO+YzyJIajhg0
/+AGJGoqWxXzLh/ulnyLplSX+c2JeZpK80qOrDWavdjK3y3yo3dLdjSYrTkzvoPzug27sD8PqHlZ
8MbVaE2gqLnG01/Qx+bEGfH3gWdAcduHbCYoNlHkpdB9GBYZZ+ZBl3eQxzVAG9uyVtS3bCg/jn4f
+egiqOJ5QwT7FYNctCvJVvzMAXcaHCkTXG6qt8DgxGZfGqFPpbD3z50gGQ8lmkgT+8gcctVm4Rdd
DEuW0Q8wBgOXv1TBB2mnZrvxI0ynl4d3xGwdgi0gjE+BpmcDMHnBym70uv9taLlkzHlflXqqytu9
isoz8esWSm2upk8h1cwBJmo4cVdBV6bLMXFpgwK/2Qv+LKo//uuHVWIhEe2GOcRPo7MACF2M/0li
MvmNpNto/f4wD4I6VXvr4NZYwQmWGYKUtq6AU7est4d6uKNVMX2k+ByIMNN20PaFpddr+QXVHe7W
goDIqc5Fy/wiFJ2jhW16TlQLr3k6+22HxJwoPafjBb0ZgUXO15NwRt0CDD6dhNlcfBbqtXwP4ziq
seI4JXGcqH21QlHcEWGd1ilDAwixnIjy4Lq/YmWFIX+DnjdBF7bbIByPQYRO2WlH/G43AdUELyDR
dsJETvm50p6Eha2LC4ruCzzeSJ4r08ihOqK2KErNpfl2gV55dIBydCE6d/gi9ITzJmM27rgM7R6m
cuC1MMG05fPm5oP5+CWSxEZD5nmEGMGbrwLYU4OIc+UaPAlhzUNC55eHsveVX5Mcj2a2QX2Jwrd3
r5p5IhDE7GvFEDpQTODpxkLRwIeipMUp5fihNe6NMvBMQuUXWuqSJaMPz5G+M0Vj/v+Vd3c/VoaQ
jWerZG8KroUwkYTjHqDSOeXgWQ/MF6a1BAap/jZTrSB8+NcF8UIS9P/9GVfcwz40mBJk+mCoIKLE
Q4Y10IRjWE5e61KvOTwdL44TmIwN/D2zoAzuXzJzioATGVjnIrxu4pSH6H8rWPr+B23JJERd3RhM
6zx87qcm7Mg56w8EUcJUrLxNqpC/aLK3piA5oirzwysOSN0nvupa2VJTLkOaE8L0ZfEW10dy18ys
/QNxip2bGiWJEYrEWHUK1izfhrV9QINNpXPJw++4TM4RNvLYycKDIvDrahdWKyubwVLu9Gxn+Osu
zZ7iFxXdwqm3BSyFZVffHJRZkKz22goOb+IhfuSY1OLqt7RJFZBLIoiOyu3w8GcnoMbuPax1o4I+
JefjBt3NmPxmOwWE9ttWgrVbXqo8Fy8ORq3/0uCsA4XFo0J/6ZjQDWCapAoG2Uq+KUnGLkbsF9nK
0yNkmLlqAOP6P42tOpucV9lAPh4j6txxifoGsR/uenKsH8Xxtzi7lDB824Y1Ixq06j1sq6id+yHQ
q+AXT/JrYXQqQSNw62erAmgLV27zWC/PKmNGp2ZtQHqLBAhcPqSncFZphsLxXLc3HG2hMkXBFCnV
qDFMcj7GgjITfTKpQnaai2YyCvRNuUz2+F3AC8LtajWnnwtLVV2lUEVW0of6Z8yF/1R5Bf38PETY
ZNZlj1rW08CR8ZemQQtEDiuT8WgmIIXbYrhmTqfZKHqY8L0CWAuCGO8n/N98OepSITcxTKdAMP6K
/aWFmIxZIFHIgnaAHw8EXP2Nl+jDHk1rbVT0uVj5C1z9A3RMrWIRXAkmPe6lWEUTtaQrpZae58RN
I9yIDKyW3xsKdSbRYJG8uYI+wKbY/sSfzf7bbayFrkZXcViiK0q2v+izuILblPYr3v7gxIj2O51z
LTeTs/0BxSHIfzI7jI17Z695DcBZPjxSXYuWueT0JsrB7d0DgLMNcj0hUs0KrE4ihoSoCrh/YgwX
Fepk/TXSqEom7COxKvsxTUBWiIcuDzvnqHJELsd+wXGeWN0TuIQ0isCFWbWuMND+2C41XE7/1oqK
zs11eWf+wLtwqqsGgydJetZxFkKNCEpWnthtQ19+8XZSXHtS4YwgPwe0/2wVO6ekIzGXwkS4ipDz
MqdAFbvYZRuLeTRqUkt2ov7fs8yBjifSsTJS48MdYJPixE80H9pIxD4/9mAIK8jUgfhbgm8Fjvt7
/e345seaf79714PcZsQ+40K3IvXBp+LJQuICmpj2BGjhAPD+VbpK+mmuDe8MtANKQFyPvA0sDi/3
+ivJcz1nytk+ecB8gsub4TUlKYzJ6JnTtIoMNXFGrf1fIX2VdMv+xzGUKLKQ8knovFptuLAK1MOS
9FNh0gQz7Fc/YYGMlYH3WKMJIwSACAgKemN57NojPlFDJNWVE0Z4ugHQvtw8XGYhisURDl6g3VQN
mK+266j02F333ohd+24mMy9H+zOjp74lZ+GAdUqGHU//uiTxfmJPZ6HWvFhLDxGKGlc6Nxb1aN1K
Q6wa9GgGl6fINqvZv4S5eIOpXxQNMlEyK2ji92kl/udN9QxJchiCRSdvxpISYwqGt7H6suqxsIiI
84Xl/1BmRll2CiLnE6XMvhK6D4g0v56Inj8SKeqSuNWupc6/7m+l4lDhqqF/N4zeLzptyhT8vW1n
H23kar6Az/MRW0b/YaLobAwEGBwnUxDPyiokIpQetkUZtQ3ijvRbVzgq5WPLE3ZnTxAWLLD3i5/p
xtHjyNZjoC5camhDDWJyTTmXmhngMGb2ODZVlx6OfsPAV3uSjeZP7owAfl2MKSPR6tWKP0Tuc18e
2KWtExlHbfalYaPxoSNFQUT8Km4pFrz5mgPCoOF8MLRfCz88mUXp8ilPq66Z86iESakbZ5rHUMq3
XOGyN7f48sPkJxuJJ+pz2wXmYJ9UEIqGfG4XejrDzje6ZOrpjrEAEO5y6CYl2nA25SE5RpggEUta
auTCuN+eIyq7Q4ofu6yQ+p4Au1j9+SEd2jGB9Mof5td3hMCN6wCy7TzEjP7GQL6JvNYP4URgMpR4
bVeIrl0A4QFdReB5DKy9KVtFZUXaH8TPhLyyFbQUn+XpZxtkQWOjEp/cq2JupBo07UrMgCx7ABdR
yS6mG9yPlpjq2aeQLFuejfo//l6evS0Qxj0tWbq22jdmJhRwJAq+A9BRvdFqneac18ZKmo5d7e5h
AVKLV2rsNNqBszWDd7CHOqPDD5gdd0UaooaSKavB/QJS2xzbZQxHXn90mCZx9ngyX994+g8pIRSB
FWoeL0CWE+G9DzdWY6lVR/sAjPZhUl+6BmU0cx7C43TpP0lFjOC5EQVDPjqBc6c1rYe2KfL/+OFH
1HS71bbCnNHJJrVYQhfQJpfwvwLQV5ymZZ1P+hW6AKAn2CK1CQhokrsQOeqz+RAAVixTBZl5yfn0
MA2BR+yZB9DZWeVnhPNavyHpeM3DHeJV5bVelJ6xNk6jPI43Ff1Cx2jH1dYOlj2SgNoxVI9tCsdy
kYADlqGsReTAO29GbPwpirRBS8FKkl/yEP3Y7GDyso26/gSmcZFuRTYsFoJk33cORPFisYBrEMyy
am7K/Fdm4+f/m7hWmvjHesMsQ0rNGEZE+1bX6blXytQDWIxdg+/vxGwUgA1Zp772UzdYZZTL/WlD
JtcZwTQz47ufO4ajenWZFkN4Z5i6KPijgcBPBpE8ReSOSnBRBHfP8tYyZDJENb1Q3N3jJXRj1F8B
rFQ9wPp8gIXaHYxcGZEvas50ZJu8f7IqzdVnXfrg/Me+VtCNOi+yPpM1h36c0TEhcpCtzu0rtDmN
H+vDyyVYE5+KeZ4XvPRJoaO0IGtxDjYd+DDM1uFwzNORUCWOg3iAHub1NTlAKq0jPvCGha3ADF05
uZyb3UspDs/QDlt2juPuO2S9E3qBvSJq1ergnxAKSQSrHWZc+MhMMJzFqv+sXZFvroBfrQffCP9g
mME3HLcgAUq5hwO4aDwouAcMho9vmvdLu0txh/A/qijx/WJRAiV5Mm0yKOLFBD3POipFigGK8u0i
gX1GZO7NUxGDLa95+2NTnsMPqdNaQB5qI4spGzffIYALZXVVzUap2syOVDQJBqb3tPsl2tzpQUPO
L2LMGeOKPbbGT4YaM+nuIRtjQDSROv2ZAmd4ga9aksrfQyTFj2HP76qHHmBUXgsXAg33SKf0AABd
1XlULTqZlVKMEYfVUP3tQeqP7HjuciT6ndIkZmDUrdh5pOZN0YHNsDC0pwwxFCG+DWLtwHw2eb8A
38LWgDf8U5IfKT4W5wk9N60efcVsCeh6LjA7Yg0zNuL5t3Ee/QMqh32BfSMUARJnHJlRYKLXDKzh
Jz1ZyY0EJ84g99864p8WSTvZBbvMUkuz6zwHvXp338BZ0FGTnMKSZCoHSNaMHcDASSrghn1z3l25
nHHKCExCMDo2Qn3thmtd6JDnBu0XN+dWxYhrTXqNa7BbRolnYn/zTgfG6v2TetZSksecHCvUcexw
L/1PiDc+dTxWVACZtB8YftIZoPMWc3jVlyObYskwxStjoXf563Q1o6lSni2IsyOjvWdr+ehlv05q
qgpeftotWBRbZjHj1WYhmApHzOXSGOuH1b9cXr0i0FEemYF8GePmtuso0KghDH2uVbWRAO9/lhp4
4fSOLn3IOUqfZsO+wuOB0Ma/Y3TgP3JR3zsrQvwQAzdSQ9VWzORFH3y4i9+rvDtopBLR4By5aWAm
UMj/HgE1qFtnXK4k9i+82LERhMboRuzdWKiM9ws2Uk4jblLPcwJJlJh3f5bFRUxK5hzrZ+Z2YiXG
tIVo5Wok/aMNWwjS3WxNyrC7WGWKDaiODGXKYIQx4dYy/mng2gT8XbDRXwgH3RrgWt3jd0fJ/58F
SvxYvPdGJkZEe6SPuv0wa6RT9C5CPdCfeOgvYverQwnBNChjZhPhub/SaHzYG+dd2ehL34ZZvmh5
QmjCC/aLtvKKku47oQzv0eiqpQ7li7Gekxv1FvNL941kfx/uvbzt6a/VkV40/fQAV5APC1kqtHT9
Za6zwdkJd0oj7E7VUld2jLcoQln/8wR7p53sGEoap69+mYT+Tlh6dFJJ0LQiOI3hDihHHQDQIgvf
CLatprE3wYmYBvBETkrDn4p2mEzHjZ2VkMyzYDeDf+XfXQy64vSolz+V5MTAukilkOHo/lFlw0W6
eSvUMtkeeam1LZdLrmvsjHwK/yhrUS3W5tUWZ10imC7RJJChvfjQcAGyBm7UWWKC+hKUNCV3BirF
jt8otmlTTtZi2qjaNtCmGh3bJnXIy79i0qmPw6EJe5qNqEI+mCiY6HgzLCQSYn30HI32b8Pbk3Uo
C5DDJSt0oTx+8swXpdwzlluTUZdUNsw6tbm+mANLREEtjW4I99FpJrH/89+s5sdINUuJeva8IZGr
m8FzXin7DIKZ82Ue/+qSnc13wM6Yy2c4nEC/NMqoJPD+ZOg+QdVXzhIBbJmWL/5jCfdS31IQ6PKz
jUrwWcXS1ZHOCEdD4+iAXdXiO1sSmTEj2FEdHE5i/Qml6pLjeAynw0RFBxGAujBjnVsH1khy5iUi
Aia/Cu/JaSjI6J7v9r0dxSl2MekaVnCO4oAjvXCyl6L39ZQJ+SycxN1basXV4QzjPg6ARkGEG2KT
LU6NKn8To7OjAYy1Ob7FUhwLIccmiwczpyOWibziuxzJGq0TtwRQbQGWHf5LhxA/ChXJZTJtNgQx
4XImHBfmlIhehnIqMeDW6+hhGP461HvawbS8fkzpJnCQ/GOIxtFjPW+JGnGqGIkZfVAHDkHeWGKE
44SNxg9oKkW7ksrlAXb6fcEJWbCzkV4RNQ2qRCklBWDBFcE5BqV9Isn2xi56weN8M67DfkRp1iZn
v85iPWoS994ayE23GvcfO8BBQ0nOcs4EfMBZTc4yhKXs7AZCjsGwVIi8XlUl3Bt4ErGw8exf71SP
uhpFprq9UDLmRm6FzbmEiePjTHDPjI8wXisoa/qDbINj1ytDvhNQgYcGbPTjIGHJ03YZanRTmkgQ
L7M0ZtoRlES75Whi+VAnwAhd4Gk02hAqKydJIQk0IXUFGuacbeheFcWrdQmo9ILh4Nkz8aG/yPXp
auIVuz+VT2L14GIf2fPu3688d2pIwyOsRZYvwP1mZwf6VfEDwLjCvnGD4ailIs3OFqN9sYfq1iPM
xsh9qznhdqmmU9qSQ8raN9pIj30JjCEv4nhxDcBTPV3zoSbFynnYCwP+6Z5xubqZAGRiNn+Z/8oj
1SahnNxYBjhal3W7gSRTvteT34PP35LIj8N1fe5FhaI5jsRu2pFPVsyvrPrTmmM/Cv+qvtibPDc+
m9qJUslDxkHhoiLi5qiLiuPZ+EPP6GnuRkvd0OcwCK6c5dt3LoBvY9Au7NWL08IR8D9UwC24AadO
888OqeQtzngBWIPldvlCJ7q0SurUSDuzN9CxY1n/XkitkNpEdIaHqCP78Bjh2D06KBxqcVYnR9S7
SyZsdMHmHy4GH8eZ/pXEWJ34bZIvayEKK3miV8OsulayLSiWWh526k7n6ASMd15MloJk3JPZpt9n
JXJiierXvkzBfPdgAtb2wK5gb8U9vh1d1iL0ZcMcCf3daduudaqomjOoXw3xodPDmsYMA8Qgy1Nz
Pk1FfmPM0SwZOSSnCjsNrA3WCw3BX8LvYvigtDSAAY+7L8GXGBzjdJzPcNNai0DkB7SsC2Tznm0R
cDEy+L5Pu1kMlkGdPz2uArfE2DmhPkz3Zo+fvSSWIupv2H2yeklWR3gssP8BXI73D+dykRe1ql5j
207ET6xkrM3D4wUBmRCeKtG1CTNWXR2Tw3VMNGZg/XWqKkgHI3o1icxAeaLb4wA1PobRoo1fNjWH
ACCNvRc6orSY84hVpo2fvb0LUqmK4UbzzSoNoDE4yu7bgaNwkLrX63ABMJ/0UKovVchVce8VPFwU
ebQF6jyF0sGGCw9plUOzz2by9xzgIM/sbRM9nExEbJUG28iAj0gI21T0Nfm5PvxDish6ICDPOnSu
pnE0ziDj3MTvKXD0JsMOSPHS0dlYDu6saB65mad3GtUiASy+c9CMimaV9AyXnXLlqnvx13JFVW0/
tzYmQwBVZfjFcYeqKovYe3bdNCClsRM1TZMh4aac4czS0b2IwNHbPxDw6iADLc6kspsQn0W16dLg
6o7ZVZVW9zvWNIIF5DBRzzWlXnDk/IJOMZ0sctVGLeBa05CWYSuAXdUQixB06VJcaCDiRHxEKWuO
N9gGFq0EaQGW2P4C3JRvA4KNCxHQXTkmjpl16ZJoUCBRk84IEfIBnHaarradR/zBIW1fUmM3bwzq
lcq8ubMhyUgbf2jzYKIRP405jSng2pSZ4LmdQk9Ya2X4ZhF32A54Nwv0LIUl9t+BAbqX7NZXIJfH
j2nzrnPxk9qfgkKxn3lQ8Ye8U++eYw9lvubkamKrVDZK1B9uc7n1OCJbWcpO6eJ81x8ar0AKCMlp
FxoC8oh5P+N7dgXV9TVHozU9M6P0x6KdTUbvPSB1szPcbH5MhU5jZReM29cpKmeJQNd420X8ml0C
SBwnTL42f0Pseb/vpdX/wnh/BmJtLy18H8DZzXg8NnnuDH3r7U0pYFonmEs0ZiDsJIQVaFz0Os+/
WKHhQhvYeWB35y/tBRCZJTAv9ov3C1ASpRml3HTHPeJ7wR484FNu1QO8O+pmpnxeYLGohVvYFYXC
/i3H3mKjylWLsX9Jd3LQFRDa0HSxKDCx4pY0oa/uheEhTs4fc6jJIzACEjv3QfVtaaxOfrMQ3MMh
F17iMDtezvWRsW3X4qMoRwMR+cFnQ28sIHJ5Fx0NKLTwb8e8UGpCyE/QVXZoTFH8cujeCocptcV3
7WM17hks0K4b/om/01hlNFPedQ6TwA2ZUwsxyi5BwCUw4Oz7j5Z8dyEXJ+53/b+CJ03noh85+4XD
Jo9fophUP1fQC6uVLJnUi95Fu/6ZR+iWHoZHzt37byH6MBnLtR7637Yq+BiL3qsIqEz/kkmO2Ns6
xlilr0e3KtWlXeNsSP7Q/iaNaAOkuTaG4kKaTtdafUJEko0DJ5cCMFXZ3VHtFWCOnXN+2evAtanG
/uWE2c9T4ZOk/G/0jvSizbMwtTjv8rJ7+RGFFEkBvr5TbRphrZ+GDLasE70iaXu3tr+sKcYj6kkI
0Z2LtcgUugk6MiEzsT9upoc1vj/o93NKoOrOyO9dy4catQhrXSqsbGEqqVbYi77+2psoxJNK7juf
EA5CL1dzTdO3wXo44IE7t5fBkYUbxtauUOgLM9VY8WbJ0vJhIvjBbFWtErS1bcyMUG0uE+aYF3E4
mLxLZ5pJh9Ub5+eRiIcmnflYn8iHbM0f2zUP1bsuTbV7/isbNOgQzu1Mu6j/B+eOTXTSYiAyznsW
EuTny9aLVA3cSDmmTwc3Cg6UrofRr7tID+xgtnTO2pnQH9lwUBsSkfSWS2JQm8361ZXRMy1U8Rsr
SzQ8WQ6MBi5p73P2LEZu3pKUw/QQKqlSLnoHp4jZuPOeJxnOjaY1/O24fNIgrEPVJswY/JEMpJyh
ACr0uFOMzp4rApMRlQ3hToYEfzYYk6MD26Y04YchM71yDIQYCntDD49AzIxiYq8NBvXdjIeTF+KB
1NdwSnzSdgz1G9/tPnZFXjU+B/XE+5GZotPgIC5ciGhGjrpfcKqZ0zvXqIEQikhBj9nGvtIzSp7K
rAwJh/jK/ArdVR5XTZ0ZRe82CiNzvoWFQv+LA2zsF30362XDQnyPw7JOWdoqZqLHjHuXVI3dgErQ
UegEBgWxrRpF5VwxcuVoVyD/kpRErZA74K4jUUq3VcB1GvAX4ZYN2ZDArkKG+ggzkwTLx0EnxNSq
OpcP9KGCuintKxyoel2W64NMY2AAIZjUnugu4/oMMnjiwDI0lq9h7NCjh5VeWu5uY7x3P0bwQDKT
dEY6gNN6pPjewZVvfgIcFx3nPb1ZWHmVvxtAwwXXLcG74r0gHvEQa2gxo/K3+qRqDYMwH9CMRR39
2RMBY02n21E2Oi5qOi9ejmQ7APhxw0qbtXTpiit347kl1ZKrMPKzCjg/83bXXJ7rJXWbTeLy7Q0b
rw/fT3LfhZCAidvUAanyfQT4LblFK20guOQheYD2c5PSbRFy0lJmjEM1+Fwq0bWydn9j7UPQoZxJ
7+KxJX6M5Rwhsgbo6sYmXK/kUoRsL4y3hbiyF2um7ozXiru9fJ2IFkz61y7wTb/U3rdHtZayQecm
vpUYaUSXzVrJsf6TVr2SJRG9RsrmcU9Zc4187FmSkwF9q5ntcuYCpYZsP9E2yJPBAwMecB0+GSvN
Brq/mS+oIp+cuIVlHypkyPjiOIWdzM2BCxU+1wssz8DEFJn4IpPWonaoZlxAj06MF+CZfujeizf4
hH3J3Csss+BGm4YH8y6Y1FfELCmProbCuAa06kXKxwQEX0p/t3sKM6M1Ai8kdyMxslEQNolg11vr
zmHCPtC59VOtv1fZ79ne5Wxi/z6XIiAspH0/DJlhCJqGXFJ3Sk7w/qbpa6igd9WY0Kx8ml8V05dy
mqV2kvzGEX6cHPbdNO4oG30m6avAeNghU9QMDEYELLvR4Bl9VztKqpDfB7w4Rf9irk16CYcu+WGX
R+oIL+ynQmriN6qndgiFN9DeO0gI8vYmMe513yg6iZ/WOgRtLZbTfTM5loUHre2A5eJVRfhnXhla
9JfwVuWn10nK7j3A/GBQP7Rh2WKPYdleM8Km0z6TvB54hIWogf9hBkTXiOJ0W/bvH4gUJwJ0bVyz
lYkIRDftvoWVuZkr3fgp2RaIqGCeBHa6baHoEii+/V5TjHoEkd7Xzl9+PNMma0cH5IbQ49oI0EUA
EnRsPUn950XhQJ6vZOLLikSs+IlQkZFP1lGCgUS/CNPanJEp0ZnT30ilwBg39Hmxf05sQnttikxV
VbNIWiGw8MpSpnBGPwdM3+gWNNLY0LTrtBQhsqrVt3b8fHhvwRnAr/xdhJVQ179nq0f9zWkZCJ1b
duWTwfKrNvd/8uePfR2Wo3yfcyxuJaUc48+vaNRuc6E+Yuaj5BIYhBcAbddh5okLoYzNdt6WwVbN
HGS6Jlmnj7aoTttCmOC7JTyaCJKDgPHFrxMADoKQ+urfouCevNpbzY+r5rHv1tZkGWGw0kYBmRB2
vefRESntL9nPaKBlLOI/df+mHzph3hk0Eruhyap/Q4QTKpSgLUIuyV51tQK+eUwjPkgZM5MSkluW
Ypp3uVVfiTC5vchAJ7GMC9hyJxd1WCE5raeTZx/RxU+/6jLfpj6+3UFhwNhh2/XnBDIAc9rrEkzV
kgZg0KoMBkOB6oPyGNcLsZg2tiV/q4AeFFokSjfyy7qj3bi7D+dcVvwXO1wr9WIJvfLYVt4vmK4x
FmTqYgnBtYu9JC6CDEuUKTxvoBT91Whc+12bzEso0MNqyyN+8rwYeRWraFaYx6FPnfpxENx2b0PP
T5iTgMctOhIlVNtbxwFAE3B0RfVDs3zh5bz08ia824Qm1rHJcZ1n6isEalV+kVcyHUNbhIkeYEfS
tERQWt4XUO9NMSdeE6tE1nK+SsdbOBGGiQWfha/ogkF0F0BlCR4t9InmOkdFwcLgcV879us7ojeq
rtFzgHee5jVxIVG5sBJ7Ig3HytFurQD0aJEcm6iZt5ayja3zuaZvQwhg1pKwGeUSVVt25aVmC/vx
EwAv35EIvER93jWHtF71Nk9ydxvw4W7zSOW6QQMp2arlwH3E7d92x7PsnGQZTjI82qr9KtppBlQF
dfTgUXLsNIP0Pw+4nE0wg02p3vwDVuFuXuwhT9FQXE0U/L2hR4p3MBNQDIUUhLj36+Smam7BoZfm
NE/2mHHE1QkLnEJv1eHLjz7EJBD1eu5Y8HWez6OEVkcSAge4eJwi60emPer82cAUaHNot5Di7NJa
t9K+UtJNftRlvG7F36Y+nlMs7yqxIInn+647WzL7LoRWeHzqbwo7jwsM9N7pJRB+pviL0BYVg5Fk
VobS+/T+CaLEwramzJ8Td5VtIfhoumktfIYcWuNlpWrV0qFw2UitwRtarf4yZNRI9xbdqNRct6+I
a7ZFvqhbNS+1QEmLk1f8nrV7M6iIU4U0jEv77fSx5GTCaW8wjr3Yv9Y5hKqd3BSx09LSQt6nvniC
Dsu9Ab0IaFrnMhnkyyt8Z/ow/J+NtTaDAScr6T26AjiZvN26zwRrnOGJRNzLiEtNXNXic/fAE585
ER2NBcw0Jx02HVBvOowjN554O9/jIE52EwehEbiVG62Cukw4XMSGCa3zkfsJK4WWRbxffZnJJabv
/gc8A91yPZpMM+VeVo+B+jdsQc2xiOKz2SbiLv7Tz9q6c8IuUrycDwiVIfxBwtt2ZzGhRlznKAnq
1+nz9VB5Rb/1jut2evSN2Z9XNNdTgvtXBzZ2v0fEeHWYPyH8ygDbWGXUS8fG7075FlQttzbg5+RA
/Z1xdMtd3+LhPgZtjy/6mKTmIkCQ+YhoAyet2hTxLu9CTx1L71IuQ4ITtDdGecVq+EfWqJqi/7EU
uy+kht1W4f98+HdyAt7R9Be+uOJMA0aKxj/XONAOCVavUFE9Uo84t7MlHq2b144aazbFSjm+qkee
wxdKhAn8FXQkwzsSZorcgTlCXrkGd7v2u2KRe+9Hc/yZXZ3e7Oc3mqpANOmKvr5+xj4rLQ6yf4+h
7Ptza7LlmW9ZsTHB7LeCMJ7BTYt/gvfwOSHfhohMBaquaq8xIzvuHsE+6WfPayJRgzDZKj1D+GEB
bncrFuohXpdm4MYvHbW/XiGd4SAUO7akQd0WudHR0FVtlP8wMPsG/Q3KiZmgx4ExoP9wcfHaC7No
Mo2nvIQ0puJqwF773tEVskSzIsmgmqZbm8Bsri33/lbqL9ibWMwT1cq7b2TRzFJfkFRk9S3WxIer
jHTNWyaPfTFNWMlUmYu4ZSfKcOZkdUOOObagzsF1svadWzFMv8YpvYMWQyzmzDus032GMRyhocmT
wFy8TkbPmD8YuCiO4xe3aSq6cfg1jWgMZgbg+rfuIRQKUXZCNgjseuGdHHVVRTrN/fMmlE+eBY6B
KB1mzwWHQonUwjduWJhLmt6FWJCErcnc+fd42hvKdFzKq87i4lXXc8fAiyM0d04zcCXtsmcjBprd
K95w8ZU12AyMwRuUz2RQ5v26/POaZoiJ5gmC3ivHMJBhy12RzjBCcKu8nU0Irz1P4H3zUBL/86fQ
cLuWzMD4QdoyNXl9VooRQi+REBFfVI3+l9l4Cp6W/vwjzVxwCMP7m20iS1FcBz39gl3Q+lMzOVp1
q9pmnC3xX7bBiPYMaSXy2Tb/y57tZaa+wdFvWTiaY0mxjGC5NqOdW1jiNFMKbT7VkhZ/qNyn2xyR
nDc+Gx1a7RaCKJ+kq8VL9LeMh4zT/l4XkHNCZGSeMhx0jx+IXfw3ODJLyInrMa+oZ1QIzERWGWT6
4F2CvfIW37xcmTzcY45dimpJv+u6lhDOkLHzRxlH6cXLfRoZSUbIiNQtvVGXMjD0JkHdzGlqjnbV
uKAcFeApQXkKrt54Jk7iVWrkXN5x7dXl2FszmGABQNLdyW2udVl8CtkUpBz6heWYPW4VqowTjqOp
uASHzTRXXB1xTU7Q3hzSTjdz1SpSsYfMkMLW3Cm4BRgVWLv1OWzjpL61v2j4a6aCFLXaaOI7sTqr
yuZA5HFUamZycb6NyPv6FKzJEcmVsfm0WR2tyPQngNn2wRFXPqXP6kDM2e/T30FtKMxoh52szpI9
yZ4D57bP2Z8ErtLwprGJxLoHNYITKU4zduwFaed50WU/WHNYvY372MSO9BfSEidI2e/tarAKSDsu
UyNcToBjEM18tm7iMvVCN9zMANs2cFbxLAxs1p6xONGEzOLgcJmmsLrtSZKtbl206rMW+Xep+P8t
MCotjCBXITosWOYbhJaBITJWcf03NPzQvzKSH7f+gHKUfOJkiLMZPsP0SMOIcOtRQnsSMR8IWWde
nPnPg9IIMpJTsg+//Qt5mV09yuZvqQjAJ50W2PqvEPnUovIGUndMZ/rcDPy2HQgaDaoRiihEUGkB
TBClyB75JhXKb5XK+Va430H73o/EJAevDrrr7kkZHQIxb8GrQD/wb6dXuMrET+7b/cQcufBIxmsA
SWBj5Yi+x+4XS3H7Cq0y+r5xtzzy0lx942IHPqQoEnkPYwHloMP/BzRNrPIq9b8Jz4sJauWXJ3cm
chChj2NAR0S9PszMqOh63SwjvDLfNRJiKUuqEKBTQVyzLu7MOFpjTef7wFOdjWujAQbc3cGULnf5
7JFLv460Frd/o7oHDkB2zif49T2UbDzW5PDfGAJ6wi9SiGOtrLpIxwA3uDl4IIDo25w9yLq7GjCQ
Fs4k6ekGWpnmpIUg+FSAvlXDxYqkn72RVnYupOmaQVWYxLlX0vCEK/ejW+tkHiK82zns4028k9qm
/P25tVJ/RnCCP6pRdEx6p4W0+alPwGUpcTA4em1/stxcVffhJ5Hzd+UReA/UPMoxzEI3H926CedT
kuW1JmuTdKR8P0ChqSqFXINQeQhLg3KVpgZtskQec0jdDNO6cFiuneVNXZIF7fO2/Mwy/kG6b/qX
A2L6+hw43tVpU+Wfv3d+SxeIvjU07I/YvxMFC9VFeCv3goYD4vBIxca2bfrH9hHSUenKUoNpeeN6
y0bJwqdy+GN5m5E4j+osMumfK2VVP34wnCh9h6rBHZijcRZmoTwpWcM+OlKP13MzIq/eR8qNmgM2
cqs/dUFgrM61OPugbaNcBJOdziGnJ/ywC19rZ4dVryDOvVLJrEWnObkR6aaBBCrYuGvl8YBDgbD6
XGBGfqj9PvpdapVld4FQ4hjja5xEUG2je4PJgZ2N3lOztG2dwn3Jv9sp+BRNas1Wn2KYgRVg3wUF
c4RaJ9B6ftPyBY7u919UOTzAD/RxX2lWUPhL+GBSfcqq1Q9YX5pcv4WmyuLa0/SCdjuS6+kw/T/C
JJih7XrGKHchOpos1QRE2hNvBdYiPMYcC49xD2MIMqyFjwyNljZZ3mdhDmLa3YPbiY8zewTRmRSZ
AS59Fd8+eEeGAtKUiOxGAGffgbA63WlT/TO7ptHCu4hKd114QLJIgCDf6hBOCbocNdqBgjSxxe/9
JTk57dJ3Hk/eQDZZ6C5aofvaw/1ejJpd0mOby0yDFZ2GYg4qIPC9iTgwFGnXIT56ImGoGaTi18VJ
ByoHBpho7KfIzHxi0ls31B4MiBLHVF4cZ40Fy9rPWgasxyU5WgVHscQD7m6tfnk5BsUkXPRHYE73
zYCdAzDG7+0LWAhXTqQZEYqsm9z+MAIqhOmTIEv9Cdfm4QEx28UR5QRYWjbvxeb5bkacvNiqDXOU
JGWN4DVTS4K+AbjRiI4BXEKYAEqGmTLlEcmU7yJpEeArt7ZBcIiI5jEzhyfsxeG0sJ3J+SFGGtX3
qdI9IwN/D3b98tI0yOqurlKsk7ZNo4eoKEe72pX4vSJ+bhh98VR0+Q+Y2gHPv0bhM+UAxGvIzPN5
RvGR7Y1mcCqlzLlzMfhgc7/nS7lb/EYU1x19ERQvh4uVTOgab/RF9Vr3/4jyzpw7hGTyY3pQmoZ6
l2V0H66WLLA2uB2eIOjZ2wAice4fQ3Qe7APdsPr2tLZKh601TQYtMg0NnixLXmekI/m9OnAbG4vl
FF0OMLb05Z4V3kySPLX//WCj4VjO+xmdCtfbbn7KTsQ7Bi6GfwiUYLnj1PqAt9P8OCb4S2Q9Fqgr
+IiNLbhcqF2qk7Z/yw28jJUe6lim0LTdFJnThoKTB1uZ/pAhw8Zxeu2eKj8ZC76jKfQ48201RAcj
G8fd7hc3V//vhCYpPWFOUtZZdtZuAfkHvMc81Hv2GIzHLcBzUgSnmdW8t4V0xlOpGoxzUuvorpHp
ktTY/6vpvbwchbpMn+fRFHoKnIY9vacMO/jAMkfeszWvm8djW4Paq+VGJdaNKtGGlKaGxDu3huqN
KNVbXabKfuqoSf8bpkMD50jRwfV6/L7RK8rGhi7XUKg07wma9MlM+BTQDY/47YNG8RzxfRs48el3
Q7wHeX9bnR9K557qIXFjLL7dURwB5zPHeJL+zkGIuHxS3eY6mTs/u82C524J6qf7OEcMOlXQ7qNG
SOf8c/RADUutmHtI6wqERV6oeeTLpJ3Ktv6sOKP/5NIrR2wbud3YACKd+tnZw/6K6fAY0Q8FXc5N
EfbujWLz0E3ewq/B4VDqjEvUKFFnGTgQSRphjzP4iI9knenJDpuD5W1qS1n4eTM3lIWS6Feh6tKk
zJBzd535fP1udt80pulgU8Y9R3s6cDWrn+9s+HlyzR12HtUZuakGZLtIqfae0KaHxuU9XByjS/8U
i3sZxV5HZk64+5wh4lvu52A6KncBHl/F3udBAkpzJ1qTfJ5NGe9/EtvTeXx84UiSjrYLfpbKTMhm
T2XhFGIk1Sk9tNFouzr/nOaE8oEs6noQ93tLFkE7Y4yc/aKyEO7HzkXjC2OjKe4KYrIYWbDGEk7B
Dze6FBv0IhXdoxuf7h8gtrAvkAWsI1eMMQhrDx5hHJEu3gzVvqO4ZpgwV71Qb6knXJhuYmRP8CJU
7J/IkjJeBOCHPo0/RufK/WzugiK1U9oIo5c1TnmaRvk5mNqKuvcIUFAm6DzS8TYsw21+Fq6cMvRN
F+NeOgJ+mjD8f4fr2TnI3Y9vZVqmO0Z5kjvrdgkEzjc0lIvoj6WcPig8AmsagYRBMNNvAaqv86Fz
699hEK8HMbKkKQtBJPVzys4Ms0m7XkETqUfkVQmBTrGnashYEcb/Jpxe16qruATbtdyE3Ypunujf
R9DDEsFY0W8K7jJiL4nDdWYysuQ305UfTOQDwaWdpnqyNM15x2qtP0c7uW34lByAFB1DYPe8iDzr
EI5iBBrm/ddUZ/Wns49UnTYMpHtOjcjJ0dMq5PTeCzohQEPXpfvFPPUYZHBNB39Ao9eFKG+t972E
4ueQ573LKcE6sIyl7fuTISkn8LNPQdZN6D2tvHUKcrL8XRzcQnTfH6c62YJiO4mffFzAkc+8Ltlz
qeFlpKzn/gnGKKD5ZRVLoOkGVi9T+xZQxP/By3l9kbNdIPta2A6zKf5q76juZ3aFnnE23vqJ9T+E
02aO0oelWBssgNmU50BrAugulg1mdoIUi4GI63/jsvYSKpycNdKITwoAybh/XrSEdhra5hKmFNtU
VoAl6pHc0XRQarLG/gFX0NRYhrWNG+QCzl3p8tlXWrUPvHOQtxRb36y7PdbaA/AaZjbYIV2k7wPJ
cOdVaNNbrnAz6Ea1kwQpyMYkCFBbV0U19PfjiVI/R0+gu7cB0Q6/ehW1KMtZhMkTBoiTyqBiBSED
6qqokoaTF7+l4C31ATWAViJn9Lg3pTvlvAjlviEnh2R9kBzG5KxS64Y+lIotjTiWB8aUCtOIrBm7
xy1uyljn9H4dV684Fdts8m6SNMXgjbxlkUka8vb+ljgozR6tgM9WaHYthOkuDIlkN8l+KpsSBaka
MjgVsoCgF69caSSmU1OdzRklDS9680v07Md4/j1ToB3BH8ZlrUEjDakJzUwFdNfxnxWM+eMF3uJd
aG6cbNV1TcUjyD87Smz6ONfs+Ep85I7z+o9rneUJmDBOjac8bO5jQj8gtvVOPDzgP54fjjK+9R1T
nG8vYmm/simAvw//1Q3OCZAZB7N+/WErYtZwvUtXMRQahUJtnZQhbsxMsDY/O3DGekM4tVNPk8yD
ja/fyZwC8E337Av0yW0DuJg3joYrpmC0RU3rlcuy07BhTl2o0OERksljFcmYE/8HpdKf7kAjh+W/
+Pb2m1RA5pI91uPA2XehPUPIvDUzFOB4YMa8iPo93RTaF635CdgwTUX9HOAap2UhV7QAlb4j4Eru
++Q8cQpAwmZg1dtSqkdDDsWgRndazHCIGTChFIyYTQE2jBQ/qrtNY5AKsjaqVeoLobGXxmxB0/J4
N7N+OqefujMoBF519o3lsgiC8SbtrHwQ+be1BqtFY/Mu/PigTwdUWCOohg5CegJhltATKoyH2Cp0
td0cRt6NAl8ffMr+zgBEP6XfdHaT2kVvTx/xNDsyFiH8Lic2ypsEWi8WiXBUx4FWLbftRLr8xufw
CSY66wJei8PMwsjuCgHiNs201WE5D21+ZquzSowEjLK71s3Xj7XaGSUwMe0In8ldX44o+xug8Qfs
A3E4LfncDLKIwBq561JyX3SyLMgTJCM1inBjHSQxVRKVP73g0ZKGOHDSUJFAYTiafnT2B7i34oLO
HjueJigwYR2E4ntmbsp5UuuNnqO4GDnq74SUJMaQDXT/kdygOdY1thBa+xHEaNtyL7q1Z+W8VULm
BG4sJi+ASPMAUM4yrNcUA0MMwUifl7WY8RTZMiSIpRWlAcvF4/pRSeaB7lb4NSfc7rvZHVVINyxa
6LRQHWpFGjl2Xlx6ue8vgMsCm4//lke2ypuumWzk9aTOgHQav/pbsGh7nvqtPbC6B/L1ecJ8NHkS
dxaAXyQ1TSR036YVUz2GmUCyRiWooIsXWjiRxtmhX5ffnSx56ym1vVWaN9XZDLTIawwMxsHnSsu+
VQqng6jEJjvJPDNxk9Kw3M+BK0nQ0TvN8JseJPWf/nNq4Oum2gYZcL4B6tetBm6IKZWl8Si3z0IO
28sYiWlPdvcC09gJGq0oRwRW5WD9d4JiYKaB/+75KILsaza+d5z8Bg+kINeGeVx2M8/P4lE2sJjv
A7BJfO6xDF8sd72wCqjNsDBaLEd0KT3pHTqcQZVGPs/kHxDhUcmf66M6x2OH/1To0KzD+dHfSmCl
+HYAgMmoAt/5iVPADExJA8T4GWqy6HgUzZGNuWz2iPMT68Y7Gxp8WkQVI7De4t2n6Y+MXZYIdxS6
fAH/gvGnbsUCau++xWq794ebbifHF78Nfv4cRIszHUdy4zwc+yYCbXOw8h4IuH3UPi1vB+mMIxKN
m9EYl92hs18dwWLo7ryc9k3tH8d65Ksxpi3STu8j2aZW9XvqTQsm7WAYOL8gQm1tXc0VMzBYBNMQ
xtzOSFQ6CbPvVP5PRH+siPku4aUuZxdPH1OOxkh97rLHliV54UtdiL2tefe263sRT9JAPWqNew3b
84292QFW5N37HCIVWjbeAnFlnTG1qm1H3F2qOpLJncVQq5OILVCnMZp1zOzWOEDq2yFQPgLUlwGF
Buy+fWhfIOscZ4YZ3pAVxprdbJL1/NkJsMPlCl3z4brLB9n0W2EP1VnlqtcvreVu4m12Q1DYWWqK
1P1Eqd7+CqLSimHWYEiRC+cS9lpBgO7ECEpBXA7A22b6Ycb6hEthG1ee2Jxhc/xAWuCZvfb1ZlQG
0yJu93n7r720IEIjGK9s1w/XV6+M13S3fIB6HxjY/B9JPTH3SsHVVwAWpHOB9uURSBHa2bbXXSN/
Oy3v/8MJhVSfWxOJJ5XdqWxMT0ZvlZ/Iwj3uUiVUZunX8Rivf8ZSz9HKBYwNGN9RMaM8fek/3DTH
e+cxVQLK6ywovGtiWailqGFLnIqv+mHYm8e72lhaXJLLE2zln0nNFypQ792hRBpMd+5rpRRxxP5f
U9WIyNVLswz6rlz3pzH7akH8zXoNlkmb0lChseGmuiUsa6P/CGgyWi98nzKoaK5E5NdShS6vGoN8
23J2cb/kLhHFlinAFbAtrKewWRo8miQpK6yTnLLPGRFhXkrSP5hbOxbadT6HYtwsU2SIYQwuAiaR
1FLYUrLld6AYd8Zc5wvknQsdPiSEle5znZc0JbqdtiA0tYVUH3dTAxGkhL45d9M85eqxXuC7uqOA
/Em38LTlGKgCMN3bLoovXV4V5RSmcXgJ7olBVy/alpL//Rx6ECbDf0O2H7SLB21j1CEmwnCnm/a9
cBeGTJZR/wmhg/k2l9cCVk6D+GglE+i5cbQXiSZs6hefEdsZ6+2tpTUr4HaGmHZ2LdNhH374nLv6
MJfbBeCCo30IDRvkQDiH3SuJ8Xyn+/WbV0/lgHkvO8sqOMWVZvbQiAS5f/FO3QKytxWpHfTNeO25
ehdw6dK/9p3z2XMWlv8kMbPbtWeMF5W1fbUVuT3QE1dnzpBBy8TgQnR4v6wfZTaUxLTIZ2+KqxIw
D5BJ19ZXNjdVujI3yl0Scj2xxBtbTv2RCzs0jhTBQPd/HQbXdvhDpgJ5XftrA4XCfqfII6bc7yqr
gIyMc0RbyVnEA9YVzibEFLfnDrfMZJqC4eX2kAzqjkC8w6mOyQxPpotA874Qb0N17q1aF2xB1xdU
PH6G3fc9cjP05cM2fiMrPVyaWQVNmzj2RavwTkL0BHIO3nQrrPiv8R6QUqF3QG8vpjs6fKt9Ll97
SMvSfws91OOgGPg2mPbW5oAVGv+3tB8j8mUfd8Cx+vuaiAX+44/+JgaY/fTSdtBUzoTKtf+ayrn+
aKWlZku6yaBExKnkwKVD8+hnpxd64rI2XG58SaweA2BcKjLAxpiysB4V6mEm2gyPrWWJzLyRlp3Z
FZOdx0CBy/Mv+6vYl9OHujR4dQ6jBGj7aMkeyfEJkTWLhVkcOW5JFbBsJ9idJYn3sO0hv38CzY2/
hhbaGOB2Q7Fhm3yEPJLMCxccgac6fjTCr20w8tlsN/Gfo0yuHwsdeLgQZJORdN2AqsljYwekVKDv
iCL7YT7d/Vx+CABkOLZQ6+QRE3/wZnGTrdDYB2/frRSGhpDyrBZBMAPhNXElhIQRaoaGtX1LaNxW
EZA/V3juOc2U4O3EugCxBVDEiimRw9N4XAqbSzf4T+DQbP/S7AuSVgcgM1s24GluwxgFiTHTmLbA
LV2pa+S7SET6cBMJ27JeWHUwXWdn2FO/Msl4ySq0o8NwDvVomEBdHkhXh80/Zzo0eMHmvAE2e+WV
waB2eOljlzJMRTX+KnuMdaIaqS6gzKioXj1XXeRE/cgwIdRu47cONYtNIPpN1LyQJGdymI7NePTM
5IESMWtNWpU9NlLTXIioO7gw/m7sr5rG25ARJRBP97VZaWkOZXF54B810ccvmF6Of2nKkUnIxSF0
+TlK2p8ljLzIHHMEllm10DpBlZnfnZ5LAd56nSJklF5EJ9WJTF6dPwY1cV/fK8b0sMNnPt7/2MuV
OhxaGek/owYXM8xuEUlwUffEkRNVf+W25fWLHRKWjWWHiF1pZVg87fMhjuexHbfEph7jKBj1z1ZH
P+0tibvOby47mssRDSJwEnLaEz7FuFd+q0u/QgpNmhkCqhPBWMJ1hpodwzBFOzwJIXYCPc5mXhCi
YYmdtYPg7D0wnZv0aHgD12cA/YwWK6IWQNmEnLhbqk1XnZ/ZYQZcCcu8dHINj1KrMyxyiI+WVeJN
K8V5pNDzuAzsMk+fmmhHsRtXzO768VQhWpts4T/RkS0FYc3Ay0932lntXeldSeo54qyemLr9PqnH
OvfpArRReRyJ0brb0xxzVOY4dchg5AuzHHqttq0KVhGiWhAT7BQ/m86pc8XLsQFfFrjHrJPtXyg3
f16TLkUU2KIhRDGPbGLAPv4M+wK2KCpymqAdflZIsQ3arrziqMbNQMWlLfLYa83FmqrG9F9lUwK+
yNzEjqDX9+KRcXo5GE9rFaG9G6Pfx8OKsaQGePS226J/dJ/qSCSkBRfUdFmoFVZcj4BmIhsCaRIH
8ICI7gwKTxZe7SQHqh2T/uo8lHdeyLyGke02Rr20QOZkUH/f0W9/sa1VJv9ox2GBjZgY+Ud5zH88
logFCam9hgYD85FyzD3i2pKLsWyZ5dIASpOMJjWtdfRDExPs2bEVb4Pz/A/n8xDIT5At+eFGxVsl
CXHxztAOss2xmUUf4i7TTNe/He++CsNQCGF7CY6sHEv0HhZg6xV6ZPJu4wOVf0qYgwIs7rJC9BAE
xzxkaOkeWuqhs+fR+LZvAua0JKENmE9bmqLg4eXUbI/jaiCLtS/taRRhw0hijLsy029TARGip7k/
VSz+qeWcH1a8QAVjLH3JL8hITOfwAWXSXAs+8wR27mWGCc+3m+sCvgTLnCLw92O+BCfA3rkzE+XI
C9Je2wOSZGcCCx5KYdgpGg/UAUy3ww//DTiWNaVa+ld17HIQr5x+LH0ziuHEL/PSbCkozpc9t7CF
Jd4djtOJs1Y3ZYOG9YwI2JhEiT6Bc08H5fE/32NXvn6KNljc5ZjlOIhnBIo8Wr1QJDro0sdfFGQo
oISMFgOj1YsILUYMR9KtvCP7tUOROmf2rK68Y4AwjLbqMY35Xtkz+h1c6zDJ50K5X6GCGae6Fx8W
Zh930w0Y9iJrAhM6m+RDggerMyKdzuwCExxW2j6fphyErJyFAQ4tZtShgEBxKHfBbzDhk30H41qC
IFHYkLzUUhYi7N9YVS/sa+RzN2iMFpLRmK1KeaOhnShRC110baUJ98BX+0qZmCvpI9K51vgzUmME
BB+fOOlZ7WsH6VW66n+qsaV1OPrLmiLKOdMIwfc0eqG6GsuYytMVDayiuYXu+/gzNNz2iDLOeb4J
8eQH9emrrluIYjOOsO2QjeIcHercn34AheNY8STfwYtMOYtZ/9+PkSHwtF1tPKmSLOMRahdh5hTY
hl8vz7txHi4VtjSP47bUmu6ejX50MKyMLWymW2S4lQiNOZyl20KAX37cq7mSoWodNSNuHNsVbxxb
HHj08twKybP6LJtbIbCPVxTynxXRv/hlBKtSvv+FN2mIZT8dLwiwGHECxWCY9uHYn4BIGTUTE/v5
gqBjq0r+xb4qpOtEK2a9RAhQnu7Woh6lFwuzS0m3fckwzUusAdpwoxTa0rtURX3vz1jcHLOdgeeH
SIEMKqAsKiNRfJJ8yGkJD8oO7W9adqfNhHMlZYOatctliJq1RBJnstMp+6GBRBqzlFgdeWGKC5TI
KjOAleN+BXtfbTltAcs9aMYVnkkwGlLMgXQ8TlPyCF1D+EApzez9+VyxJxjZCqDp+SA8sDYL0a1e
Zx5K+zWJuiXRSS3DqDxSkjoigndds7XnQnYOwq3v9IeW1evwISBpiDMIo/VmAXOGkVl4Hb834Fj3
OSDo0nAXu1K92JAcpAXrXCeko3BhQOmMKR/cVNaWTmRtAKjZhcDKWURJdK/RCs9YONQs3RWvQ0fH
v5WMQDWjLARw+CjZErdjlBjcCYX7Bn/C8vRLQsfsqwlOZoxd8n0bP6eiQqGrBjN2f/CDrA7pVOm6
b84znPemqVhlFvWhAlGnr0soLeYPVGnpb0R6q7UO6346OFiT1tMGWeBI2LNIMTI+nk/PeH6DlI43
Zovxgp0kHHI5gwnbQfn3SRWZB81zzwVdG9FOW8AN95OZ/itpkESkf5Prc29zJvAEQP6N4G6xAHr7
GsG41LrvJcCR3YCcfTbnXkhNHYoh3tWavAuFUR71dEYEyh8gBA/f2VPpBuOFiXW1Ouhj2uyIpzcg
26dATnoZX5n7snMI4jEX7ks6GWWjejzr+KIEkydX//sFu5J6zDE13bcc+ufQ09VajcndwUwOqOgU
GK0WOIOGT6/gfB1U2wJHZw2x8mjEUOnjPMYsYu/JFBxTxU1PPmbejYaUnZDo2QB5jE3fMkC67nHl
pYmM/zTmjx0E20wVSJrq9MB8Vtku9IkJH3nvwC54kOrs0yto5vT3T5Ji7SJ69fgmjSVKV2binHxU
UwQ4c9REiPkeEJ9Lsvj+w0Z+r8w5RTQn7EXdqelx57xJug9kMdUwx9glpPoq4VcBbpkGngGG4I04
IWNTDCrGXPtV4AT7jPQvoPIqdnIzAJ8hBAgyh3GWxbuc092uUHeV3P0XF9H0iCVMLtu3wskHu1Ov
zO6RsDOMb9PUcjXZaITq59Lsgrb6Msi4yhk6csU2tX4uc0plJAOokxLn9LlgGyoywWFHoFi0GGWv
mq0nX6PSIs70IPMU2g6AHGoCiMfQ10UVk6Lmj+X7wcyB+uPffhe5qPZblWrDHfgzoxEYEdyF+jNz
d8Jxkv1xPF+2VKGUR4/Ixu/9zYU2AVLe6qkN31mZGvgcvyy68M6KMM8ybIEGYcidffsl3gXUSdQN
boUsQ/5RGEVRPe4Q2I0aHrjXDDpzqNDqvnrvhC02aDXLeeyMy1Ayvy4/oRopUFVO4tG6bJ2uzh1E
0xBkvH6LMSBVcTJZShzKIB9lgP4DsOH/5HVq0yOtCu5HzzWOdl5sC+MR89HD2rycx7P+qkKfQhLE
75s9LpRWuDnyZsE3LKPDpW4MUfmsxNkd5AW8YamSF4ocWwj57XG7gkwTJSar4T+u22SokAuefjFf
YzWzCH3/NHnKB07qHxcp8Laac8UUq+9Nmfwmfr1RLlCW+r4zL7ZB/j6z3LJR2DIe1YTHpJ1u07e9
70LE5SjfbaZFiBy5HVA4mvGROazibGpYoMVNGXUbMLMuK6zLGSnJzM9ldAR51nVWuG94Ef03ka79
LyyAP6p78bye0gt8RE1bLlGuP8pfUgVUdLb+YolVsFteaNLAcvDaEQ1U88Kp2GoDKZSoTFWnP6io
WQ6ONrHeHXWOr9NQCElHmfqrhoelQOozUYovfDkwg7pv17YZ3MSTrx/ezII+c7pHr5yZ7PqrJZJR
pm/A5YAaaNhQLBm3eE8X08+afN63RFwII1BA6zSE8o5miOQdgS6ty9RA3VpbwzDV11r1O0CsP1cI
LQr1JCwMo96mAlm6i5P1wGDtZvRFAjHuQaodyuykVaZ1LBXPrVgNf93YB2FJf3MxL/LEOqzB9DYx
NbxrmFI62Te5YwBTO43p93clo2TV2W6gBFVzBDrRHmQyZLKIIGkkQGjhvPckKHFgZzWx2sQpyRtZ
DR9gbiAJzeOJW0QeMroa9PMYsiNeDVgJFZKlxZzFboWj4mlaasuoi5dqK8GITgffaG5K4yxY7+/M
BdwNTPgeGzZTy0ylFS/Lbsby1VHkiq5xtzzHvRJquNye6bUiiYO9KKTHJWUZu64iK5o3z7OjnT+L
W7x6tBoABh6TRAHnrc3Pa1+kCp8JrkRmHnFIv1h1Y/5qvhs5HdAYTVzXqqw39ys676NWmkKxyEbZ
N8M+Z0s3mhZzecLmMylmfjOoKkbL5eyMoF7CX5ZA917RiL+ehaX6cZhNUuZu+71AuFT6d5lNPSOY
AylU/ljr9rejxGgAbW+H/DQOlgDiQQx9NBtF6ELVOQAlKWlFK/6zbYPSlOjrTwZss5O4TD9QzGNe
xE1B9GZqxnZVrJFFpPV41VFI15eDc8aG3vu8kV/aAb2kmXBR16NBzeh+pk+ggWWmEJqtH9JJnDwB
ViHBaurzcKbiLNRk58YFtjoj7F79gt4k3SO1tu7MnJq1ASI0W6NuTSJ87br6QwgkRKkFtHTVOnWk
Q1Vf0pCRg5oZV/4MIyr9Gm29Qmec9jP73chFN8nxjPNZgItBC65d6SKzmgsqpjQdjHDXeStcjdUx
R44bjtns8Ahk1rZX3kONrKKVggeCoRUby4mZOo86FxNenKFfIZ2ZXu7M4kFsUariAQXgBl3rVBm6
riD4LT5DMkTiBMu9wLE2JGpmlbWo2S4WVXLrVF8RyYvAqw6lFcCT7DZn7scNy10acLO4XrVeTqgI
WG5ETJpDugrUEXY16mMGKVsQOd24WxN7r9F/Ei0qWHVfH/z7pMVqedSBM2JsZUnTs1Chkfp4ArVk
d+OkzB5t8m6QoySuvBie0WIht9zA8X9FMkIBUwqna2R+hFeEnc07xJAbLRkpngJJyeT5h+vJD7G4
1DAPTdf7jhXIS8a5gkVVdXa6tTLzpObenLtb9FzNiEwZII1TGD9PmxmVxTvrErjSvlJqijD3Xbb/
riZYIWk6ex7lI9ALTUHpnJcKMOVWkvoDT5mfvXNuckHV6dCy1X3qPQ5uWxORvPZOdvJj7lzXmwhm
d1dy/w/+SqihPIzQR2cwP5dJHvHu0iH4cN9CWc93cBlToB8YFgjur5gNEx2Xa1s3IOqcZCvfI0IY
ze0tm7sF9GkPwKXAW4MSC1a0fV+gg3jIR5F3B0IbXmjTHDcCB/CkOl9Kywtg3no1XTFOKGohjWS8
AizFjFRBkOIWvpyYdFm8rVGVZCIxE5YRaPEa8TjR/OruouQIRonEmsExT+WwbyRMLSxW0SiL78H+
xK86JdkRJtsFkqBKsCPrcPHbgEVDt7ITjcrwOnmG9OAWq3gF1ruwEN5fmmayb0xNg4N2ong3JVop
PL6a1WuPuZwfFRHNlmwCuDArEDRbzR69RuIUGVhbCZLXZ9HZoqSB0oc13dU3bZtxS61x6jR4MlzL
SyLBmiqi+zrHAiP4Xiry1oFnDBSMaH9u14cl9eUSw1N0HgLI7L7HleuIey6mLEHQKqCg52VGqSKu
kZaUiXuJhK4zy8+/ZVGGAn8tzmBtVGYrzIA9XvVcnwMI+CXo1ma9nknmpGT+DbduoVTC2yftSDqM
6i3bn1JgmA7j/XtnTD5NYGt1H9ASWb13FEujSesLmhFnWCs8km1f3u/iOTgiuWJ5+AfRMB+pchnD
wIemyNWH60cHavezbAt59N0eyfArIntLDwavLuQ93tpUMu2+Fa2jKFIFhWxKZjYE3XKrUbDLEL/Z
3dYDZbv7dSS13thINVkaDnsYg0PuHGVzKgMCGaY/3fmDjAMkjIY/yK2gk8bJEuq3mQ8gMvvA2i8P
ws4NPpJS9uXMo9LPg4WabLJOuhV2XJNUzGjPi7o3l6x++I5x0xmKJWxx4gXPNEYMoCixH6QxpHHy
cmDO/AOMjoGwDJiO6xGxkcdHAlTYOBv4J3EjRzUDPWxnM7QZSsbFEevnsE6SlDhTzoLxlpVbi7/u
6rUEvaL9yaKS5/cmqrU8w4GGC7Ol3S/DpU3fJrvqZRDer5OssnLPP8FxzCwWCKR43VNnadLrXcdj
lQusmTvzUeKNdPJNG8njZA8BtcCiDjIfYL48MWvAS/TTgB9CcIFzmgrWUXmrO9MLA2h5HKSyyPe2
eyVkrjZXq3YW8YwhZaaDv9nHj3x2SWrYmOMgqXZMGiRrkp0iOD43eDEr6Td4zdgBTVOW0UvdacoB
46ODOVw9Xs1KQknMxcKyUpd5EoGo4w3b4UFXpdUJM65hsRqBwvsbRBT/Py3yvoKJrGcypkVzaROZ
y1GexN0s22XCaC0DaWrb+DqzB2ERuK1j774aSqaK6wZAadFD3O7hsXNALuDPWHSavuEDfdyMdF91
2tH3khyAE0zirD10GUVkykD5Rt3wYtM1y06tNxTElYKhM6ta2Ie/YMHsmU88fKmwNaRjHRWpBdhq
mhiOBQEtfYVET4WzHI3oYvnQ6zto86qWE0MR1LPVmD18co6bvssFn/+FkT0Mv4ctVODBar4CSZWM
KOA14ccwwWz2gTSEicZxkI4pi3PnTmVSMFDpET4hgQRawvWSPHC5W4KIMpQnlA29xceOBgIxnlDv
A1rqPVDBt7QMNcsaj70CUwnRLE5NyOxPG0sRzoVANgxnOwv1VQeU4CQoQiqa3eAmvX+vriRn0ort
Dtk94WV/eNmZJCaBpRwBOmq5ef8oC9nepqAkx7Cv/6sGybl4NHE2pzgTjdqEb/OoIJuZyqLc9Sh2
+PWykSF/BVQtl08Ksgex6wOTDziOK/yXtNxfsHsAFGG5FwYVrCRs2gVLwJhGKQol6rqzy+1u66M6
sALpIKvEO0N5qCxCZ5EfDdkTVP02VPcPpIRwuOmbUe8wAZy0rU+cNVoEto/riaACj2G/ProW6tpk
Y5zhm9JiCal75VJmXl8wwF2+sRadZ2DE12F2osmoNZZNY/yOfflT+5TZZYZRcIHFKRyFniUL5NHO
d9MWhUmAhSodQ2Quk660ZosQi+gf6Zy9jHjqVkZMtI7zu0WaiTlnCfTuAEzO4FIatHqpPnhiADD5
IITmlg4uPAfBU8oxzAUOl3r89u58QhD4/PBO3AdBOYQTS3jeWrA0P7gnv7o0DGx/qGYoYK9jCUj/
KeR78hQZfc2uqhp/CSFW9zbvzHDSQViPxX/jf5YxnfY5RpbtbCLEj7mKUihULlwYi43NPAvG8we8
720pKOYjr+/QHSAEEwGagrDYqacUzZzSwpOZKNrxmAYJyetrke6JWnTx3ryz+Xs4PbOOXvbg3mlU
5V69F9WuVly1rQjCg8SrVUtO7N/lGqAxL6ivzKHuvxslSoDsa1htMlDgYOo7jlLr96CcHu7HEOCF
ysuVHDWPmKt3jOb8ARfFhZXG7JK/nHiPDwM8Pa+AawoZn0iR0Il12SgSnm/1+zDNNz3NaGXmeS3c
xh5MXztY8IUHIyqPY45GXNEgslqPRr3KxgwsBDaWHHHQhSufXm5BAP6zdSjoX09ybIN86B+AK1Wp
xx77LBHoBU+PVCCyYOb8cLgeSWecuw1Rx5WU7/vZ3o7GHfkE2uB6/xkhksICEJP9gFLJlZrW0zuZ
FUQPGRJEEYoGi7Gy040s4XxshZ/pKQ4nZTZ5nOQzSttbGbUyolkNBQbkYVpZ6hgg5jpPeHdcF496
XKHuYYiqdfR7zf+aPUaD4GOGuVSiZhj2cLgXxLnzm/yUK+wltdVyashnSPPA1w3WkH6464ZW3uLY
syIQ/BNtKXyEjaBekyuFK/e8Ph7Rv5v5VydwvkBsv0r/kGalMgBNd3uv5WI0SWORDSJhFt2D4AS4
hHPNXeWM52AQfAuF6rmsf9LNe/B3DUydBvHRwVY/uTD51kLv5kvMvTwSYlBbUantziD0KcaiDk1S
5NTT/W6Eq5E1yDXie9z+U98ZLn6QnRpx1GrbSTIglJErF8OnFRsiQDbXA0e4Fw9ZlMnKOuxW2lrb
GYk+BTqG69RPi/Mi5eH6n4Lt2uslViXW4IhWrRgNemiGF6zjSB1Jnyne+4Wwbld4HM7icbc+RgWd
XMnus4jfiEwSEdgtL6QCkyegiXK7nzBvDTD0uwEP8qgrIDSE7Qowkcq22C6Eh4WjJaw+uOeVCuvI
e2WnQAzheigjmy8Nzq9rwq2o63MMCk5Nfa3q5jz+V4BqOo1DQuRRY1XzsljNyOOxmm6GKVkPwYGH
TB4jWKbr11PYotevoI8o1BBvggvjqZF77y5ErrJLFACJeRdX5Fv4v9AIGkoONFp5BoV5cIVf5bFF
Dl3g/962+GVG7NIf2EpW5ksqmbW0ePnrQnlsv1Kh8YLaytccwkj5gduuO+6S2ZvvX1ImgTRIVVs3
AzBhcIpLffoP83AmwYsOqagoI33Qd+S+HFxvLBuPwAJJgWyMXTrjvHq8sVuHNRMe+k+UDCHKY4vT
gsZSwAPKmThMcMNpx3HpdISKHVGNyRnCtHiQciztfQjNROg+yOURjrekVz2ft7u0Gve12NGY9GpF
jyHf6Eo0wB6uFj8DusoYQPKrbWtqKpCY2aT5CX1bJSOHBoR1vO9d/+aQcXawJPWV11pRNYjJw9bS
+HqLLPq7ooQcfOrvJtbFEZoo3YlumDWh7f0rKE7LmB0hjEICe/jApuenHodf/t6JV0toMWi7h09k
/4OnRoRZ3FXLOlFIScORH9snY1vja4NHV8ULdATu9P4CYTrvXCmbunAx+GkT3W8+mQVgLSF6H/sd
DBw5kBqIX9MBzcXr0lLmvRyevVzI8Evt7HQo0Lysa7Y0JMWh9raWSiO9uJOO6JzzLYTu/0LE9dyF
kWXZVH0+PL40h9JsoaHOiflO5CYgz1ckeYPvBmcBZaHCnWZs1vmhm2Ftlc7N+3k/BHqe9hCifmPG
nblmBq+y90WCm4+2fCn43mLUJjWeVdZSFwwROkTel6fvy5FFNO0gLjtOBZZxsqr8biY0QEIzoVwr
m6dVKzFva83Yig9Ubs6WZ4X4EsTa//vQ3cnswoP4vBlAOtnMjdcVBNF4T0U2Ui4/1It5GXAk9htl
o6vMmr8IZ10H+64jY/YmLiVKK0udFWMye44GZk3khNIXhXcaB631MkHp73Z70krR6pbwm1yc9siW
7sia+EQU7jXLuQTftgv63N2uvoBn8zkCntwVLR57mHeIkNlh97FwrLFQ++EXLdjjrM4UdVO3EhXz
1gNwh+uDV09tzd962ZziJC6uiOSdrwDPzBzHKi2d54oONGAoSukyQ12Lgis7LMlB3jtdxvGv0jp9
10HoofK1FvikO32t6t+XtQsVk8KMNPpjduojoatVoo5VBiUEO9mTlYrMCUJndlHiVdUVmzOgyj1T
CrqIhkhvNA+evmMjHbEPuGB5rO7PN8oVGAIP34pnrlDQmVYZXeTay2rToPUfFC+dBZBP7i289uRM
WQxeTyDAfmBnuKoEH9lxojGhy/G93SaOsdalmhSiCbni1YmOUDQo/NOENwyIwavJ5LYxVv+uJsQS
cbATFCeHz6sbcM7EEoyk5P/okv8CVajTDQK13PaeNroZ1kNiCwtLURCXTDxcnMzTbvqLs/C8WfM3
JNHv8v/U9PqO+ptzZcLAN5N275NwHXdztl29bDkiViPpJFpHl1wEJZ9ILLjFAKws/VMcjvD1N2ZP
idD1u5O06ZenDpxRHI1zj1RWgGsXY/JBwqCT6x7VWPEHsZ121yWwA0dDts1RylZmJsqD1wQi7i/O
3fLPl9pJVoInKzea/9LGdn/wQMID3dwbq+jdtaUlSDK0FhLJz7KU92ix9SDJNXIjAJq78WP+x94h
exjPjjbF/r0/uYVDPSRdeoNbI2xjz1VoH5eGRwQwdYCjfr1hvzzCdVexQ2D1nTWg3xfXuWG/fvD6
Blq3Up1//w9Ai/v5eiYmwRRk/Ov2ZF7B26Sj9+5Ij9SQo6pfo/rDRywzZ/l80VLA36iE5soYiEh/
Jh1i1cVDqqFiEUAuMeEARBg9HB8rc4IxV7mdIqGr/Jnicq/00UQJEiBytpVO5o0CtBxvV6gBYKzw
LJ6OMS3giglBuN+n8qLTwBYbWbKxTJWPQtMcCqSul9Hk6ReZnvYbDZhg/zkrKanAkV6sJ4aGBN3K
hcgL1mYFU4MhXGY76EEx8LMMoKso+JcAUjwYk1sX1hTJKX+Pmy/vM4x9JhlQa2O+FqfxGcY/83MC
nVwBQn32O30+SX6vEnWJloAcow2HZUM9EceEsEiVurvJCiY9SWTEFAjVeB7w4WJsNKsKEbW+UBir
LKr5tJHqkc0/pf8KwAhL0Bw47pi7b3TY7YzHaHB80tmWPhLO7ITmanT/Pidg5UFmylPB2469Gpnt
Y3pWa0+rsvXEq8wly1r6ZRyPgPCrZKnnuwnrj0nXWTb5NQ2VI0DzX42SLcg4ci2pq2jMs8zaNowv
VrJCG3BIbLXwUBeRMgunEFO/OA15JeJZkrRJ5J2ePUBltzQhiglyBcJGD/8GbYJa9Xtt1C+8Jr3k
i4ArcqKuNFw+Bip0zUjHIHwl7lMnPdyo+jR0W7OxgkMHIwhu/i4K2W0Zy1ZkYweIwwS887k7PUv/
MUdN7FoVGjHjFwGt+nEQG9py9zad+BDDqlVEJj2+8p8p+ahgYBiK14eXx2VrQ5hpGl/eCrpg2UN0
hFGiOFL3TEzznPcoveW/NvMxViQm3o6XVhtISr4LEkbG2EjGYg79csJUY1+0gK4hBEVPoG9tGS9L
FVd24PwUGbgZoI2ta3Z5pUqb+kfUjirtirncUUbG8NrUmqMTfqoX6Rb9sDmSVsJtC/9O5yb1Hwg5
eXr2yrMlafiBC3EeY9BDVeDCex3bjbU/kN5FFbjD39gPonhSFAtdkqwiK3i6AfrXvdJGJlgYCUHE
t2zTQjQB64ar6zVQ+VLJueZmS0Xd2+tx5BrXTm2wBYVlviK4qFEKyfU7QDWiF7UnA7VSG9WJ19wM
YlaG1lBEhPXBdCh+HCJCvonVdGeEBSE670oUnp2xK8ssLfyaCCXHGiPdqpGbLxZXSJUwLe2aOuxY
LksZXkIIMyP6O8ONgCj4Oeb7szhdJQ+K0E6ml30/36oBEb1WMs/wBWnkDQMsIGugcZ2j/k8yc0M3
YhPTKJQyoZVric9n3qRPbtT8GohAmhDPrjcc3tNdc4JDK0gpbUsjcXB7nlJ6zcKrPAiqVmQxxFQ0
zuhaHjhh6dIiPODWT8RP3jJIn99UqxXQrFIWH3b/7V9CkYtDBLALM27CJw/vlwHHV5//nRBRdco/
D28gYRBpMgXTSky1f45Wg678M4IRqh+tsYglDAFdSSeqqm7uIjNQ0ZW8dsWQHrmWztTnz5ukdJ7w
aFMekndIJp3UwRdyO1T1KtDf3voi3qSPCX9MV4v8wlMai/0Q6M50cSHfqVDhuzF+fFnEjH5EFkE8
48nhIxoZVkpFomRuehqPGO+fP3ZLC6bKUw/Lis5aF++srEj0cyAJqKfcK4Eq1J1lutOYiUtvGf84
eDMOl0lmCA/EXieeZBOUrki6a4D1wMjQh6MCe6b8YYWkyz8/d2RuypyKfZfS7+3/d2cckvxRX4Ok
eEizHAYk7O05d8ZIHZWmNg4RfC1PAx9XOmsthy5iC12fqHLWW1dtyU6S7WHJ3VICDcf6RDfKYoYO
TiPqGIZ3uLhlo0lcUHr4YMqd5KuTNGxsgYg/tu1VbU/SEVkzDM7yfikl64ZYSVGwlQUUZJglvo8h
4npnonhTL7RwPQR18kjXLS/vermAqo0ijOo3ipQNqxKr4nWNS1Em1z5Qf2wF4fwQOwwrtGVwW4GV
p6vinWh8iTe3kVn9B8hmvJ/i63PSRNZa4lO4su1lhw1pi7gH5flYrpZHDSGUEaEa/Gx3yLpbEl3P
FeG7svLRdwwHCJkaDKQjwLQtiFXRHv5cWT9h2AAnt+jdMy7EmJkpMwdZ9n5T8ShKg0Gzm2knTwBr
jyCGKNvzPWkncZyigqQWyx11O6vUYZqK96Bt7dKjnjuQ5nZ2K6ulqdOhVNPhlMnKiPRULxfoz768
IOebwzIqFudyFARWkhZuhl+jBaXU+hlR14ISKdN7J7xBPOO+BuL2ko6lS/qjhZery4VAPwHst840
TlJ68Njj3XvyExl2Vt4V4uNZtOsl9GI2PoRc2BdyJuC7Ijet78HhDFm35Hhnw0IJcnduOu/B0yW9
LZGNhcml4Exn2TGmw9d+DmT/CNtQBKPyY1yhgWIFAmgOVerZOu5ujYbpiUi4ltcJVlXn/fpqkwyg
p4+p2SZMkm1SGlTE11Ir7cn9eFOirVLaGnNsreun34HCQsP6K9PchPjcINY1pdyE7seUSjvtNhil
0OqsQ4czBTsCl+Q+LNvL3Ztd0ostSBX95r0NmmaB0bfsY+V5DmIU7CL5dZ1pB7Unei56glSXqo2q
wiDiRc2jCS/bP/ThDGE5tP9s8mYPq4qfssEZLXWea0qiJoUW73+mLlR1uDQDtCh7fQqr8xbratSg
iDyWJQ4NzBZ+CkBlCwfPt1BnudyWgluwvbrILAjd7C66Cf+600lHGtoGBdL1sjvZ+GECljJ8ZQVW
358EC797kCaxokhB7Vy8aat84S5+pOyAzUXIjaDDEXRaacudAyib+dO192L758daXVLzSTtj0cuL
vtgL7NVPXYaCzpkFssU8QKME+71IO/zCIGZKLq7wPukmyiLjWTQxiRlAgFaERYjD5l2IsN3FPTtv
NpbIY/FQTo6yF3zJ2cX5udhyU93FGZV57BlhutDJIRO/iJGPxZZajbNEZ7PU4rzkPG4L+LCwLxuM
jXE/W7y6gY8XpqPIQLhGU6IiYBgLL722OMcFfOEP8jLgyRbbuoivFfVPg/l0w9NOv2VLlRn/rYsF
hQyjACM59sWpnpZqU/DDK26MbrnHCHUbN/lE+Se0ns5/k3HoyoadqoIaSSUCBcvGU3D9U38c+53g
Cm9Yvp7Zw+3+8mLvWeOeUrmRCEKWVjUFkeJafS6FJQK/ShiqTegLuXKFUDwfn3jckjbABnN/qMF7
HqQOFf0dvqnlttaIDLHn5oJPDgg2WAzUSCzGVR5fVsty74DMwzn6df6txzCFAcOS7ga8umDZv4sO
nvyjyO1TzS/AEzeBZ7QTiQPXHvjv9ZkIU3yslDGVnvIqPIMf+DdHa4BF/fzYsiHoP6tFQguJejc3
qFOcA6ehqjc5HkfHoYWO93HQd9CRaGxZrFo3VVbuqLuoG5ir2zd9jSTKYSsR2rjrMp6L6j6zv7Pe
PUk1GqI2THL6LmeIw8fBuc+Z3P3RT7BUYxxq98hnV9qF2L31fccd+g7h/BawE+ChlFEbhgL01Mq3
TFq31zCXBUQbQf3oQJTY/D5a0zFXjYUH19BJzIDaxk7jjZuxxmrutt74hqetAyoUuAGbVS1W99v8
1Hz/7w9KaBuPHzEAc9R2r9bRCGyDgXcPGSNYVskBj4U7HSnAemEGr/ngtYoQ92sntq3a14AeHCSW
9Jo4BB3QlcEzKlooJXdO/RJKbyb5EhwhImcuqKTj7QXa7WzLYbkmu90/SdX8og6Qtg0VZeXvIfT7
iZC7NRiS3Ye3cb2JFrymK1eMnaxW/J7E7CNj48Adl8n9TAJA0hDGTKKJcv2nRZwibh5VrxO4OlKO
fLIYQx0hbobfTLTg3KsdCtha2lLUgUWej4k4/kB83MPhfkA8Ww1Bzgdzj1Q0vmZnYqpahhLVefQM
0VUY7tYbpwcvbtyL3HgqjtLR6ptuosrXYhkzYhUHTjaKNHlFx7J5Ew4nQZ5JmNuAWliszKYZVoLS
klB/5VNk89x0otLmqQyucHyyIXt4PXSEfGo1t4JuuZJ3zLTOdqeF+RR/iMsPKmnsjhe2xYAV9PH1
q2iCXI1pjks5t6ip8fUv2iU/GMNEfWhMLvMgaArygCDoYovBJRfItpdtlhMQCg7Id6vhUvshgpvS
ohRDlSb8BnT58QuapMX/t7+BQhbcCwdkqgrLjKJv3GhwxElf73bJtMg984VDsx8FdyUzJByRdOaa
TLUTDfTl0vU/9TEyLKv8hpDmEsNH4hPTW4TPiZGDsPucR4BLR82nH+wD0cvnjRW5qFJoy4E8x2wb
o+vb5G4oGIap5AFOeuV1NeVsIB6A++bveKO6nKnYFwMs5M6sLXMZENtXU59Vzyz/aYi7oZFJlemK
VKe5lEWN0L1le6I0XX2KBfc/Yh7AnGNB+nNHzC0Cy7sFezPK7yX/rR9olCQkMleObi/htbCHS1WA
BRuxWpdZ6yv+jpjVuNvro2+WHhNQA4qzNXxCWeHAJdp9a+MeiPlNeCqfUPjVsFPPRhAI/6U1EP84
VjbUMKy7zrD7BNGr7lwtyb/VywR0F+dw3j0zqH20I+sj7eariUXokUGVOrNz7uqjJE6Fn/Fkq+bo
OQzwEmt9J6GsVIfagODXxt/1xrFLwBccKP8/IlCt91TDVK/Yr8FfA4eiZ5Se1k/qB7/lmbuPwdCu
cZkw+0IWIZ42gH2MY5eS3nFQK4GrjXIFsRUD5TvGuBii93KAJB8kYccmViJzN96rgvuE5pIfUU6b
KE7CndDEry+sPIebDijqXV3NhyJ2M4uO3xItFhjrJScR26V8a3yRV/smTu0AZlV5YgvOY51qh9yq
oxxaZGW3prfe5SiOBb0di2VB903UPMTUvY4tdYrfUY0JovyAcuEHuOOLGbhEtQ9Gx8/Qd6dYoRGr
uuVHxlaZP58Lh8OMmqN84KZG77CzD/y/aR1x9kOZBu0WKynMHczK7jf8YqHZZhQruBviSzDt+mG7
lI1HKEGJ9KxrZmQOa7pBS8lUi6m409YHgqbPsob9sQaGqNftvbrMJUCdVvn7PmoT4lNux1E8fesR
J4ur1hX2yDtE2g0VEyowzEpoSy089csrec3B7Hlx0Z76FQkrqEcFiuJ7McViPOBLcgTnQ1nuptIs
j1S3FUIFfzCnI0BGz2G5TkPCS0zniCDI//3cAiLxKXdiBFT33SiUW/gC0tCcSh+qLOFxJGzIYA1P
2NigbUSf9dlB7onNcYvd5ANK9vig50kPd1PbGtMtMX0SSGgY1zaenVfb3+7G3L60HBWAcfNLF/Av
H+VWUqRx3KO2OQVbVmapngk6tO5yHtYRDYhZ/eFAs9eQrS4sooRFG5EE3r1IuNfrs0tNzFWNY8qJ
CLYpqtOPR9uXdxZjIEbjbkBHrX7u1WLH5uz4GWM9wbLFQr1PjzYL+MvGj0fKIYeputf7KQyfqJlW
5bFxgP59iK6x3NU2vyzJ2YcgKmPaqW37evGpj6lo4l6CzJM6o77Ddb4HuZ4RbMQ4onBiQCICvlc/
EMaYO1b4kNBH94GOax+CX5bBUD0PIaPw6e0U5RbPC9zI4yKUFUwuEqjDp87h70uofHr5UzlC16dA
zJFW39fcoUBXnwwD8w2EXWHEO5N9k4ncoeYRUOzJ3Y24IotsiXcRfcFHMEBzh31tnTEqhGEXsD2B
XidIOE48sI2PwZ01ks1jTmWQkRFqguK49DGJe1+W7aJVAEZOTCeyGm/4o1wc9ny1W8qQPQyzcnj4
DeLf34flAr2kdW2HlrbMEUutPjfvbu/lPTZCYZYUfWmmO9rzBKtBg+vt+XNo81x72HsbvJed0S3n
Lmi/epaeOWFnilUm9uupTjsEzQ8ij821VVBf91F1HIKcZvRXX3XNqHAmuDNGA9QFlgAH88cgo01L
lEDHKWwQRXotUIb9K+HTrpORzQWJRnzzZFNbU2kdGIZMhxZxRhXv94TKAZUnjLBUQkBPxxPqkV2D
pHKc3lDDsx5UZmstO2nnGvCZAKufw+NpBPCv7B9ZnEAGQ8KfEuEcB4+TCzrm6RpqIE9q8PlFg0ap
ZB4x2Mm/Subb2SwOTE30mlKjQ6wDhRJdj8nnSSSK8T96pLlsN/sURUdjRYdGII5H6U9U5SiZ8lM8
J6NFVqflLkXFe8WclWTzLLsuSdWCDRbd153f8O22JXpBfR1yc2LNemdodCrE5lH3fOj+nqcWmwkB
CTR/lFjb1JDXMO5LydUuvxQOw5Sm85vVeiyGw0Z2e2NtZusX92aBhUo095uTKRgWBVdN/fSy1PgZ
CafBfccxImucYnKLZTGPfwG2+WpKpDo+/OXHbruahnfKcnVH8XXz82w+dS5H7RooaDiZP/N8dUX2
Ei47z+/gijfFwu1RQrPtRha8dptBYrhcjbXHIiySEJNzwL58pbciSVQIGLXc1y4ATsz7lI8FvDgt
WfVW/BDbK6Y//Zly4+J/vpPqlw7lL3C//xO8lJdpR6tDM/Hdhz5/j47VSRrGueullUKU0no0HCis
x9FpzXhyhAk1olSh9rmjX3y8zVgaeGnwGerocDP9AFcS2RS4sP5nkwODKYNvh5iVaL4ZYl8HnlD0
cRmrNiIuUw3qQgzX1ktPUt8BLEPwc3x9cEE0CiV2djZ41WRrX/xEaLJ4xKOMfo2jBVaYMx87sSDL
FL+qmVdp4//Ny24sX/XouKE3HV3Df5uNafv4qWul1CcQ94b7Qe6JMZk98yWDhy2G0i8LCVVo6Wqa
BNtZVil6qX1lEHymBNK/wy+wM+ot6BiCHGDqVnbr3NTMD3WGlfRVIWd0gmue7RyS9Z8siz6bXg8h
mOgK5kI9CdddyOEXKtk6Fcc/NgG+0xIpp6K+p76QOSFlOSMUxxuOgJaV2tgO8rNls9Lu2DdbIohC
/ihizBcRPpTC7nbpRckf004d0Zb8ivPrV5pENKSK65eyqMLpyxyQCDRD17tlGlIkjUv8VBT0EtIp
IEql1oBwVRpnlF5dDnkJ3wipFVEasrvTpJLY5SusWjpMAF2JmVF5hbu6pi4Dm50F1ytLvWQeTtrE
7uhWObkdVJDBs7e/9jUkjlZTweleUFUJ645dFqOimnAShuHbn+OIbC9PalLhzws+hNXxgmS/GAX3
VzdsQa/A8ldi3+Or9pp+MNEqIWftDInp8ZU/Uyc3TDGof+nCqGMBCrHi9Fq3HvJqj9hSxMZoyoXn
2ocLilk7R51whXVMCVVWvTrJhC+2nu/hbfOl2og9o4NXNu0M8HTeW69irNziQvq0ZrgN+BSGsbOp
Qp9dZtF4jeJgu8gUTy5gI+ul1rJjrTVDCnSVGbwz9/7GDJbVqIfEzCXvpjGtMQTmpBnfKJEfUsDF
jpFrHLgtz1OKceDgAjiTESGST11QwtmM1MwtxLed90DkcHiOJTrTKZQcoPiYc05aYGdXMNDyp81T
EAZ2LPprxc9gE9ezn25QlvjGyml/n0NTTxOKGiLZAJAhuOp+89KjQSrekf+HBxsHGH9/N+jz22Mi
RwSEui17liywOOXjcxe3OVK7BGGryFRrtANeVBSJaT7p8Nz888BdscNU2y8pBC5L/hse1xGoivPc
YB1rpkoxiUS5j1eMk7PzmT2kz7IYfsep4LOZ1cn3EMtEJhR/AUzgysDkV/ARXR7MpPaBJkZhkXnq
PX91B2FI46FCS0b+X2dKGfj7JXAoBbaolv+4NnjrmMOW3O76ZVEoSg+AICbBUf2FPUQJq5YORXZR
hVyGMvZfK9GzukEF/8nk2rWcGlnr19ZRwFNFf3ZtPWWnh2oSFq+d9ZLrLkpDvQhaWRMEFOaFGMpV
TyLT2+tucK+d3qgE5dW3MySLFyg0bt26QbAUFQYrRCinlAVA0bsym5o9HGVgM6OgCoegK4BYIHFy
+Fr4hMVHq2HjyzAu9t+I7povLV3fcuNGNpZR8lYJem1NlEnT1JRVp02XY9WhFlmftSnFgGuthmpb
uKS5R2/u1ZgukyipB3MRczUg4VrdlVSTdO37FrgnkC7ri314TyNMp8/G+kQDYQEtz0LNSTTsgWuz
QZO9s5yOYCCDg+xLMQOXJyITfMZPHsAjcQFcDqOiDuz4hsztTx5OaR5vh+7zrPVAc+MZOHlYvxTy
3cCx8hz4FGmKLpVtMnuEM4/JHvPzeuzLOzAdx+0/sYnbi9+AnW5OXXmGLTD6vfmHYlyyne48EW4p
oKVaOFvLoJqecTif2gx+22yuJDUKWun+qd2OsFg2uR0PQdJTvfF4+DJcqpv0bR8NBjKlatK0eZoj
hjlgmFicCIRVGNRd2ZOK9W2Kkt3bKNx9to7pwgm8G3csYUB7+xJOABGyw49Elqwe0bTgpcii8Y66
MmMShBjjr8PwzNvTxf4Wc9Di0xtI3X/CWTCm3HoHbST/f487KePojiM9XfSfhv9H0eehlHowpQg3
A1jBS+0VCzLt/r6TggXySINfRKG9Dtgi3Z5J0sdsPVP5Yg2yu6NMDjuxnlof8ZMTDX9knZ10fwpp
EV3uJcs+1N3pAEGiYg3UBKGacnxOdvnlXCdL3gq9Ck10eoOwhAL3iHryaPcQ/ZzIbcAAePyiQYAW
8DpGDgEHst2A1+mvwJpkCOldt6X0/nMITH/eSmW0NutJw7jSChyBnLj66dIGI/inYJK+vM9/SyXB
yvUpE3RTL9IZ7H0aRnyPmEhJZZ2reiM1iHJR2o3FvjmdAaOGW770TWXSJd0pEZcDBGm3AjRlG7YU
446FRFcAPngC1pzKbSooWwDb0JP8MsykQxuW0kKI63sgp6VEujFw1TQTOvImnXi3MfYg10EOa1mB
pAK9/31ZVtXKzWq3iPczKKqAnLmMiF4kC6FDOJPFBDbiT/jUpWPhqj3UPem0z65w/5BQ1qr6TvvM
XzVE4r8CAWEEHsn8Ut/4fGPLKh0f8cbivZH7EY0iqxaVdmOsF6V7fW0kFMBPNMA8zhx2WG9dYOWq
VJAY8ZWJVDQ1Nz81uFrzHUAZ0oO0Y92V5D/NRxIwr2Ie5eIR8w6QTTqEtY79X4zpvwi+IOr7ODgX
3t5V/0d8qZkT0aUKnzf/EGeOVaOl5tpACd4RiqyKEXQi80eI5FKtj3QqKrlsVXYQHvSnIE785pto
Ua2FBH16o9Qkx+vn2xEZxMCanPLY7BAxlULK+LWP4JIXB0VgMNPbnsw7WWB9S5ClrYEV1SU0C0TN
2Get9n7YQ4zsLYDZDIECN0uBFP7663wz/CeaTqN0WgxkGAvNiwxL4pTC/JvyRygwNuJPZHI45tvg
y87Lfgnok5rfmBZm8QYFZAnUCvKloBfr8xS532oM3qwm9upT/oGWSRCm1ABh3zphpFZihzytsO9A
A+Gh9eijHcQPZiGoXmNHBL3BDZnrIFXKs9DsVGfL06ldrZfa7m5xh74T0YsmxFiERTaR0z4dp0/i
wbaUouRdo/OgsVLWuR+6b9vZVYLE3uFgKvRkne6Qgk2+agSz4Y4DmhbyBv6no3j8+9J9/Ll4ZO7n
iVCNPhLAgxBF+xZjLmBu6/QgzCgxXf91GCkhtms3SojGymek+B2NMdgGUxihtpqSKs8ywQr3QNJp
sKRTXi3Hc7mGyQ2n7L/rCubluu5QkDBiuyvfeKjXoOa3hkiVBI8dik31Ik1yATV1qfQqljTQRyON
oK73Btkv2x5frHXBEvvUaPr+q22wC0omYVgksYHE1+pRWl4U8hPDy+mFCkiOKovIdxpxj2hxyjxa
S/5tgPfWew9v8pS4ooEvKdwRK++37SnvLGGy3BD0yCz4RAjm4vmohIDhI5yoM2evrAOKvyd15rHh
fzF+lKJ9rI8s8bKgpLDqrGIa/CxQ4MQMg9R+DWT9P0ATho6xxuoKVIfhg1ICw0GIzMEjd/pTraA6
gGFFBuA7P9XcWdKQhb1DhtuueoerEdy3Lz79qmmZiTikwzuRRmsRdRyBiaSCVytudERdqzApkX65
6dyBDFdfwtSH/2WDeTcEdqgbvWXCID+0DK1K+yByXKpn6W46Q9ousFeEWP5+gTFvCHskm/UHW4g5
XMgy10XjmTawsBMNbPOSmWcMCwWwkruG3QL7xeJpYliMo5xVt8Z01i9fWqZ1/GXBYIqE1t7TZirs
6PRoFM+8mIdgdu8G/FZ8ayiYNp21AOoO8fK3Oa8BzWg060IJYzGu6Mw+pXi3V7Qe2lnjvSSg8v+k
CJiycd7VhyyGLroYXxfkzOVAY6LTNrKg3zgnAJFHyb4zk5OMZE2b175bCCaW3TPaERM+OjqhEHQH
dVNbWEnlK2IpUXwfLtpjKy5euaNZPMVrX7+EAJHId2Iojg2+u+wLC+TB6N3I6ip5r18YgNadTKAq
+kERaIOtyTCo/5vbyiF7fUH0ATykBIyOIpuSr3MHI4NeP9lLRTrF6C/4ioDv8jrLct9QyW6YeXsR
/epla/Wtb3KhWFJ93SK3JBuUyu7a2HdVYM9jimw4TTyA5qPKSYrXtfcuo5BZGaA/7z88kU5h6DGl
+wKHzYWZ7IhbIkW6IFN0uzMjpd0J3EELAxTHsdhTolbcGZD6GZ38GWXBG6/ELad9pDjWNEpg180w
+FQ4lnCBu7q8bYkR/GfU4MaMZQKfVCnEgbh4qab6xjgjPVwyN75mT0/D7NWXV0fu5140oVnSnP1y
9WqTbFaOvwgBJeklyLvvcZQm8e2HzOrp+2xCr7oSwm4m7+92/L2pN2cn/ThgIsJFuc7GYZDxBX3M
kPxv/SvGOH/HY6WhAnF/RQsvLWXUU0VgOymxMQe1eRLJtSaKE5nasxi9ZzwjMYhP9RYV8TVJ4RN3
73VWXrue5ApAaN8kPwR56u0AZXAjFf/JMgeJ8gaH6sAP9qpCNjOD6h87b9XAunfcd/GYXEB8GlUD
ZR8Iel7hUZQYA6iUPKYstqmPmsYLpcwx3digwd54rUoB8D4h/Llee2Y7QTOzszGOMbdPPXUd/pUN
Lc2lEr33gL0pV4Ej1HXbsWS/tlUJezTM8LDKIoT4uOsjnRQfCKIs/dkF8scA1m2xPOKEz3QK1GH1
GWus3lc2t3aeF0kGwiJ2eUGUkQUA78jxcRZbkVLCWdHLvBASBVycP6CB4BxEt4E3IdHNfkNrK5gh
h8n+zSM6Gr26+V9KNAaLqZlGSiesikK2EaIAByMsm0O2l1ENrQWXU+v0/22QpTz9jFf8y15rAd7y
PGMJLUXEvAy3CNv+AjbrgkSA8o5xFlpsc3CqK7ZjC34B7kUGgbDx1HU+N86y7gwr30Pg2yoopM7w
Ylo8UAuLBgmPp9D43lE6KMScgRngQs3S5+OHBQL1YvECS59Ma6/ZhE9uDRMNKF09yw4d6EFj/+ZW
Umpajuim6F6PaMcyXu7AeinmcCROCvuYp+jX/TAq2ueVifWVqoYElqi2aIgIpLuwjPR2YroB+oHN
dZ1wXLFkjcLtVbzlejlOLU/XcMJk8MlEZaYy4Z/KXjAj4YtRyzs/hQbTbWBXHxgFoe1kie7B2ya+
NBycmrXJ7PIv5rCpf5xMDWFHKFdJgCE7fst6YDRtN+ww8l4JFv+WAT8K0zAdP9gZA4oPEBvaMsQF
MmO8PJc4OUGopOHjPmSuQKgg7RHHHLQMo5dWIeRtlp+YhZnXYuWzW7/AIlcYpJ4E2DiSrmPaq6/q
PIGeMvEOsyyWhWmc/evOQe7Syyqwiko02oI4cPDgwxynJQdGe7NE2ghragXABJI1BEbwpjP4vhFn
Zxd1G3nPPz1VbagHQ9Zww3oJjfkxjOV2YpTmjfA6sArMrGH5bKj/3G9GZjmy7yqSkLTlHH6LuPQF
5mGrnZZhilV+rWqAVMmMmEEbFDTilLL6qjZbT1jyL8Bnbo5ihBXWVtbXFAgczWcPmbdthvmCJqok
77LkSz8cmfcwSTd8RJokEQqf40xH1tTL4hjAPpBqy3NZWZyuqnO9kiBc8dlemE6aFgNGhLPSopxG
u4iuDIAQDRsUcTuOsF6/846paKFl4gDyxCZ29xsTbeApxFxjabKRYuW1h91zDSdXcUQhluU6ZL3c
okNyM7oW/SvyBuaeR/y7It0geopueXuokWN6dDNrVUu4uNGH9nnlV/C3/IaOA+fsFGOdeszm+i0M
xkj6gt9BywLz93FQ16ft0M77shZqy5ehlW7OYV/3+kNQX4dtDLlAFCNaLlYvcgWD3yuGRa5IOkKE
lIxscFmcR2t7RodBwYmTpXll5EIT7DcJvCIEpAr4ArvDymybOISNUS5O5SWJb0FbGQ9ID5b7LFWs
+XpuTxt2p94H+kGuxyRakHcLxMta3eMjYEL3i2UGGIupXnqY/E1aZpHGOT2E1m2ROgW3mqilB/uP
6I+xs9M2bS+8bWJFHUfYssbM9M3Q97WgpuICkagJkCTVQY5c71LYhUCUzvZczfrXNst+NrXbjYX3
wsieIBIpow39p6Xy8PbBl52EBE5eE07ziTrsvasInNYluerJGz/jqSAgl4MyTF7ipKBByxlPJyu0
nKANsQon6/7Jdt91K9YDaX1K7hr6XJN7lVchG9OijTTBpWgc/aTigYi73Al4U0+mU8rnCBWi31tx
XNY+KEo1jdzzJ/e7DXRFVJ7V8pFyoE9i9SmQzrHYx48RtddIRTPi3vXO8kce4xytKpwr4KcuGS3N
3tdn5LHJ5TrI+l6PLnYuVL8xi8/lARApYjBwncWIprMNZlCA1UNnxmzHg7a7cEkDbhfGXAQFyk9b
TOEX6CjosfLXmIny7o9V0l8ELmk9TVBr/ziYRg0e4MWz8jH9TXiteKVik/FlztgQKlCVq5dWDmrA
oEg2Vzn7e7EgZruvW6ysnH7Q0exYqBMFZvnV2Z9xpRIUW+J/+B2MJoNlPn/VKHFsbgkdJ81PPtrV
7r4zCb/0oQlJa325aB4qwhkwn0hs4lkRy6oZMy9em9ZNPKSsvTM4ir3UR/eoSnF8WcGXIvO18Ex4
fTXfmOyQ126A3EY2/p1TOCLt1RMLyr9jp/KQNEvkq8bNjGO1nEzEGyeUDHC/eG2WrrXP1D3f48/2
UTdKzSJfP0ZJzjiKSvB+6zpJviINFqaUazUhFPyyySEbSeamz86zPgIWb0sTjbrJommOuGUO94Xm
q1pFEXzCqrmwbfbXqcfb7FVfUCf66kujvOFVYzyl4B3HLw0Vt0X4ZO4vlVCBA4ZiyIIPVyhtEZmN
hiaqLAJXyjz4Vv2GfZNBlKzihgbKvvifsVFkKG9ibDGRTV3jdEBwlgOmOPzGe++cRy89mGJWIGju
B3F98apZpZKXL59nBKlLu1eQN5W4RYCSO9RC1ISsE3BLk8Zlj9e/ahjDoQEZQBbeI+AdkP+qYvxr
xk4txxHsuHm6/pJ/dYEvd/KAK2I/Yyx06ozDBDhMdT6gLvyg7aA8kRj7wh1lbhugkuWnSGMUUiCy
e5TZk9ni8+51PIgEArcmCV+Nwy8Fmvy1mr1uKAR5H43bz7r9Ut64odOFAPS4U+NcRRq/gwspCSeU
9XZipBwBgqX/b+QRnfOOyNfpCl8JA9I5ICkziSPsDZuuUsDsvFUUhxA4VFeHfp6/Qf2F9Z9Z1tfF
G3jyA5Ckg7GU1fPWK2UsKX4+pd9m0OKRECywE52+6LiH6b0//bQ5p2Odsr+uM9RGr70zvR1yc1oU
fWFR8oezlgSLf9hEeaEW7GWlvO1mLGqkV9yWyRGus0dneQCppS2pxKjVsOl8kY54hMPJJvPVFHs+
4QsZvT6OF1wLt1n4xkjXTaqRnMoMWsxrFAUCh6kW+QhI+HBRAIZvNkaQ73FV6WMwis3bKgL4xM8V
vus+tXkHKd00OaBKp7ey8grmPilm3F9fTfuv5mOlaF4BPmk+kh3Vre1DHndDmSFhlu0xx4By+YF/
GXibfH6uu+RocEdcYbl3yQekXkrJ8EsokCfxg0yiLMCFSKvDDB8Eks6q8MQx/JfsLILme5Lz8oEZ
hITZf92OFmKufzEQIHzn8nupVQcu1lGJf19UioYsqVbtB661n203QKEpyLVv81qVEu+LhSdtAYda
n7F0VQZW7fF53Rb64UuoazDzubIddiTgWRFFo4iJOUCIpej8QBojwRXmz2vhGzVGyR5T9v8Emrf/
Y3cMvXcNOsSOCscjAwxwK3s0+TJB1aeNoYXF7W9wYh7bNJ4wc2VSzuJ2BNb6iP35K6ILj5ntiR3U
EOsY3tIaB5AVIxn2vSqj80jkQrlNZrZlf3D4CzZKVRJLwX6RUA4nEhgSY6gxMWUzvVDOK5VcTGw3
tYOCzsUZlf9GZp/ohM3X29pU85NwrRPnqhJp9JhnAoKiB5Ud9Wiu3FjQgF746Rs2Pc0ej5vov1Ct
QlQPO1bZ2CtAre2CnRn6EV+CQ7QKmJB4tvcCmu9BPn542dd3X7wlE0G+WIYmboAWo2YEylR/GCcs
g2KcNnReVGsWqOYaSQZoKQkljqTJ1Ks1hdtv3WTinMs9Yo/IFD3LF10mTJOyVTLb4Iv64XND7PSR
xd8YNA+tDR/Jmt0BJOkDFN+z57QPlb9A6gfD71t8XoxbrIkkitmYZzIIDjXcWxOsmmbUdxZkoW5a
gzze2JUSa3D9XysOBQPZhmcKj2+D/eb111FeYvRpGyh+GHC0m5ERLIwfksb5v/huOHIXqNUyWJcJ
qwPt8BZRM8CV1VFr463mHZYDJ6862COoea3r43CoZDv9wCh6cG6rwuw0WDr09nBQke4zwzw5pzve
TyifbkzHAN5cjVbjt7kLfMeL4eWoXIMsT0K4urV16x+W6DNoH+KhkDz2P3cwZoOTL0wrU2sOdgIo
HyP9uWxC1LvXWm9nilmtAg8Zi+iMgaAHcb/FsTBXb9ZIuENmR95U9AXS1OJWq6lbGCw2v7zUwRdO
WTaUl5pntRNSJswzAZW0lPbgsRCcsHI/TbpD5wLC8qjl73jiBU3Y2CMknwbed3jLAVlkSXIrwIZp
LskfcyTtdFECNpmMNVshq/stLI6gSvfPUOMjeLdn/hlR/fFlg2vZQG4bhu27RuHBFMuBsLLW9og7
MgHeI2G4p/BnsS+XXest+mAZHebV+CE+iY2u24UKuQcvOlN6kj65Wbxa3Uy6ZJ+jg3xbjQQl/+FX
Mv1Kw00JcuDBPIOH3Hq0hvgOkunSCjwyyablpJjzNBtINYm6s6iMtHv3niZZTlw/QjENrkzXMCoX
4PT8Gr4qQAgi8Rx1YdB37A0+eE5ey7fGHRXUYKPv30DlMy38m1plVau7dOtiexM+0+0noF9+wm88
YqDxIlCnxlphId9iUjwTEFJ5OeBoYdIBEPT2ROfu7DygfSXZ75YmZ7vqt+th5dFJxks3LIvDob1B
HJCNf1M7ZU9GxXQOhl4XnNS4JFvnhBydUBt/YnowWmUrNXW9tK0My4WLiRH9xpF7hJQomfbYwzTR
M05AR5i1uH7yAdly8/xeX83ugW3ahvIqbsoUri8BDMpTQcg96vX6YAGODd1hVTo+CfmRl0wfIjQq
eTjP0s9FkaFcuoh8GjqfSxEFYpTOh0xmUICsNLzsIs3TN7E0q2ihZ6kVrEy8G/J119qffP2DMuGI
AwNtkx8QaBFxSthdnvQce3rPscoL2VPXGRTqJEEXAYcA/rh4Cvn32iKQyuyr3/C4i+uSILtwM8eo
2PNiqQFS/kH2EAFuamiHThrs6e/BWj1bG0hg/1r4zFm1PKe0TtlLF0jWcnr7et73O8m0gBmD9MY/
r469F4gAiSi6kghJtgpsM6Su9xWryvnpXgN5l4pIW/1NGFuhOzIhSK9g1UhvDpFt1oK5rSRLVUg2
hY7zYwWAPufbXDlqkN2yjrmGmH5AcRr3OLGCcnAul+46UCNn+ksfK9xkryRTKNPJWDE9izJ+vI7X
l9QhHBOnr+eX6TCZpOjPZmTkDaLeZNTq6dFfrizWxLeMPjESoyc6BFmjTz9trVxgcoZCWlHpJQe0
LJuHh3eRkFlsMPkpcxwceXXSTgqbhvCvTu1iHy4V3vEieFsEBixuezhOy70N/X3x9yZ1rF7eJ3fQ
AEpvg+n5U/G7QEhAN4TUAr6kM0c7s1Zadbjq36ulEwW5GFfpl7yLk4LNDiPDBbJjqdP4hW9qyF8s
JBWN08umvT3HjtL/fKesbfGicIDMtGE5jqH+q8IjCh25/44OygEnPTqN+6NDdEFTiNSaPyRifbn/
WcDq/6q6RyK0rAKoUoyN5UJ24ieVSDpTL1Wo8TbdE+ha/ggruh7AkkTx5sPjf6+L/qxvOMTuV3Aj
VwWvRYHq4wsEwoSJVhfGNRALIN25bcqTS7G3MtX6+sz+KsSEZ1/L2limZNi0g1PKQuzbsyqYXTWj
7GcwWqt+TrBw6LS52kqWk0bPPVuoqs3XxLxmkaOO8va/evg8/C9BSIdL80EPu9g7+Ur9b7L+dL4B
X61i1X9hbIh9yKrUSOcJ9gMDylsL9jo3RAzp01oQ/nvCTYrVR1tqk7O0I3AlxXh52wKh/WAY0NAK
Swkmy+13Wtq48XxRXipeRgO0reI/cUW8WYafRoejJd25NQpr522SanXoEY4Km+dehcjHRjkf4cGs
z+G22yC0kPOPuRdKbznJNS1JNCUIIWBN84MXM6RiLgxD0EEyNJUboeNT1swQJPjdvK00Mg7Omyq2
3RWh02toXeAq9PE5AdkuJfw24FT7zrTbCoC8gxt4E++DU64Bb8PSrHV9D1oydk0dlH4JboyCWP29
BIIg5w22XA/Uc5GORBRWMtS4cVAfT9mE5FgWA6++DkZ7Pv5pWqoGWmZjQJGFu9KYIK4gVfpjO/pd
lMVWUBjoiGGlTBST7wq+8LXPjlKraNI3sn8GCfMV7TcnnJZuc+VipM1+V1PxqvIMruVDC/2kpiYo
XPh/ykUPUwPiGv3P1O7p6aEMTebwNuFk+6Ct+M3/CdMJW3GBqLAoVqv9zHWyiYCnbxkcdlZYqWsp
x8lfX8YOCPe582vjVUSM1bUYcgNcLnmQuo8TXO4cCjjJRe4BzpPGz/184UPLNWVzGtm66nRJHoh/
VH5AhG96TZEQmSAMYhO0LqXmLLud8eMLMdDL60FrTaENd/593Gmhp8bZdTeOk4Vb1hsps4F1TrzV
11Fg3lj/reBVFl+9/7nQatwZhlZIwtyGderUvPuZ8yxMnM0Q8CGEl8J9M/VeDaJjAv/ao1TdiQj3
0e7LFljcrXMhKvEVXsD69CTyFKtHUN7M1XjOZDO+V8O9he4EUtjSx6knXk7C+BbVZaT+0N95mA5f
idySlAs5Kc/6Zv55LUeRBjbxqRgCbhsY8S24IzDxFqIY585bmQUqiBDZ3NE90RqlmOLhgw3wwV3d
PYLdQKyiKrflLot0T2JI9hDsGrBRK3/iOLEUKyq9UpsTUmzt/w/Uw5d4DaXEWNZAJN8EArtdw7zv
202v6/rrfTa4ns/EapHErAF1oJlrbK2jfr94TzYpKma6QsjBsA231hDnkenv/IWGDu8CvN8aQVUH
36SZvBBdTeEflNdcb8vSnuYZCnqfgpz+3VnCfwq9/ZaVb0V6TVagUpe4gTrtDtHOllX88QSTOMk/
dv91jm3oih5azuGeOGNPKJXkKz/uok6L1/SyFH/m0malABkt9NAeaBhEoHUVFR6xr0VKWXHkvn9i
jF2r7DxlP7So1ckp1wDeKFTGD5LYfutD26YX8bs+WL1QPrbbjIqAzpcrqDrDF8UFgd9HrWSWYMpE
+eu10KiNF2sTu0oDZQ5k9tRID9KzjDkE2j8SYt+E57Nw/UqeGHuCkSiABQyN95nVEW6eZunxmZHe
EyBONNNZaDxVdjqv2ThNFgGoAwBjvE2a9Fq2he4QuwDgACgR2OoLASanJn/9yPwcMfeI6Q6uKo86
yh7433zyR/NpcZxFqyhi+3YNKGt79YoqMXmJyeANh+lctarna+dNGWh9XGvt9Qd9PATs9kCFd6+6
E2MSPnrMseAdcovLHBm4UaXpM4FflHX37x/EjmZPgH9PLTSn2HyzrfPZLwsCzBa2IuuOwoEEt85z
TEH+63pWi0PzsPCCKQq/vJMFX3qfo5vZ5PpMT2Fi3xR941wk6UrFWZo6+sk9F6kmaq5mSwq2rpAz
Ya2fbk4N+4XO8oJ/CW9DqW+eW+3lZG5x9QXpTcKFZLpdPI0VlaLBDIxPe3I4CbdgxxMltffl+ZZv
J61woplgn6YSXTM3c5QQKvsFN8oyIa1hlkvoXXBWW850EET2JVAITE59ZUFRRleHHf8VFjjyOLC9
bRn+vHzagubkA8xFp4Xv+EwyH/tQeHts/RLS2L+zZwvQI+Oqee4SZyP0tEGqdIpLx+hoKe67+ZUy
0Jo00EPSmFNZ3y6IO/QUcFBwIHbIsibUlVOsSRYaA0Ar0MJnkFtzg4SZ4hauqhvdq+Pfr8sgmPLB
KqEVqWg7PTJFHnr1k4fhFniVVLHiN+Ow2YlFQVvmnAf0+JgJjBgis3EzIhDaBcFlSKZ+8wYIT8uZ
mytPlDfcAOfPTYYIdcaXM8kSQBEIrq78dC/1Mo6YCwZuMEnjhNytL97VTxNd9zxCmZlwdiZRuEPV
+ajpcLjqXAUuNIzvptm+/QwIdlFOIcraktSdkkMNm/DiXgm/wE8oe5rMYvQ/wf37YAlZetzPNZ73
8gEk5ISgoP3+kFIxXBouLSt6qSykb+BPGtWbdOIrUZXZCs46pted6Zgpo8/Iqu2eDbc/pgJeVKeX
RWb8obLx33rIs5Nep4WY2QT1fk7RCWWl3Zc6IcKRxflJiyvVGzcmBY1jxnbMLbNO8XYYt3H/yZbP
q7N9Z9KBnNjtFUfQK/vdhkdgTsxrqPt8fFOLo7FfKNjjMM7VnKJzPCCplwDqVrRTSZSRcIqNz7Pf
8gcC0uXPbKEWGJqzmuNHnoVHcETPzBfthxGgAPhvjDiZ3u0uXTjSzAR3yceoYOSAeWUmNbFLM8Kr
4CefYkh4KtmGT1X0Y5m/5zdZiNGzt8/lhlD7aCgYEEtRbwrki0FBsY7O4uv6zu4sU+TZb80JQaDM
wAJNEoLaYSpuOccnX/YGo6OAYSIAAx4ojLHMZWBmEytPSW4R2N/jpAcqh31QYr+Z1H5EC3OJ4VVO
1Kphe0VWhbS2aA+5vkd85yg2p4cP1O1UeJD1GdrMpFHkku3qTto5Xm5dZZeieYITN0BxFSLsN16p
TvXGwftYmNqDCe2NTpFfj0pgBm4AT/U7TBjBZzvRI4X67zf3ClBW/wqDpKaGuhstamBz67Ydc+4F
+AOny53FdlHhi8W0/xa+8bRTZoFH39fY1jtndwUI9MpMiW7L0U7Ki8BpFQcD/5qcKE9KdM21Hsjf
eUJeHwOesKELkprlnYynnaznlrOdNwHGtg1tWvbpImfONbiAY1rKh34jJHmSZmSOT8xmMbdPgxyA
ax9ZmZ2AxpnHs9vDIec0tAYAb+vVvtGJuQo5Cj6rJuTNRfeFZuq/yI0nq3wxvnoeTlv+R6EOVR7c
LUcQB4IH9XCWYQPSdCcvwsTQFCHgSuhnOTVp8YwFfXpfhgTnw0mI6fbGIH8tE5NiebVmYRcjcAot
HnRumuBhrAKpLinlmP7K5WI/lfUIDRqV2yUxz5j/W2f1OoAt/BPL8Re5AXtrsUSZrhJnH2CEn61w
y7uyt5GyFXZXmso0J0/N/QQWvuqnIVXTaKBryUfp3yiXb7WNw7ezCU/VGMA68AIR/TcDsIkSPgQb
t83iyRaLhasSAoEEV2ABDtwYtiTcURbTii5ddOUbPbsSU1GTKuhpYnEAOyT2NlsJ8H+cuanCKMXQ
BMg+crzaIk02BV2dwUfq1tMC8xEwStAT3FlNQDhYr6KNTzUbWGqrrVCyBRWt6hyZplsEKRtgHXm9
4Evr7pUBQfj7iFZXmZSlGp17dLv1khJCYn7CfEiobYoo6QX1278uQxDsvFcInmY0dmCV20nsdbX+
c4kJbgj9tpvquLGy6kTIJCnciG4Oj1x/T9H7AXCBnvA0sgStV8MolL4X1DzT2JtGNZpWbYOABdj6
/4uZ2QRlhEKQ+/zUmh9BdCsTCFvOuUY3Q1KXYWxhSPrcPZkyh/TNG00cQ9YFVy+2w6A+rNpysnbM
72WjmfspDFXLjPyNx+1XA6H8Qx0NWTi5Kp7Q2F1tzVsirj4QOgzelEqbNj3wdZmOGIqN3swHqMrF
TZ8dPz7wHQWKFYjMeTa86cGO5bI+9YlDlal66kau0PcdBH0WsVmNDL1hQFXzVNYX4VnbP/StR0n8
6zmftHUg8hT+aRrsApTLb61s4oATeaOM529lry8dtW0jgiMJEXKqR3xsvUVezVz/1oEsC+mx8iz2
7zl8Gh59RZFznSwo0mxeNyhXuwqmN2IQtfP8txGlZFLbAxtNtPzSgro0qvnpRNKds/VyJu3me/ya
0CxJt58WHh1IhKhf70PqBx0xjj+W4LZtQOVbQRkEfsaz9wFC0ZHEYtiBsCLT+gfvHF4saK9e8OXf
bonPRKXGOOJm8ROZIjNnO9WwMl3eQjnfkXETQ11Zrt6dWyaQ2jzMnMEeXFkSrRp6MsmxbuIv87zE
abj6Y9PyeEPzxM8U7uRQtvBhwpnbOMxNa1/tIq9OsORZBpWI7zswrxbkksKRoDtAMX0nsb9RI0VU
xJYUDOBZxd1U+XGB/o5xt7tUovbNs/kwp8+oax3tAXqXeCUIKv+Wd3qPz5K093bNeGlxCneiR2Zg
lzS/0T8bMKAJrD9jtHAqRFPUl7rrIZklT9f17q9V3g/2mfQkvV2yLL63eVYqQ0I/6dgjiFgmB4iX
TtYEG8uGYv7MxLajIiHbrMnsfKmkG3dCUYn4IRqtrSOZyxZf5i2UL6NbT0hg304deSitqnDw5Rka
9bxplKkyaHjyDEneBmnEal6xRyEXYv03zrezdiN5PBWKAz7NMqJXqbjkrSRVlgc2qI9sfovL0WY9
RewVXUwKt20oxt81zmbMBkb4gCRubP9ByXiAEqYuwGZ2cbayXJ9wcAyjHiuagt1V9zy3JG9PAqGO
XKRzKuxg3Gkuk79dYClaHCxvBHJQwIKdtXHZXL45cyqglb+I5oZBm42DYoNL+crj1KjWxQiUcH+0
GVfTiGUhkADlqTOivP++ahIz7QEBkP80o+91oi1LRF0SxZtbz9UXuUdG834jwslDiDKaZUo49IT0
+/nMrOKHRzVhMtoS/wbRAg4KrPNSPyEIsJ1s9fg4rgiP95UFzZFQk35fLP00e/NE63ttPTo0f4sN
aCsRiSfUJpknd6r7vrieLoo5vF8uRq2gGm2pgrksDGRCOGe7D5w9TwsBVeuHchd5043g1b2gyUU3
c9h+Mj5Qlx7Q/rjOA46r5j6jqoY4Nzkd3X+8h5/l6MRrdOahM7SrFwXXPYf7dUcL1aKuoqmJQ9An
ofO4Osg7NBHT0FFKoF+KKA6zfapH6HlBFquOlLPv/ZFuADV7L8yC4SC9r9ZrgzUHzwXMAzG+erZA
6D/MJDMa6uGybuDSdcby4VLwaHqsPMWoeaCABCJfMbQx/PjidNN6H+AbtmGeQ0l1UdOSzudDM96i
DZkRhjhzPfUM22ry9S8x+pELOe6DjTwL+ZaoGRGC11pB/eMSlAZPArwnh6peL2eQNq0iL9TyF3jU
9Vc5VgdPTsUWft/JBDxpcvAga87i/YKkrO0/VbXSTiRdGRapu9MyQhYz8p6cgBY/67I22XR2jQWs
5QFzdobE+kZNNMGgrvxOEB3u6ScAhVynrbWU21nSw5SR+3PaS70EcQit/R4wvKRmZaoVzRtxPeI4
cz6RmPzcvDnoUFF8Y7JJkDSioBebwcC4zvHtMDZsG7/fIZomICZ5VHSX54H6ZHtyyrwYOGvqXUQK
Bre1QQ8J5gi5dHwV/PXIkrl3HT3IM+2lPcfmEEI4j+001o/LXcQ4LeDyf6fXcnys2FSK3od2qVOe
T8J5vwufLuK3uMRb2vLNVibmD7sx+TbfnCXFGltcz2IscFJUDCa+Azs9rB9OZPsu/ckyz/sbobS8
KtxXQZbnQmozvgRWCHRVx9ntrWzP0jHU9lGParhbWG+MZsyGfjVP6UvMvDiiN2tgxnmd0CxDCkrf
rp8t9eD6My/TUjyuOrGvPAMNpUDtz2Cl+B4lr4hJMuWlUqoIR6q4r7AiNt3PywL7bTTpHLqrSCaJ
57D3oS1k9JIsiYJLe+70rnjtP6xG1HjWd+TAQwEy2xHSC+rE8Gw0mv8nKpkpVfR5eczBMxP0i0AZ
sbTBoIVhXST3vH/BAhFkJJLqLM4FMAV338of3mIdgCiqd0Dad1gOqB3UspR1RZBTPnx5CcoT1i12
ZWriy6j6h0sieytURMWnCNHD0vv8fg0zc4qI6DrCoPDHw8xXhbrUE5AvSfLFb9RqTEtqq4mHU8jQ
GscZJ1xnTxH/RRKWiXKX1jWfZnlmPWfUHR1tgb24PbvErITGayx7JVg8h5DEzcyOF6t4OoILo67/
vzd4WXma19ZpCBMXwM0rWYGhSw4NbW9o9bMUX93Q9de4u/ODVeEk+hJgFXmMFphH1hbLXD4vGGLQ
iq3RMA9QpDBvvMH/BH7XzX8UEO1WTqOROm5TH53beqVHjW0ORYFzFa98lo2wTDdxOrxA3Jzo686c
YSil0h7GM9SSjGQTYTVrfP92IIxsiUafkjO2Fypx7pAAYPvwdoixeiGPHztINic9/SxM1G5iXpMD
VGFjI9d3exj4TbOOjbL/Lpd5Aw+GUzN/qkeL6fl8rLsuHtNRdIU4/cXU3EV2lVl5kylcR7xZERir
Wy+z6gSnon+rIEgLf2YiiKpe+8ZnAjTKne4FLrmcu+RKTpgXVAAxuJtOPc6fC0JzbW+HpRepLsmA
FlaCbgNdbGjB3HvTJCIy17JQ2dADpd1araGPjfVxny7hYDjP4UEZ6WKOdOIZrnzu/oFr2t4cdPKy
xBQ6j7ChGgu63gBCAEL9f/oS+cxhStMUfZp/AujG1WJQ3IrtAjgRdPCZMQH4brwtwjk9Siieiz+A
dA5HfEQpy6+HNWFtyx6/9+7bBA2Scdkj8Ep7Yi17Tdm6hO/qraj8Cdf+HgZQe58LeFwFpyILoJdQ
2G3e8a1e41Jt00So43xI6tALmmr1VrYhTAgfirygd9JQ3cffvZSDDryV7+7thV2gs5qSJ1nMymfj
KIm/HfyPBr8k8sbXTKEVmMlnHRMj6jWwoG+jrmfj32i/yKBMN++06YgbIrEAeYlhcI0x1UePpP4c
JcVaiSvO42D4ZSEejFlXiHcwhfifd9TOFPmGh3urEWgONbMne1qkP07CSC2+GqpXtEejPgv/B7AW
MOVFLWKZvZs+aJXJv/1Mu3vqMfV8xCZ8LcmbFPrQHhtNKp797EVmila7exm7Mx+3bF4m5yXsKE0g
RuZwFrI8oRGoKs9gQ7LZdRNUs3EHTvLKtKaRvDuMOCDWWGti9dAFrmJc0+kC/WhCM+WpqukZlMC1
f/YkuCMBLTE3fZz+f0LNq/SBr+EViAmLCFeQSyY6nV8+jdMtJJlKn0picuFQpRzP9uXOGPD5Po4J
DMjsTbYL2qteXiyx5rghiWX8lA1NU5gu3LG4fkRlYf92UMNuMDvlevbsexQfDpB4H4bJ0/xcInVB
sx7eKRM0frMntHaqtXgvELUVmhOolqiFOP0l7nwwybYwy6YvfOXmL4yRPCLxJudvQePCPWirM6QS
i93uK/sOuahmJUkwVpdPWpYGkqiSQyd5Hpg3DFfPARyuBe8vri1022KMwylznsHJrPzA87q3GhLD
W+PJFua3watfi8QOTNFx+3boMt5Iuc1X6E5+Hmk40B6rkU2u5+lkVO7tny15IW38gl26sNmggv4Q
TdzSRkEK4mPk9aAlgQFiFun4uKPLc2msVzKRrPVziY5/P5G2RnSX5jyk739TGjlaFfrdfh4RHDfi
YTAdUWVZ2FY5a0S2/jHiaT8uuJme/Y487rUpWP7yBKqmT5TEtuTgEcQYQs+Y/Z1F4+dwbpkd7KaC
k7vVSAOscsx7hlRiAmvnEQfUEpkHaHKp7hAs6gWcF1y+Q+IEY9FbZ504UdlX3XdBIx9RlZpDmFgu
orIk5M+bGsbzZ+luO7tDBEfWLe0X33TyXCeXfAZZaXIM1ZaovMlxwdjHif886ykRz5EBKhmIH4xE
7ZXB/KPV4UPulQr4sAMrsB4en9gO1KIe94tAnjy05zutviF3lgXGgJp+CY1D84lvgeR8jRZNWaDG
XGOYZe5yhy2HTajznLwfmsZ6OR7TEGpw1os+wOPB+3pl1ME6vxFHh9O8+rBpO4XbZn/nRdcXR1PU
4cSaq+skZu0X6oBvnay2YdWBKSkT024TijYegJV42dkBrStV7mCMcoW3Gl6ku5EiVg+5DqcrySaW
2alNDVZRsrxZD71npMOp1Qud4dKZNDgmiT5DiguHCXHuaez2skmVZqGqOu7DS4Wh3OZQebiq3gxh
Bv5DjLE8xhfM/DaOLvonNyPTRhPTxDRdg79ikL+Ek9vzPvQaVFWH/7zhzIwB6dnP4/swu9AMW4Xo
QsvTuce+2utNKPGUXEp/VnkCCKbxqvg25af/sGhi0XYTibfGR+jodzKHGH8xuTp+olI/n5Gx6W1F
8dfH6Q0ZEIeiYAVNdD/jli12zc1Bg0+EddZFsZDVww0sCEr6FaPbBQeY7xRDetUPpxc+HuJ6DLvI
yCsM0FyeCLIGUlrxjU+4wB7FdYx0cl5hvU7BISSPCCoeDlXh+gwHcnsNL/ls3guhPLZWmc7aDdLH
iZUPVwLDnHT9T3ndZ8IImBeBvWstNYsRQnixbhEBie0C6v7vI474CaYNG3vhwNK3Ib37OYM6Davr
YeywdKKlbDkaRFI2KWtHg+JUTRTJJZHcdbFsbN+zTDljSzOCACPzlNBGO01BlJIS9KIT5tlAiMLV
Z+t5FNelBcvp9mVcukIxVRLcAD4UT8FmBtSzSik8v0HRKFbTWtvPeFX6X0sG5dKWJ6eJhVJ3BgYB
4JYbamkFRIqAvfjRD+/iZUljl03IJNIh7jZlSgzZhs8R6gYtF0TVLKGGEyz9vxxNb0vVmWMKD4OV
ZWdr9jvyEoJ2+nR1hcw6dCL+n80sB31JJ+hJcA7nTG57Kek/aEilX4kPrcjho75+i+KB0w4nKpu+
ZmwDVIcRinUNBHoJmTtxtaGd0EYtMyjXd10tlgjBoRxiSpC6Ke9YGceP9ngC6DhP+HXfdZf+2vCA
7jIWYnueLi0M3ktUoz4hKmQ+BtD/Fz2L4WHiAoFInpzNwrJlmSO3lS9C9GVbMx0d3McGPYi+tKW4
Y6uoETAt3gk2pGyQg5ivzlKoGmFwIm5NlEwKkQ/QlnpzHYqY4/J0NcwXq43be/53W+3elt1fxO/C
AD3waj2TDgK9zTt0Ew9Iv/e6HuTZC2naViXapsb+pbatCk7/gz7PKBl09UoVxaWY/ls901tNrQr9
GdXZ6fIzYtimrkzEIX8e4NfXE35FbB5GfToRaCIJFCMbu1FBNzLJ9ONWP7A23X0Kh5sVElG791e+
oR3Cim1XuHz39YwTdGYmUVGmTPA8RKavnfS8DtClqyFTeDUAOJXxmr1KMyo2NsHcsurnujVQwZJn
GvW447I7ZCH+ff4WgDx5yOMqCiewJCH/sq544Atns47gh6PqzbqRIq6jIzOV/1kSnbdPnrXQDGja
OsSEl/VtpUX2mztj8OgDuD9yIVS9Yb5OJFoA+RKb0k8b9paWZZ7YJjRSI0VBtt12i26ca/vXIWAe
jEOe44nN3Wr7xouQUd9+Pf2FjBT7bhjGTbRZOEo1w1c+EdhHw5Jidw/3cr6QwxIk7X5G2D6OQIdC
yV2a2pwwlHRwOpjXvSF/wqL2evgnglZctvBUgi6w5xmQkhILD7r4t5xclzaWugp44wZlqwyV/RA9
xSza+dXiVZ/N/juzVSdPiGtGwt6U6lIGfrH8HSKiOjpUe39n4ivrqFRAPQKnQYNit9cHces88NEv
RtmaqK4ncVki/fOIUOgzOKYmmNIyFWba8mBgne2Uf1ndKmsZu0DANplAiNLlqyKyk/UiPnGQsLBT
9R1NHh9RWia+DfWWhbMETvBnLih+7COiKkH7W0NlPxMHU4kf7LxY99v2wRLifLzUs+1BJvMK34m8
X6Ai8Ij0RHU4gbDtItthEVuL0VaYNk+/z8gnu2o0k7R8/JcXWBIlFommWeuL6O0uNqthHZm5e9EE
QeBTGerO9ifOqY2vOMrKkrBSBmK7FBvMOGE4DXpiH3hqNfrNu6gWlos5w+OdUlj24ZbJENIT6nGc
iH/QCxKDy22RvQRGVcp1f7n4VEBl+tts5J7I7Z1g+I+n2SwpG/mVRPmWtk6ZihWEc0sDZiXqt8oY
oGnXnIVtU52YPbxfQHXkFHm+OS0UFTqo4+dvrX2b0SPbO6LXPa2fD9cmntEfwkmMiXpfJvxbmCd0
Z/gWLJu3HRo8bJ/eAiCB5gydl6Jl7ate37k2NYN+sNkbrvvlrgH3H6UH74iQFnjL6WWv3FHD9ndy
Qx60H86n3V0fja0BqSxtgczM1VWj4+bkSJNcPR/PF5IjQ4HbrycZCg5b3kXtMKxyuGvj9Ffn6UGs
+UDOT3KsFOLZVfdrY/6xeXCDR/qaQAqOu1e47Mb0uKv+3HOUM/hqOD3SWG1oUoAO2RxhODPoZIAO
h/fJ6NPnIMkA4176ONfnCLpp8uFyDLDali2L2yhycoN5Y6FMuUx+vsU5VTNhvyYki+7oi2L5vcxP
h3AISFNx6+ACcbNfl6fF8fAyX+6Am1zqWkImaRz+AFFTEeqU5OCWV1L5Wot6l02fnataBssaQDYx
aX16NG5ZrggsA1QgdZCjmbxFmkQDwwu7ixjCS7EwrAZ9MoMlM+qlzbEEaSxGQk9jqN1AT6/keAtM
xEGbHCzdXuZI1G2v3EZkRxI7gsrjL9rEN21ptdM7PCSPghiBIRlBurnbF3A5moO3Iptp1MUGoq05
R/naaaGn+0e/+XhgZBO5Kf/0E//GRLfKMmo+CmKjhRwNmaoAz/XxdSxd+1NaQZ74qDUeLWZS77Ud
+s+jXkQT688uEwp6RhcZphSAJcsvmBspqr0lQTWmQGLcCDdnwpFuXXTfcH8MKH5PAr62/yqi7x9P
XrTU4vBubDFgaBy5wSuDK6POCYSZsZYBnsbhvnKwpnmEy4QjLXzLbIFdb6WxdZoA1CoAuT04tBrt
QIHt7JPxI9WdnYFbzaV018HWVIQ1ULjG23Odbq7J3cPEj416g1mlaWlNy2a3dXAHI6jCoV2zJNYW
P4q1AXimRIeWN58grvoCfiFRAar+Dok3h5D08Kq4ZagGYf76XVOByW4dlgx7BkyDRxjamxKaOYqz
b0BTDUeXxiZjb//xWv0Myr+WJlW6Ltw1m6qVDDlKbAD88qnE13NBIAG/1obzWE3hT4MsBx2CZfcn
4aH771sfvK2K3ZpHYGbtgEusJX9bn0v5vO4EMLAaxtccui10lHR5yZbYNsOburNGQ6nLL8mH3d0T
O31pOo8HrskwLOa2VpqwS+YSFR4D/lIhFHAAnDTwqB6o5IZgSWpn8ysjsf0XUiXdaPgZaetRyMV2
qGKTiSMlnvT/YDd0GG6fEBXSVQUuUvxbm1WYz0qmb6Eb4MadpkH5UuEsrXQ1+7gP4SycZRKqlV+Y
Q1elly8BlZ6ZpRl0D5eWQr40G6MwglT0116/ikn/1quGh8//5E5C12HQk8KUGJBsKGJaFX55ZnRC
DCzsKXNdc0CoYJsA1myw9Ti6sx3nrlMIlNT9vzEWhmcusHVuZHFcxvaxKHMnif4wg/ucjvJBHWZh
BjKesJzIlpCff5/zKqck6aJn3G0LVIxmbOlRTGk9/6iZiF6MzwhBzSLaMLRm8jac8Cx2eUuSYDQp
W8BIDEQ1gybdSJk5c9yksEsXN8yRItL4abR9hWCHOKTOFao32NSs1lE6yLQJwNvNircasxrDiaiG
31U1N2kqahAuPkbPD36PbM3MBCEmjStzfew6nzY0h11Q78IEzunkEtWwr65sU3xm75J8qRJYvrKv
F11ydIWZ98lsLv/+YNfDHNNuHSD6t2lqhrSo6SyzjHhXXCQBkQbW0AIF82vBc3fRwRzLFDdbsDP4
GKWRnwn12BR6C2VB++WFnzP173gyJL/ZgkzSgytNi29P1gyN4zBfFp9vmQvbRzm7skS1bpcxpljD
TuE9mof1c10r/vujLm+BC5pAknGkjioAVIOHF4JdC7gsLjlUt1iabcFyi+Z39iKoLfwAyr3f97Os
ceruVao6Jrr35sT5mdqm8id3LOHUPreI1XomtWTeke1ogtnP7+VPJQJmu77Z5H1zyoaOJeqcg5Ts
QRm8SRba+Mg4awXOFtne9sqHtHRX0uFBJPq8DvdG3VxilfW2HmLU6JqfDVNyFosrZ+1JNpJQLLY3
sW73dhzH3DlF5AFQMPy6FGaYuPfRuG2d7skKART0ynVT7yEnkxb5iqGF6vs2WsO9tP5Xy1poaF/2
bJu4LtzH2DT0hU59t/9nTKNWhZMcnzqoA2dmi1BIqGpwA+aU3eBA8wFF/XWA7AWGNyVODrLPRdL3
NQRIHj2o+7iDrw7jEzcJMHRqfleQ6vczBi11+miM1qvldM7tPb2P/DesnOQC8QwupMeqtPaM0UY6
aP+q7iXtaSy4Rul0nOmNP5f1FwUgxZMbUghK1Tw6JyPD2sXRZqwwDU2pg1t7OkDkLy3A/tx0pasn
vHf4Qy90aIpDc8tbaaXtEptqvrNjIlV2nmDGJxEmZGzaS3LTb8sPfjWqQa5usWvtASNiUq4bZmAv
i0TrZye/rkBAGioAEi4PWeB9qIJHAt7070jjCrbEJiD3GuvvRjeuEZG+ALVOEha+4QLp6HdcbIHq
KbMz/fzNk7Q+KMGA7IMDLd2aY3E7BTCYZLjRz65BLL2BM1mbDTdQf48t3MVuSrzx4BS7YkaZft8p
qkrjFbLL07HSV93OCnROkzMlWV7Qpdd/CXPN2Lh3X+Sd7yYA1Mw96Z+NA0tgfB9tyTTtdSyGcMlr
7oP4k8JqoNx2P9P0eYhzCM+cm1UQRTR+u0280M+N0mlsJn1nYOdfEeWNZQ2dYZeM45Hcgj2W5RpS
A8uu8TNNywR1CoR76tPoQphCkRkVX+jqKq7k1mZPVJQwoNI4ovVZ6enaGdERP5EUP6LBYg0tFjJ4
oUqcpjGzLH/ztLDNt07SyFC/2tgYyRYlCjoNyY0LlAFTPMZTa+yngvGPatSycE+WjdK4qMt4YqKh
EBkS0uknCcc2XQ08Cl1bgi8W16bcYv/YUQRkjxaup/rWCSHEwHSeiUCg4XmFUmoMcdPl5NYmjiLO
bB7oMNJEOATMYUwjqSJN6zYcVHGGjHMzt+XDI9I7UF3IhJZFmTUazrwj2B0dyUD+71zEO7dwrFyJ
NT1bFjiBbIgS4S9vQMunMhuURu5NpauP04iV8xcVjTL7bbdTxaqqHaa8RFkeXXMRVLpx9XwEJqGb
lIWGL4xeivOf0ZHz01wubEz5jBJP/dqUiGuj71HxsnTKMPMgnAuobs14xyuhAnuW+4SOKQdKXJtG
BHeyH/rUsRSOQ7yybvuLIxYlJTjFLdVz5gaCfTPw52F7Ygc8ei6hqu1jLbhD7QCkAqkI5m1gSGxe
NvdXHui163Il1ySuLT9JaeLGCUmopcBFZ6pWPcJmyrQ+tmsPIa+fuI06StZLHuhZJcnekqqdcOKy
muKMP43vZWki+puoyC26ZsOxU6zu51lRYI4fWd3BcBvXwweEgXGN3FGdhBv5268i211Qo6JLfVqu
d9kI2YBP26EwWp9C3tx2dYDVmu0fI+IoowjdleYpqTiUd1NiwNQbzL5BC/m7dsSm2pdt9SKsDpVp
mfDRR2bj2ZDALSVf5sRGrjMBExkejQhliv/kboIJPxikgLIC3X3HwWfcr5Vw4aBY3zU+sOCS2gqi
nScGUlFrntxgV2rrNQLsRV49DT1BPhaD/dok7xQbKcOcz8kLLhyWbCqFawVVQBZKBxWpf+kxMetb
E6bIYe0oO/ycvJiYPnbHBgxKClZqjOXIyFI8BGxTxMSHYyD7j3AiRzCZ78VWkF2jomfSmv/671aw
f8L+gmZwy46/XhOxxOCZovc4fYE5A5ja9UQF8aNtfs4NsxwNrb8GlZkCFWR1EtqvjxwP9npg8FEI
b5VsNirKMuqj6IkdYnq8wYxRmRWnP0KbWJkSis7ZOBXzHI8D5mfARuLbpDlJXKUiCIGBVW95iUpJ
Y9fdcO9A/cnJ9wn8sM32kOCAoD3h008pEhVhNXdaaiohHrMwL/3LzqrTBR4r/LpMO3RHJgCeMSi2
ViKYJT7P4nCKwBw10UQQNuzLU3lMMLVZtlkk/CmU3mWUiVATKpX+pTOWd1jEopTsZxFGnc4ir2GA
Ph2VJ+k8fYeGk57t5waT4o8eXMDC5WuBqzhWPSqOj6PnQBkRPIOEC3YevqQcjrBLt4MJ+eo3KyPf
AA+BEcxuTDIs//ihFmXaWRHnv4cyG1GSe0wIYJwzWGsHr1isg1dAmmf72mqC5+QsvgxzGpv+ZSBz
yi/Kw5OcRG0SO5qe84aU7qjKpeqUSPn9Raa0318/ZaLyGxNEJqceMGHTlGbg1y+fwpwC9g8I3LLm
yGxHLmi1hpZhLTA2UYDwmelgX3MVD2qXwHcGmdAFRmSlLf/1SCfaylgSzNsWgMRF+tGEqNFySrRQ
gf909yJ78LYs3KlYeBjf9BjJJbVV14mXCPg5rUzjiHIZMkGAgw0a5v4oPPhASHDd/iQJQlspQD2w
HRPzKnboe/GYdHfb27tIwyEO1SI1Mzi1PYRCvBcfdM+7AbtJ2CrWa0fX+Ze/cslkFGH94Vws6ltX
yyO5KB2hmXsk2qFVWdBwEmJeqN5HT18V+uwNdC4upPV1zjaZyoEjE8eAS71Qx3/s4I4wP4vy7cFS
CmT/ZYjIF3UCh4+ANoh35fEUwPbUWCvWacSzXp1o41L9UolN8rhAbv6abzSBK545jpTuP/KU04a8
sQs0olMZPEgHBoiTuPrje20gBeKxzhg2Gn0dDu2GTL0nHYAz4pdV/YjdjmD74acpW/UhPoou3hiw
4md8BE137u4LiFvG4dt5U0uvUXm9MXCbMBpx0GsGobUIheU4sRgCv9Xe3DIYlkXE0i/1F18jwFfo
j+dSxP3tAOrx5EAcMh52hiOxag8HpPNLhbC6nkgxZXW3BJEg4Vfq8FNOxCcsArle/SOH9VlSqxUY
4TvyIctICFwNJWCvj9JSGW8ttXpftLIsgrcTTbwIWtJcpfsX2aaDqeiuymJnNhkK1isz1WBHdNWI
o4UBW8H8xj0LAda7lDZcBUGhBfrIhELA2881V1cLGLLOvpXcBZZJt2jC1/qvkoWu4eZLCRIH0QOU
8XUb3pSbcBIYYrjmnWRa+ROslYLm9yTj5tXkjCD5qeNWtenftBwYsW3ArEM8i4bRufmh6row61tg
Gc+pEIWH/uItRk2QuNqikwA9p52B677ahSYrSKLbl3EzgVE3QQGvNokujslKzsB9FLvGFXj9SNVQ
vg2OwgI4SPaYS23+3CWYn3iJnTWdbBVrvExlh7FdPk7HxFjgIc0zJ9EI+jidn2URZmeaNCmxxjh3
QtrEQm9de+mkoB/tpjEsPXehAys2E6PtE3zYUgkX2oZztdboIMk6ifCpGQJ3aFzSX/AbRgF07BAk
ogNB4a6CDkD6JrgoevuTjdOdoYdHTJBdZAE6/ynYSW6J9ZFPtdJ5ZwCZqXRad9LkNyInGVHtKOKv
G38NI4X070TVw0h7ZYwVTri3/BNl6n1Q9VoWQ5yRskjEmTafcGNIdC7Q0PVby3iebX4QJp92UhNy
cMLEo858zIVFxKBsbqdhIVZ5zvk3k8j/FKOlHrkOCeBXa1DGXjSrMihXFwCFd2imYhE4DmcGzn6Y
QLAk9XspU1RVFb5tPJKnR/TXlYVDT60upEknfyxZPTPQjJZnZ3oOtl8UvLNixpyHl0PMhwDt7DA7
oTzIV8gv6KRL9sviKxXjyAZN9TZaJWo+ZeCB4ePPC6WFO2o1wj58119WgLBeJnjLWZiPfndS+3Kj
pHi//CmOj2dU0Ns/TmFgWYXDu3D4YTkXlCZo6S4Nuhn+3I27QjNQd3dcdF8bax2eVCIzffNYD9AJ
Ely2vanHrwPkvhgXv/3aqs9EzNws+WkC6/YvEz+jEfItOsjAHiKkzsEc3ch91kl88RcnqOX5G2D3
/JkX83lx/llToWBu7ov3v/Bwf0i9+DYmyC0cFtY5LsxSoEX35nDmvOspAs+lH9pQbI3B5u9hFpQA
RnKPJfQc4eqGC/p9If/gXpVvH2dGZcPW0k+Zg3JJhRoSA77YRI8LybxyDp9TWpqkfBINBxfRe//Q
SpEq+f90aBU/xB69oahYJgXZ1xzfH2qEJb+Q9XHTEDVzHw6DDHN5fl0x7pL+iyf405lhsBK/3WFi
KdALrW2xhnwmJytQZmuNgJ3/K7fcVmMwcGqFToeit+SBwhQS7ocmBqMUv0Eb3mRuhc3qL+IEvCIA
dUubToDAduFQYezQxKECYhgSbZCdP3d4nOZ4SuJCm0OaRay6IZr00CjkVGaidfpurfs649PtMVvz
G2FCzgxW+XAUMZxFhJD4PyjWXNx4ha0iV9KqAmXtlS+lKKODfIuNM23P16QvjUkAwoZN1N/3hPnl
gj7lB6Ga/ZLWyl7Ivbk6/Letv56hFljq6197/F0VHkWmk9pp3fVGuMZYGjId4TqReRmI3cTFFeDP
z2O3uqV4B9u2QthPSLNJDs0mK8gg1A8jnLrIrTh75EfQugZREY64TTdTgGTiZJAL67QSMqzLnjDs
2odTqEyBC6xaCqjUyBxauCGTUTza3sEHQH6stQ02ALSdNhyzfUvPTXlYG11o3d6kznlzJ8LpPhRU
jkQ/rJAu0t7K7hzx4Nu+IGAeGxw7XCIk+L5cgct8nHNZ4+FaMNYC7lQk09ScFJc/+N3wjjx4x9hV
cS5cQdzQ1lQrPZuSHXCDuNANYuzKgjpbYtdqi1yS7BJ8MoU9QBkAmsbO0xD24WUsBpfh9ToMYSwk
uyZXoIPPEufPFoNlEifIwotQ1PQqdJkxy1HLfCxD4MhhuGa44UgfyqU+ctj2b+la+xzE42JZDdpz
GzCUZLZ2ggiz7WUgsgHYIdtsjPlC8isuYMgJ0cl7h/P6xpYkl0eS6Uk4qdFnY1/Md9Qbm04UyEZ1
gC5sZk56+n6QR/DzOmoTk+aWyKF0Z4+g4W0OcTSjSqC+mcfNdtxV8Bn78YrrW6+s9l/tD6i9ohj9
jkYFDdefb5/laLcj4RgnCZyO0LCUU/hAGercC7hLm3C21+fwPsw7T5SeeYxMuOoo76haf56lVJMv
LVLdN/QTDNhzFGePu6gqMTj5pFOMcQ6+0RkzPqH8bUhk5LcC0Cb5Xuh9+r3+RZ7oWQiIQrqc6Py4
kM6ai4m4PiScqVvPZkgwqv4eVaN6SuGvGBQ27Z4UssyIdsgojP6I+yFucurUC4UQ2RTtHXlQXi8A
o24uZJNYJ0AQ0qQkp9J+u1U7rhvbrvBoMAVruf/F1ClDEEJxHKMtbQGciS/8Sw6A3KrKNGh9R0Hx
8NzmYHrQIXkt6T3RRfiPI1gkCHdbbnSGZEKq/bzcfXoAVp0Ujb0vwYBrcH0lm41SCZ6DLZsdX1n+
/YSzoe8Hu7c3Cmoa8DK0ow/J1klCVZEv+pEjs6iqmDO9AxKmvZ2FlxTY+KeijGAcRLjb+KIzFOEo
Dk8mRizTYJTqd3BJibFrZVDXnV4De377OMj/YL7hqkef3xonuQP/pW0yxReHHtHlSm684D0S8hnw
/+haM/vXlJqjCus0YWCPCWF3TAgn6w3xb+eipO4I9A9aZMMXCAYtKJ5w/LUgmjnOzYgqwsMLFCLE
KkKlNJfmKzqB7Pnbua34yfQ+qTWDkMJyjb7ujv8mwusBrsjM+IoJysd8ONkKBlg1mJ+f/SwvsvWu
jvLRc7Hov+cdtlz32zFzvZou2ezFWtecg/u8GAxsvMbvt+mpb0t23/8h5w/dokUHi/SBKFKlfoKE
ntwhJo5KSGu8gNKZUXVDhzrFxnpmyQdS5pNCBJeuSdk9YkEy5BLfpXc2Y8pzNc7FgOa91YoteplY
ycrfkVRnziZAvrokNfkFRDve5VWczruOY0edOE3yOggH3gOaBoQARdSVuQI7dMDsc5qD+aAO6N7c
b8/jwWymyxJYPguThvqIs0YpJnCsI7kRUqm0LFbTRydFCZHIxMIFEfB3XYArkp9tymx6xMsLwp9M
oT+TB+24BUxSki77Eb6KJserSV021Lu+n9ZcUkkzlmx+IksrWakzct5pFpoYQTa60QpHavroS5qK
bMEs6S05AqlXn2+/SCe1sAkYp7v5q+GrXYOWVOdj21/smnhOZZVNpvWtWg7wLPPm5Y0AVRiCa8WW
e05NOGbT7v6UXzLrHc//fk8gi7ocLfMx4xuU4/FbTM3TpwZRiaOwm5vj/JyTP+TeL2uL5Vu79MTJ
jXwvIyOBXYsbh1i60LMKjplbm5ZCzc31p9xn3NtcQ0cY3DvA9akByWgzkrxxn6gOuiZjZJUyEb+l
ktmnvg6DybssE3RzAaXICuPTCbfRD9V/h9g7VcHlIowFKLMWLuewVA8CHmIttoxXK6SqpY636G6d
M6IchYLwmv0rou+oSoBCAK6Ifc+QhinGtShI5+b/Vqyh21UhImwnqTDro2/cj+aoUsuNPi1TLP8D
c/J+urvhiZE2PtSeHWs9lzrxhZ03Kfv8DypWMHh9aaECUjqNKN6GVpkuH/95ApM1Qx5smRjZlPf8
IyfJCVYw60UhB8LG7jk/qMOW2kDqiVZOZ785K2xZR+JU/A1AF2NFVGfvnCbvzsW71jtOn0p0Ixj3
lEo918wh+lnrzGjGsfZ8F5J91Us6SleScHN5eMZtV7gR8gu5RouO/Q+J+n0/twBCrNh1HKFY9uVD
GbLUuQ4CkaVWUYxd9WBxyG3hlow4jEcIm0HItE5lKnuXYPYS+q7JrRXNFrAXgvMeOPkUAkh5SF6c
f3vUo3VmAICqyjyj9BcLbDHpxQ6LHZzV8wurrIVxPdGPStZTkj+nns05PrQ3Bfpcghi2mfkFV35d
t78o0n23jWnCj7WBoqW8rGWf1Jg0WIxsQPGiPM4e6fWhymBTiSzZaO0BQuzNxsWqpj2yLfp5E923
HUbg0L2VWntovTGIRrlqjp1XeLSuOSEKOxUKFkUFO/2dyF5FuB7MhgtN1OVkbTbUNbDe/pDX0fwt
emCMJmW8wYEy9CWvWOO/3HiOtaReRWK6Rl+OxtEr+3CNY2BfQBOXFikdn1z4z8zdb4VNyzGp9LVw
F6A61BnL6i7MJ76a/y2zR2lcN9/e6e4A0qDjyLlbfSj+JURs0LhXfCnA4C9++eDljWF8jX8ayCYa
kPg9lSTJyYMBYNgFzfWMlU40sXVZMGkdXTucMW3u6Nomd6NIoMxmH+Nrbd7bYmJ9iGcu7l20PDCE
zsPiOXh9R8QLIP/zfrjzEfrLWnJYV7Zoy0bcsWdJIE5AQMxxHN6WzqdKfQJfy540ZlAhUfHkXx3G
eSba7h3nZXt0vzdwP/Q+r24BzO6JsDwMLTbTsZLAqZciWWSFVNsUncbeSsh1MNdXbz0TjaUCvWRj
l6IX/xAQ/hz7XK+Ktl1oBjp/d/RKt++bFo+w70B/mOCXFAUrNsStL0XsodUIraL6qoSOZ242WYEM
4AbWiK05QI+ydvT6+LCqyYMeffbcba64BPD2mZMZaRi3WpwH+gU6UCaFQBH68L0xpfXIOOV2bxMm
o6b0Q6EUhGg/sC7xQQqj+R3kYFOCzE93MFBKL3qBLmrIxQPJbLUtBSC2r4a+YG1R+R2sTnsUJgwi
GkvspjSLM7HsgKyEStfZMyE119nmUAZ4wa9nCfI5C/r3RCNrnjoPVtSbhnrzlPaMnJ7rEqgHZmEZ
FV5dzXvXRqloDezEWOF3Tv9ROGh19FcCONS93xXMfxH8b2mGQxsj7dAxqrSAm3UwivXopDWBof0H
qziyp2p1y1IVJPx0LKKZFWl2tmnEwjSv6wgNFcBl6UUla+Zp1VGnSXLRj/UUdRMEFG4ZtVQ0AdR7
2qlLvUCjfQKWatnWBLoma9yWSXS1C4YoPdkfNVUAlYMCAtK+5of98ZCUyYhgxk8luQz/FOvEQffJ
4Ua3FoiVd9vhM4oVF8z1+9TsuFy2BQtZfO8soENlhOobD/AuyJPttK9/4aJSOwSQt1V41Ahm17i7
aMhvNFpdszyOVqV0AvGvOsGvSx5wgTqTKeqDOeJtw2MMtWGOVRaiKMOYJ2+yEAJKE8Q0wPZlGYeN
8bzZ4IqIHMbNdNZ4dLK3xLwmDXfqP/8ymxPUGp96SVVKR3bVufU/pijaENvGrTbLPvuwKh47Mqsa
tvjvZKxNDmp75jEVXRmlkOHMqUdngQ+JrwJKbZFopJo0IB3PlCforYlFeg10+nYRiGYiw0+z9DYY
F215rUAkGYs3YvbMUMQ6Ga7bDOp/cf0fSNez6TSA2pRt6vQb7D+crH/8CuOxwG7enpDYEv/tmZXN
NwWdUXagtwJGmC3YMCqAPlP8a7BsKRzmyN3mqyCP/xX9bUDbxewN/aTC3n69xRPiwDRj4ZHQtfoq
tN4p9WnmI2dUVklHG2FXCPgKPcufA7Vq17jSx/ch6ESwYkFc6KXQst7nI2XIkgYo7UxTxHKBOvc1
nixI1eRpm7BPRQWQ6JOdw7cP2itvBwBMEKgpWkL4a6JpQpM9wrXgr7/GHdwtooiMM1KY19OZzLem
IBNHwpD6ULpm/Yi/Fl9HRjgNwCYdPM/h6OfW1Cj53vJFIw8SQRuId1SDygX3rVFDLW+55Kr2fpUO
dumq08Wqto1UsibJciHG6S0wrV5MpBA/vDpKFLR9kkGK4/8jTgRaTzu+g1M3KsdpeDNRvRZA/3jF
BSpTP5B4DNTPUVjGRdpFb2Y/Jnx2DDpzLphETxEJ5NmXcuKzJx8GyVhTQj9kWmdoSTdseNFPrB9Z
tNSrGthS58QqE60gy0rA+sb/YU73CYDFDrLIcpZu7s0L0erTj9198lf9MCDC+EMx/ecXbjQ+wUer
nEh1pIjKr5FcU9Zfzvon/Sbtrf8ruGdDEXBbLMtz2UzjB0Bt+ocULiZOK04CDdIJWtjZMBmigyJa
dx38arsGdN73qGlDXRS9rwTuycnxOcJxsyg3htRAnsitQM83CEAJWuzJmZjnZ5GFKGR6ib5KuJVE
dIUM5B7GPTZqyG7GSUz9DpLJkqUo6+cdHNokdkxcBnE3X1lHDP3/N5z0JGxn84r2gapDiMKD0CNA
mAp7QH6I5uVY5C6Y5OERT1buJ9rfMkX2qV0gNkgBO6+JjgocTIixu6IzdD1REnHgYTUWgl192aqB
ZfzhsKfxwumLgUdOFRgkA7uB1dGPHp3zTXJk0LGVeJcvzE/9YRPPp23HBFVhwWUbL1xaB05PJgnq
q4ks3lUZFPoDE2LhTxqYc+23K7AVtcoxlFWavxny35t0QgHuJ4oaNQeulQo0KNiv4iKiHAWxPQvD
m180VC8f+BdWotPkg3RP4ukNJ6GYk/Xqhlw12B428vjUiMrWmOAgJF6N3Aop7yCsjz8kWCZYcjzX
5x5hR8lYIPTxfZM2WhX8ohVmPVg7x6VPQCH4puqAklUylWrzCDBUV/Nn/ASR0yjHvt8biYNAlLdm
iyRfabbhPvEdbAYT8TQNfO0NixFGasBvCLgl9Ws3633cQBcOLYGtR9WXMq7mlRv93TfFvY56XAhs
OB/Ngq+IYDcGIgyWzEU+Dv3BljenDiox+mfulzPBE9xM/Il+OJpw3QmsX+NPzg8JtiyiE32C17NQ
oH0h1rpNcNHCR4UeznhpSRuLSsI+caucQFxbwyQ1WKBfAwiuOJrZtgxMTMB33Xbmn+EyDoRekfxz
sz2IU5ePViPzm56Smdj2ETxG5eY+PxILUrxEKKzgtLw69xu8REgjPpmlguz5g3FNFNd21os1Pi9C
hkohmMh9WypDJAWdDEA4PHlYSNqgTAkPb6NajBuNhFczAD3GN4k8fbaLYu94XjpQ+DAV0/Dipt5d
5Th7raGfPlbnMmhZtwjiDMB+A9LqC/UxyUYYhP4lBBPNCPUsJFpP+sEtbfDRbWqVHSr9GOmg5/yT
R+pc9oXD2U7o0HFkRUD40ZW9sJJC09SYL6c81I8eKv4RULeF0ZaDHFUyoDQQA24SleOBeJeLCEQ2
lw376b6Jgug0JXEaE8IFySz3Cof4gYJ3eVTmrcmsUyrW6sbAn0yu0p93yNbQaqvjhD5xGySiFKQ8
ag80LKXDuyJsJFsoCui2eTyQMjbYYXWAxwLDwOKzzWKpF+NuLZILJhBdMFBztBToagYRHN6H3KZQ
COpZL167AykYiPcIOCi2IbJEV5j5bxI9lz3Z2maJeDV3F1DGccrGThN+HkVZMrbAEkly4abMaXhi
TUgJv4Wkw8VtrYm32i7LWq1JVQrFbi9Rlqwxb36S+BXzFcPqg9+bh+j4qPMqAOtbbALTc2JQQiOa
MH7iJLRR0TlMCn//yfzpPae/wjPOQ099fa//LkEuaDl/gJTdhd37ATKnUs1KTWkl9WlOnN/r1Egd
/czkGhPSDmlBuU6+4pbB3XSs9J5nxovsVDwr9ckqm8D4sbezfjJSqRCOUrwyiQp9u/8C+rVifn/c
zyTCsu5kVYTUZFNFkgjHt28LeBeaVJh66l5lpcfIHGMtgmagEOJwJemrvbSgYPzYoYwDdPu+Nk1l
jmRwwhs0K3QKNOZBmip7uMaull8kF1pyk/CBNoPzBw1XTY7SpJTTBStIquSWlVCrBxIFmSpTf6Se
G5CYQPucovlxfdOlhpq4lViIWgvS1ZNyVNMEtVCAuHEE2KrNYQmspSCQqQBJl21fi5qM4pc1J0x4
1tlwLDzMU9+XNd3QN6rmjml3KMlQaaIpb8Q68EgyNgDdAO0eSHC+3UFwI8OWYEKGbRBBb5M8To2e
go7e0kKemPM+rr9H6J6bVYDHpYmoQ6Sxjv9ORJHhzxCItzuc+FihElnHPGXdbOhYQfP0g0IZ5dtK
WsIlJfpc11ZVwo8vUOK4DCGcKfZYljWsOv/nZZfziNka0qFhWMZ4vn88apwo0wcZlCT95Gr6hDb2
/nKDDCZkGpPpR+85VTgHM8FB12ey9F0W1i4hW0PKbGmJLKZQ8VPYLeFtd4G4mHbJ0g+wZ7i5MWNf
+2QQldwjNi7q2DP18x64zFZebPvfxW6SZ8bMgZ5zGHuUsKCVovC6DIOMwuMLY0iiTOAxO9MBoNOl
J6n/s1EXkHqsjKXiUc9eo0LOTj2BIJ6zsOpdjoYr6tZRg7firK+wddzXIIFG7rc7sk4rG4ZJTV0t
dvrB9fFDz2ID7fqi2S77xFrPgD/qm3+vIyPAzh4vNzEdtcLSR4S9oTjbqj2ydFrP+XQhHYYp0wF6
Vuycbqq41WijNZilWk5y4mvOGQ/MhuXMCny2bQr98/wx3NVg9yREJJowSBHXopsUcTgbRkKy5Lgm
OuwhWRNjobnC4tuekDf4RSZ2UWMTlbAHFDFsMGMnFB8hMTFIXWHYoxtjROOT2mdULGFhEyYPiME4
eqVqx0IUcLqOtkhYqVGrzQlER8tq6mX/K26U9g9scxG3FAbfkmn1hKpJaYtoLp86csM9mQTQGHzO
sb7eVK0YOwPCJeWWf7mRHEJp2qsnD6pCfwI7SnP8WGAodYukhYAXr221MPhGackLnwPKsK8wxiGK
evB0WEkaw6m6jIT8yCGQmhAxwq3YMbFgnL6NfEzAjNJeGNLyUqR0ZEFg0VbHveabcidcKk3lLQFH
4WCtuGG2NcFy01A0WzRE94E/mdk7qzAKRalgXw6GpKqXRQiFPSYbkdisqepjtsX//bmsAn8Ruw0o
CmLA7VEgJwuLtyNVHe/nGWwcdfsbXkp9ag6gvQ8gYOfI7O+J7+PM0dAVPVB+RpuuoCvGqowknSI4
5x/9Jx3VI0PehGst7+jr8lzZFW5EvusSh8U/F7JhdUQP+68PtS2RS+uZSdFaYz4SzakJUE7JjZCC
30FO6MU7MEAgixunmQSw7nx6gjUVYM35NchT+RPz+njDuwkAucniBzSIrQ2guxYLxAqDS24tnO+G
0v3spnVnJHxubCQQghzinpY/oZcSg+TsPF7EICTdOXJpfKxuvAzaFIfSkh7or6iHKbfbOPvbz5Aa
tSFxTBk8qCWfdwnE+8cdcVm519/nglU6L2eufxvyNWjg2GRylvLtNWS6IrppxX2aLHhKWhWpts70
q2leuiI/o5QxX2SoYnPvn5H0aGaH7KETLWbbXi//Y14JMU+L+5SD3x/0KowsZPHmDlH9utRZ4tew
EqjK0Dpdh1i6zGD3gHyptzyweK2v1s4ab0l4xe5WuX2aCE5RhsYnQb4tvFtsXxFnflzKqsSSsd5l
/+XJUa/EW4/s/ZbfW7ylstUGsI+//gnX+mWU1TVAUh308CTtLTSmxRURAxr6qlM57duDozrRlZtd
7FMoTU3byVi8Bhvk2wa9uQFItCU0kxKXcYL1G/4DbpkaRyBIi6FRELyHnwqpYAD/xPUh+8VpLcuR
IzxZRjI+sv4p1miB3Mw9ky4UQEEZrqovBjCDvwBKj0TzBWbQp2UzOazpp/scmDf8qR478dN17G/O
37XPp/ZFWjy2Ii2OApczWe3leTEnKCJmMuB+2IjajZNq9Dsk56X7dXZN6vriRPdaC3n3g3eYOeqy
ooh4T0admwnm29mi8OLC//9Twxhs6zmUrNbEyoZLh3/pDbfCgAaK5viKawxCaBpQsEmEKFPdXA7S
/xyonx8loE1J4x1QtK0vcOCdgQkeOXDE1ZFXqtXdUpv06FdkqzNUfk58KxKQFCbPeOOpAutT8UsC
j9plu5oDcRZEpbj7bQ6A7MF9AWWh2A6iudIuo6M0hvPSRetm3/3zzCyv0geLQjGK5O6gE1WhaXpa
bDZ/M5vZFnSAZbgmYay9imzdEeUF9ovkYgFfiiN4INPAFixVpPMC6iIatf/MeJodMGZzSdBGXUgS
TtgRWC1fB6nKqSpmYzyDIbHHqM2CX8qIk3ZqdrZa8YSGPTngYCurLBtcF1tQfTpbQmPeNMnhRB3p
kvPKd2eHCLaujDsSRh36+amMJF/oweFQhIiKdJ8jcwTNXAB7+J2zQYOm1X4z/pS2c3DNOGsvswmm
RCuhnAbUBC5jd/ZUiKtE6lCTPRUlnvE23xv5fmnOUcUgdxsaU25sZ+uNxKHrrXp0m5Mp1pa00wvb
6n6HLyZHddtlIm4AwL8aC3Bddz2u29EeQYB2s2n3EPfXOKxZ/MGscamWRu5KAv+i5RaVSZq5IzHj
rHwnmey70a7mr2YcGzMXYwgwTc911L/ISo9Vtq7jYP+2ha3+Sp5wXRWXNTpAPTh8gkW5/f5H2Zrb
osFeM+2v4s3fupZzDd4BEq54nMRzsitT8s+9+ouOFlSiOH+5dJ0gRcvcXMFx0IF/unH7TTg5qIRQ
lyUBLZeIvNoHqj50cpRm3ATww7vem54Es3NrhDt+4Ag3CWz9Azl6c2BObdrFxpCghWWFlT66ym7K
NAw4KzEdLL1ZcHSnuisB2O063C3OidsHSqrtI+GnnoqrCaE8pF8h6fzuPlGzJHRnOk8ASjr5l49p
qNJZGUPPHfRWu07re/2xq0hH9HUojn06VIm54IcJ5hK0DlDUQGSzLc58IO2tMwDHHhIEf8QfFq9u
WXUhPSlUc22uNuutvNYbZC/wMDp6CdS+xU5mlMweTeUIjEgTamdwpakzGKpLLzCQJqj9eYniE1bJ
gaPhRvEmdFdjd6X6TCxXWNTUstUYDWlp/7dCIUI4Jjg/HgF+EDLGIlz6SNj1ftZ1V0A6jzW/5uoc
iRMLfRkQ0nNOIBfLGiibf/I+G3qldeIFW6AucN2C53okQr1pEPZCsn6uw8nC8SWR9SXuzc1eaBXR
R6pxzOGRxuvrMTWpHKQw8YI0tEyjLStYGFBLbFKkkR9A6RvXi1ShHPBswNC2fSlIEzBlNxR1WjtG
c6JExu6vi0qsTbeXvLn6/KyIxcm/mDpWRAr5n8vyBaFAiw8gkmxy2Bg7rUxn1la0OI7aPpNvhJI5
MFSpZ3gcTJQ7C1HiXUEV4JJxRFTrWG1H2tOQKNq7E3FA0dU6zs9+2xWRNPmue8I3xjcqF9/SMAd0
SAE0kQtWdYL3TYzrTCh/kknrP5q1MrtNfBp721XpSCjaCge4SBwMIouz7EjpFUMqkij90kCASta2
JHmleMqnTv1wHXqMT1tsQ9hnu4tFqqB+4Tsne/KuMo4wHeQlzA74ARn5XsFsyl1uU2pbp3c8u0cm
oWjraMmzHGzLEtmpFd1K2p3JH6/XxMn9YLo2dx6Z7LpY+1fRgGp12jjdkbNp6kQsvO22sM6OTf9J
lTRIGKI5HunLu+QVhWlf3oHj/ZkBIGRt4NOcnAbIK/Z8Wcs2jVjc+DEfYKXXm4x6+4OcjqLQXdTE
p+BV/yvi93zxMbqUTQYjvw0YtoEKplKtZUgq0NNcAL8wu4ZHQkkcgr/1QTXcdNf2tV/GZZS+nsGc
ptwbf9y+JaU5suRdFH51DBHrGEJuzNTf0+7zPactJVQKhC4ATLPqJVuhJkqBZ/zvjfpcCy69NUVO
iJqtMhr/6gTxSquE75jB8bc9mqTY/aGF8Hr9QNBRb4dylotXPFKCniga2lkwYcX7ZKKVDOO+Zcos
nqvyPXEX4v/x6mu9bEMoU3Md6LQNmAQBrlNlOaD1VKPSJZMgJVHfRB9aPifwjvlrffaUAvmOQzMe
NqkCdosT389hVARAEDItjy8Yv0WFwRGszHCbUNwU0+fOROH/fXlL8tUOjBikT9QpbyXkj7MogsYH
OjQkEbTtczKYoJ6SgJXKeQ6d/wOVwtm/22ZQKnEQQGpWC4h6UPK22H2hQwKIcHt9XpBjH+SlWjLg
obfPU/x6h3vlcHCi0o9kIsOI3uhkZRnA/Z6UmMXfbHXhS5m6vIo+4rn7qhdymPqr6FV1EIIERCTF
YQlWsIa5Cs+0ehY/yGpfjdZwa0jaBM+rBbau5izYRFPeOvTaz4TkkaDWGhnyP3u6LKu2bxV7E4/N
lWvCOEO3oSc8MMhL2oMVf+1cdCJofS26TDOazCV6jjmC2bL1gtB1ocetlx8q+UtL+LqaCQSmUHP8
k7ciOZhU+BgmykKnn+wGIKiye8/FX2Xr68B3xYfj+GrCcasuwC+67ocWALb6pgDmIMivapa2nwQi
W9Ec0dTQeiATu+cbVfAnAw2LPc7XBaBlrLKuqI8TclFoDEXlNRi0JOaomCDc48bvcUbK3/1dwMEO
ImxtIQC+4sZeBkdgd623EAoLAKBJpIuO6NIocl0vc6L0A+zLvwTiY8z0S+uz9PUdHdR/6NkHhiK5
OPMuh6O1Hvg/0RbWJMhEIK/v2lq94jVR8MG3oDBJA/2/dAvdLTBUHjHJiiN9ykE/D5pCS1oLRhFD
+/9z3c9i4YZHqLyvIGBk/hrxZv2QZd9+MOrhocGz6/NCVVDs2OsE+96b+yxtLHjI3t2gVlJmn56D
6mjPeGfO0H9SepVVU6xDLrCWDlBC0yn+rr9/si5tE94Kc5QrIRDthyz39Li6vZ6J54CJSRmjmX2s
0KdAIqk9AV1GuaguCpsDH4TDt9gnS2K3RnedNPEy4bl52D4dQurSZyaAGedh4wCvB7tY0JKazcdI
5tORL7I5LqYNxWFcg8SRpjwCV0xKoWYeBoSWs/mVJrkk3K8iYJZeE0hobdRonPi1ZAP77ju59pn/
giKdvKzmgLB7t0yd+uYWzP1dhs6X18ucz42NJ7RhU4GtCL6btR+6/W9kyRSWVOFmiUSMvPnt99Su
Bod8jKuZLMuHdmAQV7BP0IqUemkIPLkGmtotjfd3L4IZQif/0PlBlxLvnmpHbm40MwaUAEGORGKF
bx/VXq5B5yraR9mrjvh8In/72NZlXvm14M40CE74lbMJBx5d+BmlG85774+qjvfA1Zj4RJ7EqTOp
0Suq5qxv6OWHHLwIDjcnD8Zh8jGiUelEoIo4z2a4ZOmre7xdeT/oP4Rc7XOn2Vi1WVMV9wB3sF0C
qQRl1knLuyT8QPgiLEacKfE0uV6tUh+mEdRVQyBeIPp7ugQh0/WFQefwzLvKf35PlYDjbcoTDn36
CgzynfnEOXwpLtnIHjDfstxl13ZAehmdWEIHwm8uYLMQJYwFNQavT1z/8l/vTO33Y5TGEiCaDKwU
Fb/aVr9wYhdiAz/vPcG4fcj7nTr9L94i6J6SzI1op/L59ZK6eeeswjWZdUeYMif5CXLSx3Xvk+xL
sivVJQ7kqWlLVfGTsbZgnoI+dohb+sz6qCOpEkwtMcmwLxccYbDvYhPxZogBPA9TB50iEQQA4qbf
Oq6kt5SOGMSpgRsVW9oSmlbth4afVECHjo3A4FcJDUqgBtg8B+uf9B+bwk13g0ukT45HCUzvlQjK
uNHEYiOaHeJlmtATCqheruC0JGxaR1wY0S2S42wrsXrv6xtwmgidwB9TmSlZ0KN9PcV5DUvSnj+v
OTWWgt5cc88Q5RljXL0+/NVszfkqEpETCs6+SyzGPzLBI1/p3+CCI6flcnIBpTHc3Xf66eXpq2bK
LFaRF7Xig8Gbpjgrugh5VAcJbJfByO/2PHPNTYK0C+7ulcqDaTgAn/rJE3WmIdh0wRP9VR6Y48/y
Lc1J3salM1jH84ZLj3Ay4H5oXuBF0QT1VT+7Ebdg+H/Lh2anBDM+U8gwXzqdOcdmB97x5d1+pKPh
M1j/fsH6h5uvIcT+WIKTZ4QhCXn9XFU4L5NkmJbpI4PUU+jHIkfo+qaxbFp4RxptJvN1BS93Icmi
Qducu+ry19HYnRxft9tSRPckQ6OIiRNbrSYnAlNiNhBa51WKDeprzlqad926EzalmZdhay/j8jBL
Y9CbneN7Ue/m3Ul3CzUu3nfHdsrdv/Q9lHXf3r375zD3e7I9fUsmbywzasQTyhp0ik6VR3TudRq+
HGSbAM4THgXJHI5D5a7r0rQJI/z1KvGHVzWU5GUmAJSOaGk0XWqE8Avbo0WGHOyuQAOGowkLZVuS
r3Er5XGxAaVjF9WgQhzRjiHXudiQ304LjV8SFGoUFcQD2dfi5i2Rs3oZbx8gUesJ3cdIqPYXlSZ/
YCFwiAq+L9cFIjayJXzlQmbEUERh5nLN24mVrq05yqkB4y/5V5RWHY3ePZhj3xXO5oFpY48zZR8b
zOP2/C3Mm6/ysXqDflcjP68eImVr9bakUF+W/S3qhycFI7rAYgeiOTxjYdRNp95hmysDD+WkSI8z
gNBl83nq8Alkg15jHsCqI43pXR74yGOtQEOiYrpCaq/SVWVY1z9az9IAk0dUBQJm+7F1sNhY5BBp
9m691To8Hrza4Cl0w4DME/+fek1Bt/jjp55elFBbqUHs2SeuN/W8j9dwmdzKwMKMvImJ7BEBGYVl
EQeJFQ5uAEdseT8kt/o8d30DacDjHKYvjD0+12iXDFUA1XXAMnElZsAItBI/AQS1hK4Sze5elRuj
0upILY2QNXuVKucmgKRxP/HDuoiYGW4OD9h20EnQrNp5BChZqHq+fmVEO3k5evfTEEwXqeAsg3Qf
NxgDlw0kAf+u7U1dTAncXFO6ISDrDAY2cWgwLosl2CBqXtsIpWyJhR8Y+Sb20pumGSFDHZ7grJdE
jWxIoIKTOzP+93vOzjIe4jNURiZue3Xoe5kmDt2RTl4a9MstcrY9TH793fsvA0v/Phmjcw74+47u
mqulVolJ/AN4bwThpAxv4ZL+mxb0VOjJM2QhBEK+zJd6XYf9EDAFx2p5V8tL4dCSAVSeZvbWSCSf
iYQPD2F7b85a2nnLlbG8g7PTO8aRgdueHtKOVtyofPgOtvaOyX7DK9tS7Q+lsgiQ6O5AwX00jaIe
oSF0IsVqGPBu7kQ8FeGiKkU1MO9MtMz6q61Qrvu8tPVCid7+tp42SCvl5pz+xawsvyhgSF4972o1
BCu3G4O8OB1OElYC4Erec2uDa3uJVW7/6MAOqO75R0zxMulMLPGEApbfmDvb+AzlD2JIr4PRjmAt
fKVfeJ1c+N9D3qOXKoDNbqQVK+Fx34RTpXqQyhTZW8863JcJvU8/eiru15AbgPSP0M8OwQZd2S6J
3/uzbXEYYr4NU64xWRqpYHsRiCPLbzKuEOvNiM3uQI/98uXRpD5jVWtlwD3Q8QGSsWdXQQ2D0dI9
hVMVvwFXsv6gbPE+Bf+xCGg1rPlVSF3d7rRvXNQLORQf8hjYcExl400X5bkOBjKU7kx2uLusOs+6
j89TxnwikgW5whHJj3xHIQ3ajVvlovFzwPtU3QD5xM6lF/zof8JAU58gKswSfw5SJpfAzINwy5nT
apRZr54WcNa+9s9KzaVBX2cxcDQlDjClmBJW8ljTBL7oRKi+I1p2bjJPpyRYgA1lQ81zSSrRASwx
C8Q97l05/yfkfpN8bR2bbvEuFLwg2H4rMzLHwituTv6tLuogko8AnlOS11ON0TyHGde8PjCLzfda
AFn88hlwiDVp2BvPNC6wSdQPgCgvKTx6Sk6QQzFYBr2jV7cF/T4lTcN6j+LN7WG35HvApYfiQph+
8NN6Dl65r5KzOgSY08+NggYOep7ZKDfCTgu3OXXnXhwUFOi2FHwKBTAhrVGrVgFP6JQJvgZe7RDE
p3S7wAAgIqnhz/rSeOpVOBvv0+puFptmyovZNI6R55ev1R5Ew9V4xlq+1X/LSWCwg7jaBxhXKFiz
4nMi+g46C1SPvT2B2j99CkPeB7M0NT4hbBwYHr8FBQJR9lcBGmyx/tmHXIj5iIjo6SLUKFHH24/i
/Ji0v7jhlRQrjuDN8JmCNEOfM2LhhmS2ZIbGax0sl3yr9bOOyBXKNDLd963Ocvb6dQZdhz/u7vfh
1B5sw7JReFEVTXfdNLlxkbgxqKb8QE/lt/NvvkPRw45jkP2kfGoeW/x+PxSNAMoH5Z6LRkpBaEff
Q2xwOzDMQM4JZGMI2yKG6E0qjNWJQICARjt7uqvkOwPNjnDYys9pvbSYnEw78A8RUPDNp1Nysw+C
cRsyl5qy+PTX0wfQijfF7AMHfMpHPqmwDoBnMacqus3jJXUaKPzY2rHuXK1hDRbaMUo9kJkbnzJA
VUuzhBBYUnMaTpqgtx7xnRkl9QF9NPvs+pDsfCm7jbLvlVlTTvT3iGrUPthssr8iYx7K9SOKIh6B
/7q1uxs7e6S3B/1KhmtWuWd9VOwRHYfBoBxziYGhn8i5GOpKSHSuOKjFXaMF6xYzZ0GFytNjlDhl
O7U/SuwZ0HOH4fDytID/Ol4aWjTkg2xEtWCV2VzT1Dt+YX4LcSKDmEEolHIQ7IvNvz2TH38sG8A9
G8P6BqojksCSxrOpzecNV77B4lyBdiFI97B1H7Jpijo2W0QWjiHvGUr8of/nMDd8ZfgpQmMFtwQA
FnMIXqay/zMBhmW6w6B/hRTgT5xronMrqMH7Bc7twN0j+Su1H29DfbUKQubcUari4sKMlPSmf8ft
PRvZjom0fR6MDfAAmsyN8DIi2K7y1bYYoC899Y02h34Jl6+YYU5l1a/rBWJnFUqQjRw7HhPN7Lgv
Ig+8gRyux0peCd3PtqPJQgcMQZjCXQYNmTUK2i4es9zARebfbJ2S+XiRz9HCnMeHmbk1HCk8Ywd5
dil7TF1tes8QumOuV0faDp2SRHtie5L2tq0rLWkPl2pj/OJ+iw5rjFhGgUAV2OL/5HIxElYsNOcA
tsDaWnsSaZIwC1Y7AW4F509HqsmwzwwOQ5ImOOn5EZBWGhRebtpwUFsGcEkDcfjRNi8gybmBRIb2
V/+tsJ7EvppeIJBCBqsXWd0G5A+ciY/aZgUzCiyuU/WCiTFL9AhxtzFB+S9FU7QBIZ541Ov1DRb7
2N5FFeH1pYZWZgivrP0JEOWyV1ga9Ro9SJdpg6rh5h7YVvCBbUooXs8O41Vme2Hi0C29+562GeRd
8YXcwu2wuAqvxnof2xSChBbiuVVY4R4rc8bbyUlySCiPmDf8Up2vI3osnSscFK7Qt+gFg11cTVAY
UTFRQg/hgCHxxTfMMo/mkhCebrmW+N3yIC5Z0uXQDtS8I8nJXUqkDth5wFyVyBcmBlYBYz4kHxgU
YpA8Y2Ew1hQoqOfIkD1NZ8CcbRGeNDeFRfjMexd5DgzSC4yX3v1DMxzqnI8haQraIS/T5UBSsWuf
EJdMbI1McvC2PC2PSJgGaKq71RkomqN8hwmsAmheXmUu4pXgOVHOYg1tY4sZsKGtni5j5a27trSN
7+2nQzhXgPwbjAZplkNfk+NJRu4+u/EICkgSrd408JpGQbSTwLKezkCRnhb/NC1rcSj8sENLyPVc
ucdJqN8WK0liX3TZaK3OY6Hzwm+br3D7zEezBFknGYzhj1rjrO/yGShAKHTCYbz+o76Xws5BGrYb
5rSjg98HO9BPFKeHpMR4gQ8nQDxEdmtDXGNRhSQ56cMivsdmwhOyrUMbFXe0Tk1XnIBkpZo7ImUq
xhhheeufEinYe+nac3xNFNeBckh1apuMW4dwVIk6SE7KOdgAcVMJlzT3teGlStmuftzlqqUXOtjo
D3gQo2T5ntQOP2TnU7v3vrLtRJ5S3q6KLOOrdka13Fe1q3Fn1v1qcVtYNwsVLxBgduk1FgXhwt/s
+CgtZpjcstANSepCqn136qlWKv/R7EWByZ8IX87wVsckXxGAcZYYgofgNnc03ofPC4DDje7oJoU1
uC9CNKaovjNSsGHqnFA5jRI84Hmv7uHmHn9VBOdCjW0I1+Vdyq8A8o8knxLtAd4kZ4U167pdLt6D
RMFsEP/crRtDy+UntC+EfBhVD8RRKlKVM4PY/UivGHCP74V5JwuR2vvQg3Rbn1+0aRRyp7wuJnpR
X1ZIRXrrbh4PNEqe7vu7X4dYRXgZuY6hcJ8cGrzg7GsSxkSZTRltjss5dQr2oUKfxPJdxwTPQBVg
mYGHoBAOAGRzJ1xmY4sGp8TUcVRU1l3F7/dcKm0IdeCA6HobJ1QyUWA3TCDjpwbRy+5XvU6k7/ic
EsjE2x3UUD19BkfwNSjUv+fquaujP7BchcPXvXzoWtks79FsUSd3FOxnUVtEpt1ap/Wck5tmipmM
VSLkWw8H7+EjYnrfTZeiYCeM1EOxsZTDCPynn3v+svp4ahNQlY27ZWQfeVyLPZkfMEQH+zbqF9RB
hCN7E/OW8CjV+kP7Q56iGvyL3IQnOw/hhOQglAwnZ74Z8X/AQQk5mIun8LYiIjEjpge1U76B23U5
kTLQ2IofUOX7hglehqHYaYWOV0IE0ydz7w5d+y0uLLMJ+rDRWU6pe015IHbVhNpqf7+dOxwwZWQD
BonkMXpkKxWVbskhhdq9xPSiXxxecFd1OdD9qmumou+xdW6x8ViS402qr3P+qj7WK582oygduFY4
zKFE2xQqYSjRGL/4jIAYkIF4FXHoxOfR3fLvuJz8coPh53MMnUyZNmgC1m++8EFBkLBZVEgKBtvu
FQAO6pouoeG/OUtkAadNd+g8SHv3wqbGbKYll5D9WDOZXB1t374kvORqKPlmzlHe6oO7wen69T4N
Dk2Flzn6R9pG2XMBoFbFyCC46S92jCp9zsqClzg/0NCrcROmY0gjeL/bZ7DmUYS2vObh6V5hiuqa
hXXgsl+YF2d2DzoJqp047EYATo9BREpZdnn2Fs00M+a2x4yqUcb56/ewL8l1kuxkXBBhVrb25OqZ
hHVkcFAB+xTVxfT4rEqjwoDs6oLgC/Uh9DPk3VKmLhES0o5cAA6XIXrVoJFd+m04GA7xmwvP4A0h
6rW3V4GUHJGM0D6TgbRxyMkmcu8SJUR+VXs72SA3UHiSjIvWKPlIk6wI9IJ3IqSpO3QPF5UKeVBB
0v0P+IcEUgEyouykXGrxYVtRDQWiX2rZMNU06uRPk1341/cFnSKZD+dghsbWmwG9mUF7J8d/5tzn
YAHLOuPUr46l6k1GUvJVCygBdafKrHmbotHusUzLSY1/4YyLwPwnwkDAtZ4lgXhWaHJxOy9mXjq5
kv+AKmWKQI0Icf3nj9BI7LHKzdsK3HLe9AyufjDiyewl42eLz0zFE3/bDvK4MqnAiY2JH3Nw9d0i
ikirvIQDAVgc6GydSQF3zbphIxyijJkr2e4799i9QAEeV4QXG3Di4d88BUcR3+WlSwXu9vNciA4r
ftWiyBljV3HwBDMynXVNd3R2HW/6BFC+Q86Bdg1PD9J32A1/3UNVHRf5bUSHgeVem591NNNhtLGs
8qFDGQYRfL5RCSi4yF+SbP+G9O31RjoyRDZs2ESBfb6ieFNlbgdZqSIW83N7t06OcbNQ9YVOc9XD
Q9UdcqebF9VEUk2jkXjuP/V0Ih1BUjmmo7VtpkbK5GaOd35vow/PjaRIiIRMPo2sQqZuF+4pOAY9
MBO3UR5Ke98hmNf9pao0YfmlXANYq3q4lovZ2g5iLPcReTO5WegHkhSctcc2VC2gyubWECKGAty7
CAr49Y+Bv0DjsicSXEDI5ojlbf91fmT4aij5d/w+cpgU8+1s7mr7iL5KfC8E4ApmisB+YkG0nEN0
TP5fwuLEsbPw/wei/0+VuwaxGzRHu0rqlsCUbCnRC4eiQWyZ9BsWL/5yFza5CsGO9GMPRjDsxle4
NPbYl3Unu2hFxUljdQ6j6TLPYDZ+yJ96/b3F2X+H6dRl05VEpAaE5DVR9lXGFZkoCErwB7xaSjIA
MRAnI7wn4YZHDCIgTuSJVrvziOtCEY0ZSAh9FbhI7zLGW8ErGQpj3XJlW4/W4ZlEQKAyKxcHMxro
y1vORKj5OzeXsM6itDaS0fvLfmqbv6M8LjgC+mZgvZWwbzkt/+F0pwnCAqhcatHK+frNEYYeTuHS
J41tUecPWS5/L878BViQHG4SDVp+615yBfJow/4lAh/pIZwkt7k651uGK/qKszSb6aLw33Oj+6DB
9+hDIM+NdJXCUQawtrs+pv3MKsQar0gG0YCiFA/re9pnsvHMCxKznV0+GSQDhPx4B1Gq/YKUZE50
7HT16u6iWlowDhVuo4OE9hqqV9nRKx4JapOLw8pEZbLiugtMHTnDfNqW2eLLzm17EZ/0fgrVU0m6
ZhwWs1AEh2tBertbeywGodzpwxzVuAU5IWriKOJx6Kn88Xbtjcy/WxaCQ9X/VttMQCJbXa9ZUXy8
SOpC0lO4rkgW47amh+R/9JhiheJuO011aIytJBqLq3m5mjGEUkmfm4HeyZvBHtcQU59EEgapL84W
tHj54qEieqSc3TjuYmONn/m/G750J/5/jdcD3ctuTH/QRmud3OsFgPvmXW6o4rYiIcGTD+GBPoQT
+GdQV63kMJ5SkRISMttYk7LmDwA+o4hm/gVhY/Zq+gqEZem9JarDrbsl30Z0YJPC9kH+J939kZSt
j/ICPd1xsm34YTZEdoq2Z/QZUxsXgVj+1QiEAlwP0C+ErONLmcE5grogwULQwXQyIpHp1XRCqygl
+T7Oj+OUI9iSjtXWGMM3lhFGiLlV3DlXjJHOtxTvM3FRwAFjpRYS/HidU1fi9pq5v7kX9jKvF5z+
c51hoKfZDvWH3Gc8v74cwNR/Z/9sROEJOOPBtd9ief8O+LEIRw53cVnw+HcFNmKF3EZriOARtFcE
1RwiBGdyL80CV52c8fZiRdtuFxtMwO1g4K3TaxBsDbHBrfkzAQpv9WeQ3YEJtsS6iiSbd/5KBfzb
q/nfDJ8wqbxKS1NgPOLeu97E32jexn/jP7+2i+V7w1tHawTHj9Hpo8xU3WYUvrkcyUN1T0h8u2jz
nFN9oas4r/bguHn3jQDZhXJnL9knFvOT6zT+pV+03y949HgMlnFCUnSZuQPeHj8eML9/lCPM1fH5
Gkh23HBG0rTtGbVvlmVWGHH38RIh8sNjwLR/9bDOe/Z8CCNlSEByM7QJ636/SZInQp3P4fcLinz4
WZNhOayVkb1God08ZFOBsyj5EtdV5vVaDo2qYrjEc1ZhgzJaJVVrI7Mc7CvqhDy4mm7KHEmeNeFZ
CzCwRUSyZ49Uv7AmKR9gUjcLmyJT7ZUA0aYKhEXl6WzdTm4pC83EG6CQfbW6u0fnUHYXNDBdk2HJ
oBosarsyNKC0162lYvX2j1kwLGrkVIoY5uEzel4NFFTwcYsjeXB1Nm5XOC/+dpLbV0viWgAWcQlq
KJhF856UkgFZaDCdVWobKD57WDMplVUECLKzl8NYV8eX0TdxQ+VYjRLE/xBuWXnCz5YWZVdIgCxr
MSgfdSYrEQ8AOJ3c5c8wHzh+cTDXESvUhKVM4KiCqQiDe9en0qUMkZFCN9P6I8C+mAwOsLgZr4D6
paGYhLGa6y7Z+QYlyy83mZGCjmPaSLObOKaVaq/xB1GyGQBN1LCFh8wVOszzmAaavCG8CYJ1xhH+
DfEnbHfUAyCWbLcKPvsH2I3QgiiX9BQMGStT6VJSMWNV4cBlRlwGE3LObjQ0FRx88XpNoKjA25jc
TCJU5cRvBZYt1xdian/Zy5Qqw1UxeSJkw/utfBSv3BGMHUrmb7LgD0Vu5AaTOKomikaWJxNskfYE
yVS8VkJ7S+d2qXZ/ckKBAL1vv+Eqa9UfAQ6cWLRkQNAhcJgis24l8yU5ykMHVX9SbsErBuAtVtxr
JbdVYGV3R5umnIsMNbE6YgqRyrBA3SPulx0jB+TvR22cfzYitiNpqgnEkrdbYyiUVG9mJ47ZdJxz
2+b6GyC2Np1NRZSU3tcFDp8gBd2/8wHKnlO0YnL0qo0+M2jlseuL0htHnz+eOz55RFzFabjmfNw4
TsV6UDANz1N/PAPdWRnkQVBG8ZW906pmxV5XjIbVIK9ND5TYL6EDkvNp4x1RFXvnhrknVdUHnxer
ZQXTFfqcZ9LSlQPr4S+6eiuuc3+MfPX/MTpN5/oZ/GH9KkJmXksSesSsC/z0qsl50sTKHyVC2oSc
8Skg+TNjHQMv+aad9PY10SyPjZnMnvtNd+kUIkim0iCCduwxNnkddOwCjcMriF3yhufWYGwjnuhw
FOMEXvW6DMk/tRmzOSaxfePfTr8Fkostm0rTxy7SS6vAhqsOZPeMHBv23vkmSzRntf0Z95sEedUM
HFtnjbmTPgmXnLoXXdPTVXvGMXVZ1/VYKT2mvJdocsHKxg4udViSJaauaRlQWzIAfE+RzKN3Lu+H
YSiHtcJSayoxeDCdzmT+5jHws8aO6PH/qYp/IUrEmEFGrslYOuqpuzx9kF4mQRD8MNQSwJ8aXg4H
TBFXO0p0XSLlBcPkICV+SBbFwFwz1Hxv8we/3X0meYL7CwdWdu6fH5Jd3HDYW27b7bwSFuCOoC57
/pZIFEPsXVlAaWLFhhlxPpZYeGj9GH1oUL6TvWXN5KlQiKfw7iDJI4Ibl/7lV3FqanVDlyOaXBtN
nUjFJmqEjSfPztBX3Gnz9CZSDNREZ95sqcsail7w1bssi7lrTc4BVh/O6ADJIwcqhyiOsny/cTzS
JeFgFkHCUaMHub912fe0dfHHUxEhM2Qwb9YZ7Txi4LJsIT+CLWIjjxxllIaxaFhfQLqXgIcV24HR
3wj5Wjbydh07YSZ4nBb3gdroSODQhX2IdPUNh36cp7kLwkwGqFhy0eARQ/ygAGTELJk5XBHE+OK5
w8GJOdiVlwYXxBlsb+UjtLBuGtNVSy/UVDG7aD94fS7Y8p/H0VryudgWZlJvF4DLt60pqqcn3aAy
lavkzedgbKwWJJ1M8IpeFse4JuY/lwYu1EDa10DNn83euDqGfCsdyaTRGOWCtDRRT5gxjg3FSo9d
AD6wndRmE8+rV/DP1ENr26XFhebfHl74QYCi3WiD2aL1zMQTUqfUNlO1zvnflqoCqe5V+CzQY5M6
E/e1/1OwqBD+1YNCFVHY5tDDwoC3yd00b8onUDQkp/vYEzZkeKVtlNlTTy2ww19TDRKlt8+Fk/aR
TQItklvMhpawad6m6pkCvQ0mOLS81slHgfVLa8d/5WxIGuQ+lhyYigd9rZlgo6Y8mIWDnl1r1uPB
3vl2psAKmw9HaQaEGx/ttmgMZoP4hFMdf8UtH8nc9JyFAzPYky6lwg5KDnbwYrClgeClnAul/cCR
PxeG74FnqAtH9dWEG8ifJP2dWaPIk5ZQlkw1+GO4WbDIcoU5ZIj+kAM3AvONEKWIWw4K60c2NlUm
UGrWfZ0e6jAFidvCaXXscibx7M7rPXlnka5euKUEIBwfs97bzr20dEZZlhF1jTdYWXCC2MbRbREU
MwIa6DB8idH7N85wGIuV+D2Z5a9nOj/L5QE2WikMAhir2CpqBj4gWjGKlfeqcEoohc8nB2+T+lLV
5dKj6b6Rtd6Uz6SE0o3MskJ7NSTmVv9RCPkbEdk7Xwdx74Gz5wcBjnf+hx8Y7P9X/mTTbjT1H+2u
EC9MxfQXnKAcOBNFaEQ3a7dOb+TMFsmimVC4cFsJlh7Xx4W1oImpR79FSAuK825jk2yuI0305D45
7oKYRciXE1QZpiFLcoG8GnnClyVAXqR9iInrqMjJTpfOYwgr7WlXNd+cojSeIaX1fduCSKRyhVYr
jAoJivcwncZqwhRcp/A1yAO74Ho9Y7KTnOzBZ0Tjp72gfiGXIeEyAkbecVmQxkBnxcVquGnUmHC2
5uH5QqGcFkf9+thfr7zXCraRT6tseNoSb3RZe/eGAqQK8L9jHjdgL3GQ/H+nNkVDK0tj+3LryssW
zqq2ooyFZocA/uzTEjSmd/PaYiE9HtChKCGb4PdUxGkilvkay4+PE0CaMHJegVLg9ZipxIIdeFw7
YjppWhmpwYJVIG11TaQEpNbbVqEkh1rtFQ19A7eOU3TQwRnWcsSgW7KpqJsfxRl0RmbTeSWYRMcD
+A0GuoMyFzwuXDjDGim8yjFPmdHGHmCELDN5iQ1Zu/coYoI5Zj5NLfTM9KLiEReYGVBX1WmG+3Yq
MVz5+iexF1Y31x0E1yyuI8BHtk4At8x3WrAIDJb2d/2niIaj+H+uE4ZT/5IXSmiOWd0elWImOsPV
Uq+jzjmN1rihhucUxbOkd2Gkz6aFA62eiCMwWJ9/0DnWeDLq5PFRnuyA1AgY8kqc22/9y1aZMzm1
uIyMwAE1xrzrR6/0So4dnAMmeYKAyc0t4V2rA0QRxtA+ReKxVXMx5CfQ7SZisG8QAUNnIFtDOJyJ
lpsZpwFoHA4xrxPyuUIkSGQgjsOkOA6Ne6EZQKNZA3Y0hbw/Vo//jKlOrHqiKHLbQWKG41ff8q3l
6dOGA1xL1LAHyhiKldi1M905MsYM1I1rBHRd6Qgh1pLIV9LdFgvJO0upKBQ7rHGKG3tOf+1UnOVg
o833jgfXFQugI69qLZN3dvMhRR6NRTOLyFdnOqojuPfRkPKSKp99vYid4b45JUh5PUOeZBKrx7MI
nwh7vGvJVFA76GHbwhW/8Q9cZRcXTc2QdJv4kCvqhxb2zE9tGxSl5gt7MtaqXX4fgydj8qR6cmyr
oqzSzL/0/f4RHk6kDIoUBmCuWp9HWfItgsXTveqMK9qvQFdz3jbes/JqogbnsW1x/fH24fnnWPqZ
sO/P1ZD762Y6LciKV8tOp8s13sstt3qPChCo/C9b6rJqNTH1wV3N7zxxqysXOBNV0iSwLBhhVpAW
B6s07L5zXTHHtt3HJc0UyTcub1F8nzTUwpQbpvu0QhA5xsaLWqKBVeP52OkpOPTcTlPlj0DciSzb
HYX/mHCWcAob0Yhz4uKN07kiZVerC6u/tY1JRc9v8uXOcjgTl4ZeewYPtpecNJkuZ+7PXcXt6S60
5pXPoAftvWBOl/vnmQFC3/6Mjvw2P74uSEMI0LA2FSu2djZymuz7pDZ3eiik2roieUo4KmwbIOCM
LWMmTgYv1RJ+L1r1X4XVmUfLdYCMXUJbPWsye/xmbKD+niJNtPzAyNhsnh69csDhhCUoNsiKSy69
j/KkrsyFgE6CYXXfM7c5MoLLX7LYmdDd0fNd2i1tZagxmC5LWNwLUWJgyY3FhX2G2EBhzm5yjdGs
dY5k50KthVWhsKHN7LXz0RNk7owCZ6kPPZSlQYIyN5s08nhGuI4CMPTnnmuINvta1frxicE4OWmv
IibyLa288kTAvUb7ciEbnLL8EHAPFQi9kIq5fQrOKQzJYp9/vj4e+XMEl82jFb83vVpC3hT8jWoE
s4WXwxH2x0ZwLV5iShGqo/4bol5hOvxxQUwXnk/1qfj85UgFIP7J5IifR8i7B5RnsgdeqZOTUCez
V2BlGezS9lIDZIPsWwsvixYZQzy+9wuTkpQ5wHLkqpi7WA4Sh9u6lwCku/rNy9FxzCI5Sr4S7clG
OEDBrkUJK5LpGtwGlbqCSxJo4XJOUkkkc5KqNn+PR/E33EwXkVHqNVXVKwzqDjVg9nttWcyXp50z
m8X0N0dyPo6bFKPE5FRnHp7XHOP/4gVTNecEH0cdOWBwlboG52sPaKtUq6DSpzULt0QQOU/GyM8H
/xm72WAQOBdqH9Ebe0PGw0kIXnw4djV4FUxH1R5U15B6LUQenuwMsgSi/whrIxYCb3daJPkUDLAz
bEpvex9DGocDeXeuX23gN/t55U49HkZmFzlUlQABN9ZobVvBk8L0K0hSFv6AzRTv9NjJZjv/O5tz
gLavPcXquinvqucg8zkf/P+bQLJD5I+tcd+7Zw/CabI9Gb0ySuvCjpyemkTQIvwuG1Go1eimrd9l
pVP3zKfGpaCVjmuVzAr+kDN2OC6EJNt0L6j7wPtzlOvmTRs66qIt90fHW5832qMeIPqpGQhbSNlE
7yBSIhCpZLTaZ9/8h+wfRmCZpmTFWii40m7ZKXPiy8TqqAxwaOKy/c+IbA9fd3JjKD3nv+M/ZH8E
5N18c4DJyZ0+tOQBimgTTkmDOGTTlglQc1M869RQLRDsjvHYsHBBMVt+rGe+czMjUAukNqtfBHl4
NC2gtziUPD408uugDKWVEfvDy1KOlM6NGxSeLB99y0kLGhhQ5JmZCswl+qyNWLDF1Orolgp5sNJQ
OXXS3+bP3F/gbYUH21plDPRgRFVzH57DD1AcvMH+gu9h+lFHEfLos8MkTUoJzFl4G/0Bg9AZ3Q/g
7rfu+bQCv7s+nY0OrtwZnnfi9qir/LQ7Nht1nq9+c7jtxYrWWeMtkGFyigLwenvBviYqqaFqwY0m
aLkLuMyxiaLb/VrQN/KEh0T4IAHzf9FzQYBzqLxSzBKHbDVRVJzwUhcNM+3AaEt6YZybMtLnIRiq
RjNfuuHPa5n+nBBl2rZw+mTDL4i2Isiot5B7L6/bZAPoEl53jxWd8ipxRBLQ+bJJEUxegm+Vx9uo
1SR49901MOYXBTJW3drb5XcHSFdtH+wHdGzO2QwlOn/wTj/oNbn6ooEfhUj3LChsWKz3atrIbB9U
reDt830+VcwECaZV3Y8PQVDdHUYS9qIA3PJwl4ky42jmAm5Z0S0y51TkoJkTxRUOPH7fFu2pcI0+
i80dIZ2nrcWeRxm+bVedaj7/yJP7HIYwsrghkbzr52crb49Q1uFH2qwewHz1c9XibKUY2GhKVXRf
uT67uVm5RgDpw/WLwGtcXLMCHcGmreIna3xV0eq7ZobMTCLlRb4Kg9WzNtCgfKtgaQSFg0enDdzF
wtSkF8Pte+pnsJNekfG7/LNFdqB9qrJ6GJ36t/j4G2KUM314vcFo8T5XHJ/lTHF0HzpS7wMP1OnY
qAzc+kOSPP0+yAVYTOCOPOJ9sGHlHjCYkvNGxLqcE+UyiJSMz+YPxiX4rQX6CIz9WgMla7lWfcjZ
LU+NSjlJM0P6CifL/wmKKAEOd0TfhbBudo982I+honaA68IX1AO0VYiP3N1GR5Kt+8b5r/e3OKpG
X8Ylglg62OHBViF79D/aShH+PtGkQ40pZoxH7Zy20TwpqWgDuw3oIfo3he/eN8ugj/k46i/MtN5r
RPtqTK/6BUzsLwo2JUOww+fyfjGiM6xPE82yMNyRS/aDW6p6BFqPCQ0CFUWyAzXgY5YQON24Po6e
rJtqhjVj+M1ZkkWTpf5YsgYatuDix4NzThCGUm/PMdvOPKvXO4+fMcV2lHUCPiXgYx4gnuT08lR0
t+nfAr48+Bh94NS5iBFjoR34Hc1HL65vTxExlseQep6q0hon9Nui3O0A4a7962g9yekJoBWnfonH
tozoSBfL6dNjppXN+bIvnaxOaqwe3199LcsIFK4ubEpaPIGqGF7RCvKU0AdxCvgmU23++o5yac0w
+MJx5HKFdTgEYOgjO4tI8Hxma2J6JvLeUUhsSvAtlmSUCiqZvn10kM1xAH3+Y7nleQmcezJhTZ9r
pWoKuNJfdptKFznY50GLhy+3cMzdw3XwH4EpnUce4G2z5ynU2sOHWYy5B3qt/+VfE4LHVBLWwO2g
eI/IUQrEVSkQGjzmeym/gvgAVlfzgN1tihDczB0UcN+iVn7OGN9jGEkTfz3G41agAzfolHGUL0OB
fN6rlvKa5LfQ5GIacNHLunamiPNpXK531c0unPSgoYkWRBI+g/R6besh1Z0/VdqlVGb+1krhvfS5
YQP31x+g2Q03ZcStiKQe598k6bcNPvfoCLEUd98nGPqhgzRVn1eutDWKLLarNEKhjpYKIYM7Qw/u
6PIMfqK3dLDkx6E9kaQ6U7W3l/4nd/s7QgMOPO8+XDOYA7s+mNTHqRrVUrbwzaTeVth8JDPcD0qU
JDQ1ukzZcRZx5WMMjOeHlqFdjgwBSDJYxHgzJlQxyoEsQKjetvrMKsreqzb4jlM88eEuvVC9dVJ6
MigzEyukwRKBVVJOjVhfwqoKsO34y00DSWbF1OgVUbcqJYgdYi5aqGUMVR6STuxV/b5yrR9VIRgS
oJ+rb8VrIx2Z0KKnvT3ZRGmHWyTX04gKpQgAZwpcS/HPQVOdbfhmS/yUbj0SDFOoiY7RAU55qJdp
IyucCNl/fcEQB0QhSxfrG092hPBSiOgPTybty8e73FPfy1Tdbw4LackKMQ6ZzEw7ApVq1O6ATb2d
KKJlMJgOIkD2yg/qiTmsEQTzwYGAWOTpm0UM8a+8QaPyHsdn5yRO7JR+3yiwaj7E7n1odExWvs72
sp1dHid8s0QW5Mo6karJwCjFB45iy5uUKnWZcVL26DfpukGCNz6TTFljl8vtjH24dJ/TTa1Cql+Y
2g+VIH9MGDQsmBCcjjsoLoRFZ+6nlIK9lTGWGJgOSaWZShO3vl2mW+e2+mrf/rWLfxDWBZGVRVY+
m5X1k6E/Ak2uXJaGH63xESUU234LTTFHiwqeRugKzdVCJIXQ/EiTU3/jnfgZKiOt58vW50CPK715
KJETANYr4DlfYXJJ4d0dr29AlO8uEu75QR0O1hP2LiuFCLX5LuxXoSIxGv+kwfCtVIya4Hb3qRtC
4W25Nm0RkzWcEnyJmJ0sHSW21Uz+gJGREoBz4Y+lAkNQRVxL2knlbnTnlDMPe7/YytFwZi6kDR5a
hypU8GjIZaWBQZPp8VTp+beKUAmFFvrAtQxZg1a1XrCRKu1bZujCfLJzJTcIbCWhqDhtxX7akzKw
Esp8P/oXyv779sre4ShjGrQeVfLdNCo5+ttN4xvythH5bVHXYuD3m6AR/I8d0FUiYBOzpUnlpheb
PZpYh4tKWeKNF4XUWVoWiB8KAPM5d5/q4KVQpvIFDxHNlzkhDc6EKkyOAjUBpSKxfa8MHATYN6db
r8ZHF687MuaBBLOvt/MjMxAQ+5k6qm9sjecrS7ZN+sEert+brcQ4Quwi4aIzjIwzE1PeLBK6cdtH
ro+hiBX5dm0ZdGFEOzvQiF1Lz4nw+pXVTcb1RTTLYJQ2C9gFJ0vTTXYnhKNcu/3C7Q+jRUSEQtET
ry0PdlvopW/z/sF003S6o1jj5ZUayhq3+j40A5dVbSjsUnfLU/8MD0M3dTpG6a7P2t1g6GSAGV1P
7BY1LnbzYqzxmYzOZ0zKTUDH9ZMk4sHdsryEzJ15aZHRlbZQ/OH/ZVpT7D3cIqLgWKqT6+5SbgZN
oO9ZuvI2qQ5h9+4dBmP1rF//pTSfBJsC5R+3RAobnu2k4LSSyeepn5ctqVTN/qXjFY9vO+Q/rIIc
kuOpRBq7tSJcRS8n6Tyz+vYOg3dLuilC++VtWnVjqLRG3tB8/XPoa5M1YfDTUuV6Fp12g9yyFvy+
s5X070tqeQsEyy/Fd+xrNoW+V/D6r8+3rfFwcpNOalN/roG0UHkSSDQIIvKIXn8BKsBYZZF1e7D0
VwnOQam2+9AvUouDeV452O9IbHOKo+YdEp/Fv+5KHLl1r4sWAj1zTurnC4WVq1VNzFoqGnomgTNV
8M8Sq+G9Ew4EnaYCXyo+CNk0+WQSX2QMYnI9GMQxbdzTMCfUF4Hl4GLQ+HhXslOFs030JsRpEZZU
jk+zFIMtvR7ndLM+4G0mk5y0Xd6GCLYLiy1BEuQltpeEnEnoFBbhxSpTwfq0TxA0wAIK3SsUMA7n
4PEtzFX9tDSeR/1JebfpNiufOI9hwM0cthmdhSO/Q5c5lb67VQMfsmowKtN+P1cq1D9WuTuoN9EU
z15AFDrVU41e8+NGgzo6fmok6AbU/9XcEgar6gLzu7OwO1b6Rg/WjLAYaowYlBgQ/2lr8eu3EwtT
EimkKESMge6mrkNDoLhA9TsdOv6ehERALydSjmmpgiQ2eUZqqSVdl8rcyCuFHmSGTNQEKWp6lwpw
5wgpz0pPv8JDurOwWwFaZonHU7R9xj+q8ZDqWy3CfN3EyY0wu617svYDuA/z46URrkXOC2Q/Qkma
ygztioL2GjVAvH1QsVjAJixkP+jcL54Y47cz6XVCiP4jUkBwxU5p0TJ7E3bq55Evz3Z4CUvyXS4P
Xy28UvqAbZ5yrMiiN/5OsHrQZMVUJaXj9Tzt1RiEJq3kgsxCWom3Zhz3ochTWCR827JQLRZmMBu0
GeZ5TnZNIHrQb2peYq5U5cmOfppd/jK7mUO6hBISi65RSYAT4LG18Df88TMeNysL38SjjogDs3tb
uKsGIDfp3r2y3IWHaIoTQcQ0RW8TAkW4bVknD0kYLsoSMOSA7pvSTqeZJx/10gOE0yrYfdVJ+O07
2TXTowMhW9lIfj8dHOobtnl5yPeqDFSGWDDbRX8wRhJdyd2SO5CvO/ck0giUrLL7WmZ5oIFDR2wy
s+L1UxXAw5+B1OStPSdMJc9PViSpmyVo0q2TZ38xjwIjDWxqthaR2NW0xSOSDi6fuY6K6qgx5uZt
aCjc7OdjgW4VzU9WglZYYRWRu4WBSy7MjBR2Ye10BgJOisrB5KXSKl5q+yrmQ/5vwl0CwyLkgBkq
k7k39qcBroSa5b3w/NSQc/+CCvrr4KjNfNULTGOnT3KcGzKpTriUwmVX3K6pKTO2OAUlQ8UOx91Z
cH7G+s5m/gMRMxq5GC0aAxbyi2CkEGI8/uqQJe2zrAom15J7DNNyecJbTLEe1c/AiPDrRn7mX5Gn
jO31AW2FoTnPEXG3zglJWylxDUzoQ7Yvb75tEgFACEoGpKZx+aILjU0NJvvwOrom0ylZ14UcsO+b
MZAYQ1XD94/OxqXnoNaXVpG4Xo4BfpqNVHAFqmOxsaRKaQ6CbfBOumZ8vV13fc8G4EvTmpPn9x2b
1ZpXRHdEf1mE4bp4gnQy1xT+oybWjHPLbKbnk57HSnoQ4UClRUHG7lq3xHiMLPVfSh1EzXxthMb9
AEBv6HBoQVcjxVQdQwawiURakNZ4xt5ZmF37T9ToVPkBA60BGYxtN7ip3KsWbElT8EV/fbUI2+As
7j61A+7Cgm550bX7UtFaXQV66hgqe2Cppkyx2UFdD1vpBAum4AEcnHTUYoNkrHBDIfwro0HPtDL8
v0IT/sPOvdhsACVlgZjwCCF9VuLMKKAUPXYL8M/sf1DSZ2pIPTFUfNgE21mngFYIychz0gbybKdx
aKjH2o20LAEammD5PHYeY8jnQVNNG/i6Vw287GzI4SSwjFI+vDYiuQ1ihGZOoLmfA/I4ysKXD+Hv
C/DqxtmB153tGvJV6F1HvwKHCm8S9posWqaHmiblWcv9hNJ+JtjBtqidxdGVsb/BZN5aK7THj+k9
txKLFMOqfm37mbwColbnl7+mnK2mlVVdJ67DC93l8rrH4qKmbRMK8X4bHLT+rmPe43GizUUqR1Zw
y/pMSp8G4vpSeXP6Gh312HasTkItn1/kepcfCSeFpT8GJD/rYn9uZOE7Y46pro3qS3tw0nXQuMZs
RiHVgmwDv2MzXo0p3JSJ7mAEmPz8X7cjzZ1rsO+2eirVA4GHd4bRFXYqonIQkM9/h9a/Po0rCOj4
TdYqUHnu/XwsKx5dGVIMY+OI/vPPoXtQi087FpZTDZ0SRIw+I96KkOF5kzZBrXe1leNfAvoTA+hY
llKaD/NFepLMiU5Kd5MNZrRC3Uc1ZGCvESPA7/tDOnfgQnpnLYWOwnfkKYQu62HPbuhVMTTC8HM0
MacqfT85egQQ/1e1e/gAXnYCwG1cllt932O/0p6GpSo+yNqWH+vnOTsACrSoBouf23zFeY0CuN18
PA13JdxDjtOlOnQOHfTMKbnP3L5uqOanfvIo4EPFrv916NpW44RuxL2gUODqYMTsl4nuRMDRCgC/
W4Q+WjUUK218wjy/JDxK0BcpYTIiJ06/14UH7EuVo4V/mNYuWgxslFQ3QPj4rfCT65jXRN8E6gvL
3XFibuvw8dvYYOVJ91w7zKXiRWL9FcIJrhwW3onczbWZkqIn42tFj6+SkFebLRbUFBEOFmV5V59d
0hLeN9z5DzYwRr7l7d5nXYN9jFDL0FD9oh0qVsndkzLYKGFyEVb9c7YlIuQbRzC6TcYj+TwDZo48
Fw3wrJX3onSFLODlIakNejvveMMj659bwruZIdqq0shsmwxwe25/C5bh5mCLY1SPgPC1XOFZ+M61
63bNv4X8cyYTJu/OFG8QTDWeLEb/ntkm4jvWsEfK+ke/+gUhJgWbznXHXLBS3eEFV6uNtzgtavf9
za5lKbQKIAqllbW7zTVAENZYGmxQNE/5pargODGysxfoXIyi59ODaLAX/SruimU7K4km2XtW7Ydc
VBARfbF4auUwGhUa9eJ8ND3Vbi34KUGeNkc2woAio4Jr51HeShUE1dRkhHGJU4tstu4nveSuxKvI
ECo1eHn1q0EkuNFmWc5W6jtvdlO4icLC9Z01a8MG6w8Qhnfd/bkWLbIG/aCKbzAauxJ8/CL18otd
HdhrlwZayjZQPhASNqYp7L7qj+lnKVZXJp79nOaikpAq/JPmSd+8YSYklEvjBpFapQ4WOV3wRlzB
X29J6PiglhpPHTKofYiTaswsPDohjWIadA0yDuEr6h2DaDne9lKBQMS4wtXC+1q863nTMiNENIUS
UqHW+vay6XbncBCFqKiI6YPCVYggPee+IGFiVwFEtn5EopJJycD82QW/JxRgqu8PYNFnHX2003kh
RF2gixQSVgzhIx0jocrX6/tmEMx+GTlMCyh2sxBJQ/fVxwSUqP/VbJCpZuKp/xly6kYDJrZbeSo3
fSAc7+TsGJzD63NKJUHSAUQNGtHfw4Q4Bxm9C7/8Vd4BkApU5BAunTtMMEk+fDoNdHfB7DysgJrc
upwEHGwxOKDzQRSSO+yHvmsoN5k6yp+ad2ZcW9iXc6KNU7NF0hYWgo6wwZrbTelXIGk3H4CH61p0
LI2jZSo91hMwzub6jqoBO2mfmkA5CitgfTdfpCLcl8KKYNHbdNjeIWkkb86DLgid8eWO7LjvNVCj
+FbWxNywXSxjLKqo42am70qajTVf4IHdLLml2Ro+y49ocmRmxnfwdhQXUqPZOFIqscMXls4tkDPb
528GvZSAN0l/7FcaEJ7PBqRdGIaf+Ie+OpngFhqFaZzJhDiNmr3zdN4RokZjza2M9QmjBhoOVXnY
93ws+UoA1weAO58VDYhCN8msvYUbhGf2MJwfXg7lBaOSmsJkbHZb/f8/TydWL8Zo7P3liLC4lFc0
FQ3GOojDgLkCwEp2+7bWyFdSR3nm4S80raY9T+3GaUy5olJ2AD2rjlqNfO9DwA13yZ/szVRuCdjo
aKhfFhw8EueZ89W+ZayY+5SZOwqLxdYy0fsvmRsKB58PXjmUsym0OvTX7nhljEjH9qOsPradKKAm
SSI3YjkQsKves5A1WWz/4joz5kkulWoUXrZZUzMgAWTgMaayr0OuGZG7opIcGfp1XIH05yyCN5Jo
i22hqAnkq/ZHPIjLFL3FGl91SsU+M0r4enlYmDRnndwr+c5K7rHJuGIBSAkPpL1MmpWEIJYrHgiD
bfWA05DAkacTFUugDVwWYbb05GrX3SI2lmWatO4ERLk0l6n3dgbR6+/BPB0+lVp2DxsJYOSBDCvQ
api/XdinLTlHLHSXq8JMQGAOqcEDnzYJSPsTYKddFd+fGriPhDLR1voEay+cJ7EEwcfcSCfplPuE
pO5FyVznimfRKLlQWr0jqVa6UHYUvb33pBM4gSsiUB5+xkk7/xkD1uW9JlXiQo4Uc+yAW5jdzjMV
xoJprDZJseL/joSah3Db/e81vXRIVhasEzVtsdseaweiRJ0+Lwpx+TFvWqvTSKBKfparrQEwG1jF
2WD/RAv15rI1taiiqkreNDltisA+MV7sX/BCCO/ipIUnm6F/FhXgP5QG3xHlk4AdWmZqoif/q1qT
+xJ1Uwas4SWGBeGdcdqMLypjDKLwYi36FO4Lq4A485ssx6xom3u399+Hl3ed+3iMRHUIjimR0DxK
4xrvDkSnKQScy+NKGBQ8+b5Sp7FH1fA4/GJubZuWDEdx+bAadUIixGp3tmTn+LlaZbVnky8dPTpB
6d2A7VvPRgdPD9lW1hzqPpX/D2g4sCUQODEmsWu1AaSP8brUOUSkBlR3/MKZQwOJNW6TDVbo6BMk
EY9zJLJXbSnTyDnpWixQNhXqeiLUn4aJtgC6TKc0LgOAQlQNzFHxTzM7XLZh9GJJKd6wHIuKUUbU
NnM+SEgeRc18HzZzStAf+aYi0l1JwcD1bknNZVuwwlL/wetB/2sSc+Ab1NBBwKcTajkEi80ZS72Z
Gx346f8gB7NiH8zaoocDb2pIFj3l5UPyK0Wk1frD2KlwQWzu3Ua12lYbHI9YdRqc3BKZyjVhwAR1
M3/zlTB65Zw0P0mpISWNzD2E/iu3jJkuBjxnQMZRxHsE7vYVff+D244Ln/lBc6HAbbzo+v85IZLw
TIzp5KTXTHzgqaK+VBhLrPxtCl6Asl1j455RscSTmSToM2i29J/RzetPtVG0k0Ac/cBpHKztdGW+
1Aapfhn7DVoGJZqd8xeiutI0sVP2yLHMT8+GFT3VSbgnRSCVExO80gOrCwVwEidKE++SowyK9pd0
zXiRNWG6FMlPql5H6z3ESKK4WZ7bV/t3YtvW3+TpxOl95t2HE6rIqvLRr/PNa7wjP2wOgS1Rd4Tu
oDrGm6L7qJNQMypYeh5hsHvwPhlEE8FuZvr1NvM0hZ7Icx29/2wOdFlU7sfGE8r7D+74Wvb+CxLW
oM6mLtSSmVDlEb0T0F4A8X8/QnSH0ujt/Zt7xltqfCZ4hHW9dzKXKaXhzcXAvud7XTs6hDf/xkMG
dIPwGZylgGnQ5+8M+AwEGtz8OrV9flRR+0v/tEwzvRtXYRSOO17PV4lNNvntKdK5FGwqn3CQPyMa
PCuU0kgSBaxWrql+kUpnWb90ju9vhKJlw8wDDROxfjJc1EIvC299A9DY7LQ0gcduxjFzOTs8cOL9
gYM0xqxHQ2PzyaakC+EmzR7qOvV9+D7FumR1dMNLaX8prR5gGzUh8SHKFD1txJalEYjIgskKNWP5
hN7zmptGqqITWo8DuQa4+OL1PC6jPfgj3ZuMjG1btoIzSTtTUGVfYIsNewleYLmMlsyzFgwHWf8k
ykLuHm4eQRfPHgcbOHLwlYi2Q+JuIL6r1mb0n/Ww/DtILM7W3kwTkxTMBt2yIpLZ9qkflq+yS5tv
RNLQ3sR/gmKT9BlGhZlSrzXxWIArHhVkzQspuXnKOVFQckgC2vTgnkV8eGHbM4x2AXvo8oxBmyQl
u60GnSkiLu4FgUot2UKgpKDUvv1V7ctK2cdnfJmNCckZ2GrLqjzSoMs9VaNWlAzUOtr0mi/kE2No
/pOcnzbcO+jEshFwFqYr8XTfXAp3A7Jf+JtsRMqbPUgNHiPgeGJtO2Zb2SQwMiuhFXbJkcYU+xjH
d4odgri49b/ej1NPbdm1SinipPbrUD7Ln7R/JZVYCL19AZtjPr/AWpR5LDOa8hD3w17r/KmmlTdy
sRpES1B76hTlq8EPNeP19SVJiE060Da1hfjIEMCLfyskTjX9wFvtCBRO0N+8m99QpTQ+SVzNLGLf
iGz5D8gLN9gH1VRGkuAoNFfI8f0uh/FpnqjXmR8iuWXjPQzjkBM9t1/hpBnIM0ihzdbzSgmH28wh
cC4tGS1eaPMaDPA+frMmYMKxgg49ynKnEfomaMETKfJ8cB2mTrrXahesEQ/yVMqStC3nckQruoNd
KJT2qyiD8rSjCKQ/GN+vnzb1NrFxoV9WmUQHumkJAMh9U3ALl3XFs5Tq672190MWNhbBDyDN511y
ENSPFCVT8WfOJLOmydY2u5VtNrr7X+xGDxvHAfbDZRU424kAl6tu4H3ArA+Pl/s0r8KDF6qmfzy4
qTq6mC/j/PXGdOBAq2+H+3EuN8mesaG18bW/mAhvYNjd7IT6hlpAER4CAJ6+8fkzUlUuoi9elMuw
h5QQhCUYdRMEdEwRULwMqy+S2e8iYKPwmX/8ahw8iUxMbom63MsPu3t6pUe1Ebd+8xIgFU4T/M4c
gNV6cCzvaybQKLflUWJEUok+GSENjPcll12/o9L0kVtpB1WUP5uQEpi5/UAy8ixgbMPxN29xg4mP
LCNjil4ff3oHjEaSdZEoHjZh+gxpIcjefIV6NQIcnD+q7kxoJo9GQsSA9TqWhyy0s+ic8iSBlG8A
w7OtyRvlpfcXgaBXAOl38qum9DRTxR2WiUIpTUBBROjO90FXumBok5TLXzI901X8gFGmE2BzoUtn
R68q3XsL/XGljKJ8iuDrxNnwhY3j4bze5U+AQLUSU/K789rzpmuGCUtRFxtgQP52hrqveFV7ifTa
PaYk+a0w960yN5jfoowPsAaYx8aTfN16VbRxg2pJVi6+PdiGhfl5hVt9S6i3P3ppfXbdsQhgN5rp
vChKuZ2e9d1upYQKSNzOpk2VcmoGQJcLOQdbVu110fGtnSAyqisFvCuvPHaA32nUU6H7iQMBCOiD
T8Sj39ceC6FsTBe9749wB3kiRoHxvgYFyHbsDlLR/iW4hvbyYtKFeoargwFKDK4+8D+9BMzjlujy
GjzUgHP2x/mgP09kdRzRCLe2Jl3QrEhpSQcONxwdqea6M5g2nfxO6I/vYyjcoLLxSTysw4DpS0nC
4YkTfElulLnTnIbUEYQ6Gg7QKopE/OQFRby+12RsfNwuwgCq0639JK/O7ndLkZUb1ECVNQLf4uQ7
8FkMNeq4d4KuzOwePY58nhRcXkPGDNCCuglVWUOuLdQZfTa1ZvfeSP37XwylkuToNm4zvhN/VPSn
U9AgBtgklp6p5xZ+PaHvO9Rgx9n7txnAYdJpJryypq+YydE3BX1NZLms66HilodLSuhXeiQ31GV1
xowgv3BTUTwxUEUSOmv9Q78rsFxLn8qGTtBI9RyF0YMt9kyzFtwL2ljKGI/+JF/MKcbqkNqrlhNc
O+NWe12VzocmJoa29kC10rZ37y0Jn4+VBZPGYfvh5XAXtPuTdjkioW/qI7YNw9+3UbfLEpFptJsM
PK3eBAzEMmob1ZtOsusMrqGjtJSMBBcxTd5btXNHV7TI00YqQwtj0EdSRnxxYcro36JXw/ZdFeWp
wNV8qMSMRSFR6Ize1PRRcKzgixxZ20A7F3kF7Fst613WwgwwJiBwIjtk7OJ+cvecFxVlQ+CuPLWt
wB08Alyrm9vYQBvf+naQ6JgFUUP4fB8EqAtlPVL/e4cXbZhy1o3Dc0Z5dyjnB8wSPPirDpXZWR4N
PLD/wMMDXXwVh2Tvcc9YwBN2JYPJclgFp2yYKuYiY2GO8gPcuNzQDhn/rvs3C6gmYYlC7guQq0j2
FrzoAqoG9qbmJTSfIdY1TCITVf11vP7DISAirwhMPpwEjKJukbtB+FznyHV1eBMkNN2VAG/mVJsO
Ou263Qvj5qqCS5j8Y/dfgSM7piRtGKye8tVlBqxhOpsbYBvswj+cSCFxY6b7SurBYDp/DrLV1+IO
rBuYIQzMfT3shA1gVENgPu0952gusDJ/wM5YjxqPpNhm+fbIf6J++UFqaqqDaIvvtllfHOFCGDUG
Hdjthw+jCIninKYavIf40Vp3fbigl1yR/t2OIvEUFsuhCxsVOjRMG9F/dzFLjGD4x3iQ4X4H0fw+
ZEmGIKZYXOP1jJS9R9Dy1D85toaP3p8TA1VaUGPloO5UIOM5Khu+iUDxUKiGskxOyVVY9Ae1rkjs
sRKtC8kL+3FhmwB8ObOhn9LxhPWVMfbWS+2vvIqS3KzjkwXXOl4ua6H7YSLSiJMH0QKXLZr072HJ
61QLLIKoRM4T9uBRekli4Ff9H94QZg52/aa316SC4O2NJHta28eDz7zGcmmLmxXqMwEFH3HAXU7S
UvcLUKNj2HagfJwWwRsQmTkowwrDnZIhwG47cazlgey3iMVYb9hXqLjb8m1g3GvRx7pG2bJdIdTY
B77Ccn2AK8N0OF0NutYo8cLmoeap/MJxwdBpJO19RY39ekUJxGZfjtkNOK4uwFGpIO6d3C3nOQmM
EOFYsTC4NUnTpQ51AWsFNfv5msoHZF5E/k+jFUo4rRK5KRxWJf2e7F5kABrkhBwa/Ao4jkkIoq5V
WFM3W4pYoAV3unV3phF83pslHX3YZR7QvP6cJkpvn+HKSo5PKzhnwkitCKuPNw4CSWMVSWU0qWZ8
/FIusr2L96lhMj50mFZCw7wUJEyqC8aDNU/WKboA1KOvxzANQF2WyTPP5NXbkVFMkP50lnpIBFbF
xy4TVF/C+GDOz/Cr9XkMfjCsPnzEeYRXejemTebwaVjnWhBLlU+HFjjayRYV2NfO9xeVH85GWjIu
ZWpfDXdcmWIA9ShVKEpC5yx66g7373H5b5ea9Okr9TId44bevlvYptVkWQKs0zrcBTVBKeDqlHZg
lWEKHqj81KAF3Qfm1CrjJ+kr/KKWAp4xhjsHV5xFzJxHNKsm66enLKOBeOlK7Hol8RmLG8kx+DHf
+0IEyJwohyNG3lfFN/GoHyqKca4Q20kh9vMG4fDmtnQmsSoKXTJ37m0/lL3WsfgTuDYUmyYugIEN
8cmmYcytDZGFw1PiA+h2WojleH2Z43rtgbN25borSjQnMu0ybFrEf3L8u/X9D3zjabFAoRtq4zTl
w8sp80VFc7V4NjnXtbPrSuZRhNAMpoI+L/Iio21HVREEuyu6oPYwtecqPsjkspzPnn6jbCdSOEnV
/tCzHBSVOkOBGxZJB1/bZ4zOIn3z/txv0rkgJCfP7NIXx5IzaFFR1IcHGZdM6pl62T2SsG3xMnNj
FXsE5YTjYaN/MaHLOakPamdatQcRKDCVxEVN7tVvggPXKWQEWjC396N/2/znJ4KjxsyNppjjU7UP
znAxAp1tAsJdjwuyzAZRQGMwguc/b09PmBoLWzKNUvGpExkREOHs02j6nsUpQndvGJ8IV03r+/l0
FiW5YL3eY3c57esBH30u4ngCl4Mvi+mQ+f8u9dsXQqzog/5ne7sl774BlxH00Nqo5L+QZL42At93
PXs9ifHmCJzD0vYN2X5UuzrqIYHTjtrkiVFxlhZoggSeM1DXgNhxrrzTkcqtSOSPGg1PncnI/nvq
p7ycVxrKif4Q1Q7rKox+liwwVQ/KByEQHBAuAqkFQ334XEVqCe2MTmXzTejxgCAy0cjkWatabduo
gcdOzjUKad5PYi9ySvTPOBGbKMh26VHQIwrkottngeKIeBqeRt8Dzm7sN227HFmCivRMiqAMVslI
XSbY0MU0m+T1xvh8pZhN72UaSzEh48celjenIE21D/h5Yysp3Yy3tVVyiomSXxqWWi861aOLfdDQ
fKlXIOZzxIy1iOdgfVU9nABK5QTTGYNigVqqx0/HjF4pNIbV/5dzwxgU9sj7lXVI6IZ1qQ0qp8hF
EuIn1XUfpJF8ZdJYayq/Pp6mtWPvEZtfd+vSf2WxEi6lHtRnemZ7rvJ4RgZniIVhRgZUrjXZKiDb
zvlfx1q8wI9qMzvbFrjcZE8R8AliHPZxJJbSw6f6ykRUg7a5XV6liAlp4AkGUYvz6bv8lRb7CBQ3
3GZDStGLuiO/Ln+VnepndFR5vxdhxNxaCqM3iixq7afhPuPo4lJk7sB4yJtFO4YRQ3FTaJjAC69o
CVf65OdA+gyC3cvKr2d7zXhgqQrnpMNZZU8w4OJf+yTnOV319i9Y5BjVuXHR8O9RVTinr8pvABjY
/LOTyDR4Mp7+xxVe+gYr6ldl6Derf+OCy1CbXX62heaD97AV8Gz9srQ5rtSkoOy078yn0pmj47ja
/91rrixCzRG9m+asoNJXFcfkKwNg4i8Ej0Yx9Q8SD6jLEgcvEA01sk/37CORxKDd9S0O6uXwnhMn
7vGK8r9oekKzCoT+YDSDxMMeUiVHK0rqY23BsrAmrWfEKsDizYv4ud8g7tcm15jsos+W5JYPKz41
+6j+fmCpj4pCYMmnVdTnnR0GeH1aVR23PCCVSUdAIkLbW/Jhf5E8aOWmzWTJphvWXrkHiqc3PCmT
tCb2lgBYdaYsvjWS7Jo8XE6DXQhpm+BenFE74UtpEINFidpw8kwlf2jNF+Gm8pVjI81QmqWIgXzU
T+qaQS+hRe7MD8JYRpQmqhH0D0xirGpaK5XqLVn0GGJg3ljDJo1hFJjKv8F1uNN8Z8+2VVwzd2bo
ivOiNMkLblrHmK3Mlg/6shOokzRW6hMWjGEC7UvdkDdu1sI80tTiuBJHwD3UcSOHb7fComX/TG3L
4qKR4rdbHd3eHD6W0Tui1fTCulVmhc48YjR5XuJ/hGXbz5P4CMRbu3OXURe9yS8nF4RZ4nJBRqdq
BTMn0UvdVFQGqtuqjZPW6NqrlukXev8L2/CL59MsAm2f3awWswa/6Oh6z+Tsx2kJsTCTJq0k8vMw
0HR/aGpaq2f/JAiD74UvCEigIaE4qUuYZKvvsdLJ10MDM4G5uqBJqbfsfwc7Z3sd7pIgvybvKENJ
zlXr+dLPwaE4WJGXugcfhb03iQHxq6ztPI3xxIhp2daI9oUUDTBxj9PzOu1e9j/57Jf42Z5mbMmm
1qsqW8YlFsuO6JD7UDzVClYt3fJEA42I7cqP8+rQQmjX2tJvpB7fqQd8wTmEMrV1d2CSBNkthcjW
j4P4s566RUCq8sxDYw6SCxzwcDmGitc6faPAjmGLEJROiTx4q9EjxgKRB8v2FUN4xWFbZiadMJRJ
nVOTVFXHesIDma9EnfwlGo3jl2GCV1MnS9Tv2Fnis09mvlFgDbS1YvfzXY/4ry4+uGXwG/lpfbnH
ugIydGgwMFFn+Y5oq4c89P2LpwIe0l4GofaDaLgQw3xAhTdsnLYGvvKSaZPjnlgiIiqwafi7eZtQ
b5Y85zBZ+SfbhmJfxTTDIr2HZon9gLaRXUY6ECzyFxJwkiuA7iL5/Q6h6QKRaPLmJ227adhxgknW
NpjVy8/hhr+5l2j/yvbtUWO/F8WA4mYhWcH9KpzRO2QmTPefVSPo4McA1In+QDNykkCuuaAc8Ob2
mjmCnU6glcIQzBf9poljidsgkaxdiThiFcMj/W546jwkDHpO8QRAE0fxIbAMVLwpC83zKGtahMAn
QWckRDUxN2DDbhqVppL6yrElNNHf58sK3+VXfz1I3f2kxUqaEr/pGXORM8wTGwTyGXWHBqpq17VD
nyyPFBl1k1Bz7p0Hjp6MHAI1lrhfPuGXC6EeTrPTi3QWZXWbUncYLJr9fcS+YIjJ2VTZNylQV+iC
Dmhae3P1Jp8K/zSDZQ64iAuRT/XqJ+4IQJA4g4p3duMJXHYH0DLMJo+Pr+chWG6ge58fF1ob8LJ/
hvkUVSatyelDx/VCnOfCNYjmQ58syk2iq5KbLAiTV9Hx7i/ze0dD9Z7COcGNJrJ71VmLBqQNTKmd
48qG5H5JAjiRyIqSk+w9zVB5LeE0ZMV/kPHxMFLeYN9TFfvJYapnnGHpl75pEpup7gNTL17ljtbP
rLTyIV6l1xjYwiPKWWtfpA0lA9vU+AXdL+rFMx1Eg159yNZYo0DvKMbdwGI2b2/CH2weUX41BMHd
uxe43w7cI/qbusxOUGQz5xteFWTHzP7qKdn7ZnmpH+cnbmGL5xy/zeKYSCcFPjbBLqx6A1Ii5s70
0aIE6iubwproomBTTwbaMl21v9ZyhxGMYqxS/R78ljD54tYGxMIlF27DuEFTd1GXx5UT55mFRLlt
vj2sxnrW/YsAqiSzw0ZTrQqOLWKtORK+JMrso7OTm0V5ZRm8gmd8kcUXdt2J2/VqBrz4keEwlXJX
KF8/ppoh1Bs9vuc0KMCaIA31wCuwZZOpuikNM7GtCnKoOtlApzeQXiqSgxKaJcwfYlKrqCB+dGh7
vVaJ8AY8pr2RsuXXOYGavp5MKcqZwJNnvnOwVKONeL8j/wTtYKiqZkeM6PIJF90vNmseyHSlURUm
HIuQYN6nr5imxrbOw5HCk4rPLsatd/IK3FcjT2qECGdtf9QFk3NOUVvzsrRIAkIEWeRjjlvcEo8r
fQ3Uft6R1wgV5gVw0UlMoD+EGmTDJw/V3P+XZKo7HY0YGWUXgERqtZUh5F0sj6sTINGOFP8Ktd98
tqUiASPZ9dEKb6H6WhPqVH334X4BRDRW2qmilst+f/5zpPv31Eq/cGXyOGcc2qzKjgldbfLN7aXm
OwQJqn+e1JVV5I5BMCU64hnXImnRZSQkvryEZn8QuPVvMzQa6Fe6CzNt5UsVyH2eWTo25z87MH0y
ZYIhrpf0MODz6UCycvDQwkDoXALhicK/NznQhcbtrmOOQ6gAQfNFysktYZNk6M/RmadtO+2Gh/P+
fwXIp6FWW4segLrRIFhJ85XJGLTPi5w9mFnmEWX2wxBJeLQcMV0DPEQL4K9goyPGNlo0uGYn0Igr
mlG/14b4GnEw9jsXSjqpj8SKw7NgSyvJD3NLC+vVqlZGTl/xIAkeCvnYCuP0kKIVF5XnUYHgK1O2
bbEaWJlhZmZvPFz/rMhJ7NBBOQGGo2Pkc30RzGrZb+BTtCvpVEjkwb/nYed0S93b9abrn0xjMXB5
1uGI2MJqg00DBxkupns0lqSjTJiH8EA10r/bHoKexGEbCfEVjCSE+RTKFM+8a+xuFr865B4R4Fu8
yzIk/4xJ5svsEjY8kS3YDH2NSDRZQVAJ/J0/9orH/yvmCQfVBPgNHNqaH0UFPRwPjTIn/Ucsj9Og
tW5ZNaV4vU101uuHpgd1Y5rXPQO78g8ZFzCYg1RYqDGnBag8Oqdn5dA8Vn1e59nlKE2NU7OSZ0Hv
bx4LdBMvYLGt/7J9kjIsk/SuR9W4CpyKki1SbhrQIN9GnkX3DwuUG6v3EieN0Uw4W9+O2LpmKBXO
t9ob5FZvFjqcQlwCLJYcdcsyspv7d8PcyDXcHYaK1hRuWy+vJ2EsY3R4P/NbpF9OWhPEZbJh+fTv
EuzvaOrxhU4yEhuxX2GFpgVKfBepJrEzlJnUhxRRC/YhRe6MUUFo85YlsyIQGa0A+Y5qFHjxAGA/
/kt18j+aileyqKw98/5a/0rfq7QujrNnrdqq6vWF/XRPmZXDBGzfyhue60o5tE8E8rUwytbZbYGU
7+gV9WTyQN0fS7qp7eleZrf88ZHGo9hkur9cI6FPXwLGa/Kf7Zg41wKjdCgy2Z2AiaLjBmZR59u0
YpsqUdXhnGkxpAuo0KZ06KBh5GKD+jLtcqaGKDtASjKBK/ZMwOvW6WwrayV8747Yxkw/ciP2QJxG
Pjhx79qlsad9BXfUtMxgi30P6/Op47KAW0AOdEck3kW0APAMeICUUYvpztVTPCCfZWzrgpQCTuo0
lx66YO8OotGvIbcJJmY8BPOuLPNp5pGAGtYJurWgcn8rZFsVzXQ1wsmAxTA5nexetTGH21NTt8jr
ApS7Zx2yHe0qRAdh8g7I3Gnma/2M4FG0ft3J6aZIDFDvKHXCBVV8LXzPYwjLj4mBvDfnUxNH3YlM
YyFp+4l8QYpmzYFO2s1DQKCWIzz9SAb0LzwQQQywobpMI/+m1C3iv8tuW++bN9ISI0fxCo3s8EFa
uaQcOyC1Tz/Ylexxmk5rElUtpwYQnKf3qEbzC5vrvwg/GzmMhonMyGY9jktof+zKBoEixw7P/dce
vG6LHlpQJzEBRzEJVp8VwiiJvEigstJWjVjbkYE3UcYbjAgc0rjiam7N76YE7gnXHfOjfi5+vjov
n28qykss1Y/RQVLDZU9LcLoIHgEMLTznKQbkzzKpEUbk8gqfCXbSzqUt7rebm0/8gHd8HlU3Edy5
XfBcTOasfQWbBnmiY4cfvrvSaghpf2/EmEkkqwIKeusFiPaQYH7H/cFG/Wbbi000MMTL7SWP/NtY
eAjBw7oRk+jBnOA1raEKLkU8NUwpXudi/qcVfoMKDzfJb5Dnw4LqXQdtYD/ETWHaiZD1Bx5+EOn/
/7pBi6JXHtxQX55SRMAifGfLh7nA0h14kEBrJDL1IWUIlU8+sJE+G4c/OcioXGHSCosbjT2c6gYd
MUb/1KjW/40pxlcDoI/hbO84Bh1FvJo3Y1JMy8fn9mgU5DI4OjplDkR4j0cUihZhp1UfrJWZZXpu
CO4LGiaFRnDrCwCNAiXXyM4uw74SV7kTHE3FZHQ36+woHKSrc07ZLQPvOda2LH+FKwXjxP/vKZYk
w+OF2eWADwjdlfXaRGpypDT+/0H0+dWjRVsgmu6txkWG1CRQhVpsyCSq6kk6PX+GZ+QqxYkKTXg8
9Wbnm0tMwwPC+gvy/OmlkJ7cRF49sifm1zR1hUXCWQfuLQplMCslTFEBSR5gITfN4UNJqyXfjyZM
56Snxy3jtRKVtbHs00RdRO49iyRsfzPyKkspFVCXnbPijyZrExvJ3+tJuoWsrYZBdCMQ2xhSaXxT
S+DD6Fq98psWago5amokQZSD4b90aDiU/OdQcjGWmZONc0oBn95QavLnwXsK7I8FWFolRe/ygv5S
G7XSScLiWr5H9aT3TSLgthvPCkQnAhlkcgINSMlpvR4VHq74OMrg8HWnxYKbNJwdSu986pWbUiJY
bSvDeJhcSUsbErOHN0O+O4SI3Gu+LyQ/zvA7T1GFZ1Ey3Cv1A0MDNlweT5DP+H8tlNbboryLOEqf
1a2oZeIyp7mIMWCJEp1y0RM1JQMNjJthKAk4ZhW2UcW0CQRNAumvULYciR3ssbnPIhdfSCLJBQU7
0hlu6f7u+50EjJ7bRnxo6PkYVEej70lSNPf+FhvSEX/NVvX9hJsyC6nN/I20hkhOtiFuTpO3xM+g
pMxXgiS73w1zLUTfnXuzTE0WBxqTrqXh6bh7uv+6iK2FfcXw8kpWAwFrBVyFrse70kHMsg7K+fAS
/THUteHF2/LyiQ62W+0Ua26En5dZmNUuxXKwLJfU8v/C5O/PP60Bar1s8UpvGsL2GaFMNi7JIZlv
5xmB0Mvk3Z+pv1TxLiP49T1+2nnlMk9ELw4lTNFNTnw/RU2rpwcG+Sg6qr0Nj0MlWYM/ZdskPEWs
9rfgZI4N9nUrBuglKswmBQnSZMZnRVSrxvHfhHMQa+/97n1uPca1T7GWWYMXsoCKNZTONWjhsv1O
s4jZG+7Xsdjbhu7jXdZpOqP3EIezgMb+/ELPLZEtPkWxMFwSmjT6apbP4UCrAh1kGuKQnDQ5GsdB
aTZ4HhfvZP+CdQhKvRBrlx7z0Bv12mu8f7Tg/8hznuPEKOkVO8M6lEDh5sOx22yXjd+OV9KCD4pR
g85ci6fYmCH+M+yPI4IWYr7yxvmtNOZvcBhfA6L+YfuKHo4G4FFjS3blFMwXBuaeG/O9ojtSgwLd
Jj/SAyIG7aihn1vOmUwf7vu1O1GwsshFeXbTrP3TURG0swn5yhPKeDDHr6giMAs6QHkl90gNn5f7
amnNMYwmq4myKHs8io7YYCdJDzT847Gy9sXo2S3gxlb8VddP5XKyMwzJRlZSbRGBu/h+PrHrsCgR
FcVBY1E+zBaugHdqKBSX9JwC9jdmLe3mGaCDCpLv+BKK/hpy7Oh14ykTO4eholnyiLOrK+1LrSW8
0Y7qORIKcS7aZ0qVaWq1eMR3rVaXtvwVkqRQxlNeyqYzI/BYdzqxXguWm8GkK/cdbvo6dM0njEZS
/BuEBlAOVPomCRajGUMoSoJiLhZAYZabOviZtSSrBQw3YVUDotGrNiKy2XF0Yn2zM2sDCaxwTidO
1kCvuO1U6C9v5ZfMG9DdBd10FRuDN/ucYIP7Y4g+U9h1Jh9SwAB5EHGzsazkMJHJCv0NOYJ5LkSY
j+6Hx1nKSUgZiI1a3i70HUO8Ewzpo64UC6ibGoE4Ko44UmJfMj5LunjbkEb8pK9ZD0MKtqB+iqvZ
B4M/Vn0GOl6IWEsL/DrSLCpBxOpnXmLVXWwR9r3449UQA7irwXri36D0G4jTLkBvxrnuMsZb9F4R
lchFPrWB8L8dBll7IyMXi7rbGu6JY3JtQq3yHQzHWW1e4XHICTLtWixusNfHZ/hXACY95wxpReQ3
4jyg8a2SYfwH5iiFBguHOMs54IwEIEf2Gxk5BEDC4tu7CmiC5U2JObHLij2Y6dEuzWYN8YA+59S2
soeABul/a2jtyLGL4ct1MWjh1r04i8qKM+r0eMBqeAjjo7du70+EPNAEgj6kblTuP6TelNimuCRx
pWEv98+gzEtrwmc978Fzh8uBWalXUtci7xOq/D7YU+SGk00QGb5fWNiNqsIxlJr18KqpL/JTu6aN
NTF9sx4sS3s3COEFVaSYb82YpFFOfjFH0mtOlwDxRzcBozluN5BLu/O/V872opd9IIY5DxOrGr1S
EDNICd5owIRt4yO9X2CcLvIqhKbLJCcPiPNWUinQ07DKWrZ2cw2xX93hfsUT4o7N9IanH8T5TobX
8DTnKSOSB8OOo1WBOO6qrcnOjKcFGxyMp0PZFeuVO628/9kO+dYT0bXfPJLnAeazlDZs6z3PfSzK
anMzLO1X1tKiwG+LMt9V6lqCJFcgroSOaEgBeB+MXKkAbhhNGO9hwnW+WU3avMxd4U1oSgMUuYBN
zPzZ3xi/x8FljFOpRt069GdKSHkD2OJtt4jFiqX8YczR6kXw6oy/oiqa8/o+e42joL1W7iw9rRBN
skCYw5z48RtFgntvOscfSHT0+PO+gjVE2e8jAx3N/Lia1RvZBsfltyq7rHgwuRzI2jnlVrSxs2FP
eA5/2T1K7hNM5g/5pLcOP8XU/VsYKEBho4Ido8vsL6Zdft1V4hzWqts56WgCpgFrOxDG7mnCBq3H
x5H8OapOFGIpiWlzsyXaLETPZbwe1RpKoefZUroqmMTo3aFFtkzZqKklH6zIjFX79wIF32ChvH3t
H8fZ4a8LFewxdwjfqxZeB9cvAwoZUVuKHPe0vBmghCb4X/QMOe1D/CMQCA8SjhrZFWhWwT2Lme+K
4vAjYevjhJ/9NblJumAzO9LjbdmK3MqnB4+dMYJ9c5iLyLrIz5syhgKw0N7AVwdxQX8z6zdh+30G
Xm73RAQkZBKqz+cwF7k4nr12gYc3AQaRi/nFLdEdtGxDZpsCcPwn9ISLRVCjpsmkMcndmuRDZjWG
SUKAT7q+P32yw8gkH5bPy8Jp7SHSyRaFeW4rrGknltpUfyuwsgEIXjIV2hC4CBYgKaYJlzHaTNBq
FitcXyK9gGwjhk2GmIxPWwGS6K965Rcz1HnpioHJEknX++Y3dufBfMFuxu8Ftp9MwI71Pk3ox9Ta
H2Dpvftgcbm7g2hew0AW2aFXFrnCXpAGfKWglA8fnla23FTOaI4ariU7AcALAqIT+qxVX8E81AkT
54wwdZWqs0koGxr9ZhTBmOCJifb8Hdyz7t3lDw0F7I44cF9C6Ep4+ByXg6/43Ar7TITGz0iLAXFX
/TngyO66j+hZaQSSdJRhC9fRtbAf4gIOEEXmIwwy4TJa9D/E6FlWaGM6HC+a0KbBriLRV8s9aO1g
dzrv2iVow64e+xM+4SlUVP6eG1iYdoyIRp9ChVUYzBidHcoxOk5VhX5x6TsNxic6v7GNCrbAjWMx
4kAdodeBwvdMSr+Ba3G0XwbX2dD8jddp5y2s0H8YkDCXR4WEue6YXdZNtlOpEyRseOXeaNxPZh8o
jBcizPZ+dZQNP1Ljj9UR6o9iwMwFSN11VB5WVueziMP3uNxafoNjeDvhCKaOfycbu1CfXV4/JhOT
ovqxKqlmn1Huu0V8D2G5nb5K3IRNissbWaKNIjT2FiktYIpJZYYJrERjQGotLbP2qBweGOHGhQtP
hyTWWfybDHirflazNTN5XucrgS4ttRSyRbxTtowFHzo+VNbmr7yAUqBqMl5uD6hOlXgmj99WQGsj
yg8OvPzLKuKcCaqSmYvvsML9x5qa0MAA5Hhve74RNSHpBskkNd+oa0070pHvRjiACglt6qb3xp0W
ENHrp/1FS5UXnFHC/45uX4tuGYbamYPHCSm1DRao9yqsZtDW6FKm5brDVUv1n4WEpGGu+cEGcHqi
9FIahqZVKA5gAjSNJYqTJmLqLJgizH597n+5OiL7f40JuRNZRj2tdGcWP8lNaueQt34sARncKYcv
V6FG6NtzUTbU6awj7SkeY+VM9I4YfH0PWAFrNjgt4UQM47SGhEbL4rpfqGqqC+RR8MhQkLORgjEq
pfolwF7gCi64bj17maZvSCDSE/mzZU0Q6IpmbMucbmrlQhb0VYV2nb2dzzTBVKryBS+lwEAnf0XB
USM7lfP+I1pJj+iPm4xXRC3+eUKz8SEpQ2aI7AntDN+FaShbT2ZV1BAZZMqK6UgsS2nOyWJrocor
mr1vm6BXS/fbdZOOzy+gi3/5Qy8uWZTov0N038XSdRbFYKmRv6Ol25fZVajJM20e1tBcNB5XlNxh
3W66Lc0NT9OO2Sz+N8LVl6+9e8vtdhk4edTmpTOhKh5CsoW0qGPxzP++SQOwN2HjBU3ukTxgxB9z
Nk4hbrrGrfTZGSMJ2GPrlYQ3Kx3vxgoPUlu9n7HihJpYOqbZcsTGwY5uy0Exx4df4ecLoyPJudya
y4TClpykLPe17M3uIHvMPNy9Xk1RQoZ0ob/frfIUiL83xZLqQp40fnH6a+aDSM24nm1w6n0pL1SK
N1O7uZrpUZ54aDO9TI5nwcdfpyr6iNxSCsrDbEiJ117hbUpgD3d0rG3w45RwGzttJCpTyy9AmTlq
l3RL7yjqBXGUU4+1ClrcHbB4PH6/yHtEb7Ll0aLJBL9bYd079hgedsh+fwiseFKcdYVZbWvorErV
ZpCGKQFGUoCws7otLqkMF5B15oiZWhG04bGq75FyAK3CjYathkBdaOX5/MhkARbzGIK77whMR2ky
FoJ7LgVJ9INQ90tF/GHRWKfKfr2ZKPmhnNZWiytXebYVHDFMvXPR/goixgppQYgt3Ng4CwWB8b9U
E3RNBWjrXD7D8rlkvw45aDPnj7mKd7AZX8JDM4aJcIGIHrPCB1wij9mKTHJ4LjO5C9xASfuJEtNk
2D+CaxFvmrWk4U2GjWDUFW3w1v5pEetxCv5NZDNSCT5CgLVatfgE4lulkJWEMQtdQZiyeOC8FH03
NbskXy+oY1HmDrC0t3Bw2+PqJo7hss6vnAzkk9dtbWixIXazrU3xS+8I1zYOZlECAtbVY7/XwcHr
MMAg4aXbBln5/8LA/AqMpAO3fyor9gZPDtTyp/P+Jymh/geynO0DeNQBdKDgD00mehGp4TeP4Xhk
E9DhNMZ4v168uj0VxnJFx8wrAQKA3bvCqJYnTTZpKuhCqlv806nNDn9hsaRDY4Jt1+qdnGA9ipYp
CLW0MfmQiYD8lV0O0ZtFSV4lgx6mN4rQkqBcExV+ep4OztfwMVAEgdlSQX0GavEtIZNl0sp7hB2F
1dfVvGShh/vlLh/hduoBHb3Xj8cceGAQjKOL8/WqE2DU8yfwmmOQvtKIDGxI6yGP/xhVVbQ2EJac
0VOTe97h/zGeQ/BK14mIltED4eKP1AL5dlOuDWlOIScDxc5SM+xpQsfSEF0zpnvikJQ6dwZ6hqnN
b2De9ZgIleCK+vZDeqTdJRXF7PK+Gj2Pa7bQlsBJlklXecaiiPeHK799eanL8aXwGvUklyMl1H37
fy7Q3d+j71QGo02/bitgePAs+1BlE/rHpIqfDWOhPK4FBEAHjVLVNixFNj9juBpJmammZWjrkcGb
UxDR3iPN2qYwGCvgwFtiZoULtrmbc1JpHpWByWjiWS1fDE4TRX2orrfHpABOVF3n/mpWTfdjvn/K
rvTvBc0q6KRfuHrAzsXB0G/skU2qrSGY72ib736nEsd/D105Brxfu0dj9glyok/0v7Ut/AXJYgEB
u4yr0FYetHObAf0OcoYKO2GonCGqpfE6eiO9hK7BIQZYHG9x7fy+VIoG0Jk9mf4AJzlJbHzH+t8s
QiORyCfL1u2Fu9Xsdeft9zyILH1Llql8aDYJG8qX6XLqFvPHAuT1uDyO2yFL/f7ADIWQEzf4ZV7I
LChD3Ohh2vtoDPz7Ymh1g8xARwHw7sBpm/UmAeNiQzAqRbGSqgtqWFjtZ9b1Wc/05FsR3Jchr4dZ
EcajDoPGLLNTmMiTOEKSR78zlQCKWjXExAWOXL+7Cmjje3LUZr8E2ns5kElmddWPlbR305DDWDFP
QBL2J6GSKzEFkZ78vXN5QjWx3zA49M4bg5oE/9XlXwqeO3MsQ9DGfOmXj48p1ADdRM3pBInGtivZ
X9GM5OOAoHLwMbKR2DEF/vi7JMgeH0sIp+tuMeoEhoxkNnQX3zbQBMyMrcQ4oElTLBg4cTDto03t
EJuDio4R054DUT8eQukY+BWqUIvLND34Hjy5OKZ6tSJajMbEzq/JmztAryXOzqq33+EHSFF/LLZU
20P65vAqg29njbWmoVsNDSoaV7HLy4J0tCRrzS4Xdgccd2Q1iu4cfgnr/VR97zMZ5lDHt5zrVJfw
7MebJ7Na1IgIwA71auMX5X5mwtVgMYRFQMidx2dyHhEUgEx2nzLF7kRKIkuMa18sjncQoU5JYIei
MqLw0TPeU+SevArkjWlc7q4nUI9GZOJjoXmYdIwi/OuojIK+AushkhqCn/1GVOk1mJJqtdsSeBO4
KMIuszUO8FYbfEaVmLpTdKzM9V1hB4H5hY7QjfAQ0IqnTAAd5ZiWplpFB9PuIa6pKLlZALPYfkSj
Fhzp0/jqqwGGltPYhfHMRB+4+VrrXEPv2YEepAqYEIz4/iCNA4JttnpMlnN7gre00J1F9pzCAtaz
qfc1qinUv5KSrEY5KmQYtDRvMfSh1BzIq2QKr0vCPEjLWq0Sto7fNb9SxIBWAHhJ47aH0LMh/48B
gxczA0enXWB+y2ktlk0EBFgvS3pbL/Ve+kfQg7qUXvFrg6/tGpApnwwoars0+e6YotqL8I23UQTD
+xPMkyEs/UC94oWygwgKN/9UZ4hn9PncTlSfSan0g5lJTyQhIp8DGQfFM1htghPnk9smvH86SM0J
2SXPLaxllCgx3c4O6dzqU22M8e9hUO6GXrqxtVH+Y8Ib5IS8ZAPZf/TqqSj/FW3GwVr8bkdXm2Pe
JRQ7a6+Ungd1oZQzDeO0M+01hYpNUMObseiTa5VIf1RYE8Ocv/ybuWjeQhgxddWK4TB9J5xCmw6k
y+UV+QHWMXTzj9Uns6irFIw9iFK39tPuIMhjM6HFq9GTYFJcyTQmFaJ336Ce+yiPUJzWSzRvE58F
7knP0MlyJAUMIgOUqVi/JBsAqhRQBBfMhEo0g4o5ZxeaBhutJTZbRXPdxcpmyPeZmbTwcsm6zhnd
cLD45Rz/nGTSCo8sPzbvFf9g5n97oJgdW1KvEJAB+gNNP00qTK9R6Oc428zfvwMlSVKjfzBqDbfm
trFZ9zvL6lN+m6VCiFhvcNGaKTwhewzMINFLieUrryzcrTPjrT2okq40GpMkwyUQIBKAaL3OK6oF
yVHf0Nb40L4Nv/KzkCxtaDa7+jc5EpT2eRRFULWSkersXUCaUMKwQ/Hcz6XUgrPVZ77o1GYj2Hm1
UrH4JPFXGRrgEwaooLrMyonFzLsu0Xupx3XjgPbJHgJRj3zEzaFX/089lpfoFW3yVQPIOg0t7vB0
wWrpt1756rbDsbqxscViOwKqRGn18m16eNSv1h2cna6zWWxyBpQttY4lghL7fqfjh9Z/QHqKzXk7
V8dakI5nvDTfTcfAXXnDxQvYLYOjfWd4u0GK+OyIsfKUsoToNq4XeYl4MmNDMhQ7mLQKVx+rBs+9
WH+lmQ0gzr7uq2LnNCA7lMIWrgW0CRcJyXPVbyL2rtWEyl9wFNipvZWT7PnUuUQIff2i8XVvtfG0
BJUFPyI8TgsGJI6aDh5oCy1g2Jjpj2itgda/Wx/xyWeg1aFcfP7i/kQN6ubNfbx0aEpd11foxzWL
3yPMmAZUQ2ffvrAFEqe54JJq6e9zaF/WokEWf/cEuIWCROCTyI1mW+brTt0vV53Hb6yscaDsfyT0
I378LXJvmNOj8wt27w0fbBjz4ni+Qhaj2SScMNmlh3r8/qPkRX1emSzJh3awUu/cru2mkixOZfVJ
NfqZBd2jRah/fm7klgXlgYMFMG+Ja5hJWi3I8WwJ1sfuRE5w93gLMGbMv+xkpe7u19GVx34By2/G
NQBNXYiTF2k3GwXlZt5GO+kseulciRSfQHz+iv65F5M9jMqxy+86sJkakpEcLblLdWOzmfff3GsY
PrLTFaTi66PZexTHcJ1wFjLdw9xd68BiHkBvjQ2E2ILEyy17OotB7F3k9BNJS7ZzqBsL07Sh2Kdv
hlgH+Q9KA818SaqCpCJGohSp4pMpfrJUSY3egtSKmAHtgPBVwzdaFulfgHxzEbKWwHrIrDUvobHE
t2SGSH4QJZ2gOAFZxikmM2bHIf+u+r+1xRgGfjoZDApQzEaFklEElTOH6/H95J93oy8iOv7VYV2G
fYG0He59LB4FhOEfTxrwO/rl6UnWaWGejx1LCF72OGHEjUlB9iUH6uF0H5hAIdChYqNW3em3iDSx
16ZR3cpgoSgu6jYmVtv2rnkUqrx/oNz+mx7w3M95aaYfF/kH7jcHKJE+6uIQKvjGd8VXTg/nFFQ5
+UQ65b3nDGoXhsy8OO1OpHE4WRds0t1ZVWjSKwFHB3ADjyxUlFlENB1iiBzP33O3qFcEmkUv89J0
AfRkGI7OAZgTCy58b/IU0Mg2xEkbVSmxUNfoiXHXgnGMKu5Am+3AtZjzOJFIPU9XHTuzMdaa1zcT
jOWGshiR/jdHX6YyN1xJMLWImOkAamGMBQaBunc5fCHUvjbLYiX8JRw3uh8BzCduzS8x31aVAelr
42RmI5WG3CQcPJO9VklpvoeBNF7UB9pfqfY/OiTjSXaivO/nrCdfol3toc31AKXTsgIudR/7Xkc+
Em1TtSBCecpFH98ydBNpEVU7BrxdopCLz4QOI2U6W+Orsv3IKyg/3Vgvgt1gucGAplTqMT5ngqQh
RJfx+V37C433/Yk1UE/5rrqyIH4NwT1eIbaO6Bvug99aHofHHJRUA51qrpCICtMZTd+OD5lujlq/
EA4Gg974oLN7OSRsd9yL3Lrqx4YLb7cYtchfrVQE0ecYzyIkSDOCGxePzLwivBDikd4b2AWT+EXy
SPu/WV/vkxg6p3FrPgInRZ8Q2K92FLKQjlHGllIW0rsga7btRXrGfow5bRlwXHRWEugbo3HT9bsQ
cQm1WqBaVc9zOHRWczApJcYsyitFaa0eXk82PX5exjszOWy0bkdOrc4+uEZenScIA7KaXoViSrn3
BvTNHVyCKR/ktCqMpxizYYgL1hy7TkXENFLmDT+UGQA6KqO4TSpGVWiISRKZs83ITiZUKjjsfcBw
2Jg9RfmrWrb0d3xDMmumj7XfxP7ExGxDqZK4WOfEFq4gQc4WDPNgcuIErMAjdeMbVYI7NxjARITo
PndEYFG2Km408BdxD1TQYThX852MflhjZ7LfcV72BJo2GSEtUXeJoy/FPctR05HfqgIlAUuEoKP4
ZONAIlv/ksq1usksyHfr3SqrxQBrKoDZbWaWogUOGA1vVASKzoE9tDebfYZU5GE/BAXJrTR87tVy
ztziXrlNNu00cR2YpDd/mnOhHGL4+2DkCQGvXnImiYvyNLz7Ye6DrZ36uvqK3GZpSiRhSpetYkW0
6PkkEebfQzzBGZOr42fSbXdlVNDb6YVJ+FpQHen0RiYFG6iOxU4vlBvhl7sx8rgiZ0IPqWuLhNny
QuzNty6+KXoJ/n+4wM6rburLyIsEnNkzdB+hb7mmha9d6C7ZgWPDbR5Y6t//Xc+BVmU8KNIDxBF9
LR+47abLoNqPM+/PxJMI0AExznX991rV9Qf0cPZevdoYOAqtdoodlEqIiwMAdC9XtbaLjQz0bmoV
fQFbj+2ZIFTA5MJpccwZTZISngKCQZ9Nvtjm+pbzpnEW2NXMmiHuBOdvVis3McoDpPw+Cju1KHKR
PPQmgfGik/mtdcKS1i8qE53GTIMQLnWTOXURIBsTYP1dxjH4sCLzdQN2WwATs9nj9Yg6MVqW7uDG
xgDzIRdB0gdklsh6hhZ2tu0cj9uvWKCU97eNs9cAxkJjp/zvvE9jP4/Tdi4J38kQcPSk4djEn0IH
jQyLXpWQTpwCVd/NImI+9v9elBQF0QEicGxhe6AUYUq0ko7NR1voKh7BqOwzZ16M4QN0tg7aT2A3
+T/ovOPAUOVepD0kSFdfp2Q2Pt0/3RYgECusSO2QWapA2i0oHD6qNabGUqthQu+lFrvkVBlRxbX2
x5qyzjELtK3W8oOYtHYPyZGbcGu61yM7rZhwzH2uOIttKTLLlSb7TOXdz+I+tJc1ByOMxu18T+JQ
281bHngvPTmDJFKDzp1idG7e6GKzV2tWC9L26/KqoRfe+th2jUHDMtcPHwCdc7FNH3Xc+QJXDx+x
f7AHbpDTLdyv3w5wxyTMw7ly9evjpkFb1PLhY+z5H4uw9nzVfGCH9r4oZOJuab/7oU0y1jazsJbK
E+PXLCoHMkxcip0ASxG2Rd+livE0r3siVSHXePKpgt6Wv61DFml2gWJCxuJdPzwHRYt9nRxcP0H/
2IwNhy/p2G5mmLCkQ1Mx6/TR8XMKTb0y9+NKjVTTbLcWOejshEkTuGctLISSncDVRWU5Vao6Q9YY
GpSsl8MKRZEyMxgCw5jiZ5KvtkjDKKkPRCqoZDm4Hs/aot35Fb32RSY/nUKK7+WDym+qlD3/S3ru
W+sWhN23MBz7gEWw7AArStFM6JE57VhuCU4432WklqEyWI+NNcuxQhY4EPSf7SHqlTsG7fIhCGXR
hZsh/IqIzs5I/YhvrLQf1c06lx3p4/osChBXnIYY6YDMwb8Orbw5BBElAhVGwivzaIGOpsmp+oFG
/RSmrnnMP/7RH/lrHIi4j+MgqrIGOyTNWrm6nk8550+dEPQu7ecDJKpfdmnktbZRJNbUqMfho51v
t/BNOYb/tnMMhg6+5roAGRx/ayM64M3c5+OmQIGtzw/45KlJ9qE9qb51pvonUfEp2iyZ+xiDjgsH
Q7IsnxtBVYUQe4ILmlxFzOw6Z7P9ytnK+9ArvZZjTqllQtC3FRTJALAvO7+0eS+e2fFSM/R8UWNR
4YTXR+CMhQGo95k5ILrIXgu785VjOf69ZeMgGiEm02piExPQ3LM4Fekp9lhHaByiMhobQVyBtbOn
vaAp2zvft2VNY0lVvdeQ9NFt/Qeu+nGi/+M3v2gP03193vJGV1bBX4xEgDjnqPwZCvTJpGkOoEEh
b0JjrHGeHQ6mqSZOXCEPGqj2Sp9jdBjC2YsKVrUir0ScOK8iUCWuoJjIhNnhF3W3llClSLHXiPqM
Q98+ZqHmR5JGvh+2aOQMIw0ToF8DalOjLg1/lDl20LOQW7VDGrJQWSXcGFumMN5JHFEUedQF4PMe
iWYBNHCWD0YOrj2kzyPqUeXBxglGOmzvn71QFoHOR4GSwVhLSu5rps6MoRdY5FjGF1VWjyCh6QOo
NLKDaVEdFil1r6nOzwDsyuTjOA97ZZ7Y7+b2MGidjpjoMIn0FVcAJ794rU7z0AND0xDMSsajwbiA
44OYTiv0n2XVdPlmJReDa5aDc7YJmSJIqvEqcV8cQf3wWxwRYxAmjj2DBql8CrhdeaLBUloXyk6F
kbHQGr+RPpHEmYjj6AoKD6EXILc3nAKr5WTJnuB+/azhZ+dRvQL1ckBTwBiusYXoMDcuHbIRDERT
bEjo57RHB+QSOTSoPAOZrXvClWKdT7h8/Wj0GkrTkfXQyAaz63N+o7RaZI/29MyglPLrzmXUUl+V
k/AI9FbEkXALUfydnX7cVHmWrTwENPoXMvv94MPyUq3W15S5ikJqSVcSWe1hGh976gzKqUdHMk60
MsUbg/Jq/l+CBFc4qRucP97AUyKbkNxkd8fmC+LwfmlENKfRNIqNfRuxgocg8yr5pFlIyKcUN0U1
RvvyQ8Gt2N4Fc77B1TN31FA2qdRii7mHjdBtaDZqd6UGF6imuRKC2AwKU2voB75Q1kCC6NyF6lon
9hkv6Usiuiv9BE2SvH8zIYpPp1kAuUjBr9jv5sCFQd75FKCpDRqA9ve5GXlMFfxxxc1n0dDT6LuP
1ayqal5QBDtSjwfbA3qsFEe4GMdChRE/V2XMYdd8+t//4o+4qtsvPfz7yu4pikV9Af0LJeg0zMia
7eXKdCP6gjGnOU9AzW2lfnoAoFLpb0qU/iceKcwKRqof9H7wjlngxeUg0VVbbemgL77ZJva17H2n
ItQIpsvPtLBnyH8uSjfyjU3j1coB/sZ4ZYyJupmaGshUYhHBkHmF6+MOKhK9LSanavcBcGYD1bnT
EZc1hWT1no8BeK7Z3KNquuEdrarjJhA5+JhYPkVJ5M9+UYF7k/PH8RwhzVzD6ZmcU4f0ZJcXvCLx
I4/48fBDy2o62m5Db8qFmjfsG6MR+15vbr89DVTI1vhX8ytmmai6MQ2jz4iddwqZ934MduLlyo8c
bBNpW4OZGvo8k0sbBZFK4ro17DlACsO+Ha8k2HzGODaw1cn6bdwhi2lxwtyPRBfrA4YGGthy0IG0
/NoRnAxu9FYlPTWK41kJ5hXODMa3e5EN9ovXoHa6peFWjBn27IR7II/fdOLzfdR4Koirf6TJMmOV
VetQEE7MyZCJh/avS4y/TDr92XGQb2xXpInD4Dnr+8mZ44+vX2T5kKy3djgZfQmnl3jNcnFOzXne
TrL4JBt7lZ/yEu9/hwD8N11UZbh/j9XIpWBZbQwUI/KKfhqWfU36V+QrUvc/koUPeH/o5Yhm5F2y
WXfWevSaO6JThPH3iIGXdzhg7xDfDrKbeXVC66vd6sJugNk2hv0aabRV7WDo6Y6z4c7lunrxEp/M
ygvQBUzIgEMPLVRVl3ykmpEEixC5L63w8dZozUQMCkarzfB8lxWkgNKk4mrVDEbHg1wWPHsnzAjP
2wieQqTiFf8Y51nYCl2SzfWj/xXJWFxWJ4HD775V8GlJoDwoXciY+/LvfOBFKh4A9DFPd2Gxgb/o
t1EvxCBzp0SJpXyquf/4YL1FYlGuZge9ETgrTOEOQU1Ryq2IQasuIwUHsk4gnGKrRWRCj/YFGo4Q
YdyGx0kA+uIkHrGCL172B+Ggp5VYTLW/X2Yvi07Yx6C4bi28uy66te0zzf1GrPjpg3rfO1uszKXA
PmzyN6/u9PXv8Ojw4Eg19lTHGWIPbpuABYFCMW3DlVp/8TPyWf2TiT4WRvvoiAVNA4zQGnAm7ijZ
R0XsmHEpz1xF0mM+VrW6gylvTQola0zAE/q42WZLl2yzHHBX4aa9oLtR2l3aUmz/4CefW3cnnfJU
+wnCKhTlgtrdYsrXvQmCjLu4o+GEwO+GyQWFdbgc+eUrQ1t4JLu5Zc0XRAj/6JkQ591Gt84Stx9r
nM6pwnAU2POSxYG1iOlH3A6aVHC/LPW+0ok6bOAGAbkVKnD+mBkVhuI+/YqJ+ipVVlbGiNGRgPlp
f12DB/3yxJsptEsEx3YwsGp/WYK2CcUhRwiD/B/0sIe06+JFcHjHFVg6RbudgWjV88T/DT5W9mB1
slW8cTsoiHaDMmEDHeY8pliq13MzEmngoGiflGT5yOgqclkyaRRyCF2BcEmoInogAIHTMHZseQcB
zI6ohG2oL4uwozROgNGqzmu4GktQDjcKyj0Dys+2q4k+R7FEqnaxOMuR6kbjXKrNtdiVwUiDp5uB
4TofWwFhpvyKXdQmwhNmjjEc86/wLaxUjSKGsDRbm4C1xmDLJa83HgK3rnY7E3cl2GdZWKMS1H4R
xUXk7mAOK8RWuqQMqqcE292RkBegN6V/Ij4SKbZMXYIGF7u25/J7+Vf9gPmtcFm04o2gBJXCKZEy
A1+NJEnBJY24Q6VJxKRTDde6f0Eca8tnQndg91h6yJSjrgeyrlSbF7gcRbHKrbsZ5lFsvcbpsfMq
t7uuOLOEySe6mR3eFTwWs0dhFCrD/xKAL/rmWCwMNPdxL4P3+D5QFgLE9qmKjopMAwl1Osh9ZyeI
4hqsL0vwJBbM071orIc8bZQH4eIqR02o+mPbqUKGEqgOVVaN8jUqSslJQKblKKEMvYPOt/3pcmAx
m8aw9Nt/MMhV4R3MaFENG88DklmVvvA4gwxDG40UplP3c3+DMkXhTE37JAtGU5lHPzKvU2Of2z6m
7YHOzIyGpA0tIgk0iFUWOPX0E5DkJspb9nSrP/IPLF6ItRJjIEw7xdX9AfyKBQhPd7faLoJNhF7v
pCJF0zThMr0hTQbUzrBkJAZcFrbTLPKyT5geVQwoLCNJogc2woAxpH7SPCEMWQV0E/v/AgW+hc4E
wW9maFxIHJhYLzQXzWKiJ7na1JXNlXjTh8gAlqC6Cp7fGxa+/XSYS0fslVEf3GQ6hwxflUDD/D5M
fCTGHXcnv44lyLHD+ntUICN79HTplBxY60p/0ooShRyOYP7rs/2V8XpFcZJN01l1yzhtzzvWa4BW
rd+wn8CZzw0WV5Aclc64svidv15NVfXjW0F/kfurkD8lOuBOV4o8uOa0r34j1mh9sdrIbLPLlFXB
16IhOrm3H/5InmyvQz/4ID0eM/nWdOxxMvRT5I8dE6DfKSCJ5SY2cUQxSjI4xirV23n3W/Fjeryz
RP15QrsL8angbafmgL05NZz0RFTitoip61OlmYfCNnJAvR+a+SovOZZJuqBIFfAF5FYI/kKZwXd+
m4rQ1ZVcmfYGHseD4X+7L/uGdt1oIOSDMCt2BMuT6VVL3w+Xkmg5q6sqSua50fmVOmkfgYxQa3rA
nhmH3iHaQGPHLRkUqtf7K/Q2pZskU6X+xSK7ElFk+oprmnJqNZ9HQbqdF196qt0iEBmHlCLdFAtw
i2Om9fYdmw/cK03Nt3E5I6ERLkPQLJ5Ro7I210JHQ0yZDq3FXp7JdNC2LCwzf/5igUI5SG1B0lLr
+w9hFuuUcZA7Ed6+FGUlAQLpbn8X9/UXbBJ3d857nrXPl+dlz6Sx94G3MJZKirOcGZf0fvPG15Ro
/oYsy8ASQTIgDp2H4iFp75tPdM1/hqBc2m2Qi+Hyb8SPunNoB85AX2sFxt/xsPQfGrtzPxWd7R54
hOgUox3wl2DVacRrTxQ/FWkBwoOD8FyRd0Juh7rcO31LzVEPQ+pjrvdUT7YRUp//uXPcQURRb1Hg
iejVr/NSkV1UdR6SyczFD3oneDFU+T+SxLIcJ1XMSE9lNGRtiAt6AEkR3qBmeom7UmIyXBerkayV
PYCX7A2zZKYsg1SxeGEHHDAC2fXbRMUlacp8+dKDZN7oDWwuqVQivV5ZEhjq4Plf82rGtpAQp5QW
ogm5FTWXFtL38Hk1cvU3wCtIMuVpatZjPnOafQ9Tt1EEwxs9hlDPIIZt2yZ0gZYgh6sL5KCweLw5
SkQ+rbLee4wiadhOIQwpsotI1TZwBDttw7Js7afr9VZhed0LEzbcgNbggVoXjM0T3aGfVrp2T4zu
VIrHRl4obPSSY6oMnsPEmJ8KW2m1UpPf896uu43uueItzXTyFmZ8kHEceg2WgSYZinqXL//2rrqW
JQjRTNJ9IAf0+d1l+y0gH0HnrdpV5NvslEnmDTSyBYhiWiaAYXiRPK7Cp/PLQQtXLOvIJ8NNWxD3
JlkY9IVvsVqUJhkLST0UhFnHA+1sxmEKkvRuim2Xub31VdobwmY+9SE4E9Cbnq31+8WxSohwy6Dc
Q4Qcm7egKpCBwnzA93E/Q6RXQaP0jMZE57hFbGt3YsUdyiO+6eL/j1RwMNlwCitoiUXPW1DqOUQy
BBMuzQUghBHt487S+9jfysHuSYA9owVWASo5n5IQIVmQCBUAST/q0rfPhBPvRnCckPS3yIUnuaSr
Di1rk2dWRODyjucEv/NGfntGWmUWJUMbh83mJ/b2RK30rQ55jBygh8SqiuZzg5d391UXbTFxu4AY
H87uhBhiVE8P8tBEyFtSdI8Jtk+Z1xSHb4l44JOqDl48JGK4g5V20HlTI3odutXWMgH0P38AVqjb
ZZligVsKRenvNvaADL1mYY5+YzRpcKKuQ3OBXMNebS9/vp0lnZogeY/rdgrNLElQm0Y5Kp2amBVI
ttlsKzdfDur2ubUzbdKqt/jkvolNXbwzTdfEBSI6YqVvRY932fMELFbVTAAwpYWusJfFleylDuc2
FZ0shgFarN3S19uTsPy6ZFuNilHmM04fFxcFihz8eLumrYNymkJMeXSEqMrOJcuZgfW+UOkj9uOe
UQGdwGgcOwqRFw8GFXHOdVlnGSB39FiNnntKJsXGIneGCjmOXG9yPZhWFuw+hPVHzCBm5PEdI2gr
QRAsRZ4nrpWe5hthuHghp5vcvy19z07ngzn5CO9lg4sAo8FlYasGm5PiuE1fHrd6XDlrSNAQJp8s
hpLMblA1Cu/AcywUbvju8YFPY1DPnWoIXZdcTHtkIhdXUArzNPAx49QERYsinsuLaZ+xxy8wej9R
DjaNmkHU/oqHAv7rYcmamaigFY1lAp/ma6QL6eiFW5w+pAAjK6giiFwyhM7+TVDiqh+snQMqhtbG
HsK7D6LrfCzsmXT7JoLplXrj/rFCUOE03hnAkJvp00Zdyi1ceCo8WAkXe9zRTUUfR6gXStKfgzA2
pGG1ZF5uI5gk9/bc0s2D6HzTKYPpyr0xHuLwYYzK/s4sT5pEI1u9QsXrKJ+BXDCDJr7pt+Drj9SQ
pdbgz8etTpnUt/HJnoS4VMUp79e0Sv8vBNAoSok+3rKuk+DxeGu4oltoLIWEjZuhq+BkxIQI+WPZ
nkzLgLP2QdbtCOkuH9/QsofdiMLl+wS16aUA2BdxhBOhwZp2IwpWya/cLmldciTrJ0nydlwjJG0E
2LGGkjr6MyYKblNTyNpmVMAzBEGvhSpCg7i0YsK2E5drItoSr61u6Uim4RhQpw+9PAIS8dsTWbQ6
BbhvZCk5LAitDV/ZU8YFHMKNAM2AaiavQL5NizaRGVp3js+HNp863+cS3LvGKF8PbDCPS+xQgvBo
gFIDN2A/Ttblu9KGjnsZqdCS3UVdAtn4196XxheKEp9ZFCpd7RNpKQ1Jim1eLyIJO0maPtR3/39p
ygMVqg33EKVLe1Ff/t546SuTEaoAuUGuOXaY56BPgHPpYIwpTbJDnz8Z2Jrr6/pwTX878L5TBnXE
0X4HhaJ5+Uig2nBbucEjjf/SWgYWd6HSdNBV4b7hd862stiUuFW4p3BDWE8BcDVptOOpDEtmHJaG
2CtSDLkTdbpVCT/p58pkaSKAp/oDH8Mmsy8A4LMf06a1/6PZZuoIQFn4ryEjGbP8RXFswlbQS49S
74r3UrNloFL3lbVJ2RraotzeEvhC7FHgesnxmJMEJJx/I2k5QHKuyMDh3cKM3U0X0T7tqhRZKkYa
4K4ugzvY/YTPpgZ0/2JXvs0XwGYBfYlUSZVMbHrmCB3U3ac764kn2rf384TcGAyfeI7quwRD7unl
Qscha8PqK+sTvb29Kydn/NLz64GJtqIDmyk5QQt0+cQwbnW3DQ7RC+uayw2xIFf7M8aSbHta0Jt5
o0W44QPC00KGSfmMXoyz4X6/y2pz+AZ0pqe6wUMZRLB5gkRbPx6Gq2jkd3d0mu2ZGEBUFW6156Un
MONIKw9zOmB+ftEUjMSuvOlqwMhOErRBNWNKWx3Mksru0Ki6SgGubMKTQS4SfhzFl9JMdcNZ4jpK
9mjvEXXuvexBtJ2wtFOqG9zFpFm1lnJ5rv51zYoFdopUWOSCJNQ4OdeBBgJORLFD6XX+WRUmrFnS
8A20itUyd1FWlK0w8sd1j/fCR4D5HkjUeyStmTEVt8Uy0BzmspFs3cbs6XFD7x7N48ALxk0gG8P3
793EIaVouaKRAVSrZf+wI56TNjb8kMAZ52ySz1nor8c9ek214nowZn9+YxIaxur/YA6VymWvmEGd
DkN83kUVQ4zSE6OVED+XMk+KW9oIWS6wfKG/FDyNVdlJxchvy55NgKlN+AmhtaEl2LY6gp/7hocv
JPZEmRt31XioJ0BnnSATitWCnSY2ha8+yYQvZteM5EtW8z8sAi/Sr2+GmVwDwOEIqn/l50/KWxRn
KccKwiseLu6urs5XMpCYeDTBOo40s3IijdlXkSUTIySKxf0INmrpfqaGku1PuaO2e3qxndtTtN17
+IZEef4vLT6npuh1WCDKaYR+1SjcQlIqqnObEjJHkp21TLQjFqsUlo1VnPp7ggfue1y1FIzuCY0e
bJRJ7SikmxGL4NpWlNmgnLBVnrX/6IUgXspgtJeN7Rj2/jHDy6KZiAu+njgK7ncMIQn84tUz2/bn
/u9UubakpGeob4/YM04I5WBYNMp36NP5VWU7miUn+rc3SCTKjyIoMBlR9k+2tcSYbbHiAiDEQ+3R
RqMNeUzhr9eakteU8FPwmGquWcQLbFgv6nQWEz/kRz+mgDSHPu61vhTLXRWdyJfo1Yez9erKD1F9
hflUtBjcecj2fnP3upVwxXkjLr72rofWMamHc+Hn714ITULqEziyKJbHceS2FHaKUdnNeW7QEm7e
IIDpdNxdKjybbSR4ILif/4GkzWRLJG/jW49IAq7pvt3SMftU/GoaJt/dF/t8IOKyC2YkUFN1H6Lv
thVrw/sGWb+lcUdNmvkh9d6y9WJC1slp2GzmJ5YRZ2RYTu3MDbmV5FVQBlCOIbP07X7e6Q9GRnPN
qneB95Mio/GWdzRXVw4wJr3e5DrFdNcSDu+K0on7bmTTgF6Z5IkuHlugeVL9kqfgYiZFFVPRlCu2
TG8O+QJjqil+1IhzvZMUOOD+x2XXeni7IN9mtMpI8zTNWrhTkcGyuAL6BdZ5wmkb7fodd84yUL6Q
2wYi0cINdUezJB29HGABkmP/vRh/cQsNbIz1R+GzjobhN4gu4FPec1oIkznZT+OX0Ts4c8xylD9z
AbzNlhp41cWvJCm6YkIzaQnBQfXkxh045MnE6JyWQytspZeetuIXalENkxRF2k4QZcYRDgLCyaPo
HCTf092IK4Lx/JZS1+dbJkzwPxhnOaLiYuD+yzJpsR+PtGjtuW1R8yOjgCl7GJAzu+G9vF5MFuFl
cNIHrU0sfjbj9Ku3dHLglxiPyxBARX/7W91KWh33TKNuz+nZaUIkYHiHErBkCVh5bwQGtIIxAoXL
noDSkqzL9slKDtvCEq5Qkk0o0wNY9Gex1gTXJ7AMsnBuWfkUe/ehARCPnwdp7DS37C6B0rFN9gBV
hEdi0j1GDWtIWztS5t9+Jb0LAC3g4eUuxVMuGqaREspi4g6623PwhUbrhxiUOLHGR/YG72eK/i2N
8DM3pcaHsUgRAG+0v3eZ/XSHYlOZtHWVMy90fd3KbAJIZdEMEvk5TrSJrnYZdHtB2+QTrQvDuqYN
hSJdezcSsNobl8cPThiTy/S3leSzqIlJ8L3cTFjvwuqxltq3HZmE1DLtOsTw8G35Hpp8+y2pZdUW
KBgzdZ201Yky6dMCLo9kEQAhhGNlSjavYkfGS+80EFKBIbIDRsEdaDl9gjjhuGWj7CrYHMVCMv9S
60FA0ONnvgHOukSwFsJWNc3nnKlhY1twXMXcns8iGjrHCUCwcxAIbW0gJGr4IUdwf86WpOmhIB0w
ZS1LQ66bHaZfMCmWgOIJ0t4pOK1vDZpscIl8BLh4eSb6YNNDWIU/NtK1Jcfrd2AgoyHvby9b4ka+
FbwD9lZY2xhgjrIQu5RcS0j8PyYuVGb8yb6Rf2/P6U497pk8A9nAXS3vMMRnxRiEaBcuGYamigwP
lUour89mSe9GrgYoEiCpN82KXNlioZksk3fkypUZUMIo2YiR271RwN7j2Zjn2MsL47e8EkdREuYc
WZEQQgAF+ZE0kcRYb/3JzloawweGnf4nXMbw+N7XtPI732yuDAVu+2KcpP0/EqA6shKsJKODk6C2
3Jsn3lR6SzE/nq3odNDRAw5ZPBDRIyWSCAIxzJvZOPOtPfVS9Sjx1dOOxc06DSFBt5DjAOcQVSVl
p6gmwUVL+JHWKMc61l0fK1pcDk+Ti6VwScOsFpKU0n4RhEZ57/naLYqQIz+UOJ+IaDFW8Fp91V3J
HNdsTNqZ+JmpqNpnQRjZj5Gr0XGuRx+vzRMEcpmF75PDwvF73dcwzlmmWsfd6SUIKe1nuxkRDmrG
lh6mZ2d9u1zyT2584ZObTPf7ImOTCtpGpd0anAEMGhse9r7A6QizfgHaMTNItYnHsvmqzY0WZSyu
tCNO/ZNC+fFWs9oQ632EnUf07QPf8bfRxP8o1QsrD1Wbti4bsGzerf3Y9lt4Ewo0jZ11geqx22sB
Vy5BLuviHLva0HeMytuX7n5/IIgDvQtf0h/mAHYx7Fv/zvTakTzVCaFpY2ZFB2dIUirdPJS7tYyh
cvQPmTAcdpC3DVLg3V887Zcv1TlRDCVVlwiAxXuRUULdmPipMBK05knQxnqDexNX5+2TahkrCrzE
jCqU5N56PtYSmE0e6StcCZcrywk9pUMjuvP0VBNQlhMK6wTPQtLrCvBHV7GJN7peii2nMTL9+HZK
S2Am4HCaCJ/EFhSrRHGWlCi9Pu3qIADxsd6eMv+C66ndatNTZVH03+G4k2CU9BEln+QTIxFuS2p4
AfRQDYLPPI/Hdlm2N8VdiDFpJ+hRZuehx2YPLhMmaHzs8Ez8CKGna3jUiuMO7ftdKSmAnUkI8X8r
SsRQxRE5QmL0a+SJ2Iaho/VuGKRMACpSyB8oJNdDilpyS9ul1NoC0cZtGwByzULx09KhVJ8WE8MD
X289K+Qq2TAHW0QRU/xZYFmUGH4QzADa+6PNu6cRrV5T9uTiXsUa6qnG0K793O7ODy7hH4lvVZR0
mm0mbn/mqWBt5F5jjMT7IwkJilq69YEA7WfMzwPJjure3IlfTWqLCGLWZY543jebpyVpFStzKqM0
4/Xk/SSOQfjNjbIpFFqLLAAZsUz2doP5gDDOObnRanooP+5UVni6dxqu6c/gm37GTK8rtny+4ZlT
LeYwwlsadAP+AZyi2miiFDCkf2DRMIMNjQFnY4qtf88q5RrwPEFo4NIOuUWzLNk8w45rIi15wJ+f
Y5kk7+lWJwfEXiZsz23F35WttuHQO5ijmBvB60AjFnNPTn8xiFqiO5YS241YgVp+vqDj8iUkqwA3
zUs7r30ySGM566glwF8fWkqGSxFxWA8PXiWlr44mAJCm9047j5eKVV3zTxrFZm7pYWFBWIXJWbf0
U4QV74+SpGXDJgmDcx8GP8feWB1sg8BQ7CRw0zC8KislfXOVTW9j6zK3/gVYL0nfaVni69e2G/15
aADmOndoj7oh8NrkpDHzvI9G+T+52B1yGvOmPabhVDc1v73pGw40ElYXvTY5FUVnbewG5CkG9/uY
KiAPX6TdAoQseVSh+qNDa/rEcRNKG5TU4bmNCFP2jGzHyT/mbvgLrrZllL5uG35N9unZ56dKDljI
zG9/tBcim/hXufoL8afXmBsOd4efn2McG8FkTPA6fgsF9yLEQU/wbAewvsmO5lRJLBak8ihq3O2h
Ys7n/AlhAOSyAbLJK57KZ2DOuxKQkJtEmsjdC5G58B+KnMdyaGUPwyBM92wInkH23SGu46untOXX
pZmppiwHVzfais52tCQnenjTlipojHlM3bmLCg+EQ6ckb7NLZ1jXJXtLj2o0hSEC+Te1+ZY6JU5K
0S3lTPspd+pd3PqYqm/BZ70QjQKaKivIlOWp++O4p7o7DJUJhq7Ktq4SPZ7M7qTF6MRc3hvZ/Ony
ebBAT3ET2I9siDdb8DzzzGgGwGKQGgjICMD2WKuYlhynsuUvwiNXkWUMp0aYAF1KFAx6qjd4MUF6
hy4vJY/292R/HDhlCXDh2dzAQUZKS6jA/S87nlZE7bxhX1RzhJNoDHF5NrdeZ0Di4yltupaHT4sN
5ZcMEoBJysnU1w3Dlkf4cvdT6LWby+Mo5nNIg63Npbs7rinx4H+QfMy3zar53fXNLjkQVUP/Q12T
QAcJ2SgM445gKFE3OQCOByRyran13xYHXyWzEPO2o2o8SZSzalyiJwZo7B30B+QbR8KRl0u6yyzR
qN31xmE6+a4h0rg0r6w0rZJfDq1NdWL50RUAj0q6dWhMrdV9iM8YOt5GDpp1IA4ycmWmJpg4gzdU
W0nm6sRxoZgJih0JYfl7irBNwUrrwuy7FwNSVcwQQrr38P7jdyvklQIuabuRMS8N6MGDg/kxATYT
nkyYXsV3OhUawdlrFfWLJr9kKUnlMfLjwrrgNn38WI0BnHvmO8/mayFbfTGyfsKS/NV8V/LuKb2M
3YfxRJsDSPXe4KqbBRPUvxswPK8WSfWUCi7jfYx8AOTqKq8SV18846R5C+kFFVeueNiRxIDTRBH8
f3qI7ALJmcMAE6ci4PR989AJ7OzxrmK0i06h6R/3/SVm7BmyKuRj2lLtvooayzJYfsKUY+XPFNcv
fKkWG0Vbyg6TiaQbSGj7szMSgcmhMpoOACLMcyaU5YeelxtE8QIysF4hAM4PFa6aSo738waU9kx2
yKjmdKb280x8kzwbAg7t9otzz6rNCfCKpKwtl7AITHDwA4Db1pAZzXRlXunxp4meuz14MD+r25al
97jcH0L9gN4JhTGkimemoXNkde9JWZhKtBAhyYZ+fYC2bnhXBj517z0oLg0//FoF9MQmyGeRRrRj
03m2mDLgNkICnvAN9tvzJR2AZDf40mjhqzuavLGrveE1Kst7cN356GIxXrLnVuuNExba/l9IAyQz
UBxh9ozZDxOkGSJaKsVrMh7jLNMHTo/FxpLxRsT/BvfWMKaPiBTXEaj/j2fX2grPjYZrseFJkvQW
Q+1MMoOWbKR+eBSd2m1qOMQhtDcZ61/m3Uv7+emu59syLnVHTPQYuMhwUFebwvCigrnymB4JOC0S
bX4dHI1tCDbCX+R/AAgWCQS4SUzs05PuJDGQ/iQPa1PFkdKJvsa25c5LqnJAdkxIszgKcn4jE30d
twKvTOnVGbVRKzyfOm80bQhG3qQgYhanMWlCDARweL/KdTlgHr0lyEyJd+/Bc8tsHHKGFwF3aadu
kcP7S5OA3TMkeb2A20LghyaOJoDLocM+nZSH/hVWdOU/xlivyAp+Uu1+BLZxVJRWfruJshRbJigB
ZdSk7B7jgCUBrqcYVKtO5JQ1lDeGqzaf2wCTE9X6C+Q9qboTEDC6gqKQh/US6L97xB/4t2yxzGKN
kereAGsRuEe5mT9N5iNdbRVDNlJ47P3xQ4r1QBusWrPce34KHzK4LfPFj42cjzYfGrKIjqS0CgKO
9KVpNz/vxZFhnwQ7swQO/ishKMEvclAXtBnGOeNFNBZ0rYoXXCt9Iy10sy5eT8wXHErKPws3mF8Z
DyOm8uHmEyT9l6W0yIvgqWhv2d+Wk6nsT5enWKs2JQgRM2hukpZItGRAmdLYE1Hm3b6TffK4lUiO
lGSdBUwLo47o/WPR6nhcpuoDFLvVORcu4/Q9Ql3jIP6ZDSsJ2Yq80Rj9uAhdDkhyT2m/uK3IxDT/
dpd9DursACFZXEooecS71JcH1Ey9tTMH/kTfZhAWw866pepCjf6v0XQhK39DhvCnEcER0I7aOov/
WUaND1c+tqFZEuPGinuoF/ZNb1L2hbKRQCx5sPaAjgkx0c/7FavBoyRkupFynY6jwXQCDtTQBhbj
GzmI59gpcadyv/04lg8yZXiTqorvnKfHqX5+TiO746Gbv2PgkoLM6yt8QdQEpzInNuFyopkRPWpI
YapKhddinbYYUw+52SDoL+Z7TOgkI85n33xJIf5QD8YCJVJeXAXLzRAB0ck97iOiAlTQaXkOh8gj
LrOAF2QAo1FBMJNYhWS1suj4QZAGXLjKpDnYaufWRMieLrwxNgPyx9jKup64riWjOENPVIEIFiFf
rC9nvzfzrwnxtifPbUx3l8nLqyDnHqrcROPmDAzVk2ZW9Z5KbupIyhtAJz6TObQWMT0XZizGsNlE
v4AkmzPlSNZZz6/ff7vGMZZzp5zIXnV6e7L/HuP9BNGDGdscaIY1jaJGz3x4W/bLG4QqT3/TTJwa
6f9UAlaHaoIqUjcCVxPBKrsrDI6UxkOohBS9WOhWyldNroneP2bQpGdR3PHRt7bRCv9J+kvJJqKa
GBTdCb4akqkxk3gTnwWNzD3B4+PIcSo7rwhv5uAAkDIlFWJNdcAqFJ3U+BRjQl9/P6SyrpsVAuZb
aLyf3A42IiERw5RgeJyZj9K2YuG00Yflba8KDTunysKDK7YG1TCHh+ynyr70kBVcJr1u6uSF8jJ5
WOHXt5vjP5S+dz2qJw923xycdupfpiDK3ZMF+Rv5ok+XbSuS6l5e0Xo92Ag/n3gX30Ha6jDNQYpF
rAASjWBaNkIQwn+t7s/IQtoo6k/KTtgSMKGEXNEMXbYr5XLtSJYe63LrgNxvPLHgdaD1q9sc2s5w
JRAuhktOJ2Wevceq24hCr+PjshKa9MZDDvOOz9iW9gaO3+gUHTV4POYgsqh6SJTOv5DCaLVJLM+C
7+4PqbYz/LPa/0BSZuG9uMDzO0ZMo/S3kB0FK9Neiu+T3wsp6fs6qyi13AigMsWSC5K5bNnVlMHz
ZdfhZ/iQG1xrpTogwhVgecPFczDtP+cDisXfjiqmfPUQn9wdqWD4ZucnwdOYZw6SYK6Pr2patjVV
mn7LZ+mU+lasdqqmkomftFhL7McLNlyqyXqX2d7QWfppraddRZYX/06jry80kGisg5MOE0zo0g8T
LZVrxO8eOS8a7axTzz2/oa4ab5Jh2ZYzZiJBQ67hzZ68BDWgUzKxJCIy+gapt2TYBvxZjVWpSlpF
gFp6PnKIxqY5oFO2Sv1UDKzdBwLqJwQ2qrImjMZ5etXjkrAWCVL5Wtnc6I+SwiVVoEO6E/xEyUrK
nBcBNOJzbiePA1w80foySRF5rwqUqAzbK65/Yziupd+N8ByDBUfL8FTPY89D1BvY2w6wYmH6nWA/
Gfry58Ay1++EbGIqnDB0gpcCVssr4Pa2U9iChcK6yYeGM1XCn3cRBtfxpQ/KTW0tEzBLRISmU8gq
z2ae86C88Vp1Zujc3l051v/36TipmpO7gf7fWgkl6zCKEwamECqr2yJgRcCMee0jirQ3h7IVVYSy
F/EaoKnE2V8VLNpqcn6ChcmViQOFqxx3+YHVSCQYme2XyuWRO6enSMneKrAm94Vl7sdheXFEU341
hEli0YilZtF8gX8f4LW1e5gDYG+O+PJMNo1mug40DrN2z1+d+OfTT9DXnLrox+AEaammzB56YOOo
p1K3dseBttTNpEPjunV8GWh1bpUqviEv77l2joHFDWRg0BPqwpZDtazUJaCPZdEnneCrUsM3lExg
vREsZJMMWBSSgJ4/m2p7X849r3qUnh2Myqz/KLZapRynpNWxHfos4eNmUAYq16v/s0gj2emR5Wtn
rhnQ1pKOOnJPDviP0/TvLZdVBOSTzyjwP1F1A2RPtTyin1Zgf9fxwibi2ytpEaMx1lV/ntX9CodN
xHHVb3aw2Y3twhULwlZr94vzUDn0tmCsc17wSr3K1k4pkqfk1Kk6Y9CI9Fx7OWop6f68l4NP1Yqh
G72kY5Oc5GG4tyUqhzTsl6jH4fQ9wge6C66wAiFj9WguLyZ4Rj4E/+HI6HbSXnVyn6c4AZ9e3NuZ
ikJCK856Ny41mhI2X7RA1M3geovpkhalwSFk35RDvjjxMfRu35JiIQdTGA1MX18SgzAbvRhbg37y
iS03QhzocOKBIqQp+7gnHxi05gjQ8/CfU1eKqimpGYAAA/4B3pZweXruPycJNPd5wytWYscC5+6E
Rmmd6sRGqlG0NSzIQeZx3/e512+wvIXwyuniVuFa+BLUzQM5TfKUhxTGb/cbGQpHQURmfL6B7X1w
hDKLyBMTgc4FmXvZAY1eIwextYmNRu0sgNWX0eSMqcHd2xGxAlQ3CGEGpW5QvMZQN6eZhxc2B968
0e8E59LJVH17gdccpxh4a6AuZ52lRErjLKI52a31Q5x6EArZDPzxR3AQFNwCfH3jgOm80iDudqBk
ry5W5/FEqMsFBNTKv3m4DaUzIVDLUszTIilPCZjoXERrtywGjxcOVMyi7b8BGF1ZoQ87lvjUaVH2
sQPupvcGiVfoFWp8czRg4ByIBRgs2HD3OJqyZ8vZKc1Gxhh0DaYPlRNCqGGb04Bjkk+mRvJeHUfm
NG2PwHT/FZl1d4oMB4bbP3N2nlNTvDjZW5Y/yKMbaNWLDHNtenjH6jYpUbXLNAY4041xCiW6k+Sv
eFyZYSR4+xJWb2Fww17l3Aku0NJ+wmkxE3rNH06jOsrp3oEXJW1npBW9ubW8g6S1x2PpSYF4y33R
vfE71OR0kWZc0GQQQarD8SLg//zW3XUatYXTA5XBw5elGjaBwyx3BrlwoGzdE8pfIRmCHstdQx3u
Xf3GShYK85p/yBvkRH9WAaq08OHxUjVLjoWc0onvoKV4m0+/MQmVJ/52JO/ISepha3dy5On7ezCX
1tGMud1prJNaHLRK7uhBrE6xVnrgUSTUBmRyxZTZx5MjEJOt6sISHS7qbKho9MaP9TvNWViAoMTC
A9ReVQxGAUsu5vi4U73AixvVlSpb95bPc86ceIr7ojsIyDtfeBZ1hFfPwTNDXX/h38Y7Z6v1lAEO
r7qFWjLQke2ortzFElVd5yV01sy+sTodd0hirczP5F+VkF4XdYuX0CJ4hauOFFsHYb0TuBwI+OdQ
qNtXMgdhn0xCXBUKX1VK9sjMbVOrfLjAXbee4OqXIFiie8MrigZc0Ku9vOkZd5aZKsqkIa7nLssx
k8Crl2f607/IGyCzN+1A2rgE3N+8vA0YZl5JLHfqNIUfhyIdzURupuhZ2B67bhwtZp0zNvko8R0N
CgsNo/fgPgr5avfi7FN7vgIe0EcLIzT4Va3ilQFfXeXoBd1Q1o44FC3dvwjCUzaew9p8axtU0ksD
kzWKkbViC90C0+/mPRggsefxVbpVUHz7LcWDI8S06nvIX7f995Z9OkfNI4eccDfb7Z8/PVCPXUyv
JmDGW+Bdn9Kz8EGg7HbNJn2+l1kK4j/wz0bAg/ja7Ca86Jvmmtk0RdaFDSY3Q6jvjsFf9sNk9kn7
ylGWoYSybDDm+vI7ST1UTYl/2Ra3b8xuioiotxr4giVhMhqPUjQkWS26p7h5ZNzUDRyWpkJQeFLd
WsdHuNTmdYqNYQ46crm7Ttj0Ah8p8XDN6nogH9CVlrvgMY4ipIK8Qh+6bW6WpYDMM1Vh4bXEUCvb
AroMFK3Btagr+VEUr6a27hj39Wze58oFoZJhHLsIldqs2PPygXlx6V9orwX6W6yPV7stsQUhlKA8
hm1f7ITnzlABCnGKuGb8peMg2tfdXNBFppgWLfR+3LjVTlvk+aKDSneb6/IPt+UTN8R9lKc7T/qT
Syg9/L4enxlkoNXnBJDsT93DzqlKoFZ8Bu2xy7YsnDPSsoQcpz0NRI/orx8Y2W7tGsTaM/OGz8q8
jLGQablFjic/XRmu1ezxBjAFsFfoCS1e8FaAwPfCqm00co2C3SxIsp6DocC6VJDTdScp6OEO8LdN
Kcx22rS+pXL5J8DtvV3FhZUrJrrzRpMwpp1iz8vc0EsLXi1s2RlUfJvg9gRhBvLoZcfBMuFmOcvq
mF/M8iLmT/zAJvQnYyDpQU5AVc0Cm4yCrkmAIAcw04jnIGWTkjXQgZ/arnhgvF/0pkVH4Re+DP/O
ihpgAnxMW2qPr2LFmq6PfakhpkukoDUuT8wrw94A7uoS73WDXwTPsPQSQUkl09MDqBtar7mN3Ap8
pRF+jsYxtRooA0xKmhOQAk7DJ0RPl35nPIyx9RNVIuQkt/wDJq18tNrSbTaIeFzxIaQ09VRd4ayh
xMp0+vtslL41EZ6k6FijnJdqtdfgDjLpxOHEgZkJdvtqf9syhZ6l2KbwIsy5Pn++ag1ygH43Wpww
jRUP/6nk1jF7rnNIvI+syvTE3ofebXeDJucmLq8dNJG+AsrK7rQFWLmQeWSNx5lwu6u/axglz0aT
+LKzXUhntIQ6FKFkPivjszPw8vWr8qFN5FatGfs8VUj6AblxyYCWKNgenh2oAoGaqBoO3ZSMwOyM
9FqFwnV7zoruSGXnZqdP+qVH0xZourfHgTPCuKzeD6I0DQgH+OV0vk2jqyyXq9GeyCKEVDMPnB3d
BxgTGrCElOZGKJ8dRcVhSHy9kgosHNz8JGjGn8tAN273q4p6rJmnmJCupq6Gi9dIa3JNe1jNFvJO
FCxDMc0JBiVYSjUwct0opyYc0y3QWBqJtGFyGWFtMOeE3I7q/PzIc+S/9YWyGE23eUGDscvemez8
nQG6eQidehgjMm2vtSQoprpBmAabYFwH4kRfhX5tnrx5+FIu0u4RPUSdMsDQO933rJ8zzaTNcg5a
1GRMRI8mlpv13Y2YWsxKWNL6Uk2T12fwFKYYDE/hy1Np/la3c/B+EMlaf0z/VMabLue9+2r2/Jls
bgQWmLU5+1Pw5xyZexsIJ4Ik5L1V5Ia4wvRdSJxh4Z9lHaDOjcNhEqwMtYTdpfruUxjK+TD14v8F
OjlQ1eyQhxeNoD3bQCKFzb4kPCdg963XOmiRIOFnSxtimLTlrotmbJvG6qYMHpinrdFX2p1NuU/M
6dpPhgpVuPHSAAaD/Os4wxFBThFpqWTTAxn/V9E2/BTpu3zOkRIrXqbsnZ3yWtMRDcMNHlPxFZgU
uP68G/ZFsVfB/b7GK6XRzcH+4qraTE0/0K4OR6I69oKMOMS+HGuG4WAZGzA09k8adZFN4dISTVgx
z0vd1mP8YMS80nVFlsALEo8jM5crJR9r7p6zCJqZXAztOkfum6i07xKkLE0oukScQ8IK+jEgGfqD
unZgnwKh+25KjXtoqbQMf3qyQ+zLtpLioCvC/RXgIDBQ85dODOvH+sA13XHNU2ajI7c456D/oifI
LXwlnU4Mv46NM1ctjpFfKhXJegMbAiyMJ+8DRm0wsduy5KV3qPO0UF9402XGMiPML0kGbuZVnZWQ
wtltHGXMdTCercc8f96ALCJH3W2l/wfNIYA1ENCXkfmrotyTZWCDAZktCqlhMpCeRw5TcMe98NTD
JFoWZO3VipPAONwQkYPfNqNg1YEmLDQjLumLS5pKPdh63zwj3BJCFlwRI4NM/2VrUcEUAKLAJv9C
lSIK5tQllzJBLk9M0XV225eeO+Fy0N39YwpnhQbMenLR6r1Jp89I0BP+VyyqCILTL0oxL6ZVvdgp
tHGH9orIvmc/+vyX2+bVZwWM2R4VzesFwkrWgaILlhlDpddlwBThnqjig48gUUxg8q9VTie+FBtT
o1RNLCLsjRB3tMWuz71Q2WyjaZRzqEzgyoUTKx5egWkISIlygtCHfLOk3kB7NJVxkUL2m4vKFobE
dtzLjmY3wG7kS0yW6Z5qhItv3MDZEKA/iUXVROwFtv/vwCYcwfpQKy/serak4c94NP4dgnluqwmC
nUdYw8ES5xWe4qBPFKubEx7I8CKns8CFYwQsZuV1sbtEkLkrEJ7lWSN3KLS7hK8NQAp+n9OWzT7o
JN65zyvVMGN2xIgFWOHU6MplowrSCIiOtuB0g13J9OJJNTVznc/MAbLKzMlk385zcFMGPaLJY7KZ
Or/OLuwKNhMF8bpcb4A23v4IfySPIWYIW0wTAh5mTkntPjglqTG3c21NLfbbjMEXQQB+Qz0T2or2
1zblmHrqpch1sUGkDnwzQJVjFxVkG0drVxLZxaeLcqoz4KRnaNFCsO8JRVG1ZPIjFAB+wH955iqz
YihKfLd3Mug+7fiGGHjtzrxMJcpwk9UfTlpPrscgQ3FWj/4EUByPHlZWP4RnbFCZMhyyLTrDhbhj
uLwWX3ruq3xh9RpE4U+ewA2ZJtb3oRVrCUCGd5WOk2sv19us01SOYllnQiC/97i1TVAI4Ooo/MPN
xiP5RUSrKyDM7o1yBjuPuqIE/ewiqQ5ufSR/MugOYwM9xEBeJjgS13cjaI/MliqzOJqWjCS8JsNd
QjSljZ7uwFic4GRJ2uoWIi5LqNQFoOgBNO+Au9tz6fCAr3X5yTheUJQ6vRQnUM4y7vKZin9d/zS8
NO5Od8S9YwYbXTWCbGVXG5yO/a0cRzQTp7derwuDba/FZsTMUCXaoX6OriEZWAM1RyNPyPt6MsUn
YotJIX1H5bL9zL/xGSSrUX4AR3Dy3/ygBRNwg/UKrH3NNYpl+m4J8OawoUXvAmca4kyzwKyUYxcb
5k77WQcYFMlB29XimXf5UVGH9nIDZ0YTuGKLd/GFiEx0qBUrYbrpmkc/TiOFKAgMm2+jJfSdcHbb
e9UOHZ5QkJnaA8YXijLPlIKE4lbdXfnoz68DpFOMf8dRmey4qtdq0yyft4znsvp2EB+sK3xVlpGZ
2f5LDwwI0R1QpKoMWjRz04MmPdY58fMO9GKxC8/xsBB92HfzHQD3EDRwCQq2dpf7KAzW/RkpbMfD
vzU6HE9baW7z7KJCb44UTCrsiKQtvjsyCfak8bTSLeKenUOuUsVOTv7ygBh62O6d5knE1ah07F0j
eYrcEHDIsmqvUTbnx2K0vizFOJxgSiMMSgG8vp409Mo/n2RLCQ67L7AZVKbIIPJnHk3Ezi4yqFlr
zfO0EAZzS3OH7f2h1kAq0qEtOaP6GBjTE4KtTrfnpfk01UqD8xfzEdpcJoxUfy9WffdR9B9e+qRH
WXzFoa49camwu7VJPv8Opdvj400E/GNyNRHZxnRqh1M6tyhJ+1Y4jRi4rUryyMENF8fhjfbJvtSR
9x6ZmMA8skkUtGNoatUWHD48LIhdF5KV+dqhzdAYqeNC5rHbWlT4uxz/0FSe+5thq0s8KhpRSNc2
NP02Eztq5s1+vhetkgzj2QNE/TSxag2yFlJTjM8IBD4Ji0C3TX2vWvuvUBY45LY62D6WiNmZQFAS
O1bwZna6mQGX/QyjSYXp9iFp7kPx7+1P5P6L5offlEEMwo+JYJym5PePrmXZJ+4QpUlVkJGzOkly
DopSyEYyEbH0bwbdtg9Gm6lNZEjLRILZFu38OE/RDSqi99is/7E92ZsIqWkXACU+lYtHTw4UCJCW
PVHAzUi9ph3n6jSmCI7QNTzFNvONwwOgTMyNcS3l6O2szGQcJrhNxaVdnu0jT8/lYl9mynUsalNd
xZ9GfYoB+x5tMGgFxywVRJiec1bZ52Ruh5uoWF7ijo3uzC68PENP42Az1RNjke8pKzY4i9EdDN9E
c1XRy4mv1zrlSnf1ozTHswyaxWX/6RGqTgOzP7KVwg37w0csAXzbW9jnGmNPSxpx6DHHnUkidd09
h9oJxO0DmbaRQPNrnwpK7+lfsIOE4ytKV3K7DuK00eSzMrpHqYcQ+cbgPdV4yCASDIlid1/QTxau
8Zly1SYpkCWej7kVdp7Vv5e1yxEVflQfp2oWsNZEyUhCFrYsKoahCMaPQ1WBKMbKVORapCGP7Jdw
jFc4TekbOdEBSWi/rzzeBr6jJEvm6KBeXGpTUaLK/DL/QFnngNvGSB1QLApSwtleFVWYla20gjbU
h5imQmYy7RCOo7PD5E/rfcp+M1rJogb7sqqz53joD5CbTyxkx0OttTlH39DlaQ/c/XMTZj8oq5UK
9m33HLTVWzKV4/IQ1C5nN5yczJJIAsMVWvFQ2qKByW2gofmS1VI51EsecYwm5VKXtdMtMAB0+PGU
+C1E3kOQItmpsecqTj7Vq6d4bOT9MjSAl6PrTOZ2eY4QgE9WJklERyZW0dhDqE4s14sYZJ0Cs+5g
CxEfJYE54SdxJiOwUS9uMMqwDoKE2mxHUYBcth51cNjzWSxw/q3EQNKPWyQDAYGNSDtK0CjedIqD
YK210jozJ6XD9GtsvP/RI0TU0+LkgglLeeBQHNmHJIIpPwtKYGnQPi300/qeUITkbzpcFn1lV3ur
O+lLwz+a9HVYlcxRnbp5pqs2vHopZb9hxq/ZjoxJi8gYGBg1lnHaCRA/9I4WVAJpQJ6zm2+lR61l
zFpaMtQ7U7MhY/S3+br8a4g1UURMpUwSesPeXb1XI9N9F7JAHGFY155Z3fcujXxzWymxMdNTw8Sh
Nwtbc6rpsr+lO9vKw9QppzI4TSxaCpl7DoNeqTzzHKmhabDq1n36jJAcjpepgM1sizTTFifUwI0A
kXZxwd3PBNVKdoJrWlt6VaghZHrtkECrElkqWNWjx2P51kgvXx5lvujCDieNCM1miJP+cl7znrpj
FOmI6Ia65GKPI1UowIv0i8ASaMWO7XmwwVyzVrD59Yof2sO6RWfAKBqrPANXw9Hsfx3T2tyXHfJq
Y6hapIOUoG4Y0gMpgKe0DqpERSgDCHbtEZC1vabwn4S61V/uLYbFKt6mQBiYIo51e9q7rjWzS3J0
6LcBAG4dsrSWjf5iWYlnrlceeCjicW8xlxAoatho6no+evAoH1rB/RTCJ2Q29rU57IQp8CUVD4YQ
qfSA2Wpb+E57WJo8+sXNxZNahN9PfE0GsaBlAQ9bH6hGrlrfH4wUAfZ1335TZpEOhbD38+nk9qs3
ta3gV6KFWEhKP24urWUd1tI3XozEixLzSvlG07gMFQ0sX3dNtjodqyzV6kw/A1nK5pTEUxL3Gll9
Uuef7K7yh1crp+QmKHP4kv7Z1n58ZU7cPLmrXA4eMpbbNgB50xBZ8+H3Wyl3/p7HT1YzPKzl7WdP
6wdjX0Ho4r62x20QsVobek+PNVgMeZco+uthfr13T4AW5/v/QYN9qYBS4WktMCMxU1XKtNmaKq5v
SqVEFIPxJbfJOv4kii6w9JNqu5352M3rSKGe4vap0dKkgifRlXTaD8+OJuAXagOUf1Hb/aY21EcM
gqye7FU4zya5oeQVTWCRhvw5o20zO0rni4wj8MGDTrCLSGKQVNQKYg+pGtOaX178PCoVLeh6a85V
7zKOPSBMg8YPiOy1A8FGh9S2fnKhmnLXElBBIm4TF2DPjrWs+XxW07CsS1YR+6Ujlfd3FrE2wOUk
JQ84PAYzD3Qn56D24atMXdrTedNGZAl+lxURodXa38KXeo4EGhuVs+6HD4GnYlpAMWGVws40TsMt
8R+FzPAzHJu2LqAYAN9R4PUPKQVKPMW3NAXyDDZ7/B9kNM+6yAd+GY24zmOMDtPv4WZ9OdVLz5KT
ULFsp6IQKZV0uHZycsDIv5gWNCiN07mh0uk5FR39WuD90KMvKmuHzLjkg4KFeLLPan52WNmIsN4e
D6Ir4nRni6i/Po7POYMa8toPKXI7p1wPSyTNDNt/d7FsWJHmZA9Vcgko2O1BisbgUKjP68wsgqHT
cY06CO4iwc+5NUXJbdibDRReJrXnHPmjlQD/SEXWvujU/CYM5yBOQ7To4r7Q83pVhlf48TYoRZHL
keRbgN65DN9K0XkZ2VnQhQrWmPSk8gvrQTVktfaEKRCo6zdDmwlAvll1K0kaboU1xsvWeuDZVKcx
oBmcPtyBG3ASx8c85lyS5FKQ5EFUiqAWKA2x3U9x1JYYXZUazBdLFfjXf4jP8PyqvkT/6hYBZ4BB
j2wetPradVPauOyX1AYiEDnmP/eh7jvexxseCAuhvbSnTEZk7k9nQcBfKiUncp8t6Z4CntJ5cHje
9e6684sd1kG2CozWlD5Z/R4aQw1NF6ARKt4xV6W1VfKeSP1sJEfxkQfSdVFz6CO1r/rawj0dmZn8
q4j4Jkq7B5wLipuQz514sOH6HtQDFI5EC1ReSuBdJmpHZeuJCcJUrVC8go8Owii0yAY+RCwrgAT6
3+38YDXGYj71H2LfvTwC+IaKiu1QBTMMo4KdENcq314cbRBetOYza13oE5mw6y+ZLd0xL2JDPzt0
lmKn8UTUZQ3SvOM0Hgpp85UR5jkN2ZjR1drCa+oUtHNpsni28iEHiXDmTeSx/S/p2VlL7oBlqY44
A21R26t8MYCfXoM8ULUu9PB/ejpTK1XEOM1Ipw42sU7UPaSfTnalxP23EsCWD1zPIlKGq9cNK7PX
IQ1ppTM46vBCH912DJRF5tULHiFrRbC5yO7xDv+7231imFtSF18imJLnsLSoH6gDY5BJRTiQVsyc
NILUPwJJGl3+ehbSGIU3HVXbdG18rtCiKW4eUoN4NyTu24UKJ2r+4t6lRQIYcRB73giLwvZUoMkD
GGpckygnEmE+rEwVgBh2qv8XxZQqhL54RKiIRb/Ki8TFu8iLak+K7h7iWTlQskWnmd5yAH/8MLNh
QzJLkRODYwE2VdSEO4WHRaMP5heHgAMKoXtK/K0CAk0hhwtL94CtwgmYLlPJikM/jZffb3WzcWkT
u5l2IWKTkE7aQeDLV5A434bQmjns3yLVX9wFSJ/S9LLjry6u/75SzEv9Snu5FK9SxWwUKDlOAQu8
n9s3R85/8QhygS55DP9OiCzEGfwiPbFeX2gDVKdjwRdHkKEkISfCDtuQ8v0z/GoFSekqbo8cm0gJ
+IwU/rkAl/aazyZWm4GE+QEIwTS79Zfnvv6Megth5zRKDduc6tfKmjHV3YDLQjDhr7MxzWKMFjXm
ZIkNo8N/mprBxuY5MLCxA0JjKw8VYWZos68I0Uy9wnRRmdV4hxouTZVNENtSLBUjYk8ZMOx6LgBG
qW8SjHzn7LEmoRaWjJeWRDnwdq9gzc7F1xsw5hRZgJWWT060hwoP204HdUT1tU2phxQn0aDNck0e
uypvCPe5RoGPkWO9z5wkAeUBqOalVv0kzkwBSjpSFaVaxU6H1T6MLKv3W6Oqyc5PQYwsZQREToyx
uq72baQqTDz87UjG0tdYB7nte7fPvtZhBK+XIOTdi869qqCUkj0ZDVuhNQBU+0amBOjyDJJZKFW3
xt2VWoYh+rSB6DHOHUHcrKD0H9hURv71fD9Cc340ZR5v/RGhyJZIUCUEcSwUq4UtazZniSsnk0M1
PUGuq7mSVdKkPX/+tG/DHZaSf7TurAtd1nVW97jZ7H5mubF8tIyUqbkFxpjX5Vx8RL/o3GE/yfAZ
ywmbD4/tv65nkQhlCw9fs7eUCdLXljfMMVuwgHliN/rOSfkdRdTavVmPE6l6/rQ6xl7lH8Wc0Ck4
4SquYzXfhUQUupsN35BqzG5zl70hVNwJjj/1eHFBiIe7JjEcuSGRS7aNJZK7MJnsjz5LufmVVjAM
VhvIMfqwuQjx5mw1unUF6mQmU2+fewEqkvYtLouoVy87rCxthLtXm34dEAaJBscYc8nf/SnLqr9B
PY4ZFIyss61BzDP3cAreMUsvMnpek5h9sh4mHz3O6VNbD4qoR3cmyNuXRQI7yilzewlY4LcmpgEw
wbGRnWWsliWx3dehlEe5BVa6TZsjTfUQ5mPpi+L7S/0V0S/qHmhqPxcoIiZawJ0CReJl8RWYdWSx
22ypkmUrAR+KuZYSOb0ieQEzD/oYuR5EQ2Euj4JZlcZ5vUtmUatDiNv9tzYAmStEpr3iZ9diFBDY
SIrp6/aOlMolEETf1zcUNcBNsoMy8QX/nwB9iGGVjkT79Id60ZwJoEfwk4JVjl4qOeHEhsGAyw81
623k2yTJntGvti82KGBNZ6E0bna7Zpj3JLM7zE+6dlwzZDwVJ/ZW6UDsHXput9DxP8hkc+Gn7GvT
eguH8yBF1V+KSxQ+uHfE5BFLnFTBEiWtk7ScgS9btmB32z5D0ros4FqDjQjcanaOxuvozIOn0jQg
1vKqAFq5ApDDtuxeWkkQnoqhhGTAqa0/LZRapc20UQLgKhAzr6Ik0jeEMNzRdAtU4AJ5rF0dXuB+
R9jCvgUHManx/asBfdCYFlzcf4tryrtxI0gdx20T9CJBQLUqduEge6yq0C17j0ZU6RKkf7P2KR6g
6eEljTXTJ+8DSKxowV30RUaKTEfeAKlcX4G7xUR0wlDKet6ogGx0tfjEl7O3apydlSh4ihxb6/u2
hmvLIG3ypzSIkmygC3/wxxaR6ullPNLmb9d6g5bC5IHhdgILvN56/RsgcaZbENZZZTwTy102YPDd
o459zG/WWs3F+lb1fOO8KGhCGibjJeXvdWsn3Am5RBPdvNpbpHPPflyJi0mDGViV0sTh13Gm+YkH
ro+DGvoVP3MV0aSS+ynDFjx4rp662iMN0P7zFQnZS7Kj2Y1agvYvPb4tt1p6rvd2123FG5R6mJrA
NhTktKkyKfxQ6s08Pzgg5p3W7YxTgoYYitpLVDErj64ADzkr3un90Xe9GCPnF0tAn+pFtQ9pykkP
5q2Kyfgxg8Hw8TfA5BVKJidfAGohqq4RBNEiiStL16P7g7ZIUyyCDz+WkY8I3pbEpCkaOEIBROZz
oIaHGdUi9B3Z+YVbxttQqTjY92F/pAS4Mrg3OI9uPhvNYCTRoOi2xMEBOLGOZhqjLCd/t52Mm1pC
nhedioNPR7Jh9OQe4tjvD3Hkh/VizMwubsI/KxP55dvUIr8LJh2gW7FNFzJvOvySQjkqVtNgEoyl
EJ2ngGdOLfG/1rne5OXIwBUWj/sxaep1gmcmckbYGkIEtx+6HK69ddtU2ZRMAJf/XJGCjClcj4De
jzwPXCNQ72AcJs49iQuohV5LY0k9s1IKdO1HQejZGs7iC50CwZG8bzyRw3KQmdZZI51JhkzjZ6ug
SeqBaNWdkDq1eunZUTNZ5mH8g2mtesX4kA3aghRtuRXPHCBiIo7lyg3wgReKPGdJM0/jHBCCRFu7
NKonVT4UxztNht3iFRFbEM9GpDA517Ei7A9wipY046r8hs9IAJ/zzkUsU8LIVaTjVZPPA8Mkx1RH
OL5HAzm+R59VjtuifGKQPdG3KYMk8cY5WIsiBu7UKmkeVW60icOuGtNvGAYzbWAWU5CNv04cIOxH
qJmjSxLU17z2wRyW8c6Opytqm3Taf9FTUQIdRNdfQquxAvnlS0nqi1aTxXb7P4ybDs3er0q2LNNd
8L/okO8LwocH6rBE0d8r+eSf2WOGBiR8YU3iPtssa5VjZ5ie7fdGEC1Q3jbUzGjqalUmW3OONxz2
bIwiKcnUZ6eGDiZLLln/nJvs2WMXXXZ/8e57zXL1k/uCYl+6vWS263dq9c6jPNBrkXR0hhlhoNSp
yPqItijy2AFvlgjdNB5QoljBAv072MuxxINVLsqc7Y1d9HTmISaSdoygSOGqroS92lzr11+mj2AF
mQYFIFYM1HoB6t8ICpZiqzRwbcQ6L35jf1kzhGDObFoCxihhzhZvTmr09q0xyZ1UN5BinphA40Qw
was+ESneMmdhzs8ZCP+1vdIKZa9gyGfA4gycZAuHpZgkfkwRIrOAduYEiqMEhpJIZTRk3T5lbBA9
MrWQSe/ip/RbT9usW686IJMPKZeIVciRU3J6o6ePxf+4bVl1neLrlm4UUsWxdNJguV243NvthGgp
9NRTTF1xL5d9OB/Fil6QoNaNVs71rNMCdRlozwhTB65xNm5ntTNir1EeDG2Dn3Are2GUgX78g6ZU
Vu+s/BeWJJ9cb94NsaabT7m57s0dqziSLnNMLyOhNTzGILUXmTQEoj6mrD7nNjneydNlxewwZrK3
ngOGXG7pJqeOL5ma6I7wOAUKUK1NMf+KI2SnUGFKvloxjYl4PzcAQY3ZsidQpLgL7LYk9FEfy4QU
5mshbKPepar2H/wGaUTUstD4NPNPe83ogEXK8ALoFmfYt3lZC1hmDUYOzBDQCUlvlakxSlegmaER
TEy/2Pdf/TLGpz+GMrpgPp3X8S9gwPihKcG1e7gJHWPSZD9a+H4pJUnGe5+sfIEpr2nyj73JIj4s
uKMmy/9gtvTPUZzIbkKHedWEdXDU1jmy8Yx1jNPVQFMwMowiU511tuN9v9aAkvgzrqbK9dNxQ5AE
ALzPrWbRBYasdbSCJ8awfP/5oIbPG3269+mr/0TuxecBhjxAbzQF3wPQWZ1W4EJkg8TiVyRGItAF
ttiW8PURc5jXshj+dZtaCfuhJmk2AfWb4ra/R3SXa7XFuP15srZDk0RRuwlBc3e+0W2Z+7aV5ak/
XWamQ31elIdfZ/c/Fv8pEFMh/v4ZJ2ABJAA+Z8RdnUeJM9o5PEINEff1swKO1ymiACA0ABDYgXYZ
NAQu9nVZB7FarltXTL9eJInJc3qlBmSJWL9MhZchRdKfw3X+2ZOOg5knoyj7ZkmgLFqejOVFPYKS
iLE36PjG/83a+U4/I81Hm9ZLzn2495gnbSQieLecMV+O0FRIul2zIfSEHLLqu9BENt6v6fTe/Q99
cVYhOCa3KwCxyINi+/XpzEgCcJLozynPAeiigOiHRBFiFcDs4Qcot4uwCyV5RtK5QJqnIWBxPSb1
e6xFiiNHDZ9QZZ9I0DOGE70vMkCXDiBzUH7+Gw7fMueo9Zz4KvEbdocGQPC3A8ZpEMq9pqH64jIg
81YwWVxqU/ppNRpZEj7ldGB+SwLWhh6UyZtvVXvqlzV/khcW95M/RcdSPEp2SZo5vqs3bUtHXkOr
5kv2k/D8AwBEa7OO7QCLzqwjKRvGfBwBaOivfA050VadM/Trytyan8w+EY6NQotlT9hxiEx1YK/l
nSV7YpT6z11+KFSVd8Tc3x8QkWJEM+lzJFs9Akkdsek/o2d+R5lXyOcYvwtn5SQnKZRRJxEFH+Cn
inLtSXvuMeSumutBHkxTdpAIKJjQQPAcacYRf0SN2KzDMr6/CRCbNJHRzHfdmSz311FXxHCBRm+/
vG2IvFMDKsSZ4HG4JU3KMriT5aMkjnzZ476QQ61SrKr8vstBHDzKxRlVg9WmYKBxWLlQ8vYefrjE
DxQntqk9qa0ba2tUbqFGhcBHOPTdm2ayYVRxMb035qsJy9X7eR6bxLlGmk0BGStd4MvfjEU/UdHy
TxmH3lc5TrQwxrtwpbgqaHMP9fQ/6cKChV+KuBqjb7r6zjREwj9vYkldIc64BfQb3I1KQ2kitDOT
vj4A0wmH0Fx9y1sRZA3L+g3g0xC+WlYxL3xngKGLCKGOrtrW7KQ2FkfDd1mMp7i6EQ2y99A5d9oM
xmi7uouR0vX83AjJ0ieI7tKXi7pQay2Byzhqth2p4yOyM84a5YkCBq7NE/eRh2YWVirnDUe7iE3W
9yBl0zhUjL6Q7BDN8zOAGURhH10qOKvWg8HaNB/6aRZbnIoobok4eB0Qt78zUKX3HrZdWUtaOUtp
s/DE0PlFwdRq5t6Fd5/r8HsKY5T/TYp9MI7sTAIWVg20R/qId3d/a8pvvQC26D9iWLlTALrcbWPt
X45qs+tihed6uUtv0FbicRxH87NBnLmm7mYERmssnXXEoHr9MP2II4njNvF6uKZkzUnmlJUu+G2x
bJSvVzrwXFOk8mTPXxOFDpFlbij6UTyxK9AyCtvXXekhz0ICBr53TFABSu59tzfIVmmDH7l8SiZY
JgYw8EP4Y1VB/aZ5As+/8hhTrzT0H7b7RX11/3gN+NzJMbF03nuMXyPxvsEeE7n9dU/E51glMQwk
JNB2ppEWhTwGdBtzRvU3tNPsmaNhyJ+kEug9Oni3q3RQ14JgtYyUi2xhEOuCZa1s1hyU90KH07sS
H7gClzfyiBNmgagJVVl2Cw66WBHI+dQt+9bEVOfwYouSrzObhU02l9y2gfGfJbnTUVX5Rt2LZX69
1u0gRoemiPMcbsUF0h2bYf5xpRb+3rixMp6KQgES8p7iKQE0wi7JTEe3sbdZhw6RZkbAlU0V5Mid
zL8wIFOAmtUnivda28xuUNSHr0wIOn9a3MsWRBIWiaDrFWT0o/ZPl/7mMzbRpSDc5p48/vrrmStZ
eNVbKpSzEfnmy3xhCJq8Cza844rnvkCEKDvtluKE1jIAZWOOJQ2aDqRRoxY34EpR5qe6vgKwYAFp
8KbhdA97L3GSFFTnZK6ZBmyCs3UxzJFld1jDWSnWFgz/7m5cnbPCzeBxwtf+fwM6Tv/HBvHOxII1
LhqgjOTMj2H5cCqRqN1PBXHcFk5fzidPwfjn2wfF1jTjywrHy0KNYftswRA8z9H0Lu9yIjw74RSN
XF4J2ih2fufc+gOoEZ9AE5EX4LLzYUfVwKqKxFpNm/TAIV7z61Gnx7bivXa705Ra4IapzhizG9EO
yl1Z9DfuXa+lXtEb/4h0AJRQJCK9se3u8Mh6WzBAkTdC7Cf3HvprJwmgjOo8q8i44qJfkq6gpckI
FzfPUbTolP4bmcb3+lDHWcA5S03BOssyysljWj8SUMVjgNJoPyTjHgWdZIyqb2LH/0Uz2qMCI6qo
mB/wsYe80C1tEtrNixI6lK4l313jwFU3sWYtHCWUGyVb8Uzp/nDoPF3/RgQA0K2evMgj7NkxOjkm
RRrTMkVIpRp4oDl9lhc+fCUYSO5FOwaNvczBwfdusT0SsAh2rDTd8VKGbuFn8tC1h/2fE7+DuOSy
jyU+CSXV+ojwWJfAQoAwnn8k/YVzUBbtJM58yFnkh42q193n3kmfYr/c4T++1R8tUdRyfK5DZHDh
40/QhhUwm6VOQyMjg6XoEuGz69armjUHfhbgbKmc+P1Gmnsm9s/6phPD0wt/sxo38whA1fBju//r
pq7kaG7I7w4NhPQXwPuaU4DjBQX76QKcVrGVc0rwiRAf8DiLbiCeTqjXKBXYd3P6FPcxZndxQ3y3
diMsvDTea5msWVbuC5bpSUldURcN3fex7heQ3i9VVF/gLsK8j+Jhlp29PJB98kRpSn5s5wgNkf97
DHxz1rx8FsinM/PBYwAV+6rDn7oyaWB5C9wrtGMNWaXDG0FDQnSdeOrh92f2tKMYKQJvMr34rmnm
lly05yvkUrLu0lapGk8nJUKE4z8oaiqWJswqZqUtmvB5tAf9914BEOVFsAsIPxPPrsAQ0ygjBcEL
Nuyj8/1RbMyiP8Ok+hC1kwe78V06zusrn45v2pH2E76jMJoQ4Dca3c+ii8BhnAgvZZ8TCJXYnEMI
vr2wTaEjASR5SUAIQ69dvEbAWskSyPitznMRKWgOMIkjvpZAel+1dqqIwSQGb2hCazLgcu0lmmiU
2qSWoEksA/jIH/sCNGQJ4vg4TTJ6GFqBssindAUblduefSMZgF0zT88xCP0Crpg7co9zTSwKoClg
OoJ6lH2Pz+kwpyZYZkyvnX6QXVs2ZeS7zFihhHhmUzqXWoNWON96gn1+aEIqUkMWQd7wXvEkH9ym
QAO/iGCaZKGRhVN1hj9W7WPH8o1AnQkcIGpkt6lDgz4B0SSGPoczL/VDgr6Hga1hFgriuWBvYRWw
FIWKCdHr0yJSX7ai1qFSFCaFROI7AMXUnpMSjaHyHKuZg/2aq8iN0CNVhlbv64tDodqL5h1ykCG+
0x6s1cZC8KT4YoEqok1DFItBc2GZcZZoodDk3FjjTFIvJ+7WpFZFmzzAJ1AVfp+9C6pww7yUafRn
qdqJFap3EEYmznID3ON3sjurbUAw/peMXi9BlCa7qS6p9PXk0uOSamsUbBf2Cv55S/j07F+PA2bl
zD7UoqILbnt8JiicaA9Ei2OglRZ8G36e7bBm6qOhhi06EQB4NBFua8gzaYc66Lb69211cFmhcRSB
7r8FfP1iXom6IY2gGdpePIGYiGJ8Y4NQ3+Ao2gmv6DFgznWMppUiV20hYLeAeuN66fXeBnkjJ9VK
zRHSStUCN0v8hHwuEJTq3P6GXqj6+ySb3W9Z5bssZI5X2zkiIpNWTU2VnLda7GTdo9TnCk48swcY
U2uIEBVGiGhIlRsPgkwgwzK2CfpDtntlqmhMgl3jL5M76LDv1BeE9Dwv0asieHYeNCldE8NUcmqs
S6Vsjk6V3A7KxhUc3tD2op/karAgvVjFMDIB0qMBB0Rru0vfivegpx09dFbY0zRpLW9Z7f2O8hYR
OJDzAfZ9W6r9BjNJoXY6zdg6NP20plS65Z98optxWRHFWljX8Cn4kHd+A6sYZRmxSownlVFfBGwP
80M6sqpNerX7xKTvyTPd96wUlQ1Zx+/YqWoLKtdDcMyc2fMNP+LwYUsQYd9fKWlO+NBy8eYUnDHJ
KkuXGmYdEPFYu//0/fJN0AkE0PkN6ARd1Rr6gKaxM1wF+DeYJjb3TfYPY0OslRb0izzMQmbgZToA
Z3AUg1BxZInl3I7T1/BXmR5JTXqE9KK8t1smiaxjn6r/J1got4X8zs4KWnfvjxtNwlwRrwItBGDn
Loqzver811mFharItKoN24iTiOvXiWQs/bLkHbTayVL+UF8hQzXjtdsdGqrMy2wQeJ528kn5duqP
bJ/2jQXcshAhEhjqwMeUEbwkWFM+2R/Bj3KpELR6MWxNAGZUghEmfH7WHgc6VqBeHFtpczCJYsID
hRBRqaAZq2FlriGhgMray7Kd02gkAMPI7DdfK5wECvoI+q3mj/hhS1MxF20tiN4iE3QwAQeVsiMF
LlVanhXBEd5lVD1QhFnBC1+x7QolDt1YQ1GkU3VTk+vYGsxczrAhL42mAL4tOkzEuvnFu+PXmqxe
1Itpbpkf96MeP/pRSywiF5WIM0uLPOLxSWhJCoLoHYERFCQyZr1jNg8MKC6TeP0XE2jIat7WIhuB
23rzak8j8YCdj0t1TWBb02k5kDnEMLsU6AWfHYrwvVpTUsKJ7JGb5VqL76Y2i6uhJU464n0j6Q8H
lFJt9muK7J2P+SJDh3iRKXa6BDelA8uD1hc6LKpvX87V9fd/UmFLft/74FDXAwAIiNkPvgtQZj2X
hKADQgOWI0dB78FtzgQDo7410gIFNWPvsWHzQuUaE64AXx0LeXrs9nwMBRdJ8eGgTcYh4FAiRuan
F9vEvcO8mc9F6ZZPe5eMGlGUV2P8E+YiBLR5fC5S0+S9VjaXm2YH6AZD1F1D4a8N74NdHGptpXEI
jad6MX6DYo8EoxeE3jWTScMxxhh6b9CiWJ8ww1RYz3LF1VxTUbCAWuM3Zz3MFh5fLg1iGCJpjHPW
Ejwytl2jOWB5eTFL3x521hPCMzMCcGoa2VXNh3eeMY6aSlm43Vr7m6iMk4EXkayXlQVg7jr+leKe
t3+JeneZyqTALjBfEbdc1buY5HoUFIsGa+x0XJoTafLYAwnv91MI32sUrg0KrwcHAWU3HT7a7LLt
y89MfU+L0UTv5BULuPkupxfBlK0POBqu0tyuM166O5e7bLcdm59uY1w0+SA1EiFGmlX7UEpXN7t6
sZC1YmopIrbAiQGmQOs08mBc2N0Bm/LYaRF9s6PG1TV5bfaY/L1Ooo749KdBmDmHO1tX5OZfmhzt
2SNsaRRSqVEkBFcmx4iyUNoWzas+JmnYy82SwbyJxXnIhh9K6yJMbnn/cG6tky+1PEACNS2iKY35
N4pCGA/cL+VyS6XNIedF/3K617zgeIkO4txz2ET4I/rxb98i8yJLCa/MoeKodzYKR4ROyLh19f3D
V4wHAW6091AFAx3VjHwcp1XBDreDvMZ5So/2CV20t2PHo2v72L33ke9sZ7w843OV7rtwdec3+Kfj
E48MehJnnagnr8V/PHWg1X80P8xtonHYL93DUSkd7Bz79LOX9UL0VIfn5h/Da2JZj2FtTMxgiQRc
GflLsNh1moBhT94tg2iZlFN/eqRD2AyDH806fX1JsQtVzqBeIcQhqpjxzblNvzOcCLeGEz0d2B15
CFRJUDPhitpNJMyUZCkvgH/QW8EfmSt/+rL6TDbGMrTNa6co3BAa2KzpaHe5cQuWsMCwXs/vMA12
1dwb/V0gLIvuNDxgDyNteNkquGLCC4J1tOYT/33RWM8lb6avDBILhAspqHjtBnViFDoG7uQZcQMB
3QpuIp4RokwsaJmcTUx04Ggg/FpNRCbcDgWaeodCCdgy3BKGFS/lkKpw2JW0kVzi13Ebm2gQEtNH
PWYqiaS7L2bkN0epOGJ+OAI3YEP0DoGFdmonjQ+VfJZUzTIDkL/CUHOY7h/yISxC6MPxGeXcVgt3
vPW0kkPQzWU/EkL85qU6+ypldAmN1rMlUrPzck+rfb3lZAk/uz77gl0CtxLFo9o86JkUHPau3T6d
3jP9BjwCX3eBfa8ZlbNEsaPCC4I29QIl2OB+ztj1KpGPxKzJfsKHNy4kDE5kvWWUabhLoKbfJiVt
6GOyewWL5DHV75PMN9DxYDCFPCvFkBLlHULEruAGZYbluv0G11wEa46D8rKH9OE5h3RT3qIioknk
cfECVIiTWDAzT7fuJIDvOBZfcKjXq0rsttE6xhxsDd5Mau6wSSgD9NJJrjukt5nv+q5at033bC5v
i1a9Lb/tWh6JOd2SJkxUoe3b02p9va5Ic3oytF8je+AsWjdiuCxv/SxgiOOdq7qnr2e6kZ16MzBF
IQaXLFKkjzk0bAqggDhUDjJlQWIhdoTiPR009FMZvWHCK59I1E17YZ4Yl6oPHqwHhgOx5azBWV2s
GPUqepszdEPnbyb+BUya4nHBDzAallipkO+FMZV72mkSfZ9lPshqr23jt5ihgNAr2z3/pjHAv7Fd
FNFQxFns5K6dzWcDeMedMwsRANCfmZdj6Xu2i3I/OtJ5WxZ8heGMO3xFimn3OOoPB/ZnpGbXKdC6
o7djzqWcFck5W6pPrbu5Yg5GHzPPT3rWq3wDQR7L8VDtPeCfu1z6d97uT3YE2IDZ8lle1glDEqSf
aAlIIg/yfg1aiFw2GXQ6wEE1fWM02IbDF8bE3akofUf2Dt3p3ObaZMhdimjoH2l2N7nksuNp+ZGM
VGPTceBgUYRhUXhhElVJS80GnAidyCezToFdi9Q+tX6VuPQFB5l00yl0YQwhQtq0ueCfzl+UvJ4Q
LvXWRizQWZl7jPsa559sZy2teI7pq77elZadURZqXXOdr/xXOmF2Y5XJrtdZAt4kE99ap5WA/FB3
zUW4hWimYDrTrbIG851iD33sxUQOOkM3gmMGm68OM9vs5yc2S/cfNeG8lKzgX+9ZkQfnNUAXc9u0
ip/Dhf7ZIknTQY55EVQVoxNAUcJUe7VmvNBnmr4x/GD+ZOO9T79bv78oYFJqYZtrV1y08dMeOpJE
AE02HlKtunk43txrAFZ4fL8fCRwm1vJfHmUnCCBRS8gnhsC4YCNhodcUtj5lK6MdpZ+KYX961lmm
VbWWKfDXAA9oEgnkVQ171e01kHtkZlHF+RVeyZ1HGphlKHkEalTHKQknCCq2vxBOlzVq278q50Pt
/KQG/Bu8YLWwpVHVyIG686I5dx2h2mpYmEjzWQ4OmNA4KwgER/KCu2SGKN/4WsXKjtkzWhzr9IJ4
yewwGfMCEd7NadojFbL52Z6YnClxiHlEHyeD/aH+AtOobWz4CQ5GC13OWEfv1TnI4ICPn+WlUoNC
UvNVhnwSY1V8P3PGWJ86yu+MT04+er1nwQNBR0FmUC1KpgduXYUC759GOK0shp1HpirucKl7U0bf
TgxXdQAP4k1QJ1WK5swDOZuS0zMBK2yGH6fmjNv7SvT6fOulQiWpv0KQbMUJntMIQO7XfJIBkISp
7RX5c5AOxTpNLiRBsRvN3ukB+EjIm0HTiAs7essupe+cU6svOmobiNrSHn8O63I4fYREve2xjjyb
MlUx0HZ+CD1KPVX9JFGDfX9iDkPJjLIDgC9/ClwWDpLLZQjPXGOouimZsxbq5adu1Cg4fsgJCZdB
S9rWj4YXGWtEGXt9gS/QFOXDxqU0+unTzz7FjqzvfDvp4rmYc/jB7jnLj/w048v6RuLvU2umNjNB
0jfSYNg51L4Jldb4bfcvC0whS8tNAVod3ezOH0KzmxSWEJyd3u7FxqOaXekcJJir79amTA7vYp5d
0x2ahA4sWlyovw4FFh4FyCeKanVpAl1rss5efDUokpxqZhE5nCSOayL7k4iPBuBFQu3HxlY8ZmXq
Cy2A5N9JzBVwlPitBz9jZyHruBQ5ykHZ1QA5DY6V14xDwp8R+QDF5e+BoPh18ikwMspcKALIfh4F
ai/2taKHyUYodc8mDdZ2cwOyIOGPnszL9XGYfOCM7w1PUbzu5dC+UaBurKR5sA7c3R0a2jHFI4WE
qD7Wx5iobg6hMDWeLDbzaUfs67l+qYlfbSRove9l2Qa+88eBsGCaBR+bFdR9+0mvyICuzwd+Vv8S
JkWJ/RNC8P0x+QkhGuihOhwTNgAOtD/rE0HT0EdsfTVft3Gc1I+SxhkBcDKKNrwOrOqcJDN7z4dy
g9OhUj6JGzkiHAkeKrawLEG/rzK1E5qlL6mBeoVqABDADO5zIDb/lXxRE2QzBndKOCQ1tc0y8XWd
x/IqkJbu+huPOJgXDpwUOnEBEwJT3fgz8XMzHDEHZpLyTbWmRLHkg4YQG4GkGfB/NF1xOcckqoUy
t4lV47LfPU4OkN8SUQtRQNBdFhmdfXLRNSLRS813GwuJLmmGU4iHsaC/MWjW2Y2AUS4sX+LPywEu
57lawLotTBNVZoYrzVcmkmRN4GlGcVLC3TiXblRGig9h5LfsFBKjIQLX6ufQXNXB7PXVaV2zCwf0
BIK7yG20K7ZFSe4SDPBUSl7q7vlxdMEpeR8W3uwSN9G9YdF4Ra16KNRA3bkFQtprnZk9OdAX8LrX
Ko32zsVP9I3mjlR5PxSPojfyXnkBLeauM0POJVSXD1L6AsPj1kDMVytMUy4G5Me28omxhyW7hpou
q7/hL/pDGqa2Z/C785o8Wi9h4xzsfIRaQxoAx9yb/MAnq60eG2ZhWBu+KEdqYnnN/QyBv3FqQD8T
VhcSLH0/DwuqDK7SeNAq0VgOCADIrQwDbuViRFTeNr98HCXgrLudObuuOA617YX0K97ESWwRTQ/E
d3YZJdlUKPQOYE3jiAMoCeoAnicLR1tqjXnoSLaN6xkQ6Xw37KZlkSl/+qjcirETgxKLDSKrvM41
30WMyc4GvlR2FRcZoa7AxteDi7zUKvcwi4t2Ar9DJ4/bIKVVR5CAvK+vwULdMZNs239xdjaMoAQL
2qYRo70TxzjA3gWf4WLVcbN0KAr1DFoUXMWSK+k64EoX3M2PkF6m+XuCb31r7rmvYlnymWgtSx+2
Ctjv+ihq2vi2D13o/wwc0ldoRz/t2nLxpV23v2JX/TFZrH76ufMjRJ29ig43FAejCF4QhZiE/VKx
t9zOFaiCFMfeq/djJgOmZzZcUSFvgdL/b05sr+Z+mwATT7jnUQWQM/4F248RdNq56IfJYK2g4vFx
M3JYeQPP83Avt/ySXRcVdrO9wQcS4zAZkvfQyACuVE7sk6xfQ8fWjwdvQXz5jeNXJ9qzJYf9ofwk
PukKm3VtudvPhUFZLZ4nY8weJoY8S+tQ8Yi2t6oa2Ko1SK/mYNEEign8AjsEkogw1HW4o/CahT0E
CuaV5gX5HbVQzXxUGxG105i/8s0E6lQMXx6SC/nRYDuSkc3PZJY4irdtwckcKcoC6umH5ChDqKI9
SM7KHtJAeiVP6y/ZJpvpD2CXzCZ87ZYCZkNcB5PHv+jmihM7lklop9rQJ6+llsEb46V1C0ixa45V
pKS6CmncBQS83Zs5ctoG6kV7ELx9vk5u9wRGFhm4EcVDH2oCCw3AaA9No2zLWH6seT/ixbbx7OAn
a44s8r7fqsTjI3rtN9hncKE0USoRQqbpvt8dNJiJAnayOYGnN7dNOy8cKhPMWH+xU6k+5ApWQSp0
546/A/iugY+C5kE8eoa30ZHS7pcboOSLb+3UsiwgmXW2Luz1kVKF1WF3ocJsM7ZmrMLeeNjIH7J8
G3ffIqHa0bb8Sst1V85FhOOEjZ8BB4XQl2xe9IPAB5f6NTjkG8KhorAuU0HAq16OT+fKoV5R3XSA
mvbEvgy1Ah/Aq+Xgmf0L3QhuqH2wDrSll5ttdP8nAbT2s/JmTZwyXyhQXi1MuDggWbf9fDyViltl
5d8XmSkcKtE1hrYmcFE5KWIKOVOBoBKxf06SDu8v4Gp4MPZmmmaiXCLSIc57yuiJ0MyTtBlSE3mH
lBlll+gmQXiJVnfI5I9W6AVp93EtFuEJgG3tT4kek+rXGe32yJ4/GkhfYgCAZSqIUdcONGlbh4Fh
Tjwc4q4fNKwlfvVwb01KA5e8gmhQHz4CG1kp9OZBZXR15KGAUOgld2Q9wlXLXL1fT6mR3Pde9eRJ
1rQS9fqS/Zb8gJDtcUf71rhxkNw5e8tkjjNXdKsw40rk2A2+xAspe5Y4gfMmKI6UTmfHeEFlRUPc
KUmhC/cIUjejg9omBfHMlrPgYMo0cXYjzEYjEpFmSsfeLUflEsE445q8/a+B0A8dXshy03mqOTWn
fWeBZLyGKTnux2PUTbWhFCB1aZZJ5XzYU7HiZzS4UNEvn96og2G/2GQMGQxN93tlPJ8NrmZxGGIy
/uEzSG8lmimqpvDBgxc+KsNlofyKJfLpeFCoXExVAKqt8b0WY0iLkOUih2Hn6gniMG2M9rxG9aIO
tyxtcg1WXFqwJP6NmMd1vzgt/8tGvAJoN3x8FJsHQg6OuWKhYIQ/WJ+THw4Drf30l/MK1g+rO2xq
8ifX68vxsQftdJIqB5ByfgsA+Cge2jLCLK+l/mQgDkoyUWDXDpNM/eyXfkJOh7H/cCFMVyzM0O6S
PtwzO6Y71Vq4AcMJhqfGcVF30GKAajrAAHFoF8dWxcOqGA+psFDarT55FXiWKCxbitqXya3+Kkfs
5uGC9SmNrxHDdMt/kASULUDtCwEq7THQ4WQjalqURnTOzhMVSeZ7qrnErqavOsuVG8W4+6H1gOOS
ZNasZbSHYpflDuLnnCl0X/an/nka0Tg3j9P63yK8C64AGShCadB8BJtw3LakrqMiGwG9LmFLUHKN
jYq0Hg+Fm9CdtdmvcIvfRyyyZArpMWcFjO2z0u1a8y4TuFh1m0Wax50P0hzWHsrPRYYP7AFH6DZC
dGxnH5bgJrzJWjvvhloZ2xcskOgLPVHEDzfyQQvXHNzYZD0mXOnB60Itw00ajJBqN+0yiWkPeaUD
Wc+lBjAKCG1VfqKQ5nA3G0iddimuKrDtN+C5d3TPVtjGD1HVertKTl5f8A1sf7ygmJlftE2P5dZ7
1k0NGlVugZQlwyw8qruk0uFRaa+QQ8Qc6S73jkXlK3i358L4tD6cnYw2zotLcBD7J80uvrcGW6Z7
MKXDqZzdcsSY+5rEFy2O51TE/l6YfXGohhFDaaDuaA8RzAn+/olPWyiR1Xrd5tpbSDMiWNm2S5a+
ZtYFOUk3RNyYIBkzetBAffazfwjqAXfw+VSHgX8fZyCQ1Q8xIWQVUAVcDJf1yOa80s2aVHUgl6HH
VeUZa9unw97p/nNIKuouAIgHncyypLe1xDJUJ+vU2ZFLxNfLtRe6o/vKvsO8lfgXO64wpBwqeaZo
a+ivo5j86916Z1dyraqeVxse1cUWknVXL6hI6gX1TABUiU9IKaEuhEiHDx3YSgLMtPfts2h0VLB5
jemE0kz9YtnJV8tj2+ThKDH0pcYR+wFf0zpEPi+b5E3lMy2n5z/O23WAKe33OK5/8dCN+fRImbEg
8jCVarOt8+YcqZ10Af8KikWJOCUoz/UBKh3pOPVy0MXGbPX/u9g7gfh2tCFbQ3pqfRUFsNJOrv7p
xivA8LLzkPsBLnnyZEhlhkCvz3h+8IFvvIyELBT3qYbdq26DBvn70P1w0+NLPAFmxkOoJdClDDZi
C15GkHc7YWZKmM3bs74LLs5JuJl8HtAJ9wh07sZea3NEO0bAdyZsTh8nRRiq6u9JYxM0kqL3Wf1/
yN9iLKMVw6KfZ6oOxOsy/o1Eo9TPt7wiqGC1zd3cXlkdl2B+o7CcgDlxrkFYbSUa6e7WaBsxed3g
hg+GRPcA+yDoYbvt5Lz8TnCOSlhByXpyOyqR1DotQ4seyPmHBMwxlrWXquUwETYoIvEDDf+DxZCl
xTrdyV/GYcvFKh8GTBhmJl3+0hJrcsm8mRNpnpXfOyhQXYWZ4FcLKEOb9/PQLLHL4IIcBAUzt//y
2slJ23DGq/T7xGwgXIGrsqx5w9NJYQDXZcG4Nz8zSRJNKxM0RoO7HqAZVPVGIGl5qgHnCAadw+wL
SMUV/wEdW86JDFp+60kAVMBkPIx2Mpu6372Aw3XXgusyuTMWwIB5cYcIYpZA+dcL/8YYCiZP22F2
tw88cA8aPUu6Wc2lrE+2Lk8+5XbVq8wI2z8Ch6Nngta+88vedYHoc4GtrfAGlxN5Y3LyGMDKP1tw
fWwfUuzeqsT5Uj10D6YWL3fatRd5Cvqv9zBybArMDTZFE93Q/GOI4eFEA7EgeMhTsRNW7et5g31T
SPAzcpPUEMVZQn0MHoFmeV8yLSBxYyaF5/7rkzA6oAEBunkpW34Jp1jxdyH9RJY2DuBuHwOowfN7
V/Mw6wKwvacih47FtsKGof5I0yicEou/m5tct5TGIN3jdQLf6y/fP8ledga0uxQUipfDKWZ22sgK
LnnM2fPvf+MvDRWfyInEXEBsgqtKv7k4na9KLP2I5bJTZK/5iYTUJ7nyebc68dgE6+xJQaAP89WS
3wDUO/u1BRVIGAXmsgMtGUKAVkys4hSKTC54QC/H9SOWSkx5L6c2x6DMoR6WR+lDVOLJs+kH0yXu
RHS8bF98ZaUtTcdCKLykPN4fiFEz6tuRrh00JrPs8ZZo/79nV7MhJKnVU9P2uWSlpe6j6B+VZliq
tqIaCrRYqoqU1DhBdySqbUuf3zpIF2qTeFqCDnGYFcxDe40Cs0qxNIJDHHgBUyvq17NeUs+zKvO2
af/SvGqmj/FbQBDDaXrXRUwNGL8jOMo7S3bbOHp5Ia0zz1i/erwGv0VsPKthRK2fFzTCzx6ku7ML
bxTkHhOT4BaWM+TEkhgQkJmwcoRF4+/By9kdaCpa3Fl+BptjDh/zObXveXzXEMSfq05lLkymHuyA
H8VWu44eTEhBc20kZcV6cb1UEFLbQkVX/iA0txol1IhxzFTPnFs1+lEMnzOy+W8fkO5831FC1oK8
02xyxPhaWRGU5IJZynmdreaPOTCLVjGXXO+jZckC0NSn9ouEjnHqxzS67b9r09+wNNLyg/420WaA
ULo9qQxp50gS9dztn6jfi42rq16CgpzjjVmSBkr+ZoWNR9txrGV4rvBj0tZtlfNnLIyFlNjgVOET
b2S7tScVhZBNb1Vrbv21I2jd3JzwyIeDqMjDuv9m810KvEyZACbSVMdXG3Bl7+GV281ubQn/GnL8
EXwbetMyGn651/txyg9pkqIioZBcmeHeDjVnvV1uybwQUVgJxYYC52vkn/ADswbIe6dop0vKbh+n
KrXOYR+9ov27NUULKB3+P3iBOrI00ex/iYE94KJ2h10zNvuAf8Ph7o4VlNETq7Nxlj9SmBwF93ff
G35Bc1bBJRnQezjL3XzcHsfOYV0a/M7f5cw58KF26RI5JUP2n/B965zeHk2FlRf1qt5pTlGcRG7U
kLyewc469BmpnFHH2/ja8aiURSxiWcNjuR4xeawh0UW23+HEJ4YME+jPGRqnB8jvb0xfXV6p1WpX
PSgOBou37Nc7ZlfeDpvFWhcZKSckL3ZTis85Iv57r2Tn6RiDQiuHnNHoLM6DwmHKjS9zac7x2uPN
S0GPNWhE3w5uHnynEZO1JVs052p6Tkfo0/L0veeq9MrP+hQyC3FYfHLmhHhTR3hgy6eJwI4bS5LB
v0uPk6rUc/keDoeLB7pny+kJAdKzMlfq1n6x4Nh+PVyi2FA4bG1815QQYbbd9me/Wu6HmJ62LJ56
m3c5t3vBvU38zj4uiifCxjbjP7qLfXPV8huo4jsX7AFij6KnCtAASMGYlcObOEQngYmoiV8ROAFY
KS5gASKOZbsuCSawsM0HrEt4WDCEsAbNoilf/fHZC+/VPSm9VzDF9uOxnAYgOvN27qIvHn4JTmde
2WIiSwRbrcjZcvDurRJR+HzjiLFOcXDXut9CME0boqBhjd4Uo/7CUEoI5oxmHy+kw0647/c7NrKg
kE2xRg3nlurwrocXyMvecxukooh792SuWR7SxiaDYN8iMip48VgbeQAgcmARtLy9WB9Z6pbKDyIN
eGouY471eGGWqe32Ghn/oSzgqUvyUCEwz8o46SY9g2IblUxA/jif6XKrA3LcUbl6F5lDOSUyTR6j
z9b4M4nN8Fowe/cmHZ7szQjNZPuq7hBoRZBbJvGXN1vI01CTr9H710C67bu47pLmm6j6RM78BBY1
KsAcR5DzdbQdd2Yo0Va2nIi4FJY+KDopqmIAJ4atRWvqCdcnLfWOiv7w4n0Pw4CWei3fe0LUntJC
HpGlZjBNh0MIkkNcabpmndC86O5Jkc4zkMqp1rADvEWlBoXo3hypLIkhDaRVGzyp3d4FMtKnCXDC
5QXcdBp183kiyUw2Zj8STRdlWuw8/KIwyERUfcDcju5owE36lAbVd+tLAFH0xdqsTlIhLoAU8nG+
BKIgrx4ArSgoLeWk2J2MdEDqoQ2Agdf70p+ZqQmjVL3ey7JVYOmMpJrIlpOL0TZ7pHZxzSv/98me
DK/qt/v+UqJBJW3rQtcoMRKfpGVmajTQXRu0sA8YpcHjHX4PiBJ6lNJfgJhYRvSB6mykU7XSmmX0
Gj7n3u8wmcAC+lYUpQsS2OiRUIvCNo7EUOvEzRQKlSDWsaciu0lzt10bV8gHgmUytmzZ5iHPQ4pR
KKVYcWW3RHI3a/7a/dodJwnsoYwYFDgFr3NNazHiSsemHiVgBcCQtqcTy7uQcmTH8wAWcJC9FPmg
NMAP/TbYcUc4kaqRxC58XYpGZ2J3w6KUCwUE4aGzPMoTY9s1sIzqZW8oTqtMjrMzJlIEaFbUJuYj
Sl8KazMmpisAV4ZSICfhUgRmNXGvSIwPzkxQtLHhIQ94StqFMKZzUP9jOofJFUrV25PL/Iggq6fw
dqUMPwt3dy6AcMLvTtbdsgnnY2d3Wbiddw3NMhbvLR2LXbtddbkuHkeyHYQiywRIazNmDcfqzOq5
kYfr35l6zBCSFQ4kHQqtjBCiwQUBH4M8h9TAi1rqtjV6Z4mA2IE1g8+4ggrcnGAxcPk4gBJ4gWso
BtCmF+bEjTTQOwSHyCjYUiVXvduHflQukY0THT+y9vYZEponXscqZlqu+V2lIWzuSTmRnjs0ktSw
RYOXDg7GTUxPhcnnWyp41PRIXbPGUAnD+xnbkPKMfxAerGW44qb3rRWHT9QWf41e9dToRNa3aYzC
TMM0QyGxnVjNUNsob9X3N99crum75OD/F1nZS7QsJMaw7yscr/qRPlMFtMCor16GmsIRnCLf54F3
JS00kxQb9ZtuXVI5YO4ailE/P/1gweN9NDo2teIOOOblEqHnzrMbjffXKkisKSUWOfuntpN/7Smq
u8KTzL38GzpKQWECkB1WCAJ+nvk1udR32LfkbQxeLe9BAaZGJMPvYaqJQoiFq0zSdBqg95GhRV8k
Ent2Cj5PzZ6yRwlnD8rb5reV6i0H+3VH2HwGBLNhEO5qe8pOvH3sSvQHh4EuT7zmOnSVSBgLGt+N
R1UsTBh74xqXEq7DZxUY/m14B+Vxb9A3Vt6jePMsQDJfy5MmxNdI/V4LTc2KI+fmK/rRbX8VrapM
wil+4STbrEn6xHkf3rNE/WWvW/4IG7vk/Dogtb+5CYEinlvB1tzUr9CaVDKsfyw579uAV9UwwaRP
OvWAuGU4NR7wPblXdiEBIFtGHscpx9b1lrPet2Fyc+FJ197jIDAGuFZ22sHmdiDrP9cQ7D2qcf4W
e72AmmRe9ThWtsSCbj+lRhbV6+xYlIxyh9ILQRsAa6nWcfV4Cm+15u0LpoSKPgvYWeChtOmWm8hz
Fzp4Xi63bEe8w8diwFTsmfKeHv/mW2e/E2hHLXT/HeE5SWxzGIwucsFKgV84zShwMccJRw1mcQpa
cahudHLLhtNkWDVJuxAWpqHQcY/jjPQZbPpxVcVzq4f61hEWj/O9TaOce8EsIk942tNByI999xrh
fsJxofobo9c7lklp+vKruqvHGNUmCxjanV45DbJbRhfeCY45z0NLwFP+CEB3itreGfZRJPh8Hvuy
K3MjwnTQcnA36uEY4VMfBYFGOuyvX7ykbIVajJkirfKfsqVLNnkPfBF8ER0KyDz4GJVJBMK03Ois
YYyrGOGjyIyWc2RicwStR0N3yCeFYRFXC45Q77gBaeQ5Q5HGoddu2rHLDSS/x/FvO6UZVIjTnBGH
rarrJqwTD6de2SrxWEDLVGOnG6VLkJmmatyivWZSFNFBZYUl6AfoSGkmRJGlWCWwyUSvXikBIXRS
N+Q3Hbj8e8LL5ZH4xP7K9bEWez5Ka0wgbjI5tQqXmwFlO7kjNxPsVrMilMamDJcP6FDgma4LgvIE
fg9SYS9FfC4DamE0srsB1KlP4BKRRS/BH7mKAOLlM/n/+kA8E4f6L6mT5Z1B3ZWsREZGafXO6W/E
A0Ct8W4qyDYOQoQ5zSG3pi7SlDrOG8FWQCwvJCAzNHTf5bg6uv22xNVC5TgknF+Lb8m08QN55GXX
KsMJCKNV0/rBcMATQQbl3MGdam11+zLDgaI81rkJozbP+fo/rbnMAmr1w3FoLS8MpEk8smFeK/wL
pGJWTyi1TXAsDYJ3VGU+yFQG9NtkENqHvFOPJqnmuXDyAGUH/lff/XZcSPTWLwhG28wUsBLA9X4L
LxxYtxUXURbiWrd4pxI01ISs2j5pZkvnntfchgrBi0twOf2OihR5s2vvsd2M/nWA5cKVhsmGAiLu
HaWwfdmT/CXCvt51f46Hvbt5eHnh46vG0cQKmKcINmOlWIiTe47fndoenyEI/M/agAx0AC14P52E
so+5snSqRkmf/PCxUc1uxnSkdBodsjLPs3GZY67BfeIEOoMDYSlBSq/2mBi3RM3L+rkPOscKn4i2
1J5cj5pWST8PeFeNpOry7Njkpsw551Ws3d+FaQZkuvMOoin7MhGu6o3FMJEfewW0iFHhwTVseadi
apKcU9Xyb8cp3TU+bzhth1jiPPtYzEFWmCvxTRRJNCAnkgOlrcSMBG6Q58k/NbEkBQz9E7BXCSL6
aa9xESLwGrbIIgxtphXSyAz+0TVTG/H0q4ny2wNPCyHcmbZDYQmmAeuHBnoY18Z1HJaf4LXBgfhS
UJtu0/AN2DceuKFmNsT1RWXgzxDCSqzZFVthoGJvS2eMIJ8d4q3g/emDckmlGoQuObjOOmoG6L/V
VpPwNB56hk3ccDjMNHpjBcL24l+VVvFahoOOimjoX1zGHuFn/ZOrI2Rz978hg1WQPeZQW+KBgTzL
UztvGcvaM1XKX0ZpfwG+999g8L8gLXasNNoajkFsKusyo4fywjtwLCSGvGcnKff1QVVeExiPsjpm
N5DMWQNbfCecG9S+/h2ilEzkOKFAlwRtBUTOQvcgdQUSOsbQ6VyQ30j9kQ5aIRqSE0nsymw4RuW5
c9lPItaclW0HTKFvlv2vPwrD4RUmv/KZAMZffl0SLt3irBv3PYku2mCsh8PBdRn7LaxgKDc7Nq4b
lMC2Edn4WfFPOxv5FW+F9rfvgozs3JXTZXcm2i1ENf32nz40idmvNJ3O5XCiFJQa5Rfn1QmBAq+J
K9wiSR1TXCqEHnS0pdVz+DMI+5Oz5Kv2ZE/aajNOMlCAKl3ojM83acWCWUpu5cVfxH9+Qp6NRl3Z
K+wxdyNMg2irb5oY2v7MjJJ926srBO+6PRuzTl2QFl0IZ5T/RNakCy9MDYS1wjeaemWHA2GULakl
dWzw5EMftCa0i9UqHOyQEKKQ9h3mmxBi/Jt3Fxah90kecpWED+7fYDppTvNtgMNnXIj5NDsxoVuT
OiDF65dtpWLIht+pVALEzSFCBO0YHnDaMrngn9lSjLvp9ekPgIf6CA53gG2O6Au1s3fqO1Y/DRqR
TD0mJHDbEai8Q1fLW6WKC3Dw34831P6cVk8mb2T+MMbw53q6xa38wXIU+TJI5/uPef8atA2rBIrL
W6/ZzamQofP21bGbMWySFoKgEEAY/dVEgGMwCtRk+Tu+awFbqPJuAc8EdkJ3ELNxTRGCDKVf9sGn
fh4AmHHCaKKcYaJ2nu1A5nJ5eWcEAbCe3kpVF5d4IWgScr3fdO/MxN9Q2UkJZhMUPxEAyBW9OvwD
j3WxnCZMXfd4znPR/ABL5yx4FK43yFsI4AhC45ZwZxssqtjuW65eEuUNwMsCXl3TAlRC6n+E5XT7
WoyoKkDzg6yV2KTsnGXTFmMsUacdgSx0Frsj7nhEMh5is2/9G/VXteQi0CQ5ffaSPlE8KG5rZFQV
c+YC14ftRdESJVe3YunK3KnHQjzYLUwM8HrniduArrUVKGhIynyi78QKt6iWJBE9mGFt1g6aNFYY
DnHnYHHy22bKCGwK8P5UyKndsfyfjGNvv3ZzbSrXeoml/lW7c/kDp9ojDi8UPjKHT9dosJkWplb5
5moTcLFdWjligDMMBQlNI/Q7mUt4MrloX6mXaq+izShhQWDKg9inAEGaSlnALJJjdaaAv5Zx8VQl
cm8fusE/ss/IZGuYX1IKZoRtA89Zk9x6W/tkrnLFdTAk83zNokxvyTXUXJFM5uG3ijvGSNLguToC
yjRyjVS7YQLlak/AaeIy5wxiBE0FNtMe0rx2ryggclqbBC1hvWHr4uTkKeRcPkXURj2ryUIsUaA2
5JTF0H1r1iuge9T3zJsH2kbirTRtzgd4Nm4CfcaQZh8E+qKN7xKiLeZcCcF8LmbczpqfhkWwsIos
YUfwUv2uug+kiskAwhd17VYAG7ULyapIMahZ1IawCVqoecIVagY7JS56lermJ2RLz0r5YUoLZbti
BgCfF2JY90o3vyZimow0jnf2ZZs+6tSP9gz7HtjQeuxEfjb6kz5YrnzUa9WT/hVdK35Znr5XNUDw
aR7w/l6IVEf94uoVMNVG0L9UCYO4xR8JcLDy9Ib2vxepj6Ymzi+FjRBr23xR98Oi04XlsyqCH3sq
vqFE3y0WAgUVP+i7VW2Qhx628aQ+9x877WP3bNDR1fYn1W4UutT/Syn2HT1GWTZBGBVYb9KNzA9l
TbGAEBGfele9vzDnumChEq2zsPfT7dWZajHDH/ujS4kljMkgXt3yB4kYLhmTODK5lMOM90jW63GI
CQrGayHJfWnlKoqLyuHEgU/WcuMKMjcQYFOBh+wtCtfTedm37CMJdczAdta1HA+kzxmzMMqGCbCm
Z4a3D2DaoCKCoLUott373+c0Pm9QHJUFhfWNUXEVAhwuPaYwVODwu7VQCw6h2QTTWBHCciNhTMb5
adpUc+C+5woY7Pc/EbPa9+lFlXo+BhKa+cDnDMlF6UD9u3NKNFrtBtq9zuL6FAsD0o2jnTQTjoIw
PpBOTkMAbNmpABO50A6c+0XHp4VhdSaEHNv7/6hNYW1VM7BxHv5+RMmjed8WL/OgJozGagSDZi5W
c5nM0H8te1C7i0ZCW78lK3eMuthE10YYAuz9pRPo8pYL3+Rx0FRpS1tADcSy/zSks9tYHGn2zfE+
BUcB6KlBoPkRNfctmgdIgrZlQZiFO1RYHnERmjbifelZfQU2C7YS97KNOQDiOwH5SkLqktVlmUWp
irUp9f4CMWEzix6v+/AFjtvvrhokDK98N5EpktWyhzD13pp+SJJanZTsW/VU+fvtT0LPHdtkuxg7
rBP64f9UQdWNX6tEt6YBwJNPZvqN4lHW26AEnX3n6vM2Ley9apO1sMKZ/9b1YtP8+EfkD/qqgYQp
Vh44KfDFql0bCZiKTqwh+1hoFQpR8vcHCprkpkngiuNGjQvF62So8TGC8i8gJW+WQRsrfGYRiekP
SOs/PSKfQTueonBmRN4Lq1YTq2shoAcX04qQg9FN2ER4ZP0qGB+ltInCxFgxf46dcLUA/U2qr9Cj
QS8mkClfI/8MWH3vhyA+y1Jyx1bLqyytroEDSfWGF9RSvUWqeJad3lz0cjxlQyAgT3TwIMC9nvwx
oKCuEZOflVptLyenYFQtlOaxEA+wSh4algrD5xEznwicJu2R16uyhPBMC7TLw2kfPCN5mkWLUBoZ
jSdvqdiK6/9NDv3C+6fWG543n7J4lzmM0sYdIddDFCTaEDBN1ScfvNctVJlbbLA0dOH7hLDE+UM+
ec76anhQleAhjZEhMQMflJLOZCarKSOZLN6FdAV/GbGYL+h06/lyOT6PCMWgBY/Gy+D7Tev5w4np
/d5RsVRIIdvCV7VmLTwwZKnYocpqqE+TqcM9d2sZeBz64JJAHbibOSCAK9nUcAGhAeeb4JJdSQdH
qLYC3s3bAYEewfzllvGkrR+yBO3hGoivULWUfysiHwEdVU7PQ89JNTdkvpvhgM/ISmw9VNd31cJ3
VPGnVCy7R652lwOZD5lZtl2S/JwG0FYz268qEs0hO20I3COP9oSSfDnoB9S4eWF4oCAlnDAQFNv/
1OxMlPJKv90M7W1HFX8bLsSMQ8S/dA6fFhZe/ffsCjvB2hn+mfxBLx9QDCwqtjv3CdoqXRmIcEIL
+khPy6lGOftKGdfQY4B9ocrQYUdkMftBhd1EgIzdPRs2uBx421Mnntgeppqd5YWdXl2IPSQDJ7os
cLy2FLyzJsJlTZONOdzoVgYBOtwqyunK7Hp4luHyPPx/Msoj9JVDnuirg8fTuCXcWW1cm29aETah
9LECro2dTDrL3p4jIw6xA9KonEKWRvWYqEM6dHtLIFEWDcHPklYMwJBR+R2O8RsDP5F20OXjRXIv
/mYkzPrlEn9pCFb/C48DnQlfQA5Dn3GTwbMneNsnrDpTSwRSRuS13ZVW+9V9BTqd5XUnjCmSWbsK
g5KAcj5sVhcHT6rqiGbbp9Leox+1AE0YA7UMvqqtOnLmWm4/IYO7bFnT8GWttkLmX+gTmG4b6wYJ
8+JeH5pnuEKn72EJjf0viaT/lMDIb7ZU8GGninPFmzMhqIyBYsIox3nkUqFUvewSKzhKpZC01vhs
V/bkRtCcxnthIARICNHtIunhxIyCOpMHrpbmZMj49MW5nhtdr7jtxCRKx+cIy9DWD1a/Vh32fZVR
RbYuV7Ce4i74g3ENF19c31NHKV5QzG2+Kv/zOEgOqf9huEeDPva8iSlveC1lLKMWk7FPWwc2GAi7
wCtGWQCcJ9ar/AIVCMeaayahOuPKLv31/oJkdRYqkG7e1kBohIZsIcLGZ7rorKn64oHGQ8oz+Mpw
B+4t22fxUnFPqr5MZ1wA2DqNruHUr1KeJgZVDMWq7+nl0P+rYS+lGhKv+XMa6BNlxAOA9dkME+1C
ucCYKT/b46TTMF6rxsxm3O3TkvcnnyGgIuleeL9z7nTKpFUrHsztENQ2xqjPAG4ynFIxGcMn2yjQ
FYs2e4SnKsJxbfdShFaHJ9GTo6tLealxwPU/A8kEoU0BttRuIPNqmuUHEx6hue1AFMXdXk3taRoo
O3JX4mrB6gko73dV6slT3HcbPc8kzIDSbpUZvDIz9Zcn7v3Wl5uUDtkJC7akbSYmVlI70SLWBeAt
tNYtcm9+oYbkbP4R4BX7ZGoAptl3ot3pHLk72uJHf1OIBmyD66k+c66mJA1dr1uW/U9Ss1OHvuNd
yv0usjsnsGXG8DmWb28hi8T+UH0McrGm+NGPZlfUSfqHZ9jI2ifSEOtDq2OJcx5l87p0YMCpo/pr
t7vXnj6ChqI+uXgMTgFfFQCbo9PXbOxrJocHhk9XLSLtKtE9rB7I9qn8w6eH97oTmZpfmCdLSiuB
9d6QKlBAVfFLaEpbxIO+MH84I/kz6TxxfFqZvPSw9yH1k812uPPPSnyI8+d+p3avkbXfEGsTygNO
eXkI/vIjjJ7MfXcdLxmZ+IDJjJqj8YSDrC7bd4p75QqNpVBPYwaZI49xDc0yWLwrzyhnj6wc6edp
Ubwlu3f9eWNedOILITLH9CE5LQwV04OygQuneu6URkSK0h+O7+nWgSAMXUsOKO+AlJmMMFbepn4V
EhZeksLbCDQQ6YGCIiWrhkVzveFo04Edh05uaCmd1XwwUa0/1CVA5XjxhrGxtuKLBx+CihXKtE3Q
fNMgYCQcYjipKCn4/uIuFyOkTKJ6bP/DPUR2DsmqckIsp4Ps7jU5BxawMkQjE52/4Si+XsEum8PP
EJIDNcurk0vCn36PDnULb6FQ6YykCmRqQJ5DfDtAjbmx+jLf+/AhVopwXHgQ4vREDQq0QomDenEn
6MaIbyM2Rq96gufeSVj1eLlncubCfd3CzHu+5rDSiRoQX/3lgT+8oUwSr+LDJL5dvYbM4ETNSWgQ
umcEZXz0dUhtycFwwlZK4KvqhNzPcQRMOCwu6lXIS2DbTDR0Zp3h3hG9dLG6PRUHAHKs7ZWuASkA
yEA3mQywVpS3RigiXhDfB+SZoYEVz+LrxOBU4TmUkik24KwU6eSnHZLJ8IJtVpTnDYbdvPKC9D+E
l/og7Cd2P5zEkGvCqnSdnaTazQIyUjMP162zRxgcTz7ZHK2EqWD/w0WR62y4Es2Mv8MB8jlkMUc9
paXyGxci61tdThICkJMPnBsMpNh9snTcZmoUOurS41SxOZuwgx1lhzCMPFbaFyWPzJBaGcHZbhgI
qbUas13Jb0j8m0q6EzbJLVv0mAyf6k56MpI8ySo1v4EYq3wEaJxZrJh8TMflznLxuwJEgoK066uE
kUrpTaZKeUmtM6+uLIE+b84JHNWMOJu5Bx5uuA7I/qXGzd76QbC1Mp7KKqq6U7Vu6T/jNr5I91vx
iH18wphDwQGK9gLMrr2ptduzjegr7HfKT9ZoI25gebXFeIiR1G6hdsd3FRGpECCPiFzEvJ3GE1ot
lmfPX8+HvdDR6/RVwWuaujWM84Bu9JoJLxiw9tg7hLZ2w6bLTl4u+DgchcnkMGxceG2jeWCtKnkY
MEvFuXxsC0kQAbmllZTtqCHNOSrpOD1zzDV1mb+cSuevWRurFLKKhZ4MGF1B4n+42+YrMdHbFx/X
5pT+7ZeTXSyD65/r2YJA+wCLD+Bd7HJEFdkVPUQqZ+X4SYtKU9KeHNeX2fwe/rbQyNhEOzV39GoD
YOIXtEBfTxvgeUIQZ/4zQM3/+VuD5BI1C5D6BZbKSd05lq+gZR0Gh2mDCL92PIsQKcJv2WvF3kpW
f5T5WqFYxc+sCc90KRHpX8xI6xaMv60grOxhUz1jn0pr5cLVDQZpxjvoy+R+Hp1YN7+JvxRQULdv
OkXn0Fb4O1PR3HXD/+v16G9M+2EtuXjTIKg+lrlCqb24AgMaGzRMbqYJbjLV1bjVyee/nZGYo/oZ
kAC8akL1LeKeF3AeStqWtFvmw8kQfusv2sL5pZuP849DG1fpnrPgtxCFiuVqqS4QYoV85VT5i/mi
FRBjXicXzD1Si4uTGDVqpos36v7+2yeCPeTl7sYwAVwBRyXHJx3qDuFCxuUCMwSR425cGXzxgelh
Ink8DeJDPdqBufj9LSJYu15AWsfi9HYPat9gwTgAmvnnrliWLrHFNu2NoQ6hUpm7Ok2zjzOA+PeP
yC4hDbh+91b4CdvTB/rAN6vV8hCFVObMfGIPJ39Xi1O4elaNoXrRmmhStuZuJDutDUhAsvU+5sQ2
CAe7xfhcDQGynCbqcxGKlfZmzbeca2oyO2yqT5jCpPCtel9kAo6rvsL5iBcZw4eoiYoS/p02OtSw
nnanmPglw2qIerriGWYgD/RvzuKmGoOFH0mi0bJmHCzLa2G+HEshl3LsIlApOtdhKKU6ZDa8sj/1
GTgztrj1e956QYMXBDLTkjyMxA1CjKkCD7ej7ekEe+yIDFGgniFwNzYdwmvdWuqx8vGmBPg0lJGO
EOYnfMq1KruareCEE11U9ggTuJzeFLm8GOtTK89JuLQQ4RBd3tHflcwD4L5kZVRd/ADLfEV5LK2v
pFeG+fv58xQSt7M0Vl42heY/4g7/0Wv+zkA3Vyp61uKlWcTT0EWFKnNTRJ/gTMc6eLUhBIKXJ3m+
Q2DEd1vxnJXiMGy6fkMwB60N8G2LjitTsqcTqBbKXz5gwmMKExH4hRsFInDfa1bvmyw9GqSZu1QO
jYvL5HSkpWnuRR5jN+2h73C5AA4QyLtB/hUde7Mn0nqv0fcYrThLWBCfGn20bkeNW4EjU+rc5EDL
ecl95ta4jSr8i20DfUrKWEm2TzbmmkVETUS+hYG57EEBK/DJqYCfNBWohq/og/hDcqQcDB4htpOq
x0xJ1iKYzRo+2iRqZAsjQRc5R0bN3hQ9SgnWzuOFCSk5P/GigTJJjOYbFPcwrsw0/j8d1obUQ0nn
MCObKfY9s7Kmjvuc1tSunpl3pKSI/EwenNrO5TdR0y/1+4BmSxwo8YKBAtNa4lxpN1y24IuCjkf+
DJ+GZgCY7bbMx0wg7jgmjZc+C4N3xjDc83X+ymSUT7jdMAy9D186bOZJOBwvH0lUnc8t3gy2dY8k
jclVsVm3SOvYVYZWGS2jdp6FD73lQ6dGrCKN9++Au94jvgmTvfL5BmVr3OVHUARTCpTEpbU32FAL
zbXYCtyHd2xproOBjqdp0KX+79GYb+H3JocZIO/p5ZAZrKS63PZEdgpYO5OT8GBZr8ZoDWiQtCHl
a717S+kSHJrEbJOL+mo0f7WDGlKKw3GSAlDRKVQQET1QjW46N0XyJ6roHVFCketB0/8CGmO1r09o
cqahfYvk70/R7PmdGJvrAyjjIKPyTl+XkvzVq6JGH8zubd2pU0c441slEWJZdBvzaf837P2+iEnc
WXvMDNM/bCWzXcYxS1vDLIhkU0orXWPPdbjZpiR4GCR2pqrCLb3039K1OZGI/F1h2xmyiPfn1hm5
cvjfP7y8YlbnZFHZabNaD+4S/F8VybDrP863QrmGOU5c3+h9NcoZWHrikCjrjb8VltFj5Rwdt8+Q
J1ms23YTSIj3R5QkeKupRNlj62nU5RE2Qx7ib4rKtZSj8cn/8OSUb5dSemItBAxaU3Jg5Q/g+a1M
TPGZwa2iEOck22JRBxiJPXsdug4e044N7BtJCwU7L3XFEK4wQJjkgRZ3xD65UkGxvcbB+T6EmXJh
lb32QJZKdT3rvpSwCFi1MrAj6HtVkzl4X9Nfk7GObU3O299Qr6cqEU5oeWgbNbqkhZQk7ZxFOkr7
Gug+bz7lXF6QRyLGaJCUNvxevSBZaUwJY85nasH5w/ZT8mia6RPzteU67nW3l/RYUtm0o4Mp7ZeI
LQ56DeCxUMCYQqxsUpxMbwzciNzhbBFQhg7VdGMH/t+jgH8/PyHTO5FlQe2JN0hu+PArhwvVtUxn
bF5+FySC8n5q6nXjnFGRkZzoWJ3oVRJmcFS6cTv+sDaixxkv3cZlXocXeyvJ0hbjNZlSoZTze7dU
wD6ikp16xwJIkEAuHk/kHemgmIqyJjSMuAk4t+l/uqhRu2PG19JQr1Qw9AfJ7NTV6mTBjblDWg7z
a9frTrBugmGEkwD+0kJchiIi1wJ2MzFzegoawgomjnR8MT6Ja00Pw+VaQ5aMfcANs8TyiQXkNaga
qh86rx2ocWQCu5ZbN8KKlrXcdgDdImBsLzWOvFHEIdFMxejFa/a9qmcABksxdsSF5xaCi4Eso371
0Ud8udRXLFng0kalA/6ZraYgT2qv0EznbUaq7FGntKqWaSBcAGGOnS3Ck5WGwOdy5CPhCz/Sq1/y
LnShCEhap4iHCauGpJL4d0rRDi2p2xYrRjYIR3S2wCC1+lPPXkfuAASD7xMuPLFILRTxcGdO1Eab
4XSlO2IBOdZXaE9dwxhWBF01PMfSLV9eVnScyHGkfxKsKd7QHQyS8lTDRf8OYh4qTe/s7rxJSPNA
N8a+6twVe2wnJBC4FpekvBfdR5HbUriSKA7cVHimHr0HKMJv9/WvAUrkRf8J67mpGliCLkWfWAHb
MK8TD2R5TQ1q4oD3mtyRVFloZDkeLIIo3r34wdv5oENauFHY0CRlVGNk371oNSG7LXiVPpZrv6Er
2Rmjnl7lLFLAYnS6Tz1FHG3bsLvYqpqyzj+QFoighK4iALrBGlMOwSPdsPLyEP/znFB+YQYrXuWw
vhHUXe+AHFjeQpVBarYXAyuzAxKqkTepSKQA1PX6VsjQFcZK/UvpczuGReWxx0Hy7xugyaiQyuwt
U5cw9YU0c0XOqgh0oUe1JdydfUXsdECDb93U/WuTYVbf7wdaWLcE+q9uGf3IqjqazBjGZH5e+xj/
j8uPHIOmJvxTJqmdtOPWi0cSRYI3yH87WmmVpT6Tz/uskRIxRfFX/FQg5gjzWNYD1mqApcidGEVb
1o32AwPkLAvbhAwRGoob/F51snywzC3lz883BcZEl45c2PdlgC9/lqGCG/mjT/XeYoVZRori9NQu
GfZjVUC7zco36sigqlbSrVtIHRl144YCkPfXCbCUcqYI+71hJgqtaAROEkYBSDiHUFV86m3T6zlb
CpZXGD3t4Ath+f/wMpPK8KWuc7vrkCnp30MXjLxe4LmxM0ZGrfJ5aZr9mZ2GpZ57QAozt9AfJXf3
GX0zFlUV+t01OGOlQFFvyQu0YYHsE7Xe7A6j/PAlwSkEyw9rzp5Cm9batGFNe+mgPF7t0eb0dX5M
4f+ZQhWfiaSiYNIoJyVzyrjoiX2gFP8DbNVb3jPsVIKc3MDY/1xmUyOmrrE53jdQQkaojGXRNB/j
K6yE3PEiu4RcqZxzgrBtFLhXCE3XnQapGs3fu69rE1F+7RRqDMC2MN9gYZDAcrBAznU1ATushxip
MqSnChLHiLFgecmuD1EG/mbREuJHM/ZeVfDHo5fdLaXr4Pwiro3cfKmT+ezI7K/LVnKF19rSVq4u
M7Eya4R1OCPEIpoczSJH4wFXHPmhnn+2sPclDE3nVGPNJ5PZIml4VO5u0DJbKotoPjSEdqxjiVzG
USBWIWOEsJA5soT2munq/n8hD6lWvAFaFwvwKolyAxLYvfNfFPaWcfcWiqIhhZGzHCeEj4Nzw3VQ
cYhpkmRkyI9342R1rhbbwAH0fc840Yx7n+ge6rTb7yN6XcBfqlkd9l7zE/rQ0JkIzkZidnKfhFMn
ABK9CBhqCSBl2Lxs/m48b3GrxYPqb2e1W9v6enjiSOCWFXRRBJ1aVZzlkFNUc0d2EANbl5XvY55r
hbKgLFnB+XbeiHuVRK2i6Hubok1vp3V7hXmUEQ/Ws30p0Il7sJCBNXRxpCoi7vQglbO9zO1ixUaa
+Wta7pdPPW6fOrCrE0fx+YBbOycl4LqmfNFv6mtopYouySsSfcuYcRiweLPsPlFWmCMCrP4UtCv6
iSzh6d5jsNyqh7A1fxPFtA5ovKQsPZCwRcpEY4IUdNGIVueEG5ctRm9HAulrV2gJczM8DWQIOb+l
VvmPlXPaAS2dvdSdUaDHkaFfUEev+ecqbohjm4vBUW+LBlxdCv/NfexdHsS3mcv/lIeWif+6FBXK
UHqgpqLe6s35DDdqKjgLxgxaRfhialnLgBoa6CFPpxHRjIqmR4Zri+PmCDbqw15Idft/vIIyugye
EYvkI03Y7VDZA5fbzFcXCbVdoAFY5TJK7l2gqdVHvxAsH+8PVyt3xfG+CeCYKe+82jxCpkNuQKl5
GpoIvnU18yrw6utxfGxYe1aoDM0hQcCaKtA3+CNzf3nVaLE/98sfKACdKo/ZMtFlnqIAWI2/NbSQ
klW7tnSuLMj8ksSi7idOaZ+mFakJTpNye0fiVjaS5FwLRe+oQePLAj6iRL41vCUuEYn4MQzgab4n
u0wtGYrJBGT9bpQYVvXK/iUzE7wLE7jVV2VlZrdrb7QG7HYVITexbQptgsICk3YucfzQwqPj/Fuf
ieVqoa3P5NZB9/lK6x4uX9iUWezfXtTMGgOfKGB9XlJlkLjRunB9YS78PGtgfZzIOr0YMzwd1nlY
IZ/hjML5LlkcwVNqCDFgJ7FXDYGniYEyYYDu0PDkY+P9bUuRQ4BmOPVT6ywQqHYgWwa6wuGQnzQp
kinc2x4upVtFInvsDttXPxnAqpdmJ7NsA5qm2/oynYYQGWAl18a5BWIFbkIsZRNjejkYM1gxYpH5
yQEgumRnqLhEwPOqxcRB7ZO7CsAOt7tavjdpSL5be6/9pWWoCAOgkksv+WNC2Fs9MiLp1/nroHg7
GzNY6lR9JA4kMzEAhNsPgbnk6R+G5K9K0NkEsFCJ4I8+N68DEdBMZ+LdFkCBffBlDTnCRiSYxOe8
CaKH10Bm1XBgxHEW2AYUaBPax6WJ3cEo3wGcKIWUh/N6sZprL3jHu7E3h+qIEkSuZrfZUqavtSRi
99UW5C91hUA37zCWELoK+B5tOBPVDow+Zr2Kr2t2cXCLdxtc5RWqws2QDe54cG+i4iataI6GSbhz
nAbxOKNcwHLzHUNPaz2WNHkctF/BpCZWLBdfK9iQRqP/SOykjk9D+JmqdiM0356Yj6PCAjiG3s7j
GTVI1Qfb9VHwCbLJaaNTbG7sOHYkipqh4eRgc0o3Ybo70MUcp/GUPPX4w77fskfQbYHocp3IqnD0
2xtJuj0P3CbuBlAoWNi0FwsI/cYXZgGb79avWMfO16GSfVMlsqTsNwHkMU9ty0WCILhFtgn/Rf74
8Kb/FsuJeGzICU70IcuW9FI+WZew6j9300l/RZsRQG1++nW8sQ7IlYBy2wZZJTaJhKbumkmSyuif
TMz0TDRATGbeX/U7G5duLNTDOxnGlZAbm8/MIz19b7dqjjYRMd9SrVTSN1YNXSvcSW7u1wwDBd5G
LupW6NpmvYzdC1VAQthQUSpn+Jh6MGoxmVki8zGHgP5DxRDkVFzzKbACXt/yH277bPjgZCZfKLE7
gSzUXfZjGwtrQShDaE3Tt4zSgmOc6Z4vtyTvWRN6rxlLOzn0tSc+Cgxc8WXEAM/QPrh7ho7q3l4H
KGy+E/NOrQJYJECAg2cJwR//9yYFAtvOTzdK7AndeYcWTIgmREBabVjVAML4Tnc5+gq3W/HX+f2b
c4RJtfc69d2Uqy/4dsd9vfleJ94BYYgTcMT4lqzBKD/cP1hkyFZhMwe2cQ0LLsctoOH8wBM9T913
jem7AB9KqJMnu16FTNjtcKkpdAlrOAZhPgZdSd11ZNFf2TvxZe/m+awARLnurKM1k+5fSFF4bBKd
DIt5TwZ9meOpZ3fyoGlhe+b+A7NMomJBhzSBY8i6X/FV53yiydP/KcitzNoVu65ru304elRYhRk3
4O5TvvPq0TPrHcY5E0v2XF/PUGNOvp07A7qVaoxrRkahfL3+ZocAbyKnbDBdGQN9Mck9E8J0vlKF
O6S74pr9peg5x9aw5n7zdoyMR4dq3a2NIW/0MyKbCtx5sfg1n9EA5jDNp9cdZSgeAFsZvYqrx6mS
5kPKOLAZgQ584vU73/LW78uFqVn/P4HNFhiQyhHFFT2HTYulMRsYbiDT5PwtsnyT1KlnJIRnyXeM
JAE/n3zv+4sir9QxVrYh6BlLOV1ZRjsQrMxW8DSAODXGew5kxBA5QJ6+H4sYrUMUq3hHY2VbmQCz
t2QaAg0AxMs8VdELxXaxCRsvAHpqaG74nuu7xDiG8VedsSex8M4A8O8J8JD6sk7o9ci+j/yFwc5g
jf6wSBvQhWJ0qhWa8+jGMVpXoPppb4aWMTIPp7cNMAegaCEqESvgzsvcDYI7Jz6G4QadhoEPx0xB
zgMrAHpp2F6F3aseAilaBUc0HhxtKOPylmlw0gcrrD0YyQFtIa2v9Eb6lcD07fX4+IKBsHV8SzkC
cgmE7AOTkN/uoItHrGPiAKiRdHTJ1uaRloNbwooU4CsYfTni6P74ilwf2XgKxELyrpK43sd+2fYw
dV+H0HrJ2bwsvCiqFLk6U/y+ee0hyMvxYW+e37ohwasAnNvyXUqZfpE2trH8LUgoN93v1qD4/u1p
CoLO+7vb/G5ZPVoq+GDbJD02KZkHEU9Dkzd0YW0kkXiq2y/gsGN5bVa3plzEI6Zc4yS+4iy/FphI
erM+xvCMdMiiaroWgXpQANsvnhrZenu1JWujpTd1gmQ3SNwaVUct/zzgFr+AFhW23duiiKTfMF7b
bZv8vTun5FFliTkjLF5Z1xJyNvq78gRCnrP3gCTWlbu120ygTfjKP7OS3gOHjUiylxJxMqflHF6y
P28Jqq9GW/ViwDzWACATJ7j4NnflqsH4NUYsd/x1TxwXkIgm/26pdkZ8kiRfNUA+nBrxt8LIMkBV
Uo6R8QLVPRvgrnD59m4p16EdJ7F8ZwsWhyBka9eSdHii8v5MAKd16vWKY3z4gWvZ1e5si5RHmBGf
toSh0+M4nWVqHnYS0iID1iXPmhO5bn1Z7NhpQ24I2KqiyMZHWi1oQii+fMVfhyGe505Jx0Ie5owC
yLedhdCejP0rRZXHxFRbfCIUvFHsYvtBTazPQj6Tx4hOvkH5wMD4a9dPvI/06GxUV+igxDcDZmar
U3UyGAUZRHlTuqM/b8D3lq56mZ93aBxcvDUWrsgItI3QZZQrQViYJXDX8drJMxCgLD2T9sRr9+51
CndDlL8m5IeDZYjdUpKj32a1D837l6Zi4NskvE6D19gVuLabmHM8AUD9fkH9pQH6tIhYGCBASgi4
bW82LsAk6RXtYZAz3a2fnp9jN+a736sbnNvkaQR7sSkSzEsNNbm5xDlhGgo35B3EzmupQdnP1ueH
v3lEPdfjorKLcmUHfVq+G7trH7xKUv8okAY8DoNlyGgbbc6zWxT62O2YCwKYSDqsrDBPI2ChfF7+
PmSEEftk9G9GzbU8hOhtyMpgFFdQfUuQAOt74/gQOTRIjQ5bsDty09CPoSzPJajOMh/D7fhlCJKy
7Armnwhdri4gQ5pVO4MmQfWSZUr+MqWErslisoQKXop9BKr3J1qhPgPaLsdygHnPFgLSXoBY2vQ/
8ve2IeUtyyv4MFBY8JHoo4toFfsHuAyKi+l8h0opIelFeBGSLZN4yY1JKmOiATlyS3MpLRvV7zwV
Jp1fzoWBRVjGH1xTxoG7HPyW4CyMAdRiO1YFbvRhXKd3frDsn8ZYL5u6xk0QlseJIDDF8uo5mx9y
x9lmbJ4xfXkYxVAt3R6pcODsyM+L5GgftPVE9/G4TxMQcdo5p0DMUtzqFubEzZGPCH7lB4vlNq2I
+cqrEsyNFz/mclPTcGI4KvtPimYdIcdeTRFDvjclSXGmNU9ocPG4YCdVmC3zrYfsciKpnHyyxyEH
3hAo7VUGFr1uiE7NPcSMfHxEH5r53k9NwOsHQ87s0ROaCF8KFt8+6e36F8BLPdWhLthBTFWAkAuS
P0B3xpsPc0rDcVD3+E0f+vRdp13Y4/x1zy/egghsH3bj5c/qJ7GDi4vwGxq2YN3hGUOVzeszFIX3
QXW9XOqSRGS8lB8/Ml7OsPJNXEFmcIUSc5j4sZI+4W5Ekm5zcZGU4TKekKO/RUlpuVtfyZVJek9P
AlESfebV1mOFUqYJQstbOgNmMtckDQTIM/SwVtJpFfRzLlKPwNgb1uAy1EOGPp/SRx6uORz3nA7N
9m7d+cX0cqX5xkZqAIBTA2cILxx63Di6A3sj7XM+c+5OJo5HVzaGOgpiuK0VvOXXhe+PrlQeHmK3
3UzVF6a1HAboJAAWaB5xB/X/8gmYVbjZEmeSSb994l4St79EBHXVCK2XymmCdzQqEBdP1YcMtla6
XDN+CFYpbGfSi5FYHb+OPdXFoNzBRpcl9k3D+cM+No19IxrITYM+ZyZ6LGrtPDSn1LnFPuLWdSTd
6Eb0Eo/tst0PvyNToOnmS56HoojpxBujc0NB7zRhiV9ewQT+2MWHHoHVZuKr8WqlC6EDyQzvUokG
dswSLqE+DGc0yVoJw55W7qzFhx8RJC4B6xT6S5d9Kil6WgDszpugGQIF9QhRNZ0HtwkIG18foQ+H
Gk3Q97hP3ljWmqzKZXS8S4SdS1N69ZmIk8AuNcEg1HzsPHrDaJ7R+ETRPoYuJg1Zfjamz/a9PJjS
MDetvso11JLcDnd4+4APslJKNjLi35mI7Y5TU6b6MVks8mjEXfAAAGpdMiUUC6OI7a6shlC8WNtq
NK1qIO8bvbWYX8SC8Jmbkc8gIE2cF77hZMXl6y9ipySWinVXUaQkYaAo+94Q1cl+mrZ6+0fFbY7x
AYH0W8Nfu/9y5rszeZ1ZoBofF1h03WuV1tvP5SM9SApjeH1aJQVzE5K+3PIBYUzT3qbYqjrUuIBY
B8qlg/AOL/PIGHAuoB4xkwBrCSxmpfbfc5R9qAZj0AM+QEGQHhzUaxB6/AEoY0s6hjGA2fTHg3ju
59JYecfrnnAbe74X97D1FzpPMoBdb5z5/Ru0n1Zl/q/xjF5rQ7/JzCm+nK1BxHBNvC5Rt9fkoTAx
ikcYdToml+Bz35HZjFd8Vlf5OQOLskwU0l2G79BPBuXkAG7DPmk8/8QBDqatnHIfyTxKSeJJFh37
jK0nJQkz14nMXxemB+QAoafVu3YOCJz7EaRqrhAdBu9W5DLDKRMKfg2FT6BnZRp+RU5wOI8MLXlu
QVa9fgAM4ZTihM9WU1+6oO9qo0NDIYOpduk19rWqzQIGOf6zkublg1bMitUSqOcBqFRFt1u0MQGe
VfyEKcLuO9Mn2B5oaNyD1Li/y55jazF1cYojGpxDnGI528n59FmLy1OEAJZ+bb3Y76bJ647Q9lb9
iGuL50zLrpxeIZO8Df6VcIW9pSGoxQ9JBSJeSiCUR6ilJRGxXC0c18W0+XEbeGAHv1L4JShSeSEf
QknJzdEMCzSN4Qz730R6XwHn9qUxBynIjRFIW8KcYeGHdJjxv4GVM5om5pFYI0lbmfG3H3nRnYbU
PIQ64sSH6/y2Y+g0px7pu/1nGVtgZ/mYVMY+h24UXBbMHS4Y+YrLk/f9fb30n/1ICIzHpNUMdta0
X0RstGkNxgd6VbAVadkWGHyh/VhaJh8shN7P04oVHvmW4LYBWtbfeqNbT5BI4h+SR/pjZbCivppK
okm4w+NnJ/2XdIlSfC6kLIBpcB0lr2PlmuxQ6igRpDaB8//j3nkay+F5t0CoYvllZNJAwZ7ClzS2
40Ur2FCOzrUDp4Calye2QiltRIIqRj1dKn+9E34t1z5JFluqniHQW4Lhw+L1kHfcvx73WcQD2LdS
QYRKwO/6CYdGJaVML84VKIZbcoQ++0JT1ANyda8Sdln0tWr9omS8VGtlqEqGReadUTjh5HX/ce+h
gBi2Sw3Ll9Te9kiKa+3xpBJ5AZTGRHB8m8jkWEFJ3olNBoYI7rxEfu/cQHgxeYxsPHDBOmc9hIj7
WC2gSPol6HCvzwDY0n56jM5A69hAaGbF4Tu4D6k9MljZ5anyrLpGht71IiIejRVZqRHdzKrsDVNC
NGmmwhvxoBS/JiKn5wmTJ66iCOVqnm17PFJsMseACiAqlyPywzoWQW6f+dB4PglEIXE2O49GkJ8x
WydWCWmGVQkNvn0osVsVLfm0g5peCdQ1AoqP1urXhLm4wwQ/bYlAiNgenPi3kb62UGd1bHe9G7AR
bpyBvjdLYcOp67Szbl2xSbgbou8N2iEwkCYKr3fH4TlPyhZi03yQs99TJCcKLSipotYgjVN0p/Ix
c4OyCVv7OKwHrSWOqmLdyDzXjwkWzKxb67jft07pMbwBi2fwXZ5bOd1nKdP5k0NNupERcvdVALui
SNHQbukvKaon7vTRLeAjnt6e/2fHYz5xut280lg5fDtJJrhqUXrhfvRA5si0kp2GJFwSNfGV2xnB
PsE+IIGjLOSUvSsZe3DVTt2gvv71PnB17P4YspOPVdouOnSnfy6gIoxCuxsiZ0knkEtBEaQSXRvg
U6dc20UDpa6aT46RQk0ER6MKml91DLB9si6YlbXhy4AoIwHyjKbEIeNER0iH/lvM4mPR4l4pnVSq
q2DI1PrnWDqCzjrIXSIUkHfybyLCAbUcWkj4/FJasuoa74CeidItu5ZVzW9G0TuGnh6+Xg1iG6CB
ce0rgyY9C2Y4PWqllBvX+ssAFR7Nn7ettiK1UGvzo7efnebzkZuNFqRrehSzsmnQMPNWt625A4+3
99DA7x3veSG7R/UVb73zxxgI5KMQBXDcWW7EU3KfRWhWakc+PK8qbW+wowlwO7kwNQIyNs4cKBBf
4DLdz2qmv9GcPzhvPThjxkXXSNR5qnOpaLwN4XpMoS5mkHQydebL5B90H6YYvhuPHogV1QjuVtuW
9mABM14d3tVTZ9uDNbo0DLKOgoH5OHblHbH/mOxChiKQTdMRrJlr4JnpwO1fv01JKuQui1sq2iKG
xdDSVytrBqFKbHoFm3V/dG3p+RDAdxoMKUgGhGCGD5AHaKJC8LGWeafeYtlBKHA+HDpyEDmuXLg8
brQ+9rNZ7pSlA9x/cERipup33Zx22GSC1f/TCD8cwAqikDKQRiDgcFwGZzzioBoiIxy00Xn3QTYs
69oerqn+WczCdVk6c2f/ecwfjiqihudSwAplNEeTD3mBtHy5+se7i8IKyiU24V2Rw6hYJte+X/2x
M30pxRPxY4RmT+PoeqLFvnlPDnLQBMrZI1abrVLy3JBy2rq/FDYdR+NmBybB3TmofvYCaxOGcuKt
MlGXvfVvujau8k2NM3wTV2H4c+u4Wf9MuKmF6bGIaDFu6yDM8g+BGktpnK+vQUcXHJ/iQBGyQ5j5
v2dU2oMUgpWjf5emKzJBDWggl5CQyo44C+cEuY8hYAju97ritjN8++VSPs3UTa16Jd3NwzKqNQQB
W0hy9v4W8xstYsmJlMMROwNmU8QWzTfo91gyJO2E1YfQDbn1HM0NNq3C9KnP/rIp4lwFImrhEhYm
e+B0SMMSB7ajRJWuzkfiQAsGGUPovjd8oAnwQCi1wdqe7J6MyyPreq4ciWLuyvkYYQbhH6uAcN+W
zWbBHRgyJbdrnxioBWjXI3KQchosxqBy3r3gCgbw9jpOIgx7A8uqFDuSgNtXJtnmDuROV6JNpUYC
2A3c84Esik1TYy+XMVtzxVzHjpjMS9ELoLvd2pYBHMNw22oEUYyk57Jxf74PGhUIq2+Q2coJm99W
ezD56Az/wxTTl2K8aFTd81PeZ3nyKF8lkHTrlPsxfL1jhFuXZZBsVM6b3JaTwyVhGD1gf6qWzvVz
Z5mLyK+hpju2m/yJFkcj/73wX8JGJSNUl4ZN64pCFFNptIFGvnZrXxi7KlzJou+2iWFuKvzkz5GG
l+kZ8ian4ssDRMeZTB4gcijjXNEAPSWTmGqaD/hLn4EF0PfiqHz3crCDK7xrcbyU6WCqAp3ETJ6s
t7M/MYIXI/P2FV08fMNK38ZOO260r6wWSTg+OvMvB5VhLZ6MOUKfVV3QoZa7KbNGLhYqRiLiNPdh
0cdsmVQg5KjPb8Gk2p2riv1/W4ET363J6V0SqGqOI2wcCdyhAVOcLB1Xk0inI3yrw+RhPGkyVMYa
JoilDtAcnBaLaRMvD/plqu6w5KnIm3ZuW13a9l8dbH/u4s/JV7oJ9EEMjCBmr7IAKsUxo3LyUguA
uj9EbZj7Rzv04kY0lVbhh5ahATsCwAU4SC8CcF2g0NJH1JosVWV+zjUrZm1XKAtdEXvv9aAeYurf
MIAGKbJUZiCRiSl+AF2O94wsvfeupu1IHMT4YFtrWB0laI1on5RoR8RA6HXuWZzdIP80VLK/BOIy
E3BhHHFecT2P0JhjalyCMGYWQv2nXOrOqW4uFGnln0NJnkwLELqxeYjqOMldqSKqQmItN7GBNYZq
JR4GrF3UPAsDvVG//DYj2+7DM196yzrpIEvXFrfPrH9b7/gQBDDgwfPntLgEHFKBMlM/h6TjltTw
TrZ0/FqsaEfIAGYI3S5U1Fn5FywqSgCxm/ChnuYhgxdFcV6UTFZHnokpRd6BFlWu8YTS9G/8vnu3
t3STPSU5ftHPC/ypZNc/YXUxtSomvIReuWf6VwfSnzvH356LybLcXW0lRzRGSBY/mbNlusO3EST4
vKbSyqTeyX1avVEEoTkcBydapdTkXWpIsxsWz1kLNKZ09XIwISz4T120u1UQGEKlpegxio9CgMYR
ne9mRswXJBioE4c9VkdLsB0og3o3crHOPsKJcMVBeAw/zZGMixjq7rKn0ZRgn1MLzyzpb34qqbGX
xD/nwBC0rQxdBRyk1yOx/IfrOckfp3cdV58EZBZkgfTcisBsaZdZkQPU5X3gQma/odkz6SRFJ6CQ
3fwWu2Jm6sXwBtcKo7r28JBahkz8F1/PaseAf0K/vEzVxMFcz3Nf+j8VprlAmNUH25//hVtmKElh
yTxwSaeYjWlU1kwtwxVPtuWBVv39Jgd4a6Kdrgjpyl7zmdkVAz4cmJbWRGvlgfSAnhxyoreo3Zj7
wwjp20OtANqKotUyGjz9fX1UQQtG4nppuZ9od1BZ44uB0bI3tSfI4AnqeUI8Bf/EYiD9FeH6Wczz
qe4TddQQdN/3aIgwEai6XSF6OXeQ3FkmHP6+7sBgjoJVt5MBBvLPsW10l4Lnek6BFF1BK/Mz7Tz2
lOaD5sldwdrBQBenC+oB2PTdZK/YQuxLcMHtiuMXZPPbAJ3vRZUhSZ840UvFORz2d7adFf4pVWUS
ORGnbuqVuFdPThcYwzJTnW7dBnktTunmIqALI3qkcG9lK8awKU4Hy4tmMTa7U1OoOjIXqb3T1XqH
hL09+k22oePXz0Z2QgIdrgMcUMudo3No2yeWEVTpinm0pfPowf40pgzBHLGwt1CaHV28NLNdbYos
RMJlUH9qF33BHLbGZiTo/+63OOxgmljlfTVsG+aki8IrQ5/vrRJkizWCkCLMn6DWZcLi2RXYJeuv
FBf+EgEXw5xoTQN7bTlM1PVwsmjz1cIbHR5OhkJK00b645UMv11005a3AE5F39RImwVQNF8XGCg6
YuXNz/L7i0nWmtZou9W+xG1e3D0ENnAE907yGTKBGcSJz43mUhZEbjkQv5tPf2zfQAkJM1ynE1nc
IxWfczgBYLd2vvEG/Pbwv+NwO/z3kbSeOnjwYY/8kCBiB+B1gdIA84paMOd8t3FgT7dKjVXAD0SG
j/WG/UQ4AEjFjalplHDlTLZKzJabbc5ztED+E7XgAHusmCahiLe5diM2bD9EliSMZA9CPbqM6wwG
//tgehe7kFiRl9uYymNwf0gStG+D85hRzMP1MGNRACPje82RmG8WUFZiRZCgylmBGmNIiwaVvB+K
bK0yr3eqGixUhEgfMr9pJXBCBdAgo9Yp8Hzi0RPeI4HfnpX8wV8sDBv3aw+O6wbPJOUia4t2S5RF
x0aeM4sfnccGweJYbtPU/LClhTQvj0Ke1xi48Z9J5fYLgo9d/K90sI6GsRIN05gaRiP8rQELBDIn
00N8klA9LZduE9rTJd6Y5UzupEMhe3C6MmMtPJyCqv64kJkWaQZWdXqZPg8jYvpGQlmtRDMm918S
fi5U29oV2QUkAO9hgbZKD80Y6ibxZF3BI9Rewl7Icc4/AURK/EK2cifFmBpYbnlzFCWImJZgNdTi
ho6U8Cl7aqdaVrsLPnu2Mu4Jm2rcgMu/4gYjV2DXutQgkGrK2vsdPL40NA6cOmqQTTk/AknobrEk
mKg3uI1DfawKxAbePmAnaJGrhMbRJnsu78FtmOc3XhuE+KBjYAJIn0n5pzXrpgU3YTtHWgKSWYei
UggVaJJu+7aUAtLiGCQ3c7pjhMLfr40OlwM2SvEv8I71Wntibr0J7sety7LzB0s7jtNpQ4r2427S
iyaOww5b2Ny5QVnttC6TY2DBGBjzGVaHQ+06FDvokQv5Higt5lEDkBL2GGzcAMAPp3W8g3rI4ao6
9uYO2BbZI1BuLHOoGa3ndCaMKbrOanRjP8ms1T51aIMH5Z2K9psh4/BCYPBpqkFypSqNn4Jx8LHY
+7qIx/x2kGu5/FGDGzlmv5GZvE8ZAyakjwHZHxTQy4aK2aO4DF8WC/lfjgqKR5wemxPOG4deOmg5
frhHOBFo5Rnyrg1TSuAsMJqZDb8N6C6OukkReAvOlThFJ9/SEdhHV+XJ6AiirFZF7vh78zZeSBRn
JomhiTt3jTlWx8LKamgVyGwTJJYwym48qJPbmOLm7gRTfgQ+hH40+YW0AttVTUExzzc9jgogUPCE
6qwYDbSmYs0zokWtCiN2WgZs7XpaoMLHTHX6WxTu+NP7xVOP8LWUeG4KeICuCyOuAn+RL3TVCkr6
rs6Yeifuq7ooC1m04wEE/6sRmX6BxIbx9qHlqTgkJ+7Yt2826SzQE0ZjncoaPNLV2GQf0ubrJdsH
IDMYxg+wwkdDnMLpAY0bHdILhYQWu02eAu0zs+DS1EDyRxicda+6hDR5OKly/baD0jAuXo3rVJhj
KTwsDQTFQdJmBOzfa+O+cefz+3ajl2uJRboZIBp8M/50rYPWCBDTGIclKhmAsfMuGX2+0LVaJAd2
fLK+Yapit/Bh115Y+cZb5UH885W4ikOEr93xD0wGDFN3HuZV7C185SuUdjhLBdPXh+aGexgPUEZv
AYA8PYvShfwUmZx78bNGIZ4GjYlonN28JooCx9GrWDPm3+WVhad1NBMJylkQMaLMfsSOPJV6kk+w
RoxRYw77Ps5BATgiRairEBcDy/s5Ncz+KKAvqA63xS9qM9Mxvo3Z+zE8tvagkJovqLZqROHZGxbQ
XfmKVwYOI2IIrhie+bxd3jKVZ7M4oP8FkmNE+7tftmsG9RoY1mGFRX+v4Wl2YCyOcrxucIaYJrhV
cFc2UElOzm4xQ5PU/h6kS6mvxc55991cnKE7m7NB2A3JZaGfq/oS9S9Q+tUwy0XpVkCLWIGWzuvz
60Y8Ye0Es4Sq32UMeDVzr3CVCmNdJ0oWLBCuOcAyAhGQCJFwKvyII7qPldUSKIcLP/465dZrnyug
vBJwLYR0+wtW2nsbB7gnpMzvv5jX3As8Q3I0n1lTYR3h7g6zfliUBG/5ADucRYKZ/mt7nWX/c27s
8febiPHLCuhW9gZScxIuqjUztP2A84NeYM6MTVTwIa+2hH67TcNxxCfj7DLrryan0HhlbIN+AOoY
Ru5y3t/Ds25b0X4wV+lXqd7Sdsp1GN4UvA61l1UHBHECGndRfPRdDwnusx+WPb7M+JWIvSoTuCtv
i/WkTqd/YPs2uK2djINjXx+uzX3PsUgxrDfK7RwYP3qG6e1pUcp7gaFmAd+oi2pO0Gu0x0he4+Zp
+Vcs4T1QjPlGfxN8dqQto/F6f5VeIVrgZaM+fhZBk+6d65ccshzOZqyIelVHCABRtypUHoIO0nrP
axWKIT/tGqMSvDnFQ2AnNi/xrtBMsNVWD13AKj0eB84vWhxYJKM+NltsoVMjN/BFz2/8oQ0wcOIg
gswhfikutafSxFsU7QOtPkdWNCab56ogHxW0h9ySj8aM2qiTN9MGBLIVykTE22wVytyaKim/6As5
gc4lnda1prGH4CFyDZzm2eBdvplpLZK70cbEiJPSL2LzHkjJXoGHpAd7Ea6fWXShoVsijyC4F9t3
wkfJlF2J4/LvrAiHpRsNZI1YPlMMkhpTaokbT4ZBjz2H5tSmoM3Wdltr+KVAteHhnDjInKN9GPag
CddvOfpzJDe8MPwt4QHWXidcHvgjITsBWeygckF3LVoq3DNmQMaO4a7ymrE7bb+4hd7QZMxm5lXv
aUu55hjomO6VluB71Ub3zBj9L4wc+6BblP+d0bOgWzj82icm6LNeXe6rQqn+pTQihfAZ1d6YWlBZ
P4qwicClokxx0gXM0q71ZFargz9k06hrGe0/x1PGjYn2k4ulZz0pLrU+JL0lUcJIkqnuQREdOuYB
cJ2JAFeujmI9wotXXQAR4eJOwOvjQ9/ax3gby0HjHorQaRqTLsDFoemtnmU92Gt217ZZmUV3OGOQ
Ycw4Qw5zuMy5xZv+m56EMO2YJ8WNXyJmc6NEMDjdimEUZC0Puh+Fo7XklQicP5zqqEeHCgfq82/2
WBTn5DPIqj7Su12FWcMuOO4cMGmMe3a6Q8JSbtVcuOootlVhpBHC84Gsc5h11m0tg0e7/rf4YAcj
fqZg7LwJNAeHQTmlToGqQKhF0i4cA82hgPiSA3hZeKx3HPvcNabq5y7uxsTRY06B+sBrKaIaXECM
+U0toNU3SviKM2CwMkU/997hw+5IpWjq+GSW8WvDtp2vBwOWYG6c5mLRPA8L8QI7L9fBA1VXqPg1
e6kV8WIepDxpHRNFBtUjQNzqQWH2DpYF+RMbTkAQta9ULoWFtdr64NjML7R27PvWi6MeybpN2YvR
8iBgTDFZoIwA6EhGiF4fTZYY9BPG7zaSPKoO/MAPZ+4USNpdSCg9S3iP89sPTY1BlMYIfQ0wodHE
DnrMhsi1V6f2Rk4VjfGVIT8RS1KOF966QXHLv9VV2yn9v+oickBf9ehsTenOGqM4ioUjx//YH9yC
PBUSfKDG45zRqYO0+TI48c5FxhNxvdA6j4/abO+Hf6SxD/vW05HS9kJqMvtgWI32Z4eLiqqUoXaM
x4CXyqD2MACES3d7iFE8Al7CN3RnO0sxO849gPVNhSMLq1JZxy/qgQ01upaGUiP1EzG5m9AnKQLD
AsMhvo4iTK22GRBnQp9RxsHhxV0xB8V2+t2Vg8nlT9VhPlrgMAshDhyuoaIA8iYJ+ElRRCdnjVhQ
VFQbmiPYmdVCLBc/pRDcEAyImUnB8OzZsipD15+c9Sho3NENECioBragWReU3FQc6XO30DQNvI+s
m6xmtiMFp5ut9g8FXgKIBmRMsIfGJsZMLRnn4UD+/LHtAM9pbKSS9FYCL7WCr5E5JWxEBDdalA8P
LaITQDozGZA4IRRwimKjAOE5EE0Xaf5ApNRnanual+8Z3v7tQ/Ym448eqoW9DOGlGrUHkIbfxL5q
grlgdxxPz0DHmsKPazBUv2+XUKhO/aJsCj+53a3uW5s9T1VGQlnTpxT/xcUOYjVpT5PPqI93cXY/
nPloc5M4TrHiBqG7PJROjrzGCXmQfKaOV92/ykUhm83QenMU8W7JtYSAmxjUxpYE83Uf/oo7XWEt
rcCGErqiHqle1mtWsrXsZaG+NFAkLzwcV4SPbde5EHqmez2O6ggViOL6zPZazyj3JAeG3Tf8xGJO
vNK3MpYUaeJ3TLDu9OBWZjmqOlUBkkMdnIP03YX8eN/Nl9SmbufuwnvyQnQxGIq1C+LXzqt1abZX
td3EO5Dp6vTAzNHyhzI/QaUZ/iUZeEpyM5bZHaKeRqLYPQ/YzZPn7PIzz7UxXy8ijZ5wmtIv1v38
hMeQt8jBTrumg7VzG4cl31MQmXKWm/vPG5abFJ+Kd/5eCJKAC+VUhRzMMJyei19hgzUr2/P0kZSV
9QS0gMWsSaLEneZwBH6JB1OwMFerAmpK5v8zRAGExVKsmpycXbHIchWzlSGI72Vf5pBlE2fOvx05
MG7lSqOGW2cqpuT5FMHEbwaUYgQVypuJgr50GbACWgsS93sQiMCVF6z2CVWS9Us73EsVyMAUlNYF
U7MhwurtngQBt6S+AiPwUgXs2vrCAS5RltF1CfDHeTMRbvEd7qhbXHs0Pb55UZbT+noKBB10mPPj
17Olvc0/wAZBBbgopySE8JjlUT7ay0z96aBxmVOpI9aQHo4+3mm5PxS5KASkbFNL5508gABR5NlJ
4uNdMHbjasB6qxboW/ZhpV7EjljQ4yf4jyd0BlVR3h4/J8g4Y/NCA6i+uvZXdIEmmakmTMmv/oao
Y8BIQCVZQxHT4FtJrJvYK4mmi+9CfktM3EoA5lk/XTd0v5lnXHB2AEiUIV3Ca1GgUwJfzSArO/uW
JwNpZXWlsqZvUrjF04OxabiPwO8LJSb6CHoWbIvC+8EvNf8zqyYoYS7hmIbnRq9Cvr3mbucxqxnP
xIzzv8vtzWKvS/1+aNqMzaNuB4BXutf3wbD0w6i0Q1//IjWx84foeSVcz3MUtFjhd1yv4KquJ5DM
dC6qo5AXMKQrx/xNqdIZEy3y+W4V3xoR47huxQipswRD1qBovYV5Iv6iLuPNGlmTxNMnwyL0shaH
/jzN+X+NlTOqQ9gsRr4lEGlOoJ/EwodBKgS0ZP/wIE6AUkKpNwVVzGUrLWzQQ6E68qu3/UEWuxaG
DcINOF7wqRp6o94oNjUCF8WpABtlxzmV7MCdbXNT16uQnTcCUBJO7gnGTH0IweJS5nOuY+bpIji/
li8FGXVqHRQmirsAkczrbO+dRnOiYDwZVyz9TpbBk6QZWwEFhFmB9LsJOU31TvYKOleW3iyCmIfj
JkQYsilZeEhr7tV9fZ1Ov5DdEHSd1TLH1VE5XONxYLvX7qCuiu+BuXUXQIhfS/QMYGirwmpJbAR8
OHfrXdGm6nqtOWjZJSEnfWAChADqwvVa0Ls5rX7NfCIRZvrO+bkKFjCTLroN8HarTWcoTcikyWau
oLqC9SXPKtDUzQ179lQ7ldOUTq6ax5h7y95qefcb+Ha3GL3krwINuIR64OxPD6rU8f33M/ctdaGl
I2osJqiwHy7Lpu9sIY/KWjixiwzs0JnC3T6ggMTcdNdwZ7b+1bCh9xNkFl9pP67AnTDBtnfxYHGf
rMD20+Xh4FchBJcgmUJT4ERL4j2yHtAxuct8AjdwuKO3XdeuzjrqlWwU1aTLbjFvuUeMuOK8arJk
PnUq6svKgDuUeZqSbBQmw4/oAu+A9GK5Er0tc1b12YDDbO2nRtDVVZIo1j0i2oCdtKw+QArs3CjH
V0vOhS1v1VwIEqKiV3WHzOEsSzpGKxhAnRqRcQyhTFQgXxbntVWiHfYv0Pe4+VzDPyybTmQu/N1Z
LO6YAvkDBQCqj6ATD4ueLJXZpag9slmLux2xkE8LkmOYd/Zk8l6Oe/Z7uvYvT6fB0VPyQVAbvClA
eDChbVtODrxvVG/1kPFnjawuNIKlhLIG0IpnnJ2vrFTHZmFn2RADyGNBoxrxZUSipxAabzTeTcjm
8+GBBlUVq5S6lVzNT1ZxIXj05EEm1HAfwWd4ZtSaTo5p4nWk5LszhAmk3ClhVSg02oJM552RRfws
Lig9oZN5RuO+LggeaaJ5JG0xJbRPZYCJxa/f/numAq2R/geXvNhLlzlQuGlrq+CgJJT2uj7//1kh
2SNyQyjRiCl8yPPggwZdY7B7HgWfsjNdQRe7WyKik8/o9X54iETAwehL/wX5rI0c+nnuLUz0PChP
acQE2MWoR0yNBwRJKSzyFz3Kqvf9JaggCQZW5PNMbsdDRTsq04g2Uw3Fi6TDtBTiRP0wtMq/hUA+
fcQvpiZaP5Y6SPjriZ3DiUlr8/oiRQYfP2bQPtXTt2adMqDEUDiHHEql3uFZvp9FFCnaVA0BDSGE
dZ14a9ctO04NMSe4n6hO8vit7FkJgQAc7LqlwSWUpemJNUoXA8jzi+wxBVQwuwZKS/7H8NI0jDQe
91O+MDc4So0h5Pog9/0aqv6hJiUxdZBhrKEw0Wb7IuhhZ9lkM2s5xbiLfUiKiFGSCyNrLD6hT+7T
8kAWQwQKIvRXiM79JcZLa6zqqi0wVH7u1OHZ5pkeF5GsL1IyF9ueUpOuvR5m9reCF6Sd8Ca2Shyn
iC5dXy0Y9aAWRGgdWWWsb3kNJ7eY3gXPd26rp9FFDRUnsgKa81x6Nra3Tn52W5XY2ravz6Kp+38G
B42KsJMeY3+0P6/xGHXquxt/G/LHW6Lr1aSqdLG+NcxlYMhMw6Eh9KHeDyGbi507D8TAFUB+kox0
530GCWIKnsDo9ZZS1CjDhkzks5Tc/jgcrCny1d0ICvJbX2BBq7rEZ3W37yQSLMmtpELMmzEyinRJ
wyqL8gX5h76FrSayJ975lgeX8hI+zxV24UH8K2L3OQvos5ljYLjxfw2SoVuhga3RFlgCFGBTwRV6
nDm2M2zNPy27S9N4guZHeZMkjYR9ypUgmtQ6Te5mR/hRSLRjirD9r0UwGTfV2J+vjP+YUk0Laj5t
OzKLjKZBbN4okuyniNUubD/c0FRcOPVcC1buMd/LqbHsDqaY91pKgYTDFz5H2yaetAz8gjCTO1sV
uS2Bdyl6due8FlkKHwPM9yv19/Hf9ygm6B1y3JUJ/evyK5QZ75fczwhDpnEvSS0aD9IIohLHT5oz
MNkJHtcJmhxQZXZ/izOBUjDk8XUtQx0orWoksdahJqT9cacXJTuz/ayfHLdVbcy+Io26qOxFWwJW
dTQQTmCr27GpJ8eEFzjTtrPLtNHJc/Lz5uDzVE98yiKcXtUM4yqTiOQAPCADbrWX56rxoZA13dtN
gcFBKitxQnbAtuEm1Bg3tnAHCggJGESKee+07Y0Ev6SL4ez6kppHBMcCb/UGJHGf1DqYjDR1rmse
PC31T/ypUEPAZn7eXLscR+aWDbGo1yRC+78QNt003lmzohr6H1rNyLgIIGdVMGboa2KAbhRYHAXL
1il9T9ynNBFEb8yHLLJzfQpxJDQna0HA+6a2mgpHtNqDAgkmnw01Pw75kWsNHAT6LOeU1oy56ZsL
K3vZkp3J8HvODH9IXn9fwQ0GRERU2+VZWAlya8mMMAGC/JDQorEEppSw7/mA+j9M5eW4iAo+kAO5
KCTOBK1Mba5vZeGU0yAZxr+2aIlavJOGW4ogIL4eu0YmjW5RCy5ZMoLgt9kxlfd1E0lhsm6h60gF
3KI04rBd1rW8uszq9+oBo09xeJAsMoLxYU6rP7y+wsC/K8EA0JCl3sDTmZZd9qIkEHHHTqkc8fnT
8NJKCptwfJS5czE4fJuoHm60IWVIo2oxTFdoHRvDodfEpkURccSC09t2SnmOwSKB/c1Zx2yYOCOG
sdg8XqPaqPOIG5usNwvj/CxdOD0XARxvS2ER6YLAOEMVRMuTP5WFGtUMPMQ7eEMgBjH9H7ZINLkf
neNTtOl4j2/pMrLCxkco4Ia3dlwOiof7f9cxEAhyCs8/Yor+QganbqKMG7UPOtb0pbigX4GrCtIm
3yh+pciUcrgXW836QoeGwO62+2RIyCJ0roPzY0kzLw8HcksN1fY1q4sWJBYmyS9f96+xd6oOf5mm
8IdZp98SBVmtsMSDwbw8gxWMu4qB+cqNcaJqbfL1qI6nFNv2p9B/qduv8mg3fJbS6ZrGrj3Ys6aJ
M8ruVOA7zJqt6ccxmJXlrWD43DXSb5ZwEtms7yCcwqEXCMxz+HT4aeOGSASRqgzK0DcrqVtlaE2a
I7MAlRgoMg5lZW9XnS+Hm9pYyg6LCLFIICGElbcQAPTfG5urk42aA8TDOFfx4QVVhUUKOzHnFPU9
LrjSA62v9/Cf/1/dUvNMM8kvckcTwY6NqymbCZI8Q66Ykl2+dVQmTZ+rOj6jryv+q3VKbOHHrFyu
OXZJt9N7krw9uMoiE8q29rbffYIsKOV1vb26Ul0zilMvp5t3DWDtj+uKoh/kn3cPzplO+SB5Fxmr
MHhorY5RpIjfpEumT9WFdq9rnPZlFwl/U9Rp0IHT5fbiUpfwImD+kfqEStmTaUkel8M+RPiAAURf
Y2F7mjOr4C1geZlaTtbWu2OWJbPpuTSkcndEbbreURmBaubJPZd7v49nuRcKEfaOLenfCKQqdOV1
H2ZGaEEzvKP7KmVs9EsrLsxWMfE/KzMe19T3MAzCkAV8z8eN43bDNN0lJ700A6ueka/8xuFD9xaD
TPr3wEb0GWESwI/e3VCqtYCfyXPp0zcQ38gLe1lHM8nCQZBhsPEelX7+Cm1hyIU9KiiwlEJY/7Sm
OZNCisi6kqzQz0KjfCfS/k1FZ1Gfo5InHQG9dy8hp0UV47SxpLYx3/iv2L+Od8V+SXzZ/wzvzrJw
b/d5D+jrIPqLF8NT7sI03LmFkILOm8THHjIWIK5vn7keb1uiLE9dRC/u4pGcBGC+iM3sFDGXYbNd
nQ/nq4t0Xu5C8ZWixRLBWQxSqa/APFGquQWEx4CAqG4MWNBKKA69SykmXFRit5w+X5hCaJ0Adr0w
bnNIeXg2k7QhvRjfto26NK8FuFL0fT7MHuEg/WFaQhfuiRNdGD8ZndYCnwuTYZI8vNmjf9ETtVJC
6bKHQ8AP97Dke9BjcQLkrXCMrj4gYdEQd1o+WnhpGg/4NSZebin6VgnGkvFekmNmy+h5+YgjQlbm
2Iz2jIWnX9+f1OUZWmEts4f/PrWDcGpeDHfOEekUfd9lrEYeH0W6ah1sn7pIm0yi0OzVheWacdzR
UD2yLGfyZqYBCeCoYyaq8CFECe2wyRXWnEVRRukce1/sTG5gTlywgRjRcLyGL0YSYl0fcDv956Iy
QgVHwqEXMj91xa3PKLC9D/7wfwXYAW/0xyaFBVp4NaNoLvTWpqZHtyqGta7wSUGoLgTbfCS+TRyO
fuosjYC7eXReqifoey3LmhTBdJK2NlBaa79Nnx7aKHHZrViFMCNhHp8sgdKTZR9ddSWgqL7C/VCJ
/UvWen4v5vtOI1MFigUjwKbW73l6NppT1cI/PCMPKETdOznAwCYFKpcUryvoTPa7Txlf09sVzp9Q
YCU83IqEH73jK0thG4K3y35VTGPRSml+qZga2wh+maHQTUheex14qq8s3Qog6dXM82jxhCWJwSwI
CwyRtF8LtYinC2K1/YzDlQFy8QEfpjCfaBhEpYDXQf/7WqSX99+Uoty70SnxZ1glme6/wYOE7/yS
uSnFxLtbPXwJV9PWofN8ws1p6a+ZJ1vbQ5q62ZGuFHTAvjJ7wWTUEiWEOAX2E7ghm7tXkdAblcA4
6ihodVS7Ky4wlpDcnZC89A3GDE1WqKJ23Q5ZaNuV4KgU56chjE6e6vkoIdQyKAv/OThcGcP2/FRW
vh4to1O3PLoqvwMFldVyM+Rz/nHOwAGFzYx2rOxciXgVaeFKkUxWqusLQk+g/tU4V4WOyk45r4mJ
EDNQiFXiXWfUc99Y511ub08tDC9K8tyPWeofT3xSXHedQmnhpaSbdKw1fPiwJfXHa9KUdXFwGopY
7ewr49l7gHe1eae4PXZTAl452fz6M3N6gXcClckmY3LHGOy13U5cXp7yyb9+IovKCIO+fnlvynhA
fdua+TSpRGm2dOt1IH4e3xU2Flm9zznDN1RFmcrAtJJKv8EYStKWf/+XeCiieOzo7LEstsI+otOu
z8DVsQVWwUcrEMvq7Hfp2vyjT697jYX8y75DlBKQd33WOj0l5vJVqNPkF3eaAiKrP8+sgiwaqhm7
wX2H2u1sZiQdbpDNRfUyAOrzjLyMZ3VVGlS9Nt+91RoFsEWyfaqYayiZ2m1yMjQM8jo55tRngODp
khjDhqX2XzyQ5olj8veN93lGPSgnvIgfVInsjbB8aLyExRIFZbKy1AJL0KAhf3DrXE5j1vE+62Mk
6gzcQz3DUFGtKSlk173iZvEX39zBVVy9sjKeCW4JU07GuHZRzFOHigCqitYxmpaZPrBXfFnJ58VZ
XlDqP9SU8sC99qDHp44RnXSDVGqZp5vs4om1beQNF/6Orexagw9JAWc6ComaVd0Vqvf76/AFBEXN
l+x7TwWp/CTpG0Kz9Dn3/FcH0FiXQ78XJ7rpHyad1Dwdoy9aKxM0kSNGSMmvAP7l2Kifdhu+9HZT
lpFn2kblvGTHM8JNCqdRHTgTBISv/Z/RIZHu6o+akCZlEBjVct/NaxSIFzOemxL40mnv2KyEWKTb
qKOqzXsQ7TIain/q3SrO/bzLhUlO1PCUMdUCIjq4JSC1HCuUXuWpY+VcvCBQsFizjOH5GM6Uivbj
OxotURmDX3NHCcz+72Q93RInQtS6zmP5q1roRn4c2HNTvyTYfHoIXXk+6Ck2siWflN/W9f4BM8sy
Aey9fwXyAYZzWOEEQFea8uNz5/gJemor5LUzOgv68ZJi2SXRp0+I8sF+T+b4tMtqq7RpM/lNwSBr
ijYNjdjFPLshdg4ELwqIpDc5fKaW+R3dpv2Av+3H/A4/2XS+nWJcQ/QTl018RNfKklHlQzD8fcGz
2N8P4iFMxYpCNEYPPGqTUqNV1p/dicuOVCxoXPkeoznJiBKjV0DW/6FlDbO0kLuopX4AScxAYOc2
fsOPdIpmSltTaH6DH105TVzPkerzlihG6Af1+4EHKIbXWK6k/RgxiKZvqgiMHiQUL5q9lfyvJYgw
0iqF9FpgJdacnTy/LZHKORlcPIa1YFOWERy0Qvf/25mq3VHegTLu5fCsLhzYQgHlFIUeOoShxDev
7IHnBpAy/a6z9Z6JLa0sXvuYcfjW2VjEEJyLUBU+p4JcQbKN+1oWneDVAcsOO68ICd9h8Rs5CJhB
064enLN3B1lCTDVWeIKqMZw/p5poJH4QkgbCUQJuN0jsP00HMlZzoBxkNgR/Y3q7h96dix/U10KZ
IqOgQTI+DAIuK9/Kr3wEGewwrvVbRELuySZVNFNtHnoOiTIddgeaR8B1SEukfmcekVfFWg+T+qHs
ODRrWiz0NV3aCbzfSdAVBDseqiYRjpCfUmkTMd6G1fie3tWRnmzFE8l8iJDwy+Uh1EWVg6BvJpef
XgiLieFXXUn2TVGiWeh/A4KrIESiK2a7nUlG+QLKDFj3pTpp1fBwWIDyEBrOjuwwXn5sM+YT7yDm
7I8BIxJ52m7a5N5u9aA0/PP1xfMdRmtEWNifs7WZiMw6MgCCjMQUkYLzrh5PxhrzZSOZv2eyuUMG
xy6YM6TfajrkVC0Cdlzv1asMiei34EprEoWK3LJ0Bs1gEd/b50Vr9j4MDC9zQkpgnq4B1yHiKKjR
83A2k+Ed1ovKmUgpw/x4csc9Zlo0ZW10hlgEkF90YccLgag6K2MENLYvgurAhIi2cTR5bq+2mctG
lprr/kAG3OQhCzVh6KLkoQ906RVj2s7UjPrmoHW9rSOSzikaetwC7Ors9AAosMDly6JJ7HWlv3LQ
Lh/T3JDpSl5QQPlIIuuTDeEEnWcGrXWFI0FrA+8tEoG66MKAdHnCosUa0D7QBAY3xMNRq78n3NIc
l2FftXz565OPCE0uunF6iph1pN3udD/b2kEMAsxHrOmncgbiJtN2FKOG7Qgn5f5FAJ4K50ZgH+vk
qrfCGuzAloDFu9J6YqFSXl84Q2mXuR3A9zTZvmqjBfP1PecV+zcc259bfxo5/Fpjg1ISkevcDya4
W7NMTvXj5Dqbrp9P+Fq4Zwgq2KH9mlWHRmb2exfKoMeQmqvHG6w4oUUrmvmlMSP8QothoFLOGGRr
pRimfTcXLrsWXIzrsmG0DEc976XyN7m+h3n95tUoFYdm0yyxdNuG+FxHsKnVmQI+9Oq7dZJtwrwq
HlbUF5tpRcbihK6tvCSVjg7itauJHLo8Z/68Wv3d5IbNLnp/t8Rw/vtV14UGKJ5qsln8LsGwRggy
Zkc4gRGvQaIay94JZ7vbpayLi9MiHtla+0JuXh/gsfDhwN4nJ1eZLPel7cstyfmzm27otxwHm/Jy
NgXu+C/phvG3YfHpJ3Puk6VjbStrYgNnAACFidcDwB9ZngMNkxO412n+YaP0567AYDmTyEmUaRsi
nmaeTQry9R8QILPCgywbNsqSliQ582D8B+ckRqSnqZEGLaL8XNfb00KzvtdXxFMUwnl9X6MI8c6o
cij+eVdGmvjjr61AmL2YK6bkpemqk0OGPP2ICu5k9/WQ9p71MC82PDfX7QpN0wUnqHjZLsQG1nIR
0gTSEhE3ldXJ9GFqYI94zPv3sjptZr7X01fCrZOFhV0QX2YJ0dJ1xIkrnPDiNZjOa86VTNMwJFn9
DtVdhto51IsJg3oNitG3D9GxQparRNP8hxzJtvZzm9Fy7h3XdafGVQ+7fsMSG1DLRnBGfLHpXPzE
dA11HxvFnuHZ0UijzeQkcW0PjBTaB34m8R4HLPZcnETxD9d3f/qsVXwG0CNNWqY2lHg+zW5zLHMX
IrCJGMqrTVQlUyVZ1h0FAX3ulk8A4DA6ibWc7VA7RVrIoX7zw4N2O2YrTxztAf7OcOllIuV2hxAl
1gLdNFSq8Y2Y9MuLJ/CG+ULZMW9trhYqK5lTNhxxWk+zyTcK+I8jHqYsAwdDdxMj0PFJWyv+ePsK
nub5rzsw3BUd74W7V+CbjuRHfbr0/UoZ8vY28zs5XamDk5u8ufBKhQQRnG+aw9uJ49ZqqXLB+w/P
YJ7v+MXssTfHVGI6UA4zqJWvKkWReEPa6uBrR1T/gt5VklgCyX3Sf8IVFt2PGQTHi74qi3riWR++
b1RiXoFV+PpmEzYm5GPxVPNbUYoZ1aSfUvb5jeN0YSumFqCDvJP8o55jlltJRG2sSx5OWA2f1m/A
N+j2EvkVvKVHqxytCyUjHb4RBug5GVbtB+OixKfyddAVmOLtRO4Rav8fw5pGTtO6iPK6s+mWHp8Z
XoP3YqEctC+5IUSxYBOMUiWmj0QkZHYL3Xm+pLcvf8/VFS2+bpoMigUWEcUfOFwiWYvt/k3vzvJy
clh2AFJe44qlBpdJYeB+i64DjmlW+W8vIYgtHKxVAL4ag/eIxKranF2ZNezRqCAmseqhhhgm256w
Gs3Ld07o7WOs5XArdFuHc6GR5IYr6lR4cGSXHeA4u0006yI2rumNccGMJcUdMijuYSeSyrmhA3F/
x/sMlNclyoyFtV8Fe84DoeeWVR4o4Jgc1iHcwJJMnO4qoG3LWvc/IsbvL3noJKZr0m2VYj+s+wCv
tnuE0OwQGRLlWCC02ZirM5WTEbjn4nVY08QGQAWf273vwf0+bww8djhhLqHrlDQEdSUOa/WOjWsE
DHlWWNZ6AH53cyU04ILvkkRu8wyLN8sPX1flW+l4mWcFln2WFst3viJNAu6gUs2V4unNZSH6R+1H
eS9ZWkjRyl1Ujct4o7M5MYqm88Td2waENdJDbSOEOqrRt1TAsrs2hM5wS2GbZ+NICLKwOA2sIedC
V3hNaN5efrHI0GnoJUWaZKmSM3UeMo4qf74IpAZt9qr0MVvd8FQvRx9G3GYdd4gLHnX6LA1lUYm1
A6Ww6az19YtpN9w4SmhMfUGbPHR0WehgqhZjl5g/AMB07RxUgHaYEW/ArdZ6IJK34tSu4IsXDpVY
VNlKlLqAKAhUpZvEO/KgzxEXDahzoRYGtA9mnJ5ASF9es4ncTpprtjaNJM6KLrPvegxurs8tNKJZ
GB7drhpQe6N+yrqIkmSG+C/MjgGxAchYobClCnMYJTyMOWqg5CoWGVk2EJ18drZnurjWj565nV3F
xN/vd7SY2Ov+OnM0ZtugDHdpqHVG4+5zDErSs+pXuKLAacdiuSITHNdMP1JO7o+bElq2BxN81ubV
tThowiOsQO93lW7M7P2b+DT5k5C3aKYtJHB/XPLN6bsIMcnieA3As6mPi7tWhXdeIkUDITc7sFan
y/dMmBq9uMjMAPL6+uaXg3NX4exJ0BJpNrqZnFUXzMAdcoxuzPRBMZv7S5Qj8+OknTLVpaJ6KLX8
7m0+haKLXW7wg5s8j5fK879ibFpCKfhnAbN3sVKmaskBeYegnvi2k/fjFmJ+GZRFnqxU7hvRT84S
yExDdWPw97q/0mcBc5B55tEW08BnR84DSuFtFWjoiO3QNZFNdm1zgi1gux2DBrAY39JAAv9Ht2kv
gWU1LkhZEnIoDnDS8vYie1HTXSvxnQnygl2opRHigsP4MTomuex5A0NoLMTV1RCwiM29CE/vnb+v
nygEbF6wD6jrGUnOtGoHJaGY7zY9u0kca4Q1mLUzJ6Zim9X9PQsFXRsFOmorcsR8qrY/C+976eeo
lvGB4O0+PQZlvYmeEXc6AZRjVQoEcevjNnbr9xKuumNE4hlKfDmbjqoQLQzf0Z4RgbypQaiFO3yR
0SnA7iylF2WIRpYorIWpP2G0w9LmdYywQuDnHy9Fl7dbyLSsw+1MTmqJv3K9KCTzWeO+8CS+Lsx5
6CvoAKTi/kd+QNoH8GpwxhhZJ7C9D4mNlvDqO7GXg1zmIgnm+IaKSBOv0IZB5/bBgipyCNd+uowG
o+tzfTKcug+lsiuxUc+kibUxXw0wD60+/wXgV1r0MM805H5SYxXgXXB5VAP9krHcfHVGA1byl3bx
NWgkQk269D3v1d65xGyuTbllJv0lFkvbOUyw2f4HuiKtjbrNu3vgLjfQsK6v8OCQ+qdmnmvpknNc
IVRmbNsCQeSCjM/TSoaxumXv5axDVmcjS/FPCe1jmGSzIzuooC6M7tx4VesMa++riH+YBhUOwgWS
6vT8PNVRbMSevCyQsNKCBQakPErlGqcqGd8eOdBiVqyjfnku/3UMRKnTrIuN3cEbkP64z5kabV+c
EMKg1u5hRJi5wRHMwhxnfvTwk94GIQsHaB5cFhecs3ebudhFB3NxaJD5cC/2VGVm7XNQ/jMVNnsQ
gMzmyPLaAq0XGNZ07DDyQ4CRii8Rr3o8BAlAc0f3S7Ss6S5HbZ4M1hTG+usTaHGY/phQ62XQOks6
EW1hZ/9F5bOleSMWRkLYr2DBJEsGjzRKQNX8evxWA8TJ6tWVAoiAdHI7J7EGRC1TRDu2CgVEOWl9
DYPD0Y3pIWCZeBMmiu1zSVJQ9tAzDJpcnicojpOFrZoWlZo9rswqOqjMmFY1qAh/rtr3vdV22FE4
bqCsEmJnJ+/997XgNAVTGJdFbW+Mrj8OJ/D6SMHv6QniqKes5nx8AZB1mlAhB/nJOiMrW3WL9ov7
3vWP3Db1bkvtpXror0ChJ16gr+oYtgoLka9mYSA+Pws7kSljtlUEpg9OH2YrwI1c9FiRWeaseN86
+sPxm4Z+As3M6rsifgvtemCk0m2TId1d1eC0lcQo5RnB1rPwL+SMCnpF26wLPHJjhI0euX3oBljD
wP7inmRtZFOuAabe4k5FS/JWu10ZRFFTuq19FjBd6eiuhavcMD8l8r2G48kpk+2144HVvIInXI86
2/BQUfuSp2vZRwlI/1DIMLLmoDks55u8qi+qnsTDOFtX+tYqN88cgoAgovLSrIEE8I++m6ERIWJi
lKerfPUtwNIZ7zHdqiAjC8Q4lww+RUHMj0/WAVYWGvJGMWDNz9msJ37TYTaytrrqskNHlE/XQjIy
eJ6Fz2WNywzQUcORB1oAW4YszOAxgJUd8/jF3YDzi3GmoeyxpmhOXK4uEss7uzBETYWr1XKvIeQ9
gvP6dIP8G2hrUvQrmiH/cGYP9dFk+pSh1/nVUJbSXcaFT+VRAAxHdv9+Ol2abhm/3xz7wkvlg1vk
voh8rEjY8y2VsUw+BtFgPGBAMNoBF4Hl/jN1+hk5X/Dj2GwEhkvbMd93SfrZLn//ZXgIgVYxZi4j
7hU/3yFcuS59rBAvJVegxTCuI4+G2liNmLZ6+ipmWOtMnmW52QI4twgyg0ym0gNJO61YkHu1YRop
89hj4fp6+RM8RiGeOsUI4NqHLhxjGiC+wFCperhP23PW3FK0nqHHXAoo2dkI9SpFRGK21q2b3RN8
SdlkaJYnmO9Cu/AAXPG1O3Lki9gsCw5jRKDUZuD4Yfam3mdWOzbLWV29RUYtf1w2GswcGmQljSIE
HywfjKR4gqGVrgAXI69+jIgQ6RCtmRZYmfjvK2kiG0MZF3IFN6pyCzLzc3MCrIBY35XIJP0QTcpD
uNz5R5m/oSoOm8//+cZRiPoEVXNOaHlxbWc+K6LwvI5MUtZmjelhF9Zso+oTNUGpSHBRnMY+wFrd
4F94dhq7U+IHS01q03Lf/fDxOgjyd59VIMiqoYbcl1GNhxvpIY+LC877kce6xQMingPJTpydobbg
hiUeELqukM/uxdXs0E5x5aOPzOmHRkfFsOPhK1j/nvTWnQKtfaYuWwyyULilEBRcpgSVLsSjR/MP
n7ELWdwzlfKKadHb38RjPr1TXChNyfAEl0gF3A2mnMPtwN/lLWWaCVHYjMNPvfluF1//EZMlewn9
1f1csHlxef0b61Bb3gZAWyqFDMAZQm5S9T8qDHOjQQwdBv6WQxRyNDFP6XjWtkJfMBHQFGW/7bOv
F/a0QlXZhDFfr2YKFbQ3I7zQAvvsaw0sWxkmbFnwjs/8FhFczNtIINoKomXbc+N2Py9rrwX3kF+P
luhHxewHyjdmhPIigtS/vyuNpll8ecjtud2U8REjlrxtEK9YXxE+2/JygXGbJyaKnesaC8GDzFWb
vjsi6g41hsaortoYGbU7Q/vKUZLu0evGGl71FtOH7dbUPh9V2+PvkxON6jzHMw+X9VCwaE7Al/SK
LIv36vm0EXe8Z6sQJNditgHfoIwnzQHGdySDJ22CTlfEsX/3cIIdfQzRglVKEAOzd+xZ/yoCOp8g
i4Zv4Trk26T678RAyikHriwBVQhYDpkOgWzvNPXmu8iK3wcqPniur2c2zUMqCw2Di6mTtdh7F5ZC
Ui6yUyCrL/mhwhCr/FLscnXaKRwXxdBLWaOxHEVAF7uaey/I97zbLTglYVFveY/AgoR5l1y1fnNO
rumWxX6Nke1RpaE5hWKmynhIRzi/L3ekCgZfiYvU8rZGrReawjWIcKgR/Cup31tWCqJyPO/1I2Tg
SRVfzGKnEZTEBpAEGKzkSWAsZDJmauWapGuR5NVASdG7hy+C7ZAn4S7ci4Dnyuzkz/4P9QD1wddY
BJPSCJD458boqfWEzo7WF+rNNzEdpYqTi3Z3Y9ElCs3QE+k+JsNx+D650bthjPQvRJiVa+R+YHZ0
S5aDIchRacgtIfI0DH1iGA29IAClNM2dJfPkzBxj7pWTSUoimXkvO/ZkNKSPT2fdPMleiTGx7HRq
AsnUy97ja2YxDNWQeo89b/rpCIsMszYtUgrQlwAL6FxXerenGPyK/47dHYiyrKVzlr7Ka+wlUPmr
3qDK60e7VGrIHI7WwlkHMeHJyAKTPcAcP93NMj6SrxOj2UguRxSeVUjEE5WFhjWhZdiuj/JF2SF9
wfIPjpHycfdJEfpP0XmtLHxJp5pAcFITef7TK7PG8z/xA4iEUFOZPg/AMuyjnfsEubZ4Z3sYJLtD
xnRsFDQPzWSJsmj80zdArp3jJkdtJz6vB+Mt6gXa6XO4vOFoT+u8NEqUp+dqcvfMITwsY+cBxHP9
1H6XXNAj53MGPpvuw1G97UgkbYZvGPNcH0t9ygle4eDzqtKuMzW7Q2P/joWiKg4kGJ93aWZSNcOU
2E5l0yx91mEsT99nSk1jDZ48JyYpoV11OOEey+7W0D9URiqa78yyn42v9Jqy76ogXFp+RzryfNPh
QfbagzpwcY53PRp3DJUljCgePvDiNZKbtvSFHLPuHWWeL00/tXDGzVMg9yhiMCsENfWR6baSQsi8
/01eckM8tj3kp4dtO220J+TxNN2HVl0jFxWR9/PAfberZ99A5aU3dJvPjQxcXNn46hrMGW4zv4EV
uJslD2dS4mLCTlDhmEUNuxvY4Bj2Z9YY2pFtbr49AmUhvtK3uk87JUJ2H6BK03zgkBxtHGQZ5yQB
VpZkRAOlJESL+ezjMYFZ/2R+OK1nZtoZ364w1F7WNDkOQxvLmJR0gB+DG5o90JDIIqk2HGV0k/5k
rgmvfqelGFgJhSL/yzcpYG/kUY7Sgr2iUV7Cul91htU0YQPszS4n6AEXtIVmcr80TFliX/uUO1pV
FIiiKP+lf/gA4YXs7V6kUbAq2rdAKrawEtBbVlqDLG/j9C0WGzlc3jkEdmirjn5a3XsZu/ui0Em4
4zOBH/eX25BNAGdwjVYrVwBjZeSYNC0lq7aI9TSY875TLzqGUsZTlBMSzPtJhjjeYXsv3++fIqEy
wS/9o3hbfM2A9HmDDbCUQu0d8/k3xtLAssbrMOI35rnLGczhrpsIBmcRKiUXzimT27Lp7I27O+Ji
T34jtDqWzi7yylq2E2/FwFIl4Asiy17S18XJKlbtk5pOG3APnw+FxBmV3fDqTZfML1MUMlWH22V0
xQi/4idpmjQeIX4ortSsDIyQwxx7QAr3g4uvj4Xk/CfZOzDFAS97IFBUdAjo6Z7bsaWTlU1AQwLV
W3Z9+2IQPelx9qMHRhYIAH8h2v+1juvzxS0J44A5Uiw+4HUW7mWuewVJ1nJ6cudpYkHHypFK+Pjj
rgEt6TuRehwzgn9iVt+wptisEZKnLe6jAWbJKbJ5brsI1BGF2ncXAjeLYahA9XyWdwSBtUh5EvMd
2Uyd8ykgMYTgA/ny9AuZ797uiuoKniNNFsKpBbk+k+7szE8hxS+bPXXvJhzdSGjzrX1qkDqsPeS1
GtQ8tMwlf2m324SVIOiE8yzxaDJXGbMQjsk9qAFIPULBmwMV1wvMQPH6NAaVLDMdM620FLdeJf3a
+MIDaVI7H9ahNItKi6vFGbAVLn5e7VCmW+2+FhaxfXDNjz0EfhBBuxYhMaRqAPZqDu1Qtc8O0CiT
eGGOCRAkZqqSlDwaOYkIwT1NCATzS8tr4kIPFf1qbSqHypZbkhbQelfM1b/MLF5BqqX2AVX8wwxU
cOiDz0Ce2qd1ZTVgFUsWeF2cDI8Gr+Ek33wY45NT3U8SYYXNB4Fmjs/gil5wwtZJqiZMotGyPKrO
VjxUGmYcWSlDVvWtoIOOr8Gg314YhKs8zDQznnaxDKNpVxd68YgUWfTCoiPRBMMCN0pAx1evyzgL
JNO+IqTbI9OOkTI5W8nwvssov6Rt1NP9+9VSYswAE5zjY/n0tUwFuO7L2qWl7CsFZ51tC6eJVXlw
A8gG6tatoJkcdZdRmYX+jzTqM7m3PBp57gqAzhZMXFIz31GgKFaRpFf6SbMcXQMdfawC2k3TFx/1
NGzGO1dy3GtKd9w64FdQ551Si9ixKRWN6rkZsZG0+M9RyIXktMInSBanT7GmLQ4/W6+45kSc+qqP
CVTBT/9wpcSsy5ZR5G4q0ZQNBf8nbT2IDUf9IgWysXvh1U5JqVVikeIgXR/f1tqKolDQOvQZOOBY
oK21ouaWthNCDhm304rwSGNwE8O2rXmhS881/ehy+gKO2x+ZlgqALlBunTZfRowF2sAKUOzgqNKp
SoRcqs8Lp+cJWRl8k6GhiwbkbUVdcL2I1UkkOQfuTW1eK4O0fIDVgL/vCgnoERXJsnYXcwjp10cz
MczVjE/I8EHNnmq0S5u8rGIQZefP3wq1/JOhasfkIcrCURhdOyb3Y4RTexgaNQelVg29OCeSzbjD
MonhANnBWMmessMbrcZNkarWabVVVTLkNXOGfEX2aZpSZJVtn5LGA2U8uJ21XoZT1Upmn89n+iFi
H7G5t8MyPl+xSBxvZ2sReTMbbMU9RYmNQpbHW0COPuL1bZcjUuG3xBOmQIbA2QvFxTHy9skjTy3R
RuHZokFwaQZBYWv3Bv/hCb9aae720QQA4opdJuqxrucL1+ODmXXH0fwY11dz51CfnrVQWATTFr/F
3DdA4942/K2La05hLZ7rB6vhzng1x9cxNsGBowBjsN7WLKP0YVWwV7CjP1QrStU2SvalL+0AU+ga
Jh6r0xb6qercnhbYB3s+IGNMvgOPss+tJc1WKrbXzj4bjoKcedeUGNNX8JsYCu/nZTRD4pYLmnBp
JxT8+OidhqxCN1PPW6TR910cWiQRFGYUarDjOjRYiENDE4fZqS9Hdzbi9gLb0vZ4kfHI4xa06pEI
zE73wijBVUGt72A3kngS15HOQCh715rN8M0L1dlPr64uRebPDiIUn7qzBVnmbPaHO4nq4N/ABRA6
zHyZy/raqj+MOeKvpfLeKxAsQclVCcbX9m7C3Q/PEKKq8BOOyOFkOSb/yOw9T8qYXCW9AHLfBvXa
y7XaWlOb4wnDcLvNCPLZDu9wkphzS56iEXQrmSrCxOR4gy3+uS1V+vg9pgD0x+lrC9FA1sL4xRUg
yEBz+/y2aX2mtnD+hcgW2CvNjCU1nVTcqiHf1HjRWp0bxF0mZjkW7nHqPMPkIEZjEytIx5YsZBpC
v4NYC4VUPQgSq/ru5rIXdpOg6peTlQR0uBsyyxalJEWlwqgt9p8j6kx7Yf01yzYScCrUzbhkuoRf
nOpPSkqvOD9S2VkhR6hTglSLvvbIjFMIuAGomU2TbkUtIEZ7PqlqyMZbMZyY7g4e2TtlGNAE/F5I
h6ScRj6yq7WWVStV2MvxC1C0u70h94g8hm70dUoz277R4VdDu2a5Ljl+Cy3s9LBCMvyU970+ewia
iOLRCZitbDz6yneuME2ceN+9xGjKMZsgD4VkQv6Xsvc4GhCZwS3WCV0qEChsYWvDmtxBdzfU5hHs
OVD1HvBk60NLYRoVgE/093JiTMJUKETrvq6lmDzdZ+Dvc0dXF7p0GthLMgepZZ3k4WSyKNPj/nrT
8hNKYKjWMfODgpDAJiWCyKYtT+Ai2Uror/zZOwzNpGI7XE5DHbgcUQFMcR7FSj4VgItwul1bRXJD
0CsnKkXCmRr49SS/4qX3qaGV+3tpWdaNyZ80M7VmTC5DYJ26TrmaRErlg7yzZOJkiE9bMBN+HbMC
9L+UFKCz4HcmUlA6H4xHu8GEgqwWz4psT8M8YobKEGpI0OrnuHi2vT1cq0+8XO2/8BRdw9v/mWiQ
j1JO11Ibux+HV5FEssVf2DiXHKq7HFbIBZ5JrtcgQQtSWByf+uWnLTJ+lNyuEFUX6YYXQYT+zklA
Y5paZ1j41GFnb+Km4PLecY2dtjDTp3qHIGTaQ5hzyeas/pKcnKOB5QLi0k76f+2MLSSW/jPbpxrM
ubGFNyzV4OdFSvwa0QEkb1AYpA73dIEPpoMjyVtvIwbVY3Yn3ijjVq3147W6YDNJjtZ3rMLHCWn1
PvzUWkoNZtci5oU1Qkx8r9oxJURkwtB4fS/ReS7yp32tWiFqQX13GHt87li2MYzrwrVh65ee55tZ
vv4fRu8mIfR03JaB0AtN15tQu32aEYC37Tty05MLa6Cezyh5zAH/tsPsJ3VCa7bp8YvdU9TUcOC5
r/9wcKKZm17T0NxbY9xkbPIch2vxjLKjCn9izO0FeXT4elNc3J/lDCWyxGA+oM2IzLBX8T7wJEn1
xNLni1rBwkfWVsxAYqqgSWeEsqC1tcQPX7Eie7dMU/nBsUyunlP0tVq4FDdUWQ6AQUrnQwByLgNd
BTxgAVjOZGgsmWVWE6xmlQI6isEjiTiwNzlmFKrR4phN1Qm7m9zWWA+bRNuzLSYsSzoIbAz2H1hc
toOvh3C9Xt001I2hTrCbwqTUiHu3P4GaGf4jCFpFRrEb5yIIYLotcHRDUGnUzTmY2i1Z/8J/rJ5s
OSWfSu1ZcDSszAz1Hh3Uou8Ut7VeV2bdTzY+qfTgH9XcY2FwEXM8a1M/sjYAkUEZpRae0dLm5KI+
VHBraaVhFlxogZBd0MbTNaugZGQ7fPDPmcIOsTN95PUGrrVnBS79n1xdn6VxPuzkwc2va58GNXuR
jy1a3DMBHm7x4TZ3OrdauQYLXm16fEAE5d3CwirSA7ztzYUpTVD58EuVzAXx6MEE9Y4kbSgtT29V
xr6AA8gZpwBkT71r94SAV713RwqUyuZ3ueFPDHxUslGZM1kaXELlVSEYpzw20Y3gg2heUtzIP4FW
azpLQAK65QnI5o4IrJx4hccHy79DmGiUUaPv874+I57gajlCDWLav7tBBPcup2BiF98Xg7Y3WPaQ
hb76zWrkhmcCAm+BGQKY4wbfoBh7nmZ69EIpRMn1Q0WHuiIg9Aw7xETb5AEh/ThFLVWVOtTxXmO+
aIS3EsPo6KWl/aXee/Jw6COW4/kUK5PTWfYwj/pagQ3yET7RaStRxWSbL5LzivCC5bua6ESARBtd
iSp+CLK0+Gjl3opNQgLHePsL05WsGjABc9bWfK5rlOb0s+iLSiYVCLNuA/mKmf5gp54tmCIin2dD
0LdBRY0nnGxbibPj7lKcAgICLbVZ2/uHycrznSF+va3VtbEEOjvMu2DDsBtFXv0EySFUCrLtFGf6
E/VHpDsMNxpQVGd+3PfZATWw/ESeG6xQMIxidWSMb5ctgdkyCE204gShPOd6zoczVvWRLtQZ+yQS
W1H6sfUpXCy+hUzFe+uTrfacq4D8ME4x8j04T/b6xBYeAcwbeqK2yMWrBiz8JCNj9HA3CA0+rFDA
+clMQZxYTaNzKOBl61f2/dDemI/prE0xBJ0vgAqXVkNtAZ4qpQ6+3CEsOdHfz1bhQ3n4lx1yjeOW
u8nOKqK8VB3eIvAiKziudiaJHEOCyQFOM4YDBPtvLPSVXN1hq7jp1OwFwewLo+C59px939Mm1GzE
3AdHGfyfa5lpkeK16d5oQFidK8RHziaAWcG3osbuw2e98C2OjwC3AQQBR+o+vxf5mTH3Ljpdnb7c
Dy4miD3T9QdxUrbktV4Ldw0RHs22lNLEEajZVQS6uuIya7D2AEZPibds9CuftW64Zi9m4eVM5MNZ
wkffDrObLd2L8hnM8IxOaybgEM9xonjgEGm6Lk35lhrvfipV9l9VsKSmsw3TPPVARbO5IfvKE0VV
u00VQ4FpJI6H4TizOAKgU36RntRNlAXS0jvmItGJb8TNWvDypGIdLOZuHPn1imH9V8YoF2OXlXWB
SnsmCGqhiXypBmFiBg0F8X2RifMzQOmKItY8CtLqV5xN4k52Hbuv+cQBQzs4LDOwtMrjtAOIJxjA
+ldPuoPzPyKNqVfrNl5VZeFn0DKSWdP8yp71QqqA+qxj4NK6HByktnMiEYfbaLTnr/F00mfUybWJ
UIT2jWbug6xiw+ileuVdp+jppHm0ROee2cAFBQjltzbfv3WmsCDT/9y+FaWqo5Y4AUmV7ih1P1D4
Gp3vqsVgYp/SdqnQ70gdjKiDA7AQUMEQtTiQ2+h9rHqdfZgtR8N5CEpC3EJ8a+hJcs78jqaq5shy
na1DGpfEae3IBvkO7rhvviJsgW9x3OP0e0CJjtKnKr7hQabQujDN04raeB+k+d2d9HRDdnuzndZo
LcU7JtB18jLnEZS3QnVleP5vamMFt0bXU7Dvsg8/BRTNAVLR1jMCLspMMUHrTnhN38b3LQsMlxs7
dFZaqYd7Qot1673tq/P9ThVXupo/lHJrKZAW7jwM4G39HVWZuXLdFAVdRUehXuL8axJ3vBpIT0Qh
qLg6FLJe8DBMIDGzEZkqsYX675YEL7Dl/baB2yOGw7+NweCbsXv6W0mjxmnuoMcU09Hq3/ZH0Kvz
8il8X4BLEkGQVDPau7p2nECSNO3EXkMWe4nLP2ImO0H/RjzB2PAEa9Uep1og9LpaHK/3ytNQ6Hvt
vEjBQ36KV3msVlEkatvwjuFCMKvZHvwlr7ePyWkTFOQMr+5Q1Sj70kgINs1ZD5zZzPK67a755I6F
yvVCzN182XN9brhuNCIRanv8WB/jmWF8jrm6aFZz1sJDdkkqdNq92QBM/j1NAZoFYsN9BZ7vsnZI
yVCI7vBkDe7WkbXqcDOvAMUZYMu43kTZjscZH6CcGZZ6ziFAU4lROANAl5mcShCTRbAVOYwQeIvw
mCUYqrKaw53Z5I9kffKN+qAIbWZiUPk7XTBJkSS3WVvFPOkEKkf/S71+DN3CMfr7a403VzHvH/CL
0LFClXJOiS/jUTJTWOBln86YN+mfP/STyE8U0j8tp0tZh5+NmWLvU4GThx84DQxrwogPthr9QH9r
hBuGI0ULB6Lkya2Ajrzc7z2nxQuSkgTRzLH+4DwxNOt2CS2bABwwEt7mm8JCschlop38XoeLeBY6
ULYqbVcjjx7BQ8pinDqXgOfVfWLwGVds8MKrK6uGahdhw8fNSdKVTcfWEfsQ/zGrNJA5ZyoTt/Ds
2Nxr4L7DaZ2ZgD0FWNFf1f452087CVSXA1kv/JSOsnnWYWM7NYbGUoSJDy5fWuRazEwhYaJi92AJ
NI1h4GAT2uLMVJfQS6nvStk34uOilZGd7Ly95pIhwR3eyg5ivGMbbSvXpbcR8UjgiFrHhm8RbpLC
zMgjv3iZFwlULk0uclTj1I0IJtVhZGL0QPIELSDfH6KDa+kNydlZ6m4kTP6DDxNCi0gYWmfpV3Dj
5+CWRhrYn5x+5gavNdVy0BTjeE1mfh7oj3MY9CAGRrr1THWdksaX3A7Y7gg4CuFvP5Rfrp3bRIh0
FMjbnTDLTTRtuovkiE0Na0wcJdjTcqU66G9RXarEwgg/TTQjzvg8Rxh9rfE53PsO8Zt5a0TJ7JHB
wZQnHAVduXIC4wlHhD4BdTbnhn+1mmoaNoBzrYa/NYdQ4FsYceZ8NgcizgR50gowaWC6RVgkmxB2
+1cZMROq+87c/kUGUu1TqfdD6uas+mX7ub/+0y+wgiaJZYAJIWpTg3j6PPQFEEguTVG/D+rC4qkW
u+5edpgbhOOVyfh6lFVoBN0uWdZ3YlDlMFGEHl2XluDlb6DxWcTn1kMEv2Wk6EPIq85VmQPvFNGA
rn1qCGI/3+tDjqtoHcJFjyq+InRfz1K4p3gTugjMBp8DOFTWK2gJ90ho/XlF5x8AMmGQBXhpdPWt
7FH31LjDMK+E/Nzc3sHYnY5C/flsJRj5W3HIHdieGaPv+d/JOD/Ty+phP74mBhNXvOVzWr5D3Dxk
uqYoX2c8RS9CRTgJbqB80YM9fg+haiLjaijj4Z1EGgEpV9pnIcA27eINqV/ksezK/WqGfs+B+xev
/CEi4JBs9CI1H8WGBKNi9BS5BYKfNsXCa3wSWy6ajMkDJa+aQr89GZ76okTCQJ0rgcB0enf+4rkX
lvZJrRiHEhYw+H53CB8w7t62S9xSAVBFNwwJRIP48iYgzBVHQKUFHGepEIfr9nDhX8k7H528CtIt
nbz9LFwjC1ASwbghR9LQUxozqIj+1euCTh8fQVmbRbHE58E+WSYNxMNXicJVg4oV92qZ4VoBHPAA
PTXsCxdBdMdTrLrsrHHaHpktQQYlFyd1laigFf8fI76TSUZgK3OrScQzpmtVKkvj5xJwFpuSnSHK
b+Lvv0HRLb9ubT2SJCFtiq7kYKwqgSRpsc8+e31MYMSTLkHGRv1D2gHEor4O6AZTHO+NLSN0GUJ9
zZwRZH9gV8Z2o924gtGwjiD9J1r5/9SvpGXNbNvjqpBSdBFOnlE3BIOBMOYZR67Mwb+1xJw/emzY
6soVKA2Ww2ISsRwg+hYix+TC63cAprOy33SVc7WgQhr6rr1+x1AMlryDecnhO9T7zNpkvezuQWev
nEK3a9KoIlsipiPKV4wklG0/lZEf2PlBobq7QjrBDb1GuSz5wOW2aAAYwuGZELeVwQEcQNoEnlVD
1RRrZncQGEL8fkTNcn1UL0QienrH4j5DPZ9wQAkLflQ+OBo1cPKF3o4MsM2BdN4EcGIcvp8sMG3D
6B1cXtMp/h+VQ2CygVkbuLQNlr6tBNVR//7ig/ayuEpj2A90AoynXVa4LgPWYBNgTObdxJzhM/zd
//8CX13Ddoz/79W+wRvZl1bVWunaz7m1pxJJcc0KkgTn+G4d0QvLBPnaoZgRUXdTNkTgTR9lv/Zz
qqA0QovBw/JlCXDYOZe5VCgabQoYVVYFipyq7du+W4S8uPw6IE4Y2gHsBH09h8G2subQktP2Fb1h
iS1nSKUqMZW3ixD9SV2/veK56iuJHVlLk39QVRPXs6ZoZRChCyg6dm0In5FruZx0OC+0sQT+cw09
bne/UAJwMArW9mcvFsiFxRgBuZkF09aBSPefkhlRciDtjtqImEB7/OH/Ord3Gq01RXVzn5iVlYk7
z9+SOVAd0+M9PK3OEGd3gV4zN7J8K6YV0ns8nKWEsJinozQo5GSYUrhalnOLrcllMaVM/nJXbJf4
r5mb2Zz4o+ZTmUQbTWspyIMjDMGGedvUSa2Bwl7HdHM0RG/dUEobg+1pAYQHWLaYqJ9SGo+Zi0eM
ozAVqu7hIHuXnoCBRUNcq/Io2iy+N34a4Eb4QIM0T+S7QKTcwvU4NCTAqxZ9t9Msouy5heimoK9E
LSuZ9hWaVsbXWYu4JMakr/JGU0tLPyC4Iz7wJm9MCeDL8vT1J8wk8tomhcmBxYSZ7jiwcvFThYEd
Bi0a3FBN5bDWuhLzSczRHZk1fXceJ4DQdbwOC5AhYpUOWqJJT41t5ohe/939Sx4q5NlKqcqeBo1Z
OGUWNUIZcLClt5xzKOuZMqMrbY8lTA+ejarH+5U4hgcBLWem0IDODSE+ZcZAtyeIM5BWj1aktQlJ
A9pPR+hCCaimxr4BmvZp9+nj08HYv2r1GeHWSep/xn5xXJ+goE5FMQlYkPwHjsxJZCp+FPFXC2Zl
Gr9RZTvClGaJ17/5gN4as9eVNtNOkCPf1vw0jAqGvhSGRmJVYZGWXwSmLJxdcxt3+uI26vNQmXYJ
thNiomJtnVFE0mUtA8yNWe4lFTMzD1pxgtVLBaFR0+Pra48Lpb5a0Mr7/XRmfdvRf5o2lNUv9SzG
hbNKgVp6F12qoiSRZT05+2SW9nrtFR0yYerEFsf7Y1KdfuwkgtRNZWaHkz1s9o57fL8jBlD/wWSs
p6o6bUBFK5amhzzSDs+2xo/94trguQuRfEZ/LZqhk44R7ElkhOVG6ORNFntP1QFCoyl1LL7SRu74
tklMD1mHCKci8QyjNsa+IvgGBtj5KeXO484zHxRwqdHpySvY6ZsffC0F1VNapS6UPojr4vD67wsN
lS3Enezk0THrxhQNJ7QpCpi94z0aYtoOjUrlDwpb0XMQ7znGUIwcNBg7n1kQ8BDzAIhsdruFeW0E
A/B+05LUuRT8/P8ax8xoiFzFUq5jwXH8ZMqV0Ka07HrAXxdJQUrB6uyOLz4JdGWqiFiZaLQatCsO
ufVwLMI8XIU0jUhKhHOx5K1h/ZxHv7hbID8E0lw35MuflTdKgkMnSMgwju62mcW5MgSOrgsEXoEx
+o6jmPtRU8Lj0S7Pywj8pePDw9xi/tPyf1jgB37/gWzef6yNs2hfQZdAZzoCmNI7C5F8M0izyvJF
C/irIiTWZxo0FQHD2iimp4PIasb8Qz2ibSulW/j/kAVHZRrNxpsEAS2iMTsAkLaFUMbScAHnmE6Q
JQSMiaAnqC7SZuSJC2iwqCUIruX/zzR+4t3ggCI8qNdYVBlJsA8WVuBzp5viKVBItjetnu9FXM4e
hDa1nIbAMZyBYZNw2nQiMulZdp6OgOFDj7yGxeqHsLulFqgZVOIxI+hl/LIrfigRyRHm84CBZ4ca
70gti3a8kUBsmPVs3nWL+1a1Sg4a2S3GhfBjr/GC4uu5EbJHYP6eQO9I/2Ao9BzmQJIwpVws5SOI
8bLkG4g5DSO4LkDqgSF5X+oARElpmET2Io/IjMPwSmPlAcVo2+8U5mEUTkIXi2wkCABEo8jI9YqJ
8NN13NnMUW4sYoEF4uoD1crvtMS+Q59GddxibKtlFMdIJ30XgSkwWvF6yRAL26GpRlHeLHqXXg6+
Z/HcgAhnAXV1NZKOKV3KpQk7tLgGHFLdiKK/gBxcFU+M1JJR//Jwxw9q8QSews6/J+LYEgwRQh3W
TVMJm54YwRAhv3D1dEmFc88KR20u+6b2UEhxW8EsKUScygbB3BWGAp01upLpsHmT09yf3ySqWbNV
0Pful6AQN7vM7GaMqIcxheZ6ioETSYJW/FWdA21ltFV6d16PFNqSeyXD98ZKlSPRGhlTE0K/NKyw
msLZcDcKg7hsdGAAu+H1umCd4cPGFPaRa3y1EFqXPbIaLHaqlSVvFJCDPRsdx3B8mb680T7/IJQB
PdXFQ73hH+rovlKyjww2f26vnGDnBM7RfZX/SwrOgFWUlzK9DRlk3OmzLvxwB8vBugRGSOm9J7vX
e3kbr4yNw8fSkOyFt3gr6hZXsObvbgHz7HgcJ65DPYjgzhWlj6toXasqT0wkxiLF9GPRoPoINATc
qls8kXd7KumiNnbq+7jNy9wQvxU0hrGTlgjXxhFFznjtxbO0zYjBVyHuvaXtuG0RuOy6g+NDQB5u
gbFoC5ftbF1GQpDmk+2u3QYbc0rvGeFgTMWks3pGpQrYbjMfPMISPuCLgHRiNhIBsX98ULFQ1MXd
pSgX6uhjD2gh1FaksLBl+jNodAnR+nuwS8XAzw7hG4vBmFsfQqQbVOqPwyEACBFSt0264okSk32M
G15NO4hgKuoaaZCtVq4oaPq61yKTRaw3TZ7CqKgk5owuBeLDE0uy4a5Bwky14V/Gtv8PGAcovRth
WbBoe9+SHEZSd+61xneA6PuK+h4It+S5RwBKSSrw7BrfMmGiLoTYujAu8LSjUlhTlkB+kpuiESlh
ZPZOdIFXNa+GWn2CIxkWpp2ljAORzHfHtMTZp+9WuRUw3P8mX8Zzow6e2+z2gZEeHI+AaLDSh9H1
iki3q04ASnhxdxI8Jou7y0CVMBHDgaE2IS4MrBajU9YA11uPZirRbVVWpVxOOB0cDBr72EIXZmk2
gOkaBKqAcR0ycvBVIsbN3hCmzqsoTkqT6OAZ2Hym0M4/Ew9zBrcSUroHYk5QJ+W7Ze/HYIVwTO0C
ZVv/CYvg32Op+z7uRB/HJZtXkAK2G2y46MqQUCuCW6v0XwwyfdduQgacHw5kUQ7ngFb2c7ysALKy
1re3v2lzPkpQJuMRXKG8wfeR6oRYKmBDDeIW7O9gyFNPtggAPmhAwtAZk5FLrqG3vpuhvEQnFIus
r/h1X6w27v7vN6VcYEI+2d23h+0DZnPGQxKf3gA9sdpyIMoTn+MGDcCwhthAQN5fJCk5iNKUQXAG
iDcxA3Lbnx2khsZ+rGdvmAxAsoXWjjsUWVeH9M8F8xqYpm13Ng0Xil5xmcqQmXauKjeXQqJS8pLI
uMema5XB2YtC7/xTBKDLMtHh4srnxBeZEXTNGB16hgofGPxIEFYEq8CxIHNHHVw1pvHCr7Ltam7s
2vYksN4P/DqiJ4t4iPA30v4xLSsRBADk99oOFjjdSIei2JczucYPx5pXRiNQuHTc0m1RfQN2mNBY
lqTw7lqwibGStUdO8ZrXWRhxCGGxe/A6Ny1CRUTGWIV+W/VVz8e1EnKit6L33qywFDDLw0TBCNFB
ufKzNout+kBrLgk6JuH83iVYXxHZ+EDNtpqXtEo6ky9t+kXVIpC2SMRSnjYnA/D86QE8Ry+cd4Rl
wAo6vwhZGcI3qbaCTwaptX8xQFAHrLnmoCDInyvDwt3g5YAe/5IWW6evljYKvJQHDZpKRDvOO2MD
cpvePk1MF8tKNp97fp33+MFLEHU31Xel4SCxbidJvAqOWkJ0cZLwd710l9l+PKLPwNwN4YK1zDAo
VrVm3zFe/D5Y5h8XOIE4ebxKcsZmFDV1y2jn4xECY3HZ/+vlH1dEtPG2SVktRosm3ltAZ8FT3RwG
NNixfmkIzpuCa/YOJgKzcj3EQQbwxnADObBq0wutHZoe+6EycaLn989/tixwdpEVvq1sArtpMVh9
Uor2rx/IlCWDa75oze9IjPU+rtb1HEp4i461N5BpJEUJqQpDPX3Lds30/cLXb4vbqYd2/0+J0cXE
C/w8q40sfEXRvfuI1vU2Agd3sG3GxYLGb8AHtfIbdZGuLsUqwuuqmpv3xVvqtxKKSUprDZZQR+OJ
xl8UCRm9fseiEmz2BXMhxAgwNkPc7PW01sNgYz/i6A7n0tyuEKEncfbJkhqb71+O3waEfLEel8pP
JmxUKULzPr1Ie1B7RC5h5nDKhj3y5AcRadVbYsAPuQE6yYBrKXqzIh8akjFPeLEmmIawLwar6tyc
Tp04uEHQsWMd8tT74XOvJgGiQKQs5XTgcAK3dOAr2CG4QH/2hsOyadpR9qxHPEqsc4ZikLHlWpV1
yfRABv3R2HsgaO0M8n8LTe+IPSsDqxDGXN+MrwmaqSdngDegXD6HNZn0poTQi5s3eTyAorMB0LrC
deHiuSUeaOqLRCz3OsC87+tihAlzTcnR9hOSXNUQW0dfzwRkBsyWx/TNbFBvUuOpCjbOUaEGUATp
GB4A9HRy6Uxe/KNrybZ8MA4O6EtYxqH6bqb31QtPPXlzM0/RXks+EuHJ2Sde0GM7YmJvpLPz8UfM
xtk4U2YN8lhk0coXIb+8WSxLTOjGIM5VP4jufys5upK2WAHH4cK8xRS44fAcf50Phr1r47QlF2kd
yPFEq875CExO87phWFIDO66aucoPUlwaucKG4XSIGCtHiRVmE6y8qwT0YtZ5MjDinedqNfKnKiuT
AGO1pQVtUY8iGzBHbvb7ABo4OQSgRIcVD8kxD3W5RUDUztdllAX2y+HZXOisBhnHy9VNg9XrBs1u
OwO5Has815/KKu6sUdqEoCLqtAClrTWdAZEwzpEt3hh3Yjyibf1baY7ZKa6usD0BhXd1n2Rvfe+u
vPh2ofhNrDXI2DzK0pjtQ8MasWMfUcNpM9U6B0S4XVWDO/Kjb4q5UyYnTl2TmphdkOCu4BNBr+js
UOoMYqwNmF1xbGAJeR4+t0UzSCTtQw0MriIxf/wHOaCJwSiI3S/0DeKr9+BKMFKSHGKLanSe+Z/L
vIAFBJMWSi39E/+n/7arkGvM0t1TtnZdOxuDjOOOMoAkCnBy2dRaUnDZSC/4CdP55dqo4Ir5Xj2t
7NvpPSpovL3w491f9UIGfiE3dN7yj5KzIcDPwbcT0H3WyiLrmDYb2HUREcPchprN25UhbUD0SoAx
P/Z2AdK04CR/KjAsTud/bWwnRmYF4fg5I5AHhll5qR2sa8HyjIJQrkEATj+YTfbt6vhw17XlHAZl
wmA3j/LSmc8A5zqW4QLnd4EbjlmT8X8V2dcaQREh/MplE/conory9pFDGNA3BUGjEGyj6Dsz9wFO
Q6Z4qluqSJhJTK/xWQXqFeXE1wLbcIsXNrNxhuuxYO19BlZ/tLkv9o507VQkPDEi5lv8xqJ3DyG6
9r+8CJ1LJLmgxOnqAukaul6VZ2JQCjekQoDcs5wEBZ62QBHV78Vn80c5h8EWX+/DlSytGciAYsDr
llcKsCsS4BD24wuitU6tI1kzbMHTyLnjvQgppHebYQ+YAsegY35fReRpPQ2GFhPHmFqtgGOnoQSE
BojH3p7FsvFQhe20mSQVBZgwbJ672mMPRI0nXAVHgn+uW0BhSmvPqiztw8iZWofHCRaSOQ8YbWOk
E5VYO1/f+BK7rerD7lnQ1AO1HLnHwjlg3Ke0D6jU1CA3QemubRvlEWPmmQLCcN1ER6MbEIY9SyVm
T+dThr5TQO6oHmcd57j2eLxxPGynQ0kKHQuCnrz+LVIwyCYoaJPKFKhL8g09GEiPG7cySP6G2gdO
b5XVEN4BWz1ylnmkfI4eKLA7rYpRo6Facw0M4k9/HnNAfuMdiTLRbjvz5ZmpKJWQWvZK++5OZMlp
k4tbBloePs0vm3jp4+X8d54+FOW8e6ukyCA7dnGiYahT5CaZ/as9ezUBICHl5uUIuMoCgK6moJBk
CjIt6IDtrrSY2t6zbhMi6+9rccZKUSJOh9sKl3XeQ08XmmCpxm381rWfzCAXGQxA40EgKQspYv9y
MKmpQg6TnCOSw/QYqfIrZRfkyxyPo/UTg1roJk8r2cTkEAX20EJBCMf9yFdzF784Fba3/8JE0s/9
VMZ53h/3HxyYqsQ4YiKUsItYFP+lAwiDgwKUT4jkD14geL1vX0ihps1hstchjqzWlG58WpJoilrk
YmtAIka4FWTbOJxvg7rIx5cKXKFXnQ391bUL0VIHunIdy/fq6jwoM1w4hFtze3iUmp2rb936wvEw
+6MTdv0jTg13ErRHW9ZOIOIYoYl060chacrABPvMdQa8ReolyotMEWzsXw7mKCBz2dyUYSu+3erk
UmTWCcvsNNaQ3gkmNZBPWVwFpRbYXULznXXcJA1MjaTvWSc8VgTMVAALO1e7lmbSoc/A24e4YwsD
2Zqz1DRWzcycvzaX8yJuWptqtly7GzgKCkFobkTRjqmkpuykDQIpqsUbevbIdFzEqv0uIvsvNpF9
PAPEVqkDKS9tyZEj/t6gNwOEsLpfR7fRJteNh0WIKaw8PN/7Ril6AnBVC6ZJDQLprfvIMQdeIoFE
RucDeSkObbXFwH5H+ZKZCLnCSXcalKjJv3bBJJwhgVxJ+owQwCu6SDkduwTwbThhLA4hxkBvloXw
W33Ef2W/d4jsykybvQLbQI6cvOE9MabICRId/2UzCr1SSoWxT+ey+ah6LUWdborezpaSzQUJTz+r
R7lYtIipHLb4Dggc3MP3HXcul6DZxJxO9KutGlnssBv8OnW3esXMcizgXMrpBGaZW8v89axa9SPr
o5G7LEUNTIbrqxe23IEjB4QsoAfULzDS+WAMKzAGqQE5mD9ik+1tgGYa8ZTFDA///6ZSmdhTSNUE
DFg5/BT0r43fxx64SZdCNGqLKkfaF2jvSS8PBaf4DptJEwvt7bT8NrrQhM62yjfHRjNNME+OkUkt
i/4zNvIQu1XYdYl3qxdQb7HOpwwGCTI52Sx/YXmn1mFe0PGU4LEWcEzvQBOv8FEoU6sLC80YubUa
8o0R4sUhPpmuz3vX9LbpGAvbmJHgjAlKk37Zdkm9qeERRylp1LD3KCibNelGF364pklll8fECy/Y
7L0vSSEs+jGGqOR7daIUenfUlTf2ssC1JEeLGgsOrubJRcdctyDJGL+wyrvaMuDo0LcDVBCua/0F
lM1cTE/P1IbMZniXQo8AXJWwXXvgTF4gK4MdqPelWIb3DmmcPDfUR1CvkqMReF9SooEojNvIOy3D
Oa/G3i7i8JxfN4wPTRNZgrqg6jyCFCPESqS6X64eXmeYrdzFtR3mUISGWbHo4swT9t3oXy9XnKTr
mLPvyuH1W/aloXBGqD+Ll2lsw/sdfiU5Jz2WC6fgK6eJdbHH1DMNjLzDjPBNqXzD9jL/m4sauXZm
tJvMCUSu+0wDoyIGqZZN5t8Vx5niv5eLvHdPEm7ZdRJme/djnTdpyDSKfEYa9cVU2LgxnIwuywFF
8ntbQJ1PhYzKzaT/dkruYpAYozT32aOPbnkJBVWnp0U2pNE995jgyz+luH06LgvAWnWm/Y3Mxi5Z
BH6pGjCJoZGD143XqhtQEatcZ3+QjJUukEUIvt9EFc7YcJbzOlGtToJng8FEEDa1OBzYOXocStah
7V3283NRgehOi4T6YdhwaS2/3a82omGRZiUJZiICN2x7X9KX0azTjsLV6Doza4HporWdy0RfabN+
MXUCua4e7INXHyDilY/2vKapd5LuYaTDS+t1foorxYuNQYdroFzGBCSb9CxPVwZGxPA8DQURSU8A
KGWl9QZcT6jfz+keO5Ao55LaMVOCrUSV5tX9JRiM4d8oMWY7XZOM7s7G6uN0a/XPxVOOysM7a4MX
6gox2UGOvJKUOkLWn1Ja7Mk3vkpLWYXd31yWMwb9+xRVyRkY9yAMiuTk1Oy2VX2y/dckoAW+0aLu
eyjujqhh1Eq69VzgzXL5q7pwd8KyPttRLqYHUxfST27c899XqLAFF/vuNBKbGJz4DNTv0zDL14oo
cMugJpj8hJcBkNpb9KdKFWj7sXCEEouGd23ZGUs6Xi6mu55Aasr8ST73zGtCM+9TZ9rAxP9lIK7t
AQ4dVesNgrRGQrrKk56bB+b6Ef80SVKUbZVvMIfs+rYHG4tm+AfQeqMItyM7yF5iaM2TUugnppXa
mr1xFVs3zDmHK4IlqgLYQqVlHmQys12G+6Rt+0s6vkxcnEFnccfXdyB7V6RU+OOM+cP8VHrI9RJd
w+oND32GmYOf8oOwY/qy7eSDK5y7mxKy5RhIJvvwCr9XqaRgwUaD8qskqUd6bg6dqU/WUEBp5xhC
Aj2ik0JxeY6QnwgckBcGFLuxKFMVMjIVXUvkQwq19peHkUQON5o/mvAQtp25wOJunNKsTI6VKVmt
lP53chByWYVyOBVUtZ2mGFymLxTEjt/9EIFhgJr0IZDa1BsB3OEtnPztBw75wkcUVsRwF85YKgUo
cY2xy9dLTxy8yfKSlrDo81Rau5aJulxnbqQX6ns1TiBkMLQkEkFuMzN0QR+xIAbcjNtlenT/xEzg
8yuqJuEhgkxZxfFmp0RvFq/er3QQNPp7QXaxFqTMgAwJ0R0+0pNMY4xhEd1kXQ4Cmi3jNFZI2c8B
frnB2+w3iIa4d1N7ZUF+hrs/TwnX/uUpF+tobsyJCzBil5Ja3rGIm3limoormz2NgbReBc4i7fnE
YaSuYMf+ZBOEoIm4CKCZFVFCcUtnYDtoLDzFkQJ6Hdy1mBIY2Xbzn0oHIs/cQUSnUpnXTlQTz7YX
KqdE9PG8sLIyW9Z8082H3nYz09ssnWq+S2inFu8UWqiG3Bsy4r+zDuk+4NwLE5SCTndlM+xCZnku
LEz7JCcqXhNxURAGCOeKtgOaBcRPclzuXMGc2DSP+b0WpEaX/c7k628OiXDewvjWFRhRi+7rMwno
hkFQaiOVipKUvVCYQ2nWVSnKZIwAVdJv+qOAGNLKfoKBblJL7GTU93AoIRlKYcrGcmxfJqsOhrnU
A4GnDu5sz0f0LSyEJ2BGY25NRl3RG36VMqYZKQRPss/THmQ8SpLmQzRNBWsSFXSNOGGpOnvtFpNG
h533fjXabRjkny1qDFnb3kVhR23OkOUFaZLkMZuE0Heuta5fghWDMfogn14Oa3Crw33A+OX5Lfgo
dBevjjJB8ilSA00AHqU/YNaBN9k7ucUm29ZJmV28p6AW5HQEIugQ+7vgHzowyun1xE2DQvuyfpnO
v4Tpp+xrUZRU/CDKZCDkCMiiF5gzSLs04FCdmqkuhBJHIGt6cKKGzZxrWYGQqZpFprKZSfDqIxfH
2ARZAPGGTpjKAOdjZYggl8CcGwYwUzmjhx+ckgJipS3YkwfB7uMbNinEhrxMg2+LM0LCFjpvRyRJ
85F2te3x4MZZIqFiJIWnk7nsTzPeZhHIDOzZj4JsAFJSXbSMoF2SDsnuUmylPaKgg7bXThScoOo2
AllBxoM+wlmJzVMI+Lvl+5PcKpppfyNG3cm8ju+7HYZO4SAPDmPC+4JEQ3hSLn0pveqfJdh7rPKI
oHZ6o2yT3UR0ErAGgIXhUcq9lZHOJ2zPGfnNQiMKMy5eZhcJwv6aKQ5UhUeXuH3ykwlE33CbuKIG
eXkgXqqavcAaU50u1ltSNwOeJJ+NN1H+sdD0fqQjsEmdKmInL4QFFiQQWQ6S76wW8ZcSJ1vzYQ05
o1JGWGqcXE9uzbrbyzLOxinAvrskN5M3FB3pGvuC7aaYLMESf4KJ6ajvpQXHoKS8wlVgG5+BtPr2
U562JTyrYLfOre4lIcfGghMjSKuIt5dm4qRQbBxvNjUFxFLv86mynDc2u+H3CTyl/JsKhOGYZf+f
I6gtVqsxTUI/ZYa2S84HyZZGqUaJIzKGz1KGXDkn3yRbrA/3xbou/iZf+AEYvWAUuqoLsiyeFUhS
dVCqsWbDsezGQGH0hoovw9zAzwlyRsJFQbwhlhjzCQlLcGmilY2ba2HcCF1aW9yW4EfeLoRkwh68
uSj35Y8c6ayJV3OqlN7j8pfIxKKjDxwxxoFvUqhqAAr0euM0NdcWMrxOHneafMHJ//GKM0DZBjp6
HlrJAx5TszSTs846Kob1fOTTb2fKOl8CpmX7T5yjWKkCKsve/II1FTlBVJGQmLZJKgmSQATrnO6N
beRCPj5eFIFbZtOC28Blnj5LXVh1FYFNUJCixDIEAet5Eqp5AkGgNeYsDJxscIA98o6Pl6f9VhFS
fXW3i5eBoldEAPUP2SFHrJwq+UwBvnYkiGiFDKlRYb3xRwaF3q5s/1CYkbBpoXO7rDgY77ZneCnG
NLXmWR/tBzMfSemBmFmZ41cbef6U0+6Y8+cbZtlNZ+qVkX2bGa8Nmu6zkVSYmzw+0XaFYiPkpWVN
SgV06mQMtQ1ghagg5xJKqtjY+zgV73T4PG7v3QXoIc+JFwelVDz6V64m2/2uwh0GoaqaVDtfcqUE
lvNBIPBOlU6P+0XkT8mbXKdIXf6Z/QzV84k7MBrXweKLdckFWvBXSx0QdTEOF1z4plMR2jMRC1S8
W9nfA0lrUtE1mDYVRwvATqeKcRy6qlDXfPQUqnUjlL/A/QW81y8WTiHqOhVnA//opzTvFiDDzJ4G
7rKldBFnYsg3zKzpnnGvhhyvTzlix2y4+I6paEQ8XSuFXHVEbhiADTTFbpNr6wnGTTFpl8H455x+
PjXPCVEao5pCjclTprbSFkbZpuL5sCs7Hy4Xu6IYWdfoEcdfPt+3nHA/hrr22FgMO6cGyXmdaBLf
EXmoqug1d/zHfLnXHK6ARpe4Eau3S8nUdQtNPjH6Rnn170h3wKod2Am5puUQV8S/lB56W3Zsogu4
Jj5JsEZu78qLwX2BtgrhMq4G4s8B//LrJZLz0RxZwwXEKE8hTz8ayFuXl7kEkafHEeked5i96Np1
uwIV2VhzHuqOMJFF6IE5Y8GCBN022MfkiDAAwSwOlDSzzLEontQHKYKyrcwbhMNW46MuUyG25Yga
XjE1zeeFX9dIW7AkzYqZuLp18ymhxxgfx7u2N9GI4JlMmAXNZQ41MOeE1yqIfbPizueTq+esgotJ
86LTR+bIYMfEu9BX2tPJ/tQna63qBYw6sFN34zD2RCKWMMauEbleHNUoHk0PyDwdmX+WR/S9Ck8d
jtsI6QqLCaNey8eno1EJX0btcixzPLBb2t27UI0zq/vgJ6S4G5ZyebJsf8o9J7com1Z5mLRfUWCQ
lPOpiilxN4uLYej/gOZGhMDrv2PkGe6NhzwttNlIukjOg0a8Ee2gt2Y5N10BWf0BMfTyIuafF/Fn
0lmu4VqvDmcUw48k9io1H40faMTLRB9V8SQjxbyjtdmz0puY7WggsvtidddRcm3B5ueb7ItC8wdF
Bm3tbZYuVq2bbymb97Q3+n6xNVdNP8aaTdXwnm/TW9hZoKLggOz4Of6uFblgSC4z4SUHXzK3oyMn
uqxvVgzSZGq19fTsFzimZzwxn25/h7J1JYNL9BQcRJUFCscN2qRy+BOz42f7NpqkH5MZXw1PriJZ
JKbFQeStZ1egiaa73Hx0uLi+ejL5wtbkVtyEI/3u4vKO5aBU7MEgsaN7iSuIQa9QBnMe0TXuMy2b
7DoSYJK7Z05GYH2HeBvkObbBpIeNsAhf1hzdAZIka7r8DGZN7gT+BAnXwpFM3Yghfr0vw0b0ObHg
Nbka+NPgvWoADruRZNchYHG/2BXLxeUAI5R9sdb1ptVBYr1cf2gKXPOHox45CbLejE9sW/ixIP23
CuHYcSk4w9dtrYlg9cAmJwY8Copb88JVxFbq/NVXQjTwcr+8tPszkAOlNu5gmmDyB4XWuelcWKbx
REToJAij7FI7dOgD+Yh3Lv8N0IzHtAtj2rdO+3aBAkBaQ9GPHpNmXXCXiHZlWUzLZjKt6/zFMzRI
pfd5XH/OYEfuNQRkJ20tocVqisspyEqnEJAEnWWZ0qUTXF0J4Jgm323qt9CfJvgJWUPpXvatPWEV
qauZOCAXaM7sf1l6uc5EvIjSybZhVF4Hrsw/A+DHCBhbIcvqE0nWMyC3r4MoPDpJ0DOqgACWbz3c
P8CxYHJkCBO1vafckUu6ygSKhKzA2avwpX9zMS8hkP/kztI/TmUBzSn5PlG/BgF465Jy8mvn5OpB
mvc82O9j3EpNj3f9ToyCNHVps2E+7iwuMQjknO/fbOh9bK4ZYmPhyDJ11VpghCts8ULan54e6qQS
D7s8KJA4heLj5PgAEzZJhachEX+oxgp/sM8QTiEVl773D8VZqtoK0lvJxB5zT8gjDtpt+ASBUTl5
48MNAPa/sXxQcufGNWkV0NOMrDDmLoi+iXpwFAeq1EwABpYiFcl8zotzfAvOoIfwlP76SDrbY87+
wP37etuj/l1xm8zkN7Y1ZKZYWWVdJDSXWUEL+9iJbpUXImEtNMn4Ne25IieOaEtLztzHdwY+htgw
vWhiBVSBXCwg75MMOaj7HmohZgb7A+GxKf2lRu1+44sVHsGei+cGlpV94nWhZ9eVwB6w6RlUHFEi
C3Ndk3YQyOrLE5AEqO9VBZlSBaXwriglv8DQTiqVPgBjWhQYweZ/yRbzKYRrNPAyGALj9drdiSa8
gK6toJkbdfql8J71/5TMUmhKl9er/KWezrGPxp7sSe2LLo6MFo6Wq0GN2BsVTcm06mHEZR0gjkoG
7MnOFEuROtX3yfwb/JuIFrMJpySCj/FYRbOnVnrHneuHeSdtuAk19CFFICrmLNM7tIVchbArlLm3
lwRHZOdC1VDLKCOa6K48TQiFfpzbGoTTjfqmEC2NgSD1yAY8vih9tiFVsCthF4B+QTMHpIj+9v2e
ehCOVdh89sQx5g7E3SKxbR0Rl1ZAfKyiNGHPK5mAm8tLwIb32iltti8YFMW40rk7wvwXjPXcj0jI
kU7WN5yz8hht7B5hrgLECjAeROpl2mx0ew34RuJSXLRTQT5pgTHB68lLvnMcDHpi8kq7oDAY2pF6
m0r2sIRrAYeumIinyftavgUotGVxNJ9eF55KC3hPiKSvN/KSHgv3RUlTfHcUga5u9MtEUmXEKJA9
T54LKoBKZAV8r3T8SMo9rTf6/dHLd07SWttmhyDTQFug5fKnfkCTlBKTUnj89yaj1mnKniQLHryu
7/LIcmWny0sgdIwn7Az/eNAmUnQ+6DrzJVCOb7EJITYnW1nEiwNUeIC2T0bYXNOib1H3E5axEaY2
N428JxRJTYVVT1Mrwcv9RlZ8L9t/1rRjDih2vopMKRPckoBYsatBa83WR17IK+KusCOAoGuSMokx
MdtdNk6gEzjvFfomT+4ZbCfJkQ6OyV3wqelYs0sPGYnNmkrmx4hyFpdoleyDMByCFyNIdv7s0NMf
G0qFq0QMzUYaiZ5eoJPxVVT3LQTHKPnoJKessMad2QC3MBczVkIGTw7BTn8HW/Zw7rSz2AY1kSOZ
9Jvr4qU6v+3sr5UpZX4SpwQvdUIjawi8URGdZYEt9rleJsq9QW/KS4jaqle+4T+q/D+xIGbi55Pz
XXK4H9a8WEK/dSrC5v0iCcupQHMa7ryA1Z+YRoRHC/jkqKRhpMm75ekqbCF70+jprcqMjmSAPYXD
o0XURuXDVU5T8opb8il8s82XyNAjFajjHNS4wIiJf48I9gb2oo5JMyW2N4oTiqb+vAsJ9hftMIPS
99vMsP+Km5iKzystq2ZdKtzD9LdXw/a4P81XFRzkdB5xYzkS1LY4JC8pDYD4lqoGSekSP/7QZh6U
pf63LRdL/oWv0I0I323RF1TbZViTxgcui9sah8NG5EnrpA/TYKCmo0KTXcnNd49UnQvyXOEcriR0
h8i1w3q4BDqCGQROo/xbb2rM56jYnEDQ3M2H2Xjf4RD05Fy2AArjuBpGbsMvluiLCjA273IbNoA0
X7G3DblVWN+Mzj8vEfPePvFxDESGrm337yTVEEI2IFFnGdLEfcpF9zjSWqVkTc3rFrvApJZdUTJ2
imcUbOVa7kJzeOEBrkBfVXgTtHBYp49Imk+Uih278wnyfoIGQcpZ3hxA5rcT56Fxc4npDQS2RiwB
P4Wp5Wc3ZYSjCRQbnUVHE7YDJxwdRAQDscHHpYFGcucPpQQLT+qKQqpMly3uPzYze2fMfyUOCF68
OqbZakVZjRbZP8CJ4HCrfm9oQj9kSRYI11B1GZMaVqiu8KIgUs0pHw/6mfWyAKqiQrJIahILcNnB
dDGBBy5z1yB/xTjDPtJfRVaBM/DwLCxhDXg6rKjw9aum2XrtPAn3AzyS563YEagOsGGxLx3ofAsm
w8SXSA0CZEhbVlw+Eo3huTpIJLwJbNynFVp7sZ5xzRW7EI8XsYyfY0SmJVpfbDk4dutxV4BqWopm
3mhpakCuyrWYf/mUqZULZFhcEzVH6LGVvzb8EYf+0kooEaggwkx0UTXJkEwn4iOt92XOd2mQC8ql
MRdwyQzbBeXENZlkM+qAv3jz8JdxCAhoAorA4UZmVbZimUty+jQZPaDrF/MKbrNdD5O5jMCQENs8
8kY6KPwjHoeZovyFGdkZHN1QWbKmYyJOrCQa0/47JU5Fx29vCqfGFSIVZ1dRmCTPCc21UHfcEMgN
clUFVuM/iYh2gMwUYxvX4Q2i817K9mZqWIRF3RxhYB7O/jGn4ms5rRD2G7mt2k5WbZrHtHTfwn1D
piDCM5xA/aDBFzInblSS7XuSzgrVU+wz64hyWIMT/Th/nRGs+1DNDTO3VAAfmbq/ikveD9HwaEzl
YzR2ywFXsFJTrvOIVaYs1FOEcpOkEhK9T1qESWMGWg4tiJRtqu5zgXtrIcdN/y8s6JZLftM1lq9x
AiHVTxClmnWrlHwkySO9CuAcbKY93uJF56OlGQ/WrEN8fD7+UqCXGeh2DtjxJOsjj+2MhH75ipz9
aOlY9REH2XaBzAOQqagIw68y55nrKpLtqsgXw1Hx2MpcvWjC+9bNlWtxi8IvReY498KilXJ8E0Rl
vpNKSpg3nWNI1LN9sK68zJ0f92CdX4rxla/IedvKVBxQLMVOzt2LsqwixaYP2lzl7QwbQGeGPteB
Egw9jBdLggYGd733/cvFwIu79oQoDWrW5pMs2e6QhUSWSLbGUmGbU75ygwvayMkJg8hRAr5G/FN6
OJTeE3h/Ky+lumOqCGSEwyIvTM66EuC9a0YNh3adBcm5SlC26Z8LBKOdd23O8c0PHK0DEKard8oE
1j1dlmPhQx06RK7nmpILNQzDJbz0qV0dyc5/w+cpXyRAvw4iGaHzf2cW97UphZmHRShs+cSzd+d0
0Tc8Yh8BAhConX6NsbeoXZY8LBacn960C1WohzJhKWUlrotZAvvZxV9VXFq5/0bxomEI2Cit4Lx5
Lfx6VLD9JM+YKG+hohPbIHQeaQr+fzDwc6cLhrM15BdPUqbpAJl9DWie45hXs2rW0K6XwEcWPtA7
4Y4SBtwjhW462qkvpb45jU9dNJ5pcNaCClbUuE7K9TCtMMu21D18Nxg4MCHLO9HhMFDmuR5UvCIH
pe50DhnIc8QPwxEOMXYOyWIMTC95W8xhQRMiXO/BwfnX2ON0VenOzuSp9ga83+t82T7cv4UR3sKZ
uPNEuvJlZqx/Flg+X73yvyH2dSeanlGedk9/PQwe9orEXEl3ULu0bhaXW3FMG6y7NHxZXyUyJKzz
tA1IaVr/AD6eIRr7XNmItPhLMmaXUaqVmlnFEBhwhypHJfQeaXY9LWcy1FVytoMhFZv3lB8zDxXI
oVoMHNFlo2xLVSkcEjfMunROrjupUPycO3JcgVt7v3oT2fBOmv+YmCVUpg3v3rPobOPTA1RJxm4p
MRoLJqvly0XrMgcAuyh5epmc8FqE1+gDEEXPNgSvUEYwmO8Xweua4GMG6hvHzgAs/iG++Q9++6od
bDoQ9EOjidZSezW7WOJcicrohykbc14ARb+LbAU+XEkLWzOAxwlYAT6lYu+BzhGLgrSG3n3jvk5s
FfFtufTZsa1DxNkyc8rO98CB7bca5tv/IZW35Xsugy3kiIPzN5lm6kcbH3rLQAUhBjddSq8IG/JJ
EGiw1hKfJu3pPYaZNWYbI0r094KpMhM/8zOxgzHmpXr8IGTdEiblsLcqfORmbUshSx6nvE5VcvZJ
+faVJYj68JV5JQNn/xqjqak1P7Vsv5vhS3cHsBBtEHtf6KpDnG3S3SfZX6K75lJxjJKtyhMu1Oqb
EJDzj++rrjpxJcxjZ/+GLg1aGGrmyi5t2AOO6vHPsgzgWTg4dH9hPrg68SrxIYqq42mRb7+oorCo
jSZwvC0DD+XaSp726ZXaOPVBGQVqCMPNtGbf7mx6Ou60OKV5pE078M+RNOtmXtYcwxloGd6VUW+J
A+YdjVWaT/NEsGTeeLIKk0BA+6z93UaNztlxO6Gk2Jp5O5VsOAW4XHJt/KgYQ/qUh/mR8PFJIcS2
EVBedmjuS4d7e4cl8KFYwKyr+lQf+1BDjdVuN3pCk/vSaqT1NoBq3kuHrtPVA+W5invAIN7MpMLE
O6F6aeiCzzEoTYqbUgh0FnumxwTNf2u4OG1ZZ4cxmh9svn+7xyH8fIz8gGj7PrwIboseUOJorwnO
Pz/K2z0xcmATIDpkmf2+dfsOnOJUs1xpTQn/kwPRVf165gkGh7M+y9YU+eHznSvWj82kjvw9Xb/h
LJq9TskMMQDBTEYn0fhfaT1kwEwmDGEHKFuBOyb7ItKleU3D0hVOtuL+FGHnzNhOxF70hcRNDhvP
LArMPix2PH6A5SbWRZQ2iK9Rvkq8SN5iyfFWn5Ba1tUQYAgDosnZqmRl3g/LGRGKw0xvtqCzjXz3
CFzhD/qw1qvXfsK8aP4WlDhGuaGLDqlEqRNDxkL6MAbMogH49C+9ODn9eqi5gVZZ1xE9ZyzkOH/0
pHzf0hhMowzOVYxOea7+7jA/BEawzbX9y2LKvmBvH98TkqJhuz2LztqMvesMj7iGq/bLndD26m/I
i6cJtRDy04ygKW8Ws5fViKCHxu1WEJixBJrjZqVBqVLfSTIAqn/PhL3H6O3x2DygaSMiqrE2ImiK
8wF/sW0OtSzv5NTxm44vZnEAZZZIUb6MxRt7cVwt8fx4WgRbNwV1AZuoIBAJZrqqY7mlNchREB8k
Xdi753Pz8gBbBAWiuYf856/TEdyWIaV5SwKDVbXItTw1poWN2iqmxK8o4pAR7hBDSptVbo/rBmWV
84wKpJ96Z3LZfBe/OT9ELL5p3zb6bBoDwG/wZPaqcCCCsO1QzOFIy9TbpxeyQ6vZKIc7ZR0BDL5c
aZnwVeg7D5lpO1HPd2lHJMN65E3sq4a4++L+mmunOHrgPoH3y5PDg3+yHEsC6cLfs5NE6eG11ABi
wl61LgEAcpB0V4pq96bVAhZegGFH3O71KrmCrWKnsGusVGmJf3PRQ6UIzgicgbrnpSiM+LmrJdX7
7K4EXsnxhgXXlzyWaPARMRzQUQIuUcvYD14vsONuVkczDX1s8aBb8CJXSxXxFu0WR2/wUQKfCm4M
tzTjGjBjSz74vgSZeTfNm21byfrL2wLyJ8J8uBkWbe+f/GgG5AMrXLsTI7Gdit+LKJE0Mfm9Jclg
jGloGujt4wFoYNmPv8zN68g2H52A7LQ9PRXPLf+/dte0v+/2ua2yn1MAl4kLLlwuklCKF/8Hsi6m
T4k8+r1k1t9sbuZxtLr05kTd+QHgY11fQ20nmPHTAvz0tpL6Om8L+wDis2RcMyVVVD2jwMcOeyAK
1d2ORM7GP0vtkEl9Hl8yhW40pN7PkLPWipB/QrgBfu9pmkN6SWiq0HpSdKOlLBR5lMmcQgq5otcv
9zoi/tloefiStv/l8iqiZB9UxIVAD+3hSgfWcfJGq9ZHmraZcVKXQcOKW08FgawzjBChfjv0K2+B
ekTgz3O0QHzkcTz8420qrctHJCNb2rkjM0iVRyNTbhdPQXxUzPC4/srvYg4ixvZzJv/4Q3kuQHCG
3JzVjPVrv0X7+WEiTvEnvhtGAENiB0q3R7JUyOuPC2wIzL/J/gH55a3X/1oXtSAsA+w5b4O5pPyX
o7wcZyaJMlHISDSUMs7S/MkqGxOa47wDjgH0ywVMu3ulvRIEoHDNvoAAc/nkD7C4vLvMPEr1juM1
CUkgJZ8KJn4rOXlLArka4BlR7mmaVdF76xndeNshPUIk/UIm0BeFiZ7hWdH0PcrYRQdf/LDm2kMt
iejpwC/MgQKtxMuIPQQ4dPTPJuy7nceWZhAk8sAttPQAPrgE10jRcikAY9am5lNF4Kz6h5Pym+RE
k+OtxA9vqnjmgJiL9WuL0RD+oWzA/3gmDfBjykV0urN8NkvkyYo/W8NsGC3/HpeOzUsSrEeLbIYj
Q/uuMm8nAuqHByXO0UCtaFXL1wNLR/P53GSZNAT6GPhQTgP5b3Zr7hluJkzZndBRI1JTCA4pZs9A
kkftOrnwFltjO/IS+YB6jBfERvtu4DvDzUBiEEDqVq/GOw7DQGJ3sV/GChYD7Pb1yhuYELhq9YsX
xTPUBCBJZ9qj5LVrobFfcEpJggg4POqkt38acyTgu9NNb76n/Pz/HIzB1tqBgoVNonen11q03c5a
hD5zjuzoL/sOgJYI1RjIpL1U2nMOZHBqLoYNCg0I5lNODQTa0R2KPAHoM0S7IA+EQXugio6O9MnY
izvVVwyglveHbI171TPByj1blekJaxaRe7Zfh19emUbmLJg/K54Co1wNuVsnY+8IM7yOOGJ1+Bfr
KyAF2hyXLt3dzr3sk0rySAaoAi73x1BRTqW+7JqMwCTnbx9kF6Z1Z9RWIFzzLo2xV0/KMAYDycPL
6UG2k5nuoM1qNc88h1b93zEFSn0teV13JmxWUO5JDhBQcSKtfeyvqToQ7PIy5u6ugwP8+7ixzoJd
LNVSKqA0GDjSHxQv13Vz7cwhzKvNiw6ftNX6nnFL9x+IpUYBpZs0lVWV0Vs4zKcQTwMJHYlGJADH
uWaAirkzY/DOXHJqbLU6LT3CxEKMSVUhcqkZO1pdHcBqdxV4xWwgeX+6aqCEFB2WHOPho70YAxMM
/Dr/fHqrfgJWBuOlgiiZ/R1rT5hBW0JgK5Yf79XEugupdFRdoUWujXqlrgDtROEqyfke4DHjG8Hu
dTbZx/nSY/LfmHU3klpBShdACh/AWnCCqKwJ+YzbyKHzET8e+9Bu7ZNBAY8jB7NVvwLoqW0td/jR
DNGQXV2h36J7Ip/MPF7W05XUwbovEAFzPpDlahLaOP4NxAaieakr/43EEB/+7q2jssG4zOn2+gj5
U3d/iVKOlcPZAeDtYjwtHjLQBPzCxnxq1D4gKcyk0BzwC9L47M4HPYzGD2N3DvHHAeFCLWUI6QBt
OWnbxBN8iCEEfcB/olGFHCgwl6vcMiY913ZxxlT9qxsm1y/jG+Xvb6kRR8sKn8OXRbObpgxXqLlS
tA65NxT0IM310WWPYCOGZdnCJJr4K9S7oFb/EhvZRlootmlHeHta9VkA0b6v7ncLwnNfgdSH0qLT
HKrSnqPBP39KYQE7HpPSKxJx91ifDJjewhVI4gLrLnQgrCAM0UNI+XcHYwGq5DBAjZzhPfEadfFE
logCfYiMbFqKxMf13aX9PRNrt5xyuThpABodGcc9LULFhgyxrXnAVC7wlN9hMnZTgDQrJdrWEC8c
knHrDPPjIfeJeLvS3KJfNe2l6TsVbnWgiq2HF5SchhjfBjllG11/g5VKpfsg9RuB14PsglG1KAVt
xt0EAlh1cBz8ku4CJW3K55Axa6cksoPoTp15dOIOboIquCOWaze47skxUNNM7ETGr1GGlcHikeDH
4PytotN6sYx965EP5PfYzLzRiQ8ylvJqSzZwVXb9M0RzPiBKY+sIBwYh8p7IOsr7KgbB9HUDohv8
nncj1uaoEkj8boaS5QgZI8RQaAZmJwCicG1qyInBXDIeuu5aGvETnCnxqJwt9y30XmPrRHzciDb5
C1f3zAxZmMorlDshbw8cm/zXRsK1WKA6XwhDZY0Mo7j+u1b/4qNR8tC8igHKQTM8GbJcta4PZ2/K
pQEOrs60awksnoDo0BSJkILFyeXntxtDh9ZMFy3FbmTWUG2u0d/yefcSAQauBxzMFHNG06y8NhyW
VUJrkCvOJbjL+/aZsBQzVs3dWXkpYh3GIDjCkp/jt65/YiOTCTEX7qO6SmOCzdhWuM2JOfz+FPej
eIeAD3B6qYKBhmn9HtGFEKqa+gYk429fYBnrAHJdaNP/F0cNPIVCnr1EebN1+udEq06alxa3bGuO
zoO/mL3gVQqxQBd27rEpX3CZUDNdoweYfxfeC2jHGDfO9vh2hNeLFZ49uTdi+aMAB6DkTNeYAAmN
0nosRcMpHPPGO8RDt6ctXPtN1ashcBAjM3RyTfZGYilOeoTFLDFV3rFv2PBdgmDc3M9VobYMhcoE
9nEUE9AL2YMSH5Dx/2xPHQ1JMYDnKQIeaTkKTll/jpSIDe9NZloUBuTIRLW3OhF0m1PbVy6+YoMW
Db1Edr7dSJGQWovm/Ga3j6ZV9iB7hfRpWFQE5uTyExCgtDV+3BKhj/Pzt4Vkv3L+vJXhH5ePOeD0
Jq6H+jrQEe1UAFufoFbHhRuTd4ETYANlo0jp8ZT9pP2+kK/6AVcC4UULVtxv7dY6yF5X21MnD2zZ
c7xzQ49/5modEVy/uU8XZuhSHFD0UjziY+8CLqnUv+vqQ1rJhSztlWmKi0a0INAahIo5Xx30sztN
SHuT2wS/RcgERkNgFiUBYhZVZmNHaT++UDpFMC3x41ELRlUeecQT/qFOwnpvfluN4e5LLx2gqWQR
qCYTnVkBgldJOVEyHsycKJcDNhgImeaALju7WiFjJNaE5b+Gd3T9qZL50jJURjPcvGBqCLLY3H/U
AskUSqoIjVMqWoEL9oiucqTXYa+C6JRC8XSeJLw17WZRw+nirzSjEHIBJV8zyU8s24w+aMEroYs4
22tNF8vQzQvaa6rMe+0kIIkC7zigt9ZC5Ggt7ljf286OedA+g3CWgsWkJoDGKYiZsmUc5lupuMQ9
g5YzP8On2vTKfXvClj6KGViW2zWScEJncDAV5ddew45FBrWoqvByEIReowG/nVTeVxkpsAnSe8KX
9CNdVh1KITT+I4JFPAG6U/EFSPx3iebLWVF4YN70TNfSUAwe72LOt2qatXcne4yG+LeV7IT9fnTO
tW0+u2XGFRlIqQ6VLE1E6lMzUaLGPFPt9ZPEv+DK37t0mX01ybYtaerIrqPy0IDvcnOLiwh+SS73
l/CUp/X+ucvKDksw40QkzOhy2UeyH3azAycag54oqMw6DUyb7epJGfN0MNIWX/jjHEPGQ+9WcLqK
4rMpt+qIl37MX515REDXfxdqDlDRUgo1ijWxwx9QtrtbXUbVWgj5kT+3levXpCA9rgMKzTGcXGwG
EwQp+jpxGCZyhcBlu/eR3AXK4A0EdzOF2QLm+eBy0eniBDY+k+/tgtuAjJnDMJoj3AjC2uPzzeZJ
FpXZSFLKSlCMwHfeNPciY0NoxTET35QF1X9VMA8YeFX3k/EpJeYh/1kHpHI9ZaScp6DFnApD56KN
MZDx8feOCAJpMsq7hR6riT/eSzkbBf1FXQAxVeMfEeOjtBc2tdd00VnieN8XznunAZE6SoLrG6nl
/1R5R1bY7/LdewGP4h0nNChfJsftLuKzMXj5kgRQKr3JciFsPexfMJDA/vaGa6Tz3QtbfoFLg9SM
Nj/N9m/ChkWndXc5icwQxcmm1qpZilcc0SwCqFSGd1WxEu1ZBZDcWfPmpZoJNY/S9XCX8a0mCWTI
19dCnIO37NdXS7AwBTXlyLI4anZQKS5HW2uIJEHdh2aARxvOU4Kc2JlgEBfyT+gJBF0O/JVLzkZ7
U4l0F0Ne2wC9Lt0flLXavMW3KhvJfNSDBN8B2LsLbLOKHKBp0faIsmFbKggDZiDuQMbOLr8sJWzW
wjpX/AZzZjDiEKwWgdFvTa8htDfTDXH8FCwuGhmqBFums5QPNxLOCWBxuWENRgHtbMJyIsyIX93h
y7HzNLBqYnuRpBPrZaKTbhpyNiyRHM8pIhzdAXeeF0tiRldw4L1TH2CwIe84hFCOwqR/oTGHtjle
6CjsQm27ZrgK4QD6gZxFh+5jtimik9/Y4m2EGIe6wLCINVqlFmPKiRuWYWbtqAdOgq8RVBuXllwg
WrfHUdpwEhuwBce55mp3UhTgfkVQG3bc4GD3+NUzF/bUVTBbNwVVLu0i94RB86QXaAzpIambvhbm
eZUVSNF+NSja+QTiYXKIrJdXGqhpjzuFn1EwEwCjFSP31tzxPoShNdC8yFL/I+WXtTI1g0lPI6ki
k9+IAoBmwZxNd530slRae6X9h4lE4Xu2m31ZjzK8Z0dVaHYPcyI4hht+n99JGO5JnhJHNLAgyhEI
WKlScF8nOTNsqm36k4SWaAS1RosrUhyP39zKPuJ21UkWOK5CVAml9jaIdIejsU38clDK4Em1CVdc
wODX7Ir6JlB3BynEYMtgQsVBCsbqhtlJ8FujdoSuJoeL7JoH4tPAEweaUjiKImSBEr6Rf0ueu7Io
ojOGzun0YUnwFd5YtgPV39x7RrrMsv5AcjWdysYhcSjV4LX37OH8DfKqdesDKd5+1ZdWjXdELRlF
kLO7IIkkEzDdHdXcKMa4CdObtZKE69XAOudB8plbJaTpLgMODj0+CPLi6hyEA32cSNR7snfSt34U
QuG/ehSbsbZqy3JTz0TpN7PFmbIRfeqkmdtz9lvhc2ulFG3wxjB+YPFfBASKSwBIiFjhDWrA79So
xSjLxCKHIP/1x4PasDn+XqN9cW0JiXKmKEc/z084SbwGPXEN3/CviWBJQUQZ9MSxwfp3qhEpPhrT
7XtMGKIWb2A2o7EgL5oby/JBTVfHscwlVKJ7O4yrQv0aoLIwjpayyBD016h6QKZjl1leP5pgDmed
0fxkseaZy+/9vAxvFbjousXhZTEhHHSwBsjeITNK270BO5VaSprMomFO5hkhH55DzC5dK83OW5y0
yhMtMxyrutFFYHDRLxjUZ90ahpXvZr4pwcOPW9Eky4g18pNAO576AXUzJjAZ8XI60X6VIuP/VOZq
OhnKlbuwwUY44U/RB/oDaKYoqUSdq0sVxR3OD1MbaxEanuWgzC7Q8tyG8Wx+ywsB7/IW4sZBPApv
1x8tU6QPRwTx+Pn1s9JrnK81n5bMjYbyQSQCfMDpAcep+UGciHakyq8WbUmy/x7MgzTDmterSUcU
jSY3o3zELrT05KvibV6yAAkwHxOoDW6O9lB8NaoF3dSlvEd7woz6yVrnNWUZ4rX/UYP9ZR/KbHIH
hc55U3kBzNAmEN22g/C+K8Qd+J3jUDh6aMWzPieyVMpclwxB2Z3ymyAEnI2uocurA06J9U7mzA2c
UqQUQKzpLPMlnu63TJh7tvkD0fLIfya1hhqHvuz8IOtauyxNzp7b3qrCKi7YkDXgE53jM8XAxN4L
IdXJwY5D1DM3L+5dYSlNY2IoB/piQNvdGSqcnQV2YVpzWrhNYFt92idLh1D7mHOk5RkGBx4qpbk/
zc84jz9axKCCJmNiSqp6hrNYF3JzUFVqJsSP/j+mOHYFErf/LHcOahrf2dCxquM1CmdAA5y9B2Ko
Oi5/mQZqrFhVGZGyi7Usnu4L+WlOSunyQwzitrAdI/XxBkPKuuBaca2YrpItI6flwATKFUgXJwEc
plkfHPn+O6hKNn+2D4ZQbmSv/QK28WV4iiguO33V/ILgYOhGTJNzcY9yLht1wJvE0WAc3pb3ci6E
btEzfw11HBqGZnCakZ0/HwyI7U2tkJIIAsDX6yk/4iJ1jWKMs9YefvXAy28ffeemwTNvEJ9cpzni
VsZKUWl3Td8SwDFJWpsmmEG9aGxgwo1zoDTR93vrGKucajp9exk6OHJw0aPOmrnoY0Z03s+P86dw
x7LmA3gCeKU4sXqiGP7aP1X/1GfHr85EvD449zzxI8Q0b1gEEJGbbMkGiFKcVufSiD647pjYaBud
N9gTg4So5rASg2MCZfHNCD0+kVwykGossc2VeC3lS3NzWdkgd6aK+ssuAlqyKKGtBDcwWT9A4pBh
4ouHLRQEcaB25rxdKkM+9Oc4ZGf8R1mXVM0GbtPK3saMpqFVslUeixsU/R4JxIR7FnX66L6boilE
OR0rKGwmKLpCnw+uc2P/40KAvg0H4x2ceUBeJou0OYKw6CxZ7xvPoDLv3SLkLuonPYk9Cqiy/R6z
gaQiWeAX39jKND6o7Xint3z8ApSD8SasBAo5AMasdkYhUQU3OEv26DNZng7VxF8mK9O2TJd/XTqo
tMR8kM96CpAaC4QuwcrCAQZbx683ESKVkNsXLZqpvcjqElk6xKvU6pwRWWVyhCy3QbgmwqIEOL+/
uktJH7a73U4TdGlIdbtkfyHnngUviW6HgrOT+BHFocw276DHDeyyMOKP77nF5KZujhilTl8NFmki
LI7RRj8tEmzSYx1CW6hvqhR75LFVQ3ZGohY+g4ea0awFaQApl5c5fdCmghs23K6crYvLytD/W3vk
rWF1BDBgOpABTM8QLxbJFLCyfMhUFXAM5MGF7JNB8GFTgwrlJd1trKRVq/rGVcEq2eSLtdaZQ7M+
iiSXKSbBnWcp7FLsQAwqkw/hjRjX5xKsoyj90BsJXY8QuspfWTTBHZJUyvuLKLTpccTEv7PMwe7m
9sit7YyxJtfgh1UM93g0UIsxPhShc6sI08QpW57edq0yYtMlW1iIHMiaiwzGYqBgYo/E2Xb1zxWI
PzRCXsokDRUPmCJLJXA5UxVAhapx7FC5elgRL7ObruUdnTz61yNh/MHt4TfYz8aD8nQ/JLLtXcNr
KsuwTsP8dqSZg9mpPNq7zybn0WCJCjryP3emXjSX+Wba4xvxe3AorQbBDr8sROEIAq0rGrWftT5j
brEStsC7NJBf+ukjzZNrR5OhoD9duNZKdUMZpfpnJN4MSfFKW2ZIjaqcjySSTy6NAx3IZbQiJBsj
J2TTz0fekXoHwIOtYnZF5e4xaS+OrcJDkWiQwtry578VA9l71mpeBAU7m7HNTYLZBw2A7N6SHBdA
H+oNYo9ZzX3THrLh7HW0bCalguAarDIBxIjswV5d3yFX2sRRV2iEEYhGGdjH9XOKhVw47A8i55qo
YGS66XNejUkLDh+oxo7qvTOSxQ/X1nQDtyRw70TDuEFOdAxzX8qxDNJING0pfD3lWn3DtM3pkV5Y
6pMfsUUwLB1qfzqCU3+AZm/OUhB9+hZwpCaHjrZs9bt8UTVxJHhuI/QoZVdHB4aG+nYJAKz8LxWv
2mhScMtnmcHvNocy62V1GlcnKwN09s2q6Cgg1NKFxvPa8rgcBMr0lPEXPQoFm5oBGmoRzj9HKxRS
DgnfJ0TPoNKn/nGI7EbGqWFZWiY3Kp7UxtZ3vDOmwFYUGe9xRY/Lpsy8AKo9JizG91ycZgkSiypj
58qQpJmF1iEl4c/rME84hJN7VlDKOUmRmZvvVRZOD1ROd8MqKYGOLqQbsV5+Aqe3+P4pTX6IEmSK
3Y4QW2eyXcOAL2ursWmxj/7opKtvXZ+tGd5PhCho1NLSquaAT3pNES0s69E7rvoXW1wyd9qK+MXE
67S1VORAm6VjV4NHkJ4smT3SNGWFykk0hLcRcMclxvCS2BSDdVgE6eC4jl/Awaf/aRRBBkDz4tek
JR/yb3dqLboFGumDbpvnlfiT2KGzjHlTnO+2joH5AQZEv3jx1Mo8ElMNEmk/Nk/p3jQjadqtVfGE
TwUpC/zysqkljtw36s+kkU/39O5TKjiKBn416a+V876zwK8+4wxhVbNB/CXM+IBgEPoxy952PuTM
DwcBHZ7kgqjdHtU0vQHVnS4vVS6STAVmW0OxKOcVbLhrnH+rd2NeIkGZ4Y62M6LXp0nu5zaR9gHg
hvB4NdTddgbKsssW/a1IsMQX1hiNt3PzYRwpA6swsadqFC4qxHb9J9Z1updT0Av8xhMo9dWZcNyG
JHSojtj/I+084lSmaKyVCotqx9TXzcRf0ZMeoAWFaICEn3MpzOrTPDgS9cusGJbq/RPXZCqeneO9
pGyuJl7OwU/lX94e2/rRyhoHhvZ8c74lMTmXJV08YV4GXifgXfCheaiKX2hAuxuWYlP4BnJyZQBi
kp2d1Rid6C3f8IKE0KnOE0UNkNiWppSc0eEqNmZg5U4x511WaYVqXoySJ8lljcQ/ZO1UVm8NX7bH
WIsXqv5BvPgMwPCFaP22KKl99T2YgMuo6H4kh5KXYodsNQn4WWOHIAoJKpelGqTRTa+FZ4swOyi5
7RbhXe+3DqMqoGGOQDGpdz2DZxd3/m2pXp0MfW6qbeYgAu9VFtbkiRVt6WvHNVZVuMl2ZUBgdHOl
olpxjR1O7mTmGucT1Pj8Rrs8t+i/ha7AueMWP0SYsBa7IVLcru5dwYC/lxR2eZSta+LBrs/CG29B
0QgcVcZR4m2b9E9dvYK9zmyuRq8kXpj1e4OBWhRMsF+8B5LxzHO4e2yzm2mov5ZTeUuRM7hbOKVn
ScUVB8G28xVmdXPseI3R6TeXordGCy4FOEkKYitYcVj4B/UljFpEynfWUdi/5Zx7PbWYRf6+a1JM
JRvWYlF1idzMj+SYmi7XL8Wf0/YQVOcHxN96L8SVL+k+aBiHEX5wrQBwKPHoxLmrK+8w1AfijLeV
9fRX4dUw9or4jflOy+/y8mbZ1ptVkeUZubEYxgnoaG5D/l7LzydxDe8Yta6zE9G1pPL/gweJ5Lv/
fkRUdGhAaKohJ+2i8g8aFWATCvFL2kr9RvS145h6txGAwqsY735HrvN7JLUWGNz8hSxlJ5l1rMNF
76AYxtsoA+aGRCRRjICWePmOAb3m5K3W2My+CpF3vkgqljWhKUrjg4fZWYyYqfwpekr/3RmJl/Dg
9ny402KX+K8FOns03iVOStnaKA0p7iqezLYoo7NrfctqXUNN5FcHr3sWFJ7VCrvrQvU80A2g3ozw
8AseakCaGUOv2QlwHaBADgQqI53DtnHt0LaL3P3brwE2FlQcJx7bQyUJyiT9UH8LAIptnMuHx9fp
XDlY/i2RNiRfRH2UK0rXj5SRAcWq35w86aUwlhOOXfNbqLmh7kONRoNVcMd9LyFsVv6DbGK8SGpQ
zqf7nyjoMcA8MClmaYsk0HEezTPvliBHqsKQu81bkN1qzBKrz57ylaPCMdHiHPI0+IF0ab92ctet
7ljQAfkYPUHQMZFv8B6chBMA6NBJQL0GtkawYs29iZbFhAi+FV96CyF+eh8hbC9qk4jpVN70YB+A
EX/X00C6ZByTvawUGBz2zkSkzdmMzYukNmz3XOi0LAZqV+/5uGQiu/ZmU8JardqLGKOyRJ0eiXcj
Hya/CEWj7rCuj4L/mZf27JCPRUh/m8XTbhy/LEeoWCinMgFHN5uM/5wlVdw5smB5iucgnJ9iIsR6
zg6s57c+nKsW2sljwCWXP21/zT2veovxiHHtwYuwZCnBCjEnpuhEa7KwWtKvyAcARvqucJGjxUSM
I1AK660TGpZoUI0LIiMS23GzwVfamkn1vgAmbElHuJRS+O9GoYAMuH5U1khbaUTaIL8Ch5rg0MpA
b+mbOx4SV6F3/NAiyX6jhcq0i6vtqRG/UADzsGVbzTkpI/SbOOvWf33b+cnWARfafC8zaHzaX/IE
lYSjm0Ob2eqmueoFWNRvqm4Zy0/TG10Ovn7Wsn6tJqBAZR5eL+qAP+w3vwEecsfRAgJKABBzp8d2
nEMI/q721wYNSBC54n63UcNNaOjPVHJ+heLRI+gphNu8wjaKWPODHBpWzMP9leUa6tO60vNDEkXV
oHsWLl0g8/PDlvVKH0GLqNpOSYkYd7JqKGNu5oIEgvgmvYGFcqwCNEyoYq4PesWXDL7u4cKMFJ3Z
KbZFOs1fL2kYNXQhNTNBHXVaxrRVhoMrj0gT2wGcdvHXi403LaGRlhxWPPJb0YuJOiVYHK1Q0cqb
EGb0NV1z/twmzkdq7ORWvo08st6iy+ID8HFn7vSy4f47N4ECSbVsnp1NS1px8PhFvt+eOjVCSQCh
u9tKsXV4UafcA0vNXTzlIOwUcluuiQwkv+g5NWvgedAbNI5JaZqkWdMzUt96DcLjlSYNB5RQwZAS
MfUwwzDnX8ViBGBvWEqqgORZroJ4+UjLC9w77nBqTHkCDAQ8SG6wnsxXbnp6fVJyrH7wc98ot8kM
GvvoL/eei428feZgRtbIpRk0ibo0JauG0NTeKnpgIJgpb1Vhcq/aFXZIxiRqbRRrBOpNaJtvZDIq
olQbL+ahrhpsXQjoNx/r+wcKZMN4PCGLk4+z/pScO4i2UQwqTsXIq8YDO7MtYYY9a8xJnaS6h9Kx
y3mNWnzQksvBynel8GmHG3BjTDufxriQjKnXhM7x/3osV75+NxAQMvToKeuIgrJHofZFcim5hFDe
VCbZABqDWHY6OhrL8eDsR3r15E44AFPLq/YemitVbA0BhDZtiVs0OL+1ikRai2ZU5FyttO5iWNc2
uQS6SuAxp2WIj9cXantQVnzTTwBTcM+ab5VaPVg3j+kMBP0B6qv+YugtYzMNKrjaVOGW8W/tLFw6
bA1jrJ8CcXKAPrw/CBM7Vx25Go040Q3immba1pEEmwQe3kepNM+CwugFe2g+CfB8c41yvfkXoS0Y
aXUTXbjjjl0TjxIIy1vkGhOp/J+zAO+P3n0Zz6I2GyiCaVusGkEATrMT83Ja3moJWDyBns3+G79v
WTPIXA+yohLCe/vqPGfkPR6NSr0Q2mRSwXTXfgBjHdNSaT5hms2Ndk5w+fQ+COua1m9peniSoJIm
uZJs72sNvhl1obDeyfgf5KyC3eFzKGAtc0oQIp96nTXHk2wJhaxzY/Y7GKY3ypGO8Dnozwh30gC4
wHyxcoCXA9a+UYKdhQGO/QGoEqCYRig7i38DSFOAo+8XiKV3XHFLP/BgaoFAfgu3rvrL5M4ilM3L
Cccy1LNbKqWGJJx0HUATyjIM/b6xFt28DMF014H7NPtduaky2eaLHaXsf6/KJcbrJoA5UvTR25ts
l0QmRb4D1+wor73E6MSYjmgp+zGRuwGbOfaiGs2lfrrp7wr/AtqphWCWywRCW7eV2VqnvROQokH8
blS7LzqfMs3/tW+vATRSVGcwyC5l1DifNPZiarZsoOEK4zmU4mA2x+YeEAofEDbWnGaByYlm++U6
Ac/oZQD64WTa63fnsNtY8wWN3ZMLP9DF57Y8C+wo5p9VXf+rJzOrjxfzFI6yd33uM1LIQuKvQdw6
/kmC0u0dMHtN3XAV2+QrUNA3L+ajnS5YUF/sJH7AyfiNlJ8EAbYPALafgMtbfMzhzAnTG7FE5cel
nZM/ChRwXsfIAOWvS5iNVdWXgoiM7KAo3uETq8mU5MCwS8MtSMoDS9kj0q/eIbiBN3GPFUbIBHkl
zGC9PtxCHiodVJp2EwOy9XjaFOHMcpncbST8dbDJpuWjzecjbF+FDz/jdoyP1PtTHVtXOEe9T496
/tRLhNUdTn3t8FgOMSWWzVVVJ5WKyi2R+1FUfsHP3mzrscy/MIExGs3hIzrEYdM0T7Ka0KNLemww
BRJ2GV/u+ZtYuWjEIzoQ6VluE/rFftJd+IuTbHf9MRHVTO00kY4VJEwUTGzjLZiSMFYBVFoIuG3D
evuLdq4Y+2QzhIPiXk5JKbaSkRRyLM77J97QTwLs3SoauPRCjIMpw562I2xZFpLmvFfgTyaAFMSP
cnq9S7T7efGH9/HKjT80j/Zl3pwTw2Hcw/sAc1fr7h5wHof/nL54BYIG4FaIr4sMvhO1aSSIDCR/
uJFnNXR0H0+YgUQhWvosi+XAD5lgCwG79izZ2cTlgZhMw09tuwsXpiZ7xq9tGAWRaSB65mLK+JMI
GnKmq52laWnbDuCezRheeMAQO/Bd1gwbVTs88WG+e+HbsCZreM08OePY3g+IQUvvvn9nYa/fsacg
2G1DZ9//H18pv773xbFLgLIGDAT2O82PmDzkdxl6czs0zxxsJS7kBx9ub8NT9HG1VvanHLL12O/U
GS1x85bZ5HlJrA16MjuAIQO5d2AaMtnRkwiDsyoBAFBwhnzzb2BGGrBZ1G34VdS39Xo21HUuAXk3
/+sstLK1Pbpn50Ko/XKc2J7Ic/hrCHxbQA9Whyi7XH3MFA0N0oYakWnfFCY8+51xGNXnWI4I7FWn
BKhaNMBrcA2Jixp8OBx14ZW5gu2KrH4ftcC0PU3oDHem3EA2ffRLvzo+HIREsc8WlS/6++UBOrbI
QGsgapC2hRVNuGklW9sZk41R+KbcgiCqNZpGIQ10exyrbFsGypY/k8jEvsAnTWLiBHXpNyrIvy/l
Iymkk1WZcCx+et+DV9hLxCDP2xUdUqz0Q0+26MJoiREjk/IDMShUyqGnUzNaH8wG3dB93UXqcvDS
MRP6xbPDYJ+aHniFL+biee9WaA+ROSnO4sHVH1ww2o2hjyINpoLu7UUlMg9MG5Qjuy+lKj7qS4b8
6Cm5KeRWL0fp2PtTPKJ5u6H2WcxihM8aoEHI7D+xuh2m5Ne6LbnglBHFMaOX2VOi1JcAmQU6QUmT
erexMma++5sI5L4qceVZj5zaq7svpZ8UyizdZoEG3o6DLCZZVk935myzCye9JGkNivNjQZRkIPTs
HyAT7E41bQYZFpIr5VIqzrzZBEJGVR0H8xBbjyfihk67iLZ9Rbzq+XJQ+YyvBQKpkQcQEnxiyOaW
LXSyOnu+Er2a+hh1+ITtv05ZMDH4q3uyBy1d7lHn9LT+bQGYw84YaH7fqL8EonzHcQr/VIuTHf48
Da6PhFD2oU2tYhgJ/mjnuOObh7p6DpxLbEsjHOdRMNl5UtMCMW6lxjijKvCtSs5bGk4Xwq4BF3uu
wjgRrovSbavRvQVv0fA9NSDXgrCpffSKb36rnu9BszKjm8JEn3eJJYygB8eSv3c3XVL4f+m5PnhK
eW0COQJaMQlx5IjMwjfWNihvr0PbwtOnSIvTAbX2apY/KrfUF+aW5S4vZYv3zSin7f4/KQ7pv11A
PNLNVU/QRGiZD3CP8QJuVfJiFyLw2WFufmXjMcgepevOSb86P7E1yOYiC4U9efNVQOVUmcmrWcf3
Z8gPUP714Fp76VW0N2UCHv8mHS0C4Jzgu7B4K2OjrmeeOLViLzrbNDoTc0c97yzjFB1Er021/00a
5ihUiGC6O4cjC7ciOvYEO74x/jbOPbthPYNDFws72SbawBeP4sVAqorIJ1prQr6D/qQEabFFjDm6
7qRbsYUJAgTjnlNjItWd02pA+kjPCVOVdhxvKMTJMDhOj4rjrTjuD9892C07ga/k6TDIczzFoh0V
v8BCInONwlVY1g/JfY/ImFpTF3AzoSNflZXZGbQ6o+d7ev3D2sslkS38LDpz09+UhvAMGIeFG7Ju
Fswef0DiCwWY8W5FeJLtMSzPmq0lapnEFJlPU4RqfzypXJJH/wu4fzhDYAb6ObTM/Yvw15jUGgDv
X33nJVIAt9M1K8oSWLar8iUMX/3VBwsPcc+LFv+Plzm99Kc6vlyjDjE+CwAIBAk0y8hAnBzE1uvM
mor+vqqTrayNzFG6eIVLts+R9PjM/khlzkm96rGpCDcMGijy+WDLFBWQJGAw5idCjXafZQGC0plt
lFhiFkCm2jaNJSN08GUdSmIZvx/13l3oGrL86zSSEN3BSPhN9MKu9eA//pjR0NiJv/1FNOXcrRJf
hYqg7pQEV5WIPgo2JXwUiiOikec0JbFG6R9jb3SOrUr+1COEYRuXnIt58nFDjOVuJGQMzm0S6waT
2TsAqQ7wa+B9JTKSbUGOX0ow0fbhKgudubWCxtA+eKLvbrVE1iwl7sndGZ1u64YGpw+yYgzMHH+p
lfeeTT7yoIqas3vl3jWqI0xKyQD9riw4L0ZBWRMQO3sidGtBGdp+HrI2emUmB0BAJ4aB/hzpD6LJ
pJdDWYTqRoHKhsESBVeBQDfLghEdPWx3KyoNM1V1Wff9B3mG6XCZJikFeZaY6L+LpFoii9EmnLvl
YhK+hOYE59dHyNBgEvtOxHeyDATPUlFTbfcFh/q+9qtYPEmH6TG9/EGgz9AvsvNgG1PKJurOMlOF
uMFxlQqvRYD48N4G19dPaNgDPLPXhgxZBve7MjxfMhOMkndpdwHFD23BDzUV7LlTc0Ct6cgPkaFY
NKgWpVBVPqo9QI2mvmlPxiOfe1/kCyup/FVz0WZtKKXv8ObhRMfsd80yUXxPF2AHhzj7OiGpfQUj
bSaOgCP/n9ToAiSoMlaY1XanWmN8DyYDWQKptzRnl4uCsVMVGRjbiioSWtI0f8o0M8pTXAtHC9KR
YLOeHziQKiFNhlOvqqliMkjOHPQywxbjqCpwV7YYZhZ/GUjWzpPifl1H68K2p9zPL+HZGqt63qCf
QY9kXqjq35Pe7CZNx6lT27GrudZri33O/JZPKQvOcwPndRPCzTPNh4JyD5B9c9Bh7pn1w5XbzgZS
guoInFFQgMKCwjOVnLjakD5xObv1xgHujDItgjEbTCo+6R562hqdGlQgtZ2lwZUpjkcjgP9BENaD
u6W5RW9c1JfvqdnkmZVtnWhpFnDsqOBt2iJJF/7zrsUKRYOVQrp2jKluvAnE3KT+/yjytN1cLYJ7
uVyAaHuuPtkTfgz0MyWgiJdZI0Qe7/LPTG3CFJV7qCgC6sbr4eQPU231GBp4LCvxomYmII4HlwWu
RCA9np7n58Adq0b06PCgXb+KjmfeYhR3/rW8BWLT6yvH5HvbYHPW53mYtsmAzrC45GTv0v8bsPQq
X+HCxjPStvkg+VFj4XXpLiV7ldaHlj8NPRmbDG1z4AzcYDZVSR1N7LUJicpQF49wO0s1moL+ni1N
dYJ9AfweM3KpVSCo0W/q8fjNdqApMXzSR9QHW1wMOr84ZFeAWKWxWwK0aSEKr5fdh4/p6orLSaYP
fl75M28x3PldBG2HRUs7z02cOgr0PZ7+XzDX8IbKhbrsvoM1gUXckHQj2X7TioaHQNP1gpJ4j9Zd
rEUDXbXzn60jb+CUPFv1zEc3FDdTSgMXBLNob1O6WAbGMrU79y4U3RJ3MxA1hwmUMVaEvVaeHmzR
5X2iHZLlOHiDtkDTnizMpRM82te+mtw+jwHIek9QJYWVs7SvM0fd6bdJnQM8latkTQfsinnl1rRS
qHiKINL97wSB4Q1PctarTyIhm7Kuf8uWVMEEmuRnabjDJJZ3dPlENOkqMzG4ic0lrV42L0MfMJRx
rGWMkJUNSzQHlaIQKvr/+c/sz//rX5TPF4ikark3Smzys0uxV9tK4bD+C5YAHWMcEenFosDPOvHK
cuccvl0wLp8C/RTNI0t5m5QF6YeWm5SUbKWwn+aGwzMHlkc0rsF9fwePRDxAEKnAYLr/3zmematM
fwkYOX52FUYES+7tJqAwkguj7/lJES5NYQK0Dgr1chW5ZPm2TitNqfMkpOCYVfVC/uh5Ra7cKWFr
QxFrQWjAV676d0S58Mb+cZxH5LM1LmlqcUFDX3sh89PQMoNQTZjK4Z2h3JHbqVwGGiwXZ/xABM4f
tug3zuvXV9xhVYhnZKZgNfYIT5KqNIe56lYZCnIhwDgufYQFcUJsd8NCv9YFwgpIHvhfBDq+maXw
Rnb0dlrW34IxthVyuZStTnZ3C/mqrQ5Kwfi6xCUe6Z0odErIw8D+cBjT4w9NEeAFQwKpyaEOdAIN
IBCVNPbmMNR5Mf6RpdG0rLYR8BL/x8HjCenObiQQ9l4ZPtlbqrYLvT0K9QK9aFZnCfOBjAzDseAS
gf1kg9GuwQrUN908ceR7fslCyCs67reJlxdEvlPsygj9DJ7DlSNnoaK+26OVE5n66XqY9uZFXmOK
F/OS58nqg6k/gIee/MOiQoQvOFjA9wc1M21SB2RWJwh9mH+NKRDXCSROa/rxJSAbsYj1Q4TkV2bh
gD5H3MCnSp4lcDr1di7urPAbM2IP/UQBCblpi6f/KNRNNS68GNHjyo0MIr3kshCq7ZBkwQRvfop9
CP/lAabcKrCrDyvb0PLTN79SYTppEOngyLZTKM8asBMpK9doWIeAwPWBlkm8+PRujsr8FEZG3d5v
cVvGS7cpmhHvskZtZ4H3DhUZ2+2FZ2Yoq7QdTn2hljwc2XtOhTwa4lBmUl8QTo3AUCof1AmsvoZh
EioZDv57IrBzlBAyyt7uIsrwM+PgSp0+HpuwzswbO/rmhA3RQfN3mrrgL7iIUHbzpN0w5z0kggM/
VjWirxgWcN0QQb6QvSnbgr8rxedRo5+URIOQic4mf4JTn57aAF30hloFjO19blU0KjHXaS0xubT/
GZdVyu2a0qJ7zmLnSzfvd049Eu217PoBDotinbZWgyRq84/2KPZayD1O01AEP33B1UUaBGS2Ioq5
0NNFHFD+7lSKNDZ6xHBu5JMPtA9OamYa9hgcUMGXTmHt+h0nLqea+BnABvBTjkFQ+x+EOJLjFdVu
4CGYWEe/AmTOEoLhs8/98Sk3jKKeHWQPs3QNcIC0+qUO4/++dm3uCtZl73BAUVRW7rSO8wytX06b
6yHWXaFi5GwJvm7MRtAWymUFsZ8IK6QRyAlFmVTjXLe08IaVW91MsXEaMm4Kif5P8KSmFGRSUpJ9
/B80hg8UJG2JgMl6wJqOZHHtL+zho9qxfPd0nuh85CWbHBykJP0oOSwzkslXaPE9huAMxZwN/6Mz
jP3XhJOIiW2pzR8Cgnlsuu0w+LqYdnHXO7LnfOf0XAHDrIBOaSLTqhY9Z8tuoGy00/qo65TIK4Nb
ccxQ1lFkdADFoEPez9RMxDCEULsnLOG0D/fg7MYQ+j3+YkIhOHBXWyEbHnZTj5uBVbkMDYCNsquP
iRqX6M3TftFhYzZo0lTPoUyCQT+gu6gIJP5ThyniwA/0ZQxUVWBA2+N7bIB8aReywePN95Ioxep6
vkQEB8J9drlqTGFVE4ZPlCiAcitCI+w/T3wD61LIe1aLCtqEnt8HErVWEMMP+bQAtV7pjbhVp/xv
0u2C9IhfEVPmTKnIQBPZDea953NAxCgPsbtLb/CUTnIhavHYKjH/gYx8I6ueTAs79kHlPp5qrrq8
mJTIyN2EI1UxCTdaGIl34G7gRfHrmA+dld9GDZPB4mkO8IF8lXnhpJmAZIAlrpmU6DQNN/Io8gB8
3tzQf6ZZWffp45YFIU4kkSZOutdtPOUOjiUTTsNvvISon5h8CrJa89tG+Oc/FTyM0qkqQ6bRw4Hy
6lB2n8GMZvrOVVwtD0upfclZjRTouLQeCzI96thqUXQriaqKdMfg8nFnQWoioxGms9w03hhxXzCv
GdQ7r09vNMlb/URow/mOqpmBC7pFfcX8AIfPIKmxK0Rc7hT5TPbrxUwE2Bng5HFDVSPgrhMI2Pb5
Sw+xsBDXxZxdLc9DhN07RtLFP/ffdyyZu7m8nLI26VGN7oO080+Prx06UNdaBh4ccrnSNzlnMIeR
IIiuhWVuNtiZXOJPha9ncVyR6FuvpiZ96njuk7c9TeD/0bmdiMoaKE8BLovjp8mN6Wl+ezsAk3Op
2mAFYDxBagxN8ZEtH/hl+sDhhQuVXG5LC7kYr6lezlcOOWvuDwYSklXRC4RqOBdyZroxJZfL4wl8
hkHF8913bNjpRJx2LVoE/81Gh5NGeOCly2PxU0dqGVpwWCORf/nRyFGYaMwVTvI01DYDKSceWcY5
ZTTB/PEKPtbpfA+/V1SMqDHqJkH7kN+Si1R0672djewtFaY+pg5i88fg4yqttGbbPxosUYn6p35P
sWrYik0b5WWkQLby7zoD6cNF3CCMJwbSWtP3hDsm7Oh+IElBAfRbuRc4mMlTF0e08tffxspx7tfs
eWXCYbpGDfH/Mk2uS0liI8hhF0qgu8DN4FrZSFocvuriyqd91tSuIkUwJ6nyQS7T3rq6xZI20JFy
Bc91RHnjZMj7luPGoKqHdNUua0N5tw5gLca38vrWtShlIX56xyVftPHpFS6OgQW7OUokky6GKVkf
7OWxHa3wqMuMAHZk0rKrNgSHWZIAcKLvvcLTX2bdOKLEj/lSQ8/HKOQZV64GRZB8gT92x44O1tRU
krtDwZnKzRfrfeLn3BX2f1UTnpnNN8pycOUqEvrQRVqq1XFY0aQpyFMrthOyo3jfeWhnwPW6S4EW
TOv5NDftnzi2rZ51BJRqNZv+ZJabgZj5ci97VkdqpqB6RekVteyEStIEOlLuAkDP5ExUckIozCC2
RPmaWhWCqDRI17AGP61ByBXRRLjgDhH1aPSHd2ruTszZp64tCaBS87XgfONkH8X00lqUVilRvhzB
jYty9WnMfZlUHf/RgUvJxyhDT5ptQIPtFXu1coL/G76A5ia6dZqEAppiwoLMdWAvXEhE9vI0Nm/F
6vusWqG9RzWQw+2L8WEk9K6k/r4TZRbHUdomt0TZEVEo+2BOC7jAJH5ScXK04NIBN86hq5pnBp7Z
dwcwdxEmEZPFRL1QFmpItbjvB6CX1K+1IXfN6wV4rycjE00wzjonIyFVPuneRGrrzzgv+URxa4gR
n/WYG8g1symcGIpvL8gq6Ha7E6tOwVFoKV75GD0zuqAki8Q17V2Kbj+uzQRKC2r/BQ1NFUOsUkSN
bUUbVx4tnBUBU21PWajEVbeiGOTCsXgPK0TcN/Yf4ocnxIwramNgUKk6q0d2OwR0si+CKdzzGB6x
BntZBBbE4tcwbzz0g0O52IMbmQI0X07IxMEOq6kANyFSspWSyEDh1M8bYUPAo03g4li8lJpgwusy
94kdsS/YTUmN7qjgkgahFWONB+VWH6U5aeWyacLtI9RR3CyiAeTo94BLgjxxRHw2p2BWjqhxqhYT
C13UULjp+RHM6bzPPOxjhbwjeZPPEdIO1c6DG60ElR/L1Mbelpx6ccQWNyDX4U9YWkzvtZdJagp5
2KiQl1Iu/tiag7WNFzrqUxif5HrvwZYQXnFq86be+U8YfYPPmvMS1WHYwhpLpl6XswTSLIeR+D09
ixXSFNzzv2AZiZMfU7eoJZ3ejaw5T0jk9mkJZNGgA+w2pRmMc/VlkrcbKAD4VAbZg+iz0bKZndGA
uwbZw12pX0tWcQyOqVBnKuupPLGE9pz/PNJOqPy0umRT0FlIWMmWunqwaO+aIIELqFZQF70nPeof
l99ZMUJKAk/+IFmU+xbBctq7p7tsnPdEq/+dkl6Nk9U1euObx9bRlv7nTf8WnHzxpy1XDza1ursH
p4k/L2Bz91M+tIJ4MyEOImyYwfacsRbJgKaRD2zQAFn0yl0oOWS5+Cfqfnvk97TwsCsipzSu2qAI
zVXV91oCzgzN2K536AGAfMzq4w+6OmCjUevH1IQMtoCNgyKZefL1SA88GYHjnVl7G5moLQPwYzFL
ooS3xXUrJ2AQ4wQX41yEejA7Lm6xlRJsHPMvDbosCbNxaG2zOLvpgadAIvALov7nkdyLdY0PFSCU
T4X/+2DsHHTaDFmN/7Mcwk1ar0YBR0lq9XU7U5sTfS8f4EPrnp8GoDvS2Nu+BIRw1BU7UzW/gvVh
we9RuXG+hyhoPaZ4VaEZxOrFaO/o3KtU6th22DasbZ7KWkX3gng2d6hOqEA9EJYAr0bLWzHI0JTD
gDRwjtXtuYU2W0dYdVupqbB/frdBJFRbqqwYcBmGn6L0gFzXEsP1bv38v8wXx/muyPmpi5PSI7Ld
SuogvhCjFvzXj4667ndREoBrX8wYsiJG6sByy4Y07rXP2A4SuXabMk6EN90TcK3bx/wGJFvL7GNn
BZ3zLUiVlTeTcsOObrURDfPXoNILBNwEmFg+qUSnQKqzIZ3EbFbu0BIv62G5pEl0iphStEI5XWA5
4PVyNjvrwizcHZU7HPCfYJV9VRNL3z8iO8xrduL1YQkgr4yfRwNaCKUx6GP6+lRafKxqKcbIuvLG
Z8uiw9LnRisAyzTi0mM2CRXMOughV/7F9pK7w00k1Vs7J4gQriytFAqI+OggxQrk2rDvvCF7t1I6
WlkBLKQBMzaOfoS70Vc1FI08SM2tcpZIdMCaGZ07UaaIwJW4h8xpnbfMvDHyAVwVSlTJkq/F4OqY
y2YmyTNl96J/Cmo6KOIXQSPnVPV4Zbiu/Y6GAiyr5BDlx3LxLim1abs7OU6yAcKbogkSMr4Ok8cX
Nfl0W2EiIJ01oibU26SUV1fAgEDvwFC2VJq+hnQKltJG9SvKfM/Vv7FbEU/OeYA7WOnrxgqSfj61
xY3g7fvQ3fldkQABeNYuvYC8FeS9D2979ggyuDALlWK67Zingxo5IQnpgJfA/T8ir+gB4RNY0/vs
fJTDg2LcS4mGtVtiJEmcmR0SGaFggazn5VHMCHoLFsH8JW65ShyztDLCarvBFPhh456JiijEXdRa
2Jc6zXC5Iz+MoHcuZXenqE6ECUdyeyKaFnAxSlP1GWbOmPKDoU2EGAuVZzKF8Itf6MdBWbPv8Uq9
mzeQBEttw4xnlXvHVqMF2c2Dljo+OE51aySqn6RCiOo9e2ce75tT3HsXwamT+sh6XjfW7KlE8ZzS
2wfmcKIuM+nde6dcFrMqFsEg9ZGltccft/IsiI3YfrK1e7TIZaCsUMJOYhsSU71umKRKrIjB91A8
xTh3ZVKHTERK0QU0uUUJucsb9n4tAP6KSIwvaXxWMEFLyPAU7YbLkUyrtQvux6PtXdp+HpdftomO
EQFJIiqg2lr6h5TNGD47JAPW62VPf506+i/k+XkUIFRZkOx7uZ2+CqZXDkFZGLulysLVDQEPGs3n
C9PvCwoghk+YX6CTdYZgADRVTI7OFF9GmNa4/wNBnxzy4C1RnXBQ/JetnuAUXu4D8afwbsEVDE1F
nBx/59fCstDC4q6+fgqio3U2hH3Ja+vnxAnR5t3GwcDOOiNoxXMfzFKe1i7By7ROZRZncG8Y0rUq
OhyYvWHhFQm3p7Clena1RTqxrj7m0pfVaI7DkwMj5yoVtpvYYrEy+VSMIZze9YjgYVfMqOAqM3s1
KAr2LyhLh0lCKRvQEESNmOAHKUdEZve8WjPRMf9hh7p2pWzPte/HJnQxWP4n7iFNK855fvNFLvyV
rU0C4Ow7XJ0IYUG5uZbCPeVZy/Sc65LHKesivKchQRJ8LmY3NbduYTiq8hvcurS6zCyE0mT6hz7o
Ozwk090pZ+sFqTIbAs/ymQIbE+KN7r/APK3e2sSB4opIaMBKeWt8k2ZhQqcfVA1oF9tQ8cWTAAOD
mk/JZn0CvjyREGHxSNvtMQHQKkWpiWxpQB+9aF3LZmeQPAYNRKHeFl/gUIuNst0mJGCckHOSF0gO
RW8FALThZN3umlEB3jEzB9YdqW1982V2KFw5Sv0+Q4zfCbOrIPQvO6NgEZ/N5ZiJGNchIEk9L2SO
nLd9HJQ41laena+xyQakEKpSU47KIfXwOQ7r95fuaC/9dzofBl+8CFW9OCezrZ6ODhyytyuFe84W
tS2+wN4r8l7ZNjqZjRU77e1xT5ULK+0Pcq/zBYNWHZHv74P1nhGuCEPhNQdb77boDgYkP/NszNoC
8r4d2yu503PDkiE5cRh1fx31FAg/kxv2FIWDr3Gz1jnksw+ZoszV0P2xHoE4QOpyQ6Z17Pj2idAK
LRSwcZJtMCDROjHrJp2JITSPxHaebSfX/k6SsUcHIpbEqMs29UEkhRCvYhH0pOOC5/gulTxHOMLo
O0+T7Mg3HbSZ+EMlkwxRuBtOE261Mn4upJaEt/ALIIGBokLNcJgY30Fo1uwLHNay5u8ApZCO32WY
XaxgBfLbCkmgSiwgEqwEb8mHWXyY4PVYCyIL3T3ZaFoCzs3RBpbhWDsUn8Q2uCZGM03aIT48QCt0
E9eNpPRQHlkXoLRBy+OirHhBZOGBjByIAM7MPJQhY+Q16i6EXONYOQyDlG3ESnAjgjh3r+JwmU0o
ln0xhahoMLAqC/xZYb35ZVIVGNf4lMRBqZDfTxPpv+ItObppIfaMym6Kwj7b19m7OPi6qn1CfmZZ
r4ahtPc0kmfNc9qQnIOWkKUX1N4Hqx7lKObohyCOW2cMd3dE0T5qenoa67srAI8F0e76EmvIhOE+
O9nFIKaguXS8DyVJAvYNrbLgqbJYuVnvrlf2tvx4CRaVANMqWJIkaY1HXfpWSml7pJA5l+zCu75I
BVHCYyIPbOofpP4TJohEakt+PAy6m5nM+SLE5yKVn7OU7+knrbxuu4gPBHOa9EFTVLzUenhLtZff
vqHOb9/hsEzvJO0gqgg3HzkpU47FVlQPo2Oluix2cU4KGn8TK0nUIvqnq5NnFJUKjBmAziZ5ARge
0sYH8V1mg6/2azjWUXLRTdXA+3KH4kWqgNef4C0KeuhT2qE4JKE2A+aCkGhDoxEhWkPp7vuyNaxZ
I5SJDut6+tfhvdRMGZcEeUN10PhnzEzLOhJQQedpclnGHUgWwtygqdl9sOhGrtpZgI/aPTiP2drD
kTNQNDcdP6IbFRBI8Lzpbc2MbQUGnBVTRGyLF6Yw0y1voQQxQZnazPo3BHU1PZyUVBl1sV0hxpHQ
huEZ0yqP8CxXVckwz8rcywZnryqD+wPqq1Eb7eOl9qIq57xDy7UcPiDc/+23DCPgGsh0EAtzSsP7
diXTIV3hYmhANN9yiQYD9zvjGCh3WRXGGoZpiyHq/LQbkWEpL47UFER9oVtUL2LJeAQp2W0F52Ys
nUknMJw+bFOzMMFoY3Z8k3HHUpVHnvfUoz0uO7k/QjieGbDENGabarwGRN5iO5M6+efMVf2SWBx4
hFfml/A/NjRH+LI6chnR0h/sQG00EVrjvcYpd4eAMWUZIn+2yQ9cEaOqtY7KTvUnKgHyhZKdrC2t
FlUEqj0QKQIoIGXF+JJuCP2Ed+nXZX8dgxeMpqNqG6RZRr3tQeoeC7PaLZhL72uESTxJp0dYzb66
dtuLHqZpVE7ZQaVbz/Ns0SfXkjHZ6lciSQBRA0Z4RHrK/OEnFptutuUae83ssXEeM8ptbTwc3qRy
MXH5XJOCZ2hYz11maWlkWFGwoRuTYu/JJID2QSOYODBz74tNqEv8Lqnrqps6HIMVFiiKPuh2nCkV
yAi+e3M4cX5JHCMlvHh7rfAYvmsTypLwaiU3/dsHzXo93REsDMnYGN2ndPDENUk40DZQXGdOOZh5
T7WXkTuGQwjkf+FMjPDQXzUKtBUof9/mi6O8H8HtUQOKaJfuC3bRm74kH2I5Uc3mhjcNeoSySX5s
MvI6mkTzuuZuTaWU2wJJmR/uBGm65AlEPQlVbEgDw0dHFjQTm/z/tI7RCRgcDbwnMD4/fns6NRf5
JhmDqlotR84oegnk7Jsp+q6bkLePBKFx10H/uiwut9BlsXIAGTrttzNZ5J4MOJmIEFL4WxNwdMpj
d/FZiek64tKeXuEVv9DmeUJRqD/M0O7uss07zeCS+gYP2kckpmfRtnRd3OOXZlZ1kRT8V4ARNHyF
NXVBizG/H54ki+JwOseVtHsRQF/dKHdqUn4bjyLmaxvblVp2gw8EmyyczeghvamfZiwaxHjMjmvx
THCX8SF6qzerW39yrqHA1LZh32Q2VtsHs9yDfK31i0FLoQ/2agmwVEo5O1dzpGYzQ4wQcOdYLP7r
iD/gjqp89O302FBj3chnu6J7gNerByFTVPQQAGMMwWjQx5xIkEto+GkqsZicZOU3U5tThkLM/J7F
2m7KszJZLGarbThKCj3vZItIcZs7fycP+7EzqhFg2lrWEzDwBepOm0+cOr86J1H4Z1SlDgcrE3aw
d7b8O7Gin52Q18G7UEPXfxjZC1adm9HNsbwcUUE727RXF0OFLwhVwMnW8saK856YL6umGXEdtvEC
eXFOwaPge8LF5xtAZV25zjvVMXoCKtXd25quHTpibie8G2B/3Dh2zXv+63iehluQ3okhjcSAF3AM
cSWPHXHTT1HcFHk+woVdZcFLIP1Nb5zC+Rk0y0qCn6Y7U4ty2Mwr7kWlv7tup+2G7uaMT8gOGq4m
4rMWXi/A0B9V3SqH4mwPoZB9xhAhrfdYc8znATNbASXvJ1WmQp09A38O/4d6pTjoDp289Qk8B9ca
wF/IRhHgwQowFV8wPI9JDpC7UhGDEeHHqzb5ZetijEPFq50tMEOHDl7oKqvfRkLVHFyhL2BFcwao
CGFxG7RCe8y8+2MUdMfRI9SzKaHcAb2UKkE/rznDfcOoSKsPS+nSXOWhOvZlX2gZ6gTUbYmDrW8p
Kc+LtnAXKaw3OwamEKDh4DEMEaeqAecdNCZx+8ygoMQ2e4BkVlnrh8NQAZd6w83kI0oBLeixejou
2xFMTiqUXAN/zoz9Sn3hQHLR0vl2ea2q+vHkMajpn+woaR+CkcyB/gsJah0SKR/vxDwcmuNfUhB8
QuXVfGHkA9QX6TlBrhJIx71vJNFOQu53p7seUzZIQMZrIHAhgNBss2ZW/3RxAQE1yqy1d4rQ/tq0
WhUDxBdBlLUiEVhKEKZQlU3/TwR3bvTpmKk5QTTojiQ7NW9ICKYlJHqbBOB2w0TcKHta1GRTUrFp
eNWpnH6qvQbzUXPkePlq0iqaTy4tQB2f6I4d75ejfLfign6Brp9C+BraA5Cmbf8yRGGZ8rXiH2tT
IesNPjtGVmgPFjoJZuomDr2XdFoHRyFOJs0v3Kc61Jy6ZNjx8x8C7vz1BnznwAf/GCqqCxJp5m1Y
gMqicRr0D4X2bL7xFdG2cFV6e0jIEEbQBfsnL/XmZDaPKo+s12wqx0UbPjTL9W/9nABOYegz1zmO
BLXpgHqHos3Ax5C6bmrTdU9LNLXcZ4xNsXT4cYtvB+iFjBezhmJmGZ84qYD+JqDUw5NrtDCW9qJn
UZVAnTetqbD3IcvCd8V/yYim3iZ78bXFk8zm0ljojGRVaHM+x5MT9rOF5fcQxK2EhTPnDf+pTsS2
fk1ielciGymDNrTMtiHNH2SnFUEeDJMa4Iw6sA8oyx+b2TZ+39RwLroyeAHyoSibyQQ/XBbyZqy2
LX4sfr/bM+M/r/sby7SXI9ZdtFFBIcegyxkWHghg2huJ3lBJXvURb6n09VWq8wwcKMzKJqcH1cit
Nbywusq0ksMYQ8jPySAMm6ZhJqPgIyeFNO2qCl7/yKpjQZgmTENMQLUMu/P/CPLCFt0SbK6nSitr
igKPmOHT7ILcWyXLWvxEeOIplfefigVvSMU+R6P/YXNn1HNYSg0agQM92xQu02n8lDZHmY/ZJw3q
3lVl7TJqEygbmJwsitcx3UqqdHjOEuL4lObabES5P7+7IWtReSCLOS85pD7I8U/Y7p6uLW5PYE2G
x7K0G2eS0Ejx1sLTF54ZOoxsDhXgQA+4s18900BgnM/SbfzIH6M/tv7vd0E9ZSH/s3WzrIIrFgwb
AkFMHLvz1o8Xrb92uXxhyMlbhg0dzVJxwbqBb9M4bI7wA07ebCj2W0jUCP6QQ4gL+oaqQUqvwxjK
FZhhot/SDj5kZcw7/a9KljXHR/NhW/OvDG22JFd+TAUO9K+2GDwb8fNv1jkRDiONp6Qmo9jfxcEU
S4bTauX3dcVryDHnMmN6vPNQH0M+M8ijBs+p0/06Wck6RmcQJQ+Q0phuPwn8MwHNXAznqGfWKeuJ
OyedW3qrbjBwJKggL93c1d0ujmNtdG1MV5YV9ndKTg/7FUgiD9zc4neT35dQso1KY5usgR3S0BHl
Sdj47C1SQErcsxyO0s+vZn9NfLbz9sqQpsqHPVvraHmilv5NramyVj5lXePsdo5y0kf1PLH4A+ed
IL0rmAs3VReWeEg9SCsZca5h8i6OS5Dv7qJ9aJtNzGoxjjXct07KwhuMXtZrZhVzguDXqvB4XiwE
hefm2/+Na1eg4CpjDZJxWXTWcpA1vKjYnEWcbMSkRujsOiHDhEVMYS8ZPXC7rubWsBV6ZXpAzamh
KRkw35NGyTjJjQD8WnvHC9L5fjYulAEe83BIRY+Ka+72P3og3CdIXGL9SdlGTt9nmb3ddvn7RGnU
3XflaX1QP9gu9XKYWDMDBmy78tGnv010tbbs8/TeoHgC+ftFUmD/SgLqlFMkKsp8X50N3dBst7J4
qsLNfNsCQgNMnNIvDkGnMlYCCqHe+VIXrV1Sr+CqzY3nH6jXwGASfJxGEVBT7c3I+Lv+13xdZGEx
SM3le29T7CTHVtm/DIeEQsXgbfcvISGW0gS6egE3UZ7Lcazwi17rcLfCZx+iR747R4jS9rjNymsc
RkYn8Zq5D5vKvAlQvDOCZAjTPm+i17qUcxhhyxbp4i2QQTQS+VizTNhvKcbQbyHybTRel+ABSYcE
fqSZMzIDmm701K1wuBawx/6+OM+PSXsED4NtEKebrpEjW0ObapR7Bvv7bBkAcAdBbH1wt+ewKIFs
8TC6TbUxnrJqIRzS/wAyZ1huZoj/cbioy/GFplh5zC1INpzjULQCTAaZo5bzakgcFBzgb2d/6ZNT
YaIPJRa5Wa98N4unq3phKBxniyCwjZLrusxJkzc7yrrQ8189MGleUrKnP70nxhU6t/+czyMC7hcX
wRMWrLjgHfC1A+ZvWYQRY9Dpv7bKGe+95PK8BPIA3mZ8ifNlKhOEkqFDF0NFvQqBwnr1+H3M+Xtd
imRaVDg8r2tLckwiRV53Rm7xoNJPawMWU1tZltKavuqCcRz7kmACPKYYzd3rZEqO627KOrnAIdAx
T7MPcvHDCB9+iy5qOfYJsmXH54tr4+j8LkzhAJUsxzafpXjsKSftlSnwNOXr/vsrmcu707ZeP4un
fQ8mPVmpRRCfAfxDXRKnTXTH+SVgZwvQcyFukCybdRm6h0ZM12MsU3NUZtqFqZ0o2nce6VSl936R
4OzKbjDuX7vZMLqQkMJzyyL5OQZWoTCGraLsQVGkLN9B3nlmSkEqO4Fsz5ki3885PgqPFOlnElj7
oBQc1454it5K2NGG33JLsaVkF6urciRvKKGX08nelgjX14I5dw+9k97TsAnIjSr1QS+hlUyltEfS
h0orry0k0TZBgBVpES3d+u+shGbMVc+SK2IMi7Mnn77igCSxPaLZ+72NRk7o7Bv7uCPC4GLytf7Y
sa6pTyoYGLDjdMSedSDvIeYAyRQPdWJ6Ohrr+Ti84mtGP/Hf+KjV+/WBYXeQ67NHr6CBydmqvKcA
CRt24eWmjAN0o8iRjQxvYJiYJamWl8EH9Cj+Hs4K9OC+59cVVKi0moeF2AmMy5QKbqkCh6pPyxcq
KYR07WEKJogX3RybtHtK7DS3rmsqw9IOSykdKV8kDysK0BU/pakY8Du6Jtm5PuV5safgnp70aMw4
QgVPEGBpqIZPKRO4BMltLhk4H8MLWo9tAeIBDjfE43ZYlC9lZGSdnh2fqfGo4SrtQjOBrhxI6ZGn
ntYc/mz8svYeBIldleDCjhxbiXp/O2LEatjT0bkoekx04a5ygJLTp7Da0qWn+2HePadgLLcUg7hf
B/ub5lRi4BSvd4cF7UjZuCRSwCzMULqvdBOXkqBkQzQ4ITUdRYl2NGQKxH30U2MyngN7YWAZ2OLB
6OeVOv6cVfZvd+evTdAXcdNG1z5NWl7/BQ+7svMZ1mQkk9geuylGjirXnJD3+MblY+Ia5Hd1YW6C
wQ1X7Y3DYcT3LVGA5NEGYgB/q6Z9emSttslze1VSyeXJj7m8vL2d+ZnAgjIPllrxmw4Z/PELRYgb
ZWw5+yoo+E5J+ev2QhceYhXnOj+SsyfVCbtNxbljT5n4v7DuCCEkoBO+G3rV5opLkh4co63dncl/
dPeT9bzMu94tuBR0hlqenBGw0+DP0MUybsX+f0/yB/g2fMU6eolMZtV1ZigYFUNom8urDt+WYtO9
SodiONSsBmG6R69D18xv5nugbKyr1j6x6OUZ+zqNGoHl0WEpFJjNMfoh+bjJz7XexnsPaPtd4VTN
uSOCeQgLxuSPMmzlXss1M3kVYvqxdcqVAz4A5TWzFONWPz16mcRtxaGIp10kON3KoCw87V9L8kit
fi5Uk8P2Rsle3DrBQiNHyrz6SiuMnyirDE+Yvbbgw8RMK1gPjv8d6IkphKrL4ovQXS+zu8XYwU8d
0eF/Vhm+8OVLGypdP/CnU8sfOR83WKWQtnhqaaNKhmpr+l/0wmZJFwB+uc+9KIkUVPN+i9YlXpQ1
3WRI1BgvZUMZEBd9wmZwzrwR9M8xeFeRU35gc8AI7795v6n55MvHi+tqQov70MY4KRnn4W4F2Utl
WleDb/vBKnMM/AByUQcT3RCR7RFe1KvKKT+5Sntx0T9NVA0L35B6UdibDF7pZYXQBvG+7YoFV2SF
iClY5bZC38QwdHzUY+dcRTjEM9/JBli96AojxRq3HuGbmyaZ+E5LYD/6SruJv59ak5Q8jLZx+Zg8
wlX738V0IfqDwQ1hCks90WS+LTXRg84FERNK0M4sZknJELRR9Lygcu8iygfhu/1G9TsRidkQ42sq
elK6h6eT/mXEBBcacODOiRg/OxTZMLuMnvvWKYr+YFxrK51/Chx+DvI/PR4+M0uA90b4TCW5D97g
4+uwhbPun5uVTMcjf22PLMBPbXFdy7CRg6JjgkFUyNaVilv/XyCqkkBTrZKbTm4CRcgViIVDriHX
yLc7a4gdQdbYLQ52XO4hV+/Sto6QFleX7hQAGmstwtLCi38tY1gEJiNjA4oGBxes9FAJT5hxN7+6
P0Ox8v4wP+S5yll91NHeSsuiYWtaZNJKsLe6Zaec5K/bbPnx+ri+dquGpyLs37j0nGZLHcrRDeGe
cM21XfmJPf/vvbVlH0GghWsAYTgSXn8f/6ephtq0oRlI5FDg/7URXncgoW4f4bMto2K3lS3avLaB
8/sOUL/GHzywKFf8/sM4/rAbtdninV4N9o0QqZ0xyVHcjy5YKuu+VaVd5TMHWWQlwRtU+fRNCxwT
xGvhOcaOggSUqO0NiWJvsyXSICoZOI8HVBd/LISuuHn9batcAQ8GsLGPTBXmNlr3gZbBNbo9vjpb
r69AoWcIJ4dQGyTozPG4ZhvC16FtYp3KUYH1BDdJL2kmed4wN/5D/iCDr8j1/x+ASDlA6UQ1neQs
G/hInJ9dzT+Zhow0OVtFxUXZrst4oa7+KJe6ujzOFlblhR0EOz5h3njDdbHGW6Sg0x98NFqJgKLe
eLmfmpHJ65rkveOiEPdeX0Jj8xAU1zAKTMWky2wPiXrjmTZB5QU8FJ+IIguiIr9t7J0ZQQueksPk
0Ny+VD9RYxuGI5F58KZaqswDScKG6zNOvNpZstxM1gOVRyGY3cROBgqMFStGjcBjsJlqtjNo+oG9
qX+qOKMi/zpuhxgPdh8tH5tUw4bcomh8QLzKFtntsvr/OF3bsGAMq+B0xsy1cd+Hcl3FNRuXWKud
ggiGDVlXO+YNQi0viPHQkrs39kSSz0TGBKcfP9ABKW44FkzN5mtuPDS9aUnE3csu6qNLwYKEsFSW
kKgvV1YO4WFozzZ49AvBlifAAPmPaZfLknW3b6lvjYn26J+4zRqDdJNqIXlPC+j8qble9FchToJw
lbIyZOOfnDMAzWdVJIfmbA5+IKeA0kcUa+Cnq/siR+lKjkEPcipI/lWC3+gXneBLZZ3B2vKmfmaV
+MY/S9ZKbTneLmqleq6dqybL1HRaVolrervK3qyKCWNdeRhS0QHd3OkRwtp1ihRrUessXp/1nv9S
z69iLzJTTo/YnZbN+PZWjDpDKwTarASZowbMFd96p3ZXG5O0yp2Epq+KKDNBhpIzYKtLaxy0kCmp
qQx+jJBfu7F6mVqH3no2bJtQEWLWyhemLByHWSWFOIcYuoSGKycXTMODFauarY7yLCMOEzKI2Vuq
rNo7LpMfKQaDFJekdPkNhTGVtjxCUFygqzMe686O/DLQbs6b1eOLF8t5qqVWP1GE5DJZd1YPhOAu
bs30h+H9AgalkyjI42+vq3nogJUDLb5go9xhxXyeghFWbNDdBgUwFkA/+VM0kYlblzNBN61/Sb7A
0tYdzU/9Oai+Wk1PYwcj8ZXXH8zUkKPbiVN51PEL6GDHG7zSjl9IkGr2Rh62VPuVeG2PHsaX4IPQ
2bP5SyePawsDaIzNnrYXGHCdUFdwKhj0vh3fT5/QXxYCVEOE5+7GrDbHnS+znyFGlLT8HWze6fOz
YM29dGd5mgSJMu/iPNThme5PT+iE3BRBpu8aQYSnpHglUVkLWWJtbW9yg8VgP5b1gqJ6SGeFauTM
8Eegw1vQUVRTGkBq911Cg3yC6p3bURbDTqSFbP/TEiZSdmLM6GSKhfN/aEFI/YnWnRrrLkvr3Fop
V+BxLYuN7w0uQFj9HnSW13IdntAfEoH+eLsU9b0hdEPIVKn0UIkaEnj6DRzWyo8bQjznw42g4Xtl
LdUhd9HIhga5CEECD0sErmWpgo4ZoF3FdzqBUYrpDrJbu8lLYTyZjpTcFL6j2NLLjCU7sYo3E4aP
4M3ZlpOxPWKP8YagxDR031sLNnujMMdEgeEAqjqxsuj+VKI4SbPMlRkjx0w6qTw16be3Zvlv7kVc
tl/ZXS9t6OuJ3ZfmdY5EozLkVMz1PzVk2eTpeB6IkKiARod1q0u7RShCz5VqGtdXQXgcfEUK5ux3
jteoWC8mjxMW3nT6qXza9aFZmhRf4PLAKfgRo2SgNz3QFlZOm033cHja6pwTskkqgOnVbbSOqPtF
mU0XmXV6M//xa3DDnC7gD4I+nmm7zV1SczLEbfgUZHLd7hFqF24QDlW4uGypgh5xxnuQUURzUtF5
7HfRCHi9SOYbv6p3qO92wbWPwzNaNulweR29miSiZmmRzJS/9J0NpnEM/IOezaaAqvqbWfV8qTC2
+hxCJj5uBcbQk1hltLt5cfZSM5jUG6j1mZ5nBmLAfT6d7P2ms5aqjdGAcUJ3wjW8z6lCIAGjevhW
UQ7Pg/pW7CeWSnXdZoad6SJjZL55vEXh23XJCiiiQCLP2qGKFULr0EL3DrQbzHWC/gfERujHNmmP
t9/0qYB5ktTjV46wUqMguGA2FDOliONiuJD2tlaEzQeJcHfbV6+boDoSek5vCfP71f6XXrCR3hhw
ftRBIJMR9Ws+Emm5e+F5RecKm0eUMNUVjPcN+TFx3cg9v6YKH2ik5lfpAI3sPJpneI0rMy5EQzCq
nIXLTCW8ma7UHj9SlJoBOPRAw34vUQE4XRXYpivmVIT90FnR0A8vzDvk5q4BHIA24uikDFYOCu2S
Sb2ge6TmkKGHqzlsoLpPbqzFPzl1H61JEHZ4ciD4P10T/M/JGDqxuX8EvPxczDVHTsZ8oRis3zkM
cMTSSvfPuuAC9GB/OA2pigzHMQGO29ztFZagyxkAgOmfMmRxLD+VEuEeimpB8MreBlw6eqSMkjUC
zDN0OqguWMB68aO+uN2atS51aJjG0yRtgib2L+Ze8ZZ3giQt70reFVvBzS+t8MhuyUwfrlQ3tUub
YHi3tj0F76FFYxG785zj4t31HmXme0RadCAuoKCPuu2Zcbv9Aqpag6pqGks1iD50mYBVrl62wHjJ
a4FEtIRHX/mYotbftuObWriFJqTIxGnc/tUOlYf5HvB75kHbmcxKJoO1OjkK9Qe371M+/3yaNlNi
730AEze1yl+0Oamugebfgabjsv0bP5CsaPW43hSeqsVF/mFxEkeHb5dIVxoCE7e2/kaj0RCwRlTS
YWrmI7UaegLeuLDoOO9A1N3y/gqfct2DjQzT5gy/OLqg/PV4CSpRigN2TF/gEPKKFB/KdsOVys6e
6/EKe42jKeSxZ8D9JFdzoJ/dWzVRadAi78qjGDlvHjqH9Gig95+cC8OVzWXowEj5pZ/LCzQxQ4q+
F5IiDYVVLbXbXLxSuHaTgGcUEWrdnSN1amaGl9677cNEwajka64r9dkJ8IWwJP4L1ssCAy2npj+i
iy4PbnR9nEKOj0kRbTtmcl2X3qHJ4Y5w/c/paztRqqRddHpU0PowlD6VySJEEN7FUGeXRSj1NewR
YfvlXpn194f77Ec/6haNAbQOa1L6wkaxVvYLvK/+rKEVRu3vUzCMWW6PTpW1h3Eaov/L7SjSrJHd
gndTsFrkgHyd3I10nWoeQYoGt1QyQruhImKpGb67rtAXwVZpAziYZuSKX2S1+GgsbHKg+pUAua0a
IkTDj12G89Yp8OP6dQkYJDbqOS4WO05brTQi/+XdKc5u1Z+q0au1cP930O8CjvXLiNsm5N/25He1
sK5SXbnFKkJ0nsNvcbZWi2lp7Uzrse5fTUXdzyKgvDQ9pyUhla7r/D80XbsvVmrItWvEzI4z5FJF
0Q8XuJl2z2e8EMzGLae6qvvNYkBIqmEDks810udsz/Jr6wx1krylYc4KZ8T6728lqO4sqXN24sQs
j69JYaQHj3Vjtw7/ih+bOYRjc1bdgJ+iuC0A8f3zhNfGc8UbWpX8XDQHArUJm/8lxBpb5MaThAJ+
5Sp1B5LlWkAvey5+1b2j20AMPm2CJBF+cYLEBe52dOi8RLQ/PHkv9LAlMe6p9XMlcVn6/lTgOZTR
yzRpWfC/Usci0sgt1HFApv3XI7wZe9mHM5ftPscZv5uLzsSalbC0n/NeT4N6daHlU/P4tu+5s6cT
NorfR4fw3urh8BNGjD6sBan5c7THBDurLjAcMYCXR61mUFfKWTVFmPmqEu1FjfemkbG0iaSns7IJ
cTHG0E7zPEtNqId6uswY0N/Zo2QEzE+WoBkuoelUO9Xj6RGAOx6XWTGhX5gO9G3wzL1/FGUEMRzj
wfHiN7eMSwxcjvRl5Ub6Q/AEDkOxch6hKYu1bctYAx+E7iSpr7PSy5UypIm3kjDhqXT3zBHWrNPA
R1eZul/lumJ8Gc5RnSIaqReRcB3rBj/Txpcf3Sob7Asud+7eiCno5Wy9iw+l8R3gjuRp5XJm3M4Y
ahBy+p6eMxmYmjQpGf7CPpSYNlYP1WTIeK2g86HKMdWm2749toMN1oyKl8bDd0GgMgqjMPskHDSP
9n0KqK3u2XI5C0TFg1JLGXw+A9a3k15OBOx2RDw/Pa2yecIfQ0c0+KldrCT3ygRL/7cgQ7V1y1yl
YcHogGVD9ElLz9lkRTit/lX4hMwGcSC37sM2nJs08qeSoAP74hDFVKj0yOD5CgAx6DN6eN6yawyX
39QC8XdLzUjkaDlVGehHMQU7SrZI/Wpa60BYoVztRzXwaPWEScSlIHtOzvll9V4GplUiHVuzwsQs
xaAHoPhNscKpQV7ydR9rFH3IJsnDN9jvm/TD/OE4yQFH315D9h3bCTBwkNm8w96HA0ZniiVuFBzq
LyyKRB4Adf+x128q52+wM1hRaiXHzFsF2R1T/YDamK9LiZGJqzBIMinU+Z4h8OXedOun3ws/4n49
+bIMMs41vh8Qaav+ynK5Xj5e6VqtZ1IIL0d2FAaGrqVpULpCzn9vKlTdvP35agv1oGKKZz3+x+zj
v9ZAu2aEzBSyIfMOGzZhFC+3oYZUHbEJqCs2WSUh2bELwvmK8Kt4JN/JdY6sowHF4ih8c7XTCMer
6Uyg4I5qOFRUKQORmUAHstQIWW8YkIZRUOLslu4WVVGqxFUUs3MWoa/yW0gXaK8UL0vUlX2xtqi6
fyNFUkT+L59cFWHyD4mYX3/oJqsxpft+ygAmLMk5o6i7yV6T+BdUqR9hBMH6MhTzvQt/DI4oOmSd
GJRtfBQYrFnWtBmF98LvyeraPrVqDRFnYso19oRSWL50r/v8p4l7ZwmqoNXVP1JRkp/8vzL4E2Ry
LYN8/h3dH6MPImwePnALNlmuzBbFrgbDFJGGwv5laIZrFqgCD16pMiz37RO2mdZ3Ur5FAdcfjvlT
neTY2+JvXjSRU+rFtkqU8/K1+0XzPjdxdBbOKd9Nmqy6w9DoDW7sPqzXbWTEIzCXfQX+oW4B64kR
vga38VsBRJkR+Y1MUsJxd4PxqdQOcCJxVDwPYng0GSzJZHSyRQvdFih5VdAZxiv61755qJSVqQlY
ehHuTJ5vyIdFdAgKgXfR+k1F/uFKgLzZaAmz+aCdW96hgmICD7ta3DDjLpCxz8S+2/Zz1BL7fPUP
RfLxehqaR8E8pGl/CK6TL8Ynx6Ktke6RM8r5fv+2oOtfdwkcRvRi4LpGUTWqtS6BO0NL4hGGSYA0
Zt7JDMsCYPceOqzr9TKnVID8mhv5LzOWac4RF8NX8kLTiHL2IJ2RXtIF99jzoUFDmKXd1z+VkYl3
gTRHcMDbl59yuZLpQBGUM5v/vrIX+b2B97u2JA7MZNxeyDKTtf4HEDpYf7ZvbUMXPaWari7y/ndo
BozshzLa/PhJm3XltEHQEUUPyFp/BWnshGyj+Yi40648u2lF2zlnv0/EEGY/idA/KmyuxUpbbjpp
Jr5agAF4GzhbDnx+0Dlz0w/ByoorSAmweLGJJe6LJp1NCX2SCU9NDG1j+jxwVkvcugAhKUFhVgCw
CC6FJHRMTJzuQHbrF/GM/ZeJJuh4bKikDax5aVytKYsGNRv2HGHe0hZe4q1I1zq1Wi6xGU9pUJtK
V+2vIPuEr0FlYRO0ftUNHNYVCiZBR79HJlh3dPNJ54jMkaaxJzl/roRvgxfYAN5sp4oWE6qIhk8Q
aDF8Mb9r3u/g4vGeogTEDg+CwDdZ7b2t224VC3cXzpYgYTbFI0qfn2f+AusQa1QGXmqyvcYF9xmW
sISugbbHEcVOxshCQpoEX49+a1Rv851mjZD3SH2LF+dZKGR6gqiKCZ9QbRMyFpXzYw7j+Ul9omSI
kibBC+W697HKMAW3ofvvC2GjHhHBIm3ZBVF9VwdmvjfbMB4F1LaAY6BqrJXAGPbkHD4gpEA92Zaq
4ElbpbSR8B7eaXxD5Vbf5ePZw1cpMGqkJx4zCuVEcP7HDUDayTRxtpzFg5XQdP0xCS9DbluPVrAu
gTXm6HWqsrwIyDhGOU5utI76UYkXizyFCv5qKB0J8gDVClRFPXkO5F7BWQDoDKqpAf7wV+p6gq9F
Ra7qh6wI8WKIvrsdB3LNf9uMeOsDpxP4RHGk9pPDYlFj96qQCN1CZt2cTctwfkPkNO1tVaZ118Gg
tf56TRrFuxDGTYTrn2w00mDHZTWFt5jzKP2aOurMMu2TDdeAFtAu5a9Zt/iZd8Yj1ZL432rOMX1q
8J3eIBuTYDIFSFgH66vb9fFDVVNhdSSHj/m7tp8KXafUuDK5vk3e3wXOj3F7/baPNmmfHa4XrFA0
SdtpwnVrBfIdYnoDuvzkHIZZgigHkxAF95R5dPCpT3TsqXwWYF3Ji3gwJCcYL7N/dgcyBYRfKEOM
gJYkCVTjVW5Zz5lMS1pJUngRihFUP97eLR4C5q2p9g7ms+r30AVgbwPH7XEr182dZ5G/BAs3LZFs
p5abu63y6rGTZLym4j7OGrOtEpplM8gChp3zNzJq9lYp34B9i70MwCgc5cYESkOOB0zpW8+HWJD2
Gk/8lUTnmVkBgJ2XVOPVR73VjQg464OWRf77BMF8ZelQ3pbUDV6aZcjINC0+LfbzjXo+wBPoFP1Z
FZ6wBbGdZlbCIq3dswH7NNbP4yMLo3+pB7NqUc7/TWY5oWhk03YrEHqp8bIzkNQbWsD8dak7lDzr
1gwdM6UpJLx0ygrrDybMOO6fUiAf5UJU8hImO7ImhCkPUpn1NVqNYzNyr+S2Mkz7Xsw9k9lZvLNn
e7y2WFcme1Mx9NZMXZmX5agXI9c4T5z0iveVmYR6XAQve79QPzhKYz4Tc4FxbgcM9YSmGh2qKK2+
SlnRSRonDsPLR9gxY6Uxhrf3U8ykfVtxtqAkWFoHJZrkuZrCWwmIm0o3vestDOgeTdLVvpZoU+AG
w7OCIC5RQp5EOj9zBI/6etMjxCOVUXhhqGiSqy/F0ObrKbnINktUBo+a5HTV8j/Aud+j9PklMFnn
lMril0beSYq7kCaVmCuZDk53+NdMU87pY5ZRcV/MvoIBRCKPlvjfoXmxYfgiq96LCt4306bl4CKM
CKNJOP4DE3v/XW5M9xh62CUwkpsxmXQ82QeZJi1mvgJwPGhMGiCFy2r3seiPJvtJ14OP4ODF05tV
sgJkSYVP77GZ/7uFOh37opIrZwbiJn8duEL8JYM3Yd+vJ/evmDacbiXC4yio5Ts6cDuMzgIOyntk
5NQdEWTiCJC1lwkzg2l4gbpqI756/qeAoAYZE76SieT+sHV+iOBqNYrn+mZDJOGtez4F22MoY+ae
D02pR/Up4jp/XH3t+PDDmb5ntBr1qZJ1CCi0uK01sZJ3pLwRTNHR1TeFi5TSzndS+lFMcmASRIbN
mjRl5lYOMOys1yODHa1nq+uq90vaL2zw9aUG4xsYC9NH5FuKJgSnwQxfyksvWGVGyZjnbytXGl10
MmUo0PUZMiR11OQtLwT0oZ9y00cyoGLBHyGtLAHLslEzvCq/k1yUi/Stq+FXbpSR3xN9Raswja70
Bt7s7LPf2+3e1GHVSRZ/jZTP6I8/hU07csLHcGo6btN2rtUq8DKUvtxpUTHOjI8V/J6+Tlpz076/
L1dEhhn1Ld5CKCe6fsc9G6D6bcVo+EBvwpKHPVTySwwQsLGRBRH01US25y81NLS0pQoAakOnzDdB
WMznSd4yXB2DoKUV2VzzFM/zZDX3CVjZWYSh0sz5CLfy2Gv/4ZPggvDnW/Oc8J3BqK0AGxOiCe/e
HWcAQNzBB2/a5pq3SsHC+qNpH5pG54VoEdyB7Lx6XZ8vAsvLSmqCGzYGJhk8Vyu6O5tu7333tNYZ
d1FlL7ZBxdeCE7YolkHqZbHwT6aMgV/ThT40wBbmou/d05ziKeIYixP8W6wQ5/6SEP5O7Xt8voAp
ZxAKl2IKDBw52GF4DN223GVqt8XZiCD1MM61D9+U5bJ887jhhWwbgPzNKBooQ3V4kNw8WM/xyxzH
TTFObyf6WddrHGbpvLlgYWZUkOnCMgsFKcbx+Pw76cIRl4D8RQS0LQCdml/tvzw0Pu9y+ojmWM1O
1iCOYRakPFaJV/Q7wBlHDsRabJXovv7NS4D1KLXXu4XIp4d35ms4jsIHzhGMTOh6yVBwGt5r1S65
+OVyaXMiVUA1H8CGOWJpn5C4riBZWaswEkvkXMC0FP0rspjfNUHcCJim7jiDMCKRc8xIBHzQaKf4
pIrbeSHz+C8e7QMuFbPjs5Yz0NAo1Vtt7+OqCtb/OHa6FZBieKy4Gt/wxe6K8tTog69s49lej60P
0HGzFl6wLFT4u3/lOgsOSlcGlgh0Hbb29HhU0DqZYQ+YJsnVOaP0cTbd8U9yzb8fE/viMqtOi+QA
+df61/vuP2GpMfOEiwxIIrNd4aua9t2fw6gE8eqImPynO46vv41MdiBYz3sEHyvCWkVCXOG1+REu
sUsSyGoROkNrN+VLN+VmFAa+X2lR9Fg1yiXzUqS334e3rujkyMmcZnXuYdCB0YvzmxGpf6g3CrJH
pitwSI0xhhOCqymLFL3imsLn5xmAA7Gk8nXeKCkHlsvXZYWogTNbPGOHKftT+vEpfIyyU68cbZC6
BNTRlCEMQUc6h7muQSJ3e0E/KoBP5aLSiRY1PvUqns3yyvWmrVDC/I9vT/QAjwrUXRCbeTuY7bOk
koARv1HGmZKpU/x2m119cZXDYXXix/wCJCASLzLHMyaZIjO+91A4Zr+XUlnVii2wQ/AVSTM9j0Xv
H9lVKsXPPozET8cj/YOZ2Ja77ydw6L1+YHHc7r39lwRFLyKKWrUpUBETadopyquiYVGnvuS3s/u5
T2zWWhrKEgP+bQzI1nX9B7v/cj/iFqiVm7tUkd6KaPYGzE+p53mi4Og6cwfhqkJcbEfSQhFKQBUw
v+CU84v15f2A8oFxVI0O0W7MWgZyt/96QVAB6uLwkBwiGkNihO/Jj4kLFHmR+h/KTTm1lLDk/4uG
Dq4iojQEWfyB4NHgpMeM/2ajMypvaVajADWz4r/fsA7NUZ4ldSkaMPIk6i4kPffmoY6tr8U3SxUb
sM+bSjIKrx2mCq06nPo5977x0u/rQIgvWJOG0TLb7HzVCkVdOUg05Yo4XM0K1yfoowzJWr9AckBe
0LCCIcv0cZwutKrNfQtV1E4FE/X5wjM5doVts82n9cm9smYQpzXLG9aWopxgR5ePVlPDrOOmR5Hc
hciaThh3D33wJRso5LMErCOpDXBwnBSnR4yonRLiRLCiNNnTBouAgLoYFQrfzey1VfwAyHl2gbIi
EDTPBSGz0W0jKTUACoxeSCsREhqhabj/5f27oAcSw9/C222jMk2GXSJVk9KxtJ/wzG4jcwBmhPul
cy7+dO6ZXYNO1DrN9OL/DvJz+FvLZ0OBErveVcY/CmPvQRzQlilbDlfwgLd/1/jPh7FhauVtIw5d
dye7S1ZM7+aCmZkmk9iry6GXtYu04cbQvZxg5WXLYAMLSKxZ8XWVDVd6VQquMaaB1YkGXfZnJavE
wh7JF4XsQiu4Mm98DYxxXKoDSkHVY1JpJE6esdEHSA+oourMECKuYHLgKr4ZOc8tMFHGkmNsjOyI
UhnlMLnPfMS/bQkrEgTcqM3lR4mucJisIvnZlME38YbFe588ar0Kyw7Rfb9pPR4gG5h2+QbulfKT
MBeFCZVRjGAJsvnew05QR4wO/c+vwFYzuF8j2+MZRvy6BIoJYMRv4kFgdR0TKKU1U1vR5EwQPprq
2F6U9Eo4+lSEucIS4FHk24eavSwAw8XwT7B4UrJBlJYR107tMJRLZkN5101yo51LHXDxkK464EbB
OtkiKJhdLFxURvj6h94kIMCn65srYWQOFfySLJyCaaMW+R4h7dWYBqpbMOZVZ411GgquY7z5ve77
KZ46cOeOlE9rWJQw5DKmWIEzuyJg3D5UnsXdeYVBMBcEh6IlWbsF7uU2o5NJ7GuIt7IPUrg5noHG
PQknOVfFiqOctt2/DZRH/kcWFLHJc27FdbH5IZyPx7kflA9RXqXS3qvKeKNvzBetrYcKU9h2Xsw9
1gpMMomA4S0Wh3j09g5xJZjPoKmImaFqJ5nnvr6WIFNjWWxjSrhgdiCd8ypWh6haDFoWGs46BL3r
ovPL63eS54/jFP7+hjH1PxE6o+z+cLKjcpU6PM2SeAePVAmFu8q6K6SRA5DqBkZCATeo6nPDWrps
67HAnfcCFBhf5xRvzBwaGBHh6yxwWz4uqChbFyMd4SaCDPmNMjo0455y4XKQDTmWGlcbhZdH/bsc
tC6/JnwwKJjAK6Pa6h/jun20doVcvkH86ScvlNYe/6iNr0of7E0AFJR9NTTNi+u4ir2vC6KLdm5r
TiCbHRxi4OqQUCTWxHKPL2JD4kaVt/3/ZquwQYJIiAkSxvJdgF28R4cL4cjonNCmGJlhyXm6JKTt
plF8hJ5w4kG1WHwk+DiQNENkWfcoCWcE3fI3Z7MlnfVwdc0mhpYUnEnkGE4uPGmrJqJJTLNub+MU
CZkp2M3pm+gAZnYzNPLFWp6xFNTbY5r6B0eS8ShRXIKwrUPIPypkV5nQlhiWz6jg3/15YMitdAU4
SFQE7Yo5pmkHfCFNSa0ErZMvYfb77WoVeTT1Csbx5ifA0CQo9Q9Z3lTR+CadVw8So2hAUiLgJKh8
NZudzNlocfG+AVaBljcsSDyBkexztYKw0DhveWmr1vCNAxjNjPAtQsniz2amUp+oc3HRlPnbV+gu
5+kOK+wnmarPSY9aig6GOB8RCCNBpENDbQi5SuZzLcOLptWM5KXS0TQv3K3u3X5VUe6RSRfpb5+N
wQZE1ADkWOsTFKPJgSxy2nBv1SQL+fBaiY4xitT0gggHa6D5pvoAcpGdoW3l9UO8MTeeOlejO4JT
TXIuKfYESFKOQlaM3SfwyK58eWO1EdBZqm2GjLnNNljPK14eigDEyYnGUNDg/OFS9CiF/TRnSU5N
zlAxed61L28FygQl1n3pvSYHuVPiEPFsRZ3zSx2KFWZVghp/hOSSJp1byMTsr4xwOp06pXxgLrZb
XDdHQl2IFyYxU7lLrLEkZdsWQW1uqzV0Tj8mss7pOTdFPWuYzPobBGYjOxd5YV2EhPhdMQvrNwsp
iuymbUi167B9PIFjhIzulvKhlJqISxzuqsYVLgmYts0ype/kaY9GSn5zUopidIlrcKmdTT4gLdY1
QW7u6rG3rzzfY5D2UTESmRNu5IF1E8FiWRFuJHPuPgOjWYIDID9QWspcuPcOIQmKFWYOE/HqSivc
uJfdXDheia0OPSJOkrmEIsvn+hBVssOm4AYxCEzoJVVscxL5Kwr1pZU/lIhA4UsJsyvq9yBed69a
dgi0tvwUb0EeRtSzCWbWs9mdgKQfeHo88J6kn+j+Yk80LWgs5G1k5BIMhY9GalZnRMmsb5BgobS1
8VgOHnVx22W95WFmodqCZT3tPNgtvod4sYzHmWqKMYbFkpHokfRTDpqLtIT/a4lueaiwLXasmeik
fJZdTwKvd8hk/Uj1N2EPMc9ELU3PIwwxa5DPma9mxnxRJ31UsmDabJdcF2NztETryECVfH3APNcB
7uQivev7/qAwNDzFTrLJR78jwu0nrRLpwCYYxwYL1LRX/DMe2HrB3OwhmbDUIPjwPKO8ZwJA92Kc
P/h1YDIYhOL5h0b984bncFCf5W1vH/7PkncsP5sE4zepB4SOPqsqEVwgDTAFxkiL7bupjqvjgSYW
MbOpY0sNFOBptjYjLigIcwILrc7VMHGT0RKv4PJ/WS/WDx+tDi56B4CQ2FcSeNXV2DhvgRw9WWuK
Nj8MQjSk+apV0Z/eqrxElQmK7NDksk9v+gyb0lyhUOg4/ETbpanFctA1vVHwisf+kBxNjuQctVUa
2JUbwzJ3myXwgUGO2ifcG349a1cRMhjETRrbIrlq8YjsV2y3MHMLxZRCtfSW2hPWfOUyOU2OsdxA
i2oyTInp9eOSpdCFDibc5OO3eo2qvDZrXsnQKb76zOWwiv1OJzzWZC5UGLcooBaQR2nTlpE8tgzU
DjmAnZJPUWmhwjEQFiLthZ+UiJxuDTfslE6qXY+wsJaBf6Yd0xsrqgwIv6mgM1/Si0Z06NDn5KmJ
tuyOsXReIRpCFTFFKb4VGPFED0zz7/5GvPY8sBQL45phTz1G+9o99iayKGFKaAZ/nFWUp75oOqAJ
1mOvcn0jgzVEJSckW0LPgGfWe4SkEl0bQOCKBnAmj3Nea9xIqqr6dB8s6tESHB2csi1eIT8+SzD+
AA42zcz9PAUITpfYPYBs/qbTJer1nW/xWZg6IPK4wrUO4J7u7X8JFhCbqtCg2j8yhkDMvROwwueQ
geiC7pcfP8OEfbTdBXLSNu8ePOMu1tvpSdR06TGcV7VrCqHlzUeez7REtZW7r6x/Rp6A3M6C/MOl
qi9fg9rJRYHcI9AaxX3WIoI2Zj1SZH+XqQylZKlPdd118rK2XP9mB1dFvZGPxVc9VVR5tO5vepu3
yQoRDM15MKEtn5CkwP9JD1ItxXDnfqWwpo0ySsSCIgfi5OPKQQNW0VjLwLLq9iwtKO23195ONCMg
CbT0RDwV1D1F4SmD2rV5gFrtC2YNOkc1SzYHRJLdwbSzABNaIyZBZ7pe36Gm9IsnrZLotufag1hD
OlfTtrPXZk7wNMMRwrzL24gauJHz7dfJonQPcn+O0SnVehqU+vuVEFVvrn1gBVkba01EAc2InAUe
GSsut1aciekOtTF5TgXKPIHoOU4UefuT7+f0AsaPFUwZGxTKdm/OJS3HDojDcMZfKOekIgVbhRxC
13JG/cuIvak26EZybk6KdJUw2+bqzXntmUbDqjdbUhcX62DyDKT+uyqCWD0BE54Wx9UP/Z+fwZqF
m02apxM6qN9OO7AOnBepbxKiTTf8kkP/AZiFyF/08eq8MFF7eWaEm7BClBtkPe/2Qqr4WayURUAM
U0cXIeEH7BZT7V87YubrrDATZWVS3XQ9JZESo+W14i5Kzt+TnF+l70BsPRtzJaUpq43yYji4bxS2
q8ZLTDp4yjXM2B4cFALTl7YYnW0UyQGTexCKSOxhpwMTtxWYHlDpS8gG5Qh2qidDlSu7k6lkFTgl
bb5sLdYGzMGTXy6awdW/y0VMYh2iNztpPR+OhO89xHRGnXYqUF/uiggMQ5TVTfkZ5fCdwCuimSee
jk7ff9DK/XAyysI2KSGh4TWEi5cr6ezPBn2aJn92/Fjj347sjp2wDMcaCkQ0Y7phgxo+xmlZl3cT
2BjKJWGbf/zgPIvSngfcdyCXJMiYI5g4pRHTCDx5z9hBdQXIK0JEfiJGUI2D7q5wk0KA7dzxdGxW
FnsYeulB6c1B1BwQ3EZ80NzcbuBgRGBmcjWxG6fk3CdfL7rSu0l5mbX5O/gWOjOsst8HltySMRfd
aohJlOpZHVs5wyoJhl1iexO4CeUlV0jOjSnmfbKQwKAJTTBft3Xnl1OKpj62y1AmTEwD78ezarkp
f3RA6e76SzkzFpnq9ZxhtFHlyM2hK4/aPhagnmyWCUTKW3d9KyF85QE60GQcTpFuW7Vt0KsDWqV2
tr30vwNDi/QbWHCVNgfMU8YN4/7FiW9Fs7rddxgeGlis8tiEXhfRXOQqkX+txEAHZcEW9xCYpxfU
DOWStQqwKLAINRGHW+GNNlq7YtkX4HfFRHaEdaCTQ/nAL39V0mCvm1n6dGR9hDu6P6R4DJGdRJr/
JwCbi0Q1fUtfWS8aQNEKfs/pUCIogr+2pqtTMLHYdBou8N0ReXergZAOP3Jk4eaA/9rhtc/lEVBj
9JssVNZPrlBBqTV17XY8AuDSKS9dTLnHtJWownhBxjxFfq6N0m2V7u53cmcNo/U4BnbvwHgNumex
rAyjDpwpphu1PlcwpG9DzALj+Nufe1Z/SrPNrTDj6PRaPSvRowzwkZHT7xV0X56+KaX2cGOOLk/P
Jr/tT6wL3KogECIi/1w+HEYwZc/d1ubHbKL7goJw6vwUnGfW+2ohFKwRzQr+RyFLnawv/XUPnqB0
tdHgCr14iENVyNi0Y1AZA7mEt7Fmd960UpQ9rXGjLI3tn/kcde5P6H4ADBVVyFUQR4upfI3gxoot
y9gE4msTa5jcyypWUfKS+pV/6nDSOyhYxT30WhF5ryBOaq9bmYNv0mJyi9IDV/1VQwOcDS4PrThP
JUWvpaLeQ3RRtF0yMRqDS7w0BuG/Y8oNiWtX1jbxWif1jhSyfLGJV21bpVfAyya8EzOutqYEIwW2
+aoxwnCRCIro5LQ79WW1WV/Y8MDqlsXVGNivVY45jSfDgMEKuQJSoqzys+q2vepPg/d+0LcRvTYq
MtiADdBv54FFo6hVBv55pyZ+iQ4lt2/UXFQ7DA5/nltspWuF4e5uqbQpqE5WzTWOZsPU2kll4n55
uEkXP6o0Z5hFCCPZbJgFf+c2zOt2040MwEFCzKaJSDOUjXF4ayPjN//BrbBicw1S9rcqmtjEUPQ1
GcvkG27W9U/EBamuhFAiCEx6dh6m1p2OqCPqBYkLKaX942rxQOy3usCWh/l+JRGRaR0Qf/1SNUyY
z9pBHvA1D+TycYzHnfUA3PUlHiE4nkxD8tJ00t4Dfiuuy9iO+aS7Z6DH3jOMp9CMbPkCJM+zFpX+
nBJas0HXoUaSNQjAB+pe1SmBpk0Sz5Jk4hDz5N0sXsdy3+ZAAE3QfvkeC6InfpUgme3jz2EyOc7C
eeyIF4rPBKnPWcUEM+fkO8Nx40LbpZqgPfwHKL2Fju7huXE6rE+rVrbdpdJOqlodXHg10bOP3pWe
GEA7RAxa0LR5V/dbmfrkPO5X+sqtTPCyWNcMfxUwcpRjNuY8290puhyGFChdv8aHQannJhUPGxNd
ZPDIiCaIQ+abrM2lf+na1HaKby9KE9sT1FO3S/PT+b+VV9FiDo7cN0rCFa2AjRAB1s6l2n9NRuyW
m4SxBC81bVKou8PfowYCnD+72ubeMn68fWVcCcFpagjIoXsTjBgZ4mioHGI6EKq/v3TLOc7xe+Eo
xlhX3U1lovTwecLzCjZuaNmC+0URwBPKJTMuTGKm/5YJS2BWO2Bs6agaGuaei9Fppr+COuYe8hv5
8tHfVYcVTKl8hCAdgpV4RQI9zVVQ2HI7T/9b9hTR+a8MHg057J7++lLDoYfyTRn5ylktqJmPSvKk
GDJ1NMWYsey/CbZf8bCMyRGWecMAldcMxz2wH2HKHCp3BICQZ7JWv4855O6Z0TVC1K7gh3sFEoGN
A8kb5plcigpZijP7AlCpIDJT3fYS09NMdvXnQ+hoh2SWZ7AW7zy08jlLjE3tEwLfwvO3e4Z7sRGz
jzUJvbGwVwLn6xvvXYQ+8lmLSEOSB6WauvJ9G96j35dE3TPsTWlWrZwJ4Vq8AJW/kWpnGxXBFgpK
H8D7uz2mPRc+fTTksZV+vu35PVpOtscZsCeWZ2UcjDzdmkYIZy6KU1vStPjYi6E0y4qwvdtYbCWi
jomsx0IKGCUugSbSRo59V+Mgu7+sgIcx9syHLwvykQO2lGMZXeutlLpFvER9tAssq3hPr5Bz5FjX
pK94+5UP9hiel4WwlMExsu1QybhCsLbvf7pcSIgo1h4HaZn0FWRs0H4tofRnKeNHMYRRZUpBHas/
gHDxk1jS+FiWKy1jxAGUN3wUluqjzjaDbc8TVxS4APMuxMF97ss0gWpO86aekDM1nziYqwEqrJbG
FY/wqWVoQwqatu2n+RH2wyi1FC7RuzQRVsuTHg9z2ejcXXSQOphudH9bDcTrtY7d/czQpluy9YzX
85srQ1znaJ9gG830qvkHClf5pAf5cc/lcDQ6aAZPlSGJP78kasVdS588S7tXLzi2XoSbeJoXQDVb
A9eb7gSqLJbUZCXBSuldlBn5p+KFVSSfiCcvoViWRzwHN+J3WJgOdoI2MOMW2mr7KgzYTsiE2ol1
UUsI7DYYLm5a4YN495r2kqaQYFKKwmvU7Fl6RaYHEIbv0G/klyBWq+8DzX+ja/LwLJxzsU/i7Ylx
0wNVPNzPDk2xVkNux5CYVtjK/Fb3uZ2ORnxoU1R06Bx5xQv5JSfViXpb8ljiHPuBd4MysN6HG0TC
QDMUjCQgnbBqICw/QxTuBRhYx+Lz8caWNIy3J+KuRevnqdtR9mlmxVdvdvGG1Tnn2mjLz/ztUCkC
ndOCpw0j03IgWxac7da0hkwCyv8SmKngJd7Pqrt4Yt3GW0JX2/wKGbuBbFYgcVG5EyDTNTQHAvSy
JEoAn1fGp1VkSy77fBeaCJShCjIJJzo64xnTSMyuS2KaG1XAUmOEj0hYaIVqDHgSANwjCBd4PJWD
KNaX3+B872/gRVDYI42fzXxCfb9V+jPHh+N5zF3+n+ZGRiDF2FBazYys5RwSMUFpQbRWdPbiVgFq
q9Qs35tZUXYIU5lQrcmJkZ6gIAcMcgpkBu1aSYGL3DqcOjvhIUp4jD/Qq8GQ98VL75Y3xUOOkAu9
f3BoYwV5oLPubyGkR58RXOr8pszSaQ2VDTRHjmsjABwhzyKYRhmNW1G3/rjq1ab4ilWvMpU9v65Z
5wcAYAP+43eu4Wc9Bfz6cvILjG0ZLlATvM/fDXlhBF3lb9jb5s/Y9XnpFYnpaX24XbjpW8nlDbK1
Y65O6ZHRriLCryeVlGdbdoTjSp3k8nIL6icN2KHLoimLovMJGs7o5MZvZZ0V8bZQz8UG85c1bXZ3
0eGmM8Xua8czVEHT1ylyVnSFu4la6Iv+mmWzTyyPmqfNsXIBXZUkQ07wdVDgGN7b4Vu7ESU4iFI5
bq9moa/+C+G2Mvc5avh3vDZl4rng6xT37dsPusLddcRm2lRro5qwOTjSiM+R7N1jOUFNLL9oZXka
7OeawH3nb6mlarg/3s/Ch24x/LhlW/UkQnJKTRscIpBmH5e7H3lvc8uccnHWvrztuPO9hxnaXlVW
QL39lzFXkKlBrh/yhI7u8rMCWKBeWjAWFA7F1PrZ/LjtdvGwF6QPh5ujeDLsCa6waGVUV3CBYtTA
/SWGpHSBGGVle8B8QePdP7g/R9b2overflDlnQVYpBgtQJCpLWpnX5bhCYWRFH8shQsyiHCACG+n
uPM64Q05j8gRvBfjW0q31BW7Shrc/EctzRswChyK6nPkkfaIgkx9fQnndwbjDWuUh/+ZvbXeEukG
UIZB816/X1vkmCsDGPAubf12YTYles7qIHPaF5z6W2a/2n1F4Z3DEAigC0CEB/v+3j4f1PZnB79M
lb1RwkfSjtC4PPtbk780ugrBsF5aV0z4yQ/tWNsrK5znm20A/EE+LYnHnUoJcpcouoMWHYB198TA
0QT9dwlgeF1EbUWNfg8L833Lq0c61gKIVmLkAO+3rpM1iaUK86Oh1vAnlJzg+jWqJ081Vvk8zBnp
ryzyqGK84ERxmMjnQ63QfTX/c2uNyrB2djXiJrMf0zzSzr9kgI3caJzMW+NVruiF5xCQ840eL0Ke
5XCCR3DJK73a0xBMxLbl8Fg3g5uSb6mtZ/FZttvv40ufWLwk5PXBZ0Q2Njvm4NC4w2wTSFeLTt1t
U/E7DPMIYfhPNANQ8kaB/m/JHxGBZ+5572z7SXfPPEp3+STaOozgKqOV/D+eP/19PSh7rY0uX6w9
ahGXfN8OXJ+PQfrd4LPn5Gbx2WBrt6tjePtHNj+eDwqj8llvF264U7jwlgm93+VOqMEFbwN0Dxm4
Y1rEiOH0iNO+iPnvZwlwYRPEUGwo+rm1VwOpLICaidn3A/npfLKNMIiZWg7318Wdn0LQwOicUzZP
P+PNdUXhS1SW+05zdWjqvcuj3dAXi7U/QuZ/lxiK0pn6Md19WHuYnZY6wlHPX8J7+cGcMvLxcpPe
biLgC78li2P5grQhsw5BwAKclRlQMKWydQjPq35zw+Wi40kObd/EEsXhxp2VKzKIaI5bkziW++nM
QkiRShAhn8WLWKBqlNJOEP1MTHQwTu7fTYv3xkzE1mAhC0h5ffnrD4Aze/tHAgEBDKCjhsX9p/Gh
5KoXhJZwYKMlqsqZ8uAFKiJd8cfba4MA6MC1LxbXf/6nZMYB3ISEsKGTPOQD2Gig4SdbRBvnMEtN
RZBC4/eqrabu79g3Hv+v+/Pfr/tNPKYk0iVMnIDKCRKBbrD5RyV/G5waRxto02aV6wZzExpvdQvc
IIGS8+kbos8m12f1ZtJ7rgfr2aZk+lKOxg3WqefttqMSjnp0FJkdGtT269Cmz3h5gHigGX68T1/h
l1NgcmlIWgI13pYwRBChTSaoBXkxg5Ywl9wp5k6bvkQ5HYpXP0prCjHuh58kCI2E2c34TSBJlHo3
dJU/TBSUMl0V8o93jaeg4u9j+ixYlYxddUqharvVoY9WsbWwHzk8Z4fU2UBK3e6uDHoKn2HIFeJN
SEE2Vs3NK9sCu3TTkm/jwF15cAUQ+wb5hvSnapP+2PUF7OiRrB8ucyQ6UMyhad8nwhjm29PL0EcU
QkWmHcq5hTTlv7Bxt+tomUgxhfJo1pIXMjlyBr2bpjj+is0CbAX8CEkQBpapS4UbBj38kxYLuOlO
9/YItnnY+2IwGeBYzPQ2/RPUjRd3SAzemyjvx8MyPIsR0+F1OUhrRxiXNHu8/r+M+WTM4AFfGEjy
49wBj/nkhFOZjZWhFF8iSpiB5LRHkhnp6J19Wt+ioLf4LMsFezhrOmL+d2trB85MAX5XRjNXNNVS
0WVQTyQtR131P9vNs1kqi4Xfpn1hwkERh57CmvughDQ6W8Pw3c30OIbJCyqD2roAyUbbtCkCeSSE
fL5Rf9OG5r8wpfTgRosh3+rLVbCBWaozWhHi7LEOTW5kT6ZUrwZw7sDw3FRgShD6DDDPVbH6DDpS
j+Y2fuMAV+SbG/FQ0aoAQslJSDX82xs4hOAVWI6ApfEkPJrdBPqqYiFZCpm0MuONX3nHIRDrBzLl
JKk4FSoypcJvWYnOuBsa1Ib0l+m4HrfLLK8kZDwG673/B+3A5RrZihQZ0bcclm5bCNvQC8hZ3n8L
2d+HMqHPXJlslB5r3tIGURuLgLfUUTW5U8yOLgZiLNbjdx9HqIl1CfxhnEnSn9OmtluY/8nDm27e
uAXz0GOrWop9BEQbUGThIJjrTGuRIzayR5BmOYiUSDq7jWxrSDsRe+UlKBcnG9FHcl18KyL7PeEt
00lSxXq39s0tLZuQ5Y2we0ae6mWdNmWJOmSH0LJ9CeS8FIAG1skgKC4+FAyg12yFWtaRvIwfriZv
joXrfHMhmLJdTkVzvHvG1PZcex+sqTC1FOffdQXaNnBIjTyyeywzVg5qjQKkUtT+NittMxixWMIH
s79C94tZH4rnPkG1eJ/UTN1sS3OL01k7ZP2/jldEbCrgqXWt5TZ7Xt+cSkzdgxRW/ZObZfNnwQ0N
ikIECulH2xHeppfYiZvdNCt8sVn+Pzrrf6MJ1CvRtQQoIzY58gxiZVBXyKA0+ggNHK9L5B60tpNW
iydokDams9ao8raU63xItHsfqI4mYsIPCiWugfRwfRzTzbaVHxrVSLaORDtZJaQ5UdNM2nlW93Ex
9f5RoeWqtNYz1PJzDxNCz2xc2856/d2Lwi+cXIK6H3XUMk5/Rtco1Mrh/Gv3PSVXzHfoBmyHhgn2
63FdJ/FxQAtSI6aoKAnJ7NpS87L0SDNmQADYbQhlg5VBp7jDWg+jwktINLWHck/9N325V7aTf3lK
QF0l86lwlby2CTzCE2LhoA4SInc6B2OodN5vbMq+mWa34N44LSxOPyS7vaivgMSId5q8Xl48Sx54
dtqdBgc9DAImiKEAgixUZXC0TjE9Aw7yY7I0+4G4a2GIs1ZmXjyeP8eZuJaBuq1u0GwDKZvSd3B/
025Xvs4FDwQzWd6gnPU9E3uAy1r8F7udO9/Y5INgmnZXoqKMc2zoFiOQBV7ES10Ofh5v1LKQop0S
C8UhxWD+gWP3l9wZzaOaSvjtKpCCZ00m4uzTLaiWyq2iHAAcD4ePhyr0rxSf1dc8B771bk6lYJsX
bs1A76c156bteioeB192copdWMdefwf7fDnAVXRWLLxGJzIOE7Si5IxwTnU0xHDenF4kKh2iw1Jg
1Z9iefnMaZ/bEKs+b5dWW660JZfsMy9EWF2L8EGxa5JL7qQO5+v6o6yeAYAmEl10nIn+1nURQR3o
J0rZm7WmIfwsz1LQb2R0qUBTB1AW8HlkQudyvF/+LhWsdQhUj4EFNgl7kmxsDnErPZcjdMzZG7eC
6w4fUpknE64oEHLokR5jmg/uXW+cXbVcjATX9xQrqCmwNZWdXTQkVuqLJiosBHAI5npc8ZTh28wl
dpuCc+8EGgG0CS1CPYG7U2xCPRYNYVKWvpzfQCitQV13utOaAOs0FuPQO+yU1Zsb7jREuLmkogmW
Lu5SASciCNIF8BGCsTQzNnkkxPSByH3cel3yirs5RvwJ41siPIw8g/o9reZYi8n1wzUslJMex9c1
3nQqQf0afeGENL0EdUGsxjK3zCxkG9oq5+utenVYUmt5HBCma1Cm7xPRIfKG2v1OQhKiGulzMR7s
aBOglpfb6YRz7CRc6W7FKh4S9eyX91hLvDHdoGr9dZTx9cokEsBw4/rEX4hAJpWFhAK1hGdYWLUd
H1trWWT2X598YmFWJgPN1wIwugeOdaj2cVhLxX6ATJx5N9eGiHTwMB2CXwX0J+pX2M1NJjWay0uG
Q7RmQCuTgE7ddoBNwDsazXsSlzBbbFBIdMO+GbqqlNjvC5Qtv0MKFSHbf+PE4cF9YEnDIth1636r
e2eEHDU4tCZGR/uL0UjkFcwqGoiV6F0HlPyEaiig6mx4wVFmUjFpcDTbeshFbsHNqukngm6VeFVx
rzLtGRc9a4hLSwW5+gfTwK0CFCpbg/yE/mY50EAaCY9C23XsZoCMvmccypSy6cQOcSnFA/LTOBqt
cYJdD2OeJwrjG4YrRN4+6A93o9O5wkRq2xEqOxflpxno2gKj5VCBiW1R3jaT/WW9PsxcpbhqgTyO
+VKVd0fTAG5y2tIobHO0NqEP3kYtVcD90Xc44W51KYLunioP5vvO9//XnGMxcMS1Hgevz3sdTDx/
urqwXlnh+seNsAqBj9JA2nRfGX9yvxT+quniZh9UQrWEDAzq+Q5Cie1vyg2Nv0M1O7RjHumZMyeA
LnsiODbKGt/slTmaVpKVT46lrHqrn8QpBopsOHs+yD+wuYx4f0PaJJyMxw0QSc3QqlTQHtXYf7c6
LtKUd/AEOY7SsYO5nYNWb0I5oeutSa5x4UaPOMVQuLFshnT0W0nlZXPt13O7yPz3mYMpzAxjp43g
CCOtp3Vo/bJP9gBP8qXtoJJNxNtDa1YcDA4IxSfZ2zBSUz3HJWlVpINJTRg1wlr10JEXdrGyRIYz
hTlMyfGFy0+Oc69J3ocn0VjFWf53IQNIhcMsFEARq1qNHmBfkyITokrAxX4p1y5X4WujmLwZB5XI
KOxQVvWmhhVedFWSkZrh6PIsDBI/SH9fB7u2Lqsz0ZDT5frl+J+O4MhF69EOVnGVcO1YtC9pYkR5
o8a8bEhEAI5k5THMlk2N1CyXe0bsujJPlB8QgRY6WIjBR/kYcCLymmmSKCj5DIEASlUL3JySrD/s
XpDtPAm33A8o/eyWPD9o5DdqMXbGs+H3Kno5Zc0L4ABxCYCL1YmlPEgvtagPjXeUHPJbdTymQ/8F
Ll6D1oywrmCPyOZ+SLSqesNz5dYg3mJsGbS2kFmcPuxBFVUEBqT3/NMxnJt3NJW5bkwARBpmepm+
u+OCTUxhO5yc+7cSCU5BUR65CPnltRQjgd6wivAgbm1T3SeCRQvfEzIJMitoZ94dHxoYP8+qqSxy
TVvsJGbiG+pXx3TBM65n4awVBkQvmZuoRnFYucNm/CqOz3gZzOjsKE5z4eqGGmt6DRLqHiK1MGG5
rMnpBzmbjsg6wqahTeU5MO55hN86rLvkxWV52yu/FUtR++sHCCKmmt7Cmqfub+qbSmc0ReoAG39J
Y7CAh7lVe93gmC3gCxLJyURxsEV8aWeELnXaxuhlNEdzGlIj5H/mm8r/EJBo2Zi5TXuJMQSAiAk0
QnvOe/PqarL3zmbKIVsdbwv+MspKuB7wRallVE6svbQcJ7ncxeAri1jScdWjF7+JW9di7QkqSmjQ
Fk7JEiInayi8PhfrB8SVkKujS0ftWDIQeCvn8bKsmGSi3fPBlik7+5loGD+Trixhz1Bb+tH4w3v4
ExQVWsT5qTkmAF0P48bQQ6Yvgd21swq590+re6Kti0KuRdrDX3kRjSUiIf/noIjQiUbxLYGu+6Yr
Dl/xkZxxAQJ2hZZD9GPUTyJwrjppcG4XyMXTxgBNLYSH+P9S//sPpk0LPD3m5sbBowasJUpKEEDH
U3dtejuj7RdCu0V0ITV3P7eXsxO47Cg90plICMdPgfKKvwp5y9vCHWtMI3+IpZQKb7mA1PREOMQF
xu4/PoSgwgnIxg3vNhF/S4sjczp8s54ornHw58FC8VsbpbmaZZTXRecs6M4kHXtpyNv0Pbjpyk9+
cicXoPXCJ28RPy5ayqhQ8xKlYu8qi8YkEs2/ORlUCWnTRJh03HW/b0UzWueyvRj/WwLlMhAtYZff
nD5ghIfR85u65XQWwvy96T+Cz/sqJ7z6XZTVUdN22s7Mh8fFQTxtBykcaBEL+TM/2yac6CkkksYW
AexGMFnMC3h5yL7Jj7sUAx6aDzmofWLV6YIsachUn3KbZJvaD//6aZKIkHxJY87kb6BXcWI1ECpn
1XORRir+VqZ6HWErwKu4p7fnaDBFzhzckoixT7jNg3ukgcDlYTzEsjL7nkKFhmUdgzhCbf29IyDY
GXVY5UdQ5oPI7RMmYC9KlXuRkLV7J8DW8GSpCd6+G0Hm9pG2GY41g1Pk0jqp4teNXvEwnO0US1iD
MC5ubKAjHo4o002CrZHH7fRTJerHH+ZPttaZu2G5mlihZ+3GI/YPb0JWLnAtSkBbDRt2uXpzTvBp
gHfRoCxjB82ddJ6hsbimKOtnQYIZaO917Vfy4Zg5LVAF2ECCKGdMuRrDiIHYUas5Vpxm8AZyvXHW
BlcKwGc/bJVDHfnj9Q4BlSCl8c/ti2SC+DM8spMT2I1zivhF6Sor/lKDBWfJ1FIOSWvik3ExX39K
U/9lye4Wn+6MfEb/H/RTR5C9s68FnH/MJA/SXnGDAip1vaNT7fEfjgevVCKG+287djDArKHVkgWl
JMte/G66/bKEsKAC7vYOdyvIP8nghIHZfe1yc6YdmRzE4H+cC2qy+lYsCFvtJUthn8H2qVzAzhRx
3coHzKnPwTJNgO6PufoySwoi63SfA5mSViKduy1h3i7UOCaO2RmtsFfCXLEQ41V5uLkdIBVEWTSO
QYIuJ70WM8hxvnEDRnoXh9oRLrIyUvlDfhzvwxp8+yHBibION6MiNO7gdk0AvFnV0QR5Fw41FQJA
mgcIesmGgU5DkUjDXdzFNSC84LrcTV75brjevSBsE0qtdbO7PViCkAWVjAGSzMEpSWZeqf6GoA+b
ZnnXzrQO7Rh/7bV0e85MlFxqXo8z/fGymx2pq7aCXdUwI2cyUOtdmJcL+rBUDvIsOMtwfWxUUEj4
ncksG+EAJEA8X+iybGB0fC+sKZ+YKV/VM8wHidR1vtvJovwTpqERE5MPP37qbVvOEWpvTMxqZA9L
vXhWlv5zPz08BB0aVUQgrH4FjkBMpzaHP6+jeB7/fAeuIF/uaIT5baWmjuRxMPFfb3SBdo7xDfAd
Aj39br8Xx7EvhF5OzMP/+Cs8Pd1V+FcHhiIx2D/fm5uuZYmRHqK9jo5vtUdYDc3ZKSAk0iQIJotV
f6HIU82yizSxa3WIiWj074LTdV7amYMFNIjzjQ1HyyFYy2NzQruJURPYZoeFSjZL930WAP3UJ9Sb
9Fw4c4OCqND1nf5cikf7S7dJP16copUQKXsyoWst0fIxQIn11tjkraJ+tADcF4Lr3FvBG0okMfaT
U5fnDXVfLid/RzGgXuMiMH6g1IietxVmwTDDflzAwOjEDKCamS53K99AbhzDvrIdlVxKF/y7+A8h
H0iSEPi0VjRgFmunUHY24obVFafgWEnrC6y+zUrQ8jYoKH1h9LU4Er+jO9L201Dk/B8aEhbpL/DO
MRqOuCEUlJz9XM5ae3rsBjXEbkgzkjXCEdMGQ33GnyDrNQV6rzR0/9Dtr/H0i5fQhFVAO7tgJbmk
+qg+PFrVAmNphVFwU0SJcQ2ac1zacv6Sq1KqRXO2hdhJuxxkgiPKEqKM1HH7dcaZSPuCUhXkqIig
dhVaUIr6Wjq7ktxLfaFN7PRIYfFnTwA+f8PZsswEDI1jXnMAe6UHsRHYgLHdNuvNamVY7/MLd9wH
qs9eoQvgOJ3W/NWZVuOjv/7UiDYKBvCkTAD+19gXsgcyDfPIOBeCpC99ssksdFkRNdgl/RE59kJt
m+b/uNbPPrq8nl/6wAOCbRtbJIV/4liBIK7AsvSOFHWiHESlc2R7zr9XoTfA9ntqER8cUS/okmr+
Eha9hSs2n8n1gpWMnxldYEfxji3Aja7PFj7FvHbXqjDKYMkE9dsL02f25i5ebHAPGaPuL2XCAIde
n/dhomDcLvvPzLRtOpFvh1xpj/3e/jMRZISYMCfgI1TVyu5DJeWc/Y6TLbwNO+CaZZEAgYw/CD7T
L1Rp/erFWzrvT/oGH4ijcyWa1UlcgrFURr+vbhaPDMv4vBKeNghykrBPV1k7JK4yAAdiWfWh/Q+j
ak4DORkXvQAO6AKbC62v2flrK9eMOhHXIsYRlbSx3x448QZlibtYKI3XbdKUNwcl1PEtcF08vXFE
1qG0L5PYPH+S3Q3fbru6oshn+CY43ms9EZF68K8mygYniWcAgUCSBye4Pg2T6zWiPAGPU0ZHbBb7
gbCWTbr77Se2lm9OSaLsjQC3cmMWeJA/pfzvFq3OaoINsFqzwzaKzwWBWLYp/rfOfxPS6k80c6jW
G1RmY7kFVZzq2ASkeMiWgM40FfiD8JPY5HLY27B5VPjHUBZ0D6U3ozIyQWj2fBfV3TroYmgdNEE8
nxlu8vAf6U79mthOrbVFvNyZhawj8CVnqeYHIx2yZqyAAymGWSkPP1J9vphYdr6jsuO6tY37YG5p
K0r5DFkHKWrUGvHFgi3kTddv0G80PMIo0giP1QEab5Skt+miHULrtLvmsMS9plXsPov7+sedD9lw
7neqrKRAvxrQLPt5Tziemz4kJzgAWVDf6g3Y4uuhXfMB9WgUfxUg0L0xpsz2xLy4cg7aScthyXwJ
F6JaBmRUPzp2c1tpLNtExRsXmfiky1Rs9Vjt76C6ie8F/T1/WFDRWwt8MfNBacQIp/PNLuP6LZT1
+uLus5jf8+M5Xd8csKT/AsPUHACIxQOWXS0cf99XdjjJqhzwtQBqCw4ItySHp5WmVInSgwy+JWGL
7qS08STF55tptoaXv3JXOAR371lFpCfwSBNCn5GVFY9wsepfqgX/3CZqD11dhiqG3zIYEaJwtSIm
5z9szviWzfsJN6c2vux9oNcgSIXIBit1R/MaMwZoj31XdfueSuhkLTM63I+AOd/cGyMl71NDu6le
8F+lQMFdDezlvg0Uv9nFxVlxGVtYpd5SmZzIEqwcNOkr9GWhaUrcu5NJo6ndpMDAmEBZsWkadBfE
bDCnvJXppgA8ufG8RBo1QarS9p3JZRQFruRSLxzfpgXizWqRuBAOlHUXtpKNQGqVAF1OKf/GZQRx
LdYNbp3vxcLIagdUXHy16F0tNxjRVqrflqbydI9T4iCl7u2XWknjEXVbcvdUZ1xGIDW8WzX2K2u7
TZv9fg0X0GSe3UlEXsJspY5tVbOuujJ2UAgJlTz3bv1P5wqEaevinnOWYMbJukN0glid4nnjvrKd
yDZbMNMYt5z4M/FufcOJZ1wH6lEuVUsWLzYdN5rdPS7QnR2E+qhFYes5MmOJJ1Uwl3UxHg8g1yzO
FpTI7+FyiTL/7L0impTJZ+kGDRPLy0136P2Vy3qwIXPjX1kTnYndrcgiI4Oyqm84BhDiG/iumcRJ
4a865Hzw3+XplCNlQ/XSQTuUCKbALy7Ay70YPZqZXHwJwBJvtFprwIkAgTqZ0+mxFZR9BEcblmST
td2AtG7ZRCveNd8sqUUavJ9h7Ksi7Avqowj7Mjv1DSyyhYxZ83fH5+3CF7cXrUjkvwxNJG+yXgpG
rb5Avo3uMCG/EK5M+r/pFwuO9mnBMTpbB6ZLrnTTp+BYUTUWHcnz4q8aUY/m1LLUM5KzcxOIvlT6
wdJqLObIA7gY/0cUjrOSDNpd3if7fqw439amPskyzYh4GTD04fB/Ws1s0kW2Q3Z/rga+x7HTgEPI
sZzUDI2SkoGe5YOXsSTeZV4res6sgh1Cr4ZDaWWJ5F7XDKK/vgVMOxI9OcOXwbAywFxvb1EjA20a
edA9vB7nr9Yl8ErHNuaEaZEyAsVx8M9EDSL1vyC13cXej2alE8mFKXgjFsitF3V7MnVQRBynwDaV
MyleYuIVVY6RlLhEHthbDgGblfWQkKGFnj+NVJI2WD+3lVh3AFj9lm8Z2n0O/Om8V4fFgglhsZ2L
Q3JMt7ekXh1pnCOBr0GjzPh9W5rssNebhY1mE/jp2CFVv7U+UVfifNHhzCXoEAmsEnFBrh9iaHcb
mYdXUlQg/YDFfmrna4Zc+/Ui0Mz1zmAl/+Ro5nUScJSYdWT83iGdBm0eTFFfaPfmHjJSQR/9ToUO
rH/Ps+9ps3qJkKOaYKxgoSXHE2r0KJU9oqdZY9UcLsYxYnavT+Hp6qbZnjh2jMXodFdA19VGU2Vg
ZagG/hvzpgYq4+OuOhYNkhGi0Im772myIMx8mtpR0JIdDb39pU+52wdk3YCKtfJtSzgrkiJ1qE0v
QHHsBZQGhDoqeeb3MgINbre7S49xegY+AdRNqFrFjwb9T59JReCPBQWnzxQ4Qbpie944xAXKxQ//
nOqN+gz3vbZfBKTpSZYYacp+qJzbqzslhBBpxQk4fLBMzpzjhqB1dwWLfRr/rGek9Um0M7wvRlgR
M15nsnsPkt7nv4A1H86V6pDUL+zgQ0OnndLQHzFvwg3K/b2jga8Newd30a+8NMg7ocbk+dA9XVrj
HZyHt271qrfD8bqlqUyJLrauF3CVRurDFsQTYG91jCtI7ljp1YP+SRu1jq6hSme1V5yBK32fRwHB
ziC2id0EBCI3aHYGdwsfjekVT1wSdSsKz/lqA6vBh+EAh3XB6D246UN+eA98nCTFMgm2Dj7rMmd6
YqPOI5YO5VwZVvbo2jJkEJvxGMfP5ZDkHBYEMHF/LqYggHs0lv5ooP+Br8CDKLU6vlqI/tpJ09IQ
yI7Mks5+MITLcdf9dIshqZEzkmPcpOMmlWsjFwtnBqHocUXf23ir5fXoJfrK1WdUmMjb1L6PQOzm
TmD8TNZ2mcPQBGj40Opt55YxXTNNphAJhf0A0aRih4m/+DuSTsunr5346FEY+mqd6kORTsaZ9VV9
Uotowv4HTikWf1VS9CXpAhHrGTnPou9T1Ws2Rtk9Uai1f4OGG/zthOd4lzihtark674Rmx7sbflG
Aeli/uY9QaaoDhZFO77FkGXEzWLmmuWfLYNTlfe/1d24ZhallVBhdpZO27tBQYl37SzZZ3imYFkk
a1OqS/gCyakw/mwL42b0jpYxB3i9+obhZI0Ho59yfwMouLmiZnFUZG+Q3PH6SGcX7kFVKPa6QFKK
Ok7KDC4gMaZAgNyWJUtHwbkDhbeGPCRCuao1G1jPmE3eqxRhAPDA5nJvtfJErOplRG5g+v+IoMKf
HO9VdERfzDfqkFIVDCC99y3U+9yrvAt5JOdEXBV16kHnjxvc/zn2xHfk/DrqNt1oM2EK9c82jMY+
F81m4vQmef63tgT+awFghtOolbQ7Ma5jqnMveMlfDLCu8c+kbOkSJrRxa0LaRQDtgzpr2/dLcVoy
/9pXghVD1FMU+89vMwlbmPtpG9Vc4+HW1NZV6qwCrfo1FVeHrkgC6wHVNR8c3/27A2YARHmNZje8
LJ+hcMzBziRM5rJvOg8EEWpua0enG3C+vU1qYJo5T5/HocxpgITxhRL//1DfGkyr0OVcy63arbQc
WzjtMZwg2mq1MwMiCwzMKCJMZOwIior6a4zICTqX3hIq4y9/56LsjAhcpQ5vlBydbvvDZfZq0uEF
tBeGwCgfQ1mEr9tT3dRHMQoBjwyiMoqhu/CCt3vZLeNhCXULnGcWF83FUztM9HXZaFmBS8frdFD7
YzUwcqhHNBsGR3JN3NMq3sfdk/BlF8iGPZ0ioEFbJ35QUMtUnsChMBbjf2xdiHuobHsNtuin56sZ
9F/Fpyozkh8G3Pxy9uVR81OAPCZBhozoKhj9utbFfVs4RftEuy4BkHbodvL8p2wwKgQAxCdJA+CQ
ArDM0fDrrLyNl4asuDVxkfhPvtsmHGZX7SMNaCLW6QCiaswMyNOsfMMHVyCkqtsCJ8WzBxp4UhbR
JuIJJZrelLuDEMRwJrZ6Dv4Gf93piESQ1dYm5ax8HJ/EGyD8P74KoS4crAe4lBckTmCmJHGVQkBB
q0TkC6jKun+qx/R32cE8eMpdkECr9czPIJxMAIdiateikjjiA0IuorbtrHiJR7A0dSJXnJp3wZnv
sRARiukrvJcch+b/3WN4iFlf4tLNxWCYyzNiqXLlRqz/oVAwPb2Fkt23qquM55c//pQm9w6F5eI5
hWdPS5KDc8+KOk/AOTgPvyBbi1VHKKez/Ti46qvm9e1aoQtFKhBlcL/OLFO33CVOJ8ceMWgQpz3h
IoVwebLAfimy8prkLOlWrONPnc8fM+yjmr1BARcEpyuQDNOla7PoaN8EiA/uWDFPghEr9jsQF4fJ
cwOLUNtDQWKVr6Kmtoje7jF1PZa2j4ue4blr2qGZnNs/WmjP2+gAJTZBvGYOkooAcDD6dZ/Y1kUy
5APz5c6OHwMA5scAw4ChQGQUJPDRiusNY/USnvRmBmQNCbdT+W35jDKLnfoiEGGUAEiFq9YlPFeK
n8MXsyXnGbhnIDUBoova+Xg9Wi+s6tX0hyOk4y4jvczRLVIjf0Oil/ZrLE45gWLuKQV5GjhcX9mo
5XqZxtJ53z6gWqK03UwOUUtNXOI0Rsin5nln5dEGgw2DM8ZGvc8YJrUGjAFPV2sP/KIDj3wkfqMA
PvRmGTvN7d30drPL2v0h80MiClyfaWBFmO0IpnD7rr7ZVS97UDc9r4XkVJgSXLXUPRdspmOC3av+
7H1Fe88MsKRpKW4GhhG38VNjhxcbyY/H9u37Tby6ePSySjvrMUUQVwh1jPzF8rFQUtaDCBKS4UBF
lS83XePOw1RwKxQDygeA0QU7RmLiD1AZ7b7oJ7CLDcPk5gkvMDgxS+0rNz5h5Tqs4LRC7oFQeIJJ
fpJLDggwfjM3DfImd64myX4fV/PKqxuv2PZuXE7nsWSwPKwjqdeWEsksdK5VKfEubWMbyJmFS2H4
LmypCZMZXnWIpwM0x8xLYCmMUuLgf14HJc8Ucfw1DsnFe9yTm6EGBKdyLTmvEE9+q8BfUvqvK7CL
Bk6Xm8OhdUlrJx6fmiCRxZiPapSB9lllD2pokzWd0VjSKi373DOdFeXWasWxHnbGdlnAoMunIS/s
yiI8SgjdaxL/WWqHVcvNdOIOvX1PrIQHo3wLiTt3q6X8cZodR/K/hiGerPGVRxSSC0MDqk+Yduqy
/0xO0BX+njha9EeL7nm6Khz/11dTpyNSuDT0qz09mUUlDOQG/HivkfNvexT3iNHhP8wWFHTSzgpY
Epc3mMO3qCxg0SLJPLaZn4dk8L3Em+4GeJq6xwifFsMapQS55qVNO9lGNVeNLDVZK9KQbAglz9L2
/aIehU1elkBHHYGRuRpC35AZvM8CmhRz9qQXd3kkrA1fcIi4xA6HMSNdDb43RkOxaj4cvSJmKAuL
L9dK5UNdkXDK/Nc2mnWHv1nAbi14UrpMkKLA7Z6aBnMX0IOe3JQ7A05W7mlzmtn11lSib/xOp5zM
JWVBibEKk/cytVMrAy7ueF2QPawZtORAwJ1pNDJrSdfVKR42tJcQtcDQSY+RhcV17vWKj/wBu6dV
3anlcD8OXPWqBnDaQuc91r/Ymjf3aVWWtDs1xcXKUhNKixieYCeYanfBAYsc0nnTDTyMnJkFi6Ty
lAQh3OfMsWonyWyak2v4tKMH2cx1wGj3DZWCwlrR3SgFgiQhKZRz4GF67/R/fgSN0gYdS4fhm8qA
uhzxnNQ7LzyryMTKI7SEzIEqfQJbzpIgYEjztky4OszxIZSVbG7kB+BLczSm6AOPUPZ5O/PxBp0F
8QDBUgYqlzcs2E8WzVML8Oc4XXryRwlYYj9aKoDZWlQCwS3a1uoTeAvk8No9Od6CzF1r3v+dPPBq
oBPX3Yf4XasdcfuWMB3su+mLT/zkEaDDAC+I5WsO23dRtSQ6xaYhFwbijmAYwPEiVIPQ0kYb5ZI7
TmfNsMChVrqfYtVkAexZgNYZJ4Icu7TpEQ61b2/mNVZUV8aI++Hi8e/dBUllwgKicK4pkz0g5MBd
13ddOxNSFSNMYV8OszXENhImm+VbgFskzaHZYn/E3GOh4D8yBRRkKgaLGl5vt4JTUBbQBjbCbF+b
FJNvF5PxIjbTL018J8rcSF4ob+cU778SUUw2Zfe3p6ewEYwv0s9QsOSUg5Q9FZhx/u6CpuqR3YRr
todhXVty/aTpcHywp+Tu84pcRCjiDSp/zUvfSWqXI2j25Vgjn7h8aO2NORvT+UQiVg6PCVSie0JK
RbUR1ni4o/vC4aumi4p7Szilqto4qKb0wmLatlveiDN8XmU1HjqWCJp2UuBBgoDzoBiCWHhu1OE1
VPfErc3C6OOykStEbBIVPA+Ko/dPivvkBTDykXOhK/Hvavk1MmLgMDuAyxsOkKum72T7XHtAYrKC
uB9BXN222l3sgyRkc3I0jrGY6vPoK7HxX9QMZ+HqoqwYqIT2m5Vu5E4leJ7d/h4Q6Ewut1FnBKbA
I8/9wbQMSK/XB0YIOk6WNtRX4ScUPJnvIyeU3h/+TBJPr1Zi5LonRPdzHS38GRDjTTtEsUoEc+7C
R8Cvpanr2bm8TnCxO/pmLUK1583e+jsy1MfwCYfLjV2txPaNhkCmQnalcqTg5/nMr6SJcN4o7Oo2
81CdWAGTTdpBt81FWhM0mdXbZWGOX0TsCJpLecSXJ5jsq4ayWLWlX6blGuwcfbpm1oxp4yC2dkns
e2kpvewaCgY9qnpR9L9COwUEYsZu4Y3dCV0sKOoFeT2R3yIiwTROiNoyspGTGzFA4b5Imnl9unfO
69Ug4E3cVxV2lYhWF0O98fZ5/d+MqW0blelu8Is4ayGiUMRuZqhfMLg78u3nsrJoJY7BqXS6ODbs
ClAPqdum8D+G8DAE4nzwbwnLeOFohcICTjYQiU5MhLqgu5xtfkvlTTvnQZDAE2+oHKIqjt+tol1b
hD/nhn2wcypZA2iO++GNkATxE71tjUdz+xRl+wNIdgQMLoXbnG+fkoA0NBrOkFbG/7a4HOYHr1du
iZy/JSL7E1PklFdQevXOilAYkrciwwnzI+nMNak+E92gxYWqwdmPux0r7/ZaBcdCMs1Ja7MB+jqd
PhzGhE2kP/ihf8HDnST0WFQhmrzHlc7MwmaH8rSfT59EPuX1PmAjI+gig8WvES6+bV0tAKGSFpEG
6k3piIPTqseP63BllfKlKvXREtZIjGkqJaZXCijDzxkNPWrsAqGPbcHvgBcK/C51V9TFj2+CNlJn
yIcd4yAJilqf4ZL9MqBi8OfUVGKEAT3oYvMZ8n8VyuPnGJDaxUfzJYeOPlvIyZYu3hIqSlexlP4T
b3o2jllFhxcUWKfaqDg2ZgF0w9PL5NrP6kn+1a/yvqQn4TstuHy5pZLmFSQqJDk4zAjQb0HzgK/U
JLeOyHGBNVIoz6W0URo7+7P2W+G0CVnR2q3GUeW5gkmGWZN+Dd5Skgz/oRn7dIPs04I4w1qPUmc5
LQJ8L8WtTi8FOdivL3H2I15UsgYVBjge+WlotGpd5Phlc26vcSAiXnY1qmaWI/CvoYdODFYi0Kt5
lHMT/J6mmNSkM4TYEFR/ldgjdKaHun62kmnmLsncGd1/cVWicgjIJ7v6E7iQNhOJ1R2D2HAyc58G
xHNTLinqA+7Hx2j25MRIPaxOQG2v9d7iGOf2f+4h+sjtvhWcNLMTetUH/LBSO8ZR76IynVzgSpeb
x0jKgxklD8Nc6369fcAgMCYm7gwWFNvnfrElnARSmphmfMTACYu5TVINmZJpeDBRD42tz2mEJAAF
BjwNOyixkjAEez+4LsiFo3BF08i9dnBhlAw4tqc2hH+9aJlIGLQy5oe0CpZyyQd1BTvz0l16uEwm
FO91a3SC8iUVsnn3tDFzm5NN3CdVxZqKEur0BkVk+z/DXpNIVWQk7K38ig64fytqsye676kC97pd
9jRcYELefE0mT6YEo08stzPQm9c526EVoZHS76jE7AKIInjzmoSxEdynzycn/JusahF07oMHfSre
bybV4iKKZJ/rQahQAxulwmI1nnC0WflSplhvzgfLn7uwvREz8zg0RWV0ZUYeuIlyIXEVWMRyt28I
PftCJeWCoeZsS46BeRXbQxoLob9Y4lpgPQSeW31gXGlv31ApAVGO5eTIyIZDE0L21mSa4iKtEPsT
SWv3NR5F9uLlcwP+7JA2AjB9mBns5yL8RvohoVEpeouzOq4N6qnc4DcNXM7nk3UyqOELeh0qZhqc
6+ZfhL/mmUzpiJi4DJNCX0FbbGBEFISeP5Hpza1en+yaFGf1UL3gQaN24Mw47icABouFgbJLWezk
7hj7TtSGvjjn5XbbjG5u9naz0PL5RVaeZUc2UUX0eFdSXgutf3HcYxRM24uMuG0Qs8iE7HfLv8Cp
6AKRA9u649t462EBpPY6KhTw0PKnN9GDsMXFLRiyGWiwmLLb3vED9jk9LzdOEiHwvRmHLI7YLEsw
uY3D701rc/PYXGj4QCz2kMhF9xPP14V5fJstLXFOFL0++NgWe+p2ZLaVBqD70DPMR+klJdeQXI9j
MmWgxUSYWPPJ2mCkVu7BsHUokPHG+TwwevdNGPEgVwZcldEp2fMdsbNDeNe7i0Zq42ZphUn53PPn
bGy/vpxlN2scGP6zNN/93YERGHQXGZ04jxhkPkHwaqSBgkEIybf0O28KW7NZkuTSiejr9lhjyHgM
MtyJkM0m8+7Jz3/+capB3DJw8uZKbB/N1iJcr5MHzCQ0hBQEMRXMz3C65mKgudXZu1uhO/4WrQyy
CPfl/SPmvL3Uz1k5Z77ghueEmJYF03OMxir7ZUFQm7k9YDxYjURhtl1S4B/+NA1e+wGNy119P2bV
tHpH+Ud5jyuZdr3Z6Zyd3C0V50wP6IKWObfQgCe8T6AUQbOxD6TwAV+agvdirf5kkLxbzvuVWD6y
AHudKS5chhP78o19gMYkodMRtVAOMPIuVkQeeL+N+WM0lIDc6++Ath0TP2+6URIap7e6Tuo2DgyS
+2zr0CNEWznVq6VIDpBvYFwaNGt9J/SG2d6KX5Jq4NDV5owjU2n7LsLJw6OyDYJ4QK3g20X3kdpl
mlt16mhWOQnuyinakrsqwm0vxfHCStVo+27Kxzm8KIiOxhFBsXfmy/ybiwh0UWPwJEQfEAgzw0bx
DLbvz4RhyY78KhVxz8RVKDP3FwG3uooaLmQqgQG2QlQdCeNqnPgf+1pdShImjjE4Pqr05eA1/SRe
c0VM5ujGqeCxGqFYPXA8bD57NZdfKeBbK4dDsXBGESPpirbxr+/SQtZ88GkPkHq22F/EshJWe2GX
Unqlx6lZLDnEcZCoUeIabbeJYx1ZDGUnENJSHX7a+IE2Et2j/e14OUjgz1f9qsvAWtMRXiTTOVd8
v6Dv+kXP40NWxyJdLPHhA7GIxX07G7QQ5xlh0BDVEX6xqShdcjKZIFxvpKhKebwknl2PgXxzTyh/
2quMckcwXD7CxiyMOoDk3RZYUDYJqMCmOfaWLasNHWN4ZnQV/cM/9DfEq8v0LTwbwLpy79lZLhNv
R/ZlJP+CL/sM/i8uYexZJI/YxYc7DMJbfWhpY2Sm+HMroHngkPMFMrad1FHM1mWNIoOp3Cr/E95M
P1QRv/LLfUFIvulU5jUWPHwnrhHSDyRJfw12zreszjbDggkJDpFQ2ip82Y46OJe1tXTCGzhrmsyL
NHicC3QY1l1+oC9jCC77dCzWPtV8yub4yQOCSXToJqc0VdhhX+8wYa7Fgsfv4szQuqC792MH4BEu
q/sA5u6aT0PcfXNA323W+L+c+YY5GUbcxNIfWEQQ4tbhyZDGNdf8EFuO1ZiF2yI2I4ZrgtESRyB7
+uFgmFTpb/YPwXAMUvYnS3uwd0xiOTNueFZLTvbFmEcTtPqlrquYpf3cgD5S0IeAPOKhmrNUDzLD
hGa7axFrz0HEQWu1AlHiDQS8/ClTKANfrVt6IVSPm6MYGRUMFottOouZCLkbP1TRi0NvSLv2pZlY
Phdd3PSMCDLV2eN6YAPCQZbEn372zFwdoHwEHmwmyaXEFmT5SzRNLhA9IhmIpCchpbCao3bNY1oh
WEFQSW6s9cQ8j+0znY2lOEbydZBVJWn0yHPxCy64QLHVuRcyHesehlbGEFcL0S59qjPM/qlkSibf
8W9TIJsvna+WAdbnOcH39IYL576by4sGMrmPfsUS7lppcbAOCemKBz7wwgt/15TSdKcCmYgIxh2J
nJVPXwrRCgjGWCRzrJGhwb8OHqfyg4utmG/khUGnb+rSQFAaupXNlKIMf3DJZijHA1PWYKe74m53
5wdp+kWM21ACfxfHB3jCMdDAOy7y258s8qv5QhnGkegUcqM+cnh1fg/0Vm88xXfFqKIUaURmKpGt
NO3GZGbUIb0M1Tcxt5HyfkcxmowUlOc6mzfFPAgB/uSbKo5bry0QBxzo1LuqS5llpqvlByXPZySL
6LzLEHfwFH3maBdtE1yJsQH8OeewvVvHa5EZdIcEaeByq0FW+RjJXCZwmGbgQVnteNLC1i52kD3Z
p5VnvymlOfyU3H4Zj49J3aQMJnDaKvdTM5lWWK4n1ZhbrpUQsJ8Ta1XWeNX4rlLHTrnMmt+wgmN/
koBRHEjCIk/1Z078H99+oDUcmbK9orjYueYw13MnG1CtRHNdCSnR3inbgYCZwwoKqxEbKtebB0w0
tzQNJ2hyypTR0CSICRYRvkN9l7wqhB71/xB10ikw+IQnZlDoCMtGcYLEh5ju3NQT3P1GS/wN50X3
ZMNLA3DG0aMtgO89kQyRRIW/Eiqyag0tGwXBP+1eRNZJRrkIa1zWqVXhkC0z5GSBiwSzsvzYm5OI
MucW84PE2ubIZ8W90XAUQZpID3W00n93tKn0sbrGDlF3IbjAfyCLGGnIW34szkRlpDHmHOIFYlGy
RYP70HeKvjBKGX5hMpQ+tbDwMyMF4hbO8rd/1tDQfv8jTDGK/hDUW9oIzqbuxcE55FkGY75BWelP
WZx4abIsv2qZ0GXLU9tgZgDraXWRx1RIclLZbhxLR+SZW0lLLVkEkP/GTdVRm727fydiG4XTNuAQ
O4+nAewEpugEcmeWa5gsqFjJNndcpCKj3a7XUgHfaEtc/TaGtM2azh3BiF+sVdFTca55b3mvEhnT
QwsHh7GPKEBvK6uWr1dRFMkfFVkv4j6tlEkixXyEf27hOs/aUKERtYZnzSDRNO/W2vnJIjELoJ6c
iS37rV8R5VnspdgAVSl6+CviFKe6SZje2G3VWVptrVM6oDXSySqFwIdpeasD9+T0CY15VbFvxEpf
ffkULfrF53HH47QtDtT5VvFtfcCD3seuKEzoCa/A6oo8cSoa5FLp8+r8+dm3kn4gLz4Hak2X4EeQ
gthadZ4l1RHOr67Pn0yVYCSETPJdW3lyEK8fw0w18HxRDruwZ5EdenbwDL6T8rRu+weBPCKe6vDD
k0flr+PIzrx3KpukIlvKrdTuUt/1ZXlvm18ppdKaRe7QoCOjp4hV7kFj3cT5/i9M319RwIeJl3dQ
ZfSxtE93VtYcs2N73+WwnhBHcdfNvw0ClxnNp56hGkHBrIGYPLvCvYopbcrc3dyxHAIIxPTcarTn
E5vigUTtA8mLl0Dz1JqNw0Sf151AuPPEMreeF+quYO8+aYRUMPLHPW4Z9oywq2xQEn6zlofPE19X
Er+eMsWNA6hrTPPUgK2ymQTEIiCWJDdgRoQD0MFGXBVf5ig0ho1lL9iILa9DB0UpK2n68ghb7Zy9
SN2miXTysB9O3R9U704XPJ2WsErZUwQeHmm8kMp2XRe1tn06H413mfsI5FVAjNGEQbdW0JUPhsbq
GdTbcGeybk9ckDYtpoGWVMM/33ZbmMRJI8GyBVpAfAUsRtqg5f15byJtRyFKAQ0h7pCSuhSOmg8M
l9GRSjysVobwUdoSzrvzcUY063sFEf5L4V0bfQWcpsWpX+QdIarzJc62KWK4vdebd596IaQiI0gp
fH92BdAjbx5+cVbMWcxkp8vpZnh7IW+GwJv/ilWBLJgYMwi1J4LmAzvBjuQ5MLMFmQFr71wTBH9R
LbkitrR6KXSpwut5aAooTc+nplwd/qNq8yLhe4+A4kwIBZ0CBjXGkorBPJF+Oa+CG6CG9eeqcsoE
VnkodV556dovshuMQr3NysYO26Vs3yQhAiXJ8TKuJZhjnG6F95/AHE+eMtwMhV0qLJnoJ/FKblN1
F9ss31DeMczj0Oz/Juc0qHqfbg4jDGgjAzShhYZMnNrA3PtSrWw4L2rOGEBPsNLgwfX93/uW3Gv9
u+8xbyF8fomuacX1SA1eO7mooFl2PSjcV2NopVOza67uxGAYJJ4qQ9TMrAJ8Lo9xiP7RfHPO3eRJ
OQSo/YC+bcKNX2uM2I1tRKSgAFzeoKdywNDVhKVff7vKCWaKvi1iiCVSClniU/lgkP8c/VZnd8OG
co4Q0pJ1BrY/HoJqZ9sz/S7l0UF+FrG/JVxJTsn04CMKxSrqGrQNRKqiJyiNYHLuRnF4QMsMX091
KgxrR8CnQzRt0IfHmiBt/hNWpj20mp15j8/Bdkce2Qt06cebrxjYEeYK+EzElrDr0DayikNjVUp8
T8RL4v59b7GqJbKTHMOGG2fET6Lnn8CBC39MMsNTCltBdQNiqmc8P1gPHiGXevb6Mszeewr0Z3p5
4ckLbPYJpV9uGf6y9GoLdmrTP1j5XBEWFR5tq8xBIMfhDD3JnLy0LG0hQS4JSYQK38mPMYLR2v7F
O6tDYS94A/h0o0IJHZhZjk6FSHwHjbyDFJTfdrDoiaRWt5GdjybHdDkXIC0IJ0E4dA6zcQkRx4Rp
SElf/FLL7r3TV81T2vjFCK1hxqREAIYnSYYLTbvxlMFqrQmy4cTb8vXYvmzhu0WM16gWxUHJiiMI
EVgu8lnsknzH+kvfAIbd/DJC2npvL+7itwMZBwx4l5UF+cETx9uc1IioCOtI5KZrwmokSSxjZr/N
jr3MFFQcZlSJTbGbhoZQqiG9zIh8qpV4E42VxL2Lyxac7GxVlaiNOlb03YD6+8tjneDrYgmAxRO5
FFTp9slQvej+Wp0JkQxoJCqcwBvKgAc/ZQvJ6wusu2BMrKPQfK0++CyyNNIj7osZ/rrxQuga9Axg
bl8xFsyXDZhv3w2m+9DyU9ioprMt5ow88eATDAMbD5mcZtHMmPysZltKNr21whJqhbUkzYuQdwur
RBYGenzZdkraMtLMo+O6s2+PsAZaEKo+lX2A0uqc7qgHrb0E6kOv9HZtQXVze9OJxaUh5eHqfWoi
qMRHL2UuCzb4rCIP8JmM2EokcYAQm2C7SLsnPtGvPcWkjhF5+lXu9cYyc9U4/e0FC9ZfseGkz4o/
OU2gn65/ZZwT9J0lsk/46wUCgoBY+Ra/WGZEICmf1oa8KE3VSm37uI+Mc9v5+30HI1J91eaT4k4O
Ocp+c2eKtEKhsJIcMNwzlk5bcUGSq1lhEaWYzjxCTRkBTA12HpeFidUdAAF1nPCZZE8ctprT5ZkC
QdJ9DadMZmharEWy2z7Vi1YKCUtbRL99tX5Dyv7O83llxYrXbLmvaB5/i+krYUhLsXv6ngTSpqtO
+53T1fsLkUzuhI48B1PuaMdZvAkHTGhQVMxuV1senvBsSEZyra2vUMdXIkNzW9slewwhajC2FZqq
HSc84ih/AHWxOQERfLsVWu/U0DVXogCM5U/l/T4CA16YnFyt8g4LgB8amSBpEBAXjUIHuy9gH868
KPwMSbZeb2sUn3o0mHvVPfV5jlEl828Nt/gdHmn5P8H0ynbAnLKCL98hl8iy3N/J3sWpqfCrFtXi
uNbhRZrvwmW+m0epScVMKodUZT4c0vvnL5AAIxYP7zZ46p3YiL35GBHDeteN0NvX4rdfCZJDu4tS
EHojCP3kfroZggwP0IwgLJBh8gDdL3dPp23/pW6T1qtf+2fZsshxZkwaK7Bcj6LPp1IsL/U5yc8t
NYmqag5lFGi8leF5rUhinr5g9WDrIcMXDtzvF3fw4ubQYWoXiXRfUpRTI+qo9WwSbF9mNq1PVEq9
G3qo0KenHImHi0r5o7/ACVGV5zxhcknXtfSTDqO2uXQjJwbLSInmqDwPooS4Qd8i1tS4aCclJzMg
lnr//eVQ2dr/H1xbOg5v4JkobZxhCeRc7Py9ONinRLn6dGraX1+8ssqgVGT1EPCvSKRvTGMSmJhu
ihkIrPZ32+9KUmOZJlGnRpe/26GB9y5aBGoZETH2jDUH99FCCbtAVncqDV5rcHspMIta8EceMAmn
HWwsdf9x8okFgkGtefvMD3MrOWr4zZE44i0oUQwRysQ55umvrHG6aVKRtssVIPoOC9UtccO56pVV
/YlpticylMLojI9m3tFQTgqMmexS6avl2b07hcWEkHEsR497ABa4p1YqOKlb6HF8Ze7hv04tpFSK
ABZNKXB/h/eQ3qtRxSdKJQb9tCn4b2ovh5H3FQAhdkRbOvzq3RpCUgjvDJf4lFvbnI+/LqZQHXvz
5JUhUW0EXJUXhNz74T7Fjirch4VkafDgbFeXB7KNICoDvDbKSR6GmpCgQlRca23fZYZhVjOpGwnR
myxQ1+9mJZkQz1WBEzIMs39LGBMmOAdaolwj8GQkUFJ7YBRA79wy0CXVJUseJJCgykcMKX3nXrrO
G7cZCQZeTnf+ZfRQMbBBXEyv4Zxl/DQtyQRQ1Cf95GJ3Siq5ptrD+kV+6lvY8SpvawsrVRbAApQz
k3ysQ2qwtRGpqnWQoEQAp9gwgHdCTN0T7E3ltCe3NWt+GNZT/iySO6jsKwn5yAkOlV71HkCx1A1w
2W0wEjbU0H6DquI6LIbAB1x2hSMNIpdElONrqF6NaEoLk2jujakYk5xkBR6PDdjQriiLXUULq7sc
04UvEubyVCGquG8rTuZ1jhtmKrav6g35nJVrrAQh76u/zZGeoFti40bb+1IiWUOycnHpn8FyNnnz
rLq/9gYn1KQ7NAzsQNkxQaosZ5RMTbAkn/WsZdygYmWvJWZxZETLbvn2PFyDt06cpS7PGnexMU79
hjXRwtTkKNFJlHf3K/jwGVM/uyeAl10ui/bSL73ix8LVPq2FeVvF5dX/DTQIhRtQxBZgd5XQG0MZ
TG9NkT4GuYxJLFCdF95B/+lCl9r8TKrmvrfjpB8/AwwRlP4pSQDDLUwsh6aczKi6lZgRGzDYyo8V
axzi7PUDPqvKZ1lClrEuAGdRqn++EWnUfCovaK1H5iECNWN86nU53+wZubrZsiKxw+FwZsUiRvVy
9J263Gr2M7QRUmKqICJwPx2NVljMex4qlZ/yEp9QxJNZLV/MnlWl0Ib7Av4LqmDNGRrkaae3WZYc
7JIxxEz9JLxwU8U3AVXny73XhUtfXD7Jl6mifgmh8A8FrR8xKAcdeeXGaj+ad8RACRLkJ/4ENwwm
ghA0VJQQBrGM1UjgXN1wJA4JfPUPNMhEY6qQeuH4GCMmntLK3V3cR0Lr++9w7ajAHesGZa0aEiN9
+5qwHmu6GYHDpIj6XpMpVu/37hnUzfCG3dhU4iU6utrL4QgvxcTO5Fjg+NRLnNXrTO0LzI2WqrcT
nm3Y/jedL70EEBmud3H8NEj65iEbD/j3xYClh4cM9LtaUqeorCJ0O6DNy47OxkyDQzCOT6pX93on
SJPQgS3mqoVp0T3Z5W3ykIns23rJ3/1FZ6dOt+s0NIygGei+hsrk5jJj3bKRlOIJQuUv9PS1ifWJ
G0QBlmbTYkRhCLR9CBNFDDOBD6dZyrmMPD2v5uq3uu+fEtkFdY++sqUcGdiNUdt9l/w00/blTqDl
rA7EcHdp2VoQlzo7C92sBHnlPw5zVQMN8L2ha2OhIKWnf8mMwkMf9PwbfzgL6TRsDDH9eYHHP1tZ
2tD+3hXaB2DfAFHLrmWXXy1l6CuIe+ynbiFtZUnHzHBlsrELxtLetgbL0UcAH0StZIW0f2mwOxTd
dqm5DiYz0zMHicROE5wnE7K9eGSG+SnKRgikCqOOueetuW2vZj+w30G2ZcSDnLP00nep6H2DY6x8
yCCZchSaDS4paNhKIiWOipQCc74G5Mrl9I1qbm3g72KA//3sNSa4ccnWy/QIj0J566SY8nw8/k7C
bbqCRQPw59tSJJrG5j8nEQ64cEszieRhwOFUz4GvBZonLrP6YMBzOgEbPkqDTgMdXYeYVNRI3UmH
gGWNinOAeCe7kZ2qD7u5LwsLHexFqhCOk902RgktoDUx9Q0+A44yilv/UbN9gnteFn2yYzNrio2E
RzjV2E+IG55JDmE7i8W0Ci0vvyDtaHi9Wnmhv6gAhrGuYGcElVBY1Yygo2bJi63WD4hWlkYIMhLH
+Re3UB0aiQsP8cOh64ucEAm+rfG+r3BQ9GK+RQFO8DtC3daxwsKx+bIttiLjoTxiJhJHTyKK8KI5
rWGldX7zWNSrlkEDe7GNRotxFdnByrk2OTVztVH/kYkP7iQ2pbQYqBCbqSCKUVB4EI++3k2NMzm9
kFkOKz1aZc9r6fb3qqzjRmUAiEWcJ7kxZ5CUiCbzzAeoDzB3Ykyy14N93263Jald0gAAjquSiXYl
W2FaQ7XCsy7ZxHo4ZaNom7FMYkqb3PWM//eOAa/TY6kQ7RgWbJwfy26U2nr7A30ehMFopzKcim5W
duaSc8IJ4dZ21ouJI3RmVQxhfN1QnQR9zrFn2Gb1jEiTWwBWn6S0KNhG0CeA7+ipvURlgnD7XptE
c64frQ3Vp4Vbpmemeu1Rq+FkXWGGPHZplEvJTuDxjBmsO9KOks1swnWWaGiL1lMq3lIT1lheZhZi
d6GxOVDeAcoSdKO03bd7Tpq/xZNj9Oke63zedcGAg+i4OgazQoOflb2anwh/+t84xC8E6v8F1RI9
o8swhbx4HT8PS05w5XiZyCDTJhgRjD5884Gd8y7dmfqShO00VDEXdBcnhkTsaCVEHgNtbPAI6xxs
+J4I9kjSbvMLNlmH2rbD0xauNxn+G2SPq387+h5rJgW8O+bJmO7mQtHPGeCWWow6l5E2ss5b6LvT
5Iaj37nDhI7zPF8kPMtuPynOShiJ/UoIU75X61c9mn6U76GLzNLSbpMZYRk0PncNa7Xj/wzVRa+n
xCGZeMxdgIyMHWoHeS019BsyYA5isvZLzaDWIPKmX+kn5ZXVMVKEKo7cn/Cr48e3OwbHugrMjxiC
gV51JsCzhobK0ZZDSVD6Vs8pPxXfQPGKgFUXoXB5ddme4uMnQhXUUl+noEd7uYf6wbUitzkEJhnl
T1KxRlMMJGjD3D27okp5B3SkikMFka1p4AkB/emVrQ2dyMFg2u5fjneM2hI6EpsMD0nV/xraELte
lKp5YvgKk8lEZpYLX0ffZi25EbVU7WAVZJMunLrCI/cLVk82h0/F/46DmXaQDVQq/Dmhxauw4jH+
rPtpGbuLIhfkpy8UIleXH2WKs1lEIog6DJZA3JQfbA3sq2DxOTs5CWmzaYpgRuc7I56ygIUVj1dr
a97+GIo4oVMBbxO2GXU+fJf5jdZZBNSWdcNDMXom/h71mfEcil+llcox1ZQZ4UmKkC0DJNQdn2gB
Pndj/jSxnIpug2RF0kLK+TMTto0Dqou/exJKsQy6WS9YJlRl12GZ5qFNxKftlo/rauYsa/9ZM63H
Xeulwc83NXxDnbHjI65zM0vnAUJUV7+rk1NZvmTL0ikbq3fM6G5HbxKpsV5qaWLvSGaVio6ukvu2
967md8fE618Zz+0NkEsRFnhl67KcNhiH8JeKusSMsVJMPw4un/+dGfzn+Vwvhs+l+VuNx+sbbsIr
Y+FODTSLB+kP7L3qcUB91+fUt8zovmwcmHBkmLv+liwq1BYAn8zeGbLhFDTZwOygVw6GBzkigy6A
2tFsb1psr+r1o4C0smD6kBFG72twiWhdElnjbt5gW6+lovHgHk6gLX8BnegJwb7otWzhOZUdGKC1
lU/iMDtL2fEXd8gcEgH96YONxlyc3fsX6H6XJHXTllJfPxo3jshpUDHjDAEnWs2yDuky6owBzB/u
xHvHQAiAoz+xM84Cr2gKu7PoXQhDizG9fgMXjghadmal8Gcg9cT6C/Q8BnLLt41IiYwrhDCfNAaL
XMmvyvmVU4YxeyDpZqvu4jFePS6/x9xzmOaHWAcWiEoSlll5YRLtAEAXcZ5W2zZY7kkktXy0UhSp
nidn2sMRHsEzhArKeasHfuBU4epvPzCaBZk7LVd2AWEnmB/kwkP+bsjjPYm7IY/6VjdgqqvYP1B0
RLK0qnHdUV03byRuFimSNHsQg4s+Mxaldlk2R/fcCvRf0ZUlChvmZlw04J3cJv7aJLyni0LdDHiQ
o+LY8FHiyID9urSqh8ucQSZ3sBKbn9bn+ieSazjOtfPuns7XMAYMyCHsZSk8hra0wfCQgBRgwq9F
OSmH0vBF49ZhpJe3JhVCsmOrxOIMNO3S0xSdAhcU02ome/peW01BhzUtc0GA68+Sycfi5sjbh5wS
HTdfEBobQU4JhaTsncJOHXTZuBowX6DaikzaIFHCklNeKVDi1pj7WpqOI0xwxR1IHLBrbB4uNTCo
4hPWajRhEBkhOr9mKOtmsZVIMMuV+3K9oLf5acoiD4G09Nnh5y/+7G5kLoJCMIOJzhOFrmke3Vp6
15dy+O4VfkUIWlYax59Z5H/2ColfC95aIVGnr1xzTG67bXOEHOoTywgXobtpeD+dD2VFrNCWtqXq
ULYciDB/O35kI93sv964KpPbVoOP66RooxFOgvxucOz/0sGTY3mP5ZGif0Xq75ashaS+ayFnVSoP
FG53x0Da9NdUljAuCQdgOJXXH9zWGkrpRa8/L/DnzylD7whasbuSP5gSZNe2rSKw6YVYtxWUHaMs
G1jZQ/PPwc27a2U0wcN/iq5wqVCyGNGGkCakMz46ys2LQMF8AIYXwsvy6+zTUDTYGCMOOop4P2lD
C9S1HlFD5PoDZtdknT6iZlw/XvZVXXTs6s28yTgE2OHBAAXBvl6TMdpzNy3xagtRUOtB7unOxJ3C
OCv7WerkOS9y7x1H/KNmEHOWvZCB9VsBffiggCN2pz5nbRo2lZg3E8Dvh9WeMqy5fWCZ+Vej8A0t
NaT0VUU4M8+bOuxr+kTKOX3AVW590yUD2OEf4O0ZRvSXpioZZy/KbJoZNdStNWRVbCiEm1YsUR2U
62IIGnfp2KOaC/9LTwbr7dWyxhLQi1bg/m0U99kBX1R76lVyuxuUuSqbluY5XZUW+QjHUwQQurcx
/mObBOHEEV4q59GL6F3ZAvo0qzbozmPo7zGA9WPIcyVQATywSiYvdAdzO4ck6e8BCJQEYN3nw0M4
8nPmm6Aaf0QMC8302FIDbmDC6egDRSq554sEKT8NKMuHC+hD6fj4JOECC7v1UBy+2ifgxHehZjpF
vfQf7qGk4GA70aKYaMcIp2R36OmKQWSwfR9LQYfjHi8f7K6jbChcz+mw8VkjZyyipJZanun6hwoM
ZKgsMkBpeKwYLeiJ6EElKxNw+rzcL1EI8+63TZmSJZrqIrBHA9jcSPEQmlm6WlCX4mXOtEZGC8Jw
1MmsxR/lEkRXYsUdVHyEsuwAHcKgZrCIfhmwVssAOklnHPK6qqCuojis59qZhlRAVApkESLf8caZ
uOMC8s3ws/NatoMSUYoQCAdxeyuk9YwzoQhk7I9zYURqL0GVcu7Y2YwB5GRiW5DjOxiYhvzZHbgt
o9Dp5ucQ13zwp8jrDLGsAiz3AXrCg2Ol75TBhycXvL0nQsFwI2lxEZvSREW/SSFHM0cpTgVZk7l/
JgtUS09t4WkSAetu09kgc/tWk0WpDb6/GBpYyOJknUEb3XaTx4DvPXlOGb8KSM1Hjr5nopuh0ykV
Sf0RuVWcbHu5ZmK42tECTdXWr7RWd7W2Ut1Z3HoKtfCcBJTP7+ERVHqVGnbHSiPFONdd/Z0givXg
CS7q6ITONQ/FBB5uWcTfXfosTUBxrfE5/Eq9K4lgv23ZqkzDiPK7PoW3cm/W1C2AEB4HntJh08uC
aAv3gCu5U+9Y/JquFYgvPmkTppxTAIxOri1Pd2OUpld+cKhlVwu2sT48itSr2UL9znubcZiLGTQ5
NCiNU/tS9UvkNnh4w7mfyR+/y+sC1W6lyFzKLKS2urtx/GVevJn9dmG+7iceaLQEGrUxctc2a5jA
32pvaZhOGZCDTRAAY6rQvnVkOX6u//3qOUYjI5TeaSHSO3Mu6UGvkes9TX2me/9szWb+OuIvtrQd
6IOS+fsrf7wg/0WE3CmtuJGfHDyAW/u6UEeYLdFyzu86AjHaxW/E82d1RVRPlITYhvzGVLmucVbB
czxo0K99Ajsqc/rHSHLjiI72LpfNUfj9anYg1ATsAltGkW2vy3Wib6gj82PtC3oCGruEtrHsIsy7
q3A6hF6MFPqkENPEy7ZPHiXAaEAV0WWVN2YznB7DRBam+A4E43enMU8CQzqmCWtUG1I5PVEGXqv5
UVca8SJqM67Fbtq1WMT5slsrrKAlBHTvM3pYzdFBVXzfw4XeomI9SJI7Yb4tK0tLyAe0GsUO9HPd
sAuXI4ctg7vFbnRdikkvuZoQF9QA6QZB9L+bLp7iZdnIgKnvH2UIyHhbp6/s2twaJYvUGG14fdlz
kgrbS5c9AlmAOaZUt3tQ5y6pn+WkhY5pBHT8+NQNY7T0O4LVlDPf6K9eTC2T+QqnZdvFKlD7iZpV
byUoiKNPpaPX9aiAwc9pHyINdMbvEO0RLr2F84J26tf67YQbEIdPIOl+kVO7HgU/1H5ji3oF2VhU
/oEgy1rlVPqlzwSFgmQ5Sfebaiyxe5jzYo9f8/f/GAwTzu+gLKmmQ8eMXUbH+w/H5bLEVsuWCYkK
S0xrz+R78ePOLCA1np0/qjpRoifHFjMO4bjgq8kMlBsqiWDWx4h0Fewtj6B9DvQPQtBSuq33uNuf
i8phbWin1b6upovxq4SAZxwua1nY6cKMXP4oUPY0yxC0JNOe9XYZ4R+qtaWxtcGRjcVQzsqoFc2U
5TPLfhnVTPbvJCCM7o3/8fljA//hQXCG5k3hYOFdA+l2Vz2CB1De+JAwzmyd2wi9iLjZgmHPO93T
oXoQxlIAlNicWLornERhiiKYuI9LOEZ1JxbXsioOxfQJd+Sh30ZOrwJkCXF3R2nGGgk2zeSOZ9U3
cGNsSgjuTUXLnPLxfSCSCOHe8wbiIbZFBh6ug3NS9nUeX5ox5Dm9meOn2ohOmMbxgRCQzlr/9ruk
6uPLVhPZtMSnwqGG9QdbUmcBc/3zjoyz+BJZjUuaahK0pk6W8g6BkFgD2ugiJamfEzbLj4F2AM0J
bTokaR1AQUiDp4/QzwsZuzNIfOpj1sjmPNWgeuhh/zq+PapiYaqjEFNCBk7VIeqPFpYP1nnCmxXt
vSE/Wi2SBowFu2hjxf37P4Sgd+sMvR3grlSdQ2de7TzU0XVxfWIWp9IoXJ7iY+s7LhCBExZJNJ/Q
qldaW5Xv6CtX3/gQLTaQ8XPq1elxgyBLhi4NBGg5yj/7JRKWdds5fAMWtE81THbq0HWjT/ULG1+n
7sYkwY+QGeCntlLzeHYQKCNOTWQktDeRA7E7xmmFZ25GPLurvyd62dCsnwhhgplYQUYjisZQEnCu
RvJk0Fr8UY72j3a2vpFIOyeHVAPeZwR/8rLLW+QjPGZpP1RE2+dQn9m+So7cyAoR/WmUUFaZ4txw
PNMsfLvBD1ptcSe8Pwj10+3ttP3z1JIIQpywFcvmp178RCGSBlHeIDh/B5s/LKY9pB8N68QbL7kT
02SM9qZEaqLWdrm9WzIxRaFbX3HE2pbctxgSslnWSmOhsQ0rOMP3pLIS/XNGd3QmEncBIcFZz3nx
gyVfWSXv8OsaKP1dhfOObyFDihjL/otqA/F1Z+/69bXlRX+Y3nvLl+6rEe3dnAjDu/hv9ou68OJp
CfLHQ/z/4bEwQDpYtHztCLzLl+JFP2+Wlqva9GgBjKFaGG8S3rVshrmB3Ry1BEnTqh5M8D9zsTpr
14sfpj6hDNizPiQev0jjcFrZAYkH7/hd/BzgTYL88npiNI8CLj0hW5xw55eZ38a2t0UbUlLnBYo6
kToC5ECW+081XcXr+iv16ukeMhiV3nX0/B80T1AavenulYqfcs0+rWiTY5vt6YGLEF9OY7dVV98/
AggdOkU3CnKRBLoS3YVxAmWGZi5/cqiaCJHLjjhI3OYOuAmJue6ex/MkDyTfIE533c6jGhXw71DK
wJELmUYzo7N2ssYn/Tj6JMz900NU9dg+ksEvIZ+0+8lxDxNcKZVK8fvSI1BIBqlrWEu91C91Qt4k
MjQR033ISm7mv0T8zjUqSgJ0I3WvPAkfMcEUHFGnK2oeUH4N+sTdwx18ApomxI0H5jmffThfgqVq
AAr/J5+m2bCpbmL/I3MJAR4crJH4lazR6eeepm3+ZVLxNY6e4Dg4spZTYcksf9GWPa9qV4BKYxFI
uZR7hL4FdT0T6OSnBXySEmJDDeyhok2+Ct/FK/m0H/UdpS0pBc9A9YY2CswBt9QWPnPFMeqREqpJ
78lE0EI0F2U3nhDTcdgO78icnk8muyANrC8CIZBKGxY3T3/InMEKLHoi6eSQMtAIAEE1RYpYUc+y
XCf6pAAHpnjpQuRMw3I3iYA9UthmRhZ0A0jh2DvbZlzC8zbkfK44wz6r9506DPY3YdOQJdHpKntp
o9BD/id44kHOBOBknCyY0GjDY4u7GjwiFJXMOKniviKPWgv4m5E/vEtGwacB4AwmwcI7ixo/22hQ
xDlXOoj4RNGxh4w1TUQPCbNtMsNYj3XYhTJW8M4zs9S/kNHK1rTsW6G3NtDX2UqPulAS1cWqNFW4
SUXD1sisOPO3bMGzuH3LYeyFFzbTFpwV7NMaF4IyGyOWpOUrWBBnGla5u9AanzHMQC985HO6TGy/
70agw8D87XMrwO7x44+wI6KKFyNaU8GLpJVgyUZR4t3RRmnBawYIZN221NzvEXNOvU9mL1+QXRQ2
2WGdXq0h4lLr6MDN+KtbfNZa5h/q0M9OqYlbyhoDVL9At869n7YQewNkMow5I6EaQ9sCm0jJ04i9
IKajxqnCeR/FCqtuDjZjShZsitE/gPhPXx+UhONGYIYGp0ePAPLXT9ICAyb0/MHWxO9VUcp95YFa
jlrL5GTdQ7UlujGoSkhPnjNKrMx90UubsH8fQWfUy8cpStUgh8lLs/GcsS8XsbvQIJ+OCN5MfP2o
5Nxjri2Zinss2plWHK5pewa+dMjH6Y0Uk61R2R6vchneDyRdDWUhmkoLL+TDU+pK4PuPLqYNXeXU
jrFBz4BMpaaLwvRCUr6v5lffNsTmvjxOGK0o9GBO/RLzJBOUyZkX0D4WzThkSVx+S8Lb01ZDNaNK
rDWpPciUT5TiaLX5klD9AJMwEwgByKf9SZZjR4ZxvgoNSSdZ2D+m/WTNmQJiwmgcRVgdiGNcVfKV
mNrkbcDjzR/tBDZqSmrQORU3ZRp2G38DM8bFHIcNoAsydnSXn8Km0L1ZyXLSEsmnAht+9/lrFjNm
RwbR8uJ9pAL+yJd8crFMpEPHCytYtH0gJloVVJKfvnvTODvZu0h1jrESNhPgi58e3fA5WYPsEKmY
jXeMc29EedHjnMinhddd8rP0Z624zgnxcjrJ/tb1vKhLEaTaa5rbdvIz8FyxAgaLpR6tpiSy2YQO
W6zS1KTWW0zx1cFvQc3sXK2qVEIFsqSVArT2Ct8OcdcVxhGlTh6E5iHYJgp50AaW2Dy6PBHgU0pR
+MUR8Rh8grq/2tCIca0yfGsLr2moLslXcr07hlDCXUGsJ9E/HqBNkSzKe8IgrF45Om5rP/VkrB3k
lSgcTQABiWI4AzkWg/2t743gmL2mnVBEFtcCp3+m33/DapYuir0zx2/jz1xvi8vASy1MZg71lj0m
oWai552CGzb47K6NAQ+qZJn2Bn4gokdNJjl63onCwLysxTqbnhs8HoIdbAncsGElvl/0fpIBUfOX
oPlLi7yLV74IAKflwrBLr7H555dZ77v/JHLxn/gtzgw8UPwklima6Jd5ryXEFAsyPs2hwCriWIqI
fdmkpHww23zwJIuPdr5mhDQG0apue6D7HGLTtxlIHT4Rwupkw+33pasIOLCoSzlv1A0ZmAmuxA+c
0HEIhbJIcah7kf/BbY3AH0ie4M/Gc2t2DFw1VMfrkH7EJ/3MMhy1Yiz4RkL+IWRduKuiNWiofdjh
N11pyInogekP1d6vZN+BRm1IyZi+zxMiRtvwGVED1Z0cGiH4PgsYSOf8cYGzdgfU4BbJedu8SR5Y
dIpHb+JAhJ6RJ3rxurjWTQ0dKJy/doW+HJIBenpTEzsFcvgHJvAhBrzUqHkqykh7NNEVvYrf1L9d
JQ/EgIfnku4c96boatgPEdeclkHipAvZuzclb5uSXG0v5Cel5durxgHuwv0nAhYZjDbGq5SC/02O
qCGLgS9VWEJk6Hx6ebDadLVwXNUGh1L0WxjMG+sIO/w+/3EWCGc0Llaw9JFYqHUKFyCaPqNXJuUy
wQX6uKiTc2OPYL4zxdhB1FClYZuvjjgDJlEGq9OKsDDeYr4LoYjkbfe3nuX0BFf/EBMj5su7h6TQ
AktwN4FnHLuWJT+IweYn6F7lrgtyuo4aGMcjkyFAIbi7/rzH9CbsNVTrZmI7ydkQfO/1NijPGrJO
ciQzF/YAVawpGZcVjvkJvToXZz355jxsE4WSfb4gHBa3J13YSPBwCtXijg70iIf4QCLldOL+7xxH
XJ5dYorRYKR7Uc9mh8PBSSNuvuCtA16yrkXkJljvlhqnindIsMX4+UUTnwcuGcEdyvR1N0T3VYWi
Aq3AJN6+Op3H8jtlVmaYd4Cc77K0kMrOKngqVVzhO4jKLHVQ2c30FIOhy2YQCJK6u+NPyEfy2rzW
V4/xidBOgtpE9kE3qcqqIwUpvuBCJS8EX56RKxGLIlbPVyWa/9Vi3Zrbrqp3fPJ95t6+Z8nyRASx
vORCYBKRHaPt6tGiW/S42QBbYzoaU3dN2jPKwEjgDrAUArW1BjShVGWGnHnRA1bHtiQgVTh4FV8d
lndE0Q4fCUt3OStcdMSDppVqvhugVd59sAxI7aoSDn/3+UY0E9yiu6LasKkE1jqxXeZMopkY6p63
W0ag22dD/fLQhjPZcwm61smadCGDKdRbXLR4U2+YRYqDQFFnl7n6aYNHd5HikRSmghepNef8wYcB
87rg6KuxpCY8+74gJgKn2oisP+SdBr4J9FKJHDnHWyjFSAUX3AfUqc+/HxcBWM6hJa2oX8kdkO8x
w7gvd9NxKYv2tkHJNrOr2RAmgmctB6PuwyemiX13Gw9sSK812cx7ulOQM9aGD/MVRDJRkG01L80T
3+J8zuOFKeNW2eL9KMf7Y8YYKmgnrS1awMoZs67ao2fvLNyarS221DOPX8UhXODLSj2I4l/vQNp4
zsoYWgcq99wbX/NHwfVgB8NekAU7WfmPtTSAJ1H6bZPktxjOw3Zof/Cb5cGbs5gddvQxHYTpwHGL
m8NKTOHm2uiGCSoV/KaYPc+rVshr8tE4p3mUORanYaB1BubZHP7gezKa3iB3pQhWTU+ABo9T9Dmf
4GZf0J4kKJfljN4OF3EX/YiTXM86hFlZwtLNb0kH2uDdjc9uvj/qotvu3Mcf8m28KB/YLOo8Z7I/
z0kOIY39kbQcO2E5GD7/zz8c6FSEN/mKTVpA+udts9dozDQqYElsyxgh4Y0LkF+i1GHURroUDrvr
yXgx46rsk+dRWBvtio7XazQeiE/E+xo6zqH1m9RdGMx0ZfDH0e+nL3LgqGLewDWFS9tgvNDsVkAd
3tKWJYI3t+qT3D2bNEQEimnC47ompv0eMBhrGXTNHkCP6OKKgflT/n8jYHtTsSP54BTE9ke8ZFRb
PZF3ufrVuPnkp+7Ke5fZycaCVpFSffm8XfJZBpQ70Umpn9Rowp36NxcSWslrioYln/lCNYEUmowY
MalZA2S5hCb6Q/cTJK+HebPK02JbsBbP5q5xPtKIZL2Cyp7SBEFlu4HBdDoY6nm1/ZEJ0MXRCb7E
llvyOUtfhui7H582jA9A8DTJCMhZkyHKhsAtGZglZ+ic6syvyzju5guoON90PoEYT7iBz59yZq3u
MjIO9+Z78noiEURI7YpRLUc9pAtsalcIFLJZLIB3FWH5bVIDG2DhTOAZv476LsYsyZA1QIU3R4rG
VZIlPc4XSC/yRB8EmOdeldydTmYfJiuCWfRkwwRR8tpmt5LiSVL7cV+a3RMGZ+uSkyGOUnJPF8Dj
hP3KjqBvLDA0NxDZjjD65QzZoLEJCHglb2CyLHHZhnA7SlHggselOTxy7v+/rzE4YvBahnaHuXBx
qncNw7YAECdWx9EhUF1AZnNQ/zhvP21xh0ubV5u7nTcUf93xX2AaR86P7MSGjBASIE534equnmA2
TQaLzFOSL3L/W7fu/iDKgG7/FvJ+yS7OPjKT6xB3mXdKuWogxnxZoDunyJHWvf9ku05EoaLkFZ+Q
nGPYFyGe9Yrj/9oXAL4aYNvad86yRV3VN9Ns+H+XPxCdbZFmW5Dh/6tL1EKzmXLRNOTGO/LEp40a
RbAvRFTVonZqgjlAjDJsb9mGzZFrrbG/fP+aPkCstZppt0kGlEbonc/3TAiasl0MmKKV0CVXQihO
0kTn52fFAzjfi7QKO8Qt7InpuonWQXCVKQhnnpKefbco+HIxDkYtEKBeUUVjILpWDaQSwil0PJ1B
1HHbRoOzTrqegjPCl5Xs0FGiEUTSCk8YEYQWlo6DUJtqFvBU1yl2HX7VYANudW4LW4JSljjiu5qF
T7i0r7Dzx+IEWQQwrFtvLARXXEfFByXxLzx3BO18uBEmERNCYwXRcxLdKtqdnj6Td9rrNafkFynm
2UeV+vcw9ufSfvYHFu1q4bD4J+K1tdFpZ5/EZ1iU5eoxi/YaUo6pCFJc79qDHCf6dmTv0qjx6tC2
IRR1Gj5Hom/DhkCZaxaNJYn8XHFOOyaUVnQGrYDpkPE5fhUQPZgUpMDLZDn1VCjSP4a55uKSVtjD
XiMr9JAMdUdzsJFx3yPT5wQ+7pWQtOn+uewr+g/Sj3pzEhJtuqXeN9B6g9DOHnSIn8TMEJK17TCY
4XCdr62o3oSU0o9x4UJo07rS6FzIvPitzBRgu8zZsSsjaQEx49uEdCxvcjmMnJBaccy8dqvB6ReE
+7Y95tl78l0QYk23LBkjITucV3SdToHkislxdLy82KH5IkuxVpMIRYlsV5lrk7gAv8zhmrWwh84f
YTwHJjmOa0cxzruPGdP/wXje9kkJW6QNYzW/hAz8bfEl2SeNXA45Z9fRNDNHOzg9Udg6OiuMNsDV
FaIXC9hgit7yLjkKRERu2ihf/CfPl+CNpLNJcZF51fQfvsBqia1I0vVv8TXuOR6Ju3o6pm5Qp1ZO
a7Kk9UDOVqPSmKZwkrj650DxoXQnZGfYygrTIn87U8+L4Hi7+b79m7BkPGfl8az/G9Bel+nAHfRN
2aA1MPeXu4HRjPNhzyssL4rv+GCMkUezz6ur+DxWOajs1Onn9WIkS3qegTNbgVnyBgqO+ObOkAGQ
grKuSJCIXvuKRwILTNW/GyDnIQO1zHCeySr6ju6bswMARkb6BssbJlWyadJd9NM92Pakdi5c4ppK
X6YxxuyHzg9zTodq3XybJzuSUkK2gtXJd6vVkwLnmT46NHvYbL/9pLq73dWjP7tnLvRhlQSYv0+B
qMfWYVrSw9lbQlXFuMIm4L1rGalRo6KGpL1xiYChl3yHLRnSYSM9AcqD1NES10onOWOvj+WnCp11
VcWZkvUmep04p9ytagc3xGLnbzeV3mo1zpgFg9RGI1yeGJ2SALyEZyPFDgfFWizd4FIVZgMdOvDJ
5ufKtG1bgCrJJb86PIl7Ki1NsXRUtL8oDOICWjRDt7YDJoU7ZrgbWoKMSpgOJnvjposyYhnslSNm
Wh08VJRpPSLx97lcm43WnKMJPE7Os1Rd/D94VCxUJcI2MqSmmB5r5EqEU0W1d2C9TGfU+s9wiUNZ
uhXQVURXKLUuw3tIhAwiuGxNPpTDg38/1PF0A8LacWUhfX9LHuGkTdAuP2KX8klFkrwiGL/tVus1
1+b9GpdTftWqgF4b2+cOzXyoFL7IHBZFASpKK+alzXYHQ+XpsQPmkWcvfO0gRjPdHrK3EH4EUX2X
7ppMHDndLg7jogzb0GKsGA6vQ0dDVzLuLSInrTjXSzjFR7yLDS+cymdF/SYAsuy8Gqs5rwvPjvyQ
JBo+zdwQj6MlkigMACwPeYauXtU8GJRbf8zDqihCMfQLu2a4pRM1xrQAk6JQtUmAOkhgWi/hLIfK
Las4lEAYuiI5Mez/5eclxVrX0uIDcH/svRm/SsRsFF7qTdR54m67vct5N2TX6+tY/o/2CJJ0x9Rj
/CnfWlU0dnXsXOvKgYIJ8RXZhRMmInfhgqYYRlKndcejcoADQvCqqUy4wZBrxaaw621/VsbYKcsO
slOFApf9fFBlQSAej6ZJQzOI0iGKHipdsq5ApLBom1vXBM9eK/+EEtiEXl3Vt7HPPTMNgIS9yoPN
F/YkHhftClk1MHbzbsjK65ZOwjTZssYowztQo4nEuIrgP4Yo8vrfgbngBPDILlrQtFrCnPZJ/pEH
1yewhwEWQ1cjT2hyedgckvEmBE0+QwCmnCKTIh8e/gYgj1RjNdP/c3QYfJlTFdDgcyZFJkv0X9x5
tzTr+ZssDfD1/fRpbsAFBV2+1nSktRTtn+/o2t9bu6L/nFTM8PNP4/vvVFzLJqWiC9mZN+pHaeTv
jNo7/X/KoiLxaE1il1XHs/HPCP+0IQTi23gVhGAy3VqpxyMCF/eyqzoXdRTil6VYFHa1uiNGug3l
yT32VyVZwwPJ42z168jJq6ecfHLmUOsvP39aNTNmZ7V0M6q/5BEBhKmscqj1S02S4jab8Zba3YAR
yxkRpOjrgOHrJnnaTHV4hzRpCGQAwo7Q7tI/PCBYpvp2Qt/xn0t0Dcw4dHB3lzYBdBMethUDhAML
9YXe3sw9TdHEMdd1byQOQjzcW2ixHPAntBVvK1NnnHQgj0PmH5rwC+ORuPh/IZ029r38J2wGau7E
nVHGvEMCx7YUi8GSBbu7ex6+TWcGTQhVAnFc2iaNu7MWGG20G3sju63QpiQ3PCWZ61LM5MimWuLD
wzVU1QdNPFAFenzzfbCNdyP9CS7ZmmC5c2kBHixoPNGYLfoPBbmVmjs5NW3ui3ipWwSr8ElfiHNW
LEAgoasC3By2/DgpSjlpBWb4TO0DwJdTp+kjfiCltIaOY/24CI3o7s2AIST84s+bJ6s+mjTbz5qZ
+INDqUQCUvzW/nyQGb9GWVPWgl7GEyMVnLRbMhtJZxu6+6WACX29YJtFUwCHcaWtBpyrBxn/dJp8
b+EMOcS8/YcXw2+HsdCEDLWmmUUnlhsmP+nTTMZLx2IbISllqaCYgj1ljIMPP9yKDXGgygIFyfV3
9JgNYFMZI6Di/W9YAhloiGtBhUhlfRZqSEIAKbKbtX2ALhU01gPh9MyUu9aU+88VeSO5Aakyulq8
9ECu3lGg00kmhrkIDQcCUm+XtchH8DmUkU/qHkQRbWy+AnhZvPV5xfaLH4GgnGN8UPCDth0zrKa6
KDSYjAN7suul9lassUtMNpqFtx9uU4T0Wixztp5lHMXYfKSgdSa+yLL0ULvLJb+TebcMyPb0bzJL
ZQV/nVuNaTSokssc3L16Djt4sf0XQ+FIbTSFz7GSlIhsPTy5Gj0ATko/6+nqU1s0EvAoXlhVzdKc
ui2/04L2iFgnwFJg6BZKnDgI5CDbuAiWJQtccXibD3uTWfGRIlwMKLApZMBpPqBRrcnigS8S2ZeH
UcD6GC7mpJiuWYOywwzvcjVZnNbopOto0IFGt7BhTyOQXOjoaMbti4NL80Ziy1Habh7ZAUdTQ0O4
DmiuCfoyaWIN9v8GxjCtRdfs/Ia8v82oKk4Hm91khXU1YPpzkuq/kuuBeWiQ3Yndji8t/aVLJ246
XcYtBngT7s2JH34GcIDS2F62Dd1mycqiY6MIRcwmSrKv30vNO5Tt/xwMSrd19kD/cFpQ0hcFRyaT
/hoiUl8hiXnXMPAPp0oPDilDVybDaq2kNjZTX0jVjhVzwLjotl40E0h6Cz/cagiJZvnpFjE2+Ove
hZ8iOdJZTBNWIS7Qim/wfsXH2FErRVm3wxdG65bhrBCdPR3dZbNUGoOkfHoUCppkQ+e5rpD0b2sz
irHkH3ZIakAzPmhFzJDPca6zIl7BlF5LSibnXupYC1qjKJmmqI5jVnReWtjrcjgCpp7S6iriHjYX
m4GTctd8VacokKYxGq3D9hgiZ7oAefx0X7DxcwyBjUba5hPOoXb5lmlqFIh7O1cxEEwL7u2LyHM8
p3E39lkPRpoE+upocVEiFR7nRQ05WfIL6Yr+pr9qItUI60+k7ZRVSakRkNfYX254o6CFy6/grpGX
cmczlR4M4NU5aBaf/GSMyqzMrVfuQYcb3OR611Bz5GV127FcoYVWUeqbGw0XrnYOd/h7HFhbsNHx
OuUWriT5v1Frfn0b4iJA0MUx9jxyElx5mZWS5RjlriG/eBR9xJyIBK94yvGASSRicdv32FpqtzFa
wJnv3Non/nPZPdkn7q4ntwItO/BsIsVtHmGQcwaCaLRVGVmfz71yIcMSnhKi2YZgeCrH2S01qe0c
G31CbAYsBcYrah/E6wba5fjXN8s8oZawGLxOcGITMeHcMTJby0oIH6dXpMupMpX6+7Zgyi3GuaxL
vOxCDiDv8I0uCtGpTsLsmvQZZgYeLqjjCc3OilCm5l6hnb8Gnkzbn8CDn2yZP7o/lHeTmLBNm/KZ
OvfXU3npyVVkFHK7mheVMxpCMr/PaKFJjO3jq5Ah5k0hAl313tK4Z4KUWrVr+ucu3ZwlrCeuY/eq
+4kV+quiZNr+Y2NQ7nPMkyBgyCOjFCr8zD+CDb47iYuhFAEwOJ6i8jGVS3nwwSIWqUwPfdDCBP4D
W+UkvjnwOrH78fRK0zlGsXdLtKhZZWqKlbqR1ZVvEZRzI9cVL/14ybhCBhic6cYuP3ohMMBtMb8t
oDRo4rmxp/kxhoKtZx8nMlwCrfX4V5jmyQhzNDg50hPdD2zksRps3taZ6pIqG/xlm9QbCLiqNRyE
uRGhbH7/m7VLVVYa7MrK9yV4PXfrSZiBeEIvGy03m9QeEYg5+R2xP/fwij2GRAMSsuefoBYxxx21
EX+yeC3ehH887gggoTRcmo1ZNAkXwYv+CEz2XqYRrZm2At3dn4/FXy3vWdHY3ukadDrpoKQJL0mS
+pyvCQ9iNoQR4pNJwRb8P1IlTf8l7IXOA18VxfL0PhEr39CsZPwHinMsSWMCOF3K2B2n8qZ6PZ+l
BSiHfrDyt4zAwSA2ubJE0EGuXOEaBuWgh5nzgQ0tb/4RsyVupB+tNCqW4T0ZqE/w8xt0pAiCccAg
JBKIsax/9ofFBQDLlhMsQJBIgplDrMxCx62TCcZ1VGblytZFhXOzIuBUN3d+pLXvpM0rUBvHPZcM
FJjHP7xYxy5x5jUyoostnVmD7LyH22JYh5/lQJSJcvjt/ytrtQqjhlVSq+BK0DdjDyjFh78JcMz1
YAxYcku8sT+OIEPUQ4BxHOfbV1R9sSM3UniOUoRPJIKrmXiJcwC/gxWLusrl0EqPmFRNoBvfQXMU
t4Rl+6AuLIQf358D32ScrwspheKohEEl/H1fXaxaFUoYnozPN87vdHIWrjPNLLQe/kHUdcJdxZCl
uaEan9xEhayGjzz8vpWNt+pSs1zF3TzPJlZsH4lyb4Ut4GhYrrYxWnrTdxkcqdjRtKs6T998CWOJ
x0b5oNF+5Esf7CSVUHdoOf9tjN/l+zPofDdBbvJXWV3yu1HILkMMGCiG64M+O5ivHnnNFLaFwEfL
yiRPdCDDWd/XnREksBx9OZeKQDMGanUEK6B0TfaeqiN4Y7KjHF2c+gZX51vk3cDmzXk1BVju2dVB
rhWUbuq4TQkc/REAkDYnsfUS8xiRHC9+UM+SCj4yz7oe5nE8I8YCVUZOEgEOkZe22sHM11ZU9xVq
WKdqvRG50IY/BB+V/ZzdUgH4NpYM2dcs86uZ2H4JdmsPRumU7wq6lXVfsT9FN2+X0C0ywEo4VHo1
a2E2FLshRK6VArZqcOgCG7nuiCCXa27+04TcrQ4L/iK0UTUSIn0Adl4q+UYHcZgXmKE20At8ioDA
NkYIyt92akSRWQ5ngoJbs/TZPzxkgQIUzuGbyKbj70hLFymGGhRMncCTAo1KS4ivBPGkt7kqbPJo
7MfFP4C/iFEpmd93pj5PHQluUnWrLqHzfSRrgcT5WlgwOJxEbQaSxETP1FXIvrMXL/+2JSjwECDr
r0ELqE/jVxXKiJkD2EO01Sjz4alK+tKgVCBb4bF0cJQv2bu9Y/1FSIZ5xq1uqiDQpI/1BGdj4VQr
wO87MEb0H21oThdXWRzjux2xRrk1EzrPrmH04FNxCCz0epA94TFrmjtxbMj98p41li9OGOI/QLd0
x2ZRI6nj5KWQ9xBxNoQAerEwpZHdfNAiN7Uyl2w9aps6KpOc3hd0cq9lxIS0HR7M6AKRmOR6rdtg
Of0XDsWF7kKXrR8nCzZvulNacU0y/YbcXPZtYSs2gvZht0Nhm6T4zTaq6WZF4aP6973pPTC74sPK
ymNMDWB0NlSYeYo1nsGxa2pYvbRxpmiwF8Ss3/zQlA5vJEPcNGI2ej+HRWwYy5DSjyXT1eplRas/
8sUbLypV0BLQquujVHLwJ4P6rZvIGfJLEpxkWfDNBQJyWfvZzcjuwNCOYQVmEQUbH/iFOngMyTKg
3ajAaCMp9XYUJLPg5EXZF02kAN9vTTq57pbT/y/Nx0yNCEgd2dc3KvSAFItVvxdH50KCFPASoXo8
fGHzDVr1uJm2C5oJCMTSrtEW1sUjgifmq7ixyRdVknh70++6qhRvzc/UmukbPapi5Fpvb7Fb/eOB
Ar9YPZV16GDp3z4YKiKCp8ZTYq2Ne+1ANG7+NNsGluu8fqljtv5Ak8sb9IvFNM4vSFE6CvIJzcmF
dv+GLgTfJ8lq21IVd2sHyXX781R9QCuXRpvHVgOihBO9+l2g3fcOxgwkEGMYAv3M9GA5SmaCGj5l
hVg4ALLXOrmVbWhAs4kQKYiD9Nl8X1z2NdjMP1qnUICKIdVL9F4XpCdrhZRXsaVJu8WTAhkvULs7
gm67q61fddbWlrZb54S6TflE+Rt9J9vzaqol40BUg7ym3X8ZPIDfvOuF+Ob83MJWPblabsAndNx5
z702TBjT7/4wz0dsCSrvZa85m7bWGhnYlU1oM6lRTLzoKLKUI0fU+XH5DrtdU+DUG/9LSB2JDkAu
IwW8drBpX1N3uF8C1FKSmXwxKMJKj6dzFb2JYNjCwVke8w7DWJLn3oa8Xze1Ge5LNdB9IeMNrfiD
nm4ZAF4i5lRUuKVJqWwW2F9BZugEiGRFyBGKEe1A+wCBXvG1ie6de6zP1sQBUpGsNDNBNTm4b1Hl
00K8ikoFphYIv9iahOgqd+MxbQH7SrFQh/BK2dzgWdwYPLCbd2EGeZwyQZgFyZrLtpPHPO985wpz
OU55leIHjgOY/60pzwRvtwGPbidSpugItW6MQA+Zo3Sc4RQEQI2ObslYJ9M7KD8BPOUGIFO5pJxK
CEy1rLrnJEkSB9bA+AwSF7NJQvANCeVRLo5GosL+tb74mWyXWmq0LiwD4WvGqvOjn/xrzfcntXxP
fRn6oe2975WRUsBKa3a+iPkFkOJr64skv5nNAyJN7UdgSaKnaElW8HzabMOv2THDOXD3GaUXOT9B
TDnGF3IF+xR1nbzb2dYvOTbA1Byt5TrfK3RfNAOLxBTxKaM02YJpH8fpwByonORexg/4p2Fxzpx8
AbH0SYhn8EVtqQXp+Kv2l0kC7CFAfxN6QhySNm7y+VTH+3KAT/+AiSWQr8zL929G9xZkmKP9vqir
yXt2neyBfOtTNXNLzVw64KZmYo9zEi4Kf1AlyKxXpCgCDtuv72vY0teEcoKpapX6dKhmkm5q6M8N
CZcJr1d47f/Q/39VVQWeiCJaF8I0AKZatXk9Ux8FFRRHiRqkkxjT4XZPSyASz3rzLASIVqLKVs95
2zjtrTto4DAF0C+EAfrkuS3uu7g4noWO/3CxXqNiU4XquB+X+LTRMAS/6ACtzT6qPOmS9do/c8DV
CJyNUW4UEtkLbH3emtvIIMzv7Yj/3gKFPdXjx+hmM+1M+cmj7x772tvZGSze4Q2J/S45au78Cp9t
WYZQ+gGaRlKKu1yaa13SzKU5N4+yWWhzCUvJTr4ZSdz5QIjEynjxV0hBquV7lW3FLnebfvDo/Kft
Qfbc3oX22nGefjrBQ51rXZKAXfwT7RSWFK1f51ZLpOUDD7Xf1nm0ibiGCT4fxSMOK7oamg0TGELr
U2802hG1QoTd70IuLdIQIlIXOyYcnRvYQlGG4SV8HS1r4a+kvatVufHmgL/EYgvIDNuqYnjqvmP7
o5pAP+SAZNWf8J5pteMisbpttW3ydywU3WfvS1ownX72HfDTWTuG9+6cK7izfj+SO/W7W34/b8aW
pnUO9W1gbEj7yKrN4MC/yF7pF8a3PQoZOhu8Hm8ZRQTH972cW8sDFx2omk+jLP62gu+E2Wz7qVS3
omv9E0CG7CFLy7QzA6ENlBwY71wsfJw+PiykAMI4GVDZ6fjavmMw+VyqFHHxNIUZhNy9sFVU5dmu
7MGp+MGPpurLJIwaWYYgmyBPSZ+HTPUo0UJ6oeoq/3fqlCvTwQF6KnOvS5GwIxPphJk8Nf1xmljK
mLtbdexFwX2UioipKB4cEYqbHyIO1U97GwyGdGNuGpWcTxplaEaUTPPQwNTqPj39ndhRIQQdwFU+
Xpdv6/nR29rgHJPxSDRNnkSqAcl9xzYq6ByVyztLFYyXhAWACryz8AvMpXceURhMQnJIqg78rY0s
5WezRUcWefxsYDEftxHQRIduv9Mdm9NkEZCvYUKHeij8VL13HzySRa+tGeVCMpMshtlR1kKSR9tR
kpYWUzVN7+uQ/V5VzoUODvm59eajNhcPvSciz7akF7B0M8PqjU2U04vmuf89TRg55ES0DLh4+zHl
v0rZWoRRvwNOptI9433f5NFKPj6sJcBb+eQyh09NrpgnSEnFkHAkZ5YumIBbebtiJD6pHS/QPnXq
yl3Vfck18hP3x0qcWpGkLiFEobFy4+icQV7DOg+pjbGtOxe5RRX0OavQ0pl2t/8MDR8ZXZhHBCFy
fvf9t/Gl8sr8Gphai9yeSBckiE3Bfo36HRx/9aXAi0mx1QWgRGzWyGy0I/wVHAWAKlIixGvUtaQK
3npjGUY9D9UOXmyQiPcltKDhnzz90qd/eU/v2+3uYqIREHMn27HfzxogWPSWYcHWcx09uzq1AZQ1
mE7f4fOvrGExV0hCAomYgCwaQ23Slkg3U7zbIHDxNYEZvBeNpuHv5hcaEehXtr9yO6L8vuSB1o8x
w65r8zbm/MgkprqsNQ2sSw1BACh1OH2wvIjQBK7yzwjhJbhX0QEKUTYOGItHVeAOlKJ1OUkM9VCf
yhHkr9mKI+IbCM0UGmT+PoysYdgVpVtRWJd3HCW92ux4IyCANRsIKJriN3i72C4FYE4f1N87dIsF
l00ApWfSNHdyv54YHW5tUp4KMssgAau5YbBlK4vPWo3kyOnkP1ft0q4jxnsFrIJsaYXTYQfzkhfy
5vGpc6by/SobR1dl/jB1MKVn/4VK90i5cLHD6wG8tMXm6sn9S1Oj8N9QsczbAJBkYNbfLClZC+U7
xKCIFej4o+Sc79AWFOt6M0sGOVdgkYWjOYlMgacjBh4ttUMWyIv/gl5YCLLuCGAn6OH6NRqFkudp
nOjwZ/0MSGKu+UkhnTsS9hmScmxAtIMK74K3MqywNPhKZiCCKaRnujdXaz1g+YOIPIUWw6gq+IR5
aTC8xuPr4Tnn+v5ukWjPTGtsGdewmk1Vz2x2nJKkBkqmKK7hn1pUNRWaM+Xd3gINsuE8uuY9heKQ
fuHTDaTWEfe6B/eLPq81JnsR5t/2f2Te6CW8q4X++6YiA7W9lbFmIO/uDA1KuTYq2sHv9hkTq5mq
6KVbU7NNlbidrq+Pwj6cFAwZERlWPen7/AoxVQkhTE5kIGT6bh8YE8apYAsC8FoFGaDsZLag9Cul
shpmC1fZzx3Uss9RDBRUrg5akQLYf7uDyLh8qQOvJleRKrRtSTSRiNUxRyVAbSV4Fo1LqFiZeGS0
VjhlKjkxDa/gukf+3+JjbdXRZJWTVcjkk0wHeeWdLrjnbQ/X2y3RHa1tb8vti4eyVPkL92f+WqXC
mZfitSYIzBs0EpVyPUVAFeQ28SokvI/G22vvgLPHdkRmBwCkRH6Ob7mRo7VK3tYkamWj96B86tOE
ltPlNBS/IUYkOSlXGSEVtIQj9d0AuhntG51LyPUEdZRDHl3Jr07r5fYZAVptpfvq168lzCnUtheE
LTbtJoDHG3wYg9qj3kEhGxDRLsgJogK343Bm6vGTtCTnlzMJOFdN59k/zIvMKarxIC3YTGo8SIZR
A9DcX2iik7NmQyLkJhpnZMAM+ed/bLqQIwhPPtnPVG7viTvPsx/akmEIQnKkHGf3eSw31WXs5d6C
xqioP1cWDQdAq35kVz+ZuU9qa7cQTY2xNJcQ/Bl5IcMauY7EB5OWgPwxJeX3tSGPb88Wr9GBgx3+
i4of/4g0MpsNVNkq3WsJItyQQgfDKXCqZtvvgsWYZUPH0VyRH5IhD07h479roxWQ5o1UY1aUstOk
UrAkPfQT+s5iF6spsYIgcsCgN7DGoMl7983ZPDHnMAwryvoP5OuLgGS8cnDS4Q/f3IabdJM7FH92
UuWwhR6qT4Kb0TKgPW4afvDUuXCgkuXj0MAqEImFZAxn/vSsRnrwYJulycRfxhTCIMM/tSZYvt4x
t1aSbBRLJPBsh1yfsJdylvmr8U8s9O8w5BVGqLg1Udk7jbLSz7puSs0/nZiHIl2LvWXbIldNrf+8
XISpzJ4wGSk01KcV+ZmR0+Oe1XuXT5zMr3tkZcJJlA5KvtdMqpNvDpg3IQAHLwttlLvL0KvToSDd
i/wttp513qIEFxP/XbNj3FD+a9Qg9eBa6TZkClLFU+ONP1SVrFtvcTHJaibqg6A+mvGfmEdeXjNp
ThUX7B3VctKEEdNaL9X7EiGGOxF5yB8E4UK3m6u51FTAaMNkQK522xFzz0U1KzoYgn4krjXdhvNs
J9CZpBGRUWHqUZTLcPrihA3hk70JSPTo9XGHBjAy6ge1lQaEmfRzNVn9A58nyisqIuJ8WgpHhFZP
400YnX8WUnfZ6tOXIpl85r01lCPKEYo53M2yCu+qKPW/awyGa5L7rYm9hAReCaTwFdqtitxz6FG4
gRgtKxMbTIjhPSYG6CIY2sbB5UlWUpAj3ywzDIZePSuC8TFkHXc3xkZ7qaDfacqIUhj5e3/odLJw
1QpB/alJOVPJrxCYx0Tx9D5FD4Nsc4Awa+uzo/n+ybaS7+mi36mGQJTNJQ+r9SFtBX9CLFsURFuH
iqbspUVzKchizNTKLtNRJ7onpilb1bBMLcIjmPJW2r1sbucCzXcgopjW91EG1dLubtWNC4w76Upm
GJssRlMPLbIsI64GeRC219MkO9i0ZV1SR+ZPqyNywpeW+yyqc75kjl2733l3EU/7QtQeBuG2zRtr
PTz75s2uBkS4Hc9Qf2+/JTMGEVh1ZmdJkbA6cCW3Ssx6lBJatmZci1Fcu1a7ZJYkA41Iom6VSrQp
s4U4Y3L3GhlNCmIZUqJQ59vQAZP+3CIweZOC3RsddczZEEYML5c70R0mqiawaXZlLLddVdLC6XCH
yLJ2zAz3p7rhLysdYPt0ESjZ+yi/cPGAPuXZwzrZtQEcLm/1IS8Ok8d+GdjOfcdYExqwPZHtnLgb
glEbvnaD6jI1ops0TZKz7+CPDCw9ioQl5YTtVHiRndkU55bqMjhr3KoGoBEkhtu++T25PnfQF7W6
3Qp5N0LkoOsHMbL14PcIKK5H33YuRhpXs50EMu03/5Tu8o/VW+oSMXSBseHQTxneCYnWNh93v01I
5/OR45u+QxJNhoE/tw3lKmsfu+2KCHz8Kyl0VhcTvAZy/m17U3mT6u0BqIrT/Fy5ROpZW/schAm8
ZIYcVXWjU8MHfrBbxRuxne6ANsVVuu9B5ZACNLwnuC+qFe/a11IPvRinD5lssXBmOlaGSbFnL9+H
a68BXbgk7h94E17+dr2kVWRfKaxdwSGSMKIxEPWBxHN2dYWb4/W6IWpSbp0OPCcDgY+qo9r4kegC
TcSCBUayrpxfRSUKVBALFiTfHkYqe4BwttxoXs2UpWdDgIq3eXsjZq8GwVsZHNx3sPi/zax0bE6z
djdooufO56+TAflCb/yun3hSNmgE0lrMTYOVBceLVHwJVmwFIqo8TX30JZeaWqeO9LG3UoTlhuLS
ONcyMF7+NCg7wtHeM24QV5CaKVr0HJutaRXyzvCUzuD6LdQXhn/0tM60U8Of6m+5iOs+jGN2BNxT
T6Nuyr1hNOGhjyDhIfGJxnk0oN86cc2H00aQfMu4hFCVtgL1esJv3Q2hmoAKiN6MRtdcyjKW2j2k
VinNJrMCgPqG4p9oDZgUMrnn8kFi3+7jrlZCEPdHWmSmppDTdbpe0jyNLojaXy22otXSEVM/CMWF
+XiR5I9S3YeiWq2h9sm3tMFly4zE4aC/2Gpv81jTrz87SjcDu4L3cJb3757d9NYuAuQ0np85PPAB
ivdXHUActi6K/wAD/zzsTMc5LLZbeFPtP1uNON2oNiMUzBNZQ6ob14oG+kKQvmHcczhLHZnu8xwQ
w7FFROYGw6RyWxhH1eWBoXIgSV0qCBRfrFO2lzdUDEyUZ5SO+bmmoJucAOw8bAl+imEYdfuCuDhL
PvC9hy9en73W7G6KcEwxphKIjUV72yhXKCqT3KYWTsdmsjZXVPkXG+8y1Agv7iFzOvOAPUucmEWF
IgjW40ksrM5ZAEEk8xJG9TQmocB0Cf0YsEoYq/tFX/Sw1Peb2vuPIguybaTeq4ih6LC3WyH/DYZp
3UWMV/19+xwjr91kLUdRaoE/lXkveTpJQikyMqtkwBt/ysoyrvYVGX3++4RnIsPIn1G4FNpjSAqM
EwCrlDw1Bs191VblaoXBUnaUsawUlNfwyVveWxI54L02CNmDcGnDkc7nCXqC+DoSSoMKoX44X8rA
0wyPxFcGz4BLLhF7xJJWPE6/93+gz0Tgfa4FVnoI3Tu5huqTalSgz7QTbDPvwxZjpLOFHseFRXkS
GULDfK+HnzxvxtD6G9UYttnbNJMDWqZoNH5Zgxzxr7g8rWPux5Wc8L+6XnZsAtxMbEUDmFR48JXp
Dv3d+lY8xNX2yJFb3lNW8WswFqM7pkSWTTecAslhZcJYCbR4S5G1HbsWOIygPmJLNRTTzrYD4YfK
2mKn5GDwg2PlC4v17RPC/IJK8LtmzXZS9vtLSY0MY4Ajn/XRcZ4wiTadtDfDDuRU2hnTWsrc5oEM
WPgOUky0Q02F+QJtknixK+KUZ1PV64d+y3HUV9VrOTEb0rxkzg+5tJVwiKvqCbqBMHcbEfenSKna
TpyRgGwl1mUXyEhN4IrvI6CvD3kBzIAGGl3mZyz3wexCnVWUNi7NR0ENY+BlmZR7jBGo5T5u68Bo
PoU3+Y8DntkXd2rrpGxfj85AqkXXJvDxlyQIY2RE1OaZ1EYP8bAm5+qVHszqH/zF33jXdRvjunkF
cMEnmQPGyLqB4A4Cl1Vs8O04YTqGEIjOfc0LQdkj0i2cV2f/JzYQ9qwrsnyJa4Fh/iwDLpSxj27g
zPzBzBzQHkNAvqXaGhzj4RsOzQ2nqQN/DlpID4MESnCHAzNdwyYo7+VG60oSX1yn+WQAvSXut+Qg
407JjFubpVyy2ct0kk1BLyHrIiXyUOoKNpTyX39u/IqXA0bo3KGGKE5G0fAq5dIg0ipjDnGnWrPe
/H4j1NcSmQ2P/axiH9wfQrT35q5dHkrgIg36WNri8F1S7DNlJevwQJLY+3I2Gb6QPWIeLNwsUs4T
4HpfviCBKQJiS/X4d4ZZ3cygULO4U9XPAruU9bHi3DQXyIHydbmnvO2SVatWm5Doz0SJPc7nUlfR
H0Z+Pk8bqst91cdW4bJ/+BLs+JHGZ6mDynNg2kTMt9s61QvgArgZkVQbX7EDlC/ZZ3TKi5N1s2QL
nyQg0Is+TQEa+/uxwQdC+ssa7EE16bDARO5wRgQp2pDZN+ErI55Sc1qBxXzBXEg/4QKueFLZ/LRi
C9RCm2ubX0mYvBLvr8n8lgUss81IsKV7gZCX2p0GUysicPxYvLonjg+FZE1FsnqrXYZNZMk6UhHQ
iOmtEVgSxBzFL9Kg9EKtziCexuoo+OdXElnst6+JwA9JOuv/8ZOk+e93HNv6+voc65gwyYUZt8vJ
YHClQ9Bu1dY4smPH7ZANMTEFG1cgWEZSlnPy+fVUGy/Egfg401ID+zd41qJLK1X6Ykepb15VTMfo
iaPX0MPN8PNP/3NI13i/b7Q6VUOSNGTvZxTD1dzb+nmzwo8JQrhumggag9gHoj1TaX70PkPoupPB
59OwKJZV90cJbPh7jCJ9ovrxYGakk0OocTRAbWjy2wuYdauaAMEIlXG/rPejrSFh960G2yldYFIW
oDK8XBPcPnIfH+D9MkGpi40MYm9IhLiFoqkG8ITv/4iaxWD0Z6ruFwDQu2TD4uChDdnTLpSwdJ+0
smvQFDWFiS8i/K2hv8CGQ6vmMGbEpsj8jFfXyaLQx1/Ft9hPZVABAogHjs1U5tRQuWkb/Se59SEA
ijyHpmJ+J2/35r4vCWSjjG48SMwIDYQH+BvfQ15IliVzrXkQI4zNRONbQthJFHq7KexS4w2J0n+X
Tt9VaSbO5VpTJh+h3F1NXsyJtMvFZCpmWalXbVsFcOSpfmyRfQtvGzBixkq/hv1eVwGLSgU4/1BE
Jgxd7X6/Gz+MLpaY8hPOT1aC4amZTQi1Jr6TZWSWoq66bXsqiSw+jUWvfJi16o1D/OgLZFIsNiRF
4ovI36IagwobNVyPKHYFivWbQlMjd4fDizKYwZ8j7nyzkVnw8D3lLP3AyOsZI3lbLwI7+lIg3D7L
M3QQPkk55+DU7hdHMiNSY7dUEtbWDfcz4xn4sRzlazPe/WdhklAtyRKqsYbrm+B2eF0BgCcm8/3I
1owULhdWMYTZR6Zpf00/y9jzXcTx35V5ulfFEaJex4Q8agOSF/amddbqu0ZOAAh//W8AjDdyI62B
SG7Rwzefc4tZxQWwecI6KWiO33gQQEh4kTygg3TONXV2Jm4UxKA5b0hYeNstYhLFBOekXi1DiGWO
TxadPxeO5gAih6Ulk92P9OivYon8gs77u+bl3c0KgGEvyKQyT1FBve8irIaON9inM8Fu7TWFortB
/uljUND7PqG2J18b0rizTNs9p1nlVwZRlIsEjcQvKI3kFhBJwus8uhuUxH1CSr6rwSfb3oCaycOt
DK4127XKiB1znsRV0smwZHOMv5qfkRlB/Am0CzDxARTfykvD4m164D1UfsYV/oJquOhdTWGint8R
/Dzj0FSRvFVHu1rUIhjauWA4uYn8vT7K01hpSO9sEc87zZh5LSLf3/ORP09xP503tZlZtWFNLwi2
ZDW9xxqACvcT8CeOHrKyodvw50p7iGZq6jMtzlFzwmKkaUZRHJiWTNbsuLlh3NWdw3qRAN/pJ6qV
pBb8xzDbhUoVEuFJvJQD8c+p+Qe9X/wdy2zSMbMmZgAd6ZxNrsQl89GoY6XkUiWtWnHexCO1haYc
7+RN9qv4fC0C+GT/qIOgvPQ6YXhxDh1kKfFMi9Jq3U7PR5nyf9xzr+kg6tQzm+qWcOnkMlclpDnz
iK+aTf+YAGuTI1gfHRNIg1zPSYjpB+6t0DiDJspFsHFAZ+BXlUtjv84tZFXbEqD/w/0adu7XaxTN
TK5dV8crnW36Gte4KQEq1uxjyp7rlbFRBfb3VHPTrSZLcCjvUfPRUwwAtj5aNcc5z0ICHTVpYsAx
TGkZ0H5h8IKC//z+Q+JOE4pHlK8og4IWPNYoeiNEyXpSlL9XYEuy+UcASrGo6NOxmtT76j3xWRrn
otZw4TojIyFEEpIhrCQiYzfqcNt5hlinLwcrq/6HNRT6BHV1y5OKHcWVNgS6a+uevbssPw2tjC+y
Up0l/ZPB9bv+XcYeRYzA1g9lTCMqC6d2g/fckxh3Gh6NGRXsC1a7GPBD3qrHuhpYPAUtpCKmBXzP
/etZ16PBiBfMXmS1HkgGZzgWkj39Or0xEfiCWHUnh5F19RyZCp0DCwjD1DYB9zTQy2Xi7ldRRcOu
2u4APj48RW7bugwki8SLWRDK9Vh/Oi+CCL6c3ddffofT9aptWg4okxMZ2y9+6PWB9aABsk7Tfast
xrYS/4fRX+mJECQ0fDNPCQZuo5UFyN/+qhtiXnXrwcpA/B/cSB3nGxGdnrIxLmwDPI0zt4zsm6Ar
CukpRstl8BMHG9Izje4qIxihr+waPnWC/djAaG4HxkGnMAMx2cdFsAHvC6PGVm2nSGkwDXA4pKIC
kW2YS1IP7X4lK5SNHxnemZxYDZ/0kaBfH0tUVUDUGmmaI0y7yrACdjl14CVqyHx4+C0+xvilxIRt
W4NunVlhJJh8UPWVuYICRq6lisC2XxS3pttnQaLyYmpfE3JjrF9KMkI06Z94piXF9HUbflbQ7V/P
PGow0rEr6gpC9caLZ2d9pvp/XNRXtH48urpc9W5DUTvMd5BZDfJSiZ1VaD+Iehaps3lSBN3SEXDC
FD+ohNu6axgaQCCehUvlcM661bYhZyB0UuOSUEVEPupu2apx1qHda40UL1w5OGe+Jdflve47VP+W
nvuuHH0arS7WjOT8wdJgKCnftms72Kmo9B3cXCC0lstUYxFinoReQM+WvBz+vhfisiVU11s9Covl
h+CZNEkyE0zXNk8j32yEV8mfzWRAjEI8vZTPDrpyqtGwmFD/5/K22UaHFm5uOUTjXcR/cEBSgaLO
Enj3oI9KHHvGc4GFfYrI/G+OChTga8e3llJhfiJe0HkbYO6JNlcXwyls5+3+a0uyRF+taJaxkZN5
6uZmfw2WybORXrZtjU2w2Jr24MNOH6ck7ZxNf2FuP9fGinDCc4DMjdwkiv1LMaT67PmlomnVpRTM
1Gz5B87Bha/OyRqAGz8ww0kYRBkPtm/XOFPY0u0vBTDcOnPK8Nuwaald6lrrNoYeVRM0tdjKvMiu
NDhI7C1G7vGPFVXLPx8cOdxbLYR33F+HhBjWmHrrChrBtAEScgr3HpqsNBKHCdtYRnWBQBBfx4Pf
ezQkWKHsjAySRIJ+yliG65cXeW524HM4pU1BpmzyhyGwup/3Ap3RAJV2Y1+McnEg6Yx8QSobQZTq
Gk2e1llym5hoQxC3hIkwuOgsCWqCAVcSk6+itqlL0b7sU3FQJo+6nXMKW0pvVU0qrtVQjc9Kt9h2
D7PRNP6takZOeBFICnxXsMd54xYhf6fnTpu+ahFgUQQjaxa/eNJ+o/OQH6ztWRYfqzROWdF58YMO
xwXe+kWik12CtfgtsH57iDhTd6N8tGB3oyyu1nACkv2iVX+ci9iQj2gDUe4hFnbU6+SjfPRK03Jo
x3atiCt/0R8O6LuP+3st2/qsXa06VyXhm98aHCTrGwHIHKVnXY60u6HgBMMrCu1IWYShBIIAZf3n
4CxJqwfhYRc/7+b2I+Z2+i48iV4PsCquL890mZCknKeV8K19yJ/Sr9DvNoCXg/4Clr+KpYnpGRpP
lezetbzcQ21/YeutD1/5GlQ+j3eerpPfT6sWzOqT0Ku2piInIcugsrYSQ5R3mMxFQpYGw9ZUQ7oR
BU5At+ZvoTTxpXFxDBf6LvqAoQxqwRYR4iffCoo3gPIVaDGo+TFpQAn9ASlWucwI3uEP5jd226nT
fxpr1C5qQt9guAdBtO7UqkEP9hlXMXDCJRjajuUEP0hbpElez7cb9ilxWK1g2aC6taqW38d9SsKv
Cd8VD6T1x+t5vsK9fQRSiHy2+HSLbqfGUclWdzJixtq0kAb4jqY7mmHNCVFWqPG5+mz4MS14lyUA
f6z4UMekPfU6wDZOP4XFzaeeSwHGlgouF1iTr1aSuztmBifaZjfmrDja6Ca3F/Ep3S/O7a7X53go
yTY2blYz55Ma8eGO2uHHaJc7m04cltfDkXwVZk3Ncgrr7WIfpAsnhD+4uHIYyroH2OWQ2BySBoG5
OG4h5Ef9+QLt8C18JnpMm7rJKEUtxEjHo4e2tDhudm4usv6FKCCs1EXmUr36GSocr/LNZDgJZuf0
OeuXbelVfI2bytrJkbP6Q2ou90XHCis31R66HKHvitPBX6oLkoBloESdMyk8DMl+QW4kUDGOYsiZ
CaHflrA8fPGv1bHsyUbkZU5sSa/hRV8SgwhSZyrU8xQcpAaNu7UA13DlXsIvN4Yg/AvdWRahE8NQ
oxtUeTW1/uhkS2kG8wg4qle5PurksofUQmMoNqUjLWVwKZm+1HMsBmwahQJ5LbpAqtOL3VRnj+8e
R5Ackf2Ehl1IEgX3jXD/EJkC0JvUe7Opu8kl/9SHA10bq1IHvgwCHYTbAmw0ElDo/BRCTX1b+cdK
4DnqCNBJ6jDGzxFLFN+fZqXr9ARIO25fLD01HUTL6hyHQ9Ja19OmgTfMp16z+Pr8XwZkhMz8jOSz
BGwIp2g4CE0my5wn1sD3jJ6t2DftJ4Lq+RLroG0JTCZz02fUVYNVXdiItcGqu3vIZv3VV4EtuzIe
9BV79Ud8pGGfIn1foUhK49oHSMrjwGitGw9XvcJWeGoZSeUwcR+XzZQzhYIMgNHnyQm/x5nvfWg8
/UHzZ4Kls+DI8jx1K1+eyK0bA0xIHQu8THU6AV9RKVVdZyIpo5DSwvLGaGl1heai8BRynuGpAOhM
qqEYygbHkRD1GkZIvjgKw548oo8xAgjuS614E4HK7Eyf64D88SZsF0XicbmX5bDzwxm/dUtuEvBl
lRY1UcEhGNV+aDwyWWH8V0A2lb4fhF68HcvcQZtvN8IeXxmHFuRwlMn0vTdrJbB98/N092r+Q/GD
RYCgwQNUtIYcuEnSopuG8OmfLX/vK8F58BUhOyDp8i68pjxXLILVO7J9uhuYGAs/5WE9zYcl5omE
T8hWzNea7MsP9J5/vW7uMs4m7xOfAkX81lQdzVKIyY6sqYpEhhpI5no+YKtX95SPbQfg3X3rlxHw
ijtrVW75tNYZozV+PrnYMSPQYbT8IgWBouJYisj3CAGrm/Rcv7gTuiugYktjOEmypZEFjOV6QKiW
iVKnbQUjfI6BhxswHyXYt4UAU/9Gx2et/FX3xxMM6EKWpz5g4GQ1zgS0vB3J8FnW7obfYI0CizZd
tvcUQCDeBq85YUf62LMLc134ocEOOo8s/yijbj2lTw0JufmBi6zPX8TBZeOpJvFfcMEXC27+ARCC
OsjgnF6y3zfGZ9ZClzzaIXZMhgHTi8kBFHdUC5xEcYux3zy9rYNiT02+xNVnC3J4IsEoYbsAv1hG
8KdtJXvf4PN0JNvZOST72lUQh4YF8FsRjn1gK0kv0FEE+1hNCPx84VfFAH8mnInXofcMDmBszzl1
IeyJUoMocAmlgwujNwpBdnvUIprWRwklmbydGIpBxqO7vRcNMqfevEAY5Ng0H7HCwtDBoH/ckI+R
HN9xiJEj44BV70862+t+c2KkPjMyH8/XdKi/y2EFQqPOD93pZtpzzXZqz6Rgt7ubd2qBbWFBc9ob
/atMeKqGikMdn2mcW750V191aNT+aUdRc4D2/ijT+e2ITVcc1dHeP6DuM5xEYMu2Y2t3/DzcBTXP
qffDaKaoFy33Ay1kJLrB0sqauwkq85xWAR2Az7dnBqr84d8OOv5p0NI7Kb+INoVfLJ4VJY4dtV/R
nQ9bZIfn8KtOXTQpWR2/WxzgOf/xzj0j56ZcsiP2vEe2BKfqlME7DSkF8hpzSOAhWhJA1OpXP11Y
roUqkPm5SSZj65ekF/lg6OQ9rKSPkdl66VE5OOJrXi0aN3c+NK5UpaRZNk0mN3+CSvP8b35VPWJU
VpxBLlNoofolO39j9vNgrgaq/BFHrddotNBLENWBS+k3EANj2zIlkCisQWQfQ0vIiVINiLqBNk2n
Z979vZbhskNMgkGH5wS7/LnJEOpKJ0bvoh6BfhVZX1hWwyuZDOKVpgWwD2zmHrb50V9r5ld3fYvE
IqcSmFiMo7zMrHqmbG/vrjfN+I1x9QspKeJQZf6OkBsmTYiQ3PEApQXgFys5mNP1uQMegyphNn2S
PmLzy3rDPhOEcyJ9oYq9qRGR9IojyFryq347mhF/QhktOJBIxbywGUv2S4SMlaF02aSV4NFpNmuN
Rz+U1FOB5g1XHyw4pq7R8YQ6uJWKaSJ5gxml2r7N+SIllx5MxoobFzRagHu+ub0XN+fG+Z13sZ7n
tM9MdXQZNR/3xnF7MV7NRCkfibvyXVFkn4feHmc6y/jSWrR8CbaT+Fakt0WOxvNteOrWGFuDGm39
1bwbmM9mkqWDNxt5fYpkmUL+Mz+JgrfNS94tGrQLZRjRaO+3IEbmXCvV1iCnDoKp+OJAJ6RXXjUi
OGn5kz4hAFw8Z79OiAhJhBrs/D8g3paIisMUmIpddt5+oGTqh95r4AfuUeVMp7VRppbHvaP7leq3
rjnP4a3HK+6RcMF7d60I0hnykCcHvCtvsnPFPnmk8mIG45WUUWwTdoysozvmo+yxP9r+Dc2eMBS2
/fGEcBVwpeuNNIyOkTVoqV61Ieroeplzp49rPwG9dhear6i+/fyH8D9oEEL+P8CEQr47FMrciQET
aCCIXhuGxqraPBOxrx3u/0y/iLIFtwp52wGdLPcN5r7FcrpMM4S3+9Oh64ajz+DRgR6Icfa5p+P5
dPy+2jakB7chlaamdzuZ3+/o5ZxFK2baj8Y6xD2r81tK+6QY7sGNeJpLllNpKuFFNlouuKQ3HVRz
3u9XTB/wRQUJPjhvhhp/sBHgWgGjps5lFJFU86BYp/2OZi9vwO3UWi87qOpLGvTfFoDuxzxapKVK
oaJe+E0AGbardqO1Y5yErlND57Ui+aucaJq2B6hSExL4Kf+122BrjnJYe06lNjO74stnj8FSFGZZ
j3oXAPBvb5iw4Z2ZyiCmurzfCrEeZumdfApuoDMqVm0Ck4SByvCNmPYOXLXnkqYEq0XBp2AMo0+M
Icz7/AvO+/qPwDD2a7c4mFkiOiQ51wItUkCPQ7wATap1uRUYIdmXGNNaEJ/72ZlJoxBWCSNuFFTn
OyakSlOEcYg1o7CwjPyUNYuRbsYW/CvCcEClhKh23+N3tKRtjAvB39y/ixewfLNtdr7N9ukuDtaQ
NXIPu1Yi8TX6GoLucIDRuTzJEyGqpR4L1+hXHWTbgproehf6GxFj27uGVHUUByANbmA0exf2kvEU
nwu/Mp11nIm22T4TsJlcBWqU1NGUOTWvkg/z2fHJ+HMc2h6vT3iHjk4vEfaksCBVKm9qQBfSsShw
qyUFqKDvAQpP1laSRlxaQ4MSexR5VNEx/7eaG4WiDw6tpbh27mFDmcPK7CGqqv/rlk3gbPWwSCJZ
/B7Y7msgOM80kCwuYB9ASQOxsoT0nxW3RrMVGLfjh9Yp0f32Ey2eafXs4noMUp/5h9ZGmwY1O5LX
4YmSiN/ja5taDaUMIeIlgR2kFnbhrpWnldU9pjmaCYOQ+gmGIwd+wBDLokOeZHutJFura1vDkUcW
pZQVmpV4FLmve6PMzY2HdllIt7bPCPj/LFCofgJsWJRgM/rojzHEWaDPz5iqjtcsNQGEuctA/tft
b5DqRmJjP7HC20trB6ex7UKNe3Aa/bbKAb3ZTtn+EEsALubLGlM0C+59VkHF5ybJ/AvV3auqtsw4
e6bKFNLCd0xRvUbLv0NdbOxD83R8ElueDP6FUf5dVqEvhdyPwzGzCqSnulwnLLWvNQ2RvcbtbcHj
h3cVi5h2+yn7ltv/iNf5gxC56IacybB0OljufqqRj5MoEOKM9S2yR+BmjZ8YWjujx0UV4vg6g1P4
UVbnDRhY8SfkKPva/v+QQS3fRioS4Rt6QAsTrERisAXqT1DayhBCQ5J9IyghFExjsRYTGn2IEbTT
3Vf/6oF3/XqJAnS901OdfaF/EQM8hAhElKcVNm4/irYzJF1nbQtw4lULPxrp5sqA4QQFaruNWFXv
/BH78fyYgMgSMNmHu1aGrtRI+Wf3uB6BPDYRrBAgDIcW/oru5FXPjJTePC5MACC4slZSWBT4N0n5
ngH4SEDOFsmfPunkIb/r7navaLzmK0V/jhFlPIju9QKsuip9F9tApqhjcWb/VPutDzVTlJAZE011
WShNbs4KKM8dppEAFl6dlbsy5/slVug7ZPQUQaFGCJoPNHxoyN8I00rWvfe0qYmb0II0OUOfjIns
gTFni1t+MrgTK1i1Vd7XQoxfSok4bTtHnPr+2DfuTDNk7xOUjJxERYOqzkAXDDwajzs3msYbjQxW
EjCDyilaUPy7orIDmj/B/mcrcNvkX9UIpY8yql3GDf3lXybwWgH4+1r6TAtRqJJk8iy83RUJHIwV
uoCgHD6cpFRSBtCc22iT7XUTqHpp5WFlerQUbRYtMc/YxrRSxY/gvnF3AeHsLh7y0QHvFNgrtKaH
sFnaNpbMqgIUNvYXF3hJucu0mC/vd9S8UCfBtahK9XR9KxfwHL9tNBKa0WEmz1wzEDZFKDGoeDbh
NtOdW39TSFhjL2Zc3Gvj+iFDbxbQL/xW4Z+uKahGf98Ur+0OJ+MntdXBOaGPZ6RWUxPOg9RjIiJ5
UTAUTH3BOu4c5n23WMOnSR+sF0D4NWkMMxAjN/Ka5OTcdAL08n/EB9KkOafASyfEYfbvOXgzn+ei
PA83mZOBzYjMv1TPFsowkM9OHcKmLTwubKbWu06CD+MKY0OFwtnoDjDe6kbNCM7uK3DkY0A6M1K9
JaObTOPAbidAKLCO9btHENnmVX9f0Jj44LXqMUvoUzUNB8jywiO443yROzpPPxyuvtWoCVKCbGEe
sPIbjsNggaZo9NKfrGm/491GyOEhOhrI87MHlreHtxb5sDVRFKgUxyebCkZzjTfypt+NwYwAvoxC
Z7Iw6Eim1/g8BQZFpFOqskIFJA/lv52xGJYJe0IGX/C6me7UM36PDmfUwgkXT6gqb2AwvONhVp9t
c8DYQDlsmEPW6wniq/9YULkEsfEN0DU0nPPsgeOTgjvppwqPcbNCtFL7j7NNAbr+SoQm1/DXP1NP
zm6PA4I+9hGzL0shaas61hmuzwhvAMDUW6WVJvDc5zppR2O8vx+iqCDDvOo7Bkc36u+uR+2s3pQt
yILJR4iGi18yRfyAHt+fOF5VWNdeqW1NhA7yhCRMulJEmVLFD6INzKF/KJbOLa084F6cO6D57d14
RaxXtNNqyZix0g2kZfvUGmRwtdrWL7VkBqePQyKb9Y1LidOg7E1AaaZg/SHl91VTasPDUzp8zeWl
jmzvMA9a74SFUa+ELzvWxoJwVo+ngLdBaPau6uZ0HcG0pAV6p16njmoGyrEHQUnzQBS35VtIcqbI
cBCDNqlBMxnGxBRDJ4UagTyRzU6jHKvOmS8LE0mBAA+qDIIVwdvdRfj/kz4i6GuuvH7ndIf6TK24
Vf3vEUDSBYkjTdSqEdGdtEzln6yejjJnM0fVC9raV555TrPfVH7oK8Q5HZPpuEEpketG7QE9VIjB
wCVqpiQmby4sbG/XaBFz0zVvsnnworLatSHpaKkv1Hj27t9Uwv1OcHGJHUu6zjCdq+D+aZ9OY2CC
LjTtBRhWyu4+fRha0B/8qqPuEKKoi5GiQOfRbTqBR+s47bV0rWSwPpVF149kXNNgAiMwcYKEukdg
6cmf8nXy1SkdEu8vCQhZvT3Y/pYCf7fr8gEo+/Vb5j1nLpc/FL+/yIO6fSE2k4xkE+NIG5KGOjO/
+BxV6KFagxXjQrGvbp3fxIJ/K5dstPpeqMxU3v6h6Zn1RIKnLWTN7SCv1/w5LcYPErNVtUTQdZo0
f0IOAu2c3DyACyH6/i/yvQmL0u1Ln4ULAdCGGhHg3MBQUK6KWkQ0xZVDd8P5XdxQHcptDv3ozo4m
gKY065ahU/QaF0kLnSlrVGOX0pIJDIFZGqQKsmAqF5IwDUo78itjd0lKprJpbguslWTyz1Xweg77
mTKzcgtmTV+9eTLbE005qd2IduHo/ZR56EgWVNzv0q8WVNjPMNlPU5C+K3MTVf/vDKcjyF1aq9Ly
JnO4RJnTawdjlITAv87B7CPfQimySfSRhhnnQX+dC4ebkvwq96ij9smh2Pm1t4FYkM9zEHv2SvCD
IzIuRpG74mFb9LKv4xrnpmJteSnxZ4PnPQBzdutUNndVufd33Rl6tBLUivSzUXme2poJvVQIxdXg
pLloNvQmMCPZLIapNKvsrtZW0wN2Um6k42Y5THXPhp8rnbAyKVnr7p5QLD9Snq0+DjHiojzxbmy0
PZBWrIuOfkceUPyfO3bKDlVCUCFQl69qEmblPU9GkVYtXOhGbmeFwoc7TAAEbq58XSKLoHEa0+lM
KStn5iAHhVDIvfVN3Fmm1ccIMuL1UO2V9U2zegzn8RJpU0wlS7Xy8jnboxxFK7xr9LsB6CaYtJ45
XmNQWlYss88iOgCS8tTizWWTLmpe8OZbjZ+PyRjpDkeQkuQx5/3sTatc7FfQlF8IcgfehlvfHnz2
Fk2oJMlqLwPPR520QOU0Yq8XdDw+WchU7O8wSCm7y8eWcmNKuY5GbJbZ4ATKvok4djWVliMHJYxD
vTtUqhcjDI/GGKU/YOny78dz5/hQfCCWT5WSXsreeFTs0tElhB5xY1ogQt7r/ITsUGPWs2KlRmnd
7TdsyMf7ma3rQTH/UcLuD7eOJnNF+UjWCXXwuJ9yTXQuOpzCQicyZsT4DyKBI+p43B8cKGlWV9Mf
8JZE83bMfJjxgpJdLvJONq6Z9aHAYv1EZSaDCrBoIHTdVO23NeYrxuzi2s1jFK5KzUzSVHgn4q4u
oiXyGSVXa2bpD1KsP+pg/aQBRVolojiFsIM3/ulQ3iwielF07ebVLTk9tSMyeXhpbrI65MGYI3u3
5fgH6i0+ATOH2OLBig++7tW81y1bcfzrUk7Z38MUjIaDtIdG/AeVRzxSkwxV3ilQBfvtiGZNxMoy
LQHICq8BmoRQzrjtZ0PtjUcScM7Po+EoAEURUBZmxLcq6Fuv486VeGfdZ4IUKAxfwqUlIGXlmoH/
bHBWWQ2JZMLzEXizDO6Q7sAd9vCK/cFOz2al4HdbTu/pGm+SKIXSm/2k8phQTXzjT2QugPAF/Zq5
SJ2SoJ18RVMezpsD5Eqx+6zlfh5vqcud+vDXtK6idh2d1vzcHi7AsfIPqTCff1+INnPpTDapnI15
yishjwyPQd+zsrlYOO4HiRffJuSpUELLx79hf500tOJE2OOEn71ocCeJtbVl0GH3mhc4hHzNVWC1
rP0fIPoHTQZpLGINpKvRuj6bXKFseC933imqEXQmfxpzQwPufyT4GjglLAQBSfOt7odiWH/UIPgE
25Mb1bvdWUueGNB0nvg0X/KzXNFb4L//SG2pl97cmFg4Fov9bZMURxEVHPHGZse328kk0tyKfafu
DS40lqyh3xVBa1eMcyeEau8JkhGibHSzKRVtU0M1Gg/wr+DQTrNdbAJv+wmw4bIGgSQHJNgggoj5
61WiNox/X43z1X6jYrVn2j4gLXL3FXeuwrEO4tS13GX6Zkv4TGYvTusaNVMbqN4ojRtQCApP886F
29shyn6KLFvrKn+tAB76DgQlXwQTHr8gqZgzRmGxRs2K1TiPCfhYZmxtN0UO8lyv8P6dHsQ/0sBd
qFkUm7SmXUdDr5DkH6v3nWxBjVn+XJAMmElukdYUM+SBqgrBaWoAC63pDkkZJWqrXoF0y423RmPC
9ASZgET0wlVFHenG3UVOl2L+PU+oIp1eI1RUVEyP4wNTQf5b5IEDiCPPkyNB6JDqgZYe40wLkoRa
5qxEp/7sCT5kBrBS46K4NVF86E5iYMZRPZySDU/dxlMgFkLs5fprVXbMucl3gkYRWsBbuVjjer2H
Il8Z9fmX9nkLhYTAGwD1TAiPMJhXHMAo1Uku87EG8GMLxW0VWdet9x2ga6XYM4RU+YKDxo5WoqY7
iuKbqYlHoBRBmVZmS8t1lm/tpeQafwG33GpJxeX6qlYxiAqrmzyA7sLrT0AAfURS8WliWtozXhtb
baNOPGvAsZYOC43wo3/Y3L6IJhVviMkg2G6n+WwPtFX+0kkIwdJMf7QzeUIKproQpMMAZT2q24va
BtHLJ1ELmYYusLJHSxBtJIxIcFqzPQZkOc5vjSnGVFs6YKgzbWjTJyM/UR74O4Pr+V+kYwf7zuCV
UD7HvOjXIRe+CS3UaWnHHe0qfOn++45AkgS26Rww+IhT8hI0drCb6VafZbBrFNL7aHVpVYuxa4Lo
OQa4rlZ1DJ+01ygLMEc1nI3U/hdQIWU0onJNVbi4NkYNSqO2KzomDJMMZMNcL5B/wwPfbpJKfGOY
oTQjb2eiGfQoyIRHJlEINX6oWNOST0Sowf0mdEDgzGk8TW9DuPYujpxHOLglizBJ1G8A1EJ4vKs7
Qs9gv0/vBSLpGIzbwLy0KtnfWLneOZ6frXU6Ij0OHP4CFTKsilTgAAOW0RS9eXrQBp7PtJxesobC
ERyLMREscU3O9wLQDMiwbZziDmeAUgFebYSzROAwrYX1XD6obVaEhWyI4ru5F/BMIvIT7QoVqDwE
kF0Wpip8XpLkBtwgmZvz7JOsSBXxTwHvpMuRqez9UJ0mbgj9+x5dEGLNrTgjw1fEN4xx35kCcA8S
oNqew4VXrtXJpit2fKmnuEWXd2PtuZ9eASSpQNQnUbmTIPK7Dlcl/63DUXkKxQ+KHSVOmX9oYfRm
UXPLYp42maQISmbLIs7nNTWUkBUUOKLGDsfaHdDUkxrWXeFaGoF8lhSHX8B3nkm395ktKCQ/As3Z
O9LZ+ko0NfzzcUnLnTHMCf+3t7YIfcqiXeL5iY9nbbFadB/eZvVWQZd0UzJQvHBsOmrxw/FUl9VU
4eFWG0MfZwk7lVx5LRWaUGQM5dFPMAcPwfWZB4hkiXyXXELwWsXm94inWHBG7tt517OoK1Qc2O0j
INEU5pAXliPhx/jQI6MwlwswV88dy6nDSCKRlLl89kLac+NgY1Aa1qj6GFxXa1mpdszymcWz2wzS
hHYMLF7LTzv5+WNT3Y2Fe++wFhDm28o8D1HnlALmmGN6FYEJpWNSDfUfbkBq6K2GS0yoTkR3SWyt
3pw/oN1cL6veorfXsKrMIM14CHb1LVWF9FBr4XdTVvKGxhrb0zxo0DuS+gvaz+vfqGTHRu+EO5aH
+w0hAQ5SITdh+wA5WexgA+Ougjmh3/BuuYSdnf0wtuVONNXdZkV8iLBmLGzg8CngTCbEbRmyGVzn
IneEMizyKFcN8/m//nx0P+IGRGLVhmJxf7HUf2W3W8Y7tSV1qPpKalCY0rYWzeuFfpjTb6PbsvTG
sad1mz8pwjpWk1Es3axRmJIloDs4KYtVj8X0KyoSuSEW7bcpD/UkJ4Wdt+ViaPv3oSbRHLbWGEOt
2dqsL2+9RIL/mCR0+pqAdLAOuVfN5H+nrIik+KKBkwXFYjxT6wTjYugZKqsyufU02UzZJYoexfPE
F2bsNvASedrVUKyPC3DMCfLpEE/afZcBa58TuS6TsQLI8X93A4t+WKY89l3lYS6eohs5TSItHtSA
w0+gB551ya8b5RapScBesKYyem55cfd2LVNxrA/uu4BT1FDHv6qdJNKmR2NJ5U422dYMNNNvMEif
eLOrnqQJ/EquqayP4Y1E0JU+NA95qMoh+msh6obk94r32HXUCTIl1Kv5XlYio3nJbl7pDFI7cASz
i+bAKz6WhE+F4ndRgnwiCOONdYTYPSkEfCykNC4R+LUIacc/2/r65NGcNZoGyqYtrXO4hFPjlg/o
YRNzcpBERt1xb4zafTIrLHsmPnRRd3ZeYaQnzp5MvVBaZdu950KGHqT15oyh+s3CSshqSzsdPacT
BsBJPfPPqFwQU3Ni10HMkj7uFSkPOj+rEMcdCOQVRfZdrFFVSra8vd9ySXaBzV8HJ0VdK/RC/C6z
UIoycn1R/wDuX2qj0nMG7dPE+FYcpOn4k4HHSEQI0PPYCk2nwvdHYpZuEXuSF6CYhd+zxqrdqDQv
1gUmWHRumQs2FVBF+0WC1sXNW9nBirGWo1AF/gbdtUhefHydddmxPdaUKmfGlFjqAWOxHfne7prG
Cd78j8xAb//OioxfJtLwnjXzkkCMXzw95KVHoPmk52jkvisSF5J4hAKIzF3RyabyWLYEgQ6j7hLM
ViUaCISit+aVYjyO3nk9fbNArfiLFBPJkBvzbF0EfFAaQh/Sp7TAwkpA2cT1H+PyefWs1Y/8zmwl
4i1S/X5ZXKB8M4L8v2KyL8CpQkbU2w5OHWAPgell/WVNsp0pTaIPDGClDYQgDMB0GHDfDuX8kBup
KC+wu9WvMYkB7E5gYs3sTyfHHj0kr0NVGn5VXEcCfUaLejbU2LFdZz5cTa/fA/9Blq2C9V5NrxVn
oVd8CxoMaXDek8RWB7SV3aoxAOBOmuX5cvfMehicRQxuW/FtkxT+uU5PVdzJIIJZPmcSI7qaFTKH
6Av0jMTt96LDlqi2LUdGmZ6Fang10UsBDvLUbCXK9ijv7w9rmaDHiuRu5qZ1MYhrdiFi84KzZhA5
VKMGtgKnMOPD45nFxYQdUHc0n45ohu8CEjHO76pOZTy+FLFZM1zinZVLAp950Jt/BM5MX3hLwe7y
a/QV5ZFupOGXq2w7XveysErsSXHdxAS7TnGHnYnrZQB0a3iKq03cB1NV58OLmulFvPdPEYtzPwyP
e8XQ8SlE368Cn5lxQzZkD1b0kwHKytkbiz/cLi3kKvD1Exsw13Yn2Y28VgF4Ww8x1ip7mBHInMUq
z3zQk1ipD8Bl/rSwwdfuUstvRuDVF0WXpDCfQLH1VwaORxu9o1ZSIOHDfj7gM5Zby+jqPlDzoy3y
HQzaTIydB+A6YF0syWlT3CI5CexaQQmkloYGovjPRfZ3ogvndaI6uwyWDLbEWENDBnpC4JygqI25
/YYsH5T9hyX7no6UXksC2JOElJYM8vGhboCPilCwoU6a48ryBaY/GGYSGmbFINyViJ2PM5eHM3qM
M2pAzzvoN4nZ80AuIhzbbhyMh9YiO0iM5WlvSJYlrCB8ZZHOu6g7KqditDihisJ2ByMwbbcqK0Uu
ixAY1IZ+CZhmBgokO5urVEDGAVu9VrcgWUL+/lqMBIJppXPnnXaubtMZCstWSIh8FOuYkhB+VrGq
r8vuzvtvtuw+b7YsrlDaup5sjuYA2VlNcHKbX0a/3X0G7Lx2/KyHn7h11K8+cHdYP28fyyPQNZjt
zpQz/hw3iY3GusXcc5X7eFUHsIp9EpEocgTBDYearSghCrRXx8nfWrHqxgTZVtUaUWbFP18hmFPp
9jmhuTGnPC+4vNI4K9NNlgPA0YRa8Oksz3861UpliMgLq3o2egBEjQvCMfKvs+H2SAdB6MP7VIXL
y7Um5j3xr+27gXA52fRSfjn0PNlfsRTZ6oqb9+UhXwnMPoHZbR5fulDqyHwrSVu3xkmek9pj0VT5
maXEAbt+pljHdUR9+XVf7vyfDEcOkG/75uhDe1WMZyb/8zqW8ScjMMDJrsJfNvdONONoUQl1t8+Q
Z3U5VzsN+Gl3hTvHDKNjUXTPfXvhdeDIAKpbhabuN/LZyNnq1K1cLKZtgDdjbBife+h8tBI0xmYg
HfQdWBD8yLRkvm/UzpzUCrFG8dRiiWncenuPsdjB/M1dnBWldXOZ1adYWvL4XCV6cpeXbNtOHUNT
Or9MRsD65ESScFDNrkqz+UkxqJXaBrtcsWy20MJy5MXRPa/N7SUU/rFiYZXXuXG3nzfbJKLfnTkK
KBAHRCmHiF5WlKfNSlUb6bQqbeDHBm0dV8CBIC3J/9imj6ldx2ZiCWVSskSb2pi3fV8DXlGpdyBV
YBNjOfF8ZY0dD+SzPay4zm3fFl7OWM9Ox5fCdPBiXP/3RdaDF22C/7BH+NhylMa4OP1c2uiw3xhd
s5OD3lrS7scfu1G8eCJ86StUcgd+vySLif2z76u/NOydEfqXNqMkqpiFd8yRhnnFukAHXYYAa7wi
MplSa35a3egr4/sdidIfh6q5Q9bJ6v9u5eG66jLMklecZB1myefXcLzcMZiaM1tp7JhGcV+DtrW8
X9GbSA/L2sn33/mK5wPzfgiWmY3vUAJ6itlFhhET8KilKq/WZRerrk8nr8a07vMYQBCfKuVosbUF
2tIaM9wc4Ylo0mhb3F4qHqQOyMc2anrerfoiqW5VRJH4JeGBNpLK3OaTlfI5holn6sXDnqgcmRay
g5E4V1omhfxZORQfmVoRVyZGzLGZtrn6Bz565xxK84rY38wA96xrcUhABDRUCOQxBgwCoEbmA+np
AjAELChMGgruafLdPaaedqjnUJsceZVEQBd58Lj2bwGpl6hFxLVDZgGGODAReZ23Fpmd6E34ykyo
47B6R4sH2Y9iB15LSx1IFrpdL4PQdfneKxsHhZ8IrYeGQ4KMHecEiDKbkrGm99HiqdlYAPLEMq3D
EFZUfoVm1RzWgs4RxjKJ5bsJ8oX6VI5M0inJzsdeWBSmBN1eEdFhHntQB5QYRCwuPFBOU8taV8OO
Ll6hVKV82RXCUB8SOk4v9sO7dofD3rco1NGrK5ig/nGH1oDMqedITe0TafQ1rVwgin/QcYmMHlx3
y09x+EDEntH504UQfwQJTl5XY2b9bEmGT3gKIqNpJRX5fK3xqqAnB+ZC6QgyKhbcsOmrKeDvAPXP
uBaC0W4WJHJwO9TgV8PY8Cke6rqbEgQPVvPv+2e/mKTi4KHKkG4FM9AKaPH9z5dQZrNQCMWTScOO
rk8TzbYYw3meJRkNnK8IuSTK7OXhQ2VMV4XRmcwW+DorA3qZxSjjbsnAnAKFuPhGm88kPGZbohwT
yEJ99Cg0y+kutVJ9G06vuMZxSBVYq+na0nqiVgHZFVfcImQtBH4sbDQ5f3KdO0mSUPmkBfEPp8Ie
exSk2wydf0igEOPz1hrjoXL1OytSaqhBxIyGRIgpaoySlp0d3DJmcjGBt9Nukq2k+ETw54uZHp4w
+YIeLFPvOxpR+cxhpSWNHm2TFT4SV9bLaXYi/Qdw4zFHFqCXy+QYPC3/8VPV+9/nmf8nJAPS8IGo
5z82U9+TD6VdJsE1MLacD7aL4MACOJstrqyzOrovcxomH2Ra/ub0Mxj1sK38k+tJmK4r+SXvmlxw
8deA37y9l5NCdr+dgajCtmX6q6ZPe9O8JHBz+OPcX0mYTu7VbHaweCpEvrXiGDUUTRfhOwnxH1qE
FTlR7/aLtsQ87zmzMyJs2tP5cKCNjbuHxtv+WtF3SWW435V2Y4TNUBFaPWyED/aUWCT/+UEVbqQH
6IV6bF8TpOOOeb0xLWySRfR10vody1iOgbSY8PwshVQZR9ZrfzfEkJSPjqYyFLYtJ1RmRQWLfhTb
f88mnCrlvJpeRQB3V5mJwX4gUDLcZT80ld8AAZx3wj/XgSWDfg0yCvkn9BiJcCVTIBOA/AfT4dRj
ZMXg3M/taD9zm6WzD0VYKG5EomjFnywqBPXq0G3FxOGvbp2ZGtyGOauTJrhfebNixyCk/Dytd2ps
zLixpOd8WN7aMFqMJGh7HVHUOd5nxrjfQx1mhs7ENO/q6qkEo/z2pwasnSCwcXkVs7paxsgiK9QV
Xe8NkEzzfsnRJPd0GzhspWknTxDbQjfghp0qL/Oi9zfvjkXHzydFMr36dBFg3pVRIaXY4iJeXKaf
9Ku92cxErpuJeCgC7S5R1fWPQ+9YUXwa/Kpi/IEUi8jN1WS+Tkg8zHXugl+apeHUr/0rFWGeovg/
1X9T5yz/2yZAVE3cm58gL/CkMyRIGBqGJyYInZ3JcB3icKSm9egVRu8ssZIC0/PfpwsWuFwZ5U4c
b2Ctl4XKBGESTt75TCsIcnVpgXXwkniflY+zvp5+gya0CCweA+rTzHpUR89lQmF8laV3nKKU90+D
Jhw4NDbQqf3rzyRjGhKiOl1lDUi14lvev05ZP4IfiInbYE7sdTBytrWysBUwaB3ivf1WVHdPZTnN
aOFnuvgQ/PNprh68ffP7Q7Z/qLDtUg4Cq/UB4N/yXiYE8X6xc1BJvTo0EBVJMzBBnDiSc0m/tRAg
ZnVTu5nqZD+BQYvQ7qunRQyJJ3hgb1vhV4Ax0ufVdbdxlo1cyySWdPD3yQVCDVUW0PZUv5QzYjFM
qe//9gdsqy9cTabW2PZ1ECh0NAmupmMXQ9BZcYQRcnjrVg3m4UrqN+7f8zwg/pFTzH23Asx3S3q6
TPexrGM+HmHsILwsH0drhIA1tbEzHq9UhrREwMcgP+AQ5oo4s+smHBIfMY9j7b5IoekCS7UPy6Pj
rGu9GiId8Dn06aV7YbpYWdVTBLCW31zcRCHJ5+uz4PqLkwpoIp5VZyXMzcQqPsslxvIJNkWKAQyd
q18MaqrcBhsPTJoY1hauTNQSLSC8mxu3a7sPVRoHyz08JMN/jpYTwyZ/yDcn8KkWGG8HbZxtS9VY
3JTrKrmaQ7co7xzx4Rwtf2TM3w5Crr3R5Gs1BYsxLJjAhM7KeJfeKgYEeBO8kiSernM/cC/5skUt
m1YdYnR6HpzV9J9rClay/hgMzSwty3lyKSuktFVlTAHa7WvPX5g3WsOwLU+LfJp4dItPK6XgkvdH
1XTh3mWqQbcAfdqKrD6xIEK3xx2LVbAx49K5xq7pvJU98hBZiRAO5S4vgZ00lYNJ5f8qWf+08Aud
NhhEM+NVD7k6LhlFRIXpJXsvibLxheHLiXfe0FKoxhnjyZkSRYrpzduoNqefCc7mLPpYTU9tQWNe
977TFVU3Ij7Wsx7YOwxKIxTw19TXJnN4BpcBtErXF5ErjEbb32i5FevuTVvXS9YwXyiVHSVcmVN1
3ii6LdgH3kwAKz4pYgIOXdyjXrBVfKPgtal32vh05mek4E6oM1hPsZKldTvEV10OXdsLPjulXT0u
T4VQe1ROlTVE34xRzLsiT9YyOnJkLC6ykWzLRTG8H76vRrQixvNCStxXfivDSRwWNKGKLbFNgoeo
uEpWsxL1YvBSIk66hPvd++PlopJfv8mnvqWbXJ+n+audimMaPjNJQ21cTB1rfcglI1LKqN79R9eg
lZlXsQL6CLIgHWIDtwZ+GTkaLgvhuJbFSTzUtNqgjPuNzIUHH18Xml+qaDSKFobMT9SD9XJVppW4
u8i5up7hRY3wSnohzPZEtK3cVM3+VklBeumnjLa85jBrebaaYu24qkNtuQvyIurvb+5O3wG5JhaK
xykdxNxQOYc1u8WAksirEhKaa5x7nmJlDVa0jOPlB2G+WRWxghQ3aUY6FWzwl+Mn/7yWd7NJMP3N
lI9wSD1cUv+bxE1sr44uNrnLkSqjJjaZ/VdOzF0I/EOwRhYh0JfV3xxHibHotjtfu3YzNstzj9ky
D9hP2U+/28TZGJ7sA2vJxDg3UE3vpoyZ8DG+OmB3U9fttPHQjoD5I3LwAjahWOwhz5jypS11NYv5
6k7bLazUpUSjGSSYObE8pUAW1/VxCuEaF6a49zjiyEqSaGcWY5M26lUMg9WuWKd9PVkApC6HMIZB
p9eSWEPbvlR01l3WGxvrpdCndiaKCpR9QLL8D3W44cNcKsxRqFecF432rwEJ5b6H3cRlpUPrNH+K
Go9uI9eQJ14UlgvWJ7j0TXtwwtqgCsu6hFidqldSgdp0LHPg9JjTjkeTiI5IDslAc8p3UzFCINez
W6d+ynGqyErQ5TeDa7cgx6JSsLWV9RkPtskdSsNmqdx8S0Tmaf2olk74Zmrzkg/jLl1pAyeJArnF
3yXnbZ4XEFPo3CIg5PM5DfAnzPriQctwTTrkzIQ+D6w8vYNEzhqR2Ir/drkotbH6QAy1DXArTvYo
kJYNJ9gd6WzG/KGhXi87PdIy4Q9XycpNmph+HCx4lNXM9j0jdurUMAc+VQ/07WvNjfhTlruSQvZp
AJdpv72Sydfln5MSnpwMHG0EgiR1t4UJSELIxVSK/EA7N/C090q7Pl32h1bLS+0BKFM/CRftdf/T
9GcL9z1S0mq8DT5FeMEPz6iRGuWk02oNNWG/tmDRkWXzlEzuwzKNfyi0XxuE+7CMNg1JNQUZRDnR
ViGz4qYW+ahzjRAW9ZGxTNRUPu74vSswsYILCgpZZb7bEJQqCbeoeOV7OO3LqxkLNZnnVfKiqVUw
g5mYeEcand+OlwUMT6w0vcQiMLm7XHb/CEIok/QyAvgyugbcHfuvPaKDPeuJSlSB+9IakQOUmE3O
xogXdrFiEZ55VemlLtHnLz/McoPHmOp0gVVthF962v/E7ckHpzIdD/wB2yYEetSumd3YkUMY60qP
+1Bx1qdMLY9u9Q0NUeHSe8PhCQjFCB2/2w4ifxtS9+e+Gv+0DEjivMl3Tech1JL1KUpV08PeO0sM
ytV0ItUR0EyeZH/8pYiYyxlJdrmnXzks+bGwGkDpP9l1zkXH2KU7nt0g+I8/1nolI6jISSvrrc8N
tlZASiFKA5TG0+7cOznBJKp+R64bjN0c8UCb03Oya96i4BzIfHZ7v0dSRRdz8MojrwDHkBoVMxW1
eFTjb1wUaDc7XwDlxS8bHYTtWAzNgMrGOqoBR51a406d+5PYxFBy3bT0UEamaVYpmgPdFM51xBzU
M7W4PxIWUoao3ANH5zAxnLnG07gIn+rWG34bLkHG/aMSO/1MwoiYUOf9t7ZrTr9kRdjiKBwDx+0t
h0LtGfI1k4LCaU7CEh/WEkGCIKyWGwCGLqlpt1G01dSssjWaB8guw/iBEI99GLJBWoHjl8bJl5M5
SWwMt9BUoOfOnigQ7D78XdaK+hEdQ7bsPKMJrQmlAhg01g6/murpyBJzhkMiDPdQoD8H29IYR7tP
RXvDy7zphQFjJoArB/+FKc4fcAOfvf5Mm6jiBQySgVT/rdtotvwCX9PGOAY/cWBnJNf1rivRf266
OnUcGdTWHpLXRVX2ta7uyMgvVcbxZgEWhDhca1y/tzhcE0aYdVHtxNzr8YZQ4LCrnqEMtzvj3NiY
wsTfNEzV+UpSzCIwTxSt40P+0jsKgZZOvVZHHbEQSK3OuLOkg4NOHXBaayI5lk3lJftEm4FV7sHR
27Sp3cOaqtJCV/BU4U7vTBz6gVSDiTMA6um83pJtt3GhxYVCmmh4/qjFgw3Ha9FwJ6TcYwWZMJPG
qvc1l9tgYZxClzWW+qi67AuVGEFuOFEqvYfG2qnbh2k4QDmaz1gK73qwN6w3d2NmukVQn7Tj42dI
K6NmPHjpsFt8kt4rZCLrbi7MAI8Rb92rnDqe5+Jguv5Z1GbrxeUP0vysaIspsdnO7YcgW65j2MAr
EZxaZF0BqROCKH71u+rZvP3viDQ7IAXJW9h1nXUlHXzrYqPgvphcIhcnIsyNYPjEtiBPqV+7IQSv
S0Cna5f2LzBlaMaY4K6YhUz5JY6ITImS1+FzdaBFKLD61J967xQq0D388mdFGohQXRnz8E1sZeOq
xzKUEI3amV+bumOt2xqM/9NbnhWO1cW39Hoo/2UDrdhyVEwnej70lmT0kNrTSeUgEHQJNQf/LDk0
DqGvXekq7u9pPJ4fJqpxIkKEkKrUGF8yhShjPFr+aMHT54JPRUZWzP+Mjq6j0YpQoE+Lb6v3WoLy
fl+i7AKPHiqww8wa5lxQX4mjYF0Owb1okJ8k823BS1cKOxnkfDUqGqRKA9ZG9uPgxqloEzKBYUnh
kRkjC7fLogonjBGjohQA3V2aioPwJrFh9d5bhSlGhQ1ezDzkdYgAIgThqBobW3/JQLoz3YT4iGb0
eF14KxXn1SEWr+xl8o7zpBcvBWB+oLbZ8vdhwkVcQ+lsoi4NmTFZbBPoHoPdJwhaCplBFirKuaRC
8/Dt3HiwAA2u9kZQ+fl3yntErhj9juh2AE8WQTG590Kxe5//Mo5K0U6JjqIHr1jr73SRhZdyntnN
YYKkT46E1163ql/USqxOAA/xrTr3//kjgQLT8YAeCig0IKsLz3QMSdK7f2OngS/ikqJiOjk0nVTM
CjUgQVRJ6pZPtY/lk3bMcQ3fN8QudfNVq0hBsFNr+Srl9cP0FP0vMOiQMtY6pQOJPMYWfDDrLC5R
u5TlCC16KrgmtAIIfHJPJtiXS32OKAr2yALC52KWQ4IK4x3NBLXo9Fz29cSYo1j13QknPNvSJWlS
jK/W4DcuuqaA3hMQPQMVyD0fQtmGjWJndamM1gbNXpy97KTBfx6LR2et2Yll2joTT8yDBMBLI03m
tfBGj2txmUYRYHHEWEZCsXYcIyFRzwmFwXoPQiG26ghelJuiC4EmVDUgLPb4YtJGf8bVQmOi/wha
sptQ61SZttMolcRwPsyLp0MZa3HJZuHOXlrmYS8rzzyV5Hvn1kKS2UImkw5iG9aAr0dn0megZqSx
uuMb9D7tESN+8TtEbo8353iyvbMW3SxthCgSTVGEsaihafxlnFpk6H8B1BpFnLnghnWuqgSOHIOz
fED/f44HEGWdKx+G1Y2fbC06UiOCqYZnS6Wh+htqmV3poPOMcIvjNY9wwQvhicxLz1iO3DD689eb
EfB6dT3VgsbKcnq+JM1LO2SikKnZsFA9rpSn9ZICc19h4ur/D4qULRsRPRlv3uHr+S2fzcIj89K4
jikHtpY2Khy38DqCw7GuLybq6yG1L8yiaOv+/MFUQrFXec55Mizj9h2z+5zKWWlJFe2rZ5b4Y+Gg
cMQu2P4AwfkBFS4ayIoTgwuV6RSdtZLzUHaOfxpBtm6oithjNUW8S+y7LLX3sff73glQQxOQhwVm
E85GOAyUW6kg55amdtdvnKmbDhhpGfTz4raFn0CRU0zDHU7/OpG+z0gi2lLzZpTldHTDg8oK8EfC
Ft2Q0wtqYyED3b7PiWT0sfxMKgvbz9dvc1/QGnt2gEwJLSpR/elBKk8BHjGYVkPAj6/hABauI79T
ymUP+1Z0gX9dAlR1qz0Bs0OlWYAVmeAsluEN0pcL1ATt2QhILKufGi5paQSXJVDXfaxkapB0HGn8
jk4NA7GrqEge6TMUSsCbw79xAdqIePGWXbDR+Quuq6e9rDyyItBpxnl4TAbH+9jLFWPtbjVqkg5V
BY10pElt2M9iB83FT4HBpETZrznjgpbz4nFYJ5Of8fjOr6E2yHGvcIg6SwT+Z/6Qn9ZIx9ixK6VT
SPmfMVzvKhw7NKK4PC3e+UqpY+J6VGPZ3tI3xCXFXtNGxzXF72WYKZfCN1yqhkORcDQuenWIzqYA
3Fo/8hAbhbLsJ4k8lpPWcwkSJB/RIy6kyM/l9h0kFN1oYZDBgc6SBxRb22VnPPjCEn8ZXbqHahi2
2gSHMvoEze4BfwMD6xCSFbanfx+KpydaBGCGYwhJaRJaYBYGh/bwlPeBcHPv+tmYp48lq8UZILus
KGOGozuehqqDwjpiV1jarlPY4qpBb/6vCcgpxhpvHeyTCHAqeG2xCfKK7MEamfIkrvSUO1K1C5Hd
/dCwC5c+WQxE3H/Azyis5c6vRwxVJXYGN5BUeuemL6lhyFMf+6iKQ2mKMiSCt59moX49imSSehtn
y/rxkYh6Aja1/M3no3dKH50hOg9byTp6VTdT4hY+DJpRiCJL9u87xkvBJ18Sj+FZHLxRPnLcbphE
2O5G8KvdnFet47zgPpQIOJvaPA3LAD80xtUOBqPiBSz0k9fgGh9jrd0h5fAQ1nMiSWsK4+P8JD48
Rz4Dv9hdvHxjOf6eWw2zQPzhmA/H8e2QeD989hk8l/LXZ0nmePeuDo4hydgxLVV1GpDpyDn91lni
HDTyMM8zUuf2dBlO8T1Pe3Q9jnEnRjm+w1EsivMNPkDu3cD3hOJIzwxyS1o9/RUSBXfGBEUKDQUy
Czc5gRfWG30TGAAQwP7Icmq6NYdLBOsAuh6sCc6huI+vxhj4I55WdFJukgBuLIH6pTZbhQKEG0hd
rUUn252OSu/fVFwQuzKEmFBz+uNGDxjAachHGynofa5M9wYZM0wY7hywQCVBpWWE9R8ZWi9YdEcx
LayRc2mJVQMIyt2CgM4AsPRHpTUYvNsKYKPtuDKXJVxRCYeJK0TBLAUDz+S6b+bPC17Ex9RuBVRp
7xfXDq7swcGHV8vLUQ8otDHPs2MKsfsUWMDkAChp3ZlYqEWqwuxO7uTJLocyj6YePLZ+L2zrXK4K
KKHkTONvflDAH1d+sMTSrbBoBLXmDAEiAxtLKBMRgl6soi0Pbp/fZHcN59ET1MhSVp8rdxvAKKAr
s3+ikHP7FGSEmW5pCUqLa725t3NyG9kE5dzE5SOEFX5lVQDimi5sSVZPUPHbfL1x14hHhTqcbVZo
Pu/pgIRRehipNvip8eHwl9btpRpR8pj8jI8Xtri7BF/Lv8ol3T12JEY9MCo26wFHWARflRZsF3G5
C7UTX6/wrJN+jCpN53As7sf6OcQpAhdGfKSbKFJLRH6tJJsL7WiFZungo/k3hNLMFtTNwDGWNgsv
ImSGbVGHir56HjFl/S2Kt/ILWAP7TXjBFf2hL09bued+KaRbHNsqgkW6266n0C7bDxMI8/ngB1+K
Rq3v8EEJlYIv8qOqTqHX/jpo/cOjfmb1ZVAQvf0sZA3IXh6IPTdtE4d98U8FpJbxQW+hlenybCwR
d0/fN463YcnwZrerGkSAI49a3YEvwlmBPfloeijoPl53pxaR83w1YVBORMQOmMtR3KZc5JG1019F
XBhU1ymV4K9riCPp2T8qN4RDuYf97smL82fg1vHCXrgnNdupyQPFNBEliuA+L4evdAW433fZGCpL
ahNtIGAZ+o9ubzV1V5dZ5HxBSAGKcdwKQshp0JVk9bdIY2lfK5FlIrKZ53j8d7AQ919HJAzPOtn0
rP2gbDIRy/aC9wJ+s935M2Y+zkwT1OzHREaO/08inUNlozrsXijzqByBE9Ia+lw7g9RMmZlFB8Z4
9dpFfM/WQnI/LUVApx+Si5pxlLLyFT7zbyIGywsTK61cnUUSQiqbUVgNlODn2kdQVU28FNDLaXJf
3eFkj4PWM/V9Evl2jRBxI6GoYOvWcaCPa+aXTp5XYThsKJwGziPUDdXjuHzA5B8Aej8ieeXeABtg
rLIuwBg1+uoqmdtGCo+v9/UZ57K+RdmkPso9azXq285kD4mOMxB+SJyyyRVkO5EENXUIAPes/avy
vkT4Or+3aRoXlf3Q3SRhvRcfGocwLETyhNQss6m3FtQp7v8OFwLixTU+mmhPLS4jK86XwWwPqYFq
6auaCNOkMdjT9HUxWondIA7HaYiUkXZgNSQhGRo5WvfBIZAwy8Ki/Z/5f1SB4TKKc8obfYcqKmG8
9w/7wjIaB/hDA/rOWZ1R0HO1JwZOQ0L+gdO1ENKxpDiVNtmhD6oBa+84M5YvgyDZluRxgwVosDj6
Q6uS49DCwUM1DzGrpyaMh5Dmw+W+rWmQ9wKzpP0sFBuPxEIZvCZllE7v5DbDCcWQOfylYNizq29B
Q1XgEfn3Xz2VHW5n0boom1xxAU5cPo8yVZFJYbkWtIeO2VSvLyU3T3dzC/5G2qkKu7vrBfzCa+Ke
Am4Xp2CLw0L1WuNTDmMoNfq/16/gugATN09C3Xzt9dGnvhdrfFys4wvbcpx7xv8zffUlPpetCIkC
0oLSMUlWGUT+cal7UQdgVIwg9QgBQWxcSUXr3BrpuZ693JFi80xp/U9K8jSIoFLVXotMsyddYS7m
VKrThe5i9PnAZr3t+iyrAdz6i1Taxci0DH9OsLpu5lQVi5QaLDxXjJUqX+9dJa65NO+LNoZZYYN/
lrjiVpgEOPgNtuuFi9qhNVDIdTIahC1HqwAu7WBNPGTkKomv5Gkv6eiwQFx4ejw8pUlV0NKPaoHN
OmZlj0rkeQFDMewwTIR9cg9IkrvE88lGIdvJARe4Cl+1tHujVnQ1ktl68DL0a6TyEKIWcJhoyWuQ
OLQwFREG7JL7PWTuC6IngeG7fB8XAAmbi/xO97SVgzupEAmUA+QkHzC2/PwjekME2v/kv5JDHQe3
U8jeGuR3EqDtAO7+wDaVfgAXUxCmeuidUfCijYsN+aTFwsqrMkwDwfZOWeSJrg3hnf6baveqsm2O
R1o7a+TXgdIVPiGCPndOEXQkpo3Fe/E2Hej1N2xCsv79JNJd29x8PAGAFu99OcEdrSngtpkVZIGR
3DFTcb8tA141ijS1AiZ5NebthlhaS2PcUWmTTAbzkjlnViiK6uvezaJKQBiqc+5Ud49wqZi1WXig
cbU3OLeO+t8wC8SCZDB1hPCjjK5vQXTRo8gm0mwA5QOoZnkdzqod5n8NxVVGUHcQwZcHLLl5/bvL
ohWDW9KtWMzmgpbXr49vBDEHHzKU5ymy5UZcqbHe9ZchCr1XKgS1+Hd4Do/M6ET4W6yQ/w9QxmHY
+ypnldIE0ZBQoxou/YnAjsX85yHPeDYcT+MYm3wK69Hl3oX4nr4/zZibOHncPIN8Xsx8OaEgOjn7
D4u4ShAoSL40yS7Il6mNbAiIa98M+OJS0jjUun4j9ai3I08noE4awbhTqwbryn43CZjH00elA6yd
FKKzhydKWE6PjZ/yPSKE1aFCnZgwcm847OkPMY829xpYl5Ed0knrU2fugvYRhTymCbhcisdthmlY
s5gFmutXKDvaypkPsEgLnprRlDFhRBz2NWrHIXp5s+X5wbbP8eDXkTvbUi8ZDrmYWBK+SVVF85uT
yMWkRpIq71cKKausdmQzU1vUicGzwQoHnzy3FAkZo+sNdqWm1inWBNXWoRlhzi89WWqfAf47qPFO
MPEtyeAB4OjOIRMxpvpyd9dcgfqqbhqesCrRB9MVEi7qrwHr9WZck7B55JBu6WKrv3VDyhRY0dbi
mSzGZCvtQ8BQf5stwAi+2oixv1cSNyJWmgzROualxMqFt8AczWjDgmv1F/73cEwy96oFLbGj/PLp
q5UVdjI6jgFsKBixQx01tVqPuBC0hntg6+yXSSTd64qgIULWxnENa6dNJgHK22XMkNolSygacmUR
9AArYLn+hBkcmHAlOszDAa9nOrBR5IBvwb7TLe4kzCVCCj7oIITyp8SJmj6EhDcU4Tqv21sB3lfH
JaTfFrpqdJAWPuSpalqYLIjYO/vGk7TAbSs4ZZxVCcqwLrBRYF8OPfnizx2wKvNpELS3JOhsA3CC
HayyEn/HcJ84bcBhhlO2exhMqrZDojuza4MxZ5rcJ3r2eRzH3K1Hye1n7vFYQS8LyQOI8JexWUqy
uASaZQphLQqWAZZWYH98sxY2tIaGkKlVX3SvGl2+X+F8gWVkajOFyD66owpcTI95wIBK4t0XEVuS
Knla3fY9vPxOUe+HSIta7/bnYNg+f8POMqGy+BYTNfg4nAQHAtvJqlomNRm2mN41GLL4R8bWREjj
yiMggRwArzCXQyaXtDGYzTsPb4lpUGI/vVyRrrJR8tQaOqLCtdL7Yu+WS5pnF8HDQdAtan2FjQre
Og98zhEpXWE4DwbMseLELEMxz64SL5tHOjkxihG9dGP2Ww4Bml4wuo6riLO2kPJsuIZ4Nh9i356b
HUPBjt1HbQxJ4xBSM0014lQpgzupppMR1xw/9dc3FBsY2AkIDdVLZx0FFS0sp/X4zrmpJFM8ccOJ
xsCbARnFIyfrQKLDfzsulT0MPEvBEHWKJtWpMWCXlMwUhfbvqHigTkeGZKS1gj8wXKWc0ABnVPdA
otICeOrUMCz0ETp47fIuLWZthF6u2Ml/1hcArPApRQ+cFzVbndEU2y6023gVHsxTF0xzpyklO+1Q
oYZS8EZooDSn1epxc5+x6QG0Qs5+L+ehAMs8yBiMhji8P2adMd0dN2DPS3Xz/EpkOXJeVugjXO4o
wvBk009AehIPRumbbkQmXP+bOLbpct6cyPD8yQBHvQbeZu593t8LM4J53J5C1obW+5BMQHhA/jr4
KDDU4SzQmNih3N8WL40VhqXel7tK1OwWEB0CRHZqQYxz2JV1Wf4WVkdHNlZ+6zeEHsJzukc2ytY0
VWBps3LSihhYqj0SFMAhGGnepPBZcQ06yebiX1KYH4FMqikfBskZkjE7mCdZ7cXS5JIRnTTxZWG/
gaEHpCG5B4G9L9+K1plrdVcg6utRvl/liKVdOSrgRrAKDVhRdDYEE1QyIDpHlXAvhLphXk5068jZ
hhr+pbNbEJ32IMM6AOpV2hy45pR+f0DfoiIy5ILFj/Kc/pXGUrd68NNS3A58J4/zCn5/dGUvPDUY
nTEGPlWkwggLKFIUlXM7QOnotYBzzeSueT860ai29ZhetiONJeYjlJEdVTyH1oAgCJzUHi1wlJ1f
gAYxChXYmoEYrPtgpn6MbJMk3Wi43UIHP8Wu8yaU2SQ+yxVHh4LBoKJllQIW26CCP0ABmd4OX7Z4
lLpFV+vHrt9OUiFiW7l9za6YaLe7hpsBerl3CpH4XtFY2YfH9HDHquHull8qe97UkRRQOhbHEJnz
sgugrB714aAq3wPOrOXdQpzAWGOa0SvljDdVWQZAfBn4pNJAOo/DMccCiWTyvGAN4XXp6pFPYHdX
VG+clEApN1yiYwxl2E8P/gHZfMG3Ide+ItefR67p/j4jIOkM67sZppoI2AUMEw6VsHbpG/khPMTP
HuCdBDjb1bL/UQ3MOHRE7hJZs4JQ5v/NvZVBo+E5YSNjeNvP1p95vjA0Ob5t95ipW3dykC9Vc1RR
Pb3oiAA0JVq65pPryWf9vdLYOF/oFS8hOTBi2lran0v2cnbE975TLSQLzobWsXzMzerGdlxnlHsU
yWYFzeqAv/kdJWP59bMAyM6TjwE7zzn/SbvFkZxrmSDUcwTU5YaYk63fK6kR8yomG/yzew5P17RT
4LlPzF3VCc72ugm2K4Xy6Ql/oxBwV1IP0zcHw4NGvGFh/ZhspN5WKaxsoHErVSH/JKenqx5xO9RL
1MKfj8O8Br1uTmf9lvKZgKgDnJ5QSQsLJRq3rUS1dbC5hPKe7Xf9zQvLQRzWIxpoOg3erNhEcd6q
MOBcNTI1zy05ZlRA7cFDheaDF/sRggZUf+fm9ahWFkAUiL6fMc39pmSpQZ7IGAcU+xieSz7ypCxs
BiA3QNxnagCYzcmTXEwRTPxNaGGehVoFSgsZYie8tYjVrXp4wQtyQWMTsRMn1zLmPZthEppqz0G+
4ehdcCAwwbq4Rp7+FibWr33PKL0wZo4VeGcGWIerSzCumfjMVpdwGI8273NGecOM5kuY/TaWBHoH
ikyeOJGK5EBP1t28Kqg8802XEYJNrz6Q7SptNJUWQwXgoVQb463NxW/2nms/m8cbXEk4FtsJbN2S
joekNhW4lbFfCoXSuPoZXIRsYbptOPbvmwuvWkhHG8trvacGcjqxqeCpDrpNRjqaYKX39j8YtWV+
fgGHp25jAdfb6uquGhXktUVdXn1r8zK85OP+28BOZz1q2qU+SWlrW6HcryVGzXav5Z5QPjSE+Pp4
ucaAr9o8I4GOcALipTJo6IfkKnw+1hH0LtH3LhFHxScqpesu/6oYQ32OWOzZiTOQa1t07p2XNnje
S4QrB8bWFuPvT2kXslAY5mmugcYZS9GgeaTgDhJVR00JIzZWbCpSbjSiR0unpIJsIYAkfa7ySSBj
TGjO6Z/plPlx5JAp69deeTfVB8ncPQOo4mM/9cRY7A60lkdHMSietduC/acnteMNZmFxFG88Tcr5
uwQaO7naz/x/UP5Wy9vwRvyT1u6zQXKdh9JP0egLOSezi5cxp69YsrEUxe2s1x7FTHkQLU2zRLcB
NiPnhwiYOmBxcpI5yy35zjoSQlhUbE/LypKhLfrizgQ5i/VQw36jYWl3NEnX2V+BgcxROlAyro/0
0eGZSWaLue/TRpn86B/5Q/KrMO5CzW6WRar0zqPSWr1ubM7PTSFBQZgHMVtCvT4WpDHv/5s11GQC
iDCRRh0sNwgee6ugWHF2XF+qVbp3HVV/nnFF7TBV8lTN2YIE2EnLKVGBvVrx1IbJcUE80WALTaWW
JjAEH71PI4OwrQRRnL+X2JSrQ7FwZI1OVmjKVZvM5rUoAdWgluLomrFo4R+OrNMhWj83SVtXlQ4i
5CuX30bhEhdCw6H589+olVgTPJBqxWpH1ssL0eAucH4EhV2rHALhvDDgu+S5T45OhQwJMDu8cyKn
W0g9PDMCk028ZUH9isEknkyfJsfCpehvPKUFJINJJ4yvkEsYLytq6sQ/k+35JIuTDwf+ftlILxW7
yPjF60z1SsX5s0Uw1mXKAfbgCY0S0mb2Xl3Mw25zylOF1Ata50PjKuUadEQqWZI/QuvxB1JleV3B
NZXn4MoA4eoS0vHw3zwPyFNB5WJWIQCnJCAVV+yxxIUwymd9aWIRl8K4w4Q3qO4UF2gksSgoLyz9
qMdc0mNQ7E+wJ3uXwmQJlmBV1z5jZM0oDHB1fDydlH0mZiT+R1Yjdwx69afB7G/pi+AMBnqNEBdV
aWHtENjVeLJYKljA7sNjROy4Je9eMJZqeaIQKNuFsrmv0wWBq6sQgSHlGZd1G6F4BYpf+0arVuAj
ywxtt+oe+OWUGdgyqbSTXEVT0zzD2nokI1fKGYCcM23YWXuebvLGSIA1SiVKVLaY3wLrVh70fVZv
MB09LipV1kfbloPrVrDd42SlRUvY6m3fgMYae03llIXpEaSEdY7yVlJUnm7b2rjmI7ZqpHDBfMH2
+lI+1YDXBJ5wGRCec9zreWxbcxOQioIJLbNv0ZdzPXYV/89p5dP+Vs0RLFyGKmEDD6kK19afJDq8
xoCSL4jissucZDVoUYg44uIoBfz8rZLVA5ALTOWU4SUzszMvajbOBfyoswRRaEXNwDSCru7RJxhC
fTFoWITXyeNQ17xjy/67i0IU94VAEST/xUNS918Fk80h5EPA33qHGhKew+2AXemlbo68cPmm64rN
Aui4TF4TEkaDjdHS/XhEnEX4TlHhLdNb4EzUw9sezVuervYyBsARzX99tIaI7DEBo3HslPvngg7m
0gtUHpyOfRk+vkOFXyxXfJ9/010weDhTw0KlUnoLlUombxXBvWJfZ3kRq0Mv9scmfj5sVYp0dELX
yT73VMCa0TcAC+LV7k2B2qI3y+p0hJfeoKg5dC6PkGb7IAQ6EO3NRbPSYGiO/dp2QvlnW4jhc9As
jM/1m1O04bFJK6vQbmJHx/l7hrg4QGQiU/IJPsONhgtj665eqlj4BCwncfdphmm61XHnLfQEf00K
wgRUUBW49DKKB448lm5S0UASkTMIEjagPu3Y7/jsfEfIusWSLHzHxTSqDAFDtYef2h19f8PuQfzg
0YFGEAl1z3PqXAbM0gxSQSwXtQYgCmBGOWMHZvEz1EcQ/CdUzDNWvFNebQRiUs4Re6QvAy0ZWNuO
IxeuCE3N/KnZ5ZGbAUvI2mcTSAoTSCLVsILfraYCkZY4yMclQhVizdbsqYri/zPF5ZcpVIOsYmu7
wrHZY8PYW9YkU/FXoZplzgfw61ozFi6hImamL3HMpQOv1f0ZKhqUGKNxfg7lUGtdeVF5ipQCWg/v
TxUMjiEBsvxHMz2Ov5Io3ATbekPxjuoJ+IQa2Hr98nyB7fp4/SnrFs0AchcL/cei1khFOOEbIYht
djHBMvvGppFWmxLSsMUmnDg7OyosxQxsLJBsY0eIZlSZdWdSDVxIicTV1Ub0gHK4jdizJGTqDnlo
dJ4Nz/rbjG9tXvwmmiFLjUkFdNqY18ZO4uoIQ8Sa1eE8ZJne/c5+Cc5V+6nCYbiv/G4hDHaU8P3V
f9GMzY5GOL9pIdvw77erH5eQ9sCTTUmJuhPWJsE85kadi7drCNfw32CEd/f0PMrUO2sI0+sHkO3D
Aab0ctlvvde5etVRKL4B32xsLYxon4dZ/UPiA2uxktCqVy+Q9zXK757EDPnX+rhh0w9GYCB+znxN
2kfENTOeZxAYavZwzKnSAFk4RBFnI+Y7RUocuTklZiTIxnQ/bh1Ajis+WH5UY1HiVmqnIccG+wz0
KslDTNBE/D2W3MAnZ6aKyI76MevNd2rqQOmTrm/pYrN+1ougibJ7kGZN8XBlIuvBzDnFe7h0Pxck
WfNbx+sa49nNlfXBtuWG7f6K9arnR/GhyBvveejz5hysYSYwGMWO9X/YWhi6KyXvx+Podc4SA6Wl
+Tv3syHJnHfAh1ZF+DkorutOzrsJfzY9i5fsvd4Vlex+rb+jnOcFX2S01roVd3KTteew7YiQxdKg
ChRQqBR5PmE/XKAU7Ey/Bhk3GpzOgeuB/yvHhW39tUj3QhCAHNQkgIVELY9sv/PEjPqeeQbVjClQ
FTweydoGMiBTp01IBMllho15z4Zgcbby8pZizMGcq38zUQFZZ2uTZr9KFJrLNqe3SKXJwDfYPLmF
+WBWlf9pdDelkt0xl++88ZWxvgn8n6p4uNaXa2J0mlMxf/eb6rlBMVDHKachzERTWm5vWIf8of94
P64pOB7QtttmSmUUycmg3u75a8YboJAAQVl4cLJLK/Jcace0/ArI1qTZHGgn9t/7qhUJL0lnUcPo
N+B63hU67SkcM5ldPePN2iF+cwXad8unvi7EsB7ilWNiFa3mQPfOsaD5lgl/6+zPxmpdlSsOobeJ
ptQzbmR2SfUatPUOmb5enHzYPzaK1+FSxCyMeXfeL/G4U50K1ZJlcr2mGaI8HsZ3zSLddjaNSAjq
2RKwGVdq7TFQ1z/Au9Xr2czACzummSC5J1bjAobXiooloJAry7xd6jSnx7kV9yXwk3szWs5705Oq
fyGGiXMCcu83RVqPNlI2IbFlUQw8zBbRp3HQBGlREGia6ooBCaTg80vFViskyCJ7DJidt23oy4kU
rBkBclGSQI4tG2e+2XReuYg+lG1mko+L3rKEi2DqYmMor5Y02ut2OTI2D+GLfEL6enS99WWtuG1+
Dbr5wNPkcDqLkD0/kINRHw3pGeU10ENcXonkQbGvoi4pLtP/tmw2qU+RLQ7yyonR2sy/Itxn3ttZ
6ZbZsee2i5i5yccvbg5CGgY+UHFkP2J/v8Ip3Ip4Cv93g/YTuuLHNKZnURzbpKrLAHHF9/Z2e62w
wm5Yj9/c7qAeoYI24BvfI1YtgGH5Ac/ZC3fqNa2F4eCFb0CCYgYjIFgNgujLRSFvmLmH+DuqvdrH
brfux4D8bs7pPpdDQC6zjmpEnIccwbithNLrOW3HZZf0P5Mwl1UvgPrQW6a+RejE2GrcuJe21qKt
KDK6CF/zmdKd/L50zjOLoxoRwKPLUM/8zcdXgMAg9O3/8EcuRFaRwgCfbdO2TkdDHfQ+ODeymUbx
CXAfXxrBKAuLJhfKKrTlj6Y3H1Me2UW5ge5fLWbbwhXy7Ax6zJHWsmunGCwXJVr8X/p4KMWX08XB
V13dkYjluEYT18DnHnni3/oxpNNt7v2yllGra/hFt6vyGpjiPNY52lBfik3VkMNNxsZueWj2xzby
Yr0scHZh6PX+ANCWM2yEjJMO20wlUzzscNtAVQljIIKgA28P0Zxy5DZeo6+XmaOwv8NEptBwTmhQ
Pfq4UiBz/hsPoFuwUeZYNIOdPuymmFLBxHkwUXeuE4AGoa3v+r+tKwZ6yk81Bn/Skkh0oNfCNyey
5ygi8TSQh8kjNFJEF8hMmFnA83asy5NS5n1LmilSoqa983aD+bA8FahDdICjhEtytUS/OF5Y0OVI
ANvrqtquC2opdjsqhFKFFYbsu7954GfXUIpQjIa9Gld3pCFGNBK8o6SaGV383LREGVGyLL/F8OdD
xH7OaAdHjkAzyeoo05tGE1feHJlJxQ8OsapwQTYW4Z32MRUAn/C1G0vBcv79vo6UXGLOUB6kWZYD
NWXbPQXFF7sFeWjvkYFViP5WDZTeJLo8EciDsfpRVcCc3Ezbux4CN6A0vtXDNgMXQihsdpQBWNOu
j4LleFNO4mIdXChWdgqRLlNhe814Qmvw74dWyg+nq468EcxEYl4AdY2xAfEhGyAw52oG/xfC6KOn
yvSGun6E+1rUJUAEJ5xREhwIj6mA9xl3thVyufzpOb9oCoNakc45vD/5t7c5cE/JbQqnxc8FQSbp
d3tjqA1BCT5kCS/C/3ADPmIkgl2sGo3opk2EyRY2T8y9unJBL1Po9dB/tkOuPcH01F0VWK2HraKJ
QLtRw5N/fJcprxgxiNdFT4lN1LJBu23Tprm3tK0z55QrC5KaXXVjfr57B7CLHB6rYmhMl+w66Z3Z
ux2c4hzri5cWYQbgZCdOAnN9uIRBYz+EAxfgPhebDCyELOYLIqC9PVm4WsMvAptHzWraKJjaKOgH
w94RjU84MWlCxTfpAwi6j+tghUpLNazB/C0F5g0HxArbdnvLTUWTtaTUWFIUzUZCsu+to6jmx9HW
Y9OjVR0SBrGunoK2TCK+AHbPZAfUnjBjgIo5hCHo8pJwk9qk3gFyWXbbv1DUPV52Wt9+8O7WhQAU
DvFpQn/vl1HgaToL+BYzTXMiVYvjuks0WXOlVnOWjbiNFDJ045Avy/TQd0lLocpySY1Vn3TwW5f1
7qPqP0nrOWZuefAzNvG5MToHiHy+tcH+5zJhkZ474J23I2H9diEghgc1TULuzld915kRHdGbO5+1
aYyGXqar5tzQTZ5IfXL201OgWnpPb3CkAXNnto+rKAc0IgKrLc7P5kTsxMwZ6Av/hy+LdqU02urG
J8P19BmeMc6my1ef8oW5y2y4ML/2meld3GtkjWps779Jh0Y1qnzWPl3oLpQDzM3P8sHUOCeIMNJU
SwDCCOO4hBie8KRQoCdCOEJ7QT7BdxSU1XLj+lSjxEjx2XFjnEHh4zlkTgMPAugn9qM1oYVsJqh/
LIxXtFUBT+t92fxQkgY0PfbHHgiXd1q2AVCyu6g5g6W729Oowa+QCODzIQfyoTl+oLFu/Xe/g8zL
kkd5kLkwDtlAF/gRftAqTYz6LyaMRPCbzkgCG6kciLhpWneZ087ERlVayWJAwqNUrRIHxNTcIaa1
CEaKWfX/vc7XeXwE22jaD3kKhyIdfdtAZcXvTZ07zRppoPyTnTwW6ORqV1R/OxkWz/wMCGS6pyk/
Va/IDMn5W/Wqd/xHc9QDgJ57tC8n/dJw8fofDnWK2aez8h3D0aXP2ey1lJo6eQgRq/O8lgmo4YHs
4W0OJTS5J/eBXk0xG9PzzR+Dv4q3nBKABeLgJOwE9EoRYuhbroMVLmwIqoIB0UuYoAzsQ4MtN8zt
L3yjvJc4qpOy1jstDSi0mbcSAJ1BR6SeF/FoStZeC3G8I9HJoY3/kfVs3CnFjKwOqE51qJjqcBcA
ep3Ee17q9ADOqRpeRbWpJt5ZNpgreu22lZfJ3zGpMhnob7woRutfN1iTLmSGz9I0NkKDsLHHhPzp
txMRWl76IA7KcIRNNu+H7M1JZr9KTwfwr2rIstlK+QRp/BGJpCdPDVuBLK8Cy4h1pOWwLfdOy9jc
daTA/2IeFOM0CvDfPI8w02vaxBL6lOG/bHs7C0cL6xiWlbB/FJpzy1ToL72Qz0vm3yNLq4g3Q0u2
iKWVOWyR/JaZfxwonnaRrqDWTzQnvg5kFiurS694oDldimvmh1mkRlmIsV3E3OFBsCYahMPo9orD
rQQIyML2OvmRERPM++JMciMjB509resbdrwbtqbWT62SU+NovGy0lXsSHWoQR7chmKOQlCtNDzyo
3lYBLkWwJgGs57zl9apSU16XboH+8Ko/MlRhTAYPq6Gbi3xhQIyaMT8jM2YFyd7bqntIp1CKQePk
8edmyeGOPmAXi1/sWbZ1t8Y5w/6G7FixhWrX1rou2Bcqtvg3DQyf9Q23fn5jYOuGX7+rQpdD0s7a
IKB+p78ETwpbgwHZlmnpO1qyTXItIC55fTa71Grt4wxStKj+mBH9dvCuTCs0vVChqrDF7hN9cwwI
83xM9C1e9UUEPP+Sqzx9WkxbkX6WK55p4rETpBLY6ZKvO8wXvjO87zUfv08STQ+oUWsmZbr05aaN
bXJsCn2vINT42gfvq3AgiD9U549LZWUJbuDB9jlhNiEmy6UuqRFf+xldXCPeyf895p5705HBExW0
aYyiQHvqWxZZRRl5HXCAHtGoGPRe8FHik97EW+SM7BzXpD3uCszXw+jtE0/mBtrlaI2+aeDCLpfY
e34hSMC9mS64K3TuEialcZ+OVJI0VtktWbtEyYZ0OgSbLbOMLz19pZnJVWjZH4RdGvzc7JKYdNd2
RJyNuXdFYFEa5fS9gPgscyGN9y4GH56TQn0GCIPzXyq3OQh1furbZSvkqR8XjywHj6rM+hfCH2mF
CxEEHt0PBy2Lhw0Gyf4LJiX3h5UnLkO1imfci6bLKKxBycibyeNDmLQRLJoKd7TsqhZFo0psac6h
mA5JmODn7gs69K5W4otlA+ZZGNBQ936WJDdwU8caoGq291HK3woS5w1aO7f80eobTnofGTcKTFEK
rhDdTR7wlAYqeMeDXH3mNg+/Ax25tyqursf3lvz6MMDJKqXCWl1eke5/wnpqs7yj1UpWlSUpvaY/
XNWIZ3CGiMLPJf7ZgExIEwGHNQaNDSedXclZCt4SVn/eLFbxIoo+BYhm5VJP/RQK8bHrGvFf+Cww
PRcsvyDTpBipHRtfAi4PzCLnLhswWvtsgg6vOhYa7neZ94nVnKGYWlNK0dsquSpHR3CTwkmdBIa0
vkVaPxZ2NM3FVCO92mWu0iMoOODyPnFESmz7dYMoPr03R9KKOpBF55mjYYdcowGkYF80jBldwHg+
Io5qja9hTai4Tk32+9DYLt1r3Ho7eKOK2F9SgfyDe9dh2C90KZCQAObppRq8lQShNaCpeKLBxtV/
DnQhNl43bu9Tr2HND73PQo8StQfYPDIutoxT8Q4XRnmBzC/EDytbzj14ZYXCNjRKyL0xtW9R/L2A
QzISeyW/oLVEdaFFf/8cKjzwjg7cG4U5EsUrfnGb0y0u2f5RbNRY1IBSUWLOOoTklfvICdj3uQl8
1wWS19uuT/SaDC/jNiajehscECsCBcZoI/uTwCCuMi32qPCHuTolCiFxks+mr5m1Aco1IUZI65wZ
wy+j5uqxjcvBaElW4+OK+gklqeGPuO3fzADLeG2URleyJiuOylhDPC+tucMK4tSKbr6ywOcmkAEV
jDau1RBxt8Omx/wq+majkphTRhRiBsAkm178gp2c0W6dkS2/cfiejBquWIuDuDtXu/CPPOygylVL
1qObmJOpSnJWS/gOyOktXvMcnAv0DQXXgkNBs+fZ18+a7j8XgvmV+ap0ePPGu2p9ciDzBxRiMxnY
REqp96xI7A6w5AzIUjGn3+0ZXAxdGk+wTVzA4VwozvZZsd+767sw2JYSInIcAJBmPQbQpfMbjtnD
WqsooJN7lmqA6X8GpwD2I4fR+23ULlKFe2boao2vOvurpSdNZNDY6LpRGnOQ/9m27bxPKcXDkhpf
CjENpMoOBDKnTQmihqCaQY+D4FUl+42Vhb6drOj5RsVdhjwb3CpTAXt7zqEf5SQygmq2tDsDJrmw
XnbSFP5GrU01CO5H6Pd/H8IpklJir3SW271TlSJDZi4Vlh/JsawAuzYOkDoMgPxpwaafNWkpuf3J
0Ot1apAc4ZfSNiBpH8g08HWE/0uWawqzNSU0xxpnsBiWwaOS6h1OvZEdN6d0PqXvZDqkIQGAAAth
/kdYBHYRcElgbm/xtIKjBJ5trA8OeSoVTvUetuUKeTVris0Zrv++BEEUTE9eKryAvolhEvbjDFUs
WP6orwJp416c1VWW7XuR36HLjQtPAgvI+SzpUKsUDAqSTBkW/WexnbcYuoQ9AmHAtljTyrP5TXdb
6EUcTxE9qxDSNATecxGWnUwvVTcUPq2dr+SiAnM+/Z82GqMtedUeOUmKCaQzUVzmZ4o6r/IrsUyL
2fVHj82at8oTzskIKHP6bOs0dzRQJyRrld23BN47S85wK8S3FpdbFnlw+0mch7mljKlf3ShpstSq
Gp8cbb0XoaOXDnJBud3CEV1gfrrygxZzJf7odMG1UC1aAKJdFgQEC5nwLW5apRvzdNGv+pFrboB8
ZZuZjPAnZY6ZhSNXuCNqg7qoC3OgIMqUNNQRhUDaEwSgEajqYNtB87rJY0iCvjsmrqYiJAEcbmFg
yuQcWSsB5UB1Tkf36P5hV+SRmrrGOfaa9HxemUH+zD2kmedzsiLXMbjoMe61rmUoIQ0yFlrTPoCh
Vm1NZjH71wK8RHitjGhBeV3+B/jgbZj8uCHSKJ3DZMwbsNjwMq6EQGJ2laZJjVk+//gxQ2t0OTSP
tmbyzLUYU9lXw95cvdm4TMDfKUdjtljxPfYmq9g/CkKsI1hYlIZApfTMFL+reH9q3OkaAhDfMRYl
4fGePaiD7V9Bl9V2Ds71IJN9nAAnjBdK93jdVfVf/7KOJ4KCf2Qfjub2cgxCMuem5k5euiKJ76QY
xHVEbdMiiFt/V4WNOAfinkzQD4fTOdc7DotjWI2I9Z4HNDfmzOAJ23XAtsIoR7JbBT0I8S6xhd3k
1MLbdPH6Y7dYDDHW9H2kviS0l8d9doThmE32ayjTiUSollCOygrkXtgbLrmB0BVd1EgyIDqon5GC
wTIy1o8XQpQ9lF4toK990SSB513wOLwJRNIl9SjQ9b8jmm8oIgYi01HwgGVBt7z+ip/nF70ipI7u
rDUQkpdXEn7QQQNdcUFx4YBXLIUFXqDvjEPF5uFreiBSj/tteZSyUZ/0i6MRqphN2Zev57AR7xdJ
a8NQqbkPEHHilnpLt4b7J5VPoQ+9mz6GATOfQCoBYRFAon0mOj5o3RtZ47KAfY/a1yeAWeMMt3m8
VcDrP/LTLkwj2kmVcjgSVnV2yKapLVXeCgdqi2vhNF5aoPgN7iKXgX8n6qJtRYUAqjGBO9Ae9237
YvteGq6fqqCosrEdd1UvW4sIRWQAuimFunpVwf+R2MxZxlCwWYK1+jJw5LO6aUzedLgfEvom1TD6
2QdypD1HB/bYYtNhGfmvHE9UrtoyT3hPDJo8FehcLSEmC8VlUCPmvYtXiPy+nj4ZdOhEnE8VReeF
bEv46WaPecK7mxqcO6YEsbOzNwPpstIwuDAZMlnuLWCDdkdQGBxh987tt0P7EfFxX7TJumEEKJor
hCrrMolXfa7TKfLhMiJ7bF2o93xWXoy5rLN8A09jlDOIPyAkzRlHBBfECdwgzu+nZKIaUYkSQaVx
fGlEXQS+/dHNrLSvrUnKaACrYTrGYp9c7djXKet8G5qGXxPEQfP3xTGAZrpB21AxFmElPWaWgtmQ
lQlPTahb119fXZ3VAVUwcqA/oriqiNQ7ZPnqI6lQs744SS5chtVVkppd61Ys52Zu2RnUXs+Oykh3
OXThkmZ5bAmi04q4y0ZTegwReKId184NVeUHvd6lIJw1CSC3elwrFU4C/zaGEot+9JAGupPBILel
hzhYNPhrbOKiauX/zdNY/tM+WMgyFtHuBtNoSzdf54EhiThtEnlri/nH9kAKJLWrMhmi6+V3MKS1
rpnXBQ1ohzS2hhZA1GttcLOqGpyDKrYVCpJLEuzINLQje879C+jjqfUdz2EXqBuFp103lLmXDZaj
uvnDzDkbrNE0iBHgRkLTbP7gc1ZbaUSbttbXAAtpvGLm2/BFg5Jo9sHlGUZQElvqsY2/Q7xiOt4j
J9dM4ZwNAiAOYlQXW1f5KFs4B/bZzU5oxXwRn6ER3kqca2tRNRT062Z/rjs0+8ajnb03GNJIvLSe
riolG5GXDSlI50L3f/nKFNtyP6x7Zy74n/GEncYVZ5I2+MYhOzzMJxcdP0ew1HnCOuUrKrPotBSA
IkFtcYfQ0OEV8ePIDc+tXVQtLUBVwBrFTeWb4hlMgCcUa8B5QJl1hvCcqGgZPDLqdCsIIbQ70gjV
6ypYxaryMqtQIDjta2x4jhXNoFzVQ7KQhUmow1uLmGK95U8P/6iC4VvrYFn+fxeZnTmZWJrx0luI
9xzZSVGqWgVCfAzKOQlsND/aVVoXWdSjqWKqt9YCFW/4zMHgHFUYw5ABCmebLo85bFr649d0zYwA
N3YjvCio3JrFygUAxodQdzBhgmgeNoOB49F+D+bma6pdg8015CeZadogyOyGge3jfxjcO51cBtCX
vyJvSHmJAtc93frXgUcAB6BipyKS1wOadg7Rsbg7F5v/UYBqn/GCofLkU0GkgnUiSeiglrHAgFo1
v8+D2KdMjDFuphngREwYFcmECwVoElj8sGL0P5ZDc//y3ieOTbwaVLKcN5sp0vX7qdkdzelWMBLR
MR9oJAdNBXe49AtikqN++j1uxFg8xUHl+k7qCFYe0HIEE5p1CSxf3u7O+1EVXeV8q5+y87jLFwZf
5oKseClH5WcNiLTuZRBovAYrUU+0Lr/HGx18AE7N0VwNNtYMFDmo7qMEtqHJ4zUakntdCAzMkBy3
zgjMulJIplYBFms8Q5mgUZjIrlTp7ibWeXTp+KClEACt2zyKQONlsTZQmndLCQ1lsObM6hIb+8/Y
Lvaw1YGMeiwecADaVtkEYt6jYLIAssgVc3DcYbByfS2zlK13TaOuXYZglyWkV38q0mvE3gO6gNqr
tjEQrKoh3gzwsiLkATOlFwNmw/9Zl+pc86+wLc5PGInbZsiEbMV4l8TmkfRZncBZEDyavt4xDgw5
K2DU9BpJ4IralK4CxfD+tGF2zEsHkFVQs2G+7lnEN1bL/ky7Ob7pYa0QvNbsXjehJUT0LEghecns
S2MSS5xxlCLxyU0lt/v1QSEu3F3uUz4WeKwv/uw/+bodcN11SN/psEWN1y1j3LbjEfSPa8tOu2q/
IJ4M1bmfcDbJZ61riEBPvIxwrFUfYos3IUGWX/2v4YmyJfDWZHdTiLCnYYGZa9JY4LD2lxvc5vIa
dyu1tAl2ICBc1yruUE+XMmC21JOdUTuveoZZcUY6o9PZFiT9ZDA9cLW/fQ+MJ4Byh79D4Yj8cE6K
lUvKRNElZC1geEkCaAl+gdB4JuUFSFSoraJ4UNS3A73PVSCoDcgMf2y3N8XhNNI0Iz5MEzxoZEwZ
3NOWXWGudJqDyE4S1W/g95KxN8bGnrrY+khBUEew2qzOzkmSfyMCA7LIUK6heylyEcxBV/pJ3exu
ksoQ4iOKX5Ns55C5EY3QVyo5LDtmwcE5zANZp7SxC8LhG7DNfZHH82PRJMYBUj/RRPthss+5WHsQ
aBvH5O9qFk6u5VWrv86jlyS4MsbMB+H/kU0Mg/nUquWyDLA3jpgBn3ZZiYwHH0NceXxQpUmKwBCH
83TZzyWnupSJwyrPjk9aLDfNlN0QBe9H4ZkGF8uzPJdqO4udwW1aXEHAnfZGMwt0wEoXkiZPRNy+
0IHA2kRIcsAcVd/lCtck1nHcIynDjvTCF1gEHOU2f9mn2+bWhXbRuWTYsCGOPNQTRwb1q570At/a
2E5FQmFMiag/IpN39MYRHXIwvSxlvK3XAZmQfmRRmv+ZLnItrgJdRlH7YrO/+yAzyOPmfXS87M38
qyy3LUd1gZPBuQYgM8njfGoOI7TwF2T7sMAR5fQDx+3kK+svDJ2QYmuDVDm6wztt5mX/FMxfoj2D
FiGapFbirerciuMdudeJmZUThXs6m23xEQ28MUzAn+G8ZuKjT2gRqSzYdwQBXzSjL4NXNhHclBXx
aHO5RKPFhRy4h3D4ajIq3ynfacJR0DvtT0xCfFV7R7dFufGn+mlwwNyhYTwnHYu3B/XcigskRg13
wkaR5r8uXA8ulL31wAp3PZ87rcUo2Zg60BXOHoI9QHMNom/oBrxaEymNwt60jzPsgAT/b7iOX/VP
zQBzacOTBBK3iK96ayTsrooVD4lAb7kXD1TlbsoxeU81jvg54sRk1KNQzG1bQABGyoW0Tgbf3O6G
ckdPWyuN0ra32zmRxg/wFPtjfZjexF7ZFXmXEEdzo7DkI0AOJF+muluuFqLe7LzYSlcPIKYrJGHr
VnmXQwXbUplrUWo3IhtHbJq/a7iP6VKOvMLo1xSkHvoFZoP370fiXyUPeyRC00Og6e22UVyNdVEr
SdR5zduTmfHpaPSL2O4w8M/swtY9er0bmzFEhVU3FZ7XPA8Mop5X9qqVrfBt1c4Ih9ZSi6egTSqI
A9STJqYZhvBrbYGbfwJNdIg3GRKR1KVkBJkULf/H8ejee6tnj8ea8d+Wbm8qEYV72OvBMU0rSzlM
lmBXh+axd1wi24oJ1B+pzGAWRlaD+zc7X869kbAI4tvjjIHxNmJmjkUTCKN+2ARgwNxJ5ajWdHhb
M1oDbWTrLpjyLCF1sTkK3b6ro2W8tr95FAZ/wifrqYPlk6TRmpQBPF/Q5pJY73PmEJF1owk7Cx2U
zU4o3wu7c1iXiFWlDZ5nVcqiunwkho662+fFcAl1D77xBw2QkdsP0X7S4JFaeVyTfj2NyriZjwIJ
mR5UHObyarahsOvjxaTc/RbzKtS0JC7vA3ygMI7JmI985TRk5xVSpIcJ6erKp+L3EfD1rwJMdZv4
eFYJzJL66eqj31yedyC1yDv5FFgk6Qj3EzVYVC12jraBdqMVZmdthj/5sDnIcr7XmttBiWTIC2Ut
NKDqo9FS29ycXU5IGWcL0oDPx7K1iP7WPypR3hRj2n1YCwBduA8HSd4ylkGvtmiZ4TAlE78b9A9R
MNXJD0dM1n0blRmMofTT+t6/N1I8ejFpeYzHMibRYN5Irsl5JceeA2f8WjzYELuV4q2vhZy0GhfN
CJcvmV7t71F0Ox0VOhLwwW79kQn2VbWI8d7oU+oVNzgXqoN1x4LAJJUkcYgqU95MvaJhEJ9V3WH6
zlf7oq1HSwuePRihmlt2mE0SRxOwTYe2foW7TjrBt/gVK25S/KskQW6qxx7oSc6xqqvF0zM5+elX
dMECW2ZiHJN4hvniOqTbjy1atL1B0LYeK1iNW9i+Q6zgyxq4u+LsXkgmUBL6wmbIvNEhLijfbHdb
3j5TYPsFuSXGZvpHOBjEXC0cBnyGOEc4YJquxSVbPTMC4qjIASfRWl6YvSo4dqX9Z06IEzRqeVuG
cTh1m1rN6sJwrlHVtgJoZdNbN3w4JGuVOWBRvLLCoRZ/i3H+tHGbpgpZQ98Gvy00HvtoF/J0bWLL
+144Hyd34tK7hp3LrFpNyFYM87WxAGCkfH9ZG0wFCy4m48syEYZR2ujJbSKgo+NRthGcZhE9Ughl
KcTzXT4SRLlEkeOqJYMPTgz9QXAxu+YD+E1kmt9qfHoSbzny+l1JUwbsfe9GICYeDV+/S2EBZFvZ
RPVN8q4OvH4Be1gSWmELm9sxR9WuGEAOaIlqNj2UclFWcyixV/nZPELRTgtwU007KmnjKKTu3gCx
DZWm0NanFNh+pR8BcDQmEgoogasqlV3e/XJCtSaVxNqMXkA4KWUOhepsuPGoPZw/YuFIMeXy8il3
tm+IkQqQhIkWqQUSTrFkFZbSQrB77lCaHSS1+yG4olttwOGSLV/BRVIWwt4uxMv0D10PRpUQ8Hgm
hjSeOmhdMw94Rj6Q8Ik1YGOQjIGScCx0AOjA+DbMp4CrnCZ8GmrW6vbNxuGPNQ4+OM+G+b9Kr+3W
X7ZsD6b7XQtlHKYYpcE8lvhv5FUHJ2auXivbx/vnxmKPefJEOWSfAxqzmlwhPIRTiot94mCtV6l+
UK8JqGpcc2eyStoyF1TfwyeYffZ8E6/0sD+pkGOiw0fmGUJL1AKNNuwTBY0JFqukiY2O0zX1CEQg
qExovKdkT1MQ+/B1ZdA5JBxaoZDS3syfjuiSdqpe9hCIaYyN2gAqIjh5Yr7y/Lvq8uazIktEqwoI
ifLCor14EhNQ44A2aA1pi3Ax56JGz1VjZetS1O7FjPRfBKG6TjTZqsR3rL5r5AkUa2SoRrzWgzuZ
C6Z7l4lXW6+YAU1BnU8lDGJnGEO23/HM1dgovQWymaR8kGMJBomMXHbE09vNjnrHJAZ7SiT5J9ot
mNNAzA+OnlA3J6ykZGaENB/5009q0NsCLFGIQwwndorKsmkFwJnv4t9HCUR4P0OWh3JEGdm0v0Qm
6PkSfiP8ZHPOUHhV0rNUqNNybrSH8Vhz6GY9QbPP2ADqHp32SyAf27CSKXeMzJd4kRUJMvJkdnga
C61x1v/Je5thyIGZeVtnrZmIIiYzFgnkYZOqWzaDdvL/QYQrOCPwI3xBQyuo84r0IDnkNrWhPMCP
D3IF8rzP1U1v3xT5QzYdfDVfj7Iwv83zg5FC6Z/aa0nEef7o38DVmm45WZxQWUg2yA7QkLrVQNsm
kkPrQHHTc1rp1tigBGHDqKLO2jt1//U0cSwgHgqhKD8J6/bfJnGdeIcHii1MFzirrCD/OjB24B5U
SqAhUb7o/98+2ZgTdCmdMVCIOgDLsCeCpvtXz8CAkhNok1U3hVuD6ZLR68nHHDsJ/8l8jwgk4VRa
qGson/cGJxG2NyadSDamumtUNMkvo3lZV7NQvdUhUwmhZaVHLMGdVGhyDo+2P/JJJzECA67EDM+E
DvLUFoWNretcEYPk3jRrE/jn80sNZCLtiDpWj90JvTwNa+t6c396XKlsszyf3QlOrg3gwsrKIIZz
lIRZkSEtK0z8I1JCf9obbCpO9Hk7hr7D3SahvSFxqdaD/grwarjGiYzJk3ZmG65iIksEPPmtxbks
rc+e7kZr6Xk6crtm54ahAQPlwAgq1LIVYIHhL2URThnuQ/meV9oqBwIgTMI43xSuXMj0zQm15MTW
L9zv+ZuVZMVgZbd2A7wHEURNinBsWMoVWr6xF+BEE/IK1u/CLXYir7FjKlNsGY9LKm83AR7UdVwV
Icejc4DQICxxmmzDfP7GCjfoZszI/hmWJoUWSwF8hvMaCCLSoJbHcvRa1M6/srpiZY7w0/hPSPTE
meHNqSv2b53M3rFWbJxjdB9I7rnPjOWxc7+uay8Z/xVFT4iqvO+cdjB82gItm+TjbFxpPbC81e7v
A4chJEmrze2wSWlFttKe/OeyYK49HgfNrRrg6IpXIQlbzR+LW7lFzWbi9roGg55H5XEXPj4k05dB
ZOLJyvB81VljK9nUveI/1F6l509xBJb1K0IfpQcWVz0DF8w+TFsNEd2uYCzjFJS2aKjmHCSxwxTW
BpDPy209n0xE30d7ck2k6msb0ufenvooMjjmSoy3kmi1p5oCBDQUSVtKDSz55JPZ9PH4QYHlByLK
DSXsMFyra/l97fpHoLqzpy0Jz2FF5oXxEHhm3lQyDOwsTiivwUxoqmPB6e0IYUO+07EgIvBN5NFe
oRnzUnO8/pZlXNS+foTHWTs1GPGeKN7Mr80KUMUfFIQo/HVBkLKw00DFSVrxVjBGkECi4BTnftdB
sNnll8iYS4B20zmkJMYLeS69iF3FfIm4ghBDpApur4TIa18bocCSv8SI/BV6BSJSaAUTFQj7pG2i
CmJKB7s58HEirUu0ppaBH6Fom2dwTe2+lOI/JLmf15Cg9XQLZtiNOkyzQ8YdakQjdTc9sxk/j3bB
5u7dqceEHJnLt/4QPhyAz35PoCkCM685BnZfu6Cd66wwGwwk+z0oHCeYU5FlCa8qDJ2p1Vo4ms3O
sgywwL5tw1+3JlRXpJpX2SlyIaE29YJwcKkNDGrWjo1UGDlAFsvb9pC8yVtkxtFDKfYNlSmWIy6a
tDEvacIufZHVCkL+XzHLdn4ycR69f1MTr5j4cFPf2a111IVtHulZKJInRg1VxReFTP6opPhx3mI+
1mCRAj5ZH95w7U9XesDwamu74yAmCRaJgwcmxPKBbLuqDOFgM24Hs9GaB+DHQRf4GnDq+2ooCbOy
bQZqlyeqKzwBlSRamVeg1XnGZJQDvtKzjsMbvNcaETXprco7PSiI7gsjW3drFCiSQo9dIvciLieP
Z8rSmtIQbpiicbrxpeRcPT9snMs+CwmFNK4vziLP1DMZ6ALjjhSJFi9RE9iUpsvIACGhhPLMP27N
zwxaY0Ce2evWHtLFs0ozs/H+Lhr5IDmHZ3bLd7gtMTHx9NUpTqSuvpaVmc0rCO71ZiiPA4krJdqi
WwUpSHUks5FGk0DQT18la+d5WEiSdCKbO8HOinQ34JE0MD+ZHClYaBijeKUmgGlJu3tC51FpeaxM
lozbXl2kj6glE9IB5ICgBI1Fx7pblqAgUHi9NcfNRG9S6hN5Vfpox6EapN0ULFdYQ0vkjPdeuNlA
3a9pGjz1y0bVPIrJKtVQ+IJvUrRVTZw/iVChOi1dGBtqMVB6rIVVVArbfugUSa8Hm1aKKpUVucly
XPw7AxJscjEq9BJUs57KIeOYcfE5kPD73nqyCX3Nu9iqpndMUmkUC1sH0415ovmkjAb4PxOi61OU
LOJpjduTGicQsXJXsiZPCn6jGBgaQwTJ9clNHtWU2gM1gDGGkU+r1+Fz5HZANhhC0Epr515JUAGG
8hEIPK3Dpkoy51WhZ6jopXGuSL0+g2CIMDH70YkT9chlwEesxEkyi9KHy0+6HZoyRFoYqCV+wmTd
6w/UWQPd8/73dcExKLMtRSpWfm2wyP8jkp53aYUaLWiqkKlrbqzQrQX5lWZkR7qmCkT1M1Uw8uWH
raPSaRDje8+0veP/GUaJqXhR/Au0iT7cDeOeBZRWOEZj5yK5DmK97mnN8t08VRzo0Gp1ibkmY8cr
tfy6iExaD4k28WO29jYm1lzDB27oUnuvBbVvtzL1BmHLSmIGoWvU+ZBJ7vXX+ImC0IJQlMTmZa+l
6ePBCJj72glq24gsaFb2pc0EvYgJMHP19xjuATDnATnXSTOlioghFAb34ktKA+SwQfQpf/Ri2SzE
BTG/lccwL10SIHWrevuofA2oqesBq/zeu8p1BBotIygTnOQrS8K+Bv/kxR4ne9GdMWjOTmMv6i2U
wYxs/IWo/QqlN/ioixHvFtjrPl6PMEbcxyHFc1fm5ngqGyYXAVGHTTSKFmzU8W6k6CZHeld8J4e3
NsmXtI506jZWI5LrBB+PsRYPd630geSDGVHidGPmW/sokeMBwOvSZgEp3aJUxIL7K+7mmWXEkK91
wUwqdMskbSYHMHZumLr5dDaYodOY0S8fZcmfp+064Z4ilsD2EovnAHtJdSEJWQ9yXdJfDc7UH8HT
Xv+7WnPwSeGubwpz9mXH/hiejF5Gmg8sFMgb25OHjiesVgnTM99KdiT4lsAJaMlre5L+EwxYvoor
tJBAM8Ew7OTxesXdhPtVF5vlNHzVeNpmWVX+49kk3/Uugn/mLU1Jee0rsSZbOWPEso8xYAP1grAb
gCw1ufqjSgJS+5jQZHLrmSKyDb8abUSb0/cBD6osS1xM/qYBOgI2TS5gJHrXNQNtXcXYb9emtVrF
wRd8Y8mpWByVnqNUdUyFFSgKnYVo+h+axDx/3idiCLI0D3MGbsakapylgXd/o3NPMBVDxmpRHwwb
Zp3A2qYPZsJHct6oheFaakMytJiMJD1XmwgDyZLPrF7lBbSH7C6e5wgpjOAxfdOMnecI6h1i5IPK
VsdU8hX7U5RLFpJuodOju64Obf0s8TiEJt1KV36S2oieCRCWLfn1SAHMpWGv57woym/3WET5DwaP
WYi3s+tFJNj9vPI4uVxKGFrtUHhzldnygS3FEKMDO9R/ROWuR86QaLGOvRnm2W4OF5jhHudwa2/D
EGSuviunMfrfqo8vD45f2AWwaF/FI3HYH3tTriGaCNfe32kr7kZnTyimx1aoMa4qKO3N1Dxpz/pO
AdtsxKbSUibkA1ioVXxP7WE3cG3iMQF36t1KQn2FvWSfNmIpwB4LgqP26l29mMfxXXq+NNTijyTn
+6Y8/1F3mKmkhOascXoeWxDY0oJuAngA92tO7CawZDhuA3NA6U/M2A0JywER2yGE48wlZKvGiGlp
bAF0kTQ1UBbNTXL7A55O8C8+LJRzBet+qhxDg25RjwhzlmTdzXRBcqVttOaF1k2lE/MA9sNJNcw3
oD5es5Iy8OjPzyQKlFSkeV2pappaP+aQxjQ5uQt3jx/QctuixTbQA/0okGoqzBYZgXDXTlIgSeG0
zUSjiyvDrYiwUO6KWwe9Kj4F9F8t2KyNeIGCDaC21KHF16+JfEvnKc/IMG8svbDfeiLYnj/wpGL5
rwgw7lBusU+djxkZnUUX7CoUw+HK6+pLcTSfh8r/2U8XbpcWmcYW1juYvdqoRD+7pwZ9GINQ5D9/
OXwZuLOn3hl2yZ+iRPlCRS99BRpGTg2GV0zPP/H6D40MWx4JrvvngwA1PozhYoPceahVVtq4DPEE
8diExU0X0Ldg3tqbWJVhQnDIaY4hO/8vpndWgSy4dHgS99/1TOI6ZFkaAsPVOr7Z8561Y2yMa04i
gCA+QFBsGLuxMM52rPeCltVMCLeRxp++3C3yxsUMW827Q4AhnmSUjdGtjabhaJkm+esy9Dv4QPHa
NoDVWs43GJFbQDCLLeXPhbT5MVsIdVd67Bzgh5hYFgsqESQlumSP0y/7ebHIdUnviN4oVoevZowv
C4G+E8clBnBkSw0ohice43AnOHFYTik1+wyHDmxnpmvhe11n+CnZngAaCurOg28/3GxnxukpnLH0
NLKTbiDaUC4UAccoPuUQ+ssvnbHueP1Iv5e+D+zEaInRY9GLS1Ulju1pntMZXuLtkvk0G3r1pxti
OGBuQEUFZs7sJL0I4jD3QQK8ubEsgkfpYdqXHuoIEpiwpgH5Cs4jrEOxoG4v144St9Ejl0GZMSmW
QYDNChStr2G/WfhU+uEZEuDjAb0Tx33gTTSMafxdhOI8DmwKBp+n2TSkYAy3E6lrJw44CH+qqmBZ
kZi/e9LJv2EKOIsydhhWefsxyjWMRHqgcjHtiKlWLeuKdPhf/kwGo+ZD92hcCVCewDBNmFCvxt4n
ps39xjTnPw7AqnYlKYtE+ptmSHmJHouA0mDvchNW6IokgJVJ5D0Tl6h9zhRMtiKFBz5crBh0YYof
UgdR8uc8OLC1+hfsFKPyf4nzd1/hcGpQqk9j3s7cNMjDRHElFqgRUdk+W3vAClKZ64EFH0H7C7vk
tsRp0nbnbunZ5i4L+sLJ0QOyf1C7K0rUQRwuLATpYxPtvb9fZezYLn1d1GSJHEK3f/s8W3rfqLpQ
WL9seHg9RUOpyvzrMKo7HKJfk37/2IXx6Mr7VT88Nv+xJVRRRlTt5kHnQy/FwhpGYfYshz7ii0jX
JUVWcyZ2krT4MZZx3fbxE2oh64M5syOQ/7ojiM6yTeYQeDfM1hLlY6PZFAqfR22kJz9KqbCUkqPa
eUe8OFu8Y0UnpfSJJH48bG1G9ycYLC+YOnqugoV8XZoTXrkZT/vCkmZVXMHMrNVa1LZ65Im2wwsf
S1GP/yMYIAspl6sgJ4XQfQ2xLh0uoeiH3s8ux03c24L0x1b3b3rzt0B+eF6MQVPOucbtTQBJAmut
zrZW+FiVdL3WLidKWKqO0Wq3Sy2cIknwEQIFE2r0vq5nVHgQ0CO7mrelKINor9vPkyEi0tobGsfE
FACKRxLhyVVT0yDEfuDdKfJooU51KejwpO6/1wsxKQlvmCn4A4zgW7tP2uwDtrrLzQGOakOg8qVY
QbyBZzjsdiuvF1yNte19e2z1PNcSda0RPwgKicwiTUQeOBYpFysBautwD5BpgM/mpWWiwGEDj3+r
YZntMbyhk4AAY2QjpBtC3VweRN7CUC24UaImKfNXR2iLR67NKOC8auSaDAkeJco515+EyKnIcv2r
u6VF2UroGQHGCmt4g8r1myFoYnSE1zINPlQ50VYN0bcYma0qMDi/n0wKplJxGINTklE0vSAJZsa3
7GYzRGpbo+e/idmb07hDk/9h7hyhnAx0uYSnQxd4lm5iMI03m1IZ+BQHaoZTKZCXrPBKC76FPlCo
yHmlTI/PvdsDCP1OTLisr7rcqkTkK1tjaggie84tEunv6Vh4JtYGZkpB1rWanE8sQ3uF7qYxQbas
qiLZWn78AO2+RLWM3LZgF2njoAaMWS6h7t7ebLGuDdelUpgpEUYmgZnuZPSBTAROlKcrwFV4Lr0+
aXssWV51BYJY+lP5kEZRpAiHxxVP9y7QPkfwgmHsIYejyhJbZiwzZUmrp7SvlvDLahYTGBDjmaSX
BYqHZz+0cSphMSyl4io1PffPRPl6Ys1w1w5X7JxWMljOxus3jPgmg/mN8KE683eeoS/CHb1jmjt3
n8jrEo2mqOIx2L6vO8cSKzjZYwgrqBYfecmLjyB5FtjMRSx6Klijky0mVcQF2mKgghIvfToyiLZe
0DDlt/BjlSgXrDK8NqOmYLQlcCBsBN4OcrkclQk9IHFeuPoRvHlIAFiIY+QrtoL3y4VK6Y8MOsrG
awP3fw6jxKNpbxG7jBSLcMOtZOMx4rREPG7+QwTeSwhCkDIFWimXQCAwM8DBR4FmFMRLKpGWZJfk
S4JwPFu8IGVFb5z8eysfaXloXPnW3D3KQXkcaz9LwbpVA9s1TRIOsNl/rzbsOHp/AuhTq0Cd4G4K
iMyS6U82jzT3FfO+HdRFXZU974TYufcRjf/VdLpYdv9I/mDDoxbiYmHsjpqu6S0gey9dBl5LLHlR
bqOtG/HdRVWTH0lGtAra97gMlsCkO7OCm1SbIPWdhAYVwPjnIR5OGSl0xvpdBRfOHswpYKmr7PrV
dciazf2bkB4gv3ysMyhfL+kJV7noedvdFW1joFW+3gTl+B3bWHfN5B5lfVERP9jnjzGLO+WcpAM9
Xmg7+wypK7q0L9yG4/VWrtKkdtJMZb1apH4OSLzcbXBpSRP/uWD2mvWQXYsQpztJ0QhKLoW/RoF/
WmU71GuBZdbwySlEYjf0bAd6kZyoRTVuH8yW6+m9mZLWoAZytmPx0exHfq8dnqIt3b2sIGKf3ls+
EapvMrC7yHu2XvcKXr2fzCram7wrh16nWVlRnkJP6jH/thnyNIb4GysJKZ78SgFWjQc1EFrbKu0Y
iPK1+PALJVz39r0aZdLUeGip41j8dJLc30A1PkhI9sY1JPbwhzmBdoJZbr+iGdFHJEV7xvq9KOH4
WRClYvGThyvaq+4o66qKogt+c3/yR2KRXKHvgAj02bzj62FR1V6/rCwlVSSODFWJm9C0zjg9B9Jg
wvcwC+KN0twqXlTDGtoXJjSTpvdestVE9X9IrlFjHbz5gsEzhiuqpXiHOBPfkbw4kJGGC/mNxAoY
00IV3E1uP4ZAL0dMwVxunZ9oBuGo3ay8tsbK0DRA25ZYkutlHLDpzIEQ9x0pkl/fVCBO3/8r778Y
jtYzmDM5dP2qDKbfLuJaTRnHw5dS/63eyJeQ5ooBTIgx634ouzJ+YxfLdJx+CiwG0j2dTHi+89EG
oTWuH2b7Cqgxs4CA9500FINDkGeiYblhZqxi5vWZ99mOIw5uYwQ22EVnLOAMcFVT2l6ZuvWV8LcR
u+xkeL0hHjjXAgKO7gkyY+MHkzguapA21Od29Fi+tXdzNK5Sr/PMyORxv67EJw2jKgSlTtrWfAFm
83gQG2EwJiPkNeg4jdPwudPEfQ4RdNuDzBkePUmSIh+6hR9Qru/LnO+1qiwPX4kmsYBm1eQL1QrM
al1ypySnPisX7z65gs8Jy6jtvskqdR7CebPZPBSS93L4a1NDqPYkh3q/xzd02MyYLvsXttmSHREK
MuXm5DzKCKMLZRzshu3Cn7yuY2Yqfm0yDu3zWtjqWSGfP+SwJ1cC7eprpaWsbzdArhDSLrxhGGGY
PM1FNo4EG38ptZjQKwOG5Nt33D/BUeBAh4UHL4PxW9A5wX0zMFGBDTKw/Pe3iCrOGTsK+zJpZOaU
F1IlUKRDEoSJq8f00Zwc/uyPxXRYMhrOnzQNbOBuqBnks9gfy8puBDUeJn6uqASe1Vx1qRev4f9G
a4Wb9eUOuw3zkcLSbpyehdPoNWxlQxlt2UY+5qfuBvKQEaV0UcfU/aaOlRyv+Izy2lNpJm094DYE
m+sCdBYMJfETYnKUb7OnbZ+W/m4v6tQmsESJ9K2FZz4KauzpGCmwhL7pHmocow0PJpwCKyZIYOBZ
lc8KwzxMTNheT4ngY+uHnVkVb40BruZeRmgDcQ9NHKi4+iws4d/VV1iyCVaoaqN97dXpWgThp82j
YGex3EVszlkyX4vJloXpXIuRwLzaPVl2w/NbSYrB5vEWOPZZ9mRr8UiKuS3t236wmNgtr2X+evVH
pBpUo3MDDJmwnwSiM31Jn5KPG90pGZsiw4TkFRsNKkEtoVIiXR7SG6So7r6cBsv4Jm8IcZyuhJI4
y1HLo9wmfKGTG1IRYTcz+ZKp4w2ddGIID1/ZWN61I7FOVb0xOk0QtTgn+Pn3xkqRjG2Yh8Jpe720
GQp+bIBh31ul8H6fY3weLLv1ZZ6I/EHqh7BZCfaTFgHyXSHywmruR9sZKKkLyKy5EFVnlWKv/NVe
syxMvpwaQtjtsmjWlfZXVSeGzNFVMMmfYLC5BWx5MDDaGv2n1K3WC3O2hcod2oyg7eKUMX2ygZIg
wD8/5ZGybgISCHSg0Ci/ZAzHLmN3kIvdRAjNs7CBzzxItvldJlH+p7ez9II233OXY5c1TtW+hCVR
TaF0pJN9jvKGKs8NEKqoWtjwqwXrAdlm4qenoLuaRsaUI8g2NofEH20yb8zgdl0y+J+YVACCGWi8
pUNX/4x7vzIoSvipLHEJwDg9ImP5KC5VbOxY1N36krxzNfxcFft6GXdM6eJkwsygSo7rZ3xS0Y1P
7lTS23OsRJr2+tvHyeEdGbuSI2xr3aVj2yzDjoxFoQexGpVl4oSTPH94ecoA4SH73XAFY+0gR5hv
IOaXvo3QGOenI/G/0gPD9+ROY/PmI4Of+FZVsZnqLcHdfT2RcV0Sprkqa+ihuMs71T19PPX/e1aJ
1QCjQsIe6S/UVl9yvuLx+HClGxqWi0BltkyJjXiZ8AjSl1AueD1dCd+0Q13V8rfCYjcjs5TAmKKU
GXI49TMraAQ9XvxyJVgVPmMTPYoHM8C/pLNLx9z2VXf39SH/XTlHGjuO5PmfA/bmGIvfWla6SgkJ
ROeS0OlWfJLOMWswoGZBa3MBX1HFOEyymcu9mtstDyypkER8cl+UJXVKgLQ5Q4eh0JD2Jyspazny
TJPnAHHIZtU3LzRNMPOpAo6BcV74rTQQQyZs4xH5ikX4DxJZHfd0E/PxqLBIRqR3gv/p5Wnkl4UY
dq5YbQdjWQB6XhkCGbUXxCgjWTLYqFX1gBao63PPb02Dqj2pGgXasijNGD2qy81eKPh2FKQKHd6+
9xMZ+rZIDjRg/j2fqaUGtA+qh2o/NtMix9yxxqMiekwQM/k2COtsN691awa0hIA+LdoSfIe0LmzF
Pj7cdldSsWfzNswV1NWv+klwlfedFHi7hFEqIos9kK/8FheT6erZOrEy1OuxEzUFnbQ486gO9tzA
Cy6XFzRqs5vrGSVNuD9qKjj+IZxk9gzsS5ASzSQKTxJcjMohmX9zbXK3bxvQxo1EXWOiQi9BDCBL
sRDI0cbDrPSmNE3Wbq+VogTGIe0lyw2QnNtDzU1mY23vElLEjVEXc+Q+BqfFaJlkCYdW+cEUFHJm
X2O5Tn1XqaPZrtkIYgOMtWMAEknV2Q3yFcA0JdaaML6HES2quzeDaUBHwjNJE7nr8g+dyvdi180y
hMIUKWSXy6JlcWUdxVwTRLMaLZ0U36v7uBC0PRiodCfKcoW4aTPIrIeigpR0QPsdh5KmYBBR89iw
wm3utHsyFbxQibqlcmVHC1raApqA2HJuAMljAhsFJd0e6JDriD+Ogfu8ObS/NS/o+MaUyue9B/Ug
AdnZZhU0IvbgAMvmhzH6xglw3GxTSsswk4SwEzaxqLJs7nGD7v+q11N3kfU40alZkItoj14Z9Q2Y
LpTm+CsmVdsXE2k7Ai/2Udj+CnBFlV2iXv14/kID9Om/4y7LiVnMvPfqnkPmzwJxmPXQYD6wdJ87
TFvO8vOPcWXkgWylTeTgaaIIbY1w+g5VAtd0Yu5uATUY7BWbLJUa4VEo8fhsneZYsMT+UR/JS31h
Kl8I+VvMANVimvxteF5NhNdJi/p7r68izEvRbpT0zuSyX4U/KrbSvwxJOOuGQfOhGsGPdX9NAdr4
vvC3rjbxKQGeXTkdzeY2NJ4+wQ7JSZff2UkPs/srv7/0jmuOK0TUiKGkAWoE+6UITI1Z/U1FO/lm
mIy3VsBs8F2aSqPG+eNNduxRC097ZXkz12wuzyiFHNZ2sWeo4BDI6LLsAeEylXT7yGtaiGt2lvGw
yUuQ+WKEMfjluMlqCphNi/Y931Ad/kGB/wVx916SxxDXQxrpiS+V84iwBKNdAvKgO1Melq7x0kM/
38JBUvnMBl6vk2jl7NJKfORCdukFfbSPLKtWOof2lAwcVtQv+vesgRY/dR6J+PRnjLOaCV7aejhK
31A1EEVMl79l+oU2y+IU0pt/l4PDcJGDv8lcUV7citbvfgDI4OMr6OH/yKXw2yPTWJhqylGbAlig
eqicjBczDm/c3PokYYpdUYXt9jKlAu3bHzoySVkGpwOYh96x/1PCfNmr7/njLCp5M7XChHUpB9Ph
ThX372dtWQg6uPBJdloxF0PjefUlq3ykDysfTTfLekispnio/brPiCkRXoquRujhDJSouFHpK0H/
Gg7IKu9MSzOpgxDvqIaFGeiw5TXfGcydJ8Dlmx1CbAj0EhXPqmzzmDOFVP5u9wiTwEM7fpzfqOPS
LNytyaVq9voxNC9g1cw6AW8vkrsTyp4KYEVrA/do6ysRHAn3/dTP8hUWmbnYyUYR5TmLrVn63z+m
8YANuT7NeRqd0eCpA2sMqBmamE6xtCr5PEyIitYJ1fCQMxxJSbCxYC6nEGtrFnp8LbIsIz+o08mH
LVP+HTKYg5gUnYHoLmKBdad8FQh2n14DOhiCgz2e3qKOiDXtpHOPHnVpVNr95HNaAlXZhO5F3SSW
3zGMq2IgF/UGD3P0z9enqdrDEpFHFc1ZRKLXlc80k18NrWv5phnYg51CsICC83IUO5wGpRuebcZU
ljeA9f9SqMWQ/Z53gcb4/hGCTdySu7Lcn4O6UHUt2X3+p++zEUIo6At7yA9ooPDH3Ph2vdveafdT
h6rFFTdNlb0kF0U6NuCVB35IoM0/2xppZrhDo97ODVumBLv5fEvrTtMe3N/5THPq58KwC3PBc3xZ
O44swCwm3RPDlc+3oIrjrGvRgTBViwqOYgqrUYy9JQyTAwTzxNmS6vuYBJLCkEzxnXErKwJTjRwG
4XBp3B1yH6fJTBjukCpVOeWHOjBFev+yplNYlkNcxBnvV9uDJ8iYqlwLvPUjZJFQBdoli01aeC4v
6gWd2C+8DhwBiudvOo8RhTl4YcCMgdlSjhoRNX+r/7txLNmD3Chd9dcSUtokr6/ynlYCrKy+1NR+
THqD9zjcD2qsTQkVE+m3uItNAqXsqeKV66NhhkKCabkajfK4BFeqNEcXOJbyw2X5a2w/NPCNfvXb
RWn10MnShZPHxy94psCNfIdYVI6BPrED0jF3OSkuHWrUIXIqGF7O7I24QcOHiPnS1nc1yyuD86fz
nnJfYI0GpLuEox0PZF31tN193nm3tGZRhGA+XmQSUlbBk+Xy5CUYoE14KFtDxebrr8ixsphBM9Rh
xPL5iYqP7aJj0IFN2Qux3D6K/KtZLFuZ5JILnEwTYFZDxnJ+uC6QLM88u7vvqT7Mpiw5GfIVCDLS
cHkgWtC50Y0FVxn1Jd7NIWlBD2FrjSUIcuFtWm6UN0w2QAow/vxpUBAVZsnMKs7P0gNO9YiT/fF3
YIt8LQtujmbgyAqSEPDxxq2qIpsjB/5wBomfyWavjVYKdWjiGovegLQ64OYSyNzth5besTTOkSYd
Z0PItQfdvp+QxsOvCGsOUcnRijeIwpfJNjaMw5mvDywAbRbv9O+yzNwLDiBtcQe6Jgjf1XLqA2Yn
hpv5APXiULW+H+ZrUxGNJli9AyOa2u0akOFjUzfZpmlTuccOFk9ZPOtgRWpAWJeY45Mx3tvJ6Cg5
ZiTADCCuKLpT3SniHo/pqLWYr+Ej4FwjoMAeAghWyz3X+OHU8OyzGdl3IySez+LBklNJ6dREXsj9
PXHiSQ6S8ELmHx1ZFIynZ/Rv1xs3qK/crhntTvX4vnPcSr7C+ha7YnvAmxuPi2xORJuojlJeE2SJ
fEDqLxWL5y5hjuLSFDbpcim5wL8psDYIFkh/jcxarFoJCgttOgRG9har78qUzf1H7Cotec0ZOmmO
d4gKSx5yggbVtC9weRvOIy93fxYLLSEycp96t6zAJ5qJV2AH/KFVbQ6GO8SNxVK1c0Tinofu0cas
Kut4yPAFditmncgDIDfBOG3IuW0inQWnuD+vHeu8lgafrXE3ikvNExWzb1k2EwZqEzf5R5bPlM8P
PEk90AicqWSrY4/Sx5AZu8bMTKuYRQLd9t56U/CwLQbeJ+Qisfjo7lCrMyHQkNoQyGdog0Qv3InA
Jdv53oDTWPiykhW00i8DleC/DbuW2nXz+/M3L6RINcKxCzbJOHYLfYYHSiUV0WBiKt+P5cu4hgZY
FJWDd8ArtDPlCamMIj/3yfP0ZOh18jgss+qEtnr0BQH3Ohi5liR4l3VyJ0qoES1lYZbBLqnZ13xy
ALdga5IblfMlOi0CmiZk9OPzlWYkVvY6Nnayx4j7mSZU37fAO53NAL17YrnMxJ+IlVFjBuKE0GeI
aOtXFFaNAB1LMPlUMF089jpAZ0+mximCL52sJxlSaZ5+FsHWf6jn9cokhfLdAx6f7I+jCDukFIHr
L22CRfhZkOSE4J8aZpy3idpt/P+mzIyBu6/9cSJ2zpx4GDf+brmoGLxKIjRUwGEVgNWvyzxw4Q7L
S4ic6ZFr1q7GpAAdX6DD0WLDr4zZZbkWPIPeSgl0D+iYsNj4FQiLaumBI9weEYBfI6JmHXyNOwX5
yfTb3BEf8HdyN/sEQfkoikxyzODGJ6H6dG4sziwy5LYvm3Oiur00fsUs2UAgTopS6VQYLnGzrKoG
RVDIHrnNu8NAlQUXJsurXbE7xBxoPg8pehvnjY2JCs05DohwNPlKoZJO6qK3cNsqc4Qxo9t7hTJ4
mUUnHYSMtp+mQ/ZHKsZyaa2no9rihGz+lpRx21Yoava+GUndQfawkJLp7SLqNuOgHFdysqjc7PCb
nlhParJHVkDFNafvXmh+yyN79N3qLUGrbQVuRz/p9fPARtJfqlLTNZU/DlAIi29AH9xVSAK3C5R5
BSmTQVvMQjS/BQ5VEjszHwylNH8RU7hgQPqE4HmvTebJbZ8c6k+5pWXtYIcj9LzYfb+Ti4HeXH8/
z//fto7u9h2T6HLGu4MVHuYQY5nCj0iabY31PlGO4N+1lNP+4EDYaBhdUb5HsPmMXW7QY6YDJM+e
kVcceIQsBqh88jy6Ula1OjdOvJ46Nf5CYICddpiYp3YcVj+A5g6A8wkAhy4bfuKTo8s7nCmrNwxC
kWOlb1d+9ce16Ct8zYJNXGdY3Dkm6M86SRE5TgasqPcDdDLsNehmBfaX4L97lT4KhmJMFm1YcYzr
hYzwiKCw4gMyk4hLRKQ8ZpdxOJbjqrlcIvVS5p3K8Kq4V75E8VryrBsttOGVfpFkf3atTp+PKmlG
YAviUA5PkC8gM1hsMmCPGr0y9Qg1r+SYsJQ1byJlnuAedNytUKcmBsGOqnuYuL330KI8lo+y9dnr
SijGF/iw1xw0C56h2tK83tObE0pie0EcLrqvcjTeZLvB8LUsNez9Izok+fGbROiUJkjBPuk7U6jC
j9v+S4te9yL5QyIECAel/E/zMGuykG61VwtjaBOPxN4pkc7Gp5qvorXM9SAVoI+4mbGFNBdgtIxc
6QGw1faJk7xHRS++vT0xqUjJym0esjMNgUPNzD2rFHOoXyC0N6dbSqYq8HQB7rZRJMANOki91A+q
KT7fBHbkODZ/DhEZ9RnSXvRnCv+8GoG4dPE2ktMGUu7m8XkkIl0B/EO8PKXi5eh1chd5bCikmGub
4244VaALB+h3sSxt3dSw41o5ULsgyo1yW6RuVvj9zphfmVlyERQZiQGT+QbIRh1afSSkFZ/oEEoc
u6quhVyUOKejB5o2LZSdwoZks5J6P+1eQF1V5NZlgXm6j0W1efrGlBLIv3hfLrSuvUoJIMqMOlHy
ARb0qwRfhkgtf9HpczcabwcCqKrSVPbpXnKWV2EnCaAWZrMgPKPEp43B1iPuFvAw3Laorro9Y6oB
9VGJV0k2qzhNk0Hq/BgUuGv9S16aWxo47izM7QCKw4Nx6OL4cji+S1cK2nfT799XS8Ra3NOHP44h
3iALgOIp1Qbc6L0apUbaPijWUJmV0BBnsAj/5afTYmuzQYGTE795Yh/G8hSHa7gB5jMeymVgbo3L
M3TpTXIJC92DQIK0r3c4b2yfYVXCCplNgeOhbAkSB05sSVeiHic735zrWwq2cdOFP7iESL2Da92w
yIurAsMkuqzlfVI7kD2HIq3Dc0AFRFxWB/T0PQp47Ax2FxYYzKLCwl3XJQLxmexlxxECiERWHW5a
N6ZU7UNndT5sThb10wigXXfqxoj6GdUKfJc+a2oT0ckcTENt9F+x3DUE2S/Kqgh7H6IEYzz4yudm
cbEoS4+wIB18ugkQEqhbeKHVfOJ234hNp9nzf1pUxRVDUekLFHaTnCRHp8gNPYqKJ5bIi+lwzs06
WK+T5uTvUHO0jce5KIZlmj0L03XRVorz2IT65LP55j6QuSLng6iX97OUUfu0Fl1HqtI+4HxdcSi1
N5SSDDfjVAvMj5/gfk4NCHbTk7o19A0djA/weCqilxmhu5JhHX8eA4ROjYFE7R3DG59RN+1YfsCp
XWzglZs45qABF/Y55pPXzEvfWnHuW3NGMZlpeFaOAqGwkSLFukXlHHcbCFtf7HaqYAijp2rzl3ZS
EUAge54mt5EhDR7VF+q4iShzmzzNLJOpKQhbSBJrqhCeCEg6HX3SzRKLVLVDoM2B1NgdQ4KnClRJ
AiS0tvb24yiAg52w2gXw5FK0sJzzGmgJEHQyy5i5hG9WLsJEhR6LyOGspKoEmAgcA59UpvZmJJ6h
eYaWrD5HbiOu8OsUZ9KpL8uaRm0vpn6dTyZL8/jFGSXeIInqrXr9wObr/t/QizmJ9xs398JUpk3B
8PeSABJA21osp7L2TQagU0LjD+GaQcPw6Ix+0E96Q+OnSg3gy87KpVaVr6PETtVYvw3MjrLV1Smn
htGSIoke/wSdmL1Yz0Yd898/jL8K5Nskdh0hasf9RfUCbkSL8CgWEnmWDAqQ4EZB5ugDu8k8vlSH
maZTneFLCjIqsHbHEpdUqTmDjN7edawYPYJLRBta8VJl3AhEQpAAVkBmMmgGz704p6dU8bawUy/h
GJE12s/DmCVPYvkH25ezvdm+i2jTKRTkfxUXTixro0+hMowp5882g/9o7mYuNguQOJiCJKgfCdH4
9U8I0zS+y22qDtegQ8rOfTmH3ni/3UpIM38eH/sx3hF4vOJBNN/bN8pC1EYGhsdnT0fdXJIoICgG
ti98AWpubjrPRPaWBiyoV+SuVNJ4IsumzDggtSQNUc4pXC3O2e/dSqnyq20xRxudVc2OwMlBisjr
VKuxvdjVAq/4xIO4u3wp9SK1+H/eArB35Ogh/xkUiJWvitZS+twSnoHBi4m2cq9uTH9TXuerVG4f
W1YxjBJyIbrMvWEnQO/Cmc62soBJMesrO7VKRMAMOvLu7IeKzp/Zz5uWBMh88mw9Sq1mZddAEIiy
ETquSN8TJ04S90QViUxlKqvX5IA1F85Y3WsMt2tAD4S1puGTBDcMPrN1yp1aZnGTa+1wtsB/NP/6
9ZpCJ7k/I1msjqOLpdOkuIDLuPlmDKuwGXK1dwm2OOEQGizKYLoVmSVr198a0JmzVpsDS9OemowW
DU8/88nHz2KDHsYsV2tXQylttjYFzuEeUfNfnoe2MVVaBiwLXmVeN/iBzcXhrPfSMB8SuK9AWrIB
sJsfQUn9x/9kJAsR2uN0oTZ/IOkQwdgIGLXHSrMUk7jtmsFAuGsFV3VkFy/aD6sjpc6B1NW5CW9X
J5Rch45HyAgj9VTAVmq54T82ZmZVXsnDdi9k7AArbXxRH2MAlsSztThZPbexc5zciY6BZJP74Jur
Xq8ENgv+FBVW6GQXKolctmnrVl6H0DiqZiXF2BHtbwlMn9e58prKxhNdKfwLdbU9LQFPcR02s/a2
M3EPeSNVlvudG+HnIkfjOwy5Dmx1afOlsBPPxOl8mtRovEYTGD0OQIwdqEeFQIxvwe8iY90L+gVy
vpfCCk0ZQL+Pu9INCWzlZDSqxshpktxwQdzHml9Lm4Wk9AtaFqJWEbQXQdQWcCfVkmEb3zgvelcg
yFKyysLDsXAjp4dkkZ+TusP5QVDIZrcWpCS5kJvUM+m2ikvWyiLHiArvIuQprTzKdTItP7aKgfzr
lVzKLQmdRKhBTp9x3fANflPguJeqxICzXvwLPd/cA8IzdpdPtwT0aUPnGuoGS7cf6zn2YSM+280Q
u9YZ84NOBdkTWHHeWnwBNupAjmXMci0W3VJgxJGfhQhMh2ESKtNZoGLRy8miIRDoayTBHz8Ku0DX
gTOvCn7fsDUuSd29RNDcDO0s47y6zBnovgXZDxS+pLl7lV+RTOagWmWuwWV5t4PjZFz4UzbG3PFd
iyXIbRizgMFKeXMASBi8s6X0QqnKdwIBOM2/Z9Bw5Nv39lqyiMVa/EV/AxG/sovZToiihK/xhfnO
xiHPT+coEyuYmEe0QwCtw3TAZya+9Nh7tSVw+OSYz7fU+UUcA8UAQ4AKoVXesV1/DCO6d55z0RP+
tw32rP2BNUDqcNKy6aawB+h8LixyQYEZu6yYqi1tSElDmgFW7adbN0A+kyVwzDlLtpYWc8vWAZ5x
7NpJ2C+o/6uSZ+cbY9Dk/UQWRBCDt1QtC3hkt5rt9icPm5yjX8QJM1OY3cz42fHCMqWcRSzTI8nT
4YxwBJjWignhi6eRWQ8CLRvg2BLA/nzCBF6jAl82QO7R/qS+6dXBd0WfyImFFKIT1NBWQ3Q/G2Ub
tEPj25phaAc/YnKEI2VmoPW+oxPT/PRHxzic9qpiqFxfEho07w0fjV+oGPpzzaod6VW5UEj+fGK6
yahJseilFPYyQV5X3buSokQ6wJvliThRoGCsf036Za8Nu8Di4fVffSU1ZU37rfdR2f5veMKEZkLf
jOFxwH9n3bBoYn/3UqUvO+G/QU4aPu7VESYYl0x6BlJErfDOUQ4/raFUyj9ZYWR1ybu36DbWn41k
LlujdFfQBfhyD3Grp+QRB6k3aZxCZMBJWThFW5ngNi7iH4S5zogq3X9FOl9+vE3aSZT8PCDy/7PR
/qUU2K38SSufs3TLIPkQ8PLLdZiHKveoZdSRWUyNz8ncEMBg+0uQJICACqoLYWM+VJAUiTVnU+UH
SnP3457kGEkUdvu1tnMp7Q5vIIzzouPNCP0btzd7CDncNR0OXUjFUJksjqTPiAI01mCPMBnmI/+X
w/VxrmrgHzvqEjHfXucRdiG1VPaihcPJ/1M22/ftYrdNVWoJ6XqXzhat0+qhoKm62cCBHYA+aqFU
D33H3kmoy6NbU1M0Ntpx/KNnQpTJaXbm3efGdqSb96QNYwFLPDIL6iUI1rCFINAExT2j9mIN27rj
J60v98lLGJRt75xBRlWmf4weo8ROMIgQoTax1xOigswlHwv8CiF1+IiDsxJYr7lncWbTKzS1o3o5
abBckUNOUBw640PA/jDzzlLDeEEMhQFooXp4AHfyAV2Q9wESLGQhXEgsp5YtI5Pell68zyOkxbc4
5iUO9HYh52FXTCwbBQ0Y+ZOHon4ETyJeV5CIetwiTrh6Hgt2CO9RWha8tHLYKWKUfdx66Lr49YXe
a0K6Tm/we9YEoMq1qZYEP9ZxiWxDmQxmuWAVhCZzN4FGNFiEaofBInju+l0qYlZ2BM48bV0CSdGx
6Wr0wRsp+RVoYXgWDX4YQl7M5kSHSHi6BQ65DAgQudyOZyaPHNVsMDgg4OUdozs2gNmbe0eGqc5t
2S4oMdvKSo972fD+XoF6F0C5b67H1aVYhqsOpBmDn7R1c1Tvx0SSaEGrG/5TuvwrF7d9veb+XVkd
RSctIjMC/xkoGYn5Nmv3dxk7egvsG61NIQQzol9n87gASiWoBVxQAHQvjBH0Gv8K7h/4h9GrNqeu
4DqrAiwmHuf85qfWxaS43bm/iU1DkC+kgFTNNmteGd3WLXpVwnJlkcj1/WKZfWQ/h8lpWJ4kRfKj
6cQsYB4uEL0nDFX6fCDKSwzjLpyClROlGheUA6d4D75X1XsWC4fzctBqcPXMzpvJLFTSgwAP86wu
1daczVldPFu9+BESr7Zb1DqoKtGg6dMd2VcpRmBmJTzZSXKX5q+IkVaYHMYeIiPglL8b3icsShaG
ChGGfwqPBrBYpGfnMcnGiD6hmrT5mTsrSDLocnd5AXM8GRdXycEXYEGMZnq/zVPzNCwJhI9Yl6pT
OtgqxoP2bVU/nRenyXsLsbRJ6HOUUqv9yIkgX6gRYMuDIkSDwYAfZSKIjkblfQE9iyLRoaM2nmV8
0UVEkbxoF1qinYx4m7foOSHxXdvXOT0Y3nkd4JbfQXFL2EJbYfx4UDlaPAh4IYQ3eh7Q0C1ukaJd
PwHHSt6yHecNsgoycuwlMyLAiN5p+W7bFSrb2BNp0d5W588TMrIhxU676Z/Vn6TEjnIgm92g9p86
OEswefrYvwmWD1vcIWlRiXMEnvzc+vnhSD/YY6hcnwPPes0j8KSm/9EmGw060AePY9xHc1xq2F/j
lcr1kS1Kna5Kr0S4eVhX1NVYX+Dm7WvYdnjc4tC60yFmV3JlYtHqlTpyxwTGJt6yRZYnXAKQmCgs
224zmbcq0iHPFP2ecdt5rML8wTdn16XZIQLeFzJIy/lePAUWpGL3/k+OuHq5iP7tNiRDOKwzIfnm
OETG4cJRQpLyTlhw2TFQ6e34tRmWzidE4nmHfGTnRqkt8nLK4STME4SBEAY7WYacRrHvgmtrk4+2
tFVH4mWpHep/Ig6h/x6IVWwprg95ppwU8YOxbcOX051pu0nh1HnmyBBTIq2ULZUEbYgaRGr8rGCd
IZggmx8Peemk70na2URINbsSTh4k02PoqoXX0UymSzCNHhRzltLGSGo64WQWx1wpC/6G04drVOQ4
+OvyVTGVLcyVQNFNZ/YFcttQDANpJCWIE2FSxM+mjmMqegrztywcIFzH7b2it3SVRLGrKsRsyOK6
eVPT97XvsGA2j+ecoW8M1IsuiWKUR9pVR9cwxF6ygR31icZ9oyrBOSUqfDvi3rmnVaYs0le+9/XF
cKb5eqLCZ6Gs56bDPwEdN8JOa2atzgboMWNmmKf8FbKx15gdee1vf/YfgvC22ePQjxVhuj+z0kbn
KnhAjbnExzEzLIdJKug4tm3bnNlsG3tDDun7DibdSOFMyKrHruqQD+OvLN4lb6P04s1wUL4NlAhK
80Otv+J1+ZpWMoRPLxxaIYsrynyd6J8eGZ5cFZKiLO90iZiirqkMDlvKEi1uWEIJ8b4iO1BrMOzt
UD/5/l/bYiQP2tZkokdqyyFkj2Nl/ZyH4XcfvXQBjnUil8uPd3Tbjt7jCpsQa+8gbvwJqJ1sjHG5
/RksWN8Cz//HvJWAVLT7aMELk74rVa7vOj4RIU681A1rzjgef6R9MjwyHse4o/L0fmcGMtT6g5n0
T1R2ItGwiJF0m+5wN3bVlC7XXBiaxbxGahfFneqnKxF/T7hokkRgTAy1disPTmjbydSj84X8vBU1
w5zS08TuvCpqx79SYrW1PuAz6kc39XJKY+HcLd1eBTD3OpY/5NuwAjc0o95VBIFcuzzUWygyUAIj
GffXPJgql2luv0vqY/2Z8UX+ifDGLR4L8bP1ou3dTPKd70DFNBHKzBj3+w8iU4c10VYAeumJDCTZ
4zW7+0Qx0Q5u8jKIaJFcWChOvjZGVU65qQwnK25YgaGWEbvOpVf60nACSSm7/uWjvHTLLGZor+Vn
Ov/qBfDc3L5OXBKkCf/X5itA/+6aNFl110cvP33g4FFV2hTBPk5clw4GeFL45MK8p88x8dK+gQgm
BZwlT6UylEllZQhiVLnk9wA+uCoIQXT8DylizkDMdGbL4bqi8qx3zeml27O4Gobv8ph5490U0BK4
G0TwUYuvmtM2SnBMJZ92FQ7UdwsNbESUfpC8S4k7PPXrlmfweBkz0VPYYCCw9XqUyJBQ2zqLwgyp
nibFtuTby4ublVpO2jbFqBrHTEQCdnSTP7p5Fr4H1AU5JmR7fufy8tlfON9UXGvc+TuiJ6NELEMg
mVlSg7B1kQgpqKepSs7+P8La3CbPR/3PzGSO9QnMSTrRdQcj/HTJLkq0q9qPTNv+LelcSDp4V5BQ
3ySsedgcSEqyM/36c9ywtZLGdSkbFlXntBJPa0gCj7ikaaofpm1V3ZVTvtw4ktBXIQkSKhenoow2
T3DRqIo8+EPlJk/NKaSHrmURvCy9Dg/zjaVjuVtlN8dG9i2YaGbL6mCVu48MqZTejlsdu3Fxbbkh
h48WG1qHMF4iYVT4glrePvDpr+Hw6XqEkJ20PzhGQ2wuKJ+A1rGpiAWo6DJfCIl64bnoQ4Hx85SM
5cp4Oug0Tc16f+xk+/qj/FCc3YiFFUDH7Keu8Uy339t4tAA8r6nTCLoxYP4Bdi3HUPNczGM3XXD+
btOSh02ZxHC2epZipg2pucBojSVltJize+3i1AZUOiUBVxIglYpiamaz417oExrpUtr0hrp539aZ
KTbzTmsXyN2paaDKtNecldxgASVfkx0jEDNGKJL7FDXwWT6NRC+jog5x6sP6Gp41jKQ5JMeKB4Sq
1JPzgEDd9oIG0xSy1Xu0i3dIAfZ8aCO+O74KTWSbKnEiyeKwbvZYa9osfppSIS7G8UtiwF7e4yMH
1J465Vg4GYvnNwt3s3N+CHfHu37vZ12xCi5O1exJ99/weNzNgG2ur5nKP8rAei3D/NPdtoBYxo7R
r35wAX+SDYfyyHOcdNPwqZ8pQKchIVksBuzo2GC2ba1bTP1WE7bePmh0z+WJuC0mIADR7JklxAgc
4x51YZb6ryDVdxCXKwc1rBcSuP460H3qIL9HWEKDOxn4Xp5UbbqzC9ZKTuOOao1rsyY7EwysuGkK
GjFk4eOnjhLTCYWaCbehAv/R07ziAoEi9TdWQ+eT3yIaL/VEFREomVUPpXDjNC3h7PIbCxsJqS5f
TW7pB7Y3TgK/KMhcuR3AwIwbvFu5ptnFj1pOFFooxDtqic1AkKSHqOHuxsjbd7HuXTBKJbXocOCL
V0UivJTWuyhJrfevprEds7nbo14L/UgAf2p3MKe1raf09iDlVGu/pKYuTZLj9wUnb6rfvbRE042g
YqLGQD6UlsGGLsty82c93m51EuaBN+jK0V91qmhC21eiojayAPlHqtX1j9ShlidtUpGaVxCOelEq
+2fwezdAGXjR88oDBGIwkQxewThJN1rDCToVZ0Z7GptzetZC5+uTd0Yi0MVwDbqQ7DY++qX81OJD
Oq5T+e6XEypXnSPEEWk0C/Tiw7ONOatkQjmdYR4W9GSEwkuWV8NLv2mzjPS1CRisIqp6+YZHjo3h
ipftVetZNVJNhzYlomqeX4yv5YiioeXSGcjelbwaVSbE6OzVA7/fYE8sCFSjm82+MvfXXdMKxIU5
JEbRrXu5ZpQMDfpc9bKfrDdzCe+ZhJztgUSJYiCwtpx+IL5yldCJ5XBXzzDNDWlWUYRAwGwVhpWN
1g0sYb+/rvoISFTnAUyHuDl2Kzm7S2EkQNOCUukc38vV3iaaPiyvTuitrmUSSXEYgpeoawknHnT4
cevmm6xatSCcrEm4jo5UA3W9xyPJAXXb2WzoAk3NfmmmKQNDz00gy7vgAej3dxrlWLV7KjqWSCj3
2mAmKX7ZU2aluxGHIhbSR+Szx5e3j+gjdf8Vsol7wKs4Y07Ptt/5l866/TyQaOL4f7oB0lRllg0T
8WYOxPLFLQP0Q1yEo+/9paZdL66xmJVTHkyZAwSgr2WhV1cY6wM1Jv684MoI6NJH8m2ZT3SuLqbj
RKEJRCFegeT6fAKmeOqOv5pEiWxlsM/Zt7Ak+vfn3Vhg9k6sWbtdPbH9HQGAZqj2tDs1ebvaOnPd
Wtcjpoc924sAxdOOBbD8Dwcqav+QwNI8SnvHKfyvWtDcoOLoZsnGGcHuxx6qky6gzzoif12VUU0Y
Ojy/jwigY8BIoV6UvNfQf6dnR7YDow/jZt/XGxxvYoL/yxOzDdCe8Fgzadtll2r4marFEXfUC3Ay
Yh3ElEYEbMqfgzWDgdCKvcRyU59nlW6LUseSMD7L93xHFr2//1w9NNLH+3Etlsoe1XaOo24vjlZU
PbOO3MCPrcvHXZ81oNd79tpkjbgF04NNekws6SzXaIdQpJaJ46T8k3xEQEbCcWehND5/Mo2zWV5+
9HFuHPiT6AE7HDOyfEBKo0OMq7nY8u83zoVcZEqN5Du0P+qDD1q2z1JczQJO/Z2CHfK10src6Lin
r8EHzm/XK4zzjHlDTA4M5f57/e4SxZtNP/aR5xv3NgVPZ5mvSc8gzKp0tSyZ/4L9MUTNSvFeRZB4
m4IhEoI4aZseowVDnggz1WAb+UapnlFDKcVOdZR80Ux6YlBQp9HLbZeejr8ThlHYzceo83Tg6ykI
IuCKnpLhpemCHq7byA4MJEDvqmfAkESOvi/t7NHQw2VQZY1SNE+BaBL1nYRvmZe4JhBEw+Tun2Zd
JnaGlTEolfbEli7X3X7urMAToVZHcXiBheaFNMQSZ8209EVNZ+57bdMAvAzIPUngeOtj3a2LvYkG
OdJ7+tMXIger7krfpWQxJok0KRuI0yPFq67MrOisCFuIM7YknjT35zEeBhEgFKE8A+Kww2HStzNW
lx8UHr6uEpIs6LbMJcgBAPXrlHTdgRm1+JRiXsBPRncyo1GuSp1Us/bBRQlJNzVg14BIyVkMQ3bZ
gnvLM9+kpQ1D26ntbBGoxUUsJvTX4f/G5P6qBMIUUs1DXupCoiWLvcGImweCQpHQtNFOp3XdeIBW
V+3+lo3IIBH281sPHN7KrVUbWZQvRefb/kKeay1a9NS2drL6G/JlPljIOYkrw2aEtzI91ovsPICj
lMquuORBLIiAMw4PJJM+JSMa8OE4+Cye0sQUm3s9iCefmjKD0aBOygIdsUNLMO7jbnbOguijgYgz
hb5yi5R4pjm3T41MaGznhSOlzqbnvUPzLtiHOkjVjoVHz8+VazvoLrgNSOLh5lpZLmHGSAU8gt9x
iQHNWQckVmaCbwUuHN0t5ZA6nEGU/ubcgQCal858sDp6LQ5MkPj9esFK+YBr4PJCOVfs+VCrERyD
ob3dznMOMtGfkI6FAOLPUrRLfA22ZRdLHnUOrYjJGoT4OOTYP7L/7v0WsAEVSVyBPmRyoasM7vin
jHbJvtXs4KAkcaSBVpZA41lEZgbtK3FjZoKYTIbCDfwvJ/77G/Az0iXhE5MwojxUy926jWm/hy7X
BUV9gr+8TP5yuGT1xl2d2XcG4/LTffn7PkfrT+giTr9t60iShHCrw+lKiEEKjps8xrd3IGJX5Wx6
IwURpZI+DoSLTpYaGN0a64pVMWR7t2sNm4FwMHC6X3lBjHmEh4IIU83pSHNXlRBdrhOTzcDUg5UN
pAN1379Lyak1T51rO4ZmSUJX2ZBsSf+F6dWC+0PWn+MV5tk3V8a73P51Tf7fXOkfgiSxvqeGcwSh
Fv4JxABcRmEnXMrNr7vsDqBTNdP7Dvmh2lxv+rck02xKro2JwQqD7BXfSezlUuQ36kGKzlCPHr6H
rDXYS0f3eQpMKLRbA9NjljeMknO3bbKn9DDZ9hIonhH1ldHunDvjRTzNbzBC+mngeP111RPgiEAq
ZZQEJxULN+pemI4Z40g8Cmfa3IcZOnmHvBWqtIA5Kk2jwp8Z8oshjfJVzdyR2IgZ6cuOEJDyXmYU
RDT71+RNjmBh1D6KnwAIMAavcOJoHWbOdvZ/300vLeVNqzQl8FVVdO49Xfq3uAL4Dq/YNp3mnnZM
+FA9aXwCF+eaBf9D0xsn/57K4497iqRBkmEntf8cEv5lm7n2XSyqf4JjYGnNo99hkD07YNqrlc1y
Ujz0RKslkkNRCkuEAYRNQ7+LWDJhiXUsSolrKdF32Q90UyRMh5Oo77Im2EPy1Xf0h9njgWACIRTK
WRgLT5LZoiqxAq12eH0ZOSMN+mdAu60Kd8bTVhLjOMqPlIEIxzGyRwqy+mt9UB2RT8T+JFIHLNHN
lyWWzz+TnBZ0YfIR2r/9CscmUodfaealicfLzDF5N2JQ27aRSF8SACOzpz1WSYEtW1zw7wSXmUiK
kXv/Wz3QrEvetxz2jk8ZHWRMMdnuOE1SAqCqWyr+xerag/87IzVxuFS8F7v9IeWdjtkaENIKsnXw
sOYaJJTSgpzJ8bip5skS+Ry24GHCrvEZiCBUZh7BuX8+buHy+ozDVO9wXYxfpgx7omKPZJdMhUfu
Y9sWKO1vKNa+kfxfg/pzi8Fe2byqZCArFQCULirAGfcyR8eh45A8F2ur9TWWTnqt0Mq+uWqbgXDF
NSnCiJ4wy/ht1CWK3txD5cTZsc4wtVm0ZV7nzrzDoVZYZhi5ZoesIu5Vy6pKyn97MfLVxBbv9Kdg
AYrB2uIOpsioUKLyEa/rlM3NNa2cJno5zkqApZopFhUFzpzZANa+DyWCboe83GiLWUFi+Swmheq1
RqU7VtJNELs8rB6SsVhv1mQYcC2FTYIgvr5Urox4GV/XEP9qUDHpUcLELORNOY8HqGUrR654g5vK
PBjEQEfjckgtiTGylTR8LsdWikvZ+wscZOs/RVOGIrdXQrlreEAfYv8OXdVkwNji5j/x3n0HRyKr
70SxUaafOZZUeocnUd/iIk7eK+DIbLqNkeDrgWQ/4R7SuQzWhZg5u5PyqEOaxii7VZatt93WpS9b
AX325eVhlQ+EeY33NSW+7V1PdLM/BGhhdKz9BS5pqdRJ52NtMl9mZB9an2d7IDzqqfGHkKklqHHR
EqwN9azoSvsBZHaXDKvlyX1YldjlsvA+wh9h2VbBt7rAKFH/4wXwEA+FiD3WobjvFGCLJfoBWIHK
kxiZf6yoN3s9deysHW+LF0zEatFyMK5p7TOglUAAxIwPPMZ3374LMoRNY1qTNvp2Ke+4G0Q0y2dW
cBcAYQGZWlPe5MFrebX6WNpXAo/Rlp4blauZR6cTbpvJaQcnxz4BfnUZw+rqeH3AI4EsBqq0kszM
jdL6pGkS0X7HVS/9QYGJxIciJEd/djSH2RauUTHh7YwdnSbJGRDlSfkz2rDV8TSi8tbudpeLnNEp
3bpQnRaqTxqVgS/jfMbWLovftRId8vhTt0I7P2idHiYAx+VZokcGbNm92pq1K58i/s0yUjiFLfSy
hxpx+BiNrrazZOCFQZ+sNqokLdKL+bFEdAdhR2tilqT/r/hjZb9cDoGtuy2Ah3znNLt0ArHYCI/v
NEh12kvXb8QrD90FoFy8Vs0oypl8+zbiG8O3wp7xVPOkKVmXO+VkBaybbX+2gBWsiiRBy8czUJfG
1IF8uAbNcGfuuOdBrznLlAoVdbYFbuI3ro2gY2wjteplb+0EKAWr1fQpe1e3IH2uuLCGBNgmkPPu
EDRJk5xK1QLvQ3ptek/mqjtVSWgE7MXeXkbk0aT824a3ZzFSWBk70+spnD3LSJcxE8vC3mX9i6DO
gxDPcASjwkbB1pBgcDsq/x13iCEwerfIxQhTLIl0QsMTev1QyqiZ31+Q0PtXf2WgVoC8ioVKo89b
NcHjXw6BHJkVGtQeztdjkb2u42Ybsj3IkfSNVPw59sZ/+LRdyETaE4GzICK2NDS9Esh5eUxUGHuR
HnQhMaMbzsnAYeE94t3J1TgEkcQz58juD/IVK90OIMoU6WBdZKCGzH+sTIZ8UnwKk6ZovKs2zi1L
CfSfTWpnDlX8Uo+sOse4wYrKQSGDUqwkC/1L4NmbGnkWoqUPERgHhgYv9oTHc2BsF8AUvu8A8vBu
2MCNkVOO/gN5Uk+NrXgpurK+LiEBmUHeTZlyVV2nJfyh/rzH+l+6+OXLe0GzpldJuKWXyrN8ij7V
wUUv0uVkaiQC7qoOBRdXVSCd25MJCC7GeIEB+PhePzVC0jUN9v0RodAl1RVS4InZJmWjKZGN1Qn/
2GmV+xrTP0w3MLT5n/BhxCejU5SnHRMZcVC7S5quVVXbqXJIk/3YbOGknHMJHWStvIfs1Ioe7ob8
y68DFYpqKmCl+jtSy3hXfk/sUUkiHWnYZWYF04yswCz8ISZVrs37gG+lNz3gGYjiAsLkQOHO9f1B
IwafqEtrmJ7P/9uyyNf6sY+/dCq3AfjT81rQZymXlE8Vl0DigL6+DMGDVazhCY2zD+vAudkmGWA9
Nb6d6RlDNvgUhFRqRLbqtGwGnRwknDStNqEk+rkDAqsQxnTvoal6hTohdzV2q+trx8Wl4curwY0M
ybbHf9CxSOuGXWdYlucozd+VPaa7tCSfB6drdtQDhbNFvKcHQRIr/NDsnGla7KO20JZ96q5Robw1
fulVAszZuMTjQT3N3TQr516+64mZwxXshCF0Ly0bE9164ebce1DxuMTztw5mgFVwLuXHxqPcj2dC
rS7HqMjb/sZdHf9GAB4UxAbOy96VRf77/e3JCEhNWAEK/1JEkRT3DzBZrOZ5DN0Mi8Eo1zC1eHVE
trsoyiw8atnEefs63CGQl6jk1CzeLoG8GJM9DMfw/aOQtdRytpugbLWwOE8zfwatzbW/HiNFOSdd
5Nj4BsHV1mzeNIo/WJUjr0wm4vRSwHHdrDCk2T+uHlXF/4H9L/2p9zm33MEQoh6/NtXUasH8STPt
xskdL4wAu+U3mlrsePB1GPErzWK2ItMTm034U89O5taazb8/IV6ugRYKLRZZ1DozGvlHivhewwaR
srvdY+Gtp+W+XFE1Jfre0LYORMUiyAZfnWSJfMIz9m5Fc6qaIRYumBP7eEMfqncnwib377KRF50O
l1yxz9vvmdz2FVzILDeaBlZme/RMUTISlHxxZ8il8W49n8qleo7kOzdX6nZgwxr7IogOWQKgw6Gb
FaV2DwxxxrsG0thSxM5MRGz1L3tuhFITN85UUXxTVQsopbRtRZLpexKZ8CgZ3jhHd8IP386BDUP7
CYfQKmG6jQ4B9NByPS9aZ2H+P3gLEWVa5fpFAhaj2hK0OHkuuRGlA6njIx0AWZvi4A0Kvhd+O422
4vCx94eprMT2nmBInYc20jZ0x6KAZYCi2eISyoIDD+47hjAjj7uOMlf5fzAXXB9XqFzbJATCYJCo
ihDgt0F2PCU0Vu0XFvy/PddNYtiCtPXmMgY8k73EYg3gpL4dF0GIFe1b8kOd8Hi6COkBy7yMMYO6
YFSHaeGcP4ss4S3zYwEXqhmA5DbodPGLBj99+kAyo4P9AnGw6bHjAN/SuD4fC8VTuKaDZ/zP7ETr
xhtybb82Xsvpj0cWW7ukqKbjFOcjMiyEZmq8PIVTG7rSZmWgOcKNL6czDwAKwxTwXoj4lcBjbiK0
uVxH9+S7/iggpUyW/peu3zuvnIGn0CnQaG8Cjx+aWorSyTm0Z2p4z2bWrcslyA48+H0zNrJGKaeB
YL8lwwvPfBssqE0Fwi36Vng41Bw7I6m5qnecUxKE+t+LGJt8UK3GDaWd/jex8ITtm5qfpi9SArZd
EiJKoG8Nmgd7mBqxLDm1KbhaMmUm/TJxulAf5e2QfKAjs3OX7jBViayEbnM3c7ugfyomkvIXS6Qr
5+hpDHCagXISvBo0c3aQvykAfJR7rhsX/CjFC1Q/eldYx8noDBi9koaT/6YUACSODUJ+CEiz1m51
oY87PbOKidWeeCFYLwkorAUD85vGdbc3UPQsBna+SMaovzq8wO39kp1GHoVfgnc9XtphtC0nGn0j
zTNIHtH97K37LfMsGXFy5xV9Ta9gV9SOzqBgwxpo0uYy/CkNq9THL9RUGVOSFG7R7WCQuIcLIXkV
PCqyYmBXpDEL1x1l1PiOhomwgZIw+h3Z0GPF/0o4FxhtPoP68IRuZyXEiG6VEfKBc1baPjXLJ3JY
GKYqT/Jk20qB2jiSjj8WIsGAvLyC3hHaV3dM3HxecjHpyDuimytCP6K4R/t3pTCBrnuCw6KO3Hmb
anAz6uIPaSpEyYC3ernqwfw512fQfuhIU6Kq1s8glQmqwaL+i2bRAyPIF8kzQTSqOn37HKw0xlkK
tlJRKZdiea95pLs5apdZs6KvippNDPtXt+XxpBamyP2MkEmY0aaJWCeJ8jnq1vT39U5n2xGNOV8k
DGHjobwPEiLz0sPV43ZyCo5cfRVbJ3rNBbmQu/xdh8lr74N/ofpwRD3OqLlE7an4hnB4LpxvVOK8
NqM3fUCHOELnpmZVvNASBiu5etwvkHGDaWZWNTH0RCPrvuW0vFekZVIFYUYQAfliS/Fs5L5VrHbq
O6dKx6NMexTGfvnP7jIrv92yeDwcbmwtDkvsIWj4Z/ENCJ8wubG+DDUFzyZShwyp9Q528gOU3Bnu
L60skVyCiCjYlzIBqMVxRoyVLC54i9IMbtwf1cgJncmGH2imzrkNVdmxZquAx7Rt19ttZm7Ad3Z1
hiEFSt04WEdCYz60ABNW7Vsginv/InP81LLKBhENmmsKxdjRLOZ49sB3cSGlef19IfItOaLa9rj3
1bzCXJ7gDS/tIgnaT5txR7L25T3VJ46njOKIvzCo/sUnqQJBt2g8RMJtC/mZBIW8VsLvCSTqXLl4
pIL/ATs4Z/yGdW8i6qaBO0dbrcJJDACwEHTgr2x5LmLbHk//qNKp7gSzEUn7xpeJyexL9tRNRNgD
5zHX8x9qICVtI6w42VKUUmgAnmoMCSOV7JPIh/3PglLVBb5f3VDJnxsSllg1bF+m0eOgjxGyxYBM
ZvM/A57v0R5opQT3DYOijHKK/SETqjjaHAfL1RjAovaHIv2GxsxWDXL+n9UpCwlqhs03TE0RXrdE
j7Oft6DEE8z5cFO8dcXoSdJfX+TvhVOpmntRD8Md7DzgHLkXtKM43h5/v+Om65JzXTHiuiuEkBgj
yl/l3ECrhlTphEUxrTTo9EEzpUTDTsJ6Q+CSlbzGD2qu0BF6mRgA7b0MxIP7jZuaTb3gYi897doG
Uy/nUMVcTCc35QBub64QSHb8lOCpkcJAW8iBG/r2Tx/st/f0ehPVpLwwq8j7LAitTM9xCb3iO9zN
9lxJ8/jLEFroTBegp8HMRogJICUSyetjt7E2CQzbkZAw4bJExFVx041eGt7JS7OdbQWKkv4gnTL2
tnyuLrcz4DO68S4ZKYtN5ZCHSfSl6mzngNJioFFMd+OLNVsX9B3QACCNl+R7lo5aoztWP2N2VnFZ
IiKGaY5ULy4HFOhixy4bT7JVq0VspcuRuhiSPvalNdQUwbRtdrXtUpfphXPLuDmbyQfon3i7LL16
g9ntEOEJ5sGdISc2P8IUgElhM94UtVWesWfDB0CQilkDmrWOliEQxuJxflhv9C3aGIrn6wc+/4FW
GdiOK3DIkw0tRm/DgMaxGKuenWdcASOyH9S+TuiIxEFrxEreGQhWZQzheJNx4Tag3apOmHjfclzY
l4EV8NL3mBZcTw9cJs6bOknOX6JE+OkFB7xhEelH0K4UPRuif4hxxhWkfwMeluFehcF1wITXnWHi
xfzyANmstsv4z5w731+PjwNSZ7KfPk872ufZAI7w6dy1EJ6MArIBB6wvgcIaPAI/xPHrQ84gP8Ec
AVKgBLYKxnTSfTMpbgMNoSvNRdm6Kn7IyLABEprdEHmB67zvm9lWXiD0ChcWZnKXTWSCifVhmtgO
cGonDa1TehQ+pdGvR8/u6us2RGLVcBsIyDbFKjEDE5spcNXSo244TcaBxeEkoCkO3l8jfqkSiruk
i+s5VeRSctYo4ZUxN/P7o/hHAyjFIuvCHFu+2uRPLcYTtyWbZYz/4IuA5YsrqE3w5SJb+xYbsYWl
4fmQzUiiH48482Q8Ze9zhc6647jRwcHuApinWgxovyt4AE6lRePl2YW9HtaowM0G2jzWwqgrxcS+
niiIOa/h4YU1r95Q8GzyOhj7OaJj0GTSn/qv8FdZpkmgYb1Fx/ALBm9jIUuFzSux/acgTQJ2zGCK
F/KsbBjUVzYAAMWhaChJPMfOJ8ZcowG0cuP8ZXCfjdhkKGqPrqgT1yw8PJypVVI8V6w/DV6XPb/2
SWfAoX11J0J1UJ8UWuLs/sM7BnGNGN6o7r8HOA3fMh3lGlNHpZsEpDDs3TucB5jS31L7OQklzjuC
Fgxv/5DjtyZyGlbvUPPmVW5I3wkjHMU1Afc4LJ7puaBcXec2Ev9ANtn5A7QaC7KHk1FiiUmHt330
Bi5ye2kHJBqI5ZFyRzpUIWqSKAMJjmxEXBZ/PufJYUuAME6XpIpbaJSj4eVOGxjVK7biV+kjATUX
rL3m7XVhdODTVP90kv7ik7a4+TWQNK3TcK0Y77enk6MFUA/LtkxU2DTe6bQtj33P9Nrmgz2QUWlK
UNsI4sBA2st0bMYyg9uZ+PP5O4mXYpJJGw9Ca3SdPxwc+Dj3aQjEc8YIb9kvp8uWDjoZzZK/bzKv
E0fG0jDoaBFXaa/JZACW1mBcRh/55aYv5lbFk9ZU1XJviJJmpppeGX7EnmC3pzIUvL1dq7RKxl5i
K734p/myW2qAxFbQ2mw46Wmy5+9ZgTXARFa5R5UBMDjLznNdE1w5vmxRUJISEpItIDHVu2qsgh/W
mdeqEbf0ydY0WDoZWu4yVMB2uVd+ZhBUYdLGyNhAlVd3NaSx/yhjUkBMlyLO9PVr3ZJHjhffyDMn
//ywj21vrgS+M5dR/eT66alepuoVOu3j4bNyna+9CpQJ2e/XJeolFHYavPxNLcJN9ljUKEm3HDh8
PcC7TvD9RuKAkFOFdl0pcfOTjyM2SjRwiqcG36lvemYL4b0KW5cf3qZXhQu1WgdE+gsK0+/+u5H2
9teczIWe0HIDhp9sg7yGq7X9+udB4SUroOkGjxZti1bXa/zdEtdaabsPo9KFCwCkt2yeyiZccwRQ
UfWefkcQGXdmkzBdGdPMvIoCJ1BnKE7OSqBrLTDICNwidZ3sA6ebGHS5GJHiqf4735bCOy+1xL18
tHfLVEclbfaz+2xwO1E2B2DVhtyNwCBQMGwolimHmemJx57Y2+MuF5JkRZTqjm4TsxHah9pci8Sy
a4lEvUXrsdtGhMFh00BR46RSjQCozu7oIxgwoLXVZ1HE0aIjX3wxlZBP5liO14Xf4J3T5OHulV/b
Pie4D+s7wT+2kuCLPpDNjOO8ACK7fIQHcj9xFarY46JPDNKZK95VMVDPhAu0Nr+uCwZ/TmebMF7U
E6tbaXBIHZuL2ThzveRF/X4Epj8JHCjyMgoOM3Gx0yCE0w7q6pZOy1GCHhRdAFGSI0NZMjMS2SUa
tuE7xvdKdu1zyS3C6UhC0xb9kxZ4AvfgoiFdqch9F8EKPrbJ+KGHuKWAxWO8Yx8b0WJgcV0djplN
JbOrrfE7T1WR5o/B+gdHi+V6Pl4mtQOXylvoaYvN3eCy9r0ai63IjO8mn2PkN/kbFvapMMWm6ZTy
65RgcEoZRBdXxKBEH/mDei/DfEHnbRga1fEdCsxIGWaLCAU9E1XSc29Bh21meY02UO7jmee1EG/6
v99mTP6A1FY8QJYwSRWWX4oNPd+LaxxkBGFql8qTRAIpB71d075ZY+lT9fli3szFl3UolkhRwiMC
+w8porLexsOOHT26AxuZIUv0NTNnvmcDHa34ca83bGjljJKhXYpXbvn2NfIaWaDAbURheaJCalDA
V6jlwWpVqCYwvKRyi6gM5NeKNiVA8AxfByotdrWAchsZfteaLP2e+6xBY/d3rYFbG9sVSnRBCfKp
/WBX8YVE+qbJrhVMaqjk13ieur9M56rDWYlv7CPgq9+4gxGhyj/+1MvVDvKRTJ1Z+K1M6VkmLg7C
XoMd3uMSx7kOpHe1O/GkiCTIzTBL67DCa0bVNgxcTErHlDKEVIkLvnMNDuACrEgEq5pvH52wc+aR
Z/1tzr2RoDplpgf7nuDGBj4hEX7EF9rb3i77L5gUT2XceN29vI6wgeljTiiT+E1cW8WxQBMySJEq
RV0e5QbeC+iGQ0gxlfBiOjQ38n2r1koEAjhUR+hgxcudm+iV5+5ZmP4pKPCGnBrzVYQ+aXZfbV4g
wXPXp91RodTM2k9piTS4sVO0z6XsSyd1mCxTTNkvwyk4AsNQOhHx0k//aJ7q3LUmDaGXziTn3nx1
y9nUkTYyOb2Kvzh3vbVIsxoK4bq9Ve5p5+136QN53/MylDGYDxDpA7nSWqAk7dgcV/7HuQjyRRqR
nSam9hmYOIaOUI7BtCD6B42OYVuYyVGp1alemCpZN7a37mLeFSHYZqEvlUmIUGXln1bs2esd4nAS
/ABLIxIiNgA/uZOMuN/3OC/4JJUcuhJGGwpGpwrUonOSg5THuaPPrA3YKL417/p9yuOBJrT2/rwy
Y1IxIcBPmyp6iFdC2OQ+9c0J8l+So9e9LxbCBtHfrY1dH/57OHr9C/PgiMO2rPIaV/eRu5WudZAk
j1dRPsuFUqDVBHBjUfsE2pQFcbp6kY37ze26vLHX+9icmXogA2Z20xgvnMH76DgK1A6JVRUXYYm8
239hz/Fhvbuppls7bro82iFfmdGoBuDjbu6Dxwinu8DiGZP6HpD4PTWOrBkJ7yg6+gq/8NlveejF
mSY1nGgTzK4PHmCU2NY38sDLFYNkaCSlSTPZWse5Z4UK4cUm4QjWT6J1yWiWGNrp/e+iBDLo3pcZ
EGI2QhTb7VPHrWKfn4PmRmlDnuLlZgvX48RnJu5xhlls603QCpZ6r2aXWAQezhAimTpUsZcsi3/J
5ndV2smJeuAj3etIVchX+yunbBYmbUK9sr4PeszIEKveiddyKfEZ/sLaSdT0lN327ZivYseRdkE2
8XTe5DJP7A0PmhQBnrr+lyemf0Z4E1HRityyEaIRhBI3uTMujTAQdo6BLqrKMsQxvSE5ngav3qJC
PE2WTliMLfI1DiGCCylurFWCNwsJJiNuLoTowvMvFmsZIuLyQnmjj4IloFGSFG+tahjABkH/IEQO
w3Dd1tzzIV10H4Jj8DMV4OWoZNPBivHJ0gmLSA2IJX9HpPPCZOiM0DlLqcPcZp+U8ErwqTUe7vwy
XoGu9oRrOStv6ltjQDt0on8PkE3mpfrnAeVMwaF5WGjjz/WiuwOkZpKtTi3GmJRMEHkZL2i73ADD
9vLYw0sbZPF0dv0IucBb6g/6Q9lvyRMkysLx5F39gxRsd3dkSbir3zeWQaFD5p8pyp/pFjEpbvqK
i/UCcSeDCkW7fpNnd4fMLkbXmvkbi6E3QYtrwVOHEMRu+bphwep4pOMkXd3YIoTmB7uGwKVqe/ir
vLINDd3PWJDqkuvcFs/2v1CzRXwlCZQsNo82vdia7+mm6Pms3EctuNeCoJCmDKQ8J4lgMG9LWRfT
PBalNMpfNx850iDIZcRPN0UNktNWCFwIV8Z7ISVpli4Gid1LKpvKMa5uNQ2/tHpTwkif+TvZvqbF
AMxDWDua8mbTJ1rwzkpugn8LAxz3Jl/sSqKZIXGdiYa0GuCFnlckGKCi24XLLUzxV2eBfBXRwZVD
U2BOnrmB9dlcpjJUe3metLU3FZZnf/W1epsSKeojwygIelc1ofCLM+DpPbfgHH467tT+BIyI/3zV
H99sp2CLokBEyYuWJsaDdt/wyjChGgxMqnyc4KRQMasfouV6lLMkPEGiCjTXk1h1FEZcF/AzTCdG
vzqy+D0BOp0owm01u3FYTtBYpNK6u80oXP0WOa3O7/x08IyJk4R0F3owLeyLHnOvpkCrNXNiyHjk
xOSGRcEmqwZw00nKVh9Cizdc5APyzs5W9/QT+SbWIpBsJDldqOZX9xvqH/BsHTLDCG6OQoXCLWDI
E1e37CG5k+rjMJK49tL7PDFJ4bfOsRktKkVnLVT+6R2DRTwXBlky6S4JPD0KFSnjusGbfzrcjNJB
O9TCZKJi7OrHZmSY17onh/jM84SZ83tQ7wvkTZa/2YebcGNU/y7Ym0pkm45J23QVz6zqeySv5uDp
z7tnrRboTmZyvz57j63syxmeVQ46pE1jPbbjnPjcWyc65yG+B3I/FYKVNnkElxaOJFuphS3L/gsq
w2eRKbJa6f11T0QIwq8IN/YKfTCZB+IOTYnGxKitM4LN41ALYXtKJO6ytidsSA7SCWrLqqTBX2BZ
LULVuB/1E9YA+N8YWwStVtRuhvPgPUigVkUo6aSiCxjU+scG7ObQJqg/Q9b2j0OfGicATl9g0rA0
fJ5+XLDGjmKuQBI6XCNFBTlelSivOIcOFpjLPFk1bruTxMziC7QaKlJKbfU79FsCJSjhHWL5aL2P
kGgLx6K2RwVltu/2HKGP8Su7JZ1ObK9AOef46KRSkk0KjnR09K8DhVpGZA5JJQcZwxn0+UnHw4Pk
Et9VAn6pBZHJbHPlOZOypn7AYbSYgnyTZvU6Qe+vkbatPGhb+9v1xp6jYx2Vn98hPb3BOqWSYIHB
terXgPCe2uChiXLxPOBpZD937TUw+xHSxvTLbhlDLPtuK2mjEGHHKnGx6C4amxm2hNwk4zYL/9Nh
EDI2BA/XoQhpIYMPTyWpP+/cMImN5eUjkILvQOwO2DtvujIFbw51oPRa4B52RJlQHg19YBTLGRPK
/WgdVB7n65r5J/4v+KzwFqn1vhGzjUuWoWjHBEAfxsgzJ7OwYUvIh7XPU/flHntxEDlXIX7gmp5p
MgKuvqY8Tu4gRtnN7mX7/Dk/aEdgSzNr2HN68nCHWoFd7CLAnXDJDS9bUDCKP9B2LutaIlx9IlJA
JsuRy6Bp8GwMD3eSxAckMWskQ2v4VD+bjFIgiPCinNK3e8keZw3rby95DlQmVDrEILoS7Ih/mgec
J+I1W7vzG7ecokTk1PDalWBlJLTvfkwlB0/zCzBTJHgFkPPhOswkgtWeHGGTFCCpaZMS+HJ70kwO
36o5FpKItnz4fIf0+jKAPl/h+w1XjzIqdjIzvZNOujYWKHaEbc9eC1Pc6TWL11kT29/SvQvMD1Ac
+57X40poIzYzl7t2UTi0KCOV/Pq2I71YdhvkGGcvatPp0NibrZj8DnC2l+ieBv9re3oRItZtD117
iv3vT/DgE1haCY9CsF6xXYHoiG1ol4TCAtJux/tK6eihVO+h4Ki7h+51HdG+p/y53paukKGB4Cs9
CyzbDTPXNAGZTGxG2TZV7+0tkImpdk2GdNjpDjqKKLeoWFPuJYsYcuSaX17PZvEhcMbxSUxMwO+b
cnIp+Rwg0h0yjovsvjUifKHn1mfG/lFoONeNA/ZFuzTFYjkE6zz4qu4tl0DIg45muWCgd2tR27UT
+TJNlY1DKYPGBAxDee6S2FdwBFvVmyV4iMVr6b1h7FG/KPqAM9caUphMwb/9PPmzv95YY1lZDPNx
SQLHEXtnDoFDr9c3oHgAVoITiNfgzfYyLr7869x6oL9s75z1JFb8YYGPrcn9cAjK5GYA30mlEhs+
+Df+dubYgjK/IiT0c3TuW/byRPtQitsjucek1JnFNIBMoyp+B6KgwGyUjkAA2pZDKERE7hYP8GLx
XsZh7/sO7hoMPzE9MksToYuUSuKBK+OTtiQYYkGvbvAGObishXO1BDuCFSMYNrlGxV31v37A4oDz
aZOX5mMSvYsBU9SH+FhSIy2r0HAw/p275YveyV0NIXBLIQUy1aGhZkIhNzJTNhtVireZ99X+ynuy
RBvFqcX6M78vaCAopw3mepxKIgMKztw/dFi2BOhf8EalEdAtmUSy/02gsYy/gotZqyyalflVUM2I
J0aTADSdyI91EnnAoRFIkPBPrH1X+pia/wHdwakJGGtzal9p9uhs3BlfIObh31Tv7P3lBoR7TVKG
5YFyPwKWg+7Rdl80fVWnw0S5gtvlxb1yxeC6Sg6H7r4g8KOXfRNmAS9HJ0GQfMu18f4XT/S+Tt5T
v082kmSx6GLgdEeraFvEf4pKXCwCqHKMBSjJmXUqCQgBEnzpEr1lOc+r46iqkjuWbktSO0PrKuN6
29Z2ZF3f5HRRg8kyQdoSf8OPxuwSStBFJ3I346Rn9A7h97EaftK8M7G1lMxQ/HtCqzgrUK1UbGIt
X7HyDOwJN/jSeRCZfRohfakjSSWk8GQE1L9YQZQqL9oLiMvmraqD8ErVLHZcihniZUwAPKoxlxdp
wIAw37zJ/n6fCfOFQHf0ule2TrMWfDXn5fEqhM2GBYBBko1qLyURZ8DeHKi/F9/7kb36DiGKy0ju
AwZZ3ob2ZS72JRCW9r0aKMI9q6SWoi0GybAhzdKbxEr3a0GrTEq2DcllHX+ywTmQkb/8nU7tIKH0
zxWD5EWJ6Kc5m61kFLpwuJJ2IFuwx7WjiuOYGhWT9VlNzIol9HqNnhUQG1H+R68KbhfVZtT5BWdi
orQV40xOIcdtcCMGLrepNoTHGwCqVffdqhiWNew70okbi8On0DfPDcklWu80ozZ5XhqA4NEEW9Hw
Z2JyhSnteJKY5KJsTupmR5OE3kCUmKPiTm1ltCMZeEkpB7IF+9+3I9BaUR/Mh/C4ROI4vAaxM1y6
6dUa1Xzh0UGPsq0dUOMOXrRXV5FsPFYxFYhNI55SUG6nJnh7UOOzyj7M2Ru1dDTH7LKLTtBtr4Xc
O7O0qqd6IJHswaa4+e2pF/q5adVCSOJRb3VFepW8zzBo46YjCfLbxC1jfkbfLQC58lldzRIqREl2
WwQ+ZAb4l/b/iNKMg7gLAFrFLgm7VjMQb1z5vj5TmarDZq5Ujmm39sZhIxfaqa31kH9MpeF/JCu/
/8mYqharxFy99vNKfQDN5zIzWmfm4HVgHoMzIDEtn1IDYJK+LJQvK3ovHRLKSXRnCupQKONyUYdu
jH72gFg40FCfkaMnEzq1BWnbYmhHfKH2hbhEaPmyFnqBfJL2L5Zw2F9NwEGoLxXmzfM9KwA0zRJH
tIaArXDgs/E4rvzx9ttYIqz+V7w2kp7NRWOBn8MZqIqf4m9sZTceRxUDl23NB++JUl/vLTy1aaJQ
qMxDHxatVIanyeB678AaGaIeTJEbTGD8ZqMnkTqxsRgZmEHP7ViM/0DAmS0CisYxxcCApqKvlLEu
dehb1dwXUYe5J6aadhYgETwUhFQOOwod0RCNVwNx6IWPEdBzn1uwn6+UM0Fx8gfmvIhIyp1b2RE/
r18xUIjlIBJueLJPhN/kzFdKgyBgyOQ1MyYoLMewQkvB3eIxcT/o1/jyTQKhyM5ys0/zV884OLK8
r75gnWBv6mnAjR+mIlyImU+Eqq0ET01lKY6oKG60wqSYQBurj7SUgF4pLGWhotxdlpAqVmtLzNQz
CQMevMpPaFA9ZvGPs+lsr4elo5RK3eTMgCS2tXCdDL6sOB5HTr7d17wFF3XBEBlvTIpo31ECyOyC
suX3OzLOjna//D4GdhJ9ZDrEY7yOkuD7YvISQovt1fr2Z+7n19bu9l10r0AdCYWJMDdHSDCbsLbO
Jub4Fm8i3ixRv/5bLJIza6xzV5SJAbTGk4etwk9iEM0lXHsqin60+B2iUcvx2BSjW6cDJ27PA4Zv
KuFGE2dGWQhgpcTB0kk7JYdv9EAIdOmB4YfbX3pdR0wavwIvTULyf+pIpoDV6tHytCrvizOj7F2C
ttKqMP/EpW73dOPt/ZfXBQi/nXcfKrTZEwJokaTzCk5wn49aDWtf94din1jrIrmo1oUdvsShQSMU
KL4ViMXAXvnrksf2zCcCwknVoVf+LpgXv6BsWhE+aD/hq3rRztMW3IY14Nqf0DY6My9KfOkTCa+C
3eguMC9Jex6N29nvP73LQ21xcMqXb9rkPebgBE02J15laeeNb2ilL/N/ISnO4I8Xuve7TZPwQ2Si
6s0o6oo/z5UxJtsUl/UXhz3yEGgVidUri4lMzhR7jdoGhgGGZFkGXZJ67smboOJQQhbAL6DYhBrt
6IIG/JFt3iPwoPRoxCCn+2t9dDffB9BkMdGFjxA6ysjUN2ZtmlBQH3MQ6VHHSkinmJ0mT/UGFiMs
HQNGk9d3Adqo7JfSB1dA0Vu25+GZu2BNwj2uGE02EhAMf1Ii6pBxE/XXnleO5SCIunWLyeJMxZ9z
UUGU2aBTlagrdhL1tP4uVb50pjn7u1Da/l2Xbxkden+6W+GjuGKiCeHX7YrEIYuJrsIZzZv7aPAS
tGjfvnV4PxJ/syUCY7nAVK4SwKq93XAZS4HO2dY6Ed2Hz2nH75DuZatqzZvELk940GBsyYZUatnT
2y15sCZaWgDi7pPaYzeCHCu5Q8RqrpZUVRFSCZDrzKmDxWhBEi6InbQ7KrCzXIHtsh+7rbGhABNu
krJuLn/vZeaQ9RwF4Y9jyUoVkj+xl5zIiHV/CnzRJu4IdEhJ7Kll1tOQXHTvJmVX1wDvwiYj3/Ol
IR0A0eQ4D5MKwyXxsGA6Fk6pmkDZIhvTeylc24/H1zJp7ulfXEFyWQ9IY9d9P4xrwAC41LHdrV7w
Yp5Nf8kO2tyUaJT8iZpC75QU9jiyq7vwroCCsgnyCh4EDVEYOm2BsrVbLEPo1A+nIdq51HACXSlI
GDE4bhmIW5qFTtvw2kxqsM4js0kt2rJtJgi7pJmxQBqLn2EiXDhivc6JvRx9HiPzKzrJitbgJQ5U
x2HtP6u5cuOnIbZSZvG7nfzZmTIVgNX+J+2O9c49goUaj3oa63Un5TgvqP/IgB+s3F1MQUSXmP/t
GvUN68wW/oYc5IYeUr++4n1r2PyG4X7ZSM9JLvsVp3vMW/Qd9Xos59FiOOxmVWhlqtpzP7NkS/Wp
j0MFaqq7PqJLdTgQKywqTM+0CrSolQo5GUHA2aUiZ/sgLDKnVXkVkCRi1rCdJCqgOjZ2L3/Qzj5Y
lVG4eTawa/MKCA1j/q6Aw/UUe9PwtZdVofEYwqLuRGhBUcdlSJCa7MpQoAeTS3/8PwT0zqAtejNW
sqx0YgpV3jcMOE2kT7vKwFSsIDPhYWXaDsbCvvdKRD+7gDYgVeRKJFQlVfU6Yq8OdVTTAwoN10os
o5DweJaHIKr8hSisLTcU1ivjiQV2S3+9qwUEf0lbnV+KhJdetreE+X3DG+p5m9rjInUlw3SOYRVl
NXYXv2LII6F16c0dm1k09ooJ6J08oUauQosByxA7sUUGZEE2F22O/zelVpzoZQa6d/IsUlb61Mn/
XPjs+WmLNrkkv4JL302xY7j3H1QOKu5pP2SA3m46hVSs87Un8EOq5uBuWs62rBCRFsSaeTMwUaA2
M0viWovvItkkziMspz1jDE+0fz6C2P5doDXyBA38DBxoGhP/p+z69/n7YLtvcvj6ckvMtkEJeTUc
aQT9LDix4y6mLNe66aLTGsTJ3dsKvKs6N7AxzQZ88hYhQic86suSRBZLxTixob1q2BGSXl5PdlYW
XtJkQoPulJgZh1C1Q00hVTiINsmyNapTwUW13cGTZ1FPk9msKSuukwDrxtoagek41TDHoT8lj8NU
HtdLVwOKelKJ5K44KklxA6JcVQSXi0qhCORbpK6YSRGI2ABQqC0m25xroA5Di9VlcOqf42NrbEXB
BOMNJhT+1lOeDtoJJkJaUUWlfO63BxpfCMXxlF7FHhyan8plbPwBvZ9HpeUitpT/prCvSuh0coIh
3Y89qOKBZyBNS8e4WjKCwjW/dTGQiAkxR+Z10FPFoNlCuBORfJJr5hdefR1tsxPbmlG0oCyvML8j
9M0BzmS+k22l62wWONCkwvtYrKN+ErW/1CfRx3lskquc4Kwc94H76FcdLhphE4vfqf8D6JTR8/GZ
eXuohIjGo1s08uf+06cQw+gf7slNiHTwKBi4lQiy3NhcCapAVNdChj5i4JYAMc5WahhUc8oNlYR3
vruWtJAlIqOzZNgX57cSy2kvj/+2atFDH3nwXbMGKMXAjn4qtu72X5HADaH4KbOlL0TEIe37r90G
DXqEX8OeQpVJAa2EA6VnYOanPjbVmUs6vI0LAkv2Z/mnXmpm6rtB6aCwf8+8eRnMkG17RJioEsuF
T59gyBWIOWXiZ9kSvFXVnNxHiedHdF7BTaeRZobBiSsGdIi4VvoACfmQwOmHjQek/nOIQliuvwL8
YRCijwZErYYIxyoPqxdUXcUWqGfpTFZQwwhJSq1499tM0uwuc9cBjLfT4+7mdTGvCMzjliKmRgiV
Pur4VDBY7FzB4ufiYhCGy9qFeuUK0JaGfj8vVjZ+OSkRiWK3BmbU9HoYc/76yTz/eWtaa1xCwm8Q
f3WfAm46DdN6zIS7+jFfB8QdtHcmcIERCwRQ/1FsXNxXyS0HcHEo4LP8NntNkRBC+bKCUnD/1X91
xGZo/hnnNfHVUyUOos1QgWdy0j9SeplVQUlsojUGJem0hYIMUVx/e4SFTFu+JNDE6CWIzMJ4rWal
aBJETpXUIsoDRYYvfvLK6mZIx/WdGAi/qLXX6ZooIBrKA0XGBbhzhYrWLQeCQSdnodFuT1OS6/Sa
Cgxq3kE9V0RGCakSDakVRzZPU8uHfEgh/f1Boh65xh0mOX7RIWuCwU3W2RmIu8F3/gBebhCRMR7e
MESErEwtnyvkIog24UzmIwgq7BKvuw11k4vP33czvXszvCeNmyfk0UCKOoelZ47iOGbpMvqNXYd3
Z8nwBSMqiYMZ4zi1EO0/DiYMKX00s8k093dkGaYM75/Ev7U+qWW2wQ4WjANNMIgAu9/+DVzFRPvF
OAivMbS+uUc4A1D1QMB2PafAqpJeQ1HKHdzWhApmoiLB0IScgcXWumOKY6A7kaWcJoUMFV+5lDe4
/WRt8DAOda1AblmSnhVgHTJkNSXFWduKY14nk6Sr9n09QjkH+fKg5+No8hy1q/8gDwXTT5SJb6Vk
oiYz5YJyQlZ1hLP8wJ9lgpwNIv/WDG2g+vPrMRbn4dMuVp1DinaDPe60Z8KTbds0e7MbOtTFPgGa
v+rTs4rmP3ckoVUZtldGILFnsJbvHxFEOg8vWq9xoXsLdIGVNskXP+yaAWrj+pRri+ZkG8vnOFQg
H3hYKIxvqrEzAjosvLngWcZ7SLqsMdac1gw49CfCSAU/YGv6tRXqKcbwSUDp0uuKvwgq8id03wil
EnrU+7vwrezh+KEu6bR7uFTamZej6Us1E8utfcaK7nUd0gf/OLMrNm6dBSVKsVrvjJ+3Ez4hYDY6
KBWXP4YALKxxnE0Gyzd9/DvrP802UuuXpaumyQItofQZtQMF+nckngBkdNtJgVaJ/yVrtMwf7hum
WKcgbHVCECE1Hy1evWzawVf2IeUn11VB1Sd99hAB61WoDrQgmOuXLCitFrryO9WtGnGS2N0kdvfq
RjGYfwabl6PDUwRzjufGCJM4/rN6EB/kNoh7fRH9FQKNLlFyvcAccueEP4PfrW8D1NRyDbIJDAIs
ifU+M4nz5Rf5BWYKCUh4djKE97HsB7U7CmWZTAblm+oLZVUJT4TMENsvZNfdJsl+AbTFbkEZyPPH
ApQyqhKGVpzC2gkWeMDB2HHYsFdTeouzA+NJHBkLUACYn/o4MZdEnIL6KTdYxs8Q+Xv1bIltpkNz
0F/+PnorzyIY4gNRPcdO9DVT9XDcqlC9wdTwmnajFdmDG6QT+2DpddI8yTBDdMWoEihvPw0C1AIG
ZM6SoRBvMnXQYwEoOzEYnCshv2//k/coXwxzfJE6lphzxPBxKjiWCTB8JoOMvxK1y8sUVv3ExMBl
j8bxS09Tc6fY8yxe2ma89v9QJ9FbQfc5ae1fcsW1L4isBSCXWYrf+xVrAuvd5DBGyGkZUVaeZb61
y8sJ0JHJME6+9eDzGQKp8/yAyM/bbpA7myyMOpujKbZmA7nQonGwnBmLmCp+D/GZTF8PNAxXfo9/
A5u2BTzoW3giL+Ain52V9CvK2yaGbtozy1veVAb1ii9rOVG5uBiBEWc5QtYAqgKIKX4INnF1ptEb
XPpYjevFcL0L7uZ98P40PfmBtJrk87tbrX3nZUPumaCTYW8uWLAs6zcoHaKuKp//i9Nrmw+R5SKI
dfcyqX5Kw21/uFIn0BU8d+2or0xwcayrwBYyRQKNAoXD9BnkGYjHZjJg6GBHnaitxjcFdSKotQvA
cKzllep4QvLWOs/HWq8i79VJZeEB2KrFK6jMaRFOn9EELrcQbofh8AthF+adhBRSHp2wDms7stgu
syY94PUjEtvulFzutOiA0lfTttWIm3roc5/31dmZIgVKk0v3zamuR1z848R7SZyh4clOeJeQp4uI
DeKL3dxk75SwJIOlkFa0rdnuJs1iFClG8SDpz3OReJ/UgR7hSJt3O1p4FobjTZVNfz9zAX+Cm3GR
viM4Tp9o8bhcGVieFYnOmxbOWpA4OLXNuWoULv/UXiPy+JPzT6rLVWIpxQjIpkrG+zwtJ0vZ0F7a
QIYlWMXuUGOPRdlLEz7sYdHjs/1vu93ZZ+ldrbq+yJs7lXkuSSnoWOu6WTBcrINFZqGWJ0zv60Al
sb9bQ/jDQJIezmI+SFGiKUYHewaZjIohpE2tK//U2Y9LutpdL8ulLnSKealivjgvHcoaKbqBGyp4
oPDSPjIYqGrwlnkXhfGVBoKRzcIpzmqe+przu7gDE6r2BRukGkgbd4l9VtB40vHsV8GiE+rMwJz8
QnGh4v/Pwx5koE/jpmDW6J9IzlKYK+MsYY0FFZNJJYUBjgwLVXy34QGq3FF3l7lW10WypnPCD6Fo
6QG3zh2T8S6jm3EQ1dzYIlw3X22Hq2EwiGasX52AuG4w1VKL3XWPQ+Dnn2w98Jc6tdBPGOhZjPAl
vVFAvMtwRG3F8Ns0pjGS7M5wPcrnBjFSsuO2Annv6lLHLJBEnWU3gwSoBztZHDYpTf+AdMGX914u
Be9wk5QYnD6C3GPsPDs+buogUhJJhzTIs63yMR5vn+0Snr9X70bEDoDe+RJ4lEg//2IYSk1eTcDd
rzZ262hjavKO7IqU9/c//GoYChUwg+TMNYW35mN9nY4bRIjoF3LfUxIEQpVkFq2K/5kco/BB8Jbw
FwSZcXY+HHInRO2Mh0zls+3cxpnU8qvNC9pg3Hrqm2BTqvhuo81OVgFY7Da5WSplSeZhJwvzhgYR
YmibpAaziipqgIRP1foh27CpfT1ILvwdbsObH7JXjSHVRl7T5gdw6UBjesgQX3VHwRJMGQvZ9n7u
938cLXSevPetGvtWB/qvUpXT4tM4OWFduWr9KlnRHxuSmUwDFFgz3IIFM5POuW8H6cYSj6W4Y7+j
CwsCUz6zsw5+JGycXVoXFlMJYoACqxXxGpcuHkckj4XMapTcdNCYRWxtxNz5RTKmkZGlqJunkAbS
Uz1ohn8q7bR8YgCONQNsNBZdya9+cxxKUiyGACOkI1n9yEyyf5CBpmOOB2C9Jnxv3kYyq5br+G+w
FNi/tAXCRdxpeTmxwLp7ox0KXzJ03ovS3S5egPmUOdcKqBgajkFE+62pJN5MPu5CzM628RMXobgT
/FH2ILMMM67UMy92lGHWWN1NIyh1nJDkEqnco2hqVr8zSHJfH/Mc2Ajdz4t3pVcMfcHl7NoF5096
h371WY8VPrsvik8khcBCb3XgJOr68bFkHeUbzzwbokijwsiORRcWI341/HTdoIhxpXMviWEXfk+d
SHAPIZPLRxurADIzm1NCk8lQvdueomk3zu+WjNbTJRNTzUQLTuyzQLuHEb2kxG3c0S8ASGSIY/Lb
UvrOMd9yisXoXt7FrrqJyq5Evzv9Q6GrIadbQiVlRqFIzCGJl7G2DLsNGnZ2sf6Gk9vhDrJaTocp
t1TXrgdpGuk58m8SPGYVa6/NabxMoRdn9+eHQxD/DkYaAzeeOc0arrO47gqOU8apV5GZx5a0gh9s
dIvWZC22M6IeozsJ+a5R42I2S068w6hdpC7CRJmFOPqxyc/0Dhq0QkiRN8cbfZ1O2B3fVBIajV++
Vb4v9sro20RnACVOAvsJRnPzTR1T/bfwEbOXUHedoxpU0DalX/Pq9nTa/gL3II8ffvFCpAiTNTO+
q7+FJOyUoRmE9XlQRuO9TudsoisHdKI7Nzfp228ur76LgvGCQrA7WOB2np6w0wSIT1m42Jm7crSu
PjBsUqMDK0GLcNBlwSelZqM7/PNcIPlCj/QhqYEbWCclqdyz43ZBFJvlzYjwRx6Rt6U3lTZHlb69
9keqBNtDjqdH5QYsbb/QDN7n4b/FEgjfCKevFbovPreRnwNwf432Q99ameZMCd/py9NsNmH+WgRC
4r6gFC4+SvgGtfjcD98d4EsPBk9GHxnj2Lakn8p7N88+PV3DZXPfPR3VtVpyD7rIl5FgtSwLTvG+
vWahFyDKhRxBgo4tIE1YHfIWCKQN8d5Xf6ZRMmO3mRce2mRrP/wlXpHGKIB3qkS9OlfQu1SfSTmK
ogRx6F4XOXfTWkICzB5VIAWx1vl82uOvfVKFEXlzlm6VsJdznbIZosF1Dny+gkn1GAuDA1rnS2wY
CB7jq6Ny+/JkhaqplTfkjCnZN5fMabiSmD9gccMYrnBmT2dfaq4vv902VqaH0Hv6wrkuBVulVOWY
ZptVn9VrFPg/SiRBvoWvEd0bjb9gnUBMGR/YBHeywyapoLVrfDly3C77lsfYv6ph+w6AooJSP1mS
jxfh22rz0a5xXwjaFZLbW3f+Di3bN820u1ysmzMk2Ti4ICmXzjgX8/5CfoHeIQEsAtytFT2zLTVX
SOMaKU3pzcbPPJtotPdvhXg0cgeqlbQIqwTcTfxcC+4F6JBLGp/BBZtQCc/pas1+4238NXHtdT2Q
bWfSHvFVcKpOxpQ1AVcuECMEI+6rfrjyQ25XsL4lgVuHxox082OXGa6NwVQY0P9J/HpM4d45U5Ks
lkl/WFavrf+0GmbI5ptANESbwppZrGXDu2nglI8hKHV/OiUF8hwLEzY47FojfGg+SoSkzR6F1zv6
2+lnrRgZe39DxwQ6ocT4LT/RlcH+6l06m0H6GdWwUmnSk2QSwBif4fSUrNGqhgwt/rUJ0jMIZDqN
qyDTJFfCuhOQ1e0m4+GqAkn018tsyGUx//JNbpwmddG1B7ICqNEI66icT3yfCgDExdZ9N7iHcj+o
QZ3JrQJaQ/tjcn4Ua36jXyZ9dlt7hmcotDmLMPMaR9T7ISeD2y+iku1smlWvTNwS+biG+rJTt4ar
oi/pMN0tHbimumpKuWwpcU3Z7airwbX5XFsXWGVAiiyrIQ2FRqWmKTYMQKIaAz5Fj7AGXGpBoeKd
b+n4QPlx7UxqJoFH03amsGqpi2tYTeAWcZtxL9seDg8EuR0p0BrV6hTPAqBiPABi8NAofuImSpmG
QPcxLG000R217Cp3hDQ5PEfOKm0OKku+sZ9zcjuAAHblYYdrYR8znZw5C9kT3Y/lV/JVNsUjywgb
We9tbpdCJgkuF1kavBffcvrhbyTnmFFevH9JBXCVsqonqUcIdjNw4YkbvWr8Ha1KYPKhc/+AGiT5
apwLvMe2LjZ9n65++B84JOAKUxEbJyraJmmbB6wmkDxbG3Zopd8BxYm3kwAMBtxH6VkmuAOrEZKv
4yCuluhHYAKj5smYXwi5Qct7veTgtEDRZyRnE+bnahfFCsryUW6GYoVt/T1x7nr0GNa6L4n2qAqL
+U4C1R4LripdSpG7VGa+D1vfct+x6VJ1M9PV8bOl40GO8I+rX7oMtqbKBoX9KzRuiqlkpRsXtZj3
e9f1Nvs5y4M9SKlCKl83SWx36DZHJBbiW1cjQ9CJtgtl0hci/9eZwXgUyPuIqherxGi/BZ5jF0PL
lvKSvO9+BwyPrAZvwFWSc014NLhqEGRtI+YDgbSS4D6jCSrR9VQepCCn0lqfjl2kZnpoS78a/aDz
t1X/NFs+69rkIndhJIkUMboa+pm3QlofIUFx5+Vhc9tSacyZIl9MIIF3OExLJyP3gBO7K0rXaA/Z
EGEAhoaGuNAlK6lk/XO3ofCvrzLqp+tuQpzIIA0j+sBS73q3CSNXPSxhcyH/VsMRZesD43qE1u3k
oUjA23zMRmbZQ5roD7tHKUJxq+sb8P0m1sBeojWAXaRSucnf7g40jXW3CjSX8PKaPc+C/ZB2W1xx
uPWBDkYLP7TvmSdsQUw3b14tHQ+oR/dChFG+gPK+3cDP1TXxmfGzK5ZzJSponODIc8IR2ib2hvpU
wEHtGF4zQVk4lX1Ffyvt+6mugLIX0KnzjJ94TqER8fDaagQCOgk2RkGrz1j1AFXDsLtVK9Q5w8BB
EcukzIHuXAuk3B/4/yWJGuudLRstbf9NrT6+PTzFQlkyh3ftlvTaWrMnzZiZB7ndDUTmQCPJX9cl
vKrcZ+mXVFRUavlZqP/Wk1brYxuZmWKmYaLcgDGaRddo676n0e3BUeNNX0eYUCgqPw/xNYXMPjYD
xsM9k3V4brukFzLoNwUcqlLZBip/2pGa8cxmjP1zEECST4BgSqjITdINB1pE7Q5H4zIdCz4+7It6
ETDAyWHUwG3e+xj4vaIUoig1JS4hXb2Dt9LcweAXF3XZgw5TVLyMLLg/W8zS5X3GOwEoNlivajlk
+kbC2qG4TCLr0B3BkXoCQyeNi5GIdZuqt1W6PGOWarJFBd6vViuecH6dgmqDs64L/TrD0HsbGrLo
oHEEyhP1r9fEs2j34jC82BvpNdSS0LzGnQojwLMA3VdZJiC+h8/aQEtJEKvG6Tp6JddciRHQXGjK
reX4KDAkLvdtOUuSRcknoTjBUnD/aMvHeBvgAdoeAdR/w8rwVk0kGJhocbXAjaorcEjcXIHzbCze
u0e12jh/+vwcGKrycVDyhy+xMd+XgjRNHQma1TtVGRlScfDQrORUknMx/X4GL2SI6S8MahZpWO5W
GFyUReFBAMhP0XXtoCLhxmu/QFwrFVYudYqDOr3eefy755+nhRPVHUNhlppNn9KrQqEVw1Kgoh6b
MpWi+4es867gvw2K7VrcuMKIh/XNFXnqz6n8k0Ft+jmkZKKumoYKM5hZO2ZO87Qms82fhY8z9db1
fHGjmgEMACVgJpgrjvEksbkPc5tFPawmm+vKWSjj5Yjm4CgM9UOo3mlIb7cEysphA2qqrD9yOkA1
CD8txJJk8oYM/bi3H1dHStBs1wyB1oy/eK7pYDupRIBjB3w9bRFFky/ju0pNa3I6HsybvIPHoj3Z
nMTiDFCNxxcUtp6clLReGjL0K4Hm/JsY9tDRsMbmpTqchsaE6ZGYGLTAicwlqKbM6IQRXigloJPC
ELRCC93FN7492csGfQrJKbh1W51aUGhjCk+AngK+H3xzmWwGxEJS00BO+HGLs3y8xxjxed57Tumx
BBIGf9QUcZ/voVm6BOczkLQT1L2PSHah+xtl5rM14SwOUu+A3XhtpHpURUjOTkN/Ye9bTK/0ui+4
D0KksFDvQxFa33A95RXyTr223KH//RcllaYui5DMJ6OIKT5d1sqKk4vPfDiYX7zkmlL09uStsu51
ge2P89vXNS/ec1L7hqF7Op6nnf5D4wzQOfkdLAZEbtd1r7qsaYUN508qknpYXXlUPv4zpeDMztHr
Na+YGaJAqkXxrqb6Ozm/SvkzJup5RDGibCSxlm3YXYcjY5+Db2pBL4DnbnVCK5jWAiUDyXooPlbc
KSfb6jFY38L/FBStXrvbSe2GrS9GE8H2UAbLmwOaZlfgELX4BBDe2eUk/Lv3hCaFeG7br1je+lM/
cv2GpwTUw6LqqmpDNLVWSoVh043YdXRepNmn3EFX52XSXXQTmUIsQ3CdyJ4YsVyWVI9UFll+k8Ix
LsAgHsbzirTfAC0Vhh0jEgLg8MV1VCEALi+C8c54W1BlpKFnEsEMVSfmbZNcbjFTgxWqylzG+Ya4
AiVFdNXvFTdSxg2CJa8CSaaLwK7uqH3W9F38F8WKeJVAHGEYhz3NtDQa3k+9P3jA5nhyhDQYmQRP
4Fe6mhAxupNvCwfwNqSSwaQm3678HHeTC7L8GW5/1pfA2cd/Wy1Q7TEE0P4aiekLcC6yKt3zoWAP
uMQ42hJmA5uaPMyCjtYj+0VrvI7U7JgB6QE0EkUHNV3uaI/n4LEYJqCT9DRcSCZ0zLfV+uliii9t
o8qepSN5gL2l/ty77d9S6JQhpslQ95aR7W2TE7aJCh2vQjVC0UPGw3Cz9pY9ne1OFJNF12LVcOVC
fk6TSfW+Xxi296NgMlnIy8MhtX3DDHhFTVFm2fI+Q+2HyVS9hdbSn6Bw37DmG9A0QELe18iIWAbg
A89H7gkcKU7NzlRWl33SlTip32GernCkOMk67waLvKqWofKtfLvqMFEDupWjxVrpL9cEcbZd+24G
2iFO36bzecB39CPbkRlHXtyJFaI4oyWgCaHW2cayM+MfspcY4FqxHtfp91LhIiMRFb5oMU+AvXbo
qru/4zSIS6v3lVl68vP0tB5gxcoyGvVoYoZWmwHfX9OPkG6WsZ7+dCGKrnmxA7opj6nlF0WI5o18
+sNlChLB2O9Wn/kYxeDDgQxJ15MFqMQzOOQf1Zz8TdpBpNVkNsvLDic3tFEpLUsQlqT4YO7P0yaN
n0Sp8101SIY4HIYBKGBWrG7fhS7Io/7MJeTfYzucjg8QyOTdsb+AuAYyJBB/luzY0fwOhvoTuCjG
CkFoSWcMHTVFiXphAjQ4FTn+JKGVzYzC4cT7GE+U+xsvORMXaFexqZmOE/rRGHtMRj1HnbmhqtIt
hJ+v/2XMrd2u8qD9bVIfQsvODHUDooo4xDxRu7I2KdYVEbAlSYtcgW/pAJHoczGSuAR5gGALSHsD
pQxLcnuwd1dzQEx3OMkVdWbLXtibtieKhH9RVO2W8dZG0o5/AUnJmUaA9h92+MXhUccG8dcZAQF8
dOL3C00Q+Pjyfo2Q4FC98M9leGbybx5gQYYciaPacJEsTx2tOsHbTgnILzDuHrrauxXrQogoCBqz
eYcDcKY01ybBT1oGIaGzIMtbsnmdEqJHDnEoAQu3oCzdVriW4clvz60N+X0QlsyProlxp8UOVhXb
DOwjrCrff3egya/9nBNp2dn0vO7htmHKqoMbWLr8Uixteb2gnJQRubrU8MmJ6Ckdk1x4y4i6BaOj
khfHzfJa+c5JzcWdqTkr+1TRjateQuEI9NLMO7fn1xEAkTVm5pUHE4mQ/yLNyvgPlEhqJpH+LTDW
mXdz1Hho+cHqfsxpmUnm4mrNj0uWE1w/qQ+/TmnRp9Wb+l5QnteZ4hHKO3QmpwXMfJjUoAqaxPU1
H9ZeMUUT9lCc9qESzf/uiBcH85OSM0hFWU80erqQMvDv1fi4ch5wUl6+RgO0kRf58f38b42gX3g6
EjqIA24p5HWyDv8Rw4W9Ksh3BTWpPSNpkCfJUZt23gtXBTKRZeDHDJb0Dcq7ZGkv58yitIFyFeEt
5hM6A9HGqyrsf9cDRw12sVcUhNGW4zgEMlJkxkcOa+D0mHXeslM3TJyG0/+sRhdYr2zIPZw0st0t
djX+p9venR8wdzWZcZbIImYruw+jc/hZeDEh/GPXBXV0/lfj3+CYXqrzRSWun+6Rpghp/akzxwTS
CX0KgGjs1OY/b15uC5nQIA62dzcuN8YZTK26HWozy9r7KDmjic/DdbyLrnNF8qS0ggC1mgNcKLkH
R6veVwO6ahRg3tyd0HxbYtLSYZm9V02UW9ZPCylAijD2e6rAxJlvBQWEC/Fx2QK1O6hs0HGNz/Sm
22ctqZHkdeBds5BWar2Zkq1vVb/zMOlnN92U4pl2sq8cp2GxEqGtXbg7mU19uHx3mRKzDkbXC4wn
N6DCRrKYwUjZfXUn63DxyA0Bc1LwYBLeYBiwkVkjxRFc2wnzGH4qLNNzmIgP2tEWh9knBf1BNLeh
p8YaFq4UlU4DvIV6QD6+x4JzHUcgFL5V9nhAreWPS5/yl6RJqSCXz+CFCrbeGCKl4JoHsEjC1yzO
eJRZyf8+MmZKK5cGKEDf7PlD+w5ZDgAtnUqs6r2hTR/t8BAI8HxdkyK2hkrKLbZujUg2bFVGi2tN
OVIn/xpDzIPbdrIkyXdXHH0on+FXGMWl/SqLbVjRgi2ZWKyd+HUN9KMdLNL/mYbzpwWJEDqvrAEu
s4HNHgDCr8EDVZ3lU98mo1xrg5SjarsSh79/LFLda6pHhHYsCSbH4Tc57UVZ7F+DnvD+Z9rCKGnG
U6Sf72K8Ji/cdNs+dZMd1xzFzhVlz1vuCwrxggNNs6hYbcQt/1d5OhgV80xvg4dMZv09ZjkNOhuW
em5x5CHRPXGG7mMxRlyayGGjMFzaIEFDW8b5erp2dc4PBr3aMXvRUcK9DlWmWxWULwtA6i+i2/hK
UkTx+TGYvIMZ/hRDKmJjjN4lNm2HRGkPv8durMRkqJGpCAF7CLpT+rO73rPOMn8CSdcA+0nw4O/T
gVM7gPUhZXFmuUp8ABXndNES7A1caSUcDq9QmXreYNnolpeFtmTB6waoGEcOuFAzsLCNFjJ4ovjB
i5Sml5P1twZKiM2xbp1urDZ5vj+gafGdQ6zxYGAF02n54hcXg6/xBxGj+IgSpbv/JVa9Bl4Ee+li
Udz71cUACSMJ8VseesewowKXE0zzQFZJX13SbMf7NVGyrD0KandAz7YxxKP0pkjP3o5TOkq789fw
urTaVWtjrCrYi9RCpiiFZ0fblerMkR+DtnIHkuJZW7fatQGG/t/6Rxdlg/8Dsdz50RMRImdKhD0j
v8Baa+bxKf1AAaZjKUS6kDA2rDI8JW3HHmD4Jtt/nEzLS5jtLUk5P+16xlUerKsRWABOOHbYHEYx
4BD1Ng2twnTRwNEGJ+6MmXH9sChmVparXVA9lPr6ot5JMqDcM5v4N2qmlqX5mUDt5hs9RW31iEQC
J6jwIe68iYCLY+QEpQTUshmYh/vB4BHH8Ht5LiSnKbwe7dfPMReG+SP8Jqp3ZMwblFLQm4qY3VgW
SIB3vao8lDMMjs3BpDNhg1srkR8vYtXsQyKxxZ7VOApZ4KcIbl8hUylJ+FczrmasVQZFJaZB9ncl
k1LHVDc6W8UWCaLPOIH4LVF6ZC6/PVQhtNmXQzWEWSwg3CfMv3aZBcZsIHDZK2BVprdlzoACUwbl
nAPd+OWES2dVkudYEyf6nWiS4qTH1gY2jQId1ktZsRCZ+kNw0YD++6f3kktHtzjZNvdZxooUvMtM
//VQWRDKP8kA/otLQyqExKZ/zr2h23VuOsc5uB5vM5XJa5IS60leyh+tTKiUGTvDmYZsktGTdLxu
DyJksAe/6fBdCcvQSobUngsDasEEdby83JArIuVkievX8EDH3ozlZoky3BO65cyReIDDQXdg1Jgt
CQyMOzuKtdmp7MuvVg3NVJt/FhemlkDUHIg26IfcijmmyjaO3cwGn894aZehoRJ2rifw9EQqJEh/
tNVMMWJanYm87TJIhLZldyMOET/5eC3Hsz+Mwx0cEKXrnIFObDDpt3E4Fn4LT2UzQ+SXKlf8pyyY
xtyuRaKds4bJ9bA1PLq3qakt7xEnmo36GteK7cqPuX2FcZRM4mII8kfZE/qOgYQpNb8cMAZxPNSi
xMJubxlpFBBwg8MQkRyB1MXgyf5fEFpm8zYttxDan3SPZbE+LJjxgQnKWkHWC31nIoNx+QTo0nPc
ZzY0vGUpKt0TJ+N6Zsr+zPuGO6g3a/n+tBIhKoIadbOMotnmyrf/IQZyIlWou1DFLTeFmBT7vNM2
SwH49c8y0diEh772YjOS8qsxNXge+kBGIJ6fD488SNnVyYkQNi6Tl6mZLBifGEjlls0hgI9aKo+J
h6L0Cwk+HinlBhlibl5QixucE9+KKG9U9nhANFtcA9mV5J8b1HpiJMC4RTgsKTxrNrakGADSsbf4
ysPl24jxeUVlylO0eAffNeTZUJ8bZhsPy/Vx8PdsvveW0watgGkw20xXjnrpUH0mqvxC1lpais6n
bptpQ53GoGPtJoSPxo1QNWR+7i97SNEr9oklrcyjQ3gPX4gyLb+T6AaYiFC9rtNbmdLbn0X+Cp/h
iXoSUU2iPzbj0FrvKGCC/snyVU+KlvtlpebKoI0r8769KXc9/p1vtEu33YNtk/gA+j7BmhVHwoHT
hOy3pYfWrcLUBkpUgpVp0KCxydUSe1y5MDTDwLXq5u0ioHme73nsIyRdOlYmpI39Z/0eonCf86pd
Qe0pW9xn9uHd+62HOmPrMSVmjA8cBdSfaa7iIgVWn0LSxjCkChIiwNX8slK+QoKfc94gHwrH88Za
l+xdbAgYHIc4DceT38GOPRieRgMmrXhq4fYEzMh8tBUdfAreQrW8113xYX1fqqAqk2GIEk681EUF
wgI4qKrKVEfRrfyrtSU2hO0DaiZOe0aTaAUDEtmOkNwHLFr6w0Qt+2n0gPcajUZPCQF+ZUitEGfJ
DYgp+lZrQkDbAjHnKJSecZb508KiZoDTJWNK9Lt7gfasKnqcsV1eb6+2mk9110dT6aCmBKCy5HqT
KZlid/vnx5yF/q/eLu1mRMZCnGEBYzLBMsUKcuyk/98Mvex1QpK63IyNk9oMWrMyV9EoYAavtMm1
hwMCzCciH2gE6VJugo2j+v0EytEpnNK+TUIHUw6ly5YJq69L7P/JPwpkspJ5Y68bLJYHn2ZhBaBH
w0nKznlLLHQh46OdDZvTSUYpSir8WnvGzDHLUlqtQ7Nhypw6hDbnMA0SAY8rvuD0MSVcS88xEWJb
ay6eT9ejE1iCuhqphhabsFO/s8KgRC2nzye1e/dqkRgGQq8g0mRdjwh1DDBGUUWsQnqKcDfqmSKu
pWYPxz/ZNYB0Bk37mVQ7Nfyeckh1oJmhdVMPalRaGmRQsJjA9cMFYNVZj1d6sDE4QheVFFt7Q81M
mw3gZKvK9TMpVUTIJWi09mVzdd5U1B85SH/vzlTnKFQbRmwdtDyXL0PcjETkM/pbi9njHq3lfzLG
xWOIu0mHWzRpijCw2/ubjcTa4vsBwdcA7InrggbPajtnhcQJKzwK4XMA1X6/G7FkiEIw+s3DVyqJ
IRPyYy4ertg60IB2tJDAAekAR9sjp/Kb2TWvpWcd4AeK9EJUvvaWppS+tTYvJqjEZKakWcmYltKf
lK6pfkAwmXYE87I1sVINFYZ2MBp7suuliHoh3XovdgeuScJsq8nK/dyuosZSaxbDee4DGLT72NnC
732b689r2JgpZzSKFL7sVEVsbQAR0UpY2YeN0O5fc2lTDKqnxF1IAMjo8lZHZWg5xvNxavdApuqU
viZl1/cxv0WALxRPk51vNHoNkwsSWOB9Qrgu1Gw5V1MbbRp/ngU0Oyl6v1BvTsCZhtSYPIGxMNm3
RQjGrCAR9QmZd1CWdwMuFyBmBFeG4MRTOTl8nAAiMVa86o0UVE0QqnXiBK2+YsYXpi+sd2jGjhXw
6BAlaJG+CQN6BNliCfG8OMOEbQmncKJWnlVgx4UqVhGc9RAMk2IPq0fRDJtHgjV/SGWXDhXK0flN
R6ARcLFEjtAhVsmw+7AsuSDm7+A1cJaOIFBjIqQNjyT4U6ce4atDvqMyXHIUkQmU7SWuuag6pyr+
gNztt7CMrcA7g3VIAzzjh3nvkcDaoumegyG3QLF43UZAfftVK2juIWfylzsoHWIwPgJc91LGBBoc
iNAQejHY+/6U0HGSZQ19FdFoYDjdJROibX9A+Pz+4IPKLa7T1AWQIh3Xi9ZfhmrZTG5d7afzAbcc
p7LEidb0jdRafUPce2WgYCss2z9ZJ3dJDrsAmMLcbj1UKBhXL55pVbJvPc+hF3HRv6qpyWHwUWr4
duAPVU1FtWtPZY7+BuKCQN/YX558/fySSJMf9SOxY6jaA+ZEF4uc033hZfXGJWSgbBCwa+rwdKIi
ksDQPFj8lifxULT+rQUgqWTtKDinL610q7o2Ho5WU6mgcMt35uAthM2Pr4+sG3VKJA1riFjy+onV
Yd7nZbTdQ/4Za7yN47zlwLingqdUztvWEBxkHB2i0qCimXTNwwzikkGThX7QGjONleXvwi3bgpqK
RZOW3XHVt38h2T/YAXWcFlcxgjtvNETcroKPeqTxvTFPmhMtNw3uZC/oy9OF7wqJmbA5Da8b6xSF
fw0OjGHpcO/IKWSLByTOS8nG05GFSwzaGuWbJjmjslxxub2L1EsMA9+QOHTA0cY1WXOyBHzuwkfI
gXi2E+s5pKm+8CM3KsykaayxscZuM6YxCBbq100f0G/D7UZoMZQWIOWkXAq9Uv2kiHoExZWYfR0o
GQutw/fs1MhnXUGMn7mUlfhnx3w+KNK6dP7lfNrcB0Uf0mzYlVot5yl01YKn9qQ0JYqq4HvE3x0u
IQDWRh+e3ppqNinNtmmkJNZ38IlgIM/u1fIuhzMhkf6ljNL2UtAB70zrFxAji0q1K7ETQ7B//h6d
ZI6TkOgBI2MSUPzY0hetlvxlqTc9a4KgyScBJm/1P3n2TTRGR3kWE6ZzVOtm0jXVl3cnhSHWmAfU
4NEVkLP/nekdLVQjXN7ibtLK9E31TRzVWY5zLJsSNN/kvxOxVlnG73UlzzfNH6Lm5YbaSKZ1sJmy
+viK314Z5ON8xMTPjjSqdrx+nCueWhqVlpddyErkLkCsAsAcCQ7yu+BVILfkLBKzdpm7Doo1L31b
2DPZQlxVJBIgksi1JsBrBFNmB2C9DTo0mA2tM9I4J3B27YYUnPOmasJ21APDvc1gIkBmyuBYfjpY
sh9esz5sfXGqtRaYCM7AFr6xlJeQ2hD/elieE5TUHfVmiZ/N1KV1QB4yfaZpmfBM4yl45rj4Y8sb
O3QVEdnXin4SPqrRADv4BX96os+7zLDmNblPJNAH2Xnk+GUcLQAYWzzutJtlYyVvllizelMmV9+b
iLllq8AI8/ITOVQOXXgH6pHtN8dFI/FA5DMcRJczeALWRDAbCIHMC9FyiAQ/cowl7wvVxZazeeAH
zEraxYa/SLds7sSxpl2HOknvXA5MmnbH7X/mCoCYQEWF/TODv7/NEJJqBuMgdIRTIl5KM7QJzDOT
iWWpbtcWsIb1mVM3x1crWhOJLz0ALHnFJskfEt01qgwmAUH5NnZ4oOmQPf3iF2RayBlAwg92rIVr
hGk0uL0pm3zd72VTFGqfSSTphzivJLkwfZNJG+vyFAC0JOAQEU2eBwr9KHl6AwEmQ9qbnXv/5xnz
NKQQSqz4rWb2wFpkvapvOFz/y7D6RzFSXSFbsZvA1tPA6H5AyJpll3xuVngutHblYYvwdQKs5opy
9BOb7QuEeTSOgxzHEWbc4azisEreXA900c84Si1qv4S6yZUtCHFsww+PKxo/B3090TT8JY3fpUDq
VgNIkUuTvBuqKK8lWXgP6myM73ZfN1EOa7kMxf+Sypgp+mdvelbq2l4AftS7/ARQ4Hs+GZOwwpv0
UWGrB8IoOdpFtTFn6oce3RuQzQk/kh+2MrcOCXTHA4KTEjUTUGxC7VYazA5qxEdutbkhuEFltgtz
gZ7Zp3NbaM4Vcz8T7aHhvSQ/OOw2s1Hoe0gI2/Wv75OEaeNsC0GqhyEV4VLPcmGClWgKecOPKBHm
LZMyv7TXiGGjLzSZupC5MUB1KxSc1tCZLACiTd7Eo1BQzMTNEcPNjMsPX9IAno9Q3U2bP2jahblo
NA3feM4iF6oX4ibLkTXIbB+zBK+wx3H+mR++DQpjGaH6cSOtPa+KfK8hUZat/9T1yap6Q1tqf06s
ShajnPEWrMPr6c5OkQVJdLjRiPgd1ZA8DUt09R5flMBN52LbmQfKYXWNdaxZxYSzm8O0bfD8m+Q9
vtLOm/bjYhDQ/tZbHZHNVQ9ujKzeyZ8IjA3yKefzrRAT1Lo9QhOoyDkZ8kbcQ80nFTbPdQQ+uuWb
Iic4VMQZGuhTWM6BV0AQjym1I2aD6lNanVHotQO9g1xNZu0yPj1EkO3tEG36IvhwpuvwEc7GeJtH
1WYOIsW+jx0MWTVHJ66EEqGko5Tn/rQOGSVi47yqvGYnhIvHJZfI62/pjvLbxSqsuvDB67kglXPl
ArHNFrxhGsrOXpBKF/SCo8fzgvFln7zdj8JQbGT3S2PJTr8561Bzu00rqw6MHxd521vqfUXCTknV
RzD+7v5tuwQKgVmj5r4O3ofhR4ynG6Nh/+yH5X7rFvE60T1OtzAWAWjSuMxMFxXAi5jhEPounzjg
lIP1Sov6Siltg2YMhTSfMW//xtzIvM97ig34vXa/1TDGULyjdJ8qB50VgX1V8ZRsowSe/sRDJEyv
HW7qwBuQ2JjYseWB/C2ZXnW64H6T3Ol+qu/l5TCbt9iZHoQv5apvguzX1LgjK4ha57KYUTlkMfca
z8QQNhpIvHFWO/6YEYlRgSV6W0OpcWrc6dq8CNChBW4C2hLZUd6tQcXGo1i22kN/R8kXu/8I0uM1
5DQ75qkaqiHoDvdkZ7okwsIxh+DHgWYIsZOPPeLzLKfqOlsCYY4onzWFSD0Zmx8yjz8Jl4UdOKsT
KBv67KVKhwF7bEMCBvCaKuqFv4Kvx3JGT+H7H9k9MvzHN4xqspRlmTG/6SmrhPtG9qlFbfAwcpUo
H/hyQZa6zdrzr26asrdUOaliN+Rfm5tvbSf3xLc7pd/rWaEv+owq3tRFtAZlhRH57l/qcqcPJr7u
R6dk4Dqp2sJeAPYdRwqv8pqCIo5bPrxJzbIXAofDlJOdaqjLw09SP/ErWjHsOafdSoGZcmAMvIEn
PHLvFfScaJaCl4Ff6f8eedd5LIsH7EhoVY3oQwmnIIzLNQW76Zff94aMEjRZZHj9AP7xieYKfD1V
MR5SxrcnIFt6oSN7tVzYngIMwxaNY4iLYf72PHs/q8RaKXEBWCSd1CFNM2SmHR7ZWJbEv9gYyts6
lJai2qReAKjlCuaGJrXkH6vh1IZ7w22AKu4x+VTrFN5cYBOEqFPqloatQroiKgHj8GdnMK/YglqB
Dq4YAEfTP7aVBe3UO0X1HEbqGNSNP0AIV8fGYZCyLwMDfMnZIMt66s9CjoSxmiDN8HGT7YdIbnCB
27fH0NXwT1bd6pYZWHWBAeAJ9cjHXBZEH/se0lvHDt/PuUign5rSjv4H89MnQoLrKrrW7Jr7brpt
+sy5TRMgXjdDaGZm8UuuprLNufmRpIB0qTXRU/v54f742Kn4iWdimvIYL5ZN/28dJbHiAoWoadOn
4uHWwfdKelgSniTTki9JwC+fdrYLT5a1zVJmvyFpwHUDpHSQL3PooMPlAm2GsJHJZUiylfEARqfC
Cnqxyka+A66OQ/4qj2EKo3vficTHtI8rcj9pYafQ2Y85Xubp2ANZRljhc8guwsfW6fBy8EQmR8qG
uA/JacHwkRvT7iV/AmvqiFSbio+E6O0qkRPOfyCpzxvhC8JLLgum3CXCGLFL6mcVqbKu0CpFC9n7
bKafSLoZ1L0EBvqOgcFxfWv1QSPi4s9kc4X/nB2Jt4lC0VLt66VOShVe21lVdoihBOwaRz8KNZUQ
+M/MIjqs8CdNn8bMF2ACNPyCjO/s4j90rtwP7qnSxYWPSskmNV2ZB+U+h2LQeT7a2/cbFtKRshHi
6jhchcnTxjqGVBZgSK35qrBY8cuWFLjmWXnq4M+E+Sj09bwk1wEZhu4IGqcnpeG3t1964KRrLgfZ
BVv8XGNqqjKeEdUi5s414XJDT93t59SgQY5EgkkpykwyAUJjJzmCITUMyfsVeuSfxayAg1VyUTRJ
1CmcnZD84eIIRqLiQnNQ98ezgVz5D5iGTEOxFrrewvVliTXFsgPBRdbvrqYnM6zK+nI6J2N7xIX1
L+Uiy1yiOsMPEQ/IryuJSrpP87pGOKMU5Rldm743C/IhRvQkylsuwdQs2Udy88qbKDfrhoLOmSJD
44vLOGpfyTG2f6hJ3MaqgOYzS26/hEeByDzP4XY1GKeTOF+pYhq5nX5eqg5tT1mnkPv8iwOQDSTR
4J8zS+Ye77ED0ceyRPF1166FnCKNCfuQMCryrUrRhY6vYIndWM2JnhuPmKMdtH7+8B8B/sbIB7Ry
iAU3krwAS1/lBgT6zr0xWr1vRiOWIoUDrzHzvQMa/XsOTgwcn/Ip8G9u+Y0rWjKrljFRmEwjQ8NK
evcgqGP8WkW6khUfkD9Ol0tx9HuQlNaGnSSGPXVPun8AmVWK395fKl2LB4H/JoKFIwLgPoIadJuj
0em3+H2LcqJqlz7OlDzXkrSPWZnx885RQUk0CjRCxcKZvSO/Yp5jdoUppRJp3LelB4lowcbwthzq
0Vaeup0U48psm4WwzlGxOyhP/UpaMgTc9lJqvyCrvdNSyJgS5qFuCoc57TXwt7wlwijUEE9be7zk
I374PZEavvx/g3JyqqBtQx3UFGGocswBsVcZ6klC2UKaJPnC0wyLgc+UqJ35Thv7OPXVWcDvqDd8
cAxaPw2NB1grxSzu36FA+Xv7AYl/0Py5tVPPM0E58EskKUwSz93vzWdatm6c6h7O/VYXKS+iy4G5
FQ0ZPe53PlssmsyQuqtZtMjpPwO117jC/fALjPL9ELbqzjItcm8veNdq9p0aJtmNgVfjvb/VwnpB
Yvb2OEalrK0hPQxJEPoxQD77YVzW62ToXXoAfc//9Y24kccBC2odztS1qaK0oWUrmw4VLIBw27b8
9Xzl7hlvJhInj0628+tsSs5kIUDcVFkhBmL1jKr6Be8imnDd6VVpQa5oqrDnVSqaUPYJwAZJldnO
TXzXXB4XtgHp/TMdsgH5rma3EpWctQpo4Ugpb4nNQVhCK4p/uE5oLIdj2jVQAtJGdzegGXrrGfqF
WIN05DvR+ZmEaEDso/8z1K3wg2DymroDzepKn0f4EIhVrCjKHLMo8tYkzCLCONMHTFmprjxxHMo6
FOSOawcSODL7uCSuqRjF/x828XWwMCC2lMoqkxqeMq2IuWHHrYmI/YQtDFrzuG/VvDxboflvF9/T
9wAz3hKdPsGp0dKuuIsMYD6TW+Rxxh2iyEgkQYo9y2zislWM8dPatazTAXtjOSVspOQvCPVhO84K
OL7gIkIPWI2cNcx/HS6uPNdkPTSYYjft93LMADwfXjy6kAsChRInaEAMX+OSioYhHuBBk/9S76Wv
XVz9mbkHCgppf1GfFgmZob6IQtvf21T2/hgb581BY/lWyR0IiIKujJl4eaVkFYnvH4vyEcKZnPNA
gRoENQCaR/HYIVZbMq0YtlgHCNrAzI3IV5eFSANnRDE3os/UJhjDg65Mwd7/uQAP8vSVrwi8e4lm
GI4doZap5NnnSFakcrss0EHizHygfCPFR8jVDLQ+WUl89iGpdZbA+tA2tDsSW/1mlkS8R50nTK00
lHXZOkeezW8v9mwRXBALPhS3Fwd0oxAe3W4OADQ/itN2vjcR9dXVYkHGuDaIMHlCY08TJTkMk/XW
SW5RG83MC9jDff8xBSLZY2HHIjNW3an6Ic3sn2P7pIC7/aB1yaZiaYi4HrM29A22JuchAKaEMx6N
aACeQDRmy8mvm+rc1ivV8vx8uZro36NM92k6WpKrr4AxbAIULeZSQz1PRsGnjZOwFBOllDiFFxN4
y9yHMFsnzf/GvVeBc0q6uqcxIwkLDI2qdoBs6h57hopEC+FclDPE13nlyX+Twjrqe2+kVJDo4AmF
xt/pyABEhAq96RT4GhPwPYxZPN4KL0nUPT+yUB2oFXlmyqKCTVAKTb1/s6k/FoRm//khYDfVQiQj
dAMFqCohS2TvhsPV67uHFPTvITRJFhcXxZwxED4ywALaBFXpVmIDSSZVVgJkNsQLpSZhUXQC9IDR
zJ3+TCERRYM/H/bI74z6KAlEFMVGIZgv/DWYszrVYSqQbSbsiRHWTH8uh3gsTZT/Wtp6xXXrrxZK
BxsdqVrga2/meshlv/GSFr406PDoylTSK+d++Jg7F/7WEiXZCGoBtt+PSmujjavyDqflu4ZVbf4q
2n1wdVZ0nCcy/YTtesmGXIrvC2JGNbJjXd55sr9F7LqIfewkNpxc+QTd13O8D7pb5Rkc4UnxZJ7s
hdJRcBP5jBk9EN8CMUKQ5a1+NsqLASff6lG2/xtccOy8mlbdIbCN1vIAPZ5u74Lco+fDborx+/e/
U3/rhyfsXF7nKFCmnwyO2wEbTOu6WinLNo+W7SlEOSqXdSI8KbWR2Wl57P229FqCOv9Drkx2Ir2/
/o5nHUitpIDltCYH4wj0n1b0bCPJboco+iuIfWt2UEgntdMvghp+6rEYkeswb525ghYdlnIX3lW7
vaFW1jZMIl45tQI3muYeCi1b5VriURoT1ofD3XIlzg+on0iuLaMxlgufLuPV7xyWIIi9zfBs2e6G
srguF/BP71Phk74pyZ8LoApeAIcvlXmJdeoLK16NiErVaq7lihs5p9JOjuxnnmW2CGYrhyYteTi+
nrLpZ6Hkag2y196YGHhJn2uKYaVeCN5Vjz2TLYvaAXMHWjNhFDA/s7GS1CG9Tv3T5cwFKlHCRu6w
6frprvwXmWMFPG/CTYxYdivOez8Ku8sgiFJz1fMhDQW3lvrKuD25v0S3Ei4jdk1NGWhKGOMedcRY
luSIkoSFkhWQxHFh4usRtjZWYKllsNG3qIPNjvPhf9h5aULyUOFQrWeGEi1C2YLOHTT9edH4UUNJ
hOjBYKZzamVJvRmd/FvC7bxDPGTUGrqW3fMzzjquPjk5T8lPIDDTRB/O0Khbs18M/MkIKzqtSkbJ
24tx5QQR/qB+T+ieMzTIs9GHj7vp3BlR7/9m3AZPFUdB0Fi1KMXDsgUcUbGGU4/rn8kYMQJBF0p2
WfbhdLzIrA/9lYEBeYYCmZrDn9yXTebAb0W9Sjx8lOUp9/UPytVOcNpVW2kP3nQ2UItxw1OnSSsW
edbPhykuLarIkGXviNFTSV1agANmNvzlTNhHVWyENF5dAVjIqcDtglXS+jSqN3Nixj9ID5mQ+rb5
KJ4B1CKD+Azmr7z2PpAvRydNGDOrrlJx47pZ7RzvMEV7MuVbM2mrDo2Xuz29a4Mr6Ce6tMuF03oo
FgO7KhbF+FJMm3iVqM051okUZrVVIGVlWkDq7wOuomyWUzLy2yyjCgWpU8z7Lhp/W+LOwjfSi1bQ
+lcFYU03YkcBlLjXdTRkByfeRaoMTO9R9atN0vHpmuSI94xHciGLgzqHszZqXGmvB+VixtghYXpp
9Q/wVuNsqVKy5/FxBB280KAQ29KabpguOAqywIomoadCW7sHk7lA+bXSrPL7usNW2R5M8HXvDOCG
mNFBlfxa0cqEz8HzhY7d2/mGHpib7MZEm/XsJxtySoxZBU/eurGvjJJ2ViXlfnMSMGE6dRIELpTj
tdq/bUARmErcWGZMhmx1JTBLjIfVLCa4+aY258xs84h1FQeKgy2r3rDD45vjm1aaDyyThI1tiLxf
OCPDcp7q686VSjz3aco+tRB07ze5syNXkFwjeDP8iCHsb4Ib023R0GdFCa42kj2e2lTmG+bhICc8
hwoZCN27yV6yUkil3yYgg/oPbsIR+ttbAt0N1MiSd6DjdWGNvpgSQKAkrQaGjHxzHn5gqqv9zUlw
2iH5I0xWjFYSPjQA9v5kY4pPRmk0WtvvfdSxzX7CQZVXV2DtrUTKiDed89o4abRKwVeaEymAQi5K
hjiGajG2U0jdFzK3hJ5pXR9XwiB8B84+ZlklvJP6mfevpaUrVQwtkSpcIH9cX2f33hXpvJmT3g2M
OyXya7AjwWj88iEGgdU73Oa30cjuVJrshjnS1oJW5SjxkhYB1rRY4EndjWb+PkxH8xVIIm/j+DJc
3fvC+FcmMY2DeoRoykFLW9E+UiqZNnxAJvhbiNYxW6Tqu6zFdNsbDJxwMTpmFCkQnOaLVQFCnZqy
N677da4OZ1xSB4DZ0CGqjzw5XR1GLm2r41qRP6Uz8Wa9kShTlRH1Xy3DMcdAvyr5i22ha2fYCkFW
u/14PO4wCAO07PFaSD3PcpWrfYVELAvPkdBQAGFRJ4mYdfSmctO5Wdxpm5E21NHIlS6VeGKbEIVz
y1H6Jk5NnxoL+L+B17uet/k/9KPqAolbg2RQLUI+kaUDnMYaHk27bhzAFtfaKTj9THXx7yY9hqDb
vVXVfnB30zkjDNMcQF50T8V2wyBZDESBN+jZjp1L2pm9N7G4Xtdspx6yZrFW8se8YBMWrkCBAxbq
z8uvP60IjAGC6s7/OqNnr+EDX9X0SVyIQxuut7vP0zDA890UzUyd1cQfXNhbY0iHs42g2jeomfUI
Jv3126w7y5jCRU7uW4OUSyW4csLc/iCX/5xEb0/WSsl8vOMTkAOe+B12XryZ7wpTAKbm6q+M1cde
8Tvj3XGdSdZIK42dkUeFm3VoxtX4X81bR2neTFFqspQ2sc1dCPV/mCvWHnaeM9rJkepyCmCxYFoD
bhbcTO4YGKn8JoinTF+PO670jqU4cg0OtJ2oI9WmPrvvRcFsGf554dmvGggUbPvwfdz/LiQCVEaj
OW8dYuLCz4lNdx3d3QJ3x1x7zPp0iORw6Pm1Ddi5xZFNq5RSpPmd2XnTZGj8WfKUUD2Ot65RMW7+
p95zrJaP5uXC3gMU33VCzy8Kc266f57A9PajVgOhqYWeWlQJqhYa5JPAaajgmqcaDM52nTrxbyML
2QZvbrgGR8mBYQhhSkARzyLdje5FAGlnSV7naDef0/EUqBsxHJqhIqohAXSYgg+mm6cMUkgTGi8/
1G6iYeKqX8XQh6pKCcVyzyV2LryhSUobkM7jgM/obleqUkQl198Bcm6f1ET0C7Z1PzqUuk42pvML
zfct6q21vvcGXIS/fQE8dV+apGdqxE3BJ8wBPOtnmVtgVXCIz+ggfW9XTePCH0lmBb310PDVmtl1
zJzScWk16awRAqJ70T0G0GOivgM1KgsV7MVhrtDETz2I4zV35wPPCjh7EAkEKvysI0pgl99FfG8L
Gljmj3Z5Idp4v+RlBbvfBhToO4fbCxg9f4Xzg8vCEi6WzujB2wOdQb/XC86vaIBVRc6zzota6hCb
JyoRHmnKqDEHVYnX/wYv1ePRGQXmvKUbyk9LDjjJ0Z4wD2zqDHMY1C8RuLhCZ/fpAeWOqRFNOmX6
alCS03IDpXqGIqftcEIixZfky3OUSQVQSTbjIrGyD5aVYRVMNXs59Vu0otTrphwE4x+zsMJ54GZy
ksYEabOeJ6vM0oGCj/nVLD2xos9FLwQkQPfk22lOc7FKTj0+C0Zj4okEJ07lh9w6z4UznS2bQHzY
FXn1gMpoNV46KshUrEMkN8CCqZkS9Sjk060Uw7WTOJb/806D+JPLkQtNaTZ+70pgGeUWJ912JVX8
LJURFuXaxHPoFR/SDidZOmKotKVnofOogOfEDGuIBaQKV8K7IWjSh4Fcn+2tYoApg7KhEwHuwuU6
6a5cJayClV1ET3d+uuvtadLWkDC9oVRVlvRRVB4RIROPKsWJ4y8WujQwo7tdQobXK0tyW2fAnA3H
DVrpLnBe/zLXnXP6A2lpuD9Hv+7QDCCcggeJivFaU7SKgKvacGtap1RvmzSlOKtUEZfnw7ZM0X/2
jJIdc1e4GwmC87tSHhBi5z9ltMO3jPcrvCHjquax3y0dtJz3b00YW7PCuPL4ejkpg+3FF9fWz1Od
etmA9QkM2xUXoD3y4wDKR7NpT6QBgXk4gIq98UspxGZLGF1WlWmbII5q0PAKiKXJ9od5jaJVKkhI
jEH0noJRcO6RflFN3Vos0gUhFoEKvE47u1WQcZeUdSLap1RX8t832BuPQk8oiH5ipownLfRN7W4J
P7KlHIUtrtpQ84rSxz8Fui9QndacMeib2kUL19MX4KkHD3E1qz961pwCP6x3A5p6/LoH60foqSit
feRBStavALtmoqxAtS/3QZYyWIixl6/1Hzerzg0KiSOEqRX8SY5D3bRFueWHWX7cWHUkvSrxW9LG
xUMxevB1eW/pNJOXN7YHM0VhPlfX3lP8cQARIZpJdEAgKIEixh/jupE/6wgerKxvWOQXdVeQBTpZ
cugKlY6hNDbNEcTNhf5oP7ZW451kgOiMt5/tfTWNKraIi14DAn970+97goQTJHU46kupIwgB7/uq
DDAltEmyT65nyXPHLXUUG7MKzxeY6sx96L8kd6u1h6QsFeMIH40EhvOHz8IOBtLQb4/V2behOdCZ
3TZomXbraYLqyedmOi8W1HR+s69G1MUOcWR1ZNvwA65hOKynneJypin7NdLlzhwB5rQ7WdzS3re1
OZm9wIU+6UGVSA2yY1wZ/69kihh//qmhrHGckTw9qBKoMCMfO87c7bNFMAwoBZ7j0p9NCv7Ye2fe
pqa2kiYZii6rJqATkf1g8Vdy3pWXpqDXNvR48lGfFfDJJHN7aifJ5xHrn6WeggvLE09R4Z4F8w/i
HqB24kvcSnKDYvfX4VvzjDsH/Yo80YoQIVPGbe5vKQ+vYj/7lu8MzUMJqkUl/zsprWrVcw7Ew4Z+
y/2PPulL099zjOXjSPXmELXQ+LvRAX7nSCJFK7/NkLM9Ddcp40lnyR68UP/idfNjL8ognGPGb3cs
XABH9CQns6fCR4s6KuB5AvaxOTBoM0m32x+jMRVgaQyr3jgPQWUy7HRZ1nCZhE6tSCq3KZb82N/A
5ZQ50k2F0FTxJkxc2U81OhXj5+swqcRYDtQZejLsYe4g/GEkWyRIcrtSIvjPKiOgblwfFWrS2yHz
nRKUJ6M5SBHXR2AKaGjL6jPPZDRzZBNSkfoCXIYbff8ZjM4HBsC6HjFma2QmXowCx6kcF9j93Bu4
KSUwVQ1dXaxPKapyKAm86KsPeOfZ/7o3a628mOvC0OTeBcTNtNGB43J4F9VaUJXJ8b9ZwLJ6kORr
UiOPdg4pi1Kkga2ICrmySG9bo4OtER+URIFsC67YReeTjCEwjy+4SLh+7HX4NVVLTO1mRZtD/J9Q
m0/fAa+Tpao2tUvukgYPTgJrVrHaIE4fVgMwoOifGyLIJgonIRG7HmHm+siKmRB8c/874WGu1TDq
izzVtAn3lvEKxb+CZBfvYsCwtDU5oJnA7hXnTdhFEMHuflrjVXZifREtMf9Rg29LskD/0oC1lINA
RD8qVDKD0qKF0bMBNPCB2x+ehO2U6Jv3BRd7iMNAvmBZAuD0jCbpFxC53mYbI1UCWz8wSYnft6Ka
ohxEfehLMuXfazF8cjIMtB8/Sl6Vl3CQqytXA0X4rc+2gvQXx32DD4NdvokvIOj+ZYhVOkgq8CvL
AiAHn9r21rIOBgSY3IQGA/Dd3Q19JCtbRH414Ntf8PFFXZlDwQX5rklVWwO+d3yhGd9m4BuCgiDq
v9WbT3k5nuqk/h+fKlKfPKjuHGLf2rbxNmHTPdr+nof4EW9mDI6qaDEEVtiIAU72OgFRPH6aYwTO
NRxK4bUtJF/IRb9CMQb4gKAtLodgZBp8shqhh0eNqjypdk9XTXbouf5cndH3YMuJWMcbQzhwOTs1
x82zjFROB5XSSIpUn8YUBP/8jqLVs0sy6lqOeL7CNRxCR023CxhvjCFNuJX5KwEYJ7tTA9ihpXGl
jU7IdZjiA6PVJ0v7ASBWDR08eWoOBJ+eRZlZ0dIow1ZUdDV9l6mMqS52mxZgqbhcK5TX9mbbwW0H
Gz7eva2Xk6IXFA8oZfbFc+LlMBG0q0qi3Spyo04goJuGkOnzzTWxzo5lb289V9mhupyS3X3lv0FV
XBWMkwXsjjQZjyggMKB0TDh5K48/Dvp9d7HOtgWjKEJyuSEk3O+Le8JWZ4l7EBtZ/LH8WHOrIvGy
0eaV2KCFklN25qTKhhVRT/xpTDNujxWgctTy1UPmBi83tXINwgOy3PLz7NXWx0mf1T6R0v9+73GM
CW0eu6dHz7LtF8D8/At18Y1KANPBHXpdjWShZscKUCgnPTZJdSbdGyAP9K9PS75Zb7OTzH8JUryr
y6fM8qbrcvH+Pbe52L9u4yuDGF/xWJs6ayUG4HFZ9UCQDhAA1cm/Ps0nETG1WdGzjbZAX8QnWFKW
mlMJpl5mFwd6XKovpClD+IDGZpDKuHN+MZlTeyVgCEM/GYm/07eNkUSzopq77CxoI4VgLQDQXP7v
ALaj8F/C/H9lad9oCNyiXgS5k2pQAGoxbHlK++TWROIZ7pqWE4K3kAe2X6OgyR3sZqTolfESa+Dh
YVGTiQHb8bvMTTtILlmjhjdttfCqzwKg1rqvcsxnyKp8HvTXYpDm5U8XPatHqdeW2GVMCX52a8k4
RY7v2PuSKkA9yVO5GFY26Dk+KrVbPTkGblfub6Lhs/hhdTj0JUNNiWdjkn/FIuoYu2KBpT7eawaS
YoZwJdAY0zTH9Z/hiC+KZFZsBJg9ZV/Owevc2yAKz7yhijQzXjBDIaEQiF1AjpDAXl9uDxCyOqbc
KymSajDTA/9cFeynndY/kWf1YOjrGkQZ/bStIBaGvGrtG+T46FC6v//jQ3GZ3ip1QBi3f2TpdZ+m
bjhxtYa2HGC9nKnmx3SbnE421icRcc8xugZuoqtgjf0kuK6AY1lpwKcEls1MB1hurgV8umkCDkAx
pot+xZA56iInF+WVecg4v/PrH5LENYqf+oFtFKWb1XsKdCLdVOfxkJfnr2BzKv9qEOTAB68prsBX
DolVYN3YAHd5GJxfyqcD4jGQoEaJirJkZ9XMWF+qCHTSL2lNcNXa6nO3NtFIhNIgfZk34bUxy5An
Z4AyiW+C7b/0M9y/XS4NQUErgmAUV1SzxoeM8VpRgv9dFdm3nxucbSA5h055k+NKH2mCg++OUx0C
9/sI7XtirC2xQOkEDDbOdquQJPB5/QiInx0iCVSy0wWKfWOy6mkuE/RmJkMHND1zMf3aP9QLOsrR
0CActX31FEjmtm5t+D8JhoQw1qP/FYJHtD/qrZCKTUgZoZNMvc++OxuFv3rxNxAoxSZjVn4GaJyC
q9V0Uek0uNWWln6oOr+APB1YxMFqY6lmxdJHAEyd8/ALkGOYXlv0j3XddnG/T4aoTXPIRE0O9SYI
y7pfpX/Pwfp8ToShE+xHCfqA8aeMAjbgMBXg6qWeoEGEkmd/xEMFv+MJXliVcSARMmzvj1s7CAOf
xqXu5p5yUjY3rQWknj10BjDylQoULKFcWI04az9pgaeVydBwSFC1jhv/ivbbNrwjfqSwdSFJRFqk
O3rMaT8nuJnEQwjY1dYvj5gjI3bicvh96AfLiPXebnB+qSshsbN/d2gIYlbMBzTxSGCq0Z+6kNC7
a2rt2HZrxL+vqhLw9Gw08VXJdeAiQSkF5/w/CeSSHbi+nRb+Fx5wtr4TPky64Bx4NlSw+fPZVh84
zPtoRSJ/s/Mm+hwhN9Tt+yMs7mg1oUC75qG8X5v0KKW36Coup7JWcuZfU3Fg8LQoj6TCHcwieY/j
wpSmLqUNt69aNdKeVrN7RRuVEREsvP8nyOmkSCqcY3aSZzhZgLsrN7mXKIZk8/UqQrwexaPgwsui
1U2U6ippdV7RQtC+dVs2uMoV/Ckw/KuJ9QiwyFW0xgQFyyG7IJZD59BhWGIWGhlXVA2sH4ZPDAI9
ok/vYQctTPzOqpqVhTKW6AEVhEs3wsAibdv09kOCboBuTXYAaej3sd4IeeRbv4pHTnvwiVLrJOeC
pFJ5NUfRsFIY4ljR/Yjo/JfeNIZw9t363rwMGwNFG50QcN3sWxR11NB3eca6n+lIUAH9Ia2iWLLy
+oCoy7jLZmArSp3Tt70azds6SLaQertBuHEeoc708Au7cAet4RJ4AAMm2PfNBKpqX52xeBXmGzkD
o1IFNVYJGqzaBWZJXUV5THdsk+fjfzeNLlt7nFQQoqkHcETwiERLDi2OqRUGwsU5dHxVuORCDgTP
evvjq6W19W699VsUCSDy6Pjkx7Lms58FRquVRzd6lFBIRYcLqUOgiMtCqv0+/aemgF1KEBOF6cJP
UQABSLVmpa1ujsNWE6i9mo7ta/1gMlKnGeMbmm8lOO3AOtTKzwRR94PlWqtUZUNFbJOk538P2K6W
a24/I0DDY2p4cHqths7hiYDSmV+VnEUMtenwxuhQqOhM0rl0p22dN/YpMK4HI+xvCOZzYbrBZDio
Ningf9WQKoILdGBIfi90RbQqcDhKmkTiK2DkAVmp8RlEV7Aw3R2vpaFQtBtVdn5Go8xHpQNPedON
iRx1D9PdsiIOT4RH3HiElJsYAnPoOL5r+L/WY0Ok1Mlc2pcDXp7lz5cKT2DW5ExoAh0/VU4K5K5o
He1bnzpIMVYbsd3ktqFNZ/FdMa7dQ/6J8DnRsOLAbOVDbjm9+pE5ERcY7fz7kTT3Iy7DMiitPMZm
VJjoM3BVhZaGws7zoaKGJlMMcVJ9pK0pq35jemNsZlnVtEvDIsxocMA2Qhbk9qNxvq0oGXfjVaAw
Q4kHXCau+qiM5j61ymToyZ9JqIOWbqgBmQ3Igi+yjz6/LxnMVb9fiR+8wlBUHAPtIQnmrQkEBAHp
mVq/54pzNg/V2+cvQsGtql9UBQt7jqhOS1mOpn8dtI+AwKfsO4ryyBxnvnC4g3p7XlCbp/ALegeS
qqikaiGnYgUCURmbm/Q9Ezzdf9kCmEqoWqCRkP0fu6UCwDIb/RcB0fKKY/f7F2M3Ka7DIM4b2Cr+
v5n8Y3EDwSiBYLGxLDP66LFE5CJdIapwYzWLYKKKS6SZP/VhRkFLGGcLKE1rj/TaeZmp7TOT17Dc
WcyNicHiedElfi3qpvn3B/FyrG+m3HqGKg6D/BKJFIzH47RWMzd/37jV8wRxbIOybqEwVIUKUKQl
tTQPd9eOxVM/jYH0VOJGkK2w1vfroj1gzRTgtrPYsA3QYYz/3GVtg9v1Ve3LSRyBTEQ2x0Hx5dlb
EcBEoakn6bDryboA4iy9nEHj3Wrr9lEa44Mc4mmi6UqzVKawK6ceDROORbAASqAPeDsNAN30Ozok
wQDaPoXLBt4q7UOwEVCIFPvvaLBZZkgkk9Bbj5k0t1bhFvDZA2oJeABfu7TpPfOzl+U8DQLC82R2
P5X7TLw/9GcUHIveev63GfBzT9BzHLEYcrlSTlVImDzB/OrYUj/h1OASPlb3VCf3FUga1BGdi9QW
ykyMNVW5+I/dVcPMUmMo+ET5cCn8DoivAkGlSTb7etSsuXOxXgoALs/+TZ9gEE2CGNKa2yIHms7r
ccHXUfK3FQbm2rVS3u+tj3PZTNbMbioqtgereSKSlhQyfO0LxhOCQaVvke9GH2eTkOYHwTrHKXmW
QKI000ZZrlaXKe9rni/dH/EG4/9V6H6pgLQWU56rk7kGX3yBECo3gOHaQq++SSETKJszcAxVRvYJ
DGpjWhbhY69yZWC32zTN78/Z+8jQvejgJCczXido1JkHCPrN32vofebDs9BxyeTu93Dag3s18s81
WVvjWTzFTakg2NLYo2I64YlVIjCQYJM/81eXQ5wXv3LTY2yNTdVplOWEcwkn69CBTBKE0ITzi/sI
50jlWwG0QrC8k2RugsKUjd5GZY5//YKCqFtgmJZU8Pix0/sfwOHEcLm/kyLVvt+d0/izjjJjq03C
ryER6hmTAZbxLZ0J6RRTh+zIlLSVBGSUVvod362kiO/epIqhwaVRHq6HIMHkdzM8B+7nTq7DJOHF
g5/23aBaPoWvgUI4twNkJXho6OnGpRHh/pag2iL/WTLs3LkGbZcLKm3p9Qp8++tmQhP6FzaAQJpc
nxVlIxP9zoNFgTh4ESTDxzypAkGXd7H0IUMuv2JuW0sRjclFbnM/ThSSOnprR0uPnGPoSqwa/Wyb
laIUXjZLqpo5sLi6dDS9UuUJMHLQxPo7Ude2KbWvb936r3LjBRkH7yiI6eueIHnpmjcZAikUB8+t
Nl8pKs5ApkaDpY3vNkx0QCSwWILxvPC/QPLgrJ0kWD680nfydY729EyMOT1rXwmxNdkfdeGlzVo+
0oNcTBuOEoj2i3JvjQECZkU5X3lbCI2n+A5Cg3BXRaCF6Lo+mw+CZVB8opG3iI12KslM9NjFGwJS
5T8Ogt2eFwhcidj2GlJHiAmytaCAKy4TiGa8G0BgGTbQZnqQdZ5zty5zskUPHWlNX8rSygYZhhcQ
//IT49qN12MdAStkLGGVr0bE33T5bDmYR2MwC4eU3p/i6RVTyfLg4D6fLaqewcg6RGZCSM0DPtHP
GZ/qyBX380dmySrbtxOtmlK5Jyi0KFLO4NNKOTwkuExLf5xEu7I2c2tg/cRwkUnnagDsFDnGov9G
4TzNncWcZBbVZPH1L2JvmIMnGczJcnXu5cRDFonud7fXjobedqA6uEq1avaamDIsmNsq5JidbF+x
9kOT72FBTDfXUaYdrXOf0010KxuiiTUgDzYYeymz8RZuWLF2m4t8EwGiHUFkoxDngsKwWkNwYz6C
KUT8MjIk18n7cDkPZeZPuA5gQ/JSolsVZyxGfzmr7PI1M18PFdfjIIctIVXs7umjIl30RxfZcR+W
mznjUvmUnENqz7kCxTLDNYYd5Gnh1iq5bdh6E/kdd+JQVsD0lbZ9P1fBohEZ5k5CLVoQeQMscQ1r
q5HL5eHMlfYyQxzW+Ak6WO5iv9xqsb/VID/iCwRXiDzls/ezFBbS/oY3UPptjLEUbyx6njggStfb
TjNY2MFcxJKhxH6ITDCiV4eUTMw3MZ78EjnbRON0onqqq75yf8ukWfhINwCaG8H2ZEoNB1Ubt5+i
ySWqnnLkJ6gFxQr08Bd9PEaytjizyFCd/nPvO/uT334Fjf1VBUKsRdqaOKAbebNZGBUYNRwjEbSM
ChFgFhMJzxC6orQcMiGyh2Hlnz/V1IMtuRySNwLku5OrCPmEhhicS2HvTMAN3TC6wbftSAsTrVPM
0TYpioIgT5StrCMB2Y6i+3LBMQ5NBAiKLZ7h2pW3Lm57nd9XF0V7kjv+oP9n7s7YWO8Ax2F3U6Rt
vHYSwQmk/xCJLQOA7lOtxMlWd0+MvFyKm8YaPc0VO1d5VhPuT+FkeWX0rIEKbUJVV6bDpzoZ0o+P
g/a4IOazeQfE83UI4HdHkMJG8uViNzDlQWm1HEuZwUQhZrCV4EO66MaK9ppy4o7I1PXkyETrKC+4
Fi/svB2y/VpZaXJADM1bC+Vqf/liytWnuao5wAFKgL3G1issxgHDY5pkxgDB6mqy/hj9nGM7OtUh
/VblI48UX98BFVgylOCQLtMRoYpGp0AlEGSYt10z0faCgciVnmWftCDnmz9Un70iJxLwxbFuCxU0
Csh3/sD1DRTZrH2pq7u7IK4ydebBkLpVSuMJVCXM3b1yzq1n2jawuje4RvTb8GO9PZMk51zpLCoM
OqTsrDj92aZU2ix6Znsh2SyLbmfc7l4kpUrJdNODCF1zFajJS7gqAZ8VqQ6KzuRb2Zws5umbmfVK
9/7ur532SNWyyxqZNiRXryYaVaSd71+47D+zmMHNb1DWf4p4zlsfh2PCpIpbSZ9GLlNmvDVUHh0o
3/vWKc7cQef+sii3FyXUZbdq4EUGqAA9BcAIkZBVRA/XrdYRQl2M/Xo25IibdPOaustWh5CWau8/
Rwq4QtpW+IX99UftrUWJ4Ntv65/XjjUTEDwk04Mie/Q9/sOoX94EYx1GwJzyQnrsAFHlgdkqxxRk
wmB+N+TM159SH0dVS48BlthzjWVpGLoobgdcPGjcBmtWpOPc24Uy4vAhqfaQZiwlhSD2Ns89mgFn
xU2wdqTvplmCzUdlG1UMYlE04E/2pYMJmuyk7UC2Rbddqa7xc/cVJWyOXi8FtrLOCu0Mz1U1ifb6
wChv9YFStehlVXGeKgCsmSLOHIQTjj+i55c8UPW2nN54inA1XUQO0dNLaUMvP3dlCHJo3Z/ykzoh
+gpKDdfM4qImHeXBQUj4nT6Gy67uXvvdsoMnM/aogpV4fZuf5/MU736NrxsxRbPG0u3WPNndZpfY
aQv5WbnB/F93Fz9WWyNh4px+UIKXki5b5VnY0ve7sxdJSGHi7fXSz4K1DP167B/IhbEfcDICTIQF
5md8UuJ7Yp//0xZTqjdlONj8/3VnxrDz+0LDDdDm+5Gpl3GRlstXKblBQED4hrL6IsU5ENTF9Jba
shuOwXgaVAbt2EqNZK4UNZ5hlRljviPJbGhKB2kzFPXFdxyRlOTBbIVlpAxpiUzHtyi5Zq5PsGwE
+stBn2MgjB/cy8U6Ozf5J+5YjzXIC6KRu0HFCEbnnk562BprS9AOV98xzU8MSDTdsYVUq6SrWtjQ
4u0YlY3+AAf2uk6/NWWXq284UcUjySSUP+ye3uGEGklod9JbCcUSi0PsMv7ZxOzhDLCA8BJ6RhzH
703CK+5f3oZ18+5UmVCTwC8PBDcfmE4Fhmtq2Hu6ygwdvLFflxht7pN2546NU3k4GjDNBhbZ+2ei
MIc7g+uNZYyKEyHQrl21TBfAgW8PlD3IKMbvm8Ka5e4ZE6Tfrlr2iZ+i8QK1Arq7ueaYJ1+iNGM9
BmcrvYSdn5lGw3vPjehPEjvapMokK6wkxVnPtosvqNuSQc0PRVA3be/x5qUlrfCq8ijgMuoMymdl
ec7fvWx6SzBmkuYWaEfi1UZsdbWWACHT1KLGifuTPgaFfv032ETfx+xnijol+6mhmOJlccsQSgbH
79ToBeX31TqM0XkqLZh229W3ZwP+Njx9W2OyvlOjE+BZa1+CUhVg6tNFomMgWUzTQiGqWZQWyTKk
qCqbz1dfWGMIkpJBk5qRI7p+3VG5GHw1OVh3XHTsyUUQ40PpcOKHXMT0ysgm89Iqnk5W7N/1bOF8
ZWZcCzstKY4ql6Ecmwg8ahf3hHohOhF6nqU7hIaasCqoNcN4edxshWX65ZfhoFwk0m96s0l6jNBO
wgKc7enrsvo+WXxgT3aZ4NHD+KgBE7yekD/6bPTR/M1cLFQp/i6X/Vl7q6ZA+MSn57c45Ap889vg
f7K12gK0TrJ4i8/bcphwiZ8J4MIs7hmE2QNg2gVskOwBxZo3Jx3VQMYinNA05XpA3Oq/j0mXH7AQ
sEeR8V1ZA4rQv/Jn0pceFldJuF+dAVqeHBkfykH2VNvrJCo278z5C+x0b9OQYyj4YnSn7paaAdeo
2xBoQdvEDlLW53H2YK8ZkHAdAbo2zRP1GayMRz8YC++rRe/UNEHOJF1ZI2NDP5zXzqCF6vJf5zv9
Fj3mdRgCQEFsJpIyg+KyoeUj6rQhfZ3P/4py3xIYP82wihzARg16FuBSTrOQk21iM9/cnzS8IREl
Hr+YSfdU84UpPtwzjwNDTEbgsKqW2TnjX/Q9fNThiqwLAYwbmDNBH+jtQhuVnpALcb0rihloUG9B
61GWMImBKsJZUVkOKmLYJecpYzboNgmy44bWxGpI02G38Z5Z4PGWcBdpkPU7hdiaeJohTl+8EdVd
qoc87YxO2EEu2CRkNbqVMcF71K+Cp8GHWbsYeCyq2QGhg0zkDAL4NF2Ky2aqjvQA+au+0BWX79wB
bA+Sl6TAfgfWpARJFhysl5miXgmXT3LG8Vi/+6+JUZBbM8RfEysml0enbsyQO2ExAP8ERW/HnrMG
vUUVr3+7Yc3kRUkq3ZYQ5KaaFBnW5Ljx+IYByOLR5kD50E1IqFSfChpgFeuM2U9NOwNW7/4qqoaj
/JnLRDQZREvsCP5XrkmBfvxakYp4hiMN9WS1coEyYXCcW2xRjnSJF8i5P/53/uPxFTUKtF7YCGMh
SnHAP6JQoClzBMClenT+Jc61kS3mim6ltoJ0/hNFfYpfZVwKl7s1co9UyUkSrWtHUWYbzxTMwRZR
eIrvZITEa6ik7jp1gFK6chikwp09vQnFeKAAAzXXMvPWROgPgeodDpITRiQkSP/g4IErK/TDjqcb
2A51Gmicvnc8PeNCTjSrX5N5IJEo2jDXy9+HPY/cGaUxcx/o3trc+3oP2IZa3tbXTJ2YZ0nzhPKR
hNB5SO4dq68uPNPeHaHshu1VJqv1I/wcwQq2vlLwxTFb6itruThgxNLl9L4O0xmsqaTDIeKuEooI
ZAtBmliuuM63TCNO8dBz/QpQcXS1oKlrt0tinJaOOZcCaGKck2kRJV0TVs3XE2YMUw57VTXOa/bo
hT6SrMkDWUZ7gy4U74+9v3fuTDmdnmovWGgcU16Y7wSnw9WFGLbdFzRGy3ANBBcLj1IS6E+8R1sL
R45UWQOBPFxhyWwaLwkWlgWYF6Yhz89q+G9db1UjLTIgsWaM+cHZpONv2ZY8dIn7T5EfcCgu/gPT
LFiPFOVtxQm25l7ZnqX5E+hejweItJSMjZRUWGtAbzwq6CmCV6ODB/C4y5s6WdS/xX+Js62NQCKA
2QCeJaAZFX7HTIY8qXVfvtJnTPSv3qkS6agUEvLkGIkfkAEOMKr/DG6gtjZMLJNs0+VJl606/IcN
1U2L/dbbDpqvb/82x3ITCW8RjptKCQwsF6zbvkJGlrwCqcJDEcNv29tQ1CyZq2vJkLM7Lw4iAhnk
6xctBi8HRW3NIQru6/eGqBqNPqDgCpAKuE9O3auPxUz2/HJejA/V/0m1rtZmSLRuQG1+Jz++pZlV
jYuvaWo5ciQFvGt+bqi3FD9lVE5jCWUPNZtQd4NWdvL35ABckXDnpQXJnLt02OQZvw6RZ3WIoUbF
aZq8bxwvZgc/AvXPEOrPWGP1fhWxTiZX51M4iwSq1J6jMWU7GtUoUrsackm47drR8aU81AswMrs8
JZeUoOwFvyw7MzhJFCvW5NEgL8mpbq451gkqpQckJGJcUXdgCeeOsPEHjFofynvmR2JwuhvKGbsR
4dL026zDWz7jLpn7Lre+UUQdn36cGUIgrFBTVTxli2UUV5tPIrLQ9kCmM9HIYSgl8lVv/2NdTBMq
GoyvyUmXraMEUFpeSatllLUpY8eQmjEyNWK8k7b1SIUiGFOE/K72bImMI/p+PIT/1ic5lbV+lpg6
q7epqfajEKpBOj/dwQ0JrugDOEtSeOmMyt9Ef8QPyi2UFUhhlOuP7MjaHQf07l20VZJYXUJv5aFR
X8p8jGRBEn6qTU8ePbBcO8+rcXhFZ+lWI7xPI3ekD38VSjrG5ubK/wXUK+4lUBus5cxGMT/vZya9
fQ4XhRFXzOvVVumyNTgq5sLhApWT1x1KjoZ1NXBfUukfhJcw6paOGYfBjrMysRAJo7nRu9J4CHM8
UXooJtl9HSf9gucnEhLvPHuvik1Z5Tu8iWLNMTZqJ8QqigkO4acnDTDo2ou1ZO9TQXHWxY1mdQ39
2JfqYBLTzIcNVVjuD2xgKLXybFMd0pPDm2Kg5UBPIXGsLCFuO9SKZwE6Qgl/L6aqDaC5M8bmCXBl
QNcYacGK0qs+gSPAhSKs5zn3baHHYx7o6HJtzNVajD8kKHgQ2etg5z6pIa2pWkh3FO0rA+IrPgBN
kIHsWykmhUZ1zrHTFKv9mJXMBJHufl14dgqgxxtF/Ld6X1RuNJIkj/Icj6Q8jTqEC0H/jxlwip1m
1TRJ8IMVQSG1C7xDQ6IPQNSKqeEiSdZoOeOCumG7Tdw7hMBCavEoqUqe19V7M+Nt2SNQ+DbK86c8
L0fqMq6XAka/o1EqOoVTdHBjD2kvceKO5loTfOEBeT3ub7aW0XRyOv98HjZblSIgCfhvVJDjkAUF
IpQ1vvzFUFpuKBE0N5LmAPytH63nZP++yr0WrKuCTTlB+fto+cFUozH2vaQ1nZzJ5zbcadxyFEop
9OoXxLj3v3FIQnqygsq5UaunIYCctpPBs0xIUgsEco0MP/EtmhSJzhzhM+hJEfsrRk6VioC/QQqG
yeFKG0ps6Dh5YeBal2lR61bicfTkZNlKE7F9S4EuSlLR4/O1/XeZIyAk2t8/ACn9ToTqjBr4lc2G
4AVCgM7ybk/76R0ZtJtW8jEWKouPqkp5qSOulay/XLGjYfR3adyRLxbyZX7U6ie5erVPn0rhAbr2
xAQPcBrd8Gdmu5mg6LwtKmmtZD9z8/Az8t17JmH4iY9u+GEUiGsg8aihaCZkDQ2T4koY+9dLwiXI
f6QSSSi71mCK6lRn21Kdfy7UNJsnQxSQWiIz9z2y8OJYT8nyIT6XqZWop9Vr/Vg8/8HVE06qDc6D
6F6K8vyJTJHK3ANiHzTSMGvlKz4J1QOeEhNf5qjZ6KLQYR8XFsZQynjHiGPE8h8mzPn501XLPY9M
S5byYxprZKWaI+YIQ6JxgmPcmfy3EEnbOa7gxarqJd/Mw5bjdpIM+xs89sM6hAGyRChUCgpxPgxY
EOM+BruEC28WZ0GWpS1hxt6qRnOgDnLrdYatjNWdJWIo8/NE4cVBkHyPZmi346VABdWgH0wMFuHY
0yr+0vBdmAffMf5LtgjeRO6+H+dUIqb6pzxf16nKzG36Ee6z9t9kprZPiwAuLau+gFrqtPNcULYK
iL/dMOjfLZ1gtH3u/f9BHXJhMNr1zJDzXYVkcM6Z+abIqeAdu6Dh2M5ftHx2K6xr1oiHqGC31qv4
kgXnht4BDTRHaCZZEJxUQI91q3LlOCIxRqp8stEZDoq5ux6S+mvS0ggqK9pnV0npOERU35Y9mn/u
bVAxGV4ssmRxGkEAOo7EuC5WYCJmV68lAsHITYV5L/+xykbLg14bW97B22e42m/Faqoiyq94YfsW
/Wv6PwSq502ncYmmXTH+oNd/KjAuwQwlLQFaEXEUlQeVYCxQH677XzvB2kB/TUS27XeuWC7FCOFe
s5OdRk9+jydOj4wlPirpD2cI5YK5wi+1nk952XsiSKvuOe+vs7T8uvu1g9sWtkIYZ/ELcR3auFyu
6lTO8+OdawknTTOaxFUXLZ0SbbtYqjBdPeSp2erz1l3Sfas20FehT0M3OX+PgNW4sii5Bgbk3Akt
dyUAI4bwvWpZDeVV4+oJDgFd8tcsfaShlzZBWtPwDZoZcjmrlRHNp7oW+v9fywrmAbd644O271pK
nqffbE0xrkcrUgzE4553JPdJJKRtxj7VfURAl4hFPTs2m749Hu9IVFOxnq6KLCOKUo99YiFaFdJ2
3rsOZGrbXVNT+4SpAlyCyOn7YeMDogtDC9gG5kl+UgIViIQoebMv1hJdmO3q0wNOiu/gwxURi1mx
LD0rJfgyDa+B8IqMDEzQ4O9QbyY4fwBT0rptVRQQovEt9zUuV1BA/kwbeCtB1slmSD+PZbyb0IJd
v01rP1VDNVMidm3UV0DECbIbYjjoB7i3Ssh4iq1/hhAzNyGfPyEneQ2Nwqg7YquGG5CfjK0Hdm2Y
dS5yjEf59/VvCvudsM+qybOHxUB2jPEmmX+Fyr1YDH/gPUsJztvbJ+6lIekZj1IoXiRkuBaK4s37
Gu4ymCKTASflp6zDI5TltVXuUgddiTEOwzPUmrnGFD9GFsZ/MGLFPE4DsH4WnRhM5SRF1padBuEM
suQslmn9lvdg31UXp3ywAja1fPaifG7kVJO1F/rwaOgda/LvG7nOSv9KR5qYDb5dupNDfOhSF+nM
QkVc909qIyc8fu36wrtAxr36fbYGflrcqnkYVKu1hcBrW7uw2dSN6KJFRW113e41bzjmBLk8Kg9N
JY+bS7JtE8CvTZrkDZ3aeQ6vxx6+/oNqJq44oN3KuTnd0RV4/06/M4syxJfeHVJSvTH3HfunbY6V
HVJqgD58qKOPnI/9eCcnkTN/HJbn0kg0K+Qns0zQhkVSV4g1LjMpo71iiaaYRTj18RkZlZjBsw08
O4sO33JO+Gs/PslTaZe5RYo0frTYaxhpf8UVNiOsaDVeeqD0tqukHDtwIjjOYjhrsSPPidUXDryq
VhfGrvEKdyN0mDNsUpR049p9YTfExgyNgGbP25j5glYCcLBKYmj+7sueEAdHtkhywc0+JJoro/gB
gpGztaLgiHjXUXiisbeDTewG/kXSTtWBrwbvyoyn8M+1GZOudCrrebnpwpZ5VoCCqHorzD8RZ0qr
gMXaiQqDYjTjwYeazETCdVeNiBpVQvo7MGwBy7AUgcitVAtMeQ3M9Y/CP89BYHpQO3fdDbqc8O20
ypo5APPRNjNnoJo4vpCxTOw7STcGUTSHo/Q+aPA9d+fYN8tUzHZ9B0OmiuOsx1/KM66xGyVGP9rI
jICI0qaw3mV41cO4AUNbRwf93Gl4fp5Mj7xUh4cSfL817qEx06aukWYzY4B2Piaa5EE3a4wWiWsP
943x5o9ioRXz1lYzcpYqzAuW5tsz11glh2L8cmCmykJXRfPsLjGOMsdWT2qv6/38Rtc3fkZAs1Va
V7g6XatH/VoHOntI8la79KyvN5rXMicr8olOHTXB528RAhE4Mr0+/ybEFZBAd3P0AyAnxoVS5BXx
poClRp2hT69RLvNfyNK/DYBPyCDehsquGbD7+BHGoaNP6DqsnfVO9B0kJsMWwHucBSybNN0xARWw
oGdLgFMU2i3y85f1+VSelS4/YnA5kuJZhHVUGf+nmHs/fAufJNGx1VWHlNTfh4xc87A9jWIbg96A
WLNT3Pgh8ob8jnVPpcchgiHT9KUA+jnk6EwEMc+1U1y5Bt0VUZsJAYQmfL00BlpCQmvOPizMdCqy
aYXx6sU8R2UGuEUAS7AC2JawxDf+ixZy3CgUCS29Kw361nDwX3aG4PEz6Gsr8oSpLkxE97BLp70k
izHPWN0VBhoviqvk+SrIAMRoqP5bqhuPg9eWDhxnYSMook19IX6Qi8NzhwSAtrEv6NSEG6sOktNw
cbTQ0mNq8Ok6tcjr6N2qsRw9xqPMBRcfsHeJX/a2ZWtF+q8CX0e8UouIpg402qydN1Zh5WkaYjGz
+/xvyCtdhec8jm7Hf6o68i6ryYymzWJOWIs4qZsomBJwnRQLIVlVYsN40p8YKL2tHLa7Bcoc6Trx
W4oGFlLwc9/bfWBUl6142sx9HwKelEmQs5XTY6Oyo7Q8zZFm0ix8ryGDjM1bWI+Je+bivq0c+OXj
XXfIRD8usxJLYU2nGJLkj1Swj390Pxn82yKlyZF5vYpIn/7KZJfReVhu3KhL4/QIRxA+zLIoOpzb
01KPYzoKwVMFMDKFwN1pTd8OG3+wG8Vze6FVCXX4wPoMh7Ezfz0cZeHMv40RrvFpYHSMnJ6tlT96
ru9IcgXVQD1eGxGnjOMif0WoQ5NSgypz9HD/9l2f8shpi4FQaXdyHDgbX9BDwuCvHi+PmgnKmxPS
b5bAdAapAgiq49n5Qv1mgqacI1U9OlX4JaBayEX0IxQYO3bNrTtrZ9bsPiL6TtJmUXjvd64+FmTF
3jdrNz5xGc03S6dLdolD36U2XeRV+1aDc4GeUwod36OlBmWlwGM0W/dcgaJTOLNGz96syZLIuK48
V5bAvtRG0BY2xdrmf/FS+owoqwrFwn+Ng0HCMihzB4rU9/WbTNweIOlKnWXbc73lsfxM6VfcXSkc
HcA1MzBtt23b8wj28gbd7V5e4GNr9xKiQszk3/82AMc/TCNFLYY+xjSTnM4CRQmbNh4PepQ1E3f3
UyI+P1DUFXTh7BAm0hN/BghxwrZZQ5LYvKn6Z/Nmh4C9w/oKdK9V9sPhZs1kXV4QQGbUF/GZA7xc
8l79F0ZwNyKpgmhUmnzMZOY2ZSbbQpMPNFo7oxOoAvTPTCq0tdAYHHOex0CZl7vpkLmPTe5ozHb3
qsxQCcGLDRk6/1XaZ+o8gWfCBwGqwfpFFkQuvMcGwbnrz5JK6cCtYMCpm1/tqYSTYk0Z0y30bNMw
mbW7ELL9g50FuUmvCv3EgTrTBUE3zlhDbT47VdjPbodjUKWm6HNDjihIuF6AaRO9Cs1OrslbJ647
DuhvT3gl1iaUYfMEeDEbbKKvsPcvtTdcpVWEoQgPDj7tvERzEV4ubk6Cu0M3UYlgblxPNYh9Puk/
uh4njS67tqM6UqwvSVUkneZxxvZSla/WLX3hx1NT8F9nPbIyqmmWsfGtFNDXxNR8Y7BE6770kJNt
rm//ybVN5fuNHKPIukgdZP3NIQq4khhZRpqHpB/e+Jkfuhf8VjEotAp9LFVTVDr/ScHipEwCQ0ck
yp5S5bDgYV0Mfcv1E84AK3oLNr1f+9/tsXoAG8ik/EUT4bmsj19hnQMaQNuet6VmjxRCcX1Ybnus
I7igArMbkQ8krC7BgtUOJJ2gN6P45eA3DQwrTFsOI95fuSH6Lnl2FBrFXKCSOqInmyQ6xikRvsyi
gPbuv+BYmevB3HW7G6AYdfpxq/S/etHQmzLc9EWClBgBIMBsUC+gwXoeWO7cKqIgptRak6hPTjxu
o8fSGsegpH+3mtSqhLOH6FTrFxxVk8Ug9UlO7+52eYBSUUUQPReuyehDhC4L6SjXgepLJ9Mqkqt6
Y57JJWLn8dIfbkkecA6/D/4u+KtIQeNuOz/2mlU+ZrNeWWAF8Hh83K9+sv3Y0ASM3qyNlfJjGrN1
ZjZFiT96YHbVmbU1oLc6/1D2LG8pWwr4Ay6fSAgxewdgXjMATAulyxHpZpI/ekuR/L8hmSQLwhEQ
ppcG6usuccxTbXu29b2EBE800Ren/BpEx3K1yakXHFDYn93j0uFWHW64RR6/emzfcJX7iqTGdjvf
UWxOfCBG9SCIM7olmn9XKWoXE1hZ2bimzbr2ngFwEGjQcHbElG+alIHkmcCZmCKR71FJ7vxRuIgW
pwSGswHcLdosfBRNKZD4yFYxW6ST+V2wlgT0X1J45rVsWJBZSUD+GrE6PBllPAlgwVT33Ohut7dr
AuYLiMG3eqwijvYC0BZcnclwxA3fwMIoUSsDirYIczQfZiWZS3f+FvbTk8gCfPQYvB4kumZqJinX
+M1eQoEWvk9kLg0h0qjEq+vb3ePkPWOzrcV6jWFBb8IpAFhOOooP+yY7SpBdUcH3+BAkY6hUoyN6
twK+TbQuCPc+B93vy59fdODTqjE+Z2V25nmR5cwbRCxz3ZNxiQo3WXCfwE5aF/QuHTtYYfOIu2az
98ELHD5giQpkOL9Cbk1ofSX+51O/9ctQ3P+7nT5zBki2GMaZ37x1F3NQEIcH/uT0yMqK3Vc9upGZ
Nk10hfPBXGj9ZJLpkiTxpD0Et/+b5ufaYFo10OPzdjUEktmxhrm7et67ROHJwtJ80NUNasGv8eST
JvQ46L76QKMiL1NyEip69bHsmf581sjMSqiG8bDe0s+uHYwCktQpKUIbDILoQdeptGoNXwa5iEVR
U3bwfswYI8vJiOdZzym3IaAMzcZ35zH4/02ZdglHdjPVx0w4yTTs9bBbUxJ/8jkihGSYmMK50LXV
EK0t/vL1SmHeGtoKbnsrU2h0/5zXXwdARn0RscSEtmm+Os3j6m9Q2dBVEH9xtoTE2+5RYqj+3CHV
vWmT7J+7OdZtLk1XCyEE4RQIuWoERLpGkoppU0uqrQ4YFoG1J7K230wJjSdA3D8CalqkJmWCk15o
9IgBcZtfITYVr8HUbCwOifQy+CuscDSpIYuYfG6wty8lgjmxybhN0nZzAWkuu5Seqhjgc8t8uZ73
1dyTYiUEH8UXQW0qQt3UlRBzdCxpbogLeUJU/Jb0CY4EfhZ4N/+nRN9V+k9WUb1pGbMK4StYYyyR
dLGR9jNj0lM/JlqFdHboSTRwNlDdp1JZzhmp+pl+FYHT2BITx1QjHDwWJhVyofuE6X/8DV5RyX6F
2eauGHMqnkDpS0uOpwnOIYTonkL4USPGBFWHyOnQrNcKh6EOAYGqE4WXk2wHrISH6iazm9YCOgfp
GMBxNXw/ySn2bGOvhcfl3abHShbn41ePo6ha9Y7i/OmRT5lFI1aeVKKZGyfIFG7RTDtuBqEEQFdo
qnBaOoedUEioMHesKk05hcFNbMV0Sl5uzeF1F+qA/H6fwHUq7MuieozQ0Rrve2PdWpej04M3FLpi
UO9CbficQEUOlWsjB58RBYRbI5Rm2iwxUmuw7i28PWAGxs8mJRr73bExvowSa1EOt3Ggkb8bUkCG
QRPtllW4V8Vg39RC+cVQmyI0NXuFpHj3TlGxIrMUfYlsYwDJEvu+nMR5aarQRC99mEtIfAKDGw0I
pDQKAHyQmjB8c6n4P0FKR8lmG1Wku74ZKies7V8r4aYt+Hx/SV7MlhV6/X+ZEYHgwRazIxPzsal5
+H/4QbSzv8cO6oPV/hTeTo6r6ZHb5e6yeyTmAiIdi9DrnftZQRxM369s+HVZIh4w81kdW4mX7EvG
0Cgqh9NgeLq6U3S4ryDFwDAry6VpSMNgz6X52ChjWzqrtgpyKBQF/X6q3Yt5HhZfqzVc1u/phFrA
y/caDfv0fwmCtzTCR+n2MdIoEfyBd6E1cLqAkuGN1CWlGHVljPt+lpOBS/B8oze4yKsaUuS2mdu6
FFSzqWtzOx87NEsYy16HgmH9P98HgxnCKpgPhU88lMQpBAJNPlKDwdTA3l7gB+UdDQ6M2nx9XL6J
HOXXOc5FSJvz8zO+7Llr8Z9dIeKyfn/9wuRz2n7Er4YWcHJy2fj4luGJcsCdomJrM0J2b7+5hIia
AkUwLXxVUab8aZK0T3ut9YT1N7ufuSloMc4PLI0e0xX9dVsgJIZ16DOB6eBiDAZ332F1pFlwtLGh
t9ZyBiv2UHiCU2gowKceRf6CmIO5ckjdMxo7E2JP2oKsXM7OBMXfsWtbjEUyHbQPA62M5DYntWzE
oDXxNKPgSc9d6YxT/aYSPRXIOtPrggb0d64uqIQXI33bmHgUp4d6RRkEA1I9o/m+tPsOCFqlCHvm
7hAYMDVTfElHh1zRyr6Ux1PQTHUvyz4/kYAldEizaGjeh3lfnIF4+pa/VGGDttBIvv4o2/0jNTyN
avYTHjpIfWw0WPODaxwpkzTxqf26B4n92PEMcKAkOkeJBYbSCsgm25ps0Z5HLDyQYe1lMt3bk+Ym
PBrBBqFU/CKZ/CtltfhFuTv3oGmiCcs0MrVpbGc/OV27ksSmf2+bLkb/ZqjiVV4dBpY++4UMMkXt
zkhvyEuIncbyciMzoE1vGisACljvWMBmwribe9icp7odCsl9N+QVCIooxUtRQ9n1rd81gv77N7K4
EH1pP5sXh4t0zHZImMtIvsRcMCv6OB9Aj4XNQmjQNOdQ/ucfHaED9KyvWY7SpZPHiwP2+BnJbB+E
rZ3RJSfjH77EdPYudIX/i0fmKFuJpbR+Ucwgzw4wwu8V7csaEZSGO11cVxThfwPgHm7I38Wmrv8l
gsZ8p1m83fauHs3/f+tPuLCFZY+odYMRSaXOe30RpLEYBa5lJmGtHWh0tWAg0d0sfcW37uoc2qxg
99JalEz4y2HTKKYLEQxeO+Nbz1v80H3M1a5Q0wfJ25mNcY3eh984yuPDRJYGFTo/vluWgPwlsRZ1
Me/gtSPhPrDRzoWQQf/R+cRBLkGNKU9d3AOdL9I0MSCCitF99viGEkt0equnuPuthLCRy8bSA1Uh
5J0qjqQ/7748hmRWAClabEm6QLRAVTvdpxeO2NkiaRZtcFKY5BdS47lNgtIR8UgvLBCMPhaDxkvr
U36hwQdmzwj3AyHKc36G0IFBaJOJUm2xxtW4KwL/13vhA1crqWVf3GL3c8tcmZ8o9ZXZlfhHjXT5
LPxlz4OR8J1qon9zMKFCCnCduUdZt/3dUtJ3uKrRvuVvUKm58xq7Lo/qeuS5GD1a11CmwJKAyElP
GYdS5Iol9t+zsvvk3X1R24s9xplLTBxBluZ0/RGJd8FqeBFyzdbGH2GZ2na48Efzm2pODUN5NU1k
foz9ll9WAM9+IfFlWHzDUKLS6vTb9rXdB+SbzAHORRqBUGjLzNjdcionzm4Ux1HEDjB1G4ZScKjC
Llg47wr6GsV4cFDI6Ud3+YEJG8ajtaGfLdhEjaXdPsu5qc7X9EcvOojNhu4gkWdx0EF71gjZXIon
FoqDUDR/OWJ+VGet0YGDHUmX4Mf+rJTr5ydsjSLFND+l3p5aqS5aOb+gbw/eGHqQjUW3nQ4u5sTm
PakymSrkdsVosbKeldjkLmiyxglslCsg5u/wfDa0VLTBYT5gvly8qt6FTfCqrQlZlaVirJpluDaw
36VSUEYID7Nh+lEWlGOuxwGZEK1Wi3N04VnYRdyo/0RbTeh6wyw1gsJ9hNI031k1OsvCwqO1wLVL
0ORpsF4zuN3Y97RWFkqPKbfB8eE7l/xgkYZhRUw75JuW43YW+mZ0UMQ8oHElAaiw+agJ8c3eba3O
e4n5fBiZfYJX7sRqp+GNmkONAyl9XwI//G7d7+BwGtMV1On4cJtN9K3drhUzDS79rcq17KlTWrdM
1OCpq+1YvnsCCiIA2b4kDvydrOk0HV2CKTcUZYIGRM3zcQKRPr+RdPQSo6r5po08762dKlGkPvp+
b8pu0tEhpCsUVrI6ammwY5/bNhBRbrn3t9a7AEsos/Vdvqt+C+9tx2wYo/JBNFJ3cB5/FTck73Nk
7ymZWhlYlWerPKMRwgBeEiVPSkI6S49ZNzK+n32t8m/kcpH/sNU8duP4hb0StJn1713GhcWlx8gt
fEBCY2wpo2LRlEC1ScIM5LkW6R4I3rEcBNxtwyWNUiyzECgQFqBRBRTH0GJVzzkpAlPt8iQlvkUS
fASmpfOami1EG4rLKHfLrBjyZLoMXImE3n+aQ/VmpjVejb1dtYFzfMy3vjPmWkypMwFvIu6mU0yg
s+0LWWyOZ9djOMHICUs9tPUTLqqLS7HY/HfyMlsi1+VYRvY2MvcokSt8ufiSiNp/FCYCg3OURp/5
HXfL0USoPkCwP5BZwHSjLvwSukS2+ttwvIgAj3v71JckQiYn+akDT+J5vYa8TXDjc6TVQMUr357t
FJzSCPHZK/CkjDCx1AmqGoppPvqtvAecCwmPoiyYZUjKRhaVBJHXKzVTm9Nfoc8U5LcHQrfSkpd4
ntggt3gracHNx6oJkmQHekZLdOtVyr4xWY4TmtfJNu8aHeUC7zI3qZTQGrDIVklSD97TlwZ4jzTH
PfExFI/nRIHRabJqp2lSLLHasUrxVwpKetUqcrRPu6pIhOs4L/m4Qr81CXon1Qm+hT7MQU4+Sm2U
xMUWUMhzxf2mCAc1cZxUy8wS0HN877AxChT9X4Dhc2QdcEVAC4qR99zY3Q9PkOaP0GIo/a/3ckZC
FPOCiSYPeEA30icAJe54mFCE9b/KiadQO+e64u2Ryl0fpZdjdRe60VTu6OojkMA9D0WaIeuyTF9n
+zS6uftF17KTaYGNv024NCwcMCTK1g35+DzZWzKcpW48EG/Vs7qvcSAnUQqtOaK2nba+Mif4ntKt
g5/TLPAhWPN9rlsNQ5P2mRUHukjK2GkRVAtMPdw5UN+6uALsZmktqzKV2nFbGOTn7wdY5HtAV1CL
EXnekHoemYgqr7h4VW4YntDtvQVW7ZgOho3MD1+Vh67a8WaHovm+S1xnxZXrKatUTqZi3EPmIuIw
HMrzXkW58Lus52SRgKaormfkTPPxRmIP78xkvDvXkNv6Zr1/adlkFzEuUKOyA7QsNQ+KsIBQg6pc
kiT69DM5lDKTofkpXPaU/0TUj25Nugwb9R09BIAI4Axfr4Nk5nuzgZxjokhK8YPf1Trb/xneKmGF
p/ic1SgA0eqDkWLbZGwCU0XhALtwsPY7TjY7AJjyPPROxJdEvCdqjPgHXU/AOrgPRMRuXk6OXbX+
cTlvV/ElEBkDd1CfrR547aYFYpnkiQwTE9W9iNioKd1c7sO5utCL8FQ0KzBSJV5YTSxLgwVREjeh
CGPkAl3HSTGPh7FRvVNL9Rz2Iw/EmPc6eYgNTspvwUTldapFIXSlRaN3VJ3aJvxK+gni/H2GciHk
PlfYnFiGjheLk9p1D0/I9zq4AEsRAzfZ11nQ/0013ShzXWj9KIaKzkapMAC3VklmqJGf2cc1EpGS
qx4+i6a3hV0RzL2LdtO9HiBe9Tuqb1cnB8okqSl7cUsOd+QweNvPFU071/SMFLLo0taAh2LbUUrn
pMGH95tKExvNQf3RmjatmlVGG7CpVBY0ReVtroZtkSrRkejr4f5Kc8JduDFjQpbAKGVF5vvDs7z3
Fcgr3803X2jdN9csrn3a3cP0ySiMii0vraH0tb6FHXLqqAVy07rQaFT8c+IOd/9S3Os39oGUL/zo
DcEDKqiwheJ5N9d5hnlXfaTRXYcVIOPNPxMJ/2I0b8IDaYgY7HR3auto14Enijf18SLB+51f0tip
4RIYowgksr/tFYnWqnKvxYYHvr6ykeO5QIExqlqJat9d2oFtUtBtXAamS0OFGtaTa3chA6cOKcP7
LoeRN+m7nlZ7O+HvHkwBQFsISHMVmpIn6Pzx6jaMydE/9JGYh/Eu37+y1l8iHOFIs6r5a/38DiCj
TYzXN1TS5F4UjL6bdWK1t+qdfrR5Aex+jUuFUclANZb+Yh8wXadBcR0PYa3gLsPGq0uLsgwNm4QL
MyIJC5eR5U2eI9lfA4nw9gXvZx4b3kewG/mVJc9bRiojC7Zzzn68x83EZDWEwjoIUmoP/qagRJof
LjzaOm+icwwagwwly9sR8K64pSrBULU5UV6dj7BUux4vWgU+NKy4G31zVRoZLLChCMbHIAFP9DhC
9kcEya/gWKGWplZLQisLbgJD3nWFR5qt9VhCr2l+nUVCQWKjcgiZrd+3IBFcT4OHcDwV99WGrEYQ
bx1quIlHv9X/SPzb3vYdPtHE5KQqivDcWatDJqGVIESh5VL5EwyQgRnDDK92PDfQak6PwJorx+l1
I6uUYGZW6OR2LiuXg95XfGMl8Wqhi/+3TExPmGpygqKE5anJVrPRR4p+mczzxFSOFaJxNDiak2za
bhTSUM37dFXhfvJzDs2MC4LhkrOrypO3hcc2lL/az4M/AJ0jN3luC6PSdei+I4bfHPDWGNOsAzl0
05WvQ5q45xfFi6v5ViRcL46ii7Dr5FFjzELpfJAnT5pUWs/28jDeux06ZiqJz4unddZlruWfkOlr
Zxk5AuBYfLHXqkbIiHspSJD3SW43/HsA4AzRotfWqOdG7o5VinpAk+9otjlWmMDDQ0gwP0IiUi/O
CubV4WguglMswEOyV/EvKUnd70v8fGZ152ta0w3tY/CiVPZjpHw7/KIjpZKFY9vkKIn22kdZ+h9f
U+Em2eDdpw3w1EZIB08d4GM81ebCz12QUdeR3cUl1eR85FQ5/RChfuHl1Gw7+OEMgSaWak53Gn77
+ttw5A31xDdbfgjA3m6FwjIl3nLjdz/UK+EjZI57e78Pb+vgl75a3P9NZPXPHUdzbmRSXI2y2y7R
8Uu5u4lqfudJ80j5qeBU8UkWSBW+hSlh1rWY0CD6q4Yu4p3Ir5l/ZmAeGYiDVbFRsl0cgSljuqqI
7j9QHna89RsHcBsQrxbHXFtpBytSpajY/xtFjgucJAqMgWEPCjzzGqlH98z2Arrz/jjPMx/eZVJb
IsCUEktogCuubtsAM4rwlHOG+8pD+XZCWdeuVBfcrVrqg1zueopdcmHgw1lH+lZllFM8KIJ+0ouc
rwr01/GytL455ULwjOswfCVwKrnEDFeEiCVslEB3nAT77J04NDKPK9jQnQXDMRnnAUkkA39lD5mZ
lU0YzeX40siJa9eJvs/FL9b7KVstYdiYQGf5TWHHWm9VcdmnC6jMWBx5AlhH99LNQe6pE6T8RH6o
Cj3LF9q/GqQO7yoA/x1z4lYo6fftD0GT/mCC8prr9myqma4yJYaLihBc6CziSjgTE2QTekEqoe0Q
qSKpGS5pl/KeV7kYUlHbl5MKb3gKDQiWR2znCO5GD1Ie5nt/7891Qb3nzCKzG4/LtGDWR2BEFpmY
VrD3BNJDyYRxjM7OmI7nsVyCJ4jXn//3an8SEdMD/N7MSy85tMaLZWhkvC0dim0uz/1Uzb6PPqN9
anNAhL5Ur1wxT6cW1ieChFtFxvAOnPziTM1n1ST4+Gx6sSH52K4ld6DxHIRSdduZA2N+4LNcVmar
GplN6lBNlpxWvZ4g+GxTXprpXHwW9fsUp2yN5VOpZCfZ0pBOlurzZckx7ep3UTxB1qbDfGWE89Jn
knnKy/0tlV2YlkEl0WC19heasvpWk7RfGiCvCg4RzhcVdQGUrHjSObZMVIPZEHp/ahdRdwkPolVg
WQc3d2/TqIDLBQcZDoM9TIhHf9ZCTOEdi0IiV2j+hR+3iJUvHaF6A5H0iWDz8zE9747mGykUFp7A
WsilNLngWFSx1xrtTgC6M+4trnm6xAnj7yCqEUiATsq9xQcTxR2II/ZFIAABiZPhUn0fEeQlwdbi
H5SmWxu+d2mWoiqXh8GjxHxz32uOsN6HCGCUoE+OBn3KTMXxx1PBiRS4yHhniHr1yvLkTPRAAZPA
mGA6nbl6uFgcWZRqwM9jwAUE4CuwZ0tpPB6Rd5VSXibQG8XC/MXs81SrYkUosrInk+zFFICHN0uf
WdChl3z0ALZL0VxVS/dKNzsB5ejmVpVejWTYgzWttmVCXNA5xBjHVv0H4nC4d0r5k7kvzY+PtcCF
4B1Sypb78J8GUHmzstAm+YQGsxKKo42nMqnm2xnGeWFxTJMPDiayashXAIaSse2dMqwInG2zfciD
P8H/UWKfGHj7Pq6geWSQ6e50dJkzU/Brsdkumnskw/CoRJkBnRKui0F0m8ddsKeMlhNoQUg2qSDB
8OLkjhmWALNu/Xu1JtrUg2mJRvzcCEV39ifYhPrasYE1GTmJo1TMB2rUYODcopWIkTprUhda/uU9
ENJ0WWI2tDsXo7uJ1b8IfuySxTb3CKJmGwUF3XwnRdVHRoQeOGdwXM8l8j1LGCHk2RHiLCU5c40B
JRzRO76Kwa9c176IREWLlmy9EkUEwa9rkn2jo6txjKUmtGpa7meNtRknkk5CbhEO+jUN5gYQa9gR
F6FNyvXRMEXJXli7xlkgj3NncAaX/tWKDtp31ORE2Or/35VG4eCd15Ok2v1yRNLaKorblE+Y0KG5
GZxBsXYUPFzrFRgblNtRtvzpN4HrmiGZMAGqKZrZbGuAwQW9omgMv0lH1uinTQBVJhsB3HCb1+R+
Cb2bHpRgUrZbazFysFvfT5jEIY6g2YXZ91PBiyd98IWru3ZlWS8JBI2zpc/S7i1yheIbw+YuI0qc
VAIpz+0qJD3wj/aeN08OBjuRGAd4xgoABVcs+vbl21bJ8T8eygqPVhg38Xj7NQN0nD+a5kt3osFz
+tFMtdMyGBBWeCgjBrWJRiB0w2rCMvXTWz3kCmN816iqQ3yjblY9DgBoqGwAltsY7Otd4VjP2yuL
h58k8jyB0j0Sbl7kjcytb8HTf0Y7ky1CCjPRCG+eqRUlKcb9eHQ7iPxVUvDl3+dq3x+/8AllEgb/
PmBB4WyLj8ZvZNmxtZcTULDmaJrJdxfN1Lvn44fz0Pxb6RX9zF5wNi8dbbdhAwRqszz3Vj1KkTu5
O+ZnKVDlEnzPFWUYjwV7T32XmgFGG00YnBwi0dRnqzZA93ZKalFXKFr5ZkmbIV98ZPfuk1aEcN+M
N1XHP5Qh7z+tb4iWEIAOfFNHEfqR/dWr/NzUJaItj3phICnJ+ljbp+sWmcjnEG52AkXvchtuwu0z
Eotu1IRISVk16IRpHyASKpK+7aJglLy67kIIA7ryJl/an6JSW14u3njNZO0TiPxZjg95pj5A5yjJ
xPyNrKZOImO1Z2Xde/tIQMy4G95eiKamxiIPUI0x3xLxqINRhsbW4Gp6dWcIn96T5Zru8jWPHrAA
jnpGq3e7ehIVxdDS3MbaMqWt3j68tqKoghlUOkhSajGBtXU2RdGfvdf4cu4mDfcQ6lvb0XWt+4+H
GSrc80VOIa8yb5R5wXVnszfmaHt7Veo5mHrYWXBCQesgoEH/KdFo/X1FpG5bc0T91zvnpq2Vzyb5
jXbsaeLNpR1r13V7V1CHXKxf38w+93ZQcyVldJG5yYbLVKJ5/JC921eosHI5e54bOjFZI/9l6hSN
RRmtaLAtV/q8O+qH/VebuQKjytvCMoT4SQAJzaReILOXXSyq/YRv2eER7dWnseHIWCXaf6/TEJAf
QY/5jJDC1nN06V6eMjqdzjxa2/Ea+J3PmffrFb9V6Kn1hEGh9f6ukkigTiI/VauWG7tB8zdbTVph
8svD0HXbvRcxkbIG4spUEgNTXjA+Kx9mwzscrjONHMab7dvoVHr7fYid3LrMDGcOpbCnb8Ezxf1W
zIuZI/xRAg+oF1pknBi0KyDIwjyfdNzKydQUWFzvcAwHmUMuurQiDOHIy5rJBbkPwvgzXQ0RkedX
w0OR2yHjFTrRJvJhhhTm63Ym81hE982LNv2veHIaos+TkX44UBhiZczvIr7acDVodahobSkw/rri
bGl26WN7vSmWcV5xwy5MXNnKrLneqYdSD5B+nnTjwvBsOQXz2Fqw57x+sCyj4bw1Uu2VzU+DXP6v
2l5HwOm+/Sy5hjqoId9mT0p7r9fYaAsSKmxe/PXREJxwt9e+mUWW3SXGAKFz3kEIkRtpHxKx/TMz
B1XFamdQlWU+/tWzoQqnQU3bi457szLoJeenLSGetKK/nBvqGQG4kAOF8NBtwY+rUwESG3SapQ3j
YZ+QW7AGGK/brIu6fmBb5gIo0BessNoJYFC7GGE5S8MPof6VnDff2sqAXMfRTRLI8p4nOaNldamb
C9VUcznNFVpSrCyNrByhgm8Rr3gHdGxE7OkzwYgU3XEattfGuJT+lNexkVJIHmKOeqJ3A6c4qQP7
lJNq9twvpFDnrzEb/7LvUKg9ygEVRuQDP5LxDbbH5EGHjLmYB3jTMu4CCJ37d13FkdLr2UoQelcR
QfYAY5mhZvgRrTgho8ybP+ygP8zWfPtaZMVJLWvfsYg4C4t8A2070XIOuK4sbsLQBLhmweTWYzld
bp7m1f2JsFy6UE1n5O9ED5T0pGupdfV8Xa1JYg5iB78dCFeZinAUXdVEsdFGCzY8tzkI84bHdgpH
JmzoS+nnRJbvnQMsrezKDjPHAMD+Dp8dQLtNhXgmYBAzogGCSmj1p4U9EqHUEUb1Bj8zVkjgWfg7
PFatpsvnNSVDkCr4vwo2nOIwpnLDrAgTh4ixoYt/46r0VPmls1/hnKvybZ/0/THkoi+D9sNGaN7l
h+Qau0dWBI0XEszodD2jU4z9pJkNXzy/u7iiZO+cCNREBI5B3JgNGft/7RP9YBySiNk/r/u35K7I
kWxd/jDfxrUcNzLqXlwCOLD7YkU4Z96/UNJay0IHnhYg3jSlHR2QIP66PKJd59fC4GJu63cgrH7l
/3PQff+bMSo24u5fpmB/J+CzwzIzpRoyeyyzbWLzs3PfndCO5Jgba2w/lQ9Zfuf/6GgiTPjp29WK
Jz8SKskt4mNcK5aD47l2wyuQIxudQ7pR9FjsRj2WIlkvVD1B3yLjqVTAdVCcZsInd2S51aS2loXa
WZDgh14MqdcS3H6df4JYU8GwNZDsq5e6OVs9SnxpdZQsHKKq3Lyh8/MN7tbnGzsY6N3CK511oYOM
OyrujW7kzYQLamoXZCJYyAdH1X74I2z6vrFIf4SgcgX8bPgJiojc8WlaaLm43zH0gewgiylTbro7
GaJBPoO475y063JzLcAyE4C2k7p2lm1yzAQjxMLkeoS2oWau1OuS0yijKQF2DY7Fx3idQsVriPa2
sfQ02ztaBX9r4tpZ1/BLUh6K3s4lSsTDPQ+XY7qTKRzbHNzNWR/dFWy3M1Fqlw5qaVzxJsQ6hHIP
Faucecvxw9QAX6qseKFsz70ugNJYzyvhIaiwXPJScMaEgozHozOS/43nTvFkGEmkrRyKEdW/zNs6
IVqmtcsdBOLdrc8Ib7sLphiaokJbs1T9RYYrNegNLp1F667loQEcqft1SMuBklrKPlwG0Pf2hXrd
fNooLbFIkKahIODe63RKGigMOFqewT1+cZdpNLEuTVXP/hN8ULP0NnK0Uzkc29WDAKtWCXEFB+Jw
sotV8i79HfUsavlGVElHCaNc6CDOdSAJO0AcAUOJUVg8IR1AW8pIrqGfuZX3aSHjAZQhHZE1h51/
ahTBSpuha2ecwGiYG7iMo9faSPY5YnHWP15IbDcQSw47JfL6truUQEmlq8u7hDqZFjIJ5NgQZLeB
aTzs6/53bjIWMRhiZZFaOwYp9+hlrz7VbTyduErWJxToDzGgAWXLBCRoKxk5hHw890p8Aco+jHKs
GUqM0nf4A8dMARdRg4PzoA3AbKyDTKJPQHr7YecELUSL6KVWh1KzoSm88lTKkCh1AP33OJOHbSvO
hOcxqljEuyoyLkzyKvBpBw5uFdws4//zO5qFEoQkZHe9xQyZhiC6VwqrestDRqkH9tadKCUeSsba
Q+Ywhbi0dMtXuY9ynEZ2wzLKmUJb+CcscFU6VDU41z0y/tOxY0ikcx6UCOD0Np7fKrp3wB8CdQQ+
fRGkj9ypPbT+PM6LZZxTJv973eeiV/SNznjy4kZ/qwCLiuSF+rptaLqbb7tISUdN4x66V7JrVWW0
bYRPou7NAYBz6vCRnNznYK2Wu2tSBZhfOQkcJzmE00aFDxFtuaYMa2DxqXebVRHOcAVZjgyeZJ3c
vgnoFuYFU1UP0Mpa8uQyt4fDT+KnGGVdX4w2j6xtokcsbllAdKxne7kSmQv7EQOorR1gQipva3Ln
5U3HT0kJvjfKjxEZs2OwSPOvMFSwl/sOUfecBMOIQo79LM2EgHGe59KjVgprsxyN1p5TtxhGNe4J
XMUlvmFbWn1Da5JmiKBE7VV+TZPir7SfTf9ABQYBPxe/II18tHD7+r1erUgjLhn/JyI39rl5z5xE
S5v86AvvjcCvZ4iuwVIsbWYg8gsvZkDUmGtVYUczO/oK/7j0Yitjq2FHAPtNZYAM26SCZ0UOKF0n
AjDPXhH/tAW3iskXO7SZKQOHs4igXBds7CydArxGUXXrwVKg+fNl4N20CuPTTAVn6eKDeTuJiUzx
wXJelfQJG3wyWMmysen/ETzoeK1K6JcvQ5HN0cgwbUZMFzXJnzIji1hlhOIPd2/l6Iv0XHPiiPXQ
jSBTxX+dRQOeJaTDmfqScAgzqjvvMKvmSvATSb/RkkmTk4EsPcMKLMbj++kaRJ1otimODKxpJk+n
OWVczhmddtfFHrZdY/y9CDTe7RfmayAJ2EVSQp3JsDF7Xl/NLsMIKuMPX61UaR2yylVhuoWfhffy
dqjt0dgvj32cQ58fCr+sA6c51LFa/2isiEEwwLZm9Orj3Oie9JAobr/HHdNdWFFuSiTP95CYFeKu
ceATCICBJ8DsxybrEyoAiN5H7sD9tDMnDK0chdLunEsVSTyQfbwmTZTZBLh4RZxfYmx0ClW9DI8f
OfrGkldk6hNU0c8l2kMiWR/AwL/anm5HcptX+DFgN+rpa9ia+BZ3znwNT7o6JzHvNrEWDAQv0VeB
V3c0lXnaJ1XYBaG9inJfFap5ZoGyBjBQvFYbzbrhDcH5eB8U9NE/Wxp2iB0sxVi6gfmCIDzNHH7n
sdiruLTCXhn3lO5hUkqt8i5i/l1f9KjYvK8bepypULwreKuocNyaSPzqJXYdkwqG49ToehynFWLG
UrFLVvBVTeMg1QMG8DQrlfHIEzyuEXtOaSEN7Tau0UcgRpnwalTH5JEbkqhBiZLGWiV4Kv5Wfa34
eXNvUZXVDnF+cyo3EbRTg/AuAReFX3SpJ5B6qkBBHy4z4AL5/M4Hn6BbDtjhpvM/OLPLR/CyFUPt
dWuVxk+f0S+MOlVWQUnwPhD7mWZa/ezvBmk63dQaUMwqwW6p8+kDwenmXKKW9XgSiKHkSnlSLXEr
rTGjLn2wNNo3plKOyMlHrwxbNEFKlb36BhV5U7ZUst0rQITgqM+SQujlyEkC29eW22nqEHZeUEDj
ixn8CqEUk1xNK4btJfZs2Vrm+LVzwQw9oxBOsywnkUF+Mr9yTlINrWKBBkhJUeV2rmZnrL/U6L/y
0JPxpfdq/YRDse6hakHIH0G+wABHSlW/yE53D47BivHoDQfrVr4uC0lR0W/4zHwpXXdMGNVwEjcN
FxRvI/2DwdGcR936lv1Q/io7pc9p6GBXZNOfm5LSVB1XLhLo5/uCYrEPg2dPveawqCJ7mnZfFTD8
9G+StYiZrf5YYwJpjnJ+pWc+nUnJM/wygTNIxC9S6YaPD/i3XeJ3MpIHyq1JaZ3uduO2VlPA1PC9
I/hL8r2y1Hp/fKKHhM6yKkWte+LEtyF1qusIuOFZH64Ze1ZpPlNoG3iSo/mb0fjtbm322tpSWauI
7V0i3B7Y9E060rfRLTNHIv1aKE2+04aGEcs/YoeZpcLbcIPV1pxtUFAiVSua5BFnuzwacUmsPSTe
/xQd5BQukBy611EL6BKuNPhqHQoZoPwLutbLX2d2wcWs5TRn9F0txH+fwJzqIBbl0cTOIVii75U1
dDvRtC+BshJ3h83qNljsrOAAUQ6Nq8Q1N09FRBFIASeQeuPMZwvw4x9+F2wixB2GxsCPvWgE50IQ
E9t3eVQCQCKCyREQ7HKDKD/IlS0pczDhu8T9KbW0Tx7N18MhV/33Rf0LAzPlUq0LZWm5NK+jw+S/
/mUtfyKdDdNuV8AJHGKFebVgWiXiiiEvrcMWDSuT5RK2Xn2oQ8a3Oh3d5VX3QqIYJh0wVpXnyxLJ
QgqrFoAmtdRl8Z4nCfgBVvGLfaWtNuwG2mBJbRzV66/9F5F/lDMHhJ2As2VkOtRWXPWgycNHsJWH
oRO23x5zKsDLFQ/TY0EvwX/YDJ+8X5sgLc5qkT1W4aFPNzACY4txVPpa/Pkhj0/iq+AmcvHtPqaS
S9LRwNXrS2oNNIeLG/ImmNrpqb/rZxSVI1xnDRe8NNQxcDIYAvTmidp2UoSgMTyiie/iufuy5vtV
7H77h3MnFU+gsQwv9CF0bFBBjTHaQ9Tw7MsTGx5WrcOs9gMvTv7qayk/gfNIfvgq4lK5j/KjzW3/
F9WKpZUmhyMaYjIOCkbe3XOHBodSCRBvinhVE3BbAZQhJBurA77cdcodhkKAZqPMz/SKRwB/Cao3
Si/uzOdsEb9Yb2XnH53E6Krqw0nxpGCHvNA4pMKgYiNlYZwfG2Jc9vGsldI9UK9hiUqx8NRN8yQB
XsyL2+Z3luZSFZ/FxzYEexLh/wKLD94+1jXDqsXu4Zfq8foiGKIcHWPWYCRq99c4PN0fD7pkt1DZ
bKeBxhsDwcRVxdIdUT4f2nneUi3wZ9ugOdR6yY90HueDx2sSxQ9UpkL38UqTAwgJte0kBxMzjXEq
Dz/nDp/+WP2Xx46xVXK8rXon8H0Cr8qb5XhoOxw8e6Q3v29HohvZgXyctiQXJuuEEv/ajeBigO1U
IgOdHq59YLqZ7EzZwfhODW+1m4MBv7eFXnNZEKnQQkap5pGiJGd7ijj/HcAcbip0U13h7J/xm3s3
72/djQuzp0aMZsEWs3IYQl2ThRWmKxJAQNrccJ0Xwkx/PCoGf/lxGYTG65ecnq/6lhXoN+YGh88a
ESvv4D95qv4RMk7sqdYnWTodkEBlyTbCd7LDzIRhP16Pb46mwpnvXnTYHl2mVHiN1ohRLSsk6evz
8Sdrw8oCyth1tgZPvw+dBiEsZ8vW5TcdM2b7EwZ4lXe4UUEkLJC1V5riyg2oJpHw/SU1Ir0FdS20
yhAAIhy5iRdjWsFvVwebVUQhVwWjghpDxpzdk6iTifmhxxL2UfvrbVPpHyFYRUVDPWAZcPGI21AJ
BTy5QXsxn38V51PHdS8tNG9f0Z41uwiHYJlZHPZEV6kdxogNl0pEczvYfgjQrnDOUAl60Ux7Xm1j
1peiudxW7UFHmhV/lWvmM7buoi168WCkgT9UdbL1kUSRhivT84jH6zQEeHVhJcsffLLe7x02YV4Y
Jz835V/CUjlGTd+8QcUQryH1Bu5+FqE5nzc89Nk1pZ2RlgV+nnceKHTGCdVjzGdtOJ+CyrwwT9hm
zlKF6aHv6lYctUAodOMnWCNbzTuomPhtdkKY5Ed5S7GpEXfn7tzHr/r6scjraG3jkDokEVbDt5bF
M2VC8PZ7gTVFdB2C2s4/FcT+Kt3mIRwJMyXWpBGSo38nCSa//j7MWgZy5wy/XuXcFtNRv2ghtWpY
/Fd1eXUP0BlOM7rwfa11N2UeOjuWBMY1713qcBr+qdDGzUCNFpVlNpoXxWJTD4O0bgCLdObtZ513
JyRqNFhtH0GbcZNWp1GyfAGI3YVJ6ua3evEM/tgG2MEMSVg3leLjUJgtdZ+WghOv0KaNSfCEm1TX
K6KKsBmjRJ/CFqT0nQ+xb7nZmtS4GmJ/S+EpjMafuIGFxjXzhkz+Efg8wIPbizKaJtW7WXZFJVq5
q5j2xO96tDhz5a8M3LQcVX05n+HZ75CjBeVV0bhlppu9UcVD+vPHwZCSEKatZm85xEFv+zHB7JLM
9fIS9iqazSTK9yzu/Ckefw8dzPzPZpI4pGTuFVJ6do3NdSOCddRA11DVXGLIV+JpKJquGZRgwz1W
sh5FSU/aF2K6yHNLmIYwC5BoOVRKGyLf8npcEx7ujfiCb2g8LRMfgAzPWu9jNAbN82oewVDbon47
IyEeaRnfg9m2+FQs1B+iIbwEv/kXqo7GW4Q5FRwD8ukLNQ3cRM0LIAXQWdPSNhNsR3r8gqYcz8fL
+jZnnGbGZHaug0v6OJSJndkagbciHXiLRs161IwW0BVLiwSse7zDbS/ye+fs1kB8YwCuJVgtMr2N
SMjkPKq55CAfQaKFMJOgGgdUBrKwY4zn/LaHL36ayW4Flg6eUQ9qHaNAzJfoxDh7hCSkrbYbh0qp
XBGHJ4me+sdGNJs8Mcr9IMceBm4I31MSO1whd7VqyMiMJ1gggCjUm7fLhS2iSIXbXEQQmWTq5blY
8LxHjpMp9w/VTmPWAc+QANKttU5Mn7YkILakkN9Ef1CgYVFQoCdQoqzKOUAooeWMZx/VxVaGUgDh
sNWVhw+4bFUx094l4Xz5EubqBCvr3LjR/xncw+79TkJCDPrQSJfkxpqHQw8+yK1R0tjKLFuZFiu/
5DkYKTKIWRnso+sKtmN8wB2gUiG6LBWnajsNgiMvCHpZV98f0MVmITogZWvTQzO0H8GtJd6/f0m0
f3tbrDxT3WS7hVk4iiCzjuih+ka9pHV8TfJVpopJRCaksJ0JagGdIsoLRnb67XgsYSbtBmkTzzVr
Per31FNU+YH7GJtSPL2ewdZrmhGq3DBRKcoqSTVMoqKBqEzfvvaGMJ3HDT6fkW8eMH/w7zDSK02K
pHt5amL4KZ7LpjHvgf+3PkLD5uOtVSxSo6b/QJ2VmSDeN6ozntVGZIPfubUdzj7rQIuSrruDOs3G
QjvUv/OPmxwC5PyY3hOXwkDO4CKVGiqqOFrP6KhiUr6+7Rsw8L5CHjzqhwQjMBGd//QqnyQmRslG
tc7E03iVsueHdDj8zhDw7HtebBoPfcU4SylCLnoNJt4R0LUnPUxZyxrSqSaiKQxCGhVXYBa95gbA
vC4KC+8VUr3woY/7ax5sLSXGocIZC0lNAJl3t5aOl/tgbQyd0lwRjQNZ6Yoa4m4cChTQpjw4qHsB
x85xwiRyz24ZrpyvsVwfbb26ZzDXpz5z2ohMtkkXVjZsQymZUjXcwuVzLI5rZDDjbwtvHHAJTked
hlZvxdEbgN3+GrqDWPs9hBwxrdhDKIEsqJPWxnfxxbiAW/11tlWk4wJX6olTcJPnLrIPo93lgb11
8NDjPAfWJULlCMzAZFQVm2OZUT5QL2QMNfn45UPHnmP55tSdypZ+3yFSuXXdZa4r0x+9Sxkrlefs
kGhEtCXfNgVwoHaNSIxD6BDncW/UQXOSzyvcrnyOrvpx8z2xnYUpwUynYYE6A0AsQbQ6D0/1KFH9
/mugZEmY+jE+SahRbqQhWvuV6GZvA5z0h8EJnykm2HrhqS0tc7zlxL0zwDwH98/zA2i8VzfU9yYC
B403G+znFbfn5FCBl0Wy0+mRxmXJ2rcU4xy/VZ6r5w9rDoyUdVjGdFfO4J3NOH3rpWkfWFjh7qCo
JJiGtXh/ZLyJQFxzF5Bll9kFvWOVZlDDUStRwYfD8Y3EUpqZ15SyBOEO4qVR+zpjabxHNESscqDq
RfJk0qo3u43tqeNCMdFimqAPAkYOM2LUZ5BLDP0tGZg4XI6bivlSoejhkLMqkDkiag/n4u+Iv7G9
oR9dOguxooOq3tF/qZm7aSOmEkOlfOlmOfe7Xr0MmV1pWy+unyxmVQAfQN366n5AzcxuMy/Oiet4
PyqsghJRW4UTma8HTLthVDLzM6Y11A56Vng331J4Nd9vRPjMdNCNK7v6W7fLNrRFG9AxnEi7H5S6
fx7B/4ycJzD+h7t2AER8YmTkIMm30cF5v+OSMlnvCxWwC0PV6HIhFiesnEKJK47jZ+Cdr+QcoPCv
CW8+V2ClvpWLYmmAbszL7KfeL+g2XFUWuanz+8zWS74wprWaNP2lQTbqZe3zsBu+TgLBf3+opn69
lUdayZRSB6CaKkSHWuthvtNQV3xRzkji7ukalX2zZ6d2MosZr5jtI67euiI+chEEBgozxGOSz5zi
LGjVg1u879ndl/OCjge7QwpeoyJuCChZyIO+uJmLlEiUykJSeW5FmwV9+u92aArrf/B2xfXoj03N
C1Dz0e6Fw9zTip0yL3hkSCfqdYx565OeEJ6d5Uj5KlmY4E7tzcVn61bW4LFXOPcsLcVjoCVvCapu
Sw6i18hW82r45oyVaaWZSeNOX6ON/Vz+f2CMaFnIkUXwk2Z0pbz4YKcVIzUOK0tdCB/GRohq28vW
/cYF1pudE6EqtlQYtpcH+R0srzts2jAj131JUyFmal3tALgxhit5Kx/qv0sMn4vsCIVWhPUhjZtw
GXzd3U2e6zmDHsORt1bhWQooMtlNz8OZMLFQ+l7eYoL02uy5PzZcA83JNujx2E15zOm3nRzhs0AC
hgnMylDuisWpaNAPuMHpDpNHfiN/okA0gl4KqE9Lk8lL9PKyR7r+6QSUxIh2l5+LUvwnlOZCDoRH
xrehx8KwzG0hLiznCwB1UnZGwLOoc+5csFAPf5XJz4dnZdpE5tHT8bhb3gR44gK79fHcT6o9SHZm
2j8EeaXRjM4KyPJjC2pEpuGiuY+jumaVSiV+15NUYYUSzuHUJnyp6tDf+80npwlFtxLMNuY8jAa9
v08Rq1o46OfnGGEVS55aQUNa54EJUYLwHDf+ayV8TuuQx6cp+YAqP4KtdnzXK39UiZiLQMcQMOhU
uYv0tkQqczkIPJQk3x0srGcPOJgQZleR1/6h0AKUIdxrxENOg2wcjiZ7Lo/SzeGQ/UAPtdlWnnv6
fZJ4FkG4EEEKIJP+EE8tALANudULxCc2Yd4MLQ/Fhhq9L0ok0gP4bEFpRHcvnJyefwbmRC8O4p5X
11b279cVskAMtVbxk/gojtKXAO8PgOVneYtpa7PAkATPuGiUxXlodQPOgWHTImoAyoioXwCGEuUE
N3Om8vBo9KQ8BdW+Q9lbTlNHI7e5W6lXeVg17Y5Wzwcq1cI/t+nIxxsdda9A1IVEK+GOSwcBVoJU
u/1WOG8cknwqo/DyT2yOU9qHRswxAuJQVEAChK3xg9ydhCynT3QBgyBgJtcB2s9857UVSY3Dqu4k
g5OuUQHOQ0OBJMRDYtr5eLNwNPKvAPfhZeF/sBW2acsASTiodlITbsrAHbwUkS+AGpydMt/NXAos
u84YwTv6oxfR5PsAbXoaGp50bVBM69LTugAKbai/mk9kS9MxIdCf01ywo6ymPeERnxEYEk3nmJTF
R2SjU04v2EkFPpPWdsFR8MpkWPsEZEHmlor/KGxL5kzO8NbqZOgst3C0J7f9L17Dq40bjc8/25F3
4M2tN0zQDKAcURAUUcBzpOsbmLpvv48CV4hFjheJhygNLBVTDYputks5funK+CIOrspiiYDZTGXQ
Ux/wcbRvsjy+qbtF+hHRmcrppa72JEDjguPmMoqj6HWNZPqGPJHOt8cE3k7tVUKnVQ1cpTZJPOpV
4BTEsaDaSxDU9cWJl11Na4PZE9pa9mQeh9g3KBowfN0u6GQfgaXTiya9HTONNcghSh202R87pAwV
OcmLyU+TtK9qGoxrig8zl26X2PAizGWUYO2Q6lI/7Yon3EzbUL78AzsVLyc6QTl0iAF0cpDTaY69
flaxHXJkdxaUulyRxd/Wbmrgm9eOwZD+SIYEC9hmHqpw6+7R1QRDDu0neFxjyLbFQh0gDw6zDxjc
/2Thh2UPuGdUxGPzm8dUwWl/g1v7ZGRQsH50+EibpfDV8QiqNY9ohBAYyoFa7eCllFc8POPlGu7n
vGBrYAmMtgJoJnWNfi44SMFwZ1KkGJcTEchZTMQsKpU00xomip1ACdVO24bsB3hJzIrxfMG/TsOk
1lnxNJhtJrPgO92i6tMluA2Q3ybb6/QKO68RlVU0xPkLJfvbeQGVvKFQHOyvwQyk53auGS9JbVD7
wRG56HHYCzgfq2dsrEYUdsgyyTVaOkLgKhYGMrfZmYpiX6MB8uuQTtCYOwJgu/vCxlh+6XJX2WLO
7kloPd5VcafVwXOlSjVD4Xueg+4x/xzfd8Ks8PcjskZ7UhuxTwNQxNk1D0Hy8p1XZzv5E1Y7MMlc
qkO/qUVwlLPjeVvFA/9NgZYi4nxPBLbfruTltBkhDrIepicDHPrl3kfmD22x3TlG3N1ftuJ3CM+L
tflzSIpdgBziGGt064t6nERKH8rUc3DyjP/Hpio0Y9hr5lbGF+czFTg2LhNBdAjr05XjHozOg9zc
HH3V91MZgtA5QYraMT5x3mtBrMLokNHdtHClgub+MuMFArCboJoKG0IvnQayNBYm+2f1klH7mF2N
tdwfxsMukOJrqVDkMTv9f1GH7B1+0tG7lQoE3eLVtTq3pCTt3SpQqk2kplSW2AZQcHa1hTc/q/bm
KwfdnjOwtL+OHTKXVMSVg+/o0BgO2oL2IGn7G9r7cFyvJtSWawLIACwmhhjUg6G4HWfhRChImlrJ
KP4itKUmDcBAg/RTLsnJayRs1NekZ+Tf1bTNIGrvqgnGPlB2zFyt7gZLNPABTS3Yziqs4vz7H7C/
g3aLjqvZUMrIMU7Bv1wMIcaV3AZVqjGQASpEaGm9oJVp3SRLF9mhhkaVCAOMwaflIiQur7XXR6ih
GHpmG17jW+2jqeczcDBw3leX75jjiu01utwLrQSZs4SGg3xfdav/e7t5o9wL7DdQeBzw9EnwbJTI
IFwWLn5HroBxNHZmjYUbW8et14hjJjU2cydgug0+wtgsXhFNdzBFvYt439ump9NDbrqfBuluWwL+
d4gAuRvOf7yp3COt3cAlq24pIM4PBscYYLxh9wY8tDJhuQ3ZZoLjyPGNpyXoU6B1gcFwf0ymPd+1
ZfP9a7ru3MeysCIshs4hpUQlj6Aa2/S4SNScwsU3l9qExf9s0InH5AR3PZtr+VXI1c/LdGqxRHoD
kktpaQU+aXnA+0hTOyee+lStsAY6bt8wcC/v08TjTxAuhjc7Jqx2hggTxIaBEvKV+aIZcqi7Sh2l
MxKxWDgnAcgqj6b4gwbAI3NXEhLW03efwycHhU0NOODx0AmZrBcfLyCkM+zViJMHluOM9McrCdbB
PbCLFtaDF4Gc7mzq889sBlzMXmSlkZNISLdeRBjcEfbGtv0zcAKIpeKu0RlaRJKxqpeuW8G/gR5f
k4/lrM7zAFLEIo7EhqhDyodIAaUzIFJuTda8jicWI3UOjnBZfyciUw+mG0sz8yFBwPRQXH0pDT94
RVsDhPfX0xD+elBIhz9Tvf4TswoK9SH4jGirDEgWP1qSPwhTLinE+eusy19asE+cXOppg+Q/i6iT
Sg7Q0m4xV5uCgDpmJWWdfzfKjV9WtRt5+nUfYT3jmhuJtQjmrGkRYzCc2ZiWUsYoRGoku5SrI7qg
dkjadbV6jTk/rQYpuHBWV0R4PehZYsNlXhoKdOiN7gW0rcuHKL033pHhRSYXq55CxlSJd8/6n10j
MEfq4TJeybAr1977ECBOadG3/w2ikLMm31/yZ4opXlqhhIsWSUYzo+T6269w54pPp/L0MqU1cucs
ZrmQjLIEHtXgY3zxi4gYvVCrYxrrpLtGO2m3gToZhWl3bFfu+4HqnFWsf8F7j+v1HuTYisGWJ+8V
4R57/fv8kzeqUEbSFkhn8ixcgw7fF46b5qwBREmXM9GSoHPwVTJwZeVUIBxTzyWWtXdhbiOcPMGG
xDhUwImeW4vnQl/3+iRBZUC8DQLddozomHm8sBpr5uL6+Fv8zktbmrB/WdxQommfr0nuSolK//WT
0ZP4F+wmC19ZlVHSAK9Q054h0XPXqouWX2y+Yt6DCvm2PXf06hEtJIfpzfMXGN7xzJvuIt9+c6qQ
rC1uTtk2C5DIxkn6qB0Orn9MwwOquInqzUVzsnDwiEMOPRaVilgqpj0H8B8xTjApzyFOhfafIZ/S
EZ5OMZaoPW2e6MrnYetDMdC/5oKTbLIR0vSd5T8Jrw84o9aV1efAMyRH46INS1z+W370PtY2TXTN
d4j7mFjCYpRpExCF50DxMlFwZDJpELlG8sDWwUdgTiZxzTG9mDXS953JEdO/cyuDInPW3oTBFsY9
X//mDBGTr0BJ80VUhPstuuWBHKsQoFE6u/yezeiHLKJjoF/n/d2oLMr02lUjHztDWi8H48aIhT4x
bEe9rABHXtTqup5ZDKZQ5QABJjwKTuDThcD9c6PdQhlx2jsRyWWZHertbI7PXC98CnpYDcRGiyIx
dEPs4j9r6FbVapBx51IPI1K75Je8lmH1BSL7OdnQeJpEkYgIOLLjbFzVtQ9xuXxQaKRfIpRdoSYy
yQhEYOgHeyMnfVvfdxuyLm0VU/ZeT22KZbiomT7glBlp0L2bndJLTbJlZv1E9AGq/oTGiwe83Fz1
r52LBWImGt5dWsQHNlZjZA+QWigqiUiTlJI56ag7THT3fCGiH2+XYpkNTeqaQ1CHYNrUZLsi+G4x
Z6UE65c7UcExTjrCKKHGxvh0tXNUApMDNlgeX1CPvIhB46IR9nW23aOeC1vndbm/zFbRVubYEBlS
vp37RuxOjSeTLr9G156Z67TaYE/6ygbQoV6wwWSfLrpHFSQzbVSnLIn+DUcjCMPQdiyQhVNaYHYf
dS12OcilJpqgMrlmfgyReJK1syA4pHhoiJeaOEVPi0cGq7FWPEAoYAJvMlEdXcYtc3DpBygbVQm0
cQTp159kHf6Gl5alEska9N0yee79WBSqyY7cPlU4vWWQGYsFl72UTgG5IEnZ35x+hQrDQpbFD3Mc
T9jl+6J3Mb25wX+0CFeu1xyudyDdBHdLdipy+R97d2GpE1uqCTTq6RO5GZ10kn56ugTAOT39v8jG
dadjLIH//0405o1WmSkMtzZduGHOEIFe58+0vFAGme3PdFgBux5OnNCzw7ZPk+zJfW7qtMYMsZs7
zUM1cmbCk9m0XEd8yKublPq77SpS5fIH88Z2hRJeg+JFsVsNvKAJIfHfIBWwrBqVwaDsbJ+R23es
wdzg0ltlgUZVQsv1X0Fc0FM5t7VPNh7I/xR+VzwNXRRtTiKoBEmy2E2wlm8P4CglaLATkqNh1ZQB
4pLWatKX0COkRRIOc1bNt8p6YucwHG7OG9rTx0y1MiOG0N3q5wrIalIlTU4pLmT+k95F9Dc0gJ1a
+GQSbi12dNH1WwEdiUUAUNjdevgvN30cRSjh6YV89L2fFYV5O5sd1q54pQdV1BGAwa111dNI0IKB
9908IYKR1l9ZxjXzROihFhfyHceC/pv6I5ZfmRvOWhSAMxF/BQUTH2O2359qYz6zO7vnqjIgdgFx
gUIqFrDKsMLa1+BFAyyLiGIjTav2hRaLVF8xnyh1qMzR5zli+P02fpSuBbvm5csb8Zcd5EpHE5UA
4Hkezy0gbnmUUnAgnj0HMFVkHk7fwXm/ajJgZ70qPOAYR11hzMO4Px7P/Pw9zRj/jPCW5FKhH0Jc
2DICT6cB3TEqFlgeMJnKD6ds8+C8zJHocmnr8FimdrXxc0eN1NFh3fuf9Hoeq33AA4Y5rcQl2KnU
J2RqOmxfeTzcysO3GihJHf5tDM89G/zMpLCJ9P8Bab2A9WtR455/cyBTJV36q6Hd8vfE9vs0OXL8
Se5x3JPVhuoXnsX8SNMSW3I8SAjKTVCeaRkSl/KJX9C74kTNcctV7CBEWdwvJmPGU8oSGKuKLPqJ
bW+lVSe8QiTjzugwSoJ9pcpE3lmu1kQX94oTU3LrMmwQE8GuqtY3I/y1+fuAPLcMOxjbTvI6wKWr
MC+KWtKe4eIjQ2CPsF5Q3bwLeKpZroSQkYOvoL0estR5iFIxoKPoFPd1H9T9v30IGjjINEwYC2Rb
L5A0HlaGZXYOwNITTq5jlSBzV4ZE3k+Alc/ioQzYddhMrjEdad4qqE+gF5tm4ZtRH3ypGwHrRrC7
o00cs6LJl/Hv5qxrVCq4WaZEPHYVaTSqApsOn1Sz+2M/dJB2w3X9OkXTQQ534X6ltjuguUHucJWQ
J+319LlxP8i4ph0akEPvu6WHJ9mKW27FPbCUyUOGWMG46qlzaLahWTMQZqBIjNlHPg93OkT0bHki
9g3126X5dbFj6F8KlvdwhOC6/9//RpRm4OcvO7YotEmaHuhC25zls6p6AW7ZdqGiMvEJcjpedqJl
cohF6RDggjl83t/SNhie3b4/BOVlsIYJb1RVVe+9F4RtVQcZ3DZzGIRJl0gCXfU5zI3U/IfdSEiy
WgYFCY6h7/eY9dk9LO5Ws2vuAIukt0fyjR2Gr5jMQbhkXyFgjiWwwxJfUWRNQqDtXCCa4Q98J2VS
G7/4oJDgbpa+PrKAql/MK1JbuepP5Td4z0zlj/ctbP/QJ3R/IoPvv34DI3C9I2DF8wF61VVKxkb+
q6jH71KtubltUmNVP8/OKUDyPBWGJU45qb+s1tXylM2hG/UOY5CKb+igdExq68Ck8lXkoHDmlNNI
Cid/tobjPqvfb1rFdyXAmw6wjIZIkP+45FCCQ9p6Hf0lWanQYP1aF4jhxw3Bxwpcbt3ZuhBcFtUt
5DujWHf113phFvyFyDB4/VTKEYFA24w8f+Op028ZxynwIXRgYcB+gKUqE2RGLv+TEUmh7R5L+pX7
W9nbNpwPUQ7oOa6DXiO5BAkoPNAzUW5by1fNTeSpIbwrbAcaS54O75X2C73xB719SNyb/NVTD3TA
sovIIvdIv3xUDS4+1Fi0uPMTcJZQSH5BhJ0+mIlvEJ6KHGQgsX2jgmcbcqW1nts6NRfDw4Epzdje
SzyyPsvnKsaVVNLYoyzIFNlZUPZ8X7iDUW3uDDVRXXB3n+VWJtflfElQk3n/PMwnYH0G5xZbKfaD
G80T4x32Tt4VMvRlqWpP3sO4nM59A4j5Ee7+hqKmSfY55sAIl94JOEOW3+UaQboxtdKLKLrLk7Mx
r1j9XKRPfAttW8ZMzSJdYnmfM6IUSSwd1iGaM1AH3LJ0ThZmvpEz+QODQBzs9FO5n1gX44hyGiXB
ThH0u8/GicbWykPkv0DvBFyKq67qk0/pwJtJT/IvBKw3Lt9K2AhkJv74i3ZGatF6abeY1c0AYJfz
Oi09DRcIC0VMzrQyHwr/RSWhhlou2P4BdYTIQ7PQgxdJ7zXIrAss34GydNLmFZ5sUFd5UIFp2OPu
chvubPL7rhr9PZNmnndE6O4pc9q+YlOOSPNSy6JhYPkBxYhSm5J3kNsutKrVr+K/KzojH/4jxRQj
xfunhYRgeTNazRm82nhwfD+QqsySq8G8u71bvRd3wFZ/FJuvEuVfvEGRnd/A5GJQx7Ld+Pw/P9bO
f0aFYR7DzkpLHPu75xTyKcUdXVtWYHjqLYyRnASeBOyCs6EaAzNQ8JZ2/G6DrZwaBmw9lMlYyrlU
u9Gm6IYlhgbHbpENmBeLY4zFdu8EjZmBsKy46ZtN37aXfDDn6oYGNMf396bTbPLAcn1cwXuss79X
oUZOZ0dt2wa6R8cfY7N88dE87iRHAG7E2CIYo5ULyPM7gb59QD3sFKBvJX2xHRGWyGDKVmd6ihNK
D/ZvwpmvtgQgqS6OoEmPmThN5P/80mUBrdAATrlWmrxQj59sLBizRiDUzcFDHp+PIemrnkYtDQRG
pKBDXKjQfSxtaaU0xVc0ISWxUF+tXlrXADG5di8zT8x+QC9i1uF4HBG07Lf9KBuHwxbLDgl7AQz1
xAYndJ1BKlUJfnY3XVKEqnYYhltlU+Kk4yRxn72PhVZsjspMuPxW/gVxjT3IQYWR1aZbPxmDdPUS
HKhUp3yntuX4RtEjnCtMLOIETsTJbasgx8VOJD6K5bG4MrI9REM8u6NWquRPVEkxB5Z3QniIXWQa
MxF3ThDeW4C2w4SN4Wm3/78ko5a6D/KdOT3RtvhYLGL9En9ZubExBp0UiGKryYaAdXZT6nejhVKC
GNAowQOG9nez/FzwDYPRCgZjwmF88awLitxV1cgGQzkbkScBCuLVmDXkmNn0Tefe7IpW0z4ZtVGu
+Ucc0sruj6IzxEmU0Q+lesrfVAoA2pdMKKKdSdJii6xmbWqhq9VEoXMQFySxd6gNAgIJ9Ch+Gpyf
WWt5v3TEmET8bPyeVRSbD5BZmviKGmmUcqhtHxXP5KbY/r1xFPf8o4fDHsil59QT89Hf2GCkCghr
g+DcxzoUhw53Y1Oam/LlTEh1CVfvVsj4t5zQT605NUmbVKBoQE6f7Bk8Twuoq5vA9cGJ2HuoDPZt
NupJ0BMX3voVYuqaSklgguIDD749g6QjDIbt43U6VG+12BrpZY5A0EC+QohpV3tL8B7PrWVLAg57
cIIz8zUsX9NaAWKEO8fx7HoLTG1MxJ2gpFkRtzVCqs/pVGmlndbDq9xPtfVTtbqs2HaztMe9NPeB
BEn2bSBGUX3upd5flbYuFKrQG4Lsa39Ea21tft1iK99NTdBbuRdtbDqoGTIiTCyyYN3kGMaVYNM7
Nxzo40+TvI6DKathm5rINhL4d7zCc9Q+vNg5u6fzrWJ5vT006LY9qwxfh3+Z+hhTJ/cgMcevx/NF
O1t86bYmXRrr2lWM2zbY2IAsDygUrSSjXp58UYzQBkZ+jx2bJ1n9RMpwNQvBeB68DyDJuQuegvkD
B3p9t4Ad4QSmUuL5Be7b4kWcePFOBA58oz2HNOE5tIfbVTntv4M0/MI10Nh43lKp6vClPDx1jsOw
SpwUIU3cL4IQAkJSfHLpKEbZzj8/8s1QndFlhC0TfxELZMYm8PdguBaoWdM/7M6OUFIT9nrQSoXP
wgMxhhYRuCPvVKzCJhDpRc90aDn8uC3ZDFrGsCrDZWjQaLCJPie7ZIi8EB+7Jd7VtJpN4k1c97lr
nIrlXJzQKCNEZ0uNEk6UbtyXqbNeQ9K97VEg5S3DS3+icqz9TyDC6CWhwZiy2GZnrw+/BmraoUXk
mWEsIrvX4hkSz6+98zFDR7A2IhBy1gBAMnRqe+uh4IULuA74wIuc23pK51DIL45fNnnEYai8myMk
JsbDhcd2V/g/yT8ROMsSiShkleUBZxfhZMjibZ98rycrf0Pt2E8rnmTGjFQHd2qD+NYrF60W2qWo
J7cyQsphHIPGoqCgo+EWaynscHki6JcjKKaLxZdU5rBopdmO1WuM+pn1oH17RvN5zanAdGGXii+/
8GKuO4Q3IlCKRsWL65Q60TpwjIzE5itmDvveGhh0K0SbAo+mlEsWuVIxMt1wJPUcrnRKET6Q7IMk
ceoR4v9hIV1o/HHZaeLCkFMavhoCVd4c8y5+xuQmeG+uNiq09HDIx+72mrmcvg3iEq50HAoZczZA
aAFMKUR5yvLfsHcjRh9OF8DzO1PS4dcw8u//UlOdielzPNeWGt37ke9t282wbAkGJqDOnjYE3TSq
omNKlsYhimvFXPZjNjJxr5MGL7LruS4HjsqKwzI2RWwQXB6DPKEf4YEpk+sDQ4og9Q1mQAj6Cbm3
jmOp/64hwQOyvgeCzHgOka5BP1V6vzvsX+LJpg4nYBfvjOiXD2eCzMe5+Ce+uZx2tg/BdNMZC6T/
y/Zgt13d20Ut+yklT3iHPe13ktcVqaOsywSD4tGnE7x3VuyXr85OPV76/WTsQsNcmfIBo1aphMXL
m6fOlVeKWfH1h9f0t9PlfQBIEFIlaJFE30VgmDVsPSljt4OW9FGdXhXq9maunr8jR/esqBkvw9y1
UCbfOPyO1N1wMM3O2bIStGq9FNuddB9DRAYYcLWa5M7CKHdqOetmsEYczI1K9neksLnhUqicRC6G
q07Zfi/NlMF8hYo8Ogr7SNNqQZQgmcP/XaHsP0u9PHRWU8bWHaWhQsgJeZUDPcx7e0OAA4IKoz5W
ODwqfkvMg1Iuk/fNf9Ua5VNB1tEnN1hO9h49wvlG3OySsvR8+iSG+tyWCDnVcQJvJ6fMX3+s9cK5
sWM0Jfri8+jxzlwzxhpX/ciw7X4khzHA84ZEIaPUC7B4iYHipZFONp956USltN8v8/Y6TZql4Cjm
dJ13z/rG4oIkztBM4aa2UfA4lZbUrczgCOS3yub+v0T79B3YbHq5VLOkcOgZyhv1baubiAXtOdr/
ODQbU4s8Fx5ZFpi77pzQdoBjz4aNh2SkMTUr1SCRmSCBV9Bn5kf2j2fconlPqGrpwi3XhM/AZ4Zi
SVWUBI9BbpRzy+DcCxrlfiJvRecTDF1FvFpSF/74XKgXFAS2j/gYngcTzH+g+cXs1RB/uBsc0Xpk
dhWLqNlzU038VWOPpWekFFZGyU8qvFTth8ToURLakBE1DS8CcMsJTevfA7odsacQ0nLGKTqkFuA5
ibdAWfJngh09P71ijPExWPfj2v4GTC96zMeNeYT88n95QcxggGns/LcpAz7JSqRwRNOZigA5iY6W
Mfi/TaitLFJJRO/VAS405c6JzdKP3zSq1R5HyIKOZEWXahWv4COJmx5+UXzggI/P2Tv5FUCy7szF
c82MbPPILEPvGfhTbRWMQQf7oyleBDS8c3ewaYBFl/FrCjvMAhfrm8e8ZiH85Vkv+CgC680rDKUQ
16ktu0n/mRTCchoD267BfTOUsTuVFFLTVbRUN/t7u1sRymUe5w6k+ErPrmtciIaqU006IoUfDbli
SQtLjL/WFuUUNGBQfeH5JGg8iAGrGVsxZyY8Ml1mst399pD1DZPfV15Bi+tEiqzYsPGjAZj+HLJx
InuImNOxbFR1up0u5fyIhAZz4MTgOWAg9+yVTjOewSgrI32HHK5IAldAM954b7ztpap3qB9gHSWD
tkKBeNEu5ju2N5e9n/VfN1zlHNmG9gGnyjOMRqubJSSvVX+BPQw1DsDaTbBhhGnp1RGvw4FR6Q9S
Bi5htldtmj/i6GwCjreHyKNQm9e2SenxRa/8KfNpZhK/Ttsrz832nU7p/oXaRtAs8kz93TGAk/xH
BX3DnAmIcewNCPuUrCbjy738B0Yf7igKR3ILf1P2DvtYFuVLec5PnrbmY4yJ9Gv9vTZT3SguFlOB
+YCQ8jaNSYUrKuoiWj6B+WUkXmxKKHagJewCiJbMbeu6Y1Ib+QDMoASKVM3WHw9nHxB6ibCcbODU
qwJO3bZ24arGRgTcnKIodQq+yiDQb4cDfKHqZCIv/Yn4eRk4hh0y4tlTpAsUuulfKvhHp0U5N7qy
h3b7IhWUWOwmegEOgcOx6DgjYdttZUjXkrvTc0gu/teOvzzjQ0GiEIYkEOL4LcD0/q5HblAqo69J
0+ef1RvWNDiCjmSaHyia7bH6J8JDN/hw7pwIBin8Dr9l/ztbMNc9TV5irSzfDCmv/eoauYq9Mnmk
TDe/TQL/xumTvFugglgbmjAmGAtYGAKQ2ZnSi+mBEiZSc1AdPplCFwrrSAsdlj7grjt8QH/p+Mhh
a2m/4RqfhadpkkG0r7Y2R4VV6KQMDVNjW28GVX3qhaYuUQPCKQUuw002L1fysYnO12P2gbV5rLvH
cECIYaQ/KloDA01DhWj8ruegEQCJdFTX5MDdoDopFJnGCcV6GM02RVOzHm/bXynaH3VGFLgK9jUy
d6TXg9sY11vMyTI75yg5XBQF7jZnWC9zL8gcHEtmo7EsPYWFLODz91g11oPPUe8WXUyc3lxkY5Hm
SceO2ZXlu5ZXRs9AQJSTM7oLb9bkvHXE8WUKhk0kV8NSIAkrSUlXvHIi0Mi0b1BMuM/MRw3r9MEF
myiFQGrDhyUS26xwF4fP28SL6OGjmcuEQBR9+w4XGgsFeboMKOjr6lHHjUhkXnypYHRMUSdV3RoT
MKA5QOBp7sQl4LcgxZcw3JEmwr9dr7T3MT769uV0N/28/cLr50XDB3Q9AYuot09GhFXGjOV0Jy9i
Glhw/S4jCTcByKhhlpmKW+tqch/yejMlDmwKANBwkqRaRZsP4Eyf71I9i8sgVC1HxwggWeJopxau
c+394bcblXDKOqGC93WrWIv90ZISjSIASlgYOjf8MI46HrLkebbLcVhuWGI6RHPtH9sJD+lVYetp
WJ5HDfuycPxRu49eYFZ3nyyoXYnWZqETaI805ljXCy7ieeX7HXvO1mjYAokohuYiiigU4CGkP+G3
jxy6UisoXoKlCdIkXPFC8gF14WJixD0CemNfhY01LGLByraooQ6m3gHNUR9mPPPBDc//Njs9Tnru
Sdx0E3AJKD+GX2J9rqsSFtEVuUoRkrbbyadVfWHaBjDRr0MC6as0NyIPEf5kRk/+fYXDzm/vAcLF
8jDdf0CayO/QEOKWPWx4WnvirdouUEYBBo87TxpKe2RMIcQ184fgpTR1lC+EZWnp390tTbbB1AxM
MmB9koDdROSQst6XX5U4sckr8ZfTKRNo9dOW/h2iYyl/+H6DD+L+6E6DMkOP75i5ZFm7wcPRlazX
mcq7JfasTimBlPZA2Xyiyi7SkH2hKfOU/w5IwOIcSGLm8BfAHaNuP5p/2ngC7JTPvnt+4tZ61YHr
FlxHJtKBL2FmxBg5EGAZYjGsNg43lspOxkDX994FB8b9SOlnFgoooQYgkIum6Iy8eN7knIZx1ymj
95qyACZSi+Xn5n6XKtFWMBjBGjUacNZeoBpxXOXlhT+5HefllsgVYLrhTtt76exdfWXKWmfCjaD1
fK43EOaJ2dRhX78X299Ekl/qNeTGvr3EszASOpY+Fly1Z98AuL+/pcsahdLYbAh7QGWjHgCpgLTB
eCWaTS+JHhP1t5PAaPCrou1gQcQtDUudp0eaA1JtWDE4uK4NSTlXCzySJZzAaXcxQnXYcaER2C9x
DZx4rKdlC3Y96N20srm9RhgRFzkIzxDak2zIQhYFw1nVIBItek4YIkEry0IIEVtJrdOq/1bTyikG
SsMXfWurpUvQKPbj81s7oQmOAaMFIGKOAHtIIjeIOpxYUi2uJ7cSVg3bYj74cvigPYytQZmm2kNn
qBm2YI3SKasNRMxVfhq8XqkdDnG9OosYl8AoW31EkLoWePCfDZJrID8YEsafuh2sXzBud6NkMBrZ
G8FVl3cu2bXT8pz0iteThmlNjj81MWGzhgitv+6/18Mk5mDHCyxv7nun1tdITrpSJVOBd2TfJQQM
gE9HbQhX1VSME6bzuvYOEPx2p2odwZ3/LRr5DleGYLllEMqxNnJnOqFQoHDnO4BIvEuDWqkr734/
dWnAHPEp2r+LkDNtSCGP4g5hLcmzWWpoMjhmALQl+/TIY0cEZtUT39NxPZFZ/j/QM0u+u8HTJ2aq
h8aK/HBzc0m1KWSLJnJa064cCOyPXPZuKh3nqfTSFixuegoxYZZsNsUS8mGca1206kDyYquSDWZ8
ljkOjpDqsi8TL9eBebz5juwvOvOSIebc8bdA4pUvjKxQ9VB7tlvaA9AVK4dJpuZfxu6hq083eXy/
qrGaUnFwXej7BBp3/g46v9BIC6AG2AtrmckpV6c0GKZRzGw2P0BJHe5ot16ilm2OaoAes9gIv+t+
ggxRlUvc1sWsjlr5bGREeDrMdIUi7kQg6raoIMGDE4MjUvKmtHA6FukTBXPubr2HM8zaatn7XKCz
c0+9/fmz3/VglTWvTQp1hvbqgdRATjiDkEKgeoWvvaYaSP3q+BKwKZYPq4nePXbmXDU1RBGIy/yW
qCLw2Y8TvwJ0cTrxi41d/49vQEhA7wz02j7nX/Q8C4zbKaBHlSG+QqIsrDjRSkiTvTbNF7aWO6VM
8cv/tdAdpfFpTvUQj8J9azvnL0ACLmc/QYfzk2UPNEJNRmuq98epHokfplN/TeyssFqAEePnsvLZ
NwHYuEF+eNRxx62jeVUPHI0moR7x5VOcPXgoiCSrLEckttjIaaZLX8CjLmNNhYMXq2BF6vMtBMbU
3rehD+foqm7hFCFNkyVWKqTt8MfFOqXz9gOS5Pp0cZmo9ZBFThjOhlEkVuLBWawgj56f0LVNtc3l
59vdfI6/Kg3JmeZ+iqlEx1gleL3w+y7IatsAk6/UNy1sefzdIrQqU0VehYRPAyWQjaQ/TN4rM/7b
v/FfmLe1gVWttDdxJN4yFxHOPy8ExI8n4mPq3LQS9pUYBL8wCptn+TOk/2aYBIlqf7f8IOaPh6HH
xyeD+4VUXG03i3okLS3DuiuaJag+bRWtk6hDt1K2csYX3tGk202gLyAIF4C9p6UgZi1jSE/Iwu7i
HgKUSbe9g7WVe230jJFY8Nx7iUq/st09LNgM9pewStjh42+5VqGWcxWJ+0q8w4wWPd9R2Hqj+YgX
JOwDQ/zbR5jA7rTM+4jRlRBL3FvGe27fbA+jdcM3gL0q4T8hlvNoEwM7TEZb0KNkGuJGh1PuzTcc
AJCOR/DIH/Lf5pfFCJOPgCUa7aCpbA17ay7onXYUZ6wbayWQKTaHiAvwjVn6yHWZk/lQCUJpnHso
Z8DVmMyMBz9zpSliNJd4B8CpIYVXU5MEhhriV82Lfnv3CyuFmuJPHrTlmRm0n9+obwQLMonSJja8
kTeqbdxJu4eL6x+Q4lbpjD1sX9f034bRpyXzKPpicJcrt8fp2pMXHiWPwiDDzP0tj3RF14NKuD99
X9byckKZSvLd7dexsoebKvK1vVWChYJLj/M5mzEHMnD5L0Y/zjIZxSR5w0eXVZMKh4fXkUFbGzuf
M6enX3pJcIkQprrkrGLwZFLpu5Zpuh/finR8/oGE+g/qdVa+zBIJdAM3pFyu22yPf9JTJslGU13K
fcoEDyIAFoUeBfBV4nISGpXsyFTIW4kWp0+ePlVR3ejYj0ejN7MUgFAuXBmHfC3V6hRawg1/bNme
iNFSEb0LFvFQBJN+sgHzQ1lFfVT0epdwzl+R7XLIi0+BWN4Sk0iBuI4X0dLk5Cohe4IlJXw0d8X8
44e77Z8e9ItTVR1j8HUzrSU//OuHixGBYotHV33lZTTODsdDBIJbW6H2m/+FpBYYRsDTnN6OLujq
YzaV1p6UOSJpvGXJ5TWsA6KZc4MTlxfS/CqvBaetqIah6OEghSuDdX9+G9wnXRvPEBiHBHIZUtYL
poeVUroIhuK/Ca6fbxzF+fx2egLmjl2RfrOZNArUcovLY5e3mlVw3zoG/AmAzyMoK5Zu2etyNFXa
Z3xH6TrMhQhqMuqU1BOQMg8cOI3RPMF3ve9N3uEYbrx4r/ZuXPh+CKu1oPuS0wATPJE5kEFmHptw
uvyYqff8vSJyGO3l6GczwaHKse8/waDTQeDCbixkiVlshtuZNY01DvuA5E052uh7h9sdguJDcKR+
/BeE9baUQiZ2VMNRj+hwUqEPNRSWUlCPrIBx3XJLzBF55KzD42kolU4JsVzi9slitg857Xe9zkpx
59JOYjBBHnL4BUvtOGiIfXXZdHcB5ZVRvwqM4VgkpaaJ8oaM2iOlAQCsoO2ol++ZTUy1ILKWTbbQ
M0AHBVt8SssXgnj+8me0TKjemC4EcOy1jXtucrE5iAzMs17LpyfYoSi3yxjpTOjdGltZTInik/O4
4tUiLs5Mv8ZgXnf3fvaw8LcSLGdN2xdu00O9VbEJi1u+tdMjUkyJiec4F0rRwuGyD7ggKrZmHIuT
niaO/d48R9QhuI5cosWvTlA7ume7CGWP/bvZJc7co4ctk0G2w18DECx9ri3dQmTNTPudtLIpP+ZJ
rF9E+pzMa3natcGZdzvUQQAiqKIemud2b7V3ro1/mrDcf0n7SJBtXEvQNlrs2jMLpUeJKIH73zyk
D58xQd8nmWQhS4K7NTi8MKiAIFvkHFHiR8bDVbPcht+g5DuLx+du37SeWuvQtp1uf2geEJ6yELbc
srsUE+oRGvdYxt8754xxfgKeaIT85N3U/2xCljDprllpOSqhsRtpO41AXowh8p3Nz+SeI9KcSbN5
R90UchyV3OQP7ZVWdRmFv56g0VDMWFXjRDA4p2VTXL+Zj4MJf0vsxhjkUz8+L+DdpcGKvWqAV8vW
aJGT0Yt5+ceMSHvKBfRNc7eR1p3gd8Vg/5EOKdSilCJy6AOxNhAoD6vkrTx0ARtgoqMv+tHz+gp1
+dxp5CmAW2BpR5V8B2d4npn11/Q+FoxISXMysNiohP+BNg5Jl2Czpo24HcshlnygepWVFNEseYvo
VTZGQ+tBoFCFQK7Fan/wU/n+4i1ASU05T97zfVFGkyWmg3W+FGPzseP7wGChS9ksk5vTGDiPImIN
grDTvmTRoA/OAPShRqdYXNNy4RcFdrZZA1uZws4+gj2cTxuS1l3Z8/UxKZPZ2DN4c8T5K5qd/i17
J1SiQWiYTDxHud67WC51ALWmKF8ekw+Kp4yqspOh27DRKpnupAALr/AP4r0WkmcD408BD5bGLFeG
CPIdX+4hZShkXnjYl2QEVETF5peVXMzqVk5snfMEDp+owIACsoCjFswECHVj5OTdUjkvgAGyHq8G
JJcktwVvuMTbtPHAtVqbMGJK2BWV/ZtqJtKo73M1/jm4eMsrHtMf0OkTjZl2o+XZi0rzLPeU882C
yJhTojg8qY5KBjKRub18eeYa7v5lfiL7kIfm76snKogihbaUhzgj6ZKCmmg33E/EgHPThx5qzc3F
XTeMxWO+XzRUwpnthgZGBmqNFkT3hX82TmRQ7xz5bZ1fAzEOn8fdVzK0m58G9uN7JbGYnAlD0rfY
SyoI436Ze34gaeQjc5OHrFN8w7OOsufkyECSAhgArmbecYe7lgMfTkHpjaGtFd3eguUpZW56qdiO
jvsF868g8LXFO5C32MxvwmVutdS7X6y+Vm0wxl0LVbQDLJ3srSk8PiZFQ2tdgITt7s40bRKWReqf
tY7JRuMEAcGLZOm6/qbNJwzk9L5KE0k+xC8nj60hVL9sjXFev1ZLiwpNVli2L+ioORnUeG1tmYgh
L0GHiWyt48vsYffVXMbgkxmzcOkFHTM0AcGQrFtkjtt/FBo8ZJbHnkMCLtSv+RpwVvBs3OncIJo7
DIA1AsUgEBCpsMaAGqDYgVtKHQCHeUas4oVIoDnp7sqv7vAb3OSI47kU0w8WcHBAoV3VwqlPNMO3
j0dc1sMnLWtbEiLF3EhOa8tbQWiQDZbrzJ5ZszewEO3lR6HSGRUokKyU1LhbovjJNbLg4/Qv8h9q
BiiiJLJ97+vjjojXBem6vd3NZM3pK4w2ghKWWIjAtsBTbuGhRi6UEodX1B8Q4zR8t2UMEJMp/zNi
6HpJTepNWOyB60YvtCzFrDMIFro7Ira/r0blFMq115lijbevUG6WHxAZtQHk4WOQ6K0kgQloGm2B
SWXk7kWwt646IUnIix0XEtobx7eorw5krJgFO+8rcGVLwLM7HmPkEq3g5WAIV6erFptZ2wEjxiej
VUykI2lMGHAm6mi5ELX1K9w7gnRjSBj1pUAWcZss+kMYZU9UdSwz0abM8CLvKV/r2BUn6KmxgDcG
cZJMwwPzug7Q8gsDbnlyus2A32Xfm7FqDdEZH3OlEmm6BzY/8Y2UvU8jukX5y/Qfms91WuaWmM8V
dCocNRFyTYFw84lucdD+AFhGHNSEQiSW4S7Bkwr1M5GvRlyq0d7MAaBFW8DFFGu5C7uHIs4DZ+Pt
L0JlpYOgpX5p5vmAVvWc5gJ1bOlcrChyvztZuu27i8xQ2BLwo1pmZ4U70HAdo8bPxq9DJyk1hiB7
JcJ63w6FksiefQZv/GmPmaSbdQgyI6WkVeQqJfYlA7+xIxfQ0bskgNgsOD/zKqUi3JfhADpkSskx
OfHCuzbJ4UsT7SuKq4Jf/Fwn8z1ssscHkh/na/C2J0rhxv6Tb4EE35wvO1QUkylssGXoeg6J9vUf
cQhBkE/ScRjEWC6Vnsi05oedsAHEM16I8MDSCZERXA8pTrLOA9Anwl8Mh6in8P5Kei6ILhMmD6eU
i5IkAkYpHmvLwnKksOSWW/5pLtTF6IydRzwKkPxvh3gOzcT1G7GJz4Pu7HuUIUUTOhn6gUBnDscu
uLktpjkCXx+0ksmlKo+/Kwwo3qNsEk/DZTUFSuuy2fncwldyGM76V3trHmrmM2ToILDxoLSGcu+T
0l3xR+51YhnObcxbR6rBZyXqm3dY6dhtyXpnttc0cFi8y8wgrt0hKzdXXH1gqTYfWxjBb1nLZdko
L449jPSXVMhCSeh2Fd3IXXtZrmpU5rbUx5Xy0uhCX44Z/nj9eLJ9mOgiXNrBMcsNgHSSWSg09FfJ
a8cdRQF4gSaSonR+tDFOaudzYZAY2PLWWxJNTrg2A2sGFqA2yc2xb93u2Ily4CDEBkbrHVHYzkTG
RdM8b6Lv/15IVIJX9fiZ0R1B7dKGS8U8JkUa7Aa9i3OmXeIQZ5k/PZ//nXXGW1ILuivgncYfBsTe
NaQE1EapROJ0XmLVrUcM1wXKrdo+bz+EoVTsLKa1YENh1c/ZNUYwkr/zTZ8zwnPxoTeB2S53Z+Dv
3T4v56Idqs93ghu3d4JKQ+D4qL7Q0+xMInYTkkl6PGVYnwVKuYR4pOMcQjcmVXkAL+o863cPEba/
VZnIofvVqe88WRiB8AgOu5KX7mb+ERS0KFyEWmrd1boNwHClSD78C+I1yBipJcFdmiyXc47oQfbl
AsDj/dtZ7aKPwESTsmDav3J6VpeywPIh11eBTcTr0GcLPmXtqOsnqeCq5AmZxqor0EOgzuPgk/R1
1MuDyMPpk6AHHbIMo/EY9n5K9CD0YlMCRfYT7c+D0uLd1dVe+nWZgh5ReY2NdxLuxy81hkJtMf+w
pPYccluAAupKwMu8n8cC3eYVCXd2xnvpBsDtn6s0LpnUJYp5wFwdkmGj31wWOzfsPA+MjC1Re7nt
zod8WmPBwxRxwbHQ9GVXaSJxUcXoNuRMCmn0puJKCqsDPFDBZP22GoNob2h3ZV2Gb5AISpHSG+J2
4qgh1m8/pXEN2RL4EgCUIufhTA+W9j3sig6A3+iey7GMnTX6exLXg6Zg5HSzRPTXP6uhPmn7nJgV
T4fjd2p4gzwRxIuXHcrfK8xvQn6UdBTncwzgG2IC0WFJAsfGFsxioNsYRMkwDcDVYKAdplZcqVZB
fnVDQ+r4MNEOxZS26H+0uwwyN2sIn/Vq2E5xd5xGy/8BnKq1ANXPFDRUT8if/sNc+YXjWiTq+n7p
aLgmRr1x4ObZzS7G0wo9NTEifjB8xOI+mH700HiJ+OhYCTxaSvhyDSMVnyLlhq9FpYLpzqJ3FwAM
y2yfisXh0SQVx/86H2gO/30jm1odxtOj5gh8Qdmb25uAtlLzv98qLLdUII1sOHbvxHPJ9ZJJFXm8
8AmEmVW30SbKH0zMj1HuFBSHNdu1XNnPHUsNX+xSRh8gEeaNI502nXIUMzGU3E/Iq2EBGjaush7z
3+IP24gQx29Su4D4cAZPnhd8R2BNhjDXRDI5IJIXAtV5h5gTVDPeC8RJCvkOx/rmeUSB18txHXx+
3arm1FDZzYw22E9r8J+wQvLC4RIxeSuXA9a8BTpoqgd0Kybx8CWs1pxC5BmJa2QdSVh51URUhSxk
ZN6Y5pPKelazlmn0J4zSFRG72r/NL2ne5ujutyUajteWXPTzwS/wXLkUuRork1c1Xq1hMnrJ9N8K
MJ7gmbfEkaQPFR7UsM0hYRoINwBiI89zbggv05TyhYtQGuF25ODo86ThgPFR8dsC+kRA1PX/b2kQ
3DH7j55r0gVpM84fFmQY/LqsuUjzbq6wIEHF2CmeiJRbRF5KAPv8Deok9SF+7czlonmKJZFxl6Jz
493SUpFrHNL9CO/gmWq3qAX5NDzfrOypplZizm/3PwDQcqusXmIyKnrdTYtzsuzIEqyC5iXNVZdr
A0dcSC6XD1PuXpshg5UafxoDzwWx6VyxlCv5GUu9QrcCqRxXcmlrCmMbXRfMFlVBTwFybCiQpx5r
k4NSDIc/3hQau/T6E5VdaMQCFHbGHOqJw2jwaxmBNNFjrlQXTH8pSXn4RmGJMvmAonEmf+q0jRVe
BvECVrbchfpqCGQH/ooXU78Oa7zWZPNKXj42l0BYFI0WwCxQscyj6RMws3tDTNmF73y/MSBBdRAF
PS/A48zP98WZTuPyLxfID3iXLilEY+Ki6vqzwJ2Gjtlqqq1sebfIq3HfHo7l1unydc6K5wE+Xbvm
T3K2iqaOwDv+XBUeaV3N7pQeY4KbL44+yEsSCYSrSlcPNlcrhXpMbFLv6z0EVTb4988F/AdZphN2
w84owtZSEnDhI0NDK3lLkwQnxZ59rispSeC/TFJBrP14qp5i3KN+DrFD+7TGis2Uzihi2834JdUb
Lm1LbwSRDUHaHkbNa+00P0MPthoG7o1kLZHtd7BHiqlfHTvn1YhzUYCZDEcaFP7ZnKAKCcZbCsh6
SykwX12+Ioh2dfrVr9P5LGespre0NBcv7EQRRFtgEDfJL/pdubGm/OysJ0XApfIIxgMFTG+RNdJS
b6Xh/voH8yvKCO17Xv3EkLv9aqQW2nBecz2DrF/P1zoByQvwemNl9HmsaezOjFqnQDR1qVsg+4qG
J42rOZmjoq2jEByy/hwwht+I6DMOF0Wv/far3GV+hdmAZypd7JnmbATwyc177LX/vnAvb1RM3eEx
UoSoeFWuo+OW8MSJnxgHozkWiBmXhyR+nNu7ui5iSaHcsa4iRsbHtlPtlbjqW0V2RQS/mW6qxsQi
pc+iSouLwRrzGrTkjT045XZ+WpKPwnInCKb5NN+peyXncBytNmHlYxSNQ3EjDd3HON9ZDCvd2tbK
fRaqulquOz5RDazEcIWjlvd4gZL7c/Tg7mSKn/e8UG4vfsGwPwOaJ0FtKEo4eYH2ZdvsQUkPpkr/
S+qBg2pfLbZePvoBd9aBHSiB6iVD8vc/HaE8EHyLtGqQ5Jsr2trBgPyxwojWEQzePk97gqf2vLPZ
pux2eGRjQRMByp6d4lCbEDyaLjIaJh3ou5aIH9q4pC1ONKELFpcVy6MH3It/eX7pG+KZBZoBNgc/
WVX6jf/wEPWlsOaKZ1X3CAFXO3DhZSg5J5DNiYRUtCHQ2/dxMS9f3s6p5JyTxWsTeUdBw8e04dIt
XZ0mHsCP0f3M8gq9KbT7ThVTJBttU8223I+/JE2o5DCci+RfiNabqzXNsH1y3GQ7z44VeErcr9NE
wau70YNDPGWeHDOgXZTGcLvRKk1cZO6cjvUt5qTaX5QF1sU4vBzUmgagScWlZBpEyMak5LKiqKWe
SvnmMRIKL1XyIHZCKopoNHSdT2OIq2r/EqClxzB5NRC8Cjk1ri0FLXxTDxoyc7Isha7bmMGwSOHZ
jGfhDU4+18qVYtKaJFBwiJibjvLwwGvfgFSqtpBfLb9URoThxelTC56Ot0di0TMjo9wbxhwy4Pcr
Y/SWIhMs1ZN3a2qZfHATr2kd6e2be6XiIToowZ+AC7+CiQuMydUpIs7En2QWOzE4PK0bP8G3wkMh
gGbhhyCYL+oq0lxPVVipkZn+wXf1NO5ECCcnOkBOWUx6VpZ+bdjlbIkNrtruhZm/mfEBZ7YdZCoY
TNzJzflFnVm0wSUYxmJswPTydDTEYJKN5SuDUze/Llpa6mWh1+yBUheqtSumG5a77tt6Q+5g9Jfv
yCMSgtDqJjLU0awYyaOx6G9fZOdkgKO/oreqkX1F8FRkP/hX50nuDM7EHfluVGGK+FKrhCUSkNK0
m/7MzveWj4dQOGZOuMdiIAQB7iFyRUKusPSLq9nkHuvqDU4ObZAKxhmN4ztvOI8nBdUZUOag3xiX
YWj/yqBaTxZzlECIc1Vr7bnYE0e8Y/G2g+uW12nhdQ+eBY7Am5cymKgj7+zfVRogGvZq+uNJfStV
4k7U+G5BNnCu0sAmHnY/0iDJ+lj5n/MoaBsxHebXIdbinsDQXwyr2EZC6DrmeEGYMCAB8KktAf1B
qXBjVeLPQ+0CAaM0Lml0FvM6No8rg/33nEoKmiTI97JByUyUdGqhdYVjLwRYx0WoiHjy/XuXpWI6
n2mJE1/jA7E5jbsyPjOfaVVRybda9J87gcQ2V+s/ROxWW6Zg+UlC43egAgTASlQvfDr2yfCfwviL
IG6x0WRmdZRtTdJCpYoajTmejP2zBJfqkfYqqCNBJv2T2dl5hdCnGxmBaWLu3Qe0xOyXywk0Vu9U
Yg+3in9JIQK2PtA2U7zR0iSiDkg0D69fmp6er/PNaWPKB/CDzrVUSJeT2i12+WobVUgu3sn0hHty
gANLW/NanMEAmS6GPZaKoLPxZK1YLvHFnUWId0IFscGLMx0Fk/LfU3ZSO7um5u7pwBBW8/wUmnHl
f9Ou+cYZKV3yPIGuvvQjK2/fcnrjiNXDbmjtVaBMCheJG5cpZHzO5bErjv4KgUNiJhemV2PbH39R
os7WjBOpaVBEcQP3Vnvg6V+lc7iYKKtANfJ9AkWvPHs0EwvBu0pH6XcEbpVihenapX1IVpy8U2ZC
qKIf719RyyLTsQVVuHtwfyMzeL46X4a/Ne75vT2rn4gE0iW/P217TKWEQ7LeX8Fj2/W8ktHqapEg
T4b3olyM5jEhzNA1Xg7DfO+TjEWugxggDe5V4CaZdciomNL1hL2hPr/5lqLbrkJs/3vcdebh7+kf
NQ2oS1lOV+QtLelYhH1CNleaInGsW2jF0Sa5BIW2kVk5UC0jckV+KgNX14GYCLSufFuyCPWVfUAs
RAPJfgjBYjE6fkX6QRynHbG5U1oJsmyhRTUje1mHQOd5O15lUTZmQFnsfvYEOUs+/UU4v1NkWTSi
DSXhTZJ6dWMMC3Sz2WXf5TYftt9/AdUiYj1vfuDCI9OGHeWfjdaU0iLmNCTU128hsAXZhIJ7HKx9
X+bAI7zAihuEZIs+ROkIT4p4Vktu3s7lfyNLzhf2gQ8Mm297bzzY2iv1UV9v8nRm2uJOLAj3NLpI
YnE8Xscjha7SffOptJLN9t5rDfeICewkBPkLUHFihb/2H1cVLtYeCPkv+qH0h4CXtHHv6KM8CT+0
3S8kEK6Y7N5RQFQAqXjoXuRfQhUM7JZXmOTSGnROv8IxsgmJcom9dRsDIewxTjo1SFsxamst7RUi
iQrMRskT556WoWRU1yLxqBLuwMoZ0Ej71fTis72KcDE61YGzh5imunCdTbMITMz0HEOdTM3Kp8kK
+gResvBdq8W0WwVnMN0p4cLSr41EOaOD5Iz3cGKgUa/gbZy+ftMwmWtngACbOqT3BJJBBwMkCdwJ
dxGmWmN66iVL/gCPj5qRf0kof3L876nJUlYiA+SixxPraWHI59fNLOTJXTgrB+A9B5TN3BCJZBtP
z8fBS8N5/Mgxk/xABbj6QhUXx9R6pRB/bCP44PoYizWy6IvDMy9bK7zI8dgizJyQzz18D6fV5bmP
NNtzGjRSNSoobPQWXLDLNq2Y1IHOcrI4+GrW8hsnFwLuoMyXjZNs7apVwIU54uRRjZS6ZyMiN5W0
CsIkOADe9FOdzROyHcFIjOiZVDRftc0pyC1VaAFMnuh/xaoeZkiy9rlA8Ea7yIUSsLfElbDl28lc
fC4F6kGAiJYJ1VFMXrRbsGUTo/Zh3Afw77lBLnQSaqAnI+Hno2p6B+3HG//8lWD1KfWPFIPUDxKA
lsoeWcw6UgS81UvhkfvBgApEZaD/jXtuEEoGI1utRixJdlE6L+ou8zSLStmAbfeINkst9UmGHYAR
BGPFGsxtz9RNZoaCYA96jUb7hRLWV5f8nlilxqnA4uhAfjNV6IfTV7aMwxF9LzHoRnSt9u2Oydh5
8SegsweIrOlyh3dhJD/pcgpWTisJ0L1qSfgwvc25dGNv4JAJHc1NAm7b8qFwL+2CA5bJQBQuopt5
7y+hKuBpuC1KbQj8jMgVUC6lLKAE+MfuQLR4rT5kzwbHNBgiWxZ5zy9/ksSTe7twwuJBn8nyu0sT
IwG4I9LW98H67dM5/y6s4rlWqu7v20T0NJ28YxVXdnsHsM9WzClqBDVkzCJaw9CaptSVPbjE+cjV
dFKkjLFGH+FPUVH0Sltx67yWxOUbVbw3T79krwGJe8T8N9brss2osW9dehmUD2gfx9gTtvIkLjlh
XGolLfckyjFb/qtXrOjq+2emcvC6tBrotNEigmeZ8p+PHKTO+GEGc5onsJF+pXSYghEK2JwUjcp3
HPRkzcULPbYGaXgFoWQLXHzSCz32MUWgAGlAdVl2btyYPNoODoSYddjHL8Dm9zcWFNyzcUsyORdM
jtZVlRXEY69yRvmREZ7qDx4ac1Yx9L2Y6FQghL179Ah4jfBHJvFL5oV4HqMuZtJWUIIxHzYTgwLb
1nFs6tXraaLcdw3PADDuNE/Q2XZqXdVsqNGSNJ9dtqCXadjodWFiMAstGGlHQE5bpVRdI+nwt60e
KgHzfsiK9EmfAWKimZsIwIFTm/6DcEbEkZZ88bzP1HZ7boZ5uLkeVFB+0FxOuaEWJyWr3bmdkGA9
KFJZbTTEdky5SRTXcCDqVhSsmtTgFmHSgq0PVWQOJPfXrn6dRty6XAewezDmIMRzoB957LyouA3t
TzcUcGxe51Z7RYxfiAscoB+jq4xvduzoe+Yc22kQl/Lb3opmbUOvikZcZ+mNGNr65gdRvGDFQv+t
9hUu/7KK4HNbJAv+moPvz1SwBAnb+YN7CszfBK/DUIBLNBr1vjIjDqMieCyydf3aAHmCaS9pLZzb
0SyD2q90U9UgP2v4049aASmXXRtF/yX1zAV64QO76lAA11E1XXxQ5qS9o823esd5K4HDXH2ZZqyL
4SGiKQ+DyVhMmmpSI6NsNfEEKA5Y2qs3pud2tai+7XSZUeC/yeOFNtIcyewJHqAzWTvZ11/PzhZu
9789tfGIOre8TDieHat54R9KqTlIRp/rbRglLMaIhMNTQKUvBIBfejpK5UJpJVf355/yOkQp9foS
WTvLImq06SXAMOcuFfM6kmfI8mfy0xJoWygzp1bIWhWRN/wCjDmdk03aVycXUkH3+RqcATWy5R+2
Ru9ZUe4STWfBm4GFYK8Nenid+NGHMAUGYrwgYkgDicDVHVUruJiCKfZ7KLnk+Cqo0afyhgJJe8su
51P5MAYqbMTEA237ZLZEk0Un6jACaVqMmwCHGM0KjGL1K7tv7/u905Ep8OFe7Gs4uRoDxTCkWOYJ
O79yg0dOMtPnjhaBfEH7IwW1pSG4OHIIT6++u1kcdZo61/may7Gnp0UCVNbRW9otKVKN5MuCeAIn
r+BQWeFEI3etlEXA++C02tc/rJxm2E0YqoZ86VcwnxOkOORp4/inkRGRokJuFelkPoqX+pxwzt5d
E+soXy5zRCryv9JJ4X+89W/IaR2Cb9UCHORLxl4HMOSvXVGRekqYpvj4KmEmjyY72AaAEWkVU56m
TWF2XgE4h45hNPBqI2LPU099UJKNkrGIMpOtQ2+qQMlkGPDkTN3BoI+9jsEmwfqqjdkCP8QdRVId
yME0dpJGDzuqz9G9XkN2nB0uCY2nb6/y6wdGG/0Bwvvt1XZtFUvNy65z7zLJmFlCXhiMJ2nNetZc
CzVprMy9/W9pQTYwS0TITrcMjoVNCBrdlOlx2/4oFG1HDdHlozwhpgINt6QNkU3SLCs+Ln7n7KZB
7xgHsIaEFWXZ62slmlan0fCGcQBkf3BOEzXf10Ahz75O8Je8xeX1swtO0NphyDgCLrFkx6pFqOF4
OIkwyk45zLORvh+00ULgstedeurmT2FZowT+XZNCHBnhurrQchdLV7qxT7iaE2RUabuhSqi8tL2l
5D99hM3NCmGwcY14mqiPfi8ERUQ9ICXqCLMLpCa1Coi/rhI97nmpMsQqMUE1WkDu7mmMKWRUHEmK
18gQiTJ3QaS7FW3pJlwecndV2Seq0/raorqd65zuCtHYF/z7C3c5E58NxcHKjxGviI3jvYOrFevw
Trx7pE3Os26/pPWqAsoMeaQ4muWwYmNijcFFL5IRy5laSxgzpSchN4mm6h7ZeG24v6aJy6//Pj/D
o/NBu5h9jB1+iUqv2tvFUvZiiI3noagTTMxpvXSxTgBChSN2dxy1Qu1wdxOTZaQrEkSzHwFjDUMu
lyLvNl+0SfBdHzEuj+baF26yeBig6ZSdSjC032+a8Ro9GRrLW0PCMMGM2OiiOIz1sFT32G84Q1+x
1Pwg+MgOjqx39woeu7ntMBx0lV8xLUttdsLex1a8pbP4UlhZWfi1f1fQsWw8BqejTWqR+ZXBbiBU
md3dyxAqR8eWaNo8s/6HqcDbMkcvltGThct4M8d+La2of/W4CSIrrTrEJbOuY/tQjhYtK++ECbHH
hlKr2HX1hwsD5pABGbvPzh4Y9qMax7kUHgLqnujj3L3KhoMu/omIk8yRsT1mD6t7QtkRgCxwRQaH
Bcf1p/UF8SQkhcFWXE/H4nBRLiiYr/+1d7WVpdfnYvw5sNIoyBh3w+YikxdpHkRe9vNB18bFMwLs
8d2VnG9Rzu5/PeGPFSy6xfJehlaz/pH4FERgNBlLxoCMvpMwFVnaU4yPROIziE+6rMlqyJVg6TcH
JmthMvRJ2BeEZLePiKtd/WyopCNyrhgrCQEZnXwJF6r7zrztM77wDVBgOYI3rt1svJ5tjwk8wdNw
qsXcP38CNyKaIoxHairCivzHRmDyYSGPk+3zkjcPaFLuK0vu7Xsyr76LsHbPwpHyt1W2A44wDlaG
nu5mPDlT+kEUX6JHMnWdLufN2pyjol+qoVn7GWB3vi6q0kd0tVXLWdDkL6pQ5JA7aZyDQiLGu0IF
EZNcIMHtWETj2p9L03VMqJmF9BTZuN1nq7Q6MuHZNmK5NJtfmK4pWR0wJBznlyj/oHcmDkjjTmIa
vLRyGaOZP4bOxCQqU0/wqeLON3BIRxI6CZBAnS987cP5x5e2d2EYeYb3OCnYj3+YRAcLVT1VuIAv
FapTLrA8hoRt+1UwULcLC3/NQBCbp45f3rBQkQFfHp92vUP7dCoc+3sTc/7TMGwc9DM+IoYxoyBO
nTRT3SBM4wiySgS0gwKWDabX4Ypu6x/lqgxOO9OZV21mWbOAYkD6l0lRuFI3cWbbUgDikxUy51yB
DARYAMx3I7QLMlDHbktIjLr9A3i/FE8R0+tszaUPQrnxRjqyQPPFdYOPZOE3AkYqm02gFAp1adbL
3/6ZpSZZrVw2GuyYTtuGKYNEMElJ/8u6K3oZj/8fNQ0c85Pe/u1xLKA3L1z2Asvy5BMDOZnFZXoR
GjSGJv4OjtAXWbbCXeDSDkQRX0E4rykVofBNpWz1LVSX6o9HdJR7agA833TEflVT5eatixMPyMdv
jSatk53zoWlA34j6HDd9roYmrLziULrNFVwi9+p4cdgaqwfvdkEAMMLY2KKTtTT6JLG1GH6xIdR2
UrORtp8snxvRFHzApPvE/Vh5Gh/eJ9gMQJ5O1RKjDWs+5uxXfyCAkbDgmJV9ZoAXKcHTMyXEyPlM
UmGR3qcUdPfSXh/x0kPfqnGMps75O7FjpIGmJalgdepz3OQJ5IHqsH2uMO0yqoolsrGbimQJJZqf
KrwqEqloNQIdROBr8/ZKqcGPxHLlqBmKM1EBgC9rn+EXJjTDJE3Q/GnNyUssue++DNOcj8bAlhXP
2WWF2EK2VNIhb5D5/aN1Ofdg6+fRydwxpmzX61tY/JjPBbndz/6i66mPIwJe5m4iZEnueHELZOSC
4KsifGrb6m5zB5dfeEO6VOhEET3bDbRzpsTKYjVWD+uscEESm8ELqdWCowJf8ft0g9Ptj+EBCwiB
EbQ2DY+dN1rLWLkgruPHX4d/WKSrvblMGSZUihHZ99f4zMUM34Yo+k/nZ9no1e2VhoZRjL6W7cV6
1uo1cDByTIlaBu0q0Czt353IzurOgW45XhODrhdsR1OrqvdI1pjJAKKrTB/hdnifmNJXyngCjPH/
Us1dpTmEjSrAlJGN6GtQa+IF1CmjlcWA/LURW4NctGh/DTz1wU/oKWQRbn5x2mYWielbutxyaXVE
I0vEFT0pgHZhIrX32Jz4ZlcSuVm1rnySeI/FslVqkMOqN3PPrH3PMPGKHvogHAZ2sg7fVCim92Eu
mxa954p18mUZpJhXcIlPkORgIn6uOfDRbFQpMBQSiIz/kWzcrPYSuqPyY2rLZncEZctI8Dal8yAU
o7s3wtC4fMhGVghRumpOzsEG4FFFXrc9Ue/6dPv2ng+lAEcaFj16Y8pGFGmUtcrWV9Y7XgFICvNn
dzRaG+wTeuUWcfJD8vpXn9OxjCLV/OP1DPd0JVuU1QTWUu9XvEfD4+Rs7PpoSn2dQ3UTLYyovTu3
zw7tRXpQqWuyQwi/kLv5YNKl0PV3FndlvqpEhuurwTgGmMnMGxNcEpDF9rXs8INlxk/Ytv6pyJ0I
naDDGpBKcbRJmnl7hFnwgIeJQNEANBx1NgAS0ehR61o9urkmopTIqTlociMyUN9H9zBFcizaihaj
vx1OjIcrlCRlgz2IHEYPHtUBZrvL6R1vzePAJdhFq+OAmiXY7McB7AI2T/G6tSts45UmaXTBxDxv
Zf8oZ5pkfaZ1cBt72e/YAJiBS7E3qvfPtk1mqOB3RqYFpI5wfemZU6N1naZ0DSJU0KoiM6cahIM0
GpGkWT1gg4671arAQxMGryPinUNcJGFHq4OvGwWQgzewe3uOkuQDqTxpA1BxpICOnXBo1dTPZtfE
jWCj7XrfmsSzN0Ww4/Z629rJURFMr73z2jOPol/TlMmkebZsJ9Cx1FiWQDXAa7gA3CTZWclfRlun
OuvaHHQcudf1pxLStgucBvSFX2vlDkjDu6ob24IPfEQWAqh532spGOyGz5qCUwPU5A6vVc376u8L
57OHNS57om4g5u/94MSh66hZCkI03p8rTH4VxP5oHbYTglRPhdFkHoyH/PogyBrvMwEIV9kCFbBR
1FjG2mLwiSHBnYzjqf/cNl8mzP6LBvRmI71dzc2jnYasEQeDyZb8OUz21GHXxayjxUF0pwNOinbU
5hBB5DLahQTKPLhI9LbGrW3agPZ0RApzZXUbN06Nbg8zT0iUP+4Jfvde9lodA+P2GiPdYc3Iiudd
CbQdhiFUnIatUQRwCuNuQccZl9gNuKIYJ1Tzlg/46HhnFjXpUx6a4Tc8tBr/sBCU8kYEDkBKax9L
9o2rZjyQitRRlX97QxI6EuT4FS4u9jEjkhVBIXFb9mj5otXGN5hYu464fSJj6n+DaKdOWSnau/HB
ELGPQZ6d+UHqReob8J/aQxmNrWCcUEyoU1UI/z8RfsOcR8In48X/+VpVPa49jjBJAgxJnANDyxof
MG9sj5I91SbKPZeTcwpPhCCrBEKXEFoinExfmhnk41N1TbMCA5P5+OnXRMxKW7U/RLG6tAN5qQC5
JweNuDzHKfTttCVqPnGB6Z97NzJUMVKBYxJtjSXHLKDN0xm7cEFeIcPn6l8CJxNza3zhZq7sh7Xv
rx+SsV508s+95/R9MXXos4M5/nXKX8d2obuxJjYnV/l9ZSVijbmodw6vrIXYYbZcm0v+MHrip/Ci
5higaCf35ETl0OOvg5ASC6zZq6tlryuKvRVZWCJD6SrxvlVbYf1XmFEN75J/r8MIGk/2uA7pQNEs
hZKQ4UGlECOaoNWnrG7/DxdeElSlcFQ1ryB8ChMHT2YyyWEg+N1euB6p8FekefQQ7mZ8rfEwUty3
xPkgADtbTklOB3PVKqGoo50IpsCrtE/5bMzhPLzP1ZFGvhPQQ9idTYdmcZOKA6zCVTcjv1cQur4O
TzSJJPhaRt2I47aMDwphrYYYUircLyM0At7KDBK4YPY3pFocDB4+/F5xFhGlXUnIiOMssOpUDEa+
vZMwJLBQZQ+h6xVGuxPP3M3MXDOhiOEpNAXlJfn4UBngh+yltpkZv5krTCutRyNsuuejyQBzfBWd
HRzg6M0Ddk3sp33pMQtuad/DJNweFqESkrPmsHzjeYg8ciTZArw0yyUfLv2PMXOb3itFb17+2zZN
5uPMNuzI1/eP94HhUqGSvyD5wI2e6sPBHG+g5Dd1rykpuNfnkYhiftcMwFN31qSXIVQfwntIxvnm
Uaoq3YrGCgtK7PLpGq0x7P/BnnRLw0jdQUYHlH9ig84SGJmpY22/3Ezo/7+k13AZFpPLZHC7J8AY
vH8R8dK4na3LHZT830uhf3/TtUH3QDPx6p8mIvvTGV1dHdHcgIw2F4fzE9r0hz3mbFXZXbJkV0c8
IUucR7Sb4y5lUN97RcOiBJ+6wSScaM5/tzgcemQdxxoRQB1LZszanHtBIKCudFmSNxfa2wMgdiL8
suTjFTIRhEtS7oKduBYqPZ1Z6Vupk/gDbecRXsFATxNiOX5NNdBqV7WcJVqa1mD8zdcIa2isYWRF
tuvQHIRfaX71JaYBhSdVvyDFcEpCiP0cGVXQUGErIj8MlWJeCLS0ZxX32xHTybKS8W+x0sPWZXLD
m9z31Ju97AMeaG3dSRC0M7G5LFm3s4F0wsBYWE0GKC+4h8p9XD+I/zbkkWZcA5K8qN+hb1Qg0HyQ
bHbkL+XwnkDlTTei2bDBZ56kE0d79VWL6k1Echo9ZxuH864IwfNiYrXETG2DfuKm5xopcrYy8MLx
jVbtom0sAEi75vSZJhgdlvcH/vLcRiGLYxaK9xPnEBPTKwDZO77GVYdPcFQ7P79FL1ARojsGT3LJ
/5yJa/upi+ZbpGf2ODSdz2EFuXWoxD1NPGdp1PNvtURbvQkIWIS7P0Ik7xUhd2VFwunC/cDFQx96
4QMABtHnsAJZgBGjsyABkMtVixpBct2at/m8nlTU/szMEArSaEDMCZVXCtZtzrpI2HAfN6lHONPD
8nUxZ4Q3s96A0uRfnS1Wj5uDYP0PtDGcF3N/Y4qWVFYL35OvwNPtmXoXqxqfytx5NMuHYeOzh3kP
cF6xnzizq7f6E6/WPNkX3t9FbUup97J7IG2rblBklmNdStCPMlVbI9DTyqVcrWJ5l87rcXvFIKnR
pAeVDkZWUCP7RWgt7R/VH/S/UkPEwrAvki3ofSGttn9sfDfh4G7PoJmJFkXwZpS5eRKmdLR0cFt0
5Ycd2+c84scwzMgSeUZnlhS1QXjyCpQdj0l1ibECOf46R+yauUAAJR3FH3RkOfAjXproxpO4Ct59
CsTysH3Wz1SJyCNJdDQMSphn673Oo+TS20NWOkD3UxBYLQ8ULhKS0v2y/KCBIfy+ksoSBBC22/IL
X3cXbpZ2xuukICWqOmI90wYc5iap2FBuzaQSct5QWMEQFhwXsdesJthNj/pSwCsXCJX7qoAyMo2c
n8t/yBzuCaws8iAMiNxg8/irICKWEaM/NdWcFi/wDguFpWOx3NFGVExucq8w3re7NlqCGovi8SHJ
tA6OJgCeETzceZNUgXSTt0H/dlzIVAig8gCKikepX1W+5wBdYJNDqlz6XoaND/NXeXuT/NGhc02Z
4cuTQmvsnuYvYqt1xBpZlmunAkgMAY2spJq6aoH+OegRoedFUsJdqfjUSGNa/BouOjN6qqQHceT7
dQ2P7Fef3HH8NNMX4+LoLCNOiB1IZsXoF645gnGZ3nTK4H8vFHEbHD0XrlqmrEv6VaaKMBiIugLM
qcZ9EVmxLTJHb5IbgZWTxdjZFePWbhKLhEkHDKupCqY8iXKwVp/m0cOUElIUd00ZQFQovnj+5l6Q
Lasda/o5tx/n65YEvXECc2ktR6GgrMTESJBMYtExdNrTcZZ9oLUAY5iIS+aXvAcrb1b2ZcJIaoSY
t1L8vRrh6dxV/SyX2m/oYVvGzUORU2QwUXaASo/3KZny8QaXS1OTHM5UqFW2cyDeFuk7df5li2eI
YdhCeJ/HAXWutJrh6vFYEruvcIRn5il47VxaB8AIYQo4wXjdEGw+p+pCG6WLMZ4FLACY2GcNf7tf
/wEFt7YIKRILYIuqP0Qw9u8I8i5C3fkTuWUsGQkzlD+O8LJZSfZV+6EMWkBWqn3f1CSHDR4/6/KK
JytqncWhkZWf/HGL1U6XkPGAnVWZnvMgjnYuDw/g5HNraGuIdkU7ap9DUxViscNMWaUS+Tnl2pz2
f7cF4KkeQJbjKp3wRP+DKiyeE3tlDpBxJoJ0GkLeYpHJ68g8TOFDg1vFZdaKnILLVTACLex1W440
1pv5F3WwQNpFirWrhivvNTCcws0pamZqOLNieRbOHK7AjYu+N4Dzl9ekoRQquIv+Srnn9xnRFf7r
v02Qg4PTeZR3M/FLL/UzhcVRZt0R3nDqfeaHLb2JCCVcLDd1c+pxNeSZlLkOSZvyX5gxay66y2KO
pXP5lWKymHB6Df66NxskWeKfZe/kziDaTjAKfZCvZ21vZ4ly9BXUnowCghgXMSfIhLFQhx+fFAgv
Qljj/Ol5XCwYNFsAUsRmYsqNuWNlUgISlISoeeduhPXhHohiiOypMwhXEi6gqqq+XRPEVOHUGn9W
wjbaWmMPjGLdXIp3YZnlYMjUAyGidcs8aIS7rIDJulffEmoTb0NXkI0n5xoRbCmq0ntjO+kE9uw7
h6TKxG3itBqVbRucb4aoVSnk+kToOsvwC1skUlj8ASSbwC1S+Bw6Qc1gsTif630oFjuQv2qqzt0F
V2ADrCEGZgqGjkH9++0TpmI5Fh0eHSK6wkHGqrznVm5CAEo96XkQCiUbUxr+js0ve+JsWOCR/xa7
SEl9FlYw8EC4N4tr/aPQhb/aQYXulsuSejOCUwHGrsIZIiqogHQe1n4YoqFrp0/a+vvaoSA4XsLx
yRxM3OUPisr14RMppc1WRpn5v5nigqmbRq9dO4gt8di/thZ14qpyPpInsZcvTHa//2TYBkpp1jEb
Hfr13rBf0SyFaUP+KSjVlRI1JcOZ31Uy+h5/q1HjdogBBv/MCjx9oKmQGRF5N+nFmdwU9Xar0SiP
JL8E6CJkBTYt/B99De2iZKCYfqXE+KMnYNk4hOcEHoOBQO3Moxh75tiU4GxVqeO3irxX4GIFwpQm
HAaWePZVmCbZHdfhy9LVIAVkhI08M0LfteJnZVNdBlcRQWvyd0dXzDeapUQ+/drq9BP9WP/N+LDN
svA4is6Di8c1eiKvOFWTxP7qNliQwA1bn92LmYHEqgfmPWHyZgYb+bAMKjTNgy6D5YWxnFl87zPF
MV8pv9de89GClTNTtjgyyH/7u24NVt4TUvmNN5bBkH4otwTh2AqLgupm0yt+JyjvgsQFA7RiVoX1
YeeK20i++Q7WgWzjq2MGpfIoqNYDm8Taj9ZmWGgZULB1it08sYDNy+BH5e7GRL48R5r/hvEBB+1b
OHZYZLaKWksbPf+Kg6P3oWwJpO0k+KTpg+JnJstjIML9pm37Z5HsmWi9pb/F/BMKUI5n2ghnu1ja
HZG79VCcb7WV7RpTHX/xzsdi29pBPwyX264xxUd7o46obD7pfrx88tGyYOlZc91HlVCj4+iBplZ1
a4Kp4yUtwQnY1mAL7GCWLohB20oXoWd48dRpCsVZ2e2GgvbPD/aVuvSnL2rj47qsNGtthdIBUMJP
JtmlIIP0uVus0rDPZxFcgtml790XXXkubFd3Ra7CuWtZs/AkrpDMI53qAmIUwk+hvCk/iAGdjbfe
UDf4mqheNXWKQbs/kXYWUSWDMQ60BP0f1uSq19PfwiVURAVnEj5SIbZHL6cZZV5jra9Ty46bmpdX
Qj2S/av7BYjxte/L3M+Ur9YgR4LdD+r/uVX2R1cGMAUsrYpg5CQNQxgGXpMUx8SdV+Rhv5wIO0lj
CtzYY+EE+lxwj10l6mEQWFVBQgoOnu046KPKfVrom36XNaAKDqPkGbp0hH04GMd63oi/xvW0lgQ8
4Gfnlyl3yg+EAqn3blYeTsxGNc2p4HXWJhttYl59rnwxm24rWuq6x1dglqFicL+qhs9OvxC0kpAg
c/H6ak9nrPsWK7mJgf5q6P8JVtzezxHJ9us0s4qA8vIZmBZjOzLyuMJzqqrvchT8YTz24Jt66GSy
A0kcbvD6KlwGOtxmkz+PPiXIMIZuV7nUyM3fwvhLQX/8TB7zkRW4RYmigfar/D9gDU9tPvCvE0RC
HUBGIXC1mgtdQG58h4GQlzvpHFh2mxxCDkEBfFFfNOhdqtGapRsMpR1rcS0bcGqUeMZZyQMnmslH
mh7IvU62qnwyOjH3joQ1HNWtZOVgT91c2z9+BD9dMHjoSTK62UIohHTbkyt4CNarZGas5J9yElUe
GXw4ES8PY+QxBgWMnmFv0xZ+dbBANlVAC5m20jRGfRsK48XcYzgkk/P3ZsSIp+jm8UXwNUe2CzZI
qJazqDcJaU4ehOoet3vvk3Kq/DKGpru11wbg2cutbatvDwm6fCjQCW/dZhv50OsaxJd8XMa3miV/
60OxN7H4kfYB9Jfe/ODTk2wVjFpnf/G3ajaD8ytFuPhII0d4CJodFWbjpwtCrQbqKE6YEWEzcjbn
YZfiK6LYU0Pnpvq8e2qLVNsFBDRxGe4VVbZEwW8ogOPinzoOHs91wLI6Pk5j/sv15Uo5IwnZL3gu
1ZD+gctNBsUbgH4j0o1otbIdiAEGh2SmkLP4bDS+Mxl/aneHkpfJtkqslTva1NW4FHM202NY/vAi
W2vtwHD+vUq8VkH2arlP99MIEzicDWfTaa7PCrnZYjiE/xcOwaMwBYqJhlV/Rlo3GaihzSFyDMez
2eIXI4LGgHdKGDjiXmOcPFRxpXQtGzhKCGIAbFZrFrbsGgEU+s5fctV1n3dlurk4+AJp1NJRNFdH
cZE80iWnAyOLxhhNvPW0MvmlGiQKFxLAk2aT1cnCSm6yBDfHRQN2A35muUhgRDong3Nxfe22yFcT
eNULA35S7awbDn8jABCjeEVkSk5I1hkAC4TIj8Ojbn1HXh/UMcCm8a2r1fu9L4vWEagwavvDeCQ3
GBgk0i/vj15i89gS7Yraa5oGCiKPoPVl17kscurDsCpK/uZGuLyk9v8F2i4lCMzrGcoZoz63T7vM
Sx6jUFSwdCpiNxcYA4UnkyobyiBQjBVny1XBLDaL7+uETKsRHDOkQVJGn2ua3BgOkDjEyoM8epGs
hnVCm72WZB7qenKpZF1E0Umj8rLqGdX629eL9Y8brBY0eSsglEhhcLvxSli1N9BYV/E76uZuPO0m
w1IZ2BhSBc2PXC7mPoDkveN9cTJPdeDB8zD10uR6/oTxOcoB01SToAklvCHdIo8293shkSyLAh68
WjKpKol4srJlSvSzhSu9dIQMvlp/yVZohCU6PKvVKrAJjA1keceR+qbZO/TPaSF7MLF35Yg2v2k6
/vXVhahjx63WzFm5b1+rkcMzw+sAsGxciKGDhKUSwzNBNLgW67YUV3Qe70ExmZ+x8WkmWyH9mWsO
WX+x/x/ansgYjI9KqjQ1giPmpTtPVCwXViMoSd6nDNk3GkrnlHCt1aM3nXtBmb/fQOSPx3ll3qZt
cAmlvUJuQj+FkynmVXa4pjoS75Qb2xxRQ4QVZh3pD8F3HKKLTbFUgmgMIlF25cYYiKv7OOOdxlj4
gj93mhh9piUKaNdQYI6qw6jXMCbfJzpUvrT+MHmZtHPEpOKKu9D2AFtvD9HsdqHWxujtYvadMyaM
rWbe3+lWynP2U5dTiFEFiE/Tri0qzqnEbXSK/3ST/norbkSOlLNwtzHyaxTS4BRt024B0Fo/O9rt
Td1T3vnJCFYUa/IiEalLJ3eZoVZs7BQKm2+VSaU/0U9QsS/+Ln3IGURmUcAay51nlxH8RoKeIgNM
K0JJDDLCRbC5Dp5Tqehe/0f/La9zUvRyUF1itQEomRbovjG1VkQOh4bBlKDI5PpFl9AXJFV/1Nf6
IGHNtwqTmWxOnxF5rZh9+/8uqFM5qyYgk5R7bSrNvO4jlIEx+QgF4OcagE0h6pKWcXtznHjWoXFD
4jbPd/f0CpAJjYNoOEGMl2uyTTMV1Ye4lqMQkJ6vMZ6H3Ex9hDcOgsPQvnHZvcNJvpPfJ486MLdm
5fQNvOVzKSgazPPCWvcrLBmA/mEYKTWbvSztXsmyKRzc15Dz+hhqUPGnE7SDohArSFNHa9J1MdVH
0K7C/DyHVlDrN25RO3MF5RmBpE7A+sYORnvKUNnprF1JN2xzQZIvyFrdcSU6VUo6BSOSwt/FMycl
YBG9ISDbHyfsp19p7qEyTPVXG5CUvYq8M8Obai0V5KkDL9jTyLnpxofcJLNXZ1DbnP6FBaJD7dW0
DCfPkQ2lnYUJmIQvI1SFaF0atedt0wea+pyOMUNDTs5KtdZ8hK9JPDNB6ltgce0eDotrOv+dJ+oS
WHoViuMx2sPprGlR7e4d5Kar+XjLNLmwax8iUhP7jXcUUyk1Z81JXs9BE3llpUlHO/L6VSam/nZd
D03DQo0l5863xUZrSKDgcbr62nBmLmon2YBSHwELRSJRkK85wBr2Q2LNQ/ySIAUVAw7UlJA84V/H
7JllMFCARZS2h6fYilVNxgaMgaKWCFmXpmAhgrdAEtXYzK5/BfwyOQRuamiXwZARK2rJuHo+I7Pf
bY7ZN2DveahHGl6AclLkRo+HoVOVLWkj3jfh8Gv0eWU73z9nROpSPYPCoNQjfQ4rCX1UX0ldq+Rt
Vjo3pg1QoWO06EUH5egsxuohGCKwPPiQCRqBEz5yyAH2LG0TkIsqujYmcp13yUecQzp3eXappB3k
c6iykm9lE0ujiZy6AZwXHm1mML5rpJXfgLAeGGxVmQq9tzgRjlzrzY94HDR7nO87K8uNqZDG7LvD
kV8n2a2wYAKLdy9dDgwOhXYDCB52otsSmwxCF+wbTsSzdMe9QfAbe5mtSb6C8xIfriJyW9L0FJVi
hKfzoSnCfGH8Y3nWliVoOSOgRrR5IhUivNhv24nq0dhVUO5fEtmehoe5hUSa30Obrk0WOwiNZGVf
ryFaBeXzMDvA+Li3xxUW+EAyhw/Ug12tNhbQfb/N2rs+DQnezqUmxwiUXxRwDajbIaONCxq/FCzy
N0aTHkDU0emfLfyKC50NMB/i/bMLHpveCuhe8GOcjkAtpn7VIMhVhoGqvob3RG1xNjEgzx6OaEJz
db7rPNpLbl0v0e7FVSp6YYvR6C/0UbtXaPOy5eVNFpa2I1JhiQIjhBiZCQrpJWizBH1IXLahN1TJ
yTmzr04Pt+OVccINnFX/Dl874rskGCSoJZE+Hf8zI2mEt5SVz38Os+uW9fEmQQpc4mkswTmV3gL/
ey1AQ6S8SSz7MxjTfbMsbFFt14JuJ4IN3lZqzt5svBbo6eX6IEFIBvhIBRCXm7dDqdDNrsSNx6FA
XNcMg1qUmR+C3S7ATrz7yed/4NaxGyt1rS0wfK2Ro/etonyIfLp5/11mN8ajV9k4Nd7wUmSUg9KD
AebhcT+2Ed2fSHqkcaBXwmTFs+OgPkgWNntc9+eYcDON+3u3HsiU0fP3okSWM+3cqFFV+EJs1OQh
Yk2XSaguJf6P7BB4HaT1cBCXdEJ+R2Vr5ChaTs5St5ytMwyCTPf7SB+0Ndlr+gGjnB02uBAMGvFH
9O4bl5Va5Tb04o2QN8QWEu/nQ5aY/XzdKb7D4r8UzEVZx4ZvoOveAPFMwKTVeqk9IdL+hDdQQCWU
zjTiaQO8ZNBtH7HH2rvXAW4lVJg0Q4zB56xEFtvmcfi6IprcpM/nArHzmAQN5O5X4VPctNjROboN
7Zl2jy7SW6Q40u2ciHC5pP3Jsb9F+sZvPJJHu6u9B3jQRZFT1W70pVZErsh0bY/FeYsTeBeHqEfa
OwDxQVb8OZvvwvsGBeBi1q6oBSh/Crk6vUpv/kR5TWxkU0CxI9XowPvcUvV5nLrb4x44DqgL7gQq
b20BJeZsjPqIoRyMO2GeQ6hhW/0fJD07smPBDHaG8IbW8aYg9UwOzPF8LzbRbaZzOluizhH/LGms
usSy7LL6et6TIzzV3hk+JSjHPAJOFiv4BD5RItruhKGdhYKwx9LNw6pTZJpr9CuRaDaqX3f2uGVY
0kaqQ1EIdtUicuNumo2pLZz3nmwsRCp1sKddOCui85wLUuXNX9qJwRU1MZJmX9+6E6YdaWg3kWWq
obPCNf7t3kMu2rg2eF1lRCnk/2Twgi1/suQghmD0HdoyzgIoLM1QcQeZ3tuGe+OmJG2LsBXE5Jej
NwWdPYhoemGE8KfVmOYQXp5qudIoQXagvADdj2Tvyun14aMoeFIpol7tPnx4gIEsQZg6NSlQeBUC
0ZJM26k9H6FKSys25ViTuDKwZeIGGTPnSmiB9T1ctdTy3f25EmAuUEmlZMc/praomoctWDVrDkcK
XJNBGaIpI60YsafaY6/bh6pDy0kl7cnhfIdTDpXLQh9uaZ8H7Kthx65ZlZ/1Lq43H7Mjf7jNhlN+
WdairgGtFsmhaR/llvBWUKJsKy0VsitVnml7QXa+ZmpS3l4N//sMAMpwJiOVJUQcPsW5RhzJldvE
Q/6q9A6U+ejsHM3H7rxf1Zr+47NCzpCM+kAsKWlyGoWpQsgPrYttp94B+3I5S+ufQlnntL3AtlR3
fLBi1a3H7OOzCR7EnO/nue1Gf2E6jmkRJj6mdqv88NQiXm944x9I8wcKyWaJJ5ksIlYjJEBLVFll
d1Ww2PURpt+0hnkEQnyeQMonwf3e0HISlGsQGZJyL0gaLAW4nqMPjqO1UuQcwEpIOJxVS964RuOz
G5tbkoDYMybpyGhKYGRjt786EFo3i208aQcYJLhcZV+iXe/5raKme9nLh/GBcuQUZnK3COwrzIO5
Xo9V85Vx3j2nugNs82MIPzr8Bb59+33gZ4QKR4RaLdtvpiUSytXNw7xqWNpNyPxlOleNM7UHRQlP
kkZx3LaKgNd5vG9eI+lo5tEdvG9L+JuX8ZHGFZzez54jJVY30G7vAxNXEgAYC6d6SpesZw6pe0tw
rUy+11oh25MOceudrYHpPA1KUe0hZvezKUfCS7FH2AlUlgH8oCoJKjhN1gRKoQPllioABw/WdnYs
H6+87b4w5RTNNh6xy2lArRF/wHNg2CmxkYov0v+FHZtlTBigV1wLd920DO9sR7Ipu6tfXfhxatj8
H3WaYTHTRf5AwNglzf019gVV28GPxqYdcGd+v1esDZegclrdH0eDBbUjROqCBKy7x38Yr/avXKPL
S73wDt0I2yNH6Q+xsvBHnbpsEO9CRC6rU6AfYknJvw+CHSd5AnqDayRV4fy5Na4VvrjLLaib6lab
LqTho8cKrDS9Y8PI4Fr1uwyo+PKL48MYF7txXV+QjkXbAlCI2Gf8An0aV59cM061ovsTma8dXinW
GxNM2xUlOIE6F6vdqhlBiUHMJBK4AB0x4puWBmY4PeZ8KhV5R3ujvgTYGvGJpteV5pWEgte054si
gEeWiKL4DBz0xmpUQVoTzTq3mLkyP10ef6LQ2pZsDEoyT6VSUHxVMX0s8YXUjmwiQ6zt/JmSbnWA
+XKZblwWOEQyGzpXKV+IrVfTNIjudO200ysmb3whFLHVQipa7GiiUWgSfRFEU3F/ZUPqYB9rR5cN
F61Pk9JU6v6lDGMVFCqsXtYvrGHw0IFS2bqoYS/zEdoiXQZNQK118njuLVS9RGkOjaL6fzAKR1Q1
1Pl5DuoJIDm1nWn6UgQWqrb76hqLfRAvolteQry6eYSoBJ+u21I8/2WbLht08sSHN3I3Jh8c2GL7
FJ3olIdFzCDzB7b27HWJvsjQj8SN09jZOQbIB8sblStfAfQC/u0rSEkRh0N0+d8PFF/ZjT3ajAJI
AOJxvyyRWovea/bche9nCIBfP39pX4ymL6OLk3rRU7yCVG6xhX3Rfe5f5kbi3hSDnHkceiTpWAhe
rr1t8prVLDzpkCQt9z1gj1iQk5cYEABSaJ0ioX/Wa6KWXHxhKzanX5x75/NSQAIEnqMhJlMhjwiz
xZeC4oIivU4aJkhSTfbJMgDw1kJbGs7KnU89jS1XA7swqabQCkwncz1g8VNGgs7EaMHb1DLjV8bk
kw2jtMAyiolcgGCjIOtJj0WM/4itVkCGl7xLeurvSVoFT03mtlSfgPfN6VpMpyRE9jc75BPeFkNN
76Rgp51wDeWwO/9G1VBskPngLWWDlaiZm7ftna9zCNxGKXE7l7Q34Q8g7i2GLph8/Lcc+uRMVpbu
fa2L9E1PHGlwzwmc0l9eDtfAd0WlNmCQR0UzQi6k5YHuuHNWO7ysUU6hiLBhuY3aEYXdMfTVZiQd
MPzOLXBc/gqm7NGvYQrJZFhl16vCunFW3/VZtJYMhC9CJOwpm0Fh+uOAwIjhOxMwCDDJ5gsJoL46
/O02U7Imdgony4uRGC/K8D+ANg/wyrosdOsmFZgZtAIUk+Maz76rNY20o/UXhNePO5ThCGV0Dtn1
mEqK6LHAKrWZgV6yZd1wT8HwYgKSJVVeHy6ViUWQX91GcX8vsdFc6awCYeDBnIQpf5zZijscRln6
SbO6bdz3jcB9eJbTT4GDIz0Ice2JyQAN9aGL/Dzyd3wgyUujUo69tRXi2K8+YLQaBdtIMjyUZsvX
7V6MvVLBTLGbYzF+tDV2+uGL37h2sUmidgXoQNlWSmJKX7mZt4QE39L/9mC5ydPBrh1xOllLm/ud
tJCC+XKPuzz3EQBe5d3rHVac4VXJC5ePKSAIFSGRSyTmvk9wCk15J46Oni98jwnRAtUg1tMkHqMx
vl2SL3Ov/vjM8bUMGaMZ69jgT3dsGibhpKIRVqYVLcDJjDPQRLQlxn4MExb0CYP2OOCGBVqg3APg
lvb9/7Ffz+37H7fYkvl0Oqt60m0cxI0aa8PARXVPpqUmACKKp5UcpOAlzOgFAf2oHFuzntPvwX75
hli43fPEbUFM2AzhhvLrNm4qh2coimOlR6sgaUi0zPimBNsNysl+nyAdA4iLoQNLC4csKhpNwz8/
q+5wWgKJNGdT5mbCT92ielnm016ebJy4hf5V2SsMTkdP8dBaf6hPkxO5SgLaPoDj4K2BDHhyp75P
gHeV1Ue9pGoWRwZq777oiZjt6qjiNkUjPsZUau8vG6uil/fYSX/Mzh/8o5l2gWu9TSTJMfR5auOx
T1Eigy1xicJMSeLqMj288RCoKHOWdLiurMOMjWqYaLwJ8CVOj+ncMs3SzELCsMhWe0rgINuAWMU8
hRQIYi2GI9GQGuASO8pUICJ0BAHHybtHMm5UoNnKhetQlTIFq/29hbQNK3FOBCoo12zeFiD0xyto
OFWxjDj0NfYOoFt1dH5CuH4YFzCpRfGM5nD0EnStZUYVRZe5hfd6gcPiC4MZnux7YodD7Bml9OCd
Jt2fSyhQa9P16Evwkrhw9rDDNOYK0zWbDz9OzSNIwopLLZ7XSk+UsxL/apqosFlO6TCTqdubFR/S
oDgwvYvoCSEHts8hpKHfA97vthtu56ySOgPG/YYe2WncCQga34pZZydW/x+D/yWJJbJvyLxiylvF
fR6cd9E3j4GVBDy4rqb7rTdvJZD48O5DwTZZutBHk9P2jr3kkUzTLD6xxXx8siWkJ24luy+evgFy
4J1ZZQ/gGo1sQjy/CqJL29RXZic8OW9Eja0mD6ePq0tWYOG0qMVUVfKuf9oNuKDWCfV+ivJG6ivp
ms6ceJj7SZWGCXUECPBHP+OD0QRxzyQe2lvorJFpGxcr+AOZXFe3JStsVtEuu8iP5aQ1UzEMxKCX
2u/sKwgGxD+Z1QTKHsmF8/QsNat003KvtQ+kclcaRjjtkdIN3WM+QUo+tuMebb4P9TVquW6RPvyq
OC5goX8/prVGFF++1MyRduDj2B3IrQrHZBfFRRAEb5YemFr0/VcbupN7pC971AkLozwYqjhd2gHl
TvJ10b+ueJn4XHJSzipe4RUPfUPBDBY8uFAikgbrJni1TGorSVNmEpdolG7tuqyzopbuPh0ldK4k
8SZO/v5bZ/+SrX1BIX2/T4Cv7Pa8kF7qGQi358HvQy3Pr6ugZyz+2t2xySliwBJRylA2d+QTAj2H
9sULoD3SSKOws3YaQDCOSf5DgsiOQghhyEEmevP6jqdWho+UWToYs4ThF80hOABIYDSwf5zYvDej
pPWBwGUbiBtmOdyNiIieJoY3wp9WldmO9GYS6mLnt40/P2ykMLpcV04grHCx+ng3Ww68jmlSf28g
eWu1qKU4tVYV4c5DlR01m7ulLrr2MiAlQfcBQcfiSrdV36CUZ1HQPAPkARbSFCaalr7v96x2+XT0
YL8vmGe+nYPdrsvNh27Ji8Wmg4SWtbGjYvU4vtZVHwjLyMO8HnvliWEQ8vdkJk/xo7kiHXHzqK7O
TOxMx/RojUAcePHFfLF1dJnuNm1hmmRg/B/GN3tnyYpCyT76qEG0nfSAU7N/maRQUmleaCGtQYwu
Xyl6cBPK4iVVqNuSEglZi6xBX/ysE+Wk+IXE8jDGJBJ8WOJ1vAsbH0Gx6NDip5y3nDYWxoSKeg82
p7iLtUlVPxGNTlVedRjiY8b2R1EzIKaueMWI1i4jcUiPtKHns99ufJyc2EdElw/VtU+mj1XzUv7R
BX8YvICLG93y7yIpceu53dWeaKfXcXxKTfVo47nDRLLBu56qrJ/F5CLuEnzHaYiUSfjalsbXvHzp
LQKI+zVRZAbQl46BQ1Rnq02SArQ3VfwzC2K6hlRVsTZv5CQsClvrCPVJefFmTQYHB2V/30j5Vku7
VTMCmeQmQrc7CcccbvJ5rTA51ol6yuseBaHZl2A7mk5aOKGGfSpJ9hksuerxb0a5Ciujx7FJvNP0
BjPgEQ3x+XTsgqXiuBO1cLb72gqm5yba2yy+/Z5XIwA1FNAiSG6CMLIID9IOV+NTXBVYCUzN2c2i
kbQXD4GWlCzdJQmLG1c6nly35ZSxmeX4rPqt4dB0YPV+g1ckUllsjEJr4YZ5YP3AmOlxXMZLZZJA
61eXqNXFB7PbczI+jmFZmu0qCfOsPFh1DjZqtSNHUXh/Y5/KNwONLfIx3pKOo3cea90QdssTtkyk
3TgZ/H5XjPS+bpEnLBYgsczgEL8nM0bUh2VjXngombAqmBRwuLukNigsSjjhIjJ8AdUHC0t+bnKe
kJBfHy/MZPHsV7yy6LhIInIw2pzUp9sgzrFC8deVbbOghS6p3vLU+SsZDjnzpufVgxw8WkHZkzDO
3sQzcj1cKqAfSXjua6vkqCNmCb8YDvUA0Ap3jDKY/SFifbu+65UoSMA+46nJWaJjsDeMKlJmvvso
OuNErV5Oohq0PLf7cX7KT043tE4EfH/wdlCL4Ihpm9H1GBX3GDPKSkjnhxGGT5jf3pLJxqpb9v/n
DKuR1eh9ubOwrhoUm5QiZla+NJsuiuWjYxCyvOPLUSv31wjxKekzKIhKLPqcQS+x8QETasXzLfzp
dtv4zEwzTvCvEyj9ouTSxy6CuzeKBAkRvsNUiR9ugsSU0NBHN3/4Gw3rXhsI6DX/JX/gX5g5fEKP
S8DGtjcYkxL0QpojlaMR/EWC5aI1eLohywzLAK/PcvD2l/vNtF/9DVYnqxfj2LDeHXBbRujxR+Z/
d+w6n5zBsY3q+dr+3D7h18Tw0OBWF+hw47CzCH/zXN6T6RUr4zDu+IIc1djQ2fdRp19rO7VKA1nG
eOau0EDQNLkl0Baz4+H0NMlCgpIto7Rvs7DzugGjrtikB1Cv0/zAtzkv09ZdYPrF/2r1icLnJ0cW
ctggT+EovQ+Q/q8Md5YNljVONvt6ejz7Dh71Hfkvj+7ytgreM/Tv3SJHArHypfiJjnKg6jkzPuEi
pry3EfdXBZ7z5oIWmXQjfr6UaXPtM9fkaVzVtDrG6HXjGR5YRZg6RJ6IHQDV4n8Ck7b1y52u0/N5
yzH/JDa2j7xktDrO+yPC3jDqoHxdeK+MgBxgP6FBp8z13LeY8dHbM722ok67yidwSzjimRfdp2Kb
Vo6ftpjqqt6YeOf4FgdGIj0AOrde/0Gq40iOUxoJIQOBvprNIbLdZmgXko2ukfLScJs9lvMxYPpV
v6P5npbpK8mK1JSp+cmrPTNo8zZ2WZMFkXDswDoozX1/nHPDQkUDPfwQ2+nKyyxwc0qL4FnrkM3c
hYelF5gAUeip7rSPbj4scas1bGixlCqkIzmgZUapbWk0qoGvW0PhKxCZTV6bUGLhOBmT0PI2wS/x
RxyZ+vZfpC0l3vswMJ5t51vGWp7IKaUssif5rEFgQuyzie1TMjPVQrgPZXIA51z/hbkj1VWbOdbK
/75uY/IQiRv4EUKP50INqslVFDF/8BXQI81sdfvngRCV5ZgqWbPBjAHHkvGNAjTT0GdOAp573dlt
dqIOf1r/x9+IkQDRcUFktXV0vowAlkquhkuEKacI2vYC65CDK4OSh/FNH795i3K45pt5V+pNqNhb
205GBOfa8nJeoWiqrhp23CPNWvEY++IR+FKDuP7KRu/YYPu5TOLkb44k8cbg5/ZIo1IM6D3/Lmct
x4PsFUQ1NiCY928t/cOJJEGh5oH9waze0nFXQ0Fyd4JlSDfXw+i8hKui6+/CXVXDkp60lgl600F0
pGE8IoTi7j5dFt2j5rziCsaka6e2Rxd+85qYfVzHy6wywr7rHba3nVo24FTI0adMHNZCuIOMIx7U
etWo3h23Kv7uzMdkJnb/zDOU8OJSZlOw31vJ0ebpX6fCgcaAJOdL+aIhg4eyGeCC2iKw6mpY8rpr
1mi5Q/2sftXLC9h1oa3Dwlxe48XPJ05P50LZPuXOzYlSjMaiSVYj+rr3rKyEdg5xWDYsYiesSGDO
gx1mneA00yzmsSPLBRjtrOwBvbMtEFVEJ453KHJx5YBZkFdCPm+k17WkYqJLaQRQtihkmEG+I3aB
HqwKVavkoInKd05Z5vpPl9oQTHHQYz4/4NHJUR/hUI5/g+bm6eHIaALwC4y0/BU67Cc2X7AhVN3W
TS0npqtgTHEZ0uGXxH3CrJOEG0UnCzU82DPQ+683RwUYYf2Ta9BS03IX1kPoY1vy2DSYUV0/8jwC
L9y64hIu5KmCe/HiO/QIuGtYQep8XyRnpijWlSgvH93bEcUeT5+XL6nEQB+pXssUuauAl4TEV9l5
J2iM9CZEErCkW6vQOrkgu6NROPIB+tcCCl7O2VQ63OvUfZPkXinFa07FCGVTnOkbHLKpy8AN1PPe
kWxrmZnErOj5NLPMY9DmjbPvj58dYxeYyB71mTl4UbYfocB63jqorlT+Snop2rkzkJhwY+TH0Xgm
NRM0yzlIZsadtucNMAWdrM588+M/I9rNsk7sOXB9CM3+MwMRHdyTQdJ2e5NUI9pSjPf39UlrBdKf
6tmonMwM/yWG+F/HC2DGp9Im21KL2D3ulsRKG5XyMa6OWOr3Y7nhmprVUuas7PnBmVk/gFmH2rLA
Njxv+xVUtil8EeOTl5lEzfmNhWntNNcxHRXKqhYX2d4JK5rTdFZ5QU3W8SFdGhMEDI4S9zyQAzf1
WgZFvbw8MrfneMddeCM+98PvAMMEcRornzTC2fDhwafMTMAYrjJKFx+I56IM4LWJYBtpFSxOme1z
p85JaSTdJQr3W4v4fhdGdmNG4SWPE9BK6wYMbwW1zxsssajK0cqLfzsA0csco4WpaJEmOajDE+bX
50Bb3+GwTK3p2zJ2yRyaijjXBoHBvpq/AyJjUdCrb6TTYBRs8c4y7Xl1/f906hRKQZbdprAFUUcX
D5vZRBJICYcxZbNZ/L/awzYQZun6nmxNWlEX6zl8hIwUBvOiKj39qEhNxydxEObAyFGJBaUR2Aln
eXSS+0E3WDaWq98WJTTXYMTkod4GkrwwzRuGwJEnc9xxG4BdM9AYiEVdHUHq2o9PPencAggyAnwP
lAckLWdwgoxZEG8XLEkqIE23fjvFSr5/mF9TPx+SOtosb+R0qEy/CQ9+FHMVvo3bRpp2g+SRD0rc
LpkKtRLYufXftPfPt8ycCevvY40ogSeYjTVEIXUbq4T94hA18pEy0wjGHJC52eZrRM5lXVcg+0nY
j0wKKZEDoM02/XZQKSbw3qtgbBs7lJbGxRCCuSx8TOTpnt3sTZertVYI1Awu0VBjmagF6fGiPSfC
STOnEA43AUYp/gbm5bGvqbaOKO3e/ZsHVI4DK8kOFlxIwpPI2TKI1ANxYj+rPsTJSv15Y/S/AR8+
j8gxPfVOM9V7hwNkTj0ZeNvki3sSaAynd9RRRBtp59bBnbJNP84i4okPz6vlIewuekZWCA4eRpZb
+pZgxPFlemmwPlL5Gto/wEUjh2ckMi58ro2KknzLYAw1f5q7TpqJ2KCJ5DqwteRRofQHRkp/xwuV
5I7Tn9QY81aQhKJfDbRpkUWLyw6kWiwA02qSPycB+dbBGcUssp0mi1YeiKBvNMxTsiZ5xqli5GJe
bJJWzcJl1lbAJZGU4KJ4YszAYEIw3nFdhqURNDmEtFMpHLTM6aLV10kly/CpIm5DrU7/SEZiV/ze
U5KPEpsub28GGoc3fT/bvIBbIKXkl/J07Hw/WhG2VpcAF+f7TJAVq8ZZEUqnqq5odtPuLFCKmn78
yI1DwRkVXtSKMCO23iWWGhC6/f4onq+A1W3xKWGBW+Pml6kPlouQ8WSEhA5nnoQg2HTvm+HrqUQd
2fWgnocajgdFh3L1ziU9Ek55Dt9oWRKHJlT4FyFGWZw3ZhPXuVeEJEWv6emyM2BKyiLFIglBPR1r
/rEIF4ElphYaYmRw7ZWNE2/CsLbMP5DAJiXQf6kwQ2icRz91EM4v1042P9iMho6tPKwHYom0MX27
5VN4qzLRqXZq1TusyvYdugBqbfj1YzeEYCXaCGVOmvWpPcSQHOUctz+91k97FF3uziyl+8K2d9Ti
9sAlTlIL0DXFaylYwRqCimDKkrh4XH8d2krWi2vWSx5SUBm7uj7WT0H++G2utZPatsJR1nvvwLk+
yyWN6OagDTDNdlHYDwnzE8bvEa1RcMMqMSY0zvN5INEACtRMzAO5++VrcKwWnKEyOH6xPscvbRaU
SNWv52+NFAno+9sQqocHuFIRylucbJNxMxmrIYQOeG+C4dStvtfQatk+Sn3TGVQqauXCapyWqpPk
tUllV3ZAVsNdRBVa9KP83IkE9moRFviGRgFwm0gJcDqO6aYWiWM9gCkKrEffce7D/AYcsrag9p/D
wszHHRyoUaFc2VuyY1pcee4vtA9r84V3jWk7vTMQhT5HgQa77yn9+NX2B7FTZeZtnHRPFC0dSthe
z7T1yisxDYHZThybWQf491B98Vs42EWv3HoIB8EVDScia3JF2jWiHB7zTbb2BGao7cDFaKVhGUe2
i01Ya5nIZU1JwvAhAuTYaFirqDEB8QRA1MeA65rYhnbCQMQrcaQhfJffpVGDBCPnyV5pjmbq81Xf
Ns/MiAuMBoRxnVueODeGLoK5GmLXT5sE6pXbK9GM4d+LwFWvRpIn6CNQ9rQVbh+/TF2bwWkAmOYw
1+5wGFQHXo0iA4xVC9UaZIzNZJxHZmuxE02Rpr1OWwAL+c9+n5IjvbqgyzDpFQsCyAkGSI6+b665
KzOF80Ur+6afMYLfwOgudrwobDxbbBVEzJVN/7JoqIJ6y53bgd7XuZFTZrF3l2mvMDgtJ0jXfOtA
1uEsNLQtLEeyHjY9EYR5JEJBL+qinQzV3haQxVYz1L5PNMhSLh58lRFzavg/0NKhxnHChdY9weAj
hF9EigtKujGd79vBNFSHei5YIiGuk7u0/e0KTglX/SY3qm87MHFoAUCdywqeTv72cY4YZMpqGCaL
N6gYUfIDJoPgo1Qe4vP62tbWl6+Gp7kZFtbcgiLP/hX78EDL0767j0wdx7jiP4XYsTrHsve72bhX
mQt5UxSWM0R1UpTVQdciJJhsy5ZdS+2cc+TYG+4pk+5EmX4AWfLWP39O30fV2qHawMm7c+Qcu/rf
UWwH1YP5+Hsv/nxGGfFfE3KT3T3L3gxI1M8d067pMwqDUx05u/wQwcd5RZ+WB5tj3jzMLJ5pDzQF
vh5+xjtny3gpxFKzMwfNlr2zveOAN6Apk2FPru8lpjKMQg358eiFacdX80NwSQX0cWNmKO5tUMqD
atavI8GbIE6O/iVDkUDf7k4z0b1GJ6nxVGJVPH+HZD145j8WdNl7vdZCy0fhGr7rnheSUUL6/xLY
LGhgMf2qU8wCzJs+iutFsW4r2BCoBTM9uW2j3oDxRV7BuyrGkyGp3pSFw69nVqNrURRM3CCIqCj5
YcIup6M7dAjVn8kE8bH3+konpa538dr3+s0GlBRW+PqwULBRkkf6goZyUqVhhSUMCpPP8zG6WvkE
HEKPbfyVZaP0le0Z2J6iECIdRYEhG1Mj9gnzyf9er+tLmAPmE7I/PM5VxRQkzjDkq5wp00uFAW7s
jcJIJRrCwlgfjBoYocdCkqddBlCzcycEoE92Ro2jhLaLhqsj5SKl+86ump8SluXtXrWSPlY67pt0
swhJOImg9IKWWAmpt5Rui+9xymPyGausiCHXWjYPZgIdD5+xDcZgOHbrvH+BFEKZ2pPkZbcU2KuE
ikFf7c7Qy2OIWn53kcw7NEFvvWajKxmju2IDZZYfFkgWeqbzd1BIXYftVLA3N335KsTIQe0ttuNI
d0n7Hlq5Gc0Lw8nAY2gU3zcWBL4Mn5gPMo8Aag8hYEsCAcYx2Huop/VM9YauCsiNA9jBD6mZnwl3
1KgS5ryVfxWUYOgTjrB3Nm2pCFwJyNAaF4RhTaYub4RwYky9d3MYfuAwzdYvXcvtBrmpAOjW1blV
IvpnkVyLhUTTMXHdMPYGN05Xgl86Re4XCXsjrh3VXFmDFFm04gt2x2XeBnjloxuUOtRdsHaUqypo
eZI+k+XooYBDsKfNYyiBPpD7vWKAMhulcblnsxIBOXBHhz9cFAfshPMypIw99QjYNJkfe6NB9T+z
W73NrGrNqWzkibH0cnGzK/Q/L5ebSDP/1Y9XF2Cb9PX2a/fEW7c6JFOAfdgWq6hPKdOLJhCfGOnH
cFjpDmtQ2yO1bLng0a93EwOGeCzdOBhiKu1YkTprYNhK9sHq0BtV9mXfkTVt1G4oMlgRPFJ0aXBC
hGwGa+5/RIYv/T3nw7cojUfMKb0F6RjUMi8BVgmBEH/mRSXNMbNSVUVUC2d6aqXQOhemDfuDADge
K26p6QLygAxxssrus5XmU8nNWLfrnD3xHLMitWHsU4iu40tDZMQoCpg60n15P4Pny973gtZTEvRI
moKXWSdKPZzaMgUUkK+1qdTVmFadOilYfNe0KPir+IW6xSr9y361KqgBwXom2uqgvR/qSttaxwos
RDM9TY9z6jnArFB9bltyFdchSzl9qzLGDlRPekXD/43I3GZaP3v8KMi4VkbuSLWzAWzdeXgElcvB
q29YcDi/uO8HoxyoHEIcBMmPUaWuI/dZ9WE3fF9wgI2MLYVi1HY7k7+6RuBWTc3zVlG8MI87BZEu
cs3AnpSp3vusGCsyuqf8G8ebGuhBk2QuRS7m/GdWCrAVjOzy5dT/NYXrsddHMuTZX2ozOjJd7njv
gwqdPre7KdnP2NHTWstDZaL2UU9N8Vyu3K6TFNjN9KO0+Hxc8ZmPhEWP8VD9cO1EM/w+Og89Kyjs
LChmzDQ2hHDalJqWcL7DTC9Cc8ZOwGI3hUoDT8imgbaDHC4gll2jitK78//Ov6kFHc+8ClvTfxB3
pXLxB4XNEM1QsxDLjX2HhbzH5bDG1x9LeORju23hOBTfZiOD579/tz5dlz1H/l7vE/evLgPDUM/o
T5Idydn6e6fB18CdXZ8ly5R4L4olg6rYcowFjnzpADDdtD4FcYxBH1snWGWcO/EKnlZYY9rJX+c4
GFPX66S+cEQJNJEm1g0hG+QXEyNiir4tSq6QNb8WiLclYeHbe3NY7NY3FoScUzGtFrckyOtph5/d
XaQL/NmTP1iyjVClqhLq85TTqn4cdRfHLVJZu4SUtdIq1BqhCWIwmIOfvWA44BtDCdI/NbTLGWg+
4MQADog99Ieg6J/dIrrAZit12axQkwRzc1AINdX1xuDGeSpb7CfLw0fEBDhs8SPWlqiMgKNdC8Up
WqkO2rfXuA5AFHVhzjjlpEK06XJ7CbVQsAoOTEPn3XJwwUttdV+rdFamOgc/6mGP2SSNOROQqK+d
9jJLsHc0ZbO/1mJHd8UAIElLcA+c6r5jYuFm9Vic5bL8MJWCOImkG2yOIX16uOjgZt5PvK2YS5O+
HsJNCvqZlA95Y+pi2/tM6cz/g/7xvlV1uOfUR9R1A/1ArytVAeJ2gHFiTjxpUplVQ3MmBr3Gohkh
o5aoB3ayVv/ZOmGckikQWHCKjs/GnDSKKo2Llq3XyrwYkNUZDrMnNTIuROlnvhjrMakuNg+PsVMo
jEcrIvl2VDeZnlKiW7GdPfLLVGPwOKdOuvKQ2E6YdinPq5punVWE9oB2ROTrN41el2vFHOKftB7L
pbeyzMNL0l2wWLKuwTt3P2PUI1EWgJsUwIapdPsHcpvhueBoGqQr7Mg++HechgzuZuqoGFYiBjgS
0PK91VIIQ6p5ZYLStSFDYIjdxdSni2dNZq7p9DrorsQy1Ax1l9Mk23bHSow80vfKRo2E6/C5ffRG
OKBLZSDbQ+VFZ8wWOMUDNUsnl2+HZFlalq3CJDMjecWZOsxTE8pddLmJ0z1N0T498YCUHdUtR4NJ
G5IOg0rJX+38YnAGkzZlkHl1G8xOQq8MfPrX3aPDS0c4QPqQjxNN+oFU180PMWnI4AHWHeUcokSH
zCDIen4PMJaXvfDxGIfZjQd05g1MzMWehMcwIWVKmg93q7QfUrVIU6BdGqV5Fv4e8o8E64Yotk3r
uRA/okQ1bCsHfisTlJnmxI3eC63wacM18EVgIhMtj8l3Gx9EzK7hJ3jilLYgg8u9cpPFCksNT+nv
7AKiyea/ho8RI4Q2RbFhEOYcc8DcMdF0+1g8nxZD+/rz3P8dSZfPwSpIMoknPix+df8V6kA2E3DF
v6V0N7MNBMr3FfZvkQxRcBbVdXXvKnRAjDLM7Lf6ydcGmU5BuCZEG7tng+okIYiqmPK6WAb6VW33
JN6rJDHOrrlifBYDerwOgRpTYFFf4K1QXFMcHfAXCxXkH7K34Fv0BoNeZXXLhlvtBp8yGXDRzULR
e87WUC7976EPAd8nNIinuS4n45mrogWNv7p3MCLFts7gWQmUph0r20nYOgxUSx7bBHA/LTepX7W5
pQKM2dRL2UPUt2ZSh1EfbEovhFXBDX1SokjewxuRKKAvgw+F9AbquAv59gtEGDjclj7U7WWqrRpE
CMx8cjMRqHGq8PFgKC8NkSXb3r6VAdu1eu7AjPNRERYj4fBiNGJYCX34eT4MAYzAM4fC3fUFGcDD
OHZ1dKvBsv+XMEVm4u2mYupjwPH6/tLKXeneFnNpjHDZM54LUJQV21XYKfpbUFx3Dv7/XTmoyMka
FmVYhxtMZKSTjNE6WGLJmP5Y/okboHNVNu14KDOWiJD9apwV1sXmSvHEyWAJ/ENFy8RPMwU01/0g
7uSFNMQXthyMsjBAIUYhXXRUabQhks75++7NSPkjHOYVZL6hefz0PFcUjBsfzzG8B3d6T7pwz8N3
DOODOfSJvblBLO6vvqHx8vQPeYkZjk2HRXSGuy8v3LCussx20C8Oj76BR6m3lOkUHacy35HPPxKr
OlodCluQlrYfqHyCgYmzROH8sj8IX+3ny1kubo6zD/S6QkYldLJsphaOT04KjfDCQuBjUB0cXDkc
tF5mtzEJjyc+GYmgKWYFXEo60xrt5QpTilddf/FcCirHv0jTQYx/P+gFcRTPkJSTIpet4A096k05
AwSAKlLxovkm6roNID5fwqSkeNxW/8VQmMV8KBIqFzQwkYvAggqOBaJB4w5H6HVt9h/a9FDBzXGB
jEh8HQc6FNT4C/PAS0bPFri2DEC3WT5zJ+RqzwSoMR4gVeIvFk7GYn8cBnv/y3XXavMzzyG6dnII
htVGwogOw0ES0FB8CZfS/ev5Ah0La7l70MzsE7YXTTlGwKWVi+W/MJxuzKrkL3ql03ZmRH2CnqD/
3e1sJw2VjYQEEz5l/qRHMwbnfRKN9tGkQurisKzq7SRa62GKtuLlJcNaRH8r08Zkl0OxC+bx98gv
mkLpwtC1U2v8LS6dRogx1fqHfSxKpZJ4WAzcZnEyBAF2Oes56Ve7bgZ4Ldl/uI7EN0Ebn6NF/QuQ
Fnnpm35mkJQK6xdjMcEvTWBaZ/BAgSe+jq1SK4bUhtAe7ToHmv+cPCSLRdWJJlLwsGFjIFH30uzz
DPdePdHQCxmr8Tkm45nPK0+ZP8jm3rr3G9gLDawaGrAal7USdGNCQtTzmc2eT4zpdLd4b3w/hY3/
SWuYZo4pINDCVcs4m/YCwi9QvphFyCYzEIk2nsXXmWY7cfGEO8JnhUATEaJ5riRUDNhOeGet22i5
95JB+Msv2F61gQKp8p4l3YeoThu7L54l1knYATQ6uLbrF+IPbTHLp1nRuO9HT8VYJ715RWoeduKQ
fDYLEblweSNUlRzwWK0ImTDiKutz3GO0he7vlTAMSUyD3rIeJ2X3hYq9xcrZcfiASGK7kT+TTx3U
rD6tKigG/M2LUO58DJ7rLrRYFHuuzfT3Qp40h9O9IxUTirAPVd2JAtrdGR1gNUWuNAYmrnuDRSWV
f5sXHDgCGxOqLRJfqcly2pKtVL3EctAlwKbM/YSkHlbWrSCFrvz3Lh/5QA+1nkdb4BRJywVFbYPX
jlbD0D0dltkSGfp3FnQb0oPm8jeGX392Zh9ts8Vut9TreOLqmwrz8I5LXEHDZHnSna+mANIwBjfI
Qi3GQtfEC4KnvRpJK2qMUkXr135RBJPRvnxO1S9pvmjCnk7tJDr9zaig+CKGlpjIrGKrdkfaQ1oB
ckq16oRw1w6u505GrmX7vX8TzGkfW0wRZkhnMcaIk53dsEtJIKp+ODWTx1XIM3wSWnnw/Jq9arh1
ZXE0sn6rIO6eiqWKq4LVZC9NMOZEhuG7HAmatqRkQTp65Hhy5/o9bLNXDheBteS2DuEiKw9xEx+P
dLnatA2M7J2B4LMrXRhWzxo9Jb2P8HYlVThuKaho3t6UjeFz5LL7XwtXMiD2DssMBMu/wSJuoMnX
bbmfKfGMYjVsQF+MIKAS9ppqBqfJZPaYd37+YYTAE0MNf0fFRQaenkUn3SEY+Nyxsvn0Q5RD+Jgo
F/QzqttVAvdfnkIVuv7FCtKHIpHKG1ykME2E763fvXnaAKwQ9ny6uwLG3V0kp0VknmJYhMCXkD00
eISKIEEuOu0R1l4DjBhL/wPy+gBxyQiz9mRbsOsIAQevzAmx+cnQZU/GXFGo73lRH8YwAM6BQgOb
HBG8nwyBMj/QyIrPALrtnunRIP42yR1SWFuguvunj+ou/NQqJJwCmlmH1PS1nGwsvVIjQAmZBn0O
XGPogiNoNZSdEs4XA1G/xWTA9NVbLKYQ3bq3HASt7+LVIMlY0iP3sXo4u3tjkSHNkfppN0d57pvQ
93465z0IAC7HSafYAj/K7uXdzqzo+cUOpCkO7tghMAKqwUL61ZfcdyVMk1Orw1sApn53D2ZcnRRg
EGuL9CT12xetdL5+eTCHMi0NAYVCamWNZqruYz0x3z5z5e9Uf6GkbZSfqklgjAS4JZCv+td6wtXA
X15HsmMChBQHANBE9FDsoflaHZdqcNSbLKfV6xyItJPilGDng2sMo5Qu12I0Uy9bgDSTdkYpcMEU
nZ5SSFheKgLE8eoXKbDZX7IQdpXbrnJY6KIG5xd0EmJXGMtIKm3UkcLOdvdmmu7IrfNzR79ancxP
+zfmyAZJbiUHenySOFJtdjAQCfr9GKn8Ls1AuA/9sgP4eG561dQ1P8dACffeKyd20WGkPwfTKb4O
FKwmMsD1UU34i8K52WBVKyyS5YM6/RkrpejlCgDnUHFXPT6NvAbL4s1sj89aH1zfqCWw/O8DilTr
R2ET5FmvjU4LFWAQ7IzUSIFYBVx+A9HTFQVkULzaZ/1jD+g6gP45ID+817P8tk0PWCVb7frcSmPB
BwMpL1KDT6jJAR6oca0BhUnnmaAsFPhdCh3W10Z/PfLkitgrrxYWSgBW0gy3kmPzrCJQwcRn5mx5
KoUWffV++8DYwetMWwgTeRJxAsK1NXyA9lfFuKNhbEjyA67QLJ9Vc3ImIREIhC8pfVIEIm9V6rGU
vtW5+eOstrzKEBlEPkKlO6yh8ED7qhHgvFOQPBKj8e2UY2wZJgHsjh1iYmCl+zpHHfh7upgabTCS
K1+x1PSbiiKkR+hSVCS+3sVx7+td75CuqOLr77XLMlTtL2wlBqYJRatjacS0WCESepPm85UcjPcS
Ft0dV73o9tRr/lGJ7stazwyArnjy/12Vyh2rNUFucWMwmhllto5QJD+WRBh6d6vIgTLvrqH30xts
MmD1wixiR5FPFNHqot6wpdqGr9uMTXTaR9trKHn61sU4/E6M60FQMeipuk3XMLiujNitLBauxlEb
OHBQH6U8lezhS+zYn3thGNFjYIJb6FU6TQjxgoiArAVsmwKdM2unFqmpOU9Q21WUaY7VQHww0rj5
/cWPm+5gRWPmIH/g4HNzfy/o0lB8197YBLJHAXnB8cfDEQLs+gmeRhw/5NE7EmDdRxsTzF8wpmWi
QjCwflT5ITtZOqREOSrErsdd1Dj0Esqe3k7IcXOdGl9E/gDIZy1oqUTyPBAfSJH+xZ4tovPpiP+n
AIC2/Dph80PrWKNWr439uO3xMPyN8bi/e5f4bO0EFGEkzjXaQZqfP1zHPDvCMphhE80J5PP+iw9I
RZjOQn3NckhNB9v63h92EbJZNirv4hpyzIkk9CCrV4Pck9nZ0EouM0VFxo24kb1DFLk7WiZ+HVpT
llX8yuAxNDidYTb/YUcOr4NXZNTIZJdxGIsQw23e2jrOAfubwusVLs9dQ2mP6WJzKnEuhtZ/k/P/
jRNVOOPxb8J5BiY8TJGIg8QmocT4StjPwqHkY/LLbqiB1qOUqtxs0Mf9EEZa4NfK0juADMpJicv3
Q+e0hZZlk1fxSweYeeiVOE7Y9RoRatuwner4vWRovxMl26QqY4ejeEFwpvWTKho2y3V4nLDt9QgR
XY4pyVT1d1zu6Y5fIpQoeAOvFDsG7Iyoi/Rr3rgWSCmZB8y+LnXbrH4ETSeDXagPtGrx1DTB8MYA
Bl05SrcJhQCaULx49Y0xfDCjmuL7/szVExGBcvO5iqkFMvr1nbJY0t0NwajW2p8xvb/d9VKMYt2s
utOcgDvDUJZxirhslHUDoGgbVV5rXYuRnKudr7xsxrsEj+eVDOe1rpMpOtsZqOV5pBgPYc3jIhky
kMxX1UTRLjkTPo65YlFTdlka/qbCggAoEDe3aAwJRcR17x2BJCuviQdMOERl4Nm7DnNca8WSpgT/
hGgxaS0OuP43bibHMxxV29gAKifVRZ7tgQLUxLiWo16mDmhE0Pic1RG3zBabY/D4dns6IGRKHqyf
9S76Cw7eOAUX/vHZ+b421q9m4/5wp7+isr35os8uFYY9mwsFItYiaazCGKm87akl1Q9L7yPhfRg2
9/CCPgZcZBVRDgPxXqzgJ4ZjhGGq6H00FYdBiA3UEAoOJiuO+Zy4hqLyFcGZX3t+nes0uiZ+0EnE
T8iVHg1s9Ha/hkcGpF7PZ34+OEd2TBlwj020NsZJofNtUL4mUPmrsDmZAVVHc6Rxdpp4K55jS2I5
17HdudR7WLgoCNHsSzezNKGVYQ1Jkz2eRpvpJMdMG/zqizUlz7lRsY4gTDDw0P0vVZzNP52yIe9X
k5CQ3v0c19e26onCmYll0JVQLmcgnYNK6gnE/hEx3Ds4Mc4Nd6dhm/ekeyzmcEhxlnSsRy96vaWu
aOq6qrGu79N+VBeFwODLuDlWTXO4oqKK5p50oqo25vv4sxOXfVXWi8HOxuYUSz4YQaaPk/bbLDhP
dIA2QQMs5HrPIbs+X3eI0Sdp6d0hG4sJgKqQ57Feut55AbURzsHS9LQciTD78lfVmxNiZqEvreOy
QtEnUd3Jpq6aET0sZIoWKzXLzNskrW2LDZYWpV+B5kR9zjespn+k7ZXfjJkSGcdEzqU5Jlve42hf
odK+vqiXQg3md/M3kxUqt4ahAYR1oHSWzB0heAVVcd5z8wUVw8xUGJTNswsKbvnswA8v6nk+ouFb
dUVsLn7M3Numiqj+NZ4gjfZs12DwW8bsHej1Uln0n7LweO54ND3iavMn3jOTgUJ7NXyXwmRydMqq
yabEmRuiEOVYVYG0n6utfx9qAMD2hfvjzalg8zB1RPNlaYToQungI+1P9KUaXQNwpv4biWErsMA1
G+ERHPFctmIAKoWXzrcjI4LeSqBtbfJwvSFuq9+32TUe7dlSnb+HdT8v8t/90jLxgwarTVELgtil
PIQZ131blFnoIYdBEtB81rVAmjltHJDXcay/KwbNYPbiJzRRKQ+0fnj/8zdTc6mHHfDj1Bwf2CPY
gpKsydSjnaF7sISjML+2BzMvjH8BcciQ6YNQkAmgB0+L2IFKZ1m2mCFgAWA6mKskH/RZ+FcAeAGR
e1nZ+2m+Q5G5HxhbWx2L/hyWrLp6+3AG+Yc51ffm/ZeX7nrTtGiYmUNg+jHU4iRHtO91T3ZFLjJa
kkTvOHi4vGcGaUGCURlxNFeKqySD3JEQHmHNR0qLoun37uAR5ZUgJgc2kr1kZizscEKzh7vvZOeT
EEAsifNBfkhlX6mPKfSlpzb3PS5Su/JqN/iTYhQ4cR7qa/CQYkqAR3OgwO1205ZgN5O4I0u1SVbX
y8gl0ToFuG+vgLmorf+2/eDg6S9BPf1+bsARKBSuqv4lA3/ANpccUTa+BY+WKVi1SCzMgODl57CA
u4HGkr4fwdWv//MPbpkgJxer7Lwb81FLb96s0mV5DAgPi2y9ELY73ciVgrwuXZa8S/lMjnOtBBF7
HNW6+GmA9SDw4BoACxKK7EazSz0VpVFtRvEhlklDkbG0oE3s1nHA4p5JsKKb01kYorqJKh5aezjP
UIRM7QkNkxH9rrSdHlAw0Hv1rPFmVMczBoAgJDvlM7ZuzqLpggKkhnrrXVEQi8uh6Qb1+YEIclfa
sK4Fvxk91OBS6heqQ7ANSALUv9lg9SjkrtgKtJl6jMKEjmU8emrzAA0Ff1fV+ezqXQPmK0rlaWsd
ChgP7OFTR8gh8gHvbtJQfOHMjn5eeFJca2xYNl0+GiGs2rwZQRk68EGoHOF4JVySkmLVA6foxmUi
f0fzPPCx+PxmbndAQtP3JGh276xn85/ZZ2UKLWnB1mLFaRwI0bqLXLJjts+gPvscXHMcOVQqArqR
dVnCkni/R+PiTwFU/+uIxG32WqTvLGe1tCSc6Fakv6G3XaBswqZkC9rZz7sEvEvF/8yKa2pOjALa
zQuXouK1VXLei4Ykje9mwQKkKXbFL3K4A2Gd7R7UyQ/6v+lFZgimfYHQDQQ35oF/fnJvuyERSfcA
QqkEfNwXj4As7yYESisEFZJLxdY7cqDE/nZfnJRnVc7TKiHnFce5I+42QOlQ4LqjTg7qhqse88y1
/Bnvl7EVP5tMM95Poz4wArTqVVOK3pg/GrM5k0/157ywD5mwHR1+7cUsJRipbkU8FSBayfxVKYq1
tlgHlwuZ1XmEl7USa/oA4ld2AIvV+nsfvOiJXPa8+hfbamSXUiuwjRx2Oqo5vgJ2L3nNRRlxrXzp
YpzKiUcYhZBSGg2/qfG1NR6XOEJVGpRdE2Yds5kO8z/KRDjAUaF3y1B0f2z2Qf1nsqY0jFUJrG/O
grsy7I/jBb8othc+ZOKpUZ9G7IMn75kgIHnKeIGpPrm3ObGv4ZWFHT91I2bKWduRXh41PuLMvito
qMn14hPoNnuZIBBz23Eux9d8kHNATwtPMhfBxthzrUTBPsYk8OYWZylXJb11rJuBR2IOmhq/qtWG
i5neB3Z/YxjOO6AvY/If315XbM4nkGdcNubINfmJ4eGad/yizqAGp/rIxfuSPFpzaiXDLAmJgYpV
Zsuqla7R0D1GnzsNI/It2KpT0W1CZ1t74AzPZbFqwYBsJ7+4uyrYN8BD0iWjSNMoJmpGkqksazLg
M53rPMR2mksbZuC5ILudKsvkiDcQY8Cm93YiAikdqhyb6xIWbUMXCBeJ5X91ukHLgP7nFU7kBk0C
7ZYX8F4XhJC6YwU6OFm74T+na1XhE/yFa14y0NSa3jDdwhOOD7dAwEQ4rPDhM3Qkl44zU509WqID
8gNne+lkLA48p8fr+PbOzTUjPqLCRVqLVe8KviBuV/nMcVRC7dx6Xn+c9k6Ne3yrCNpXi6ZjhEE9
15cAz/tC3Wu+EOBtj/G2ZFDwr6VAkliQeIJGn+3zc3RHW1YpUqO0BVWnEZv1KDQgeCiHlqEBeFgI
Dcrem6fKpqIS3iXqyiGH3S7yfIHYqh4YK5W30iVtrU0b45DEy0m3NSke1U02h2GdhcN+aejBnP/o
J6jwEbX9NPM2/hV+DGH/XTdIjnwCNdRqLfmt8UEJn/8OhnTv7tPSi1BL1TkeiTse/mcT1ycJxazH
Ux79duxaL/wuCh3IzzeBclCQzTyA+m4RL4ZxZr3hmBf5UqOdpbuFW+c1k+SimIEMI6kxb9JVhPAs
SWKDbUm9YEJeJHYGkz8rzrDf+fK30gn+hoV7zpgF9oAhtfDLrZiTRiRQIV0pVPCA9yJstS0lxHYw
U/c8F9oqe62wxVvum1wlmddI2dWRM00NP0ESzFoxN+Z779xxLZEROaQfEivMjcXoI3R9KJMpvQAu
kpGozYjWOqDf4IfX6h1AS5/Oxd/p3SwVLJ32oSdOt1HgdmNx10rsIgo0Rdxy2XHSHtR/Zde+y51K
SMQAJvogUCC+TMyn7Oq6UP/FNnMXnXUhczVVMNd4gQ93QwRaKmRU+6pRAJkKkMAy6ygGuPdGwj/C
jFJQDb7LT5lu6GNCDr/7fNHdiEaGtODzCZ3ui68a1xWC8x8eynfLtAxePZXqsz7gmWmDI7/8pWTB
HaGplJsQOnGEgA8PqjB4J2ehIx0+RXZfeGkQFiz32HeNTd2LYkM8UShS741QdldMszF9ZMCcj3N5
dCWzmzMWnjfDEEaQSIuNGcECwFijKiLZNXNxVw+XWevYAjd3QmC5ffk3qc1TwAwTIXTqxx1XHeei
AkSLs9X/O9o6svjmR4zbs/dYfqImYphweig0e4TiRYqd1ClGeheazk4/JLY5QZXnnYMWZp6Awx9g
MQk0tpXspC85tigqf/wOHSw5SWgCDOqANTioVpDq92sGdLQqmnjDSUKlFmaDr+o+p2lExJLnUMZL
QjeOfCNNVSa7aADoSTWDUUvB9MgSnxDJIbsQk3EpcdT+LdSvKRXVnybQ4wjFHB/KuWPtpvq6g4LH
o/JzQkfP+afnteE4dzoToClknCvvdCbMsjL5RQSxBx2bTXGV6TixoAn2GXGCdnqyNsNEqPv4ySRS
v0Djfc2V+nUSdRitf1PwSXUvrBlQalCe7pm/tGkIuJSSiypRCR56CHsUEf/jusLKHb3dS0pJrOEy
C0CdFnoX6H1bUSJA/71pvbG9oBrelYUFwDyjsu3WSSPeBa+ZQrv2aXkKH7q4PVaRieT7e5VG8S9v
au+9W/EH4HRolkh12MTuhYzukgly3YuwR0Ooj+sxe2GZCdPx2MRXx0PA0AbsrcmEA+KyzusMQtxT
jnfMYmUquZx8kEFCX1rfRtnSoj3lCkk39ZZqe2mw7YXxahCVHqf3vpCtbAqhQ2iatqOyH7rmsXaj
ccDftjbPCe8H9z5222fI62YJzy4h00h9ObPB7YwQWFkWrdb2kTPo3pZ488ezKyQ19XH0erJ3wpXu
RClHT7yD05j0Njr/LG/vmyjiVNUeQIw43ESwtQ5Hru7IvVyFJDgNIMqn2+xf4IbOj1TXj+HhkNYo
5l2Tysp2S5LJpy+dKKrJFG7w0+RGG4TZ7sYav35IDvi2BdKlc/xK9t51NyRUbb6EAINrEgCz5Y46
EklkXw/tQ/Li3DF260UsJ3EgPhbDvAYe/WDqBBd8ZtJ+ZTACVdjHfEn8VB2uhk0WBhWF5skt3lUt
rjyBDTLgnhylnqcnZkith/0G2xmzu/5RlrU71A6TTi2qDNNYRGpTVsVPYN7lMeL0GvryQPBIwZwh
IAR3CbbnjNC7lro+Fz5nRo+YlfmFPiz+fceMj34k2kG/wLjBHLndwSzrPCIfO4v/MXOo3UbUn6wg
6Qmf09fnCbge4rQ4Nt7TShGo6y4SNQ6gkGTQ3BG9KHjXcOP2ytl/3nQyqOw+aP/iDYNrj1cJ+yem
QxsGv65udmOQBVmHLdLC0MTz2oo1V6uMsG5ZwBcJkKHpRqqwjZOYfkXvZcFkfHhzFEunY5Cnt632
5tPtJXqe5SJuLsm/yqzFHZjD8AsmrAMou5pNjwrlhH+FXmeD+N+XLme0zC9huRxUHoBGJmGPhsx3
cD0P65yl7sqvJij5aGqGR2L3DnxnDLRoe1iWZXXX8dSjKzRrQKAtyFY/YGPmJ/gnyO97wQo2X9UL
OkUboisQUx5D8hw9dzhT0xP3n+0k/TlvTWVTyYa6jZEDhE08nVC3Xg/ZRkVrrVPCq60ue2H9YArU
xw+4zrctXnWWVWrlhZlJDtsBg5PyxMi9j7OSQX77bMkEPjuIkG0PF1xjga6VOhCZNixWsTDbF+GX
fvB0Acvz71Vpl20gIBI/qmd8kld6b9/hEKVG3RmeUKjL9xcjQN0qEx61jqSCaDLtM6QgI1l1RqIn
9N/kMbBZTAIRGqdOTPvYTwU89ChcShAuGWH1hFcMBqTAneM5z1WZs7R32reJrQaRgwy4HhVVq9XK
jwxxZ3tkKwRnv/JrEjb4dOYcB/Wv2g8gq3Hzm9y1ktXswBEYUEeWNR23OKvLQl7qlsSnPMzs5p/Z
cCicwiyYLYw9v7CEI5yadl65p7eT0X1NiLD9aV3YBKY4Z/5sYtNzD/otiO9YPqYfcRttRiMO9yF8
+KpZ32zfPeTJRX0mxJ+hr9Ra3LgnunTu8bttovR8f0ahXcqgkNwXNC8n6A88Q6frjcMLuQG7woq1
tbcVUHS70TT6iX8iZB7sfdqmQPLJz4npqwjAEyAP0io+AofVwpvQkgDCIuNM820fbbtbyy/PQeNc
rhdBN/0uonM2AmHB5g8pnHKDv6KAYCL2Vbalstnd3NaeViybjDXdXA9PYqpVDarJkQWRp0/4X+Jm
mfOAuUVHFDVYeJaEDm9wr84EslEk8gRQTl631a/ylaYRL6a4bOxCQghWd8wm/fUMzekiig7zqq6M
o/ov8QJpRkmf50oYniwMKHgt+XdwPUq1TNSjYmsIh1yXXhebAQpRlyvRqPKyoTVYKDzp8YeVmYbq
0W3q0FbpMdYvX0rWs4kJ+wxU5THnlqPY+McPODcEUdhsQGxpjuhEu1rAQ7MKKeAxwQQ3zJrB2wTc
8c2rhIrXyBheoPzjuL+qo06dprcNhsLVPVZPatbmiBUzy9hkXdEayy+CMonku2oAFat4oyZZDK5k
uKaGwG1L0ibMxM9mMoYJp2bxqnPJyIBI1efeCSyUjwpDPET7ZPs750RpU0Ch1SOBC2Nk6zadPLo7
Jy+KjybiZVRROE+de7o+pTi3ud89uQJ4zX2F0dVNIHIN2/jx8BgpwTy0uCSnCrYeNsMPns07UTQ9
yQMQKY8LrI3fAGZnSz317d2YWjHwst3e8LMsdnFumqF+4xqdtU8RVjIKIcCIh2jPq6DruKSb5Pky
Vh/6reZpf/rMmwFkSNHFiT6Ig35ncmyKtchPPPpOLD3MsHUFJPzsxRXjQbmztzhw5mEUNm29pEVq
Syr1tJNJ1q9omFek5P8BZrSuwTwRi0QtDHyRZa7zfidKToxunHmgN9VPtAqzjv3gFuzNQqjp2/sp
zjkxsI7zX8OvWZthrQNzojyFFPHk6tumzmKEJyLyS7NIMw9jKkGiJvJafqb2yl6vDKNQRYGGRO6H
lsNargtHgBzTEbv/DqhmiHJ0gNBEJE8AWvqTWRYsnY6G/KFWE8rFBErS2rkhcl3g19hF8KR53aww
rV4P+ddBxnDC3jt2B3N9h7peKFHAK77A07yOjZbscFKPTCniRqFLUKouErAH/msyNtuFC8MsUkR1
uOoaZKUAZ1D9TUamSv2ChFnx17Yk+6gMz5Tou3sh5VhUisW1PY5z01oKEoBfAokyScc054e1xfW+
BtDvs6dnu6z9RUDVKbVpxX0hKVZ1F3Dwe3+yl9cl6k84i2npcd5lBCkL7cVPBvSaPZsnLDho5mfL
ibR9GoMgTvZUNv30rdAvYlPVn7nPCT2qXWEu7w7/bGBi0qHbladpMVGc5rX/8PYE0qplttxGcA9I
XcZCMgGsvXdLH2ht+9qofE3fNSsGw7hUtiE3DhAFILN/uoZyr3WmxHaKcDvx4IAzNnhn1/K3R83W
X7DBEBgZjTsShqgpEc6Bb6iFFLPfLzXVT68yiq9fltMSRBIKxMM0uPu5FP+bA1zk61iLcNJR3kA0
g+06g0cxyS5I/GdR/FaKa5D1L+WB2zZXWmC1tRD3FAxOQ+AqAINIExTlLafO4E68A6qhU7opsR/W
dn7PhGVHzF5xoIT7rQVTyffMPPDqi2QRSnKKz9w5C034fsGo8KP9EUJXYfuARmiKruBGHM1GPdtY
wcbwcAOiC2DKoKniX8k349OSlJM2lfDNbz5xFmsXJmkcJgChziqzfW/1vEvhnpBeG/8Q7wGvwHJ5
YtXFd8Yk8JuLQAEBlNLQ1G7i9nOLxqywApPgG5BCSiM7IPY65kyDukxNY2vxX1L0CCtdzrBG6/Ac
U0ni9zl4TEg/OZ7K1An9QVlXJNxWJb24mLnx5O8FNEiLA+/RFtbjSes56EE6skw9SnMvLGdvmVgb
hzIZqJE3axn7BwwlD4d9uzC4WMsBw4LKKKop0sihcUgnYb1GO2Hku+9LEumZL2eHFMnNSyDJzWTE
tk0bubTd6E6qwmOPjsk4sjiY4z3oikH+VrExnRI34/aFtMORzrPJVWpXrzDZLWFvV4zEbcnfkkeC
k869HD5iEfyC1+oY78ilIKWnsaguhrtafpdh3zdM5gE3ewVLHCHxInskaiekTpylLCOgzdZqgoOC
Ni7gHHDph29Bs+HQTkC1b5samRm8LYhdr2GW1XtSUfHHdlxyXiiYBB/M7fCC/RYWUVgR6nUgv+OB
FmLysfMo3R/vuDmhYnuxP6KHkog1X1GzW/my3+FVg9yuKtv7OPtyd6J6yV8xXUS5YVGZdPxZX6Go
bkpw2kmeOduaQtmhbTbQNygCsQT9pcaJWxk0LJzOf6FRTU2r6A22kmQ6jVrxKhjxltniQF00qv8P
54eZP1S1huY6xWXoz53RJZwKhbiN3futCua5lpnyHNDlReBieFg/ahDvncFC+WWb97ZT++vvpw0o
sPh4qcT6bf0Eq7XG/6e7Kknxkgl1d/j8JyC1fq3WG/x/hyNGhkQJeiPJLpTWKUvnZJOkIYfgcGeY
XJSPT4oEQt+GMuQaTt+vcE2omsMEXU9d/c60dljbNnKASNJqA/m44snJFcOGg0wZ9BR0z1GYwA/C
Q91bwwvcX8xj2chXiVXiuD9L4ZGLAHYG5dzvx6Mt2TKymSFX0DioktnMCiPArUCBCXDQeifzwNGb
HFmWgOt5/NHzDCtNVpLproBokLA6G9eGQlH08y9egy4wzKnXefthUd3Y2JSRmWUKKNcFsp7gEV6F
UNALt246dqr+eLTej+8Jc7uwIK5VCCsVdPOgE4zlmWNuHXz20L8YNyZ2UeNp4tIeoWe7WuZjMhac
BD7RhXCD4R1NypFK8ar6DTvl9EVipe8JSQHyMMVUnezq589HJQBleqvVaAtDBCBrzC3n0eVKOAD6
FgEmU8xN+2cXjSvG7yOwnBI0sCFnS0oHh/AZ+LrKiAijRzTSjUpbdM0oG4ZknWeG0X0wawcGBTUE
+j99QbJpRcvL979Ilz/vrel/ESCmjMHcrHZ+WhhQnqsXAaBBLbBP39sWJWZ2W6M0r1rVu0oiufWt
TKNkELZcPIrNBy2Pudgy9oeyhb89QnWkLH8cSJB4sdgTrI6GNmD6PjnqGC16vTD4v8GMAlD2k4iY
QrB6cKqGnSi/PdCVco9XyzuSFgqlxTNho+N102LaGfaba2OWnhulD44Bcllhd+K+Rds46NgmDnyC
ohUs71/0cTGaswQmsFRNZjfsuQ8errwPmC/vw3ALIyD1933pGW7Chs6v/CKVtM8diwEQztu3xCHV
ETTiL6CHzd8/3k3sK9XpnGsmOj5pbSBYjGq2qwjj1lsYyLn8xCh2X88UOOLw6Jxb1RcrXZGJ3pTH
2brHBzgr6fADv5Nhjwpqz2qK5RiQpmQIqHlqqwSP6/F0WWEqHHgET6nYboAMcToDPNt69aeWHN3P
WnbXBEw6A41qPJPfXC0fHP9w6WAeAATjP6fzMHOF2oH8oDohAYmSAqERV+hGuCJENu6B3suo/QO4
5wc1Bs3UnzHXhgqQpXUURposS2uNmwtYfxv8zNOobQmJtqKOekcz5iW5a7BLeNwCm0CosHQoUE+Y
dHa5eJdZnmygBXXH4LIJeVu64Ji1URVLJMLD3kSGizYemr/DoVUf0373LkRM9evof7jluRWh+XD3
FjHeYKgH2mu0vJyBFKa8lW+gQQcbB6ldKZ1QwugagH95zmU4SIHCxAFzNCeVIht5XCBZeFJQ2Pxp
dRBKppk9/l3DNIT+ScR/KgXIYKQcpx5MJPR0qarrghC50c2vkbxFkEn76TUZj38q3qp4ls+NH/sw
xhJDBwwf276dDLr0OlIYjQQn8ZiTvhWECCw3bDjaibO+hLfw4RzY2jiONF0vHFLWQNnr371yxrKc
cmm4ba1UGbQpUMNg2lWdJUzFAjDqx1/eySBMZFrJ0wVjwMWlWZp5PIF/+dZg/MqEZhzqIQz9DWaa
j4/Kp4vvQWnsk5HJwcFwqdtzjgCBSF6/JHDXJk45GlXFYZAf6uUshZ4B7sDas5B2Q1Op/em9j+g8
Y0FOKHHQVnFgLhWodzgEXjCIsezw8fx/f6njZsa6c/AAprjH3P0+4BHOTZn2CqRyKl82h2p2SclX
SyvQVgFkvRsjD7iWA+zsa9uBmjraYgnrvunxypu8GpTz/n89uqK3VpjdodI3swlIB8VwaRb5s4oc
c7R/UayWiM7Sg0gdJqxBq6SnIZisk9cEzkITcZ85XidGt50PB36MYTx3xpJc0uSgOoyYpS/MPtV/
bbH7wHfQUurL0zRavcI4prBcyz2v2/HxuHKIClP9mIKzPKFSnWzx0jQ5zUd+WfgGEMWJ6Y2FtAM+
J1UahaLYHZWp35p9SvEepiqw9dtAf2ytFY7u0SnzT2lHWYgI6jEpeFnfuV06z1Bj0gBS1Mb3gZLY
k0yf6uAnXHQOEQ9NCW5tF2R3h9ZvnRgwHl6xPtWeql+Echl9vQsEf7RsvuDaiHjHWLc00Jwo8RK6
YBVeRMuMB1wxTS+DRQrR53imyPFbbzWet9PtWMFkAr4iRPhWApQAaA0HBpehTUU6yTXA/RabCNaA
fFgBROsRlns9dNaEeXGxjEsPbYhZMNIZWsCv6ANBAbrVAqSjW6L76QYzu0utoguaIcDmZy8JaN8f
D0XEO5fIlbiYCsugqgow3sPPKeABI0ySnFFDm/5yWUizqBGLXi1A9Hm6Tj/S0cL47u5HHodT3Ggp
Gvj8s0EGvNLQIvvGllzK+ujJRAsn+9f9LFI/gB+YQXCGyiMct23oe+s0tF/HJvpNXtr5eaK67VS6
oFppxiZWK/+U4pkR5JnhKZzwaqPA6jGFAQJBkDecmOvJ/VdmkVBxGXNeBAQ9EZFvmKhjK5D/s2+z
uoIevbYVd8AN1JFbncN+UywGqSUi8FI9/R829T0aT4eXzIs/dHA33+FEs2Tdjz1Ueq/m82tWH+tQ
jN7UFq4sE9R9WBiuSHw+hqEx0Pu/owXwMWzqyc7i9wJU6ZkIXAZCmZCjDsD0axaTT2kHU1Sz/Zaf
8mhbRLoI9fGxp/IuTRgY35/a7lWl2cmRozTO83s/PB0jBHkHX+d/LOgFF1F/XsLTDrUJsd/n3I4F
bI8wogzf/wenLpheF43rSZRxeYsozq9OxmN8p+2KxUfqbMmsh5WKdygFnVSGaz/867pOPSAekpXs
ukBr4hQdyVr0EyHClThRbvbrvwHgrQs/Nz/QCEuxH8hw5MtY93Ktw8uG/hWer9JA9ziCXOjAwgSy
Ci5aKYh6F4zQP6qw/Gkfa0BXFUH/sRA51FEDsZ4gLLGU1CdgAVYmzkCv942c7lOYHhg5Z1udyOUK
H0w5RXXnOhjtXW07XnGvUuDxGE8b3VzGHedbxTrdgSNx1Lry/7m27eLGoLa4YnEIaiXTofyNjUsM
k+1TfxYdsmB70PlWaVbbbRlOUeeD5WzWc2F5mQtr5xFwEm2AHNZYAG0SLXwk3kGrlAnkcDkOl1RF
xYVXjpVN7CGoroZjNbiuoAJF8HyMSDJHWVp7Sm+9vDT7i6p9o4k4/f+ycgIU9HmTQR0jj+kfHCPc
QXNvu/k2bEXdd21TgnGw+M5+kaCqgcBkVt3AvBsP/FWMjLlijLq+Y6RX5lgwypyfFfb+prSHBTMW
o5lLApZjwdMsraLJDvuG2zsbp9KeQbfF+3P7tp4MEM74TjgTGD5Cwqjx+KA1pfz4C+4rPeBJRL/u
BQiZOzPbyHUD2+v7maHGcumToRCDkLPVY7gGf8AtrOB5gQkbCYCv0uY8LcTOb/+yKQ3IjqsZQtxh
H85jP3dFEhVA1c4IcRPtb+9h5BHfSTdcv8Nx2ZTZTcTh4m+eSAmHtDj0/aLf9lxlujZ1rYiSL4mh
2xm3sA/Oym4axM37jF4C3R/7T3UKBqyFcH+PeQbcEKSocpzfUfc2gbDSh8ffMTaVqX1f81McdfY1
pCnFBHQDP2fBM7SAhYG2PSOl0UPa43/IBBqu8+se8eI3w6UXa1OcIOvagTLv2fLvYmSjU61NXNiN
yKVT7k7NU0HIyFUQoC2I4JxXtIvq8fTyE4xZcRg9VfL+dN3QxSgcrNBble0/HvF6reG3Vq/8IU1N
ckom8IeXseZHjMA90mvH4GmHmkKFQTyX3drSITO5YcD5vA/UJ8+11a+7Bd9rvdwomrrpRe8I5RHC
3oLR16i/F6sogAoOZNer4yQZJd77mPx0xUr+aEYwLCcSKZaKOHZ+nygo0BMikR3PJRgSeT5iQDYl
b3n+7gCI75SkOVW9tA62n/pDmH5fmcwREvx6uXaaaCEOrcw609vIfrSYRR7QZE3aLW4nR08OVKd1
ZZiw3FoiaO0aYIkgmhHbyZVWo3zVYPoQsXLTyrYCaONBpIAzsMICsb4vSAEzFoRF/bhlkY2i19/g
oIzL38ResgpfLLg8/hKHEnsDMNpbwHFF7u1RBplQYmybgsMQR63sdW1JSTBSgSqX0X6xlXSN9bLG
+oToZCqQrz+WsQu4P1KFi8+Nxj1P8XtRwMQfKtFBhUH7j/naAGRDF9x1CR1W6T3JHTpUYAJVTsPU
g3XY9Ta7XXpxUGi2G3DxB2uYDPLbVj8Z61Nql6f+ouYUPvQy1pAXKBms1PABHxiyPqs9PJgw79ED
onIw3MDRG93QRDq8+rM/1sj604h1hWVyS4uNSyHfrUCTpReAmEobDNrNpWAPmCa0MjiRGhhekyGg
xun5wgLBNDQQfTTbLkGvO87fbe+n5HIljGI/Iuu3o6Jr+kVT6Og0y8XWsPUncv400W2djZYY/iuD
7sZH3KPALWhJcguR7mhz0YM71oy0YEnZx63A2QjgqzOez4e46N+G8F+r7qXBkqrTUReO2M3iECQk
YLsyyDLsSvrXM9DOhetbd4gKmAt7lO6CdIkiWhwqWWA01G1aObo8+6zlrBzbfrAyAzJlQ9Q9hQwP
fzSuo9xLlXj0NC/wYuHR/mfHDjXrQVdOi6e1pQoG6n+heHR0DYqc89AD8zgFQuQUhvaAFcc3DNcG
pcI1V+nyCX6I+wVUmwBt7ZAroEPka72Mvah7ZaEicooO/QcAOhR46FKaJ2m/Itl+uydfCp70hzoo
ZoYrgrMeyq1T8CmIEigkNieV4F0TtVMicfRUAck2Ui5S9SnER8b58EQLluPxMcSUaLoX9cD2dIGX
SsrVxucC0q/3Px9oGLutTvDkcEEYDJ74BMR/dwRt3N0F3vJQ4c9aFupdWfaH9gCIA1p7w8OgHdEv
tNQ7OnFOaiNoeZRMTEL4nSyXyq6+CKA1Nd+nRxEWD6nb6I/801sv1m4cGw52pcjVKM/MQlVt5Qxl
Uvm+ajK3ZBoweNtwngoJ2G1UP/WJpvbBWMSekxy1BIH6tHAOx2BfLFvbXe1fBu5a2rEaiJoH6o18
SPSDmGHl4W/DQr2Qs21FVUIuDRAnbpou91YmcXpE2cnmcMHSGHRq6mZJgEROnpaaA3tQuDdzDp7T
IhOcz4BsabMZFr6WwnsJRM8CYnCnwFX+xWhr6F0AyRqhSbnsvmHEYr7Z4ApcA6DQJXPJC/6wr1EA
xBq7mqpII8H76wBHCCtl9lQ3lRW8oVL115FhZF2u6m78C/FmJqH5PnxYygEOwvrwnFPCP0daN3dQ
ZEEcX7LAfZOwedmBOe/4y5CiE77saOeiQefEwlclfGPTGu6b+xuQiOaVMviI89LsC0ZGclfRpQQ8
NYbV4CNxW62nHLq9IE+EPwa0ALkxdprsi1BX6iOJSBavTQMahY/pzy4H7o9LjiyU7LMZ+nTV8lSB
Iy90MqJMQ3ysr6TQmOn4Fq+XkZspYDJ0QPAWV8yf3lo2TtQzmpcaNua5TYhQb6VDMLGPB6c62d5S
EpBLjkUCO8x7y3CZiM6b+9idrIc1qtOIFwBWb54cp1DwX3/gYcDedusjcSfoX1ASWGDpWYjkhrdy
nn+41If3wgo1mRLbFsnPc9R18SgjsfoCmkE730MQ7ZTVezyi7R5eB4vQHpCFZqStcak6yqCWXByt
jNWlZAeiFbRM2amOyYIPC/zeJfLUJmnpBjY3mSKgsVHoyLjyARbpwhexYzX4U0+eXRu0NaFFNVCV
FGUtppAuGw08o6FY4SZjx42377ixxrmI5SmKLb9N/gPRw0a49vg0rQLsy4JIdAL4MCfP8Ricsflt
a0uzuIXhdETHmltVFO3xjJX8g0JWtX4C+o2rTEG+ff96JyNr5qO7g1b8a58MKXZrWU6t+9MJIQ/z
ec0QetWpTO5REUepZ0zWSOFUprmcw/9u7IP7YCGKmtZPvYQRk225k1ptHptdxAHrYz8fHq4tsht/
iKKyDpyU8a01rCt5uINxeWFeCMmHYEsw5/m7GSoq7En1U00kHLhZDWq4TCg6vOo6pQlM4v8UBxH0
ga94Y32eGLJQ8ORwW9WtWQQz8Es7Fy5KzjDM6RxBUI0Tnwe8YpLdK1SrG4ooYyqwusk3XLGR2J3Z
p23j5tQMKo7sz6Wf2vSm1dux6PJhbZ+SVSNj1qGkrPTXLkIXYUjajERjy7xWFi9tYzyN6iZdjOSS
ukg0aA7AGF4BhPF397gKLpF4b3KgG0KJrTuXiyIc5TqBcU9sgH8kcIo++4YvrTsoI0Z2JL6xfkw/
yprXKEMVaggzFPkcMtVdTuwFY0um3cNG+hskEE/OqPa68JqPGCYEr2FlnFeNyIMeH6+TjqK5Ug9N
9ATp8BmHL5LrB5pf9d5MM/H5XLVRIZAfVM7uKPwC8ovl+paF3L842xykIs8N+SXe83LzdXHoGLRK
xPhPRhZzSfX9A7VputZrMbEgXSBx6jupJZ5EuHlyp2E0V45V1V6hPgk/3ZtjnVggbEvu+Qx++4KM
50dtKBX+2O5hE9R8vDk9zaUNkoiOvHu+QfOFJmZ1gVnO9stbALbP2z5VHL78VsPUdtsKBB/eXoxn
iCWj6CRULQc68l1oxcSEkidrPcdjAScINWIkEJ4eOkbKWfCGdeoYl5aDdTBNinXC/BNGjGGWvFbg
VpR7hHPobbLfyhu0YD9qDCeaSash9abdrZiC+4zJMNpPJk1CdTmYpqUWZj35m+TbLBKpS1YQcr2z
c0HkgvqkfEcCAoFz0/2w8W3c6cUrOnIOw9ctCVwmkWeEl+u6FJGRCDAampLAPZ8c/qAREZjTkn1g
EtTj/HoceJiRCMRcKFV7VmKBEeFek0Y53XG8yISATxsdKzl5pRwVFGpnxjMcPN1CszEdECvbwRuV
dX2mKiClOwLMc7qfUm4tmkxb5OBD60IqFjJMv3cqsTB1aps7c+JFO1a3m2OLp4p9Jb1S4+1DIFEB
BVlkvVkK6sKGdkG3h6k16MdJG6XCwJOgdGbGfTNp8WroJUbrbh+DpgiN0iFPKZ5Ig2kbdyhvZasd
SuxW4JThm0k6Q+cxqcUERO3IHBW//WpAn2NTFxNkc3a0Eqm55FBcaJSpkOmXxz2QHtXU9/mQ4473
QNBiA7pZ90WIFcA7j1nv9GchvX6jdJZHE76sKrJbcF4Yhp/85dJN+U4ZVXtXvF6Vkxx/8UxxZuRb
TkEzDYDAKxJixOmb5QZoQFK1dxFPR6rYEB36xDlSE8OTfEBTrQvkNDAjIaOtsvoUTuh4dXyhkdvh
D9/2iWcHEJ1ONrVdypxHSpOJ+vpw1sB8M9+M73eQH45gNuMl3umlcKZKxHWkLtciRfODqd/fhLvv
tJ+obvi8/F52NvsK/2aAWeZC7+RwCPATITCcoPxia46hqo54P81BA8roR6LkjRVzBqC6Oy6X0938
pKyEpMhtenaLXYWCH6okYnU6ajz/0aVJgr+BBIiTYn5UmLcrarWhjmyd99z7AL6q/bOEkGzBNZrB
6p6oN9F1XpEPzJVeAXfp3Cpa5IeYTgiZCHSog1XjlIrytqGwCV/4cCy6zem5mJZjDQx1Z83/QtzZ
iSN2jjNxudYTyA9qgp29X+4Lu3H/ZEKgjhzFPV6aiXu+NOQGSFvf1bpdtaqA8XXnvVzjeORlb4vE
EwJaJtXl1z6WuekVKkTrVsacPwrkzwI3aJ9ezdTrPk2QFDuni1b8x1vG6EDjDpRgdq5+lC/O23av
lDqKRbCHPG899gIalgqdc1V3EawlR7lxn/ydERWBn9LsPuvBuNm1JEy/3iJay6K7zbdYw2eKpc91
iNd0UmbU4LPejHaWphWqzMy4BSC5AqGrXSdarT48yeuuNm+GOlHENqB+8iVQysL1fTwKvU2tSqNE
D6ZrkOCTaqFqXiZMwK84+UY/pSoZvrRfqaa3fa1jyRfpia1hKtstzCOR0Q9eOlMQ8XMPgn/P8pz9
e04Y6rVm5rIhL6NnlwM/Tkps1cI3C9Y8fKxKW8WGhCjKr7QHZkKf3L+VNNj6uqApjs7JHuMsmhUd
hO04+E/0e/AsSHFKojXVo730ta16opIRESlxJ02LjEykWQ0AEOWm4Shu9TqDAApFqNWVyXE+TvXM
0PtJ99RCJQYa6XjwatOBP5vxFBTrsKMPCiuTSpwHXz0A2c8a5RO3/5v5dNNWa2As/o16a1z18mgy
SR9TdEHxXqjn44PBbXTpU8iMxc7CzhEAUOd31fAcKN/jJc8NJln8yi038/Rh1X0n22mxZgIyIZNs
l1PN9dfT0bPJyagModVjJf/CR1XumjMj5yCrOJDmU6kSfv8z1xy2j2XlCM9wELH24xRpaanlMvgP
/GV4wgxR6qu0go+ndYGVrrBe70gUKVYSeOtiXm4rW8yf7KLcY4YDRLPNYywHxsMjXPecaGnuzYim
pU9cPkJRmAmibKOuqCc2hub4ZzdrVUs48xLbdlN7bzN5mtWUBZNdl4qoGvwcFPfL56hvWo9zW+GG
LZ3vBpG7yDUDLYIuArIJk1G5ehn6cR1hLWbLwLBhzlrxblBLGVch0OQz91YRuE/029QnA+jT9loW
9qVCsnKRNgVd2JxHYg+h8GPx0WfjNmhO6Sw7u6jj2wJyrrYpsqUBGPcPUICsvt3t5jNTTPEvjcxK
7o0UFqUm06iY6XMBevDI9COAtjLYt44DcwKAuqr1QBAx/qaGBYplG/gy4ZFDfzj1B91ok5M1wLnr
NC11r7aG2sFlBs3DmRUWC1ehchmKnEehZzyKTxT+iLoYcPsaLSmsODeFm1vVGTw16CK5gzML7ly5
W67VuF/alEobft917sau1hrUxsz5rn1xmuXVP3igB2ryurPJUoWYzfjlLUuNM373P+TJ2t7zKpGF
HM46UuAniB0dFnbnI2DBjWQqkktWjnjJHsHFdXE4IaXroifrzoHYa7lVxchIcFYcGwfHFFaWh83u
HkwaxiMnn1XlHnTEWFmSnZUG6QQdNdcmvfazDEOAwJycE+uMC74rvaGOKk/bDOmlJ2ZduZ27PlGu
t0wycoX6Baxi60Amw08+t/uhjVopWtfmgUTZVfQJiYU9QQT1ZFVYdscXZzNBzfqocV8fYrwUZKsQ
fw8euW6ujt8A0hplHR9A5Cn68yKlVm1oCQcSNlb/+9jmWmCAKtMsMacpCfO6d3uKc7i4j9Ibo2Ix
KU4jlGD+7fI+ifM9VUOg106q8xmUOdp9kT5pRodf+0uWoKwQltbSB16NBaIzHTbc3Z4h+m1LwizK
nlU3NjFQxKuKxKev7XNcdb8AhbF8VkOeQZkSvn72DOb6cCfLbx1UkN35uaH1mhXb9j00veomWiZM
uwVqk8GLCGLEiDKCosH1su6al4wgOvcGHFggbyRAkJGlmHon9wT9NXaBa20hMMKCHndIEq/0Yx6Y
QZJfjDRKgkvWCS0b2ly/QrmJlo51fHjXupbRD4IV8bgIMHjdMVUbvD2q4omcONLOwWfHCjrp4z+c
GPkmYxFs+Ai2E0GHjdxSbvGJd4ivKJQlPWUG0KNq0/8g+XEdRXjMwdpkp1aQuKT8sJMJT2K6XIIZ
iMtCD28owz++Au5UCQvvJfek/bUdM9awqNbIuDc8EQOX40XYjnhqjopolc3zV5CHcZMN2iAW0d1N
MeLLNJxQe+AoUeg8gBXEnM9digvUsYGj1qxPxtdJizxXHh0XXXyGXUKEC3WAuCIATBHJElZ0EOxt
LE9bGOBQRR0Aqf73brgqEYXnNW9vJLunfTZSdA0q3aXMMe/dCos63vUTvU6kFEQPTOLPTvzpG+23
La5HpB5mppNmmCDhzVUiZxu5Mp/sO5d40fKA/5G7ap1DJdBBVErmi+sHgZZXkgni4hJ1Eznnxaew
XKo1w9934CBjXcbf7PoFLOrgEWbm42Gd65d7bJjRBgOwdGuf5w7f2nibcKtAONucjFhalEROrh1Z
ia8u1AFd+OhtoZ1mZWPUYzzzClbAo3wk+KXe+iOc55s81HtxphI2jBMcVkaZN0Cx5yKbd1Gfhclc
Wg7T+1TvL4D2elrOknGIx33RwwQC21GIZ6Suh3hmh+d8qdsJ9EoQpLdNSuDoSa7vzFLEqBMd4pzG
o3K1I82A9e+iL3w+8nT7kKAy+mECeC+VdTy0C4cgBWj0uAgdtQOMvHqYvbl1XZvWbkToVsV5S97Z
pHkIAyLmZXIy33CSsstwlWPxIwFPHISTKOIVtzfsa8gFM/166hLhRb8hRzXv5/6d8VubQM2VrHqw
yw9OWZNuvsZaSGqWARe9qD366XuAognJNO6L/GjcO/KaFIyRbJ+sX0KkvZ+vQzgZxwjU7F0WpoFk
OScOXaEl+jfw7qVs916qHGD2RqumXaYQM6U9mkKJsgZNmV3EySvrEqNZ7DiaxAaoXDFaDc/MBpth
bLq/5q5VN9gC3E7nTqdRggnL/kggU8TTteS3cDZELHLq0T0J7Phy+fxHpUbEjHQPiTEkXYA8rkON
gOHzFlaxvxJOhiZzmUq1OoRl+zx/kWdbjA+a5xceUYnHS5jL70kQu3NxrNuO+eakMGq4sHAGSqLP
egn5n9Zo6M6kqR4IjO9pUUMoNOIKQaQ3ps30ltusPYLaV/QWUsRwfAJeLXiC04DYFQOP3Tp8uGYd
Jyiz1otJb2D5OrELXDqmQZbxv1dvkRvDxX/2PFn/0fQU8tdEX7yLe5DBxVKd4oa1lpaPsvAW6z+i
VqUeHYNW/yCll/kfWwh+pZjkASXmThiZA8g0soH1MDu65OZB8ArRxkCXqXNV0PuPLmx9cgZdA/3g
I0bAL/km9nutZ4AgxrJKu4r2XMjdKTj848mmdwA9HN9OVdB4jgbDTYxvinLOxdSNNaTyGRJ2NoGl
D6bpRgWhULYUBFwpps+r4KTkXHAEbP61Nrcox65SiwjzuZN1a9MnKQ+DOzV10nHO+T7AOLcsR1P8
G4NyLaNs8uU3VkU9PffEigDsrydBaI8NKXHuIuIoK4RyHAlO13CxyelHT47qVQ1LvHWE5SSOJimW
iseDQHH8IWnRUcIlBZoSKJgZhzcW4V3HgRgSuc56x9Wf4H40XNgr9UiqTkS+KWgSUAPMKURU04qV
B1C0g1RilGhNIgwh561e2mEzHhXx5ynLuQom2JNijkfgeYbCNeHvb4G+rKQlym8wt+b02RNiLVqt
uXDX+uy1jdemRR/fr0p/nNPWPMwMflIEHg/EcOvErgn/q6FPrBKct+M9cdEXt37YJ/2j50ZYkGju
txaiDb90XknqQbQDWTB7da3w5FLCQoGcGojmzcBhlz0smKo3wS9CBlw027mm6fz6a8Sfrn409Y7m
bMB08QFqf34EaSVo5ChPqpls+PdoV/mo80PwwK1EMmo4aCnQCwBdJfH6vdKBlglikjsJIbWXPrN3
9+SUrtcZp0fxM4tsgAGXm+933F9E0cI954SOWwH7HFLjDvQOxsNwz8cR1ei3pYnQLfZerSjf4vel
EkimkL/MLT90zGLSCiaplUW/oruWhO7wtwt8HptJDIjJ9n4Uo//EBwb/d8RcNIlfNOlayPndkQOR
qMVmbnt2s4EzV054WIKhwwRzGbBe+jO3JBsnXsdkBD0Zz1Nf82JrLU8tiXZopyvksPlWw54IFCmr
0r5aVVYdreALAPPl7EzrlRoL0RW+E1ALB1crYvewVxc8nfZkQr9pTrZWNbJLAnnSvdzdFiq4OVzl
wbrT4rjhpa2zgYFxUjod8Q3lKPJwtVsXt4A41ZmSOQKZsVHnvLXS4G7DBHjKGSL6BiOEiyeu9c57
fVB/s4TLJk4GHJZzzFAA0MfAMeuhrQmguoLRiv/of59yYzm64tSXfC1gHn/GVXMWzBQwCEBglK6S
yroeUmuvEWxtfG7U2gQV1jwpJMRtdEzZBCMEJUbngv126qCAAS8Ic1NgGT5nA4uTCk9qt7iAvAtb
e7WOLXYjus84cG9oNtUNvZNsBFTkjldYOGp06j6BFropYDyJ3vcI1jTpaJsVDEn/nG5kNC4Kucgn
wkvDFnq/Iqc0gjTwhGjTvTrdOlpjk4KKftbFhLdwMliOIv4CDDm5s4IIxKuWvo+jtYG0Whx8fqAp
r2Cpw6b9eB9tqJMNr36VkvQ/1rXlw3PXO8sfe1cPGMP0mM758/1KpCIzNzZvZUrdbsKg6M9WwUvr
hcS8PeqMn4sl3SiYFJpG+redppTq06awbTGeBYrTR5ijP9n6l2rvLlGMf9abeRbkOC1CF28oTmKl
CsHMl+DYGvR2zhYyl1UtmFApffaLpQ9YUyPvmYOIlm7xYs15RN3O+2h/sdCZkHmk5shOVOoDVhp5
goLwbAw+Yyw8+T83eMJ3Z5jiY8rRAFpUFidrUGaP8QNPEy/jdiamayLhoWVg5+ZSvuvJGoPO+2DK
W/HATPu+dojFopu3FY2KpTTnfLKnLjGX5zM5R6ORCPfmrNfso/EuF8aXodHzHzI+1RZzTy+izfSD
inqzHTbvQV4OEwLK/79qr6s/pRGdT5Q5pgUjBArNeyGMJK9KbBSgPbkbY1n6ZOsBaPQOTyv5tic8
annDb+Oy4ywxqEhEMl5zmKdnQGzYZeG6eTqVLJYCe8+KFMbVgZ/eXmfu5cR2YlzM2tpAdcdudtaD
+JP98zdjofBou6RLbOpyq6dIVgWcMt8Z06cHVvl9k6lgPCz6Zy7Ft0R0ybmX3wM14mxLWIGdQbC2
nOYSiK2lYZo6zbeqdXgfrb3GDn+PsnhmjXL/7rkDxnSFwGIWFbn/SEHtNN+Ht2FVnIqTHzrpV0oD
CPwSLMmJxhhe/jtfdfPEcbnfoNokCEiFLJE3FprXV+RA3fx1n/fCTChJIHZ8NeyMevs3A0pLPwiU
fAKWaveduiBg2zn/40urWMnYzHfeywlgRUEDe/3VL2xskkIIKEoPJzXFDPKc3/tBvEs0jw5M8aNB
okr2xiD/hVmyg28ZITDxZugOBB2x6njujLA7KhBO4yY50RgPOKqTgBGi8kc0+vx3HtO3WyCFUAT1
Jcya7rhX/EF6puFZPCE/qJNfXz0sDB/BHZzMpiy/9QbNvgSantWl9ezkAa//IxvyPiUCupwI1/Xw
LKeP6PpOSdP4VyFk1y3E8rEN68j6Lql+7Uw68i1vzfFKWST8fenO5ztdEHmHIPuN/mxzd9zEnkmt
q3IMsSug68B3jkW0aa4HxzxDaEbTqsUUdryUcQegEbQztiID/9i4O3/1m87vaYMyn4KTYSUCr7Yf
XAXkMSyvtavVzjISH9zyvn2furwRXf5IFx4DHg/5a7GyC+FZ0zbxVw0JVReV7YJ7+EwzCWG8Pvgi
64LlQJiPqKw947Hu0NvnjrMu+HiztQHvdvTiD95p02bsvPvotJJNFPO3kIKMjkny/7jqf6Fguvgi
gsdT3jVavwlNPiA0XCThgWKPEuR2iu2g3zivbfRSKS1Uy0Z1aBEXw9adyN1PW3if/NvM166DE1xW
vI4n6pAggky5JSuXGYp0rF7Gf5cPZrL/+3C4LcGoDK7JZIQRh/5E+L9o7dHfHZDQagkJG3/f9Ng+
hhU5Dq1bVpOGXoofPYQnMhuPRWhJGv/S7+0SBgbl9NhSxss6nOo0Aes2G5YfGeDSbK9osX10soGw
rH2HGyi93+HAIhz3epGddWU4e1D22wCfOia1l00ZbirhVRVbnGB4W0nz0cj2H0zl12nuNSrmXQpj
ffbdQXaHkgcPMHi0YrUi+AMhTcotMgTT9JAC5nqHhH0eMnhSuI6RftFnWHUGcBgUtbr1wHMZxzg6
Ogn7RWR4rzg74XvHrHGIM3RBEvbzXLZ+n/tu0idGOWvqg+fa4sUYourqhjyNe/yrHDeC7OisnG1Q
2FqXQvYLpVik0g9v2jnHfuuCUmuYW27xl6Z4aLeC8QmjRbz7OM3nHn9LqYoG9RY3l7a/0vbaf8lQ
NmICkt48rDECd/4Ur2kFmR4dcGVoWLf7TFi4QbXxhIgCQh0aQJRQDtGarcSdgTiCsw1znO6XrdNh
q7tipUbH/gZom1jyuryspvZiUvY4B6lsL5R95iVc+kupPL6c7N9E4oUVhEMrmz2aQSprqZxtmEYW
bk5ueO4GQzAnB360oNzAW6GbndX34lzXwWBRoUTMzgUNgb98saEaKK6z3KV73/VCIfskPI/YIQ8z
Hz4ywuVj4N3DzyWLpcaJK5Rq/InOT+FtK7FErmyZhLhHJv0lJmj/uiW5XJLf3sJNmxL4omTWi8oE
rS2dTcHDxAZf7z1c7Vh2hZ959dkBZJnauL84ImB6gdaKDuuom3j28k0Yoz2dFl5xVOWeVnbcQ8WH
gAIX31F/4Vay0eIzELOKTZ5eG+kJfPtXku80Zf8GvHW5Tzj3tlEPvX46Q/Y989axBrwDU1Wfr4OU
UxpfVVE+t38J8XToq9w/M3ou6CTKgbnaaueSkyOuy5WU6yuiaJYeZ+V0NwVwCPvsJf+hHRXNndgl
cKvDyvWAzMHULJOU74rBmlRDsF3iRx1hozRwdDlhJq/P3dmEflyrd0LVu8UL0WISIS5wO5r5jDsf
UBf/qy9balh8bbjyK3XTObYQplwoGMNM8hvYAHZ6gbgXil/ppyGzrbj0uJiMnS71hprE7ptXXxue
NfbsVOo+Szwd3vIKsZbsu3pwQ8iK5miJl84oLB1dL0G89Zzpzz4jl/6UX6tAGiIg7qP5je0J7tPe
lNPMGnHteyJGSc81JuhDeL6tbxJFkcAV8OejIn6D17o13fsr17bk43wa+e2oGEYLDc2lJFoYLgZm
Z4nW/D4lByfb5JaSSlAajlSen0zosJ1tDzbPHwjg2weyakgBrfedjE6pBlpVzxg9jCAPFXXONbGO
NQGl/n06/K0ADfVnF8gz86dXBT0+RcpTn2uqjHHEHTaynZziDkFHKdT98szfszc/Ir7GFjCO2Uvt
6kP7upnbWfMpaC9uctx4YaJs1jDhMG5GJNcfE+izFMfVcGPMmVTqrz5ZI/lRSr7A2rbZ3OKRHfNl
AGGuiJ9LK4wNJYGI6/xMeScieq0Ep02PfeL09mjg32p/FJV0e8U/XZ2no1VR4OvKmD3Kc8uLuPH0
yWTSorCNwS5YUKp5etLB1Qq1b2CcHoYtLK6g8m9XnNajwXxC7eaSEGpTF/eXFKYQzdf4LUcerTv4
UjjpZ09LeXlUKc1eVu4zMWYZK6/Ra1o3JawF8IEDg7SKvFvs96H1OdvQUxX48eE7/ekegcHMc64/
9a/0RF8GLkWNmEvXA7Jao43m7zw8x78bQpH+TePXm6ZlprRKBT+FqEY5exwJuUNlCZzmyecBgF2H
6IQ8R5YE1k0a8mFzWzyJm1OlihKYM6fV2NK2pelZSqzQBYzO9k9+B/l8qM+ka+ve6B1UrVSa1KPe
wmQfVUBsujfksyKkRmQJHvPR4TZR3p4kchWYZZIHkvhCWdZLBJB3S/YuY3xgn6nLA3mktUNPlgxR
wKNhTqCAFb2rAnchI8JtwpWQ5NWObalcEdT7Mayj8JLYnTAv5YBY5nTNZb18c9ghcNRwY513IWcz
QSdXys921nbmgbeHz/PKT0hB+7Pnf979SJwIV334nUbIGXD85ShScGYOi7DsxjCNBKv16n5gYe09
ohyHctE2hm/Vp1kOcO9TDcYfUVNcwoYgy2ckl8NBLOjOHou6c84tKZfjjPyqUImQxH0VOkgbXuYS
GYwMADi9kVwI9i6kulatdeGq7Ds+pnuR5CWC392vs75tAjmHgopHrX3F0Fwj1tGTaCMhJZmFKgc3
tkz7/Wltkm2bmcjBH+P3U4GegnvnerJOUJX1bWlre7pb8GUURZw1D6UoS88w5S3WoTowWun81XQN
10lN0550B7aVl679mxSeyPgHqVHSU7cNbP04mfDc5woLnN2yKN1Ge+UO5VKOeW1MqUEulAqyDc2Y
BbIg/4uGLtE5rq/6/dNwlODowQXNWzsX9/LKcnIEcYOEV1y4CG3n+m939u2t6pNNBQOWwwZd6z6Q
KzsLkmHeO+hPqiPyKLDuy9TO3c3gJZyKyt/yltMss82/f7btYUqyHK7PEBqLzTwzDs7/3dgvJqEV
v0VqpQaMS09OAOMbLG9UptHb3U5YXdy5uYXG5FYgClMzq8RoWd/ev3e4x41NHNlsGNAnXV3XUrIN
WN/w8wLS1yJ/quOYTqRuzaqFjS9D4g77TO/bF8Uxknrw+vsrzHFW1nw2AMwsFUJuJuQkrgylxLk4
5ZvaCn+i1eIfevHP4bArvRoPvseU0IGvnhrAzO+QXTBUnee0NmjqUa1HU1gcTY5JN7OjvbwDOWV+
OTYKh6/mxe5sTfhTXXDyJ7WShEl2X0zWV/DFuWcl2onkf5TQhgqBN7Vq6QiZI+4RM8nQnJj4OIOG
AthcBOKjhx4GTeX6x5LNyeR/v0kEWsY2x8PY8o2V5WSyUsjwPmUc8OEnll3l9R/nyT1wX9wkCyEQ
TtSb7D/TNrjeerdUfEOYvglkM3QvULvVmu1rVUGK8jt4gELMplFz0mGKYcu5OGoWsqkC42mijT0w
apXIvpGsYWvw2fUe+O0MQpU+rqcc6iCtXlV8cFj1+L9LaJPX5INUC++9bpTMUVw9ost/7XHakdL2
Kd+wkFwNkK8fW8RM6xNsMA7Fwy2e+FLx0fuhlWQ/PoyMSYgxG+RQm7/13K2Biv5dX/ECtGHgty21
KcWVAzr0e9lk5TJafbQmcYay3hoRxLtqKxV1PcrTt/PSOf1NhLI4sginy94Q7Zw+QphzlL5aiQJW
7R0DscYbuwt6bj8HZWHOuHIJ+JPNFL2NvCPd3Lskfbyy+8ffLvW4uL2wx6Z6kkshWk+N5xB941Ni
hIQ8S1zWqyLOoZx4biUfZY2b2dMPiWN6mOztWcgJfper8D/Zk/XHrDlvvmnDyHjeRNG5kFhrKqJA
tUhhXzSmxXib1bxCBo1MRa0ds0pDk93IF8P/f81TyPc9zUUHAAwcJuckLprzRIM0TtA5RzezkeOI
rXfbxxY+oeOdcyh1ASUksDYjCld/s0r0zmHjGZVx4cHAsZCdBCjUSsRURtfIKXkXqFtu8oUCl/qf
ca6ePxjvw55JeUnuxiZTMFeGLVLFgtfdW7uysn8U+1yPyzHkO6ThY3vizwKgYpVCHMtHHTrJsXlF
6tdp5Sy0QMQmOSSnC33+VFL/zd3sx2B26rMuT0e25eBYc5zQ6L0OGckOC4ysU67YP4xpYnOWRuwp
ZNv9fKzqka6eOuLU2T624+SeePTQKEtEfKpe7iHtMVKx6Wsoatc13LbiPOsjiyr3qzdSPr+WVHfT
tUGHvL80jP/43sACT0MZE5i1zP5Hrue0H92docH6+D2h7SewL/K8ZFQi3oFlDPqa1PDG+kv9M9Vk
fXvEjnTjcKlW99dWLwb4Qh5EpxLU+cGsbli4CKZlK7Xfg8LMhGLL2wLEqdeR95kQ0SuHOOtR2WRV
je5vNDMs0svEm1BU8MY2Rl4dCLIrohBVTNi8Pyyr63eQ3YOqwnV2zZNm2TBBOgZfOdvevzcOtE9E
7x5XqemwtHAVMhzoHL0X+W5YmtTnWmeMQr63j7hVIQ8jGusaH1ej+YM3pasg5VjQzVWcDadDCwmB
zFnPWU5tGImLiULQx8e9HunlkMRxYsZsw/vM4fjY9WWwJIICW1bQJSD6PEkO+Rvl9e07AYUzyBcv
jlgLtSYyEJpFz1/q9tNCPhduu/k9/Q4MH/ziOFORSKcuRuswZfj5OFPbevqOxhgjkAi7QbZWG7I/
4eSEmWB1V8PhkxhNCQINUS/R34CmGfXkFcj0toAppL/RYacRwKZApNpDhoaEbpRtIy2eRgFf664F
Ki/O3Ur49W2jPNwqvUDYzbllbp0nmy0hSxiC6su12JR7QuD08zM8Q4rJDoszMQPc/j2W5ClEgiRa
6yQUtcllnFmZmpq4lVfirxHHs6nXj4uPaIDe5MFAvqn0d8Ogy3FTnoH5ez3wy0THCBJIv13SEOwi
HiV2JvqET4o62lC3fPnt4yFOlBH4p79kV6mraN28hPEKtWFJz/1GTkZPhssDhjW8ti7ErUTxd08H
euT+hrE3/WkX20xkzY9JLOLlndTX8j9tICYZwET3Bkmda/3oTD5FoJHbNMkCfaUCOIK6Dc0o3R5S
fQSA2o+noAplJ3MDpN9gpvexCM+N2ASrmIOg17h4ccyWIH1v3cjSQr44TlrhLWq3/0N/qqHt7aMa
miO+3F2rwA3uqzyNchEnfvy8BZ5HWCUF2zGQOurktAJyWKathSmekl101/UE8lH6hmie3aJmg4MK
uEoc2RuoFeuCok4MAWlVRWxvtI5/WgaobGXCCK8BIzbQz5OK5KvWS1saE7siKSwozUGU+gZN5eMl
ekeQXpvF70W3YdeIVhHOMc7EDfqGRNCoYevxO/nTsDMRhIT1l8plRyEHEYksLgRa3GmgH8dtJV/H
00cZBuHbNyza+KVm/xWi434bYglK/3NjouXV7uPxwKRBaxBO1u70zF7I9Jc0HlBUeziIRbIz6rMh
XvCIHEhU427ffln7qMFuNoqMpa41Nv760zUUgpJpfoafS96dhNxxzSBEctapIVoQCe9NmWF27E8h
LGvn+TlPYZm/Isw3oWqSVl91INTZn4ejT5XhHfo+qBqUultZZs0ht4fTlpof93KBdc1a4cdXb6Ka
fgs31TFp2QyQqDvLpJNgUXeE/lIH1Lw+i8zZRg+B2mmo/hga+I0qBYO9101QVYKG1FMFhLEYuQI3
K9rAIU20msFsxA0s//sB7EDSCB3StikNOXEyI0eE+glplsmcKRCv7syjsxHEFTFa0YMpcJsD+d5K
98FhFcSiSOIfBUfTSFQVnw+1D8oA3B2agozvj87g8GtN+rYzszkuKe/v7zLCKfwi3V3TmgbyCd6/
Sk0aok5oHGZNzlByLx1uZX1aTM7EGQzeD2z42Zr1JEGVk2OQqCIagAVbUdgPmY+Sy9hh5yj1rv33
LAtrBSKc2C4BCf+4B8AvdW0hTnFRuFstEkFFLt0RfkKjVwKMith4OdyiBrHMph0tG5vvMbf3tCJb
8/5lRSqPpCd9g9eh22VdiiHjYoT0caWrknG1r49NlyfjVdUnmBZu1kjxLHC28meRQiPwJkt1qAt3
1e4r+aPUfiDGzVO21rTR0HKasQyl1VyYPgy0yUWIWQW7Inj1kjbs4TwVyrxzRLVP3O6a+w3sybdh
E92od2zH711bumbaoYZETv4Al8yL7a2FowbOGIMA0lUMp8xMEUk35ao7hWhTUc6VZQCzf+/ftdhq
1pNMKhmWok8sSr5dMe6oFZLxIxaa7DdIfdETdWVaUpP5CA4hWGYqD/g91V5UV51Ljj6JE5pZaN4A
jTubio8sKYSjrAiWv4Pdybv/B30Ak4/tLIRqB79v9RUahmSyH52c1YR/5kHnUSUJgiVZ1RkyBU7F
4vsuTbd+Yvh+NRgTHsLbclaDiGrwwLKj1eLwjKtHS8YU66tBh9KibeQetNMgyhdyWcGloIEoI4Wy
TzqH0wWRQGkNgurDdcZz64nJ5jK1mvkFKIDoJ+FmBnIXjr0TjHLodiz9JpjQmkBz0yjPz03/3XOt
0+NidB7VyEgLvA2WBzOTBTx9s0Zu27/ecwsuK9zBmuz5tDNlfsAxKMU7KcDgvt0NTgtghk0W5IZE
qJfTXtVqup2exYcipKGGZrIIbTOiTPDOrX5rvqqy4K1tujVcNI8qac5yu7I49H0U193HGtWsq8z/
gwtcWAWLRNkgDRy91liBznAG3L5kJ7wDJF2ABncb39GkBNH0ik5gbJ4DOlSGw/U5dhDukjQqEyRh
+7+57Zf3Abe6Mu7GYP5AERy1NjrSuaIIXhtbCX3ptCy6Umae2nH0CIpKMXTwiWI9fesTMtiCqCfK
Wouv6PaNiuS0IncOgFlbDqDtMEPILCD9cRBS80vzo0gW6kx5lAIGfKa34ZveJ6cbnlhhXiS8J+z1
b2wMlDBpj7NxFFJ0NjVyasEaRQQg4UBXhPV0IiOQSWfU0PFOl4mzX1yxXBd1Sg8b+ILx+5sUxdd4
1dUyt4cveYbfxMEFcuZQwzUuhLo8mMhJtFyX0mKWAV8FFYwdAnG/pF2+X3QF8ZJSABefV2NNXjcU
I+z47tL81C3ff0FO3WMxeGZKRP6KN4V164bS44mX0fD1VExThpEMxoUu+QxiXilj2oQpmNKxgldx
valdF1j8SdZZWyWlRVkOPP61heTKSrZt38psOClWi7VC1sZmkgD4+E7X5Y+bOTbOjMQ7UueiPyV9
sE8rDHWh+3AyJnQPFQcX3iwRmP28bYrnjNDidAArzvS9Yeg1deOcIvDdJ+U8u8JDGW65x5E78O/G
KPQvYFJ07tbIWIZNj6w3W2oMc6UMJmvGFy5VVFi8ZZd2luTzqmhxjkKu2KX8K8v9pBbrT1eM+4mx
Fh4XS0jViwTnc1cX++hMFUywRo3KMYQTNjV+XdTg+8WJrqOCUxlKcigWxCOjKC+gal5rxjg7t67q
B0Eyp7TVwgNs4ms6yoDkOw4qDrvxW4YbjYCe6/M7Wf7O1v7zGdS/MwhAUr4x3h6Msx9YFbUd1Ywq
l/8L12MytnJN6n+hiKicx0GrrDd9mEkE68ntH4K2qeSV1NwAOCQHwRfbVOO88C82I4Vk1r+nftgu
0gCWmncHHlDR12zlLbShy+cHl42FZbSmjgD+w5HGJUvEcWgGppjB5mzmZh/V9Mz4/bNhmCtc+EG/
vayAgKlAfKDTRWM7lrI+9b4lP3Bl5jlk+4SPss+JFVuKdmgFjvZmV2r2aoOOHTnug80DMic5wI+L
AqVhY6QXcI9DHB69XI2VSmvOfezdSS3zwXNx9i4xL4jEjPd5HgNWK44vIBwrWKK5agA1yZ5W3RYJ
Fy8RK/l0QhH++3t67DHnXF30eMKeYTf69K3qpAY4Lc5A9wCii/61TFEcOgbB1WhY+lYuUN7Nr+gz
Fjm39BvzimX9E379P3P7lfKZn34riI8p3z0lYsSIGufY8p9NdTF+cVsEo17OS56DFeXFM1vF9qT9
+G/QaZfc35aCaeIhLIqdlXACBJcSm4xMslJ6zlPzIQ4NFgEJNhfFl3h/kbKgBVNcuH561QPR0mTa
KcUG3Oi01IyJqBlOGF+/+GSXIM9BcSjphOk3dWZhqNdwCvuQBn3wRt398hC12EQExq57ERQJgKZn
wSIk6mEz4jlRafsXDCnSBfH2ikgxLi3wdkSgv5vWHZahvdXYqel1cATOGj2fJlXWzb5FufOl9IRy
GVS95ww9deSmTANengBplilLixAo7jffm20Nw73R8GKFt7hQJealiUJgC5aRa16NXxQrr0DrR67c
V3Ugmh49tqIjVfXZr/jY9QXtC+fmUcVJ3aIQP4zpdiil7AMa7O5bCSKAgLk/mzxi5kV9EIutZ98d
GZT2AlAR0+sKe6iVX2z1DHPY2EpvdEBaGrhrreqt9hkpthyThKpK+6mxXmv8ORA/vD+6G1pFhjPx
9JZ5KK5gqPnCh4xAKT1zOlSRMvbHWfdxmz8aBfNkFVWHpG7mGhdGu/jbyH7lSN5Vm6a3Sdd9LpQt
232GbQCgd7A0uXcNZXc8AF/gNywS389oRT6sRJhGAPRMxNoiaLeD54OE62PBFSnG+IAyIgbeHjQw
ca2ol0yF2EeWmYMCJA3VSX5UmTSt3WBt4b/NUt3GXecHpgtwkBFhV3y6S0M02SpKRDhi74eEjQpr
axi62qguZqRaYDNSZK3koJXZQXH54EcC/KV0B1EOo7ZLR28NQzyB6IWcZbIJfMKAp+r+V/TrnNhg
dBBfMFtdTJZJsriLto8XIBB5nIlL2+pIl8BOmB0FvO4C58DTEyUN84Sb3vRmlBBtzLvYBLTMpkEn
eDyFbBqlGs0mzlp/rfCYbhAPOvhYFcd4UK5PLhLg80TeJ1GWbgPjiKGMF562kGJswkpfXcwrjBb9
ly6r42sSP7kiyVz39ZbhMbdWEzYSHYcJf4iZUrRfdUfZ5R5wrRQT+ba7DOrlY/ljAoqgnBFnm2lb
WT8b9JW6K/ifrvfGc47rV4yGQNKvWDfLiZ33lSg9JijBVHzmDuqwl+AaCMkzLKeyXF/c2ImRWy0o
O8nEnYKyeQqs+8NAjAgVKXYwkXthDTG3937kKS3n76lpxVider/8uIIxgrxB+n3ET96hHpy9NmpS
isVnw5Yaxz2zVNqdZ+8C+8fAkrShV/UggRD60WNzNHxBETRXbD+ACt78gwjTAaJ6thJhDt5YBxQx
G+THichh4A8HvD3JQbfmRSCbjZ5Ufl1aoh1uGCvpleUuT3COHZJDGpDA0vZ3M6QhtLbICREcHho8
nq/FoDLKJZtDwAS2cVuAlMl3eL12v60tT02tvQDIUVYB+st7a6t+DncTa1F8m/8yK0T163prABFM
2M2PeU4y2+pVANhWcsfGhZjg1e4Hc98E5ct9xX9NXfhrd5cGtolzBv7DhFa9gkhtXnOpLL+mxDQK
+wiNEPjMKcY40Gsy6yxW+WGgcoGAjQ4XVcIRQQoT9tvg5wQbf5OlrQ7d77qruixGATTIcW5XmnQq
EFgFVSJWxD4udBg7T7xmbkJ0wkP+6Y/6rMO//kHx8wCtfkV1hYwHg76N72Ss8EFQ+pWoaWSfTc8r
mAhHWyYnaPkuOUEjzo/6ZV/uS8TONZ2rGi+n5ni/oPJTbkMkrQSToZiJhdqvkolvKOGhKmLFztk3
ZwwmP6H5VOZb/XS/PMTfw8nsdbCW1MdSo2t0EW7A3GC6gUKs2tVvPlRUpCvc9KZMpRCg+p+Wx+su
S7IsK/Cta1VD7PXjR4ymIS9hgLhQ+SMgYlbYETbQCpEFyfMewoQKAFbnsmM9hfoQEafEc/Xgrhjr
V1Adgv9tZY4nYTaYUdYKZxT2/qWi32My9XgU89A2/m85tSOGJ36prsPkpoMHKYs/SEKM1haGkrxg
yusRVxLU1Ypaksv4Gv+0Cawn+DNeSd3JjligAdsQqRRi/RRXtNu3LIG6eE7irnyWVquz2oPU559h
0CMTxWdOfPXzR1K67tBGWclNkAczuWHWD8/J84wHgAZbasWMG16otdQdhStUUqfBke7O+Wk43vQD
RvsReBvkRul+V24M8pe8hwRExOiDsvEYWb0erGO4/w49bg5fOKLgspQcnd6WB9ev2/b320+U4fZ2
LPwhVbVjttltwGqnTC4+b1UXGPv04RuiWBxG7KwOobQwx6pg3KRc1EKqEtOK874DHrRLpz396HDV
hnSZeGaaPrA9Xd8lmEKbyNjGYLfK1JYITpoP0uw0Ipkwh6/1oo3MepBtHh6eXrAgLBw5h5Q198Ia
c4WPiI9rsWCnQYv3IUyxWV66Nu10WqIBT/dg/6K3hjism68hvgi4JfrwpD91hvXUKQ1+sE0apEdw
BzWI7452jQEHjZuD3chxu3WCIdHVOuPjAfrqkkwVdiSsy4UvE3iN6gSog3xREpj+b+tpNZfNjOXJ
w1fOmGcKTQx2kCYwuTq8Cv5FKPtolZxa3/iDSp8dSADWdPHSXDniypT6kqWsxfg/kBAJQ0tRNzT9
4oD5ZtE3WCkc5VcdeF+Mfi/EAviz+Q+5Y8FGyC0uwaWPWAh5uwejk14s6vo+Ink79GYGjpVjvW+W
KddQJISmJLpPefm2F41K1Y0YOCFKqz8Q41FwdrQ2z02Il+OKd/wXn8QGxfXRtkrsRxn9leEpGln+
0P1J6JMI6pTuFBs9M3CX/xGA/9CKncegsoQFMAeVcwpi4giUVT17dOoGFmvvgBy/fp/Cr27kV/od
NR+2EREfU6wttAlsMAheCrFdgu60Qg9Dt5Jym1KC5FMdr6x/Ff2Ak95TXZa4Oz6OvP/FQY4uA/2z
Uj06VKm92j2mpEQeCKaXK69zyh9Ty/VoVaO7/rWU+ewHmy+ie+taRlGL34zNTH4Rg6Mj7s9RTkyN
l+BVPpMGk9xcU907RvyG3nAR5mnhDC5GGoUL3NTR8Je9HNIFyB/DB/UjgorgWaK8JT7upzlnwMmG
LumHy6KSfBtxSavGS1UtwE4/vQyr6WJAM8TBwlroNf+soEVt93VUNGSqUqs3yuf6T9BjJZr7wPnc
cclzrOv92Gm5HoZYvaiLVhJEJf/mT4Qk6spyeDfYMXXnsvBsv6b4RwKlWZ3Bg5dQRbnr5I32s1sy
3fri51A03XSJfmCSTJtbgYQM7hHaeHxhe3GP3g0DcD+MyLK+sdtoeFg3StcXOyoj0v6KYkr++Qqe
hB4B92hCtf2htId+mFxg6EwgKVMhHedq6MopozT8gPr4jt+CGafkStPA2TZEv83GPXBcSsQ5/Scc
MmZj2MUPxu6+AyYH9Tyn6kc6VHOKkAPkFO/SGOzzpK8rqCE/QUNIGzCjqfr4i65oR65jBvOMcRUR
gjIyTl3lBg0EkKqMjvBMIlUB2ECFrVSzO15azYfNUlzb5Mhnvyfi0mHd+LvDPNpdWKX0ic5btQ48
SC88pWk9UGV+syCF4tCsGs8OAO/OLn0xznBSDosvb4AapQp55441rUwZ9mbys8hnJVfzPGUiocSk
lyv6VN4JX0McWi3PaLB1mog/ZRYJfo+iun3JF2ZAYTqowoZtkhKV0Uo26gxueJEzmcnDGH73BALj
VRQl0mf4FSc5jzfK3CPP+CDssJaiF1hD+UbRipAFtuKjx8kWXKidipZj4sXT61IVC325SCZbsMJm
8YvzF2rc3DaggqSWKOgSvAJbFgGAIaIR4H31IyXFX1JBMQeGKJZbh6XBs72IIe2uHS4X4Pf7Acwm
49G8utusH2QhCnK1RlibjmZXB/2DYeGzgUixHwepG1rJsVER+akUtvCm/TqxW7SREXy23v60sQtf
1FNE6D6hqUcSkiSpVx1GCs75/xc6De+F1ek8iUAjcUiUL0zgm7kTr+cIOY6sh4Em+eNc1gJ/I7wg
o42YHIITJ9ZfbbHQjLlPHC5jNIZyAkfFjhqGB4qvqUmwinwmUzu98lO7UGmw4oFvtB7JgciSYLrM
Zb4Hzzzhi4b3ESxGznvrd6RIzTjIiNAyvEXPXKIHp3WtOzSDZnm4WXA7c5RjiReShAEj6iNTmDUW
lm0l2RHoS9zi0kyi6BN48m7NMePTXhWV/fIDCcxV6lzQCaORyvqIBlzxbE+C2QQs8Yy+CNlZW56v
Vz4tW6IdmQkUmRYgC+fN72UJnHtGd6CAsmj5ZxMJSj9eF/bSMhLB7VkxScWQ5pc+9p+ZZdmOF4cj
zm7TzdiKiEphFMytNMSN5I4Uj0/7wUGaAiasSANdxMt32PfD0mKryYJTdqiwhzPWiftKdj1UNr8f
XgHniuRF64Jjh/pgSMK7UN1FceSDcgx/rIKNeVbWjHSMmS2dOauVKM8lF79jW53uzmnAL5uYyUen
jXyGXR3UUsb/Otd9oHEgBWeYnq/GUrgqrOB26yStANBWXlcoG1xOABJiamoFeTRbbJbNvZiSGTIr
DvA6cvz4AlV05skt6YF8tyF2zMCqjSVxRS49eRIRQBRUBi6pbkIs2sEE6c3RvJa1FPaPqw+KRTB9
Fm6GIAbitH5YVKLj0Vd1aoulipZSk7u0qI/SBMC6mhUeJv07bEB2XLGy/jYj1P6HMtidPB/HJeAu
bnK+eE/nRgKV4bSGPx3Q+lZ+MhZTab4jy1dehZT17X7amvE+bONZ1hTjmF7Yd5ahSAb3EKD6RAYi
cXjbsxxRbOtooh4bpBj/GYeIOjU0Kku5rvIYZuYFubjkCKZQNvzBf+i5FRrPHDqBKvUDMOm9sQzp
pRFRbVHRT5TTdCLN4GoP08bn2gqLM9x69tK7xac7iK9PssVf/JBC3rvpccXZ61E2icE3S7VqoM7O
RBLzSLzVh2qhQNs3GRkf3UAuyPCBOtzzc80deLe57rv9tw8p/PTw6GsZjgq6EXJSBv80vdC2+/Nr
oiNGTA1Z2pv6YGL7RHzKq0ivroWX8gjN8tCyONCCeFNhWcE2QGuNBPl4zifeGUBfNzPRRibCHtMd
hI8/G5w4o33HpHTrjKKBhQrhT0msRRhcVr6r4Qg/zkic/sbDZvKAQVzEvTxNwKHBkmFgffdiUxtL
lX+wENbTLgnL5LbaB1n24l1uCbsoSm2yM9M10CjdJpB5NvoxMbuNL42bLNkBlzZhO/k5F2rYVgdy
z7+Wt8xlU/09BjKKIiQeZ5lxYfxxB3zui57R1HSrx5xLo05KGz0C2FvEA0xnSHPCuYtApp9y1E+h
xEIR8iH4lyMQUtl5k+5G3PYsr3IkN3jxX8y1/79YbINWJzj4Iu/wSX7nO8k3WS5vwaTJhuoAwBoN
yNbr5aSpFLW6tKM6m7w3xvMv1/09bSyizSeY4uSI4KzTXB1EmeZqxReqY9Q5aEoJahx8vxK28KTq
PsXoDzEZrKPuUp2oyZFXqS6BOaNqv8+c08sV5xKWUgThP7fJs31WHs9hi7pFW9IhqRIKjLa8cme+
/K9W7FazIOpacsash5WTGDWqn5DgqypzBHTCkG3jmgaM/yi4jOsOHofXwazA5Rc9fylLewsxlE8W
clDHxzmv9pOSkLGILp2um73IJ79Tkz17ukxi6Ph+SjlaQ11mqcwGy+0UdBmsXaBnq+rjJw459w35
yr0DUFpPA4azl1e3jTfW0V+cYVTgSJRcMjAZXxMHJF6e1ad/fmEyGMMR5KJCIP0ezOlhCeBbNE73
E36ijyBt6tnmJGMpIfhH2BRKc+t8ywgmcA1jbKvK+aGFSXdPqFdVL0BBNeSvSugThxbOV2Csidwt
MZU6OEEHWbmqyO8+4/p3s2VL15KXSDASeibR98LC5Zlxj8ImkTwd1y0/af4rTPCDCUWqSZ8FZGDN
C5JGT4wGovqPmKTHlimIg5jp+x8iEL9kcRMWqqFpbfp/ui5sJzy9sturkzfwSTbHPk6Caq+QMzjl
pZD/1+XZ6KUa/K9nV19rKQQb3Hdau5rKGo3G3fO2A5xzUEIn3oQ1a/CVVACDAHEyY7by5K9o69ip
hc0/RINIbJZUh7DPg2Y1bjJjSHI6VpP4V2useUyFY4o0Qhgyxa6/zNemBP1/vJvRcYqAf/tm/cUY
Yt9YqxNCFCfIuwEMYWdOPMRp+TciYrkCHZM5FUhNqPjBcqYmaLqp6CsgS9IhNgPKAnng0FlWh116
ZRFJgm/cfwuO9jd3NJKVZsgS57Z1FfYxyt5CfPduYXcgmefK1WCxdrE07KHEJTWK1p2tFPLrWAoL
KVGRDGINKM5eQXoi6Dbid4c5UDMfo+3zZK30hBgBZjZUTXyJCWuYUb084PTbNyrjggUBDYwPsmLY
tpGgUGP1psLmXp8ZMk7lFVLnTrkwkDc++rq4gcLCYWxrQCO0SCStgd49OdTURFi1YCNNGzQZFBWl
Ii6hSJd0v9CqaS4ElkW7xL3JgaaVi9Ed+IfWx6naO0xkkhNZ5N1SWL78xUVicf3i/sI5ZUSgxgpB
K+DnIJRVLH/ZaBmuvC8w6RNgdAyv8dlOy+FCyht1OKzjqtN0M9biug75BAmIXcgNKl0jlZcx335G
xfCZvB2NpV1oM+q9h5vs9ypzWoO3uu8e7USf/qmnS7+D3x4qGGV6rLx/Qxa4N/yCG/qX+x7vRnZr
NVO8ClbIAnA3sNEmlMUpHqx4bCFm1JrL7PEFakZ6C7fduencYXybmzdM7wuutII0Wy35v8ziLR8h
49LRjGl1csdz9hb4u48zk4ViDZTwmhyJH5nYj//+B6SHIt4A1REzdTZMkK4ayhQMxZmvqSbrDdf/
/b8dDhIMbKtgn99Lo77uwPXxLXG8GbDC1lutvTXLKCe3vbD1VSP5VOqrD2QRoQxwaTOQm23Ff+Y6
4DqlbgN42a2yj7R2oj8RL0gNaN2zq6Q++HllBmIx1AthjJYNzftDxKI9iQLyp2CwCByt4tcLckG8
uJkzqp1+l9k1j6x2bvPqIwfShAgmybE3eUmdKGTz0wgBnqIV8hQaG9MscUUIeLGitpUJw/w8/2IW
n25uSc3sd4bu7BS+UMi1k03SmhkB25295Huu1O9YBSDlG+As0wT35Wh+QfysLhrf2ivnYVQydXuW
idID6NjYijbLHR56eDoAQtSZYnfB0wi4NO1Q9W7blzoov6gU6a8g3mQqCMGqgZnFCkJCfuPHLheo
hP4x3VL7EAbFAyjo5TNZ3iGn0lJeZ/mawhmySmCA69ndTEfSCnH/sxDGMCgfhyGp+3N7BeWFNyQH
VK4vE7eDDXqJQhKLvX/xpnW4ROw7m3hAnBHpmG7v6wouS+VjO1R57YA+pjA1wp4NxQeCDcbgxPV+
tGXymJ5pQVaXseLe3qQWfY452yhpohD0yTtpKJBjP4Y24J/durcFfgmO8Ao1Er/QrFWmu4XlDto5
Z+cyeLb1gKyVfbAl7d4K0ZT3XKyM0Na6IQCo96I/jxxs7/6bKm0CXuLxOzHK+hQgQxHg/FogdQoC
APqhJDbYXM6DivmzSJPbKZVBnYNpgyEOSPkNzKhHkpuwtKWnIQzSFVjrzZZiTmjTITzhroO/6/DY
FXVA44h6MHREUviLcwlVfaFBXsjze/HSfiTJc+t+Ffhk7+n9JU+fBZ2ifQWCY/51oRof8gg07Dk1
5qEC6psLiEydboQoQAda2rgBOe0QNeMUrIsXEpGDKJ6nyWrXGUcyK18YvL/5vD4BTlaMs95pkIpD
hyyoScndUHJU6cq+p0+IoIE0xN+EbH7hc/kJQ2eb4MrQI0Il5nR+f8UoarylCLOxrqzZHmIAcJhv
uAMqRJ6kaNTWDLFdr1N0BirexlCjwz3WMLXYLpLSh/jf2/Xgsbae4FpTp52sxyehVzhadXyh/xh2
eipNWwxjlSbAlLtk7LWNP1EQfJ86D6N9GE1K2xPwfghdul/yZoqlkfoKQxZMEfmtwXRHjfvVtUKT
lxOfk19ZrM8nXulbCu7yLlou3+Ob5Zeheul4SqTh9pprErEocJpRoxw927BtHpFHBI7Yx+7b8Kdg
AGWMILVBBLYCJVjuqA277/S/wIyVZ8cIafQOXkyEdmfCoc/vtmjPBFf8PsTgS3DjJ/fRqsaepyUq
mm5rv4XyPwvA2A58/k8HQM2OXnlfS9JFYjd8dtLJaDhv++R/f+NlsZYBjmlyCJbG/3WlCNxrQGqz
wCkucn5+O5JePvZjNyF3wF/8bfvIpVUqg9VRvznN0tWTr7nzU1BjOgNgUZSN3pfy7J4+FFKazvFp
Pv5k1YM8EfG8WQBl4nQNeMQMPmM/vfmu4j/iMDC9qXnM8Mo3vVOQEnQZTdGImukvhrAdW5BjShuL
0TR6s5la0G8+hVYsLrghYr1AanZ/Frba+iBv4ojUA9Mr7Pm0Bb2/9fMn/trwSdprgkYqjSSQVIMO
G0UHSeNmyJ+KY9L93oGn6yDArvBbB01YT6AXA3NqyHdphahrkuNNGZ5jP2bklAn/VITdGyt8Z38H
DsZEWRXvzjllKDhJ8SFTcdPR6lvbVvbV+r/15HVtHgz9ZkNiBXSfC1QCy8mvrk1X+YhyY7qel4EK
peBgM9ZUHN5KrwCqjIhRgeHPdj95++6ndv/OOlij/3SfedM9EPUbz4xnSOF4Z+xNPYR7dz0Wpkgl
QMp1oAh+sVY4OnJ6KgVQp1Oug5BbbVInj3gHGw86sJglJqDgnUeT6npVYFJl/xZZeP43KKgYrZFi
8LF8Gijop7V2CffPZAAkB3FeY7JqKEaK/NO1eqNzB5Ih5Nnp7jUNlw68RfVw9VtxWK+6Xq3FoQPV
xX/7FI6IWwyL8kSUNhS+AAtDiiJR+wL05Rp0BAdlT1UMCn5aPFhE3+zUoRQZRU9IISMnLNx0uREs
m2C8dtJ2Pew9TNsLlpjBfVgeFIbAStx5bxZhuRa39XKaw6UffevmaMXSev5CJq1J5y9ia2fQxyXF
RZsElIPCgWsPaUinNhxaCUpTA1kzmRE/X+EqjI1fBL147uib7gBDeomZ9AOokMHIteGJ5T1vLkvW
INTKQyBiznFhR9KjTqdkM0PNA+JGA+hEPyeYi3GJQnxhjYi7jl/MzLIVj6CQTrMekd+ZSO1PLYwZ
MXgh256ZS6YPZcWQuYve07Xksd0ro5zL/XH+ldrLld8nDZK+wQh9+PchtJWoJ7uJldTHefEjVPN5
MkccTzAf2uvxsefq9xpxrVz3W1WQd6td/wIpKw+7DU/EfftrOzeVQFsmutw70DV5O1Y98zJ/mQVc
Fja6UoVtAPlfv87oI1Fhg6rDU+iRnMVXQttuj99Keu9x4B3x+g7SWQgcGu7q/PN9oC/uiRTpjEqO
PzAsz/V9vAWS2vlHrUrvj1Uw8j51DrJFKrIWzbt+ksJfYcUv3YzjnOI26IBMJHZKDznhX7bH+kL/
z9u9iJ+D5Y7EZiGtAl/TdQWAWydVm1n/atIe6hdczstF7KWiBXqwrQqFqlWBJaO5jmsLHwzmvz4G
PtddEMHBf8CjQVgG4tM3EQDuurFOOp9krk/KbkbbeJyCxcaw8H2adHYS2CcgBg8W43DcxGuRI91M
4sIsZM/PPl/l6PT4E8HchCI3C4pmAbvDiYcSM6ItUl33CXZHG27e/RNBVklcJZMybBteAc5NXs/C
Q7ACw7fonJteizChlUFuRLNxJ1EXTLEVJsQCLshGCjKyzJ4+iLwSosXpv4ds4irGT82p1UA0Nh8b
8M1bTFeIasYWAC1dppghTLW0l40gSv9Y8bcdTpcycad19/DTjkO9SA3zPRw66RA224/TTEk9zuDx
3mgO/tYFE4chaxFGIh1zwDZqf84WbuK775akxUMweS/dDjDQvsce82rzGq2oSMaJ3gCScH/TYxhS
1Mk5MDAz6PXhK1wWEuTZE/JPUYFJ6ldt4Y1IqcnsJ+C1gJLY2YCvsL9y2HczrYHF4EGOBMa0z3rQ
OpD9wUUXc3ZOnGZR+fPR0h04SxpPHAAW8uhyqOUzcHbZrsEZyjDSwT9OdGTiU2GJGFEr4LhmgVym
Cs8RxPCbBVxeoUrSpCsQbu/zD+xVUmOgMl366FCe2sVTA84Y1cuKlTlhW67cWEFvwG8rcIuN3I5e
IfptC8E+/F5wIKYtAHlt2uZpXU5cd759QG4qi6Vi8tTn1ZJsQEKsvZG0N7JEoF70mOvILdfXad+9
EpBXfKj0Yd3q5tSV9f6eNOUdg6Zwci6lUm3qV6nt1u6PRGGgv/FosrsO4aENcMGatJwfy4FaWqIe
LZQp4nbDzCQO1Hjkzr6vmWKsfOUTohfU5bbBxy7QpGMieqU+9wafvNxkyVWL94pN4x9DD2BytFu4
ssISErrCkBsEc2ZQV4jOtKkLXHEsMqpKAHBw8qr46M2U99ttuMHD5n/jtTwYRlbCSPKUXPpugfM2
UKX1aDlAui0q6xNv9aFIG2Iq/CME2hZGgFZ4h6vo4u2ANPa5KmjAtawFRSerHiW2HGxigfOtydDL
hrto5QPuESL+I0DlVVQ7s0yYYsIYaUAqzivq/JFAR7IxTeBPcSxLsn8re9idMZYQEaVDeiD4njBA
LBHR/E4mnCgN+hF0w2KetIBcyohIKoCiGJlbywUMMU3EFTEsc29PYIK8eKJXlqJ5cEuNQuFWq7v8
BeEJLDK5/bxDam/xoI04oqPAbiY1cDQVyO2SrkzLHq0pAA/zwPiJUyUjOzXj+GrCzoc4sjiGCu0v
a7+x86DrLi/laNvXto/sc8F+Okn42sR9nLqVBZHhBminP3V2bT4rDSZBrxFaqZPXnM8dn0Loxl22
Uc1j5Wqu96d+PK6+UQWwSwqxIGfNw3gEbsehLocp1NrWv1ulG02X4dmxLGweIgacxXBcjQxd+G44
S7TPKF4FHTJlfx5xZmDntAUik4z8VZDf4wx4DAKQiZm/8nACEXDVC/qQRGhD/STMHvwkatKEiK2L
X7JmF4REnA4w9CK/h1ojqeMVaG1ZzWz2585WV9xmH/rLzqaQwFf43pk6cpnHGYLb7WohSOh1cUAy
cGK0vpqtR0LRc2nESpE+bDFnChXgHEqzxVoY/sxusP2r4J3DHL3NHTiAQVziUkao5HzStlhnxVSj
cB4hES5bXSaDA8f8arRcol7orRyJwkyLwCI7vzJnO5VeovdV12eppf6hAnS5Sizu6TCvg7lA2LWf
C5bHqPvQPS+9Htz+CqcqG3BzO3ezO5xdkvEKfZA+M7T6hNxdimL7KDnWkDCcvjuo/kwm9Aa9l/X3
lagzxwsRBPnR5i5E4QXkDsG+eO2MihYumOJpkT1shV03YsSsJT+oq4lqt06glNuEXkWgy3XwgNzL
zsU7cwbFas1lUDD3tnWlqfjiGhehO1RHJUYQAVXZR0btmTNLiBRZ2ealzy+MjT3umkudgulV2R4O
XD2nvT9IQpNDzvS4Xv2oxy8XjWXuTKuc7lfZJ88IYeyjIsdHk7SzzTJ5mW1wyeXszo8rjVX9y9Zw
0HM7B/Xtc3EWKsy+gZpOcc9Xf5YgR18p1cDeprrdjPlZfbeZseGxBDUdrWWca0aqoTlyRcOCDXCw
hxHQPy3/YI6efFHJgO1RL4F3v0MYbZxyj4twcvJBysKoYfOdIyFag79DlY0hYa/DoRBQvRoYSRTT
Be/1NxgCWsqcw5r62Q3zFt6URLEJ5pN7Vi8SKveJCZg5mGVVaXZ1VKK2QECWxyZJlkObZ7ncckJV
ancxBk0MHAhkCCyL2qRnX8reI/nJzjwl7dMtIaVeiMPKXcbQYw156ykRPXdU8fCB0fh96HTZ0KC6
k+/o7FCJ+m5Y9CeFnNBGQgxTQS7XrZzc6b6SmdkG1a5Zc4M9izP/EnYt6+kRh75s2LY8hHP1YUrV
2CqP1f4Cl52/x8qvJa2MrHjbGSdDDcL+i4gbs/9shq4JpoPAk0+fKSyIAHjA/bfMtwuAMTS0DM6B
ALOe+ZhqA0DjKtDB5yWyzvNj9MtGY50UR6f2r2k15z8QGVAR6FjKjJzBnT/hgEwS7/acCAsfagpV
o4By4mPj6mYnZbxzALkD8Rk+nQiG3EJFsz3UvhFgQ4CMcem25Hke5hlFu+du2+nmfG7wLOVQziO0
DGNLWImO69kOgj+TWtDPDs1mkNUAfVMg/1X+Mu7MqrHGUeVhYWjej2SxXbJERZvkKUD75JtjQeQt
deJsOftapuNZe00RTzUM/CjH5arp2DSjtYC3oOk51KsuBoWhCmQ9qjmbvG8pVIJksfj/izc+MvlA
39v0FyL27xK1sAfbNwY+KDE8Tk7RSytFe/8jFIm1hwSKNAJkPsWhFmHVmXXUh0IY2KQHbUIzkcLu
ptjgsKUjRfzUjeIZEaofD30gROJK9W9mICN8VD3FumpPimkc8Uzzi5w6cUGJNaVRyoYxCOxRcfgU
rf20q//ZtfL3Fu7Brk3tNoBZN99g1CtKPgIfnZSN91OMcKecmOZJ3cAnATLksuthSQSiaP4RKTqJ
EhiwDoAbZFaz/b+ySUiSooFjfMtowRfUFBEtL4dA9WdV5u/kR5SyzOFjTswO0hhU6wTR9KlHjheU
X/CQZZWdQLAY3C4aXDgoA31CLATNhkKY6E9YP+EZxCW5/H9KjklPpbt7Aw0Z1+9GSlFHdV3JzfBF
e+UJLWzzeo/snAmB1m1ipWuh1/ckl4uW6L+6FmeuDL8OnSi0UyNGq5UxZXM3y7i5i/kzylgklRHe
v++tGWMt/AzovjwG+xxA61VWVj8ag5Oxkj3aVxSIoEAMGs6l18uDDy/aQvrlMlhaUtNr/rrcClmo
4WNenOndl29aTnmwrzUGe6RiP8+XK+6oPpxBQB2mEbEFlaiTcu4eGFGh1R3O8ESuDIyOr87095gf
3CLTTKTZCqKAwb47jZIc4y5+XPMKbw8NXmuY0otTIlwUCPYk2nlNgs3s4gIa0oRl4xcJtrz2Ce88
mzERi7WZLQ9EovgYoYcxwT2WWknnj3yuLD8XKLlH6lXjWMAfakTWi0kikg6LGVkJuNwgzJkGr0YX
hBMZD1sCMBFNKZ5yW7K9KqQH2pxlOpkc2nGAuv40YMCdOLBgMCnRgmK0AND7U5LbStrG5zPfCFOL
Ok45t86Obm7C8eiw3Cz4TSkafng5pwUv9jpZ++fqx/epGcCSkhkonRIOORrVUxqIilMtNXDWyFxL
KugvadtP38iWd37ds8MCXLK/opaMQnFQDEF5zBojAKu+tziqgHEjPdW3svN0GXGBfakIi3RRKK7r
gjSu81+YgmwwecnKaR//03KMmkJca38jJyin6MyqmsFcoz+S5qFHGwIqXMgX7wifGg2dVJXwoDce
y1OjOjAnIgtwe4/+mkoj9+2S+4+EN7ERWlSY72JPu4sepxgo8T2TajHK9z/srSfitDl9jZFwidpF
xEtyaANy3YUIK5DorY3BDzerj0kPJJLL7u5tvCUMV270DWSLGz1pB2l1nAMg+J8hlyQ/eNiRBX0h
phJYlVRjXUY15Noi1MH1t/dqTtOOlBuJ6Cyqq2zOPNviejLZD/35Sl706eXgmYjY5QY9Xo1PrElI
eStsnp1gsJCN8IZtF6HzJ5fW1O/S2Umq1sICwS4mh8X15xmvfCrF2p3nXZQFBzSTH845mBF69CS3
ak4OoZFkd3EF2QyaI/gm4CcLBQvylX2orK9xNGi+V2wddIFzucZcTW5XqckDJwlAWIKhBNRvP47s
1UxiYYqs3AZ7XIAScH80tQEpvBx2f4Qi7EyTQC3jcoN3gAIaVuNR2lcEQaoDbsXL9jTdy9scJ5qU
EK/U9ffqG7TnaYjvItvlUIXm71AD843iMAwPTZS/AZlHjylVeCHAgvwNqwsQy8R1kFF6JyA+iThD
70Q5cwcnq01ywZDfTCtIoBCXkf6h1nVZSMiHx6pK78Ec1Jrv0A0jDArdgLCl+uXhEnq24YTnCAu+
Zj854eD6g4myVFwk6zjOPxZiJ5PTZOtd+gBVq6jh5CUgA68josrT9XeEyx3rAQh2LUQ6NDXrQflJ
+Wm4vuKhymx2XIiDf+ff0+z+slnEPTtc8HKZMYbU82rQ6e985aGEyo3rendH5vx8L4VeFww+o/Fd
apLKUq8NMEijfqYqB1h+6bR6A1O2d/a8n+Hp5HuJkjyeT1JYXrz7owbtcxy64iDS5vhSbKGfXUw4
Wldvx7jSn7WGzSmKT/bKjiha+yaggcqMV0+3gnaf+2RBCs+2iKsOC5htdpt2aiBvNIiFTqT0C32l
WkyCLjq4H4VhfZ6XeWBTLpPXZ6BjrdIr0PXDnjxSilEaxhELojPBM5fDeqf9D3ZGUpZ32VbsDh/d
xrBoqsNrhp9q3AYxFC7OaH6ewQ0Bo+PNYojaablHeVHAyhNbHqH3eIYEGhMpuVgDQmrnO3iTDK9A
bIJyQYQOutVkC+DZ4G/JmL2O+iwQqTHelogUIsE9Da11EulDivJbDtfos+6fR4L9dso8U8yd7fb0
d1FNSUT626Yhcg/nRUQc01fSvGyZcftM7fwSYk0mcSvp3YxFCmyblCGKIWqRSmeYoBpQzwBhjiUw
n+BStd0YXpBeIatE3tavxnWiyr5a8ziLt46wo6di1boauSt11+/6YwLbr/pnEjxFrRZ6S38lY7A0
UdThBxkeV8sn0b6augE14/cnvZ7CjDclgtS96ByMM3P7NhOUpHAdBA7lN4ctsXH+LM1TbQm30Ael
eCxw434nNOM17daMDrwH2OtemssQCvnyMo2CfLbmenjGfk1YwZCMt/kT1Nvly+gK0ox9DTNNYl+r
CVg3EiqjiivDxuCVfLNKCW+THRjSniuTjMLidFIw90Lgh0Zp+pej2+N9qrDPDw1dqYeAm1iXFKYa
8z7cJ7VFEC0XLYF5n/GxunU6BDVDut/azcnV0y1mqUHr/bSaTLDgwxy1+mz7RlszwEo83AnO/V2h
H4/bUaCc8J0vPCGVhkYLweyJ69iPGAzhbV7a6TeCyQ8IL0JFz0d7WGwfXLVQZLsE13bJlTRcx3Iy
onqBRpm8URQpNVCxvw9VREeEMWo3utEa+yzRlRtHqVYiPgk2adWXGZ20O908QJe9WiFX+Qmy75A4
HusCUsnSlpknKrt8yk9OljzNXsAeMNIczEBMnBc3tB2DP9Iqk6S45UakIGEci019bFRvmBFL5PEF
yFNdg0yrc4GfYGNaO+bJq0IEeFysKak/Sxix37zt0rsDKuOxJQF7c4uqE8ClWEa5dRbnxl2brQuc
xYRce6dEiAS4mP+Gii79SJ4rc8Pf/XyBaU6Yfm0vbTKU2yFw2settxv/AVzy8imoLPA3AQdY1Zpj
r6g3UUytuazRXMASg5R4HY5a9pdfOAerSG5VRFMDMOJ3KB1wDNCRH3lR3DxPNRA8XmTJTcAe/UnG
RzyZ5Eek1H1uNcVhr3GNrOfIVHh+bQnIPlQiVjw/oFstVXHK7Gg2gaDulEvYXHmgFFTPyzEs1+QC
1EXbt9/wo8044vXsNofE/vP0zkerbW7e9rRLF91Hptn5VjG91ZJn7nOgWqNkt2MvmvqOdebKIx5N
yXXBZEtjMl8wLpmk9RPLR//H2Vk2en2YPsOnsyL2OS0W+dA9vddpfMibYD60dsoHiuKMH+MBdv+p
1QryloLJTcZTZ1CiLajq2jMfutyXtWItkfN3RNwquf7ZFRJjgOi/HYus7AJtzi+nH8ihHIn4dLTJ
Ks2ZY8XYAjPNO6+o5m600FzXtfM39+wznoBwtUF1d3IJel0jyvP1FH+O4wg37qJcHXifuCIC4DiE
dpg6j0S/1njqURzqWFrd0Iuyj/YPcFDcNQeEhRWC3Mrvq39KBbKXgK8DKeZX4Qs/p3V/36Y1Iata
FeoQJN3DpoyIIp/RlIP3b/K9Ou6+CUjv6agVgs9rFra9u5SIImRnlxlMwra27QjpAqgAAYPduAiD
2kKNBtLXOSnZXISPmrIEe5AB9ZcrCWwLYqJNNghudYwmMGkuGsdouoXuQQqCfljE9FDN8B56K3V6
daxTGYL2SkE+sfDa0oBDyRgmDdUKgvor02Dv38yzkCc87NSD1untIxrPfXeAvTyxqFTH5poenKaS
EXj0kojKNwFBu2S7rTC91bfcYuUOJOECKgKe0l4Cu76o67Lev7RXcWRFrr69RqZJCut8Iw9p7xD/
B3FytqI1kUUjcpcwtKbAOz1/16oM+wd3BI5Baq6DjAnDRyb7izWmEMm6bV38s8MOYYNyLpvPQxJl
LtrUbpepWoXnG9DI9Km8LbL+LWmOT502LP425jxDwDJZWf4szcSJYNozTlt1lvHxNs2QEHX3eubI
jcG1aZhQbVBb1AF7bz8/FNVVe6eejHx+YWeyLCN7N25gtrPOxhkVhyKwrihxBB97H0gqnyzkZXlG
ZsmRa8rWOKt11W1GJyXily7WdB8q0qbK8nm+z5Z8W60KVVe3s0SFOwg930E+xn3gCUOhz3G0dTg7
KaabzOECOfiFHLeppLSXUZATAhjYYRMZRAOOvBj2TSweZsq/JuKRdi/2xNVuqmSNfLrB5x8Ls1Zi
zDfsqEFZidsODPRjUkLHefQTgRUycLp8oqJ7UwmP/reFNGUg8smgwF4GVzDYUcp83uHV19im2JlU
OXuM3Py1cqDfbf4kdiqawPZDL4UxZVIwcDEi8Fgq8UPMR2KOXDYydsAdzhAQZo2cMi4FU5uuGTj1
kPntjc6U129Wu5+NxP6KWYqX+4GgVS5EIJwNMSMfBOn56mlrnHrxNXlFV4Yk34rcg6s9o8fHT4Co
S9k7LyIFkOe/tVCpXNhQAjAPHGOJi89FRL1ijG/uWTrzDYDdXayQ6p9mFYHBBPI8U7CdPxSdDJik
qzJDIDnbHPaaRvXvRwNPKrxktMAhIqP1ThKtgXfo5iHNN8OU87UYZwTtPM2FCvq9aNKrda49TZIp
vlUpMZk6icbL6KivNLD7nxiqr4PUfNlbJEnN8KKrnbvY1k8TA58E6jHp5SqTtw0Wn1SjUVepIhuR
W2K1ZgyMQByTj0zZSxh9zcGIzcIJtlgb72jt6U/Q6acU/wDzipnKH575As3tEnggZfrl2KXYlRyX
+i3bzE/s3kfZYHeNOf15pMFqZkI1vMLwLHrw1XcFuvSH7LKyySLxUVvMv70eyTFa9fxJxY3yJGK3
2nPRzLTQZMiy9gzJPTUrRDuYTmcyQf+Cv7CFQlt5wPy3KHHUD1DFhGSuvaLJk+Zir1u5bLRNTm2u
vLBlwq4ElAFfqqUsSMNn4AMJG8mVPK6/6/xz732Y78A/2GEnk2F0yYml8768jYZs4z/lDNwRvBb9
c7rIuzra5yhb2hZEOEi5TbPvoOFqq+4cez6iIkpdS7KOQ29FxNtMI/FFSYYUzf0afaNh+LIAVpLc
UEISptWcsNq4T0KqvFqASECW5LvnRJY8ugucuWqKEvKtEBBHnmVq/RQ2/qOAoHJPZqmtNQlrW/OR
NGUKNLb1KynZMMZYk+wrtTt17CNikvqAj5hsZEcW2RmcsplcxWmoVyusYTCbAFzv5Zk2XPx4NZ9p
Zf2zs90hrXDLtkr9lG9YgvUXGtgoz69t+gmtfTgVQz84KS5vb0r+esAeMwPSvHtrMWwo/SSrCp7o
yAh+trdre2vDUmGNiN/bYm7r3v1as6t8AP9pCqk3mMX+stjWRu7/0OGYfR6ptDyOGjP7mqtgNWm2
o58hLRYqfDgY3/6j4MPfQ+c/oO2ySt+VDABG6riWEfBZ5S7JZ13tkvFjS4G9+buusssVnNMR2b3B
mLMnAja8KZxpCpkbCpuIZLlBpz1tD2kIZqXFghQR585ibKrSX/Oi2eMYEmunzQ6oMSGQNgiRXfqE
Y7/MHX7rVqoAhyOs22qU9sSSqZvjP5961MIY4Hvj2UDPRT69fcUo/5UBx4Ja0/if1SVLdFI/KSGo
lqSJn9B3IZTkf7N4tVEOlSR/iwu5p+7sKgWzrhSUuEPGevjb/Vy2WoTe8fF9Dh1pchKY6teKa8Y8
8kNhP+arXnh/ShXkgGHdDBdsZVLBgX+tYI1lxCZ5PjxWr1GfyaNQ67rPBw3tRp+URn0TS3dDhnkp
Cduf4Dw3m1T8ODQOXEsSQA1Y8Z84sk3y2zEpW89kMgQoYKTDbMCP+xtFwv7pq+EAO84Pj1ggIbIH
/s9Hzx6YQg5IkV5nHKKBjrpV/dFYMyHDka4XAe6/3ptZaotxfzdOx2CdScFh5f0C2bxAMmIMJeil
I0r4RobbW+j+lOEQqjwkHyeivne8U7nkxy7D9RB7qzQQmj1a38Xz6TGAM7cKsBVFsbSepXUdhoHg
FyQlROot3t9DVPj1rRCCJlYQq/9ySAmFI+DMcI/khn+MNMBFFj5hllY9kRYscpcXEvWICMTv2e/q
8WrSc5k/pxhbjzviaVxE5c2ycKaDb8kH8n84G4Ua1O3Rv5qezZlT2YDQ6ITs6B93MLztCXQfTOto
4Xv+IkIM+rnAjzYkg/Wx/tmWsq12vBbpzhX0Lhtp9BYQoNDjdyGZlTEJsFfBURnPyO+STTduHhcG
e6hpV3jGeqhqn+q/a/sp4FRXzHEMqKZgwR7oOwufjYXY5539qYeyxQDmF90eyfnOkcK7a0t30I/W
/dWeLucYOpjF2uIHzbFROTUe3WkW0Zl93U07IBhDhGOirYJrkM+lirlcHFh6wppsdEDFo43/WTsE
/tsZOzkvNhdBTKohL9DE246v5RdmYuQgMXpzpF2/p3GcAGvpaw5i5MRG3xVH4lxi/A3QTCqhiH0M
uaiGneaZmyKA4F7hrdmGnuDYiZQaCvhGYpBnk0REf16fJroCf7GZilZRANFwszChbfpNIxstt5SE
rz5ydQm4ULmAdfLTztPfutiWmDzeoY8e3x9AA5vnCkvBrrlRSWAmHFjshPxckzrkJxyZKWan9KYZ
etaNS5hjAeG7shfDSc8U/tq2SUH4u+kf6CeJ9l9MwNIucP2uriiI35GOXrgCdvK0PefRN+e/JUw4
2PEBaxbTeC6M7/PzDBLnyU/zV+oEPdOCoTvgitt1axhj5Uda9+gx8qssNdtCAetVUtPdI/J67xO8
YGlXLeePETKWeEKgGzR6Qo1ChvnR77kg/OOD09bS15zf4uCKkgdLy+73iuzrdsRftOLZ9H7mJ44D
iMMhTGyxRT8ly/jhdcmBthproBUmedRuq9j0MhOs6tM9PxGmOUiGJbvyMgVyZ69XytRs2tjGvZW2
KuTdT5svOiEqErYfabqizSo4XjBa2hn4YWqIbjbZiXjRxSJyx1fWmBkK+FqW+uJBUArFm/Pixg1g
HlQmJ0EQG2QhQ4uyEzFXMpnNXe2k3qqQYzbBuzBoESgWZCqhfRI7T/5nxX2ZU4/jWxblpciaRJ0A
beaXfxUkAgAzwXblGTFijw23wDe6nmMuPDZqhxLEq54TrCKRYiLCJUnDC4u7KcYHDeIbiEWwGNK/
F2zuh1lUOkf8P2uza4FWDIbd7mqXlls04UdPr995xFOoXt1P/F8o6x01TCNBxEqeGfM2Y+/3gTTl
FteloVZ+xz0Tf2qZO4GCmRyKXuNZxFW7XCYVwyn/2gGSlYI9W0f/b0Byv+YK5VDdk7lHkFIxk1gl
+4/Ib5L4cZc43m8UfEXff/K4TmHeG4NlS9krjm22KzjY18GFUBuxXgrYzUYndHqkWSvd7PjPLfK/
2A64KZkALEOHF8BX6jYuKEJ/xg3UP/v1bsRd7XjOavkGMxp+fWdklT+Ycqp4E2zyTqgXk+xyr6co
3EUaZ12LpQSomOqpkauYUtNee3dzgUmy/R4+9KxAbh3qmjEpJtNjRnEveWBqhylGlhabkZ1DZH+t
C6bb1NmFNKwqaNCHOSHnhtVPINWyqaXQkxq6wf7X27RRcC/I3NtOtTayaKJ/PgKtyLsAQrk7Fmhc
zyac7MhqzrzQw0yCjT2MJP9szZHFdEIu8EaQS090vG9C9v6i/QXGOd2Xk6REdFc6gNxTojH2/xyx
bW6ayc9Sy4gEHjNYtVRNvYKM0/TA3BNUIX0WivoqGyic8nYzLE6wSI9jdEGyxe5zjWawKIJ3sq/J
MRggrreCzfBMIm8k5loNTGIDySGe1dS5tERp3fohVg6HzO4j/bcN9yDjcdNxheKbok+nSZTcdnPY
u9i7jRheG8nKPUPM89Bf6AdbpFq9Ojk5vjufq9JsFwpGW0AchbkUdcZuFlG8bD2jA6DCGlOY3QNg
yl3CBy61UgZmBEJYU2NghDTih8/38ME6HAm3xTzDYtAQlxx7+jOxjmXp4Z1joe1lwUhHCVpmWnE8
+yhbHQxBSPWDnlDOOEUx/xeNOVGCkbMNAPGWUguV8ElgTNbXvD3zN6vJ2xIha8104XBB6P6rj5rb
cQpcDG/0QuVZgKofSgUVwz3bYPo3pq6/T6tPKmQhNE8Cjl1y0UDrS/5Jzrc292fe4zYaNP0zu/7M
sbx2WYUieZkoAEuO8jb4F18svZlK1LJMP4zxJtApuM/HvQgXJdUpND5JDbbNdv8a6kcQlec7Arqv
3TDfoqDfbwVWeFirEzI6R+pOG1nNF7stCVd08CiXf+nYLJnJEJUUa1H9ydGy9YM9yWV8E0sdWp6B
zj59MxAu9TKXkvcD7S2O6vr6RNjTSgc/EAm0RdoRfnVsV2pAf6Wog5KuttCoLnrT8lxUUeyafdnp
t4CwplXXpreX48QipF9dq8alAu4EKEuSlkUpKXyGTxF4mTxt3IJBoCw8A7Ek1mAI2Mv2NAcRUfJy
1Ieem36pOUP9z5UScLLfzwduhbUGqqVtWlwVABwqEyvCbZiFju59do5/TCa89xnS1fmwHW2Jem6U
GMEEZTubhTu7erXEGWbwRNHcecrCowzUGXPvI2VgMzna/nNuRFmoW9XlLLwpLRbOJQ3+7RdDkE0U
Jn4cILdDsppditq57M3vVNzHNQUDmvyikfuX8lO3aMQVVpromK1EtQ03pvtw+Xv2N4t+DSfRfJF3
5U8eys49ynszXhnF5fUmUl9LEco5EHjDA/zpKKT0yc4HZBUcE9Rzq44v6z0QIEv/zz4L91AHPpW1
FlYaT5Ow7GiuHctAJEUdeV48QQtY9MPU2D4dCigp+6LtJW9U81FImkH83lmSQtxcfCVaqRz9C6A/
gm2LQwTkHWJGJmgqO11/mIxjylIn7vJtA0qxsmGjFoXET4c6UBeZQxsVGp/wUt9LIY45P1ErUfHz
xgR1fIj1Wou9SMhvGuZR/R/F23iZiV0SUm7fKAlGn6FJr76oLCTtNMonqG9ZwFYnU+Dp6CuZ8Llm
N0QLfphC6L4r4OdhFcESCxrVniIUJ05fH+6Tm0aDJaJcG5QX9yalP7idEMbbdKfduZmmchft8fMl
Hs5DqZxASV9FgL2hOo/of7aTHsQgzDxSr6i9CCG9lPHK4yq5rev2gThQqvpAbFB44wnkaqr4lja4
ZJrj7irmoFnBIyPrcgotqYrXZ4ncbzYy16Ujb6XpIg9vW2jnO1dsaMMaQpNz/ugnkd81oo0zk0Yi
S6OFZo0zzI4B11F1RC/XoYaurVqlIljC2r+nNhP9IBPoXaOKc/erpmJ8YBAg5gsN+gultaonFYzx
+8Gf79Dr3vU/9kTCwOiA4GmE40GcSNFPmVPCOHu8VYXQ+m4+XXd6ZrShqYePBERwgwoE/jp8TOts
T+U/WOQ0t3xPRni5CAmaG1bkwRnbYqhxaFI0i9BZnN18C9dW+HST01ZD3/8w6JID/AEiQ9in5Hwg
qQMe0EqLDcqidnTaBAWbCwy5z1Vw4SzlgZCX5qMrdqN0YeUmLT0nNVj0iwIilqGLr/VcEUAa05m2
l8LIJgWx3c+nLlSIUbwsckW49i0DbEhgEz7+SyQqjRKIDW6k626LfwLSRXxndfIKGQ0mYY3QmiMd
Pm7sflGMSormE4rq/SgbNprv0JN9VjgXJPL3zrmVKwcDE5vQuskspAicvWIBJlEzx8EKSjjSqNEJ
qsqZEqbJ7EnnMyKay/crl185ADNO29bfei2J4ffxAAnbW9rRyU2mZs2YOs3lAOy7ThorcG6DWUPd
DGSoFGAeiGAipjz/4dnF0caLZjAZ+FZSeQX06wxkfhDhaILgjLHZ1jOFh5eN6hWhP6EqHZBMJExY
fEGNwApXORHZ4TUizL5gZ9VYp3N9XbileK4XgqpZyLf3K0qwuaxXeH3jrtwf4qvAp8cDNi0Gy7xZ
Y0wgDqk9RCiQCdKwYTJjX9GF+b4eEuyC93mXhu2kRioPpbOCdEsbmAfcLZpaYqF2fnCQ+acJ9+Y1
yNgZoPr+01/iKDcxEypqPfHgN5uziSCq3NJB2hLWbraIJ841fTBapWN8PDrf2VIOCm6EN8NT8d/w
zPNGBds5DSXpPc05341zaAPu4GOeoZuOxJ8NyXTxiBswbH+Z5HdAAX2IMHFW5KNZYcgq2tUM/ewa
peJua78KlA0/93GCxx1vu+aCKDjLYRVytysfgJ7JnRGK/a0B5fFhQDEHbdK41QlIWhvsJmOJ7WZi
xWwgy4k/GskZdsguQnYYKQENDfVRmiyGzZ5W0KZlnaCY7GL8M45QWsb/AW+KhEZ8Tsku3tEdkO5G
863rQJHn0iLeMFVd4SMNm/XNb9tHZtksQpkbxrjgp06ned5M3gUzJ6TC3+pW0aspldshWD+lxQ50
Q+6pHRS0DLIz1gqff9/Zw3RnmmeMwvCvYxd5p/02sRBDxkMcu3DLiHDg7af1ctZ1YEqdi5X6toia
v+CRxfZwj9/OeoCaieKmKtWKEORxXteDZtb9YlaQ+/FOfxJw1VvbQZxBdoo6KjcJfADUHaEBAZQz
5OCiOrZIevPnbm1b/ndDc1v25grd25yfB40+ccuUa8SnwYv4XTv8G+gHsiOaG7spQRlu7ajgkbMj
LZKDyxPf4lTGN3OvAmTuJgJvE2aSvvi5qh/ibKGPcHuckSenUy0YbRM6BhSpUej28n2YuJzPut43
EbplO+m2FQq7xSRBVOvxuVKkJde1Zi9TbGT8QMz9LXKcqiioAfnkPECASGUvr3opGlBbsTYU+/BK
aeTAbJUpTfamHG3P4g7QCsOv6G3LviNNE5Ux5qklIeXtwu16rU2TeEXC8OXF13Ggrj9vULUCT6ww
tKMeVOieg2ohulA9afScWxNOvlmvQyw82CsjherXaRg3ZlJVAylCdA0RlbejqMDx5pKFV+V8Ysrf
YSnfdNWCppim7eZtew9IXmJI88QHhPKHtVtv2preIPJvN7sfazGi0INeG1ri7H6ovn8qPFcgzo+D
W4ghrOyEhgH5d/feTJqAX9Ko1hXv8xhQqoIXIgaFpX6C6dFxC3Qr7c/1Omn8QfsYleyX2jjBzKHy
XMoyOJkKvUR9dZpd4dHoIRxmdTjJQFgKi4NnpdjZShimNLFlqeCbNbdH2ldLRHM0arPrYL8OCw/t
1KmUUcDuq7XTYOFMT8ytnYAP6YUIUasbvs/+zSzpXWLS2JreR2LnZgQZawHnSmxKsAzTljxS3VIg
s56wJjs4foNaW/pS0YcGQJk+rsylE7qBElW7q9vY3BQl/Ojo7B4YK/7EidfQROIy/ltlFdkr+bOw
WwyuTlE33RaF9KDAO2QwnMOOQmfE2hrfJWuxeVDePYMLWusGNrdY4GyBw4ccdRi37uJ/Cn6Pj5kw
6YxuaS2AWfR33yJf4+jbA5itk06QX8Z2W+8Y+pZKpF2vOxM4QjhJ+FeFjrKacFy3JHOsPIyeivhM
DoYHX3wLGY4g1XDvI78aFqZULuOPQfciS40bPN6X8Q87V6pwjMSv5BP05Ow7E9ec6xEHOmBDz83R
uWKqHsCRo/5SVzk6cFfXwRkrSynQ9Ade0VRR6z7rTZ7DZ8x1e71ws84grbrh3bCobgGmSTvs4s10
KWjGJrKcHXfJlM9HYYqZ0WWVdrE4D5hYgisk7qFs0USc+5HVKvtB14iR6qnUEaK2DqFilaB16qRA
OvdGGsH0FkAyNiViazS97kZGg5MuAEpAkCRKhxZEcU+RJTjjvbcCSfwhehe6tt+8m9yHuHzCjGf2
YILkkkVjJJTYGHsGnf2MJr/hFJfyzUzcg/QzcghZgWMA3nRURKItLmhPsUpgwH5G3PcEe36wkBKo
2eWS3wd+HdVJCwxHgnsIq8vPPmHnFDt/rye6V/68Q8MSNaTOLgHz0aM9y4ogC8+hW9Yi8nqkkZWI
biA9Q8eL8XwMFHSWCifcDgC8WM1FnAFgLgsnewk/orwcIrb6s4h1gyaxGh5R83mRXpIkbpot2Acv
AuCIzf2IHVB6kSVWJJLLg1Y4jE5VZAQj355ZmbODwUEArfg02qBYYbhVwk1BUyKiQB4Pw03MUX5l
0TjyniQ5iiRkDq/pdVERRcuzVjUvYcwhRKTv4K4S+wvGxqGoZ5bExGPhsldbjKk0dS7fNsr2xtEp
ddN66E7HigiBJb0XgUP5IlW47IoWEb/oqazNL5w0ResgM3QBnHFMl2gpbj3AGTn1E7QS7oC48PIs
F73ZBgJq2ETEySRbbNpA0DenEFhuEVEI4wgpiWyDUponDmsOYM9uDeuztCH268nkSyAd7V2qBSlN
OTthVEMWg5GFJNJhCT3GppkwDcYuXbzuCEVPipVs/BuFp0Jl0tlaIl7U974P4j44sTzVIKuv5HuS
9a64Zv6FyPgoXaiekRNuXrysdYrGD6fF34QiAu+pZMbVxgYMoi6l8sSMi7P3fPY57su5rQbHqC9I
Kva0TMm695nP5lBPVV7/BvO8ZzBi5nmAZrSUmd9GT7weQGJpDncmG5L1lE2rUfoAQUyCwXq6iOqe
EC52jRhVatwtrnOvoawu9gx6gNtR02PdkNvNMdR7R8X/fkTx8GfbhZlnb264IbRWqpKKauYX3c8j
3HpwH9+FeZJXjnWl8tz6VQArV02FblfLNlsitMToEbpmHZW3XSmnKFjTmSg87thG2ozPCQmg914G
OMJzMhdoV+AixPty8j+mfJG+CeXStOM21JSEa0ONUO2n5N5GxEftgiSDEZi4zPlMc09L4zykEKUe
2h1NmcgWhZmFyGw5xvO3TTFT/gjmZLcn4EypJjFp2jq5so1BNL5HJ56MaCTiL2jlVSWyvzlXQSyf
NgHqZeDDJAx2yL9rZkpUAwJd9ZhIIeMt4/9En8PtLYXtw4rAHUOgQb1ruYApiBMGzXezOG0hzxIa
sVQfKJKJyCHRKbfi+ef6OYh/Scwl9+SRjf93EAEr3c6kRRiKV2AAmy4tkh5KAaE7p9pAGlxH48W9
gb+7rGVW/S+rULsZ3M1e8p9nKIc/V6rlbj3bLA350QidlFUzX1x4zo9RZTmQTTnkEXexn6Dtd1tZ
lldQ2af0NS01/z2ZfgzLRutBikXb45g6kCzKPnRFwBi2l7kaT8W8Ok4sbBDmcR44HBue+CYOzuRz
251VSJXyjK24Hvty4Eg/RDd1XCOQdnboRXSfvnInbo4AzSxRfkZT3Pfp8e0bZTk+pJ+Xf5hcbeEO
bWEzf3d+qElPZVOhokqZbMT0Rgr9tguo5yiOortwSFtLrZIDlb7AXwUKcUSbBWub0BFqKSfKKlsc
PMfLSQoXRH41Tfbh8YI9YbyYD6Dg688Al4cSJO5uKn0PTZlzSncorLYkdJDSQ3r8Ir8E6QyhslWk
uSyo++aYaDEgVe2o2+uhAVylX5Pf2kbnu5hSGoiQ+e7QrFZhY1mYtVU2trd99etNSM0AoxunM+5K
KdUdjmHK9gw2V14MpC8lCTrbRAg+Gz3zhqsm65N/lMYYAo+Cwnme79PxPBKjKw0AGUD7wDhCwsIa
fLw1VcnPqFqrPoSXSQ24/m2ZgqXmGaACsoDtigd4jk7X08mR8s7SZObLoiSztP2RWLATG28OrQbQ
xZqQc1Ohbj/hqRkL2cMYRjqHos1EikuoaX8fl4n7/I7v8j0K8YTI+XjREodMjHvUs1cRxfgq/Byk
gEkUqVGAWVGfHm7No4vhRVnjJeNY3b7aTZF33ZBO63PmzUhLbWpETqPX1RrxFtcAsVrDTHUF5x3T
yAmTFaJC2L6U4myfbZdUTh5/6hzR5JiAxML2V764+Pk9KdRAZCHX+vvr7V/Emr38/wRfa6lfr75f
JmEN9EXEIsvNqhOL+DX4MHoRHPpOv7Hh3fG+vyRuy3YhidnTITahyYF+l/QwrFMZnAUcbSDDOy1c
EUxzRoA/zjGz9jnwn3rIKl63mpqkggs/ERlIwHKjEiwJMYTC0bU12VJLkC6up2PwAE2XeKUpETXV
s+NC5UhEwCm//VOAve4wXDvmTIjg1SgZfu7kA5bsuLJjjyJiWzjGVyiAsG74u+aFSfK4JwSOoNOy
Vr9cvclkm4abBe68oMkKIQw0SycwMw5sG0KG2k1j2OwptsEjesSih+hOrPyRVIsq2iXUEs/CCygj
TJOVuNKyEex8KUEudDihS4IdnnLx9jSq9V+ivDtfPTD7RRBvLjYzZKlGMwNMKLfu00a7CV0dRrjC
0jTN8j3lEkkm96hsvWif/WnmUFxu9fVzuabdP2f1U7daHp3g1JD00KHfxluAqlpUhyMNsEmeNyBQ
mBmjIY4MvRLvqgpAfvzSnPNtq5MqvVMFysOdOWVe8WqBqBEnkFi3FQzTE2TTGD8bMoCMtLx9Mg1a
kUY6mVSXIEGqQrUimOsKBc1IoYAiCUzQtcRX/JdQRh/b4QbimuVMsmyubO9yYiIFPjbKqM1vGU4P
uvRRtTXph/7OOH8lJmw0WytdLpgOAXhwUtvX/okPXzz0p6dewIXvBKyMd2b2vZVm7ZN/LcKXP9MQ
QN5Dp7dFDOis215r0eNGWndXzAIqZZDi2UstC/Rg1yg0NmlbJKtoLeB8gP9KU5Ahpd6l1urLdNr1
NiolXV7d+dg1rq/GUxHxhU+7VaC/xVWe7QNI9ZNGOfLGd5DDF2/+Vu0p8VDPbN0J4+GKWARq5Ccx
FB/B/9oXB07POzQv2vXQ6JvO+UkkgQzmMlLsNeMvuJyUvhSHYPA52IJwbCMGYxGbytVlge6kvQ8U
M7SsYa1O89nEbBjIzL/QdNu+91YGhja9MZljdhKlIa7ArQpfz5CZRnkvPGvXNAAsVN2q1ZRYEK/6
Y/QjKMciKQAXAVP7QaF1+1Dzjmc0LPmGDYawHO1b6UdzAOE053LLtf7q0UWU0T6IhE1isaxy/5RX
JplkE+LIjzuDUBQ/SlNFnh2RPIaS0oYgCI95B7ooI9zH4x6L/nQG0pKkcFbczrW2xeLIq/zAOSab
m323db2EjOw8fA5aABu5d1VXYlr293NsQvpnTraowqQIz9kXydKnqAdqI0XjzJSzFiRMi1iqVzr2
AosBP5eaIeOFDh3vpIl+Jb+vX6RENbBUULkmCL+fZpsb8chF8fd/fW5SvBWZxdQ/hlJSp42NjEdN
xFvDjkszt3JX8E4SPCtOxyt8UxyRnHBe1p11n+YkyO7Zi2dYarwXr747Q/9orFiyxhZIwWI+Dc6/
mlQ7Ix+ESsv7uXWb8Wmc80ewilGDDv+TCb+hh44eLFDPTEOoabaIJ4nOi53HfPulu4T4AyOdhAAx
KjNmFxCQSbq9aQjfx2JgKn8/Mqj5MZmYuTzqhyUXWK5lD1t7XU+2a7EkarqB3jaGH+NvaIp0i82k
ywe3zJ2axXhFKU6xZtYDGhTW1uO2K0kLPg22qIf8v1T3EIpEkc1go+xipaS3B8CPR2/jmzGcOlVM
gpeuVcBYHYrLlZpnTbrZm6VCNmuVm/ZsfaPJqsV34o1hFM1QoDSx5dI1v/WOQnfya5DEsvPw/N7t
+LkW6AVD+DYPeroFYV4N3ZuiqLzdZrtxWhZpfbUL+XVoxCzbThIL8ASMqsXkdyMx1+EX3JZ54hVb
SmauXBAGbULUOlVnUafPRi6fwuRyc4VRRCZN854eSD08ib9havw/YH7PDY1w8t+StgqjIniKULIU
V8MDrZz4fXeqa/o4rIpHcK8YG7GBIZCsQS0x3JL91ZiB5NrzNecESQ3mb9GhmpNP0wRB60ljd4An
EP46tCGQI9u2XnnNFvgDph5lCYqBpIkcbM5MDgr62WVL6IPeV+cieJLo9/wXLHcSJWkhxorgu/z1
PYNwR+zyzn+O0LQPImq8rcV4DpH+j653KPDlrjvfA7qFTpG3SCZnZg+7EfqlOu2AmfJz7MIuSzsA
LJbaafABil3lBNA7e4h3eaOiTXbnun6qsZ3dugNADle2F1x9rhWXXB8ZiizkIWxftNZusYE+ofx1
KScea/VumP2w9BT6yOcauq8HUn175diWpX8X+A+zDyEnwAoeWFbEExAN0z+ci/uALEfdx/xqMah6
45cN8kG6f40HdAn03QjEtx5HqrsXzXWjWlt3pIqJVMgUZJTSZcc2mfEoN+f4H4yo/pNTffIrth0X
zVv90KUm1pNLrMzGzCMbiwS6JpfKZ97LgTl7fcU/ITohKZqfpLDM0KkQD1GbEQWRjNSIq3O3lD/S
K34eiGvZtHsmAXgXjqq8L4HKFmsvH8L3Tc4cd+uvEYA+atGDv1O3uqhvxmhO+zMoAw2uvmiQih+r
c+pkMDfwZRzd9gcXVleiGzzbcSHZq1TAN0jOS80iSMAWhSpraByrwDeTlN68lKWQ0+VHMF25B0C0
KnlhaD5MehfyXfPk3ycsk6YhrIdJN6LE7EVIPG8geoK3/tuc14UGJ7aFxRnk2kvJuYKE9wrjrcYQ
gKDgwWr8PMIrWPME8CPVpsfukvUcB6wi2FmEp6uRjccKvlylObGRB71Z9xaQsw7W4uotu6KVutJb
am0rNY5XCc8CrS8QPDbSLf3vWyxbDCif/3iTI+31IG0MJnxDKrHaQR3Sksi2yMTZgmt8Wm/+n4XS
9FO6eRopUC0/ZveGALmyDqw5hTnc1rQzpmu0WbmIFE3B9ZrSH+QG7vRZELkqfCER11Ak0mUl6YZV
P8Twzq9twW5Z+qJ2yeAx8hmwk2QxiZ6ZWN+yJcfcbI0M+qCtuz+Tswhu7zeYUcMenvmbrn3edB34
IrhmO7wNdVUoQN4dGHynrltO9A/Opz9dtTPCorhWqdrHTsvPnRsfbgIrA7IWA+3xi34jZJ46JL2v
umuFMMJOAntPUJWpHbsiK3SctCY1uMsPW8dG+JIpQo5dwe0N96VwIXJYNet422l0bdaOaSxF/Oy5
NXlGMS65NicHd2B5pwkI+MpvzvX7tqyQLB+ZJDzxMFgpxmaKZCLa4TCbvsAbtEhuc0JUQoasNWo2
MjGpQgxnU7DQDWgEBC8ATFnBVxqwmqDvGABACatJYf33CBwsQKoxOEgr/HJhkW6pGUXjPtXSGO9d
LvHkParF5559RXB4AZFitNHPizPhZgCwwkgsTzQ6r2+FL9iYbyvGHq8uXcpeK12Y4LJcM9EZijXM
5eS/GWhX5CHjejjQlKN6C1tyN3TdyLyeFAqx2xdGeQ7OqsO/XkbT+Oik9TCXwRn6YlBWY2wENofa
gPwOsGbJFNj6yZ4I9NE2NKdm8N0FKAZ/b6L5nbM/ZtoqLNMrxe17/pM0iWjm11cdQhnuqRwIuT/F
0hB4w9F28X3FuRRdkU/tETkLUEg/+5hDfff3O5rn6rxEP3E8EfF3OG/EYm+Nmmzf8BM95XdcIwBt
NSlni5oh+Zj7YkavXNW/xhaOPvnSF1+DYzTntMPWttvo1ayQxnsj/4+dow9HrHfXoaFY4QyCSMkJ
MpBKbp3BRJYnPfepcwOXPYptY6ixRZzv/UYxaaSuQU4htx9DgxfLbl8AEDqzaEPOnIXXOcWPHfqw
hp5WkfccdbAqkWR0pydl6Xqq6gH7z5y15OosxmoR1pW3m8Sg+swNzCi19oXsahuyEynivJoPtyHt
3tUCVlh2fZWZmI7MJomjTgVFbzrnkSiLpvTYzr2ZZD4folDZ8c1aATd/ZTtkgRTBjc9CHt4ZyJNp
3Z9z86kNG9oRApVjV2m6Yx5GehphagGstBOIy3+w8dzNDDW9ypnYGEWS5sZUS6Ds/Y0orTsTBSDF
1dKbgy+D75RnUjEJ6ssQEel+aYT8Or0h1jU8ux34pszs9pK2jmXpVzXg7qK2iNwc6A3CSpgU3iqt
dqvfeLouySRAax7eDOtoOJp2SAhSiZzQkrdkurpreNI4o1mTQbmwhE7lF8o5AeSx92Z58qpEwk8D
R7h25Zrjye/N3PtU2ys66Ry4WAxxJLWc+MeAb3VfUlUnzTFeC7JHbTtMiUgePiCWvRBAmGRIZ+Ua
H5eAGR63vNxuMcyNHE6ZjNK/FJ/2evyQkZGjPPfNpWuo7i1pW2pe2xEi7c7p/klnWxd2sCHTkTsJ
tt/6SlQ7Q6nNmFsTEHa6fnBA7E5Bq+aUqSpETb/TwPlx4wvrynvvjuQAq3xAgMyGAspMPetmBa9b
wSWIs3WwpyUhD7hSUAwQEBBE6m+AN2up6U+1Z7LarM/SwsSyhYyfonZX55QbwbhRG5SRJatK9DVr
VGpTa/HUV+Vn51g5mv4CgtbRPA6weeaBMI2pbt3GE0RNFu/Yowy3qN1+nufPErCfsr03PulXQyRb
AMqhkgS3Or9IykIcPPxchCrz8xWwSU9in5QUDvprr/IFm144g/vELi0TSDl2eX3zwYwaqmQcAMhx
hF9+pBYzr/SbZAhJkyDU1D8ywgSx3rxDWFgIpBClVGcl15BNzWdUlsswtVc1fDPpVfS3bdRG6+Or
G1eiNJ12u1QQsQZRc8hrNcweKv/54LMnM0fLbU2vtkVbjxSu/d+ZqqRBxugZKHfNZfE4wS567UO4
QrxKxkqggrmaOgjIOOHeY+VIYXa7XLcVHZB9uDF74al9UHweXE+MwwxvRB4sSp9QHGufTuUIFcis
TrNwxZ1eFoT5g/Pqed/RLzV8VN3z9YMAJC37j3XhT4hEn/a8hoiPiS2Wx5ZyPxZAf1haZSLUFPfT
G2PktfysBAujhweD+gMv0OCLlROmzDxepn7Y3j6gNIKvK89DFW4gjHGG3M1gTARjwV26nyXsK+9e
k6euxgctyXkoWZkMANOI0ChhVXaMKD5uNh1+W9AcSKSNitkrS/3iIY2jWWW5qncZIcZRw8VUxLLt
lfgb3dY++vX3nkCF7PjBSay3CZdSmIOyoMJByx/rvMTR/9mbPDgZNcHmgndzjU58Hgi2ZBnHcIxA
KArusfoLmByrU5Px6RuB6JFkVGMwGXZdbZkGjiATXce0UhvRTR3YYOeNs7AhFGoWswBEPxce3YX3
HWI7av28T3DfZ2Xlnu+gCwDEaHicu2CtQYfjTRAHSyuE6+jzM2VdPDA2DsFa6WxCSpHYseFpy2q0
Td+5D0fHiCAGgg7BUElTOatyw9jX8xNbEo7SGZZqcX8FdfO0UuqfC2osTBukwFavSurTpvAQTzA2
SocJouOlebwqVlKN1i5eGoD+Vt8l+Lc3crQ0K27m1fUy89hWNr8VNyTs08EuSrOzCWDKrmBQILlY
ajjMgcjKWvwzplC8IwtoLgJtX0eMTC8ZWY5igSA3KwGVWDsB/b3nzCuRJc/4g0ONAMXr5fIGn9to
EJWNvN7snDzj3bP69bGazrgCiJ2YhKF+8Z6x/IpqVBArEVYffyBQWJzWEqh8SHWsNR1K+jOX5TMq
mejeBeEr9eCW5WIQWDVSOgCNk7QhZXBZoXJ64qotHbizRAiWHspiVL1bCRtrK2Ru8ijezbNqJ6Ax
+AWl2y37eaBwxnLD727H4txz5D94Yi6dnczDtvcZP0Lq5/2puykQ3cGLq+7BPc/Y83TaMunJhtNs
w7pggH9NCFjc3Ir7f0h4wlOlTLw4bTrBIvp2AbGErNEUrWon1U+Z9SFSZVm1k450zSIHoB51JWuk
2ZCBCzLy413ccJFzGLG5emBJXvtEJUZlFIYeeeBuZiVpSshOHQWp4XBrRl7OtM3yS575eItd9tTT
gQEhVtGahcdLjVON1sRRDnhnX//dOdMEQ/VisLLrEpqZjeTxLwt/qLcQKXNsTvdxpIvwfT+w7kNR
ThxXgoXbBxUKRfzfhaGXZWY0oLgjxAtr+1r2+jk/GJXmHexQF3j+NPr2qzlrFt9g+L+4D6ISr2UJ
O5jkNK0i/dFlJYQblVgY+1iZPozULAMoMp4p10S5N1egZBfp6JETOBzXCGwrcC/EpbpKAmzICWxc
mZh1A0u+39drITfq63gE0iFBZ3x+sCFJbHcvIfl18b0CFI0fg9ljh1YUXZN7VjwO/plB1Oi3LYR+
zkOKQMVeWpymlvn5EzvDAb3vQ3K+/qv139MWc7IZzYSE2S18vOrhErLJxMyr6VQm7AzfL0P7odq9
G9GvbSqzi0L/3zTq2ZlEKrOOIRLGU0j39FE/hBtrOXcCWEd8gaX1OtsKXBYkUtrnjxjBoq8l3jKD
cEMdNaleluDykPON6KDjTZ2N587IpnxvFu2dIE8MuJxS2E63msZ41fuqd+RF7GqzFmiU+FGfkc7Q
Y9d2Kw84Vfqif9qPn/ZdE9HJxTHY5Im14uq6lqhWKfp1rjByi1ghYbk7x2MABlXEm9uD2KJBuVQC
LyaMLYLNsul5ChlWv+9r6XWCgJr+ret97hIBt18kh/iDN2H6+RM6zq4EHihx9rmeCC7JcZ89/7cT
FgGzfIcpykmx8My1w0XJNsRI6AuGVpS6mm7X5BZbKyz7G2kfUWb0fn7smsLzdcifXLAowTxYzhMW
8M5XHoRWyN2Bbqw5i7uKbeILmaN2DId6JFr5zsSp/li2YtWCLkSfjCaZBGP35byKo2V1oqMg9zYm
LKYOT4lK+eZwpaNnQRJV+TI274cuRluvmpVyFCn2rW1UU87ba9gYJOrG4t/+c86Kuco1jLQ3Aj+p
C5goJm8m9oasdInJJ6iBTiqQtCXo6UuPP4AI1EMpomlhbbqXubWBChjhXToH9JEbM0RcBbKh0mj0
/xTmk4rrIyKFqAOHrNKIlxEhTMvOse5p5QX5OMtGAlhoqZafGdUwc5MJxrJxrUp/7bqRBIpWdkOa
iTYtbdoVjIyMXfhmzrbhZFn4FEqv9yZO6rIc9R7uXSnvHaoFyFfx9uFz97rs4x32GoIqa9joI+37
uERKUTmfszpO4obHUPzlsbKUSwpdpfWttf3wbtDIvJfuXtnWwQEFzr3EyUUOXMvbZ5hSfN/CZGI4
Yc5QzvOsPTxu9W0858S8qfwf/9KdjKdRCcMIu2EFPw84RJX4O2HNlfx/YQzF+rXdhdsbQvtKfPKX
j/W4qHJPFvPO8GMT+0qVfzZQ0EWH+nKIlcLR5x6F8vETVsOoVMNNKckRjgSFWTMn3W2OO9gJ0wC1
W3SubV7Iystq0rbZxgomUJ6othMtpg1eEseAI8gOXVT7+4A3zPUflA2LR2DRUIdgmdSUClufDtYg
Cv2k2VNe//rxaCBdsBKgwOAVl0g24EjKmkisnWkc3JOTxnsbkFsMIYO8c7+9NH8O3KBMxOaLSSZH
N1nxl54myWA9JUg82fknt0ZpXF27lcYO3E044JWEEAZcA3FvjZ+hao8Pz61L+PRwjgh5UtJwLK7C
JZM21fwwWf09dTQJbJwMbFS6bM42C9uYKBaXbUPi6wzdfYb21G8Bo5wG5OH/tF5mjHxFBgZcR0ps
KLcAZiHyPTgLlpZET0qUaxR7pQ335uqDzVRZIj9AAPBeUFkB1TvwkhZ5x7xZNULFrs6NqaQUXQFt
G0JrDm8zHtEZR4FRbUWOBudhE5pI9lL01DNf77GZZDJhmrKW+NAxtOBC0LXDAe+eOS/7a7Mk6XXj
pP1oITHVdNt/cinU/VDT1WJLoPQNYyGTBwGg7BAvJl2pg5v3MUdxQqavwLwa8abH28HtYIBdRbv8
BmhkRa0NaVS7ILGR4dnjkDPny3VcJ/yXuvcnq6SIr1McNC3F9Y+iqWHbsCYHZ9Db1oBdEIdyT+kN
TyRhPHDj7ukmMC+FHQgZkLeK3ra8/4xkmiwepLY5/SW2nX+hnKVyoTTYY1XxbZlRDS3/XV4Sml7U
rV0N13b70X5YvUdZdKcNKNJO7GxCvYLQDRxWE35dLtLII9sSGi+Ow41moO3yQu2iHzuR+cipHSCO
NCbP+dhjYiGb9S2aL5PM7KrUiv17Y/Qi1S7CtTIRzr7kMaLWkakMDfOQRR//yJBYx3jjKUXMB6A5
Gt7YYnj1QAKaV/+HpruLjX3YbOOn629+sVTMrvI6anwgD6O3vA59HGzdNgClSDi4y27kbt56cCXM
X4gyVGw7qhdU12mb3kNzd5lW8j4BMGk3Pxy8OpzZDmxR8ZQxlRenZzDRNNwcP5JNTKpB7HeGkXVb
/SbT6PWI2XNMzdcLF/iMCOD/zQ5PoUJ1OVU/+SMkqJteRsCE4Z8ppf7J1EXQRowbr/MSjIPDmQXX
BOLSeFf6M+mF+uoacYtvVF48uPEIjne6ZuCIE2p77dlogqUQ6iMSY3cq2Pi7AJn9juVzuLnVOebL
OZyFMygsUwLBY8rHRAdQg1DtAeuxfv3XTHxLBz3LnxnUh0mNe9ulTFlLNehJev/dJPTphCPLn3DS
EO8+tb+hB6nIM0a9DN/OmFtvZvXavHgqY2fm7YnJ+mZl4upXph+ojlXhNtl8TsoAh+GMe/RoYyI2
JbrKLbJSFqQXkyBc321lYJC6F++mqVVNUe9W8p0T0ncWwlBdK8cRn1wRznqdVWt7MfcqAzEykpxA
tURv4lYlC01zt6IDYBN+DcnSE/U839Yh+qTfO6+ZcWaSjA31HfqNKeu+CF70cHaVevgemgNC1Lai
hgkEJpgDie36GwrVDq+1WIZGzatfVix8XwZdLCdfXl0CDRcpCRKvzhkfkFv4HK2uu9GOHSiDeP07
a6VA9+E4Ys+ntRxBNax3FQ8lylAXd961Hiw++8QbBYtJCkqNxxXDzVZAOWxgpSa8gIe/2xVM38vc
JgmITe6wvtuYWNTKjlB9+ll/eC9iM9iZ6Bl9370B/XSzvOywsGsEEzWi+OGzUFAcBUypGIZ+6FD0
wFvezDGgznfS4fmJz2Lkyv/XQ8Yxey1imKeBk45Xd36pob5e2QdLs3CnDx84gPWnDS/wC0MVqdOq
5d694md/RBoVRRa92m2ZdzrYaoEejnxpvl30TD/3eZaZ4KUhqmlQrcs5TnS7HeGQM3AuOYH2o2XB
8dpwwCrHsy0x8Camh2mM1ARqkFMxb6V9CqDs7QnYQeISU+NJ4OdgUTCj6UABVLJae9WClsx6Q3KW
7KY87jWM4yw+8Y4MSFd+6aRNpqR1bnkNXwhzUSlcFFJ4sO88KUgSvcLrHuYto0MSpVURT5aBAUGS
s3BL3jxvbhtk0ghdC/o1vJqwWEi9bQLuBGwLHMKdu0YC+hk3vNvHH39yHXqGZzmLtKoZ5dNXEIMq
xJjjoH7fCK1VK/4O2VSSeQm3gSjQXN5cCsJK7h+0jtQ9gnlW+krq5bGeMxzRBVkRA1tq6e8c5yZQ
9RrQjiXjkB5IDA69RsPsfuHu/PYDJebajBOUbSp9c8VAl7Q2rTtJTIcsYIwN9oF9SqBn8zJGgzHd
cee6dik2alnx0MY0XRxz//xvC67fDgPciLQ5tospwiDi6+uTc/hQyBRDN9XDtggOsawQthSDflfp
7GOJBtzBNDnK5hI7lURh8LgLU8xHcM4Qa2PrZRLeRptba+3LF6z59dSiMZvvwhSMr8DSujFmrNjG
P1USycJ6C3lnwDJX9qJddZGdhyfvmu0tPu4E5n/Q1z9pAmkWlL9yDDdk1C/QOvUeA5t2bBHQzjF/
JsdM7W6/bYH0I3n8gp+CsE/uSDmsdMCm1zaUkrM71P8MJtmQfDDQjrKE7g3OygCoLwHu8yyW9KOQ
FtMPp48WDlKDqf22urjcC4BVSutED0MBOKfGSjoDm5/UPTBd2mREWuokXdhMWFqPF7bqzNdoYELf
350+zwsOTjkf6F0ERCaEoOJU9fEVqSh2raZX9jxicGVv8Ak/JqfuaSkkLDC5oob1uBgI7tdlPBR9
ENj/VmK2tHq73vDdY0e0Fg0gs1kFD5aDkv5/3aisIs43BfzH3gULij021+8hw1ru5x4Tn61UUoMX
QDelLQKttnkpvhMEqAMMOmAx4s5udSkVD1GqVPsioKKvvwFzNwbg4QwRKCCxAob8TqRVogwmJnef
Dj+i5ejHZT2RRkUxCfbg3loA/lBgoKhT4xZJVOD4hRM9VBAXni9M+yLvDZ9TD/eEyH7yWhuKg8fG
crry76XEmxpWHZVFmGyWrAyT1GUd6IKi2zqvtJl+EX2cPUqEaYQClqpuM4o/Y/IrMyiZKpLvts/z
bCc+lO89yNUCRxt2PrxgMBOWA8jVUk6IptkVHyFiwfjmZtCYLJbiemazGKRMVRhXrwi3bGwa/yDN
EtYY/Qufoz1ThjMCg0oUecsp+X0ssa1IcpmPmcSxav5kyEd/mx3L1cdssLFJDN0SVXHDuABGjKyg
Cecx5G04Ilk0tGNH/MINtm8juFufg7ABh0KfFTpd7MCBSK32JjqlMRG4D+MwWqIAbjd0CUi+LVFS
9QaaerIWFSyRTd0APqnEkaJbPspYXaw6bcm8fRPleoeuSJ68tw7H5e0zMCH8sbYIPA5uF7U7QTz/
WIkjfgQUs5DAawQNgIsd8/kjnbrYPWWzmMEf5UoIpc5TkGv5h0HfVyXpDPmM0cqb68yxtMEyWvVy
SBKPF/vIkwUH2tUaRevvHfmKDVWek4a1x3mt2JxJ+5vP/z2V+YbVpoNAQNB6npdJsake3ucWSFE0
zBhtuKTAh2sTTtgxaXS1Vwyy0T1vRmUYxpV28FyY3RFdLXxMTb2KSOf08WfNneVLJX3HMruBbM3u
OpHkfXOMxNKzkJ4BS6i4E1qWfa25pYQgSsrTQLtGoz+B1HrDR7RoXZnADEC2FhxxW2WCWKctHDxs
Pwqb/YJ32tqpBetzCV3eg/IB+HLPRLqbvtY9ZZOi3R0qUqtAPq2vP5HuIOYohcYQRaEshqykFQ8I
iAmykIXB8JbJkELvrEELJxUKsH4o2ODB16mWk/vxwP+0EVLCLcKkSTFlvcbU9fGtHquvQcLRkBJd
6Z5rPPLqOBvCzPAoM/z+X5S4goHvMXvSvp+6y7nLnLK7pmM6xj3FLUVik45wuOi1xFbO2KbAJ5k9
m98zF8HspodovR11qJCyhsT8lbn0SZmI01SBNgiqyDCUEnZdXnFhiujb1NO7daEv7FK62I67gNZo
4aGcIRW/6SIvVSFyUjo0NM5Q4GSIM6fMHs4CZsUIo7MW7m8AwzC1WduXi1oBxjJ+mhoG6OdnQajP
L9D3mUdrjiihdtg3s0fh8FqW+vRif3FXMQxQ5ogwd2TaknCNQ5Co0Bc5qWevTCDHs8lMPBL/Htyr
pQcu/0xzFFDJs4pgSvpIuzib4XtA726gKn62Te9dBYVzrSekceg1MFKqeZKuALlwmDXyqysmC29E
0WWDX8qM0mHK2gBRmEV2OJgPbUeeCFZPX1gnVK59AJXX7s5AVSVEqUW+XXBvK1K1SqazU9JLNaLy
/H4YIkxX46rA/SRPk7uWoKP838DmbhlNZrKVFJkyiU7IvXwbfChNVr/RHyw87Vymcuaa4ijmMQQu
8dICgNUMBpLYbMRMcJKx2qMclLtmdEOQAOb3tvFiOPA7/53bXaoqep1cp+ZdbiBUfM69jYvgBIH6
6Wh75YsbLaxD4ShlMRho8TT/PXVbuSGgXLwuzK8huIZyhDRiyWh8vjXKX8HHvOSwGK7hk0cCLWKB
pULtwyssLK8VBpR6l7NexJz9cIQ9bC5Pw+UeXRoz4mqBNniSwXBD3k9tfYqRY31yQDTzGZmKypf/
frzezdtHxRV7fZWOmqC622lzfitXSu4uwtH/pAL1dId3v2D/LrUTWpWX40z1HBwRSYvW4OfepK7e
rpExWBHO2nXZYgi7snodUNIOJib+V0pjr5GP4uOzFY/1k03Cy7EiA2ZFAUsTjQLyetfmcO5Q+Hyr
wbjtV/7n4PbIHU8yAo2hG+eakJfRxAjPcdcsdlCTpXAzceda+k0AVTqHaSH83Bxjod/Vpu72/Dig
x0dnv/tjtOa9nqBoyAon0VYkwDrGZ/a3qM1Pe3O3CDvJ7eASLwAy81og7J8q+coYp/162qD5EuT+
GCSs9OSqcWShvSIzl2SEqoWPp81wH05dkQ6gQrHSqGzJhbLyBFY8tooY04ATntu0D4PJXl6ZN+3+
QZpa8NmPapM2jYX4HcDy9fhqtdZpm3wGHaZdRUeodzc25DijKP0geQ243lK8k/bmNlEUj1a8Qvmr
/d9ePASwJmJ+lTdEtxIpNPQwZfnBf2L6R1LxK9HSHxlrEQ6P2e1Mh7+L7+VK3euUOq/Rj2LqmiUv
FzuVfToqn46+s33JpdThvQ4Tl7/nsGXfF1MePuQCklIvoxRlE9JNwNsAfVAY4gDWs8GzeRdJ+Q+m
mGtW/QJk7dz7SApe2IoKeH4nZnwFLimMgzm92CyO+vuhQwcaJNroTNrzZcCPOEMjfk+6mrOiKii2
4fjsO4Lohfa5HrInFimH7KL1TJ5qRqf/brgp56plyJK5mV8gFrsx06zdk/1xlIUDUtgungRKunLN
ZzfpUFWxIGjYatT3NF7eacJuWdY5oQD65nCGOvQAxvcNiLbLxDsoVzMLCkeAw4w19YZqIy2Xabku
aMEEcRsIfximelPAYGzGEHBwlOumgQBn2oZ4mWk1WrWBafy+0YgE6PYN2Z+ApMLYrppdfutc0E2h
aJ10mbDPKVwBVThjVXGHtNglzTzFeeU/YZ1i3tglzVaPe3jW5Ff0W5GWZxdAS2z8fwryqeNIEhDK
4mXKH71Eo6h4dsrpktTdYqjNHbeX47iGhXKBkgFYL1JlbFq7CCCaYMhWkQnak6vOhmdBuA3qFzUJ
h3cVJUAYgKwgdlly409wYmaA0MEuicJFYBWAaLNqos/Z/RHuo4rZuQuhZlOvqNd+sDhgDjar+N0X
gxP9RQHi4xaxvP5syIVMLfkwPHtza4FcPl7Vs/KLMjxlDIepRyByOy2BF+yrT+rkWD+rcYHSB91r
Ae5dAvDDAQKkIV2UDX+OUWWOD7REWTSo2D487As6kArSuhWEezjPWoPwmmqezbr/V56EnxmsC37c
rZxVbmp/5IJqpe6vK0NAhFriXJN8YSHDNEYZbcJAXv+tsJ/mr57lTT4B6rmVjyLgZYyk3Sg1Bqvt
s1u3QeZG7M7REch4/A88n3T8cxnGkhjxInc5wBCLrst3E6KqPiJFhjpGivfGD7HGx6SL726Mq/if
Top662wTDrRbHly0knCIDUXoEv+67vPGbxyDzDGpk92flaSfeEngQJ0WHuQAp+n0Y/k3OSMESOWH
Ha+E8bGRpHalqqK8Go5agAjTp7ZDppS5wrZwozycJEA02TuTLovzv7Q3v6FPhTwwDlVJB0NHHahH
u2VOP/E3SbdJ21GF/CEC04QULDkHqh9HClXnSa4rvej3sTnlj7/zg8VqHW23GiLJw0E16WV0td/d
5MFzgTPB/T5UmCxGXf+PYwIHRvNUZI0iQS3qRbFKrFAV3W1m78yMoIduqAqATZzY6Qqch7DVX42k
4z3I1u6J2FwPeC53GFuONgPzh+zqvD9KLWgmhGcD6hafFT3pCmZeclnie1qpNIncf043m0NJmc/i
7IR4Pmy8PU3IA54iPQvzc7YhrVmUZ3A71Z+EGk5G+OCSO1IWB4+fyJOR8NFkh5D44Y6Bd3XqXxkQ
EqoerCvPwkfDe/TVxG5iJjP73eI52eVTJvy1WIGt45lOP/tZ4L/dCp6Iv5Xr8eGayR3VDW0dkKuD
14F8Qpy326tBgvile6bkeFT4LW4+FV+GVyszrPzGvPJUnW678SsS49ow7Z+b08jH55TwuFXy5Mpp
7DnGxmzY7k8W0SkmPI/5FXjDmdOWB1/UC/6UCSJfmGNyjwdQGScC3zwEYIIHhPxq+f+9fFVTEJVH
Gq2zAchiPg92E06mkbS+oSXGuBMOAqjOryWqDmP2ImVeIzueQ781U6hCbp1mQVMyda/f5jKvCPjj
ru0YtvGVB6ZgiIsKglwrpz+oRLngNUnlgFnVoHdlZRiYsqCLA2cbRvVXL8/cMEkeAviHjtzVZ9IH
5wRL3x0E7qLBYprLwPYlhsO575wPfJv5hfouSfV3UYyn+UYC37jSJNlikDySRmGHK+To3b0OJY/F
urPyyz/lsBAglNKuE00ytWIiP6h7xDeDW6QgrYOYbNCiwknKDUDuBT/G33hcd052Bs2M4jk4nd1O
Fx6hvEJP6iBcOGl40jGkbuK72v7LdSX2ctMb1ywBaebLDKCYGNfPlbOZE7m+fru30t6WExJ4/bq8
KB7rvUJxen3ngJIFq+CehYbg5gtnQXBGlbrjUlfufYaTU9CbH+G1LEDM8gBFTFk5OhA1gFFIDjk4
c+dD4E3npDEse+94xr5R3z862odf9zlU/EvhAoolL28C9j6/er0J/fNXDQwvEJLTLtL871kFa7X5
sOdmqdLqoa7gzXgpMEMITo43kTobaRXtSLm7mLkjaA/7k9Pjzmd8t9HWP/j3phxNFmeGOPFcpVb9
oI9f4T6ZPYww6KwPmTUb0GTLpK2YbiyKTcZtL63J3JBziAPL+l3vUo5bqWXItTY6p2+qG/HZeppu
KM1/EzEgCDPbdIiadsr27uEjZUA1DnQhrYl41XOeWEGnFfdni/FPLVCDUiToVxKQelMBXWRWHY4I
F9US65czWcRhc+VaPhVYjRQEWnoNcRbHwvH2/JW9lREYZgg56HzMDyTg9heIFdxRbLm/GHSbVNTU
eAci/HcmrWc+h7xRe5leq3ohy4eIOYxjECjVFxfcyFdSFPG9WRq3Ij1+/95l2ZAM4q4WvyL9Vyxa
/+STwS7r0SSVCAnWN5eBShVZjCnB16zgt5gGcE0h9cPgVUIhyaSdNITwcN2zAqtE/NdWBvOMsb/Y
o4xebY2OZFBzbCUUhpQObmImKFlKL3Iax2E4wOpR8p7VoQnG/YbZ3RTY2K57q75Ns180Q2wHFQTA
7e8Ct6MFOLHkWiLXxG4522+dkQAXNcrlsvfaStoECaArXs2pHkFQ9/79o0fzFn//YayE+r9svorK
5DfblqLVhECHg3VLsnvnNa2uZGV/q6cCxdlMTkoaQ7LVOLCy6KX0dePZ9kC5/eq9jH9Gc5GZHqGG
AUHDLaLy4NipAmyiPb4lyGvu+WS/vTGV2uMXV2uXxjl9Cm9+Dk5c4IUZMU1wiLbeVyKkbr/yXVjs
vxJUIJcAnmrG3pQfGCymMTI9QzwWLYW4kcMhoGxdW6S9ZkKYZsOGcF6ETKK5YputpJ4FI6YcefRJ
OT4/+5tzUcKiV93Xlwfh+aWZHGYCM/HcynkbvPDt/kQvy3jcwRfzdRu3yekILwtc+QR9NiGP2pmt
2M3umC7vwnuSwO8OVRlBlcm5c744twqGY9z3bDmcjBS9EOVsgDNkkLivCk3xjy1t9mmH/T7JQyea
PjqVCSxw/zO1fYauYuRyp8KSpDBffWcozZOgos8UsVQSRNZV/h1FwUI1Zm/y+IxpSUAN1+z+WFYH
+3Ji6K0pnQELMRmSte5M9a+eqNJU8wYHvqQWz+lroK9EzzcUlviQhd0bbVUUVtcim1b14r6y4/KW
o8ttU6OtW61ijYHKi1ePbtetpu9OAtPPZkGDXfZ2WicspZUbMac0dAspb/V5jytjkPvPgwoDCTVj
pzUDnbpnxdJorwrYhyKCQFObYSDgPbIQ9a1pIWjn+3L5fTVfCfXksF6F/059QdYlyO175N9MuT6G
AvM646ZVps5NIANtrMQeUEw78zU0+A5SFT9odzSJxmbof6+KvIH57m2yxXrGy8P+J6ov2s7Dkz+X
JrUCYUumwM/kVddzTwSKNwhVu5bD9dc7bUnTmtFgXf4H3TDQklT6GVC1DMX2a6BabQi4zOem5mvx
t8tEMJj2cbzfcjFbK/a1pPEg8TDxil1k+iwXd+NUZhkJOqJiRfGsPbVqhD9yEynKAmV+VbYdQGwh
keQO+aEsMLWWyZ4NiKmMk1pZ3n5Q05i2V/p9jb5KPT/tM7V/HPu+/uAf8CdQeUekEqDQHJ7OROx+
2pmY8vXt+hOgxbSqQET1Ud+hCZnQRRvkxa6ikCKZ5xDu5+I26JaHVV+UcKm6G9BgXBXP3Jx1eeIb
MfTk4wxjl4z2osbVXMgoBcvXGqdUQ9HunE5JDvWtSh/8npeU+3Bvo6Ac1K2LJ3jHkHoIf/uezqiP
MNillEIsLDhBTyOvkwjT1I+JwTL/E5/jICS+KisnmtEdIsK6wlqfLgvbY0ID4BEe8fPZEtimII5m
y0glQpkyTs75fuxh6tp0ffyaYRkLfWLxh0G68YHSfQGloQZxNPfmoYHRPOg2F3rO8VSvhvwNW24/
in8YvxlpKTHH3utlhMouO9KJTkW4Gb7rgPanGbGoktIQ+DAQwth3bfcvzvqqYt7Bv2Mxj7i+setO
zMwuyW6/5LRbmm8/uaiw+/X6J33MVfM8VpwE8g5yzTy4+HAUBTofwAExCBgV+A0HHYSdIstRLrQ8
GFXBnIYo7o8KpUwyxplvlVUnvqNaCQ2HGb+a25N1iZzTpRjz4oG1K65JJEqQuTkxSjb5evtNtavn
Mg7JdD2/S7B5JptumU/mjqXe7LROucMmZT/JzOSKS3iDbInutyEin+4DBSiBX4r8F3t6W7jJVJSO
Pd3CM/k4FhwUPqmk3s4u+thSmxbTTNjsnngh+3UNfjdMY0tJiMWa4etsrrSUKwbCZe76L+HlNA+E
buFpXPK+tFMupOPuK6PF+0zFmPnnWDl4V+JB0EKZALJ3lMskwpawxNGMXNe0OTxNJq0UhZVFBgni
1NLE/kIkN34iwrDcLIqMYpwsUucFk0V0IPcvP7XlLtDI793Yt/g67q6Vdgv/noCaENFHL4fSd0eE
zzXjzBjXsZA/4/y8XJ5d/g6Y6ciZuzYobjAJ1dzmE1hKHGJUwIGsOQOCf7SgWbzqqeN7GNz1DFmw
E10te/8yawLIHII9aIGDdJiF7JwCmL1p3t9bESdYc2Hnt7pnX0dKnQ3f+QP2Y6wo83BDlwgEiIhz
dgEtbkmJwz1lUQEIq6SRmmlAjxcrw98FUmg3JUD06o+wZwukluSKC4BAQh7Bzsme6M3as3KUeyAq
Z095gq/lOQ0H6lPDOyoh9Q2+6yCCn2wJXj5CfnJZi0MDputvuiSwdpk+qliyfaz6vwuQ138Y0dBc
iaS5VwvN/z9muoyFPR3Qjal1QYBel1ojUV6aZtIfRxg2kqOMezbMQWejqw3M2ESGHeC3Y0phrA5v
8obGBAOeGX3nl+wXTifpq2vayh7Yx+TbBYVUg+g+3iwKofCg7GNOAs89NVbGU+tFjTSRNO0mF+lc
Gdpu2w3N/fFzKZqARSZZJcuHXLoRpk9JJCJSru5Eu7Z+HnBR1YSg4qbV5wEeo0s8SDr9ERCQV4oS
xEibJMeFPZIBsBCGuk3ZOk+O3cQw6Lvf6bRegbFn96JSZXKX+CCgNtTOVfyMQ0M9YwFJ8JtSnquw
FDIN5UuzckgfnipvG/8T7ovbMc+YsYxozR9WPEA1LdUy67dFaKC5llM4KJZYYW94n6YAv/m44HaR
qCKTHJnCgebIKFSX8DYDiavVtUx3wm+WXDZ9ARvZ7H9phujURC2J1K7wlNvndRheupEnJd5b5jMD
68Me84D7RuBy8ZeaBvoTkqgCSOcjI9IAsPxWcqiPqZfLEh7Sl6OG+f09mq5o3Ez8aopz38CDNWCZ
GF31msJOQ8w6jS3CI70pyof2N8vSPzisx/wcI90alc2kS2soX65Q5LbSPlXtIWD+sq32j8cZO8s9
N6UhXi94dvJal6IKREvFif8jWA6HSbYYcc1LymLVAsXg/Is8NA7oOmjNbqOjclWRMrMsIPJhGP2b
obeckAWaBD3K2yiLopjmy/6oktM/BnYxdFGRswjczKQ2nX9OZWqbyXTIwsO9aRfu3AtzpZxFFcIs
n6gMi/jEGRvohtI4NighXrlNgP6PiUmNapK/UIBy6UpD39otTANPLPuBnZYRb79HkfXMGRMcx8px
P/jSomE4ImZmRR3m56YDJ6WIMk9bYDduFuDP6a7BCWje0sZt27F/bwd4FL/cHmQIkHm/2LCA69Is
vGX8e4AeqtkDbj1z1Zp+71hKLWFjfbFX1Oe+8kEWi28cOn/uMquIBPtnsYpp3f2znn7VtEbbDin9
NIVdkm2HhczMkTvaRNj4b0LLoasAoIuwY2cw6bNAikZHHZnRs9oNPfprryiu5wUKow8pVBCl67u2
AcgOiJarUJYuObIgMNz5JfSbm4AQ8klvwAmyxewv3pdhu/iGkhFYXtj0yzRWxMqjcgZkOccNfVUF
GfrKQyvtPvsHQ6/rdf/sT96or5TXm+HqniBsc6dgHCY7iOIt/ruCXseuCKjVk9jTuLcJWH3XMsEq
S/9UzOkmmEXTmlWQJ2zEjLkcXc81vRCmVcJfwUGDixxNQkFN2Oalc/f5QEalDgX89y/9GbHC6r6G
rAVDyeGR12FRoz23gUfjrcAtTdXdJkGCKzdbSNsDhh2v1bTHBJlidO153T0djN7OK0ZjcL/aqQNd
vkSeuY8oZBcE5pmn3tUZzdINMsVNRu4kZWz0kN8WXVEPoBHi49hMv23Zh7MbK6uF4bQu5b3zLcrd
qWuif3NUkPHfEsmS2mT3jriXP950S0sFo+x7pdqPU5GswbHkHJlDNTUiNlqr6LJlsq2Fy2tpGIqk
jx7ThLuRYTOG+hLuXVFN8P/amKG4bsU+wk5F6oi846u7ytFsVrsv1E1bq46wX7QFq0q+jzuZfh6B
WwYI9DV24bdWWGgGcCmm6lUlKhKuOCxk2+M1BcVfZSsCYoJ3uFv0OZUWf15PIG6VdhU0ezyIsR2V
bbrjp1Prv7PubtemrvkF9vXfVNhE7mqMYbGsxrGu5VnilExcXv38ng56QVPrwXBo6Lj5/m1k59s5
hl0HJW2IEuuwRkA06BR7RbZamsqr7Ydnn9ZZuhuHUQV11n+3YntsIIOULrIY3L1zzwf8qnvoNzxA
iRtCX4XfVwxd3BD34SiEtu4N3Odb8nHGUPwOGUf3PNWFBUYTbCsxlgVo/xMUTbBWEw0tAl9UH9B3
Jgkeoe2lbfBgBhm8daMQOjeXLjWfLW+fxtpznWQZ0qQecQ1xxmj5OdUro2oH7C16i1GLyHOmnDzv
/VbbfmVHWRQx4IIwT0ecIxX1J4QsnS2HwJn9sVu+9muxQilJgZjjoIWXQ+1WRZ/OTaNROnb1BTzQ
1eoKxA6MJ3UCrehgbZ7Ms5Ps7DgAa/t69K7+uaeLe3NQK7uXFSsD5urfMcoWLGp1gJ+nKhuG44zD
mVIk1tOr5KedYy2+eB5OuTuhDTdFZCmrcgccvN/qaQZa8LXynqGcw+kxyaq9h8ROe+ic0Jzt4bzO
P+ofDWokvOfQBW2TgsV6rtPlaIjCnCUHa1L2OtBtgK8dK3rbw2b252zu7Wsc7kcMRt+HudihbWLA
l8D1HrEpk5c7IWsSfnc0UowQzO3/eiDJJqUnKGAgtVK8ODMFJim99ygNWv6iQy461DGHVbe9pzui
t+oqbUCh2bqW9l8rFBXh2ydEsC6Ib2hG6hjvTv5NFBm1E4W84VQvDos7g5QcNq8WYN9pIBnLU/rL
F2P6xsRi/qoadp6T0wIwt2vXO6Im0zmMovkKsIKcxVUqbgcsXGSF9ja5c646bH2OhMtS9rwfCZFH
PaA5HcJnAqLOe+4bbbefVLEmKN0oNrknszB3MIrmCT69vnSfnw+YLDfnqYsDfitlxlh7eF9S4jZl
+wUUwtzoVdbJ1Va+/PC6nYF/au4LX/OpvQ/8m7e0nfck5AEz1mLp/lmIoGizbOM2cDzfGRrhubqB
X4+ZMITsdWw0ALizPAFqI2CwTbZ7OXKmz0EULXHgP104eBixpbM5zKReL6ZLIzCVyUCiLqgyr7Tu
2L8KYWyEW8pd69KbXRkE1T9oVtCnwH6lBXZb8Qe2km+/OyK5QvIBwF7q9kC1Jqa0Lnfhg7lpCTZ/
ogiUymylompAoLdmm+ecZhykD2i6ppCWBrKEuJASYr3DCjNCCkI9u24rWXsmTtgzMFIrN/tLZnG6
5hEWhBfW3QENur9Xoe5Cj6yJU3ymxjCEArwtrwgBwm8kVCLydzxlRM66t3UJH7rq8YAMHoMfG/NH
ciZutcZpC1pwteXUVDzaWWVrRjrbJCWX+3ZrKnP0BprnDFFUU/kuMqZTceWnn8KZ8ROOnFE/aRQ6
yslbSvgv7pin32ErID57Wa9XJLPg1tghO6mBUtBFfTeJyamfHq9t9qZj8hr/MN7FJw5dJxJeCwlj
0LCHU7tJkMxaRTtqjy5LitDQqEkdonGEBDyHtLmpxq7e3LxKb7PzCh00eU34FpZBng1lUz4Iet8z
FtKlXduB/27GbvAA6xyXy4Yu+os+jOVCenymN2S6rjlV7VoQcbyN3YV0xq1UjjLp3CvcbdzbksS4
ShBU4M7T1bGlS62Zw/0KT8G4TIyI8p0l2d8TitfnidUXX/bTxpv4eQv6wgH4AIBZA29Xzafcgkby
519iewPMB4IPKaG0eTBfufewVkAZSmkwimQt21w8sm0/61/2Jhb2jHzH+Pl7In1mjmalRkFoQyfg
1mzkTmRegrdfpoQvcoNliOSpykj5rw82+TJcdmoHmYCBowHCVSWxMuM+TJnQzJsHi7p643/ct0Uo
+5ffNHf/dHasmjv5d51sMCj1uOKXBKuB49X4PLqq0nV+KxepmaHOIOkkx6e0LTtwS3VnKZWuDD9J
ORMQMIuN63hzcGI7rcOTO4QhYFAd5eyG6Q5XswuTgo3PsNsFGaVfykgH7quUpmjnnJzLYC3CdnOI
zkulmemukHuq5NZMtxe+Wn82jw4xwMCt4+6HRZraRrmWcuxiFSW0kZrg3r4MRgsRIcWuPbmfSC16
AXpDTP+ZM7OY+T9jZeGYFwqQzNxW3FnzeyzB/SpPa4XM/mc6O5UmnRtIapagKrgCaPGQ64l3A2Nu
up1ZD8Ov7kJYmNW93BNfzbx3UIGlEedCQ9DLWfa4BtX8UtqrecGpeWerkVBUrHvdFV/vxLqYy2oN
c7L1iEPN1ckDOIySKIEls1TGmDyxkbGN0HpdMDhfTxktL7XlN1tLubALTHpCLk/xYc+d/2PXX+Y0
l3+PXXTjmP5/SPDISA7RU+gD5CrSJWYJyLNXfQsH7bCBEw7E4P2jI2uE9EabTELoIxpWXfzXXVRS
GhONnqFUi4u8adCFis3JFZYL2pgIbvRnJ2COREwlmNorOzP+1P0TzqomobpHp3XN2kDkNkLeNgXs
EDMJ2x9RztDixRfKglr6MqRFQ0qSOkTJEPMfVxBJvW4/Ku3EifD/ATnwFs7nJr6jE48Mr8g10qfp
j/usmucbhdFRYbCK6MS709E1UbIcc7iz2+H/rgTWFAllFJHmsDgFj4yBLEPviFnkPZhCbRNWqevi
0ZNpVtDNv53QyiLukjv8IWs/1FScQDZFTMInsUcLf/8A7Uw3CTEor+F4+yDLDkv6sndfajwFFbO9
klFUBVUH1sR+Z6XNCdCiPwi5uTIpd1hNU4ZbbbhXDaL16KDY63gWBCaaGj6PWImHNW1qTtZ0ClQ3
1EqQZFVyRXeV88Qc/un1FX2HInOohUaa/v8MxP3fgI4HVQKg/ydqpabolNARE8V2UFnl27PuUtRz
d1WTEnbpzFcEFU1Wp6zEDVu6X/8wR4MKcZgIVV5tKsUxYcFXdOzvJFeiCusKXmIrgnlONOV//F7K
sokspqOw71X2BcKj/EHAInG8IbPxDGMZtQHbVY4NfVpGFkrDFVXPepnCYe644VFRDZkWgA6pZjX2
/bBFRobswdZUWP2w333sXBEQjXdkLeTba0gNDgAA4cDDIqg1Xq0cUmzKFTsKFkooiJTTd9MUbVsR
+yDslPmaEJH/R8nXdQ9uQLtSM1IMfjLXcDJtwyCLwQEsqTAZlsS6ayPmbVspR3NQ8INWL+ZjTdUO
ZPJBEA2Cb7CxlQLD96zDeticdvroMSn9lWOAJOheUNodZotWxcGmPKJo+4M5WtApY753V1/57Xbi
0DeJ8jel+HzylOUGA4vIXfIE0VUhuGaArdTEOb5jToLWCKGIgANvzBjHKNxdyeRWJaeNqzpwLbMR
SYyBsJalU8/WwMVxrW6E00/il4U5U7pOLdExLuJPMzPNVSnTQ+R4Jv85+/4feaV9ROtO4509oGrM
wd2iuUN+fY3pDOHD/+0zGrz2GvD1ygOI3iFt6tW4VAdGQE9BHA0gTV2DM8xYISNeQFONkdNdVdcS
Y3C21hPgervYrjW0GAgvDAlTDERhsAe9Qlxut9DbLdPhAFY+xgQh+MjF6cPyas6YJ2DMmOem/HFp
kN9UPdEAeFq0M6POmDgUsQM84TIYsxECh2+xrPXaspX7XGteanOcjKoR8GtpwxfklN0v2aOXeVBW
pnw2QurOlPbDgm5+bP1FIsi7NEjTvzQhYd2DWIx2WyzCNCEYy0gxYgQrp77gAGd0sB2B3RWsKVRj
AXnNxVrIyO3KBAiBRUK48SaCgPiaAAO7fiNpsJt+uCJByRzcZ+1efWDpJ5MNYQ5MW5Nnk6CZR/I4
OcAB5Yi/HbtmFnlRYlx5Nw6SO9fRMUvm1pbNlO24Jc2a+3sIE1qpWt6tYPH+ZAqYfnAnBjqVf4gW
yhIGfr/JvdGMuG9iCCofHllvz+igOceHzR/sEoaNc29jLNN/NsnSvHLtPy+QhPRPtKknQjrnfvYf
SiLnrwE7Qz8lpzhO0jRVeANKktiBPCm5U/fIissTE/BBe8ixCQDGRiSB+T4xq5T+yDMTUmxmBOb3
n8h5q4E7X2WBpz40/TTTmNb5OdVa0RvZcoJm3pm5ZF7DpOLf9VieLOI315jLeErYN31VtbveB5qc
eca58tUw2YZklyezZ7IERhspKv1oFcU40hvY8AMdXVnflKP2DhJF18R/CCeuOW3fVagsZYYjH1X+
bcjHRI2MHZz0QuTdVMpdAN4c7rVHCGabvBz9A6PGqYBNIdinBlYgDFmrEKyM9l1HBn9ra/XQFtK/
MTHZni8gg1/Bhkh8Z4GR64GfRWY8OLX13mxmOh6dkOrXKTH3JIPVXwIVKV6QnWu+UGZQlIGlyPfR
JN520Uyw82t8uq55qgzx5UEKbr73vX0LujK4WUtcqKm5diNDjGpMFCZb93lX/PfkXx6yEcTXs48P
WvoEZmk3GhnjAXlfY0U2bCdupC5fH+eCNoq6n2VfJDubh96eYjvz6zNNNZqLjrdgX/ZjFpqrvcgq
tbJbZ7qJ9WuKAC8Nlkh0L6oPLGTynZ1m5a5hGugWGyfVVtcm6Ckl6OKRcDnONEvdllxZxd33TUqV
/H4TAfN0+GGT3PkbrKdxNxm6mTBpu/e6wmvGmJqwkNlxT3n98asQrwbP+TXC9HcQu5WQfG1i3pRw
wuyDKJTBIW5YkpXtrhlhyue01qeNiwXuD1IaxHtOci7ks5Gpb+aKCjaupfvIWrewyZBv3zaHIMhb
gYJniEfu2QzPNCT9d0ckwo+668OTgvKkNHbmrupuc8+gZsXEw5F+lGVU9zKBbptSYiFxHEgr5hJw
QWznTqaH9K2bYP0DdLB6tCUpvMITjqCu+yMJES3xrLdGTAYtbYnDMbqaAp5CepDj08Hh8fvY2Ups
W+ONxBKV65U35cjq4ezEXuyb9Aeu3ghgfVEW/VWP9zOU+MHkatzOy5rlv75tv7Xi7lkroG6LUrbf
jLnTTwCQR4GHQ6n0Od0SlbJmrdTiMn+7TF3336sFAdIJoszQRi+hMz4wEokVTL0Px8p6GSlJ82XQ
5aAOE8+HCoPR0iaR17+IUxrXlLRiHEaUWZcNZ4MudddAc6vBM5QGm8WJ+ZSr3b2A4a5M7Qv2eB8W
9UDZsou+B1yBQEy8duirhw2PbL1dEB6FWRGIjjYcMQKcFlDG23l6TKDDa0FJgjEWKVb4IvzwuhW0
mkCCsglGJp3/V7eKRhFLVrgb3UyznK0RMZ3VSAmMQR78oAOpz8BqVsBHPzvBD81gZudl882ynMZ9
N23Je74HiAUNM+niEew4F7M+pbuLvlfMxeuW3iP7t83yM3ok2H0sEAbKSPOSNHGR8w8Q9f7rPTKe
ukPM9nKeC3B/751iXsbfDHdNRgJ4U83qX+QB7mLR7g72D9ZYVSzwfxwGCLXDm0UGOLAxlwhtLakD
+s1aBcRyncr4h2M0aen1memc+4lSUzcTW2bjjnIqGQrbhSeTLpfEBwfCOzeRpV0RhPK9Hs7cmS8S
7VrcJTQZlUMAS0+cRErDKyZVmjamnei7NX5I3xe3wUEOP3Bz3a8Vh28et8S6XGgTgvB5ftwrDzH+
d5aOBTwpkIEgaTwakNn7boG7kPepPJYcrwHcFacPUCcPsC0kBPT3UZxz/1ZwI/zf3Z9D6cKFD769
Ly+vKAYc6aBlH1faYaLSX7g8qm8a2vrpgEG5ZSmT15dFXe2Yfw6nVJLjATDx9wT15Xh7Ww+x+bzi
+Uw7TovMzQm9CtBgi6rgZ7rD4zjqijBzh+ugy2cuPUJ4tUtLmXXN1DtiMtT1sQ3M1AJs53/rf82L
UU5ApUSS7WEnxqsY4vOtFxCtUc5lxq2FQSTLqmqtFu5NSOwqpeDEl/05pP7bNzItqwmX9f5tOF0u
73i5pJUuIyQ6kuxjejrduqNe3ND2f5s6mRbqW5AVtKZ7FtXfCu5NxjNZCefCbgj6UFFWflmbWkah
pjZzeE72tVWLcxMYzZqT8NBo1e9oHbGYnvBmKyPRfc44iUfk8u7nhlkXNXeBAz2HQP1bU94g29CK
Cc6KA1q7kauubajLRo2Ve9D4RMJByE00KuPYbh6izyiiLpn2tKRn5/YubgD5c2TmkVIqZiZ4hZmC
jnIrhbmc1wvyAwIq9TC1CWxyC+29CaRtoSZOWOJa2A3j5Ctrvte/I+HyrF5+l75NgKDg8lBSK22Z
9sGZj9fA+SgQaGoNlGEwkLYMGO6eBGUb+aAn6bi06YCD/4azWqVYN1pJ/Ow/izse3Vyyiy1OYr6Q
7uPEwVp2sfJSjOaDTdf7uPPP6T1opgvORTNth+ni52hr/URhRk2Quu4sYf6w43QXWhqOnVhEFdRl
mJ4jYSI8XtAtHjc12ioM7aUVy72s/WhzlhJq3D3CMJVnb7WaoWZF7Ixgv8mxUcaHWQVgHfS5YAIJ
J3iSwktvfNarllQAbiJEvsxZgRYdH0ZUHHvMLSi2eWoM5leZPDfcolnJyYv47OykwENofdpbHUpa
uD9g30tbtFpRmYNF2VBFncFQqCHD7jSRW70l97oW0cVF3qkeejmcXLh155VuusRVsIcxugRhGLjC
5q+lcrFVR30vvvytx0IOyFGTbG3GwCIoDpJ2KZINypI1K/03y+kV0JEjhFE9hJw9sVm3TFcsvFIu
vFYCd+lrg8mYNa5IXVMu0gTXZi0FNpCybS/fbVeNekclR3c/HvFDHV0fNyhzEX+E+b13Fxho/7Pc
A6zdf3dgoSDAEQmg4ukmrVMCihMHu7dwHPUOqu0egfOVfYI0aWM6azwTtFMugB107aRm4z64D+iD
otlq0aWUNSng4E5V25bUDmRkdkNLpWg0QafFevgSplB/OlNQyOGgMODS+ZZTEz4ucE/a0cY+xK1g
KSNY37llbY1JZiIKuLGUce4grQa3NrcTneidfXA5NPjvqYkCts3m8rwSFYm1AKjHkaAZaClMv7SO
4GswLilM1qwn1qLPjlhwc2lhQ82aK9yZPnQqEJhurRwPPFBPiVyfSfN6O7kTxSSD5qV8uqGtliqn
jgGYpm0z6H/HJpyx5C2ERLx4DGNMxJHcbW9la+j7sJdRKFNLejMveFaG9ZBLX7LW1aW0iBs1qAzu
CdBUE4LmSNi14/FgvrD+4Ebj2GhuBfhzPPHFyQH5hFnubiHfg2//KzJnsvFcXh/N5fx8vJyZQet/
23IRjffoOUfu78EYOb+ejHrf7c+7piUj9RcWPVdK9fGCB+EahKMMPrVKjE6MnTcDw5/4zK3gZ7rN
Fh0x09YcA1XhgUM3M9KmuEmCJ8/8dLFFym78BYzXfBx8tBUJTbi0Fw3P3ltaE+exp4+AIQXI4Q2j
tdYJWA2mISL3arOiwO8uuBsWoEJ1NMtycZNqHrwn/JYg3G6Qz1eaqwC3qKwcAXChuK7wqlFDFdap
DqYQtTBzEHhRk8LPn+G0cyqheA3H9X0GxSUYY0YpBa8E2rl0WQweIXlAtr9woH+rUO9atoYHQI4n
ZaKKu2EGp+9UJ3tvYLvZSzZwllV1vsjpPlJUm/KC+eyOarat9Z3pSWabb7lDlHzZIzrynqtUBe7O
+Jhxr39TdImpE2T9cClf4a7QmSW6cq5AHxNEK/hFSmrFsLW+UU8z64ZRMN992qr0Yz65HYLHUKJ2
vavs5YbGc6dtC2/tshtYw5wpvlJS2EmBfcqvSaFvhG+VqkHnOmEtr9otW/boAMS1DxcVNr+XgIEW
v95LTebEeicfbTEQIn/s6soWnXI2OC19eeSM0izvOX/dVlbUX8O587aC8syp6IDTCqpd9L00a1CO
4NFgTBRFQn2x8kM9TkcOu4EHd8JEhds8IwV8hL5h2v8FGJY77PKU9oLSE6fl/p+QptXwGQwf6gto
hRUBtcKaFwgtWxu7+3A+qi1qAqGhFAsT/6zAkUtYVll5bcQ2DCZCRExiq0JUhp4wFiwg/kSuI8bo
Bsr41FPT6SWV12dTE6f4hyf9yvRFi2bCyAS5QO19Gyju3cMamMNxKzUTiRgO+OHaoR9dqwcKEJHm
DbfkrUReeQyUfOo5eo4Tl0ixuIKz3dEEGFfyNLvwTbpLKrjl7n+TRayDJmLKeb8FuaQLSQxtfpEc
H8WFluwdQ5K9a9fovpl5doZ6IVkNXx1tknAe8NY5QGC4E5HBBtK3o+7LKPArZ5pR72XTEaaaquVY
EhUbNX81DtnSDAGahGygEsAlepYTLfaQ5L/gapo4h3SIkYcNvbXJOrBBeVEWVIE4moYoIZYEd7OB
rDwArXwE933m56MeoCUBPigTsourdkljeHsbkoYlaed1nsfAZl0ZH3aFx6q2unjcCbHLB7K7xmUE
0DONN4Rp5FZR8bfI/reGs/QkUM/DKLeZ9FbzPpwsGFG4IWF1dgDFe3gw6GR0TIZ5oeCP9jlDfI3i
fIQrmwnBe7+cOz77wjhTxR9va7zQk6Z2LQqQc9dEPUfEZaM0T3tcqJmXEf+AllbsAgDNsjpO2ogr
b5mlD21ASMNeMvvp66PegFSNxJKbgtGvnKN2U/m7CsdBJi8y9gniPIOu2zc6NFgAq3paL2uXFdOa
WStOD3t/mxfbDEXxFY3b0ozL8IxKzk0LjITcUpQou8jcJfFTHzwCA98hgi7yt0rH71OAnvp3Sz22
kclJcxev8XF/y5WjfP+SjdFZpy/XBtnuy5E44dFBBCOebqN5X3rXXKY3fnLzjPK6M8HvKUS7//Z5
CwqXOTOJ9aPqTAa7PsvN+PQNMSOwAOXpKk2xEIAREx/kxAQ4FKsy2Do4+iWK7bkFsod4XPJ5bif2
u/trw0AxSSBS9AvUTwez4aEhXo0aYyax1EeTmR2BwNdA0OHHrbMJ2F11fe5Ik21drd6pFBqJNjJY
iCsSDyOd89hjodQp6XatSWE4/4diGQ0hIGc192ttLBrCno5LzbP6vcjWn5SiFYpf5Ts7UzPhA+Hp
4TmkqpQs3sNNOy7shEEG63VxSlfQdaq2jos6aAH65E28ghL4KYntfVEg28K2z3RAZYBXkUKszW9Q
Bk5WyM3v1+0Istb7H2hplS9Ls5eY29R17V+qGMCUfO+xhrs+FkO665AS9BDbQjGkzRmN+HI6elfs
tW31kaCiI9bh3QmUsC3uAh4VT9tr1DKNCl9crbl7PDOcxP3pD2RLWlu60GEeWxLe2/mI6pe3rC3p
9HtTwzW3RGKf9f1EwuY1SgMmOLRHM7Q5Hc1BEazgNdR39uyr4SNUHd71KH9gpjmjgr1SP//RP/lp
EQ1RT/E8m9YsbZurbJ0u7r/xz7QSW0ClTcF+j3HTufmTfx78x0O1WAzW3fR2AvikAEoSVF1XVv77
tj8sxjCCnC/fa5+o7PRXH3JeLieh5C6lpJKhWLazUPgqkgluTXT3WS/g4Hqwnyjg3aIO/OttKSAE
WuHS3riYvm6C01zyGS62zr9rQX34fOixV3z4T4xkXouSYZ/mgJuCxJdMis+oN5iJbom0p2OqnDBa
NG8+fBhKpJ2U3sdeann4Y3sQ3yp6JcX3wbIW/xbaBHz9fI5c9CjrhSjRF5YXkIEZK8TW6iNu6/11
uezkW7WY/MuR5zY350HNld/7zf1dL7vi282lWoBLcuQa1FZBSSZfOdcxjxPhyd7jyqQRSQatc+9J
YN9AeyMrOYhOhoZQbco3eVAEi2asf0F2weU8dVrDlEFsMh8CGx6wkCncBtd8ZDdY+OaBl02EKIN6
mhFOCIpLmL1BpUnBnAguKLbLrZxj3HJa4kPjLPszZJEEgosCz61MRmc/gmgEUy7MzwHDQKBvZ+fN
bShP3PUsoyEJrFFtPNtiGZ4GlpOybpwLylPdUsTEEv+Wz4HX0CBAWvP1Ppyw44esVYEEfk4A9/b/
j7Nqf8BWvr5DIIACX3ltpnb26PzK1GrAnr2Q/qo+SAob0BOfjEN9Rsa3sEGxuCp/ZNVw9+Pk36aS
QMEOV0sKqps28Bsq1OB/eGjyV0qeg0uVm9Sq98LvwEga5VRLjcKtM+fWrVCwsihD1MPhVo79Who+
RiIjXSRJM/ot5AtXygUE7plOLsAzmR1+eGuP/eLJrQCqGV9AiqW1eQUUOMTzRUrm5sPI9ZfnjhDj
Kz4PFUIDsKtFT6h+r4JTnBwfwVzQx5m7iy8OYQi/UW3oqm1BfPaqLZTihKLa/MFa8oGqwxN3cu5c
P7zokT8L6igEHYBwsACob48G/GjEFjbHQlV++yDXrZ3SUnlc974lh4wa2dP7WcKyCO/wwnXAFbX/
OTH13uwYvE17gzKXup3veLLm28fRyug6K7cU0O/mFy5+z75D8EItd3SRSOSz0CXGtnlXvyoO9Aah
QvmSP+atRwINersuL0qRWq+Ojamc7KHMWtcG3sIccVyBUjQ/qtprxQjsGt6t3BUTzmMfN5Em+iCg
uYfuF0Er4C6nkgCE/RnRls/Bo9heOFgJMAhdVMM+oMlZcrpe3lDU+Za3PvUZFplwxp03HpGEp55s
HsFx16ODnIZdofJZcrIx7LHvHjIpQyFp9EP+VzWZuzmO9S9gcb9MJSXfgEu6Gk6JZUwHTEka6+O+
4xWqWl8SsoKSoP/rIHykbU+MZhm7saQvscK0/QZQTHtGMvFRLEfLL3I2yrgzwfz/rJqastfHHEIY
kRSLGmf/PsaT9jU0tk4CssY3LaLWGV0gh+yWTQv5A0Law+BtIMqpD51Zja2hecGFFfka5akesevL
z8eyXJQC5+umFqfc69TVvnjNqZbvoX2rJwqRvfygEJrNZ1/KM70JdrbfCKB5g/C2xzkBVajbE6Gl
+iMeF3My2ylYtqEIU6tAmECOnFNOixGrSlnDoEpXvqWsGaKd85kr9tVvdr5lrGutscOwBRenRDzb
KkaLVnRzdSzPN1HOYSTikjHUYqpwkSK0yAl1VTXJjlGCMLM05uQUcE+hYcsetBlEY5Ud8tG12LZO
Dp3Wyp5ALcefsywgHz0TTB9MNJzS9jMmRwgYO1mvfXXiIB75L4IR4jx4rmEZKq+5qrCT5ajmXC9u
BSbsd8OF33Vq/AexBgtOoOLvpIZGw1efSg9nw1xq4Ny/lP18eh4oYk6VxnWtUSlS3vGWX7vM1g9q
ymkhK+43gIgM171uVNe9NVi5FYTEe60Cy2DO11U3ryP4rgqqrKu3OWXU2Pr8aRynBdCA+UvYHLpp
R34LD1FxBWEqAxuILJSsOwfFQ3l8vUXeccGVywcSoXScxSVt+7sZWBc/zkCvDe+Gm+2uyHq0SW9C
sF99MAQ8zwEUivfIY2Dg6g9O1ffJs1AD7HAMURGbv8FIKAyyf+38MDgiTK5m9XPTLRDo9fZq3DtE
sIcMiL2QxYpkTwPEGQ7LcEetaLhw6Dk4PpMIAVhRQjjTxSZWFC2gKCLnndkWANTwHn1INEzOvZoZ
enwQ4PWGz0cFALsp5ARKJTBwWPJURvw3Vz5sKNS7hb2Y2si6RLdY/t6NsSR1USiKv+qvUjIf8fkT
JqFVs6FgXE61Ax/P0wIM2t6kH6E61QzebRrznRJ4W4bg1qDXtFbzjprLeITX23a0Rdn6B5dMzJrd
WybWgxi/KSSLv3wZeHMDJfMhzKtN3UlYgvVegeGY5dDtGQiMhU3X/Znf51nlWAuDebsakhPwzGOu
XaDYSso7ZjAzBtxYON7VY/QEa/rFVMn4TOCEKW6bi0Y49IbTWlfQb2Pgy2RY9eC2TM8dyNZ8Ugxh
RadwDhTN7uHT28driH5+6SGpN1UB7cIaoAzyZNDbHyMWwrHTnJT96gCwLtccEstKb0D3SwMgOTwO
LpAXlGYWAiyOKXKAzV0if0yrsJSru8BK84N7z0tLJS1VRXCsQMwmynjdi+jefevapb2aNF27NkvH
pUFNRUibHcsBQgYGZonEhYS2nN+ON66pgwA06Jl8qcb8zYlQVy+CAKuoTrNYJkxJdRUIrHzvpONx
GMzqBYXSKI2z/tYCSvEaozitP5sSuvzsMCaWmNqey2rncuY6Dwf/gEx+U0oCqu53RVB2n13rysjV
78ZcTfcruzzxrqK2W6I+wNGwb+fbPMondLbgfeazq04kQ6SlWZfwtROS/igd4WJDatB7Wd/gJ29X
cdgG+lVb159GgrLh3Y4QeSYaswqvom7h8f6EC8H32VQD4VsvXb+L/yExpe0ITiktpLEjjiDLL4uz
0GbXo5vESz7HKotC65tNsaGjvfDdtFvciapK8sKnIOeJveQC1eNht1hhOjWIfcIKNdBezpFeTrZs
PuRA54y0DIrUJNrC5jxO1xH7So9+mAQ/zdEjazAFo5p65gOIrIS+46O6bK12F02w4kwB5PU70Th/
5StG2zJdeATuTHJ48Jw2aJf4kUUWSkACrbbzx/MQ8vSZ//c5W3R/nZ18Ak61Ab5ZyhayLWpNj142
MqItI4c4I/wJEqrwO5n5CZNP3qDX9878GMay2RK6C5AusRUOCcRVhAr0jkgqz/l6AeKLXMVd783L
3/i1jMkimZJvNTdFGRYLvWmrBesrHZpJRC+0/I7FC3xs1CycHozLV9uZewLQ5uWflGH6EGcUbe67
mrK4r2m9pdRF4yZSYdRMAkz/LGHtkyJLmrZjPNI6CGcSHc0yIyg4Gs2JUbxJog00BQY2KxVlNNo4
6oJftQZciSam6dgJTvdCYnPvHT+RAFBygyxwo5syeXArdu5bXCLn4G5fDLLkr0AkEN/dwvHcKlAX
toL3/Rs7VRoe3N68sDObS+nuBD49yUhuA5NyyMCe5rf1co8nWGGZVMphfVTftGKf29UQAfCC4U8c
zk6GvP+aFWHTE1t3O2zuCpgQCiTOIS8Yc4ppSNiI8SavIHVrld9gC5lQ3E3wwZEUgjCO6ppVqp10
bZrhx5hTnn4VtaqBzjlshrs6c8IYhPv2H5yLVj2WxPCQGV/dH67cA/QLebMtm9PgcOniymdlSCvu
8By/u2wPB1dntlBf0sTiVKZu60Jl2J2ZRz6Ab03AoRRyYJEslFXMz/ntpe4M+Uh1kBvi4qtQNP2L
OuQbSL4g62+MPVJGelxd92rqqJw2qnG4DSYjenpy4m4F0xQBqdEwKfHXNxJcDXIUflqcZK47TVg8
g6noWXutrdkXaBgpX0DZRdhJImi79F9u03RYOSWikdMswjmIAc3FIcx+eC9IzQwgdMPzS7T0Nkf9
g1ve+xIspulvdGqtB/lBtwVa6Os9KuP0y7arWT5DPw4pazQqnExcR3RfeNKIX1+bjFyG5nCqtdok
mW/hWRAUOX/M4ZGlNagYPeKO6H5jgWNSPPgVylNL0PlouJqcV9jeWtXyauEfem98erl7ihzfM+kS
WnFvaNR2glzxFXf8YklnrzPsDKxZc37mcTkjjTuqWqwAvWSN3iOaFJWPhZApz1vl4QS/dYjBCT6N
UEyChZYAlrcLzL0IkKDPB0iCO9vB5xLwKEiUIuuCpLmcjZPUm9RcjFpevLVGybv78kyR9yneX65X
vjh6IF14ow1DIlOwx1iR3N4EnSKs1hKMWAI/yuxgQ1zS3Vna4OEDTig3RwEyFXa8TCXC9H+7MfR4
jE/UtS6XnSYnFtNPLuj1cKF92PSP319VnW4pYiUeVSJvQ4TtwuMitY0ph/doXPUXMSFhI7SD2gDn
a5f/eBdOoH4X1oZ0QjoCbpsqbBihB0FK8N2Ke2TbFLW3dJB8Msusw117RXVaPDZaRGFyy2YVzvM9
sNjLcrlGM7SpRZetbmIzCF9GyMzGOykRr418qb2w1nbAY7c8NFipCCqtGvhci+b7B+VbVPUItvbQ
87sXjTox6t6TZMGeeif7pWIw+YGgJnJ8x8yTi20+UG8YOUpfTWmXpcrZ1mdXv1x+DYRWdbDq5Fwx
5y/VB4QLCWPkW+2Tf/GGjtaVtAwVreuPK2fK5hGRn6rRjsRvWUaUsl0FuFB3z+dCXxULQFw0GZ+d
kYGQdCM8aPwHqx40Bob6ERqjAONlEXGgY+aFPg1y4/SL1p0W4hrOTEQEIAtWXcGBYs+fHvCPkKZr
5l6fA/pp2IorUghdrdamUuKziqdqpQQBKgXKaBfYuZd8dA37iOhsFSkkCOLJiYgxDz5gwdJpOZCZ
7ubaAlV8v+lLrXZPkOm4YnHeks0u1OZ6VBj7qiGG6ONp5s0d1aPN+6c4P3PW6C1DG2zJxV3B6IDr
6h1inUetXVI2jIaM2lM9jEx4FXceUJoQOu5sEKne9btj0iDaCaw+Fd2Q1lxVuA47MMQ2TxRDaHMe
XGSbZ0vpNcyoIuegHG1TKzVhcBiGFcrr69WdquvU2CREskO6WVSwQC0WJBwwvkp95zqIuSq5coFV
/23vyjYQlKwUgY9vx5V0QMJt+i4MpPVl+MfNxxfClrVAhkxZkunnGNL+MJ0DzqnloDOLzB0tAUBX
LELPztFzRMkwvVVA3skBt7kJluQKnGUxoGPaPPRlCZxFgtXMyhK3wbhxbuSrXH6dSQD/OFPXnIe1
710xXyG2Ypt79+sWV0oCDuvk6KKsM+WZqUJjEpK+FzvxgCNQ3ZkSAaq94oXfEiC2VlZiJ9Qfefa7
rLMRu3hKEwFKR5kf5Cw68vG1AkByY10UTDXXQU1J+tGg9F14bt8KpWKUzlE0+t1hFEqkGOnaHOXv
bM+RWuy9maOqeVeFkBl4T6OpxOWqQoiaIlNqhLyAfo0fU758RjtTIHffh904Ot6D1WVXAVaF34RJ
aTmU8rux+V3tRwS+Nte4m2abBxyrXpXwb1nXLywv4Yw03hDXecSzgkM+8vSVC5EH9JjYQMd+cRr8
lEgb1WOBF02MgMCywzRU1CuOt3LgLprfaV1Vocx3fGC3MoBwbU3QvU3Kn4KSDivURK4NYXPkEXyp
zMBoyjSa96Uzk8q+Oc9ZPhtXuYsw9Y0xTcksNjtHhwirhGrfRMREVUsXJOIT08FnXTq5vsavVw/f
SBCH9D7KTOtYvMDvwH7lG4oquvhB3laXh0LEcWZHPfmQCQgNd/YzwrERY+lWg4k414f/YoZzb21O
ELE3WiF/dy5lzGgnsOyaU86vB8aiiTUm2Z0HVJcMbcIs8Ag3noSmKpWcZdlX44f5msazvkP7Dc4m
gUuI9j54QnOqUAT7XAjJ/EtwhjT3SDjzZum90MmJl/URxGRbr6gn864saxww38wRli2fu172LMeW
VlryGzk74VsW/cVApILX7LMgXpdSBSutLkvAompgDg2KSqQSpm9PwFRt9+Vtcz/NSRaULOruKmfM
aKX5hJC67LX3YRGTHigY6APMQeTDlca2OhfnKqaH0az3HAaTh+8KWbZny59Yj7WkJFh4rSwMYg9L
JmYxiOXbAFFqojQ7vulCB/zzDj/MjkuLaryWlv7HhTJMfVAcqD79F8almEWqT9MMC+sZXaZwRXdF
7SU0SA8YCOfbCAACh07ERvgfdPxJIxuKR3eEnMYNpUjWXzXisMHpbQFWDBvN2mX0qGMIhGPQYoYf
duD8l0L5R18xvBrmJnpRvMJSI4HHR24TJS6gGtoBCrr8YuNGSdvkxo2PftngN6lpW3SZ0NNCJFLO
RD8UBbM/oeovrC8F+M+mpCVOEweMOdEzp+JCkUkmljrGIQeuNpB9qmu6T0Zm+2N+9t79f1d98de+
8PDs6XnG65PNPDG3gk91TfmAzua7DEk5n64PmmwmLcHFP+7yOWMPkBS8KNwwQSI91C6o5CyeLSei
ls2kbEdOrbnEOUIg1K/3WXQvMQ1RnjZZV/KZMszI+HynDmjbdpFdRJMnLhYQ3SxpWlnOggNR8z0l
aQDQ0OZFlFYvR0wIUouDJa9AeeahPHqcSynyyjvFmOfG5CNfm4rNtMqbRP1m5A4zsKQh7xGT9FAf
Gy+iAVLB0Xgk9mR4sn2Z9GjrJf+TwF6Nn2TiuyXz+lvCT7COOTM85WjfJNCTG2bqbjhFlk8ZKASb
Ih38coVBtVjKNCSufB2uiQjMZFbrvblq9H7dRj6lSeQ2zVFeYRdSou0tVsuFNrmAeLAx2YftPfBm
tkOsCpxZeAzUNCcmva1M8m94VEgFu34qp6N1NvKFkHA3/MGRie+ZSOnN14Uxa64ZRunCuFHJ5LXS
nnHxH6GvXZ5OQQU5eZozQUsTur5deyKiPBO2FZRX3jjOD5UV5OR1z4SoZO0+xAV8jnSHjTzXCpiv
huYe/+EWj5f3tv+vydAG0xgP9flZev9FP/E4CqPt+oZQFHHIdAy5ZuEMNIb/CxTUz6uDNZMSFRji
xm0DrR8pv3aZLYNxMGlCcBwAA+LKWSaTOctJ9nNZQoZE6iiOG/8MbPb7FW5q7Zw+N0QexaOR9v5Y
HvOfsr6JU/PnNDO+vM5hk19Loy02wB28derGHHiVZfkmbD893etJVe/R+7U+8jREh27xKMHjvn8R
ZwoxfL9xXMDnBY1cG5rE07TC38y/+CIAPN94UBKXnc7WEfDEX6wizFdhtE1xkZjfc2i6axlarSlj
c6gWSAZCpG7uLIfuiyy4ggExAmpJtOBeexnS/IdM1+ruwLP8TjxOAQBEhLMMsmYh+kj1Klc01sd9
Q/q+ycQN
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity i2sControllerFifo is
port(
  Data :  in std_logic_vector(31 downto 0);
  WrClk :  in std_logic;
  RdClk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Almost_Empty :  out std_logic;
  Q :  out std_logic_vector(31 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end i2sControllerFifo;
architecture beh of i2sControllerFifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo.i2sControllerFifo\
port(
  RdClk: in std_logic;
  WrClk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  RdEn: in std_logic;
  WrEn: in std_logic;
  Data : in std_logic_vector(31 downto 0);
  Empty: out std_logic;
  Almost_Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_inst: \~fifo.i2sControllerFifo\
port map(
  RdClk => RdClk,
  WrClk => WrClk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  RdEn => RdEn,
  WrEn => WrEn,
  Data(31 downto 0) => Data(31 downto 0),
  Empty => NN,
  Almost_Empty => Almost_Empty,
  Full => NN_0,
  Q(31 downto 0) => Q(31 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Wed Feb 14 11:08:35 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPADDSUB/data/FP_Add_Sub.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPADDSUB/data/FP_Add_Sub_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
DewvQp5Ob2uTdfrB9FOeXk/wbKgam1KBVW92wAknAIeznHFCxwtz2hYwQPnoDphgxe7N+TivyLSw
nEekWVB8eM6o//t86plGlpnLV999UJ2qzXolsjX8qAeowBBAfAEc2k9XCFW/Zxg0vjXEcuM8/RuH
59XJu9Rq40YoFHBMiRwO6Cju/O7FwMvzFbktsA/g/ecKh5Q57xneZB018UaIU5kyxmssTkBqQF7f
IGKA5DRNhuFZNOtVGUJidLB70JNke3WpXix26cvvi4ryuH+unqYMPxdwSiM2L8UrYh52yzUnWaX1
k6COu2oYDPAyaQQy6qPca1NFZcqIHn5qddNyZg==

`protect encoding=(enctype="base64", line_length=76, bytes=272128)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
ssrXoKvHaJcGONJmtBizgLcz3fFlyS8/b+BPsut57MDE7mQwQ4t+MBIe3NGtDZAF16YJJ6O7bMhw
hRUN7gRWJlODQljaK10NZao3p9h5NxWJ031iSKofSYEcA3KzQsw9xFkBBj2tFqEwP1rsQuC0qYnK
/0wng6denFExtdSlpbFey5wnjpJjky0jvImcvnfQMj8p7IbfSKSUQ4VVHK6KauIsyQB7GxslruHv
+7YxVvnYfOYc7XhplzgEO9wj8KVGbdPaRS7ZrIWXC0a/lnT7m+MNdbdZd2V42ptOxh8l9wqPS70T
eaVGxvh0E3/Ntc37HdNyi30Ik8mTkzUvwpWZ/pZwCtPIhb94lreHeh9jRZGL8TSswwTbKcH4f9Cw
R2QBf9nf2EuNjITQBtikVoYNBWyMASFdLDE6VHY6K6cCo0d5ea6X/HL0Z+jEyxI4+6Hlatz7YemV
OsPZnv244KH1WolYW7OW43HmsyfkCPckz6giF5ovVneNYiKt3DIa0Z+sumi5MpGjD7gDQkLGZvL2
3A7VtF26eHeNIyaVv04UoIwsz3T/+tsbjM00j28EFlxco7Nw/fFsv0opKVB9KpYOkK/SQcCM+1c9
u94niaOQIFAPr6D2NsEJlZN9TLUPM+5y5B3+QN+fzI3cVDMuQJ9/78/UDSgoy3yRSrwnu3XrEQ4C
Le7yN9R+CQLjNbs7pVRVL7LTLgDTx8blSUO3Dz1Q2cJJw6luUfc/x/QufO22GqWfbvFWC6vxuQRO
NLwSfeePzlfvvt+Vh6Bc0uj1jb8SXhs4cyR89l8nWnu9CDY2k3ZMSBqdD/YkNF8VezsVtT/7fhQe
JRsx6j2GAKqwmRBmSjknbemVtjDNOQ6302fMHmQ9LytxFFXfn1f/+Imp5ulK2csy5jgivZPQgved
3zehutI5zqiKhSfHqOT2hFmcHWzYRSVrveTo0ecE/GRNFv030fX+FIIsoy/j2ulZAeFMGmM9IYTz
g1sZMem9/bbdAoCLMMPgzkfh161q2HVR+Xyum+LoT67vS+C1F1nANpfNPn7vMwG9ezTWzMf6Sqgw
XPEFiQvo32Od1/BN5Wyn0Vmik9/vD4KgUUaS/unobsrN9j7tOdfcNm3sTvdC15m1Tiqs8qI8gCaW
5KP3TFmjCBad+tSnkCM6bOkqGnkM1j1xuSCMdXhXxhuNeVZ2cAna4NL+SI1Z9MrSdgZR2BF+VihX
32WIUdvFZAQ4aeSqe90Xkj2JNOjLK26vMe/8HswbxFCqS7JY4DWLhfNYo+e5eyAuR3UAGQy/9psE
kBIm1+FG9GYqh6RHdLJWg5aTckE8C2NhBvbXMq1Maj8+BWLpyc5dbm9hQY7zsYDyrSLGVMIOt/co
Of6MiEVGl2w1Hymi4YJfMqqBnyWN4QmzcYRDm0tqcRlYgBzW1/X1krUYEj0vnJj6W2yM66/lsWqn
s/jkpPxdWhvQQyIdhbyHU90C1WVtic0yiM85SQud6NVqJLyjE/BKhB2kFrNrtef5IQKso0lCeWkY
AHTgYa8uede8TkbVj65f61U696h8atA7cEIcgrr+iEcSysMZUEeXUJ09ybwOSBxOvvgZDdbpjitf
8UtSZRBIoIAICC9PsDPFHPF6dd0wgbES5Z/w8N2F3h769J6rZjLlvkGnxhNAQTCgGecExY3/8+5k
+WSE7THFPx8ZwbZOVIm1NUtb34ArEEqeA0gLZoKKGWS5I+wfRYxqFQEGEj2jggt+oU81Gak4ZZJ/
q3J35oDKUmTjFKh4SHvXN3hdNwTdyVw19AnlKes4R9OC6WTwf21dvn045tBp7bo8Nq6CFnV00IRj
RT4VhQcVRXjnF2JGr08MwoCROdKhop8tTU8Q6jxKnyQGxXJyippIbqjWyLBdNlNTA/QXSWZ5xh1X
XA07cWA21sV46QcYQ67PZFzNcID4tLRIjDaZ3daJPds2sg1BxTZGvH9M5Eoz1DxNCShVriciFHDv
7XL7cXuSaBLyAsv8OgfItC4UzEWnw2/UZSim8robQF6ra6jjDgi/t+0AcisuYX6vQF+i5ZU28GrD
odls3pk1BZ9EWu0nOYU2ATRJp0HKmVHfKF/MrLyJRg/SUvIvM0H8GHy/G1kvtbXHzPSMqfR5HAyR
dtg8rCIxGyIv20q/V6dlDAhWoZ/pI6j3WT7/qKESUYP8Jx8ntLEWfXjCG5IrNrB06omN+ZyaaKzP
KUQHPbMH+44fbef4rTRz9ZgML8mmvwMRl4uoWq6tA60n7bl2kbHat1M8+oAmnUWEUbz6n9/ZDEhP
Ir4Fp1mbyksCG6Ntmyn8+fOD9PJBouJ4SWa45Xtbpn8pLj8r59QzPmBteadIrQ1/oF3eUqTd24Gq
oarf/bH9wCSy0opxptt02ov5ElfEUMAdjTln/ir323621Dvh3e1IxSDTdvsFwfTUmV/ZOg8GwIjx
m8wVRDNR5Tnte/pahIT8Gve4GqbAEwe+1Dl4pnrwGokllKTd86xG4vOOFBCyvKEhkXYgoXPpZs6A
cIZO7xmoRje/OI/unvRWVCp6jy0iQAPwhf3w/D3ch+59OTP5FcqwzKc8PFeh5cXBbmmcmdRPauFO
0k8d76bS7ohz+sZba8zriboKlMEXShBokcJQkyUXXAVVQY/e8fSofbnPRooFu9zyzN95Oe5e9+Mf
QZ2KPEIrlb6fLpKMjMP5cI75lsb3x6QB6gcbRXHkWonsJstbEStb8GoAuJnznjj8kzpW/N6qIZlg
KrFb/Hm3H8gFhFxOhaG4LPPai7VhhEd5eg8pHdnNG+XqrhbPAbFjY1aO4VJ/+2hlkIHO9HMjt9/V
93Wdl1izdi6HDoPMEHlMhAS13/ZBBMhCQqayEju0UuXTu8/rWjF7jSpKv17FgsYVuwtc9OzXDdCD
Ku8St1IUV51mpIn1yGctzq+Z4muKNpA4+9bSyfi5ltQph8V+om2UXQt+4wJe2VWe8vHNQ4sFvt4s
jAeZYPUmNCV6eO5/5ysZw0DrA7rsrF0fBy4YJaIijdCIsI1sWpNyqfmO+TdIfranfBRsAxHjlj5g
KTj0jj0zHVOMeLuNb5h8Hoj1VudpPc7j0Q4GAeUB1g6V5bjub1tVTpF+7Wp+Hhn+HGxv/ERdwAP1
8/zvj1r1jEEsKr5oCMafn3m4TD7s6h+0Wi5Z9tPY/sL8lcAsFfNmGQlzIhSmLLHtTGlKLwleCPxB
Vvpb/Sb4Fpyw7Pau0cXOK3LvdEzShTeuKkoWZaWCqXnQk/aM0dbWdGUArPIZ4kXEb586MO9WuR3p
RhDh0DYac1rZpgaSuEq+Vk/oo20FVtTf0hCoAjHcOcLnv1LfuM7ybEoo8nU+orS+N81em8U0UfUv
Xi613Xda12BduGyZSqksa2oSlB5q/4nnunPZGyMJ2mr7IwRtgm8rbP5eR3VJ9cEBSIcK9d+l8QJS
jjic/K8pnZLIEMkiZl/o4m+4WP2mFWti4ZVMMHA2TP/MhbpPDpKz/32y89CY6lrBZ2dvEGt+BzoE
dLCiX1jwiQBQr94gapMtHzaM6At6E3qVija8OM0Bk4AIPGWY8SOqfntsLEGJdbeHYcpfrAXkja5x
Ry4tfh+GwvnaJgybJEun7hGMopKTSNJyw3+NYtqXn9WYjzRk9lTxQCRLDolCtZ7EgPc1Yi8IbMP6
BCH//q/KhQUpvQ7lutxqLT7C3o4yT0IZbUhLtNGQrWLozyVE/eaDZzn4ZNCqnH2YOhikH1M+OpPl
IxcasZj94R4jwUEYVKvEyfMQ5h3Q18pCJy/vT6wXiQmypJTbZDvANRW+sSQOfhWqUb59c4f4a5yR
dCbb0+msM+gZ+LFdlpzYtRSDFLd+D0IlwzQw31YqDl4usA996VRcrrCID3my1LL0l7rgKpoegg3e
EPBgJC6PNGwtbfK3PDfLBSgu0OJtVhlPYu9CWNyo16THsAQfa5xBgVxLblUhmVkOHMuSG/4cU2vs
gh4JhjRpvm2uaNU8YnIORbnejhTxrstNcJwHi18DTjwwpYC/OihSYguRFgl4o+2g2aMMsjyM5vE+
IsRErVXh14VLvBR84HxUYYc3x4VERgB3IbjK8JiDlycn08fnd6fMvooRLP/KsdzQvQqEKB+KyeaF
hcUV2s3nf8U6ZZPJFlgeaMzIqT0bbSAst6fV6SKN8PVJvF+aj8+ULpKcAQVtB8OKr/y8lZYpge94
qkF7qY0Nk0zMESAztgFrzjqvh37lP+OhtELQJF57IqqdxBtfCjSaoj8OGLfar977L/Dhnoi1Kaou
PalvYIvuebqwD7iLBRLayCKXYYhRWk+MYWBOfpbvQRyeJNBhuaushePlYNFQEuHHKNnV8TKdDYdT
WNyuywEhOWk68+UDDibY/HXcVt1ANjUTxH1Z7sZiAYCos19I30UlX4v8GU18zkuFEYuqLutlFaqY
N/VzdS8EYDvBgSxBT9HNf8mWOnWZ0B9hhaM57syKUBvIo3fMcsdzhLqBJmeLcHpwq1JL5BxAcXWi
/UQ+KTcxUjGLOgQ554+wppszrrueX8TGBBRY25u7xFO+D6utQUK1vPHVGpNVudwME0dXqekaO5+e
1NXv885RqO4MB4V2uRJ/nr0GnyTUvAwG8GU0m+I3BchqrF9W7hmdGIH4HtOGAhDfV9HjAu4KHbyh
owt4RK5ppbqs7tayV3amC8yVNMSaBANP23ayMM8FSxinvE7+zs4SK04/3MYXtD+0P88yJbCdXghQ
4r+qYSuaAYQbTzbSEPxhVdGwnUMEnNyLBVhWZz/HZyPY+g+zNgDh8pHRBxbG0oHE1EkK9MOh7TWM
zq7XZKVlZk0yJKEPTNw+USj6QiZrWSYKiwweddVElYwYKjDjwTNW9oUkzfTOMkt/NjI2GZ1hc5pQ
iG3ulyQ3jmmVGe5aEl78AwzOdU5fkhshEF5GsJ8BOxY4DVSMwz3dP7aZ6UbJdH5SD4HhDcsYgkkY
iGCqaEOgR+jLRFwK6H59gfGdxsNpJWt/87VmVNPimPimvCvbyqfIG3pMNwEr8hdpHiksJWTSN1XS
ONb6A5NOhg0TcV/+6dHQq9thqwK1TdrV5w5HYK3EVzWc/yLGtSXY5L5/b+m5g72RM5eVFDeVbhmo
5T+YUON4MgP039bL/Fae3wMXufU3X/Qu8VDSz/ScTsdvXfQsBMhDbb0K2tSon88VkWpdjfKDqbcF
ethIYPNxU/+4z3nPOgOMMH+dCAHZ8uJbA9jyomijYP+Mm+01E5A3LCJyOSWzqaTGZBMwOCk1gW9l
vI6nkXvjaFcd/SynjbxlzpWv/g/V0/TDVcbBZ0tKziLWhdw+EHF4my87WZtYJKQBfqVFD6boAhbn
HNVRqgTBxqzPUXl4FC6YN+wR93SKoI7FuIr6sjJAewLR1MFvGCQfZUttjtBfJgz8wcTKmSeGkKa6
F9L9/V31ZG1e9Niddkd8m29SLvjPrwCPFv+0iHvwU3woqRe250a0bgpgruM88AIBdV9NKXqDmAMg
B2Dm0ov2fhiKxtbWdHrYXv4sJI96vRdCP12L/YHskzhMaoj0iKXm0byWC7DlwKnCwZjNohaTq4rG
IfMr8DWttTrls+ZA297GBV72dnA42B38OvulBIiDhlPI8cNPBfbxUCaN4hiQBd4A2NxW/5PyCP2/
78CInofxeswgN3o8LcnNKgqto1omqZahr+OFAn3xv75XQ9WfqQRbiQ5GvbIyv0a4CWbuo506suDD
CHNl8COGgnuORS6q3hIfZgi1gONscqWRE6/LcOWJwtAfP0Tcg8LCJmnJOFQCrJYwNRr7LnQ+r55N
Mj6fi7OO1JICJ1yrLQwin9ALUrtY6CSN1BL6d65TodB/PtCrxmm6iscGSR5tYEzhHu82alp0UgGL
XEveQwytp8GSJ523+E1fXh4cSDB7JCY790JijxY/m1NWRNXDfzk45cuzTQMZloZFB4imp/lg2sIz
iBnri7Fy9aeAx2JItdr7A8lyG+R6PU5+RFQd3IAlVcK6ZJFJvtbvT4VUJ13u8a+TqXTYj6tzQ3hY
LgRJUYg+V1tBXaMNg/13paCJ0ccSGmzFBCqLHZ2RIFoUiXXUwG3+C7JZw7asyRbSsB+Yc0wLs9Iv
6Rh4+xtx22Xr8x0i+3zcZesLBHL69bljjoVLn9TEmKH1r245mU6W4Gq0QCY/IVK62hBDQlz+RXeU
+8szcAkVr2b352UtRwm5DxYZ1sio/mAcDOSXF2l3YS7GYanM7aShzOwQ7YnDD0Yvzrt+FKmO0lmn
+mjRoSztUkYofuIO3PuhdTm4jIvVJYBLKKrrh6rNGUwlS1S7vrmS9MHBHuIhiqUPzBV+a8zXoh4s
kdytGcPu2fdi5GcfwCpugGHqtaUgWnze66WGwydj15HgVfDohFcRn0ZMasJR99RI6q4v9RFaiykz
324W6cJJQyklbyK91m8gPEXRzh2KnriKi/BJhBWpKZ6/kB++Y26Qc7DYROuCTDyi8nwHQktgO5P/
bhoUL8vFnTxTDu4VWdwltmbSQQav7c2c6c3jasD5f5jkVHT2IxZqDzry4MtkyZ6NJKyY0APgz0Lp
nATUU19bqVPJTmoAaa9e/fT+mXana42p/dEmczVz81T5rz6ffW6UnmaqgIb51lMdD21BmMjOepIS
/MlfCLF6U9G+9dTtILTf3fCzRYVhIhdYEFdM7ecfPfecmK8C7FzTumIYbNeWph01m8vZlHY+JtbL
8VptJCa9C5X7wnCaVXQDPC8kzh+x6kqmkdz/Cj3FVsAEhPVN4pJ+UX9eVheiya0OquBoG4erE4Xp
G7aLeFa3uWyrOgCQottp+qRCQnqurzJ7b1ExQ4i2sWsZrk3OfjdhPyxPjnCoPvHPBkjLn2pTDQ8n
YN1yYlGqeIetQJuP/x0q+LIWsry8DYalSB5Xuig+mNnIvErIPVfp+rnRYNGZnvXa1/GbQwi9HyIV
e8VeJdeI9XGy55T8ABFy5tZLemAFUlRScr6UCt3JtElzTrPJ+HxHUaA0oWNFZwTIyXpTXJo7mFUe
7gq1ZSwysti149B3u5zQIEbhCwhi0aNJPLMr0257lVXz2QofjjZBkNY/ftsN3Sx2+2F4rMZMBdD9
ZhOqrjSGcaQUrG1SieCua9rTHrKqVx16rs4a5ZumrCR7T+3Y9NW0ykxICHI22M1xDO1zVOeIkXVt
/Rrx0bQXGuVEKZiw9IS9a9aSVNwUC/aGqvgDhKd0hoxwG6sKwj41MQFYUdlC6gFusNwmkJaUN5qT
rYZ2JsX3FDMW2FXqy8mYvA7BC3VmVVnZrT5XosCYeiokODo3fzbmuGooFSJYb1ewmsND+aMYUX5J
C7n8auVFHrIZZGrVF1ZwK5aijpXqZ7qqNL9q+a4vCXP1bc4XEgJag/7YP8V2Nxylepdo5K15QPpD
bnp4RTFyNN6TcL2M7LxLrx6Bn1thYb3z4Jks/6I0CWLATTRResVKUFbBG59rI+eyY9OF21HM/V8l
6Rb8HColcE7KIwPC6T083JhMMyM+F7jyyb4jzhB5qGz5K+udioYYXbYgfeikv9KbHVuwimZI6qhY
XJsdgKlPsfXfvcFkTLCg/per67SfZwa8TrXYghr0YF0/peQOzeq0QRjJx5mXhEJsUeJMWP+a0e7+
bHBmPoFD+VSoJXQmq2XBEkYbSkHyzVIJuKK76v8RH9QCZcCZJNP0VFUqSOzL7kbpQ9/bdQZnbbrl
zXluzek19t+ZhcdekNKZ2sU1TgwInMNGwd1+7k9quJ2EFjs0thWu5/GD9Tc7IfNGpk1TCs/udFCs
OX4THeIGLpMrNNv1d0fylSkE2UIRUlC1oMbBlxk0kcMO50vv7YeTVtep43Gdx+lZEKE+SLDQt87Z
cwhMQmwXDlvIT4NLSysOgSIfbR6YimvCdQ3zOKGSzhl7xc+Bult6IJO9BwNjXqueLFY9vXUkKiX+
FbE4YwZ1d7dIEFMsKxMiHdyCu7En/VCFQ/lavPYiKPTJBMP4h8ucgVbfGo1k13NcUqEpX7OhMb1C
QH1h60tvPl3N4zxquT/TR0gzFijrRZf6FDw0c9/SKUr9YTUh4UxKBLsHMIjUzgHjC2klK9ro9850
kz0fjb7zhG17TkpaiNCzeHgXqz5PuTPRwgd5AOlpgK2iUm06v7QboH0nNqGYyQt0xExmOz1H+Jcr
yZV27FF+urFA4SdP3uqhZSq6IkLFzLzZBtKBZO7W4nGwrzJbiW/+KSQ45nBysIjWPUprs4XHjOHF
mBDmDkL6cVrrYEjv3p5gTuqYjyyLToW1vP0bWVf2tD6/U1gf7yLWG8VpeasNreKahSbUI2uUTbAV
npcu/izrTMNKGkowfyFR5Cjob10cWYIdrTUSvLyl97+XR1aw6nGYBaNnEpYwJzHXZg9QyaQG+Ax9
IvAj+k0VrAhGHikdpT9bLIe+v4Ayp1a9EJJc6ry/z0KtlrhUN4z076pDEvMV3xmNdNsSbRL8xtrE
wX2gqZwHMx6K/c2hVMD0+VZKJy8lWGLs1//2IOceAGB/k/Bm0SfSpnLIW23WTsu/gB4b3ejvSXBF
FCzkyXYfpLZ2ly/wVPVjTKCqrc4quvRahAih4E6hLgxj/G7qOSMyXyzB2VTWRPI2tMm4HF2fnRHR
Ctj7UXqLiVAdo4yrOfQRHCkLPbUwhH14azAO1Kq/UahdxBCFnHjN/VkgqOYgY6MUfLxca5Aom+vJ
xXezv0LZU10Qb3Qe697WDQYPBaSRwcKLR0y3oS9yhph1qeYqrcmjvSl+eVUcB/G7EJAQq7dIICDQ
N1empSFPPXYwGrl118Qpi6hz6S6zBmcLj289tASGpddhRhkHx+9XNjUp3XUZ6QPsdgEN1N7dABqN
BwC44/fQiqVwby5CrsIRQ9m3ZpjgOlnwGLcJYV+ggBVk8DtV3bRKQqcA3Jw51l860dGa3FqBxJfh
arHnfrbICDj7Q42V5fd1bShYg8tdzmH8mN9aAeo4qpgRwROfRwg41keMESZDTX0brt3c2vIyfJXY
iKO1jGO7qtdwez5fCDfh1J5gnNvqS7UuHi6jHuqh7Nuxoka2qKnyIWf4BY3VER4SQGjNGVqlyVcA
kN2SH4bPTkIKyGsQthUC7GBEaj7D9sd5MAPQ+I0FHnwg7pkIJVUFUc61fnm3de0vd0GsIwh3AiYu
xS7vh21II7bztJUnnQVnhaKTaJ+AZ//okz9V2yruRn8RMXd4I+iQxSMNE/RIppuXwtmg6/UjKos2
dlcXCP8Q03I6hIWgJ/uSGFrmTcdsRjOsuu/u8RsoTOpzeo0Fjrs+Yz86f4X8Iba/BxFc1a/+WIuO
Xfiy3KBeJyryK9XapGoEyRDoNFpCtilX+0wKSH5IyjNwPJVIVSgsm0HWKuL8UO6eeA9paVM8XxJU
ElN1nH2s/hIlMaHfAl9aYEMVWhUx1ZTwuGOf/pXzpgPfi9qdn3gztEkOCuq3u1N+BidlKFBunqoc
kYMsLQ3afLioAP9IEKEMrLW2FWLPYhqmF5GNhx3HR8+ZtiXOK5NCYNw2EdnF6B47QjMN2eIsDiVk
dZUvyOph00vvgcySgRjh0LPMsZhIodDcTYCogYr3D0s9BK5Cjldeiy6Z+R2DdSvZ/4bWd4U0/Obv
Gluw2pwm+fqHihPLERe+6rXmp94XLGh4PgiCBhjzvYlZlOb+wtL3W1Hhu29dMNI0pGTQ/yqnJsn3
9anp2fr2qIDrwRsjqTb64eSXcl/6fwutqnlHaIFtpH5u/qPOcQHaRCMOqtrdqIFY9c5uYcwvVu8z
Hp+d0Tb2NzF+UcNh5k0d2BqX9ZOLzedKTCbwHekn6ZjEBcbRjAtV8NvSAjpTUL5PVyMKp5clmRd1
AbxqfQ+8J0zyB0jcf9euO8al2qWqPflxW4THCEaJjV6Ak5ErZbCOwYmevnTCa/jwfUDYINirY23Z
5YGeajpF/U10g2KCyrubZdeWIvaag6sDxjBDCGXv3VOpvsSoDWg4RApZ0lRtg7zUn4R4frS7JRiy
1/RaQiVendBOdjzjFN7ZQ90ggQkZLrvS2mIz2PeSbueX+O2hqNkDELOfx8UTwrH253VnXjXmLCUC
N3W06sDMckRm/hOXYPrZXopNejfL37xx0VIGmN/DMd8pt4Jv2jlNrXppLY5JAm0geYCmLw40c+Aa
YmQ5wPjRHV8LZbU6kVxPdJdu0LUJG3isEnENHCp5uKZAA0e5jwQJAysdFcYqGMc9v6S+4iKgKLEq
KAR+s42f2qTCItxdfo6wfGPWSsPcIL6/X75gK2UQ+Ks2pMzC3GXc/nbJavgRANDSKea5VFGhRKRK
mkBg2eXM3V9qZCEIHTuz6ySXkR+KfuswWfovwhRopfMScA4a+Tfvlkzr4gadKfKXIQyjQRqWVZ1I
zMrweM0pirwdfR37BFKOig5MAUdIrnbRCBM5ek2jZ2pizS1fe2ZVFOfbOG3hGmJ7C++yL+Ksjo2s
aIzwHCGvgCr081Uuq3Iod0OcI3P3cySFrPWfIaG2gPFZpyEB01Obfi2q1rZLhvKqvviZLwmROWY0
kR/zd+PI454vxuxYXG6YzoMVZjVsbelaYlI9AUuNsn9Bml7VCXFaShXqvC5iYJdijfYhIrUbWiDz
0n8D9YvjJJxbrBGnB0KOzG5PA9r/2oFCRVaNCYJCqT6w0/fVmHSna+mQO7mkMwM6ue8X9AYITJQY
3ye54vG/fyJNByC7hxOdeLXQxRIvff5tg8qlbyCDfsKKBQ1lyPyYkRgnMDRuaL1SAIZ2kzkwwwQm
7ljZMhbLmdl+4hY3ZHtxl9UHVVNNYNg0GKfP+ojZptp4EK6qw15SqJebzNLm7Jsdcw289uRWLdOk
3D7JLOOxa/9LZSXWAkaieNnjlN94IbEmqUaUk4yR+vtAFBQuP02oI0bxclDc0Y6KQcZeiGrD+Q9b
BniJCGURYdeJb2Qd6oi2mYP9RLyVIJtFylGpaxyJHiGed3EWSq0UV3aBr/bMjf4+nRkFN9U6xYT/
abYDh+5BU+y3JloZ3x6L83+iYfDhzfCSMrYml0pD2IkVAgeVFLOM9E0rvnKy63avTOPsNFP7i7Rm
+nYhDf7ZGJYIqBSwRZRba0l1PWdLe/96/2yX+ji3npqjChu8bXHwQvk+o4eR8a+yNuTwB1Jws6QU
C1wcX3FjrbLaA+yTK0TN+1T2T3eAji+P61zviIVreMkRd5UfwoQVic5EKRXKCrwVWviium7tvQmB
6SDiLF73nKvfGEbmifUwMCTxFttY89//lwIMGwSvvzy7EtgIQ5rPPKJlaqykGsuJE64xGWOyUx5r
M1AyjC7AVyy3VS9PvsIdDaf0ICM9LqXhfrMHF4x7Sng5aUyQtYCDwJaWD/o2QwEQkLetyRnoFN8E
V7ARM0W+1QGDMOJYYPznSubCEgyLGUIPkMmDDJAyXxlIKyoD0Ig/8DDRjxhuAIoZJjsXD1s4GclQ
FqMXsfSzRgc70JxLj5aLLbb1s1bWNpTkqME1rjxbs4+qCWIR4fs7eLufkCiiaKObnK3HiODXPh1u
inFQk3zod75wPtBjGmXt3NX2uujoynJ1w9bxk+6ybNcqR9i/M3/R/vgRrULN8dQnlS2NcfqVAUYa
phY+t9jMODW3NCAy3AeicRvTEAVa1Prpg8IybpAiDnenv7QLMxPDs0IfB6573sh0xv/jXGWEnZuf
6Nlwyy6eD/HB2DoukuhCfDzgq+dboFwAvpVzz+9q38aGD9ZH5+++uk1WDk/BmHjsxoC/13VMuN1/
skYT4rxLmn3ufY725uapONri7uK+GL49KObe/TN0n0ViwJ1QiS7CutjV9RUrWCsYmGUHzhzKSJVE
hepj/UX6bKJ8T9Ufu7cZ/kca66DWNeau4tESTWdshPrsBPZxuv0TjdBUpUseMNw/z+O9Y0uZ58wT
t9ChL5nXhgdtUJFED6IzGcUFE30q8id28tPRoAdmSLZoY1nVmlM/8uzl3PBOogJXx05QL3tc9qAS
IR6w0lLHb+3VOqg5N4VpFXduJY9wmo+jr618oinlr1nJ8Xdh5c9onIKiCpAoS/iUrkL8ctNSY4EA
fyjzf5h8UG9cNidMklNBSkHHH2Xd7x5edIi84aA9zSg7ZNW+fvlj8704DLXp/mRJqmehsNn/pig2
AZFtPmkq5N5+q5T3ay8GpJzRn7q9msR6AQrUcloNtQk7VNl0WypUg5f3/GGqGKX4+oJT9E1izisl
IuPJH8oPC4z1zqBVQz5cKBNw2+GIfcTP3vqZWBX2+xCkMXR8z1/llGtg6Guz8vsVydwGhJVOPf7v
rEviMcojnvX0g9wvOnKPKpWF0HoRwamwjjVDY4JK7mIRvNNmynXlPA3WBbCHDef3yP+k5+Jw3EaA
YqGqdJNUccuMjLkeGFVQe+iYGo9T35+ZKuILrKsg5JJwYskGwRdqzDSvTUnTqIaHZV2y/ZRgxpbR
uJb4j7ZT5h2mZL0djCw3tJIkUOJFpTICgJsJr4gZ/a2gPvd9pv+lRHw3mxDZ/c2vpKzk3ijdYkgV
nBwCmHGvH+KbAmjDMv2aUvtdRCIWmcSoGgAuDJXKInATzDgki+XjtSFuEJ1bvsq2PXxwzz3wBIA3
mUjyDA7/n71oZtaV2s+kzWIr73xzspPdq+SVZ97SV+kyG9JuTrHK9Ih+1HcBlPh3W+FuFjcL6kSY
6LSwirg6nl5gKh7zHbhqwgt6CeDfcFoaVO1bHwFFsWaruWSFXSWQFkaW9A+9crQtDW1b9Fxi+rsJ
/5H/RLRMofVZ4lp3oT2L2pnJyisyy24u5xGDMg99wfIkHjAPrqHS68mfwRNFuQl0l7h7xJdTJH10
2Tz2BTYzjK5ZeDWG3FT+D0a3PG+zOMl+ymu+eU0UoFzoC5N+DzQrIfo27riOAizyI58BPlSbeX1T
lQXdMvUvJuML3oy1Ncsu/mHR0y+RHPkpVAtyHC/wZw0Aqpbjbv0jyNzbJE7OBKC3+fCdmRQigOBn
Z1vW8/FjPOfQzNyfrK6QfbCGJXO3EhbrlpKQT05E9o+PlhwWWq5GkODHHOcGvGUu2UegPGvVtO/o
PmcJQBleU+ptfOmMPCgVS+ToLtiBupeWSF/VcHcBK8NnxX0G2iA+PbB+vXYXmcqBFCS6TjacRubL
J9RpalvN9RblCe74r9beBwnSq3roi7WYrVnlWMnHYAbuFBQ/IBg1uREBTC2qbt9GHg/AkiAG/FeD
pcZrn1KMKnxgsu9IJSW41y5gk9Wpf+AGnvurUCc3EcBGd903Lb7Vplozd+beJN3vOAIl+2mvJHia
4jXK+QeYp+6JxB7JeMIhA9/VlV8Ky0nFWWt5UAHpCsRXbLWR+I6mOVUphlhf9QzierO1r4tOu+oW
HsA4ukTRZe9SgU2V3H5jG1LlJ9RZ/WgOWWkDmECM1ammssOxNcdd9MyZrTEus8sXMrG+8s7G5T2n
Pcis63CL+9Q9rcE+uQPxQddxP1Fk3akrDaL1gAgdAwDbEFYBRcnGLJx8HZHHT/pVytIOBtORjfQR
Hr6XW0xYTRkbf/QVc1fet6zl+I1Xe8tKmrG1yPvcsh27SLsVzrD43XdjyIhTGfI5Roo2w0s3Oopr
mYvls3bj5xdq1y+8//LKpLJO6GdxYGzLl9y5H/XZQXFcoIItEnKw/oHWEUaINlPYLPEpSAkyUhGc
O0Q2flvXmmL9vXcaOtxrJQDqa0NZP3PlMpKmmw52MKdGJDJIc3Dbgs081tUceGgowcDBY3D6sSBC
TY8LVcdogVKRvGGwfGDIDT7Ev9FP732xF6swMIJYDqXwcn0NNVcfWyWwGd1SJikEQkxmiBtptWMa
BMkAT8fcCAlcxRjIKHNkTtjFR0MJ+ojGgImTtoQGWYcJKsnEM1aS88gSBR2WTUD+Z2MlWbDtgtfM
SonK9OMB/EhL2HtJc0eYgaGvHwcgoQoMVunj3DFYw3Mde7htWRXa343ZVIuBEtRDTFUWPSkRHtkT
0yUnpTWOmobQ6k3FmXoYO361KxctIVEJ1Y+PyUFiFKAWxl/F4u1juMNJKTNcCLP+LHdMQd6s7zIQ
ItkWUcJTWa5VcuMcJ2xoD9DAdmWq+5Wa21eg6XGiG5STtPNkqKips6PNARU7jwE1UN7j/1gA+cL3
0QFI6m7MtBKZQFj1eaww7i8hYz++1GOkvJ4+qJyUAP14kvZyJ1tabSVNMZNCE7RMeCN7owfEhAjA
nZFZ4aSbLi4FxTiCjwQc5gfYI9O8LLm0xeufJuHnt6QV91cThsdhRt3f7VCWXLotatnDzlGsthn8
fzX2ISUX/UyacatiQo6o7CnFDh22qVPy35ovlH2xAbTKnTRRcvYCojCpdUY3kGXnRa8uc0RZJ01A
qWlJedg+nxncuQeV8GEbedUjTPTNDFyovRUmFUarFTogvZlMx7q+8CIGI+JlUUfCBi8zVfykBh2i
Q0QArjQeGRbWlROxj0l06Ca8pY8OECERet8JbEVGkpFacJLVfu9zeLbit0ikjuM8aN6EAqk9bYui
+WmAuC1joportqxTMzJ9R01WayqbLGfDAG7I3rKX/5XxhGjeBVH0ei3ocwoal7o1hdbpk4GplB43
B2gYDHigtWxhUcX2bcuImSlfNWcUncL7XAQhHm7VFVgBESmJ3ZmOfvLvHEeaa5ib6ehZEqFWh9Ix
1KwCXaw2ZO+p2ZEUHp952Qi+DIlEn/dctzW3IHGtEJjBC/x6BTCt7icIsgsOy/w6aYfssiNZlDS6
XEV6THGVgYCLG/ZYN4QxZcDDXCkcFSzPZ+cd3d+XSOYB4/xeBRdkps47Ccj2e/w/vaXE4SK99O7Q
ruzjV6wY3iQdn8ErK8osg2vPAGGc/ZyshV5cA6vz6fmxNE++LUqUeLdlcdx2z2ACBQEcVzT045HA
gMG1gf9NhdleDRo0bVfyv3mwohHbIP8n5omeKwy9142w3TzhkVQ+afEExk5ZyETx6pW19nYNrTpN
4rVHzkBjVuh28LI6GfAxXfor4VexEUTRlrYPyZoiq88vwH0xKuTSZ6f+gvWSYX9I0cq6fDSpLtoM
e306p9U79bufVv++w+jPjZgbd7PKiTuyErsrbms79s4mPh1YxDIbjuszXB04KzSZshw+gvIqYpjb
hOQ+AbBjOjZ+wonJUqkQwSAzgRihrB1osU5sbcAcMpj4pieAV+VUfthpSFgSDpAfED8L5hEDp9cx
AZqXIzzKSQ9s38smMj1cGvjI6m46BfDDNUrcMWjbmhUMwLnLnfEOzKrgGE79T7kmLV7HOk7rEicP
qqi9Rtj7F+TV8SMBXJ7d+JX4iuGgWpfzdIclv0k5q5iKfK/eHDtwe6ar/19MnnYRn1ywxCBeNtMM
T/oXV3O0PEO63LWOSSZ49mAJyBtSJ1GtZs79hZY6VFm+CR7IKoXVHU7q6wZBvMTdXliBVBcB6HoG
WcVSA4JEqacP//lxPqgvvIwZ+ZCyvEtc3lqk2ZCt7Ol4vmxU6C3qMQUQye0h/CAk4jjYuE2dtvss
qZq6HtX/wprxreGHyEIoF5meAqao60+NqZBoyAXWkxoI+shOuUNYgxXKFQJSrtwUP/JMxT7XAo6b
SOAbH71z1toTTWiqMQnQ9W+2vnlGYAdNLV8ES5nPzKydPN74AEvrPkjvv7Ck/EWlvTHift7DmFWu
jHvJTVUYvStJiBPQh9BPbcG44nqq00QRowvfSRhEiFlkiS1gaYD/6qWsX4r1I1HdYpBhDyrTWA6U
C02gbK9U6FG8o/ggs6lvPkTDR3DUYf/DP+vjz0Mu17ANyiGa4p86IiEZAQE1Tc43BHzDfRiati9z
MxjW0oV/DPpW/KTcaygczEUZ5UK3WgU+QeBS6Ub2UaZrcyfr/9ifDtz/sLgl8kvQraaxO2DswzdQ
Mm+GRfEHbHau4EuhT5dBVMnYk7lp2SdRhpliquB0ennmvlrBlTREo71tF0Vlh6kuA3NPJX1bufGV
2H2xX5fwcJABE+dobd2OmAUcjejGUz7Q4kKw9PWIQgp+OvHAqmOlc+GeroQQ6FUY0C+g4qY5Z5Kh
qQVVScUvtKHZi7jc1qgNCZbjMS0uyHHXLaaU3EXhnNl5hYtni+63o7OrHnyVGpzGQfpbfLuTGX0M
FmrQ1ScwdrpyPRSbGWW04RThMGHdhoCJQ7JxIT5LuaplXF+HraMF7UsodQPyvQD4de8hIZFw3k4Y
2p+kMhxbE4JZ8T8uGscGV38o1cw0c2PAwTyIGEeNd/uFl07iRTqUgdH9ldTmIHdRzjCGUsKXmKm+
qwXNGOJGp/fFfFsASRpkfgB03C/8KcBxV4g8Khy/F9pvAAk52zuYGbU8/HgDTS3BA/svf5yEnJYS
9EdRGcjm2c+1c7ulGZFzJGOisJ7MCZlHjx/pq1S9d5J8LMWBtEnUTCcAEUjolPu0PUy7oof1T+cp
atL4K5sYzb3/cEalEXoqEnbeeBxcMnRmMhw34vkCMsPvOB/433L9QjCxQVexZJO0SuqxBitgLyIs
zwhuH4IpCRlWU+0qBzk/n/tNdJdm/oCjd2mMGZZ3sAiFb9QABZl4o3fvJLTWicpTfE2v/GFbSVSC
FtZemrZeQv6SbNdQn6dmLpfxWpokHAJ3OS+Gnxpr3BbI/iP4g/j30Zg8+7vXjBb8lPgeJ24CdctU
GfnTzlZz4eN1qlveO4SQ5s6ThgrfoKkAU7LH7A0R5hdHMaqgVdEyClPCZExAj/NIXr7ILn2YXwXW
MNz1hsFr7K5wOpqxj8gGOMk6nmlnGOFJW8AtnyDtLUoTvOpIBnKxcqax9tTPzBUDRrvMEX/qXJb7
Qjk/SpcUCwS1yxxnjkqDdSe8bmd+qLW5QokPKBDgqoiOpLkxvYWiOxIu7B3F/19kJ12J3XPxz5C/
TnJBgc4/FyzsrDFR4u6VV2rjVr9LoPGtza0spuCzeRHy48jM0bOIKzaLV0NiOHbwEQjvuhfwgYNy
Lqs3LiZfKHIxJjHxIYjP0T/dAiT6XaEvGnLNWrsAkpkB6tkdJOt1ctDMw26D61EwJU7GOSYZ/UZT
0qPKsvrR9MLUZJwWWkQ9yeLYbVoyBMR7X4dy2KDdwGd4NQLX+vnn635915KI8B7lSPB09n+2H0hh
luihRSWg6bLYPGjxnq8fkEhO5oKRHgdzCqyRluC42hmhxOq5BQ376Qs4b3BdPsps8Kp5JqRVxHyx
UZXJRptiawF+YeTpPzpENIVf2dK8x+XPNUhJOUXFpGxZOhJaL2Ozke2OsFGRGpqwbtLri4KZazrV
+PgLsKGxMkDGa5J2S0wxNDDdC353dMl/LPvrUtiBqbjzUouk0+0YKLY422sskuEfi0zFVqYv3OC9
XDld+IlF4eiSi3yMppRl6Tezjk4upXjfY/jn6s3Q5cJt05C4UoaIOuXzb/xtOo/5+I4okpn8AuiR
u9jXtft4/ZDBM8efcg9JiSBPfeeWi0m5/eHocPAXkyUDMBj3zYnadyGjfWmerB/af7Nv+StFhqeU
rPf9QLUCu3hxc1zetJgTiML9LE1mmxLJZ7pP/IYE5kuyDlQQ6/pnAYNIjonT+8Fe3xl1yxYe35N6
uABzc0W8jSDMaROz8Xe9NNlobeqk2nheWTjzqvTTrkeyMLlB/aTglsuN787E0HM5zPG2/5FVQyvY
fU6xbL0QrpVzvOsUgy2I6JZuQAUmjZykwrDBfMHZ3jPrSMqFbXeNIATCKd8DIPL4PKSC9483LQNR
C0Doyyy/CZpFYcRVbxd52Km+3Cirl/K4uK1HFdF7ipbOFK7I2LQpAWACEuSiiwyuKNpIiRU47sry
UIsP5ypI5n5ihJcKZ4fbuMJH4Hk7saEEmtoNdvMXhYLTu1y7X1CnjhmwPhCnJeXXzRVVNYN+9fbX
WypwXaa1NTxQSN0oa6gJf7BHv1KckH69m+97soZiU5NASJXEdpsFomHg8Iwn8/u163bAaU51oN9I
t+I/Gz43i+GtLsIRx8MJS0pOPFL1+J1aSN7GpYQ1NuGZ9VdktqtQzYqyW4+nQzrtTr0AaymlCWK5
JcAGv1dOBnZdlqEu4PyyGR719LwMhrS4j6tF32HqVvs9LDGAiodawWUzFMAkg5wgRoV24ciOjG5T
g7h8sjY951M4u++y2SSaJFbqxWgS2j3orV8umVXxZkAno2+YvJN8wXVwl6V/7AZBt+n4k7IDs84V
bZ1GXbmBDDZuTzNAO8CDenla+BU5YVu8ghMuSCWAFuu75T+rsnW1Wnryx1WXsObNv65Ys5kzkil7
E119rmi0nU3DVWA033sV58OhyKF9EG++iz36cvqR+vWeTilCPLbBIzHOYIM7v7p4DhZxkpExKQQR
Qq0DVAP3iuMXs8KdeX2sndwffMiDG//6HD0xJ32Q0zM7Z50EjOWguJXhKTAW+fUTYwuwD/TL+iy6
A1gCaw8IWOZ5PW2ha2mz4Q6VEbQjZHWqp1e3cZ0ggE1JoP2MdaMm71FSTcWL1vbciqr8x/PwQ8t6
7MMJF1Klu03OxwS5M8Zpikcu8x4YH2d12mmeBo81BOK4ARHP/8eQ7t67MNcM6QkhPKbLyg1Tde7x
+DAs/eoFN/Lwq8qDyNEpToLk3ZlJh9EB3k2eta+J2S1pLL2VmHB5I4qFvFT27d4BXseLhEbMtRr8
sOA/GqvIbhSbOYaze6TChBN8WPtQYEJ2ObNZhTdUKKz7LvmN9GiUqdLh1rrGMnG0JV2wDnhvJRIj
bNq0WvSZHo+dOWa3dqVgci/BNOtvKLTOaxHaWIg0wM6zRKZCq+pC40uIrEzlf8F8J4tbRgvxoxVn
4mm3oU9pWRtZdEF7MRJdlQW0lN1L66qWJbgQgFtzejc4s9LxexTlqPGDumO34reHiBi7gkdvsSOb
XP+zdEnnrjEpBZc483wBh6gCOkGbo0P4IXZoTEhkdifW6NJRQplzS3mLUwcl7PdcbIcoJ2PhgWd2
Ba4kRQV4zCxPWI8B9XcjqbgzBPD4AyVrH1dIaxMgT1AUvfBDt6tLX1aqqnYFjujdX1JXzDr3Jhm4
5N77n90+QBMxHoTtzaVWj7RpR/LGQxe6K2rr7kOwjxpunH93FkyLfYAr+RRNiEy2g7j/NhjR7yyh
FObnO3O7IMhhLRHwT2kZwr8GEO+S50xLvGmJJRfbBxDbxT6G1XYNzRPW1DPy1pELqX6YEULiFz1b
dMY2yA2bjdAS/ZZTwI7plI1grpGvvSH+Igl+RXxxwJGxshXsYfbZPTyB/cfX4tIY+d6eqhfRKBqB
YnlNMV0kIDQgpPq8i9tAFPaJEKIcHIcYSSrvgOFObXRLE/msULTjbHifVZrnTMwydRXO2u7IAw4o
aE+xTNVYBN/EVn1YDdheUpltEgvXIAcX5+QLgSRc7Mei5fUh+rHniwoCVfC/RTAVclLhnrol1s+M
sMiKeFecEI8FDpBU5+cCRz3ImCPUww6RB0+JDTl4pFZfD/G3WYTbqppUCe55S5rFRHJfwusJrHC2
/y2cupsnwgnu9ZsHHQl1qS32toy6IMJSx9DfUKlNOnWLHmOaRy5rc6fC1RYUjJ8SgdE+wIfQ1+cj
rcr7b0YwepSFNb0CC3wyW9AdWRstqZIBgenK5/nyZqmqnE5rhN83UxKBrWDsBZR4ACFx80KTMWtS
Sq0AKTEhs747TZmtUyi4yOzFVnfHy4AS+vjvQrvgOehhrfloKrd3DIVD4a4scIU9huWe8aW5EIZe
kc7SfToCZy8k5nhSrbn468QsdxRZGbP7glsX7qJ2DDA+kj36JlFIxnShbwyuHEdFuYQeOg6xoYCF
5RG0TkUrjX3OVVWfbiCqSf24Pt0tuL5odjVOuJTcn97BiK5AfTC/1sv/yAVyl8MULB7/q7f8mcKE
R58Qvkk95AY9Z1C37ogf8PkqlCaR/s7MKjPTmg7Lmf1LpQItVOxkDwp1o7IttcMyW+ac4yV8eisk
AFLXWQjUYseY2VC+W+UK/Tn7QMpnzN11eDzTxEokfSZerguPF9xz9DRa/rotaf4n7xAkEAKs3Q6w
xRtp1SGELLY2f8yuoAMlpds3qpxbNzfT72BqL6GRtmeFNTzbr+Y4NME4uoECWCxU6GOBSKyBPvaj
kJGvdovTGKHE1WrflJWr0/9pGU5GcvXX/hBHpzLvwAw9O/xVHClOr/I8YNLo6k169BZPgd+GJdtb
Z/+/mCg1bTbgHgUCk/09sq67BQAOh0hcLUAwIutbW9TWaUmK3VDuoEuuEsUF2fWH6cvI2IOwX+UM
FQ+Poc3by8w+Auldl6r7ITkzc4YKytxh/ecx3Ih3+Amk5JoO/igVn6q2v9Twt/g9RnWH2Z3Okayl
wcSGlCwzT3zl8AZySQn24dS6zftssnXo7oYVronoIspe4O8T2lGdrfzy6NRwf59CVmtd74X8zmL4
46WbkIlz9cjsRqo+mdAzSSUzO2wSKqgYJcpd2lmfR/ZlsfONStWAmQtF9kFYL39G6q2exKHOyqq3
x5NJ4aPmu6GXQFFemLsEnqureg0cgJxY138jp8tlDZbcVMI2ZqdJgDG9BLxXtKotkkrV1xv/toPl
M82zhHHspRMocZdkYsxywZgvsyNsdf6HVSEP/QjDhsaJQFHXx0l52mrqY7OwWSpgkT/unNZdRF3O
BEGvzfWZQE7buz3wXDI2aT0P8xaD3ZqiriaXeEHrgmgvNdcTW1YhhLoBNx7SithysRA4eUBKjZFP
zwuW2Dz9ziCQ4UEmFq0NFI+UpX8S/67p1Ly8q0aevswURg/0llnF8as6rF3QLFkxo7P9MO8NFtiC
F9gRYVx9mrb+dWHhTqdWNCsRUKWbTp71W7vzAsID8XOlMewY7EEzB8zuGQOcjxXg76S2Fs/SGSL4
JAIhYk0/aRtC8JrI0f0IO2pLdXOnE3+T3U9JW5GHTMjXeLrOS/qie/OwuuQxEyfHr6LkEvPGhyMW
pI8xGXZ/lr+yACJQOODkbDb84kisWgwiAZ7E9wb1lnxqtGpKFVKKR7IcxisbJa1ZAZZcWhxm9SID
RqtDJL1QDYKhiukbbXZzu75bgjuq7R8WOctriHIEcONn/Mr3pp7F3xl08nCSs0cKEEex8RtC7604
G0rh7WKrKQpiYtWqnC/Xvbz/aQBSzy0WzIZ0M0/+2iaBscppkoMTPDAlXoXpvDqPi4eDeWMNT18U
0dMb3PngQMeqxEAjXAPzDVs3Gl40aoXiXWl7wfJHaV2+nHxMjRsDUhgmd/nzIFL3l2bU1ijhiGd+
pWGeRedjCulWpJY+cbxM+dUv7cqWbVy05Nabm2ZMk7PeVIlPPU21UTvV3clV/fL0lX6qQa7pZOcu
yWTT24YVO4d36P2EwDjcxmigsag1oTfZIl8Cjc2+ftgxv3b8aRu/xUO2oLeXyh5TUG2FSVF8+aBd
kA8Yf74j1jM6xMSc5Gnfb3ViJ5MjdJ1emXIKEWg8aNZYHbw5E7w6puuWgs1xEwYg4r22np1biyjK
VCF0zZm4YEHS5sV1M0QWayX7JGDzMY4sKQELRXLTB7eWtiCvk9Px+SKVatBYKO/UNwMiqTk/GBMu
72DBY9yR96vv6+sSoJUJWFrWwzU1cX/Cn/e720OQ4o7HKeEa9hAomWxeP99rgGaTH+iET2geO9Ql
fblWSth3YyZgdGg1rt5nHo+PnsC5b6sFy+71BTrh0x1ibaTzLTA1k15kh7cJFFNxrCuPFKmi7gHy
dzUNwoZlGIvPl3YAPtqUNu3BMpoaQNKJC3vnsnwmcfyQjws5y0WlMXYKZoEu6UoVR9Q4LjnHLVwR
iMIKM07sxILsCaq4rDgGKYCtiPnyZuX6h0+vL7Qc9K0DwSO/Eat6FiYFA+YhZZGIKv6zIzoinE4U
YEZKNuo/DIB6agdglBxbYQyWifhutBkFP7clxPTW1Q+edE91DXeRk6YnDGfjgeAPGUhQxPkSexa1
A5YJPpgB+78YZJv8CiFbFs8jYPPs2Ah9BBb3pEWvvdl1tWrDSakzGAstQvaMfc/dcyGLlHWR7WaW
J4PekbnvG1ApZ18P2FBcRBB8p4HpbxUM0E2cMp8X2xNEywxNlwenBuEU/CT/no8PuY6QCUYA3tUT
XsGZskdCDSeAkOItoRDe3FTePzr2fGLcIqEzsmGpny2V9vF+jrqkQuHrgmyzVNDtwaZfMOl/Kl1C
CNPUtmKnohRoiCUHdQIiarxgrYCl4uYdD5dBg2z9mXVsBH3fR0o0kz7fREzR8XjcINn/I14TtAfb
3cZecNbAP92W77wASvCUxkXU39rJSQMIr2hXKQ4lPsxoJBSIQxphYBz9xwkokLeiUcWcgxsGzxtb
KhIWImLKUV2vCCWAePxIR+7sSOVIdfkpSSfbClskE/nFwfBUxojzKU/6hf0mdhQ4405EhzMV3sCb
vSjY2sXMKdMQIveXHoEnmnYcsh1x1S8qoiNSAUwzQ7tKS3KRtF2YQZa7Vzo+izKZhTBF5HlJYWEh
mC7eL9/6FbpwuQIy4N3mrCSWKzyCcEhun2GQ6RyKKrEloAiD9ZgHQHf3qH/d1LpOfR+3UBBBfFhw
Sgsvmch4vvbztn0iA17eBzO8e8XuNWGsVLh3niR+LYz6Eh/LFugG7dpzpQviYHBMroaW44o6mOos
eOG0LbeMCEAGww5B/BGrxTqjjmM1WW6OUx4Ra39XNSpMqS5SziRfI4D3bn9RkmetjHqAqoc0yph5
GhGPI7zJq5KiGdXtj/qipcBl94Fc0N+NC8FLv3DSIyNs55+wYYM6p5pcxv2Oscg8fdLlRkBGJ8Ts
eO93LPPNBveeD5M3RkpeUb9mwAzqcgVC7A9yhJjQK34h1kFbYtQTN3oUziTmC4ixWUzxq0cPg+zf
ddkQNS6NMwMIpNJ703FIW5Uz04gsHhIBzwE8NoJ6djmyrPaBZC+IDZWroYu7+jXgahQqLOI1WTyw
6cwfoTTge6kDWJCFSDFmJqCTJsysUTqg53qdCO8EMInUsaaNhJofWbAb+3K2IHRZwIEWx43rCW2s
FUfav1Yly/4CC5dNBU1xVTAkKpX4/yV/S8HGGUJJuUaYYIsd8T9j+W4f/1qFfAyKtjvBGMkosDf8
c15wAcmM/u8JpumRW6i/eH+pSRSXycD1XVpxSMLC15hKe1pihq4QqM9+fgS6bs3BJCLTxP0jtuQG
ZS9MFDqiEyB38hhV4exetXBSOTqCquGwKJg+7bjlY+75/FYYtIr3cyS6fwCzjEo2xBwv76bTqP0o
JjEP9y2+Jy2sRbHtkP3kOnt0XL/3DkNHmcDtAQYHsx52gK3XU6CRpdwCMkyLWOHG+Sq2kSNT/6f9
SNB9AI7ffdxAgqr8EyRrujc8UaqO6EtKYTYcyqVLt9ouArJbNrnQM7JUJuDD8jvUVeCBFUlG1y2L
hH9b1GU1sRcqWI3qqnATXTjzj6Zuv4uJ9c4CppfE/UvB3CosE4Uyg6uG0dp9TK1rQ18mOR6B+RH3
hHcb2W3DmfyqhdQ9kuHy8opivnBNuRkqR4GpMMQfvK2nOTQ9tqceTKYB8YBheViv/sk39RDecIRt
ijQmZTWvugZImqRmw6RbhkyjtBfhjbjuJ5wspsfFquG/vDNlqOEwHWM7wo6v9O2Lt4iJuKs3M1OC
HCNLJ09bNuUgd+Tct7jNBXjRlw/Lt65o65ZRV5O8PcAHl06MHyEfQSpFYPVv4ArTRC3K9oebhNFK
XO2kfIapJR/0wwmnwyTdXQioW4OwjPQgl2OHrJPNSMMNEdsFBZtWnAOY9N2zazLuzee8QyuvWdyn
PYzcGm06LqT67HU8QPb+YwjTDrrFQhtkiWkJRZ+adabV7kYPe4PfJ0oIDvRpm2F47VFk1P7FA6I9
Hmb1ZI4Ze4aSN1DTNdYckgHxIH+fZj3ytcddnwHXM+iQZvAAGN9qNGomCKtg/fTPR5wUaKBzP/Ug
ZFKGA3nlwYvqdMrp6F+T1kPwSWwRfsFkjHNGWdSLb/o/EQXVhFZBOJv4jLjeRNcZbrMJHJuscBk+
jFY+gjABp7BlC22BhX5cORosKIsrJIS/jH2pbT2WAvpDUDpaDx/ubYVHIJuunjCHNE9+pxR/wn41
dYkTMcluD7NQLfqF5Ws2dCDfpZbFof0uorSYiyBY8TVST/jFxfia0mwR+LKRd0PsNm5pp3t7jqc+
k2ZN7dqsRe3rYeFX3de8lxqTU+p6ulbr3gqC3dNWiXsWQXrSR/xysW3ZvbgCtEPG27HisFqqftG/
9V62luN3ocftZjxxrU6Tx/v5osMSPN63qf9wuQ0IS4MPc60guSxd/87ss2jecSWzWFyql7mUOVpt
frE3682ZHJB4+aTIRd21pm7b+cDwthr+mKfr6qmN4k9Fr1a/RxU9aZa3bHfJCnea8zPbdkCiLXMK
e9sZsGE+8Ys1my3MyiW7SSU6erNlStr8y4Jc7+WIlOVl5xkpGMQ4cOcZcZpUGwukShPCBxVUKiEi
3kmgPachQfELDUPcG+TB5EDvId7ipC5IjWHHOobryHHebzK7QPqJBfwqPItGJ1BIi8PoqQDwehWA
lRbyqRqI7ChrkWsDqDT4jCl651zchkPAk7fRa0u5GY3wK8oz0JyJBhHyS9YqznWDBQiZ1yEZ5cP2
LqwMKKUtn8Ds50P/AhA1TAqFHFY/7/tv3nMIZLf3lbbpcwNkkUb/maT/9uR2TDfVa4Agv0j+/PAP
8d0URU3i1znoo/Xu1BOF2glUceasdfZHbts2A2nze+c+Gi8ZjlMmE+N0Ye4FG1wSMYgS7Q7qoKKM
TvU/ubm6rxUdQGeDhT5Cnu40PIaNp00donZkpSVoNY2pMT2R8jqp6RW8pJLOTlXR69xYXzonjEaA
QTQ3VjJHxiTfAfjxQymzC+m5VG7D1zORZRpdWG4Hl2uZXz9rfIVDJAB8DidD5aXYisI4JDs1gXIB
Uc+XDQ0vIfmIZHtqKaioxzbTkDEgPQpnXKe1AhRoeSM1iy0SrOPUWQhmBi64aZ5CcKv/6k2fKQE2
U2JPQVu4dLgyFaebsjPYHtNacdjqn0HWbrgg4TKZztpBNLD7j+/FSrX173ZWLJiIMK2g/2ka8Xee
O39cP6ES0XGzXnmI2nmGJ+zdbYPDKWTRLrdaOhzPg3I96eUxw2pAH+X8SmdvWW6xpsHxf2lRDHlz
sSfF6lg6IkyKi4yWwNMuYiJLEMSQBECCugZM/ubysruratUlWIvYJQdDDWI7/Um0rhEtpLuZADDj
OP1K7NGw5PBq71l6Ho0aKT9AabxQDEuRka46h84Vs5Hvhc3jLYR2lliJJAL+4Ellh1U4VTac934Z
BH6xrSs3n7rIU9k1jZCj+LYghe0PcV129d7bfgyHgIfr/CRCCPDyTBXdIzyEAVWkiSCleV/zszK1
6ZZyX1urI2LybRgeLXaZ3DntEg6HvtVe20wr7qTvK6m8TgXa8JWeysDXjGhV5BoNJYjVfHpl66w/
FggbhBM1/YVZnMfwwnWTvG2J/Wyp4+10D5rOJwfzmxqdxd9ByVHO/9tq41x7SKJHzB0je2c5HhQX
UYEafRr6mefMbkQwbt6myUmI9l5Unfzur6v5+07eqikfRA0PGbDXYUOwFfYejJ542bnOzCj8UxbX
cEIvMM/L90d3OX1ZOv1qY3UvLnY4YDC96KRuOSGkw08P+1ZaykaKkXDuaxzc8fEEzL6JYjQa3OvM
CvA9dY7rDg4XbvBVmX36GJ4n5kY9v5Wr2YoMULBTOfJIPrnmu2f8c5iLqXtnYBvb0lYjZXYf7tbS
Azpy/AR6+2Dk9oxhe8B0YpztErF2W87QAhHmDqzigEDTBQi9XzTs25cL9rZRZHyymfvPUw46snDb
lGp0b3d+0dLdHD1IMMhYvPya9PluYdzzS6VRj5qxDb25lQR27dceuVdT6rDDe3BdNz+pbZJ690l1
LmqeKuBodCfH3bCarfk52kP671qDgs+3KY8QjtwyLfDtTvNl9HPUisXw0L5EmvBi+FMQpcmaJZJh
cpJF8+/MzzLASIsLBJIgu3HcBgID0hVlL8MdXlIpnkzwicbdKO892dy56dAL1zvj9Sa8gK2xTpO7
oqjXlrfIg1jClUhaBMuYozhr+GIFF/zZYkoAF9OIrqRZBz6ZJzPEuH/OW6q7SS4m32lOXxVjaPP7
hfyrahdjqBX3wVSCmchQ68+xzyv1trRAJVXZSCs5ngYApefUuFzxZxo8DSGB9QSRpprKVyxSxcFT
+DwzDbdfKmmIzndtEGA+xDOxIiNToxnVBpIz+DxmfHqpSQ2LAJn3+PWFJ9/3NJXwqURcGmrvgoUf
VD0UNzXMZg4FkllJTBPHp0OGNWyYLXzGrqDZ/ObYmY3rkHs2IDnxxouNxDcVVHqouF+Q1c4cD0sc
EOXqoHqRE/EN++vncBZNJV5wQttVY5iDk3SLxknW6CBKNcIzQg0ZkbPbnzotP3eTtdJNy8Q/D+nd
wZfgLrmRGfOq4153f/+JhLxCul042d91kbdGJXWmObcxfqhyQ2KqnpQnJHrwu4QCPiemQ1uKNYr6
v9rEzn1ozJb9rtcc1mLtp7hTPc6w9/9X94aV7Iu4cDWEubGS3cnOt81g5eFpZg1rEUT1jIMdv86Q
Nbi58v9tZgRrir0tvZaBJUAPXWo1P18uGB1KvmQixn6LLPU6BWPRvRYFShuNv1MqHorVzEhxXxPq
5Ek8rJS4cBc4J5DMtvp606Opc/ZDhMaVyP2GxRC+WhPRh1QHSse5Cxn6oXRN9Yyn2A9gn9UwidGa
9xrRWeAqqJ9l0QTZqbHd3i8bTNmy8H0VzUA2SXENvRypm/WV1Z1mUyx+ci5l812qi8pPExY+obh4
IP1TV6PuVD2rRP1UoCzsnz8i9POkLrkIQStcptkSfgqYDvgubLpJlQWAdpDJfk044JEcRofc3oL8
QfxaG73tZzvG/krCdY6RWBmKWH8uB01eA7pmrKaV2C4QLPl38Xyt2K4fJf+YtFqnjF2Yg7sXiuyV
70LPDGpucSSTGD297hwN4wBLgKJ7ksoSJmHjc7e8xkKqPd/HSvLou5HruoGJEgApbl7qSPrBq/2M
qd2Cjhll/nt0cbwOt97WI6Ks0omBjZDAZaL7GbcM+DcV6DK19KQziGJgBHemVjPZlWx+D4JN2AaF
az8FZec6NpAaiU5RmW998xI+OPh87BpnPhJvB8dROVNbkZ3vzX3Vl7uaHJjeG0m1vb6L9cC0PM+e
fS0TfGAbt74eEPQHbBQnaGnQnwaRI3Yt5Ue86knperH0mjXFgBYowGTzZcdZ0apTL1/bdgTri6gk
GMRZAlWdMLOgadeULtdMvJaMofOou1vXY9QU6YKjEph+KI4mR2aOK/UWUOmSJmFQ2uwH3+rDf9ng
B/5b4qWosDB350v6VRaHRH60OiePP2Gi9nLAZgO+E83gz082nCb+kRQU02qXR5V0sIVhIG5c/0sK
Ii8B7hilLI8/0tdjB3oPVhuNPMMhVovxzsxBEsZBHEAVhtvV1pOEOEXxwHOgsn4NuEFccs+LI9Vm
nY38YlrS+8/m/pzcUdGvi/5V+njOkceee4e9pBHWc90NrLU1LTKs7OJ6C0XVrnxnc+N1TPiuAvLp
sBr/J0jEaNSEQbmFDCWXpZ/5Gkeo3BIGOrZfOpaOxDNbDwC/gi3+u2234VNJR0u7/h2PTTzYh/ee
DgwCXYklOM9tIL3DSi2K7WW5U2mfzgRNtavY8KEwjZ2FULXL9eN5gLfsHvuSuauCLRMzzQd/robH
Ub0H77mPWmBnBPIXB4Nxb6aWb+vr9aQsyIqjGCeSrh89hYN342CKYItVap/3rEelkqidSgtNFApX
T0rh8gpX27weueU7+NOjh3PECvv6NuS7oJSfptAJ63xuUCdu/n8YIo3cGnIrriZdA53TqJr53Y8N
3vvemX+8b0QgoidRvSnZOwKYZeNMJmwMFo5eOXg8lMrF3ZlfM4CARySUau5ICqJXorFa0KWdZMqX
Jm11JMATLnHaWioX4gnKGaDOqmM6iWZMpE2KfQIWcyFUy6BgG5w1ZK2hU4TZpy15JK0xk+tdQj+8
sJPTzrdnW+vcimu5SKGHCAbMLaQPpDAREsPWJHvT171IauEhWftBuWywdidMTBRdGvlVED0gD0kN
SX8RizHk2Q2DbMS1WfoaD5Hp1ybWKhxiWFpPazZpXn4mzQOjHI9gWlSDF6scd59Skkjk0+jOKZJt
ASViUJKHbtqpX3LD6wgYqBxWK4GlFOsKCr8Np+EDovtqI4xy44Sbkero/ys8Nf0ii19N4CX1bYnG
gcRB3Htl3o0eqUcg65lrAhzDhdDcseirdOfB+E8AOPPRdR1agLQr3GDtz2DBNdz/hMzF3UYgNlt0
rvUgiyTbwSINqPU9IJVrEg5Ph6orz4mNJDfJ/HkhiYw2oINIUGTEf6PL38bYZak/NB1PxyPQzcal
GgL0kuaMoPx5hLT2DcIqHLMQnxW/qFygoDUmNB4X7CC2Ozh+Q0C8sy5moo1KoBc0SqYK1c5crgGh
8W5gQ7fuuBHj6kI84fvHWJUi987485bYkiTVSkLBQ0AXbgFEV9xt/Gm5w4ICL3MMsjLAk5dW+X+H
jGOuZ8pYPgrjvkOmr/CkAhQMQ4n7sNyzEwpNGXZov6qIinwB6eNKYIW/8ZLG2dAhZBto4kmcLRHV
/3BmSXeNkJfuSvxQKS94EtyNgjP/tp01x41rTeku9fmkjhPHPEFaitC2u2Y8xuMRXqOhDOyCOInc
giDumMqq+wgQraj9LaNi9dtfeeIFtfrqIdJ0zKV97LO5xvhzOWNtOoJl5kI47io+XX/7Hw2Bwg5N
vaOFykytz8USrCr65ein1yxee2rpNGpKQ0kXWrdqqKSsvnEvUZPcnUfpjh7mPs/+yTCiYRmmmjrE
W1sAoNy0sFN1IOcvTo4M9Ylr4DT7N+GMT3EfEzfMeljFhrKym682upIqi1ULdF2fzUaGvN/BQjvi
WMkQ85scllHTgK56VQesnW84tdb7icwov+zGAqmCOM47Egzb9B77DfR7mt+mGI6nfwaO26D4DQKo
hzXrmNSlKA9c5pfFDeddI+bVJg2hRvV2stfH2734H5uMvyf+pbkf6D9ZKELGlGP/YUMZr86Ya0tO
JsesRzAb+4PMFtl5swxoY4kZ7euX/jXcEqzoOvnybH6TkbvvtbLjcTduUWxGNqbXG6l84ea3gbli
BObFFrDVAet0l4waEciGH+yoZOJzJT0NG7i5q50qYkYmphUagHlsQUguk5FUCCczgQ8EfcMoiPby
CRWM5lTXeHakWSPcF6Ncwy91wSr2oB8Dxx4Jyk2zYgt0tnUQ21h4Nb41ENiOn4YFRpZMxK9qTMS1
IyTHkxyeKGha8c/X75vCZGqdhSFSJafgIUwmdHh7TTDkSpUB1i9Lio/ZfbTfp28sUwTRftB+UzFy
Pr+X7658RIZ1lMXSkwg0vlEcTmvqpCiG7AYgEFdVxMsOseUYrw5bljF1lDubel89SBsajM3ecdPf
C3PUsF5TE/EQ3Mgfe8zOWErCM+ozAfBefdPeV+XLvBQPsz+9c3qJQzZKZolnAFWO1ho5kctzAS3o
5CXp+HQK9mQmT/JN158PXQvc13XpvsRCy3dNt93JibkIPWqjWqpAGu1vjpQtjrn9Wv/ar9BhppLn
lumgd8mJp+I3+V9oWdeqctWjunEa1QmAb1SM3fDaWlXQRx4jjQyS0uUQD9FFJZ0YejY/JluqQ0xA
7ZK9UL4ouCr+YfGdyjkphIbGxJ3TJtR34rbsQlasEGR9lVQGzRxo8vU5Lusz28U5AKOE7KkAosai
wwlFg2q9rXRkvcV+ChWcboHeWVzTUiVOHI6/fJSAh294zZYynC1r4YInU5uaM0y3re1bRWe3uIZI
1wdM6a50KGLNi8haHBwKZQvqhJBkzN7EpZmch1gG6FuIXDIqPBRlGnT2xXTcDUoryiGex1YwMmx1
nY1Li03vxULAH4h7awsL1zI5qA7UdkEzigZOrhhku61Lj3rG4RxwUna2L+RDVMaaX1RqXXMWkgGt
ELPwhdI46HT7Jx63Q+Id2fGvD+1TXEf4jAfBH59G5hHvAddF2kgovT/UIgBtZ2cRLxdJKVScrz22
MESW7h2AaPsB+hsYaXNkgH9nnwrWBw8uBiwJBK29N/mK88MWWtLnUwNsCcmfKN9zOL/gE5d5iuav
Fx5uLGQgMg5DppaWEvfDy2g8UYvzkftO5GnQP+61bBH47oUWhpTQxHPORMiP4Dhtr/VTF+vr2yf0
d1RR5vdiV3YwMyUvqy+nPQGVran/SqOQDiYkAwPtalJAheMGtTZCeFk7E/B0DFI0jiadfhy8m4HH
+TFX7g8SwgNu9gsMatoU2Wqx4X5JAWIQv2uWpjkTYdpzmEKhnB+8AZ23yJwdak+3VWniUfOwYLvH
LHg20Eo1YRFwPThK1UnuPkfJZqHF6mHfwfavZxu2b4PSmfJszzmFA7Z8jVNlWn+p6+9IQdA+JPUn
16FLbenGvupxlAVIj2GimYlP6pRMKw5bAqsdyHJkxxEJfzw4Bo04FSCemzU/Xk1Vp8M8GVfXK05v
wjT0G6mJu9ic5qvLW0d7Z2NP99kh8jgQ4yUhH92n65oup5ye7wt6X6vCS1+p6DTkiEaywxHECnYv
DiyMBeHyUg3/eQ1G8Lx5m+agT+74Y0c/A/1ylHFIELcoJCqLAgt68hmJ/78DgOMSs6q53/IHHYq9
fI0EsjBRbmdzMlRQAwAdh600voiBSVdBRuk0s9HGqjT5KvjvhfcWOxoAirDhBiEWHFo3sWJFm/eR
KuBKnat/kUYxtx/j5jvGmvBYMV+TQLJ0s1aLlC6Mw/V+g7akFRm+7n/RNGMammw2h2k6GZmoeKct
AJQHMVC7MXGLX30dW0OpWVYW3PrhvW+kJeIdCxcLP+yWQOrai4e9YS44c3AHMBlflvxyIA1vecua
rrB5TztlEhjI3J3se+y9XFEL1WX+sCDf22tgAoc5pn0dAvvXrqaDc+hOfYuV1IkMzIgsvLT28Atu
TbbM2OPD9y77FlJzQTqFhSlQig32iWH66MwViY/kelqlf34Adp5s/DhtT8LV6zfsPJiMpmRE7PKn
4nEaXojrr9Np4kY5b6tZ1HLUROQgjP7WiAq9Q62p4qXeH87c/zLtA9CkIpMS78C9yXcwbggUUpeG
qHBoffw49HICyQXT5x7fn0AVvD/KFCgFC0ip1CAB/Bg9xUAt70aJxMjSJSMyeReUctgzAstDb2l0
ePuyOt1eCMLeJQuiu8x6jrh0he0DL7beoiFCQcjXIMPTTkRiE8tc+qZh8820RwTRCJk0c2pArSRj
1W2M75nCzEaLRzXPxwETpTSYHDDZkOb3lZ3hdu3gATjYHrpOgOZdKF3OWiL0MXletfxOREDOkEOg
t5e0WvMKz9DfFo21rE7T9+etByXt7cOO/7ljaU+Ee6opgRyQq8iYyKeS4g+qwJybZaME5Bfc9c7e
u2oT9z+T7RZrAS6w4Uwt3/sOOEDp6Mn+RCwtnK9CfsdNWIz2GpAKg5dctprbsywQu3l/NngUSRZv
KCClZG9aN8l0sDFP82eQ35RoS057TQ/V+j7MFCnpYlHg0qnTvlqEer30YVbIUQ7KaPZFB1sjD1hf
FoPmCoddrroyCi8RgjP+xmsnbGEm4a+hS6o5W2Ap457uShi+jZ1NVteQUuFzJ5v+ZoOefIkt7YKH
pE6iicHwvom8U6j/gzXClstU2t6DKl04Uz+3XqX9CihDcbSEo+z8XtTtkHzFvw+U9RzfqGgd6a1Z
PVqrskQJpwFZ1KPO0V3XCF5EHBe8qdNhxFh/5EBnN8m1pbC/Ycnwnt1LeGcjvz9v3uo4hkOh7pjp
XbzH/eLCcofx3wn+97t9B8WbcBKUOdTABiGlZ5p06cK30h/ex2CwlIe0MSA9MCbLi4NrRXmpyw87
rQOnl/uZ54V3GQzC9kqyFVCqc7eHVfdmb9Z2k69rgHwxb/RJ5bjbUV6r7QvfoyNgToyRWI4M78Tm
BCw4DjfKh2BXEGbTzu8g3eSzTT5WZA6qzT4Ec2puYMI/gDoPTWnipwdecrxrgLWQra4Z8RAiiehR
AVAjHhW41102oqNOwpax8E8B4yM2J5V7vKhoKKP60RZMVq9Zmhzy9hnSJfRkNJpLFSAo0TAX2zx1
lXdD/4AI1Utj+FokHG4lfR7jrw6dLywAs/EwOO9P6CYl5Obi6bAT2p9GTHR/B2BY6g8aZ/E17gtF
TCWb7r9RcLFFp0T36U5qKLZmLMWtRtv0hatIAYKtxaMCI+Afb11laiC0wmTPEB8GqrVTDcS+ngNP
Nd84sbPl5c5i5gOus2qP2hn1huncg9sxQhlVE8l8RObxXXnnPfBYA1t52V60VSfWYxTYvhJRtAqf
3D/74b0AQ/b7g0qFcsrCzhqf456SEzHaqYDb8nsciEP2CWIAjqPZF82mqwcLh4CFMEnt7/mWS6E2
dPdJYFFBM2zwwFLsqrykYWbi/TNjZZONn6dzV0TeNU1KusroG/KuvW1LNDmi6SXWGE9wcYn2av81
fAWlVnZz7KGGvMAfX3ZfJ4TXafxg6DDO9mYWCwt5xOzKa/ELUbv92NLDqT3sUEjAXl4MLfJ+n3q+
wShRvCJqsJq7fome3Eq3rVtjS6bMZjMgtEODP4HhvYFUJ5IuUKGiFDq0kWZ1XhxVlvzXCgp4Hc4e
71zayU4OSCjajKBIP5FH/5SBJWlS+S80s91tyzNFaUgn6biNz5xGYq/1L0oWT4KkFDps/hvcZXuL
pq/2FhLS1DjYuggAj3lpIeiqjdJePDp0NGF97dyOzdTK9+VDUpcTtkC/jQT+lgMPb3t811nUNzO/
yUQ9KueSA1+GaMgZZjR1MklG8+kZei1zeNeHCLW7txsSzmKH9hQm7JRuhmo/NyucQD3BZCjj6OL4
/9T5Hgm9KhcHRkxj3jj/wttC+63tQH3IxjB2mLOJrPm2nFVRCbk5gxu/pRcGwwEfNk1KagUWFNmV
PWw686CF+LkAo2HLJqDO1fLnHKafdqwTXESf1obOoqs6DMsClQUr1GR4xGlfUOXn+jolyFFl98J9
YGdHn9AXkL5SCx/1c4/a1ElYgeNL2g79FJBXKEnxE004C5f/pYohOOaCnujkUZOLJYwDHDzTio4U
nd6rdJlryeCZhQvxt4ygEDeu+qVkth6h11flyjUeFDRvYsZXwr6Mkuv7Xx+JzWU8snF5qxhUn52B
5np0/BcG/k47mxTdc/h3XRfgqk64j53upRt7M45AEBF2qWzGD512lEjGGuL/T3peExd9eF+0EhDd
jV81AF3hejj7hQT8q/3gRE9NKd0F40Tu57PtKyI3nhYaGFPgUKQr+vSOaBkcX7UkpEuUvOVbF2Se
rnY0tQk4cvJ9bdPe+qYHbZKzkmFGjX7xHZFUwixhm+9Ij4A56Pk/D9mieoVZ3HsWHXI4C3CehUUv
J17OuI968MIiqWeNeafPZrZ5kRxd72pKI24H4n/9iYSPCQZi+/QCXtZeJpepZdknBMXCeijMLRP5
j7ScIe1RPa45FSCFBvdDSZJerYSVtcDMwKMQzaMmjJnrx6jP0+o0oUh5iAWjGnU4D8ygEmshIjAI
tJVx26YP6JyT5kguLcDRR8ORMGpGAdyFVdalOU0G3+JFV0rICnaTxZvvits0e8QXjHeCS85zDXDP
wKJokZVYBOLqcBaO8Wb/JNH+jMfUk70/CtkewzPi9rC7Ak6gaBMlieOLBcWuBwXf3hdkycltGLlj
kh6aRcSPwM6pa0U9wYzLeTzQROaKekX+O+ZchcZ0QHYlZ20/0ReepHUSBrL76WNfD12Ubkiovj8y
EvFODijKXA5IyNdAc1rh7fX3FVDW/QO9kBoHdjQnqgfOMfJuwQ1Bz1MfoV/dEKDi1BLk50orHPCx
xzXN2B6FeYYcnNg9Tvk5bvXVRwT77MPXsKRemWX0fI4dFtCpE3EBz0nZDioNi5zTrsVqaVwnUyUW
IYU2L1bnIm68rQgfk5w5ib4jSsaCuJkGwS16YQotibt7V6BqH7HDsvvMK5rSLj9ktQJlfwLci4fA
Zj+vOQXBIQTgQKX9Ts0tivXRM/ts01HzlkZ20/eCUbA42G3VV3yYTsdaOsWAYfnfVwnTM5rb1+tj
ARY9CsX5x8L45ZAeKECdX9nk5IG0WRqMU6jHel+aiuydlAos2p3jE1lTertD6zALFatQ8saicmRG
nAEa4vGjXfrVaPVwpNhSvh2R/VSObVk+kcGzrMOSFJA1xxPDcRQFtxLltsKZY4NCL9lqD09vVxVt
Ne3RmGnoAK+pw6Ra4C3lPT0wl8B2cwZOo6Pd3SAylzf3Z1kQ+shxUqgEQUyNQERGfxQZU6L48O0/
UC4TGu3C7vwLPqZqevCeJDeTAxt2wTCwN/CvnV16+LJVmSZoQTn/gOKGHplEl3s5emwJ5bW66Gvk
/w2vEfjQq5On7IGLs0iNlQ/3oO229qSEAj8syS9uS+mJLjcca4ReiuT8To24y1XRIipr/AsmenTg
E4KWEIG7jxbzN3cy1WskxiRL6P4WOPcbAaEL6oMYqhvM1DiCEkXaIobksGBPnt4PmPeLqCPG4xok
2q/yuF+e7y4hLHDUh+zW1gUnYUWLJv4g6BwUapjOFhv7OlLEBnhFDZIDrunXaKzukZB9Jq3oHEZ7
5kCdR2coQcc4A0LDgem5CYgFD2FTPUM+zUlir7MU93yRehFnzwvNx+EcEffmXqyP1u9/XXPKrEP4
OSPWOCQ0ENlgvonbsQJhUy5+ttSwktuCIxozpFgY02L37mWPG80mHwT8oKcxhC8/UM2yh4ZhBsN0
Jpksna5k+qsLEk5pwwEBCVVjDh/MVwlFPY5/BU6NyS8kQNk39mIgh6zFWQVpWFl2IkSKkQucL2Px
8NylFgeZaZ2o9ZEvPvItOEF6zXCIP1VP95RdXpyThUJmjREpRk1fNz1Qk4aYZCM1iMWUWeAEdhHj
bE3xbM4TmpJJAEisprcicdZo346vw1WcXlRwOFrmgnobOgtGqO8Rmd/Y1qRr9tfMyJAroEXhaKN5
V2DJ06ZcdktMoLrVZQilyuNqYoFvVnkk2RVoE2otUTRrry3GmR0CRkX1phx/kiMSJHr8A8NHYYcD
jH/O5nk4BZ+vIFjkEqWsmf+IvVVYlHv8y05WcMyDJZprrs4bU4EtCELVbyhy+8l+f/En1L/cnu/s
/XKNR1RULrVllHVAZoTHNaUtC8itV6rPvpLWkk9cHAxThGbvm0tSkx+b8BhoXX1J2Rfj7143eJ1x
+Mwy/OVH74Bc990KmK9EbmK4JyJw7GnoD2FDkgXvS5ascOSc0JmV9ljekPD07q8nsWaUbqoXZvFx
Cr0G8xtyMXxxT5XfIy/0cXmg9SCdcVHOw09zw8szhVIU5lB9IDj/CrtmenC8xblzzUuYNC6a1/fa
Azzd8tFIbmqtVl8tsXQHJiK0MdyL9fi9wUIJsBD5o1gPKeCVaszVd7WjEymPIPb82C4EQuiXEZ6y
Y9r76t4Ky3swj9PS5zo7TZjjoBjdfm6RUDbW4cZpePXFoT1BMCNp2OVTAAWc7EiuSpjjpHfx3GM8
juvjXC2n/IqD3RQ/2HP6CdFH3zX7xp+1qjQ6hsTUm6J9Wu6Ohtwu9o0JkAJd79cjJR6K9BtXLa4F
i0Jj9xz3f/bIo1Qlcx+j4ytQpMQuDj6HeI3x2pnEk89PXn0AKIIL3ElZ0PqD3MJ6gWOliqzKVsZg
XuiT1OA6dbXVI3qyvP53bap/5kn5eBMrsYlnMOA94cSWI+bInkZENwCFN1lScNWDymMmdN5MAiNc
nmbtPBnfMTGISny1lxPQ+XGzFCmR5AU8eMaUM+JdzyE1RY2p++EH7U/VD9UvVuSClB9GS1PawaRr
uNuzLZ5k441MMcvQ1LqwE8L6XkmYkSL2ysKE3HeBsKCwedknxlsCOELXgNcPawOeTTYRWlXiOeqK
GuCF3hQu+TP4lcvqTa8j6+XU8zdDmPC9XDrleLgMRoQ/tkzRse5pQlRmXcyIQjz3FqNDd3RpdlaH
FIMQWMtAD2f1r4Grb0sC/L4TM9w27hmRx1slQyAY2BvlttKoRgoxhS9jH5JF6V3jbwnxf812BPDM
n1ZtHa2a0ByMbuOltwJf6oFykjqv15j3ToJo7oD4KQ9I7OggncmQ3sbqSRE8bSCt0fCDMPZKiZ9i
96O4UozJMXN+36h1onGEiBG/nkWZwqvr5b1ldLAFoJnWyR6ChvVBxWul/qoR7D4NBixYcVmq/31D
9zA6yAuYpDGpETkeG2gya7Ou8QuHDXgWR/ZlZrhke13wMOcBHxhyd/lMn+2yCFe/MKjinrpptH19
y2J+8BmoUk9Z/C3zaaRG44Cry/gINC1dcTgRmMw9fSw3TTWZZgDYUCOiXz0gngEZrfeTrHr6slH5
ihkup3t9RtsXxfirFPh/FK8iWjO+tRHm+QkSYr0NOUEBogNiRRAedB6gC9DcMo2BOq37ASgTBqzZ
bYYTKoUUrBqiXdada8DD4g4S9vhf3SilLeKPgKo+psi/EsiIgs5PrkLu1I+yg0+diODZUmVDrQKu
LgPwHxaW595eEU7s6EGp/26Sw9tzXejjfq3haPHWB1n3zylhC8KLQ9rtxgl4/RNgrXIMsKwGteFb
fHWle8aSkrsFneu3ts9onZL0eutn9JFuoeWxdf1onWS3Fo1Trf+IGz1tD0t5Yv1OR1viAZf+vbi4
9oSuf0X0TE9MBwEXwbBAxAICj2jNmHbNtq3CBOd+1yS1SCdu2Dm5D5Lx0aOy50JrtGS4Ajv9xyZO
eG8MCedvuQ92mj1dHyNLu84pz6h/5mCAzROPC36ejTbhqMTHWTURRrxf8iJ0OARSJfjAL1i1erpE
sPOVfL4B/xkPDV6L8r8vB5dT72YZ03nlrHW2737iCKz9CecP9uDTviSTqZSU4/85PXJ6jdZgaVcu
ZBGTswGK8NMN2VS36ZnbvJUY5FHqbcuIWbgjU5mxtaPn+1r7MI8nl7XC9UmRHp3/beKZWJILhK8J
HOISNZ2f2vHVxFa3gfgtcozeUE5XIaK2UvH7oi0Qz3RHjt+uDa0XJSqZrjhnKQs6L9JGvx79xjAn
hoHiPU9h8n+NimbuOekZ7u/XdKDZ/mqQBBWMo7IbRI0qEY0ZcjmjS4/qKCSJnuw/qDZeUhplqm6b
q3dTjv4CK6kiOHYQiAoPfIJT5YThhAyRtrgZ2HPKDeFJaID5ddqdmyJd1TI0WTCkKA8q6Rhbyrk+
ThLf7dqclDUO9HOiauET9/luIeMtU1SVwfTnWN2mbtafiHULONLov2Ycp2AsXniqbHxpcmkkDXay
t//LF9OoDlUaszKjo9AjGsrbFc/twYOGXIyOyJ3eyLnOYJhbTCIA3x8z0F0uIyt+jn1WtE+nuzwy
5QmgkvkqsqBN1TOU2+PtGxVjpU0nm11QKdFEpbTHgfJLfSijg2ZlYVBd3fzkBPlaeg760O0KGuwT
xyDH8pkO+L75nhrz0sshjEVXTyXYGYHhq3KxdmdP6VWVnPtWYxj/jrZHZ9Azk9fr9Pw3ZdmAGMmT
JAwZDgvcdmljfRzqbxkxG8zki7SW/gVkTbeikiS27DfXp35MsTksxPhx13ZqxcE864vEK0XErDr8
VXzOuOHToha2deyjiiT9bXhFupWPC7gTCiB02+P9Zuj5fEL/HTDmzmycTdx4fP46251/qb5Z6D06
lK5BrWTvgcyHMsRqYZG/eyaqnYWCzTpztAHKZ22DAcJ6Yw+B90L6M6KeLDjoIB77xyzNSbgIuDyf
7CXmNihL/QyiIlASRkQfYS+/yFtHmj8Wc1+CaZJbe9bkKp3nd9t6rsP0N8O7TJSWeGoDo02NVI3Q
XXvQmeKLk7s4VRdEtIAhBw2TiXD1ahD3bAK9JVng9dnXFsVFvow1+BGA7E2HoD0AqaJxsyPqQUyW
dBxysXeI4Y28O5FBZ+PsHQSf0ate63WzsfbOBugEqCFTVr4iWhFT0PZJDU9A/AV+H0eExvsvcImT
eiq1HEsHCzKUYLZVZmHBcoAVCTPcyuuwIHzajXPWsvPvB+5XIeyAdOnhbe+NuK7mMCTslSi9+O99
S5m3l/ewojvpzwNbU6+w1BrBZ0C5sCI4/1dlb/v6nGS07TKX7s9f5G4qtpBO0O1YhwOnmPqIMYjG
iKhR2PxAA4gEfERNnJzTFegizcWKSHyzPFOCLc0l8EU1OgP17EzTCCmtA/c6f/GUKOwNPGwNOORp
KtXs0MkvG4TBxQDO1qp3UW6cFtCuZPTsl4KIf//m8k89WQDKtH/BkfSZOWElTSJi5Ji5Vj2/LGWF
7KE/rx9Et/Ip5olPCzkNv8a3ZDNenqZsqr4ib8VN37P94oUXRgUnsv9mGVB3s6Xpa7Nj8UT1Rq8c
DHRprFXSTw/nLale0puMoRaw12WT6nbyNIgjLQYQlLD7VSPYQUEFVIe0VTZ+tb7l96Qm+tyv+cWm
yl7jMY2KPMbvR3gEPsr6odY/hyeG5shgJdxKTcek3y9UtYRLpwjxG4gOjia3g01Eea4NGc9NvYpw
i/bG2/ebvUk5cW4o04uY2YEIlOYIaIrjogIkPPUMzLiTxEA/Yns91sOVgffMJDbLqGOKABQr0+eP
K9C6ixkQuyu0/8VuFIK66EUKnpzZGiVzIzLE9qFT9tS+uqpqwWrDBfufxLXne3LzLk1RIaFud877
ZKasyz0mqiT8+o5jcErnHUa2Lybh9dGJJBhZoGwpnTYwcwluZJfNHUJXlVmj0DF9wW5Gvu8sTh6j
K41b7XaCaW++DPpR0XRD6/t/0sC+euDdUIYYUngk0KU4Fm+ebgAP4GjFlkx8MtWo6qPhCEjn2hJ9
8K+9TDW+OaCxo7oBLh8E1SMEyAXFEzJvUUhnnJKJF7RYhPBYQz3ngEwqW7M+NDlh6m9PvZmN30vo
otkIaCRF3rqCdCUK/bpjm05T3aneD3wnnxUfAXaoauMGoYv4d+IMcSyByVvugaBqSMIbYjYFBejn
SXDfdd1NxPJyrdG6+EztIssiXxGBEn5SqX6YaAew3G7xiQZJoAAQTivor+uhZhHxTZsrGO9OUhRf
HAAahBkvsrlV0MWTiEvWst8SQSYIG3/v+BYo/HZRHYKP3SVFQJ50i6b5MHfbsAZgHF00wd4FiW6s
DHkXm0ctIOz/xahqC0QnAFJtQYe51fKOz8oEF5jaNdM8CtzN4MMqSfcQQbHBmRyYzQ+ZbSlo0SJi
90hWVro2XBQsrgIvQ6RD5XwAHWVUhYcpEp2LUywP4We3Jqyt8e2J3eio1Ibp/IxgsANWl7uAVptT
gD3Bn7HXTxjIrRdy4Mx/0Cz9RaPpI+B5lTNWDGfU44V+/sy7xG5ZEiSU5LyHfdK9GKUif28kGKzP
OH56JrX9tY4nG9OAY7NOG8HPCa3gt4Wly1FLiZxnY6vb0Pk787i5uPTqJygpyFtXwjOJCJP5fe0j
v6MuvCHUZcchlzZbTrDLOnk1PksCZY42PquVvX8JkoxcfJdUv3v9sAR8bR4TqXYEP+knnpiHjcKm
qYHkqFDg6ruxIRjo50ZX7KDviHmEunWSS71O4O6jjFgjbrlYO/asO/cz7tk55JX/FM0f4MERPng5
f67qcFFZNDY78GtYg299Zv1jDVV8q/2C2VZGxGICKEgdn3UPXRxZk3XI1sANzLo+0QkpoAJyEbik
sigJodRHatM5dYOqRWLtLqeGVhm+Kgr+P5iBIY6MR8EygvOB8iTuKVbz3OqE/zoDfsCNlkA7NX0j
/KDN/LQhxzSJYzv8yGRZUERkQh6xl9c89+xskUZjsi3quP55dq0Jh6UZoqZfzK7w9n1GAMjtLn2L
Tfh3ikYPZFmXIh75sRMbijbEURiwVSphoTQqQ1sQjCNE9z3jL0ayKEhIdNwgGnlD0e6rO+M1/mov
XGYJoYLoGl0X9nxaCXw80EDqQAQZ1PPSxJI6IROvaxeZSCnEGrAo4pKvOjrbj2yYI/7M6YgbC7wM
zT3MDAsPmyI9wzzd/yO6h0KAivqozzxqcayLDajzBVWfZnKnruZgwZ0Jk9k5yFSJbfpmKyWFp43K
fgcknz1jInxsOBA+FyslD8Q5bb/dLNn8YMJDXRo9oAkIvJQrY2GHJF7xyHws1L3RVw5m0vmlWcK3
hiXTwIoaeIatxV6wdptfInegJ1fjjP3+74HLowjaa/8JvGCvdagJtLZlaxKzS5sVX4yQLGnkIL/5
p+7xATU3ZeuBk/J6zU0KCaVI5pa5JkenUcaq9BKzrLvCy1qLiXJf9CpqOMst5ijMBg8Oj13CU+mf
8sVAORk8c9w4+7vuFZLM4wB4l3JuQcW7HNq8Ttuz+77dLHDmC+Qpao+YnxYfX65KMFs7SYZXTq0A
t+ZOrfTtZGdw6TtwiRt0iBaSOAz7Ptp4JCI8PKn5j/czStYGuHnwHWbomosevkD5d//SqZFZsgRP
Hpezjd2AHW0Ba2Vab26We9aMCLzgSbGijH6p8KQo4yP2irHaruQ7cQkj3OAYmnTyE0FraB+goj7U
ZYbKUshxqDwwuytjD7goUIotA0gqSySC7h7wU0sdTfaMlJXLwdqaVHSkvfhzNay6wnZybe+pgF7d
13DCYZUFTluKEjvBs0SG0CyY8+ucBvP+rNyNXj6OHDQpaSAYUrJmQThyxWhu2kd07AOOnCLXcCRL
dUc8rx3vxpLKIIBi7VkMkKgU1CRkFoG0I34SNCQLULvo26mOtcm1Mex3xMEUwBWJfReKKOuaQoTh
Qb6xMI2QRNt2ZynUNbHp/6GnDrVH3zegeoiAJ9Ekqn+F9p6PNcLijuyCb7uSCsvWVEhyHN6a3Bi6
0aHWxtf2FEKKnGoEJZ/mcpvgAOe0eJWajiFY6VZM2HpBqr8KzibVUtop6l1W8+NbZ/ofFE6rkhWJ
ar9fHi5h7OsGFVSCuy/tBb+8oAdjXqzGwU6FgLJ3GseKnKC2Pv8RW5fp/0ocn1qdyhKj1M1guSbS
Hf/s3bFayIaxavQpqPTgFmTPVdbgzh26TBggeKis0BPvqIbGzLCkguSincLCVFDGoT7DCvnBGFSD
Fxjs0OCv6itX+dPphG9LzTtnUpmI80dIW9m6DfiKPoY2kyxe+ozoogFUWw37m03kUgFWT8kAFgph
3788SIfwqCLV2sJ09N1QV+dfwMBuHUjJJsU4RstRQdVnqBAv3LbaUR1b17zM1NuGQBYnnK+RuL0e
iXt4bqUSS++wV/XcijlWaFIuROsxKvThtGTWLZXNej9Frb0aoFsVs9IGEYWuxtd4f7BjSW26U3ri
3/U2j3LMOlPeFJM6pLzb4ANX6SNHJ5xlICPdXLadG+a2m4W+Blri10lQyTyR9yQ8+iLIkI1cc+gO
peFBLW+f0bNZniYcHap8+55cbXS2mx2L0LZuicfHO65pi9oDiSfme+mGzTeBsJaBsGYHCmHxqqoo
IpbKTOnOT42XGdX57mxf9UMooSdalhXu+hiWwi4zCICSdogYqsB7hr8bmQ8aO/nACMWaFwmaDnH1
rs8fHUVFryKjQ9KQGFZyz9he1Tz8I5cmuO2lo6zDhYGq4A8oUY+zQyLygGckR9+yf4C+tbM1RSgV
kxgyNA1hYOe4fcnMd7W+hNkmnw3hAfsv3/A2xZ8azEmCrTIV36+W3myrO7nMXWvU2ie1P5SgLYbo
dlhxCtx+6fYg8H60UZs4rJv2SVe2FaGrEepP3rg6SV1NUgz/rCiQp/spIQ8Nn1+AhvJ/eklNRZp6
SdCCH/3LXThbiI0u4DaYlaR4ifVJQ+0V5VrCWcNcReTAGagqYaFeEYbXrs1D6yEBfigk7zX0dCFz
jw4Ft29HL6q00rOEXfk0OgGCen+71L/nZpQMZ+9Nux2wYKm7Pv7vDYRHzgtRbwDCgZWfF+HArrMW
mvctoJH9tQMS/frvfBxJiBExNe/i+47dQpc7ucfkiFHTeoAcOTz0Y4M5h4PSNhmavF2NXazonSfV
GK/LT1ToKGAo28UXYIn3JEE7xIgCDDqFclz7KKQEirv0hfVrP4f+6XdCAj1JgAAap/wi+3LkQ3ZV
yNXjWXgorgSAfkFufAO1SfA2tscipI0kN4VnUwNCmbDJTiOUnljOR8dgJdkcFGSXJMh2W69j3Pav
zrnsKcAd4gYBjdwp3df+wNAXxMjwF61/XCzoVg0HZUF71BQEBSIlwZxQVpxNXAxTjT7SrUefYToa
8vfuRYt7fpWHAc7s0Yl7Zyj6rwl3Vgn2wV8uQ04Je4N/jQWiybsiCLsJblZD4RpRJeDNaUYgb0hh
4UkUOHlwn3WjQOQBgVF0ewwrBcya4Trb3uAtvqLbBEPNRT4LOcQtyq+F1nBTkeCN2WKvP4wCLTgK
XtJ5+6nJLdVLsMhbnfVrcFyZ0B+xziNCyYNq5sfVPykqvezLWMM/2VmlaV3gJh1iv0lpZVbRiIoR
84h69MB6w0uHke6B35KUXwXgwyizx63aJrsX0RsiNaeXsVyFSWx0SL6V4R7bdXxpbp6tWUqrVBFr
y/Yr87furoOQXbIWJKyvoXIJUlDYu6ymf9KsbJOo50+zrgGEWdu0h5Om3BI4nJCbBV3J6+kWW0OX
bu/Ts4tBW+PGM3W0ZjCNYsTSrtpLjw9vOr1jv4/Cj/TmQrsmMWu8WljXdnYjshMGpG4xWkC15IwB
OGUVpvHex8Zyqed81CtsD6GI8do95VX7n7/oON5044Vn8vlBPUVOnmseDUJvO3nQ3BcrUeZpiZs2
aPAj7qPRjPLan+9YmY2gMQYWJRjByXS/Fec07VwlcJy00kw6eFColOmY4KsREKmdbDUrwImzknme
gn7nqBGB0tVyCyTq0mGbvkm50Ia1NTCsuZYj/gEMwgfMSpzyx+SLDiDGyB1FojmiCKarSQu2xKCw
SgJDksqX7q/c2tHKlm8AfHTAmq4ApWtIawyne+aVkQJ3z8LvxjfoTaMxAminqptX1tbaMbLjzlCe
AZI8NoV4y4O4y1jW0JNmk2ASj7D2FhWNs288Gy2gPaxZmnM7JSsIVsa4jVjUITo6SEkQie3vDO2P
0wR6Wk6C1XsKd6RFnn0jxm4MBXZ5ZwPkc6X2ydhgPzfKhqXAJE3zHYuXIEdQboSv2CDHSM/wsa8L
8Pw/Sq8LyOezgBV9lHdCOhgclQLQMaN71pZxG/vGm4y/RLdHHG04UKtZiPL9sBGlYkOTmOPQPozV
lwvfkcpmU2oOxE9dW9da5c5qUdcqVcR75p8nG5NPh92bgSwfWxO5saohwbzecvuPtttlha+gX2/4
3bZ9uYI/8wcJ6xqh4Q3v/XKpDgOwGkxPutkC74HwoM+WwdHG0AcGngwPZe1FeK9Ge0/kN4XNPLEl
S/bEv1qSWu43Y+4vjgdknLBO0hLLodYKweNTGJSqBsSbPHgzweAbQylgB8G+o9McmxLO1AgTu6cl
YtPjNgWNicgArySVzNJ+Xo16dGBxepDVEz2VBvwsuIjdggRgaoLRVwQTyPiJb4N7v6X2T+VNN/Hi
rObwv3sNVug+IQAdtaJV3SWEOA94OwmcHQmtA0LSEHZjhIZK0Sewh92sIQbQIwcwD6NEhl7H5t7P
BHKuZia3ylG0BdKMt0wjMD0yL4lj15bQYjZ1fPBYk/qJmr9nUAeIfbxVK3FfhLMjk4p2AgC5t/o9
761pd+1TNc/tNOpsSSrTyfJIr8lNiim2kJeKKVT2gkeO8OJAly0rOqqGy3l/Y4s17dzMS+BD4aIm
Mm0CWxpXllYsDnUqmNW4bRGNqFen5po8a0OYkm8EAel4vIfSZtSwylRdyUTZgIEtZGy+kaINXDB8
5xWH6gDySRfi2RqxHx2MESg2YThjCq3JGiDBuje1C+ZilzRefOsloJKNqra1Rz3/0sODSgC9aZcD
0I0jDsUJaSAW36vf9sFOVW0WtBoZhGKOQbxzv4o5WoU9BC2WHbqi/rmvOpU9cv6utgDJvEp6scWU
f4DBjJvdtL3Am4yfwHq350NXIQVj3EMuxomViDXh7o7K+yE9BEgxvYc7n4iQ39e2/3EsuhYe1w6i
6RxJUfiPKW4+E4LJE4/8O7BC7/eGXtL4O3Pbb9pfTDoHBobyziUGmy+0WSR81yyW4CogwN1K5glX
MJAISx1gKgngPQLB1IRtHnNS9ql2qzpPw7Sx7bSG2AsyqU9rMaW0JrYsX61CNoc0eEetbrY12veP
/rs377MUh/ZuLC0z12rmIy4FTlPYC7xzj3GLepwuzPgGc+6vLjqj67DuVpsTbHR2mjmcxq+Pnf18
MrmB1fo8BFyWMR8q0s2Xnrx5CGyQnjX950Au2GmdjKAJo/++hYSqXw3r6cX28mAva/aYt7u4+TlY
JXr13L3Q3c4N2jhCurZrxQIpC8t1IsbVTBysXa5iRVruhOXuybxcXA+X2ZdHzDZWkLjU7XEBtf1z
lqLarOcvajfH+wrE/8CKVQbFruUjWg0CeqXoaLcc31H11ygnMLIdJMhwq7sDLLj+AUqWmNBCWtoP
QWMx1iPT5wDXssj29Vm3gGfyqhHKyKH6qT6hbfMMMpdMLhDfIBgG4Bgh0u8X01Khz6sPehzYwAIJ
Inc63xEaYhM058R2kIr1SmRm4de2RSMV+9Kj3vIJD1tpRI7zqsjYVpYbO8T/whG0YV8kgtwU/rAb
Ea/0WaQyy8zLBlaGC6xp9atJRXJABJG0P1Kdvu5IxeyPKAPqrx+9ERhGHH3Jpk9HI4tu/bD7koXP
EZctUHa0Jg5D6UiGhtjAeOMJTjkX3lREyW8JYc6rO0gvPTrCm2hbezvs4VPF9a5GDigWLeADiAGX
dLv3Djcs2Q/rm1vZNBjT7lmG3cVDaKD1rykXHKonFuMhOkUC6ZJhTXC3tTl3yOBbj8mXFfgoQBQQ
BfSz5kXPoDtERChZ5pNK+dcEY+MuCv9KQu4MxMn6xD4QHCRuTdASWcr3yMGwGJwjP5NdL3yE5ptn
CpB4/k6JSPlh6KBVucUc0T3ipSpqwYebP3IPtqfF6R2lsEHVU9uilYW/apXSPmRlIun9Se2crA8N
5V1xn8keSjyf9h7/GT/iJiPaa20xRSpWuyIhNysD6hKdgIdYWnKvh/m4CN29yn/fGBuYyCL1U0JV
zj5vKJjtdtmNw8tyq6d3trc6EakZvoc7c8h/dL9IfnXXOsssoqwDrbO60K+6bEngcHCtvPB+p7I3
lvdkY5sX0O/XQ/cw9Cxjq1DVjlvrbK879qdDJTt13ezJNXOqS2MZlVE4vZRipH+QsqWKlE+4b1tP
KZntIDtW3HB3RaZiRaclj7UyORSYD2t8HSXyA7zp6CLDE9MmDlWA8T0XxWQjRH5LpDJQv76HKjZy
W9Ksz88hvhgcyydLkmYiBuczONzA4VauWjDPshM/Nyt2gW5yN+Q+FvzeYcPHL/kxcUndFDRLgwNj
mia3w2m08kuYSrQPRuR86ROJIRr+LZVVmPqOFgrQZ9I6+xe+vrH6eHLhkIJIFDFMs9sU1zSzKdX1
bPwrg/ABVPd62jnD1mqeB0ikOexMWe9I3I4qs2zD2/UOour0EFtmBRvAVgjOLSyhvsi967Vm3rgJ
PwQLbNouUTmFnm1jLCru7lCta79zifdCbEddErac4/keX1ZZ6YGgrNWV+aPf5H2DI0VT1hOwqRF1
uJDpaDrddwYGANlGJL8mOkggu0phaHXJivIODcTs9MYt6suvp34l1soaFNyfLUSC9yDCYn6iotfa
R6x4x81Tizonf4hD6dUsJivhyr1qkqyOd6gHkM+1AzTMQk3lxxeR2K6Vw7mAgNi/+VUXdCT2qqwQ
26aSFxL0+urfjbDeOdDPEH4zRCJeeRuPt9pIET26aZ6IoeQcRkSFrm+f3x66M8+fDU0nuarLnBCN
Cs2emSMYhjdhwAKgrovhmyVqEmhHyOdd/0NfZRhBTWKZ8Ugyj8DuGUowNb4FqiKlkM/MsBRMcfXN
p6IZJGlqszHOd/cC66MC+kXMDg3t4x7oCVxI8HxVs3k6nMqS89D0qvFYUQA6NNEZqHLg8liQyGP6
OP1r8iOOfMqK9hdzOejRG4E90y2bfjiOI8tYnWvA+Pp2FPGFlnfkxf1Wes/+e9MAOyOxiGhjm4WX
9SSIisPX7bBldR6gN89bZERg4MEHapM1jeN1eai5UavF+rbTClYwYXhwC8Xsgye2u6uLfDAuRwTP
WewyKTGMiFRT9j0vNQIuGthMOfVNTenkKsVlzgYeitLr5TqPxjXa0T37l4HJ7lcb9F0WVWJQaY1y
txDJ/PE5MYze7km4nS27irhTl93qaXakdpZ9SC6jj1nj9I1wK/TCQjHknAPh5qlJJ9f36nw8YEdJ
4dndTClLxte9jjp0bLnXV835Pn4K6RLHMQPQE8MypsHa38spzCm4r10DUFRhCHcP4J3ktn9mWdtO
URYVJUqMMuD7FFmvT0SbXf07Aipy5Zk50U8mm3fCldDiJljGkt0+cViYabzzq9mt1xqkp7dCUdY+
k8dyRRTENb4B293AUbLJ7Gwr/kSGzhjowclJgCts9INLMifGdjOXgB/uGOHBjMw4LeSD5vNs2rpM
1vDXTkXdHAUYdrOT82BVYpPs29BhgIN0tVmgWtEloVdJt8uqumRhj6dZjidUiiflUUyXV5kDGWTB
3NpysJiLkON9S1sotK+c6A3R1SM/n7vinXuHbwO4fMYyGpSEqHF3U2cKQjA1N0BE+jyTG99HjGer
fdhMm1FvH+WNUqXcIMes1RXcTGIx8rYisdm3TDiy71T0gBLCEyiLTcnaWBSQfv/u8HjpHBgAYmqX
4X+Ullf/x003NUvm8eJgyOesdHRhHEinQE3+gxEfRmmOZqiHUGwoWKKht62dfdVTHEYQviESKkhW
S6jGmmdXCJlU2JCWaf4IA4WMoOgszyDtGe/sYx3nTIZNKviJMeDwlsD0sTisBVAQwY9O0mNHnxkP
z6QXpGF0eoyCWaFj1CZqsfL62vRG1S+j1kxqEOI/2oZaizqaEVTx8YvrjDMkjgh3ITVIz7GeCrhv
lWaJi4dCGPxAEaGiX9WWMydj5mF9/dnS7oBLDZ8YM3Axe8JceRXESaHalaRMEHdpvA5vtJm2JUi8
RY7b24cwKFPSMCXFHlA4zhBokq4q1IZe4a4dF6O1lrJUcoH2j2FtC+fXa7s35V6m4g228CMMnr23
DQkWpo0hkXEukUbekSdCkfrBiznp08nn5D/JNie4P9d0YmD/0ombQHeemdNMnir7i38nTmjvmB0Q
pT1OjY/yXTi1Vw/UIQd6FBWNGxIB4c3vHa9aqfobgrRTMlnwJP2rs7/4/iySgKAtgS2Oc7rDGULH
HpLh4OB7Sj2vVetoiCxcqlB5DXgKiK2E00kJY5j5o20qafbJSnRgO/p+nGfNk/3m3rgd5Qwwr7vJ
TlJu+x6m5fKoXCm+5xfTuv5VjCvLnDrvnF2MpWv8wEJa8hGIRg9sx91ORcEkbmBTlfFHKJCnh4FU
R1cXsS3vMiG1l85EEzejHzaxPFuHQLbiabU0X7Y4Dqh02Qp3PDvf1Xyb01aTlOtEB/COKehWhVkY
H0sX//+5y4xfIpxaeL6Oma0h9hwfirqiCR4927ULeRBIKWPXnHc8iJWQ4hsbBN4ez/sP4t2i6vX5
/Sz4LlcU4Cns2pvv2jsIpT0FHLn2VjDD0uUWzPyKwjtX6N9Ad0nJpUnGHRhhwBjYQ3zPbgd158FS
+n76znMT9jnpa9Ve3XLTi9lKUj/SVeyq1bxwuffWJhYr93MpRRrSumV5DYUxFgpQOnAGVghp1h0C
6oWQ4dzvQgAAZFlb5WFXuqZeul4jvllty6iDsBb+vU0CuIZCouIzZPMNX5WM3KRp1xB7KY2y/uuV
sbXy1tAF8BuUp2OK7VrgRiHICz4Bsmtm836iBVfFjwVQLMNYRHa++3+ncUMrU3br8PdFc+Q+DqgE
XlzzkNMxYSgWNYlyuvqLbexVsoccm5+Tkp2U9qUQX/mp9G0pskqCEPIlsKljixAdBmAbbs/YmGWe
e1KIYoaDkRvC88P7xhGt/yMby/43Agg63q1vLulsBwa/lz/kDApM1UcorN5nNxSEHhhxeEu1io1w
5AzNHwjU7tWMFFzJVWiA54HxaR1hn9tbPMFfnjsHAUBsY/mTfwbVf3B6oaLbOGtiaPLIYJijIrwj
n1EzJACJigwc9S2N+xz7ywfQ2fbqcUqlDwAHW7beu55FYHphVOHpmXqPJ4TM03yXWNF12ltrpsHp
r2mfL9TL22cyVRMCUp7TR6SU6fDU9hW2PDhK6VZCPkR5RFIVPE+fQNNveKyhJJ0QsjecjP7kR2Da
7VqaL/4WiMYS+URxJgFsZQgQc6e9eZ5cgkLIQX3mNJmBsHq9eCebqqgWZG8NkuJbndRklUiCBTBH
9zHxzKXqkM2Hau8+zeFMuj+IJu+DRf2N2ihRVQA1tfNPkoqV3IKiF+p4RrzOMOFttS3Ezt+dlFLi
OIn+frAZ7H+MlSvgukmFaCWcxSb3NsTT2JR+fohxXv5RQKNWh6/Ilt0FU5uoEjyYCXiPyKJV1jMr
gc/zaOTzzy1bDX5QwnEjAAzBOp3rXFXQ0gFeu8RFlIxQIchye5/ecvFtfYZIH2mDL5Ynu+ss7zA9
7ggggbuvFnn9yTwZZXaKynXWWtzOdw6WNLPBp3UeBiJyww0JjB4dSo8i035X8H4KE0o1Vk0fOTIt
LmGDl9fjGCKqhuVU3Cop/S1LU/v6yqwzBT81mNPRNK2+TMlGj3W/nVP1bWoYuwSh8CyNndUkp9Bg
tvWQw5aOhPeqB/sBCTyquKMxgWa8bS3Dch5yYSzrQN82DGFVUMKZeZdDUFm+HwBRXblR90h3bxVj
0I8EB+JOaC7PJxs76q4epRj9HF43pnsWZvLiVb52EjFb9WoX/1mQLcOfhIrXc94oM5MYQ7GhDvGp
mTypMgy6J4Mc2IWXcTuldZxHmDqzIprMWF9fZtElG68cnJpUari6fd08YATPNpRzrnnjRPDV7yWl
6FNqgrkfnGwC6yNspAdw8ys8CBhzcQ9mBNp5/iXaObhmGKbdToTqE/IAV/FxCsozbitZ5eRFNBTg
+TMjedAbApO9tKbsOoaGupBAak2wE3A0udYpYt4MfADoWEygx/BTCL4czkyFUmBFhtgCYeC/91R0
N+3qOkb0WA8fsLOQHP4L5Wsu49CIg1pVkj0OAj3fLBnc2DWDkAubodEHpfKEb17S2NzLNheHyc/f
Cystko0KyTi7QIzS7PpulshbVxA7sIAZKzuHRyJp4wSwujajlGxkdQQDllfoAAYgQh4USQa/B4P4
VtnVO6J3UU/CY0MMn1gZxAwNpqHsdlHt0u62sKFc/4f72/LUZVWk3Bk8cqaEbqt2Hza+m4UCDQhT
6cDV2Zo0LM3CpO/atIuM1ajWL/yHs6Frhh45obTOYBQ8RtHj8HXScS83tHMSC7GuC8lRjxsmsKBC
lnESeAziMd2N9ylFM2WIU5GTlmy0Ci4O2S647V3mEMrVPJ7Ehjr/pH9HvfaQclSuaJnCAqo/sYQm
cRgwQGwDHMSBWShW0h51u/Y3gDXNz2wlLtLffHEgTLjfU1QfbcXXyApSKP5FIhJUk0QtREjrv8Wv
ERiu2tGtgJQlagbZg4iVU1PGYR57YLsU9vaoASZBqgJSwVYJRMG8QBGfM6M9slQXuiJpeVCX8Pcx
CtX/73uUiLW6UZROd+SZaLfV6PiQyqq72JO5hA6T3oShqIs+WT5flfNie0QWTvSbaYshZ5g9F4S2
9MmcTR90dUNI2eeiQSIwTVv+S2iJrwQj6YsGM02bnxSlEqhZw0tZ7DJzPoPiQAm5UdvNIEwYt774
/r8JfZ5x4gxRlNL0bAAIFVeehIDhNa8rRl+m/Pa4zmQ/jGLwmBqAGuOynScIBcLo5+wi5fK8NWi3
VdMfDlT7atrZFMyoToO+e+FcxCrd0l5u5Jh75WscpFro6+7fNYq13xGeH3qQaQM2DfIukwlGUmly
MuY2/NYuoFliQYI1wqd1iyr9MOqPq9OOQemQuIg6M6OCLH/JVS/TXGpQbZGFcXVhV9XLDt3gU7S5
rR7gukyVn762wcRtdAbk7p3qfe8pQwEWWk0di4UEkNo0B0gfVrP0syxg3iuKPqi9kQlTwSMLXfIu
eWTadKrbZrVEtdKYuQprFULka29MdKGmGg1i4ZrmaMetI+XuVvRGARtNIN1BgBEoIAl70RtnsuaZ
/a4nrOATGFb/JdI3EGv3aeABo3hzxKmgQWIkvp6UfiBNaz9Rmk76R14G0wrRx/B6VQKeQZGutiXe
9lqGvn8Yu5ud5PSV78/d5q7VzKBKiDHRQYNK6PuCoPijtw4lP8qE/9IAuodm5R1XaIqxyXko5eQC
ZTbrCRCAUKf5v4Nd7DbUynpK75iv2hW9EYr7JtRUOCZCD7UQ+ZCx87Fd2eTgKbqWGqm+OcOH+xeP
rWYQt/7COogYsyuoH1WFDrcCnilS1MuPC2SUNFo1lulJ74NMty7NcfTdOOXLNt5lXNE3NmBz9Mpa
b6jswkP9KWofadalOgv3AbttWOh+IZOZDLzEYGnbl2znYc6A2eDGAGiAvwuMJsCbDUfkO+1h463H
m7iH389ByKng8jgC9KWS6bXfDsrkPbMRyHlIw6A4CWcg7ssjKmwIBwKCE1bk5ZqdjK3QEvxLgD2E
t6Ngq4KBebVy5RFh38+SEhODfa63p0T21/99SIfWlb/1pHtiFiLMXK+KY/1hO0JxPP2RSsA3r6Q0
MAGWBfoB6YKXaqAv0qOoCgV3X1NkrzjF/ozxtqoCIJs7AoHEW1rNMLf7Uqqn0ODUnhYu7lGy5v+8
1dTQSmG9dFc+nF+Vfk8RV/cB/JQC/IuxY+AF1f/4LgBuaUJE3ZcE7s+kJp6YTGCAc/CNaWGdhsFB
BwTb41Hph5awxVTOH2/EWpeU5t5HdEraUBUxUVbe8TFz6PKeMZlIXZasD5iZDMYU12AAg1nislaY
AP6wGYhv1QYnDrtYLj/GNgh99N5uYcp+BKyiOMdHA5jExhKVCX3GCcgpkLj1fDQbknolomfTziFt
6KPxQ9E1dNxB2Ez8m3UXoLGJRsN7Qi+4iNtjSoMrwa8yGjP4zcIA8bhWkqV1hyc+8Q8NPeiQ793P
bLPhPTq+6+TeLI7mL0+Z8FSpfgqACTFw98dTPEp5erWgyqz6QYYB2ruuqEnSisaE7tNK/f/FPG9B
H/yQMIvMUD1qQMyTd9d8TaTS16NFNBWhz4GOi6LJ9GywbbO+aWObpSct3TlG+qCUihIB6cibQFce
kSvpOmUYpzCd5lfkfmoYA+dlmaoMg4G780L/TBJZMjh2o6pcpUN8UEgV1Eo6SMMShvhoqymzhDjM
JK+EZEdqvdDQjqxk7hwV74jkzzJwKrdIydNB28e3l9DepZ/ethnCmgU+ZjbWezrHnhwzVrzRDLvU
XY7WldqICKMK0za8Sps0k2vGOxcR5r4AoLA6xEPbhHi1Fjo6iLiS3cpbd2DP7YMJqJWSRJOwiuB9
jiV2rpelSry6AqnuKiOJY0lllsFNeVQ20OJRqw7U8s+I5LfpFj3eYDyorDw/CnbB00Ha7NfhtYFd
fqd7rr/iUI44l3cobJ1JHXaVtUiG/1q2w0UC8wUOBrjMQcWNFkdAs4X7MZHSH7pCXBkHwN6kzjD4
L8a9nWjOk6ssmGn6IFFWNMPEUZDd7DiPAHoDbBym93ZvNpBJK+hWlvZdlks79LnfGqcf8RlRzaJ4
IJYjBGcsvw8fGG7zH/NGwiomfQ7M9RBpAe4jb/C6XzYiquQfwV/zfQhNAO6gDfa5stbdZXKBU3Wy
VLhZ23g9seW+wuXtIxPbHmxg6Kl1Ryngz/7oVWzN0lhIeHTdgJVseZqCQ51SJmd6ic3+vPFH+LQL
7HpDpF/c3HVxWfkR0sycKYasfjgtY5poPE6sAcBDQDZlITKVpy4RMDdPzaCGZ6G65ecCCZsMXned
sV+cpQgtyz1lDJD1DoFZyXrd6nJmobTHnJXEvJ3xspET2+d5JRM+/FX0pZKvh2J7DbKFZ3P7shyF
pYCX9qAHtaByUb6zEWRzIFZsgIWyIrJkBYQX2rIMnL9LYA0tZN3Ac0I3IjyOzB7YSrCzUbyYRYKi
uduwx0YhZy5u4aloHOJ6TKaaBpTtuVwHL3bHK4GI2Z3goa1xrk/T9RTc2rsDUnTUdqQZNA6e49YV
0tGKXSD3zr1vCGTaZcmcym0WOJN3JvQwLgBR82XRjUMzC4rnS6f3ZXL3hpYQdN2oboIyOgfnCEWV
GD4SNcbSHmX6pcoUCRAH3bH83dCGdbeYS6FGNTyJIZImxoh6tjdiPWKAsjxohHwJ8cLJHpMfsilY
iFbB7N1Kxj2b8tlG2U3SQBeEbF736qHhiONkYuFHAr1m/l4nbMaQsILl9ZXGQ5hAlr3XHN77ue8U
jKBfL09IOAIHAruBh7gVhu6gvAmb0lAD2Wct6LH4xW52nOhq0ZUbmHGjBzZXw88KXmfEqFVvBHsA
E1hx4QErWuy2rfuktKZBvYNHNB/OLY3JojHshfS3c1hfr0k/AvBizQLz+Ale64BYlfG6o2cHHndc
lzBjLh8Us165GFGHUuuBFQXz+CnIBBY3/PGnatiJjujo3qLFfSN3U5HFylORVwu+HdLXDLRrA2Hc
yKBg7S66EFFUR3Wojf44gXg+j6OYTr+clRmDMKQh5FW+j0fNaE3GVg/v1Q78BsBS84KO/l7Cg4gY
z2r0a/mjJlZW7qbI+IPDT418HCytQhcYg6qUwN1B+24izCDYEvfflndU0cXTus7t170XMT5z7aEW
noy2LVEMNKsMCcbaiSye9GCxS8x+BpdltPRgbdftkqQln5OZ4nioU4kCbwsksw8H6s5qsZMJvEzy
lP8v45nIgGIjXNEYRNONXUHGtMRf0PZgE4dsXvOc5iGer4zc2Gico0OyWfJhwnd3ass2cOcT673Y
notc4yAQY1v3UDhH2yWu4y304mW/1FwbAsd10TVUTeTJK8vyWzoK2ik6lQq/Rha5ViSX93TVzw24
enpHUvqUOOuiHGgPDGBOFj/FVkz4jPhuNymFIZTVP13sGi6OGodH5Uu8TxI1D4S2xLVAWxyXtvfc
IHBNImfma0caVr0E0JD1i1FT19XO/LgVBAJSdd83YchmUMgNqDaW/psghlGTF+kMuxsvu+NkLe5a
/Bk87JJe6b5hwVYvnyaQ+7IC6eu4kQcU3nk9N+xMAfDqTH7M016Dj7U8gvIEDinzDSijqLuDwJ9o
u0kqzBdvOZATIx6pV7U8qDwNmIAIBb2D4RgVLgTO21C/pCAkHF4E+5mjiPO1tU7IGrz8Vk842EdI
vK3ygOj/rfH48YrLusOirriRTt3dEp4guo8Yovz06Np28uNlGCYfkRS2shMPbK293qzKRRvzh1Nv
/Xu2RlqQA+YI4PRjrNOTagY6v1w8Gwlezu0IDQIhCk/ZnVuAJx1bqN3vHM3vcTbRIKEY5rtw+k3J
udkYnutNyKnGX+p4v8uuUfAmza+zMYBCwUEjXm7THj8rk/kHlrC9U3wU2pAfm+2kp/wrTBT2d2F9
uT/73R0zNHmko36lotjymGgHw78BjsDWZGxiZrRDg0sOP9Nww3GLP8U3tH2nh1013yfilC9hFbSY
mA5/TDT145xw4Nq/JFlsmCenHN6MtCHYsS3yIPBc8shQC+Gi10jioj8pNFOXVvvqTPn/L3BLJW1/
w8LUk3SjPyly7ZgLnKLGaqb8tGdkuh25iHmWWJYti8l3DZYJA8K/d75PZc/kwfMQcpZYpDwYUhhl
NddG66bGEJkts0KGcGNQjSIA1ahWK9X8ZHmH9tgBkFMpjzWJTRy0smyW+0VTJig1El+JXExdWOWW
lDlKcIjui5uGwPoxFdTekO1jX1nuGV5EIO5aYMddZD/S5j+hyoAmHfE63su++GhUNkuke42T0U8Q
5ypnPgV9Vzw/s+VGOYlzseqk4o7duK8DcyHD6voFfdiCeUAoh6s+SJwXJab9+7COInTDiGW3mSUf
gKYOw57VdZqe65PjM2HPQ69ASUqaZcZqqNmMr8HhYrPryfGhM8HWjmMzV38LHW98RX9AZ3Ulz2dn
kJGPHDgNqCgdsZ9oJGnslXWd7gidmzZAvNCKXRS//HEr3YwSY5GR7+YImz5NK3VjJqixkNQ0PVWW
VaT20yq4TXjlt6jZNhRXxvPB8Nrxs79q7k1pz8M68EFUSTO0nid2mTfCzb04b5sB9YruxCGSgDcB
Le1HCaKq8v42eZE3qHgtXl9vPKJfYswtgta/pvrKHhrGPmXYz6KxggQUud/aTeQB3CPtR0yECD1y
1q1P5bL1HyCvkiQRA08sSHXJxvFM/IdunocrfsjVb2yZFnArNRajXD3V//WBMZJU2TTmVut5J08D
YtFa322m1nC3upU6BAUh8BuTDtZK6wG5ysKaL2rzflWPeVQFOtxBLYWnOoBEABtNbpX4AIP+V0eU
fyDm6hjopnN8k0ejxhf26/7jtZBsvvurcfGTbKcEEEhBKo95jhygTRqW0LlOHl8JbkWwohRFtAJf
431QMIsaOaWRr6QrPKjFiVJjRWxqmjI7fk48cfNvKaQxQYQcieBStAcq9UkST1epKqbiprJN/2N0
RQf8DAABI3F4ttl5yh93UO9bGA4wsX5jULDI/IDH5mgEJShfBLANNpqrnnBB3zrTKampvuyKQQfX
M6saP88CatxrslP/r0QuhH/B8oQKz6YHKCKABBlYuvvssO8Ul+iVOsNruDcOLYsrwGGEi76tpaRG
ZgTDrN/rHpVwYDoEbMK3eDI/eTJ8lEw7R8+m4Fzv0SA1M+KY/r3Ty7irMqYBZsioEN58CBdfMv/W
TVeaS0or/MfkUayybuBpSc/gb+fFkyBdzQqFWPETZeU8nZwWrCwvQfwU5a/YryHBZuGvLASP2MYl
vMuudk1M8DORqf0nIOOpjXeOgKVll5JwmOHhREGjH7gtomIiSAGbm+6cqD/xOFxOhZpMIGb4ls8N
43plMQ5jc6AUE2uOY0hfXsMpvhCV3NpH1hRe+vs3ceDOJpuogFBTjXuMDxVXbAoaAC7j+Ah92Irb
CnEAU0Eo0jpeD8HkA2qSjAOeBpPATukjN8hqVzP4FGByrMDirGHk9zjDgwc9gAX/nF2WtnWDOK01
c27bRZ8r3rBhwO+R23y0r3zsQovLIzA/MZJLF6wrWsrU+pevNRaC0jkHmrQeo4rt0wbojAwwTjAl
a4qOSsmRvlntufjDu6zfio2czLTIO/moY/h+6J0idDUaynyEf8QxcCYQ9yzHZROI/hMa6+6ADIyw
veqncVeqNMmmWTcCBqUw3KB48NDc88OZtFBuxmVOnml/10QynaKiWLILfAUN33zzqyxcuRKO4Beh
eBjbYSN8EjHvJkYKRXk3HAjSWc52egKvMT4DEFOMJytoaGU24KLa47uG1695D20fjg5uZPzbY/Qv
mF2F/te8FRViU5WhYWZB4b57rsx1PpJlTnnMcMXRlMJ8OArHLRsMmb7LTqihMSvS0zU70UuIoPv+
bigPCsrwGohqYZCXW6JtsMVzWtrF4+nMBk9RqTEVwQljbAGTfinwGEbHS5YzOL3F2QRj6MfQz+Qv
I0tNDDyIR9jJh76YhRnqg0ZmtCtBfXy/lZqeSmIMsIVpSgTENRDVyTL3lCfg/zNgGphmyqyebKZg
lDCCtiji/+nczZSNCm+WHt7z/xw/WscWDJkwnvC1JbDu5MVMP9sI1+T4RHiFOE5j9UePWG/agAot
xwkMkgWzY8vZn1H2e1ErfauSiZZZZZg9tRx3Rgx7mri2NjgJjdBApsWyPV+hi2nRh5wwSiWaPZ+X
XfWYYh2IsnUXdwzulnYpC0iUttwhwX3I0IEc+EKverjkVfGkrSnV/gpetzvVk6M80qNUxFgfp3f0
AiI+WbOa65v6LWoxwXNV/3dmkGjkWNT048fzaF17K+XWKb6XFxAdSubl4VMEdiORavELiP0fcr6p
apFwFYYmvqJe6glogos5iRXPQHYcP83xdxn6jEz9CJk+CnSNSyf2fG7/m3Zmd4zsNm8BT2NiGDJQ
OQN6h3+qXwJt6EkF2EQZb2+IzfhEv5eLFE6o12i2lifvn9o0gb8tD5GKX9Sxqav4CCSrWglKakfK
MEIS76vhZTc5/lxhKlATez3LrDvCiZ8Mt1tNAg5sp57yW1irBDrr/Grk3SB/hHYcXZzW6BIBVXLT
M9z6pXpqjnJltQcFatOOaR+zQL39tzYh9tiHEsPgo59fdcnbz8GxacrlGJcDJvCIwwIf5DC4af63
U2xOU7Y5ZR4cpyf8S5aRqjgyxqlVoox+RPsRTxMRaGMw+28sBwGtChsUcRQ44j+tY9q6PaDeEXxw
tIuOQclg+YGDz+QP68TIRSSQKwBC9l8kcJIjezzXzDq3PV2jmgpg/bOH5I3DZznH6IV+mAlB7gay
wfp3Ugua7oT0QErr0+CqPgcxq1ZHY4wQ+VJzffjzFMSIhufyvftbvbc2KM62rB+hov1tQsc/twmQ
XNdGxmIfCT6yc+oPrH0ggn+3bsxADIyZsh756RC2GWamOs7VbpT0/o8NLLtu2bo5/qChHLYmQO0c
0vLCVUWsHAh57+AGLRTe2If2pBCKtWKAQ4NzDqh0jXo7gzjJqxEYG7Swz6NM/zc7Sxr/0p6RqodV
UMhUD01MlujLl7/pJ6YaOqXvzlb8X4quv87sGAW/mGIMZNu5XdIHxWdA8Ip+nk12dMw3FswjE5ZO
tZQ6490pOFOnCGlB2tNEpxq33kqoqoK5muA4HbrNzxU9fzdj3MoUBYpwExomN1oIDrTuLFbr4wtO
BMAJm3JHYJfy1XtO5O0DGsTILUOlFBXh4wev2svmIlULJadZygpVpBezYC9OvVksH9FuxZTLAYBV
6LcQBUqSMjfYuOfhwqiLbJYAhHukHeKXRJsfvZqPMGQbBlQxHgTfth5PXpkUXZBGMSZdhag19c7F
6rCjyG6jZjsVsO0YkamvK2dAFyTNewujjWqks+Xb+hxXQfh99PxXI1wTrYjDBOcrDalkknbbdB2U
1f6RQG+4SXkP/Njd8DRoqVabXhSdC+YV+9/Bo4iFVofrKc2rBlJvZX54B+RclENPvV9Sm6GxdhLH
HPbCmbAuMnJIPFKztJEjzUvPOQPJ6VEAIMaVxJpg8v8ezrLeoSVy9bAy1vYmuSvw0K9m5X7NguUi
4lo5DfO6qmF1mt0secbapxULhz15LcFRb0tpJAPDqWhPGNLqB7E4BfyyWJqiKMa0f855OqF3tNRM
qMyrLVxZvwj62jULMiqHuO7Cih846dxnb73XWp3R1ClWm3lFz0ZneWsOah4LLTBLkfzRMnnsCIMT
Kh2hdg0w/5+lByWygdLnotBOhCPaIR+rw3KAlAjr7R9zbnp1wj+C8RzytzQKn1YI/9HAnUPIXZAb
H//nR4RzIa8RWZn4JWLu3W6kAcufo6jC0RkTf8tKcKkII1yjr0CfUWiiDIvDJw/yJF6WRxnxyW4c
U23mCE2NLSZn4E34cVOK96Y8vE6HRMqPbznEVlkKci5oSIIuEwLIn+BpWeAYmZqpX7pH0gcINx4j
A6eJ6cKcmZqOnK+6uHgSEvPWQlPDcMroC/J2WZVYBGtFxRvX4bCQanXfQ+W96xUOJlx1zJiRNAWb
pJ+qhVfk/0aEzyNDZNeGEctVvAhiZhcPRLdPaNpV0TlyCR9xhPzOSTisSj31k7x4zJIkZKLCkh+J
eiNPHQxC4JOcz3f6tjnKysRDBty4BXf40xpRf3Bt4/TMHRdN8p3+YGUNl4oF+ucUZmvFJ8bKWnEO
hH9J7SqeoQM/WjoMUiuknhQBvhs5J6BrnTS7TBjAAPit1fXJ51J4BYgpSGbc/JuJnDafy9ABP0KZ
H0xXXzoU1CNBoPKEoKE1WwpQ2ezlpKnsNYPP4W0i9++36m0GcpQtQ5JWBF9A3jOkPLuGTHxoo20H
XiGPvoJrtwdd3mGbHJbtVr6kxWD7QVeXLq1sbx9zqaxbHne925J85aGV2P/QwcxACh2+2FjBUOuQ
mVQ94H0s7Pt6hhvTiM/ZjLyTVCx/McFClbkcOXQA/O9YaJyVGnPMVtX3ZgGiceWzB8NpWDr4eByT
cTT1/+fuh3yFzFQk5LaLEFpf4jSoQeUTi13p0/3BYnEr4MdZunRdW5/elKYQloM64g0+ITVJmfis
JEFCG6f0XzDdVDdC60dbr1CJLXrlwRTvb87e8OdikuBkoqg/G7UH32Lgm6XB8gpA8URafvZX0Lo0
YYCMQla437JTixgO/y1qg6Qz41gm9PD/kg0uxPYpW4OHy6ACixgHn9LoX3ng/btsDKFk37mf9Ao4
PyxLkhxOpBPYo55Ik6lausO2cgsEyb1UfEm+86vJ8X8xvCTtmO0pLxos91hydCQGE4rmq4ZgqPBS
r2GCPmePa1vYvVFCbIAgyqrXCOV7WSlcEppxZIhDvuaLqtDZFHREsNcnu8yEz9j4APJHdKZ7EA45
6IjBgMi4Ii4VInA5A4NNJRY4eb2qqc1QgdO0ChtYZO0aHoLSil4Fjfzg6Reg0ypLeA3Mu69Iojgc
rPY9Bu/s22Y7FvS8jNMDXGFVAtVi/QvhhpciFT7I/EwWtyoMeojBJdRpcvLrqmNjwaMR++BK5f7h
Roxt6s/W4URFKath65XiL385QsO9U03ilGczGh3GMcvwpG6xU30jVZJ1CbEABoTEPsIuNoAuTiRV
7cvOFPqNOJczd2cn5rxWPW9c+UuVaWvNtCsWIBo3Cz/Vwenrh7/8evx6oCREo1RG0dUiurCxfUOB
Yu3FTpafJ6UhxLHrXrFQDcQ1F6F7r8NDb5TJo2d33eh3c6+X+0ISl5pZ9tAQlnFeikhS2b/ZXxjK
1lenlPnZEpvq+SmQuixwWGIForZ/xCcgC8qF32ScJCbuQWkjx6CpZYYj0+tqETk/hhnJS8p/nduw
hlNtpt7y6KTXoj/MOZXxDlUr7T4lgOkWfffdTV5zca6vp7hqylPlcOaVSNGGHE+WO1w7AYOHKmtb
Bo7MXJSw4nHsZB/tES7D6Qs9TMLkkO/2ZbruJF7YNTjwYdtT+fs2bWShWsjKO7aVh4CK53lIv0BX
sjMiw9wB390BTLtlxhG37xnfDqGqjZJj83nawFhK175fwNz0TsY/jX9bhAQYgR/a6y5PPAEzjjRM
Jd+W3yor2KpF/quqHNdaML46yiyo5lrgoxA5lmbXwLj8J1/3jW5C/c274YWBTUvBJjwM2vVOOa3M
3xRjUcM0IqC/vcKRrWzo597b8ae2J08nPUIl0xv5Pmg/BghGXsbaCX9SlhAB8gnSL+KXMuIONL42
U6l+rOPAqqcSHAimClfTCg8PoDl2gmqd3Vu8NNmfIpOxl+1RwxlrNYIFx2wh4T1WySTiRzqLL8AP
z6GlwBA22PcHLf5nWn53O0QgEsu+loO5PI5iI8q6y1CJL2bJi7KoXeK4PxWjFSTsbdh14maJ9Fuc
uHfw3z+CqtS011EZSVBy0PxHZ2Qku4juZV83OdLrVgIBazK+lJlfsMcypAT9T9FqMW7Q68DpHJFb
1TvkFV3/SsEbzG3dtAQeDSJvHIZ78D0/wGX0BVeZKGpFKEOMHRxXAGxskpEtYMuK5Sjd7tjCiR2j
9xNwLOL0+lpT4rSXQcrN1YMbWYZ8QMNR6YhC9d7P2yUP7rx0A45RT4TRAwiu6/LsKs1BExa4YY11
ESv/dXMZ5toG+NJ9i0SAiBjVPbOOHOrmwt8BFGswUqcEO/SeHYclxaUi6QY1/lS0/JyWgcXOLY7n
2a++u9kFh/rUBZD5TXjTJ3K1JhmIf4ERRMpYt1ZYaIefCglu21sLGQ9n1u/ktKRAXYCSikaNPyBx
IXM2gf7E+0m/OiliBKDrdo44ImX7w6Zn4Pw8v0FQrKzA+twk7YT26xg8lpejaAUIyQ+d1fyrfQEM
rI51Z2vb/CgxzW1SB2QFwq7VtVtZt/eKuAla+q7oVD4hVl4Vl1rLNQ/F6QaXZa+hhIbcDXu4dDfb
8TU/J0wA1JDgYhC2xY8dvfl4hoKEWWbbHPYE1oISHEQJoCOt8aOaIQaBHajh1yFCOn2hxNkYwPlN
1+aWLr4ps/T97BAMQtrpfM0HrN0xehodHJPx5RdzdSXbSiE3O19EyBFUewOzhpIAplDn/6DsvGnI
lBShvgkPCOVQuDmXXuTaXZtKScICg+HVj9H7XnvUMHPPcwIBGUHxtAsZEjTwwC8KFDhJutfFxNLu
G8sxfVwYj/EpiWO+69gjV5XduF3YjY3TGGsRz5V2o2mOKzIUmqbq6wyjqTDCFiO5miugDZUqJS5W
yS1JLwqV0EDmeHQlYJvArUzre38G74Oyy2E4NfFI5ZsZ8XD/AROvBfmqwFgcfZ5mkB3AZ39sY8ZJ
LNTI6SFI+OkEJpCHwdtoyMwA61+PtlRkgNGs3F1fQRTG4JbmxbaFIt0M7hVnj6W65yhKVYrDCBV2
PuyqouUDtnAdmFn+Z3N6WcjfKjkpAXXavON/Ko/9uQ4A62WkgzHjxQZxGE9uBa/Xylc8Vfxojsfi
+51yVyeXS06huZzuuq2FclswJ2DZdJfkloRMTRL1fdDKgW/22ZalCgQL6b6zUdqtK1MWRic8ViTv
HHpP75FnNNgjfaKRwa3FwtdCLgcj0u9FUS15kZBrIHDnnb0abBhtqM6LOGBJcSTsbEZyV8QNcLB7
LSO3Ds1hw1dVV4m8x/k58o9pidatjBMvqT+p/EdW2ueOx7NXLoUJ8EZXyhryI6DDdClLPQ75zFWk
C3UCK1dcY26OLMbQrdU07q2AtrXotv8ytH7wAyY5J4xFt2r/hOUWIxzpcw6bCrgraw7dv/F3H20i
jcgLPL9VPgBR4ED7nH37z+HbbrHEiFxgrYfBSKMNm894uzVaPBOqDRIYnF7FGO3qG7mKhovaEArb
FZMPIBTsdAMO0o9ZEXmlz1DJUNjj2AoAZ0aAChVM5WQVloTAKJT8GrT/UGX7TXvUKQP1812LUFYM
3XpDgItBDdf1hjmygX1w664YKX7w+0/SXOE8i3EEBYp6z6TaJSjNPSBiksG+ADBrxWnS2wDvz7vD
YZXXXM9EtxoHgT/wW5I4G5g+bND9kqUS4u8kiZQ+IkpsyBsX2PhXsN8YskVGYzYCmiivA4iDbPML
e3VEeNWJntyh9XxsPBw4QG8IDDYSVvc/KUm51bTHyKAGAdL9H64jJQiSBwyhla6Rbopd/19oU4cJ
LqKET9wSXMgU/DutmMr2BD2G0ZmhntnlxKWeko31oU8QwI33u/ORrXG3OSs9HjbVqMPtT94IU39B
owiZKSDxaz67DRTE49FzycDOq+YVEHjzmbD2b/3FYxKiio/ovsrepkZo7y222g840EPN15I7Zy3t
L/lBS5diiWylj1u5FGfsKipCzVd0g1vyzyLD7T2ro8yaS4WMmkE4hNu/+yjbtlHAaosaDxOZcFeS
B/zmFtSxYLFfx7XrfClpP4iJ1X6zBO2hkCd0/ihbSc9pmIZ6+y/HnR/+q2EPCmbptag5kPe/2s1x
jyTXoACipBtd0V8euwQW5Ylqxs8uFRaVET3DdTGMw2al+Wbe5lg7iTDiCmSHsEZU3Siba+T0d9BK
Pp1Aomuy7jXRjBgJ8Nyc3gWmYSqvMEow6utrV2vv0mt5cog+ikYJISBuv2owCToVdp+OBoRIKLMx
LgX+wuCc0wQBrD1aqkXk6whQRkhzn05GilXYMq/3tfJpplia+PYzqDBUlaLefh3nKwwdfgY5Xtg3
PGOWbrpuB9T28rsoxQ6WlK6An4S5UlNs/EP1sHNFZDhcQvViWCj08tIvXEeEy97RkE9yXIVUgCFf
30cnLT7Al3OJGbqK/Mz7RnG29mmKgRuNri2AaRTyJ2rLYfr0Ur1HM1/TTcW89nugdvP0nzLeFmWV
kHjKwzf9NlBnl2LwBF3FDlymcvR8JPxE3a3/4kE/gR6yVrM47nSHtkoVtjfo5ZqTjxOB22CFi5CS
KXjujeZvqOJ8kC29w0SmxjQLLyIJqB/JytH9uub15iL3LumvC8W95AC5e+VUK1vxm2arWfjsHDnr
nzRPwSr9oWjntdjXQ+rBRW0Q9CxfpbTFjo5g5bLNuiTl5Z0OcUIkzyOWVcSoWSSZgJwV/scnHBR8
JgyKdDRIljAfGz9qJ3BQQzRG6sedAim+PJN8JZgQ/8uRq0VJeRtAMH7Jdu8eqJGqBoCFDWhCR/0e
KwLYUCrYAbr2bDCKl8mknIkUyP6dVH1y5nfe0iWsihtUrhE/pFrqyL+WsfCT6ezb8s9qmYxCO+lj
6gkxfhOz/oRnNpDNExyym5waB1Bbi+/3YLTZ/ZbUZPR9bQ21g/hTeeeDPkoWPXcO3rnOUyYZOBoC
y0+gcommEnEQqTJiZ0igT23WSTWQfLeWrcoWQcPw0ZHfSghPIKxaFjfxGXmswEOWEcrHGDv2NsyC
fQPhJNU6l5+baNd1iwreHRXmArwHKWCuqOPRfcalp5aE2qsVGZHlc3KqJ4ulIIotoo8P3VqRIoKz
LCf3f1kfGCinlbXsERhNHUg+tAh3WCvCbxp89VYU9/nQL2ODTikEIVriiiDsjk36cbl1GZaj28cB
aUhsDPBgoABKTf9FKc9+pC7HINRqhSYuLvu4uOUnMJGrJQ9yk2HbqszdIteeCfgV1P7FrxjqFPWM
1+zXk2S84it44eZLgGUcp/Kgz842nm2iWg09LLgcPdr5CSsvYNl1rBYXnofF9E7brPdctwlikXrK
IVR9+A00rfIYYv3S38P5B5U8WkHO2HMr0OLM7etLvtGtWTuv8UkTn1EX/iHOpS5I2v4VzptQQcva
YnQHro4QmMqbXzHPY6tsUe7bTEO+cd4P2TzwfzZ9fJn/FquDSOSnA5nSHd/slC51lt2fFRUk50vL
wObNxztTS/KpZe+FX2nneIMAGpTXO/HX2nMg46YOBMWaUC2dMN4fVk7dRMHH8FrayAAIJTqpaRUh
Hp44aijGwYaTBGrSSKxLItYuQTKTGG71jd+YTvcMFYQocLnmsQoS0onjymOrjmKFX0oAGkd6CQQ2
UFYrc4tQGR4cYG07aG/j5wTvc8HHlsTpY27rlOhUmiuHbX712RBoiKQG7i0CndsWIWgTtlZ4hQf3
T60F3sC5h5RJzUok66B2jSBBRkioXeFp60yORhvSqdoW0xCGVRwKoBJhmIszLmP4jqKk8HBUfIDJ
QlT4K3uD1I9H+iTkgKgFa4Y2C0ENgzszi9qXObhNH5cD1m9NTFRB5j3wQpgtFla740Wq3WGvJjQx
uRLTBtyHBBW2R6gTATriRw/sK3R10Jq+F4rMbkEqK7Jlx4GPQgWGiYGt27VvWjoZ8cBgP5usZ2D0
rnhzf99YGJNi6JhHebFTQ3uxV1CnoBo9SOAZx91DBDkZhFKDWc5yztQf36gCFFYNJ0Vcj7Z8GV9T
TKrak9tym4ija6Og6IlHAmIHaYTREBpKU+LE4pyUVnQCeUAjXN4R028KT0x+OrDjPtiQvoer5IGl
BDf/yGzT5k4r9asG1xS4ExqOvCTIQxRy6uCX1zgP8uydHERng8VT4ZCRp2Y1VpbCwna4nc1FCeR2
YMs3P5zPTT97VDNW+MB9qFRdNqQdsTvmoy3yropgl2uWCztavEkbI9XTE4OO/TPnVoJ2GfCAY99B
4HVVFt6SkLygHk/DQhFt3qgL2A4eFC6eQBCfCqcKaM1LFxBxkkzXwUdAYoilofeVDR+II+M1Xfuf
vRWCkzAfLliHCloANrKDIgxUuh00BUFmDiOflbbHTfG9rdIiahNO2cTea5C9H5sHLHxUG6BVe/Su
e95qGcPMdmvlrwt14ddih6A5teySl/Lw7D2Glzt1ERJAAGcwvs6a6aXMbsVuUKwPXu6q0D1mLZ4S
MR+QxND6BH1BkSRhwmsSWYWPMU2wqx2La3ozHnoqDU7vSoIxKESukVy7ZBC0FCm6K305FOs+crGk
yiAAU/0NQjQknfbvdS42Are++yh59+laHi7wd7DBnaURPKWSyewJyJSoY7HGoim+mZX1fpbXPNs+
lSlIZsU2IkmZanCf23I/YITTH80qL05HRyjEGE3FdYdSm6rIjFMRZlKXSfDFxogbFRv0ATyZjKeI
0Vz3xHIXoQuzE2AXGMpwij6zUa825iP87J0Rk64xF6v2d1MArBmEdeIahoOmbC49RO9X3l3MAbM6
IDM/h7xulSbotkzI6/eVFK9YDbPvuxOK34pNv8DX5GmI6OUs9wJpG73fIhHQi7a+5vrLjoAhiVrd
J6hRxPMtSccl0MKKxVkQi8xOUp1RGsZq/u4ac5cWBbQsNmKzmJp4Mp2xOYnRLQDVsyxljN5FCGpe
okM1pZadb1r0LvNN0brus7P2I0cW2x/wdRJ1bF68ZMrAWlI27pTJZs6NNBKpyGgtL//Eh1Ie87nU
nff7xp9v8WOGJemoz/RNoIfOUFHBgP7fAF12HGR/HtGkLh0CdGED6xnSb2vJcdW3btl7nxa0E0Hu
KbjxQ6a3dPHakUcprOOwT4kHxM0ipu4Z26iaequt2f4EnJ6OBnxKW+pENUkBwXG0/0tT9pFc/dFH
QD/Xr9XVe/7sSZywJbHQR8cIOlMLo/ZmpjvCSHk8QGuAj6GQEoGJiSfq8oARTOhFfalLSPt5xEVB
JfKKw2sskxB4zi46ygAD0pq/TdJFt2oSR6+uXUp5JEpl2efiuMtgnIoaCCV68/GCnHn81v1fh3DW
hzKYc3mLS707DV+N7BbRqs16mxoYcwaXmGvhN3zwblSnTcJKOjR/+ruimMSjYgneW/papqjOOJ1i
mhFDIN2Vm9MoC6ERGSUzyDmRGs3r+jhoh7WP/XXq/WlehU9am0bbZg+xKRUAucQ5gEb4BbwtFTA/
Y9gpyPwkFYEjHl/Q796rexQOOfLjJM6j88Utq+5GoFNq+UtDjTUqT7UBe4k6bvA63tKjbnGZMu0K
HvIqSQMcenOLQV53rpeuZgSOtu8WixIK1PhYX6Y+a4wMotluNOHFDUGE2BWOVDHnhezKqPrjrihH
gVlGJm5qUtZrra+oLdhnvHOYbsrZAEvgDYXfOol2Z3YfVnJeZY3a0qlI3VUfQ0TPnfqYUNpjQJeb
PyjbBJFV9wDk7ERSB4c8+VIwxfocSkUgfVmXiwwm64UIxxYem2wibl2nlln1yvHIvzmNEkPoIwe5
/SfF7M4K3nZ/6GRuqewuaUdThhgVBo/Dpdn0dUHcVqedIeWZqrBkLX4SDBdEqIc8BCCicrNbKJeU
gwUQbntOhOPZPuFMXoKCgwnTjZEJ/othMWfMk4yF84xoyN650hRyf/uTbZGZVvmpsvx0ZmEauyXr
AIaT82m9StRV6LzelZpkNi35HCrhL8ddi97VDb/FCvYknGJ2gXs58ZSwPY80TImi4nzmlOWgzYHN
C2+h5eyBmFOUjYRdjTkKrVEkdgXQ11CHjpK0z+rfTtYWo+9C/NbnpY0YOEvL5zHCfaEQJVLfE89H
dGhz0wJmph9clMBFpYrCTZh51tSENr1d+MDzgBP3uzy4Jzgp78iAbhKrLNAEXDExMN1xn16KRWsc
ZC1nZCJ9569OxEGugUhlpftXKniYoaLh7TzOCplowG8STa+ztOTpJMhg4IvAPLi5tzygYos1KbGE
BLU2pbrcsCBh2qoqppfzMkc5hSWN0TfZJuFWF68+ReEJi06TQVkVU+gVg4Uzsedix/ruLjPui/Ui
X8cBZGqPHtF+VNRetCYRWr7YhMsXnO6eFGy9c+6rlYrk01avOPvC+3DTJ1trR7GCmELSL1oXSN3/
xsWqp9mVJAGWPImuAUCuCcug8bUHCdn6uhOVG3HBZQfpR7hOK9+eccf/pTer+CPbedM6Zxzb4Rr5
bYNnNhtXCSVclfsKQLazz9liFIQPsSdB8wrhwopkNeMcx/jJNs2wZixiy23/Qg7AMKERGiZQ/bjf
uH8uigp9JCf/Zmblv8fKJlraIF+Yt5F7mCROCzSqKhVJHWTv4igbRPIMai13ppuKRzCBzYOvLo1J
y2NZnnpa2HjCBsg5UUhZipzkBNgpLdOC58sJYwDS0rf1kOaXpGjRB4Z6DfVOxbDjvgHx4k9hV/Iq
cOVRQ39eSSUgHm0MAEukv9mW+4hWrqGtz0LT+JpnafcJjXqaxK12w6zaY8XxpBhP95le3sjPdanA
ksfL17Vcw9zk1aViapU/aAjDnX8JRnGMBHMZhxLuNSmXi0dinVV0BVYvFxMaSHVMfofuIoFEB1Ej
er71D1dpm7mTeMDKT5GSeUVTAv12xNJ4t9IppjX9H2KKJxJH9Ni4UpKuQqOFfb/FTbmPbwEXS9yV
IiochdvujTjq1PoiB+NAznTOqsdROfHCjbupaCeSA9B3HD8Apnhn3PhPaqqIu8q9li12/NEJC0eL
JzJlr3j9YV7T1y4/srN8Fhlold2lTKjMt/1WunQpSNpex3LcqRjb01JeCBC2Rn04PltPNaB3X4Wf
vogYIBvzG2Jc0zy9XSIqfIuwxhwN0BT69QkQyuoyM7xKx9lcNlvIGgjlTnLzechkDPP+QJbzmSRS
gi2jgBcw54gNI+h6yaZR/rCv4rlw4xRbst3/v6c0kKOcE9Bz9tnaCvlEez3zL3yZyCgWNlPU+IFO
CyH8NA320WJelBEeLo4SOtUhD1SYp6z0HalLqrB1hH3VZB6kMG2px6NkiAed8C/SXphK7G65K+5Q
72McytwyVqWEoF46BT8olocWg3XJq3kbOA4ergyJhMqkv54f5sivQ4LCDoiLRJA/saimIbnM9UFk
aNi3UNkewvzs/3T/KJsNqQtE5Ybyf2Gi9Jo3hw6FMO+GCdqKvG2JZY5tbq1BC+LkRsxtZOjn0j6+
zXy2il+HY7i5SfFpCxwmECtbvuFMH3+SUKM1f5Yak+hNHygxpeaJcEcQABDE8NnguAfIPaXZcDLK
B+AcZlr3pIvYJ7v+lrVbWIhEGKPi3xRzgG8LvQ4kpCo4Bi//L752BtgjFOI/GNGPelKJBn+u/Hkh
A6aiKgpEZ409YyQkNJFP+t55ZVE9PGiJzXlexFauvQGMbjcdeWVHJhWycvzqpMrcqn6kHl5Y59eY
q0CK9Rav0eiTgvnUxl3STNZywlmbZ9UeFbfYY9nKnrjPavDalbBeIYCI8bSJplYx27LqhrpMSM2C
QDEuCD6uSp5tNn6BJkAnNxi0VA8Ihpru0t7PVh/Ht693InT7MFji+gZ/+eZ4k+NzSG0ZIaTtLrHN
VYk47ix6dJ31NYjLjo6e8cyG+DwTm2Lkz71bivjb7ryb8IxLWBhqrhWnSW5Q6ppFh9j7YJqL2N00
66c2ktPqBX9Wt/bf3VySig/JcibU/YlHLJ+x+hKZ58d3RJv+orFUl6FStYMLklhgbKwjcnzF2C+L
ElymSskYyozlRipNMvcNSnWGeOaBUuyO/1b/T2M69gx+1lkjTez8GOu+A6RDQY/xjveumQ5iMb8w
lX6b59NzJXULf61tT+3cPtQyRP6wvJ0jCM4d3ooMBZVm83RgwMRLfh9qj4M62GYFjaX7HNyj+zYD
Fpwikl7tAyTbptOxv9aO0rYYfPi1UAh0XVR76UacXI0Bb+pewu6TYGU37KWKXy1kAOjFFi7QJwnz
xxb5FMhTFTLrKAiJRboz3L1ff/Swztj2pqI4uKnDW1MSKgI7myvMu+IHP0YbZGiOfqMzJAp+TXX6
xuXFI7BB8TaMyj+JQcKoZ5aH/OP+mIFu6KlKm/+IIPpBZw/H8ZXBLoUhPoZlZoUDGiyQN+6s8dwp
3r2OeiNiFGAuiLs+Fdw6j5kB/swLQFtPlDb2a+NRQibpni1+2s/Fq5BWZA0S+XGD9L/JPNKSrozK
9r8d2tSBySzRZhrGOHvyiYFmh8w1ynEK7Htyo9Smt6KMezcIXBmmj7F0sc1SrU+uTcnqBYvJedQP
awEy2WaK9yNzVA7HGnT2iv1MHwk8W/lrF5zw6VhGvutqDlh0gqbN4NxmbGP080cTOdv5sO1pdB9C
czNow8YXCOCyrXuHL08JBhCFtk+UXhlvR0La2ERkRAOEevSuAd2jLyAO69Cf9yfebR0+sv4tD3GM
oyA2oI1/jF1AvTmpaD0Ju24rhyLlmeJepDDGKPQrLGv9ZEsekXe8mG4RTvf18yk9yWN4ktX1zymw
LpuFtw7kGURr0k4kUAdDWuyIWWfT/tmeJpP2jr1PYstgQk9osJMkfd8ZxMdSxQUKb9/4duQwWcYd
fh6tpf+9n3ow+RyM1kD/xMqNV1nmeAQ753FfmameGO1OrI9OwpMiAJoQ3ra4k9Vw6q32GgLkYoph
cCp7JoU12bWZNNXxKvNmD61WHhxpgNozX2+ieL/kjiDI9VZ3L+4JjAkX1h3ts+cvsfhd/SeZXSlG
EfijWdU0pTH3/u7wwkk4bHwDoIn1ixX7LqTnoEmIQDahIWbMl3rYkMPMlNXiM9ALLxlSMdXt67IQ
l0PLqxfFRBAK81OsGIfeV8dyxXm4tDhiyw1QVmf4maOq5OzpfdAciceXwQny501e8a5s355ZrvF7
GSXU5QjCbySDsPb4bCY0Tj6FXCjKXbQLdsOZ+QgqMNlMnC8WJ6FtpgEnONvajlg1nUThnavKDZo1
FtBKAkCuyyjcDM0OHY3D0GYHFc/b+7nnYpyASK4N4j1d5JvLVeKujEtPv2JyW9kv3e/WxrwsGCOg
tHNW8FGtV66OXDFQtofm8/FuzfLvDlpWRnzVHTAl6ICu/CfBDZmHZT077nIaztC3JTkIg8mAnqtr
HTNZTO6qBjNpWKiaskbwmAEQkBlaB+1c7u8+mFGuiyfcdCuN3cMRijnM2VMHBpHdwPQ6r5WfhfnV
YyG8r1mY3iaib3hjdAk16D19XIv5NA29QlarZiBmF5fUJLPeRajYzka22d0DLlXouGuWvTj/u3qJ
iO9BqoyTasamnLUpS+jy14MBdaMAsF/PKAGlqC2xMubhwrxjt+PtSSoq7cg4CRmGcYZL6UNfqGPk
OuJFZQ2Z6S+rP2UGjay0mN1V68YoJnz0PRVLMYWqUqD74f1GB7hBVodJNMiK2IqCWqEP4esJNA4B
aq06pKGXotmftdHyrEBC8Z/99jCNvbPCIuXwqnvgUOU5C+XV+6Ugmb55m0XBEN/vKfMg43s5vOly
Vh0Ft5F7KFbPvlN522aM+GNb7EGfDA3rtEHDnn2lYIivvmUTfG5Wx6zuDxjZ7Qp0h+cVDnc5E6Zd
M6UbVLF5MApAMis1/mA3maDmbUG/I+kgjnKwFd+y4zRmwhztz05qrk8tjoLJDVzRQ7prC+zjErfP
FXRd2kVoGzvFMNpIvHeBrcbtIykK+d4m4S7o4EPGt56hjfHtkYZDXId9ioXfEe+W+Oz9eImVg8KZ
cQ6DzHswLP/yhDy5PNAVjxUMgHRATsnoH9s+X5EGf5AXq2iJJPdzLdqpRNctElzMHH8XUBFC4hjA
Be7YxhAk+BPCXAnwEJ7u5j9t+lNnaQdw8X04esnL+qOPe5ykGsuO4u89RDPQ5aef28HpYcjEDPqA
KCqoIV+88JtkJKPyVVsCaDI2zjtgCqfh2bkKV7v5KWafnkI1cWPpD9Kwykji7ehjW+cB6gfiuuc7
1i+Yv5cyROBdeFc+X0jyWrewDScLRvmfZwsiAtcCJ0oknOu8KWrA1jU9Z4cCra3eIxyv+89acZR+
0VSFvgbaTQ6Dc2ugPFwlhji/U7MbcqbL5yhDRERDuSh4M+C3tCOqVjGJRPmkOm6hLDCBUxADOpos
bud7hFs+LilracWrXtrAnsIH1Q+hH4FpitwcqD7R5IYIcasLWDlOQOWv7Yd2MSPO1w+Rnq/tvayx
SljkVMiX8BbWXMz/MrkpOBPFzdOhcgV3QIq73dRWDmI/9q/AJJm102P41qjsfaxeAyerZSiyONZZ
4wnljyPdiZ1gzFLMjTHVFtC/E6R3TaduPnuzFXzigfvw3NEcjTPYMNqJXXt7kbHktWZVjpVy9nIh
fMQm043Z7Kr+5kUn4rTjl3I34mMf8BpCJuRIC5HfR3RfxojwwwG4KJlbkaWIn/2UyEofU5LKcmz4
JdmagS5nDdpVTMMJD6ocHxxNZkZ/mBqqFh1K4L93KNfqpN1OL8BVB4Ky8RYrIM851ua56IfV3KYO
BBPHPA/H7uMxXLPewdG+wNSw95VpkzukcpUBQu0kRdlxNpac4wSlW8be79sRiNWsvREx5bueFYvi
bX/UvLJzZpSBNuEi0B5yVDC8lHld54O31irFBqAgbCtDP8PrIrbAHN4cN/VEjHJ2RlmrAH2w2Wy5
3qtUB9/q3s+YLGAVvzRBmVrrPACMfic/WafvrX2EyasJPj1qaSKxLrQ2KpF2LRzgfsnRkCYKS5Mj
klieSDHuTzwwgSQrgTsBadlq7H5TgJH6cPdxzTLHY45AJjV1OJhOX0JCc2Yo/JHpyMtca9XTC8eL
wIYmbtrHa79pqYLsb35QpquAcCCwC0kqH+O5BF+g6w/SvePejOOCh75+hmg8Dl4dwIktiKT1oRsT
NFEbvkJy91uH4zJVPIsGjnHm3ay5Ee47Y/W8qqmKd9A6wOoZ9zvH0VKhFPwC9ExUfGMUt8o8urAX
bwp0o9x0IBbcreUBZk/37IgXgnNq4GP9/F/P7b2PLtcgjS7zgs+3lN4MiAlxPFGJ4SwLidTPHmMt
DbVWrNxCG5p0NsLnJLs28/t8s6e9yDapZkw35zk7Aj++TXaMHSoX+dOSJ5nF7MiUkxYV8VKKsA/A
lc+og9nzqYPVcTuGroVh5Y/5BRsZYmgsCliz1kEJsxWbt+YPKqfeBnnsGR2bPmKoiwXDIIEkA8eG
LDUoy2T9OA7fQxlxnLrCauOo0iHMcaCtxgKPypmnqYq/2U8dahCJ/Fq8Y9ZtPdKPq9CxlZUa4Fgi
Zfx3EdX94rXstTPzzy6Fc6sZ5g+3W8bjqdGhHTjYTByUW4yuTjiwQq7ugkq6H56BTQFJLuLzj3g/
U4cpfdeNSVmV7KDt1y9tB5srYmE7OJTPSBgWn+hUNEA8J9v8jf3fQ35FLj8P5e3ewlNvcwWQbKdr
UyBTFKW0uzzpR2SdBvHlr34dLP0+/6gq2E1nLWPneO/fsvrVqFGzCK25058XLh5H9TNhGU03iiN4
JGCD7P6Ua3YTggaj4VkjFHD7Dvgq/X5KW/2yUbOmZH0OM4vcEb+XTp3Bp9tS8A4Hn1ngxUsET5pP
KvCMUumw/QbpOTgGImJwAOkbBqSEjFVULlpBzAfgDRdb88wlLHLReTIxKMIGgrYM83p702AOgZDk
JciV7UUtycdHeq4A9DmaqZPpASg5jqP7WiLLKqYqrrgxE2aAJq9wNE7dqvp2bcwHq3IfzrTJQKIe
rmCZs32FG/vVsXdPkzHhS6y1qT7dRqVqGl12UHvTTjdYwtqqs9dt/ozQlVAzwQ+k30zZp7a0y+0X
aCte3oyG6PQ5aQiS116GdDXvWJYwCl80rMoQWYA4VdrLT2vjGjYLN4nvhUoKouWXWp8eJ2x3lr0J
Lh7U0BOXWVFpzy/l1/bcESZoyra8YW+TL8OhVvV0h9Osp/EanAI6aEDBCOyS63RnWs6JjSxWb9Cv
/vOsXMJFEm5oOUfJ6ZhqsCQMVmGQgtMlqp2LxCXDfsAP7xFoYSxx/Wv0uaL1b6gVz3o8mMrohUmz
y2sl1BDSMkuv0fjjXHQLdQelzsuS3RlCPxUTJVtS6pTZy3VzPVbrlR+APj1uVwg4N9STCX1jL2Dd
sIAI2K5T+ih4yjtxYjuNpD/89aRc5bY73e7fWBPHDSrHZfwAPqh6QAhyb7Cjg/nk4c1ddL5veo3K
x2DSD96klX81E7W/hww+Bopwlv0Gmk5hiiQtnpJ7rjD0pnm1Mjmatqw3cVRfAI1R/SJ0lnpmxNWQ
33Hjh2WS8aFm26I8I5nhpZ7HED6TjNygfNKao9VHssZJNqq/9RLp43lHUwv2aqFuwdCANXZsjIp8
Mdb/Q69QySKi400CH0Wnp3tWHz/QWfrsMs5XORDctNEDk+6Pn5GcIQS5f448nYpjNvJrylYgX0Yg
T/XANCVfESUOKR9vi+JLnLQ93nGWIgANnHzCi07TGAvuPuqGiTfFcHpq2nRBM6iKJCStZWvnHwRs
a4nMBglw6DbL2yJF/tNxWy5yjOGVL2vagVYmCxWBrd63yl4PhiwAKJ4hEeSMra8VLqS7KcDOjWF3
maPHKZUTi2egiWKMYpedYiVzc/NhgHfJljgR7gYc2dMidTttimByP6iqHfOs/pm8VzbzZOYHkImn
qqBXkX+4mgAPNoHviMTxoYoxH5lMttpH/Y0kAMYtSqiE75Y8pyGa9usj3R3Yi+xaBlFen2LFqpLR
3xCErVmmQYd6jgEyb89mzZHti16+KwHSHadCQBknqGgM7pst9Ee5wpSvJkGl0OH7lLigI/XGYBTF
yR/umWfb4e1KX8oLgfwPOAE8CQ+AVwHy5KmSESmmf5encpgBC1nOOfW9pWrmdEo40vaKjiuIeyT7
kxImQG+kd4jAtOnpc6P5RI1RXewQGmmMR4lEBCp0xepujfNknjYEFPtdRFybi5+ji7Jl9qfAgWFL
zIdC4rYqex6RMA/5U1XrrhVb2fvX52R2pydAzxz/EFstJsV0RKpcRk0bJqf1w04EirAfxRWOdp25
oiwF+xvSotX013offq2NGl0NmXb75wJdE0rZofPZqmr8DLu9KYibAy3fATD7Cim9FFX4PBz+rNX5
4pboG9LgE4J8eD35dVHZWvYWv/0LkH4n6/iclLtPYXGSHHb9+ULatnPDXL78JQFspumKmBa84Iwy
3aICa3/NdTBLXSPpmYUuR75jeq8n+/lWBV84SxSvYjEPeb+c5sigND8041XSEDd1FBN/s3Kn0dfS
eoI2uyfa1MC8XJwXgVbd0h8ZJfnzeUlrnwmdlPRQczAJIocL+j/w5+jiAhqZPSndNFLqYkoU4FUW
pV4m6kFsk6ZbqdPEWgDjKXtSQUe6ZL4Ze4xeyvdAAnn+bPD/TgF+eA8E7AFrvAm2DNsWrqHp7lYu
LyvLVCjYJmqwVX9PLezfqB/RxHcRj24tApRu5icc/z3WLakLW7pT6QFv7SDcehfL2Ia/mq7AnNff
cmx/Jt92cQETboUsOCaWgBWlTPodABKscRzrSywVQY2Wm4pn9kDIO/HBQxdKTVTVLdL5jWTQcss4
Mwv253jWe30FVa1vHl28Ijh2N9HsvuAcLfECsOY9/JSLFZC5sqTEmmX8NkGrSwU2HeN8HWne7hWk
v/snxW+u6SxQEmIjFFSgipKcp3p68ZAYw2cMaW2cCBXEEmE1/JlDcLEE9V7/zfiYPegdlzuTtf69
R7PhvCj/t5NE99xUw1WZrKDGOargrHjcKKhBHHztJFyvxUugmbBPWWiZG8wFjg055RF+uNzScITa
Ptj0Y6+i9fF2csyNiqQjhyCWiM8+BXFOZ9NrZSvJBE0YMPMuPF5WjyHFwPTUIDPTyUuPDlKEps2l
LHgfokMpCWUW6ZRYlqJ/Gvn0bD346OGij9bS+UqIAR1+30658WfmpoGtNDasX3t+Ntfsw3w81ILP
yClL1054ybDCWxHPG4VJZyBv2O9ZY4zjKa32eD/+BzszlZiy//YEiNHwl2q2CUXosmvl67LH/lCd
XfB+2UkBQGCJJGUkli9+XKXgmRobCoqc9SDEwzk+slZV23JGVubbi24Npq1Ip8lW3NsDA3j4NgU7
rWc0rBKWgmz9m6GgZz2I3/01CjB5dTkNjnufdIBOK+rHE1KG1LOEhdUSu/2IE+pJag6BafbxHyT8
7j5rEp6tz34EEMqC6imXD2d0Sd0OhTZG728Lpv7etgsMzpGH6e1nDEG/DOBluqxKSJxN7JhxmYN1
M9T1qBcbWsEpeVuDisUOdG9axZGGYgiRoRN+qQk7rLCDtNHOhlaUYXOplIm2RM1sGeYh6n4lOHBh
uW8dnRK11suWPFuX2KU1pQBWhh51c/kZ/aravfDmbIsIdJpLWgPEnZzAln65kNxX3j/jWQ8bY8M7
Vmq7NnrC1Y9Ew1eBweM7m2v4laih0JQHKuUSzuNCaUSR5IZQ/BtLw0yAFHLkLDscUS1ZodaBi7wq
XE+aK9k4xiZ3jXUVKyKtLvyRmMl5d+4WBXfyahAIVZXcA2zY5KqYNWWO3I1gh9FbTmiwfW40/kGN
DVutTyd0SYr0fzA/aP2J5sqyHGvOIdddBg+XB9Zj6vcXuw+klOfoxegUvTizubPVLe5pjsMeJEHZ
iydBMk4mDj009wL/h3we4zY91kFrICNlK0LtK3ZxNqyi0zgsK432fkaJkfU0N/03aSsAq5CKYlO3
bysifRtX+hDJW0oQZMeoRWQU2QqmMKnw0KtnPOUIjC/hDd3u2WhDp9f+QZhBAAWqJFuXItA0mUXf
nKdSWCEtJB7dGL10D7nTvLK4Do/0XNmRSDRSnXhud+TwF+tbQ7zUs83BZPz3mhDbemeN+m0fZtFt
38lNZ22hjbwL6E4B2j0TNG4sdIEsCjPh14jbb8T9HaPGu8SpxXsSZKwROrnJX6xIStzEq+1wPPVo
JrRvsW1nvt6nz/2+SxAiYo/CNvATRExdC7lUwqTADcU1XxLsEQQyDGpw0KZtuMwIabfgQGcj5fJY
YBVX0cmT7ziLlDQOu4DDPOAjVAPuQeatRRVsOC4qkctkStud2Hub2Xjag/wMJqSGc4RCq884PoIr
DCNEDCnjVdRuiWCkVeuoBDJrsQpn8Vx0CL24VFAURG1weq6vc5VG0NKuZmZEqHxNrJX0HVtw9wnE
UFV5zh0BKPZ0yaOGPv/dD1iHyHb1VYgvIvnX4hyg/EbhxnkZGWuUghwj2z29dgOgK82USyFoq350
QnxoM7RTWfF6DYuxcKJWqjdqGA2C7P1b5Ox3v1zi9OQPNlnPLQAvSH9odH1m+53WS6lHA+SRTlNa
cHk9h6HPU8KoddsebbZANW4MUv08USEFKxrbnhjnVXis/J6QfruNSXgjmo8AF94EIjWa2XWWIJtB
NBUOihv5QQqOHj5LT51cSXcYF19YTSWQ2mPTR8+EZlkRfOjgL+3rcpxUmtcOhCj7VW5GKiVAa7ee
A2n+to8CELUek5TzRlgJhH5YiI0Iz8dkL6Wbzs0x/yBtSckHdYCzSEI5JpgSnhHOQiB+IiWYj3fc
FXrTkepMwwpzWUedoYrt3guIXqn969tNFnVALW1w+RQ+rYLShlL7VFifWCgjBqQRrkCKSFJYvtuv
tPISsSrFVms6nmU3OU5vzud0O6Qa7upNdzVgerAk3WqjOMfeOIYZKCuQFOY3faduqs4ll4Bg9HiC
yrVeKl68sQr+22IlAZapL+m9dqsUo5vHteHCvZGVN35ixlBGdPkrkMyYJD3dhA7PdVzQxa/kZACC
UYS4whg0AtQN+eT4VoPXDojN/+BaNV/oNepIDTkQp/jFhkizz338aN5ilrmOPwaV27kB1xSAfl7W
vTPkHsbg+5OJnposFl0IvJeAWQuDUqCAZhTZET+ZVEBBZycd7duXcNwQrPYL4WOcVCbUs1/wC2MD
1g7I//Sc16lpG+AcWptzhnJ490hXIXzajCPKJ8hEy2ooy2qo23PZWhaYRW1V2O8y+IASParYFArP
myyo02RKpj+dKRqHEnMKVejU2wD5ol+r053flPXdH4rILC/EJUChD/Lf/om2YnOXzMnguwkJlJEV
noJKk0mkxWT+yhHyOqBPdJp+SDTzn4smEz1aRJduJrz0y45ovtYL9LTTq0VTJKrrMKv+q8gICQ6E
G53BQ4DPuY+kwvf9yMsTzH9HJBcJ+IuANXfW6Nj1a7m4UWdmZWkNOigSXSQRyTfbxJVkcRErF+oj
RiHTMHHOO3KvBOebnCX0f8q/Nqn7hr7fZd+ksvKtqXN0/KNU27DHEENI8gS0h8s6ytVHHRC8hQVK
9MyF3KwsJoYISvJkk1tvhJACrA1EV7cc504AhNEp06ucDDVUnWyiZ2XISzjTu06eV/qmR1qxsD7o
QGJik1BURiOrkfq85TBcsbPef02HsylTcCEDswK31OXrW+XAHJ80EWe9tFv7Gct/tnj9Xb5JlB7k
7ptdClLoMkwnJJivPzFlPqR9QOdFdK3I82WQQf9/nv/ED/3CeCFWKZPfiA3EFShApH0kxR0dhsJE
iTu1ZhT8jsFYNINzEq6TKciy1+X0XdZpmk3X1Jpl2aKGNHYQNTf4ZOx9jVB9h6UriDJV25o1Gpv1
bRa5zG0QVmP0QPe51CEVFkboC4Ms4EzAIaDUQGE5qEorbT00UbfauduBNB2k/IRtVsHLN2l3SzXi
9E3qHKnDmfn7hcFMGaXsRMHtEZ2h9Cy80OxXjqwyhP6pvswkdBTH1Trsi56q63/YLEo/TpdDRxT4
PF4nvXqZTeYctiFJLEIA2PWqWY0OczafX/1iybwxieiXOzu0p5pOip+6DHFqdNU4d91A9DySNxtM
yEryKxW7eJXAAFWmYPc0dL0/parymOhBaTAOH+sGltvIkUK2QYd2Zxrj7pH9HV8GFN/q8AsZ4oo7
VcHxVpW5cBlUpHvt8E08cX+qQWyZPeuvK+T39ONWZH6RBu/7u5CQuwELkD3xzzxiCFBKlCao+W3V
X77D5661mrvOaQSbvm13KMwSO1kDGTPT20h0c2zARDZuFAkcH/kj6Vc1GZGbm79rDsGenPsHWpEM
wWBsD/fHWFLbMUkV0TaYQdY2eXNKoIVTSiyGRs7chpKdlbLhEYen/ZMODhdKZPGs+WOzt9q24N2G
BRQ4LBe3rUIZcwZHKAMD34cA/6R1cUE1PqLgP/bdDuedZNhpYk4PLwBAvGR5iLZcdH68GwWAuLi9
zxwSZ2HH52TRi8IZdPgTsIE3j5LyCo11CFgX6WgGcsQJB2mlX2X5sgxVlakDAkem2sXD+DcKaK3a
cRQJthtjGukkqSfZhgHWl5F1Z8lixFKpMrWYzPCq+aUnyiavmbbIW6ZidHNpgGOV0bQZMyECLmMn
S29wlWcJbhS8Uin3iSEBKqFZmhSy233OlR6Rvi44yyFvWjjyn3mlPe7dvC8nuzkrl1sWyDspPmlR
fwK3af8amPVUJNbwIP+ULnXLKcZqPFOyNDOhKPpOUt31TiWyFWq540CIdvbMn5uo+4g/WOMCCDH+
UCD10lQNUCArMAbZVA3Sb+p/cx1CtTvwQ1bHgbmZsGMttdU9XcuC1y3CDJRe7BD3laliP0F5KnRv
WxSbpQdaJEZnOaeBjTqy/0TkM5XiSsm8wN8AFIRZi+jx2MIJhFKnHIIsda+QzqZTeLUqD1x1M0KH
10CzsXpopk1eWuBAcS2nU7EAxcAxmufhofhqRnmLVCR00k6YAljNvBd+kAr38rlqm1mMgSxUDIhy
dNDdnR5qnn6xrfLzQBwIwx8SVfJt1iECO473fTpjw+BF5cpVZfz0olBPVly8DuJ3d0pl1pKvfgWv
nLqNAz8PHfEwQL+Tk1pNu1fF+WDRXi7qBAHZ7UJeplYESMZWX+AeXUg4t0e18y+BGS0oj+jDNcpl
CNeRhhQILTvb2UomZz9qr7Z1djJqBwDFbhijWy/ujKpVhYoQ2+nicm0gI4frPzH57f1SSME91UfK
LrOke9MlndixOrmjXOmpZvuEPadVoPXP3nLqSw26+PrWThhEg168TsXSpHViVpFN7SXzmnU/Owbd
NoQdZVjOk1hVE0iZclqyKuahhTcKdaKANiHc7BNkIbIK9jpLEpKZTnCvtmASag45Lt86XPEAIzM0
PyChZM0wIg4KHX9V+7ldWjNatpDHfKv/aX/hn/OSEHPvV8OdW6clDoGxKcpW6NwMgk1hboRTjOnD
8hAJCXwaSi/R2p9jtJw2uixIaFvJTRglwb9v/s4ABZTKT2ODx0xyQfu6SmWeLfgHuGBHoSh/nY4v
Ck8sessO7zonYtCrfFmYwpH6eZK/iEnRs/jE6AxY9+0ItE2MxnYhoyqfaYPCnVXMEQA0CmOZz2EC
U3ILjpY0ozkNsjGFv/xo435ZQSAoih9XYHw0B4sAM7kOKJcUnhAnJkvgbBt3tgllE4lhsVOtW7QG
K/Z6QAWbgGtOUiWOULG3gxnb/wjpkg2lwLEluvzg2lEhbW9MJErzOlE58wSfUt5pIsg/teHTz+Or
CRUPP3DpzeNcXXQFIzrcJ0ylmu6/aIV/GXPLStVzjFZSIkx1IMlRN9/DDBtkR1T0rcc04hJJ4801
1jRME14BvG9w92OR9eUds9386q+qrgq9B/tMTSKnuYXTE+2FIvKvB01KxgLIFN3xRNkPTcelIMDm
SuDpLCmyCnhrBUZ/DOiDToczVgipqqRCKNU4/OGGkGIdPMoIBX8snQzFBcUBYXKKpfzEsOYlx5Qh
G7SwQlT21PYOm/uv4itr/bBvyuhz9ehOjYuK3PS/7JZnW9pgQCiUHmxY9O8sGwCkRjqWEUWvmIII
I0gAoo0y0G7atOek/y9UgA8mg0jqDEUKbTuSZim8jsOPvFMZOVxMx383O8q/xE5XHHuPrxs6DLmz
nNOpyNtWl3iek3UpO/9GADE+yL7Nj/kpkD45C6uvm5jZZujlGE+N9Jcdbvvx78iVidVSfsaFfjQ3
mq4vVDvfs6F4Ny3QTKFQej9AFZJ9Uq4xcLaHJO7BWeBHeSOZPuzn/RwxyQcsUbrLgx6my234vZa6
usRvp0cH3nV4N/iM3hOxgsEgeAUtbcvCktomdMtHaRu8EMw4WxID0LuvnsXqVxKk4R0tnuQv2rbP
3F8ehMk41WeZ/kcemIYuDFEk4DsEZ5CRv1KBavfTC2BUVMQ085mxuY/WMlApI+mrlLe18SAK/A25
MPjn0Xo02GGBSu/p3RfGvZ3xq2f9WIV2tXuEnO4NI5poJKNKTtYOrKa34cjwB3Y9Yf5Hv20kufDe
F7TnPNMkAk5HWqK3yr2R8aiHzYIKo6Oz4SuH2d0DfipriaWoAjaOVSly52BvsEICsHZYriNfXHy7
qUuP4B99HKgx5HRk3A1bDv1hvqE++5V7La/9ZRG3PHcAiBK3uDPsi4GvB08EJq2rm7Nr8PeDpln0
WjOus6lrrx75PldVjBoG3SC997mIw68dukPESKqVJ2w3k3EBrw0aIu8LHTsRMztrtMJHjlWOwyZj
KEBQZkBqQO8dn9hjiUzP3IyJ0luAxJtJXYePXYkC+7fMBWxRlzkZC1gzH0jeAHBiRVQXx+MowI59
nyvri6J3tUAjR8eV2XaFXiMU5ee0e088UWamHCdet1kiDmOJP+5jGmlFNVOB4+oe9xv2AbZyhMYR
pfI0bptStwvnCrVqVAteJ/XZthu/+ExnKsjkjIp6oOrFS+BXrKENVQUWCZVd2+bM+i0Ym6CX3FI/
0iGXT9kUh5785fjvUyRzDLVNT5RipOuGNRzITkavhWj2yu4wmylgwLrO+EZGD1THJV96GLG84ywh
gIMZMK5APW7k2OiAr52baA09G6MYX9Wv/t6fbuH9KGb47tSXZbpsSYxmYbpCGfbpTi6h6OudY1iq
vkvOYRuGs6FfN6sEtfKbImUlXwsy9y6nySfOaPSKeu98WDINxOjYmJ5wq25M0x3b61Q8rXb8wLRL
UPpcVgoLFemZD4uVjts1MXWL4yHGW8Y2SAiDzunQPARFtct9himEc3zzIpifx+itzMQDo6xd8Rbv
zmM9LE01lP38m1MqW+qCHM/+K9uv7l2EKPegiQQ2Hx9FQctaA38ifaeZJAXqjQBPmpdPfF8CS6ux
HtpSzv1JUANTbmAk66oEdZDEYiGdqdkqoi389LN/KspxNGYrD3rN6iwx74iVrP+FZZ93ekzUv55m
LDsHR+8tM6ybyQX8/aRnivenppldb96Nh3WUm1jMnRQmzwiZcTpMPVYplngiSRn8Jiq4TC2dBCjk
xTejenk/2p1lBYYFcEazHkmA7bqo5fWtGi8Kw0VQl5Ir9c9KRHPmxvkKHf3VEbM1ZhLH2M1V2zcV
ZVm2MhFYgYlJSr46C3XmNGb4poXTiv5Ckeals+mxNWuX4iSPlHtc9Y/CnFy2kKNsqmL+KnDH7Sp7
2s4maEeIY0LIqbIDWjMC/LUPXKy0kSfZP4Dzj0TA1THybInCKC5IHgivjFK2j7iLebeti76rLdsk
URdt/87qku/1J/L1tVUEe7WWm8H/GVOM6BfwEnQfhMrCbJF/TvlxfG+kuMztZiGqYKgSpz9eGxNb
zLRo67gSvaK5nybJtH/fkZcDNyN8xnpbnX/ltiyjKLXoEowv9O3WnP6WB3pQqB0emhdKPQsW2qnF
0wbzIKGBFjKLHkpW4dKc7WgBNNFBqh8q4ivoU3zFsTznBVKVn1cyRdVmdAwccGwfPiP9EFp5QCZB
fAqiG9YQP+dlKZ7bP4wyoQ5MIUdl+QJoPLurkwAhZ9cD4N1CNiKjdleXxu7s1wDrRgvxFwWbaiQN
E8acxi1a3lr0C9zmfQpTusZV0iWJT5S+MsnvIWX9uZDqChr8FYfxKY9fxUy9QJu64na//GadYXCC
KbIP4NgyXCQIHYCW9bKFS7qXQb2/abONFmaqGblh7TkRfo604KItHK9eK+u6mEMzuwFQIySsL2rt
IqvQwmZu7TesFC0SOLAs0nvAAK0SyBxjUKOb3xZ+PbNZHkktCVxovYg9UcHDQ+EYWmBjT24kKJb8
aCh5kmZCTbcqdbctsaaiaDq4qLLnbD2EzjtY6HjNxo8Z0hlzL0XofdzPGPI1AfHBckKJWSZ4jnVg
BP6UAUTqfobWltq7Jc4MVI5Kv2FB+vVlg+f8JexkjtbiELU4Ec7WEX5NN95Ds7V5mshJcqKiTthT
UpbPYtI5M7q0CVPtnk4ivU4uKfVDK7KHXrxSs4AYb3xIadVwa8ml1Asot2O7ihH49RGcyfIPa30I
Qb3jvouLdS8RU9oNStiDdreJf+I/m8idlZ4nGzfx+xKRLtk1cBu5b3pBu9CpVcwi9guoXooFQrbD
KYVAQ8L0Mn+imWSusahX+OB2vOft9tLHxRSJjg7PpveVsqVeBs8krdXF6DpDvyNk9OAxAcVIwxMh
+qfLMFY7+Nm5P6bbjmQUZpqRAJud3u023hnfxcSROmSKpgItxb7zN35f3jXbeelc4xEJLyDBNsB5
jVVr+4MlJhLiFucRgDnTKWafZTB9wr0HUVGn6c3TUWoZhszJCcH2R46fLK8lDKdx6EPdoS8O9kNO
C7dQjHa8YSnJ47hGRyeB3eTOelQCY9/kytAPivPEdbQl/bHe1wiLo48xG7cYT+o+LWU9qTwWkWkC
2CY3yVa27sSib1Q5xUdiNBPvfCK9tJ1C4V5KgwkPYRbPSfggDChz3u7/JfoqQ1WU+3+AIGmHlgq8
SdnIeXtUA8rapptpEmJRVDdxN5AO6AG6rq5jhT0YYJubPLJ67qu9MjEYEShKOAHmOZhIU5AUn1ZQ
+o8yOMI5R9B3wBTbTmuji0FuZPKjDIAu/j5zF0zINDugimUkaJFwopnfb4HZlMhMrNVb/1Z5CzhO
y6HfBGbfr4kyuR3ANXIuzZS69bsZH5JGiSXR1Q/VwxpqzyR8zw/kjc32J6aNx0q7H328m6Zww87V
eLU/PlDnLMq6Pac2Pl3hty7mVJDSVmYDwR6asr0cabEXItAxuwnN7EbSRf3GXJ/RmqxHTeBttO2X
iMClYEu+kh3I36vWxBqe8CAOPSP8HTO0ZbhjvWLiQLLcLTADKCJUJUsfeKC+FMhabea+zyEqv2/z
ab7LrCqJXvDG3u+IjQ2tMBZyRDgLQZ/uVq7u01pvu4UMLNtu05c2YX6KXjb1R/lAfoApApiWsfi1
dVWiJOUeLgzhSsRMFtffQnFbtMWqYMxBOV9K1IFdLGsbbpJJG8PaM0T4FgxeWcAAZPLfwNKBP3V/
FCrib4lL2Wqv2JxYV63+qfsD7UxIm6EQoCmeo4NKF0qdXqO65VkThwIeHTdSLT+KSHFt4xkZGGye
uxwc8H6Gj1MUiXw03uAXRJctHKENsgvOftVDb3vL3AUEjZHLA8+UFA5a2zbJcPyMX0CFt6d6y+Ip
yerw+sp0f2W4HH+2ap6SWFT41yO6vDlJmQq7mPXurr/wZaHZHbcpWqNomWMheITfullrrc5E6ike
5rg1LPhnDu4kOcMrewYpASb6BIQImkTvpIotyk4WaG24zmKBKWY7dHUc5D4ax8YXL5kcdfTm84cU
8aYB857X7lBgIppwXsuOp/10a0l4iq+UEP+uG9symTzaZcvf0c3YauMI2C32Rp6cfC9f30sEjVy7
Ff33DtWTBlntapmIH0iu8PE8An7Qs9iCzhExdZlhifPl5ryrCHS9VJpZSAWxlBQVXjxFN7cW1Ngl
fMYCk/c+FjkWviJWIitoRNKBoyFUvYOBgDtyb86hyTuR0ob/wW/N/mzS2SQLzJTTLCQDP/VDyGli
chTU4GDnBTyhpXYe7U5xS8w+wKHrCYu9AofgKsGTbYNnT1u6wsh3JxSVlAHlP+mq1P6r3Zhjt7GK
O2WG27ONVKaSkO9QooWGFrgBJRG5CCV1kHuSXKfm1wn93VTGaEwPzWvWHzq1aJD3+E06peXlm1kA
9GaILMblTBDvEMTl5CzDSSePC2QoE8+J+CF6PLfKu6PqM2+pB5qBYdfYNgcSz3kpePB9s87hO8fw
7R+CAYrsr3kQ79et8tdrwcQa1/8BPoJlAyDN8pwUnjAR1FNS/oogem/gxqqRgKt0/X5L/b9NjAD0
2TKpILITBykLscE2+5brJTnCyhy17rb+Gand9rQOiWlHF2pLv3sFW+J0051/+D4/X/eQh9IHaymL
UxfxnOsadoAOH2X4R675iyXYEQPCteLzKe8SWwyaK5lLABxEEXS1R09dbc8bG1mSXPrPaCL+aLIP
1i97y9gPjsYKeIiwmnGt2+cygp94Wwzv5IsJhxICHFVhFCwM6d7fMgrveXmAGNk+mnBr4U2mud7x
A/DishssSztunqXJgUlqMRNTPIrtTaHbt5KvhhzlZSZG5hPpBg/TsV7YqDQnKFobcHOD/qz+z7qz
1JDzZlNuCs/gpyIFSuR3YOl2obUOSbOsuxdoJrIgi+FoZVceDprQXJn5EnqDDE33VGctEc4homlf
8c66J1jhkH59AYYpXcDOho4+X0wg4Xcr4ETR1XDcZqzaXaEUhRGcRp8/WIa1XyXAK3bjiHqTnSDZ
g8PdMhNnfHtBTX+8AeCV6kLCW8JLWQV19S8IkVp8Ulv3xuw4HQDvgeuyM2GYt+V8TYFdZeaXw+L4
XmhjeCjC8I1pMPjlQU82rri5YkKhhKFkZZga2wR/vhYyLKQsq+yvVmTftAg5m39E4qvcTJXHb5ve
KhaWC26dXu1vZkIEfdgsJlQrXq+mZbyQw9vxeKksnyhtOdaXmfOwjp1slp4XHUJRYFIhtJYPWrRl
i36uoFLkAS5E722wmH9AcNEWVNoFjD1MBvba1ydyGfCYQ6LChBCHGRmTP623VRoNw+n0oRJYV7JO
g0dkh1g8QwQYM/2BKvx7h/fyMbvxw8kvWW3WSpafoCuuf5D5P9JmorBhwSs6G+rnWKlqF0Y9JWeF
a+CEgPdyjlEVhVeNwZcFNBes28qUjhxOFskNzkJAvFRzdoeaugh5hW9Ua5Gs2/tnD94+lKbTyFRM
uHVoYBqkK3HfmJKJHhDj84m0/ZFPiEUtL8nwr2bQxKIi3Gj6wdTMGTcgTChvfohxLstKF6i63FkN
NPKqBWn4we0UHiVUcAb5WAdsTcim63Pjt4A0IKO2avKhyJ0C+KqrIad1Jyd7ZheAx/Gqh3xhjqxU
PLlp2RUJqrJ4NmxwcrzP20miY0F3Q0Kp/TxIsAoYx/ZznI9K6Mwh+The3m/PQQFVAuSVRIE/hoeT
GJhZhgwKBDfH1FyangaUObHVphfYkkZjLacWsw1f83c4ypShCWbAlnMEJ9mkZOS1hWyeefvF/BhI
mKEO/hW0t7VEeUTK4wdBOzWmFzsL5pesbbGlSpbgWUESdZliNX/1mWZDM45aEu3NWM1ZuAgarHBe
8W9Ri9g13J66HZyNq/WApsLofmG6WkelYX5fOEYXhWsmfwpaHdLHYV3O/fEiJH02Rs/uBBPVCcni
56Trvh4VSh6bFn4IW5tOyicHMY1iukhHctnrkVnb70+uxdtsGoyf8hT7D0ws+9ce4p0tohtNgDIc
C/3K0MQjGntfb14R20g2e5O+C2rAfV9not8FPN4thhtUx1+YmMDdvUQFgMVP+94KdXMXsNsA8B2A
G6XXHYIvPrMb3ElL22kweOV28fOELiNfGGSMULB/6SNt/P53PRmsARkZlHhoEOxasDO70HaDSmGf
tlsR+rje29AICl96nwAQxQfjTctaKEfKf5nfareyP+/mNn5xlD2USjagE/07gNonY3EZJ+FqhOkj
TFJRABGgbFgheHclQpIxzmDMTk5ci7Vct3eLQpkl2WtS7XmOsQmWEXKT+r6LZaWomI4LOTixPnP9
jKeSi5vEt0GMyqns/TL9nPf/MQk8Y+lrquZAwk2iqf9SJdwQ6p7qXL2DbpYs85p+Tlu0NfzKbGCE
4DIUeY0PnLrwH55xRlBykV+MB4MUddGu4qwxDCKtEthoZaXbEMk027pC9kOkvtoqO5SnYYoVyxt2
P3Z1MZJv1NVXxKU3zChBlqwXSLKJ9G5/VEgtGisSCcmm1zzXkanQoCSCwR4hKVSnfzIz4Xs2ek7s
EBVhfYPn9VXnBRBM+zx82vm6aCKlgi+frZvJgEIcMXOBR5hOQjAYAfQXAFYXh+Pisuee1lDxXz1a
zAgWns2qHoIH4876yEQRLnkYX01d0W8PVcVUWk6SFUutzOEYepTDYvmqJQZh01Vm/rtgK8mu1v6g
hKZjdeu58x4uO0uwC/yOF9iBFWSHvyerr9awCxW2Zu9CCXQNujE/4uS65cnwAVZU1SNzHzDdbsMu
S6mWSxhYUkUqpU0zeBtJCIYcHTSZuV4dbemZsctxU0zXI+2ZSZJETpCDe8xh9qNFsp7af4sIJKXa
fn7bwRlk6QlCGX0FIZFQl5d5yKfKLMHjjsNbUrhSIFt3AP+SvJMbi6e9UPmsNlY/IDuABDs+bkGW
sq5g0+W4u8dSEk7wSGlcvEJrzHqYt8nFqW0BrfDosAKooRbkO/3+KucqPLM2+pxFsZ5FrGdG9KNt
epwGfL/ZNcpjHrZFHdSD+qkvKz4IT9a8dB4kmXUHgMVWqFi1GKjnvAY27Ok2hFbu3LGmuAIbdfMI
PHl5UGtyAO4zoRbY2PH2nro0Xi+Ade5ChV9xTYknalZMcxq1JOJgxnqyYDJ7/Q0y+v2jpB4cu4fA
TI4Vr2ck0ML+LfWxuJslrgOvpgHqXwpsv9FZh3i1KA0vYAgTZH43jlBXfo3MYKPoPXprcmydvf2D
/wZqqTZduvIuz3mfiBDSOyIvjmocNA/re7dDhwPmCSrjh5FfJr3Qk4R3cIoXw1LX8Qd+XmKkwlzh
gTKHY6tUZa61fvuT6Q7Pkhi7KXaWqNlHPVawKWLMKnszjBR6dzlYrIFkYxzTNK2xGMSG+JFLZ0aB
gTFxHYrFRvi48Cc7cHNxK+2D+gDCFUzBRaL+JUCWQgXCO6ktNPUrtqeZbnn/W2PJtYmockS1M3y5
2CKAbkXZS43HD4xMhpTRCf4hHrxdCOH8KSQZGoA/QyN2Qadm55+vK9IICZm7Gchj7urVcgQgQA55
gllX1WaZCfwD1gVnFW2zSpAGBhOUMJVfHwKs9lPSdzDLe3nc7T8kamqd+qm6aSh20SlPTtYfMOqt
wb3QRgYjGFJ1vM8EZNqDiOYh0NtORT/Ax4WoHBNiMc3FOYsrkbEl21tETzXNyYI6MNuHdmY+iEKC
LMptsSL4diZigkHa6olDptye/lFaxceOg78arpJucqgCPtOkY5csalAAaEY2OIojrtQEtfQ6tSbG
43UeUvAezwV73paK5mk30MfdWcttJ+ihmGuLMWiApVefc36v8MnvIKGZmD1wlQELwIDOL9b9UlCn
T9xg/gYgeNCFqvcwEWxMeHlGXv6ipAZXDRMQmzq6l7ZL3g0XSXpvxj5p24MRD9Vc4qXCT9F1C8R8
xCmjGz7oW98xheynobGVD12+w1fTm42kS4GLSYg/9uS4t653gvHllO2tLV4chgBsF0Rv0iyqEwwm
TVdobU9VqQiipUKzvVE+35ricrhy58eTn1gVXMKna3Wp5keqmeFTr3Wc+qn1wBJtZFk8cuodhLfC
002Annkcefa5o1dHJusgNVsBrv5IO6gnDXWRcg6L/fmHhh938+m/smaCM65k5UNWx90IQLmFj+d1
G0uhYcjg7ESJnPetl5d/VBWr2GG/8pdalK54HzDE7Wl3Y7F1vbrtD6YAAMiBTGvXrYxdXA0iuM0v
DwlbOhj3no/gzCwR4MrCD6C/soH3/EgAWTFCPfQw7oqKfmKkz9YCdoTe8714HpmECa+8e/Ymv6yT
iu1n1MTzlzr4VT/GMwyaKoFvcP0sO14pael3l/x7fyTx//UJge1oBvJD6OT67Yy0mZavHvlwLEXO
ahKl0abotus+E+aEG1IabGRebhH7dxWrcgWIGm4CZrL1TRWs8Y2fO96iHT+clyhj4hNFjV/viINs
9THEHOxqokbIre1e1LWnYvIgKPSLzm26XKNOeT0PJChQOWCDoCOy7YRZSh3CHDtivORYvk3QyEtz
r+4kWXEt0ZxOaokandHN3kUH3CUu8zhW55TKIDUlcVqnBplq442FUwd4C/IF7PUjesmNhvUuPV6I
QBa0EiQ47EVYaaMLHKo4F+kZ2jCn9L4syHCVPsjurcx3IFmxGp0a1TvfQbw1qeBMtjWu2WXKoXWZ
ZV7XMmJpPJhnEovEjnrrkgyuiVzsEAUKhsTTKk3vTztDTzeBrFbIWaXmbZp65fPaci9OfIBf1fI+
vRbUVAuXDB5YPlQgSYsfN98DKg8WDi2ZbiBnX3ZzAOUit7H0L5sa6Env0J9YfTmV1JJRsNBLxKnW
NtyiDsqIgawByekTvnefENwlD73HIv/TXUF5Ghny5XE/jjle+7opMHGnqc0fKZSIly4Pb+CXPuQY
uZlb6yuzhON0vsYZmQlx5o3IAJd6/JMyCWIOc2Ed9OEd/rq/Rx2dkBl7LwIXJZrzNLy54tLJDwwN
eiPtHWhl5evxLmjTh/Z9/8ouInRvwdfUfeol4k3Vm16Q/sipsfh4K8gxmF9QHrUPtx1bcFDHKnas
wbdOYTW6eQS7DHsa7k1MdIOOTzqQihhs+v4Ppreo7KO4jn9xxadOYYGKBMmalsYqAPy0ZuL+pymW
mt0GKT8KWO8gWW34V1RM0zXt6GncIeMgf4VAcsEPNBqZT2KaHq45sSXUhXbL1neoO+GSJa0PxLm9
1Zn5LabkNfNSyFtQto/972Wmis63d1XqFup3EfrFhjOTj7fhMM8EdclfZozv0P8ycZbm4Vgy8qB3
+3iTwXNCbCUqniwMrCw+1fbLTRMMPIvGwVnMErRmgi1iIT6l+NR+s/E4GIfjR8IR26NkwlT78IIx
liaVD9sV27eLeWMZ94qZiF/MVsOgQMcqNGGdsAtpjT4/37wiil1xcnXacz+kZVJxbNIB1bCxfzVr
qlOUN3mqRWX17cyOJDmqu5Txb4i2jJ1q64EHu7lFwwgzT6Zpix8qhNCl6VS+OTowkpqCFrThresA
SUPcgih5j/mCTUm5ogJjxxU7QQG50WwjHG9wrtyI2lnVR31uFIZkm9CBfqth9EvWJkg6E2z/C//d
3dOnZMHGgxgcbYcrGzQLX7cmxRpikoDuyE6GoWLmo6lqqBPrD/gxrnDv8e2oG9dLBHgQTYAYZyDc
PqlcaG5/PqymckHysnpKORX4Chor2LqKLePjCf6iWRo8SI8lOWimv+lMn0TR/M84Sy7pDuM4SQx0
OrBqeAN5W9JnlY7vCcB7azsGM/Jqr2rkABjE7pA8DCEhmKGmufrc+VlK9DVsogBUPxsPaOrlFxTe
T7DiVZN0JoVFe9YZrBLAigTb5TKIFCK65HDO91PKspnWTUXs43I1yf+kMfLT4rV4UIc8APUgFcTE
YChd5c8KABAlCvSG/vZ73QDk6noh+v/xKC+stBRZRK51XDZ1Eeok/QvM60GgLmbLebwu1Q9rcsVO
TWKota+zlSsxlwyzRi3PtEPGBN9XvlqI5XNKTvXmhVueArNy2UjA3DxqYUpq3TbdAknGhUYeuL8M
i+IRYFrKeb36uc1IDVOLO+NhTByr9sKgY0xXjQIlkb/N77qnogUIn1NMiyOIpiGykKH9WKpZL44+
bgE1t79v5EqO7GGmCHwxj+MnrJa9gkSKDfw8GQnyZvUAz9fkEZlyQMnp6wQcIOZKP4SFfpTknu+0
D9aC345Iu1pOF7dVeBpelcyjE8KD8gAByLk/Kvtl9DaVEjJIo6k+hccgxqeYUcOX3mSqDCYQWvUF
4eTZuC70zrQyTUp7Tkcud/1V26ama7Xjp0bvMuWCX3AQiTMb0kkLzOhYKjMCrxO7qWMOjO/311dQ
I8cEAZs8k19prxqyrisj9tKEX/ZWC/KDZbHZ3tc5BvVIr/wTKUWeuPVM6ezEI0WDIa1ud2ouVTE6
sFWg8/0QP/Zav430QYXvuHSmNTFPRqCt3qxLUlvP1l45vD4XNqgAzlwcVg/PNxXRK+8hscYAjfjX
8hDyw2OrHh/ld5Frfaaz/PT4l/GKNWNpAa3EkmAPSn0hNdqfNUZRLLb3Ed46U4QL+qhxXzJe8g0v
kD1SwN4eX9ZDQ1khx95HwDhiGqEfUoUl2aozFn566LBrdUdhXUqwEgk6xc7WJHn7+eQSEzkLM7iE
w5rNwF1/ZvGb9QxNTu6HXVQ7fbYvgIckokY/VWe0Uo1bRSfN8heosDeG4iLnZUCVSuuE+4xzi0tP
A4LCg8Ittbd62ai2yClc1j1CGUq+HQf/YQZB5jmYZU/uAUEsvC16TPPJrPFDUMq0B67+/HGF8I6x
UXIZD1w0/kYA6KDkSmc259+Nct+9A/dATE47MK3uq6kSzkk6FQay8GBgAk1I013/kgTGXdUfA0ze
BLeJI7a7j+1mU/5P41602kx/tCUNSoFiUWu5AKP785oj+TQsRdLHsybC+vaNBSaw28/4tsgS4J2k
X8Nl+laOeouInYZPKoikZMEk8ILTiP87r7krLR6awXVfyrzD7Ok2x9grUkZ/msIILbD3FV/tpBuE
4LxPfaOWGY+rSQfwNKYIGljQyGlvzXsw/z04luS3BP7tiCbqCkiQbPRrxdo3LnoYb9UixbMGijkw
hdhUkCsX/vDoyDMsPvTFz2gqae8FPqMyXwS/vSOHReNsRQjkjkLWpfzCdv6dlQDORhXagrZaX2wz
KUQY7lM6qOoKeTNyN9JikrUbQjSTeMlwfpq2MUAPodd9U+OeIZfU9aC2sjXgOWP1cAsLX4s+XTqU
bFV0A7SNjIPz8X6yAiS31imG7ut1yN9OUhXDGZAVwKFt+yQfNqdrNT4kXpkKcL/mbPG6bM0Vngwc
314WwKJ+ITfoZjxRc+MjUogoxTBATQ0zPqunZ7How4dgrCElylQsdrJUNPMcpOZt3QsqpnndgU3h
VG+jheg6U0B6kTzUtum8mQ08tImRxKE3W3xaST55Y/CcRQvgqQXcDh13cnGmaRs0RNyy7Ic+5Fk3
CL41+F//UAc66NSoafi+MfzxLJw9/VY7XgfxKtdBSTXDtfh5XmPwoPZHcdPtDk69kMT/eF3IjGGh
V4C4sQT4jLkZrZSZ2g/YKKOIvUGHSNgvKAlRp/Zp4k9fvN4l0KEVS3varzyWq+FT+xu9Gd61bXxf
K43kjYmBpigJPPYsPso9OtpePMKT+QOhEiUEXGzyJ4z8HbvmYSmNBaJ31yWTYaEQTj7QR6bd1rlp
f/JRuHiHcWB1HIZDPz5OqoT/D/GKHyBBqE7tF3U8RjavZEyuukongYy5txjfQsWhqlxljn2v4xUi
zRpz8oZ2qGqTUZ58jF0jRHELHzT60iEhrp08nOvvM6F/cjbNjJhq4fJng0eou7iDBd6EAgSoc2gl
EIja0840cMNoPflQbxCZrVtWqw+13QMKrZyrdo4APQU2Ip7i2uOIcgOk7wh2dyYdP5iMrToNNKBO
EJl315+KiZ1m94YQXELZu0Widhq7NK/w3Kqaeo/LCFPasGxZRsQ8TaMPVMGpRXwl8oZjiwEiZQ1m
o7l/i9aP3EqXYG3X0nAlrbJFO6ayfzj1LHra4nJQ6Ek6V0D/eii/+r59YgeE2IdzYnCy8l6ojKde
Unwi07TmZ+T3WpQmiaJyDiolxTnQk+YoDBNYGX3NUuTTNBBjUB8+JTCyeKy7xZrEGPqWs8lkExUP
Hfl6OBBNwdJtAnTcsFCKSKRmkOt2CoZJUpbv/DmSv5jPL35SuxhPdZJNkqeCuyfkOwWq+m+c7RDO
IIE1/hgL1bbKKnipaQ30JkL5T3lmwqjs8ekwYLxDODfAmaIrxD2IyuKzuEjE56qRVPgt9NLIGNCc
VOeYuajpdNF3rc/cF8JGXCFtAcJQgOXEcjeXPK+wwqNz4vJmmbNhxejIN7kCZkoZe5fRJnf5sY7G
U1X1WVInMYtR3jyK3jn8qqdlO2/qJiACVGJ2rirbOU1fKngujSOEmfVxxL3ct3oQJhfwuLtU5gyi
EbnCVXu+R70FqYpwbJicOuQScH4oq5s7FAfaYI+GL5sKd4884wa+Hy5MaxQq/fRWR5+nL/RckQlM
xMDIXWk0i0UEeAmaCRYWsX4KWnHN9uBXkFjs6rJMPTdhMNAT4Rv9x57BjltmSwgCZLBwNWL8ymHj
oW97PhnnN1OaByUG3AvbIweqjTn+PE3cXXpG3L9ouKu6VI6F8DSGeOMW1NEV6NegSgEJx23Pwqqj
Vl2A3AEv3BDw4//u0hom9znf6prfuLqF0pjpLqLEZZ6rjeIUN5B188VvnVnjmfaKc5GuOkw7yMqs
dWpJ1nA7hWSGRUTTCuzrrHa+27xEHaJJldUyui7DVqqXI11ZK8sVTU8u56gP6F3vdd7YZaNsKUHH
QbX7AAN3YzGOuiD7ZQbCv0zJZXRe9jn3XqHD48N30sIZ6IeLNI3WG0xDhuOrQVmbUEgfjtcmaCNU
DWrMJWFE1QVG0a0rjnIDJmhSQpCG0GEvl05D28cdY0nvReySLhcIRcxYJOeIDoyxypFqc+/cZb9Z
qo+WQaYhc6j/UNmmvAsiQcy91rCA1TRJzcU4z1hPs4CXQDZHX2TIYYtom3B2ItwWftOpl/OiVI+p
ZUT8Zk0DNemhIg/h0YISMfkd+5y0GLVqwurW2gPnHzFiDwXxQSXnwMb5LGccX+Sl4azaxMBklzOn
eNjDlvGStvDh01B31m9X6IuW7krT9jqNTMPwYXnlnIkkvJCfU86FrkvRbhcodyVd86wq2QxYsYM5
TQK8u9/8TrQU4JIeZcPdUZ4kyrVy6/fFgwVsxXfnb3ETuiSdd9ZKgc568QWSo8PaqOUcD4Hv5+9J
TUnzhs7VK8+LqJgJ9dCSJZuEEtIzqAxTWgtR0Isikp5Hpfbn5zzfNKKK1gQRffuTyV8driLFbloS
miYpe9JmpVdBLwH+OjwRc4ocMdtxM8+h7MplD4y+qCTX8Hovco7iefbtEA5UrZgxyIkREk46DXQW
VNMlifTlxVY4m4pM2NWMjmMaOcpd0ZvFxtkVJQzXZr7P8LPeINPtdDYvYj5lEp/vrxxMvg6y2ARF
HiESdPSNOfxlHVG6YSeH1f5TEPmYdKCHYSPWLk3BMl+FOD4rp2EnXwpXxoxVFSXEfusKDqik0ce7
RUeebyw8+Oi0iVm3lsL+dkkU58soNlTrgzxVu9TgFP5YIIrC9vCESNqi6LH9IvVyvnuvoigrx1uA
LqTDXI0ie08ll0QRmUIc97RN7wlmuMZGwHBI0ZpR0WlO6iR3FuUc2X6ca4RtmKjyw8u9ILFBlpGJ
sDkdSH0VHYCtyb2ITPQ35me95/VSWLLf5Yu1Du73zz1JkQjaDk2pwiOKwrzsHc9YwHLYU4h/j4QU
eOApBhYajI5CSaqdRlhZSAg4MFEbqpRLg4q1YNdhNgId8KsoKICQU0R7u4uhDa5rSKyFIJRx72hZ
nsEUeqf2l0HF47pwVsYDoJ1UYMHm8S5H99xg5DKZuWA5Vvp2K304V4pPD6RQe6RPsesKHQ7rPid+
CVTLtWWs+C/HYAg/YLs3vMRAt8l5ObYH8oTb9YEn1epwebhwqqjITKMRm7HNd/o2Vs6o4Qg9fwtM
+D6t5g6HB5EBlLkKHCkVOTR0e61Z1744bnNcoj3GobhE/3JcBh2+1T70TXzfgb+HlneCQJFHWDkZ
hzbBNzIw9rvhPkb87HOrCZCYxhQkE/zMN5IUQyzI3anF2K0SHfiNrAR0iLsOCqxjfb9njtbSKbBs
AHaHfig88mjyCln0MHFlmyZ8fsxLM7NrqJsD/dq6m7wBU2BGPxSED7m7aKE7en1cmUUA1CsKsokF
cjxMMeMEB9f+t+xP2KmmDsGGi7IkIe1TdA7bvR3koa/CIVXGHJrdyMVcRv4W0vJlpR691e+QNLZv
UVaVMNS3Cczjm+qrOmDJZ/gllIEXlgpxMynStF6qIVNrg3Id1fpAqxt76c+lVWVo5YS/dL/H0Ust
OddDwLCRlNrHT5Xj/8DcS4vF/Pjw+44udaanZU/qUACPI+g7pElzsYRaswx9VNAopJDMdDljmxFe
jj6fo1jciP8UliXAbIeYr5uo8/gaerDODJU7SORbSpl2qHMVfFGTR34nQH75ffigbbPt2n3QYyKd
wydU0SprXbafpIOV4ipfNsNXXtDZzt5i5k/FppXdOy3oXCgUmz8BrPjhpJSVL3png9SEaav4vXRS
1GrbvDLkNjUicNVN7OdWK/0OlIwAgCbFPaJCJUS/OlsFGpBD65ZIGjzaPMuiK5wmAoIE7ssJ9I+l
ggp/5s3fyJcCESdhh89F/f6AQzWPniM8MZDW8ovKqvHQzw+FkURofuBPEDmnD8nwa3ju4xWCM97W
pFz8cGmm8bM0wGwz9Q4ArtnmkJ1IJa0Bse72ausIBdp1MR51KHn6I1C08MYamEfHx6Te2CqtClYJ
m8NeN2JRpysV/ajgJbirQDJSLwBzpHPaLIRzU5ICeH9zWv1kAkGOjMGonNf3xusi9aOxwmgR7aXJ
BrIiKYukoauxddk4bpTqKwqp4QQ/tOLam9EVE3u8hU1XPHvqRd1Yv8YIi3bHF3ECetaCOXJUgDLR
BvkqfqQWevzy4Ib8Q0P0kBkAMFX0uW6qoEd0b4ewDpGSJgEpwLU1r1BBSg8XfR/AKC9liKh5zTo1
XPL+v1l7cqC3Vfp+Ko6xrr5bkJxBGs+M5M9cOzynR9Dl7ztSjbFe7x1sXYDNXZEaX7iPGtb7TA+h
obCZDoL3rJI8YmLf8XdPgFHnQK5O/wJ3uA3Vz1Y5azbaQtAnItqgckIRaEZQmuOUn1N8XjCDWL6O
3PkK+/9z5Lh9Al3Zhyl3R6503zK2lBkEifp+ISsSlBfOAijt0+OSg2cxCe/wMhWLmA3Mub1327ET
CqBaBd45zVv2uPwK4RfgUFIFaYl0Anl+KsRSMQYmekTmdZupmgXvjLQEBPzUsl5AsvMv7lXI8Qfs
xDFq9TlHMRJGi2akOkx0XZOV+7F8ChNtajLfFM1HLt7gUzks8b325hWmyHFiInskEyCNQyN+f4BB
VeNDO11NKBCQxW40HlZ/19diKBSr9cKLzvGgTkAUXGIHc839EcBC+2qOHkNEM0tajvoK1vInvjnE
b5jNHYpvFWmIssUmDLvK/mYpGMQr9Fo1/+1zwW0NkQEFZnHNDKaBkrY2kJxAq5nmlhp8iC8R6Wxu
fO2J09OZ1CTZgwkw9fT/2zIEtRgwfS8EEFNlWOiSivs0B3laRDGnCp69CxU2wTsLU6pubrqJO8g9
P6OmCSSdRvXZCkjUQz3v0+vTFjiceKbW7rPEyHPC84/mnTcZLUrh5K8V/tmNL+/H5w0K26HkwgR7
GlSHoZuwh/BanHMfhp07OKQwD38Vd03ltsTZ2s3y7BrOxSkY9fkX/nkHRIu6t13GBaUDo9mBQ4zE
BiKJa3biTMBYLSlT45VpvoeEXmgItNMs7JGCKlw1cV4UWHgLyKTP6SiUi3IbKeoZBD6LlumrSY0p
09wmkm1Icdd7AeiH5KaN6KMiwFqqXuZ9o15t6asoFy9TKwcK96ma7OQMRpsP/WJSWew1zepV4Yx4
pVUP4o1fdpSCDCl0kj+uYa7gWWiAVFJFaToHnAipgaP3ZnzuhWrMRH2LZyPEfoSlFRxKafkIJp0f
vWxayMl4Vhf3hEJJdVjsKb5BjnaPYTeJlFwjI738FXm36T3bsJV5NRXqcRygSGYRRoLXAXILOBpy
nuWZDgLH5xocSHBz/mQ0K1N3rRQPykiTMlioghskcLp7tqxPr+8TztTi3rDD27+0icnSX5pr+spb
ZWiNFQzSMMAG4A7MYG4zzZbQ/SDxTiz6J9FyHLG933WJoH6bDh8e1LGrBjyydBexSAFni1CHHm1/
LPoQzy+qkPNbgGbxjhw4klZa3261/v0lgUVqI+JUtG02H/yzORNSnE8wAZMjR3B2+MI0QtJu8ucg
ooerLeeizI8HCpRV7lNrrEZHwDqjW5TpuLjs3DBAVZOIA3kvFEmNJXPp4rwV3m0WDVgeLXLsc9pS
YTj0UujmYgnNbgfNTebYSs6HKi7/p7HbBlEGY1LA1SNkzxwg8nmLXhonaUlHaO8jEHy1B6nUKedo
FGEfKI/LieeX5zSsSJder0y5sbAPvHTcDKbLwMvie59GEb9gmxmUQSaIdgMYRues7U99qfdLnMb9
HayIXXybwa/6EHuJMpE6y4TKOHwfCJe9rrCrQXvBNoO/pM7I9txgW16kwhrePnBGJyv7hDaju+Z6
GTq3wxP9pVID6zOP2t3qmDNY27Q5D2FtCmb4uOExAutVER7tloAzi4LoWZNtNKDyz8UyyywRuSB6
FHgSQXzBHdxtg6x40SSyM/1VSFCvye0mGjPXgbRdzx64qgKnB5Y8nVgfk2Cys8szBn3L63dzDPvD
IYdI50rsuxZpV64D9QKD/eZWRo6UTLr5HDJvj+DzmvF3MyjuBZOIKgJ8d1nenD5VBpYopkVPb66D
tdoFuolI3CCqaFkAmsyoLLvinPjt1+7N5ZyB0mk42ljktleu5hIou+Qq0duDOpOHQsqR/H5X9Fo+
pBPQr+xotk0+vicya20cL39n1J7S+iHzlnR19yrTwdzhP7HXx9AyOQKME7aCVulwY4URukSWjZnx
oqSU/9lWx/g/GcsJmgpDetGM/zCHeOuNsVnAqa/JfteMuou4XbL7Ed3a/cWrzIj5Si2bwmvoxL9V
9MqbWIZt8WWn8hrpC3hjb1hezka9rsa+kSNu1+3el7RuFYNnBpi492+o422zwduxtzSP4oV/qh/K
Cw4PcoGjFlUavk6KgEsPaRwV1ThoNxpyRBcgQcmaBwJ+1nS4Sm06XSlxGgaALfGFUh8QWWREbxJY
msUlFKGSfJlhgdh+HtpQ+JKGK48ArdoHuPqo7HKyfZ9qx7/k9IvjgZ62Z8Pfn3sHAve2gc2bWoCH
oel9p8BhAF3W2p3BjETu7Uao+zDKsdl0nUbD+iQGNoBIk8O59fahmoxx0eYYE4WhyxGVVHRlH/5y
vUVeTFuQ3ijTrexlmUtIFgNhziy8o1FfDvWYayTBRgfP4YwHj5FO/WIocaPdxuUlWuMX0iM8Nt+s
oXfsQjghxnVLFDNgkiImnWmlpemvSZ2oxBWSuULPfNuwV8gxdjJwirB4rbP99a5WMKXqkCkAiOT0
0MCZhwkztfb8UobuoiogYPrQD6UvOBvKU0dJEnsqV4utoEd643OhA83D0eOaqF0zemrcTB42MzwV
D3P2dkHgsPFem/l3p5pmgTsVxUSGyR90c+GZSNNib1sNJTCQui5YD+mKOSvLywjGwuTQR2EnNg6m
lQS7624VxibrMf0exkWXNj6y/hsDAbxI+FmT7sPFS+zULKE24lMDz4xDUt76i+gTlwPMFc4Bw/RL
TX2SMCvdUOv0b4Gec5JEYCiHsPFPXk0FGjB1+PTCgT594VMh61yV7hn608mYU2hA8PFv9Pn60AOK
lGbD7iBP8gEA4VRrassWHXPHQT+kH6g8z9yj9tC0jl/5dj+hJEjTYptZUOqnGZuK9icshoaajXew
mpSEPIXHi/SSSJdutErAw2a5iJBqx517XRqMzGwfK9+jlAIMzOy88tk1VMtYKf777ckTJ11HfiwM
LYbQOFxbRM/FCt8Ow6Pq+6utUD31gqaw2ALSwSwgDtOrsT0JWj4ai5CrdPmpt4Pdz8h/liBBbf49
FxTIpbD8dkyEsOGQjt+OcRddWtPU/NhBBjKnawkCfcfF+xgl8nO3djHFNKS1DJYrF0a1rR44MAwP
f3IquvU3CqlVE01Ztx+i3I5eZu2OEJ/ZgYtoS+qvuDw7Af/KWKM/nunIiZFrh/VvFbSyW0ZqXD8d
nBqxyEO90RJx0tIU+L5EVa1JiL/EeUUdMLma4h9d+gKkG7b0H0bk1axqzRycdArSywGS+2Njoplq
EHLuAH6OLWs12Sya8Zz2WY0E1Vf50i0QZ4MIJT/o8iO0HFu0UIZ7IP6mo/oUx9sxPUIkzU0qlPmK
LnC3WuX2sNRLZsgFyiMqdWK8fJlHrheHDn+F1R2FY1qi9dgjCGMZ/5hrsgm4SwzP59FAzvQ87KWu
BExjL3vR+I8ItJlcoe1a6BBqsyYl2iFaBCyx0ELzNPKNUBVYi/zuHny99ulAzLLvEqcIX7z9qYWl
zF1cVIv6/cJMJxtMuBVjDTZQagcV4mi+X7NEeeXYLKWRQObavaMU3xsfc//3kdMHKdTlCXZyfFr4
r9JlwfjUfKgw5dYKcBnbTz1mPJNPxhW6pPCcd/uqeDRUuCAPqo8mcPJv/ar1Qyr0m7nzQe0i60iL
z4qz90NcA4os2+QS/zEJ3s4k+LlV8azQPYzzILTmKU23G7iloqoCPeRi53kfoWiiC16EO27zeJ+F
6JptZfHtZMTEofzj0OPK/W0KdzQHdswbsjsnezWPZHeLHyU5/gaic7yZmY4BjCBPfdzYLEwqE6rf
D0yRfft/2Fn/sjt8vvIC5ljHDhaJRex5ckQlP6AzgMemJ4c/VBNPTHhv//dNG8XkAhCUJAnw2DdL
Rs+d5Nlrn7hVvZqSfgCFQKILXYwhz6j7CB8tD5G4IbAuhHPyGnRo3V/Ydgc45sk7FiHVJhKDIUiH
6+BiU8gfh5/tTuJ31UPApOR1LaDpUm4oOwkH0spIJLQeK+y65LzC2neOcldZ2OSFep3k5qBXtgpo
P0JYBDYGlJd1ZgBYLZgBRirisK7dOqygoWJgEbZgEFLjGqdIT6wxhhuzkhTXVMj+ESYASrv0mgHU
SwUwimEIXn14CWlh+n8cZ5SLSl1TorHJHAGLtv1ofq8hFL1tocXgVcJQABe8tPCGY1S4O7H2gOhH
EbyvXxlJnf8OMkdWRa76rDgBkTrmsj9MYdErRDKdowSvZqOBVH3rpSHBpLKncrxTJA9VLH0uNzmC
4PkH//RIctMlvvzPiQQ5Asup9/f5uqpndCrLzd8sHrpZ6qGto4f8FbdVyJtXCl72s40GtF6TjgWj
YpL6bNaUHGemserYihPCSUL7SOx1X2JgMuzmtkYlbFuLcFtQLvlDq8qSuFzNS1atBMN0KoH0VVwf
oKxrRDycBz4r8EcRRwuv2p3dTQbN2ZfpE/QeL7tlmmxaF6IVmOS9/maueTL2gFT0HpdS+mKevhNV
LiTUnXgIhRdhnpbsgAV2ogAXsyS/rCOkhLyBo6KumPY952qJU2jvNfqgTmabY9/Bzv3wpgo9yMBA
Jr3KyqCNu7tYoRCWgxYLJSdAm+KrQfC9lFOMzLuDnef+xQAU7qwBeT873cggiu8geveMDwxdCcDx
79gLmhLvfjDcelmtENi6orwY7g9zQV0oPFkTCqr4f4Ajo5S3o0vTo8tog6xLeHSCDimlbub3WbuS
U3ywyEAdpSqbqJ5l9zYrTFlOIUZ5GN/WHcs1efQTcx0DKbc3T+2jajyaNJVUlIJJbeXiN3YWfEpk
Hu0W6Ahb3nQ7Y0GlmlMCEBv4rPxtqexiPZW0X6bB2aHwfA+ZsXF9tHYoJd0lgt6F54jmWt705GgZ
wRt0tDuT1smMjxfOjRClcc5HcgJufmFEMwDPFG7j0bwor71WTxCtEZl9DjD6qbxkwkXThekgZ3Dl
GP36zD4zZ+i+Mhj7Ab5uXJBn0H9hNQbw4/G6tGskRVLscGjMQFycb7xzrW+vEbvH7wdS/VGn1V6N
rfuwMA2GZaja8aU18m8VWd5D+b7takDsJkpNfGRWejgK6PyK+yg+drVxMSVo/WEmeT0FNzWWANJF
/n0TN+VOLyjynoM+EDSfePsWf7cmT3s/J5bANhNWowZYuR5lM3zjpbRM3IkF4fCTJcLV+EyTFwfT
9OY8orXturZ/KrXgNBHaPp0AOlVXWXTcW2NTrCLC3FMCltWZUXB6nDg3gpycgQldptQLfVCRj9bm
3gLEBoBQPz3YL4BO5y0tfg98eZGtwfM+Yy6fH+BuimLT8YeWq9GZdl4WJfsVx5Q/sK8IXuwpCzJ6
B1TC4iYxkJCduDNZizxIBPoeiO/05YuwZUlwjr5XqR0HXDFPO7FOAEeoy91S6ZFnllCkUhpK3swz
znsoOsecd6p+iTeksq6ANYRWV0ar1/dgbpzypnjxa19bmwH4PNBYKnK2WLUy6Aa0SznRvPJ163+1
OybJM2fBle1OmE4xqTGNhWg+zG2Bjc+GsJRMMK6ixikz+8R4TFnBJPbKzIs389AXKaI2zViAGWFM
DVa9rzkt9EYvoQe0WbNdzwxcekDztoTMDYjrwIeoNtMsK9lTs+Kch5vtXpW+OddFe4U7GMEg/IpP
7SNrS2/kHzs3SvO5Yy3Z7MdPPxc054KtQiYLKDpFcUW48kFrbYuqa7xMvigH9UEvxo8aQm7rLr+x
Bw/pLGqUw1+6EgIPMfC5hj4HydIOeNQf1pPQBQNDTcMU54GCd6g1csbuil2rQVgpq3HbyP+elnl+
tsa6y3Cs9A6txr3uxjca8z6/mR/rVEO0QRYoDLK3NVH0f/nOfg4w28uji5P1LGzXMmfQ7kbvZGzy
s2KSXYIhWBD9DqJBGRo0gv2xNr3nZ7ivZrDdA7GP3pR5rxYNP8PEy4lF81kgMEHVrEYu5IJy/DIk
4F7n1qaFEgM/hZ5E3y0pt0sIb4PMhWxGepGDtdDTSKfsxxUbE19dBN/KMII12uvx6Tqn7ovtcenp
kKUo2TVqOW1LvCLbIFO6MwPrAY5qtVu7pLJIk6G1EZCJkz1bq5N8NXdWycZAk4iqed0s+44twiN4
Kfmm+scm4GJ3tqMzk/4rZZ7tK6aufzHJ8hSYRVuQwOmRd/4fw5z2L7n/pQTJcg9XwyyzlhkQeSyF
8CBNzh3TQnxM2VEBSoayCJNtwfM7pY0W+BtvaFIZEdMZ81J2UkMZQ/A+G8a6OeIEqtTP9hZchg88
HYuz5HSFYu12tjQOayAbmKG0T1Amyi8LlNddQQXr/lw40VuxEDI1nGxZEQfROsAsU3aLxwczNgjc
j4Iz4AKznWNc4o6LyzxyuAVwzEtCDTk/rLmDU5317dcl8GIo6GVd+iS8JU2ixaSbGHg3filP+fIV
SvT906p09b38DLL9oXOr+TpogQwsQWgen73KsKUjiG4pFfDunc5phTrqVXEKCleP75XLiD+5q8DE
Qtkw9G/0UrzL5ar75kjfjX6TDSxsiJcd08GmVeC6MZLI5Nfop4oAAYDZv6eRt8vbewav2oKWrMvu
j6XblmiCeZAKA9m6jduWCHrzUOXfXjlk8OpOGZklqvT1BMAYa8/TFanh81cw081orIq6nIxLAiwQ
XiL+t5hkJcEMnCck2v63H0t1fjqbYCtZEoXvQ+sZrHQ68/R/I2P4V+06kI3QwCksSkfCxWrzctTt
2wroJ6MsdePlwpkFPlRiJzYZkzCTKONnPum5YQsrh/9sDVDrewuZ1IEMVchcoILfnMRJUV3gPH9w
NsMbplE9pRGOgqFsO8yJufoVjF2cEiOA1aPDYK5xw1l2YDoLtvEKq+Zb7XyAPa3RgGVEoNik9CQu
koFTFgJXJXfqtaq4b+CoIoeOsul/NwOry8yXf/O5oqm6GD3V7/ro+dxFarANI9OYgzD+tO4pnGOg
wrZJfI9OJ9Osuuly5PEd9+hDSbz2LqeVIIG7DwmfJhOgj6w7cFxQj//O8L+N8YzC6ZoUMFk2J6jD
x41pl0wq/a31eBYIZqp4Xja2gUYaVQGTfrxn1kBSuHUW0XAKtkTqkyYFtTNRrTRKcfVmXRV2kOHU
puKCH1jGSMl+09AOyIpA2FdY6VjUSfhY3RGlZebq7Yz1STUojTczqjLYT/te44Lpmit/9YZmFRpM
2zf/NSWhiC82FC5zER+hzE9B9eB2d7lO+Rs2dUBtd0ApSMVDFdp+LV+Uj2cGYpLYx+Ug7CmcdA2P
MGYIj+FFeUMSyplUpyvIOB4b3hQNOPbCOHsrQZIFVx8gur7umK7DNUA9TfM1/iJWig4IiXmlHl39
W6ji2I0P7PBisBzyE5yfS5Q9LFbbyvhovN470pKBjTWCdbJN8uNw9EOiUC5T+zXkWijOiIkGk23V
qx6rjyPrh/pFIXwlAvkmdPTLc23vlD4N2kbnD7fAeq0fjOjMeCeuOgl/T5HTmYM4j7hbKE374xMf
gjskiW/Iqe2CMtsZMp75fp1w5r/P98OR9J1cRq3QFGhyNF9Wset24M9d70X08ft5KDlHOuX41F5g
neQ3et68+zkVzYv0YPGb01QwwB4laUoSK/2J6WpWZPA9Af0Re9rTAASlZTuYtcAtQgAig94Fkz/f
LM8ZC57ra8VAEFWrkkVd8GUJGW2oSg/6IIuKUg0imDsMgd1ssqW2V0Tou8N9MR0yTy7oEgriwSFJ
QUMMsOLD9uqeOPqc7UtlsAoJWnvwHEtvLFYmTCITCQ6ethAoDUxgI++O7qfWZLbHwNTrxRlSJFsH
S5nYEeTmt6ryMOGMddu81qivf88mKRLbPoB8fRG0zrOREO3NvSxDiaa8D/XbueqAZpXvbV8ln/L4
EGmEkEqkBgQQQNcLoxCcwaohbf2hcFStdNAR5dAX2qVcsB/GkiAH6lEF0Xce0HkdSdV9iil9nwWx
nuc0IC+/7Lpy4e31VvBhhNKbuerE3VsVYDTtMQcDIAQwjBIf7wi8SQjGpwtWnKOBqNGFdBCs45eF
6sh43m5+ca9gzHLHz5iJ3GgJtpZeM9+f093EZNvzmG0L6ohjA82roOFv7tlTbS5pacg83T/uNkLC
WHC0iNJMwvlLycssoXkc0yLuH6ouxShLbggukdAcbk93Dt9qYPdY28w/pzyYSvNUg0Uw32La8XTE
rguMurFaIBNgBfcHmnjwC8us9ToWXzSWicQ3AW8q681kcvYkzCkpH+1udVmOAnbpksWMijMAUnQE
XnAizd6FlQDcM2/uhlFZD3XHCUzpvOUrAOQpgO7HBzDYhliIhA4RyH1ASWLsOfUmJ42KZW6pQvCn
z48WDF9SCMkMU9NAc+L40HB3Q4p5jaTMO4uJZ/fGGbR4/WGiGHycjRIyq+KOGvOT+4X1neCHzZFz
ubnkuYA9rGWti1xqFMeSrWRHWEsAaYOJjSeyovM4WARyfGphCkdArF0eCtQt1Sl/aPSTtlMSBuB5
ZdHcDoAvKM1x4o4xOr8RuImVgqSRtLX19vV3KvOpEPUjeFaSoLnW+rufexWYZ5zlyh4OGfH9cUvW
LW3oD3eFnyeE21xR0Rwuzs7EADTznBv7KCP7qfVfaQ7q8b6LmotNEfkwbfM98fF59CSeDC7/4ZcV
rg6KhdILuZ7EVu2+XS5B3XheLaedvClnrXG0Hc9yIo7xI4KtqzYOR/ixjFFzEg+KApz6kwEUbMvP
Ofn1FzaNgO8sBq4iySDw/4rIuzutBj0MGUtWsznDJv3/y9MV5C23jRmRycdUJ8uW6xZQe4ndh+UG
uxxGG7UHRChORss3Ct8D0glWzGU4qJaie2hUt2Bz/ytcJFTDwuWGOJyEnmvWxsCoKRZW3I5rlhxR
+Td9b7QhdkBrt4dwdo0Vd29Em0ZsGu4EfUcZDPl9Ie43TuPAbXLCS9QftHLHFS915GN++tKa/r7Y
89sgpP2zOiPjDW3Mel007rHGMjmY2TY24+Lz8E/TRgAZ7uSys17vWXOmsgzySXXRnz0PR49jAlyX
XMupZRbLN6kFmZezzXdHCGxWoBiC3/dDEW9t5jzdcbobRFq1EmX2pJOL5B4Hv/8lN0wTvRFVGGZI
xVSn6fpYoUgYSNMth+B0t6rddEjN5yH/dBIQsSr+94j83hZvk2fTRaRwGjyMCFRilOKlzdfighfo
GrOaV6uqMLZfg9cfKMWSuEheryLkWgsmJA1MpU+xo2Ahezl8/DKg4NF6v+YwxiUpUWbrnbjwT+iv
0ygJOv7g7Wdcmo48grS+Vtv/nRItktJr595z8gVBTOACBuR4NaBLKd9SQQkp+gIeF0C/+GHozFko
hHw8mYMhxfhxGXfZN9hjirRLxzUZqbV8ISoCoGF/RmYJ3h6YxLs/D0CEKmIuiecDExMJFFAMp7uC
jYtsquHHX9VTCo8KN6JgapScAXN8DMgXmPCT7f+A8FvcV7ocoOzEiIPpDJze2H7qfZG/cC4KnYBo
IOt8FNOLEVvY/urzj/5T7o6j1EqcR/CF8n/N+/bkOOPNsW0W0AbGuE3+G9z3euXOeRc7/UJsEm6H
EyAMKjD1ZSwYgPjdS2sU6YI75mlR7KGCNbsEpvLDbyeOgEqh+3pb/sa7rS5vKxrR/FD0ilP3In/t
C8rkgxljEG19wdG3lgR9sRIy3lA6mEBz/dOMqaq15c9aVcv1WDSc/GWJ6T9mzQhzqjacy9DQEjzO
0+3rymIAfX1VPmemIOHYiLZ2lmreG0MZ83qnRwhVv0pY8dJXqv9Cno+GkBhhhuCqZyl34idseKTi
DoQ+PDgjIeZJPZSRNpdS0Zatb5yvADfh/a7/yGD/dltdVnW7i3dGIIRFMdTOJLfHZEnlLVnfFcyD
XhPJ9zCJYO71cRnnYtDDN79E/5kWtx5yDEvljk7Op1F0OZ+p9nsYPxtZ26z6h8FD7gM1WRlNRpCF
HHyrcY3q+cJ5fgUIlaDVVvST05tIROH/PwrWW1jhjJqe899Pr2+82kgFhSM4bq7uT/upWDOZ+f1A
Qi3TDnk4XE0PQFNDwy38mn6+416Wad8yfXvZuoInacxAnOE/eK7lBSzIofahpyOPnrt2UF5tuF+2
TLDOaLrUh9dABPsWS3a2275y5W1/E9/IWPFIOTNSFcH/3CeulCVD8brfRrLfpF1RypTiZBeXRBn5
FDJfS4klhAIHJOh2BNNC243oQkof1WE1yce52vC6JAJrhcJNqYeOduG/EuKmB9zIVkZAUWjI3Yx4
eID8284LkaAl5SHkeh3IL4c24qZXwOpKs0qHdxI6LcBt8ZkT1S5uYXQ9QWO/TICIJIFUG5fgyNPy
Qwx0+cexQevvxvJS5vR/yxnfyNC3LQ0YVGSi9yh6HfAHLzxYp/AjcuYSbPLAJFYbqMsMSA9au/K6
2/SbSWwyqfn612RitBIhdBTk8p3r2gyy/P+S25KNEn/xW64v6GqdWVnntskEfxexhlEqUgV26G+C
Tm4Uq/Nbc8ToJH5ScAY7GAfCnVsP574meuc4RIBdW4R1F4pvfzDE8BWr7wsWQ7wsPvFuFOpHJuKP
q+fl4oDIqZ7MWKyTrKxkqMsvjYbSpdtfFnl6YiVPRbIVsXmM+9LbsVQOagdBKdKJvovtzh1HGpNX
rOC1fHDcLdCYiDSxbOS+hJhvk0ItAzZVUY0aoo6zzZNmlOEzb2+7djVjJmar6Nss38EtusiWSaeS
e3AMiQVtQq+5oTOKMHpXicG6ErCLQpO0GVG/TF8656tasNnAaDSRmFdzEuCEZYFOeepGuTAKts1r
lLHCQ+nLHEYHpkQ/RPoEO0pVeGL6N3Cz6eIpi1H5mvgJ3JhF351GiK0eYal6M20lnc/2BFkn7ydF
mYXSD7ytU1igBdCagQIVVdRFoUuld6qZu6++1j2+fyAWfN+ydCR8mUN8WP6nn/2dieCS2xeSBMhb
vYi+TI7BirFmh+gRoONAznPicIkTLkGg8LT2QTQYg1rQ0CFnCGNaPMEm+9ljJMCBjD1AmnWNJQxC
e11tnY24jk0khjaLRM1j+VhPtLfKsKQvSSXhmgNpXHLfWrZhrxpWjNfwLC1yairlK9vTDX4hSCmG
u3qpY1JPamUQeAdoEQQ/6WrzU4GSCw50rCGpmr5Cj3PjZjcduh1C8SsfeSbTmCmw3MPUdDvyogRU
VZHRSO9V1A5MpBa4BIfHx3p84j4dfaoPWLT2JqZKGbAr1mglxKLCOmS1XO7ElDY+NbmTG1SY5gZr
q7kiClTaZhyWtLbSApnlbxKDHsZ2rqaSy7xNHPM/cN21ZgMANVXACYMgGY0EyzbXKBYNalQHL6V+
GFyehHNQ83fNsCIz+hg7dCy9rLmMX8aREsbqTnPZ9iQ5eefibMLQEZLTxmROgN+XCZuCjvw0kZuj
Ajfrxx/Z0Sf7DBgpLyfA3W+/j/A1nHOJf3zNrPyg1PmrlH4h5/uYUFUVFW7zBYn8FmuRtVSjOFss
V+QPN+s+o2IjFkWNLkKBBjv2Kl/n87sgNH0WJCm47SkhMhJ+txsYnCwox+Nu7T0CvCKCKJyVssg+
7KwkLTcuzpM3R49O+6Ey38swOS0zy6rqgMxRiWqgZ8ciC7Sqt0pbt06n4masS5j0z59ywPbmuBqH
Dm08v5Cj9lEeUIZN/TxDpyAY2leE7WzcZG8HiB1eGCl5YJRccmE3VGwvdaeqG6v9mgPTLXTREVNA
V0QxWNmix7DWRTzGnRVMtfsVPDcSc+GUFDkUhx9+bqvGIVHQT4wkLRhq87BcxH40nrLkFcFrDeR6
hfLdXPIne3wNtAPRDwdzpQrpVWkbPRwTPSu5LxIyQzTkfVWpoBxWTujKmXqwAIANMPoJh3gTiwTi
luzU/y9p9UgJUA9pTzvVv71o24dZgfdRzv8+XWM5VAGk6McZThAIj+0xPJ8KsrFuwyly7klpPSe9
qVB9w5gVYUxE43C+1HWGusd+obelmf7o5HtlR3IgolN3jswpuv3aoJmFkQ6Rt8KWu0rhU2Dyb8pV
KdjGl7tpGozVyK1y0dAwlVV1kvShuAHPxPlW+XiJ19aoTod3RS5xw+TC7pR576X1NMqWHVLwM2M8
9aa3wK5RKg1Ytvo35S65R5dRwJ0bmdR37v3aTdYD3QxJ/hIAbS/+rOqM+d0c8scU468YaJrxhQLe
G2siID3VPz1xR5BGqncMEisnU6RMjT7IkMJ7aAyntPp0qI/KLjGhzKDA6q32Z8I5pcTx1N4AdGvz
e+QUrvO0et5jQxXl61sLMWrcblUcn7qmNlZzopUdsIb+BJu9PDxmZYXZB172ZtvPiCdYdb63O1mF
yXoHGbBPTVO9TElkaZFDukdT4S+eapAfKhWljaTq7sX5rqlOZNFbXSDh0LqWJc2WVGcGeAggGUXx
fU3ry/PF9rXhUCv2j00h86dxr6cQ5Ptnk4eY7qvOL78iQynEViqhOhWex06KAlteRRhglYC65QFl
IKSnK4m9W0PnYiyucAcmrEXyGaEcvbCq/khEeHofrn+zUZj08lKIOKkoUXgJLaMrMgkR/quac/v2
IqVCdGvtTfxUmnRjVJbjCzRnlmuVFH1lVrA3p3NjlFbFhIBy4bJ/rmZxsv3+OZGlNjuLHFcGuawZ
/hVSyV1xc/TsKDEdHJwyYpLPqr1YI2fY4lBxlHUi4x00x+VjJyq0T9F8XcLKeWsJi07MKfXH6efW
ynokqT4R1TgZmodmrcuEGsVzB1Af5g6GNEBNuMmrhaOkq2jTSuoK2iUaNMPJw0h+63pVl0oX0Fl9
/GymfWc34h1DJfqaQYqVjB5aGKkP3xijaEfsPvBxAav0juh0GiYdauP3eTUr6j0XrH8aVieikC5m
fYObYgWwhpuEMZ6dei1zS8KKk0sLKzdKt2cvZcGzeGmL1BcJFq4ail7XMvuLP72/fjqLTP6tVcO7
sDUm+6g78zWJ28OePFHiVUr1+IJ3bfeLa1hlqhKndw3ruiMqB8rSPTcgEycNQ8X3xArfJ47/ymLQ
FGv7pHVyRSyzZhp/78OAayPUi1M2BEe2mcMWNvEt1yaAVtX8qNr//ors9h0JN2pJ5QWRXrY5WHmh
4GdC7pE26wHYQhOmhYHuH0C2adjEh/iE7EAKBdAr5AEcFnEJOmqfdToXROmxdVvOQxdPj7juckrn
R/pbqxQVVlAGNqI3F2W9HRrPolS0DHPWZBIycI97jxb4ZaKgE+AQOgs7aqBPbegl7N5b4vn6jlJT
FdAnSHku8tuHR/b9UvLNmBwMK7Sv7gWZdvH9GdRngwGUSiPrh6kR9vVmoQXhAj8gcXQMAM96aHRA
WKb/0oZXmvQFex7UngkQLMRpqA1ceg/41oeKJKK2hol36O1dDV6ey4S9H7uIEh0osX0uM3wPGEra
GGmmiEijwn8TV9VgKA8pjX0j0UHC5NUaF9gz4O5taDfzKRrhR08rQtSBTCJrGeLUQ3cWTpuQvw61
NserTYGl6R56bKpaf6c9iTtsINhQnMI96mIeQLdEl6ZHC75FDpdEY3LmcQ5YDfK2onLxlT9fpl1M
Lqet5xm0WLG8hJXSi8Ju0jliK4wbe07txuh5grorP8tCNGZ9wZ9i7kyz18J1WXnmXVQa1Y5GfrHU
52d8pt8CojrgwONl+sGJCoTj5sctzViUqF5Q0XGHWSZmT5eIyIlkTwBS64/lkF+NVxvxXh3Oit2p
ba3RzDqBhYSpYwEXyO89foxkSwXJ/CPfdhMEq5sje8g9lZ9Jtu6k8l00bj1aqQIf/IQBA82IIDjb
GL2peNxvtI+cvfYdvA1/nPeg1kfOBdvbQ4taQrpVBfwcUniDsOIzGMo1L0V/QmXfmSZa0cHK9Q1g
9ncnjhga8Cb6kqrYIGl6to9miTTvYzhGuXhYrstH0hxyrX0JA67vPT9c3EmuP6s3EDiB1ZlQ4FlU
Ro8duFQSk3BYUMXeSmO7NkblQvakXJcxspnv5v98rLoOzH1O7xO7/kT4lyILjS1nMu/IBMNhHbNK
QDSFTQuh7iizJiXOB4aqysLwsV+bGoKP14RU1pTMdEjMGHmtEfASY/KcHtH9XjTajohdk+4QFEpj
qzF/iX4P36grnse9jVUs5uYkpON+rMzwQ0tzC4yi0JI68/0hjnEoqQZX8phRnPeEtcdJCVrSSZCG
Izh0c12nf5a3CcMmdFuziNrmR0uzs+ch8EDYo5wwekrLgwKPwH7WndDiNPc11ejtmJ7f0aFRXdSL
ZECMeyB4bVp+GJnbETYdqRZ9kIRN++Ny0fj1r5U+MN4xqKvQLNFodTBYiLFCx73xsESCf/7tNA1f
OqpCdsz8OTBrZXpYpoZe6w5vYDpFaDJ2vVig5/BZk0kVY19lvjpOoWOAurAR7BRF6ieCHSIchddv
BnMlhV0hKbcYp90SRSQAQXScjQ4Qcbsv/n/X0COh/RsDoLKlPorEpqaIJyo8uxgvr9A8HEZnTcJ7
nxtd4k7dKYfI2LsWJp/PJ93gadl1xBfOWVvOQgTX7wFRUm0W2k9f9H6+MpIo5+XJIU6Hc0d1WzEf
/MFxM1TYCIchGM6VFDzqPk0EXe+04qj+f6LwlgVG8psK9UNOi2tU0X9CUpLAcbQ1gKZD0S8gVBaj
w50UxJmwBbb94VhWzVK8J2doNo0LN4zOs+7e+h9qovVVGE+QSO60KFZaPeZ3p7iBuxxsxitCspEl
OhVMJiVNvicyxw0z4fylzUyoO0cVBLfmSNY9LDTuKbjsBIc0gnqOCs7ZHUnG+Ufb/uKfoH9Ik7II
F83m4Jnb61cI3Ee7FCi3LGTpcndT+ih9epWP6TMwTQIxoUGBFYlzLmN7kI/xlo6hdv9bAjW0e55u
lIm6tJ1A5s4h8T5xGBDhVeBBdYGrpur0ctA3H0aWUSSoQ6e3+Wjui1fKOXhxRsIlFIS0K1sur64F
ugEybzRtYj9rx9Q+VQnNmf6gP/57zu6OF1sVOI7Jzi6FcpBLBGrWXHPmzF0DP7zAsPW8CCUOLcDT
sYiaUeuob+anchiKlWAITSHHwCwTZ1XaapKMBprBJb/bo6G1ag5sxXfFzXepFfM8HVc4EtMa9vUn
PalXHPuJVBq6CTHg1U8SZAl1hEYXIQCDjGVQwceD731e0fBuTY/TxgPHv5RL0d+RJZc/JIDDu6jM
nO6nvINAevwVG9/hshuK0TFa72SHjRZhWS+4lXaBMSzn04peMqNNYeQi/SLP8wt2PNPrZozpyCob
GbgclYL/r6msUMJCYzRM+vgkWYfOCnTfuWHE9bxQPMd6s/I2H27Ood8YxyB8b6cSvhTy+y4ftb0q
IWhN9OBaZg1q2415cjtBm3l6aCkvaOel0so+YQiOwx27/nHZ+ejQ4iJ0OStyQikHKgOhMMo+u8nr
abkoleGA0rLrp+9GdNs5mnz1for+qPoJW1dliPcBNrh0uHp6nhuDjNXVqFffnUavDCpBtghKPP8S
1mMR6MOksNllv10QYAVzI6FlJnNrt6MIyOvLc2coJRDcBLYCoqjsJg45I0tGj5mRqK5lvV05UGNJ
v2kEn1to8p1iJdwHdWLseo6cmrJ1oe9PPtiXcusjvipHInaaHuoBD0m4UAx80XyRz02bVA2dfNti
0QGo0/sd8sfqCfzPZ9Ca2iXlBq38jUiC4v5opBf1QeoEZAoXV/5Lezbt6+2ERNEWjaRrBbBm1vKq
Lm0rPkjSAHYcE6yxPYonFtX/bUXwBOXlXeX0sH42E8aVdZvxg+eWz7IA4Yd1FCRm2bQCiTnDTE4e
3JNUYzrr0ssAfo2hNUjy0YJHJ/+9jABfhdSYhMPuVLIHsUeBpge8YBzOV1f1kMJKXaYhpiTwUpdk
UrRV/Q3IkfNYEZ0IajOBv2c8AHsCI/PRlUxWeVTv5/LNZV+scesuxxAx1vYGIoL+kUrsr01XXZJ8
IDDU6ZTHt+eOb8myUAD9YhR7pyN+oZZQb3DAffeDZQsmujdJrqEz+iKSs3UplFrhklKKdAkRXaxv
99bC02np3f5JmDBKxwO/OZpRa9mqXOBKeh8Zpvq33eS7ivCE8rhM0jWjXUT01pyJw7+In10r3ly0
RNsVkr4IOSLhB5QVKKxZhnpnbM6JkZGdQgG/kaqzMmMN3QJ4A2CfxDA3gc/ulkE7icp9p7dALxpZ
yiWjD/Go9cokB5dcIXgbC/SygMBNNwii1k0O6T/CINW7noc0lH2apmBxpYl+EUQCQILPmfp5XzgP
9OO1sKmU/TabXf+KxY5X9S6zQojQJ5cNyB7OSdheQ8UT4hC0h3MNILjsmO5nCbn2nCjuCkdbdJes
UzdSSQHFPHEShd5pGhqmYapUetIr5g0G8O/H4BgeBHokMTU9QIwdkOMREnv5ev+siv85aCOR5dvU
+D8inMPPKDoNlONAb38WaNDnvhC2bpTRyGMgRiAJ+7BHwyiWVICM9S2uSuHwP6petw4RhN8Xwq/4
xUAlgfXsAhtrOw2QblzG6clFznEJPmXIBSV+ttL38UPn4qTMYWay0VvI5SZ0eOucU5i3hbw+I4H6
U4PNgPCP05lDvoPgESdJxHI6PRfH9RTwUPV5UWz8RiqvNCVwNz6Ek863sAm49Lxk7TKaVwDxNbT4
YzjCMy1cQUU6uvkfx2NK8Eu4KP9FARCo8GUnWhAGg6Zqj4lkljnX/RIllv4X7KRAKbsaj04BCixd
+3k4tSr11RglxEtkg5RfrqP2WxjhJUeE/YlN3e46AIhdnhbBSPNP0jfeBJT435fEgAF1pOpB6lNu
MqIZ2VZheVM0dzcWpmpTAVNBrVQuorVze7JTRIx+IJbsaKLXIERx3FBK2FvFedbzygFmwscRa/oO
5HvOSZi729fVnCQX2T3c7+Eeg/LoxCFoTiKF/CqBVeCUHQ97ASCkLB/vLCSTEfQXU5xmMBlnabUL
bNdvrlX7vrAHwV6CeHD6cgH9C5+sSHIkyfUqfgUeE1rXZCH9oeLLEyVKXXchuTocps6ZuKFCRJXm
BbCUxRlgZ2pbzwIrB3dvK3L79QIBYQBGCxGsm+UGIlJM50ECuTC5BAyqgxwS3X37bcYwLX9tZrMl
w029YFu/m/v3/puoajnoNbkjxWRsF3IjX5zVqRjUwrvk7qA7EWiRDyW7XUhmu/V8QjGCzLCDgErr
7F+QLodwz/GfwL9A3pXK7QtoIKnYKOZsUFjEFEV9LMcAKvSNc70rMLdGXeCO+krH6v5rvLgdMXqP
8GPSPU4QQEvSqpVovBZAXpDY/vUx11AePb2gKeHPYe5r11AkBhf6MlHmF+KAtHz8+6O1cg3AGosM
8P56a6kyLZTvwSvV5ALvqt0mD2IB0UmBB5211vi4twjCATRuBNCRgTwUCQ+oO6K+Rb3MG5/9svUX
KxftFqqO5whWrZGUM3IyBoxyvlj2JiYShmg/RsPijJFy7anmPeQ+mPhJDaOszbGTY16QMYbDT72y
mmALFlO4EkcIbbHnafnngGKo9rfTrgl+lVOqWyRceyiuIxC9PycyI50Kds3QZb1VXhnpH3Ok+FPM
vbQrMxuEHV+fHboxq+sUTAIFXau0X6gILcQqORTbSqnknmP6RJF9BEJLNdvVPX4eaU73WleSIXG0
6qrK1pEZeIcGWZBOGOkcnpnHJBAU80srxmO9TwW4ltlGXS+nX4bWyjXRqJafg+UCi63N/af6aRcE
urbebSd0WwJniOgUk/CPtpp9VAdRiQF+9f1hR0j73orMIWfEca3SDI9yq1LxaxBRSawBMV7VDdKS
Dz4YLEX5IcIq1LWvfqwaKei3+dtRM/QHng80rwklIJpfhY4U16B7y+ykjAiZckxsieN+gmGmiG+U
674VjudykbTg1is71ZMrQyFal3hhh9XzcoGq29KU2YIyx4dFpdsvLCsnPb4CL7Rqx2SwiEUSqWSy
+j4BgMaGXwy0mWJNk1YW4q336MBGS4XUQ2o6XJHNZ5wUyWkX5SNZna8qRgM35y3EWnulIjRKdDuN
/pcybZVdItTxQ7WFxu56A38WXvTQVmpUFSSB03Km6cbj+sPhDz21rgmdpF7am5/uqsKmPNtrLl9Q
ycAEllAEhhjcJfInBs+uH+e6kxlrkiTUuixHI8jefPg13IKhDNoHHos1xK9p/k66BBl2X/D7EVe/
u7ysBbKmAnYHe0z8XPpeW5fBssxLHyWBc4mnlZDzsPZC5gRBCpnSr1AR/L81I/aAROfmAWZ6NfGN
N4n4KL/8k9wsKIAA+9a4phW98UnHBdGc3nuNbPo3RiGvhzQCx5eg3wRqfGCUvTYcuVcft2HnjOm1
WAGSY/83ERORvwk2nlznmXSnGAdE5dPVBBBXGB8oUlFKwHD0O9y0fq6LK4fmjhgdYGgg/LpFnr10
m7IaDlgrNkpd+LYTJjPN+/yxVWHAxjXS0ozaoknap6a0DhEuLY9l65QqilGS6zf+dm4plrUvzG9O
zlITcto4wOMQGEQG5GnbmNKD/yzr9X5Xa5Oi9HD0XVSm738NQ7HAp3pdAKMqC4BOs2CKq4ic58vX
SitUhXr6AQtD6o53d35Q8hpRTWeuUHUWudQu0b/tCzYgHe4I/Tb5IoasVx9epsAU0iFAJyoUPajs
gi1yWi+aFxAaMzUDWTXwulC3IjtGyLi4kzLuYvXg6UUxQhkCbec2uhTYOxJr/iJ0Ehvi97fv8tX4
YZBHm6x/W4rb6sL5ExwrRPd2ZlD4v9Fx3PRyOFXhyCF2JZCj7pvb3TimUHFFmCcvQlGFPkZWOI92
gysE7EG8BWqxyR5sPRUCPr+lFWeglP0qFcSxAMm+V8NFZx2+zw77QOmY9Joj5/xHFs4vPSZn7ah4
09lgXydHIhlcpo1klwJGaVf1LHqmxtpV+UYuEUCyc1AZr2IdcgpBBY26XmJ31l6SI+GMRb3HANVq
XNqsTukzuFMoIlqP8FYMOzOoORcaJcnp3nUCOTgNQ1o2u3z46U4Wg5/zh6IfjMoXa21zE8phvkKr
qAYQSbtJruKo/5ZnZyvnmnKt4TTwMhSo3JXIGThGs0PpJk1yeVHD7OV7CbPBGh3h5Yjiy+2ouaux
OrJo0vJIPfBDiEfsuA/6IDXJO+SMkAlVy9/HcUpmWU1Jwfvk7uWAQpTEVaZC0OTUFYeJM2vPMWIi
n45WugYnO+ceXpnYk7WijQr0LBPVEWunkpKYO69xhyTgpJto5R/2XGqZYWZLo6Jyyimv4bEWeriR
IyOfYR6GQPcnMuBgkjydKYMH1GgfuLvMWumOTDfcahBEMasT0UH/CyFp5EZYTANXpf+C9AiABOEa
igA+NcLrIWCxSNQNyyM9F5xhs1O6YdGrYOPtH4Qk2UvmX/mIrbzrctmK+w5VLl/Ec/I2U3wJiLYu
aRoJql4dmtwpG6S3QRUb+3XnIDAYZH5JFy/0IsW+K6W7VA1KBnu0MatWmsnRlWumAZquw+YM7rxc
QIyvm/EYZXnFG1r9R1tGgWvxdMDFCeyoIbrPjA8n7W7IXmSgb68Rt0WVA8n0oV9ztxWxMKxRrR77
Ikv+80jt/iJQKXWOJ2MLUwxkF6c6xJ4KNl2dE3AuDhSiV8E+WFLhVcOSxSg00lgDbb66rs3sNEZM
dcgVvn68QMlHqF5OxbW+3fgttLuMjTldzhzLegSv2flQzYgZUWer6uluAYhcbrktjJgvs3GrwFRy
p7ppKwn/SOk3Tes/f9RWXz9IEBX8BM4eqWGzf9j25LZDp3aEvRSSoPiL0loPce5tZYJq3Di1WOti
rx9t1fXYtffvjW1Atlj+tw/i6CMxPRD/T741a+8fcv5ucd0tKVQ8+TfC6uA8kDtNk/x4aJXwDpZ0
0jEL9wCMdBttVQX1/OeQfe8PYLUCh476FF98BLfKGrYLdc3/zkpWJMGblx1P/4AdsQyOxtiOoyZ5
PvKMeg2nCK9wuhKrv7+l1thHNljAyYLJg0kUZNC+Sqc21v4z4RFwZ0bGJ3ueb4UOIb291527Yjw9
9N83st54fqEsW77qPMeXxZBPfVu2jrp8BfGDfJ+/NjAfwl527nsw7/Hlbz9swu5kj5REnuw+i9uG
GkAT3B/N0eZhzzZ5+x/bR93KRkyxoD7o4LDPt9c1x3RcnRKzLeM/vAtFkSSw7KEKumCsSei/V/sG
EHdpsBOQHAZHXIem3nh1bHoIZzYaL/sqFTR6ytOuLbC69rotkrhRX85xSdh4HJ/wh1hILcChaMNu
nFQOuhMTQUrN1BxwGpHu3AgJTd6+wfx/GoCLdTGuF956Sjt0vTCEVcp/phXvWxgwL5WKz2Iic723
Ku/BuLiFs5+YNxxRW+kWp7dvUvZukAhmIq2c6xzEo/QUDZNprZpHIfPBA4zOZxk8+4mWlYwB4Kww
5HdRZ9nPba/Ipj4NvC095xHJie2b99vNT2q4si422A/ATwOejojrHW6a9kC//wqt1iSpfRdtdc8y
PC4XcKYMfCfwV5D3oPGVrgNz+mUfhwMx9VMwLmO55qbICSJIrm4b9xSVOVimnHa4VX/pCg6IZsyw
zL4d8km2UgHPEWzGigRBs37iKiG/T3ucLfx4K4Ef4Dhawe3y3e+znIBpvnO1LeWwbUzjqdGRgfju
Fvs1MmDpVL8Y1peKRCQt2i4dFCCvJY+8TtHq/HjNBz3rV4JDoUwM8E3OeU8t7OhdFGSkn4U7pxZf
yLCR65kegJWpGBfNM85MRGhRmaQ4Y5qVH8RfBvK6PDAP6LP0IGv2EzvfjznBWIwF7lWAXY6cq8DD
R2VxqeWpE+RbAL+iTcBxCgJvR1Z5wNIzAAGkiKFigSAWouK3P/ZMJlDm1J19LPqpDPnTyZJ22gNL
c2rmvTmeWNp9Or7tXzsgwLjdcS6ynDLaz7KN5gnz6A8OZKZQJ/EZ2qW6ZoNHDjoGjJuSyc0P6hMt
nFvy8FUPdesihYSZqP9rCqqC2PjZiRmsUcfpXgEKve8T1YT/jpQReVavfsihkBYaZHVxL+CLzXGR
uKEPVb3pf7AiGJprMBt5qA/L/FjIx95JyrwvJW2KgPsxEF7+ja5TGwwYr2GOOBwOF/97/wrv+yep
STsc7Ica5k5ncGEmdx3BS1pEXmlpUFaMI1mixBXjqb0Wzi2PjQPDEvDFcApEM801EKZzIT2Vw3UC
9Q5JEmLhnjCNF+vCeb6SKW3dkJk+dV+3/GqSaQAbk9oHuhePXSnP6Qs9D136A2nIqyY7pYIoT6KQ
Th8egfgvDSU8IdR9dTUVG6gO5MEP8zjxW/d2zU8GSQ4js2MnjX5bz2XUBVbCOWr5d3T7ukKt0J0U
SOxfTOgSRiaW1nyth8pZECLVta/vPg55a9QIbYP7RkADLZFpbvqf+L/3rE9IcPHb897KpbZcQs2t
tyMLa2hMsT7DEA6D28553wUX/ddheMJl5Hkh4eBErnH8XHcULVtVFgtqmZxS0zJJ66pvuzSTJ8SQ
56d7G5crxU55hEZ+lTe6+FUKvq3yVm2Pz+r2A8Go6UZme3DotSwjaeYBga4TNn2TuCWRm8ceC6vm
4uG7Og4YaBH3FAMSIFMVneftMpakTEeRtPsCX/opMZFu6pjg48j2uI/+blOvtMwRxm88IXqnUSl6
lqWT/PgOUX2pq8f+RvPSpHU2re3Zs3l/WE5jDkcn8C6LULEnNnhtMQxqPJzcoYPYzQWrzfJp3tkR
zpxuaMkEN7+261eWWXi0JlOuLS9Pqpw0CK1PAEbcRCmju1DpCS3uwOSr4PN3jrA+UJ5oHfIi9bQe
abXlklOsrW+MmB+VILWyEsl8lWDx3+ckhHwu3kNQ/4uVI124yUl3S+5zSjOc6PtY8oCOm6wnhUUA
BA8wI5PFXWzT4o9w5zfJQ8QyzdAjssmBSLFfMNahVOiE3yL7gTi+QgZ/9JGx1H2Wkasm0hWCyqlW
8nYOdt9VmRJ3Yvf/ORZvyXmoE/fyAb/H3WDTNtHA9jkebvpmKHbJovc538vp8KM3MIjF59TAR59t
T+6XDKyAho5ke6Kt9IQusySBNhGwG6FityRu5GrZzKv5XDfC9AqyDuA7RAWiI8mOj41hnc3sIOd5
FsKFliYYH6LMYmuiVHK/29fRGMl3ISpb63wP8aoUfOOpP/9EGqp09ubMYdWCe3lM41ks7Day9uEc
ZehnjMMOKWVslasNShNdwtFhh4B5L54gIPAmJ47TFpr7UjEGv6iOIslA5t0as4kmAXKuh7PNc7BJ
Oe3d8o1f3dUQwp/yowdsmrhboVI1fnPSprTFZM9fr2M3VoGJ/cVLgiqz/e/HxbP4Tr2k28bp3IQt
Ri14RlxNqYbXCa0AQQTwPrXCfDRehQky4t405yCWpiIeuLMHRFmNQC2lnIK+pARcN8yAcnVkjLTl
WxG5gR9AdHE+7MlNhQ2Xd53cz7YHcLuh58PqaSP9l+zRCIFT/kfjIrCJDZE9+c4K+5ANSPjSKEhA
iZnUb6coxH9b8HoQPqylh7y24maiOo/4vm/uCsvFxNaWKp29vXxzOQPR4loJpw30aM4PFPVrMKvp
p6Cnrxu5vcF3IvrUzEnDIll3/3MyrN6wZZRdrnR8+fyu/EZY2JbpI9RNjW+5Jg6TuUyKmE7blP3l
AY4khyx6Jew3y/XhSdiihBqgVF0yzUwIIhg1sknmUUEdidCMoeB8Lhbz4OO9Z99/+nHQg4pKWsTZ
EAVqh/HA/4APUaXu7GG3/OW7aHG6XHf03tD34t5eO+BkRAxWa+Fm9rYJDKjc3fUb3OQbQ3bdPAFK
mRIlnvtOYq8YKd6B4+t/WrUJmXU/U3Q2NbCKvaz8LBW6K9W6+AKHcyWFvQLa6KyLSvpNbhIHSHSr
+q8TCAegZdj5lBDZ2EoFKTayng0jdNjCVKO+xRD+lSOtfp2pFQiipnOrzJZUot0NzdipayA8dxiQ
7KBZ8mfmNS6OiO/H574kSVq63wcvAPfd+OLJ3+EgFo90PxBFOIkUkpErIxno0fak6dHvF2Y1JVEO
Wq/IuAqX49CYxZGf4dtE/ZKkJtSOq0HIRuxDPlpcQxHJKgTT2lbABOD67GK2b5cPuJmEUqNMh57Z
DAwWY2VBqrijsmf/UjN+8rmscvDC9a8N9s3NPW95uFryxxPH+LaWdVUaS4lYtdRTZxfcMQGtkHsC
u/N+zpqriHu6pFPjq3WPnheMjyRmiK8FZm+Ueyhu9iYcZg+gxnVrtfQ3nbqHvs6Hedg6FGj2eRbg
UBDvc8Z3Jo6yRFYk+xmHGxbrtVUmAwoZDwMZpnl3lfgE6uJ3e35y4tRt9ZkOJf/qiS63TB3Sq64k
ldchHPI0KKJioE8KrXZWxzzNzxa6paImHhC9ySn1+E95gKixxRRkqx5XgiGvjdSw/4U1BTwlUwLY
0Eu42W/mb1857zGG55TVWOwFouuRVOyGrkRFdNXd0/SHPljaoAGMaiXfdY/znUm7jnB4MZ7Ywhaf
IkMe/MGARBN14ruWVtfTGMqNnwegyp7uGMe0AWNB9N1JQkZhAdBKZUsYCypGtTP7Bp8wp0aqqt/4
HiiFfiPgulzGNXT2H+/h6oZgdO/oEDO9rkRGrHJmKfWDf1t/lneFUSpRwjrT7aV0nXw6ENKMb12w
su+A9Ij7UPzberwrHo0fZJ+r8hOYs6K/Jf0tUZYbKCG3tbS7k+Pl0CJJ3AWGUbyafDdxZS8srSJR
Pp1YFWZEzSkWC9kdEmBf00w2LDWl/2K03rP4VLuxYw3xpKXR6E28B9uFL/9gYx2TQCo79YCd1L0q
GfBTvxpbPOdfxv3FUnDHRBNCTa2wzcS4+qWuNV1MJq0h2fNudu/SejIgo0rONEwgDgaFyv+1nQ0o
+AFzWQFeFre4y0ZR7LzuoEsNMNOWlB1CeywTUM1XMNmzLOT8CclQQYsv/wY8bkEyiQueQBO29s6x
FxrYidiaPnmWKP5MV7EyGgc23KbxWQQVHk5eoqHBTRB+5yxNwXuZQ4cx2olBZSv4aoeOa9grLsAV
hX4vUcdiPTTeWkbaPVofwmkK/N6Df1bdskEwdoLC1xw6DoOi2foGVMjYZBQ0Dx5OTiy8GhJSv67D
5AMhvEaBrw/Q3ezfld1QP5hG1f9q+U2+OmkYaVZO7E6zj2Q8FktnoAV9Ev+EYz8COh6AvgHzMlOX
tbOz/70Lk85o3ME9KppOHkW6q2agt87vROsjvSmYudr84w4DKu+qDRan29iZIfzDnwvm5CPtE49R
d788bbIIbrwFHWyuzEs6OOQaDrZRHXgfGil9eZ2dJFSlaVJnq5rkE105C10km2rB/eUjuI4M3rUx
YL9O5s26X8lYI9v5v133YoCh6NRhMRoClLALdKoo8nRITLg938c5UFuQISmQiUX09/mjlyywv9tm
wUk+WWwPsqG023leWwDZtTiRy5MlHq7kPx+aNghxh2bg3/J6v8LifhdqrxYbROSRkr1nPS0GCJ8R
AGPkj7l9y6PyRh8Sd+0cIP9Yybs+rmtP9BrxNfTIzhjX0j3e6xuVRDHyt6j5QiYTeQqQ3VSBSXKX
cqDl6Ck/pqu3VSDUfaED13IukWs9TPau0gD4LVH+TeT2sImVnhKUyPHPdomeKejGGNK1nLJIIA+H
mcN4DN2oIYC8NWyCq0ibKO9Kk6N+vXu8+RU+pSCo4DC2LWyD0uSnpzD0s+Ypr3TKYkTBGFde9ge1
vTOJSiZU0V1H11QjOrreonwlw0Ln1+aXqCyAwzxwfhkOyu8FRlHIHqfAosYNls66GLFwmsGvtS/m
w407N3CjwGhUN229SD3HYUAdYW63VKNPeUTmzChBbSQbcy5WoHxwqCi5h2TxwLMwohL6+UWWtvUL
0IeuchlYm/aOgLhW2xpG4mX0gAyYUCOrrns7ZrmxyASWOtC/FwMq/XRDomPaXJMzoUpTLm/5KW3h
5LTD8c7J7OgnGwUPkhDJsRop66UhLncuSx/WiAXPvuLtHNsVxQiynujtBiZ13OmFUQTmiSmp5pxo
wR/ArVlobipK+nji2kNlHYBtHi4FyBNZazQrZpvA86u41z9wR53X48CdtCEl8iHa3/oM5FMn+BwZ
P+9l5/YUpHLC5i2sWdz4SY7E2KT3G2B0TXNFPIF9QADJ69EMXdqANeulLOTIIx0Y4BFh69vwyNWI
ulpwgsXYINZ1dFBNMQwNuw7eBdO8LffH7q9wGVaq2/TnsTazLGZCMs12WP4TYpnK0Jb/IDRcpwOf
zKJhL7a4wvKTGmjAsR7pngBRfIMHpi944qnV+o44Ciru4/GeyC8yEDMOEbSxCFy+LxDmFx2jc5Pd
7r62L9MQyV1v381FKz+ZrIOuCBbFkedB0uLs6uyWBw1tK1wJ9LoP5lEnl7ahJlSaHwSkZQWXLtx+
fceJkGBRaSKgawZ9qJ6WhQWP7Bk/rEDwIEJuxhlIPL9T2uTomcfqKJG2JFBXjBA617BWjGb1VB2j
2CZPdj0ufORINnr9edBVrVdqfxcZevY+ridF+LICXA+AudGxnsBIPSoE5FciusohYnrbdeFoe4F1
EMd3HsFr2ZZxp76Uflb4y6Z6T2ebd9Qs/Km6i5QR/GT1l31wEWIUVbYyNVb6jj46pq9Zrq2SYo4O
zctXOlUCHyKCykb9sNs6EDTlJFc4M/K+L4VL6VPDw+WH+djfwuGDy1Rakt67rtSSzRVs8HiBwyqJ
FfdUVUJEULRV9R8s3iC3GAUfWMwdkvrOqXLLIfxGhepliQDbJZQWhDnd0SEy7zQl7DvONAnddUGh
6nm/lVQt10/PdEAU40pT3ONXtF/HUofGo6nkgiysSUIZyItTB6ixx/4e8qHEgu1LtRE7qj2XNZYt
EArnvJOJj/OMzWG2TXa63Pz6xg32DMsQA3vfE8ONmGz4aG76fndzOxmympBZT+PwJxCGXkuLVm5i
jOw3Z1Uu20M/qq4I8gNO88NxhzKhDjKmca6zI6qwe52w92ASlhosBQOXhQY7Iuu2aaSYIslsn7GL
CsiCoFdkDWyffYf0ZeS44zK5wWl6Y2CflZ/PW7VAyegsc7wwnclNj5EY3rRhNWkEt0lKO5Qxq8KM
+hoUNyA4IjtwHIfz/ym+/S5qWP4Mtld95vb9pHiRhE/XlxRyIajKlF7joxtmMh8ApBa7ti2rdNKS
r/tva04x2lfBZ5gSIpb59zDtmeiUA8pA2kIul11BVPKeZFbqw2jWb6507wpVt/h6D+c487LwG4b3
ZMlOGzbFNefoNPgCS6oBREssl1FnLuPsg8H2rI6G1DtWvV6ITbspUFeYz8mpj9q1UC8Ne6DhwXyB
C2grDFDVanYbG4ss+boZY2ktJS2YEgKViQsYUvYo3nUQNuuItLRxskzYMOYe13J8YS+PVHLUBswh
tZQcM2hRAd2udYByN2ql8DErA2EcetMVD6h5cdndxjxZAII9L/6j1UyNZ5pEQSCd+hd/5sd/k5V0
6I1dJpqZUu57hkj+DM3SIdk86GqbGr7t5qimhB5Lu/IhGMAvVk8DwJR4oUiecbJ2kDwT7ZUXwyAW
7xFPeFq6+hBC72VMQnROVV6AdEJ0yNhiwE4yaXSYzknP/TFNx5nP/mh9oDUenkoLjIjvfMC26eaL
kwY6RQS46j5NKwBki0atvvKsFvYDaRiAimMxnTBr2EgF83nGsQ0cmDsMeVFeTwEpwzDGto71RD1a
RyhNQmJKuPFRLP3RXNXCdtwgnMhATHcZX3W/ULK0QnLDGv//mac9/vaqENU7X7AR8kySc8uzxlvs
uS7aueeno/vI1gE1Rj0rT7/7bew03aRQwdXbZv82ruyAhaYfo2OVBmyzwdxtBwUhz6iFUEu70Rj/
lQmhTESnkfj8tET08bb4qx+5rR36qdQ4yoNlWINkSe0aj0hPLstRA130aPTALLyakUbAvBlLugku
JnnVO3gApjeHgPEtb0+QY1sFpU6IO7m53kFgXSa0vGRnsl4O/iQ3ZOAD14FVNHNiwj8LlD7oJDk0
IpgEnPBXDKF+mmS6BdvAazwuPJ7CAudkp4ZqysFJSuCF13a7h/539cBfUssEMaF3poOgorNnAoYf
a/UFJ3wQPY2XC1VRFXHJhHAhCsxg6V+7aNMeQ5HsOLu3tsoAwfZXtK3FUdzTQ7RZIV4N6mRcCVvo
oiXcm6ryZa0u0nVX21r2SkvxoKjwqyNM+AQzWHE7DvF7cxOQo4K/0ogzAr3EqHw5m9B7IcKNgqQy
xH+YUxWr+hfTy5/s/JnCsYrhqzMLegDHfd8NI1dYxcFzU5ngC+2hbL+iARpi+i6d4NRdDmibdrEh
2MpwYkTgCARIFRpAm1NnTo/0tUiZWmbFIpPu1ilKzRAA2oRwu13uYs8D2bwC+Fr4EqDBaRiEU3c0
tN6IWI6WejR/hyxtcaSwTh0EnEaYtMOup2FIaGkyWm/aMtChC927NORED934vFZ2J9TrpWOhXAJ7
YvYUPwwpx23JU4x6AWRuj66f7jMkuw4hbLcAYh2A+lw+WePDG1d/r1AnDHRZ+jpxOBJg18FwN66R
WL1jynVqgUQSfP/4LKLqvxEvxctOZEwnbGvD2+VCwk3dhQ6XPO/n39wKt67PZV7MmZ3xrYEbjQ8/
jgAbIQXlAMAVXYlK3UNaldpYEqbMYqjOeg2sLaOmEOcMp8E4yVz0HYC+y5I3d1x1FwR9Vsl8PWiz
bxDDUK0+dmLESWMSA8Wsuh2O/Im3zcoggj7hUGzFAe9pt5OaX76dB/aSRWsb36vjuOmdz6C1caZJ
IwQkuQ76Jbk+JwUTbqOLft8mxo9NYQA5U6g2loCV6lcUIbyuXb0jSqeohn4bfO1adi0bZc2NNk/3
6EEEl35Rpx+wVPBnQRdY/YkiqfXKsuxl1+aYrL9Fgz5Y++jK+i+fh7ubxikhXBCUTM+QnuEqVK+R
rR+Is3MXH4yYx5SDLxQnHgeAT/0/LJYF8AdqT21XjHaRPR9qZ5llapWS/Db2lMrhVIPqGFfXeadR
beRXUj2JzE4Cr9/Y8JmSSO209IgcagSQCfiBIEEmlkJbgEyQd4oXHJXNWIEP92OQy1gloeHR+mr1
W9gmyqQHTK6g1z1oLwMSrfBfIDpN9Y4elOVJ49Dz8v3xnTDuV+zC8xvLkk1yE+X+59/QPviEbmTN
wuVyKiaJla7iu6nNpYSCPuvIzuP/aBEukWphOuMO1phpHo8e1jrtxh0LqOvjskQfA+KXkN7BXJwu
BdRISyJ2kB7rF0cvLOQEZZSqaFC/78Qt8XrDHiU7Uf0xgJHC+Gzb9y5i4a0HKLPfuhr4RXXzPA6H
viiLcr6eNu7ewdXqxhp6FlE/k2ytwe/AxxOjY6efIAZscuLgL/Wyg8tTD8oZbSuevVIg0gGt3TG5
cwEA8u/DAFOkj5qVpMj9/zdChh4H+V0w0LoFonMIoi8X7FSTB/Wvd4KC2E5eZdeIq1uCBEQe9wPV
bmZcGMNmQdrpK1gjFzxOws8B6mt8fGDVaF6uzvxYa1FmihaUaPV3uS74lPebff5ITjDJh1JvLgd2
ElqunRLkp1iPhwzYD0MeS0xigFveX4mTJlaWxZdwj16asZ3zDZgR7aEjtRRTa7uhK7nfV5R2ILVi
ol5KV8XuitNL6eK1eylJKRH34BfXJrSK+WUlZBHF4wMyfQ8Mr9IMtXaRURrrCmKpvbE1e+8bBirj
YJW3vnr6qTtm/6O3fiEEJIzkMP+KNlkbmgacumMopb2/HX13Qy65D6bEqrsrA7yXT/gve4paILQq
bofO1tRtsE4q3tL9Z4j4slXtUcAyk0NHTTxfjCX5eGY+/1YID6Psl2LeEpZmCiFaV30Sp71chm/P
fWFXjvgIhmoZZYrm3sjwNP1dJNuyCHTgGZaHrETpJXARPvxeQQtCMtp8MLQUsOXYlr845Mexz+pS
jGtpJTCm+0dqyZabXb6ByMPwZ1ALOEPUR4AJb2dOXagEoFtHW0SbktqFAKbJlkpvBoidFBVHn7b6
w9eiTeHtnMal7ahNgJ8/X7uF4A+iSv8y4iHOVxH9fX44V43NUGnInS2ajIG0ehfA7as3z5p9NJQP
nlFwoeqUQJwMitiIjB8MjWgBLMmYN7RtJdHFavK19LYv4l7BkrcHdaYswHQWJ6CbodAwiQnfPhDE
bJcvzM59+wxhT/6/jECTtiucYdxoD/H7zLthsJ7/oQZzUjTVoSLcc632UpdhSgfIRqMCGuIpOo2E
rp4h3LWmqXKvRu/jFxZr9KohfQraimXvopzxKxDRYF8CUtC5nnYb/KOHLpFDwC3RN/2/EatYvcSc
57aM7ZPNclZ9Isn4lkaVHlfjsH1Qn/1xrNOLiWyRSTyteUDpi9GJb5o38z+hYzL09EHokb4n5QcX
ZfjVLUMnL1uuIjc0lwQfNHHWt3oHgZrE5xLWnmleYT8uzolLWetE0U/tK9fcQMfNo9yaJ24LiuJ6
U7w4rXY9Wtu/qvtOnnxJlyy1Z8cjdYm096kYE2juxQkq99bsK40D6ScWxeqr32N/Jw/IlmUBSnbw
KKF6yIKqsj5NIAmqtO/CtM7KugaKWJsAPoGN2CvDBiqV+6Kzb3VVAQbMfYUab8tqJn4VCBf18A15
pIi5n4h/KBcz0IAfByjA8/WqjMM/NfrZylTvI1bsXNjY1qgjUqryGQufAZH+H0ViXvbNERYGdUlq
6IgxN/tz502Z+eiMnfeLLYwfLMrUpKr9hwH12PFaJKYDN3yK6YwYhV3mz1dZb+/ylytaNb37Bzgp
Cs9jnf+cWsRLmgWB+yEou02ZAegkU8WD89DjTV+OY0AXn6hs92dw0pbjlG10eU5IQfGy522RR4Wd
8DeXcc8gKhkxGFSuicxyVW0OG2SL+f86shY/aNbDmJxkn51xkXRp0GS+b40BOyrQRMSmlzFNV+CX
sTwEwqIdZ6RgmSRvZiukfkpf5lxVREsdqLrfnRla2ITkUhuNb1kEWEZwmeqirwmnCt2QaYBrndSn
3FNjR2NW5wuzb8HLiFk4/u8jBUqJQ1vWnESoLWy3UH9e0GiYqCMyLwYlZdq4mX1uILP6AGMCXIDP
EYQTiMR/q5emN4bR4822XwvJRl81b2F+UbY9hNIdzsTlzUYzRSxv+dPvrcNtSg+wZmFZXSeQ2SI9
hzMmwL5+BKIMV0HQjUII0LxbyR94zovNjzsDOMI/pdwRVDWXAL9aAD9oCS7bkc8rXx6mqeRdlyp0
i+mv4FsKVJNqb3fPk+p+9yrAbKr1PRXaqw3KtmMJ/BaRYBNWxxSIBHBk92RkIcR3nYsSkarowQxl
o7kw35lTXWI/+IE/5CNzJA8EVwi9Cqj1G7fWcONMao5QQmm0V3YQi72n4KHXOx1EDhNv/Hw2l2Xp
OMv3O/5lU1Ck9QGPyKiGNuCkgpW9ncLMjIBkwX/8Oh5j9TX6zAGxQd7UPCX3i+G4XsO22O1X7gyO
gEVzpY+nGDXIBu5dJM/uUxzFoSCqbe75Azy8VVMzmhvNMK6N/DSrq7lXKVFwe43wY9xUr8a16LOC
F/lWU5whLmBQQSXM2NF69p60eKUiI1KdVfATNYH9RVzLY81zPibHYCmq3tjtkthqCsrQRioHmwIh
QkHctWx6ZO4SqeBQ7vAKSwLiAblADEv8bgtL0tyvCOL8NPdE9CpA0/O7HTrKTb8W4KpVX3OJQSOl
F7g9IuLUB30oC/7r6zrhqrR+cwrglfne4R/iesxeZoA65GjKC/654OS507qhnHf+G+XwmtyIgW/k
Obvx/KV2Hms8xmfXaM4mjRklkUpEY1sFfNQZx/3eHXJiACM5td63o6rQ4WCTnIIzY/8Hlm14aIkD
0ZDsG0PUV/D2YUCKotMbLvYsFq7Kz5/KuM0Kttrpw6/mKVzLu0ZFJ3aNsAwRrO3pRNjOcNjMqMzg
BJ6p5X7lEehePYrnB2LBuubVns3GwxQjjywel0ecnqlhgLM73+6NEcUiLPzVQAwq+CIiKrxcj/Dz
qxcxlywp9LqoiGq9uhSmkLnmOjFcPm+qxM+z+hDvZOKHnPuq2cr7SjgLX+CW72y4PrlsPKnS6yt3
cvdGd3VFE4ft7rlKgDB6alIDp6jGcJjP7Kd3GzfjLQKAA14Z2sbuGmoMXMBJFiXXIRlIhFFAOJa0
ONzkzUIyf+j7krEpSQLZQcH7eFTtBwWaGfmczlNuagBzJkmbfa42pFLkh48vzHNeEGBj/brIiKmQ
Oi/uS7G3PqNtSQMzWNMhTEabbJ6x6O/P+REkUGWi5K05Cyhe4l8yk89dJaJ4o0xVxdfzLqj91Vue
OXRkn0O/xBEyfmAoTa37/KlL3uc6RzBZdag0hwm3UX6rO16e1zJyZZ10dpfvQ0N48q9wYjLfOqst
O9w664EnzX4QT0iOv1uNO61I8GMnRJwG85l/hdptvMJiSZYRgXQyxRdpgEYdxiAnMKaHJblJxGCy
lX39F2RyGTfiNvAF8KPiHZqMimf1PBBC7fXK4heaLLt9Y+srdll+v+eQFC+cVA0tmfrR9RJ60do6
bEWRf9/MjmVDKEsYFgTQJyhGLJU7WcUbAXzSXBGjY0sOO+G+3ue0EDKQzYO6kkocUkYjgWSueh5e
sxI5uRKp/MD5TPzA+AnD4mLYvd8XtSYKbcj5j5+KkGcz2HBT/HfzXvwYh2bUw5SBwLhsRFISltgs
4LbWjbyQQaKoRFL01uo+AvSB9xdIeI/hANEUQSgt8jnmFym5Tcnlw9VbX7dNFWk+7WsGUwBDd5kw
VXArQszcC49iDzxxBy/265tKYWgHZ51QZVjVk6cJFkbeh2r1THyImERXTwYmG7uEokYvUP3HCGL/
N7IrDIWvKPYm+l4c6+jTnKfZoQ0TLTtbY//Of7FBLq459T5xLf/GMg1krROBVp2S2GSnQ6jU+5tE
mBPbRRfF4XhdFo9egefB+/IWp+84PnEh7o7v3wOmeo/CzvvArJZU+f/QplfwLeccBcDqyygojOBt
hCAnLuQae3dnHE032HRt5oiI/H7exdX5RiktCK4tTOB50sFEwMYUypJdXjQyh82AnJx6bdEFqVnR
ndr/oJZ6T6t7cDjQWypmeDkBb73phehzur9SBlu6G9ENEEgO9qAgukPa4kv02RdgGp0zbGqQlLwc
Id4jN3TxIHPp9k+X2Q/11xWYse1XVNJUSQWCbT2gQxFPwsVKlRzfHpmJhpHY8xXZXMgcTWqG0dD5
D6cx3Jl64SzDmClsisFWL84oiGfd39000zWKCj23LwB0IqE/yMp1gQ6O4++p5/cMlg2gpDd7vBdY
rAthHych+JFxk39FG3xIxyXSOcfVEB8c5yZVqVZ6GHM4uKyy5sCSKwJ9biG+WNvW//ogvbTNvmZG
jQ2ucrF03kGtLGKi5xwmocDKquN8uQF1H1MqMPpdaeDqtXPGy3kO54qRuRnfvvIypZlRmW5Ex7x/
YOD8Phb4DD0zJHtbrF6ygUqvWscJK7RLV6RED+YWvUgEsLb4yC/BpLAKQ/NplNOSrKQ8RNmODI54
zFzNzxQB/NAoC/FjJLi+1nI8Z8yGI/PcSG7JEgjDpMg0oL3Z/SWpXCSEtNnIlwikX1w0neDBgPxW
Of2OGSyE6pr4LlC3UFSwjPHjJqvVKyNApTwwPPeiQ+5YX3ZvYnPp/1UHhAiQnA23yQyHKJUIPomr
E6zvJu9PEpT1CfyMSf5SW2EUSAwojnfV+GwB7eOdjyjtwOqgOpV7tqoFVNxWUq+ejp4keI4m53NV
nMfFGWGmaLhRx34FdeVavduWSCBVjj7T0Cbx6vqTHj6B94R7Bi6kq38Fj2Zhm/o3IZoc3QxxxB3u
LNNdBV6HTXHqlI7d7gX7Ewogz+jZxbYMB1dilpT5E2AiVi6NLTHojh1qNm2HoPza+Wc873E7mF0Z
TBYwesubk6hykQDgOEfFOho+rLgIWUTc96ps5APs52KZDhp9VWulbzpJN0KcxMKkMDCsBgPyVfF8
EsWtlSUt8kMlrxa5Au46Gurmj3M1av+P6qJdbJ/3goK+sSKb7Z79wfuQyTxileTrHbObED7ZC/oK
AfzfuDay0Hl2p1gi+tQ2FKHaZuq56cOjp14mQ4I0SRZlmbKLsoVBalOGCRV6043Dk0h6Jhn3K59T
0WaB2qfO5uRPMy221qAEU4qLSCnn0UmFo8eA5MBs7H8Ht5UqPG/aKiCQC9kX4tH4e0W7K5yaslXG
DGTHnZM0FVCGMUGe1j1IkH1ZFM+FHLL5lVJ69ElJg+YYyuWeBs3/101V+UCp7CGWhZF4kE1E+Ico
nK2ZMMzNzKV2unobQVlq/Tpa6v2A4e1E4Uu39Eheha3tH9R+4eGykcm9AV5pyF1pTWGCd1iEvyq4
fSLaXFh8/DEU40RLxMZD+c2gbmQXxfZTzk6bvj4E1J/77dnIv70kbCWwfTiRCAK8yumGR/Pgy3oy
T/P4bnxqs6XuWbHmAx75nLhzDgsr2QMIQQ026ELw7db30KSituzKzVd2MBYH88IJd6PZ/kPU7ZLC
j7xOzo11VOMQmmV/Lj++q6xNIhjyo4u5rKRXrPrGSX91yB76GAlCsb/iv3FsMYoQrtxwxplvllq9
jql1FpZD4p4BtuJ5LptQMdu44ZwxgPYT2Y/HOD9UsijofdZigZ8edQwZNm8/y4I/YbUOgD1dQfbS
k3adCh/cryNckYmqkr2vJWmSyhuJCiR+VJPxfOIOJnNlJtiJOGpgvkLpR+bMm06YeMs8O0D2wTwK
5ewd9R7QkfmNHXirf0oPWxS2woUf49JRBDHgUgaAiV8WNRBEygZJk3eHY27meAbMd1WO6Bv4/uQ4
tBJ+gI87GbGHzvzC9WF2w0qcaYRH4eTvw2lSqEX8As1OWcXqiMDK1YbpT5eZBIbxmCR7x/HG7Ok2
2cspUCg+Ck89VkaD359g6SLVptfv12Oc5coNtNXr/d6jCQMnsSCC6+KpOsfcFvcrJLnCMy2tr8Pf
xXmlHgLgvC+IZhnU0ywH8HlC3L2q8yYkEyqIPiXXlF6bPlhVkaucj22Qku4n8MuXuCk3F4diarKN
VWV6Z1P6cSKS5OB61UfjFlK6lLghOqOctRnAn+gZT4Xh1WK8NSLOsDnkYTOVYNl780zS2K1N3NmN
L/7S+I0Q5N2ANZeRw700V0zPwt4sDxDevSadpo4+Dft0rzd1a7libJ544FIG0YBxk+M+Ui9c/zYP
miJaFuHJ3nEVCJPYGry93urRIac3SpUcxXwBayO32C/teECDCoPu8cjOQVlovsP+mlZIf0GiZf8d
Fb/fFSGdY2eA2Hee4k6WQ1oGMD4iTmDGwH4i8s+3mLxdfkmABLEbksfbXzbITMb7mFeLQMWu/XN8
suFIJlHireykEHmhHm8frFtWy01/shnlAiwBsEXql88xupUWrUY3P5fRWfQmHAbumbBp25yLLGcb
qLkTr0RVtouxfzEXg6mCjkYNfVMfULyyfh3mVzbUiCEygkf4GAUNT0yt1jAGlfThVz9haGUeDy2s
eI2aJTEEs6c2eiO45K1zx1CDpmg8f+QqcEq6N9ySLF3unHiQBk233JohqvJVQH7+ngabSZTOUki4
jXLsbvCeWyYidr0MXFSmDrCRO9HW/e7jQBqFPlawBsEuNutsOby7bB5V/tdsr2unojy/w2J+RN4i
B+DAA917tXxvIQwje2yoCDFKE7ygZ7NcoyQ8LUlxyNxTwrPgf6M/7qgWyVXcPk6BqPI/SCkVbdLX
k1dxeK2fb3dP4l/uKzpENy6DaajT9cg9YEhydWwKoEydfTuHChihgVj/F4MzayaR09k+fpT+9bFH
vrG/jEgUSd4/mP5wC0A+1jzVG3FgRgN3BJvexa56TrdVv0ZWxbg8jnvtRTry+q+KvshNCUaCmJ5L
dNQ5RJLZHmM2hBGpnmuCcJda2EDXWredfQpVXk3hBY9Pv5ZgEEe5+wg8NE+jERi/3skd3bHat5K+
Eh+LVYDD1nUwvrUl5wqMvg70Sp4KN88QgEIdbRJNsVwtKF/O3raTsAVk+MwxGeayzHyZTS1/DhMx
2pBpOmQOspAhhZqjb9rN+ypjkPoLvaej9ZufCVHppykCDDmRFqHDdq6RhnGQzv1IS1DyEGDZG/Ns
5N1hFCxzdVA+MJA/YPXSnLC6SqVn9SMuAtG8ICfDNSwBFPzqzyfqbyV4E+sTLZbuMKvGxSpQyrEC
q3qx994OAa4hWqdCLx+u9TabOSLZw30GQZldf8xuSqvYw7ZjI//OpLJmZFDhiwnApEZMwMdEHT24
X2d0cvYPpHB0vyvHoirwqDwJZEV1qHNXp4K0XTCu7EtAo/NZzJRkqZcw2xR79ULTLgMGKk3N8xqy
wLekOKl7s2ZyW8Fe7oGk5Dw6WX1xbRimOz7SpwSKS/ckTYw3pqv7OHJvtjWOIoPYYamEG/Ycd7sT
CbClpT/zILSycVeQ8T7pVddpXQ/T7h9vU+32P+FIgxTAZEzypwF8i/FyluC9sONP1f9om9k3e5jC
0nN9UJqIV6THUo672ee7TSmsU7jxylxN4eG3nnnYEcBd7XY8FKzn7sF2Csb4qyB+ZYYlXAHbcItP
EDa3/IKH3n/jrwtwgNGdSmGCRB5seX2G5FBTrJhjM3O6KaBa0DH7p8qWSx+HIR0yQ/CAxhw0H9e1
a42ye3MPDFKHuZMt8DIYSODOTVa/ZiNGKBeBxsisQx7iSd6q7HASDXP8pESrJ9GGnvcmezHUUabz
HtY2fdOfb2wLaVRPZ7fc7LJW0IyALtZNUcTkOl2HVZZNs0b1zoV/Uf/XYjbLywFe5+Upzh5yQDwY
5471pVVnaECWE469EW5QtzdjWqQdEef7lk923G8koBzwGcsYo1PUSMKYHEGd5xCH++zbRz/9yh+l
d68gf4E+S+S39x821MrQAt0mgHEH5ievY6y6ROUftvrrkYKbqbHEgSrOCy9/anNIKN98oRXsIAJE
j0kygrpnYlzdAA0w5peMHpgnarNTCkV+AVl0ePVmBJOszJfGQjh+lteUgf3rNqSd1JU7hNZKMM+7
/TPCbU1skf7GZ1lrRIhG2cBZRguy/f/JjUidTmRjtsZX7QI+kwjKkmzBuSzYYeLZUir11/qP7Yzt
hupelLHcJtkH36MVkIACNzEinLSWl3WLrPZNSL9dmvc2hdDP7f2VJxZm2ZEeyO9v+4VoDnyFbiWS
vSOJKaUb90TSkAZ6f1nMhHFNRp+DpjYd2ioNmr3VaJRS5JTzyLqWcNtzD5+JuOtTeSnwMBt5StvS
f8hruXK0B5pNNnIC9kDrrQupsrX8llXaWAF4Esey6PHgyEeX1CDddvOIpQhRO6ahSjb7u4fpcyov
qxJnKWFHkCpMbkHewUyfp3P0qh5kRrKTrWwbEUo6L5XIxjroiOqo9H4VKeRz0Po4guPbhcmljX89
XA5PyLl6/s6D5J96NhglOjxD24v3v2PKowSKbvRjLS4HIENPXHSO87WpIQ37H2y2Akzh1CEicDJn
b/Kl3VBBORQTgqhbLjnocKLPf7S+eoDsPBhnrr+O4g146UvWzyNxXkJgYOIgUUlJ2CJJd+NhEOyU
b4QWfXgGcsHLAxwY9b+/xMxb78HQ/c9yd1Xrw2Z5eY6EwYC4x0dIbA2/2ei/q0v401V7352uy2gl
wDaAba588YJOMtERqsen71V4n/AxauxoAGetw57XvNIMAocSfLYrdclnm0Qi8Qo0B94EKL5oCZXz
E8mqehRZ+rpzKHCyN8tr0sgU9OBRFqZUAy3K47sSzO/Z/75zMWBYmWNGjLKUxN4zoJpIuLu25v9a
Bl2mAZuygmmtOf4HpFIT53TM1Uc4Zjhf4cMc9IEzEn9i6z/oQG9OvVbHrIHTNZo0F3jCiWZEr/74
8XI/CD0xphRP8Czt4U+4RZJLTHldo3agOi+VvxSDI7QA+0d/R86bIc8eaRYxOgxzqyl2npIqkGc7
M8hjgSfid91YI+9LuT7pokUZ4FQWsB0Vltp0geqrSQkUXn+U6+gehCyavB4LhTTpUjS1PZH2wGyR
uw1Ejnqsw1sokSw5cqqz28FFdP+VxlwvKGXm07qeMcoWqojcl3UoufSMWaKQxgKaVhQmiI+YJf27
1kUZpvNOjay73pGM14A2626gP6JhuNQZ5CRIUZG7PQie9+ONseoNVnUJQKWxpxyppZnVB4yj6E+R
3B04aUeGZUm3GcLkT9Yu2tXh2EabTCmEBDbnJHmiBVIGjhhTAUDOZ8E/9TlTbiVOYsXTONhAS671
fie6OW41CyzC28pmU5Roz9DFGreDtDE9DbQ3jfsoSzVSvqweWA3yAYUGzTjAcHYfvHri03jou+XD
dI0BKloHp0dj5OgObQpX65Ksrej4X9fZH66T5/yk8c3ZQRHS/m/Xa0IPuIMhzUkw8pKBRl/8UWgZ
TE8o67ZNEIGFWUvaV7iIM60Cg5z2+u8RRJ87tYIyDjGAtCMkp1zUGYEQgIpQxe4pqZnR7EJqFT3W
aUyNLsZI4K3/PsQNMdaYppcU54pzLtCckAYid+36IZkORi6oFvk/vK0J8zRLtk47uym6gmYeueaX
KdYQkxH0fgUjs3661TuYU3JuyHG6DJ6e1dkYP5fOSxnItiEhNE8uNqksn5hUz9PI7bxAY5bSA/U8
dpeu5fgqS6WN99XBtYd6Kg5aewbjUQavLupZQsZGm7Dory8tadOw1eTssZw0co3P5kEd421FoI4k
ERK4QPz7dH2CppWa4MMgMoux/PleXpxeU4KpTAtcTCF+nyjAHQbOoNxOtXchqsmBdDm+03zYEgWT
uWJDxBcD8lmSoumQGJjM1D648KGnOLapd9AKLLHm9KlFTwRXeMNJ1sLQi+ixiNMwvgvdYTTqfmT4
x/sdoFpY2kZJ0HR9FM7XTI5cn5WX1UAuDxIb/FAv5tz+je5YnlTu2iQ4CVyi5x3FMs5ezjjYAPNl
20iDO9zJBHcRnam5jHwgD/FDRCzlqWELykGWsFmez9VXBSm0vAGP+X283mzbmaZv0KIJuUltxYLW
Ceqq7plF8ugi5ihSCrMPu5+/C+pcvUDk0pRf5iTNkb0Q370jrqHsSrbB+YTdzBd6j33YYwFmKO8Q
22hJgnqaPG+gfqOCMR+lRatUUARm4h95JBigxEbVE2PyEB0wcag+jCWyLdONbFdk1okvTvE2Z0fN
CNMe8CUVUdfxq3+4CvvZAa0Dm8TYdkMAqtdls47MsJtgW52lqxjc+7Oof/cntewbct1aG1CgGuDt
cS/bHxvzQTMRh/ojB5gXPOVkH9VIfuiKahSRZxyGDDyhZdxl90N2FFm0aQfTW+tTBaNi9lQ9ZXja
NzR7UzII/AGi+yy8xSKvF3Rg0pOd9utRrnMCDmwYeMXBwZF4K2XqIhG2Oq5pXe/sBKQNTLC3GLXg
p2u1NFWUfnDHNnyTmcdEmbq1S5lzWS3OCxS7hz1z1z43HznsstWGFUAtDRKSPwjTtIExPZAE7+2F
+MxGR8pcMOiKD+Zmsgp9zUCIUvSZYiQ0c628hoEbAhmpg9vKCsUEsPGv8n8DM0/bQtDMqyHLj0TJ
l8Lnud9CMjKiM5CrQnw1xg4xKuN89mqcKKCtQdXg04h0HpYac8e9X7Eln7Z2slnoHyvbTsu69mI+
eLOcOlfclCkzPsW0insotE+kYsO+ooLVpDod4hmk+8e5SNqEFakU+BYTKCmN57d3/6TgxBxjcYzT
4Te35qw/t+zaAxQGNdBU+AN/FevGMQ8fp3W5+wQxsI7cdQTgXE8NeDEhLQNQ+F58HwuvzxAwy03E
PADdZnoaYXMb3zdYjpbskRBh3HZf2ex1VKDoUsyMz0k++83KRN5u3MNtaUg2GT46w8QDtG4E20Gp
OEvvWAeKm9SWbYYXrH1bsWVi+X+fVlw+eDMBgIaeV4LjWk26pxplfs4BbpD29lk5gu3MvOF1bA8j
2HyZyi+LhRAKM3EH9KkfbcnIc6L6fbzHV0W2nZQZ/Seo9oCJ48aKZsROFCJWBGJo0znqRNSqEIJh
Chz/GLJJNZUDlmj8dJRaxT5SNF/xUj5RzBlEJsxMvZFQWsi2O1gzGs5YhHjotjXa3SsUCHTaRDTe
VGz77bxLktvkl3v6ESkAvaJeRAb63P/lQK7BJrKaNJExY45TZZNbaCiVUoJz85626uhHim9KtlJq
fsehr/REZhz+H7TVZSeij5sg4XOXl6XMVcKbTHtS+gzMAriIu2FlmzPKuLRb8QT8XKgKpFaFvTos
kBK9bE5E4ccvVA9ynfSP3+5FrxFJnN02/2saTQrzfsIAzPCs4mb9TW5RIL2gTGGV6SroURCZrbvH
BF2PyFUj828wTCF25vnSoDbFfuQVfdgAaKxvRRZNXb+Ivt3vdsuKy81IubKXr811knm6U7X23L8d
STuHxrJCCpiR1ORlk2IQAwpi9WnghUvxCtuP5utuxxOUH4U9KbwBqX3p1va/hCNbhmGKdo4ZYy0Y
xbAnSj60Ku3/269qdZwO2iG3927gfVn7JFyuxO9hYD1oUGJeOIqPPmBkWNlYFblhRO440UaFttlg
I3NIwSTLpSXAaURG9cwAiaPjYc9Sp6TijdAkJSTVapEpsw1RPiYRVVEJAqh4l1IliLeRZUNN43VS
kpVgpdLfeYo6Xctg2nGGY4V6CyIOB6J7yfnt0c8BGkEyaXZTDMd9KHsVuYHGpbdRWcca73WhpjFX
iRjrxEqNuVpPK+2pVe1kyzAIhzfCvYJnrmibQs/tp6Vo77nL4Vhw6jQpFvI2zwUXWo+A7aILL12e
4mEuWkPPTjDLjCy1mW+cpaa5+WSIqbkXC3V/eI8VP9t8URVZkZAloyVMxZkC4V/LWDXRcbfgamPV
3nmZDbHNZ92vzpmwxJ8QRspZBizB1xq6NDLZKzPp64fX97HOmaAA1MV+dJi8qyI66q77Y5bhSkIJ
XKHDQJ5vAGc+lHNyJ8saKP6Closl4q9zUT1NLwwKAJCSSfrGHOTi93JMGxE7Bs1XSU8SQYCOyBXP
w8QqpENnN0jSnLZcc+7kb/FkJOwM3rsjUkBlc86Ez10WqxBlUTRsDFB0w1delRDI47MfTnOHH/Cg
TJMrFVvcmk7KkbctrmDabMXm/PE5pF+ZfIsMtAgOi+OFGzvSA/ZbZ7PEgACSJ3DXEQRoHY4yJ4bT
qHQ3ZR0dZ7u92UUpMpTsrI1I1TZYM/FjA2OK6Bt68XtRTtL+uLixrsJmeNBxbKzwTgbcOrxFsvj6
keuWVULJh4szQjqcu+jUIopjyvK9WM90/gBj4qCMKyK9FoMwMJN/u+va/Z4TgbrRpir88kauN8CL
jp3fahdvXdFsVudPv+24qAjO6rIE9+PXZu4SGDZDkN/wHKFYpBGeBbILNEbJaUWQRvDSV0x3pYQ7
nO/SqBHgNYR+RkWwG+RpSnZvoI0WJxI6pd4RxfKeuXqyqU5aZxNRVmLbFe/FqgdF+zvKSUwICD+4
HQ9yILxcRm4ljNGCk/jLnZDD5Kc62NtW+ziDMlriOOwGT5zEGetUtvIPwo0sn1fW1AA7IygiFxqP
cQ3MiOx5QVYgRY8/as95piHr6h35r9I2o6eR5BBYR2x/lYYpYu0DzmG2YvH1JkDTTucpnd+gRuJ3
0QTUHrnT1SFoJTK1taN3aDovKszVghBbSitJvTj2lxIHJTKchYO9GD4rOwhxg/vX0CO/7DU39Zl2
10wVKxZqUGzJtTxHXep8FzgqER6BqdyfE+B+ghstfuAIjzzNcDBB1LgkrNhwHqXl6iDMtC5aoSxi
OWA0qeWw/+AuQdhWqnwPPB5AqdJSzF8S+7exRohmToPaWbRyLDuwIheYyiXUjQ3jFzNo7wwaMzAM
5C73JvihC3mwibi8g/NI6SKJIeLmilcxSOK2YrBToazEbODzGqtCh35+UCTGEypsSOHAtQGqQnU2
IzRs+IEIQws7zoVYjSzcwqCtnAvuQ4F63NQRXU4HQk6RL0DnRfIMYkG/Zi4mdlV0EJM4hIBOSjK/
GbkvcrYW1nlgetgGziEx05+D00yI9e7m3il4IykpM3qrwAwmcMXXHI63yXbD5SeJqaiWWp81rjBM
ACRU/kFbfzTzeqGrSW0AqHyTRjvx8/fpVJVF1LHQb1EKleulQi7oVRSOgrewIGXOn8AvAACncAcL
VAqrJHPxVYRGmjxnboKLJLzhukTK25ixRK/HP+hG3KRY1+d5JCZJ7TlAhbnr8x3IjkVzSDGSNAhL
olqdSVTDtOrTzN8AfqC2k1NgYvkOYgT7QTiCddN8wwY1WKmNLITOBovHra/oYvhQqZk/MxeGiA4o
e/rwhyoHOxV4QCIn1F7FgFkgVqnQqjS76T63MlqwUNcuqT87NU4kv9iKMnYXoJeGlYmv7Ix8I2wJ
MNBQe+OliMQUDJ+Be741vaWEMv7yKtx42aGJLIQSa+2ndjRu83MVZHAZrNOqBjPBjw3wVneKuTDC
M35qM8lxLdjo9qsQqIfUjramMDxQWEAw8BLq+SBh1SnuMS0Mhh/dR0Htw4hLiNCCi1WrqC7KTFcA
y5s+kGweuz3YWXXoIiZTDRnXRgKPner1Hn2hLG7DknmACW+17Q6v59UtAzjQc7qgcM7Up0lvaAWU
x84pct5UYxCk9H0ftQBjYxxsaWhJvx2FStFKOOnrK6Hj3tNDQU8Fwwc4cRoKbYH10+7dMrkRdPY2
+j4gfYGJr6M7nQRXxzCd4pzuyp98YZUu+Hj86zpYavvAvx2zTmVzNt4D3gj5qT77WDOFitN+k4od
Hym7ftDaZBwrHu9tXYJ6WYXQmcmP8XLzl1YgPWCjGwQA1IAP6l9nUxwzLNxcjw+W+Lx7v4vXrKMP
YhzflHnek/ofe++d1hM2UIDWsG7qfta1vqrc0MDzLIUetgvMkFWKevEdMwLBX9s6Hxz0OM1hEt6l
rXt3K49FIF+n2+xW6cITm38Hxo9m8UifMWikia8VRlBhD0Ee89UMsAvpecx9b64g5mx7dqq4rfcF
2cquhBoxC426Uq1MnyjBun0F0eFrkXlx+i/PSovz6Cns3KIy0WtnEW4H5qZBVSpSqO16QExedRVW
Hafm2OWzU3F0lAk9L1rPgO8r+eMOkmP4A4hBcxYrYqZafus7NadVsBVDHsgvbTXrCnr9E2oSi2Qd
TIt+l82/a3NOyF7ppJvdNeFJ3ja6/gD85/GE+XYWHpUQaAei1UpnRyc8rUEX/gm8XrEGbBTtXDH4
0GjKXGsSphRJpICekKZcVh5cQkaDn+n7feIq0qF2qhIWzo1/XxPPLxC1p9r1AxriVznoxhKu3QTq
mm6np5iBTMKDggfsehOyqf9tN/6JOVbMdCHUb6pv1OgIoJUhU/0Xn8TPgR9/N3q2P+a7W8ZjpBk/
2ieQ1BJvaA1EGGu3KahJdCd9D2WJJZ0gFtWhMYwAnzWw6tthtCudvKHEu9ZCJsioDG5hR7xwqYCn
BlI7YhT5gA0AF7LjEajueDrrXQfr8z0JGkGzT4bdciwLoGAaMYmV8RT0gd7Jcx2HbFPi7Jv/aGn4
qS2GWPnTcVyLfg7qrtMhCu7150fkNvlwaurF9VhBOpsnMrLSwR2jbiPrfLqnMZaK8MCeP1zPIKHJ
9yAuSyYX9iV8Df28nKCrF/HyZm3oulM02WnRPDeEKk/Hd8MAVVd8j1WhwEzfuFB91Kdw9AuKlrub
7b6EFLcisdOY4xKGvIgDXxsw/OoV3V2a0kdX2MsW9rmR9lRQP1iDXM2zYY7TySg7mZQinMyksRG8
F+fSBaX/bbFd30B6o/vFo9+mMc718fES7BOpIQwj0mdp/h/MddYJ0JM+lj2VpgaOL3xe+sI0P8Is
CjYS0Ssm/RfT0ENUYdlR+CuMwZdwrOX5MSDfUUaURRcC2WZN/ddxY/OnMrT9h0WXCf6ZAvDS+p8r
lJmupgWnvIz/issVngResbt9ecEKqQHii8LZlvl3Z0AicJm3P9YIGhnjpZpXxaWs6ArARGJftHDF
27T9SHsudokd/nsZ0olC86ocSiwqtcirDlWUiLRU3uY4Kow6czOTafVuBebl7vUt8rwDVa7Slq2b
kibMAvDYYM7dQOSGXV8i1tzSAsIcaKZQXar36s0Au9Im1jtJIKIF1ordFrBPoXkUw9zDXcZiucu8
ndPenX0zzqORGGKMSWZCkfAJDvoOLhSzZ+p3KSMCZ90DO8BiruWy0VEwnNyPsE+nmBdwgGee3z2s
8vSVHJA7P7DCH5afkMxvDG3Ovg/2qYdw5M1u9hfIXkZMBaUthqbl5bP5ZziQCyxwjNSPiDvOWyy2
gItdYWuyYYnqICSoNrl1s74hXukQun/tkvwg6+CxH1yFKsUlckxdFGgkxGW7LLtyeANTWEEKlXSM
WOOKZF0hw5bF64M5eaW+fPR1YRxYTdTQ1kyUU5q0zoBwI9Pk6cjbWWZqYCGRet3FzfA56avSkTWa
VN0roXeQynlRMOkNsO256ife5mRIgwxK1VJjdfFNUurKJNCm+5Ltue2fCBktB4/IM0OMsittA3E+
a0ohUlKPH5byHJ7w6NVjtL8aT1I20/FKYoiYd2oeVXg1wh+Mq06WjdiTE8JrmPqec2UMaAJ1sRKE
agcOfsrv8A6qpOQn8+ZXQkVlucK/Amp3aNAJvrru1pK5Ligcbc5ZNxhMZzjHtnfQumXd65YjsrHr
cWcMqVloEUnTs0mdsqfzBVNhn8Zt9y/2MzrwRkZkaAm8CIM0H+5B17XLMRk1LEeZ0XTR6wYacVac
ESS5vChZ7W/BztqAVFIyp1Tg19gsTfyz4pJzRMv0gMxd2ZFu7pjoxmiDu3Jbf0629PYGIWlWCKr5
PwzyuhEq4xoIBDZDSV1Bh7wpTJ7aBK3gyEbqwcksVnc6qz3VadBieKNqYFp1wV3Cx31mqgFeBP/b
qISyyxOARwIHWxKuplhhSlg27R99llqJirChva4YqUNpHfCVYwYAiNTGsKsmHSIGWuzGQwPO8otz
lGOxsjElkgBs4JWs9J4n3Iqx0oQNQWRliKxvOGdXVY5jQN16HjfGN/0QVZRVXHYGqJaVWEvbBqjd
W3ZHak7QjuLHoVE/c7zfbhiL5407wb0KpAwSiL9tX34WMPuVe09tekWUgDmxqvnWL2INt+YO3nIE
iZz5lnvj0SjDVpJTKsA78TVyT0TEJyH8FbUNJJm2DDirIAOfFRQcOdsaOODvGwWXMb9esuO616PG
sqh0xrsbfgz5maqfMcbKllP8Z42ZP4vqLgckw6JBwF7oLlU5ZS+V13Ven6vsIJ7XTKkbLXB5uxSB
ZwXIcR8eWPLUK/oomYBNir9pLJQcKUh2pEZnb0BRKD4YR52rt+rBYtCrpyn5Mzg7ulWtATHn+Pg7
1a34BdHwN22f8pwqeONvc0Hw7cC0J0TKuDmIuymH+ISCuhaKKWCDzysE/UsDL5vF/t92hPsfnawf
BPpTldsJ8PuD8lvqLakPI0hpJsaxZrrTGDRztUauw3BZMTQQh/epVZCCqRpqtXpITJd6G5hw320d
VAqXoUpPfTx962getFMleDA0Y80CJK1g2fpBHaiD8hPNvjxcGI5wwJ/YNdkNSSxCEMBIszipOzob
MRjOb6XOKDzOj4d22Umw+lqxEffqGftPq6tIc5Kqz1L5lQTcYGWWF/162fTQ3f3GacpcSoacyCFv
KauEgtfpSjG8uLGkLOv400iTXBL8nstLzll3jYnMtYBW1Xanh8dahAcFHfIz5qBZ+EgUahmhrmcV
8XzZIQCHbRWiI5ecB6HNO6NtEMxBnLWtJJHH5jDtcqFUdQz0nOa2niSev07dMsHxfmQ1wKLFT8er
fJYNgs9mqdKExJwBJRh3+4lNiZ7gn8j/RGuAR8V5v5cZH3PPzIpniG9MXalPi13DmSGk82dNKdXF
DKbizuX6m0YvidwbgRIs2j1lO5zRS2kRNN/AUcdu3a/u9VCOBs3D0Lu/LWodaPMAxRtw5mZzdQM3
4QAMhmU9zHZ8j5miYStj+Up9c7RhZeMehdXoRMklL80I9iRXsG5rNC8WMFBdEU0b0P/Hvw2COJiH
eSVKQtVRFOoFEpjwF1PI7Ptis27q//8Axk26zvuHn6rJUzIXm4rcMn/FT9ErmSBYyQWI5vLG4xXy
p1g/STSek0SfEzqwMo2Vgn8paz6v6UUSF6ZrE4orzl89UZeFMUGMJSIgfK0YG5PRyaLdDZk8meG+
5SZ6NB1sqy7PwAzNyJp8f1TVBZpxOow9ZGTjdoQtw18tx9fUKCw28RhLWW/UBOuSLcSo9DKrLtpV
SRFihKweWaK+LHFsgXEvxP3ZrMeOqegHbm/S4Rh4McGIt8zb03wnXxRFjbf2x02wTU/4+fkOQCY3
jvOIv5l7zirNntGjSiq7wUW7ciJ45z+Ot+ff88rGXfZNrsux6GjTkzqBHOy5WBy32Zpywc7D7W+4
5p/aKcQgFJ2hom8X51kWgOf+ptRdHtyLn/Aq1N+Z7pi30jfOr6y/RHSzKalE11q7HXF9nhu//bN4
YffieoAFfA68vSMNGCjV1uGhmmwN3pvCpEYKSTqKxztxArQeGHQ+mWK5VtD9EY+dgZr5z9tvEpWV
8lcxd8CRH6sNxdxv7UL6vnSNLB0uBNegSWBKbDpEGJklDSNZJw47K91ykL2SxECR1uAX4IfFwE43
ly8P6CpqHrkC3El7L4eAOnJ+/VesrLoPG4ETUlyW32l2WrxpOIY2fbs7BZ5k7ayEWwixcxE4xp57
maNE0A0CxD6wt+gPLhDKCQweuR9+CbB4zBnG2MyG9sO6TyAujwiEsbqM8I9msPofeslfbb3w8M2M
7sxfndK1f855BXgzyTBU/JsI7eBOkrZnypShlQhwm8UPAca4EuRNaL1VMs24nuab2sSyYiJjuE6H
X+61NzDiDP35JT0qY0Lxqjjs4R5KU3S848LOQ56d/9nCnB1MfRouuL7M7rQQvZp3d+SMsNRqe+03
yDFdAdL3aEWb9xFvZ36g30aMD/R6WVuWuG11LYxdXTigrbJXAddN9qSK19+mJGUvVetF8qTtQD63
I6eLoC/XNpXOJ7yYxRdOnkhS65I1mjkGSZFDeQ1fxXaxw/Lp3087HOtPwES76/1KyYnB6hjc/SxQ
b1zZxjhzi7Uq67tNpj8jTGXdhhos9oHQVf9GkS4GPRPfitkFXO56l6d+l+2aLgJrO2rVrTOuOBDN
5EGyYtV9CySCX8wIBST7D57Ryz+x+FYFeWpwWC+m9d2/7kZR5tp+kTNpVJauS4ZybL67G0FMDwnS
WInlJxqXJx+TLh3ifLFrps0CAbLxmxsuvlt8hl+co63Pv1ko1Wsitop6aDgHjA4DOH6uMZT9UttG
vmcOVHIO2Iz4ZZO4aiBgtLJTrfDRQv3kdoy0Rmy1GdcuIfrkqtxbbMEC6TTNJEibns3DP6FkFuhS
wIloBh6CHV1NFGGw9LcZoSycCOWoqzPMdTnLu+FVQgPRp6Orngd1rqdF/6JmNy0lDnuSwPoxulgI
7J76amKF0l+gUORWJbQ78IGrA5YBhjtKzvh1qgfQJ67dlaTZgYh8RgaBg5MkKTgF06xVXresrroo
kNe97NCMrHjM4tNf1ZNy5hKk0GUsdt9RXjG3XFKqhubGGJ0cupCqNLB1yzXNgx4xDxoPuaH3Wgl7
5JvVe+4/VuyvlniMby3TRvxBCN0HFN7gWj1IaLAxeyQvoxusoI4Gq7DNV2pBtAo3JhsC1UkD0CQB
G2RN5vEFDdWFagoJpFHPNlWKRO5dlrs3UdcK8TH6jB33NCQVgVHbBV7BQb9QEbKPuv6/OJGjsHrl
JV4h7LhRZSG3q17rMm76nXoay3n/FOy+r+egdQIlYyQZ/NKVDnLBj9Jf+ef1qI92pFHXSzreSewX
yYyM06lDsU/ot5D0dK3zTdZfiGjFYh4UNZpPt7wR8D/dXgBEfDyk5pJifKFywUhAWGMDeLTsRbaX
wss95pjLW6mWRn9Fvg8vw4FN67Rnt+DU0zQKtmIHz71iGRdgS7Af55TV2BrHcvZ84c1mh0IvovOY
Bjk91iGdDK5pWjqDegwN+HYYPrItnVnVPZZxI4BTsvCsp+cltjF4Q+mN/8Wqh4JQ084pMy57uxUx
SGjgj3I2J1iI0ARKmQhnMpuB+dErSYeLkmMqqFJKy79HFYxiB68PfObqx7BEsss5FYyyooWPBo4j
/aFMbQfu7z6WJdVXZ4L58ylOx3bbw3zwW6+t0Tmtw4MtKxK5SQxy4eIJ9NqJ5dGhkETm2EX3umAi
7Nv/LZS897x8fwBef9+p++fG3SmwpF5cPxhPlGAQYuC/A8+JXeQp+ciBi+uIY+YNv7wDfSjDXn4n
xCCLGNELyJFJGJT7TFOC0bZ8kHS4MRoAe0kgpSWTS1K9aVxLRu0sTGtX36ydK6dTxRO+QyryWc/3
4BCPj/bOmAvjoHojQiM/f0FWx+RY1w8w5OVpfklP01fuy+LzoXb/+3gcTTM+vyxSc9VibEAe8ITZ
xGVlcabCn1ciq3A2N16YjndSkqRxAptN03s9rvb25LE9vzg1TizvXyWb1jp+NR+a4TVrqMwkkCpD
nQBUHhHrERG+fCxUNv7AJ0vZIcg9Kd2MSqGJh+4qWIXTdlrJqzEc/mdcn+dgmL2/pPKI5XizpM7m
8hoyHX47uTasggHKRryfADg9eD/O7k3gNduf1xZRpihtvUNOzDej/wPmuN41BOCe/jkI1e+DBjVg
1xqyqQGtH4cxguBuvxaDACYuwNsE444nullifRBwp+JaFR+R0Cv2wjwvunFBJ7KaXhwChBxVbRvG
bAdu6S25p8y0qMaZdvDvO37Y+dkK+nzNjDO8FVpGBxxxn8roHrHWUIkndEiOWwzdURA9OpbZIvom
i6i+5fkslNIHMJUMciC8X1FGx225mWriwi0h15Cj1Wp/eG4XJjIcEFQUCFTwZ4b+RCkQto95Vmc/
lG8N1nGy5rVbqt2yVzkMDPALCeYqqIYRLKOvJPtxKK6z8WdmLYhaIRmpMTNDcNcuVkpZSk2oQVJw
p2hpn4UQx/ou2Nw1P3ln/P6TK98c1K/Mn61/cjJw137Py9r1HqAgscTqYD+cC2aTTxpwaXaVSc3F
9x4K1VFaKRjBXxeqAI5zsSxCGFaAEu9M1O2L/eWL7/fQSdVQcqfPg9vg22L5UucoTdcDJiuD0j66
ij+Dtd4UApAKlzgoYyHpx+eWepR0/lSrKYIffnRd2Zl0i4nAhRN8wU+KbHDIFpBbqFAMZrrVAAww
MbYwcov7/cPvYElsl/fYj44AEG3u+ck5H1wxDPSrak8P9CzGAxBGUi9/9wQF2h8sQqySLmaYTIby
7m09xZilKjJvswoVgsD/wABcpGI7tL9aGSNK/p5EM9kWXWXB5A//oka7JWx9r+44pPm/p0cBs04k
TjWLHHPAaAkL73Q7ToLZ+r5YZ2Yd+U58FfUoebz/Ih8vtYhWu6FXABjeGlnmJ3A6mfVMwSqeUc37
+9VEGEDbRicMg3AshV++J7wxUl5O3xVj0+IqXmWK9vtnKhXZn26aIxN5naSmUJVKeMTVZqoQmULy
70+Wfcg8iVP5xzUT/iDGvbkHwUUKpQitFLII714OrJTvkDTeIJe+ePTZ3jJW/dLY+GlmL3xBSFCL
OwoVwLWDK8wFpyzidXIeIKQLtJ7bKRzEJpCyxB+kQ2IyQtcwkkFE8YN3Y+qyMt9VsvI4d9Bxrrct
K2qkQRZAdVdvCVwAl2J2ZCHXscIjgt7jYOR5+E+OfIrWuFNIbsvTBjx6inml251kDVVuC27jQYG/
R9oWyxxZ5FqRsDMZjqupOVPksn6IYpWt5pFo4qyZHbjcQuYH/5wpKPODfbY4ClB9/iBcHRTjA+ss
o5e07RirTVeQOcDExx1M7defn4/eS1Yj/dyWwY0dD1TOu6tNfE0rqtPi0DbommGpSmiFdzHzIvhS
xdj29qoKMpfFa8MuKyS1I3+1AFSQ9vyIYwlvlIrUyZ1qRBccPYkB/hrH9iQgwWm5V8RFsyQTCJ5Z
A2v2BBUdMvgxGE4WLtjSAZYwGE9C5CGLZ6qHYOF1fg2XS2fYUSP8OcJV6EtBide36IbCk7WT2k0U
YON3Et9v3QY9cu2qVbdrkVTfJoqavKFplfuNmMZq2y3Qf1Xbu6KlPdytF9lsclCMbyRRlkmpPu2o
LxqfXd6D/8jGj5yVYeMncI35E8wI4bh34cghJNUFd91xGug86NbpCp/P2pOsjW9pgjwdmOBQBkki
CCGVJeHhfmB3+iJQs/ydxYcH2XRL7fdp8eMayFRw0u5NeASD9xv4YMKARXlOApiw2SGQ0L7YvfxQ
ek2MCJKkVbUV1rq1PlO/vzrTp/iu7Jzy7dOafKgGybjvgDfG/B2thM0ZF1nXVVWRENpewA1gRMrb
HLDT8o9+rsIoQ5ZjuOFxp1SRPVBBVAKJt+/kMEhBFw8xCSFsc3IqqeHpMBLRsLqUR0nIdJNCvcA+
wienv3D+Hv5fPV8Pt5Eyl8xQR3nwgFc9IEMuvPjFviLLifud00/LHizUDMJPmpqGk9LVhM7/ZKSt
w/rbO4LjecUwhPnm0pqWG0YXTn1PMOCtYC7dEEcM7WAgEvZKY6DJHNd85ic4/KJtuE1YS2l9JQG4
YS8X1ZJPCBC/nyq7X3HGGYvYVErk9bC6Mj1RbmLSH+pV1ZZqu72G7E+rKTYxokhp+ghv/CkWLm0H
wThbZZqAoNmWheWZFYHeLQGJDYh8SioUviYdxkMN0EtNsr+xci+tMT4IbeLlOhoA09+r+LvFk83h
Ss/I7eAdUaGwwJrberavSByVpC6YQwvkeWB3osSxTtA4o70duLn/LsLBBKBy7O8bSIgTprNBU8cu
iKCwWoU6EMEEbV2H8+LbcopIHkPBGZPfJrdzgrHmlcytue/9jhMWPa97OCC07Gijgmcd8xpdzfdW
LWtk6HzkHvCEQL9UFcn1ojxd0g8oEA3XM16PV1bguzoeWJdyk0ob8RrWPLvFTl/WyrL0Tq6QsbaO
Mq7bXTWD4OxqcvOlZ2253GDXwpyEQu1p13C0WWUqHRu+t7DWDeFvhCA5en9WgYv/a9VDL1Ov/cJh
WDJ7EUgogyi2KJmSoKiaoPtzEhpV8tv1REVBkaEXUaZNOoHRFF+WzvPKI52ok3/dbfZHx0Y5lNay
61BMmuLpMaEUaKaYSdsyj1f3Z1zHsgjOe6dNCoU57GUUdGXGUp8Izx4BIEIvWbEXk+KQ/4rOmL4F
ASgxmtDQ6dY6NLJDrh10tLHNpjcTq5viQmkpXuTVcxkoRp/Zexdt/t7F0hB1N3JZ88FDf0cf9cAB
58FJxpqxjFwkEsXw/nVVtVoQpVHtVYW4YI6Pc20FkDBszkrp1OLEssWpyXWlmKTklCPY+HsVbLc5
Cd7yLhbQGn38bbHtjuRWSkxXtZ5p/jG8I4kH4OSHPMh9DXF66jtcrZJdE/W4Oaf9a/EzDrsVcXlp
L1adfxWdAmvfiikSh8XwTm2Ly9AwvJ8/PAh8IfF+0Xpp+q/iSb+q+bm7TIO9YLLBrgVCD61dK9Qy
MVgdPFcAxEVbz9P8cDxPhjkNrmT91BT65JwIzIfN38QjYaHKDv1mRtcCop5JIZu2qwvADYFYY52N
aTP5+ah/s7QA6dxTluguPXALDFt7A5eajI7hMCkqZgIlnRD4iiufBzaRyhMV/B/5oG53ypP99VUW
DfaIDEJnvTQwlgURN873aQTQQlYjqEaEcm4G/Jq8pcmgkIfgM9Qn2fBqJXywLHZz1TbV96trLQ1w
nhHFdRT2fc5LpwbpukYJxKdViqX/GF3hT/MFSkD/iPYY9zDRswmzSV1XTY42fJjSHKclBuaLPefH
tCDajQeDVww0GqQMKLguOEJY/xxQCLaWd0we0PZeg4KLKUvpxzUZoB6aslhAs+OoO68emGZrwfjr
1+RWGgmFtj3xcg8oh/E1uNd9JusbV8ohNes+VnpbH15zW9VYcnWcEQfIHmgVClLcrMs1G152B5Fy
a5dH9I8MGpGeZureSE+mphKI/+BjQHTA+EtsvPeIpGAeb6EftZIVeCbcRop4sARxeL9AmD+p2k+w
P/9EzYGfGXZVeNVaF5CIxsFIXSFMyphab+rf3er8jUlwFh0K9MJZEgMjBq9Ql+ksS0iRH+GIv4Os
eR0v3qkCcWmTGqnLCrDRpvpTQtOqbHo17XcBnQFR/4J0QbyGjbrylPScDav8B3RUt6hhH34njkYK
V9GdRHD6PfUiumaBOSm9/KHN/PxCvGICP+EZg7gPOjoSn5ol+Qq5xD+kfu7fW8PFEic2uWAd6M9b
+Bq59WBKwouSWbPVWQ+etNMPlTJo2vOR1EZRxI2OGRiplpAvj8kmAcQPkT3oIUwEypgPPHPH49TZ
6aUbv4cK6L8Nwbx8gu+kT6LJ0VOG70ULotbnN+i+x2Y8e2g0Ln174bDH7NJ9iSs5x1SvEDSvwQMa
T+Nvh09pz0EczpCv6HMaNdyZjjWZAKw+YX7fBKgNW7xzz6oV52VqiFTLgXb4gDAIRLiWD5hhWlaw
9PRV0NDhz7zjf3AmK2kf+DSUC40mmaz5Ena5DHX64uoiGkJnOzmlDPUce4Hrg2xCNsbh7rdmW7Dm
EUetZuWKW9UFOYJ3J2B10CSKnzLYLa7IW8REVpjmllsPi+iNDugiFsODwL1VaIiklfkC9M8UEnyb
eVWp22SmmSasdMayHVHjtxLw7fvi+UR6EqDTnpDcIIRMMSTaQh36sdtJ8t++g4+Xjly2WfwwAOGU
Sv+kEKXBCUV7Zod2qus+Zp/Pjl1yaVRczsK79awjdUO+j5kxDQqGGxx9yXvrM15PJ/yW3WE+841a
ejSoXk39Ie51Fj81TrS4oMUdgsqkn1TaiesOLMErYwzI9TBsEkL1ggdFsA8UJ0xETbrNSHrNjL7v
o6jdWB1b3MXkV9H/nOVBa8Lag8VQQyIKs0IfJLwFvKWASh9yTACejpLRpJEKM8fADmZwWWcT2jGB
gIzroN6E8L2bKxkzYZd2E04e8kAc2KgheWsbtsOl+Ylz9uRkPuNA4L/a0Q1wlohQo3MWF30Pg93S
MhbtjZmk1X+gnnyDatuG62mBrEyN7t4ht/FjEAzNae6PsV0UTPR35h4I1cFLl8X6RWBSZbkCYtDn
gzbCaYouWaVyq35J0uUDfP7UaZkAXxTKdACv0cqln2zAkMdfDLnLjKCLsS3tFGwC88PLfZ/Lj7cA
CT2XOn+8lWx0UseFMZDVABzY6FeO1y1IxRKH97hcVmNfvQdRn8xY5xP40L2zzQE4d2hKx1yxTXyQ
oLlvrukig2+ifI72xrTXUXU36csplSsiv9+MbBv7rc9FBFeyS1UroA8rFaBRHmMLvu5/Akk2bdkK
vwCvsbScOOSVliHwygqpWIiJljFFUx2SXKDOb+PCwv70QVMH58RID8r9NDzgxbATD86uWFOXM5VH
TXO5pTwBjHhFjikgj8mHE99Ac4+Gtlh0TT1QkXhwD3U/Io+NRfrO7zFKKQMta+zJhXhrRbpfIuAE
F8JwYf9/6OaNvnR+M3d99AU1aL3nSPsmCbwr67Vvrd1O7+yJyxbNmuAxKg7Bm/Sct+JdLyIQt1+H
YxZGHvqVE5gOdoJbz5AjtYzVQBCJGGr+msDGUTpff01rpfjsYfuNDLp5WL47d/EkuV+TuXfEIfll
b2OtyWoxbAngXq6VnQ+K9MyrFVWe3R68t5FHB5c4k1YCJU8zMd0SgivVppjFSlluLpgykjpRO3SP
YUfmGm4ZtFCEjV7mX4mE7bD6KZQ+2wOBzJo+4wi/kXkDfNyyL4o5qZx2Pow/0oFS/7XxaeCzf3mG
T/FKlNBXkYjeoAQqfWzBxEHVlxdSfc+5ilZCCe4exN43f2Is9HE8trN8aQWC5xLVM7F5Gx68fSwG
4cYuAqmmtTVRLcjGDcYA7gDgA3qH2XQhG7TkwHUEvKGwSumfhLLllaTby1oO4XoxCK3Bdzo9VCXP
5JrcVyuH6xuCrha3NJdY9iufstld8AgkSDp03DgVk88d1opkEp6vDKXHCAkKVlZFlwd0YroEggyW
LRije2xq0tY8SczvjT21aPQCwJw0hOqICG4gMoBbcBG/kRIjlxIhzu5I7YoWItjghHGgLgr8nf77
klyCgZb2h9/7DF3FhtYVecSCgJQXTUdj14emVsYtD0YBI7iqMvEmTCrjWJLwzW2xPhs9GpmhfxkY
cZZVpNUXLl4ptKgSutgoJNxhK9nCgFDEtOh0mEEdRc3vf3PFhhZYU5AOAXpZU2eydND+6zaytPbR
/Cs4BZ4oBqMx7TCSEc/kMkIxmYKRm+rvUUS6FvbZLS37zdxfOz/refNe75zFs9uoAeCU6EG+6Pmk
J0rA29gF8TOChRR3YNrAG5fLSe6ohjqvQ9Q/RZatUnp7OXnJ7MtLzkFkpsYRgpVNnEk3ee3hzrn4
ifVkql1i0AVJYAwexAfyVGHC0YJ3/waWT99TFkxABM966rSU/x8eeILgsqfAVnGKKfQYXbe/vNC7
vnlnsS8lSuACM4X3uEx/Erk1q988rE3KgI6qCvOgbHSfjuZVFJHVyN/NBDCKHvfQyCVA80q1p24D
DIR0Jda74Z23tsnLA4Fsqwq+01CAr7B9rf4fq+cAF3caRiS0EqiGCEtGp8N9rbQudUEA8vXJd9j4
0QKWy9kz57FybJQVzLETTsmcvUA2MiRQftZdCJdYWiix2OlvLyq1MF6WaVuqP4U/m0D+J895Ry5f
u967KjtOieIkulbc1m6cOK73HdYQopTW5nU3UqXanDaBaIvOQoRi8HETIfVN8ajK6XghdHqlVr/y
Lb+v9f1uXxAldkkwZ0mm+n3btxnzcZH1G1F2MSRLuEIEL8WjB4sBISUgkB+nvV7loXEGaVyX4YV5
6nyQKUaHjQuw9mLPe+DSLUE4N9YYVD98uHTW5E5xOtshPzXrnjAJDos+bSsrPQlgJcQ/aaEnUP3Y
e7nqCMkB3I7LDymxkMU+NKwUzvqP6yzJB0WGNpi59NU1fDcXwipN2NuZ30zJSgm2SXyrtD3wY1HT
0BXs+5kbz2R43By7vcm2vgCc7Z7/2mHjxZA/T16LcXRtBXfT/ps7yxT5gFgsAvYTR1odGsHo+M0W
zwoa7YcDvctzUV4pCHlUnzfMUlHCwJ7qehWRNQOhplbwZiwWbI5H0wCht3VgZHkHSm/z9CbEBj7B
R8e+ioDhAtNkBoo8NEM7x2LDjAzjfbE+fEM7w4L7U3NR4Xx4UBkxXvnsPUSa5mPG42rz4G5XlIzX
fAnGZeJEakVeCDpQDi6U67tQmhBkN6SYNyUdBt1iZ2dzrx9ay+OqB7qThqGzPRbfvYt7xkIAwC98
DnZ0gylDMnR28NtOYhVGr0dZyY7Wd+xjQtoGDhzwaAvjgun1oqrXhI5n9fy5zxKyXIXpcVcMnmvS
KRek1sEPyaghTWHLn3OuS7juSwlcMntuwHjwBFu/7lgLpbxfoA2Ipgn8ZiB03OE7+uP30doiVuRW
RJqIv+bjhMi/Igr2J8CZHmPHx0iLBmE+FvHgwX7y+gzLFRNMFT5iTlLXvrIqE1yKTI0V8lLQpNlu
nSguAiXuG2hsjqomQhokqeerbta+xuz5sJVQhdX7YF6G/74IyMU3/18EsZsoIDZYiBE0+w/oXMip
hAYuc+pW6j9MBMWwvWZ3ATLNAuAeeRAcx6mp1i1LGCC3JW8wmyGSRNN0P5n/Jy3rPz9LV5mBXyzE
x6fBpVgb7VFTLsttyS16XJ7ejiedxXBUxUdG9L9SARzfNEJ+tuNVW585ho3v5pynbbx8HEaJ/X6c
dXutXIdxCsen8nyexdrGUki9xuQsUbg9kEopusZqPT7weEc+g+nhTAia3jWsJ+PdA5Jxz1ZDnbPz
BlqNX1ppmnflY07CPFqo/rxgjuwj74R8AKGvmZ9oetUou9Th2/4U4Sy+eY2vm7mE1gpyLPPLIUVc
kZmRpnTGo+7F3vn7GdZKOwECpyJvWxpA1S+g7yxbo3loaYXeL5ieBRsuq0icpFDfAhvUalhEU0Dk
rXjq4g8k9dttJQotJZvQ33T3mIbG1FYO6+GfIEEF0s5/N42l4onpKWCx4oasMrJD1u8CoPyQqJuF
sIKxz3N4H39LaEFUpaC7ZD6p8cFQsFkojdZG/XIjXiJIUCQcDa3Mg5MEriZqUOYWkEEzK3oJQ+OI
9krs1X7l7PX2Ot/WbqBdi9d8yyIGCQpdxiE9VNxfoBbzbvkUDKGLlGkhG4Z08oXTGGl3kUNncckt
dkY1YIY1u2bNDULnoWWDWOIdZD+NliqMpjwBXfk9hNqafMMKyk6H79Hohx9WcYT5fOZRaU8Pbc64
BW7IUoZXcQrS3DERJZTxkkh1Mu4QZR5N44QtJMIUCs0r9jKQSxHo3PrsbKNaR366xBtZea3OmGm0
eKinvSfYN6tnlttVmHc3+KIURpnT/k2XpZNCqHfyPoqncA7oEaHMJas25sRlq1tlDtcttqA+1wIm
Vu0qdj/QLyQ+pCvhmXwvmQ9Y6Z1ADFhXrNbw7/1FYxxg10vXjEiW/Kdt1E5raFFysCGVwDs4T+m/
XRPQL6RuiQ4JWCqSNisxZmIPAE/dlBvOgmKlIW0bSo2huDJDRgEJ0PiRBvLLQmbj0AxN5bC2j0fE
mB+0VntGdmbPfX3d0OrWTmyQC1zywbCIyVv7/GAJzz9ElWAtBGbuPqDAqEvHVLNZNLMFhsRxXful
UnJcSaCb6Hp3DlHEcxFa3sfUOlI+1avAptJC/JhdMDSVTNXHvuGRhvKX5CIyOl81unlfe/hmqqgR
Q/lXyQlYBQ/wQhePLkKgh3f+RnvpFYC+e7JrsxH429zhlIXaHrPwfRPS5ARGUSJ2VuOpFoJ9+vYE
HcDNkhLSj8YluAFPSmqMbQjOgOucYTGVET8rqjM1nqhJ1HbnqQbZmr4tQpi/w8JE6Mhlo5bbsVhu
bGsd2XKbBr3uxE80A2MWQCJmYt0HJptE3tRCnVFdgvhvm6n4/3FjWaC0UfwLsc5qDAA5zbxOkgS1
Jrg6o8gCJV7Ku5n2NeAEC529PZurNQY6Q/NsHsVcR9MeuGuX+vAEfEAK0bW1Rtaxt+DqkQvoryiD
xf8sRU7vvJ2Ix9SmhvWub2Av2SCA5B2FbLN5OnPnxpCbBc56IvE5Es9d/WY2rG+UMEHAEPqM6wLz
8QGmS1Xj3GxS/Ckp2XyId4WjNQYHJcVmlJ/Kw9xJIV8PpfpKcvs1KQUhk+PBbF9tDB0irQapDJEX
AJDElKoClBCNxhJCFsRAOQaMZ7zz17pLg9Hcs8QnUu6Ic585dTO+awUyLmrv+l7O4/mB9Z6Qs0da
edTNKBGp9065duKb3XkwQI04+hCe93+k3qG2KFlc7EcSPpaQhtCWATFMDx8JCgzh5ZmFc8U9La+U
Gro6Bp7MDQFLK4WGKvxLAyZS9+9ZMaOf2iI8N1kKUkwdPvZl0IEjpkSokKbS2fDBCD2x7Ufng6LQ
sVYFtYRhtVi17jEQDEuoK0EmCfbOcwdnSUQAlR7qqlJReaHT2whryBDrW+H+fuN3/kvtCDxfjDiP
OrCA9/G1Rjk/ajrn/dmT45OjUM9dV61GFn7NmE+rAi7MNiAqQx5Byk+hYhoNwV6y/m9nNakcqP7q
lbEDzqNRNlgqYfhYr/FxnSkfD6M4WMVZS6g276zghpAm5ZNDrLn2g8wob3tOPgY1hJoLg07F39BE
SvXvVnCdXIe/BeD47mdVIo3qzm48V3Wgw3V6rKLC/7MleP7aFjNAdPWSwOzoc6mKjoucEECrZB//
M2XeVKdhMjzOKYqNA4y4muq+VxDjXaSnHSsUC1VJ+cHotaufPQrtiO6Tu50jAigm5GH+SNR1J5EX
Z5CKGPj69HfuK88SZsQiEfMqq/8j6T0qgAgppe69KReXGKV5ucnwCLWMrY11fE6TwDSYv4MIOQQz
HLPbNkhmkfzMaJIwfu91D/GDsa+cxXNm9O1bSILdHGnVW2DwFaMQbUbcQ8U4sHuaKbJ0x+4g7yyh
FAc0rY/sUNr15F8pEPMWna85UPSHqcWmFDW3oREQkr/EDr2EBx1Rhmi4d9KKW7rWHNRyoO6ZiZ0l
o7zgqkc3Zy/fili8IR0uTo7pZnJ08rnciymheL8nNvZHVCZEAYhdyGOBJm8tNuHwZq4c5IHdM/CZ
7Nis3vQFUQ53uWbwseknqKixRAWQL8zDsZF2mn6sdExyuvWMkrJ3cvY//dZZScAXDQMS5N1WHFs+
NsEOmCpKhFzODBiuZeAl2R72rb9ucrRpYo5X5AaaQ5kP2GBrMEDkFDAMlFou5N0FUJBfEvK/k0RB
CB3jZbcP9rdV+x8jBBoVm3MeMMawGwDZry/EkgHha0A5Ffv0R46ED+ym86N0SObM8l+e89fukHX9
ofJQlt+PWmI0kUVHCGzJlFDHDtHJCDEK6BZYVGVi1LwMnOA2WJWE83pcSxcoRceiQdMj9H2m7c0l
rSiQ8t8jblxUhTuEBJ6Um/lrrp+F5mWtpDtdeY5IY0syeK1IzMqA3i7LJvsncBXxB18K4bJvdI27
/o87o+fGBLU8MMCvWWvm7qStMzS6DjgS2onQtg5OIYwuspg4vwmeIb9zUFecuE3fBZlhnhcCHXVO
n8v9yBZpIKRqQ6k39rDP/byrlNjxrdMryFw84kc1frJS1ZenSTqlwJIm/Qkk45GGRE2xlX7iQLap
HhIOpR8PhUY6prJUs1PAGbbYgWOB/OGQWn33qL8kfALAFM/XGfg2QXgyf7Lr7eFtXqxBqx+Bo38U
Xuhplb5R6sbZfaaOtYycrC7QKsHzCEgCZUPQeevIqay8NeMhJ2+oFiThaHI3VE7x54mIXrqN7sYD
AIpSN5TTl0i0m8LcN0dSLsGZGDYRqk2pbFfClB4Ca3yZW3mfdqZU7Bp1l3AAfXw15dLnYIulmmlD
NMZl9AUP687lUgyF+iyVgyjntskuE9OPUexs6lo88kKSiqGt9XK2QsKUXWSOTvMrBj4HyWMMrOaI
3+e2sl3X4QFEj7eMOFnmkH/zKokKakj2q3zK3K07L12F88+9xXHlyrkTImiTpHDCiNc4fbtS758x
WHriRfepjT7fqCITtxVo5YTbcMyxiw8IoWKyoyLiM+kYAyIiKoa0RzR20bHy2iq8O7z2tB6exjVl
wkX6aEJQ1BMgZADSDqKmLrDPg5ElGn0Db3aykZqimQbDvlkwE+XpqPhII0MLE/KRtlOekF29Kecj
O/dNeCA2FCKloVYmjPQlqf8esoxOTLBj5OH7Q6C4lpmsttPKYP6QwLfNhQ/biqH0//2ep0qn/GRb
qd/vHL0RcBdBWfqJVUAwgb3AWQ4X2c1HFtDUm3OSLr8jXydSR7TsKsCn/VUiiXA269kMxXDw5p/x
4D4LLZicm8Jjmwutud/opKbecqPBqDcqz4sEt9Jmd3b+PuzdEUNyxAAfbNr1Wx5OZmqgr0RN2AUs
Y4pvzzmUcvXsm7NvnmxorEFv3c6yW3EmzZqlcw1MvlXpNgwpQMUbNJvrz4nNR1xuTnI6//uWtmhO
UcvKjuN1cF0v+DQlgDIxA6iQpVaSOUyuIChoyaYnycsVmzwyhgxzTu+mLLAKGvSl2bgpm7T1tJZH
mhqO7y62vMghDwqnE1ASfePa9RTN9KxfaeINJUL+5TNoBtob6SQZetd+PrEuphSxZJkcTHiraZjW
8ltMBz0GowKDomkMLVthDKF4hryIBIEV5zBAI9JB/JRUykQEu2Ug1m5w8dsnqbhfpZnU3/DXX+7G
iMkBupOd5qoxf3yleijbjEKQm3b+5s7UM1tPCMw8c8G3VeebpfeLLPgkJIMXtsx/YzLz+F3D3xam
by8x/NUBXdgNDvpdv4Ycz1zObIwPNGtqQN4vG89kv31kumUC/K6LJcZyqP0rnfdBOXIqFnfZD12Z
+qdkuNrdCtyQNDM5wzeXRzTEKz/RZZPpcTkRp7J+Zox8LRCZlRi3MYGJ8G4P5hNjUFlwXbOvENw/
SSFVJUaeCQTXUpANJns6f7Uj6PSrgbkNuY9eFe4yVMdYoIiVor97gOhbp87ieJzQABfDoyH9+GfV
Bxdd4XViyLw+F/OCQOdS+INg82VVnqmM87qAMpqbjMi+gLImPD13XszwmwN56GN+xMWFFjA7XPRA
KfOpZTT0hB3/XfGsBnpmG8kPKA3tOfkQo46gz/vWsxaztACDrnAC8J9z4nkgVtT3jzuqQSKUCNC0
lBERlxKkGsTxTXcvmuYRXqwh9qYEGs+HFoWClM1bPnnwoeRTO+OUgxaIPOTouUV3eMg1MKd4syBB
HXdLqRhgtv+eqsfYGNkB7bP3Xw9dsQ/v+Qzwfhj4xshl22gUbwe4JynWYPTm+r+TdqKn/pb79B0M
JxeSl+HhBsZWYu/Ms8JFwYE6xEyqSJf5/dk9C189DZc8arrIdJlE0VnKug649lD5+bDUw4q/pcyO
8G4r7tD+RtHgQQ7igqmTBQyf3xH7sejOrRy+wQ1/qYIJKp60JlEYggVbDNUgzLze59FLoL/aD5xi
Ni5WLPmCrFrrEUQ4yRDLfKbPbg6XcuUYEAO+9qW3JVw6alsD+Puo79htnXaoL0J4QH6b+bbUbaaC
iF+2Dq+qGDapGre5pJfnS9FVdvSfUyzCsNsgKdEzc+SUex/N6gaY1jL3w4z8aPL7k8poIM/6cw6x
te/3Lgjt9QDlDfclueUw93uiuKoJsmtdPPvosqQZXn5MRET/a7ff7DNaQyWYlKuzZrYIkGriAikb
0t/KFK2t2pg/5QIhdpsnqEvTzu8yL/Q0LKBGQHSF9mwDLYvF1xkXE3lmisLrmYNjCqN2T4Sqm8ZW
RbMI53wraJc1mIvDqjOnzoJaINn4xnF2IOWJ4LZf5wEotnTmCB+JMX7vC0nG+ZMzOWAOK3yxBGff
NFv4Vugj+GFkxlvRtDspd9NPquC+nx2+9T1dr/k6XJyw9Qk8Gp0J5faKrzdIHKlIydAYCgoxjZYI
biTl6LfvJ2auaZbWcMOTR+mPAmQyioKuUsOsstOIROPXp72Y+DuIomtWHnvetXNX2oHUelBDR+ih
641N27A/uxcqiN23+QRb4tzsnjQlhH07wogmGrO43ODyxG+ICFXXyM+ap+AL7MU6T/G7zAc4I/iA
Q6mzJTqLQSwBO0bkeShAjIR1lzLJDC1/MqivdlH/05J97mjukC1aDCDhrVNS6kENqDKJ3iSiXEum
Mg4YYNA8/tkClyrNp7pYnZ5zPwMftlQhuH12ulwBM+blT0fayAaxUOZMLj/VGkNTA52m3gM86xOS
QhssMxC2NwHfDjf71tzhfiev+ddraJQqbX71u51NLvpCl6ZJrzUyQqnTQi21vmPyH7le7l6sdkQR
mhZ1CB1yThawhRnWe8nuVCGcyIO629SHk+Rc58Nx8I/tsRX1o0MGzaJlkff6LExGgeZyNopTMEfw
qlk9IlJY/NnuYTOW22d667N/D977OqtAPSfNQaMfPmYkDzTzxTW1NttH+PBEhW5gcaSdvusBz6Vk
Sf66SuVy69tmhKw/JxUi4qudYNzwOr+vb6m0tVO+jCDSDWNa6uQ0G9KFwAgpkfC6o+v/QFihGy3A
8j7o/AzTjtw83XANVYJrwjsZA4tAMtmogwbrmOrsvhTaV7S2W1U+pvA+Cy41rFjTbzQRB06VUh8h
/E2PLOjNhmpZra4roEFPbyUyQmkoFUX8WcRk0izt0JfU9ybnYdEFVowNBqo1t+2QnsIYqCzqgjBr
+rP2G9giyCZavMn9XnWPgpEYV03B0kHOY+qmwV/mY2tgGvFzGsU7MmDmyYRNvUJqn8v9RwVVNF8p
F4YRZqA9BLSEoEjxXBAcvMnIQQn2Cp6VASfCdeZOOalac+i10E6OoopksH7N+5RK6RKBUzrAZ9J5
O1JwdOx0PUK7xjnkRDQmyLmc4SkEfzQ1O9XkUSdGdjBCN3vRVIAlT/eZ4/rW0T+Ff+svCmN81Yfy
V5tmv/ZB7um7iighONHaKlgZtfcDV4XXYhshn2Yg6N/pxGoCW/z1svhFbsI/m4kPYQgT3MiGiOIM
SKizqlcIuPwUN59ovrW/Lr1dJIC2nfoeR6JECW6+C70hvHr38Ol063R3HilhHDe+qYlBAPuOSEY2
aBAHUIC/lGy7AkEz8xcUoGJDIvKKCqznj+4lihVRLI6jlXit5pzgq9TuTnPFl2B9grq4mzeMowQG
Ayg6xQeCoCPdCyXr4wTTRGR3syAIlBco5S3i2R+n6ebskrq9cz/O/7k1GdNN+Qj2bSCwSjrstlF4
I7nQTQK8gfQ/iWEET7zV0YOBQ5ZBAqCv/EHRxf5oafPKTRnWlW52On1ICnlkZX8yYDkePVKlRtey
izQjDjP034WLInC2+XBZ3QQzrbMuiuJesC/ZzmT3ueB13nMpKnrUnaCsPmjC4xPOqLdvHDNjjZz2
LpAPZU//cGHmeg6OeYKgDIK2nR/zusrP5+TNXPUfy5MikCo6OJ1O44oQEJpX4Pr6hQhnlBE8gMAH
28r+QoIlpf6h6FYzWvG/jtgyZXtSXJRrl/2OtpkKuqwOPgVocdWT2/njtGn+JM5cmChUTMvI+NFc
cLnLz6sl8lxuqvS1U15VY9gA8trJc6MeQFlIOloSzjlPTtFzAL/Ykv5riE+AqxqdV1mwx84aid4F
Y8QU8tk9XbaogyXtRD6XW4JJnxja9KkyXLs/CEoZUsEyLRspj+klbvl34UqeyPJIM5wO/3M2/p/X
s6vFEyLNmG68ISi3pMcGQnM7ct7vc/RgspAyt86hoTD1UDdl/KB0yi6SA15hoiPXGyzCAsAFRcwm
xFF4MOKh2UOLZ3GkwENvznhf474AVd8luG2umOOE6Hnge6dvJEhQ1fS525YTIQHRcgPkRbrKA5hH
7z+GbaA4lnZpZkQDJmiOi9fWXLxzPQQ4BPZBUJhwpV72B3v/V3PKF65vw2BRKKEbHwb6NsqICZWI
f1/ietuzlVIfWszMAqzSsRcbQc63dW6FdMed4Z9YTUiWKJ4BvrPpOah872Y2G+hCskOtnBpAhP1x
0g5qb6bf8CmQQqxuOaaoxn4n6Z4YaKGurrGWaCHpocPHViX5kHkbABmbhumavwrmcPbUk8Yuq5fL
pTd712SHJDKohvCp6LNgjjhFX2J2FiL3LEHHCTqWttjurRq1qgMkjUxVywE/eamfKD8vs7hGRg4w
tkpUD0y6Mcy2UZ+MZgaqxZV3WlaNl/FzM5ogu+5pvg6yPFPlzTMSujZ/qXwuppQVRRXec2u4ucC/
RjTtyHlcm+ueYElkzv6cnBsvBx4DiMCBvMkoH874k7xpxJZaNiXCPot69OhZSKAeuWsSodClMwnx
ZXuZOFF1DquXFbRk42V3XKPvTHLMSMlyOZvZyVeUuIEKcHXtkYXGRU1yqx3FwNtmIBwUXGSooxWB
CDNhqosuYUETjsKnb96KPW0eyZfnz6jKjLlFOySbDtjRPV84CMsID9wYwc/W+5b3+6YOe1+vDRaI
mWHWO3xQV3hVqVUMuUABoqDqEp2DvgSXAieaFeDNcHXD2FdmHO9K6DUZIS3kkoanlqlTQBtkQmep
V51GVE5bVE7x53soMOAJqV6Hok4dV+0g/+OqGVXseM7ggYJhxwT2fPicN9hrKtQi5gGnOxO3AH3N
inK1poHLFS6lV1IM0/b8ZBwVH1EkMnWESOck+na2LSqBDsupTRgG5CPZQTH+R4jMVXluvLRxeiAK
XNTVU4Kk80kiquazVMNViFUv6M/R176fMGMJeJPMXtPFnZX0n3jLy6hcSYih+JMhnv8/7o17JE72
uQ+O3eS0MJnu0hXrQBkNuV8Mc3ecFyfd/GLsdVMb6mWTb8RCAEtrIPxyfXPJbc0IMT7s4oJH/jgR
cilZjW3X6ROWSYzcW3oAN4rxBxOHmsD29puUrbO586MgYeUCZjdr9tLyWSsJrI1/lgi0gD1CcZqk
0gIKQS8xRV2UUTFwUQPKn77/OWmeOkiDGopD1dmkDfLbvx6/w8BarObZjX/vGb5sVwrkeFIcKkq6
2rQUo6tMHOBEVVSSlp/eMNl9YqIqIqIiyhBBCNPXMPHrdJlyBxQIBqNZIaid/81d9CS3mn7F1f5A
NuvVqS/gFbbAWPJ6Aa5c0hQ/pzimgauUflN6AN5uyt+wjy6EYz9MqrjaYhQIPcBwb8Ocl39q8dTM
lwgFEZid5wR6MJKfJ2w35431pnFwKsXST8Xt8ndngnRQDdVV+A89XJPnQ0MDyVe+13pmK6pkplRo
8NtnCm5YwPoxYQjH9s37EqSzWW6sA0AxmuQmfulnNbTcQVLAQNNIW8WL6w4+RbfEaj7HtzLUOWFq
ayDb63FG6V8xbmEtD8iB03hExMNe/PVeEXRHo3ty/eS3r6Bqd1fZrzgyLeBRLmCEJbP9kIXUPcec
C82KX5dRIHjmxI0RwGF/RGv3eRIHD5jnSxwSQaQ7ZmRFoc/HKqW7MgZh1JfUOns76iyV5PN9zuMI
WxeEY3iLh376gjyVahjPVaJEKBirVbjtMsScJZwJCevLql2wKPv9rOwhUx91/sMrIEuePF/1sXxj
mvP+DRFF6uyfaS8I5LPAR26EFoJzPvpg/ANBii517yo9/mrk25Vq4TcmycNRLoIoAIe5i9KL0ppt
CXklHRXUsCM+A22SUj+wq0kLBQtQ0kzqR6y3Rblk9cbu3Yo/4T9pC+oRYiIluS5OT5hH4UZOVxMh
PtidZroK360fJ/tRNSAwrldfDiJjwWV3VTswEOMrZuA1wk3+7DTejjaZ6j4p0HZagqlwuWQ1iEQ8
1/ZH9FD7xpQK9mRcJkSw7KtmBKbT02/NHRH8IS2NgnPfKatiwzATIrogCbnQEKeb0ITLy1OXm9TP
HSxRVULYbc3B0MLsODrdhkDqt6UFj5Eg9YzxlEMntG1xth2qaDYJqkAa5plgDm7rTpao8cg0Mxmh
h1Vo4gmu1A6aZZQdYaIiaOSS8PHY6qe0fP5L4nM+J1NDVi0a/t9bBQ3JrWqWX8XizdCZAeWsRMZD
6wDPprdB+4gEwmiJ+gI4ftTTcb43SSeUYa1jcBfbaidj79Td9yQ4gQ6xHoTCZpj6NBGTy08lY+Vp
bJpLZZx0KpJ8vHlhHgKUIEWcBYN58PUM4U61vB5KLLnk5ilEmzuOR9n3Pwna8O/U5SSdeebPPF/J
PChLq6An7uXV+t5VwAvLfUZ1G034zEQkMA9Pr1lTdcCrNe4OzCmMK4auOmR4yyc+vi7xl45l+rU0
VBC/6dSYrfw/FVVdYulw9sxPuaeQc2QDSQJugDBAn9vflm6F3wxi7cxJrVQaFQE8J4pDxnsYZKTw
tR01oFmgscv5k+KIIhPoJ9/OKzThQzxbjPC33pY3fSrLui4R/KQ4mZoSar1WzVdUy4pvkC+GpvXr
GDuImPV/oIOeuKD/Tr+Z9ACxIh4ak4/PdaL3p9dHU6Qs4NTksSA3AGNEpaG0iIHDKKAshFucISYF
3LExIhru32OmH6KFKKgRhMm19b+0JV4calBySyf+leyk/MSePuzYNl52oybk5SquroQ4hCMjqJFI
vvFLU9uO64QBzCKwR1FAdKMl60u8ufjaw+siWWmm18oA6QDiwY3huCGv0potWYMRfRP7jEabfMH/
zsUhqT53aPU6QLv0YJmZrelL9E4PFHrWICUJhpNEv6xnAeZX65n2jRoLUH08AgjnVkxOvqWKOiSN
cDWX30q2fQ9PI0546pM9Z4xEYO3vS29WlrcEKxeOdQ8hP2aqEkWbqz3SxrcBPMSpXlsax1iRizWq
ZiNSrRCkxfKL0XdIRBk/ciKkOw2LtbZZxbEMS8mELupDFO01m1H4AbkzyMmr9Quhts/Shbcgs/CB
UX5rCVl/MQiNu0sHM5x8R9L6/kG0RY+ApuJtIqmNnTm8ys8YygCGY7rAdScFB124toK2U68cY8nf
ZQ/6XXg4+GvtabcMOikn25ROsKh5fV37GpzB70QodKkN4JIi5fSDCWt9K9tAPsJlif4wNvHwWc/u
5F+n88ErekRryzHSNea+jo05NeORvh67qZFd1LscynRVrUyzEeAeoxvdh/edHLI0WWVDyMmFLS9F
MTl6AIinfZw2qY1zPtHz9jBygOaDxGCsZ98OjP9hG2Z9EZZNLN6b+AYgYLrOzpIc4DQW5Wn63zNn
KtKDlmcLvnM0lZW1PenqtLqP6OK4fODA+5Vh/5D25UkF/hctZT5FHO1itoYsdrXxuvKMpFNXn7TW
VA8hlrB0onPhZ7QrmhJxcNwV5r/m+sdibw3BjK8hyN8NbQqjio5asTPURzj31xHfsbEpe4nZopHb
rv/+Ny06WyoHMfJr/daNKNu2OlnnCwHhmu9pk3/nCbnb5YKMDO3y1mpUCt4l3MNX/5Xc6JI40frp
6X+DFvkVlfNKg+6UfyCpFB3hcHnrQQC7sAzCmj9M4OUx0S1FXFrsb7T79hsgUr1EDLHtQMbFl+wM
GfuVQigqOe+Rr9VS9svIzxCALxsnqZmhI4A4MKFS3sgPBSX6MfGZLjt4SrBcYY7CDhe2Zf4g+w3h
8LOmmXxqu8AIptLnsizPVA4PSQvEFzfBeFOMzlfM0Mz8mK3ayiUkoHQmwV8IS3cDtVzmT7yemLhh
o/VKWYH/YhIhYqJZRuxdbp01nTMiEMf8BcW+b4kr0y3F8UW4oiegkCHUm0SjtyHkiLQ3GNKxinZ4
u/hx0JU7JVssP4F5A8WiNYWHwId1CMnF0yxYH38dK6JOM8CGlnzn91ygMfrnlNJ/fePrNUIIhWE7
yGAAHnwxBw9boFJbK5zUOADuAgLIJvhKSk0ndOdZOT48E0STJ4yG7k25SnviXcHKYiNnOCmkCKGg
L+rrRo1Ak1fxcawPMUTXO+qVja/DVcWcQgWzD0aDZPfnaFnzasB8osMNFspBUWSM1LWCD24lP02x
S5Fn028u7bFZN7q4wVRA3uMiF4xhIQeTbr1mA8xZfURaP2BH/YIF+UVpWbcfTB4ZrwBTtTtLezJ4
4iKEimVnLBzFcQLY+SVMgC4jTdF/3PwZ903Q1wBHQ3Ct0o/nHw0u7o+crZwYXX98igmlW5MJZ8bh
vt17d4/Bmxs/S+FufhQMnGPgqj0ocYhlvwSVNGdF6/77Q1mEEhTaowiShS+VLBbPqNUne6SpJuw0
w3FNM6bS9iIVTaAixS86RqqufoUN/eqJ6oRt+um9DTe/zH92bYYDO4i6fTBRBCzd9KPmlUIkL6Ly
r0fjFA6Wf3tUU4Yz9HEDgCIAwrg4V7O4hkhUi+Y8EdZP4jpSe1GvWzKPUXRDgIBJ5c9j1CXVnXa/
JDIuwMyjf+g1LNGwLzGrQhrD/VkwlqXDncqTyr7Pyn0gpoqGp3wc4b3N1MYxB8yobegP8afI9i4p
i2CyvZD7prdyytCperzIqMAReKamoLafvJOf/i6sseHuQj1gB0HbppEnr6ezUNZdhJn2mmttcsrd
hfHYYYyWXffGaU1qYRowImNBftD6+Isi+H/2AKfOp4tUJ/ban2vIjH7K4en0dTpyoIbztcB2Jzvh
Qaux0/1aeJtaAnMa6VXzkLxaHf097y6XarVUFqVvh1+HgYZbTHQfI6WJz0TsGhl40QDE+PeAJu0b
tlp1An3gWwLehBcnr8b3nOrcI60TN+YjwE9CJbqX1ZCj//LeKrpJOHSqkINAUA17vXLvkLJLxQu3
gSy8w3GONhHkkiH7Un6wDhJ7PRq/k/vMqJcvG1kIAWPji8vDFw37nUUeXegj8VNhF/JegH3MQuv7
RHIWmwtl7PbcH96JJV4kgNCzOSmwzTduz+keuiUxRNjdsYSCNWobAGRaEC4z+LdsQSGhdDbRC0Pa
yS1NbSFzTgcRk1iC3SFu9aoJV/dG2OgjZvbQVUtBf2mjRJuM+Bw982lS5kAm0jTA9bo51uVirWP5
ua2drTaNt0+6gjpcQgyJ820B+BYNqRK5237jjwPh3JGRx1A4e6Zpceh3+Q+2kvomlpor3vcWFW5k
+7bznua+oz7gHxck3SW3xM5zc74o7LfQat8MCe8iYJJZO/5647wotxLPS+0znau7nksMdzjsy8Jn
gmWawuDWdML2ikXo65absYvtlNf0OldypCJRmiO7w/6BfCvguI5kV4Fpgo1Kv+BnXnQ3eJKM7x/R
mIsNo3KIwyGYYIUkjdrwc1iIdFMzUpjSVod/CTU4FQRmodykcltZ2WI2LsI/SP6clA00sRa8/COf
qp+sG4SogFJ1OJ6L7gS080mJaX2IT45/M8TE62ii8K4LS+qIJczG2ds+zHuwjPMsSS6zsIL55M4/
C8nbMmYwE6zexel03OXTz9HQXTRm+obXT40aoIGSDbhGOtZp4yzJ3886f3DgR7ER+g362JPzQKi/
xna5tAsl7+tQEdcG/AzJ5itKNVVPUKrcZAnoliW0nYcwZdo3rp2Dq4eLaDkVfuYw+E9xnkZPReSi
CL+2hy3B3kiIw3OYwy9uAnzR1luQT/AgL0Hyoz4ItQV421LDYAAKieveY3Tf0/DdPu0mWJsIHFGA
BXuaGSe/osOtlAAkh9dG58Z8hZzrFodycO3rG3cvSJko/u99cwStxtSP4YNjkysfELFG/HBGUIts
3Bq14nAxoL/5/RzEJhXycwn4w0ynYRfnZHKTuGvYsl1nd/6EQ/4TIhEGkCEIRvCwTy7cVZKveoaU
vpnRMlQaLVuE3wN4OudIkm4oKzJTT2+9waJ8zXaCm2xbcbFprWk7URA/tdSfgxukj4jkCKBwdNDW
Ef/j5ClKvr2gj3hG+nxAySgzMGuhMOMf9YZEI70redqPCJiqsMBdpM0pBaTVbSD6r5jQ1rYGJ6ia
i/ZsbhYANQ0R934YlMjg+RxGsnPjsLdEKC/quTigWL6EE++WU64uG6ewOsaPoHEV67lDFCgcN7/e
6rZu2FogzX7azFIc8dCAFZMJ3kNVdgjCc/cOtfJ4WSrB8CHWDr60bGUkIvtZbxjJ9w0+VW4B21JE
UzlJuG9uqS5hCMKEf995AbW0vuTK4t20zxNr0SH6B52cCycXStcRf0HcPbjgCyhm+nV4MWV/ytMO
466+5O/XXH6Db8p4EHX0+F6GNcm2jUCytTNA5AaCr4ixMWqjd6GO05Fq9jPF7qhycA1mu6s2fbIx
jHR8rCuQpHVjGpzPWLStGtztamhcIEsgjQNkBOkhjQCQwsVs5FmkrxqnKJuq1iIkKlaqLvG0YH0r
4GNcu3tb3wa3hldbc8lrHwGNn650OD1uqaEWSCWR7cBHA0BiNRxCVGe4QclNKThHCuE8iKmdhO2S
neFyTr65B+mni45d6ZKf8DJcgZHbqA98NcDL0AW3bIPlkQw6oUYW3NLDxcxVEs3sBQBLzsbunvvw
TYgCwugJOo7j6WmOS/sGKiCwsrk1Kehk1KjEUlgud2fgSur0gm05NilxdoLDJYsj3YbwsTbqMmHl
KEJM+sigUlNyLBM8YdmeeMjAfvCJR/CHxP7qXpoccBujzjnk8NEeJG9gh6E234UN2JrOF2irRmOa
5cYVaFGRnq4Q9sff6pv5jC0o5uXb/qNX9pj0BEedKrFWlIPGAY+pITqQ8gvH+Gj1NUvMNuF+yErQ
x3xttzU2/qzU6tsdktMK9QT0+xLWvGvClmj6EbOuoUPLOmlErv8zckgb5yfqJfIwxGPX90KngEZ0
OjAYqnavFKj5H7C2zv9468XEkLNrn+93KGGAGUq9VzyWDkAvMvWYFJgjNk5JsDkHHJs4v6u1LGtA
upPsahi55rsvhkfEQAZolqsI7me/mkeAk4i6k4jdwFW1jn6/Eao11WkJyIGuAF1KC+lg9CY2kwcg
AjDJ4PCqs1ViYBxG5+kzvvo5sJfbT7x89acfnwxIT2NKKRZ6kJ15seK8nm0A6zB9nSEqeQD1pmP3
U4LUt2tmVEn7ZKcQqF2n3oi5LGPXwaLTtbkXpVpm6Jwbmdp8H6SLGdbLnZ/pd7V7H+7darLGoaSS
WvWJnq+gtbhyOrf+y9ksj3HIi30/ihbsiK2fHV3BFbnLo/mpe3pPnHk/n9xcVg2I7Hwdk1qzi8XF
y1q7dda33HnS2my7s+Af5zmVn+gKLvjBOcczJHYIPnF4Mr8dJPc0fRj/HGCQ7UV4Ae2av7SDvhhb
iiRkWp0Esq27WoHjIJxdM3+q2/J+JtXQxidFMA07OP3eAISLZln8zUW9c/AY1w3Op5LDYXh5i/sy
2fB2EQYcfYYBFHxTvMcIubtBwBpJdeAhbRempDLxD3aAHl35gnrDsFPawLzICg74o6My4G2B82Gc
v08p4wiWkjTAxR5pFfvM6ggXcBVwI55WX6CijjsU3kKmw/ny3qhEV1KgUe4ntKgHFlQGe63ZM94R
gX0aY+T9s87RxbgI4kFihE5WyjjKZbMzLcs9Yv1cbPbnW1xEphDRAfyUu+3ZP7Ue4DiRzs1pNmpB
KGGkr+BfT4GWInoAXIOSWoQOZue6dpWCfVXhAwUkWuv1502aGCYUb2OFdQKnMTdlgcR+Z8Pkv9MY
4ZR3dRoTW8EcILflMgK7BW4eekffkHMrrYGyH/cwkGQlZ6BC+UFYrw+qcY3z3MMj9/VfEnBuWVp0
hZnrXCvtrBommf27r2XmVTdYS5fiPeeHCTFF6YUfrOEEX68UnTKgqz/Ten7Dtnce/ohOOOTC8Fgc
ftju5mP602ub/8SnlhmCZp07DAv04Iq9lmCzyhrHdiMgjBh2nSUnW5Pojk4uE2GRtZ3Oi7GK7IWg
PUrUxLrOCW/CkXPncCDA+gXxaO8L+fwkibIYdPW3Uduq5+xj6ecHLpMYxiyKt4yq2b6/KduUy+fL
V+O17VFNNqNRjxr+33IiO3YOqZmZVQXfl9nX+xL/cl7gYe8fv5BWTPAi0ViqyvvC01ER7gzWv76M
IoKYzOHGAKh4vuAOgr/qMkERKJuBGG+nlwxxLYCJ3SEunSqP+B+n8xgnZHxswyfnfoDoLkJK7lG/
giBs3St1zrmwMOkBFHSd3cBJPko0P8+/iz6KhPbc7oFs/8YqDudOpupe9WMmfnA3niLIG9XMXdT+
s9RIJdaR8bPVjksRrwuWnSlGc0tgN2zNE7g+ldKdqvUFyXah41jsES4SCUia31DwX/TecNdxNo4T
/oa01U9fxIIztXQ9oQaJLzvTayu1Nx5Swl7V4ZsrGYet5E4iLeeAa/Xra7L/rpDZYSqL46GJ0Vc+
q2G+Nv1Xv1G6fbmOI7bjAjwMMkMwKi4piKhd42FY8avVKnXPqt6OFWjSXipr0jfem9vgLRHp9lST
r1CbF/ElP+XUd3ufcjICKFkfgvfC+Q/MK6C5XL3MmRrwXLItsgHB/YiGUGNqMoXR/t2LV4YXrKQq
sjiK9QsiGxTGA9JrHfmdBUaS0pSCNELGWa0SBAwHYnC0dhcrNOCEWBJAT6cc0gzg1W7M/9QEr69r
0B28DduPM2ZZUQ/tNgdu6cnOqI7FriSCjolSpDcF9Eu+14O7WP5zq9KwstTIDQQCLxVUWYTkXYer
VS1mywAo1sOh+HW7NuMUx864LNAjuTAxkzmz82RzUkUawiWIRHypsFQ7utQ/MH+Xl96f/walslvv
BNBUxBGF7gDaWPOMcdF/6roVwZhTrCNwHsKZLBY59ePE4iNPkb4gIP6jwV2ZMQO5DnzCgZQSkxfG
y/c3qxMnZchcFsDgkshtbmSwl1jdc4bnQrGVghe35uqcEl0yoeOmdn9EmRl+1sZabzdu953jj8pQ
wAed91CPilj/B9E+KXEVtK5juBQ9DV8oNUk0v5cX1W29nXLQ7Fw3EzF4RKH9J8MArqthV47baYEM
u1eGItPrtaktnU0HKRbE85EBF79rNV4fepr8XCuXjFM+ud8DF+mKsEMRgXoAKD4dJ8EfLuajIJGX
lb/bFP5ayqGI6CFKPj7dx9Nok3hnjqjm66xjOHXaJLdfZtfvjj1LSm42or8WfP+zeiPhqrtXicGf
/UBe6Mf135eipiTS9KmwjWGDpWm3fr46ioqRJM4F0lmZttk+otj5QYBF+HlxrMlossPlhQKN+g+t
f7nsiVPeUPhOgTnJIcbBSqa9AX7Bw9z8eQsmfqKHaeWU/xerCDhJ3r+gYutvN6HG3gXORmbDbYdp
mAXyIlYiN7rI+yQc1yCPZ5o0L5jK5DJLDx1gpo7Fl4spEKNdaSLlaXoluGZAom+fDDugGDoa0NX/
5J8kyEaVEewFdG0RrpjlWKVDhLLftYyfwd1JoBPCJQGeAG3U6Tz1SYuJpk0ws7McVCkbJNRRcJGa
c8jwn8GkOWoIzdCyuZHA06LKEEH+LMeVP+9LBewLLWtNZefCvsJE+JTzYd2w3Q9GIYzsT8t2FNCc
HTN8Qfmga4WOwjbKeobB5wdkXFDgLkc4OuFFlREH0r3wPXwssoA2aZ5C01syW9evxbLPawOfvi25
7LyEv+1y0d53KJHALH0HMMvfI3Py59Zlq6Nrw82xIVVNG8zp153i02J4KSTFtxD0BIvGEnyCeinL
MNRzBuBgUB3SRgk+Pa5gMzEAcoN21U9ClMV+4JkOjGb93Ye7lV6mWvMRWn2AGjKfBz4ZA5ogmUsd
1dDSeatR0nQValgqNoYq2zLX1khrybi3mDHH/SeAiFW+5ZySrBt3p7C/+VPxeZoaWyG2OXkhqeAp
z0ADLbx/BoUju7xWXLSLFTFzPSaZ8AoHe09qwbOeMISttpTatg/9D9gzbAeC6iofIa/ymMWyvpaO
gbfK87uv/PIQxJxs6BQoXnQkJMQuWekEPpUGj+bj+Sd3X2o21Wk8SGERJvYLeQNv+IO9APS4zavl
vdDYryTDuJ/apG/v0YDebx9ahMvUbjlXT2S4Qqb4CU09ewnNEIIOwOTPvBGU+HF/T2NlKAS0eabX
DhpbxBKDOSLssSZul/d/+oMP9GzpUr7O+UBtqDP75qrc7rF13tiyrPRAnvyLQepC8i6iAUeeFbMi
kGd/GzCr+LPAbVhFlyRGNGUNU+/bn4ua2HS9Ozf8GPWExgCvj3ym/FJVDokQOmabqcHC+YzYfj43
yko5duUdyYlh6eberaFBXwj87C6XDFsy9IGgFeouuJp8DHI6wcTGP14nsftKamqpLdqPMyRoGkZg
C6Nxg30eRFEaSdgUIqYROZoODTsyXkbS/btVhFgvVVTv5t5P7t8SF8oQX8ZoT+2KifPKobkq227C
g+AROiUFwMGR92C0Wd+zYgcp+wwDPBgReQvkvcYBCP8o3qpOULLBs7fxzEXJk4n9bb5ctK08hajb
mxPmJjTJFdVven9FwohA2sr4wtCdUDhmIlIxbzppQQltjogUArlC+5g0bNreT5foIEGr72yohyu9
LjV7JwMHBY3vjH3ySEO/IN1/k/PRx5j73PYe8NeDDeu3t+9qmKT13KqZCkaRrZk43dlVvU3KjDW7
kglGiE7uwNEvxQdaGe0i51QdVTm0W/4kDZBSHyz1oxJ82fqw7GfT5en++sehIvRcSQr39OkaSqtT
hf8mRP6vvYP+i8dBVjXYcnlZlUT48blPY5TSdvGZ5lMF4bR28bNiZfSIgkVqe4BTxtiuyz7ImVDb
cXPYkzWM6t/D6nM60S8ldVvccgkSq2DnJTjWI5ItpBft2QcEXsY5cZ3qqBGxcEhlyleViiExaI7f
tCfidegeiuJGhitSWyhMLW8hxqJFlkUFVo9wowB62tmJmmgz2cmST8KawmfNk+PfWnMGLsdahIxQ
LoQddhvpALCln3xQDzSNStAlBYMqNKMLXboEzxLVa9cVXCxgLCWYhHy4CWafX1Lp78VePR6k+De6
jv00xC5bOiKtgF1a0lj9HVWxOAy8qlCpykWMs7NwQSdMPQWv12DHpZIOiwEzasO80jkrI2FM8a3h
opIW3ou1HhNBjPKNDyy+fZNKjr+FPRSraV8TI75TcHsobwZ5hqIVDUOjPhShoi1rLQIglCfKCCfy
sxyMXGSGpKz+MSREuuWTcrYmD1oUXp7hVSOHpndcsEpmempP89RI1DVtvqg1sBKRlg51VLHf1TGA
mhEkyGeRqVb6eiPtf2pg9/SCrMI9LEBRXSZAaaKR5OCAE8/iCj/mFuelxo6buyNZkFg4lvyvCdLw
yY18i7EAK728pAAFlvioZrLV+zwTC4Te555MyH04U/PjHBfv+FtuP7OHa/kQxLb5zLpx93nIp8fs
tyQjR8bbcAp+Ltm6LREUg0Hhyda3lPFCteVnSmV4+NJQQgZS817Vdi94A37PtvhWeer6TtlK29oA
WnK5ykwYoM4sHkTLCfq0Gao76JmXAwvylGU9t4U+UzTV8eJprrbwnCLf1X1Yal5Dd0WG3vayyMkl
/vMzbuIAwVl8i2lpsVEYD7bF0b6HZhy4agVZS+1J3d41AG/sq4Rwx9elMfjXTv0e5AmAODfjSLyH
IvgopzNEHDdY++3d5WMyhZhrZ1dfZiHw75Pe84T+EMwJ0GLE94y4GMhD6DfaHWCmnoOdk7QytByL
jF+XRVrNMR1LTUF/zRyEXM9W08J+AAcq6FHd8PHox5gOjnWAvnuJYpWAJfU2duJ335lOctatr4dl
W8p28IWsb/2RxHM+red05zcjAKXgObhIAUGogArJTKnRaAUcvFVyKx3ycwtfB9J9GhahCin8cCVg
ebaYv94mq/YjBzRU+wUmkxcOX2G5G8FkANVTntR9kp2p85hNxCRiDmR1XWYT1HplF6PfkNf6a5Cl
jk/pjrXRgye5dLrFslIG3PsqTufFZiCOv4dfl67PXMoeBaoEe6pbsK+vjswfql6R46VcuJl5d6Rx
KTv+tDamyTnAUS5w0aaZBeP9m0cuPdvEo3GruJaqHk9VS08r6Bk+FG/BLCrr9rXOTEp9Xab6nHkW
wH5YtZaDKNzOdVdxDzhxzE6uIz+L6CY6IdovNUBZVYb7PY4/8fFKROLJRvxsCor/Pjz0QHw66h1/
iwy9h2b+z5+KxKjZ2Geba48b2AEHB4xCVFtuLM55GviMkztB9sZDvgqdgMkaTqtx5GM6OVYfD3Vy
NDZdHCjHD3vHYhGPh9iwcHixzdN/qGMFmD7nfgQxCFSMQlp3+R0Ow8cL+Qpj4kR5c4voHVtyC0iS
pCI15PurDSffxsvISGDqt7C6SLZ1YqE0lVhP6lScX6aug1LA0si7uSHbQdniajdF0GLSCCeruogx
9qVJrMz3CIna4AMZ4PzhFSFqT3Muk/O/SuY+GZ2CfX0U/IA7auGZqbHQ5BhOR+dXDJvuEbMNSjFp
Rb9/g2Y+pY2Iox3uMAsL8CxwduQOvaaaZj5dmM5WIwSgqXFjwZ1VGysfrTITXU2HDDYe2E/5FS8L
Z+yhtJgBhqZg/KJQEfDxfpuj+P0ZlSWVLVmJpOevN07UWaEUZoqfBQJtrPql9Khc78OCmZr8ddfS
khFsc1mm83UIug+HlKRvbJ/zEoxM8xIlme1ti9tfIknKjo2Kxu8VXzWFJAQtRAnqT+yXXkjNteNC
UFsRrBWfl99DXMhoRvLi49myS/r7UqYcgohI1mTpuXnvUTn7O12mVH2IDwiRa36HQNNH3/DtlPn2
xvaEqbQSfB6lshGEAsSzGQMVkaSVy25uUO6hyO31yPrwyGVZqr6WBs9SvvLsNM8dnVIODTdNhVRo
DXxvqgMtkwK0FFMgt3s98DL9K2i90dequbl/Wd+dn1BSTvdNwQnGQatBPwqnbn0Tx17ZA2jjR1D4
dfCerUfpi6zdfUn7C5z3XDjq02j/24pEEjpxgrC3NvrqN6GnJeCdrSoyS7Oys0ZTKjh9oahiczB1
Jwnd1cnjwLd/xnScbGGEK5o0NrKi9S6OG5/BO7eH7vs1qwXdOVf8olFfrcYAGbZgaRyfx0AEDPln
y8W6ZW2NOeOWf3RNPy8hbOlpuz7dM/8j1FjkJQgag3X/dvVR4eJ+cGlS8oXo212TFsVOQlVF4D+W
sY5WRpq5+9p3OInufxa7MKXuN/dlKC3l3Q/XhgSRKxcxel6F0l+C1Z2hKOAplyR2kSGUKXYTManP
Fe1FUfoaSO/5mcisD4CmaFmLXywgpcLH+UUZg76GNpubMg8xVQjVS50KYiKyCQA+jMu9ukcryH7c
psdg3CkkIwyuXUaJEM96I1SYaFQ2S3R4EDZISEjsy0PwAhswv6sb7DShBv6cMBkKTkBVxEWQ+baB
Ql+wqEnAhvp91A0b/XbV3SRAVmX23uak963PBGvrJswqgAZbUmmUeFUppKoVDlVxTrixlvPS6AT1
ziBLSxCoXZZwHxpt5unl0WspbhBNEhML0u1qvCTjtGTjbTY2cHvnZp4XYVIAf5HvM4xUv6CJpt3N
dWZThlD2kpsSjpwfKi/Z39YN5a/PDRUclj8kOsjFEj95k83okXXlsF8RoApLJucAJ4NSVWkx3Yw4
ir6lkqJPRnEW0D/bzuBZD4FTq3LYRc49HxOXsmbBtBL9RE+qsAigJT2tKMU9i1hTrN8MNMYgyz97
cBt0Gt+t6by+W3lUNhEXd0y835jaZh+DnFmVq3pma5O2ksYTKk8rGA6J0pgcJDiilQoDCNHipjQP
sAswFRPcc9J9qBLynQsiqqdIZOuG271H2QmXhAbSe81JVHBgwW4Tm9XmJGV2i6IZvGb7bPYv2T36
QDgN5YEF3vA4DaopRS759fkdSBzqhkskmLrq+OyUDIKqlNS+BBBQAf/71AycE+eceQx9sxM0J865
TA0uRHlASRjwl5ttbPowIFpckdHl0P0ML0CYmXf4QQT6Pb22/pd6zhLBwIpgD7aKTHgHnjqg7XJm
bQVTc2IzFhFpHMhEvtkbo2r7KZQb43/MjOQ9wsq+k1uuHvHY1NTy+hUmuHRbU7DX/Ag2/xewJpdd
SAwNOzHJ9Wp7op2GX2kXdkY2ecBNLqSiOazZ4ca2euDmheo66X6T5p9DiOK9zsKPorCM5sRXl611
zj1LOzg8j8o7gKqF7zF/N51kjeqI2cPwE8SUlUDXAc1wMqRk08YcgKkKzpMaOgdwrzOFIjKy7pyk
8FSjsv8g5uJyBpfJT/uxv5ym50E6hgIRb/hh/94xtvyoLo/wYmcGo8SFzB4KHdpI2dMHQ1YAfEW6
xtJTfwyFozPbROd04cfqf82zN5ch3QFInXkabAGj32SuDfcvXPS4EZT6Ux+ZNLQj1cRFbT6h0oVY
FWoOzWLezG9LV2lbXc3rCo3LtANtyGNN+18PgTLg+P2XjHtHq8+c1KnDRhtvhv/lkwqUxRHRNMpn
CykSVL2d6bV4KTTRx/GUe2UNf8y9VwsJqiVBDiNQ61x52laWtYv3kJJSy3RIpDPnk78b8XPR5qeh
MZv6sHRllAlXPm2K+vNNU6nu3/vDh7hBv5gIc+eV7Qu7SC9im5hbH5auCdrnPpSf2j6DwpftQX0N
1OoQkFOgTEUeDB1cu6hX5t3tOK3sMBbottlsOCnNF02tqqCVQpxCkoFTM93Qgv8b9kWF8PODcHrS
StpHN+xK4IHeK0HZy6qz7HHO1QB9JKeZ30+wi7H714vY+37pLAOemKssQtV80hm/mfvDwvbqgxbN
me63ggqpPe+amFfNfZ579jAwTY96YfMlR8Ot/2K+I2HUkRkmzipnRPuootGsmTsJZdxTeO4X7Ah8
O0rY2ebg4gMGO3M3NPZ/t5p2xJPBA75AEJuygwebTklRI0ooLCUlb8YA+dBAz/Wu3MIayvmi6nol
Yj9JNqZBDrNEd1M3ZVcsL24lz9RS+FTrhRgZW7K3bLFv84apl1CAshzxVDEEuGsEVPUrSdTY4WLO
7XhQLg//M8ejkmBM/n71B30qT3a7nxMKisi7AyBcXLz648NyLLUDXxxnrybTf8DIdFhP/FWGj36X
4lWqkaXcMTEDfkmbXtAsVCYFElaJFlRrfDXEN20Slh2UUmxauDT3DvGgGpdpznMO6ZcpprNWd/cn
tcaROJ1OnzwfjB2bKUZjluScD0WMkDDP9zl+As2SJ9CrtlGJBLmI0t9fYGH+4ThzvNPVjJn44W6S
ZfFvWvaUYkHhYRB5gmExmcFfEfsPKpcsCaSz/8Cyytd9KCJK7RVIjkxM3FPwW+jU3gaAPKoJbyJV
dRWBFgk57mvQLOKH5g0X6X/F75OYoNo8aBULK54TexunoAVm+hlD8qJzWjshFxBM+e5pMeKNl4KM
2Vij9cbZE7SK1GGiU8cmTGKHmXGq0P7Dg6V1b7b+U3WUqq863Hn8X74bi8wIX4TAXgHlXCMDKse4
gwgdYsFppXd8pnFCOe2WIt41G0iqEyg6knDlqEyBuUJ5lE5PdXE0fJo2z7pMwMbdX0GpSM9he/jn
L6g7NOrWIznIIfuwJ/DvHMJfEFBv4A8jQ6XK/tK6JSy48LXyymw6W++XS52cg0ZkMjiUu3tGgCvB
WkaavmNXaZ3ELhHt6tWcC2MMf49+33uwCDrz2YsEQs65qiBkQXKmpsAYWbd9nrFnQ2JWZUfFpZeh
tc+CUx0fwovrUX9wGQY1jAsUL3UGiStQ74lbRot8aYGEovnh8YNmGIE0+omBNqcz6y9EMGPVI9Lr
O1/YVRjKhubc9CaXpyhzwCE+uHfzJh0BOGCr3WSGesDrguwQBABQVZGigkQqpi/Ty5EZglIEu72k
DZnXlSB5iFCbihEYYLBb4nqRzhyINk0UVRt3YX+Xtf8QeakaatdNk9uybSbdgLUP4kN/YQHyZsiY
Z1EcquY8+ohmjcFLuXHJa8n7BJ6TO7gaIUMK15phZIIS8v+W/00BIWAjFIl5bVaghrkhUTQYSEUN
MlKI2HKjPyBay7uI8s8whC60fAGsCl4PXd95AYaT93hmd4p6wnxM/toWXAWcFj5U6N9uzOWqsw5/
zNUJNdMtELircvHtZJ2nHJcaLSKXj1PnlBGSUJlsb7s23gxbyZikW3juIdENCTiGC71z/HkcdBEI
SqnjeSG9hDMflUXpqKAME+O4YHcEbQg2kHEZ2hMf+VzwuxdDU4UBWpcIMRZXStQZiGMYr70kwF15
XAGvDygg3rUKbzTojLIYAv3d5rNqT2+0Rmu4sM/2rBGZrwkLzeRN64Nm/b+vCLZytdFciIgMPNTJ
HXtf0QpCA1j6wFDovE6yuTU8y6PR8dIbEUiq5SkHZqrY0dqPW96rUFqIc6xz1bttAokH+mn5NuM2
zLJbfb3Bm5OZSsR2MiLX5jdkaliUEqAYttpQTVSyEqUvvOTjwRjkgiJELVztuWxuz27rm0oQmUvd
uyAdQ91wcap7ykFcw5xUMce1xTJAkkfrUEvX1D9rGOzBYxQ7rtlqtXXhhwal+lF/E2W0Agu8HK8o
h7KwZxkliWiT8NF+Qr4oUWWi9yT/M4vEF2K1Rwhv3dDriklTrIJhZ5iVE2vyvm33rK3JbUEuPolX
jJnCypvdS8Ua7ffvUtfgGTh7xIAcH7Od7YZ46LQVSsIuE/CDlMf133V6Dtx6JbbYYDLU9Zv7zTyU
8t1R9bNVtRdr/byA4d2YYv6Cx7bcqTWB3aW8C1EvdOMxMv8ybSFv42BoTzD+fegZO67eT0YoyHl+
N31yZeTMkqCSRb4bXEaY+7GLL2GFaY++kmwgfmse9DORzYQ2vwkKXeIER0VXz/r9K3OQJYpdCI26
tlCHJA+gBSNrBGy+nJr6s5O6GQAVbUZLSKS9WayDcxycz7fKzpGkwA892cBH+4G7hrAWKYGdnGpc
2Lokexj91QpZnK9sQPAFedQ0xalRDN4Lo+Lrl2LzqfLbUdy8BZUZ1cslAodJY7mv/XI5L9DmPDLQ
zk9Us/Ik4i8QVEDgzmShzXdq+REX+MSrV7nVrIt9JZTxwAtU42eVbxcibJpFR6kivmjabGRztl2b
O1BZDACaTI8jw9LgzSvJQCftxnQOykvwevsoCAVmoBhmkAWiK2gNhMNlhhtREo4+dFX/B36CW+Zh
iI4fRto8xhEK7mMDrMsEjSDzqG6hCKp/99MuOmhWCbH9I4ffgXwD6k8FpZmjjD0soDX0aqw/6kDW
+SvQStk0ZRjYXK7y51GyWFWdzZnzdjN8dXly/J0tQap0AK3h7A09ahjsCe9ug0BASNx9Mh8WqUDl
WY0fFQDw+AzyDBk6la1cZJUeAP05SW9/qhXybatgmTAft7i0H//r8kwLnKtSgDyzhTKykNWdO0e5
/dNPPZwHRqaNTOo7cX6he3aRw02Bko3Rjt1VomHWvQ1rw07M/nHPEml0fOGqXenR83vhG2gpMYIO
BwKJs78hm8nAfefe3XKCN5uCaPqgeiZXkHr7jwrKUJecjRaqDYCtYyhSPd4bOxuV4qvG8kJc3qLR
561iKz3PvizW6ScMO8NGJTemDZVNsJ6AOLnhGVWaIFTqh3EaRxLj2wryT5cF/v2zIucpkJl35LvX
KzwFYDdsckE2cvGLBSCgrLruMRAVfsHUt0GkcooEVLiAupmyrLUPUF5rtHUkRCrQRTTDPdyLi4ov
L1m9aann8xVlecmPam0JPYiWVhcwDRq2XACCO3Rjy2Gl7C8+hR7lEinjwLckMlbQyDFsAXDgdoHO
i8FXjN/Kt0CyMID5cUOQWJyQZ0T5Jj//BlgqmunftZYJF6AsGW+TiSndqIl6hYdxHpbsIz8G7iza
O3h9WLEv9Y7EtdHX9wgCiRBoCHnkpTqezkqMP5NTRa6dT4PyFznx7XKYC7LIpuFeWgGFfKa1WNDu
ErnIC/Kzu6DCeianKPDxids/ZwehJbC35p7V4uNqKOm1HLVkjPeG5gO/K5EvzI22TpPacUjFJ9Lb
1XjwYcHm8uaERxmq9LPkxO9kdWA64ClHYWDIVln5NnjhabY5ODHJX6+PzpF13EumlVFXp3JDKZxh
9ZQWnm1OY2faKbOS74wbaWYdLaBNA/ZnHA5U7E0xpDlJr3zri4cDSfu+soFhHrUcv65ijI3Gh9do
IRGZEVY6Lx5YOb6z4oA2OdzUAqDrpwUbsvDxWsE+NSjYNN3+KTOJj97J2PdmfdbOPeuw6eAsPYfT
vciutlmkR5kRSGCKaImExM2Vkdr3dUxvhvXKQhyI/MBIzbRieYLtjooruoTeTZkyB6zq/HREu9P9
H3cvNsG7humFxClnOveu2R1f+W6boD6Ub1Po2f96M/M87swlVfFCYZ++EI+Td5h1LpTcEZO1ApO1
iKx+Xoor3gO+B7Q4nEmJXimAFCgCMQuiwhSrvonu0qopgTDLnquSM+eteLtyz+2hiWPBNK87cLfj
oKBf1e8irx5MBuBRzO4af4MmkN8RbDUpqzbMLegeQRyoYejorFWPDNmJzIl5OFLAvDNLI/Io5FLm
QhY4eACqcpbCICLx1w8DDzzyGon8DibuTjtFMDSoumpEJPQMpJ8VriyZg3dbrfNXdIJA1wqJTqBc
OOI7U6+xwLvhNgi54bTvThVE7cWy0r13GnfTZGZPp0NErhrfhjBZOjue4lA2GCTOdY8O8IEwMadI
HoU7dxO5A2InPGkGpPXpv/EZ8THXRyUmJl1RLLWgd5cN8azZ4PXrrWYWObARyJnTisuq/wS0fXXA
oO7AHXLaaGpfduDjAcRaUjGrKbotbkKZJULopRqqNr/bTXNPkO0HlWqt8UJgXVQ8kbo4g4zASlx0
ZhvqBNJcpaoxmiQLm87ULC2Y702YNPlPf1ff7bC7WuwuarFTdRxAz1M2fB4LRixXMF890+ory+3E
+X4kEGNeXoX8dRTDsnja6tAGScLby5nSCtzxFB5ZFO5pruOUW4O//+ortjCOuprZtzhbL5HFj23U
wXFV3YrL1GSL6oSa05Wh66yu2YntqzBaJUnekrxfQj71RQA9dCRX7iGwjaG0t0KT5cis7NJ4wf/j
tigdwwK6FINOz74HN/GaqBafjEUpY0NBP5v/bIZC/n5rlC2YkRYP3+4oDiLMm+1wLiZNvX4mJy5V
a3DY5n8nrCcYntK3LaG5mvw6XhyT7mJ15zrlkwNDf2b1iIx8UA+xGUQDALh7oxbATvYWJwMqlVFV
C8k71tHLRipm4cOA3GO5VurA3SKCh5KYNt87cR3+yIHdu/H2J8ENKC5UVLMKe+rNds5glqUTtv3H
sHNrdl99fIwKOsei2hvSOwhXzDo4vU/Ejx+BW4EqkGzZZJvUy44PUl9KWF8VRUu/qWq1JjI43OiP
JD5xh6lmaXJjUVSv8qqR1hO3spLy569GdIWmalWlfC35VT7fc0c5038FrktWTgNBkj6Esf17UOa0
R+pFtZdMvL9kj1lpb5Sfl1EnJQWcB5OXu19RZBzUzBqZdjFg04oqirXYbGTOlCP5NPfvHUfFewnR
lnO3fsUYbCfJ2Amb9yLgw1MYpfOIpLbnySlBFXwkziOV9+C2tWxM8fdsfD95kbxONFDpWBV2cA8t
dUfGPwKhaYNjolGwyRBHqxFTr3yU9jytJgv6EYpZdL/lxAA1QW5dMoc7Ca2fOx4U/gi67KLRdVPn
tCP2Yj7F4gz2aBaypHtLOddYQYDmBEX56t/hdwV8l8NENBond5Hz5rFLcvVhwdUaKQmO9fdSK1PB
RujwT+ODDTelooy98ATtNMKwcMau7aBw11OABjaF+Ts95KyJH4/CMN3Nd3o7A+jbHMVGqy6LZW5c
nyGoW5V5ClTUI5PfuH4PvpYmbRc6aQYh4Zl9gouuugaWnw2QOXo4xTFXBJC7i4rmtE0qHaNekXCC
2Tru3Tw1Ul/2YW1WMYzVehuO92wCAk0BeB2+MrKHIMppaA2tIzCPKV13KcX9gstz9Qh51+H9a2lh
OLmdKXhDrw/gN6pn1T2FzbQUSlZrx+F/n5wQGjd/XHgNtNEnil9SkkQFu8PbYYcfgk6BCDGo0a/q
3cn/WycHYdRMKODVoiIcC3PvbGP0u4b8ertGzdT6TkpZotFA0D6uXute5gU/8qw31lmd3gWzQTzf
vUQ+OrhswLGhIQoufIIwvP8VMfs7L2una/cldcGC955p4D11NuH2CUXLAI1oV/bZI5Ry/rugQLyG
zCCCBfYIxX8STp8J7Xr9IlEMu8VUGljCn6arzlyy5e0z5xs/SPU0kzyYasTlLPzreb1lhwmHwlHV
LiIB3OyJ6JlHk5kx/KifeGWxGbGGAA2X+35sUBHtHrn3zv40wIq1n30oH9kfcRbsYSNxGHDf4bve
LPITftLoGQoaJrYB9rhv4bX2j57841GyTSzqbZ0J1F8JxVBWxmZaPvJpe7sHi7c+H1P9Or0xrJXA
Mce+y2PEMzvxCA2CtKxMD4lIINa963so7C62HUtwExBEC3KT/SExKObrIAsPUv5GJYGOske5DfRy
4CNji94u0Kiy3IQ6ke4yuGOi4FfBXmSsQf+u2iDaFgNKyerHm8hiCMM96zmsbD7PZMbmE+1RcASk
T8HyiVzUi2u/UOxIl7HicXsaM5rmwUcGB9f3quKCC7KQFpwZcbZtmomBTdSigSVtUokEhEa2m+t0
93GaMSTzd9SQg4OEVIJkgb+opJaW2Ft3IrExDtFvtDmXGKS45lQWgc0W+rXbgibEHrnzWqwZdD8G
wnsJj3z3cdddvafniz+b8w2Yru1cvi2358MVFeKalKeomarSWKl4HnOjnrHwB85dwYckE2bjFqXW
YNtSR484SoS0r6DOXugr2cfm6TOaWrp/ncGgN5YRF4As4JGU/Zcs6PYkE5rG4aFlIfUY/XOuE8Z8
TQ4oQPxhoztfX54fA9T8dAMy4HOFKGPzpqzUiqlf1wswCdBK9byqw+rGkJrREfFwLQcCSqh+J6To
z++xdLYS7Z4v9Y+qX38ujZ2B2YJAxoxojAq4LlintQRqUIhTadYDWUPzX/Y+E2B/4zzpw6anfZUn
sBNWoiVKuhsUOYZ/++xJqoWmW53c9CPTlm564z+RZpzhLk9YPGVlraaXD4VvYrs02laS0cGjJ64z
plcBKaoUAOHLo9ooxTg5zH53QfWWMyAgJLEgeHA8iR7LcxLoNikHpAmQOp6ppg3YFJ3RAP4q3v87
xh6jHCn1f7iAKn1aejo2VaxA4PGBRW58GX0lFgfJmTpm8183S7Z6TduqvIz1GFWNSMoBnAD109x/
SCZ+isxSKpm6R2Yr2nkUMMvqPNy/LpNWvZSB9gb0yohFkUkyVLJM0hGg3Na/Fn4ZnI8mIpbnmusD
Y3JGp5Y8SBwzWJYqcu7/m6sUe3hnvlimdrSe1n8WMI6TdlNIlSivGb2Hcy/jxQDLMWE1c4/8P8FV
/2uZzgfMZoQth1Rv+9VX4rGE4w1mv4zwruaEtJf6Fy2h4U+1DsU11khcwAy4OKfQRzATGu3FzLOs
S7Fl1dMVB1e9kk5Ja2Ilq3bi0SkgUKGYCCARlHf8Cj4Jo0ohrrC8eB8retsJwfdqDLrl5l8crokn
worIV8jkOByedOVQE+uZug6nLareKSW05jpckrACsTzh/yK4RTHxqklLzriTRzBWL5GtnkS/v1jc
7nmftolRJujDKUztbT+12ap/cD3Tu6Ypy2H3XshMgC18qF0QmRaQTVj7oJG7fT0NU6mG7uedndRV
0owkAahNZqTKVk1Go91f1NeDWcUA1eoDy5SVh7zYorJElVshn13k24OTd/Qc8p2lUqMRnuael9F8
eMPE/d7g6QgOhL0mVfu+aEm0pDday9onI+1/iPPwg94ZmCEDzLG/g0YPJKZlXYloBItN8Gn8Ft8x
RNersKE8W+qDvibMElriaqYI0vgFegpvVoNZnNYyVRwtlF6/PJ8a2DC9lDWy/DsMYvJSFgba+0ZL
OFfZF1Sfm/XVh2pFivxhl7v/Gd1DWWpcu76AzJId2r38KqLeay21e0WNbivmmSOSM1NRhB1vpphS
Xq4E587gIzC4YMpbvDxe2f9pFqe/teb/IN1fU/YgRmTnF21BXco4NIP8oUTtutk3ZhOhXRnvkXXa
7Dc5gXtziv3Y4BvY6cHEQPgs5ndyLD9OTXiZaiP2ddmH+K23cloBo135nqTqarRBfRZggdxcggiI
t4p8JWklraBZmLILaeP3CT9hKjYv5qcnI8ZBvE67XrEtrrY5Z6/pNR/IY5F14p7faG+5ac9pHn7/
f2qUxq2+yK3f7O6E8PZcM0Ln3+YSImGwMPcYaMvoDJChWmAe4StpxdNkzJ7Iulqil72Q9IjcWDuA
XLfha9X/97n7F8Gmf/84k8X0DlarvAfzan78WoXZIujDDtaUk+Dy58oArRVyLbCvMBabMTbRCxDd
LWnSOF3D7fJwDw9qD3fJeEwiZHL/HzXqu49PmFsUK6WrMtO31GZ95jgLLBwuqQ6kzAOLeWCLFh7u
LVfHKQXukicNcX5J0FmF0J0ZSuB2vXDZ2v21OrbBjkl/T1B93VusLknG+ibVMPi5mOkVIRec7VpX
gyYn05Eu/RbvK4RNVPgjkJm8nHJushpBL6g1LLCzqxUDasI0UQUCrrcy0iE35RMdln+vcpDtV0kP
lpvPaAL7fmMgDnEy4JlOZWH9HAulTMiIToR6ROSSUbCXfrhHz9Xr9qH7OUztfMAyMMuSvnTVqLQG
A9wmv8QJBrwJa1Cf8yNLYu776G29Ur2bAYZZBEvedTZ81sHAtM+O2/V2LvFw0ptFyOwo5j7XYFiK
JBzOogF+K9GFWBq48HAF0rGEWtZ41y0BXilXGs/mnJ0TVd+A2rKIu+PQi2zSA7fBpf9Imkksxiyp
OIMdAyRYLfuNYD4eUKEbK9gL2vZgDmv+NJ1ScuWm/NcBPorv2wxoMw0VoFr1+/edFwrEocn0PLhY
duQkruLUlQUOSSQ1lbie212umsuxI8D+Wuzb7Ei8AI/3pbNMiVKckUxfIvP/A6KD3w4FD12How+c
z47LkL52CooXb3xtiYiK0KXMwkFpSTpn+QLihbgRslG+JEHWSlCwZMfR+7zdTjelqv6d2IHBRKqq
oNnv0aNk0/1D96I+KF83LHxSs7hQ+7Vqw1BT84sZSKNygDo7rzYTU32TwP6gOk2qaQRLQ+uHFc5h
9gr/JuJ/SI19Qvx9mT2CueYzPdp/788mHVSTyOEXpgu+/iPOUR0J8kosDRRqzKzAs1pLjI8F1lKr
Hj12Be+zu7p+7AFiU70mwStcXznJnvIIdYYqXg/lWPxRfpdsiVT9yKxIh80mHNpvt6KUzk5ngt61
lbSIO/LxN0XYrt5VbEwSOrgowzmrSoZ91/n+eSgpZXfEzJM2oPNmIpBFKnff7qG3Bc8cOG8tzHTa
MpcXjPGPYtv6V13UWzXfFYtTSsPMrCmoa5aRZdVXe2eEEm3/z+P/B3LSi1syDrz5kW1+Hy55jJ08
eXQo9Egr9pUcr0l6Lt1wFJN0WocgxlDWBfaJsk4VtA5uqtjEH3V8XgbRShZtCRQu0v3L4PwiDzsb
vtZXJY0eLNJABiVTHn9KsDa1EUnl9PXzyIvyV+nOk0vvfukoMng9APafQkZvDkZmeUJfvi5jBSMO
Oaraqw/zRVbQzDF/86cmNKAJX1fzzgs43+xwCpYQGnKF09CvA2bCX+686YAgFz/xDgqnzbYkJ32k
+yb8oyoKFvcRPJadA7uWvQiFrvolyJFyFxxABvTMDaji08yClJbBvtm+15xpPb1pKYBvqirjMebX
QIelB6hDxtNWxuncVjgRPAMNky+Q1Mv/HOlduNGBDIsjfsm0Fxz90TbdkCrUgz3gYL98P2OWrrPU
Wd+ggRJB98vedL001WFzp5vYU2fBRq8aE8RD1NPYjF52O5oR1BlWeL8pk2nQynGNphGqZkFKpTZy
CwqI5/JfO0NaAqwztK4zBvzxk3jI4DtSP/ijBYOaGWuKRW4irbioikT2VTysTkiWTV3sDw/M0EzY
nHJpPe/QAfpRRUU0vQ3SUUon+ibWAsoay535RaBpMvd5sjq3iGYGiTll+HKaq3SPrB6QJzf+4U21
336jGrTVw7LJg+RUWHg/tDYhoRP6N6ibqwWZzd+5Re5TQRi1nAxsLhshM6BaR7NOjlj6KdeUzHGp
PcAqUGHAG4k6cKvVq4lB9P6DpI1nCAH8dB6/5xw0g+3VmvkZbKgqEaC1kgGZGSNd4Z6MBGvSeNBG
PaSuykhPdxTl6n7lr7ierHzTWLCkw5xmMO69Iw7FKNTAk1oPnma5gkyQxLuEJz8yIw7iDo2kUgxS
FpW+b7B4BPeZS8jpXupdmGA23oAZwjSaNek6W3LnJAjPZwrb748xDP78JK8+Pqiwe5qRZAwuLc7F
FCsPE+Z4csrj2+1l3TfaxVVNA8eNRB61MItsnEYHu/eoaTLKo0BvkiA8ejBxhoMjwfU8kC0HCKxV
LLM9Z/bLqHtblU/rR164kiLQHSqUyZ6iXnpC+kSwAMqTw4R22xZmbs2HTL80YOQOvc7VeNUd4scJ
zR51jEXWEw502EGSHEOvKR3gZag490Ch7rBn1o+J7uKxZVdOXpRswBxQrnANsXgk/BtBzikn3r11
ZOPIHCv0fH5qH9x42nCs0jU2auWn+hGSTPJj+IyyN/a+nSEUB0oh05p60C6XxAZjiyDE5ZNl2YgG
qI0icFvS/SgxLfyUjZFK8VG4NCcznjwuycXE2UjXw6EXppROQe3P35jGraU3Z5kwTQafe19xDfhG
S/qpMqWVH9HzerPphP6bz9bTMtEFF2YZ8g524H2gnXcYfCZLamHOcpsF4mJeEEV0lshLRsZAaEPT
C/qLSTaSbzqLsm7p+B3LgTyXVuY9PaIOHxKFXqB1Xdl1mZ5P6W0VZclAYRZUB4ITpBdI+OveYkUj
xllTn8tezOPi5QOzKzO7DMYRolxyHi3fp8WIcy67dfLB16NGSxBvJ3L5uN+Lj9qeAf75jlb4tPii
28VD/zJCnvKRzZM73IN4lGQ1yKGSw7DakshbDiPjPnS61MkmY7QLWxxz5ZPFRQxP9yZmnL/tgRWL
qLtUN1/sYGlTdSaQyHawiNlxJBoTLUJwnuogtRO2N9idmA03Yjv6jb0ucupQtVcuKSLQ/A0KzhZx
nj3krYk/k7NUCvBHuzjH9cFiVxdSqgxMkcwsloZUuva+E5A8ifrrAA4DI6vKWkFXh2AqkZRwEio8
byWMyGxek8/JA0Ms3tAtuldtuDUUrd0W0e5vK9S1OckkVjs1uV7RPU/7x791ENLqH8eR+enAlO8G
w5ArYWeZW78gKsElpjSKUur5pPcVhY/JFV+5Pg4nTN+4Q8HNeegrsfpCAByBuPhUnTi476fMwys7
f6nS91DtI56J2jZdM58Q74ZpFVK7nFtDNGyE2yljwSwHmkUqiCPAHZuzbxv0SzUlDpxojcbat9pq
yE1sge8dwhjAkWAScpsWwIhT9OH+iwBfN1kx8SR/t09XmQ+WTzxPIq+8upGtkFFDtdctIenbILBo
xQ7MpNEVEwFXIZ+A6YKPfiNVgMyVLL/8L6rUMsghXh6OXtPF76mYpYTy3T4tG/QKniW9T31mz6m6
ll5xOfKblXGqQ1Q/2N8iSAVvRSd3UCp7VjdRzNhagZwzqN4HCkaGw8cXRnuFSV+0YYnsLG7uqTly
OcwBpr06i900r2T5QM9SVhx+oGppnKOrhkJlEs7eUX6VZkb20KONsnlc/i7rdizdtTHu2BPjGaH4
4ryPkX2pk8I9EVeNwirTXK+Bt0W2XO4He506orSLFcvS+47GBfcNa7KUsTpA9+OQLKL8hENstlfJ
LwDq7U5fRhv0qH3OTXSJOGtxtX9SnuWBiT7E3i6dHOEip9pY8IKgABINKuMH6DHQtQEgTA7eM5eX
TZ1YLY/n7JcsqykddA3HdPM2wTx/7dx+dIEFYo2RQ5GUT3A4HSEQu5u2eP4f4SNfnQUR4xuu3m/V
nNmBXq+MexBUXTAWyGbyJHVm1u8fvtOQkSn9+t5GCVg59eG+a6CyZpTvjwfJdsrb6n+Nee4FnmoH
wgMDQMse5EM2HFGHumDJcK9rNGS38cSKX8p7MLJB+EJ22dlkykUz0Wfp7QHUTbfuEFVTg1+YeqFP
PO73AcftZ15wMbKV3wvAMuqZstqlps86rQ5yAgLK6agU3vXs1Dr0d01UlJJq1l9qay9WvRjrRwbm
Q/dj8rp0Ja9qhOHzjU9DX35lDvNPlyPwRJecj3t6E1thhh/fu0bR8OhH5P5uxJ/7toM9bvibRaqG
eJE9aO1rBsf0x2NaFm47XYubIKfXIi4IZuYEJf88eJgbXN+kTa9ttHu+sqqvKE8skjmhAh8s63W7
hGf2dob2vTZePtmCv+/OYNVK9z7G9imV4iWIeKU1KygAawFJllsq8ETbno7cjFHYHFKltY+E2d85
pYXQw0+r+Te6J+IXdMtEW/djTKIQBWF8eFJpx+wk0OKItjWbojkZ1mtC5MeaJArTaNO0d8gjhVtF
cfEeMX2fXNdgCUTq8c3C5Rh2woXbxLEzbPnPv1RWQ2q+NbDKrv9wK0tfnxpAg8m+sd7g+zb7wUqf
jFxxr2wxyBr+J1R5LpMoWGYLFzqyJ+fPJOnqq17yQupl5hiUwAsZwOPVVePwAtljmfYJ/scm1yRX
culzvOpWUzrTfcXQDBofIH+SoLjFRG0TxjkBARmJJiOMQupUvrIRHEh0fmndAR9KrDdrYFytXfod
2DHSdLofO61i9Js3DktKldeNHw/Ri+NgqIZ2Zho9bmE/Cl1PcszgbcnzK4V7bhz1BoDPl36RsdOr
a5OqCBd6uZApgwsVWz/5+SUmjIRh2wh7blXd35hyuYZzuo3/ylGfNPYn1rmCm4+B2swBEB3kIdPj
rhvwFrAZqVrSwgsKtZcuruBhevgVhe6PsMOtvRULOy8Em6ImjNQD7kY79OQG8afkwHPw8sBh5ZI1
Arx5EPErWMMxEYD5jNGTxuovjHiakGNTRimqek30dNtJGA9Ki0bTTSYRkdjE4gzAKcdgwUeEr19V
Zupa3+gTctey3HLkL0KAcVsRdXdWqVGCtV3UKYV+wz76oa28PE3Zq9lYinMdI2to2GjzEh0aKaay
/ZoUKHIf/XA8usEMNKfXds44a/VBYSE0mvxmYK8pM7+5rNQC8oeJUiDEBsgCCB8loW1IJLqdhrO0
ocIYMvnlehYl6A//tOKV3QklC2nw1mKrvo5u2Qb9MJ4+LklwUe5FWlXZL2S0uh+U+nU3BjNfs5am
GYv2MbVCRuxA3hd6ChvN5OqvkLD55b+lTfTgOBzb38kGwg+ORDBlrhsCDva8YqSAhiwp4lrBw621
fzPmp4EwEzdAgXe3fGpCfU+PbDwPS/4ebZaJMXvZ1K8KGYM15P2n9FIC56SOvgliYrU3GBSA2XtV
ErqXx0+RKyhAx7tkjhskvzdgDf9k7M6ZsK6ecSbqvZP4euLsovYzw7HOpncmzN+xVJABG3gKGxHv
MSMoKUZ0CEtOoCH6IpCk0dboPXgwqaef9nQ2LPxV/7ixKWFvgipnxu9tZRNNP6Ppu1ZDaIUTWfh6
VlxRg1PSuOhPOoNlXiHSnibG5Du0hoYUdhSn7PAjPvoDXBrb6pLQ/tnDNiAH4FfA4uzoUcMBiLEc
mUKN0tj4xTseddBe9kZFIj/2+SlXKJb+o8L/wYFS4//Rs9B5lK6uFCdAKk/5uWwt2o/1PM0XPvKk
RLxk5Ev2FtyAQlmEFgR5tn+obQU/hi56CY+nNDrJvVXsGcWlVxtWy3s33vGuhp/FPbGwRp9T3/Hy
qTLzDJY4NkEtIP9ZTfZfRgpkn6djAMNQrPSHKWbX7y5tqqvSJ9Kv2h0pbcv+q3O8+I6j64AshMnR
Ne+DNFLvYzWAAjrqvQ6YEk4hHVtni4+5pDAkkYYtF9tLIAp9LvQfklNVxNcLiW1ib1rAPgBr8/CH
av8f7o8e7bfIUfjNfqI2N6IQB1kgJMN/vwuJ8kyxEDcTk1vtzCD/Ir4FYOq8yBEHyxO4B90XAdEn
azeRw+1tgWgiyPGuM4bj4VATgw9cVAtNYEsRcD6J9E30kW4EmfE1e5PKTuqz2JLIG6qT+CF7XHKn
SR2xHK5sSfGAc/3yUNItaIT3x4duBLQfwj5oIJbQSzsra7JN0wWYMEEs9jonZWCWYP/U98BNXUTj
hDv3Yls7C0uuubPdYeMmWtxZ9KjjUDNbzIHdGODHhtSLkGe36aiKKbNutBRmfr4zU5CcA6UXMJO2
eSnSyJa3kdU7+y8/d19f2Z7qvVsRvK9DUKvoCZqrQLG7FcTAm1I8OiKdXSh5t1p10y0LQENz8rdR
zlHP2xcrUvGHEID3T36W3AprdjQkHOVRSvgUrrDfGABJmF8DtKWFPWuGu2IfU8SD7LARoHAggrrS
YoOkkxrAFNCvU5PI26cQOST6FZM/o8gKA0tgmJEK3BsHSbJxaByTLVJsJFrhMl7cbX0a44FNn1PH
TkRhvlyS311KtnGVGvsmL7XktPNP+1/yEgHq5i3/d2Nm3F3snza5jJ4G+ovh16B7ULSjFSOduH1F
A5BBwJLXtPXVZwX0xl+vk/FiKXkKLVX6euBxnSea/cFQqLkeuvHLTS3nJa6aMDHVprUGvor+8c3O
i3r1bWbVNb6lPr2GD9pS5O1U0cTPBE/16x0hxSSNL/US9/2dSAkNQpFKLUNCKi8llVScz6Xr27Y3
GA5s+hXCswPLXkGNJ9axylHalvhvSMnMUuBD6LR6E7kqshM0RaXN/SRslWoqpnunZdLqpaqGJkII
Gvm3oYCMNJlLVZro/GN91mYyNdMwfu/yuTwGPSqPkBw4h9v0vJJJ+fvUMXdJLR+5voJbcq3PXY1A
F5SSEAxb7W1RcDxF4RyTZ7N7hNwBqix5rY9nZ6AKa4WG0TiB9pFvlkuYZkCXRwibk6eWWPrbr8ey
Kb651DMR9VunniD3aPQa+TXDBzJySLvlKrLXHJS0xWcKaUy6ES3M0zLs0na3aoU5KaGn4XPXZeX0
ziRMCKJ9S7Q072JDiFOOdzA9uOXhcH0LVg81ZinTJ+kx/jyCDg2k/cDJ4xrX3LNGxMwZ8w7cgqv1
mzPghfKg2OmKbKGKlILynd37jcuRaX+ANiCpZjf0CkdaqUpGPMbonIXDq8+QID60RwHMVa4sMesK
3XIGPytFqEzZ3TtT/aB3tHIyUXNRgddTCKj2iHFS2BOIzYz7gOyJdsClBTFQ8HIirF+Tn0ChADxu
3KreRRIhls1SLbguhk/rP0EByIxIumomtIDnkyRFUBqj23w2R1GBos2AGSZ1/JcdmkauqeMnRmtG
M+KmeDg+AwPSw8UehA4DQ9TRRk5vUp5tmD2eSosHPY8jI5U/NKcNyVF0AXFpE/ZqUyN42fBparDi
f6j0HgmQwdlNO4SPng9YK35kkEeVK2V1DqY7qbU2o+16riApex8kzoMn9yTN6ETRI+zc2/sP3/i/
L1sILqvIgyus35jX+wrpAjOuGAXNGXDPGY+Q/yZtonFekR1HfFdQqS8m0dH8NaeSfEZsyf2mKAOh
bKtrOxMvCCUoEvctVC/FaHaE+SDThD+oNNn4Kiq49p1RX5c2q/AtCDPJzsPQsrvhqcSpOIoYoVaV
AhhiXDfYt3atRdhfMXquRXM/+OdSbu3l3UYxiVoHcmRvcAXijAvECCgdwnILH+KzqdG0ox9VIWLc
gQueug/7cCCeEty/8Byr3AChK5pTW0LHenbPGx6XxUgrK/rtSHZHawqqrAMqLmUAd+E6MKbkrulF
yAEmE9Fpr6vOw/ZxKm2kb+4+U2IO0z0+6cJIQI5XuXJ+uJ/jrP7srA5ASdjtn+qmTCGdLUQkMZUV
V4HWerbipoaSA10R5gsDOjlNNV7qLkJ1twU14cTrgNUbuUg+P1wCll8HUKVc6ikcyVxMYaFDO+vZ
eq/JGFqa8mk1QRoeVfT2KlmzqaPZRUlbRRN+6yr1xITa/L/5bQipujlx6XpMUBeEbwLL5pBS3xeC
sQxlsUNsO6PPmoil9Odj/h5/gs3ZHszJRic2UKw41rNObV2hw3yhv8OnXQHOw91MzrY/n2TNq0Jc
S5JllnX8M6MalTxeSTwocxB7ibg1w4zsLt3ANHVJW4JYHfZ8EDSsyAJ/19j4Ck8QyaRpTQ14mRK3
fwOG5gMnVn6XKysbglL4yj1c1YVUxDtvVFxLROciMaFc5lhKH+oF3cOyLhq2CQtcgCrySjKx0jVv
1/51QXSEOiHp1nBu+BBnNwoM4CTjiYL11M34iUuH3ZV/SN0f+DdfH7azScxg6aoTa8VZDJwOYv5P
qA7Af7J0uekE9LCi+nrdwOW89m+CLsbzGdsNa3vFa77QSACvvIYTnYwGBCs+Kw4OWpZd+sNnkBDI
0boLTUXl9m2fEi0ZXxUBVzUEwAvO2rbXWVhhWmfKLtLagOF9L+X+yXxMS+Onno2a+D1rsBI81CPX
aNoQ5aDwkbVkX5ic5j2Fmf5uCIVkI5GAlxU1IJN08r7y45fgVo1fUzfh0vs3z1NdkSK7QHAscGDv
4JOCGmGm2pu9Yyt/YwWWV8OZmVbAamYH6niLiCBU55XZEeLWRlTCO3uxBuzcjs1TZd4ppdJ/tlrT
L4FbU60jM28wSGBdhetHw11hofoqGt+BtSV9l0roqPUAhNEKYYTLeed0DiUrjcRy93C63k/OR55D
8hBuOSoMN1Pe3o2zKVJJZDT2m0vFov/BtcbsqqRqADc/ovAknH8SJm0lBGjZkk8inT6/lCCHpStE
rE14oDTWPvy1NLcGBt7OUW+EoAmqRuMeK7WD7yAX567a8HRFk6p14vfQZJw7GAZVNjgkwMfmaUr8
YWtOhrE+e0pjYxEZ3PGNDBEN4ea2xpmojvv2MJdwKuP1bZJGYp2chZBRYDMTW3Zyx8MeLeUv0zq3
QSPr+rfUeE+T7JnCsFqeBIil807LL2ZYCNk0LdeVzs4ohpygvjBkrcYJjhZLo+1X1uI3phdTRUHv
SLnpPgCEOEDfjKk/5ez4OpBJJTfGviRQYtgC/Kdn3+LM+k1AOlIvbVCs0BxP/inoDVpEi/+HvciE
fviwuL5DdiwRIqP1cfpy78nkf6+d7ZxwINF+LEa6Rf4wsPXLj3JJAwh0s1obfSpTsfQQCd0Bo1wQ
5DKzpk6bu5XLkVlQkVR1C9GaURayfSKn2FpC2TZ/ULCabgCqRtdSQY9L2kmAxJrTRJGaKjatUkdv
gmPgrVqNHrTaVfbAJeKwAm9T/X/JRY4AEwFG272GWpyDJSB5i8Cse5QOmFooJyFrCZaWph4O5Fal
5cHSxq9KNtQQMUHtYbQa7D2POavbKX80WV9rk+lCL0YjqZJ7rf0Q5WIWeuYKTaVPHctqCxIBDl5N
IiHQppHXCv5FzqxVOUcERSYA0RTJAEeLpNSt8QiBr6INT9Ckxqu5EV+v6UuO4tLx8nJEi4IU/cAC
DQ0Ua8ywYGx6mXpb18724TyqULL4gEvj4CvT+Lfqe6Wk1smnDCizTBtN2rj+Cx/I4bTyn9EPOreb
tvzXsrUFhlbpCuUqr/1bW8ybN8fX0ieZV6jpYaxb04b566y4ihC3A75qQjuLZ6coEtRjB7ICR8LW
aO8HgYLpnsfCpR5XW9ZUKL4dBBTZELjCLPnzwL2QKYOcV67D6ogsZSr5omqVMFTfGJOHJxm/N+6L
D8WCHAqinmsqGJ0jAmF2KmXWHd9S6lRUPQVP+WOFVXAK0o/yoztyKyOLQoTZhxE5EcEPEq8QO03K
mHcZcAZURih7/wr05thrZAEnytoJ48Rsoml+W2YzSiW5PzUBuVQOKGjkB8gqF0i5r4E2L2sez85G
7f1HbI/faME8BP8C6ZezyBmg23T8nUFlXM8dQg5uDi/pDGHZMUG9wL6eKCNNIKPiM0hV2VH2JQ2+
X0tQRYLsv/NguL/rIJARI98axzgJ9n3CCGHbgUgbNPMfqTfkbU7TsApdFo1/RdyDdLjjDyMC2l/o
lET0jCx963yp7W9qnaf3Um1ItEOu9tZvwl+2LCIEd/ugC8PlBu0m3ieonajOe6nQmdnpCY3e6U2d
PGRQQtZm9MNBU2TgPqS6zW8yXC2YUClqPq/e53aKci9yLoXe9sU+K7JFwhyxylCjMX+huY7zvHef
LpXOVIRyw0W/fU1othm5yVf/c5SQUzvZyKNs23iRje3dzGsVkBcR2ygYDo9Z0VL9hTi5FyK63pFV
9Lw9+VkbVk2y3ajaNPJZ+tbVJZgSit9CEEV2tH07fWJJmkW9mnRFypN3WRvKyYjo/OCQSbgVvHiG
SNmUHf9dlt2AmczQvOJZJuYYsIQ11oHwe2nY3F4nZitsa6rw+AbxjZetOLnWicXb01SettYvjwON
Cv4SAhP7WZCjD6reiyXmhtS8DTCvzmqpR9OQ39GpKh89GPb3FsglHjqJvtgCDxRyioCbqkSwW0JI
0FYLO0K277NYoaLh8rJNOHIfqHgMT4/mmzN7rMf2JBo14k5qmkfyvOhqSyzxGGjhW04EdFP4YdV6
hbIw46CCi3py41rWxhUhol4SUDR+eCoFkcxqdab97RV5uHaVR73vhv85x+rGJ6uQmchfBB7WuObU
kL82fjuCuuLdjLRPH2p92FG3y20WE+eyRjLAEBG6COf6urOlB67TAFodpM6AB2oXv72hrGNIACjI
arBf8GBTzf9iCSHC6TBoR+cAxfC206krBOnAmtDjyzaEOHb8/mxj/lzX2X2XKOGuvuKytE9PpDXt
8HKirGfBdtw1quhRWcuTGIglh26DHvciE9/K7Ir6+hEUlMbZjSOgYJ/kv6z9g/hw8z2bxBRZeZac
3h23BtsMo7/uneknjUk2NZbYX7NJDqnqpXcG+MH8iCRtkBho40TcTumGFt575fkjqkk3iNjPpvp7
Xpd4HgD9oNqDJxFQ5aC8B+3pQB0Vm2PCIknxcdEhDAovZT+2wVUuKGpX/sbhN49LCHHzKX2pCAFy
k1ERApTly8G4fOhon7L0sKS/p8POi3j2DOoM46aHGiq3BdrbjIdnhqUwRoveQtcMzW20QaHVGb61
R+A9o3yL5EEE16P2YC9baZPk3CTKtY1kIjf9f6yNIszAau9OqBN1FQYYKvCWEP1jcqkwNU7scwV7
JOKiGBENF21UHSVNfWe+QpAeWRQwDXiGl147L9r6Aq8GtuAKvDB8pKOjFlIRKfP9Nn+KF14nhDRD
0IikFyVTZYSS+RW1uLsEKEqwkQBGF+6Z87o4U0kTZz0QqMCzymZJwB2+f7W6Y2ajKhhQW21/bIKG
CVabT6hRMMJph7OWMNYNDzcRMONKFtNXI3BqDtgFu1JHsmpNpdspv72S+9HVGptHJqZ8mNHOC9+k
RMnuF1/iVn5t35kdgoFJ/pnPQt8ADvJbcZ7r6HNiA9u5vo1UR9PntAlriLJ52NynU9bKqauR0mGq
/W1SDQIaTkvKnBrWA83CzAHxfqdfi1NJXrn8UQvh2K72OI24swibSbtRC++CN3rzmGuWi9dlHq07
vHrNLouhEoB0W9zs89BEx7+hXhbHWH6Q85jpfKRTfUIGPvxUsOJWim+aOy+47vf4422JF+rNDH+R
CIWusOKNS/FGI0Ba6l6CVoAwf4CbRwvTYE5Zpg8tvljBhN3yBjF+PYsz7UNgQd/MluaBrKTUVTvO
etoS3mixlc0DlGxnt+SsYtwQbAtaSNQ0rto67Qooiz3Z3qIUN5HO+KPCzr3wQ7AaO18c83gfI1jh
HjN/WDWJoiqkxKLePfI88HQbHVgjjG4IRjRfoAFfi9nU9jWHRJPf6IwbfcgVjj9/CjI/i8Sp6jXG
OvmZgrvtNOVgeeMjMcbUWeXI5HvO8TZ76pWGt1pCcScJZAIqszu7jRQFRSZU4aUEmtm4omAToec2
Ub2qC+vpsJOzUceaKVhPYvKBXZpnR7BMkSFx0iIUn+T3kgwvX7vW5sZIMFXUmjlGNfUQ2h0AgLum
6ztQ1S7Jj6iidMEt/xX1oVNNkx5Ex7zAhAcGCP5x6MHRKQZV3LW9hmeLHz429ZOdROaZwnhIlJ8S
eJyw/HR00Y7/7i/nLNpgZ6Jjvp+4EAF9Ol3yNmxq0NlzSCRvFdYyjiLsP1wxAjDQCoxQVgtN3krI
OQj4Pvtw4hAg6Y0mDhV/0GlFmMrWXAVW1AGy/aDMlcXyYc6C5kfFp3MMUNkgz3xRWMsRuxYQit9r
OeAhHmgV14hi/GPntgl4JjXuQiJfAsLr/z+cR6yf6+8nZHjqgAWmFfqRa12AWOGwO3H4YMND9TNK
JgrVgUymaLO7Tv6Yz3B4hnz+22NsczdJZOVPbqaut6dPQIRhS0KQtpZKV/qxR8BVK6SXb+3dPlIx
bu4nzZP450b+ikfli7P+ox5lzcuJtbV64wZ+gWxg8qJPjKDrPSkptrnGmEFgGEGVl4+PoO8/geBj
7LmWFwbRDWVXzqzpbpcOyUPgck6ODQ+fPRDH47zW6+Qx30KqnEmkSH2x4K840erSCkVlX0aZT9qg
slox+7YPZlS9V1SsluUrCdCvzS0RqFSDNp6J4nSLa/7LeOmp5311/3d7KzEBsf8hMwzsp0jx4Ea2
5dkQGjmnZKU8Uh9yBxUZ91YancEX8ZkshzcvYX0unQxGLD0/22WCUGHOAKYUGdIZA0txRjeB+l+O
incdkqcIvu1q5bqILv+U/bOt6wTfTQWW7mMqf5G5GVSoS0zcj28S6f3Oi3PskAfHmoiOGHbqNiBG
CFM/qBmwiWr5agNWilLXMhlomDCcYFTNnZKQzwaRTkPkryEevOqe3bFpzniW9WwOZKx682kAhvtc
99r7oMpaxANd3IiggyyfzfWtAtFTnpKKGGGKtm/KZeCX1Z/9OgEhrTpv5N9jgHRvIJ6y2gbtVFO2
yp6LviCE97v8wJ1xSl8BSBzWqot71JZ++vWlr5zRz/AWqQuuWvnpOsgAdZ4L+Y6jo8je463IZfBi
Immg3PscYuw5zsLvBDZ+fcsCKIKYAuwhGUo+/4pEHitLN0bX6cgQn4EYJ9qaLemZTrhGj9XadTJs
9cN+5lvyhi+9Tq1I9qCV+7ssBF335AzzHSTbGAUh1mWsEE/znEkl720zQeDWNZWcsh0L4StC+OQ6
oia6aeQZ8ROAlYHt+uJM04bvpK2BxAW/Uprrs4bWjwadLHipBsMfuqNRDpLmBKjZieytXM9RtTaH
RKhsuvVD43+p9uHL2/ZFpaljax850cJHTe+vR+OfyIEcrebtzcVKH8CbTP9JEIBD8Srpupge7RDH
sGWmSOqmluYyiY6MoVdD1lzbG9qlW1H/ibHkXenfYzevjQ9NIVL/akA4GaJG4nBPv0vACvP90Usv
eMs2IQeOOe+cMLrMF2X+xsWNWXdKTAl0INolGo3NKwnVHx2yHxiEicZcFPzuQb3041gO57r7lXak
uJy3YvpyMse3RUZF9UKp01czTxt23EE4F4dcy9uU0IbnEL4gvF6ON/NqCCN58Bo8yXkKTAR+o8kJ
bVlpxPl+hd2s8vgG18t9G8eOXI+9NzpufGxj6M4SfmzlqutDS5BoVhF6+zVSiHf6u/FHfHq4MC4Z
Il3xPyRrj81psTthHNEz79kb+evCChUah+YvdqQlpOCOxk2vrAHbMdqc8QQha9dMSJZHSzauVhHv
DCdsEUroF96vC14Sw3u0a1d4OO3I1mTCE/AKwmM8v04GEOFDQ8FGmRnP4aXMqM0bR0foSDiaQdw3
9Jn0OW0Q+RfnZISGThVyR+jyIQCgUzfEe8gACu+SSMWu/9YsBQaSm1rSGQWsneRruVPu/ts0ZYVh
V7j7c7jCJ8682EyprtMIg6iwBNvKt/rxvzbpDpSCuNx4EkTKGMC6YfziA00T8MRJSkJJRcPYUj+w
L0Xm5EWO8/8WC6wt2fAvHWr+w+ACuxRGfDdwCAYZNiGwB19b/mIsfJI4mtM11gZho/kMw6oz6AST
Er1y8CNsicVGDE8jG0n/PUZiLkatIDGdVLqTE9FxmESsveV9dH5/KH1sXEd7YQ4dLcfAqvAMBBl0
r9XEkrd6SXhvlZ5TGcHH+Al0XAb22vOCh0xH4lRdAxma/2B0fmPMchiBcfAgClsgv2SYIJCgRY25
8EJYfzAsXxRnNW5TNQLShjwJ7cWnvDPDH6j0aZqbgKwDkUbk4Fr1RRX0PXPJNY2D3iswHmuYslPH
tL3NEVOFhxCtLgY01wNVcM2BtgsgQdy4SQJ7T2i1lWHWCYauccInavcDBewuOZeT5solb5NST/fB
Q26Lv7UWDBQzNKPsIBFPecntdjUAHDrHv9OyvYn9omHoO7L0/cPksQX54mUWi8/Gexet8GrXKoI5
LkSIjKCT223bSYdTS74tvelH08hg12eMuDrsYbMbToetZ973pwUeIdsWyZPbcuyW4g1xuGmdaGWK
Aips8FOFXB3wcWXSFI7QRJbJFJyTMmiazPeOkRrvMMnbziWr5eSTUjbTT2Vx4AtdLCn891fMf1LG
vLQV46xXXJ4+E768JFDUCqSmd2RassqS2HXSHREZZljyEZzy3mQB0PjcXWEe+1DCrOT4h0HZBpWl
adbaqJpx2q8vixz5kxUSXuUM4NefYEKeEMBiDmNGOhkMmM3ffg551/pTg323iwtD2Sur06eOwRsO
JW+xo7vWSHbDVxHOKl+ncSbZYT+USVoCUB7PvQAKzWgDNDGmh8CLSs+sCodqOItqSjr+JCgJr0OG
QkAx80Laf4IVTNYh1YFHHlqSocdMPxvUIQcgdIHYOjmj8QjZTwufOzrmrAPOCT+OEcp95KGdAEN4
9UX/9OyUIG1JUn4RQVOJpJdkhJfJ8+TXHdXBYul/JSgLPW0G14ZkXeEcPrNi7nNQcCvxYymu3e6j
ZX4sh3Runw669qucLj7NFw6JjZlxUgUTocGGzLIh6wbmzcxobE0ZOHw0h/OoKoiSpBSEjlYG36kh
tpblDHKoMWEfIhuBpyizIfGyqkA0UhbRXjjxd57R+eFV2zjRNAlG10yOUiJez0kuKnh1KNQdzd1i
AO1AeQfLXC2TWZAlpMw4INtJwtfuX8kwtITIbh6nm81tVsHkT/p5/PQYpuIe8tu8GEtgf3zDxVvJ
TcMTCdU0iJfwpTblWew8bOK2+vItmHUOEjzFDsbB2K6xt8BAjWxne9sqQsSlquS7WV3nPC0/ssTB
nJQUGOxUShbxXNNU2PWcEQ+3aGEyu7UtnLUIGgtoFQsBnBiQTSdyFRlSShDCRdflJ5lUlN5PeFbd
yMbf0JacCijQj0t3sWMSDNiw9dMw5LKUbU2YhSF4vMVmUjHhODHEBN3DtwtsdYESu3uypVeTdu/a
8yDenhKe8J+kKwXyfcBxOn+PSrnx6W0HlxcOP1RlRdQY08fV0fRSl++c1IYgXB++AKl73w8oOqXv
W1vxgH8MXuCTdaKcYZtz17h5HytY0xBP4zN74Rwss4aK/dsm1yf5jdHL+frfNsQBn3Wi6uZkFWEW
TEDeVd0m7fKUIdlAGjHykF9XwJVD0tskNPlqXnWNnYntBUl+aJtRTlrffbImKUml9BlQkZtgWCIC
VnZuW/FRp+k650MVyO4BbuKgvf5JFT6vzbpqCX85lF4WQNLpBXRIgSp5BRmM+u8RaJkGJer4N8Pp
ACg53lmN5SSVFjE6cP6DX4I90KH+rR2N4kQZTKN+JVkYh5nzz64kje5VeQe5l2638lffH5Xyyot2
5LIoGoqBTO9NeN0BZl9HXA/RG74YVC9OFjt6TYA91gHRn9ISrHQpvHRp3mRCYyEdxA1GNagsSHBl
Z4RUHMNok9Dd/7cQu4k3WrH9MKyqHffSVgRi8uYdqwJkhYcxdL+KT1I8guT9Qkhln0fyGWs0PBRR
hl7c4t/3qv/jWhQYuKA9HZayU76M8xGcU3ipX728KVr18sy/E3Ikc3eHouRL+9sqdd2j0xmiUVd4
5UnQ2p6QFm5ZMhrvzo0tZY+S/Gr6drZy9UJJc4PcpBnuK4d0hKQrLr7V4OLZ2g+bSSDyfVUvYf4C
y8wpdIc9MIL2+paBTgfM5eyE0QhS0RbKqQk0qqorBRMLz3f3odYx9fTbvhBtuyL7LVXcjgBWLH3O
A3YOZOLlDLI5vNgiIgRPh1/P9XpDHUIcFkebQ6hFVi92lskOJkEmJMCG4Axo3DmwS6Lk5gbiTdVc
eaDNhH4BxajGN3IzlIZKk/UCzvpQCGf6lRq3QmXGO000xH5FWGGQ/ORSXU3mnIgY7fyisrJjpmL5
/uKhbWJKRvpe42zOdJSZl03iknXOoWrtu6EE1kR+WDnZwhC4xm348GV4lSM76edxVER8qv1cN5YS
IZRcO2bw5Aas1j7xN6CNnB1c8R8/BG1x/XAfUAdqbPovviBU3mobwCPzGUXHfPjcvXwt2pNDbqPc
SOz05f4o4UrMNVtx852IRwk6X+j2qSY2pa2kdQa1UhslKJoevsqrleCrLLCiI0oICL7Klzo1hwbU
Ukvo0C6GizWm6DhN6GmyYJI2UW562S1F4MA+0eBxtZ+ApHVlIsXiPldVmjCdBjx8HrHSvVoCypqJ
KkvG/AaMWKoTvMPJ9LGixMw9HcnNHNhuuBLKlUfDiP1AEuHqNpQfmPbN+TorwjVN0+NlI9kCxBts
rw8ulktOXhg8owMLX5/otpNFmyVQF29w/cVkD+ayVQ3ihPQhB3atJHaIYGBKG5r2cjNrTChMGPjK
6cva9u2qIiQQSkWgdjrwFUs9/k2HR3OpeKlmrRIAe2+ynEfvR5GX89V8P87OKC5ZEY/H+ULZVmVL
j9OHTorX90Om9+JJwCj6t0J4WYHv1TiJp+lcr+RYFYn2FKwzAsM3hmvqNsdEuM159K8/sSTor62t
t4kT9mMFcheXzMeoTCfYH+XuED/KPHGTCjmrfaI8k+a4f520Y4OcFFD43w9C25lPwDUHO3MpdQ8c
D2C/8R7+E/w4AyupOBugzJ/WQuhkzA35aBR+F2WBthKLxdqv3Q9eTks+BCVnmr8yc8aSfkX5ChIn
6JPMP91Hol/MLZUolEu46i94r4GHiu3aW2qGDhFd7hRwtGchZCVGuMQbUvomSvQNb0XYvIBKwogO
JaEl2aoObt2YZpO35fnghTf7n04c94wl7I9ZbyC9vp+9zd/dnRyiTeB9yNznJkoQa8PkK63TXagS
MlWIxV+y3vls2bX67kIzTsbtuYFEUa6YPyE0PwuNs1bn04xj5zRuQflwEfs9GXGp6qW5xuLmhZVK
gbCXauQV3q7aYPTv0j2WU46f/riXu1cB3PobLUfyAYhMO/wlWKhJvnHrsZNWWxQ1I8wf6/MSMSEg
fliCgJeFi1X41AW1zc+wF6kHHS+Sb3QiPlfH8W8DhvME6StcIz4qgcSjq0lUa4abCuMVPr+Fmmnq
D+USAlSfaI4MwAZtggF2wBPvkD+diqPaqMDxIkCb5lYUQaj/QvP97AjY3IbKRUTkIAuu6DEjkf2t
6PaPcL16GSZCmNnNLYFvnoHszvgf0l7xJQUix2jtRLKyAdYQfY+miyIrBF2IUK2yDx2bnBh69Rza
87SyLzKI4VD1EXyZ0EGemzBi6vGmqRZ5ZsaJwTZlTjrMfEUWTctdec3De2GEMqp0PezW06YKGTal
WjM0/U+vlYXM0SniiT4j5gvyZ772HWBgQB+Ge6cfq2k6WJM3HK/fsKAeZDKlC0iRuqKA2IgxESHh
rT9z3Niyjbctk4jdl8/GSUrVHeG2MgA/gf7pzyy8WZoBlUnkwdZ1E9Kw8wWfJ4tCrA7TvPBgKTN0
YOAW2kQCcnhkvpBler6mJ0IFScJ3NibBer0SizEWTsKyCi3XgnThNys9pPjuDPKcb/ukFq71BwxS
qsqpTo+1j9CKHQQg50ms9GHaTBHguMPs6l+SoF2hHqLKdLcySOySf0D5fojHZVTdYzNIGVJX7ao2
md3nEobK+2gAB1QcT7eaoKok9bGktZRkvVeG3U4WIsjHMuh4hCMucri3b6l8NlDMfV0BDWN8rucS
aTPNh+IWkY5HHhnKYnM5YZPbif6IsCVPTsfW6r3T2JrY7zYzf81mwlG+HmJFzQ5edlem62gxyKH1
+cwRe/RfsPMFTT6fFY23/tS6n36fzb6XsnYGx2rpXrUw6uowJoRIHmQHOW0P0atGHh5QeJW9w4gw
5wY2idO1MAO9FQ/F2BbpbJe0fnyBu160XBJtjT3rtMKTOQj7U+5VKB2YxZLGPFTLJjgNdzpUwqIJ
2kqfjizEgNIkJqzV23oD4ZpfJJQUf5fLlsFFQwWNCcEKsKgnyjHxvMtRVI2ORhmQ+Tbw7SHCLumN
hO06JUejSvJ7N5XeWWCvgCYAJAc3K7xRw5+3rhzQeSk7/jUSrICoy4glYf7YGH8gris4E9dvTfkE
zfo+Vl1AAPKygPVuhsoU55GLISVGxN18MsBWS3PIMgUD67utxIl9JaK4ji8PcjvzXQTHcGczezOC
DMlJActRiK9e+rfevN6hFQl86AycsTOLvaj5u8fWQIYyzbxzttUAGFnXi9G2TqvRDyn5O8oH4B8V
QpMHolkYbYZwpDeESF7kpeHe0VAo0weQlJECBY2fL74xefCxjuHf/F8k95R7Jys3odcX0f8K1fbk
kEpdEuqqqfJNQzfS3EITDWAqx5+0wJR9BakF3H+FAZ2mVFwkpuxpr5w3FbaUPbgwld/Dx2hj0EM/
6Vs2KguvT5QcDaoK1s6NneYKJ8E2A/VYv3xzARc4nyPa15s4MAkWhlDhCFH93DWufdoHiigFg7vL
prRST/py4QBd0hIaDEhjhNDt+IKU6ZFfa9rg6AytsuRfdc0jbO6nlUds9Ifxcs4XM5JDlbgdGHrD
ZTPAz1j9dmTh+58rqgnhnlgiCtbK/+3FW8cYqv9ZoGqt2CxVxxdWs6OoUx+6O7IM2uXt6gVqb/1+
GoO2byKTtF4FNEwO+XkTjlFIbU7KI17TnRS6/c9E16vmS5lw3nbJH7iGpmu6hm00L27SPaBAN7BP
PlgYFJPmDIT3BGkiHXjlnipHSN+t25A3mfLiOi57IsVNdLM6Us/Ne6mYdspsdT9zX6QiNHH6oRx/
aVIWs5vLwEJpq7u7JRn6zNG7DJN7V7T1pfx8DiXcziqoTakrPOkVSzZBumUiph+/n+QMTms/OHgt
V4LP8H+5TqZ3YXr4iVfx3LY5fbiR7BrmABE+AaeV8Xrhx8F0HbvR48sFhYCANpwkRzn7ZIl04Ayq
+D75jk25w7AMkucX1BnSiRaWEsb6bUDplXyWa7UIjWbTuuLKN8aWC//Mbb7cfcfXFfBT07v33O7h
4n0X/AfPCVP7Zf/0ZCnEyfSYX+Nhc696JJfxlLoKpzzmBGoDnBmQeKdba8L1nuoPuQ696tZr+RfG
B96FZehDbyDYoIe1XrddGklEjSbq//8VsvTgNkTEQzopvLc1bf749BLJYR3xvffjnOZKv0C2h55a
2DRr45xeUckNA1OzRvUzUzaQN6ifNeQCzxD+IBt3MuVLJQ8NMj17ymD8Jneg+kao6QLQKDpYnpRm
nAm6vqjxWtfmSINZCjk9c7FYN3T+V3ltf8HljviPa7tqe5N7HHHbaKHmPli8moQI3DOChF8/3hlO
EKdWt0x2GYAKDO+2qVH6GNnbVfJVqgxdLfOTVb/CRzAOt6IFpYqN/zwARUGT9yzjS4NhrQBLxdPY
nN3H+1gT4BDGs+JPCWMWJWWpPfh2ftyQLf14mDwHTiwXWbIOi36+/Af83Jy2jVj3Mq+v7dRVqQbs
3v04oyOiA3eKg7byugB0AAPE0CTtU/1Q60DZamI2hpDk6jU9qH6BiajJJayO+aH2wzLCp98lknJ3
4oRQ5lQr1Vu1eoOipX3ng5Z6uOEFO0/O2dYTXmdPHKdxyLWXXhmpvul1OEnnY0DkD0xIL0M2A2ZA
xQmTOC59ddhVaa7L4RFNimMvNwrc4rSoUfNf5zauekCQLfjBaouC3ZnISdNqoeEEdzFki2e14NMZ
pUtSM/9nHdnPPgK26ooKqHd0wiJmP6bzulwaLCJh4KQvyd3CxurXUHbyzPB4dQ36NvqnRoKV4eqF
uYqAz60+TXVcm/d9B8S+u5hDJ2UZY1jn0XFeK9VLrwVAs3j+2QRHNC6gD4ZxQlAuoCIDwURkN8DC
86xdiI2AM/a8LLCLx8UA8oi+HRCE2Re6T/W7yENfw9otiWxvT32JUnWMs9n2bJOpFN/SmMuyM6L6
/p9RrIjlPwKnBgSZqM+t5SqTjFA8l4LHKdqx/SPmCYGg9rCQ/E+eaApedW8goTYdSis5novGSdq2
S5f7ew0YuPnrmEEcFio257jvsY1KRJIrGrU+1nY+JkQ3es7m/ZqD9KhBpNjeMmROKcbD6zRi7KAu
3ben1wgWZGl6neVnelg2P4Bi0gj9+EKrAc2kLBXAX0Jcg0a/7qEikk0zMEMqsrL5u/mfipmSsSw7
qhCglGsZW9kWmEPNwGuNnWhAv21Ebd81Dw2LOvMrV/EprXC3fhg7PLmhsqQCEEf8s/G9JiLWL1c1
71cwSXVfmW/vX4QeO5Es+K/ZhEQX9ZspEh4L+n6qsE6pYS3I4VZf1aXRka5ygM/oeGboSpAVbMgi
c/scWMYQo0tGNkGH+aEenHPUbjeQXFkC2qHo74zkN9VX9Fkk08khrimi9m/Z/9pQRb0IqFMt24+T
ZX+kLTeJVZhrCD/QaHNto5kwCBeTcOq1yTpjwDxTkMnQ8vA0a2/w2fLFkvjvaAFbIYTJbMaXza5D
FYxcARR/+SLD7MN/Jmn7BXitP2mubukTOiP9H1hxaVW5g9/Ob5G7EyGi/7VUXIJGHMse0LuJIrux
0NjgrUU4b1v42YQGRiW7/6916gb7v2mKCiEvEB1QQGpoXS9UvH0/0PTCPiL+wLlY9sCK8WBUdtpv
WNwPkTgXb/mDxKeWXNE5ZGR65lZlEp8H2TgUIko35meufRf0xaPKPzl4RLdoikVNhE+9espxBX+p
A+kacNaIBhGsNRQBW2Y54/KcGsqmoiZjEK0TuVEo2JgSBZaHj7k48VFYYTHKRLGLgQSkeWf6SfkL
qFjHwe63KmB9ghtBz6I7Q76w9fxK7liuXRWuVfqpLiqVXmrqe6hnWPVaStFr2dE1XghW7hdAAY6K
wq+FL8ZXlmq/HJk353JiVfDVW9iUDKSVL8z9qTKvvJJ7xxqqiFBg7cWTiCU5sWZzcWDByEFf54Zu
CwDuXbg2cX895m+j/UMXKjsC1T79yOoxaXMhtud0NzSC5fqOmaT8knX4h8+UQ15UstkRMtsELkbJ
V8lNfde5qFksG3dtU0qbRS4H9IFo4hCBv2Qo61i/8ltqlxw5QbuJjtZ4YwfG7slSD4OwXPct4czN
Ht+NcnSygjn5rLoyXI0YpTWJBE/jpsr//Xpj/ZYP++WWBGwZOcSk3hlNR5h5f+LgUzLu+3bMRTh1
lDOBGzw9NADWK75zgpheYBF8Km/4wPs8W/vBIEqv8+ZZR8iFSvHjHiGBHh4aus7Y/h2EvATh4Dst
0ZWJHqWoWYK9yYB133DtzcHXBpeTKiWb5l1mpMUSkur0sKjbA+BrCk6x2ipgn9ABrLBCmi3lHw4U
iMklNbql/mqhjR5ZPs0GZwMygJe9rhtc9F5SUAl7/t/otnFTeuxL8PY43UlVQjFcuHl4Xzokb0FM
2WJ1fsoTp8nBj3ILZOUZFMVRsnyCuPCZKTqHSgaxoHi1WF0QBQ3gvWDyAAw6rWdFFFO8GHbtSFB6
Vs2RCsM65K5Gvnb2cNzep0TkszlhgU0nQrmYFVMbZvYQLuEkPId7fdwc1MBNXYwpQPSUHkLBIRh/
72I3bUnx7/6rh+KrUzPeZnm9G/CcGziyQxC3PZ+5xi/yPwrcSjqkQ5a/wkSoIVMymjbCJ1OYBnii
mUg3HGecin5lO9Lpz9100oTVNT2imvRiycgVcKAAVuXeIsnX4zN83fbhOWkSd33ctrkDwVa1NWxk
G9ronWbiEQp0yJwcvRnfV9wSfItA1QvjihUdRQAEkmE3PxQxx/YChB0Hg/zpxCzFTGqBPVBunDI6
tvnB0yCRq/5llGUS4nR6YSbdt1CUifcpQzAfaq7OP/fW+y205LzZCQu6nlz7YD2z+rRPFP3EZZqs
rpcghteYPZtJZ/WtST4OKRZCVnr86r6Q0n6z1YJYclz65KvkP6K7r79F4fee+3MP1TE65721YA9C
v3ADo/aRrxeeA/eGepiMaQ+6FnlcUqs0oEa79K5lFF48PHqD0nz/vVba3CbOXAyeBxemsDP20zUi
gRiAC/HgP9Qm4y/TWcj6kVbybpRp+pX9wLeuctQ4WHhyLPfTiznOIZy40Ozurl151cDcdaDIkUbq
bsBdphqjArzU6b/MPVCYyhjwVFo8k3TdN6sMKqDWdhFJMqlrIqj2ajs+axksdfmNjei1P7RkL9Sc
eQL3ENi/QY8yVuHmZg/HL0r4BPOu7nwSFLSckIuN5S7LChhkpvwGlFWC6yFdDSfwFCg8FQF1CgTe
uHpZLTiov3qLKIQyJQcTIUHczQ63gnIcYpRDZDl3tv6Y5zwfF0qONE0tV0V7WTwNpjh+Uy678nd/
qj+YqivWu8x0SiWxmLQkQlN37YLKY3lmTqaKBvTraUTGVQNcFmYIklqAhqyQYkbveJ9LixtFUtGj
rCPs1KTi2GoCOb86NJZd2PxdtdiZlNy1H6AfQtbTI7fnNo+/NITZfKeMn7mqw3BeYjPy3H8Z9euX
nuEsxWDCBvZO9i4+yhIGtLFLK9S3UbfQs061Sera4kVdId7OGvs3Xfuh18uWMdN/WHYfTDGlUEp5
d/kKYdcNeGoVt+S6PGoAXZDr5XOJHIw6UibI8oFq8KqOQPQYd+Oidci/bEvkf7+M7/3fAWIziFhZ
33LGKSx0sR2UEb/UwmyT2ERnaXzBwsqeqW6ufXOXL2wHgrdvhLOo8VgbE9QnSqj8q666OzzhgVsR
l/wM56UPu13qAHgz4icPCIjKcJ78VoyGt5GlfAa9Z4DBG43jkyQzi7KiFV4FiaQCTaYzkBDzsfzh
8d41ePlzo90/VbSIAIL01kFhEOFrqPlfaDMC45PutoJamk1XSjH6p6uHvDgzKQeE8fk0OeJUo7I3
aljW6R3iiWm4ix9c9OTbigwr9fUnnmE6FRR3UejvsvxZ/sVBa60u++t3AM1M6+eeQdA3OiAP+ilr
V3UqV1aKFH0neGQpU5/jp3/JdfLdI8aJtEHHLe2NSPR47RUqkckbFF9dU50HZWGRVLpW+/Zk9hFB
/U0SHf+XwJ26jvt6tLIdbdC/ogQAWbPLuDKxJ3ocLeaKektF5jG83QqfZeNFcUL5j5DAnVf6AazS
jpCj0q03Vo3Iz4KAjsDd26NcX85kt79Jgm6g7byesKXb2XVCr8fJS2tO/nmkuPwPPjx5UQu1YVoX
x2pAjRKMxFg2GKXgMgiiosTXrKyIC275cMdp6ELZEwNr7Ln9DA/4UcV0F35/7LzxzEvrKISUW2ze
/wZ0bBoONVvfyna9NlqL+pJtYFTN0dlm1vPWkWoEfdC0LqFMqZpzpBBz+4y1+/xwLZcAR2tYhQKK
0afh2lEuM+8fs5z2cArn5QKX5dwNrrFGtQtvYgb5/KDqWk+hoxmSuCxXUbPW0P3qWbQRKoHXgZVd
yteVAmgzTDZf0Bwn3BifWvsWH5tOkHhMYQE8viNUuMCaBepyNGWr2CR6b4l4q9BLZnoFNEepxLMv
sVny/CA8Bi7Oe4nZbzxxIbq8Pqvlg3YxzvWm3TZaFPMQJ6k6gxYOGYe2Ygo5irn/BWMUbTkDjSQf
9ka7Cm7qz7qbvERGAg5nZgPQ5nORH/NPXUFpnWQokt0wBnF44g/yLAMl0tS2MHVM5UtfNKnP50hG
ubBzl1Nie8sei/WYwcX3x8pP1fJL7yOTjENtWNumycGwsnGQ1oIGW4tzV3BRHNtmGsWneopG8yBk
eh/mmL/cp7LxWOX+PSrNZ08gnPqJb+drUcJqX9K0H2uCNfRTsaS9csvFq/0dhQOHSXZ1R1PZOOoA
pW3WLXp8nTeD/HM6mV9rCa2Z70xeTd4FH+d+Lnwxmt7VfdtfG01N3iYKEuALrS1H40MtJiUpHNI4
k2i5kvbgVDjewk2IFzAFqs/yKiNRpnEp5wDhDFDE3yZKRDJms+NPtVxZU4f0l5CEV+D6gDxk2gaM
r0a9XHqJK9kacjV3pNO3RzmfudDmnQWuX5/68kMYwU3RX0kQeL4q+Z0QoEMeqbHK9UuhIk/YEeRv
14fH6fY34S4E/F9m0p6Aqx93fnaazTpVhGzSyVzN4tIUiUeof0Zv8ZNghbS4wkOT15fp0anLQsO8
m3NDycsRbjtObDbuKm8jiv7Dk9DHxYsVjN5eqdVXyM+uZQwIilClR9JisfQAqO5YNURxoHfc5MBm
VO3gYh0DQDNvyuujTm0dy+hABVwPK3wRX6ccXIVMf/3zhk0aVhsBEsMeUs7IfFWydEtVgUmJ0OnL
2FGAjJsnRZQRhP4zuhyu/AZRBuGvaAvB9UoeSwXC8L99SuIi1In4cj7huUCs0YcWMxKdLPDryKAC
dRGPdWO9DctPVeO4tzHg9wYWXCGW/MAl4nPnsHapaZ9OcG7Jy7kJrlhtXjbyBIDakXgIUqGDO1Iv
cVgUUUNiykgcrFwHtiwj57s5HFMPSKJL4f7iddnxsenSZw2lWK09zwQqKz8ULP3Cab7PXfpmZ/OD
CyOEQU2S8zyK3+VrXZAu7f0wb3GBtr7a0Bqd+6407c4C/HyINMZEgWXWQpVsQRf4dCO+lR1W1ba3
sVKgtanD2WKzcCAz7Foep3rvUm8qdDE5OM6yE4P7FDzjXQR44+JwcF0wFKowtosmwpvE1g6YHTvu
Xnjg/5al/xTGDQbpydBlpstVm7lpKOZXFOopxHJUH9kuSq0p1WJJCJ2C0oh86WmNrxnvdXH9J++/
leh9oXPkbO4W8ewI864HoWJziqIAeuiNlL5enLWoGgy3ysIiTb/6dy+dcNqjHzLQQWSq5o0OvE7G
OM/1ZnTJ0EoXATI/FwnB9skbwu7Ng9xPWd/RzL77bqlMAdVlliRvFVXtmhIkXFyepIBbYeI2Xm6W
VACZe+t2MKlIdd2Es3rB0VMf/3VIjRFbvTMo2pznHIdPZjKRM+AyhWOT/aZSUd52+NQu4mNi4M0P
WC82iRIsH/XHdN/61QfGULQ0ZBqYv5gFzT6Kb+mB84+WXH+poQ0ESuBcsMH1q4nxqpAXvIKjrA3b
C7fvABz49iIogmo3wVtIKZOczbkTTRpiiblU3HJ6VzY9Go5cabtRS+N0RZ5ICmKWjQbryoRDECpe
lzbfteZd/oSqMUB7dN5JYK4PKbwdh64jEM6rg6BLrhleY+yQcatDF2IEeEaZGSluYzLXXag+j7Yx
vkEVUEgUnRZV/ZehUwYx6WQ3RbcxJwmYhftqsvl9Mz00lvG4NeMu4YIqS9KxYZ7sN+9aDWWXOJuX
m/Sy07AEU5HDn+ZWHNaM0G7w1ssEsXiVBbcJt/LblZFnpbX6F245gqBueV1eyfmJOyJDCHmLQTfl
AGGrLXfPzfauNLAayxlMZMwWLk5SeMZXNRJVn0oVXcNcyQ5TP0BIx6Ry14Gkfh/+yZN2WPqbl+ns
pWjFHY5UIOsNqWm7QZpRdg+6z9trC6e6DyeFaRIuSWolHo2IU9Gj3wu3zaJ1yDIBZGnAx2mqohX6
PzOhCsTu9xSnhR5sk4Q5p3UhSJfeYrz1Iv8sDyCbX1ODqGvMJVYjO542RYXVZeT4fjxzC9+phbyc
pU4LonzkB4ruSscive4IDJti+BdhhoEijG+6AQdKPmVYzngCzhizpH/gc0DXvcjDDRvs7UE1cCl5
P1POjfQp3395T2kiOObeCIMFfs0J+Cprv/XLbZtl72q2dNQ+BTRlik6CzG9jAXMr/yNqe6F+JVrK
F5pwM++fTV7mBzKx2vWxRw9hSDhzI2dAeHcnYM1Uq4VEbZKvbJz52fxV5w1DgG7LMEBcW26GCljl
TvAvwqDoVh4sDtRgHY9VXE1/HCVOSZat9DpFk5i8URbOq39CN1yjl2zeBK7Usiwm0ARphRM/XgNg
WEBDgSsZ7M7A56esO2sqFScKoKaKRccXK1WbZmhGAGehwNM2BI3EupNTIPaVi4sRcoGdaScoA7jW
yiFGFn6m937YJklyj/abTNprQ/W7/dfzN4A/gC5QLBieZFIyoDr2/4m+dPJKzvpAHeXzr1OVxKeT
4Lfc47mpRPHpHmI0HItGsOyuUs3pPYiuOs7i50wIAhg6cTq5Q4ufWfFBuKjZrGTYtnPppPA9JhMZ
JMWiJgfVsUOczD0G3+ewIFooKwKddIk+JmnDbuZhg+3UO+qWtCajqBoTxCqH08ddpkbojhSn/3xW
ncDbOuqJxWW18i6A4Bs7ao9FBp9hVeATiywI/c1bCAgwatBLjTtEDIX3ktQM7jU2H+jkt7T9wW4p
Ym0AGjVHg8ovbq7QRYmuyz5BJq82kZvOQXNHqUoCaAldxVFbGxGWS3S1YBn0Y+et9axteSUbwsq2
MOZ42N1BA7aziqAA9hu6dGS375rnLqloh0EN3lizo05qwFPMxA4e7TDn0KvWGySlQwTFre98Atqu
fOGwh5iRGp5mZj7Ex/PirY/AsZMFbBipl1ETgtNsk5u5bWjiXHaQio3e4ReEKdehiwpO8FmvNXwY
VTuKusY3u+HBrjkxIp/EhOuaCcjljnzk9gXLVc26DI+HmV6h4ogOvrYq3sYCOCwkMdWm70oKE3UC
fMDfW7gN+4hQ2raIdXp5K5VQZXfhs99jrzUM07O6fSBxEApzW5MoqRX0YHY6klh/7OJ7Q7xXvtHF
Vwjx+bzRjCigLxGXdPEepPjJrTK0C7fYKaqhaXD4qEBUPzlrVE9XpFTngTFz2vjB7AQJQKhRSGDx
KzJrCopvjyemA4B2jB8lcWHPv54yAUMtoehCbo4fydVlK8iITm1J0kmAPC+P9nx9yWXnOb0sYYbb
kHoChsvhbuMOdiffkqXbq72uu4mTbITfa7/4PNAhnndc+f6hu5jCS53HTVq4DOo+GDDl7aUExYbV
7E6RSMMV3fHYP59lb6VtiHSvIQ7mCBjUPmV7Cl2o3XF0IRTs4o66TEW00YkUuYrPpsxqKhW1SHKj
ovh++Cas7I7BSlTrSna//o3TRqAUMk+XdZ7PZYlTh66tfD8eax6BhCAphUAikmPJ6jA+1Au10Awf
uLIB9iTi/LfMwNJqiEdabHcVXH3JZDiI+/EfDTnuN6Vg3kEIo74GoNAWN7BEyziUeATOmCt+0AJb
cK9WSRAssyUsSqZe+Z0cPSEX9QqPa6AhzNIniK/gVEa3LHL7YNeSkzzHQxyQhmFD+5oLVVTXOlXc
Xa+NKtnCth0AT2+VJOVbYjpmRrKubuAchq+RauL0IooCVYr9aRd+tDsjw5z5Mb5Diu3011zxwtiS
S0R1hN3EImn0uQyBfvGYHLThRXp7Pb3NUJp1e6R6AeXQEjcun34845moVyvI9jO880KHglucMo4r
Rt6lBRTAO4x54fypT3sliDN7ym3v6qQqCur8IddquUa214xgjn+PhdoUNgQnS7MTqCuAag527zEx
nEqao8hPGDHHLJccUq9iWhOPUexbvUCJ9MAOIuFI9MZ9ImDC9/7rrDue9/OoOlmFLpgx5rn6RMiq
jflzrRrbh8iUbw01/CCSy8ddp8rRRyC8oGsNLVG7dIzc3OfLEhhVLvFOq+9bqawMysDC99mDdLWA
vYBs408bJa62KLRBNqoX2PzBYcSHXHu6C0QrX8kuUiD6D12EgKjX17B/gZ1cD6sHcrv2/j0mdhQF
63Mea4SF49fVJk0ibPxKdMpm9YZSv8L1NTs0GuMIDwbsmbWMqtnBgZyxEuEsl+3IyO1iDKoBzQ5V
LWQaFejRbhDBpbC/71l3tGwVAsF8N99YhbYszOIaqMCCW0A8SAyhT/NSvRryyZM73sKa5P21Swml
Gc8fx2u4Y8BfK2Ai64bnU3yS7ZaUqGLR5FSCHTtmx7dL50n0zDkYub4drh8df+9E+KyRGEVmF4B2
kjWljrjSL17W80Be3Bi/UkHOynxwY+wWPWG8li8RL/WRQbQxOvo9b+DvnkZmhSjP8K5SsU1lzecG
SPFdQ3kxLwrrQFAxALvarOYvW9qopDkjhm/0ErRFPAhOJ4NQN7P9+25lLiPgHLTIWv4I1SSzQcpn
rSMkktRXAOJiUSqp2ESIJCXRGhqzrzpQlffr3Af2WnoVIdb/Eca8v/SoNad4VbgM1Ew0QfTir+zO
lPbTy8UaWAfi05u394c9f9+pIDuX1kDIkczFcQlRRlC6a7JK7vQWbx5j1GV+ouzaKBtWf3lVPNav
nsTz1C6ffSGDTJX5PW75YCpJrMMDB+2Xge4juMbhxj+YQkJQdNaTUrW6S3Pxb7d721/Eq5kOJc+R
r1I0eJTV7dCNWGhww+zu+dL+15okkcBCLRJqQoZq6zJ6LRYypBLcj2uY6RD1YemKsdGjwQwJX9IZ
R6YRt/5ulNaxFvGtIYRYI0MrOEmcbb8gIAICIC6+PjXCTyW+yO028o6J7x6aj4XOMD2u6YEm1YVQ
FldX9e80ui1HBHisL7NmWXhrI399wZ9B3byhloMCTuVYGlGeJ/+J6I2uKw++2Q6tjUHFTmxNtwhN
zo58ZnhlU7Mo3jK1F9UPnDMTi9YoG3L6pm+/TxYLZUfshvmBuCGcFodtEbRffXTUpiquOUnx/Onk
+/xh8Xf0RA1MGiQotA9kSn6X8gOa3soTWwwfq/Tpm+TcKCQKqgSvTmSRRdXgk3GiS5WqCEnxFSmK
HYGlMJFHII284noz7NzORFMOs7PMI6HKkUuJKZWSdIybDnwaSOBeQQpUHgqDe5aelX02CTxDWjtL
UKgStP8SkEX+bX7X3WkZxmLdjpAUdPmrEEH8HVZzsLZnhIKfGx/nHeIRRtUdDh1gSdqBnsIE79Bw
rEnjJH9vmkjr9IFxJR7fII/gTiNzJIWX7h3+V/ZSWWMrjVxEYQCgysLKZEz0JnnLDONsTSQa/vXl
9adq477eWIZdRclC6SYgD+5WuSllSNzaqGDTarsAw0V3wHpHg3HSv5Bxqm3Z0b4YzaEQHAqNfe8Q
TlGGsN/EbpKLL/a+rDs91IA1EZ+Z+QvnBq/d4/rLcocI5fAH+dCtiyD9Swa4+F0yq6Iqv9hyfA6G
NHfP/doUitOULgo/Db6+7FdSbaYHzIZtqssM4vP6uF0R5XTL4EFXv202xm7WqvxaoaVzDdoLxfaC
xZRAJxPKM6vBizGajg5NJJ64DdJ/XNZPGj+G1pDby2+tJVrUnUoyXC8drSGdAGWgbqnmVTpN4swS
McJND5DL1jvUIa0tX+1GcDW8kgJGDuaKXWpZytR/o4RwxXVL9pwtZtElG/xLNicSC4qcuQqh/xe1
rq1NCfmyArRu33iqcUiiNZmhHvLHC+WcBvvqtky7nF0Ejl0Fw+QCtMd5PSSDifejT+8zCvt8KwXr
oOhIVnDtCXcJfGxH3dCx3jc9J+CGcrfBSe4CIIqDQkKLck2ttvtW91zNozAwDgzQG49YmpKScC0G
gt8azD0qX89BnLjCzzVhdNGkf8i/4JU+ltYqB8ftiIZS3G5jaMQuMiX8l1nJIQzfPk/JQ7o2fzyB
PIC4c0SmZIVq+DDmRY6dBYt9Qs7CFKhJ5OmDbWkCy7snMXw1xFs3OjZ56ES3OYpvdpXtGo+B0bf5
QzNlYIdVWIGz/BhdxqiPys7uRndRckpm5j7usuBYN4cqxAArXB1Qm/pBxsZCPGin6VLDKSLAxBSl
pGvzbp+Yg9+icccN4SCiYTpwQuPtGQ5kE3nwAI5zquhel7ARq37rjGVsqnAeiwfWgS6b+bZlXHkS
Qop25aQqtYZ1b/MatBu34dWZ9KrwuMb1AR34xLmhTaDDrvM8qDqVtGWadB3KMT3xp4lBUbyNgc+7
lxlumkO70T4jocRA1m7m9Xv2OCja9F4eSFZAqXw9XK+nLFg9w+BNATlJk1V1C4f5T6YEubVy4iKx
do03Kh1gqZdheNr++MlR4zLdkLODdrjPP4hWSdApdMC/JN069q3z8t9jZpEhWInNajuUuWc/uRtm
61HLRc00yHJ3yWhmijWuq+rSPfEjpFep9dvVP5+kGURQy+ItrsBC32cThqeglA+IWQ/Nzy6rN0+z
lJ5MzRQPN9A9iC+q9TVLNGmpWLXXu2qiXujf2GHhDnCRRjPHg+J4KHdtaa3LnFEVZurnkzjg6gbS
LZd9TNMeFbzTc8IWBq9uPwC+GO2qDPZXKSmvuU6lRn+3/TCrvPNDH5+0fP94mEMKRfnW9un0yQsf
GE6cdIPyeX3YLmFdnP+1o8ZusP7IdFTuLBqutYMnqr0Nt36oP3LSBzYRUzvlccio4Z9Doru3vPiy
VZs/4I/j2vwzq9vT+gTESCdfNPf4C8NkcyEEmBKaZT4u3BJA6R/1nKmXaSPvxk9h9NNiBcKd6rva
yjL6hrHVYiYtVGcfw26JaWleNsAFMDl4IoMxElZCBbK3Qm+eqbuSlEsZ0umvY5KZWpBlM/ufFblL
m1bj0mVSw3ptFrXnE4F4dJC6t8mX0/jH7UBejmjjD5BpIo4VvF2iz7MxEqS9MbQ90jx2mTop7+oR
kvk/5BhbOvdLkYM5FzRMUF3CUydj6o5vC4Wy0j0+Ty3bPnSSIP1CRTq6RVoTzEFiIyu05iahvvfq
L11CA3PKhYdOSj7A4stDWfJq8061Kj5CujwmnGLRhpV7DusAuIBwmEYPhFHFEAPMP/FtUWPsGsP4
L9TKldwcYSKLKiem4mPj3Tsbbf4MK+VjYb9l+OwoPOyvqHGOuVUTg+SHqrk9BXWdwJLqoOhE5JQM
aJhL5Qx29W6wu3Bfv0gbBWeGu6Xjo2mF8LF13VTnmIC+AgUskqJycB4GjhQ7qH74Q3JtAQDr0LzD
bDF1PJ8AYL53a57X3mwL0Z0n4UaZd4V6cppHlytclHxXT0kSPbsa/DYPyLVASmop2XtrMpkmxZb2
U/FQS2Q34wOnUkn54GW0nYOvPbWhc7i2Lz/g7Ja3PDvd3ltsmLbFbuEi1it4ezGeaVhMZC3kkcii
h5yYooBnoCZ001VID0vZnJ8B/xDGpYK8WRTQ/1R4U80eGP07JWMcqUmi+9hGkCLEKh/fw2qbA8Pt
ddxb9fY9obh6dMSDCpiGuAG5q8OMUWXboxa1h8XDCqfHsZom7kh5TgJc1VraoRUQnnB2iGGrlCls
qkkJ4izxYctmyIKOrZ1k+/pN7a2WvDEZkV1Gi9o2brKqZptGfuBLGmVDxKyuw/w8EhOuLQFrNLk5
9+Hp6Dp91TCedEy0Q31T3PKzEfoYqW16uYArLUmZ6yPqzHgchj6lY63yE7HUqQp9ssPcSPVaZitj
h4/L7kyNyXbHEsBJpsgN91QFp86tjwqip4KzEasT1IfK7Xl4MrPpNX5yWDBVJp1zOEMldlHnNThb
oNFkTqmxxUN7SI/61n0973+vGIDU+YyAV0DqyFTSKI3qFdlOYMDtLRZU19rP7Ah7toeGCVIMewO9
YDqmB2qSN0y1yhwazAzHqeJxUX12+8084R4STMgmTXs8BSzF8wF7/qULQzDDxmebniOZ9fovQnqn
ciDzJ5Lhle+3qeLABePoI/8F/HV1pSGDhp6Tjd7ZpMWLE9mdq8nw3IvZ0uG+gz6Vh/d7T2CpkESV
fXOd0b03FrojvIBw6lCsL4vg4MfDqujQZjsj2a+zTa1qrBcXAbjnpLpQfrCF3LX5NM30t+wL0zlz
aByd3vyP63O4uAqAzih5kxfun4/P0mQezYgBsG6Pnrkr6A3LMl7iw4YORlIdSuQIYP4NNScdafOz
URxTWBQmMgpk3Qsz3KbiO+GX06YSVM2nDWRau7lZcYlyt/vgsKbYS7Xp8iqPah7Nmq8xeQI0zYiE
HaJu7FAFNMTrNsM2UUWHY+N62MO//6+Dut+Lk5D/C3iSZco2r2iNZ2GXwRUgF/3PEf4iBW7mH886
DX9g58kuia3wsY6u1FKPFpyY4+R8dzSPRl1LMfcqrbLWQqNvGdvMbGjb/fCkKGls9SXcfQKGhzZD
fcUDTaV0qdFCUnkocISKQQdAXCgebVO7a5KvWkWEoAf9RNa8D9t7D1dXeY6QzugCayxXw+gg0yeg
uXvzLqx3ms8UPHikGXFos0aDGKEJwj7HAG/QaYmnZ85fd6c/0G1jtniIxAofnMjhx7qDM1rv4vBR
If8ZUxyM6HQCyDV+oUnCMq7ms+fE9xzlHcPqtUCsTUqWgLFCfXm8XAN16h6h6oZmFHisRFKrmUyU
LESgRq7rqA732KH/rFqNdommSLNC160JwEMmRheuPjGUmb39rMWeaUEddIHPu0gf5w9yqNbnEIyA
10W4ym11JSdZ3mPpcZgmyNK3WE1oT4bgp71Du1gNOLmBV3Tp9liqz8YI7t8a2uvJmE53+KOc/Cp5
PbeO4gt7rb56xAqaKGGvo/PvYKDGwEQlmozddl6tu+oBMFzX0qba2euQA534Ro76e/Y0zCNsOMrk
jU+tSZhTF9LYRGeCb5NOmL6uKrV9TkiVtoi/7EAQPo9+v/iY+0PwfGJxi1Tk5csb1ZnG+Ommpv1e
rGWqCtTS3+bAT09r5bYU49sLIrX/CCvW02aU9f2gX2OyU/N+Lb+bHETR8IddnpgcoHDReLkVYNS3
PICpQBgyX7NMv+jX9knFVLfKwKC6Vu1SZIAa/WZIjXP0DEyoSjRGuFe3xj+l6m79L37UIg9c3TSa
wPTOZEDeRXqjIDRf822GB/q2y4tDn5xLgWGnOujXJ4A2o2wK9XOcBfk67h+t8Osfv4BUHNPBRHrV
BdM6NTjDPUXZlFp1WxzfRzyGUaYEJq5TBTNcCe9Whv2XK84sIl2X84Hnkl/2pXtD/7qVnAUlj2sW
x4NLYXS1OUWHXXJQvXUN/Z9vsYU+Oa0QGq0QHAZCzxeoWc2N4WM01B6Lx3ahRHMrYqyCGV9aanOE
nbYMfkFiCZo8oeC2uxSvq2gtOp3ZtmrSk0JU6C87Kpx7lJsTLIRPAe0C15ktbjDOLOBX53uKkzIn
i4oSUvCnJmfrGfWpsJHN/2sjb1UaQsQuCs+1eQZnjIoQwQCBfKgzDpuiavjUYyv5FTyK3V6Dh9Ej
/QbZeHEplv//dk88Txb7Oh80Y5YqgV9An4CA1zPna4j4O/vAXNtrJ1l9Qw7Xiz0nrsf9Pu9suDp5
8Rpd8TIRpiMDgrudXSeFQpfezSiyLTeTt8FDGzhRX+oz0bfzFaIRVTZ746yjXKV9nWNDhvXIhzwF
3oSnq70WJ4zYjk+uk9GdQ1zLOejTQP02N86HCssd3fKFSzIBMrhYLHBIxy67P3AaiVNSbfbpf/lu
aF90dxMrfaH9eFqgHXxL5dqG28VCRRBX/BkO59cIMFmOqVWiEpbCDB5FuRetLxCBKve+yM13dTYH
D4QkUwPzSbsPxW7TNpfSVbkJZXXl5tGHPCuzpDJ1G5BVN/oYJH+yrK8/AcLrIoen0L/3ECtEtebu
MktkJn2eDrcI2bIT3HGq6c9vM6M4DDdkATCtJa9+9ABJgBHxZU1NjNMawa+5HTFGEwYudTeKoZEC
c9RV6mr4zFXt+eMYG96pIHSuByT4wRQRzhvLiVJyJZbtrsNW3Hpc2Ly25YMNnSSv67WoFtFcFWHj
YyN+zXpSz4jN7N1KwTT6YJZZji069LJW8aJ0+Z8+HLBeEYzFNWs4uwtsqMG2BOtGG756WIqW0nkf
CMByoaU0UMKYrg2HxomSducyG5CCaKXp9DQpeDVaCqcDKxLFEoktOkwDjKS4YwF6m6SSFGRdSCn3
SL+NzJaFugXWnZYuFDTAWvSigJi807ULIgYpCXTpkJTLvPeOZ2IZoNCrJx8Umqi4glPFi2FBb+9Q
NNUIRvfCg1ZZWuKvzKhqqGfNk3HoKb2B6ik2kLQO6lDQQEQJQ02/Rxm0XE8J/b/kILjrfkFaQWaL
fPV/FojonS6rYcD+boZRl1MRMVm42JTXp9Sy804CnIQcn6XHSm3S40GLxKg/TxNpx7A8fr+qYI4t
cAy7qztoEh1YM0AQCT+CFrNh2aYP8gndQscVOIJvyt8G9DVq4v0Gt7NmPcvLHI/rVJCS2kUQ2KIG
+R1wU847BiUK5/j8MYlbkt6/U/R7du82Tk7xXUTKtVnfUzYMse/ONN85vBXbpPe8IARNTSJ0bGGI
+la1k/uNlgB3jg4q5d02Wkit1IQHT0FNHZCB1Oka4SfuJm1uumtRPj6OZIrmfrTx5IZud4tUeLZM
9V4tKf8VwxWja0yA8mhfonbkvMSXze5LF31KQNe3Ee8scFiU6iJsT6BQoA4VGjMWJGldxqVatPff
BgRcpBVsKi1EHrWGvuRtOnMC9gLBdnzOGxIDXVKJYnH7j7RWqTZ892Wp5tjNkk6m4B84K/huxYUB
dvyeJ7+YyTA1/KCQlmE2qiJSpaEGA0nA5lx091a44UhS+UyavsLH2Xs8VbdfwOe+03CP85Kl2VjO
bUQprPk9+/j+1ENtCdJUPovfcGCB5GP3P/bBlh1YLw8jvPIsiG4zB1HN219panxV8oFyDZ28lIOj
xSQIGZG9MgaeO9aaExVAVF0O5tPnSOALeCyGHDBXjbcU5LJvLvj2nt13jrm3INrZI1fH0eb6Zgi6
N99tOpzvdsJ0Rz0YsYW2Bjjeabqz5NLcsW9H96OuLOH9uIs6lOsyCHXPWKt3Kx6pgby66wIhBr1o
ePVSOWCtVT2MJpUytq68D3lfzrnh+0M0YnQJV2TmK8ERVgSCVHFunIz/5lip42RvGsLmjRgXhpUL
NloUiKKpNOjeX+y5CGLE0qBB1a6sRhflAOYeJIDuQRbFIoBRvDHlDqHhxsI0QNpKgvpynzkZ1igF
G5D/v3lxNmGl4mxWGm2N5vBv4745T4aePeuGXPh3QmsO0GZ63ValgKHnMPn31qVzSJNXrTyxEGf0
rv4/udwA/W3tOK4jKOea1t+NM/iIU9h3TKw5RpFqgVJgnS99WhTrB4FOLBM5iCPcVU2pRedRohG5
/6ucJsxE+wv9C8MyQplCvyoQvuJSO1J9d33TysSOIaKobE3cH3VO1yF1Y2D2teXkcAHbH5hKvvlL
ratWgw9Y3Nc7djrYwgMUoy2OlviLfTNbeNiQOOOiMdyaujkOoxPsE+8zjEE1am2onlj/jM7OFf1Q
ZI7ZP4MvrwbI3VtCNsP7PW3UatIb+u/JoZvRuscwMmNLjeSt2Ddu+qlrrGKqqOvDUL1wNFt6qr64
t5q7+TNVvMjWz0OqUeF/Ys6p/8n4xdtq421g0wOwEd3fo/L3DzolgbKGAMAoKzrW0SnDxsH5s/HW
WJejsdOSkCSLpSe/RvfgQrZMZvQ+cWcM6VASrNdrKS1SdLiGc3rmUV6LRh4h3rrd1fjJOhb5i9v5
zTLsGm8GWozrNas28c2dZJUB5dbNWokJENR+TR05eRE0E0lNFGvzAMnRgP4tBtZIRGTS2cMdE3vA
8aLATAwdaNsWL7tL5rOFGxIS5Cw3fvU8luRkkJCi/KwqwdGB4np16A2KT7ThoSZ/KJiPRmIheJSR
KaUp7N2r7U/dIPFroKHc7/sr2PzUOTp+bHXPOrteuvbu8VE78btZhWNE6eXc6kPgrTLVdizAoRSI
OhFOSi6MaRAu4hWkj8MMBsI5nV5y9gd9NHbagwZTrZxGcipuNUZeyGfbyPhn35gi1pQzj37dnko8
z/v9rgoNwxQGHh0LV21amiO1tf9w1rDyq3sG2r6AjXBuFVI6jnzojronjdaVctt4Th2lROYDaPiZ
yO67yrIY5RcvGb1tB8HqdmktCQnMaj0SsKLvPYw55v8lOHXmyD6HaC6lMtyh1ebelOQIPo7c6TPm
YWrd/fuoWe42M4/50RdyraKAcoB1fsQch0yO2fBDEWED9tBBoZRf09NH72xzMwgnIqsF090vNFg8
+JxrRtXxOzqMd/hxhc+gvyybV3nboPDhQlaPsewNHS2d1Y1AFbl2I6QvFgK9T1NKNOieYSRBHG06
pNfiyx4lCaeXeoiaxWa48aQ7bserpvLHQhuXJVZwZd5HKf2Z5jf3ozKVSbndh9vwf/NUtheiDAfQ
lA9R6MioR2Zh+b/ZiIYM1Aqe4lwRIjeBiwEj1FT4SAxMe7NWzBonOEQrNvP/hup8WriAQNsl9t1G
dmkWxJLyqtGNTDnEq6olzZaDizezcS9qfpb/2pAnjt2sOJnel1TXuld5bS0kzvSfcpjHSY4S2i3A
5kzmxbXY8AYo/U0D2S16OEw6VrAeZ8SaGw1wblp+aenvsDvq7KuiAAXs/6rQPW3zo9yQwwBOvg7f
E6JGG9GV7t2GNAmbf8P3A58nI4ancHELbALsxM3bmFKJFCh8MRVvfoa1bdL35QdJkEu4ibZ6rvWb
AiqQ85XM3s+Hoq4IkUMb4aOCvWvYSRW4/ezfo8eDbtiplwsuYg1u+B9VOFuNTXfrvfHlUSBDCZu5
LydAWnIbJ03YrM8GhqOASl9zuEJTvO8PEf1tUaOLpESOxa4LO/tTAhL+YUWPUP5JBJ7kFVbY6s+0
NYKpjCeBB0/lIz50NTPsf2wuxZLYRk31O0GmdfDdm7+K6OoeojexB7zUlWV3bCDROw6byat4pcNh
VglTrs3YmM5ysYbEFHcgMS397eVctNrk5chczIt/xjp3aCrnA2a0B0k8MFKTFvSPXIZGrJR9fDgP
NtEkCLKsJaecph+HF4n59QRLAk1/knJ3M30ppyx1cHnYLY2qa0W7gLuFXZlLrpTKzsHry31+kubS
nNj2Yd4h4yDkHWyVZMDDUHpZu5WN3I99wPnMzW9vzMB74cOhLbpFpMt/FbPQpVW1pyT+7rdzVRI+
0VFml68/dIdiSB9ylpfBrl5fUjyD5dik9HukAaGJrFlq/m3hYvmoDulfk++LbqUQT75dsR1XH3Zx
I5lGqKknD+FUVxGkVxQ1JV6arXXRAfMaLQUNTWWxjh2hgCXwVQDlABMWv9SVq7eEUrc9GhSZxmDQ
ssfVYXjTrzIJ3vYPxS8DuIIzDCFQO/YmDPqKM2f4kJFvACRucdrO0GOBbyuJROXXU6yxC6OMdurB
6VAF4OlbRrHrLSIL96lTeJ7Cxtyw+Ooo/63f4WEj13GUKbWi/vWLnhz2ClPUd8GlyImODTNCRYZA
Yt93xx7MOE7euf0Lg0W5in7yNDGCj/E9/s3FfG3cXZ4pA7OAgqqV1ezcw5vaDIFHtA0k3cjFp9IH
Fx/PZwP420rsFYINQmohk9HVB+BJD3dtcCG9QzXNj13XGw3Ct3o/aJylvOdvrrKq+wHBhZJSeJDe
cdgSf6ncDShFSxue5SgkCLpvdvmqUoAYrE1OIPZmY+i6Jl/KBMzMFPkf66HlXUqRp0rwT4wKcGaA
fn75dEwBCm9BTgEf+gGPRDt+xx/KGaSPdM5qdkd0GzKY5qrxTmuY0LRfQiFdhp9SxJ4sC82H5sel
X6XAVM9CChYeaDsErLihGSsewVLM56KMBpy6xL03WhRf1ODNJgiN92i3HQbNmMjrsjFnC+I5+h7P
TJzFjh12+MFVFIEmUqvVXLl7NpClM5Kij/TV2zsrMMTchVyBukJr4HbvbCLIkaOL5q3W2MGERqhy
xDBtWM0vZlfRpYOikfkVlpoRwtFtrQPs4kX+HOMmxlO14xOH4R9ATj4eCmEvZXbvv6e0uNhYzFaa
p78KpVlJeyPry8I/vHzesV7L0OuO2RMwAlzLYR8wDxRhAt5MucUM0p7v4fcaqHOiFOywszctA1ql
DZDZAIi0SS5kf5hbVdsRVl35rYxryFcR+yHoGV/m2EZCe/pMLOAhFy34QvQN3CF/c8Kq3IgtaeBr
eR6OJ4UtHA1R/RLJ/rS1L/3Sp4TFcuc9C4OM1CHnyELKMwr6TKn3zSbdcgJ28iMMUyJjZlX1bQdo
FZVpo0hkRzEpk1SB87uO2isQoS+dceZctr9brlcslCxwENFtg+s6e3wlj59LG1gpgfOFY65CgSi8
0Gr7G4vy8chEFixe+N0NX5+40l+dlojRFN3DzDVt+Yl8EW/Cn+/DGzchcMFBWb4mjT+3fzMiPKwz
ZuIADWHXmn7BURf8pm08WQz6RFCqR78gc/XN0Zz/zG2B1o0yTjPXbug397fMuh9Ks9dktpOw7JCx
6/++EN2EpqlMeTbB+quwXtlZWxPijudwYswmJDJzxGzUYBXVMCoR/r8exMgpIc1+km1TbZ+UMwSX
BxDTJexzxNx/X7BGXxBTK2j2PtLOh+UFB8hArGsuRMVC6xbYpw/o/t3Odq1GbhXMWEffLCa66mLm
J99E/L5LR2kVDLmWSMlvWuuj62O180PKQrV3zeNI4fySg+JqnaR14q/bCD+O56BWQ22bTRaHs2zK
NPogw+AtR8l4cLjOgA9e7AvmOs45NUwokzkE0U5rvyWGWxSjsKJdHSW6tk9DzS3KurogFtTN7wwC
YOFwgorssA4XHhFNpr8nMXTAHyz01mGO6G962Y9rRktECcEfxUdvG43VQ2C78r2kwvmEA4XjoQ0i
KSfBdqA8ZQlGezwtxgT0ERd3+FDyyQ7n9rXliTcPRcT3/aK7N7OVa53sdYbSS7kIZUDbejBoNSZv
EbDzqTfoMQ9je3Qf8UFKBqdOJmS5feirEyjqfulA7gNFdLPP7yDbwyMXjkDAxLgzRNSKe02s/c+I
5HfswLF91S+Dsgbr0Cf2zzhRD/GZ4YMH6MFDskZKZU9LroQ5hfyA/izG3A/LRR+wUbQye66LpduJ
0HnGou4CMTC29KE1nxmWOVdekXUdP4Ud5ePO/436DhSFSYp/COGoMnYwSUNsJ1qG3HfmNBDSkRmq
/0nQ3sg8mmFgHzRMwGUTt2ZoH3l+KsgdxZZWszmcgPuW9VA6GgDResHuCwxLBj+5o3flX3mrNm5y
4GJ0A7VZJSDOI/61yiduw6BDfeMO7JDq4KZCQD1/xgyr/zTOLLXRrjswLTUJwZUhX3gS+PW1m4rV
4NYPtJWKL5y/1Ghe+UAgew1ZGoKhjsZBfEdK7lxeLu2xq9X7KJw6dhyQT2+PB1DXvk3NtqNnoEZX
B5OSnoFXc9i1xeqlclSa7XDxUNsBXXcd2SJCNnrymyCzoDRwSBr0F915CLxB99ERdpERwj/MF3q3
9yOxISaXtiHVJ0inZkjsZUP6AM3HUfw454PYxDe6tXrkmcaeO4cnOr0ZPh69v3Mn6f0sqsDYergc
6F3onP3bLCYVAGCn+c9Gtgd6L/5qvtljCiu+6U9PDfJCgSTL10SPM8crZO9phoACLAXMCCPjyUcQ
0QqVBBnDKINN87Fgu/Heqi2xSax6dOHyhw00vkKpiXvDk6lNyzwol6caZa9RmAgAFuEFs6oYYG3W
hcUe/wMe/Lxb8SYbYQtpsx/QQ1fjTJzXHl3gJ8FUiDAnWNLQohRBXDCrcAJDQnahompNkiozfm6L
88YlJsK8awUgxizSn/k52IC9xbhe+g3uh+0swmSJ6DHL6aZQ6zFB+atrv14I7WB5DXr0IuL9vsrZ
BveCSvPB/PhprYZlMC6RqtFOwQtUi7EjYbxWp10N7RnZZSUOUJMh3JSY2y+Q5lU3+g6rZwfKR98L
4y2sQdfmirMojBcq2JipX7F8H7vCWOuNJdev/zk+Z1uhxEYHY3OnPagKB/Q8WTCr4UJivCCFD7bN
uvXOiQQrSHSIRX7VHMgu9pDTE6wMjjp6wKIpJTEd/4qNIM6StsuE7J9IYGQbnhfoM4+f38qWsCFE
UQPMZX7d1D5IExDvXm0Du7Ic/87P+468b+UiRMRMpBbjK/6wHKdJndYLzem98+v5orCshZZtoe76
fym1eNpmEow8l+fc+Z8C7yX/CLnn1L0HrI3z/vnbldrQNXpONfRoh9Apsn0V4kOX5DhviHffyJmg
jYOb/p3Ceiv3RDz4vO0i0hoxAK/LH5cE1Vv9LhQEihqfj8ru9EIQNhkAw3evkc2Ba5zitgX4SNGZ
RdE0DIFh7eUh7vb9WH1fO9g2HJoRUioek2gEOUpR4TUtm/gHXbZyw04gsXXE2HnBQyp+v5RAxQDV
Q6lMzaaApLRwMtykJ5cz210xyunwydXgaK0GmVtNt95eylc4i5yyXK+Wjbz4Xtq35sBs3neCSnes
bwEgx43mcD6/FA6zgxAfdxHO+NkZoV7Wdett5HmCjhhjmtxIknRr3s6Wnb4eLUBWjpP4Y+PtUTh/
dS4X2T3U/6LgPb7puofOHDrbDBT+NXsARzprJMJcFwCfsFqNUg71BJhpKuYhGZuneEQOWlQ/Tn20
fCOuPvjnLMRDiUaN3D32J4uY/pSBN0KUoRc4Vt0I1doFEfdMvPtLFVM84Uh65hGf3e1D2EzSUEUb
UvwlYXCpZ/eF+G3shf10JDtX49b8deDgOlGsIeiks7vfZMHPFp+8Vz7aL4D9ttGjssF8n7QRbEk8
FkeNmjau3brkIN3gvKtB7dL6sxoviyp7Kt0/fcxrEOFLLyGUJHWuBil8nSFwVyRrXVhFkToQjCsI
QsD5kPTFwtI56qMSUG+Y2/B3HUIzzsxxe1HA1AL1VTwguTju3zO/gcN6dioIobqUzn2zqOVXVyER
O1HTOKRigxX8stsDpkzUFInlHE0ySzTfsjfGQVFGye32wQYqKEeERDfh/fI1aa3buGxmJfkscuCa
ShUY0nhi4ezcsv6vpdynS5PHfXBGKIlM0K1dDSIQ/i7N1W7wZRL5in/UxwEqZ6WLF4Usvo9XmdG9
xOVQBwLaxrn4NI5BRWFRWdVUY8au0T2OkXNJegygkOUrDVnHz77hWvvgDVA8zlhhEZ4dnm/kHU8x
vpDlhqQE8prfQ9nlSg39U2QKiG3WhfA1uEcJ00tnOiBKg9Q7S7FfQ6fGdYBU38hrtknMewnVfZLF
R7/QiE/ktLznYmMl0qULIjNaUyGSUH+0yf3ph8jmQ/myn4BLNbxHZ8kULQlKKJKCrSJ2NFcQI7l9
aBoJbf6qM7e74gTf90alCcmNgXphbRIgrcaBH4feqvW+VgkI4UXi7j1ZMzp8DKXu6HtfSC5OxWad
oMFwVQTgFifh/xdEtk2Y+h6sBUmSl8hK5p45azY1fSQVTC1a5klijNdunJW/uAT5IXxNUw1hoC3w
TxvSKDXN/5g9LaSBl9Ns0mfQBNCC1D3mQ42m/Yzj/5+peTQV7/+8dclv3SwW94GY3IAQe8SkVOza
k6oCnsfMZ2uFbCyGYck3AMrViLrgV8poCMPKnJXLixnLexVE2I7FRtoPgi/EzKSZej3vZCKXZFBr
isus49Udim/WIjD0YWJugZuBkMDjRvDMXd3nbBaOgeeqVRqd9L4QiHLhBPVNOV+CCraUNwagDI3m
uYqDW7EJv93lHFi2YnyFp1jjCIGR/p1mTAhUbUaF3GvuQLmjFOjLI+g9duLaXepNwpdLRi6YShtV
+m7vLjYcCKY2m7X3G3UyExgLMGmWBvCzUG2B4xnwfyTDNehztHtGGGt+7eto8ADK8knYnob5/fKR
PH8Uom863auG8dMmURU91UHQAz/2ky6ReaKfgwv5czl85qdOgScYsqsrPOGBsleZYJO/Z9OozRgp
NKEy66+SArhMux/4tOu4xs/C3VnmLEkgkgMmpSfyOyP9qyK89KNABe5UywQf1JaoQRQBHL/8JWYS
EzH6k7A7ZmQ1L3KLkwJ6scypKrHOsKyrxJbFwWVKt2mc6xLKGM7dA9+7pyuQHphEpr/TPKzI5KqT
hUV17A9X6klhVvtldhMDQhSc7aA/T+Ukl0cpm1Z0WA5wAgy0xgUGfI3L+JrC6tTgdiRQ5965q0no
DGgIC9ijOyI1GN0TmIqHolbg0NdW2A3r+Ba4EBNo6WcGUgt/dqMUfsl6H26ouul8W0nwfFBKGVMF
nn7Him339PEEtrhm7ilnwLYIomMI3FBFoZqnvJzNWHaeytYiRI97s5pEUVaOvJYE3flMMDsFExrs
KllgnrYrJp5ljMpKPBE5RjZmGhLO7Vv9GuH/F6EHL1Csv4COBiFIT7fTnnzJrB5y4FxbpNxY+XYI
upUktpH0g6yJ3fbpvw46FOZCZ9FHcdTM5scMeDnqjYMWJSvinn1jo5NRooHd44YsCQ5rcWnaDWcF
QsV/L6d+fL/eh8uNgLXpmDnXwIexo3lch4/3klnwD13n2oQyxB4jC3p6mwpxteVw45GKNk93CZc1
+e3CDlGHjg4OIekUlF68VuMXysGlViNU//4ki6J7EKpEtnQXwb3G+6aD0Bag3x/a8KVtXMW2lNnM
B931Yzy/Y6abISLq4RkSbC075GtXUzDY9kS74F/DUMW3AS4QhLGLesUsPS48JL6WIXCdKEU/6H9L
tJTiMHnEnSsSXoTIkxjowXrsy+PskRjxelKEfb4SXUvUU9nKNYmzMIEDLpu61v+aDs3GbljShUkz
/QokK4GH0oZ05EtB0HJ8D9zzrvwKJBv1g75nTjKwu/hkAYA0DdJqevBEryVMMw2TW55g13TWr581
f3q/ZVjga7K4/MAhOCYA+4BvAfuLC+/197BQt+LtXyDogUIRJnvWeS14KjdYfgVMUDHEY2Oj5XWK
ekAV0olyNSCOF4OksiHOwIHM4O3mGMl3Y0MptNM+7jBENqmRVybNKfxtpHkcAFQR2EWI7EaHPZAS
Ipn2J4sjiLkgGPq4W+yhy1SXvDZ+g60VsReiUgLcFxCJjZVnndXB/i6ydVSCCg8cc/LBl+6ELpg8
PtbRrNKCnVivvm+KKxExJYjIu5GPF31X/HLfDTKSlzCN/9htK9B6fN5KTXoGh5EqOuBZXRDI8Gg1
8AhxKcai0QsLfUROU+ipNMCP0UwrdiEQhSqwQQ9oA5QzoLryUSvTrR/Is6rYuUT3gH8aVrSiw5L5
AURVRqPWqx9j1oniQgeDUJU1Qeqs5bbAwO9TBVfvh7bWYt91FfHkH90CbVwWMM6P665J8ILgA2HV
ohV49lgu4QnI6Je49XsBnNxSImGYZOVZTlXXoIZAzEdClMO+DNPdKrQsz0aJmBAOiniGZ1wTSIFB
wgnGywhQip9d9c2BhMm5MPI/KVBqOkMqduX3/kzeXUKdN1GjuLPMHQwztLTgqW6LLHWINu3Fh1Bv
uD3p7hTwuJmtyY2z3/GnaLfP7D3/jH9TeJmKlD+OytRAq85HFpoIEsKaANtIQzfT3wdtpVV/rYH8
d4zuiGCyQZ+JOuWuq43F9neA9GqJkbpvj1YtHJ/7kP1tb7C7VclqmqVLBL5TAg15FPEM2PPMW1aF
QdIS0miERnhiytwEs/3nmQGf6+JWpO3M/MhCxa4UbJU2yCHEv4fY4Km48FXYgs7FncKCjCKfc0u2
w/qYqvBsrVVInJfyrThPADnSo8CneeJbdgao+7mlOIWIoQuNpm8CStXEBKvieVhlK066KOIrbUwN
Kbop95tLW8fldLC7F1z7G8No5R3I1QSNt5FwObU4TkyYid/XrucqdUmf/T55qDwHWmyINj/A8Pj3
JzZFBokdV0wzkeJAYMktQTlILMc7qvBwz6WIb4YzY6VllEIobIkfljhSez7spRt/YPhiVvGYSdpA
uMil4UdEZeOgCQvzs3bR1jx71ePjuj4jg0YyUOUwUjP6xpWLXUVXr1S6Nrikb7GzC+4yv2axLcnS
KZ3iYRYPi/5pTYBrjCHWWwtwyJFC0efSKitzkmdNXvkoW7DfHN+jSk/4roPiaqbHv/wkRYGaUYGO
0l742VqWZWRwh1Syo+RIb0/Z0Jq+iRoxK4I6zPlaplMLdMzaZWSbTdZQrgAmj7QqxTXuJAbTRyzp
nD0xDhKg4GSLEs0nlE+9o4vEGYZNQrQ1iCXQM5w6uaGPGlzegADJWCYbvHs5JEVYnZvQgUX5jXLd
EdGrEbpinhiE5PdFd4/Nb7w0ChorkvPOlugvOv2O9zfBCoVczvL9Exmjqn8aoFyAdG+v9hH5nJmi
UlJ5VRcdC1SjjrLM8E1RJja2ggOmciomejo6ILMPPtWnf2tdMcQYqx1LY04shfxmtjYpf+/TUEBV
2UYUPKXOqmzPjserNXq8M0WpjOF6XB3M5JLIw49Vd8oEBC4rSAPe3cSP9MhrECyfhvO0JvZKJ4z3
utYjR+W5VkBR7pg5eR1tAjpL3oY7mKj3kIWAkuUmCGE5bFqgfWTkOddqqXD80vR4OgYd3EcTS0AK
IX21+1PancMm0CxARo4gJTWsYDVSRBhDCQplYhR6uIWaF+F+6sMqMvoYHjhCnH6RRgUQW2qdTzcr
BXGyyU1MfkKHVgX4uXxMnoigHitQdgQh09bULeHpkJUNyz0r/8Zon7BSZYHExRQ0Wdruak9Xd2pl
pG6wgSjBIuahfXQ16E3IYBGs0nvXx9zCgz9TCZnMMgYdTEjcZXBeHt+K4wVIVPkvzMEqo/prxnM9
Jgki4Tes6UVz1qLYy2PCiLGU6RXTBTnZY3owd2IyTwqyolAM8+gOChyVw8I4XBT0ouiKtbLl2dMv
Bya6+MO2rRyfGtSwYubQX6TR9E9B0nMyw281x2vKu9t2gjvuYnst4uK+OwDHAUxmEcbZnPL1/g6W
nQCeZBO3foWwMw+dlstp0oCHMww+GbiQMke8Se/RkOeDpILuobD6v+4C4Z5Iatvx5/ReWa2ga8wS
xmcnUesJT25xtT2vEUQhLhS6yCmBc1rbUpQ5tlleg2iEP1hesd5vZ3CQMKwpenuMHv2RZ+jnTugD
1xhrooWbRppo7dm0HgcL8TBQ1pfJm0t9BqHaX8ON8VX9HCIabOyVVzrTWt2afD7NIJEAW3eGKhXt
JvPBX9YYm7ExZJKblncNHbdeslJvVL8LIg3eavHA+t5/EeYUxIu+WgQaLMHuN1/Cq0jFzfSdT8mk
Tzt6BhRPzGQrsqIw0OlHm8BSbckmdvsMpIPtuRUTzgwOE7JsZ1E59RCqXaeOA/LMiDhXLBmolGLE
AsIWml9ucsK6H/BpVuiUA3Z+VC+DuJtJnDbyyOLLmm0hmBEyo6BD7Da10UYbrNxOwaS0vS+WsniP
5cfqVE+Bk3MT4+CKhPb4ZmsHhYKqut757vqnUzK4Ix7r2EU6P4Nl33LqeKZqZ7ph0kyCsADHiK8o
eLDTcG1thT97UrSZKrUvv2JszEzUYM2aJYV2jaDZxuc5VCZa79tk1dULfkis17uiJrUwG6rCVZsW
JJKRSHA6f48WFOyJ3LuDy1QV2ZIxWEDaggwmY9Ad2LDBwTENIHMtkEqJ8BhlWyPr4jhw2itzLCrK
MokEmEr4Xq87xne/U/vtklnntwOMfzTgt6hgCfR1Tx9OBe81jeK88yaDeQQiwIP+EwybbTzGDQ2x
fnxQvhnudxjqTbLIij3YiZJgc0cOiKHcQ0oQUWuWM02Ydmp0ScEHhZlIFvVzSiqiksAmOGsalhao
auta7icMUxdVejNgeUlViXcYLjpQ6ms29ga8RK5WUnsedYoNja2er6IewNONn56zo0XQsfmENz+S
omCW99V9PJDax2cJMe5DQke4wa15j61YpuA3kYB/cgZ/Mu+Zcmd3A3a7TZ+8YnWKGV6m/p86ZTKz
ao3AnHccnBW0MFWUHhMs5UlCkHymOj8rHyNP7DbvLG88U0Peck4pXlr6NqtNN+93t8D8O1TG4B+Y
RShph2YtA9R9bXMMRuKiUcsYSVLUexlcD3EfB95htHGB7SPVoF1jd4HY14aBUl589rC8PiHEU+Gm
x8hCl5zTQSKc23AolJa3TommnBbUazhb7QfQAG1dMl0DnNjs3mjgNQeP89SzlCMPvW2SRki9jyHm
D35q3lhhT2iuWGxxTGpJCok1PGHdbTfBwictdhktx4QnCtBmsZPw8WUeC3BGvwff5NofRTra61Nw
sesvjaBCr3Ve8dqhuUPQUeN0CDCCfz3qieKcnqSGuhLwDN+qpktPKspx+6y5Utuq9IICZ5L4CBVe
yD3OWQAC0C9PnUXxrevxUZdUojzl20o+JuBIYJ4gO3/29pirTpczdHzHImPa9HN/pqDgxNE+SSvo
QW6bGn58AcKbf0zoDFlvlWIFNrs/M1QoONHjdqsuJMHhNzxvj/c0AFTydAhcRpj6XMVfVP0RdIdS
Q5gyIN7jtI0W84GZj033LSMsXTnAg7kwFCMkWAYa62TjoO3LK8/95Aw0Qnl7trWJfXoWU3isEP0T
/g6V+FX26SN5IL2mKB/QZos2ONJbtyjNsKOiQYWpjKr3OvCXkWIXuSNxsnNHWKsGXRSbIpjENqlh
Va4yikIP1JCOJhslb8syHKuSlBAMPBQg8Ce11Ub4ISQTpjEQJHc10O+fZmHu9ne+eBFwF3fRbbcS
XIIsy+2TWQmkHeTCCIuVR7nte1p+Fk62eNspcipoheIelvx2OjiC+t4DlltT3M31oRyo43RdXh6J
7W2jLClBK4jOuhdcbWllWMZbeyWAGlAHRAJL+hoHF09t1vaGosnhyx2cjSCqRYTk3bvNM2PRFf+W
vuSMDgH2Bm6iATdX6KJ203kDfdsFceUyQ8M0oF0eKZpDw6qq25tnfU+OdYb0r9AqAYK2V37YLCy7
JjrTB4AJU/YRA1j3tuq/NTUNh+hotrpfZCp6pUWlzs0nv1Sn5g+ALVs1inZnzxOiuEzepZdILiTQ
3DPdJ4INsyvs3kHWNoGqT/50o/8tu2+Z/t6t/6bFkF/HtbJ6IK/n7DCQ6jXSRWzASAR2jI60Q9WJ
25Z46atgrVufhATf6m+zHb9mj/SQN2kqH7zrVQjAJHfGESOUcf59mcPVlaoQfLXKrlmlGkAi0oKW
9f/1vylxuDGydSpNsAijlxyS7oUEv/qgrHxDtqfkmOa8IYuDfmK01KUncdlgYHXcq1t5wLJpf55W
gvdFr/iMyrWvUT1T9s0cxyeQciRNJKQc+wTApVdZ/LqQgjmwjx2d8aEx8VSFFUYBmG5/yYZKVXt+
i86gdMIVh7m4pNpHe2pVtzNsK9dhj2pcQHLAG0K1hS+CshnvupwsbETa4vaYHCoOL0YxJIL1UvQW
JaLz2ehc70MdIGNbKttL3vaAytSbt4rkrJgLAgIi6+oZeSqJL9JlI5W7vXOtnQuUAjASGDlviSGt
Z08rtv2fEiwx3SslxLK0muxR4Zvjq5nYUxqCUvAnZsHRvTc13mecQWd5MDVD4j6sxPtqELF5wrQa
sIMvxiQ9RlewK7IhfrNN7GiShHPayp9q29qac/kXI+rhW4G7w4en/LRyz9c+HMCSZga9GV76/IEb
ajMxC311S/vJO1SBgac/pTzjPWsIPoOzXBu9tX8zuf0Ynt7vn4yPaEAv8hsdOM/Diegv4PCKzVFZ
/KsFI4zXo86PzN2npO1ZrG/cAbzdKx/+07Wbcv41+RL1/v4N1Y6hlCkugf+FEYAvgFUDhUGr3mDP
BO79WFNxV4QqX4inoae21u5dtebDPBapGHGljencZdjG5ffFTERzHPPvVxaw2p5gcaeMNk6gb2/F
JEmGJR/J+vwhgjdbk8J1ItJxSlJ0a55APD7Ur5k1zC7dBDcLto4xeoqACP3nWttYO1524EFNNVXv
CmS8Oxv91ry9Td3TgB4FsO9IEVA5hy0Wx9fNF+VC6JyEyB8TBBEqeHSvKgN2GsQ7EyMI9fv/wPu7
pV4TeWF7IfV4+60Eec2/08kaR5cw0bbBT8TAom7KPboPeK6B77t++to7bYWfrtrwUjUnXDDVBMp9
1Joa1o763cwgSiXKqLMNgDJ1e3wsUxuktOtXG3Nm978Wb59afGpuAOka496dyNxGnAeWE7NAFc+D
4eth35wAX4GlCqAIVE0MO52VhPHmeS8zntpWiiqFIEDjDaffJulrykMcn9rU11XXCSS6Hsgvc9Fk
GpHOYu3/IzpETTjY2h0OtPR/xWjRBToD/dwjxP5N8j/no7jGUZhYcESW9DvLyxE7N/KwmWB7jHvQ
LV3IwNdYwiapnvYVQT0Oq56C2HhQRV154X93Y5Ov4zjsL7UZLkO9ZoxGlkTBzWRUEVpZiOVGSXts
Jek+LTlniID1z4gtko28vM71Yee45Z9UmeaJVaoLFMdeA42+vhSRF+tGSHlKx6I+IvbwQZyLH6TB
aI/3/Um28mkzI1n5G0YF/kzDDkJjYzwRZA8kY9Sixr3elVkN1HMyLJgeGcCcItzj49EbNwF+eZ+w
DKrpH5jiYUHTvS/fJpLDDOxfuEFyTS6jGw76sj+TQCdm1RGihdter+S8rotNgSNDa5RnGo4aYaF4
IeCGgFEVEHb9/BR4763fakrESQsxKPEI4Yr8b1XqMiX3eacFu26ff8ro1aVC6W9j5TNFTlVJ9JcX
fjArkfiBT9tDAnUwxVGZOh59nd5eP4AgZWHUIEYx2rIuyVuwDxJm1nzkFCtHRsoAj9PBihbke8Fm
AsFfgcTTf4USS20IK1QKJBfxYxw+62xQk1w52fyNc/5ZSNGhadAz5tQCWXpdez6skHUfwnVmJjZJ
v08wCApPw2qM//k+2kC/b3Y0UTdEiy7/CL50LGHwZWxsp2zqrSphzqA8ihMBSjENxFwQaB6RrUww
eNpY4lp91CCqIQsC2G8/LAbiedv0QmIcM5SLgp/AgzhUBJW4QBM1rSDQ/vpAGZVt5GglqXvyrYML
6QzJHEOee+VJ0LcdNQFyvhSi7krTTnH0BYyWYU6i0l9LiAeShv5Hqt5LfTJzBfcjx4vbY8GclySm
g0Wb6bLGtKqLpo8CsBZBpwe7bMbGI7DloqdDqXoleKsRhpB6D1o7lXfojP/oXrs6ThbSx0dwjDpn
yd6v02DWQlK3BPLUHEW/M38tnfz5HBj5Z6tBgwCcdB1Cr+B5JPzM2Gsb+AQm8ydu1q7FOT0gqT0l
kLiA9GUEJOh41cq1RKmIUniyovOE++M9H3qV2s28iLSWM+lsy8ziA7DyAlzzKJJQY2XjqzoLbUZc
s3IQHDN6H4MfN3+CwDGQY3gLJf0Wl+yEhiIGKvwTlSxjMxHrtOEqiD7NG6eCEhtWA3JrdqYJ5D6/
2KUZWPJ1+wotvWA9NGNifozTTiUbVcaPW1dvo73Btpv11MMlCeG2SrTZXpr7eWp0hDKsxZB84pJl
3bsFqoY9ECbG4Xei5XTa3Gmr8lWnDfr+80oyKmLq+9jbK6FuiOIFfwy8Buv+cSaFRVjmMa0CUg5J
bEuDbPJmwkWcIwHQLeYXHg4VssR18Q5W6sRv7/4AipRQi4xLFN9W7Oes2PB4d3o445Rn3wSgkQK3
RoBtJJrSdOiw+xNdbR536OYgGaL43jTn7CKwYUFdxUWNqnhy/cuw78s7OLmm/1pjC+nDS/Blagz0
Kb73bQH7qKNycEF1dEthGruJGKW2ut95SH8DMOw+pk3Cdb+fSs2lvMd7OzzwwLma57MNQQjylAUC
D+4LEYH4PeKcK4QvolKkizittbWa3kmnLPk7IYrEBx9/VZak6CU06hdtIWA8e3ZItjC+UfhMn6mj
SZ6XvGO0fcOcX+8QDRE4THQ/lDNkI6MpxMw2u7O4VkQDTh5b28qDstJXi4CUBCeoj8bfEgOPRral
GG8M1bA3ftkPRLTt9YBhMS3l0xu2kAfbvieFqRHWktaTRq4maj3nE/BPglmTTZsRtEpPZ4+rGzGF
Pmp2GYtpzw7aDTwLeVNWfJuF5v7tFojmH/qyYkMF4zJY1MzsIl5lL+RkaRayKx6wIYAGOXNJvDZk
7oufEawDAXwUXSesliQlMSqZ+d3nvIS5+umxTiGN5+zJFjJHiFA2mboLMZ8jHTio2J+BkrC3O39d
fjjkLvzWETcAN42xOq9HzMpCih+jfH+5o8Vpn+yT8uFf4go8zb/BBqAm31ScdeHjeCsUVrKDG03K
V7dVOVW+/lAAetnhD5yJfNKTJb9g+f7ErZhe5PLCiP2jVFlobvNPJOPvFAyTDHWMqPR4ZMSnJ47l
7Lv1VJNY8XQ5JqwIqnTMTA2HOEjGY8iBisDtLY30a3AglA2S6wZn0GweExHmGStmPbt9pfaKanDW
77xL9/E47hYucsdPL0uVpgpFZ08lGeWqHiuzJIro2YmiCGtdArQvaSaVIvryivgOw7fTdBxAKX+X
go6B+Cmo6wjUCXg9eeYiOgkrH8HGYOdJmGDyoTzZWipXXJ3thXRLCnAvqPwVTO1/3gOPb+xPb8mn
19iVpFb3ZUyem+p0gLgfyyh23STpgM3JCr2Pa6ZCXGCxP/6UsJzYadf/x7q/MOEIVl48yJnlxB4Z
X6dzEcGDdDlFxS64+OuWzyEFvRNWD5fXSBLx82YloD6BtLO1FOM/tdj8Vmej+orVnXS+M9I1GfyC
f7oaKscfH2r7WDRy4KuVtkcePyNwDAJm1uFoV2JFVuLc3sNEzJDoi6225lPFg7IJFXDAmajGufA5
lfWnKbuJcINWWBrNUb05cLgKSfQkmwbZZWgrdduvB7cLHo95tmcc4cb79/g6qmEmBab5W8pCn5Pc
b6ZS0reMzvOd5L6kYFM+mGXXZmeVNpzz+U383Jv70PVHYunPSJsC3JzERkWkQI14ImVIzGhHzMH5
LPoKg9t2MRt+2NobocJXDe7uPkRP9c63/OSOYhImIRXtVJ3EM7dOI5qpy3HmJDvrblr9Hevs1if8
ni4oJwUCGeYiAKku2JD8MkIO4tzc9ml4/T0rVZk7uYpnneBV2rp2kb9wEQNb9LsDSPPB+WMw8W+V
gqVlBQuD4bundtvzS3dL/cW0XR1hwiC5qnrbE3F+60gC7PiSvpKYKCTBoKfesPllkYQNoGxybh1A
+Xx+i2fYhzvOAUzn+oFIg++zJG659OVkTX1JhfwY4chpEsTY4O0je8x9qK0yGrR0dhsuwxTOpx7f
b46OlWIr8P1794H0OfcdnzTsjgsA3I4TuQXBaBVIaTOo3bQFHHl0vfB5HJ9SNcnRh/6zfWED28ok
Njm8WPdTnNEFr7BBxcCSLJ8hf7Q6OOGrwKX1eBGp+5atvxC5OYx/TObqDzhVSUFPUPo9BJZSN6as
WYsBBmNEVkRCdLwnYq5vxowbLxBzKnjjDDyNyLKTXv5OlNtDR6PBNnHMAEGG4M9RZomoNrjOVrUs
EAQk9d1H7Fv+UC3ntbHBc1t6SaeuMwTowNDKfzGW/vuccuTc4BU9aIX/JIZVFe2iR4PZ41OMxNE4
lmi7016SPxO33nqKOkX3QXkpUXsroW1e1XTgc++t6rb7XiilL4m8T9FzH2DWEGIjKn8qvoXXwWwH
UTDOkAjBk9WcrnPod1BVwBdgHXq5b+uENBoU9vfDYghfmFIWW/l1yemW+I5jXZBKIXiMB/+os+vW
3BM0Mimip28SofIPa3kC1TOh8U4ftLmEdahz8xxn/lK0guEAgb4dWyKANSl+utNbWy6LcjmXCjcp
8PxVtGS3fuO/ogXhtd/F0KjHezLkdplBIdejzcWMTSucOOKdr3P6f5EQ7q4eK2kEVgetTbrsb/wq
jsQfYGti1AQGOKuUi6Xrn0MXnC27f533Osi7ZrHV61tUAGo6aqsDa47YHUN7HWlBvKJxVgcuRDYX
3L3AnVYdVgOYgfBZg5i0c1nDwxti6FoMf5LhDHF+tj3TddzpLgirmR7hYXYGHTgja7M3e+ZpvPNi
owuGYbTW5uw6i+Gz35coWsNnDjKYBV0o8fk9d6U0McPb3eIsBScCkj5weWAd2SnFp6kl/hm/+QQ3
45mMwqdWnbuRYrwtKYhAuPbS996W0hipcsH+6c5QOAl2Ggu+N96dRNvRrCPKbo0zPqvWuaqkZraS
n/dvc9dFK2cSYBBGlHcVYsa/3SHK+iz4MZABG7P5ZameQqVztWQX+fWiPYpHyWYKCX0/oXm7GWiO
fxaaogEuWi9EnCyVncQZTA8VFU2V+9GfDtD2VNEPwebpkcEbsAURh529hk06usxIF/QHuJJMPUn2
0wuZ/0roZjCgQ5yks7QBbcRhHUnmMma8RzdpN+w67DD7Y5u3KqoC8yt8B2SgU9bmqsFwYQFOjdob
ZHB0h3UKPxoB24XNdOrbMlAZAL1I/Z/qz91N7vtgbLDhhTFrcFkoyMHk3XVK4aeoPqPgu1RnBkMC
vEBwp+h7aGJqURK1ZD+1SRR8IvVUpRT6SXpyAzTwMJjZbxNHxptS+kzOu/uoUig6X9v4dskR2x9e
se32LvMq9e2P7/h9ng61Jv0Qq12lbUYtyQF54g7q2LgGHalofT7cUnHatDxskArh/9saIzVN3vrv
6WdaHvSpmjlXgDu/HxvxN/OmI4RfVHuk6lg9gx6/iMbFk1cMedi7PnY8t6MxZTz6mU0oiE22dZJx
5Wa9GhdXGxjnFAZCO/pGjUg6KvJat9kKovOKiX8rCNHPhRg56wGQX9x4ea/P4kF1zHhCwpF7U6C5
4N/eAd3wuqfkGKiJOTR2bMMIt7CcqGFKEgmAjkpwL9EwbXppHJ/Yu/c1YJZHUHkITuHMFGIib2+8
/fH/PVXI16Hoc200Ja71TeIAZo2RMmF7dOlQ5oEISol0+N6mTZue1TyM2BjRkJGV8IlzGUkLLLlY
joe17zTXMbwlfncEstVGuZEoEx8wkSFMsfdFqFCB2rHww9r5ROL3FyPakpiVznLSx3D3LVvYJBbk
0KO+jLTrr5cejymQEFImoNkPQGuFyJ6ejPg1Wg4WDexsV7Ehkk+o4XJuRC86Tz4dAwRU9XrrRqDU
ZHGZr7B9xbTYuGf1sRqAbKMrKxewmARh5e00PIFHvApFFEFAJfM7MNWJz/FmCc/ydmSwXboLsS1/
+dqHNZmyA+qCk5uiIs4x3A/mV94/JExV68JiX/FELw3bPX4FKCw6Vew0xCpbqtQjQdtwRBbbHNxL
JmC4D93ActBia29L2rBaA1Dp7hVrS/UQHAY0X/mToiMBmUxupAn9BphV6O1XK8yXC/usv905zL9q
+onOMJRXG/uZXIa9EmvV+s69oWZrQtstPGXFzh2w87CFHGKG2RPVxcAGOxOM2/lDZzpx9PQK4ep9
pqUXiI8olMQfLbvFxUMQ69V4dIbKYBvuf90PQssx5rCVo18m1t68OFOILykYXC4YQxaxr+FJe4+J
6N/taX5WMn6GSbdKrjX6m1/wNg5WAxm2XO/M13sxqZpyUsPzpRwKbdz+gzFTQYdo2ACqNV4w4v46
qc4zg8498wIVYVoxSXoUDkbN0AIMZOQzgcuG+BrkV98OPoO1wgrj4/PnOUG9Ssc93EOeLU5VTwtb
h63DizKTHeKaL94JmlM6k7KDomuy/9RUy1nPmNiV+yaUhEWaQvAVXtXEtPwCZXqYpaVsUiH1yFKW
8gCx11lmv6saKlN7+NK7yYplPsZaYOlaUQii5aaFstCTS877yM5yvaZgyaUpmNHQH5emtf36GGiU
b4Xb5M03NP+BNK028Ad383P5C9Av4+Cl7mzp17Y6wt4rsppWr14RUoVxIgZQqCijy776U9RXrcH1
AGoRWVa+TY4548AGo+eFDRmGW7bDiT94motlGtUz0/7SKn4dp7BGLE7JF49McMKcJ/5QfG2TAYq2
ONFVAkOUPyIHTF0CkjLez7HsHWysRFtEK+TEvlR9HHrMCMN496hVe3fgz0gp7Cy9O+esArxLLila
mC/bcq3irFefnARgzIFeEdaAF2rGOuEMe0Q8tTR75Po2UfSLMUV5XR+oQsbH9uZ0rkZmBTLkOVv/
JpzaKTMom6zHd1eOzPgH0fEjP5Nd8LRW7zKsYdKLa3mh7G06kZrkqPMpeTY9AWB06QqXPSscu9xz
vPpRpKgYj9BXkQAsNBGoib3zkl/PwnNfRddlTGecOZxcoePkZUim23bLiwa1morvKwm7MjH6HKUM
F2CwyORe48smW/xp3j6HisDeA2VIugzU+HGPfz9RO+To6HCy6/iqvTFd7lUZfp5eGmT00nwtvNYP
ROUm65YBs4734HmkrwsUzbbqV3v+PAX1NSDJUrFxuBZTE+u50jr499DP6loT9A0cgTaPKBdF3Iw8
fcVGUaJCVxES9CtKP3UlR061cprkf0A7SIZieDgoBhDvgF/wJ1YNXLK/zLVyduuXOTUh09Ybq2G/
n2ZpjtuWZ+P9SLz/Tv515pfhS4G0PGIAoLEU1xNC5/hTrmty89TXUfMA3+vX91UtVsRBSovXV0F6
OmxQPVFtZ74lffa59mW8opudUUuX2fPbyIEgR4ybURyYbFl5X4jUqDcU4hasH0AFj64eQXlo8EMv
U+CBzArm6eExH1jxDiDHgLlguro3mC82FeaZt2d/ixVlI2bvZnTZc0xQS+mbosDvEpxe6NwWPQ6a
L1rSxODKDT19bNKN94+tl6uwKK927Y9hngCWehWq4L0HxgzjBIUkhdx7c+54lUmq4RWQ2cIgFVrL
U3MIjkPzXxS45X1Q98VIIZeBY2ZYTLZe+pHwxbWkFzs3zqwBaH/EUrxINGirWndbw38L1S+LFRdE
fY8TVP8nz5K1VDzW+Rrm4VlBHFfmiJ6E5pSZDSIq6CpQJAft37oV/pNJ4bhXfGqFIRXMBXvb2HZw
Ce7Rlo4Y9heJ4JJMt4dJh6I22NU5IUAX8rtThh7rgL3xaImJhQQsGWJHvJMZPojcYcWHTBVW0lOX
My6Et3sp1mtahJk2G0lQs30LAgteI6DMqrciPsmLPhD4g1neoqZ5DxiY+kb7+T2E9go8nRPUlLLk
vD7kk0phqQecOfHyeQI+8kxH67exTMqpb2Z+cy+tFkbF9T0Y4vmJPObkJKyCxKhNlXMb8ILHn600
0jjCo8ZkLA525E88ZWz/Lxf3gtMD3xQhqy95PwEhzwdKdkJM8cEMJGUaJ9xNS/4Q5ayw2U7JYK+u
6ckZkX5imW4FCwqk/HQ3/hGMtfxfNWq0CUTixNVveRD2ib4FdIs7bIjG3LkFwasRpV/GblthMg3E
6d4DdpbYfJQMYX1SLyOOnFxSiJ3UhJsWTd2F1ZqXyDTIHXlNQJFB/XwuH1+41Qarfd0PO26rEE/R
0eDY8sd7bgWX9X7dj4how2QjjmQmdNWdtBIGsl+PBtI11zR1AxIQewHz11Vy3yeNDCy0T9u4SlMG
4MNEPgZxyu2DE2NHBMdOdQnexp1Tf1oMglKUwjZqCT202mmqjwD8rwKt26u9M3/HyOoHwdGKZRd9
0nqswGAFVTvaSipx7p04hi22edNnFPhXK3Uula5MsgNhfVZK6opo0EHs3ym9Ww1kJunOZW56ppRd
fz0qxOWoPWXJ+ifB0hwHWRqESlISnXmzVs7KCQASQd5vloFsduCkOIXoqiOguqiUs1tozbe73saS
vliPIHUhxQSdalptL10WcC+wg8sIi19PcbKIbA/Gz8oRGh1rJ/wx2DzQSWIqb4x6zmaWGIR8YU46
nb9o8d9MkXoysUto1KoJnQdL3sCXfY9gJfsFJat0ztEclnW4mcoKZabCX+ckae88LZc0p85ugdNc
e9K0QKlfwK7aAbl390QbvZn+P+oX6KGmSfS3vuRENx6OZC1GT8+ItnGdG18bLvZ8fSAx/PYbduEf
g+1mz981ciHPzQcSgcMuLHuqVveC7875qaHJEXlUbivcqd9sAcd6PtltJJRFeb5Q+LQ77ZC72OJE
W7rjsZ+YGIGrk9g74ZoDtyYmfqVThvOnS4+WZ4/iHhs4kXwaz+A/y1fll4gUHsDyPWNzMxGKe9/o
0P2qV/UtNB7YvidUmZXhPCNlkJ/IAkSLwNja0HmwnXzIgPZao5YhOjitXiEbJaoKrqehp3cQ5/Sm
YmyNfioGLnjMaIGed7h2m/SCNAVnaNfG/qsjJWOhGRON6fKdOaQIObctIOi2nCdDMvUMlIJlCHSB
WgoOaDWbf1zLaCjs39PWgWwB04XxVXdoCbwUH+IV0ZqOtXbPfN3/97t5lD56uLhDeI4HmFvQo/y9
jVx5hMSQHYj/J1IN1QY8I0Pxt1m2a6RfrWeM7Tl0O/itD+Ix83y4fNfXvYD8KsjS7ouSetIHnj6P
JE+bDR2GEj0Uje8IuSMOVnBsxvqhM9HDGLekEbrvrkrU83lXj/pChbFabYoZH2l0VNS6wd+8CTz9
XhE3932YOAdSmuKjpp01aE3gGOa3fwgxEV+01/V4uuZpkdqeTnFh7eWCbTiVUFnQ+Evkv2pkQykZ
ElxSiBQtm0ZKI8aFRcyy6UUWiZ0/GSiI5dpFMZL0r24rXMrFsY5YCf2bvfDUWoIILp4w9ildE9O1
od+pTykv5eFj5TRmzcmySp6W/b18fAF4iInrnTA1kKn/CKWh7Oi2L7LCFJe4WKM+80cEFmFMcgH+
H1av3K8Q3mMreBAFZxaCOMrv1l8aDcffL/fW/oOn5RqJ5hfFutS4l5dhX4jJRagbdJn9yqaZVAG4
nHfZQDwzWwD+P2Uaf7BBQcGhp+8l6ttO4RvLfkA3+59HjQRJXds3vN4kh2nRN7Ipr00KcfatCNnC
MKi9SVfjYbTyc/cu9oNnTvaGLqcMFHtj63eAErBAIZLGARXlNB++JXChaZkDxezRE8ed/fasGzlm
xbjxp/PEKPW5+IKzVp2Qdl/9JcrI0tQ0K1qmsCfWmz0IJmfCUbcpFJdcpV8IK/2BAOmeDOXgk4xS
kNWSy3F9Pmejfp4v4C3+fQMX17qFFQiR6oioIUzR0YIIfeblpaNTMAnGr9g7yZommlfGYSEg+5L2
txViJ3HB6bvinBs2hIfzADdZiAYgmnZASLIjWM48bXGsB9wzccQM5AGoIy7+M7MwZfZJwEG/zCvE
GZdajItcfvFAmgeTziKSp8o0JQoeHUKKNsRxWWNTKq7oV5jk0Lh9FO8RctxzuIzQ+PdtFO7zA6Vj
BmS4hVZFdtBBUeWqbi4VGFM/AvgklE81Cj7Ob3fClxT0COsa6nkIXRnhIV3htEzWeUVzIJNTXH0T
4bytD9XrFnoHaC7DxRg8QaAvZZTJeYXJzOWUWHul2LtGxkTtmcFFHRb6sFdVDJO6JtvMghqUCRMn
0GGu5/NNELBH8z6LjLBxBD77VMtj/YpJsQE9rzQWs8idgeCYI1q4uoPjMm8cnE93QYQ+cQGtCqkq
aTSZAiWufevR9HJal21IPUxmylUmip56/em3IZhpxFO6j+IwOTFB34T207BKFt11OKvnTIfhdKhf
ZIqlFt7VTAEPXKwLvISw0SxWqPNZb2LsyicEaVrwNhmTWm43RUEEHzLsw4R3UZ50hCEhQRFljP7O
yHx3RLMcnH4HgUlxU0Q6L+hFMoSXdtz8qK+Zi3pkFa70zKm1sebjVwVjXZk6E5jKtAUtPyd/s2TX
N3LnZ0iwSGWXqLXrtZ/ue4w7RL0IZs5PPRDH97loH+NZxc9uVEv8z9hWQ0r0vTiq4trIW+ISHjxp
u5ULoaLECkRHgPtIivTovgte4qECq70JS9Xp8hnDtJk6b0A4r9JBZsZNUqlOs9YkQzGsKcE47iiM
PjEkPmAo0QI6d4Xmok6NAu0vptaz78FaXeskBKAnf1hWKRsQaQD6EE8/T+l746bgiipK4PmnnVnF
D21MpdrO/LC2nyFa2Hld25zjWUDiYyifBzUKHqJJqC3tEGFzBWnXL+hkpz7sKekRc9fK6TC1nQ3l
hAzZzrNkDLKz8+lcDAQdsM1jR7tY2BUFslG2vVrSk2jC6yeoEpjUY+YC/EuiYJ3VQ00Xo9z3pvxq
PlAtjvKzyeoo2dp4rrfOATmj3KewqMO/R6wZnYxUxlFcxNrZn1YYy/ZX4Wh/4gicBO6YaaPA6oGL
aC9vh2xTxuEJYMGoAmBh9uaOjbOuh7bPQAgOXH9XI+SRzP2av8ZuRh3W4J3GzuoS4XFNh8RgjEu2
KRfjsLLyeoDOXucYV6V/NqkqWX+1wJY66I6p+q2y6sHciCRW9otQZB9HLfeLJ2f33NLxuQ5knb78
5IcJiWuTI0KwrgSS8DJkVcqL82MgqVOrueb8mM13aCmCoZp5CgQHxkP6uwjw4INUlTVJQKhhOeVP
CLuRgB5iqfid2992nx2iOCs80G6aJkheoEXb9asY8PdCASaG8oV0+c8kwf3aO8+/fYqq9duRSPMD
AUZUlz5hvlfhnTxLbH+q7fV91HniBYLiN2q8SMmht4NKZv2NxaO8/6wWl5/0LWXP+NKklCpOCHcV
7jto5jepGk1+k3t1dPF6N1zE3sZ+miBAIxkzfiQUG112ksj3aDStbC2EbYTt77RuEWQcI2nen4sj
WsVYotXl1zueQYpkZ11/cODu+v31ZYewoE3FU/XPewLxVvf+ygcxstrrlOiHvI9N2hBWSoq5zx9U
LB8sQNmWK/+b8DO19zKjsQ3m1rzT1gPLa/kheugFwr4/KeZdcAMPkR3usgbYnD9o5fCv4pDIssHx
2B2BcDaLmXaOxK9AhMciHA/l4/vyfOUlzZ/bd000iRisLxhBH8Rlf5KECX2KUN5z0IMB6sx4GEjV
xgr2yf5TtqqStuscZAzFeDpIF8WZe3buXDeak0qlsWoQr9CvFRRk4EqEdIPxWx5yr+c9QKfbYyZ7
vOrhPrbCxNbfb/VGkup3Q1KtlCmLjQ3iGXpEdBVOqgtHuub2+JegEpIH8YmfbRs95MHCajkJtgOX
x+rKPwft0bK4qD3tEQKwRomnCBEkDlL0DEaURTdxWKhaUCDl5XVwD1qvLKOtq4LfH/cQeXzS113t
M38NjMRmonsG1MMvQFdZhndDDyY6VIoZMIXcEeotrEoaCCaGnkRoCjOlZ0St0foohs7YpqRgvt85
EvSUQNEQJFjE320zLbNJzXbwQXs2UaHBnIW0F8Ng4ydxVOSiJtfMbrPz/q1Eh6mhBh6uk4sZiA45
qdDa8FoDZZG9+pZ8uTl/2koT2Qujj8rB5eCTyLJf4SnyTNBxon/Lr5XCYpULtGmPnYpvmdBA2KPL
p6jC1I/Oc+k2TLytuJ+te2RCoa8Ouia1wTY/jfNyOGPy7UF3AfNpV70hNlRkuzkX7P8SIClLj3iC
iXVAhvQXDhqUyKCtT0x4lUptZtJBh1MtYRt1r5FYqjf3ANwt7anvT4nJtPIRukB7NCT+Vn7WUyCR
X4vkj8S3Gq4cYgrH9LlBhNNKo6/5DmarcLmAyjoXUhXxgKSsqnl/221SLA1/1yhdSBsdxA03mBOn
oxym2MacA6t7yniUW4j2V54bLeDKhIDGgzUbyq6R2SkmGukPgWOc546pJH9pC0OD3I/ZCkmBl6h4
TeyicI5zeTHnmbI/IODRSMO0BupsM1u5E9neaMlhTMs5zAuHtj8q+n7s1QGHvDyVsHcExFVd017u
Zr4Lv56yPqsgFvmSjyviGT+GTJeXmwGb/cKOfyN5AS7O+tJtBwde8BcTdnGxMRwY+pnaAdZbmzTF
tKWaT4FOogVcH90RiPWy90vpgbYVu0TzDdYvqcp3grwFB/1wx7lgt4/hi2RAxaq2i2Cz/1L1XR4v
qVdIgDLOmDVMJ0PLNVbHIO5nCQSx0e4yCBhFoIBOgGxUVlT7ueoGPsFv1pdKrrIsTTgZN/5hRpdD
2xmm42pxAEExQbrSf2gVKCg/G1mJeGalMFOu/Cn7aTSbAskOI3DEAD3SOxSZvvQo+RD9fNJtB8QM
N7UBjRzaEB83YA1JOpZ1vROTO4P+qbCFQbzIVO/WIHiSKTjRCheTmIssmR0LEUrC7TCAFt7fmi4l
4aji8gwUTbULK90lXsG6dbvTcaSjqLPTWAu0Ndozca/k8GbrcMhZKVw+tZ7zntNSybfbm1d07Uju
I3Uv9WdThZFKFKuUPV4sQMZE90agTWOQBWjZUPSorr3JnRViWYUPZ9+qhGoyZk6GssakIRh+OEVF
qC/YVMnOlqF4MGlUoMA1KXki3aOQktNJt/stSNdVqusOaXEzWJ2Tbto/OgBr+uWfKHYkfpoqfcCc
GD5AZEKo3KE/UXfiIe44CetBdxP7WvFo3DQcAv7KTDcP+58nle63ql3QM4YBbksOToRD3PUgrF57
5MdE880dJ5Lz5p5+j0yHQiZHEvSfx933tgQddTkFbgrWaX97jkL1qbC83yl8hcZmYJkZENQDIqgR
ufBETxqu7KotHQZlqypzaqKGCzxItmJCeRjk+Jh27v5dgo7As4D5CQstVLwFs4yUQhf1Iv/gtTNz
aln3FSE83ddZKPB0Ddqd5kxQfPCcduEQDFnrHJBbD7F9T69sBQoCpjaUrNWhhZnWq1HaX3rLwEWr
FgpFSlYw/SfAUPguHMuZ6qDs70hpQzhP8e/MWVGYC2PfQDPAZnBJcD+FZu4hxzlQbfLCEHirDbgL
WVl5YLe7ktFxhESUqDCK2o9iFP31fpkhBhQfbb0NALyT8RMdqHo8xvH8/Gb/6BQzOiOa9Bjnyi3u
ArxwlGb0Y26es/5R/QoObOkgTi3AW/D3RS4AKbH3WPbtvaC9phd7zEBJZwAOJRjdormgFzUVXGkS
SbSPfguU4YSQ9AY7Kdskzx06cIJ5DbQUe+ureUPBZMKEKd9dEeNcybrp5vz63Yrj3cuhb8ert9uD
lKQj1ZG9YzbnIvrb23tz3mSlL1dg/NRjeb6k8YiYE+HJAEVZrzNEZLgjdRAWNfIDYqWcIEAYcoTo
kTTnoOc9Sythbo7twp1OmaVsF7ZfjxQRHJW6aFFBhYLJi+TPIW7D01xolJ2wCYrjmlbtNKz0Dp2x
HHmqgAnMnshaQ+3yhEQrX5ZkCosPAKhEwOENxaEzi/WN0tr8d7tEdioSTaaeXSjTV8pYgVMwEN38
Bdeyuoae6AaaTWtc++yyO7PUdFZyV0jdQ019yrDMAbKZ4y7Q9iCvANpbX2M6CTaJA5unAsIjj/Rl
1+xmhHzF4m+W5V44Gu+SpHBBSi2VWzwUrtHI81gFmnChPpSTOuDRZm9dJF4Du/dPLfgc+Bo/OhjU
GOo5JXj2/jk0xgllhjNG6KGU8/K6znk6m3yz+RJ8peS04Fi/d7WjBNuZj6TvvZfpUb3fPRfsv/s2
NXZLacZedo2dXyA4jsAQBigTtchr4Pn7YqZcm81bVgCUZRDuM4XFo8L+TCa5MmB09pASm/O1BMki
OnVzFb23qntR6y2xP0OR76ieV3IShHSgKwVEsdYwNSI9Gx6XPEoSWGBDoDwd/B5jXUaasq7dyowR
8ZbWzlQ1kfEPxfdQhMbRH1FoX7tL5feoLRokxlSQ48EfjaA38Vyvz9wgK2sIprfy+4HZFR6OFoe9
fbCJBqiFGh75l+f4H9Iv8KLdcnQfFNLOK00sHdO4Vrq/MVrpvp02qVe+RZB58fjq9cFV1i0dwzEp
IUJ/a8LNKWR+xFGX/n4bLeh0gSCXQO+GqBJYPvl8foHnbDtuopITdgY47mrwopw4hHnMmwVh1opS
79Dod4Sd+yKxJvGhAGxhUb6EaeYAmFWx8HKI/YYmxmCG6SbPxPKrDtOYcikR+26vDmm/gZ7F80NW
Xc/xMOmaf4bM+kv+eGl1CF3dVLZgnF/KAQEF31dFq93feidXwJrw1we3I8lS3L1HFcyOcjvWhp4T
h1ycFyjlkiJkv0U29JSiTnCj9xruzeK00v+TGDokft3cy58e4n/cMH2NrIXx4B+a+qO3iSX35DGp
PPA1zyzcwkWvRIR+xEBiJYYHaB8JLcjkxFDyybhjUDF+eoQOgIGN8sWkGAcxwPPan3SpJCpe+srE
ae6zbUY6cDco3fnnHMuo1h2VSQvKJVHaeniw98aBqNly9XTzy1sGj8Y4rEaLjc/mkY+NY+mNHEtV
iLvhmyKxr+ts5PdblS+pUcGAm3Yk0uldIMJdu9KHJ33IhJP071fRt5q8Z0sky3F8oqthgEhMkNg6
1PxhbTYgkw1UrUStAf2T7ZBPmkGXF+Q7ovpeyEtK/RUc1g9nkEJOK6ASEV5qcYjnNDy19n+MZqH9
X5mcjkWyLQr/TylEvj0SJQJrGuDWjTL9xewbCod4VEvOpLB7cduENIH1kfKwj/EI8FPwZWm/uhjA
Zyyjs1W0Ghz+irUVyhw3sU635gSV0JfehPoFIok4sUp7iY/TRRQIzH4UsDQ8I2erpl9rL/xCU3xM
LOHfnAeZXYFlGyocpjmZxRzzzxMHYgKdohtjXnZU3qymkB0IzfDoZVuZGu/WBQVPU7EWaoz7yfku
8uQ/lVG1M2d05fDtHUMbO/NFWNaiyWYcDTadfZyfRNgwr/FDb7IUuZxsOqU+KP8D3qdm8KkI85FZ
zXs1KCL0SQut5dZsD++K3bj+4DBcp8AFngYKsYXtx/hDG3VrwTEWebo+7ApmcWHtNs2jvSLlQpjW
FmpzMS1vM/gxHkK6H1Qldl1oym5qwSd3vb1at2adMyuMwqtC7XfdQaQF5hEPJ7dI/eW4FsC2Hr8e
BX4St67Z8GQzwKR/AZ42TNwn0WXHha16tnkYUd5C7njmUpItYxUq5Kk0fUONLXUeB95/h1+gG76D
sK4bUM9W8YLfwq3z7juP5ZvNkBIRC5PI1/YVV0itbC7Bhw647ezoppkH/IexS8Hca7eZU+dF05Rj
7PknJQbh10+IySyxXlvr262C13w2E/BFZiMLIz19EmfDbLcGnCtY4IZIXZpqPVLWnx0T4KBSCPQ9
XmPdP85bDSB/yy700pmIMA+q7NNX3/xanu5b6M8w24Vi54GWFNNWK3DdXVKlF23KKJTtchMkIH+a
4IF8uLPvyG+TIds0jjuMv/0mk3++j728Kce5IRze2qhiMm3A/D9nNELRjWLpngNADR7j3MQI9ttI
n32s+egFJnzSASjH+OzmR/C4tszbPCvCIweYiwhWSAh6JQjzBiL0LJjBPJcCQCbf7Osh6c4g4GmH
f6GUwhUXNBQBRWoijTXKt2OqfTFEHXOD0fp1IcC41HYw5oBKVQDEXotnm2bJ9CFdLSUMKJEZaXRK
JvLFzotzE3CQTtutzlJ/qBFJLyk8w7y69o/L3mjn96rX3UYlGE/DtPQDdm2rC3wCD0AKi7IGCjsc
nm84EvRtukc/3awQWkkPymXjy2RTRaYaskgQJhNtXqCDQNZs01HfOiHeS3kf11FWZgIGW2JdG19P
6cY8g0vS0KfrL0+3A+l4WyK+6bIa1GbL/xiSYwc2okzPA2SkPsisYISrAdz9BvfY58hbGg8VC/3j
rSkRfnSAABKMECHQIwA//Pg5gktwtWtIlTSEco8WMgb/yJ3kN0bJuIn113uIk1bXcH0Qbq9EpEHy
PtvUUvWeL4/XmckWZiijEGsI14tKuW0/3B+5J7+sAZGrhGgVlk0iL00PWGDDFng3EdSP0RuoCeOG
TEz6hVpwNwrwCNRdoa7mTIhh110BeLQwPrstJzk1S/+B0NpMdZSjEw7WXpC/qko/Z2iB+e60EZGC
r/LQl9kQeX2wzUsFdoFyJJaq84l7UAKtyHRBV6aNgupYoNCNb6RW3HAb9vp00qP+nb24KQTz1cpu
RbJzIcmdOax23XO5vRF+bwhevc3lqEHKtlPiTbIAR8iiBDhdOaGEeZTOrwJrKdXV6GWE44gjVnQz
PyjJ3mFgOxZ3f+65maDJFClWCtIC1WCxsoVV/B6YkN35Z4+k8er53qQ5PKAdaW2USJmWONzKjyEz
Fhy1+tlmHQfZaRhSrMzTLWpEDvFKX06IAhh3n3zkLOcg1qTMLQLQNzQDGIlb7sGNo30y/mH13OC8
mGVGwOcjJc/Gvf9RZ+P6U60EhpROuDAqfYmEsU6I6cxABnUSk8GF0osMBOalckhmKiuqxtqI2c1I
ravXQT/vTGEgFDT0SmYP4nZxfb1YxVYVEBHhv/x3K7bVKTGS0g4+40bAlGPNi2Bw6taUwdYrlGKr
FOXSZ0bGYh65Tz0ceBVseKn1CmPyaVTDF+VZN/FkumTCP55C658C0yBnMFYz9UdWdacjv9i1NcUJ
DssWVreW6hvPzoW8iUYb9E5gcGQJtUT0f+DWgDkDRbN5VM9MAdSeSroHO5Gxye2cJAcUcZ4Whlsp
BpRb+nU7sV1Uyp5AdDtrvqj1musOsoH8cQCqSXiyaqbdP8zglZZ4hkFW/YflBr5QHZ6yR3u+nir3
BljpIFZ6tGStga7RKS31twGJJniBztTCEUmIM+oMlgKYj3QVuCyHWhJRc5d/frv4YvSuxKzFuLNe
L9i3dgyCqHoCJ+L9/qNfU2nh65QNpF6mr06AfBeDyH5RCnkd91R/F4ztTiaxIHzAB92jaNznIzjc
mmCYlQ6AtMhflzu32VACws8Y7KPYH/5N9rJipwznUClnhcPesq+UGIa2IGjWZDo3nCBPUjLFmGar
joHkCE0RP1jIfj4ZUo8XKa+cDlL6OclpTydtcQR6q9Uw83DKECZqu+cPwtWfq4cRw9srDGM9ek1W
WZoXLcQYVUF6Ah38DS44i+eBZ84ioGf5iSp7ciwKyvwWp9ZS0fQOdjNi7opVXarod92t2ovq36We
wco6PC4PPmLyq/C312E77+5OEVxdKmvUfaGbWCeFMSF3PqtCCAP+wjTEyHrk92mY3D0I20tBAmv+
DFgAYo9JfrEGJV7HyhSbvjbZDi/KlvAkPS/6TPLWCgHkqv3wMC2P0bkWvHjK56GSA+IngifxztlG
MmTUsALs8l30ux1rrBZp+lwtXTsI8nQrm2PAAUYjhUxoTy0Urbn95u/gkpMqQsBQ9589i1QvJ/55
1UpYD4UpVuzmam2q9CW17ALVB2URuIAQkIHpBqVzRYMmreB8can+cLd4W/Dw6PLgP7A7Zo8fr/pL
Omx4lFEXo71MBpTXvSCiJlF7DkGmTGZuNlfEK0OtoTIoraTzJAlZlg06JIkVhcBeE/iPAhmR8k48
hvIX16X+pDDYgnDGa0sNz+3ZHC+ek8kqLYp8oS39tR3Du0XVX6HnpZnKY2zMAGOEsvJvx+YXlG5z
3SOITjKPf2VXklLPrRyVFtfEgB5FGkNi8pXSFyRuT6uEFfePJmzlvJJ82mZHY9IjfLCHvL8PatdM
H9Hs1VQBXRRJ+8I0LtFG35cS1urPpAlN6V3NP6kFzJ0jTSslFQTsrXNHhmP55hR8OfWOYU4mMvcu
2g6C4M8Y7Ch8v+7/HVLX/ffEaKD6RUcfy76qDYaE5qvFBhdrVCSM+H7zhTMMiVtLk1G6weKMez4B
IfJN5aIe3ECWv/7IRx3mpX1avnNbAXqovGmiut1a/fs+dcFJJDF1mSMHiRh9J198eXaoQJF/ZZmO
bTDwrPFhP5r58QrRV+5RK6KryIo98sKRx8l6oD5vV70rrmCiD3AFYRHRPl4e+/31EF06qh6qt7Xc
Dl+Y8omU8N1WS4uNUvXtqpSQOisSMsS09daOxiJHjp4/Pdfkhjjo17hufwe1kkLPKe48HxM/jrEY
PQEiDl6bj2TXcNEqG0w04IwW9NdF81n2mzuISl664d+CShtFuj4axpmWr2q8okx7MwRaDP1abT1o
LQ4G4CeAqcxMxR1zLQqzbgakPjalprD/18D3tOiYnQftW8dO/27GBo354+9tlK/IWO9MDlbNxOOW
NSRU5t0mPjJdV3KHT2ArRJLsQjWsR5uTQYi3E1W9pc9EaKv1xlYo8yvlN9gY7Z312fffLynzzp5M
f+mTreFd6oYsiec7Y6O0r/dLqGDtpxPeso/Uj/EPdk547bz8c5GQTIBBe5k9GfKgPcI94gEPJZdl
2F17Ff51ACMXiO8umfOoi/cdpPJFU09IeAy99lFGT1eeFVY3zJz0G21TppzaIgYcrykvpVvLjPdH
T5oEo9tIUCtf7eAB0ZSCHY100y1jfY2M8a4YlCkZvOrWwm4hXfArMFf3TRFZ2mOo6Z6SO430+LtG
JYMREhHc0quvgdO6dBTRByUiNA85jSr41Z6zB0L3kP5MV7mW1RkxibUi8W737XxuPVno2YZwmTrv
2cgtlChGQg82AkVt0cfyhEwVDL3FK19T2wj3792nb1iQ3TIV1oAFIw9/t1CHBOxnCbffEL1GQFYE
65CRsibi7Fb2d9KHR769q6c0IGxxLAZ7cypWhGV1GxNINbPiHjqb1cDGbSR8nUFDhZWSw4YpfLT2
7q82CnYHrqwlu9yz93z1bb/m/oTfTK8kHsgxNislARESaeNxrWkPDhNAhGEaUmTxLG4VkZSth9xS
+sxJnIIwkhcaYbTgIsJuF909XtRc+kGkoKnCCIQ4eW6kfrzEs4IRaGY12L6lwud5Vz82MKKRqpsA
muwkbqbVt8iNbye+h8s6LfVg5ulq2YOkc0zxtnuJcsbtNTiMCGdiWKnEyvJdpZVaV1PjC0f6tI4e
BQ8qLzTMRgQrzzZncXGgs2uhVRjaiQrYlk9/f+r5qFXK79bHS4rIcDpOuurTXAZymBHekaRwwvhB
7sEJK2yNq57EoVm+eY2KuLqITUHAU2kH9OkM0W2EPNE56IJTavzxKXZujRowBcc5BNvpF38roGrM
kuTmIy51hvCoyRKH9ONWa8hq7hnc6S6ZVerv4eaYd4eEmIqebmCFewcmTPW8JV86xs/V03ja1Qar
FXfHbUP9E1f3x8oYpaYUQmk0v3sPh+2b9E/x7ghky+fYcz2Gd9W01gCXrZ42fce89Ta+SvxqTYlu
zsJbRzAmr8CC8KnWgsx4rmO+hR3KpNiZ4tl8tYddBXBXmaJxUZEMVPVlOQs4jAI+35LkcaSwxJcW
lgvX4yuuL/u89XTfJen8Q89C3C2v9NKQEfnGBZWKv+0jHlWhe+8RB4O+/HMKOTipmT0xRGKwNJSh
/Jb7rjyQHyOI/FNR8lD9i0lKySpuWDoaXKvzPPmQXRrv0OsRL/y0DZ+LEJBydosBkM/lxBOhmysj
5NukIZp5XEP/Q4GY0T0YE5X2la9CP8gBOgYM6sHKjY9j+9/g6QVSrdnkeaeQVM1qOC3KJW3MuEe2
DBzHsybGqowvRSc+35bwdICwen0eqxhmPQlBxdGRU8H8GKFBH0TDRFoioGLEjv+I3P1a1JVmn95R
Zhek0M2k6m3uDxM/WJusAu/t4VkLln1yuyjDG+NlPyRDnC8tVxsFMKMfy9vh1LjMsPROV5XKuUuE
SlvSDM4yLZYrxyJl/rNcdLEqaMfEYtqCCpwmUxWyiqbXEqHJr61b5oCvMg6Undmm2UVIy+2SS/km
a0lvCwfxZj7KBfIuAz3HiXB/Wqm/w/NRpUVhHfP+PlcblNWFVhgie5IR2OCKFBjfEJs4Bm7RV8zb
4tvxEeg+7B9gkIWbZ8MKMJSQ5ieO+1syYQdi3crtctXS/u0o/pFAumomCMSXuiAW6OCMzVrby+A5
N+sYEy9RHTITHbPP+/IVv8zXCuHyedLvTJS5a7nSXJVHXAo2sUsvoUeIhR0ohY5nHOCkxCb3NfjM
3qbEBXUpVwh3Jf6KvngAyYpI+av8OOi03usb/rKjlhmiZwnkZ3fkMvkq54PNgtdU0W917hpTQpdk
KB9yZQvctPbfRqer1RmCI0ib6OMkpDXsUzHBOcrmzALrAd9Sr8fLv9B1zhqJToSAM+80HEv+vwzy
VkQ53rWX3hbhSlw9AJinF21oISf3ZryfkcrCLDwl1qe8OKT2dXeqFeg6GEG5z3ubhodPElWZpNdF
Ba5ImYX9QWjIromo9XkqIRM1uXBXQA8GloM6nq6+pJGtxjmSXRH8le146mL1hnlG8utlynvz8jwS
nGVS8+d3WgX/UgIyvlfg2zQ2CONdYbKJYrphCh7lwhJHocMbZ57FjVPf38ScZmo8yXGKSsdRD/S/
Wik9ZASPnjIspnxlUo57ptngVqHBdYQfxXuyZsVA1HEyD2Q/pRIvmKq/Ucnpwzoq689noGuMVWRx
CpveoTUnlYigwwi/YWwwhyr5w/UHrGBPefcksHYJeoFdBjQncmm0mr+0tlX5zaKBC/bmG/zT8oyt
mhOuYKO/JcRWyK1BkiLjwLm+vOCdJipPO1K3GjUjZVnMYbW/1e74WGvp7M3Fa5KblCTTF3SfNMM/
IxKEC5JHCniTp9czausAUt41EeR8Bujr66Fvdel3ACozNhU1yu6GffIqqDgviki4iYEHWykuQRry
N3yrj9JUjkwbS1AYSltTc/Fc6tpuys9Y7EEHP7RciCtDFiEO0AMLgrOz21pVALrqRCT667a6wN7I
P3TCX857W3jpbbqNHZfrpVA50XmjPvltsqFeXcCw3ljc+OwU0bWYCBAx1IiA/BHDDMSPvuayybGh
0h84Oe+Bo62HX8HF5b6eLhPzekzD1jP43d3MC5R8Rmi9dagZRCwWxLhirGrnFkS3Nn939UAB4oaH
hANG5E15BjAWjwqMdhx26lF+91CHpz87J0bD35elpNlT8Qpn8lMm2wvSR1s7nP/k3zQmi/POGXxm
f+uQ3pDoKQu/qiWyjFgBwZ27cfaKgoG1ANb5dyMlHgTCSy8JYR7fXPkGPVIkyUQR7ZqV/huOO6tA
99sqYZKjdIza2nicdRRmhk1LC/DHRbGR3VvOYQWAeyao7aJRYvIYMell0Cj/pfFCkjGjK3Y7dr18
Bnquhv9nllVcyzUC1Ho6oyjgiWIxriu/M5lgaLfOQSQBXLwKxJoIwqe9cLVWDmkZbp6LkLiz6ioG
QPKfw8yaqifNpaj3t4iKXjQ0DeUkj9aRddCSn6t6tiNYTS1CVstZ9bqM98zOrjs/88mqznREsbVL
jB2mUbWv136jm7WLSHyzJsB6yWsV75ep0eAhN/iTp3HtX74eEJk6iovRzRzjus+lPWPe5dsd3RvO
o2HFXrV/XNoJhAi/ePXykTIqa2H2z1a+0ZeOYAhP/TtwRlJe/x3tr4Q6f7whWPt40z4NO4TO/6qV
E1Ejt6nwWt8V0E1wQBlU2ZU+B2VIbozraNTLjJ7rPS7kBOKJ6dezIECE9qLFJDkRpP+k/NB9H1yc
WefIvfnMfqNczwoZnaaFL36AEDt3cwKCS3WThRswJ4z72fr3qKCgzzfAHrWEOMIfE1AXi5dQ1AiQ
9HmzuuVNbvMLo7/imzUNfFu5MEQ7YI8KP+v3wPSbfO6fxt62JBceOrZ1jxpRGrpeFJLdtN31vOdO
CAfFjcyTm4wQzgNlkQ2BxLUFCW/G0JZBBExaxHx43An/cjah8C/cLdKyyZeu9Nyq/E0BvhNq3kWX
VV9MEcz0hRoiwjfeb9dmTXGvoppgqr/yQvTKyyth4xf4IL9zhCa3f7s4rQ/IW21icoGSKn8vCw3H
SCV7B1VozvRCemXHAD5U3fRVVhWHfVsY7o+Acv3Yb5Nj/WUXrN1OJm2wDS+Zk7+dsSTxfIAOzmej
raM5log6s0+roe7OoSHPYrdGy6u6GJ7odyeXHUPEdwVRRfFQ68GgvKU9HENlVDpWfDBIWMS+/Bxo
SNnI8S5ZuW/iC93x80LbcrYFXooOzUxCbhmv1hQCl3xtIezYyl4YKMu51YXLHlPq9G5F88JA2eMg
O3OtdXVJmSZ64fgVNLSRmDkEvpXGheaPNi/jmuFlKtGviyg4psIyHAVx26D3tmH+rQx9kiL859JA
QS+vXBXkkhuLm5CWaWwgaFojzXwCcRWXQ7R+EUmkHJjEtN0NlU9xbDrCMA+aOMBvuA9kQnCdhlrS
9V9OFrRAgDDHr6YtOS3NR1I/N+xdt5LYksXqRG9gfHr3iW4HfMdsmKVfVRxKNXodjchiozxzbFUS
nD2ZXIMaxIbswlpAlBYDoVQa7HGDGhWGHfkV5n75JI7Sjx1AFfwjntMQJpqmPpBMlPdPQBKG6QPc
wiHhaRoMwdRfYp13fCFc7S8jiuJEQhz0YaLeRMgk3mPzRNMkhXz6HbM0KOEWBguc76vVUGlZkuFI
4ViI87Qf3Bv9xz//4Cl5EwKBYubleSNXnPytjO8g9rTayxbsm42rOWFp5hEpy1uOfJB2DL30udos
PW+YF6OAAuumLWzRXsIYVOuz0j7auKvjuGGbXzJsVC/rrWikyAyHME4YIACxMzDzh1U2sNPQkJYX
299hsL7k1Tj0OTSMqmI7o9tchadoNu8XsEUWMT3Hrk+9NuU+bekAOUIgBlyNeNba2mWHGMIZ7c73
JG1xWZf7VK0U6n/NqNoGxNJXbgeIKWMU40M6GgwlfuWsuB56dIInC3MYVmkC4WkOa6knN6POBU1a
P7XlgRHXXreSPX0zgl2EGhpyQnw5eB4OWyiOtYDxq+lKE/jhWBXOPXIFD14fJKUlA7K4ur+7ZVCc
2lvt6I7RKQhJcdYYtGMxVQSyjUZA48wWgsY0I0tzJgqYLM0MBmFLE8+3gvXIHgyR5CX6h8mG1FiQ
hzOCU9y0qfAUyzrLjBpCbK3bI+2hF5uR+yD4qbPj/oyUbwCt4mZdEKyoa94sre2d0Fd7N6kkR3Ea
hD9iQM3rxY7V2OVU2L8kvkrUChFmBNQg+FDQrXHah4gkNvXzjJKt762w14Cf9NJX0ZBEElTWXkY/
tZ5BCs7LSSJXOdBRXbP9WhffjOxBP19i/c7QVg3EtmPobg84r/OkP7HXHVlAgZizUjFWQskJF3ia
SM0948wej6XiVOwMCAOn/zqfutBtIZtdNVmIxnwRAnZRNllc+1vG2/zODgdnPMKnc0uQYzYW1lh/
090xJTUm0nCVdpZRY2Ja2DEWYzpslpIiRTo4DfT6ZHgzg7BtPu1KKb1hqpIAO6Uscif91EtqDBVs
5Jtc+LKMbmHT+CVgY/y6G3FP/15dA/qXf4R1vpX2EFhG86U9RqgNXJW8jxAGaCbB//zHHUi/Dc+8
iPk5EPk9Je5nfUsne4ynJHE5pInuTit7hiZFPYBNRQnjnm6KT7Mk2P6ZmkFaQSD3rc8lJUWd0h0F
y1tEiez8eq3aW6s7N9etQE8gsQlOrEUdVoJBXFxvhw22WJA8QzSwB+SDcJ3PvKvGq0b2dq4TwS54
cyfqyDMWpnkyzyLM9NGaBZhTAR8UbDGunkWvGfYCRiCtFZH9g3D5tTNTmIqpEyA9IGHNlGRC6+MB
MtUbILhaHZAVWd0scvKuBLUJi92FIJJXwrGqfJ8MTim8US8pHOiJ3L/I2kP+HcAX05Yo41q+K2Ou
C6+xl/JJxf2KKATlPa1kZ75M8cl+k7TYejnptasnDEDLCh3pzOWigqUceW32E+1L0tOQ4LjaESaI
3O0vthhmnzF3gALFLeMSyRVgLNaAoXSGF2ZHeyBVbsWCr8j19WRxGtF3kjlxAmSOCRhRoPfGdoV5
9fDkb15Nk1JfBqj0O3Bazmv0wxcqPj+7D9EKBeyB63vnc85tGcX+N97T80xRX2eCCz8U0bnl2uBk
l9QkBZA2kFoR1sprmwkrwfZK70ZOagzI7srXPCrU8ydrkjUsKlGOXbVqQSl/pseERQVDspcpF6pC
LQtjJMapORcTdw5GKiSupAe6p56vSvO8ne0iHaWypJCoxGNWLRq8CyPM1UONZJGrfvYfx0t0YXAQ
0ny+HpikXb+aE3wkm3Xk4gMI+cG7qOvXhiUrFZknETx5GvNhuWvazcUKJMZZ1OdFtozTADBw6qi9
YVv6ppHVnUEkAbKxp3F6YcjxRe5dj8pm6jd7ncFl86hLW2AtPOIuMLfFEGBrC0qwQDXgvf3HXfZF
vvJpVKuWRRP2/Ep480PUAUO320U4WXGK6d4VNvDzH9NV5ya/1R1qxBpqkO0qqI8F4hiAdJpiBXrD
AABrBKEJGFFq0qHXdBRQtZIxO/1qcTRdadBX7+JNiL3vMTtn+pfY8h+JEiiDOatVs7i/OhV9BV7G
O+QFdy+qKy4nkkRKH+PflYDQakxH3CiC4H5zMXUuRseXvwTkMHGMB1NQW/z/kFp9exPr5wynsTgf
79jSTePRP8UyUxP9/MBrpV2g/CJfLlHoeGPS6X1pSBBKVEuLc6m3Nrgo0EFazjS3Qmkv9h3C+96I
GdfrjJWMqXhXg9irVvz1iFMA3T5EZaUMDyqX/1q8BoW9red6wZN+iuFTB5ni3eoDdTAz4xu86WMK
ZqGZXJfa4/Krs7JufHha9MgilPGz+2EBrluvDMuFw00p6L3atHE+Ee2tYCEhHMdK6reQ3BAwutTY
LkmU1GxnBJmjwsD2y1g9JI5PAE4ZZWdJwPKsP9Xb1eLAVDqG9AeHiQgafhSYpnfAars215mkdV/9
TzOqWEiIFjRBSdTrBvbLUR+BK5J2p+OlsK4Qi8noGvWJdHEP5iNioUEk0GkETrOYF4oi77JWTB71
zBU4jAJsJ/3V01aMd9ivu3sIRpGMptF/WRrYz8UZrT6149/W001itk19pldPEbDxIXFlOCKqs2Pg
ib/al5xgrh3IzqQmIKxNMEmoTkgRgSVhFRPG882k1dRIZ4Se87jkzrtmpEhvCszYq/EWUp7ZDQaU
IvopHl4YSLSNF36Y9D3FdfFb3mgRPHtDcCExqInpzS7QmB4eSOldDqgageSX8kwgPVq605sMXyI8
ha0xcz7qU1UeR39bhtFrz4WyL0fsR6AH6Ysbgp0T7eGIWHjwRBIJpzIScZo/wWePSzP7Pg35NU4h
o50LFiZRi7oARlcYNCsSB+JqCS/o/aTaIBp5kFyCFM+u9I3nMW6oWem+yHhxb2S8pXYpKkpAnNkN
haxL5Iwxt5c4AAKZSqRBiO8RFF0GyoE0AhmhwFhxwEzpeDfxD0JkHfA65ft+q3qz/UnI97FtVrUg
JHRF1hulbjtRoBIV8c2D+pdl8Njuz2DhODtCD8SD6f1maZfa8dVrKL2G7VWurK6nYxy7SadYZBAu
dx9Bx9s53U0N09Z0uoaeK70gpGlE6jhMoyC57873D5b31I5ECbyr/AjyorlebzR+WTfyhAChhrN+
dyNWptfvfa/ct0KRmKC4QVgoBSvr3TMBX2aaQTtSl1rfJToUEmE/j54oeS7ejx2HP5Oz6AUOiN9I
xmNCch8edb8sraA/8eNtw30SXqJUGnoZaFJ4ZHn01CxIGrkOdzb0T+1JKq14g1ycRw6XkZghZYyv
3ZcPdngb9z3NiZjF5naFlDRbAN2V2msS6Sw+gb/7wSJy+qSqPgTcsjnXx2XfMirBYnRCaYeTKYeb
84otT4etMoP8WLucuB8Udz+VioJ5/LvuLfRjTYA8l/LhV9g4UTl5ZnWq62mtz9XkOu9w0Xv/mF1s
bEk2K1dOan8UUSDCmIJa/vb6vGcXlrbQIGQweUnpfRqvfshMFkKcrYWwkOArsN+duQbcHJ8Mckpr
3QKpUGdQ61Xk9GxpHYbaoFmZsTBoY2BisrZmG+cC+ADjRapE+TtccYb0ctK1tacAWKOpFy/h74Wp
s/+XggE899qz63DaK7GvuTHOQp8dftOqABBRVkigQOzGQWEqf1OM2AvSN7SQxXD5WkbytjnBMict
mEycBg06x6YhCxDU2jRe8fTc9jyJs5IXk5HUso4CEs/zezwJkkbFoKBK0XRVt+wpllOb+hWKVwpH
2tqUAilkjr7ooGQxjclEZ56Ue2pvYMtwbNyIAqkINF3Er4m8wNu2jaSpzT1m4e1bknR6bfErdwZZ
mC8cJqt4qxxdrsit6SEfvin4LeIGgWL7pyaK3D4ucrE0UzrRhuHIyAwR+eS4sPjCz0T6Xf65Y6HL
ysciP9eUBgmZ1vC73DO+BNmE3vhe+Qsm2+1uM2ytRT2h2Pd9b5ydrjuv9BDy5tmQ5aKJPSsxNPCW
ziTUDkfqqmQlcZyNlYHtpZTpaf88AbnraMi8n5YOjf2vO3k5EAzFjSOJd+zbQLm8gO8B0NfbyRcx
qlEl9Vru2XctcYqsV2FAAf1Ke+lHM7MU4O0hFmtXek23JZBNyyxte6a75emjkkYjiEaatJ0bQ5zm
WthiM4Nr7iRqCIn1f5QIvm8MA1Upx71v9W4Zx5zjhyoQmFLdMnLmnnVFNhkrVfKv/e9iEhQ5b+W9
X1Iw/hgYEKZRSf5EtCqsXIDLn/SWJlLvl2jNjcg27h3IiHxGmFTaO2KFfzv9Av2ajcPqHjGHFWXC
xZrl3kuc66l+iL7EjEXKSyyv9iaS/WhYYHY8W/J8VUWyB5i8ycB1I7dp2FeVqB95nZU4sxk8zPgR
IOYrgDS/LO7sFzTx7a93Xtsim5gW9syT9C3pm6z9PkFRCiEn+pNpfZCEhYm0njq0oQKVF2YvGITa
yH5B84DdavQ1bvSm7Unr5xhFMLevmAzvlLDVFdFLEJTp2ij5Jf5AvQrZNFuEL/B5goo8jSqe3Qml
GSxfA4HsllqlJh4fAKAVMuYJotvLZoxk7hbfQRek/BZk98ukuUumCy4tLYeAGdna7bIJ2yz5iEnv
BgxokuPI9qqtsd+l51ZuNV0gcxWLfgfesqQvV+X3hpVThMOx40O30xrXW8X2XWeo2jD0UsYEFmAl
Ko/FadqP/ffYxdlO4D/6j5UoHfs94KCuHt3fqOMkNFAS5UX168c+OlK44H7+J6pNToryNVVi6HSe
szunjYgcbj3Ee0U5IoTv9DNV2g7j0kjc9qobXvj/yznTGiHlWPwYBu8SSuyZ1hWCRt9RuJ8GRBeG
Z7daerFHzeYuH/pXN4jBjsTmUxR2oD81uBahJuaAOA/1fIUXq8SZb3ZsV51H6uqQ2+yUp46umzlH
zvAvXYWvB3zy574jbPyVWwb7Ps+hc+x258mVvuqiVaxIHtMoc2s7be+/My1c8pRyMwuL0KQ9fU0+
NEAfvYM5sdAlGBAFC3+oKHn0dRdsBuzwaqSFSVUlVu31OSgTRj1oCedYdyurh/MSQLusFOVv+AMQ
c82wKCa0wNr0JWqS697fruXIvIArID2IR1Oue4AAeVFdG+U0+iOgXUGMwhWzzd7m5U0f6S8ozl0Q
1F9QC4kvshGApUWYUNW3Atmh08z/IiMJpIYyOQyM98kFgFuZRCVU3RYNRhBxiv4VTygjNnz76men
NG/SBGvD8oHWvxDxgar9M2uVPbUQnvnzh6ieVCVEqYcholjZdzfWtL/kxpHlRFdrwdiXFhi2CmxU
uVc0QprmQw9PmWM3ziWbeLzFhhYLg/+6xQmGPcnNCe8+l0ALAt19tt73SP8nhZh8WHPzVT66m/0N
ejeHoZWvkXX5vovmSUxKreTx69OOAoAqR22/jZmvPni1U3Wj3wL80eBOh7srJZZHKeXIMUGfByPX
NmH5W6RON0q0+73AHS/h+hmme3QouQxUJ4FvsVxDHTMaKPul5v4OpgfSe7mY//NL/ux2CgnkiBAe
ne6YhKPBDnhoFL4FV/q62LtIFt7jtfeFP2yrqEncoGjypZtS3veVMgQy4JoYuEZl0KF7TrU9DRjj
kMapV/rocFjsPGKOY/Inne44aBCwOBzfF2KUHBDr6P9LdRekgenGZ8ae+Rl5Ys6mRWy6Jn5lsvUH
N+Qg6PvHFicXrSm90p6GQ9UerXkq1q4Lt7CzyKC6tusvOwmxKtrULOw4SAuZGHA7Wfx2JQIPqlvH
Z2SIzfGXLk5GCJug9/kHD2jmDT5PGnMkPO+oWDZJ7ZRsMrpDgS5yYFytNO+TmJFZm1Cn0W/SUNjn
WUZCxse6eLZixKei7Fudy94FpX0incuKKP3+T8cUjtCn82+dNxUvYq/fSxnXTcm/pzkd2kzQM7Gx
Eqe4KrhsvgdBkU6Uuxr1PJwaYeMOfFRN8b4yd+X5jRAbE+IOGmx0GVUIDroOA+KNMlPLeMtGHIWx
5qnMmrQQ1pQSd9g1ZP5kzR+xiVboxbO5p6NSaVG6hgaqavsYJgIlewn87JyNhFRZaz65lTdj94rw
NVOqSuZzJp2Y5eDHcnBt9RL6W7KkjBQD9S+hewmFjp0BsVM5WHAkN2ymrOPqVbFb59/YtkI2iGRw
tqJuAkxTJ6d7YZhhI2QeMuUUXZIn8JlkY05A4kN+1I6+k5RfTs/utX5JtH8IJ93O1ycFa/2ipkwB
wSVv8s0xzJvH1Xhf58dJteppqTuTYOOcuwNgSvkuhwR5ToIBiICabQqs9rWpjOKX/YiOD0gHnIXV
3fnICN1Gk6i5Rxf9vdEx9mptc0HZDbM/fHPOxmg6kRJebEqYydvC1Zz4a2U4G2SLhjvxv0CUUVy3
U3+ndwiF1XvKjf52sRvIrt1ArcNmk/Avj6Ua+n/TmrQtF+WLS1ExfVSJk4MrbOyrlNX/w/aOdxgv
nYagjlh0FTFd42vIQ1e5BcTqBknUzU/4L00dgcrTtD4jU7zOT6lQ+JPzsUpI0Da2RYkPS2CP7Syt
LDqCbE9Byl11XLHDLZJ3Diys8t34zNeCfz572SBkf7/7rSw6uWhEguECnVzq6MdRpIsNKcKd7M8K
qhQFIDvvIopqWx18bd9lBSXSoDjyeO1lWrT3XnsDvzY9zXasFDgrYTGsHRgKpStC67CVLUyjbUhb
L2XC5m/bzyf0TpF3ouA/vV8wxuDlppo6wzGjzU8SZmPMgREjQPyIOV2ITM1qHoA4DkFHeDnE3iIh
Y3aaGm6s5JOb7PPMb6E+hYPL/SzlrvGyj3ZAFClNEzpQA8vF4vNBqh1mRhvaSXaFXrRO2Zvaj0XW
h91yXgjALg46427EzegRU+bSTAr/7jPMTGVEJdQ4m9/dk/Bf9LmWXR0Gkgl7LOamNvODVs/7beuI
HT3zTy6fbQWP4YSSjBkEKwggOxNyhhqXRXf/ASbwzEHJAlOYwRdolx38bw0ZuhoqH4N1GCNcokUU
d3T9j4IeDfZ6uLqPGzHPZaKZEYVcIn9CDwJl5KIBbzIL6CWecYvB+GYKVYOK0ba/DG58JSk+mvsk
CMWIR7HIaBXD3nMoSW7naxpxznfS30/l16XSfQPUbjQyYtqryuB9IJ3J97hO7yN3O+NeQchucxoL
Nm5Vn7aJxzEprAsARO/6r3dIYA0DU1/0Uc4lyup1F4MXslTz9ZDxGzMa0CKpWJmC+o5nxNWVc6tb
/sMkmL0wAK7EXmswkk4gaPuEkzo1MCW8YcdnE1qjBKo0k46UmhmSh/wXgTqd6SYysZisbkwQZHWS
jCOTbZ3UdrBioV/RBKQ0Ipjlv3ag4NKxCtLxBYlFJgyIv657DJhyL5/7DRc78jcvm0ttehODp6lr
I9Kwvtn4jcl5Yf0ggJ2git9sx3r4vlmoWXjWcZAmP/LtIyTRgf8K9NhcnCqMV5GOa9GwzNaSwkwF
coMJKoM1ucTTcXBO6gI74EEdYnrGHjfGn/0iGt8vvylHm6+1cR3uTXcmnBDnvUd4sbgX6vvtbaaG
XvxVygOTBoif3GZ9TeErlA9tTjO7EmJ8ETfk9pLTR5C0sDxqDsD4h/sbfXBPr/TB6+QUoRR9cUu7
Sg6P3K+jRldwEiM9q+5r1Uj4AHRtO5x5asTIbzzNXYnkxSLsoPnsEbTWKAgpPuuyLRsPmpiPQixp
z0AKvMme6NNdd9bnPkwbcf4Ca51iQB8pUdlS/0oURd53bboZTYqoJY+X4g+ClaMBc7npllei+i/D
kXMD4aOid0HmmFFpE/t4iIoVfdP/jM+eSricacmjGSRVsNhNKgYj1+NM89zY1dG9y32wTY9oJIeW
A7QdhO9gmYOx4mLjMyUH6YBrdXiW2ZtdPXEwgOITF9J5YeE365+vT9GiI6YJgoEr4N1rPZnStlFk
RnQYyiGg8EX76tYqUuCVsPaoHe9JiN6KpL1fnm9HDeaWk+N9I9qBU0eCmSRWKwT5CTpgy3SUx/cV
qDoWGzHFUXtEOsXpsWXrCD3CbPUAd15pRxXtFCsRgVo3XeJDKpo+zhq7t6eEOruDPEmSFffPs/zW
ir8CyS+jwMlyc1gFBRhvk3GVWeG311rP1SfrR23cQnjrxA15f7wvsvwUE3T50FJuyNmldl3/6a6F
93RkO3X4akCKuBXZF4IA4BUMOwlMLjhKEruoTQL4dUIU6b61eXLXzgkSLe/VF7AX1MA6QL8nhPAX
1n4NGTIL5VDUyojc5D+cJwnCLE87LkWd730D44PV6ayKQQ2CjRM/iSs80O0GJSo1IGl17l0fhnDp
rGOT22Rphh7xB2eqG7dnbO8rKzHzNDOACYcRIGFEfVWtdfjKdsI2Rwlw4xCfjI2dv+6bOyXPCgFR
VQ7IenccszCNM02JySNJyW+cAk9JKYAaHMe3tOoEHrkbRqc5uMqchAIHIs4hSQa0Lbdun3WIO3ZG
bUxyEzGzpRl6eEICKpSgPhMgqYrGnjCBkuTEn/mOLXZtS+azQndxmzoTQKP7mMU4GREFezuNI1Tm
ZzX5NwSq3wLOOUCHk0hjPW+UdnhpeEcDGfvqipyGeq6podDXynWJo/CnbhR0AASWYHSbP1s95qvA
8nugrxOo6RiUBqYWtZ6W9YTDlJstClNJ6Ne9LvXIJ6EIWvFOR033JnnTcVQ4Jin0CUQ0W0xiqDVP
xOMkVaBwSWp5H/U9oQEusFk2pWPbrtAnptWiaJttzgN6Z3D3l0vzpyzSxa2EJqiiqJ1UhggdGnIf
VCADbtbrPu6YqsSkKoBxUEekCCRWdeUZB7q8K0Ev5ETjaVLiFpehupRM7xIw8RGl/fOttQ1PJ8Kb
jP2z+o/lGlb6Qhe+gR0j7++vPQV/XqgPozeYVK/0NodKzZwVBA8ucaomftX+UfA/06fcfL3wf64R
XG3F1zSfWMtkuf7PxFQheS9/HHswk4OC2WspToCIK3jGxdivRjaMI2o1Sk/MX1o6zCbxy7lVxGAY
uHzmV35RB8pw6OmVxLkThhAxqpEGW2Svbu+4GbZRiXJpwW9f/CygetOlr+5vBpBXj5n02Z0gZiGI
sV97tvGsduojVk/UCDB2yxp58HOnWgga/P2vajquvtlcIiEyXOcVkaIwIF9XPavldPgr7+3GlGUa
5BYi/j3dBqTP3YLn3czpMFUx7nItzXJ97+lJMtqTc7ou/bx6MsAdyOSOuAOCK1G2o63Ew7D3CkZ6
o+6WlzWBWPjfrS5ESCrdBlRoxre8Z721wiOVWuFTMP5ROMpUFvfhaa30ZSpgfNtow0PMwZn4obMt
Kmyw6r9QhukQ4aQEYcB0DId4dstbIvvQKxKLD3vSRHWQePdsXxZDIxqMr+uJwJ7KQ0sswZs2fF7M
YdoMiDF7vb25xYPlzMgJNGKvULQ7CsTy6cLBgGODEkwSWYwaCAxCu1Rnmt1fdwuN+jZ8oh2zv453
enNd3m0UllZ223u4jClRSYd28Qyv7uJGmr84bCZSy1okb3pVhAuBF1olKxhaW+Q0INs2snjR93O+
aoWUFSEmKdAq4QTtMEuGGNqobvIibpJfii2+SHWt73+g+uVUHc8RyRKHO0Gis8ePx+yVwm40syUs
ylYZpeZsgGoRbG53/ZyPml8yAcB8z/5ut4l0qTGVXqLcJr7DeDnltfB1jUzq0Wxz67gRRc8LjXNc
kFGnGFlimSNCk/q/E5bMt6lg7Sku9L9GIp9qfb9mj2fcMH73V2h91SKbfqC7WrbX0MR/5Z4e8fXJ
JKpI2slKB6WUEeo3DW9KXvJBO8sCUoa5Ft1aV3l6z2wwnjeKTu+LE+Knk0ynJC4mWrWfR9AeFz3x
RmtwhUqlbAHN6JFYDuHxkBJ02cTCIH+ORGFMkN5QwzParMeuq/In+nj4dCBH1ZuJIHQsSXPHggJ4
QyBrXzRYTvIEzCPLVUmIr2PyMVAnR3w3UQg5aZOu44e8pl9AxPEXCCeq90sD6IM4LafpeBxi0aJR
dQCWA+4uAOcUDztgNVyLHRdNLGO5CXvZmwF67FvT55fLps3baUEo9kqWD32bk6wJLoGrFazdEjXw
MjEeZQGn2nP33SmDF2GSC9eXGS9Y0YXAFjyIZGu82u6TRqkE/dwu+hM1ohAefbpAJ9xbqYiAiaW1
bj3qLTSvPOvQYd4by1k/cjtZyipgkwUmr/ijReanAeZG1qMR57h++CAoRVb8qMF8D+/7IVPrZrfb
AuNNjzB6gIvM/WFnhDZVY3av8e3zzfH4pokdZIyzqog65Fuf/oAx4mCc1M4xa6++NYCGo1T4InR8
IxdoYx7i30x+wPLTddW4/hz1M0tTpvlzr/Zvj17ZtutXDcN9/y6UMmdt5FjDWKDqd5o/lG9piqrB
5TzBvjDZRpshwytlUwv8FgCHTTOcO1W9F9VIYOEPL7TSPrEmgHn5/bJsZOHPk98/lg8Z9c4ZltX+
62f/JoFFV7bvdxwBixrYqp18GSCrn+e+FhptdzsXC2h7U63MCuJ1VzkbV8/UMyojWUsRsmJjknQE
Q/kW82Oh978ltDSk3pWmY0E5wPBT2D+gCQ56KP6QEIO+lrMk0gvgk1aTc5A3U4jtKVypVDHaE3qJ
mgBQzvc1TS+3LiBFPkxuoE+hwf0wERiPxzEMt3900ypzOIpOcFsva4+NnzyuKvadujBSz5Vr1MQY
II1TPxCAl5HWJmEz0vPGPDAvNIRAnyDqOdUAdVaPtXZn2WYkt1LxK3o0yT6RU1biGI9GGVC3ZkHS
pfD5OXypywZUG4Zk4azEkZFOOYg8Pom6R2KZFjTHk1VyPGmIihYeQE1VMSGaYXjOOEfS4Uw0L0xP
FjEfzf1XDl4KvL8qMT+Ufc/jd6BvQWI4dIfi2f+/RM8BiVpvHqkBNt9TAmiORvHiM6lzUCc1aYRU
WbhXH7oMI6RexobJNWNHhvKlBS0u9JRkkodptXDLEVoJSgr74VdPta7SPvLYxMLr8AH3JCeOMDxn
9GhT9PajaxwY+RwT1oI0nq9XWDdInDH0X6ao+PDzjv8vqgPG8MpgQFNMHWtUjTjdcOyF3y6OguAg
LQ72QXpOQZTgmeoMzpAJ9p99pHH97n60jF26CDkppICnZKHwiy2Wz9fKke97vzrBTFhbOy08LQcC
DVaeY6rL9UeDwi8CcncIkh8EMhxryZMx1w3moa6yDzfX+xiJEQQgR3MnItAFOxmOKDZqnKX/NRbE
hFpfSpHNW7oSvxz3K4v1qJq9J9wAYoeC0DJhsyU/RvroRYk7AA6YtZnbi5BpbyQLe2jQaAc3eRNc
tbxy9FW2EOdXzXOpea/ddER/rzb23pqqcLgPyxbIkqkAChJqeAPxz5gVieGCN09CuuzWKSJJO7u8
3PESpoKCZwIvXaIJ35G+qbElFKg1wMIromTcgSICAI14J1aLNFSUbAD5v0HguvG9rR8FUcROqA1q
V5QYL7+7JJEFtVQafPdnyC6/CjjB2tRltLNaf65VZoPJ9aCMVt72KYhDB2imDyra+p3Bfe1qy1gP
j5/UpW0DSqqcSzREydjh7rohSonVJUXB9upf85CqDDV0l7W29O85WyNtDL5x/oglCEibpXY7si5e
OmjYfkdlgsEsxEXlT1Sa7uQnKfUOJ8bxKmXwaAcHhqrzaiD7tqhCTJqwsknPBiqElskqeFEJXn2T
ykmjFx9OXfWzlv9Vk1xeNwD1HiTM8MrRP1I6VkaCrZTlpfRY5OnDpjc07tMq2ytTGsqLICnzpd0k
iGnj8IaIyKpks6Xbu7uY4sPQT7XQ7O29UrJ7k0OhcuEqA+OfMk6pLJF9FjGacc6SQCcg+JaCZfoG
BQyafSai3e+EqhQSQt5dGcDK4nPrS1DOPTSBhvaG5Lj2N9HQU8uLJ/VOhfp4nNTVWtF+I9H7HGkq
qHBY7jmu+ATlIElnjEdWYg0eLjj3KTe3CmmL8UhqkPmcR0+O9yY0FqCAwxuNtfrEt+aaMa+4avYg
OOVgN10Wv9xe8xbGYtFu7fRgFeec8UkWPL8CDq4PKpmx1byeLgvHrzZKK3CfG9c8zVAvGxt6pEma
dLRH0CxnW7zO91LgJmnebmxHOx92U+kjpjMYpzCpbohf4oy/478lRDyQ82dqFcShGzvjSRoSOryh
hObpu6wa4nNwxbV+h8AHxOoVqeQQLrgUbWA+EHbs49H7ewjaGClH6JH/vYANwUyO9jjPejZHvK6U
uJbYWvpOizlGhXeUQageN2CvxMyWgcqjXJPEOyyMpYmpg3W0Tt5JiDIhidgDCEEVSU5UDo9LQfIP
HYOf+Srq3jaf8pmqVSpq8E+eZYvvOYN0kRyH5nsY2eA9gaS96g1URkmERb5wpUOpN8saoJwCe78G
SMs0Yc5gfXsUDbnmPqnOwMRnqRNdDuCUw7We5Z5uowrCCKLPHAo5Ucel3LmDAi/QUP8NG9PGghY6
wQa6TQTGzHdeNdpTGq58borcVcekM/BGRDBtsyqsh5eXvnEhBHzkEjjmaIqd6XABz5jezAQzKTBM
lGXSBwVvrEDy+KfDSLIDwtQgvdfALU6JB3geP4dFu5FhKM5r/KW/17ThPFidBIVG0ssDDPI4yKiN
ihH6cEaPdU+QJcIFMd/SniPFHOQa+RasmVY9m/D27ntou2XxCV3Os63uEBOpBbq+C5kNLIZTZ0oM
VA2v3/OTm9UiGSUwR18zhTsfi1shnp5RS8RisoH3PkpzTXLzLZ/1hzRmY5VrFJVFfDwySGnqWvZB
GT0H5fpkrSGOIXP3xW+hJhmGtS/XxKG5yTdtL+fNqIBk9+zRR7OjogwyJkLU+udN7JQlFyeB+y1R
QoCW51UTqeZh6q90Ldi3otF7ZVx05kZNvNr7oUxBUVKahp0Cmg+UmdRb/ymx3I5MjaUwS76J2neh
SbvxkDuA1V0H1bCTCvMcnPwGa6tvxWvD7KwZztiHVXnYMzaSNbc3QgfX3XS4NqGjOylfwI1Tj7RQ
knJi2St9BFxBKNbYzoPmnRdYNgbR0Utj40us9yc5npDD8pLaHJu0AG6SKm22m/92ovXWq35D2t78
1qpDBd/dDt0QyFbX0tP7LfxrAqid8yzk50zz1EvUX7JWG/d7KfTIb2NPYqd/XwwLi+nul+1Tv+Zj
FvZci74EnRKFlM6gJ3NqFfe6hLo1Q6PvR8SdS0SQKNDeXimIKlq4VFULTG67HGJ4u0mvNBPZhcG4
NGmySZUh3b2O1dSrUoZW6g8zfB6nsDYmPlY5dfTUnITDZyhoU8AyObMhH1KiilDxJB6SkuQs3ruM
9dY47cwMJ2eeNdCvBzglJn89+n/zq9szpC42wGR5qkSe9gvnfEo8ltVVHQ2X3QVlhsnzdHymraEh
5UYh3egDqQI74sf6/YG0YvIUa6M8IoImednLmXmJOAQTRFcVzo/5cYNZkMxx9XR0pDHdagJ+vfde
eYg2rlHAjjfrzMCRLPX9cacItHhiKcOES8mzpRHWbVcwJTp+PWa3R2sbV4rIPl9nU1DVy5l6QQgm
AdoBM7yIpGBueCHBajmF2Tvr+ChxqtjFZPalZjGdJH2mtG4YnbVOj/ik5MTpl+AI4W96gMie0YFH
s1gAM4kn9IoijyU8awKtL6x3NS7tisSPdU/WH6KUXTiYx5JPt2bYob6MdW3kD0ysyKnYDU2kWZ7n
kW5+36ZSCgEP3GR+Dpe1H8txGGibl7kDXFGatnV+aRSgDMtHicImgdFeKO9Vd14EWqjJ72lZ/SH4
A6k2lkRh2DVY/B5yEfPJk0aCGngEujJp8hcGWzn7h2M9FfdSxKbI/1tfWfupLWOhXQ4XUTM5AJbN
Cgw07yE1P3UnRZVOFUeioMmvSGGmyC6vh+axAKA7y82CcRQHg5a2TnumOMCOHykffJn3RZcJGwhw
r0UI40LT/VGSi0RzI4g0HBby3sq96qyEIRE6L9DG7YuXEHM7yKu/kw3WRTAxQjEIDgpQkn2QNVMS
sm17ouiSZI0zvzdDUiLAguRZwLUDwmh4ir19HwAeBnFVr5jYt9b8asfVSE2v48MTZ2XZl1v4FxFk
5563cSAyt8dXzDqtjrYImRAjT+w+EGpXVn0H/HQiD0OcYr6cabvX/zapHzyDYKeumrD600rE0jtI
4r2d58TYTj+wGYCdZyuq5WFdocp2siUfotR0Q2n6gmguBYWxNyzwYbLw96hlhzJGx+yaPH3/phVI
ENN861M1yda/5zb2xeZsTBe9vqWI7ykUSIaqFAWg5u7oYFeYkJSuxTMthk8NDorCs0mV6+UaMGOn
5DrWfcsWJIATFfcCVaV6cc9fB94j40A2aXFiq/zvNY5NWMfG0o9y0aBMeboYivrnwUHYZyZKgMuX
CTAKo5SO0SKHPOTBWVdkg7ABmm4inTc9eXzXTDZxy7ah65abfPjTdwalQdzL6agmzuak3vMKf3bH
xpGhCr0IVryMTO05VqJuXsTEYza7sBcZznmn7df1rtLBFna87hPL8ep2wRsCWqC44OGmd2IE4TO1
mZBFaFKcf5G41Mnxg6ZfHYHA7r7b1chz5LxWTyhR5gvC/mEf8Uic/EN9HPjH7R2HrigAaKvUTMVH
pp14DzFrRKv776IGqpkZv4uQGxsnPK4enoAdSSIm5CobQaUBcmwlgDvvAf6FaVEVJiGu7edHs9XI
lC28zozQELBDkqp+C9i1a89m/AkKXnKrdaMQ4ZMSwCOTpF/uEC7ysGrei77HZL20GF+/ZZhW6Yvy
vj6Xg8I96uig31Nv2tMZHRVYbY4Nv6cpzvhooulyEUiDWc2bHHMm8dlFaZORqEJRN8QRnBbQIwEq
VfH/9i3s1DN9KuSuq5cirBMI4GcK0cSWGhQbsOzoTEXpXObc4u5QI0V29F6Tuwv3Kyl1Tj4UALvt
gVb0cNHW+zUgL3eLc87eXZvwdUJ0EkqfZcUmny3j5wPaj5lYwz8kn2OGMpw7fSt6080cX8ptmGIh
3/UqVUCzGKH8PMu7pJH8vHzJ5XuG5MuSqw6MPSj05xNhsRBC72AHiz/AYudL03GppCUsAGCNvArH
Y6rRlQN2l8wHCcasV4CHAKMWgh3UHE7KnR+i2CvXqhGYEtAA4LvD2R79YlqHyqxUeAw9Fu3A2DRy
IgwrgFRIpabqDU0L8LsGXXPLk8vSEFXPE8waWc+cB9XJL+sUxoPelxyOYOdc1Wih4Ivq+Y2Q1izo
QHFdlyD+VdseTbZGtMzHeNlLaHtpFguHdUGVmMIppVBLeR/AeVPk1ss7xnMulS/Jc6/pykkxYhii
N4vNpI0Ziqqg7kwLv9GnjblRWX4KzkCSnZfKt1F+IHNcVUvZbDGwRFrRgOMkM5/A73lC/4yoX56U
Ur0heKzIPtlWtCtilvsSzLDHMu7/QOwgXDVnOPOSkpqnR3QfszUImLdBJCfSiY9G2X2emsS5K95U
Yr4GI2jQtUZdY98Ab/wT52q4Lg80uEzHKRYDGBXte9r+A39YTqAV/Vz4nWllS1X7QsXAYwkRym1+
djKZ4sETUbV4rUIkM4+87HX3FcD6eOPZxaOD6sVTXaBNQ1ExgwtSFhMKbwvIowHA7XmwIDjbsLCj
NmhKeV1//6/IFcka9eyFaToVFzI4oiorgT7bXRk1uDve3YL7G9IRzPA7yigwG1APu9juVxrk1fMT
LGQHmFUSfoQyUiTi8JUhj8aaqJ/zVFKz2P2QChS91DvGjLp4qh94oioLl61TV0NFFKXF3jzU7r8P
YEcHc+ZRk+1CpYgeicDYvJLUGaDelFsQz6YosQGElXHXYVqx5GbpnXeoCW9os0dDBO7bIoXMpTqK
0pbqFsgzCS9l0OFw5/LRNDBevxDQhEjc/Wz+ObPXylWd8DMdc8SRCUIKIKho1SkNi/aZSdeaCjVq
ke9nRP9i5i0efYaax31YIglcqCPq/LMJQOxWhG1UT0Ma4d5xLbJgg4tlafPBYg3h3X47XgAh70jP
Ij1d6j4vnKMJpVJg6/9VcdvQaanDKHu9cqLW3ftnxkVHeD1qm3FnI5mOhGptZQtFY27nngTTW9Tn
spRHpTMvgoVn7DA6e3xxoc83MNOGp9eeSej7B8hI52EVYZ2N5NsQwcm6KazE87tJr5I+wqH8wLCp
VxIV3cFfQ8epQL67BX36fGXSWZyjOmGYNlFY6uL5gshwwKYNaSvuUQhZl/XAfBia9KJkHtOcndRi
7qketFu828daV2/kw/FfH1yzZ1tCGAQBewQYvQcVQgBBGMg95ZEqRh/RNIh6DyJ5ls2zYiQp6IgG
Ju0f/E+a1D70FVcEELJsND/5EcU16MwTuhShE5EaC7iPe3En3ljmJUCWESYhltln4QGJgxV78Pfb
hAABqqExTrPap2Hf9CWzkhg/eOA2UgE9Ll7qNn4ghmFtosLEJwVLZvWSrT/ZJWazym30B4AHS3Lk
ynvrgmHb9hdqA2QuKeeEY/bLAtNS769hZSM7/AV5jXbZHdvMcklQ2svSoe27HpFfZjSa/OxxWq7c
NtZUc3fnNuyFQEMA60ICWL9SrO0gTEles8LuRF0F6C1uAVitXUaTSuO/mK4YkiDtF14k7dtfqppt
yPnmPmsMBUjfNL8pgFvoDeVQet3LiHB3xi/boZwJcWeCiYo2114wjQTAccSMRVcZsDLunzqMk0pk
+UGYUl/0s8DCL9VYzC41R8VPZS/74JpL+k3g8ipNcFaY5oLcAuJS5oJaZiNGDSv1bPDZl5Et26+p
eLCwb723jeC6BPOSf14CFYRzmvSQAOf/uJ9VbXXKMVhTO6EhgIUvoGJgnGAzg7jfihPxT87Z2TeL
Zxke4duWdgqvnPQaA+E6mZJQEiBsVgcGsWIu3uFToM6X7+ufaxUFeNu/h5t5tMKIfF6zCa061K8j
XG89elkAsqjpWaiasZk8hTX6shEXm5eHjGirafY+hy/+IqCe0n3Ox0owHeeVID6HG+JdCcpk0njV
dHM5hpYZQXVHliI7tLOHMX00hn+vO8qWmWLzhnYBejcio7Pp0T09sRQRLKdgb6dAE29f2QBX70W2
gpfMHHgiEaZoPxlaiVkJGAQPFebit2AmEP6vziJgrmq1laZKXBGqwXppzPRlkvuJg23Kl/vIZw3i
ipKUQESxQDjhZh/QpClrBZRds2naAsrpMvGmm/kiUnqokiceYcu8tVaTLUNwu2lmDouzyTVtIYt/
5wxFisgirRQpNaj/JPoWJoaOKRqpI1wOpMb+xIZoZGrIvBUfJ5mfc7NCQA9uZ9tIc134kVwt9cBR
zPYs4u7e5SdPN3Id14G2FPFmZ8FzJVQdtkHc/OiGgfJAJ+tgrkhTypcgAUX2erleLxqwPqLUR5fU
BdrrrO1GB5j/CLy6epj+BFw8al+g+j+J2fUyMKKdqAMtm87pycdp7jYRj0JeT4PSmQ19rv63ECDd
VkSKMa16bGYySBsKlan9jhd97wbW1rsf2X9d68rGToPlestjwpJjgfuWfGcoqxNmZ9C0w15+GsdU
BWPUBncLrX+AAKuk/8bFx3pcpqhXB8GmCXmSVKkFqe5s+nto2J62vOQDqnz2k6PC/fxshTMchHVv
xSOriK8vxfoJyOy8ZZ0bSlHjWAFrP0qzyxuOWxzlpPX8kJcw2LJJ1vyct4TidUl3JmEyiiQHu92P
nt+rXYhxi3Qsob5KxvgsXMRlHV9nGyXTe7aNmJ+FPxDBUBABeUAF0BTciRzNPWiffC9NDYFLed7v
T7k3FhxUND2s42JUDwm24szffT2pEwZGOd6z0lzI4flMIwzvXqba5daAv/kZfsg96C9UPDKs7Ssa
3M/L8JgDb/efz5DR2k5QCv2BRkl+dgPoM+MZKjKhdz6LqWeoNRwA4BVK0+dRllYuHS7WCz00HqHa
tL9GRVTgVU3XUo1cXZKx25n2l8w0qoOKW5p/UEZW7kJx5SMWnRqRBYnshvQl8m5UNjZ3U60N7BhH
NktnOt2Qd7glL544ydplF8Iwndt/O9afKKWvhEbWazdgR9OY3C2ZnuHhGpC9ouUgtgO+hTk7d0LV
uPQC4zeeGW3fumhlPB/CXaPyAAOB4qGqYJmNTPTf56ZsH22Pyv0kxttgu7+0WOEoWLWXyn1Lukdw
RTty9jFuFqwpJiUjr9xEd0KMx732ugE+8BXuArm8cwDlhtKvRTMp5gmKVUNsmwB34rPHS6Ndffgb
kIASxVcbhiV+gFpGqWLacDXke2VeizEzdQaMngiPNBN/2v21vJ2dvnvHw6O/sy4XMUNc1of3TQG9
RLBDGAEKJdPEePvFSiy8nwdnNexMGla51JDtaoHWBi0G2v7C8gBlL/VVrRPHjoEoyRu2jVfLpXN2
45oslP4Eb1ghKpcoKVY/N3+bU+lkAibmCxZBkdx2I0uVEnlM4SUC6Dn5+3RTBKXjmyhUeRUCC7Lw
UZ8N9r7DlLP4UfCiQZowJIwrfXoW6HrhftbcIIdaZrD6O0Kkbp0USzCAcyidmeLafnUsf9C/HNB5
ORkthYANEQuVW9pYLqrp54binsAbzzWTssmMCwG4ge/VA7c1FCgqaZrhoEPZJxHq+AH+Tvt6GxLZ
8wGBYwWc36LTITNRuatKS6lFHRmJil4IRIErWMxTzseetQM36BaCYvyZQowMFlJBj3Ep6bTzjBbX
wV3bdI0TjU+X7hKbSyj93XCNn0o7oEwnCMA3h9GxPRBEfeJu4ixaMu4AZ0UvNzYtXZyFEx3JN6Aq
5fvBbIzw/zZWVh0/90hCB/Phmvhq68MJGPnk6GqNK02IfBXTD48oCif6SN2ymqW+rCCGCCs1iFgN
PjnLuCXLHRrFoEIw0Qpg1quXkS1/p4MTdX/umz02694HR5Ijype3JlUdukW97zBPUNseMSffSDwH
/qW6EWL7zlyagucvjq++JmMYu3eSN1VcDZtWg29UgnGX62FV7YzvOcZ5vagVgIl8WzxwgUN3UPBP
gsIpIcyqP/TPw5uGYzppTUl3PTKAHrG6ha9i/yWjGdXTCD5yjfSmscZ71oHOgeg2kvwsEhJv79Vu
eP9Ub4NFoWwTjywi/fDwMvYRqN0WOD6x0fAdkjvSTXQzyjzp3pLN/KSXfzqW8K58DndyX47Kd5FC
H4h72UtkNQWTrZqdeKUKbovJg7MolJaOLqppKXZm4BaHqx34QT7p6B5vYth+j+PSGN2kYqihLiWj
ZoSMRlthxtxjRaG9oQqHilmRoRdmdM+BqizUcrwwvWgH4b8gDw0oQDjRnvS7tVm0E08IypSnrR/w
XvcjsspZr7eVKnxNil9pR+KMK1pGcIA9SS4QzSUcv9Tc2owFPmC1W1ozc3HXgJBtGRSTGr/7A1H4
AUkg1h50tR9jjPt4Lbg1dS54vqhn/6gRMBePbaWydeXqiy4JU8dX09wZopBvAzYbrAF0T1dUAQ04
z4+UJF7hFy9G37CXC68e2reZDMlSut6+RmYdFMFuG9ZueJMCaKLH9fOQgHCsXrV09S+Fna6hu77w
3MHA8j9PoU9kLmGwY7YMvAT2U3XASnfcHQSG3MZEsBIp9mcG/k2295xOLGHjGEI3xqCRLhL5+YCE
kJvPl0iyT64txarOWytsQLzYcd2j4l1TwZ2hffljJbMQXmEpKkeUrTZvAvjZITsAGp2pQ6Aqqe4M
GFGezTFksrK8ssNL36AgdJFKF0zE38hPd2/G6SGP3/yoD3LCtvenLesbGXByHxUU3w4k3JbTYhAD
n89Q0OVIbAG7jAlSatp5yPjgtLlxfBtflA4me8/SMH8q9CVCVGcPOIreguUog6Z8LRnFh9KbWnzx
8MQaXv2QfrRuQZgRyKMkoHscsGG5YtFGbTbusDnW+M6Mv+0xUDdVz6xZwtbsbpdAf0l7IujjPnbk
L+TugBonRix4E2kXMq5baWGOOTza+QRb8nMZJvjK2uEgphzDZqMg5iNCAkyxCySDHIAd+p3kvkH5
us2uxZaZ2dsBOO8GBVQzQgbR9jrNtyNTrAlgWqGcydDrnGtY/TyGYLe1x9OnSqYrldWHzypd2A6v
Jti5IdlP+zD2Og4RAJy9QtJOOrXtc585zCjfNuaRZqC/hGSzXrBTy5StdE5185MhGYV/2tf9XQj7
5FU3BIS4hKY99mp8tktuRxOPcsM2GMhTyeIl2Custfurx6rZFesrfaRX++i4LVtvnhCM6Oye/tst
oWOz8Z1PVAmFtm3YXFlhhhCnxm9J5IgQcawGsD3vPUd6/BlqFecxwWioB/mJQ2+WqWiyHFaBaUWt
bEhBlgZk0ow79o8rf/U350AMUTLW0yOfwWygK5MtUrU04fRA7ObBG5lcgt7YcMWgyCwzPsPbubdJ
LEyR1XFhOdthGHd6pYZRv4D4AZTX/B5yY4zroRVrycvtglLhgLP1D3TGJ8vp8nyrALhUI5mbEcPJ
CWUadeeTjyMlRy24quiDMVm7+mFPwlJBmQRtUN2jr0vn45QEP6VNxej3VsBMuurxgScfuLBo+xRh
dewrPwmyg9CZXxrvSopBb4bPs79PJ0cA/Azc+LjamWsLm33pxrTJM8yzjgyMZztzk+xMHA5uDeuH
o0/AvL2vRmBIkWgOo2kSAEDoFZJeOno3d1C/U3IqoLJCPlCnFuUifsOHFejcyObL1Z8CYsVIttph
VZ9mMIDh3nKpfaNhTSRMmKX1Vb31vI7LF0f3C3qD01JPwvCBPQPOGWhGY1LYSs8XuUszWOd1iGAn
lo9OtjHffkUwvdmUvIC+IBZ1KH3S7lSbXkxxpjdbjLjAQIMnEnsQPrnMmFJmiC7azj9+aANxR7p2
h7+iyZcP56zm9cm4+fg2PQXMQ644Ie/7ht5hGYzwGlO/Gs0TWcVu2LMpYP7jN/GqBD7u5uVrVt3g
OuBwyt/jsVXmH31vLu3MQepPItqSPdCUZ9PdmWY//7nTZ0VraicXvy6zBOariewt/0P8rsjJ35qM
mBTnknq7Goa7W3/38FOatbRR0jfjZCrI5LhidZznPSaLSIxZ9v5dEx/1BFXq4Z1G1mNwGP8NsAU1
boglP7kC/luzuG4YAbsLpVAgJLV08NszEWzQKfOxHdPrgpFA0WRSmgH7/4PG1DozogJwnYRhYdmE
fLtTlWl7vQIlkV/xW2Xh6Ue6Z7K55psNlc0E/JqbNcW03NmM5+xvT/ih9T6e26iJSYZ6lCsG/bs/
4IkiuYlrAa6LpoOQsCBdM744NildyrJv7nrHB+985oLjl0uDJawAHniypIW1U7admZ0vWVlR8t7Q
CEwTE+nqbAlFPBAtOBy8BSS1HQRKoNNGN6msBTzCOmbqzMJ887F3qS6v3b56xZRA8BpWpbIE7N00
6RDIQRrqIbJxEwr67vQJ8NNUGkRt8Ozw847DYjCfb7CfFq8BkmUjZ2fxoBPVdyHgJ90rGLvrBiSc
s0bsQldzdPAe9r+kj4IRPeGdqlOkIi1SOeYfdZYpqYw4+tHYGSjWDTdUxvJnwN2/LU2cCDEDwIMW
6QlSIL+cY04VUojdwUD43Z3wZd1iAOMLPi+L/SVOc2+SM7pYhn1uw8m82nngbtRCVmTcuT/nw92C
auC2ei5MrPHpPFLJg9m67UvKvciuVF0kV8SYC89L2ETMHo8mpI7xEz2kNYR/ekoJBbl/WnTGhvkJ
wMwjCRSWzDAugZgpw1nZ8731+S8m94inFsf6PmOZSOmLk4ALsKo4Uj+s9s9iCFuXbaaTbZWvm3d/
5waOq2WvGOHUcBIdhzwKt5s3hF2QK2eDZwtQpAN7vC9pyrpqTwzSvB1qAHu8tsmSPZwiXUmF62B9
IKbUb2nhX282KS11kgEJ5E5Dh1Gfrv7j0c6K2f4dufvOr4JrXhI13mbSOogZ+r8ak79qLxC+SmZj
n4E27eijfim+z+jGdwBUGb6IAbFzo8ybcnHDrxHbRSqW8jcYoP1XlAGYWlDNiy2MGgJdgd0CmQNE
Rzyrv1+rg4koUVK5wsHW7kdAJsgDxhH6lRfkYX4U5EOFccTdWv/1YloHsmPdmafqYuhTi0+oBqhS
b72oQY1xQFHd+cX2F5i3cfTOJw4WMGiowyGqKCHbuWrZeOnEq4fLiMHbWFCHq/2tuOhnhd9FaYg0
jhslaUr43VffOYC5TgCZNz8ojW4KyNJzPyIB8K7mCmOrbGNBv47sFRyCxebo0pyTNV25l9tVfHIO
SrsDxdkA98jRdL9kMsJiLZx9/Jek9EHhGRqnXU3KaRfVBAs4SD+/DcHnm3hBnICM8R8RqnCHkULB
1N0Vd9ZLgBwIFZzE24ezgK/n1lsL3nOBLZqNip0jAbd4TdbO0/VxuTfp9T4Q+9ZKixendBbmsrQG
emFu8jfokD+TxZlbukLxNMNCdZ7xU5q9ZXt4WsPPdbtlC+79iDBApSdjIevp3PPmv/UjPp1jxqJT
8M755W5CglZtEB1nLUAV8Y7hQ0994k/FWO0dTwkn0r4PqOdc3H77/6HeVLWZBzq3Jc+04QLpd5H0
sUqEdDgWVOdpqAOVJVCMyaqkSsMdeds+DTBJRF91Mb6TXlEptmGdPRup9kg3zbUl6K1XxC7WvmEE
g/6664GHddkkGR9E1jRYdAeAZfLTi9bKHnGIrnC/ktVyd0/Cx+r7EHKFShM6sUmjx25Pnzj7Sgi4
qUJHVyqG4FYVaCHocBcpBZ/E7sfCOGXA2Yjkrcb81urcEmTZOJEk7NWRjqgoQ/h+i1AaxrA3kdix
mGqZ6CRNGCbz49SV16IlpYBQknG2/4CeBB8mdtIOdEGKPY/EAfID2CRVLQuhcqyfSEx+2GBmjWDB
D+ZgZErcvfZQBcbOcAmi/V/c7NIBGDFzI0v41dvNeE9Fle6VugiGd6zKzxx+4tzbNsW9OhBgC5tQ
AQnJKDehxR3YFsemTyi0kF5fMFBupg3j/adZYy+Jw/VODn5j2gQQeP31CX8DPK7tFWxWtiRRPfzQ
XP6rdpdEU1AKyewkEF3+BhfyeysiV3I8S3h8YxCY/1Jh0IADzhcogHkQqAuru9IynMhfUtqq/Wz7
+OGkCKJN5PLScI793j/F2bOIau7gT169sbNuPRX4/7KmHzn9c2K8qeUWA0NUVthpGsfZG5aXTXAF
PzRdIVFbsuUcanErLfq7YH/eFEZj+HZPpfPZ054CimBtBEuhE4Zm/5J69IN6/WxMtQeToBn1VxeF
uAVaLMR2VVFLmGCixM0gIYcx1zeEy7UwhtYXW7wLN52T14Vyygi4IidTX+/C+LKiwXFMgr4N4g8T
6o6Wt3tC7Sk8E4USqTwV3sa2Ou73fGQEQB0Wr6rBtANaY5El6jfVb9ehwXrgrJulbwO7lrKEhOhI
ASjmGtPPxCrYMWY9EChpmkI4gEApD0TTBYBolWxtqIvh5uwVfGcFpwq3NQigY+ItoSL0nHRYxBTb
SnkY0n2sbSAoZEUKYoGUCX4hSk3AQnKQxE0FG0YSAYfjDXXbpS+fsTActX9yGy6iVtU8/jRns1VX
nnimhzeB79MD9F/zvnpBCHBuIU4EK33luAK8Knm8KQipV604rfp2uuhjcTOn2AIpE7BslPk43Cap
HEB5dv1CV/1zbVeMZkA2KPlW78YlDmqNlD5lzx0lZ1v6uJSgsRazYeC7O0yboQYEJljVqhEV54jR
ZYBkGeXFTlq4zxChmpCCKw9Kv3SuP3yuoMW/FZAmsZlVoURCBuYIgoOxi/8PBDABnOqv4mbMf4Cq
gtYoen9xk2tqk66BJ+xAEBG1MMcPyU5/HD4DxIAPLAEBWxZh1NQQ8Wd6YBllMcl6D9EfkPw8ISUk
bOuJCtBXYbJYlJEa646RrTCltGGVgaw/sNl+KUqk4elwVRGHSzYJj6mgp5+U075x6iDW9Gp9USg4
28JX0WHVC0jGDqXbbF2iUlbJKYM0yDefF05Ae1U0FIbLBeRY+1oaQ5kJnCB/ObaBB0AMchiR6Bwk
uacU+FKhctwGeCUvGMUDjDwyiR3wYy48zBVS2j9Z41KuIf0+UrkK3Z5KMwErPO2TasW9VXzqWyX5
i/L0AFm5xrCYewvD9gq8lMAjxvTKYzYapSY4WWb4lyWjx3aDXUner6zs7xQqf6eAvvpheIpzFueO
7XKgakurpvyBprbcLoQBjJ81QCh5g9jcQDeW45zXJzEnh9m13RYE5o8gQP+3LLeCssE4QNVi9ZzZ
i5m4Q4DJiR3EUGpNeyXxF63kPEzufPmD/CpObOSOc+rUdefVWsJ0wBITH/uE4nMFiwS/I7tlS6TX
qbsOTnZB1gEr254ROPzAxMoPsDH2Ku3dQhIaIZ2x1HXvu5iP0FnEa0d3Ea9kmO7yo68/1mZh2we0
FTl9cJ8LO/3fKkfHnIK31qovcu7CxK8QhJ9gcjA1dNWcMqq/yUHLq5TaA7bBBer+mAdh8fpr7jb6
FvQrV3l4TF8nNVNsFMysOdcK9J+L7M2RbxBrY/U0524q16ndy5ffiMLU3lq9ugKCT2AHOCqMRw4a
QrBQ6onecR5ti9kFWxiky5bNHMMSknfGhmslfcwL3Jvk9ZRHXpPjnKd7WYJNcyDpyQnO1xmqMIny
I1yNn9UB9EXtXyb2hpsMonewiyA2XMFd8V+RG5NvNmXzu/a17Au6HVI5M2G2017wNxcNMvTkxZzs
mSnCqzrl/bxhU34wSJyZNFb4xEzo0ehBxOPCY5AQ5PEsP1sWK5WJdJI6D06GgrFH1OMcfT8RHNKc
8xcnXeZ1fj0ZzShhqlBD/Zt92n0ItBsBsuX3xmWgc74Ct1TXd8CiVf5gVDzckbKVfS7qJgZeTg6g
22xjmMmiKxA7pNXs4N7JsdfgyX2Oan3JKFEIcbrsiJ8kdwsf3hXRGborCIlC+Rncr9kXIaSYEmQW
k/rKmtjZwsHWs3EbbciJtOIzDdZ0gDH4G7zl9ToJqDIYUvqgh3rjDPrkm/LeXsiPFXVdWMkKpb68
CEFS8jy8D/d6rc8IOBB9152VzotooOfhefWoN3ARi2jyPWY4UaxHQEN7cd7UsRuE6rXbAJo6qOWg
f0hfPxysinkDfdP32nPdoCDgD5p+SBqrreiKwJsQHALKiyJ57MfV6S2IKrjr3sc4COmvcumAYc6c
hRM3aZ5oZBzEcP5rBtmxbImIm2+MpjB0Mn1YCE0Bu4rw9ZpzFpukANgKJCpNKPtdW+Rk6nk7nT8u
zGlprJPv1+e2GbME8wUogOayh4E4TwJxxT3Wy/v6ppiSEqrEcgfc7okGsKApTLHCOuvZktgb3wns
EJamBWbcHBmz5StE/sf3BhMp2KnF7oSiqtBkqNsobXG8Ac/CezXUVGs/I6rGTKSfdQibM9/L3iCj
SG/6xanzzghKFFUg6SiCmKnP3Wauz6i+uoBYK0JFRJTZKZK35wE4F0b1fqRly24ITyqIBL1YaE9n
hrE072Qm9ADaWHd1AoOKm/ScOTJVqhXMFftACsQStkeEXAdVvjrT2AiT8T0nbdN6IqiE0E9Qk0Jc
BvSi6Xs3X44xn/DoFvFfCErl8dPUttHZfdXN5h3iker6LdLcoDpBjMoRYe1zFXCsVJWsBdCm+BAc
7aw79K9Y0+LHOqGAe6rxAAnK1wK4QpPaGOx706kymQtT/v6RlUuwVydjinviCF9IG8bR+Xj6jkGo
Ycm13Ts5FUQY72ViGfre5O+lu1edtNgXZPHDBm1mL7E7dpVQGnUiQQk1PICIvmOGxEAv0i3MXD12
2z23O8V34z4LK4sph31lYLhWjhWoHMXNji/wPiOGGWjLiWG8zyDLwO/BmCjf6I6IY+UFmmBertRU
iCgwrVMOe318lEAsw6mtKxORqXW0J3II24V2bgbd5F5aGRMPngkRajdioHDYrWiC0uSuJXRZsnP6
dXM8QKny7ZZsDeJNRLITgh3Vvg655jECZDWM2erlrTCQoqWcZaJBL58V4sM3o0XBVvpFRcLXJ+Uu
FwcrzydnuAVqBgLpT4+tgJ/SMjPLxhYkDwOCTwqQKpiCDhY2tOgtyBQ+p+RWh7O6tZ0r8YPTrERL
hyiFw496k41A10FYrMGQcCJDteipjPo735QAV/hO1oP2GG0krYST6osCOm163REAnZ8yE1Ogjn1Q
Ml1Vfq6/kvb6SYPgoy1w/ay3IidXH4wTEzV2Jf5q7XKmBGlJXHrwcwZ4ioD12ZkGICYGBtwyTyXN
mLdx0Uvv/IaPGVw7xrsIICfluso5RdHa2G4qmp1p5WVB4kZYgjD+5/kpZCULFwKb+dx+sSgie3WJ
C29IRsXLFH0zscEpRkPiN6WnI2Q2pYo7j7Wkfvy6ECx/pQoqmtTNY0Y2yLDvrmEgLKrvp4m4xLGl
zTmaIhWiplDUO0LW+7kyV7PpMIjGdstz2RQ4HaSK8geSS+FZlWc4NSV6boITl0rKz+f/BJQ1Ib/Q
sAIuRjUaCAlIXv8+61iZRnwkpBdNMpfJ0Cpn/ewqr7YbT7sHmkWosT5sdz8IizVICy6k5aq2o4Rb
vhVq7DRcqjcX42LTMer8bIRIgBDevj3raqUO0NHrFf5PW8WbdYFDXFEr1kAxtE6FcpzhE7nn+paR
tJbZhp2boBThcDfTc+r6DRD+CnosxiIhdjCZmQ75gTYBv3keG1Ba9YLIxJJpfFW7U4h+jlTC6zvp
FeRikYIlGPXruSPWGCmB3ABhbfRyathz67eI57XQ8eR3EZo3IfB1evjfLUsepXtdSD/Zrt5Lad1P
A9oWEG0gCapMZwrfHERMtmuXV7DLmOhfgW1HvvrkSos+5k4E1NR4fu6sKoJCviEKPnDNFbA6pNhN
61Yoh0Jb4hfDCbaOU7+aL36fNkkWEAoKlBt7zITqCkN+ZzhQgKbon4ZgVg8nm5jSFgkfcsneoNR0
4mI8bDvm1A7BlMSXa1n2KAa42ARuCprqZBOpCGt/R7urTACVhIURz+n/JCnP5ZlAJ61uQHs8N3Nt
Aho7BWGWHg14DAKZi4izO2SMjVjkoOejqGUyPRR98y6PsgvreMMdDlEhHHZZoT3AbictG2f3FgSx
QqN9oMoYG/IkTv3ULV8iiPLkaEEJcQMwHt2wAgydzh9XFBUXv1/TOjU9IPzTzKtur+X5+Lw7mogw
MLD+GMWmUpDs+ACemZqztGeVSZwSuiykzKx6K9k5CEKI2UjAGM5DggfZU92vSlsFum3q7nPNjeig
rzJnt/xYKcHSYhnVZxhyzXI0u8mzwZD0g386HvhFRL9sQ9RKXg/xdIZ9IP+xbIwmYCHGXS6m96qh
vqm8yBl7isghfO0P4MeNdrNhM+UdC29cJfDn9HfDTKx3Nx0D3kbzdI39jfskQJ9R9++vO2sUDyHv
sf08+rQnMMSxF5e4JQcnp5e+a6BxyhTBss/JPCzjtgnmUQFL1wdWQcMBqE53zAolf3FQ7iDJtIQ0
YsqIlzXDutWTbNvvLMzmgBZ+yJcwyu3SVJ6d7gnZ5PDwXBSiKjDcliBzMGIyY4/lEHmCw6+ioZJX
3DD2VwYxHI1DVsOQWgP94FCI7N5p9YNJ1hg/ROzM+C7XRlfnueN24aa2o9gUfLryOh1d+CMBi2xn
xbyesIwsQpyniZeSDXEe96cuTh5we5oMNpxf8bTFaeea597M/SPbYaKzntBHoK8zSKz7IxLNYjaW
fU0emX5DWQJVuJfbFw+fILwXg2FvlBiSVYAG4wbAaerx+P7rZ2iM1LLmm53dF6eInSCS07xpxeA/
9OhCnVoyAEM6WJDd17tQntaH7UmAYzX1Igpk/nTtL30xMb6XzLu3HIGktERMipc3AtAwI2mU2ua5
gmgnVgotET/HWivbPnk1vg9+NNlPIe1Xz8FFG99xWsoTpSjbtnPp46gvH+56MTItnIF0N/5UvQHi
XJqRPWMifHyZN5pAH80SBathikelmXHF+1/dvok/lRHv7jZihsqX5ro724UR9AsTWOMmdWAe6Iyu
TlRJ78fUORluhE3LyxN7jn8b1H1WhlhCEcU7R8usQZ449tcI06/J6ZJOvc/DgqGninDuJH21t5N5
MndNHmKT3R8FbrafdVkzEiiG67ViBe1rdcDFSCPS78NhDktK+EOB5LiDJG3xLHht0nYbk/eZcxoI
eBP1MqJKQ3or6/0VdbQhDgdMtt7CEM9YGaNYahfGM+21Rx3sAQxhFSr6XcRl1aAUTtwlMkEugUfF
7miUDOwn+92mHqjJWoi113ZGzTboh0StnrwsyaGO85HznQwTUn93ah3z9gXiGBLGvbFSfvoTaIpI
cOheeG/jq5rRgAdTD0+uLiNpQ3UbmbKB+KODti7a0xbsMwBKj61NQFl3YhW8x3VqdTedzkn8ZRCK
O9B68Xk5/y0BX7y5ASDMZpXH+DElbIC9fz3AwL4B4tBNOv4ssJNzll2OSwKPIBt3XMx1NeAQaYwC
bmEqNPmKdF5Wis/7SrVqdJU2rsHzQTvjxuJiCpdUd0BSPYwUge8gd0MqDTr1CKofD+Oqb4HX6af/
MYHhal6MoKhzrH6inqR1MnDJxJGwquEnLh1uhXwNYNq2CQOtFrgh+ZorUo/rWpyKIAS37mZKgCYK
RgsE6l9Bhfv2ZJ1sVoMaLcMA36uiGnty1aZizLvgRiV66Uj5p8lW28ZpUsvQErw0cntp5Py/xVD5
3KvXpE5lHWveopVswP7OWfN1TLuu9FHxlEGrkO9yBYWjkvUOROJhtE5uAxiZpQpjxQAKq095h6aN
XuXLPkc3wUJe49bI1MbDi33mj1YZQnE4TP4ZnXZ3XD7YoypNT5huvMPz5LSQSb6yYcR8fPyNpJe5
1S990mnA8I5c2mfJZs5BOh2/n1e93d4SoR/PWpbBtdcTwiz73/fVLY0o7Iwjabej8G/H3HEyy+u4
A8eknfDjx5fGL92cYsbzSMq9EU2mWVaIgf02wucr3BpV479PUV8+3tvsD39ycQAKHaqTwStddLzt
kJxB4D91L1d0TX14tGBKhAIgfRNkAXFA50+I5QxP5mmw5k5rzp0wBgI2bdIZcEbzDkJm3ixZ81JB
vtdHyCwnrzz8D27/gNO1Uk5xkaFuK57noM5WJ1lDlwF8OTlsw2OsInG5MRvdQsyYlTzuLipYMdhh
oy7ebMUs0J3bNhkdLa1N63Fex5OF6sroyI0LoZHK+DsAuHwqsfR7RRxYCTYcEUn66KsLfs0Wh+mp
HNnWLAZIFsPL8nsKuWd/0PMFxoZ5meq4DoYaEiwLYCmIJjEan5C3gi4JpqibAVB9jlTCAawAB4fN
JM43a7qrIHGyayn4xifAnOI2fPna1GgrBdzpZd9RxzC84Hu30SfZNirC4THHBziYHG0qoG+KzoXW
ytkyFT6ueqQD4R9ghmemtuCdh69s20YkH0blmdWvG8aFa1Ha7ttREe/F+lspuHTNArSCA9KJRQKa
zdY8XFRGECI2H033dR8D/n+8fxLOniB5/vF8HCgpzdjsbILKgLBT6CPz7z3YC90juNaFdUg0laY7
PE3esMS90nFUMjqdPxOS+tzQnrLCiyj0rQ1QJA5AC6sN7+BdROsbpUEZsKsg9pW3vs2OBXIC+HBM
f+PhQwbiRtScagGx++0dKqJYTbdQe41YEEklLz67TRZa6p9CE14ndqBhIFext97l4jNlrH43Ycz+
vY9w7H25AYckFiwzlRewiN/tCLC7tURMDcvtGefUI6SR83CXmXPqvFepNKqdTBt1/zFMRGbVbRar
dQyiXNYe/KVs3GjNJKDI74zmnr/di98Te19evpP35ZvGY1zg9yY5iPyp7UnrOCCN+svRLAyQPW4M
AQIsahtxTZjDGs2jOsEGQHC0X5UPs/58h5Ia6b0C+XmYbVc6LcZVk68T6InZ+l3MHLsjzKSYUOwj
jeOsPD9FV3ZehM6tVbT/wjB2KnAVmQTHpWL/xy7W676Netesx80UkthLgP8zhCfV4I04Vg0f7azb
2WqDDbKXbJhaylInOnvGWNXikgdZ0Pdhlr6cxOGP1c5G3Ab2KiPaazjc7xqHrCLo2FGIlTtVG6Q5
zD/ewWLk8zDbfkhuG+ev+74W54kt9krQH7ySQ3TnYlWsv4i4/INdtXGMFessAKTBOXgV2LooBNm7
1GEyG53YQHQ98JUs/IWZonuJ7jKsXt3+SKAGIIvaY/WfO4o//gAxmLiBaeQVtoXE6PF6zkSNCKrS
P47NkVSkK9MWCfYA1YrqcYhFKQOLdIJXbXh10nLOdDMuVp3ZD9RaFfFsY+d+w9n2E+LsFf1v/ev0
7Q3SICqHy0KrL/hBrzJ55QamzY0FfU3qF57xWiYnDgrB466Zqo16HpRvZ4FnTkE4vLb6bymmGlfP
GMqmtigarRcsJhMs1lMTr1k2G64J/buJj1a1/FC2tXhUGKi+ViXzSGV9PALyKEtgGSL0tMfVteI0
oAdFOCfJv7fiWn7zV0phl5ssL+prbjlq1egDpOcMm7Exp0lw4dgYfRfmmATkaAdcYpDVkmquNeBE
Ije4h3d265pZ2phnigJsvZoNHCEIvs8tko5OFQfM9DnxP/JJlePBJPOWcr91H4FMU9r1m1JFnzJA
x/vxXyOQH7bq0nxiVgGU46VEGk46+b3fqlYZizXwNulRGzcfy8jJwSaWwOW6F2ByZyxtE4G2mzCs
RJd6l5XaJP/cspAAGEQvdiBUTbdUKfcfQBRPObCd9QZ+uwBktTkZuHcCALnRZZ3k3zfd3dzkURvr
NrgbFloAyTgDJN854/gmNWRMtQLuWGC7FrPs5aBAa54EhfysOb+ohr4+4Z/295jQDIGEzgxCa1/R
UqmFdQrsB2VZ4cKyz7RMq5eUCmdebXwfk55No6509h//PrJNpg/OFHbCHn7TGmFRolblyO2PtZXF
SBOrPYRnh3EJanhaAqKqIqVEwJAHY7faRSqSxTEg+R1/gLhI1woUlFSNz4vrBErDpXzyHvneVm2Z
wYCZplmaGJyfZ0dgC++Jnz+ctjZlEHjU2j0Tz376+d0AkMpyIhTeGzx3TDE/2lAspZhAr6cwAw1q
dnU5DY5g8AFxZ2EN5kY9RaOQueLBFPq4pRSGoPWiiMjrdIOVhaVp+xXAFq/VlN2kkm7LlI0urO4O
1yTbNeZLD+Nr77HonPtl/gsPKEyTwCDXkNIrZDOWGmG8kmC8b4rYOLZgYuMcuTEQNNwObZVL3z7y
g/VhPqa8NXl5orTgSWaT/plfpWlDPYTUfaey+Xiui14j+qxHTZ+GR4FgFNqv/a1ifFyzycBmvG+O
77g9hXYwI/G3IQzf2gCp4dWjJ+4JB/4HUEnwlB95XAx55pQKh3N0Yl3g2W7s4SPfRvbrymAzghSu
kPeku7LFDbK+L5To2+eOwWoNsy9dP3uCoveqDucPuyRknTSkUSOXjgrJbfager6RQvcJUIAa1qa3
mGCUEesD426dNhiqM2nBeRyyqzkMRm7w+P3imysMNXJV6N1B7oUUbAWYGi47WvCowo1fN6pK9Y1k
Sjx1Ku9472jgBkMEtvT6jv1kWWPzLypT6z/jGhW9ZQEFDm8ATqD111YFNVY8ka7vrv13NXJlYFGI
nOAn+/DQ3BK/EClJePfFAoEoW4lZz3jB83Y6qaiHieDfIOjICnpV7LssyUs3q2EsVwfzeS6FRk8e
fD++ALPkfuQYMTDHqEg1w1/nAb4i25iSHZKQVB0M0MmIAAEdpQkZNASfvw8nrL4Vjnb6s9aZ18aB
muskh7Qt6wrsl11y67NVUgQsK5sQkUpsUp5S2JHS2zMydBjTvq6+9u6YG7q/NsrURXFlwHbAIVKo
YPWaBlaMGvuOZka/RYu0idGXu+Bw/zXNRXpRnDe39WfPmBBpto45eTurLHG+4kLBuvIu4L3UpDbk
AApewg1X1J49NGVza/XhAfqlbuKC9aNctHj6eGb94ZdONMGfo7QfUPRRJbnRJGgQkL3o9tVvP7+O
Ib/eYV4jpKeWd5iUUIG1OBB7qreWWGfOSEuexo+VDkqTZdjdOm1lAqzGBGWlJFSncO1VzHzFa10M
I0ZLsS1YiN2L4SdLHmE29s0HgHP1XXKnm3532nEToOOz71+6BZuNRanHU0MrCKeXpiFq2x4/TdhS
F3ITggOPsWcUPh1XbARWYBo3Ca2iqObudNadnypbYIAmCoxWedTWAS84IRYaGwlMyUMPUCsgrODy
QbL+eYAAe8N3mysmvE65f5yYGZ6ULu2Y153Y4Y8gmP0LC/9pOQSpxdBKPzC8hXXvDsLvBuilSiOw
CtVvZIYadImDKfH7g4mi853kErM00EJZrDQu48bftO14mufrUfDN/g/XGNPlc9vhCHGwc6a2YlnY
UbaA0BAZ/JMu1zD2hZ3gmjCYPKuBXXpUzE8GhPWEWhNkptOP6K6b9InqAQqCT6Gc+us0kHWR7hXI
8R9pboxwdWUPti/waw3uPPonUI12tWv7+Czu7TLGIcq3E4omwAd7809gOXZ1IQ1cpoll8J6U1kgo
XY8EN78TvagYcCbuBEycGGQkDxnpGBQFi1L7h3We/rPru7j+NToyaphbRCauj8j8EHlslcxxrseK
jCYsDbzF7srt0Dh1m7/uOkyBqtgJwFlNNLSGC7GQz/om6Wchx/GhIIdPdjHA73KwHbTFi+UY1C4j
aPcVGjJUYT0kxvDvY4AoeYrGsYvj5j8XGuH543rVEp7jfQyyLhT/GqVdd9S1CsXyZo3rHLr/recj
GZHu0ZRfYCF4nFH2KWPgi2iYzO9/K9lRqyW+JYUrA3k4tqCILl+4iArMLkkFHbLG/1SK7iGWT4K4
yzJET7uzWXvMIdDdUaEY2TKl9y2K5eAFIqILqjzIVNrXRqcG+Oz9+z7qBzYUQOeD5Y1pKIGDgLhX
yTYdmOYB3nRg/3gFAMftpxl5G/GJ5vZckE0qfKxKnaqyxy8JZGtth9bJocme+I0Gv2xWwdgjjeMS
mK1rYx9+siT5nO/LAHrYjfukSbhlI4+uARUl1h5EF6JamQ3R6DfOeCAa9jyt7QTGL0jx5KYBEDsD
sirwAD8OOzwJ+aqAcuJL814b671pjTZmuPUUQUy/nMMZFGYkGdnviMeGKtHQridBgAQR7G6Q3VGW
ztMYKsj5+uwFjYSnEbAv6Xyizj3mXXvcnUmFaD4dcdmNx21XJxCa/qUdjOC/4VXhQtn0q+cLwnwH
OU8sdVy5HdGYV4AiuMnPXeJwei7pBPHNojScDbrSGd8yEbCKSboYDMmZ0morMckDFfmzli+WLUTr
0y1aYYaP4tDUDFS7sdkSXklHZR41x1mf/eTJqRkKFenRHwmVWKssWiW0pl7QB67b+Qzsk8PD4iSg
vITFvfo4asFsaA2ea0T8Pjih26l+2pvZGWeh2BpGdZeSkHd9djYNLTBdUTZpWKEV/t6Rtn6tIV+8
5GaKekENo/+WXDoSbWrLy9yo9OoKdtG+A0C4CXsa7F3Mt0JVVLXLjiPq0RGfFz8YabcXmw/vnySF
sRZcDA703Ua1T1+lmQy2O+Q5jFUc8wnmX3smGZefkishJATLBVIKXmQHXLJr6mpiLDFOmVUhXG97
XZbBePw3N80VzsUd0FRv+0o3vYD4cfzASkPSzq/EjEO9P1KSf9vjXazUxoGUSgw5Xm5Rma1ARPBn
IRuaLpAzLZelrv0sE9qwiRuDU4KZ2AJQgUHOjUb0Qz/flu0ZwKUxrj4+ahzfMO6b5UUwnnzK4n2S
LUg2bc4AIYVtrmqDMG1I2mseXmTN3i6NjsZlfEpD21OK87jy5dLRup+aroX8Ze3BaYqHy/epPt91
m6V8stQmhw40h0nxFeRfAJGAvwD5vGIpegIqSjl2qZWf4A1MLCRhV6d/LzWhygoN1P2Yt5yBiviV
0R0aWnNNyLdej5DifSYpywEiE7wpinyr8cy0JfydJvJJ+plWggMb8/nZ411k0vcxtmTrshdCEauI
a5lgMIh4oT1mRdCniFDi1yehDpePMmYUAAD6pg9Ju9kl2cSHxoXjRoLhjpDOVWm2vfWa3YqhXH6b
k0GreDnABCl2KARsqajHiaklyUZG7YiS+0Km+z9x4qXfjJ4PzVZNjAxb+NjoVix5eY4jUSwGQZiC
LaxTMRC7ERLLXgJ7Ar0bzzRTLpGaIS8n86pGwLt/nnfUz1BYwQKdx+tzn+mfLBwkvnEhoI5uB47Z
GGm3SnBss6Y3lw2qBgJ6wmmImlZk0nN3VK7l5KZ+cDZv4yiKeuUHmUocVQKQVQnAQEPPy8652SU9
euepfJT6+K7sTi25o23FySYmU01iPZUTP+amIPRCdS6mVbY1vSW+J45RIzethgMum+XAIbfwRjiQ
fVHFZX2TP6zxji+KttoBmmUUvgsEublwINtXcpin8edyEqsFs+wNoL6kwb3HYyWKfEHro7cDsIGY
8NO9Jj4FRBIQk/cARcGrngcDTAa0hFZz37BEK4p48CESMgIa2FWQj07upa+28AR2+scOG82d1nIF
Jht1tKEmZCp1XFBcAMOfy/2x3xmwQ6TKcAroo4PcsHiwQ5Crf1cPuAWB7NVooMdqoKS7tTlrVJfW
vanZGlowlVwGOMfzjVH3ll11y4Q0COGHaiP/pP2Wgy8PWMOMthqWrEClmDR1xMoM+oSrhxuLXV0K
aO/hFSSjARpewj+62WqzV6Sl9Fo+ZL7GpnfH2KNW0sS46buJU7Lp4GDqCTnbYtLWQWizSqG8g5WM
DgjQ8x53GC1coxsyv8w0Hz1HybHi1nX9e7raPa0NkhbvaCEoAJwplb+4JMg2ea+djI4uF3rHMmwN
5wMWZ1nSYmIkilyOVJfm8/wgyCc4uLfCc26pZzOdghyXa3+rFc60jPWEXy4eR9H/jL6LgIPLA5yN
LRj35hdi7l1dZboFbSHkgyLTo8mhm9SpN230li8xpxGMy2J33cfBrWoux1rAUnfdIqbfTljpspJL
QbNWwm7aQxXZMc0e6pGqy9289k1hJf96UMvWJHWFAb+S1Fd6CSS9UYbCIAqkslcNd6FTK8bXdiB8
fdWU3yA6Ls+eWwhjtV+Ca21p47Fj6DVLytmDajX8rTukyZOu1/sldQF5X4+qGM6WcTx9lH+U0YJ1
cDKuRQb1kFNptb4f8DxXkzxtJUVdvCZWbVVLZSKNfGoHKYWUAnyDuApvMc1N4AzeCVL8hf89G2zq
UkrhU7tEaolB3PwZUvVhWGXrowESGEcSSzS+4KPnS55jfP55XX6ojoPsEs0NcbwqkIsQTqevJxma
j+JqMvkZJUU+xYu0Ws9BUUAi/mb4dm8QtnjPdFGSFAAcVkn36hlhS36BKQvqZaWbcKc7HOnWc7PP
B5la5PBBbHotX3wefLz7lLYj3sKjlYn34olhYPEOCrDg2apcqaE3m8NIXEFbzrgEgg0mc08Pfw1X
a5KhTKx/COoI/FgYnoYn+k1/4IKlRNDEa6B22x7ZhTW1KYWWzV/ozh3+nLHnT51pWD9qC80u0l/9
zqF9xk7rQ6kkNDfMAe438l9LPxjEtdKit32skQI5wEwrqCOSXBYFcY1beEBH/bFtasgkvj4rxNx0
hYzJGP+ts43ASGJNovdnO37Lcn8ccnDXAsr1SU0DV+ZeXK9zy2fp5lMf1dpdBLQc2hzgHw93djCo
O929iGShk9g2bRmy3YAACTcwZciYsNE884D7QRZmN1BBMLAWF3roCXQ4DDOGsgdoMbvBqjNEOtD6
gpA4wBYDy3xWKV/krbqK3IRS/SgxNWXKnQgeG3+9ht1vgIxkBcmceWl5qOBJsKWkN15SJLL0SjYD
WKRM+YCCf43BSP4BLaoCRTwluBa9cLxjQOKJMaZ3W517XQ5hz04bWDhEzQNjMof5Az5sFbKYYyyM
/zVwIckOgzSBNTpT6A2u1dSRIOF7PWKGA8tNjRTWmDeuoK9OObEJWAXe4IgIFzNCn0oGDjQlkybh
tEv5/K/0D1khOMOa8D4VsGGuVXX6VfFvkA4OHSp/BCmZdboqzJ7PloEO5aNlEjMbnXALW3KbbrY5
l8pVgOihaTtaHul49Pzcxho2vzBXN+VIk9ourz1c+/dOX/VM6oFC9FboDtOdu2Kh3W6DJPKTp62r
5kNLyF+zVUCk6c254WId4uJkPFgWO7/6docMfuCacuNonBYA0hYCsI+n0GXiGQA21loJCaT3cqWZ
GuDdg/0SwSbvNNWn3rOLxCORo5WQxV/TNMj+Sa7DwREC+/kE7feFJhj37tEeZFZDqpFay9Dc/j9t
oP1ZHl6BUKBqNDOvsjUMa0nvA6WcfHgGs9a8XnlLkX1gS/xqIBff3gmGwa4FHFFQrGsHMhCdGYMB
c/MR3JfX38cqn9adHejzrsEAIyLMmkWfYU9699pFYV+ptkLp/UW4iMURjQ5NKO3E5MFjYG32RFLF
Iat0ayBH81Lp1kqfkRauwSN7yjG6oECOXB0Avll1TV7JjpZxagqjtP3qXUi0LvLHzg/ydXERjsY5
wOQyE92iuUeD6xsNoEdYkpggq4SyX5Wf58BkAE5SR8AygOjR2mn51/bZZe2Eq+xAcg8oclhCcB2T
9BVRYtf526EmZE0T6WgCYRuVwjUFyFIe+Pbo6KT8kWVkSjbyafpVKLKamxOk4SNNUS0lhEKGixXf
N/gluLtBRjBA9Lel9Yrsa2l1ICytvS12NdtQj8JYzsBvSl5qV1XN09t/5IFfy7tKqcWP/NJs1bKG
KdH5LcVtI2ih2eh/ZcJ79JWwxn/apMEMpPfucRGWcZqBfGWtQdp7TCJKqb4KMjsZLUfu2gnikfqS
NxruOGC1OLmtZlfAdz/KDifRktd2ovBpYuHnL7Zc5dR7/7g6WjPJj/CrSVMQwFZE/G8er1Fq0Ev5
dC349H7q/Qd4Vmbpzl59c1e4MRglBex6K5bZr1t6lqCpHQiuURioB0KGswuN+C6u780+6my03x14
5dprzWpWb3izBegn+ZLR7wf86+vek2dBG4K+LjLg3u5hpCAXE2dK3OaItzEe2OMljxo2WXJ8WOiU
LXFV83LhTGnp+JzUdrXGV6bxXcT6ToYXNHHl/uvI1iQfmvOvOBEP54IWEU0jRQk0pJT6nLI8WxvX
kw53mjiTf88Fv9Le44DNwAn7/6Q/jpdrUbr862NTmpPe9xuj3vRsmzkTQn0fIvovXEPdW1jd9HFF
7LsW+3DxEG6/hx/JbsN754CvRzsks640A7hAr+ltNNIqHuQFHVThZlJreP73tSghtlNu0UDDECkB
fIHuFRJcQ+QZkAkWeaHe1qIOjeYgev50Z3Ckcu+DgmZbchv6LXg8ZsqJBUujlEiYI6MDG8kbOfru
j7lEt0bjj1xdYuKoBvT9UbkhLiGFmezRe6g/2KbKnvB2Ar6JKzRPxKjz1rr/viMQrv01HfrqgA40
FlqfAAsdQ3ylT4LGrXOcAxEyYk54wgDHprW9/gIZfL82kIq37FT3ZDtk5oEcBT0BuW6Am4nWwbAm
xkDLkurX10q47ZO8gZpSzSwMgfSQ6aj5Trtt131Cnzd5v+KGW5T8pTwtHiXPu1FGtS7aavD4nzI9
ff7mdBGwys+KMu1HZRGFDG9X50IsLolzSBExqCkNEyfFpD+9ljCd0AX3AM5Foi967jCHWH5MugCt
EAPc0m/y4Faxl9UdeNiSBL+7QquCrcKG/RtUH/Ymh84AVXWPU6qUTr0Cedp39yxQrZbl7bA0I1O0
qtLPbnbQ+tdUGW3Lp9zxWdrfhfTEXauTnmd5l71CoJRSuZva7vM1IttfbBaFvBy2GlMf8XpR44oS
xDFarKmSOYss2H/bnoPHO9smJwMxZTjzC6fIknFNE3dOe36dLxzIDnpHqH5tPhV3Mbtj+nxuPuYD
ZH65yVcLkX5ce3gHN/hIi0TqsuK6JQWM1FMdrAEfKZYNcefuAy/A/WP9y1yZmuE4nLPtXAZrufHT
q8r4IRHzC2x5Yd3uuAedkRQvjSjQndp/hkn2XwWUijJc6ehKdbvcrklY93h/ZeA7p/7DpwtML8sE
Dv4O6cbQdaWZhnUi5Dzzy+5GoA+UzzktbUcfII2z3kGS68kyaNRk8knyTSzAakLyG/GtwmzACdy9
aw7TSEabGWr7hyyISK0H/jOk7y1D+dSp7BGJTKioZlFsUHvs1vkWng2aEaGHWrB2pJJYWHhK6RaC
7cd8HYw3YDqC3WuFD/QdzLIRYUMyi3GzNmH7JFiAjJidZYN9MRMn9UzAdhq7ASIpOn4WMc+/oqRL
r+o/8UJcGawprFHDvVVQ4gTE5nDyeVqOQhQ/tTBFA2Esb2KEr0YS1kGrimNGUG89ClPuOscItYsu
yn9eOwkPwatKoHIqrD9traWMmq4dttb4b54JxlZh895ZJjQ/LPXKKLKrCybAaBZod1BZ0r/Z1Zy9
p52DuUcggZoZWH4S1MmeP5UU2Bvn1cmDzoEldKU48bIGhY49rqnHDB0lmTOpbhzeS2NHdY1lbOhI
vLkTSCyDdideTrr/RoBkcQB5n+0Chk1GTRodlD4h3D089BRZnvll8f9ts2wj3lEMvtC3tMhzvjlL
81+1lAX4255BfzcPW6ohtDvNt/Lf5ESxFWnWwlvm74sDXw7oLhNaowr21A/2QiKJvMBA8pLwXS0l
AKf1RQkW/BZX/9XPDzgWqr7YLIFqtH1sFNZpJBSffyod0Moj0ah2CMYuSi67RIyjZLGRBwDtwQRq
7poX6WxtQEreIqvWEd944rJtdAurRIN65WLuOxzjRwvp/m9CbKkk0wylZA23nidqwm0z6ZVgcJ0f
qTmrU4joKooXlPpVvMTMkCLuYv1n79ZnvdNdYUWKdWGID58Z9qDZ9/55I+GlQLj7TcONbRLHnLRO
fT07zVH+sTqGgj3Y7OTPa6Sz5EFrAEVNhtwyFiHdEB0//UNhFJ+kyvhRynaBE9ZeOhPuIHsdp37N
0pAkLei0TuZPezMMBV9MJdUU4f5goBM6COvC0s4hVFmaS04jX1sfTBdMye6bslA+l5eRT2F9rKOb
5GgE/TZh3oeU8EvuYBEkHCRWlOszEvXVV413XVzB6dWmzn1xYBR3NzK4LSjv4l1md4rbeonrgWfz
pxc1iCrEGGZzlsQ0Oi34roYc/hl4trph0wk2WaWGtf4uLXjEbz+MN936X/Ok+H9oJ0CeForEE/st
gukx5RX0NKktrUI6WTnsIzDpVmyKS2TI37P6PKETvQIrp7FKazjoil/EMDDBBK8a9R4dsvNwCdwD
HEqUx5GeS4WzPkIQUSV3RlZGOySvTinT2P1dUUwbGds4sTZoUkoOkfT8/e7ax9JEEDldLPx8JNl+
54tNsLa+6vZow3Po/WAxr3VN28pkNXGtO1IArdtlrTrxISnADcKBAyaf+x0T0hiAHo7vJuGMf7/i
MM+rjgaO3B5xWi/hlnS2LOQl1bOK3TDHy7KZssddhIXPk9Isshtet99VCMmI6ejLYmF5G6ueC7GV
5FAUtuSOMT12zXkxBu8oYqcY61g5POLyJ07TqczTR3LmCAszgVvlwFl9x8dxgiVcCQMJbcvzdbPv
uB02er2T/jqY05fXjesF7Ke4uQwFH10j8krQB0wragcbDxheIPyRHvwv0y/+O8aLIWYygtamM4n9
Wypa4zPid8YLgSEPMYmh2Hw6lHQlZntVjQ8mnL8bbXKrAkC6KRY6ritCMWu0kN5eH6EJFe0f3xWQ
cI4ozx+7piVgtOu04+7I8kZacQi6IyZ5FmBlN2gAAHyfhPYBESVwDM5Usysuc8dkAr8nVhGV58sS
dulqHGNGeTCCxzdNC29HSoqYLQWU+27CAfyzovfH1GKdh0PojDcxLbJO8VY/7DriWDydQcV4Fz0K
kmJDwSrHOh7FF+xVe2mG/XIFVm2tyhYUZtclQlg3SDviRWpe1vPSxJ4OoRetN5lxTOu/zVl4JY92
2AhQJemC6TPO1YVjHnWK09WyCoeqB4P5mNM0RQyfiu7aM+B0XY6a3m77FZhchNs2kA4llKkgw27r
Ef1AEYPOiK0IqoUp+ZL/Q4lPrtQF7cVR7M18SLujIhwW0Uw2WO3+WSG/NM6ZcscuFzgnWXuzS+mn
lldylmHu5ugp4M5Ht/ALWyKQjnFK0i3vtIOmW/kTJ+TAs7b1UYWzjJxLMqacJZ/FyF6oHB2WDr9N
4MKTqOhlX/i0/GvKm8n4Pp6ZggHW21bzseB2SV0HzMzHJoVjZOCeAfesXr8xzzM6oRn2YKsjNyK2
Xo3bG9h0wlgoVQ/4RA785fYTWxh7AOzJv/VzcOVlcahH/ADpyovZl++A8h21kYX73M6uUE0giE9c
hNEuA1O+XSJVWYiQo4l6kYTaCvousZThCynfsOOzub5Xcfua2YTusrA8Fk/7BRjod3UU3CIkt//4
0IrO434uDiU04qo3Ej6LbW8ntGz5iG00+BjxXgkwqFjP1JPaxfu52CfsJGXXy3s3R2MPik+B4+Bo
+CSjYSu+cG40pETlOFt8B/S+TAR+3SABV0ljfmc67FifV2W+378gSzmzWeVwoEiNecyjYLgLefjz
OUDcPPosm+QsRi/YeBzjSoP02dKBt8H4WsN5+8/wumWKvSUzA5nXyrZ9JhAv6S9617GuDgveJRIJ
TC51VpXl0dVR+JvjgozMAfkHHe9eNK1wPXVJw1V8qpgOq+ZJpSzvD2QJHDWckbhrwXzkiMf23SVV
l9sDP7H0nbqrB8fpfnmce+780fjYxTw/LTza54hOqflEMOCIcBsh4CtqipjfiK1dBe5fG14S32SV
pD4tuYGrtPpu+2QlcP+eVP3xLi1bS6LUcp2HGjcb6YIoP0oqPhdTuQF4KkfP3UGXxLcjZnPC0zav
eaIxJ1AppYn421esDyeA4INchbHzHx19zru2eyztpGZv0NVWo4xRe91fKvQvD91pPftar+VLW5mN
EDJ+SRxtIr/K86wZBKJmfwLCy7Cq877an/QHNIa/ZWPowN0KwSJPLn4pAGE7eWhzOzoMts19aj5X
TJctU+Y6X/3vm+OFnq3NC5ZIvt0JseokirOuJicnLl9JhAXl8W9PZ1rrEHmiXi6l3nIoFhAI274M
WGRfckCK4l8VectjpwlffKLEMaEhTc8gL7hu7xcbkV46KQjjXRSsGpG6itHMI9rDmy2ZYN1ctH18
iVH7wUhZoKPAhDrzw0mIqOIlSyuSEJ6mAqbt3heJnuOKZvXcl8wJI5gNyBsj2eKVPeauyrOzq/6A
BPTyikanS/GN/L10rli7rNizN27guNcomQCu2yRvYc0ukuSi3Z5hHiYtI3eYRqETR6F5UwbxvLLe
LPeFszSbvXmwtvhoep+vcJ3RuY7gZhipG4hGHUnCPTnt8+2WJfQCBegTqT7ooJrg4m0gyxHFPXf1
MJaLocj/PjxPvBsP0hvuFqi3xa7y4oHM5YgjOB5xy4qyPebNgyI3LDu+G7xXvZEKltgBKKcpMpgC
1fSnvGRxrHnnlsD6BdUJq7Cmvzz7pMIe1vSUk3d7udMeCx+CEIHNTQQiWQYPm2cDZcoLtEzDBzUX
NsL9b0ZZ2sBGq/m2ajzz8ZCd1GZbMBxgZBR3p7nMIEW0qR9ILHZ8sodztM4GCP8Wf7nuwO7RSpc7
5/bnpGNe1VnprmhXVZqSagbVOoVca8P8ZQkPZxiH3fLLgP6sJ/mmH0ghNCjmVUCBTJXdq5bvw7bT
/scDuZvS8McpYc6YrAbkdZYVTD5gTbx3Y+BJZCGolfovI+vPrM4Na+zN3W9swetS+3+TJMwYqBDB
k/+a4muGfFyKpRy60ZK27XJOH+A5qH7K0sdQ7L/QDeCkIZbWtdIEt9kqaCNLu4hOLzyHd8r9c0At
ftuj4btga4zNwsjvulOKOXfnAufzmsrTppBYXb9d8wtxqjTu4RTxe/nky66IIzY/zKj8yB+X6H42
2LCufr5FG5k8xaeF3dCZPfqxx4HYqlbpH4v+TsXUwnjL15mQzvHK86R5/XWbCi0KF8PyEkHmLaEQ
+O5mGud51MW0ApET6JitGTcWbYiO1rgYEpR0QVSwCO4KO6Qc+Xoyi+BmN9iyS3Yfy3601GGfRfhf
qCN+Rnuc3fWuDn33npCsJlCJWgY4nrRlX4YIMo+wJSIg/j7zQnIK3i3ZlOhXf6XEAInP78fUafxc
ACByHjFlCYeLxer8pv5Yaf4/tXzW/C7fubnkbedW1nXSSi3Gdzq9sHRnP88+sfaRECvXCGzvpqiy
glUlR8Sn/x9ROe4ULMymGrzqLWnidCOV3FaySHkKb1bePNsdVLfzntnggm572r3L9e39Bmk83X8q
jkKCifv25RTU2XQRBR3G5bOKGEuLBz7jQFQ6iMdEbnYC1IrT7AwVLT2/7y2Y5Py4TOZ2nhjCNQWy
YTOl4q6xoE40oaqO7ko8TpePk7K/FFXCKmFXK7xSqZKe94HpX3XwrRhnuWDrfcM11DuTg0P8n1sz
8qg7uKCDeQOD+vzavvgjEQEKbV5hbANI7tx9jO05okcopTLoOxieIwrVmMz6xIs7P+K7mozkVk/s
rVMCCknztCiveoh/BWIedt5tujxlHs+sZPNit+dQlh77YIYnUfX5xRZTX/Iz83b+0sfGzZiLSXon
dgokSDN0o91Ly6GHWIVJcNPbrgiDMK8BGNUYxwnYdGVlCRzdYPn41kQl4C9LxZYS2iN6maeevfmR
45/ZRpkq8Z2/gDsDDWSeg1YSn26J+5NNXn3x6QT+k7dfUYLCfDeGfMT42H8ZXfUJls/bcc199hgY
jtv7q/L60bJhTvtEvc5G4AA+CPh0feR8ca/nT0kx94aSm24PfUdLdocQN8/mBSxSpbs/qkaXspCA
QPBMI+DUEqnjg39plLswBVJA0pe/0eWUIRSRjYwwqlGUwYlG+R1KhPsXQIPqeiTnr1L5RiN1X81j
i2Ss+pyEg2g/DtRY2ZHLd5h2J8cbUAxc7MRh27fbpzMWIOAnhFS6d2eTjfKcojJmoPuxSAjpKKqd
XZW4TSOnXONFEnB8BQNvew9tHhC/eAHk93qq/6WIrYgkQxv/2W4rxlem/dx4N7EXdvxtWBbyLIV2
6IPuYOIy5jZ2EDZt2Y+kKxSKwzbG81RvIrXaQyYjf04/flKMfVHp0TOKXLMk3s78Iv/ZfussWssP
9XyYtPFoRs4n+uLMxXBHv8r0TpjlwLO5a+nGlmehCS49dB7DVmMCqTqbKTBFb8AKIGty8jQHU5Fd
cPZdXE6WiWNyKElsYIhA+5/pEFDnwmgH8pdWv5R/Y5Pt5Z4ssZWZfN22sdUiiEEV+m7RR4lCjgpY
F1pJoxhffDreJQ5rIRQf1NapQPI5T+yCOv9iesmjZqtBapaElBu+hwwM9Sp7UTN8eGNoXnNrinZ6
Z5e1s+iUwHkPR7FJD39SpUufZuK+3Uc2pFE3GUH6m+AIkHfECbpNnJioNIzRuhVKkHEVjmnWkh7A
6RCuYP050xq+73VZ2NieGUCK9kooa5hqcwk1sIhI45mDFahNzUVlZggyZp31pZKQN0BNFIbk8LCC
DTlVu+Vdj9QBFVoOJGBs4STiq8hqri6CHl06wwrK4aZnU4s6g7j5u1I4mdKfRbl1MFYboxArEit3
+7A0HGYDKTPw88tsZwC5gLLH68iAYWTwVnHmGj53iulls5nvBbDOoP1pwjAhdHuvKVSKX+U28v+q
JYbetTiB9Qh5mvaETnKqkF1O72joYSzmAX1FxzYh7GRRreKj47pQH1ic+b2tRQpThQyex+EmafYQ
hGEJpSBiAgsdH7w8uY7plzPp6FuaQY55PZ3h3SCD+NxApm6QeVRqRsb7NKB4xubUMdzQtOLx2oqE
Aozla6x8rGf8o3CU++vZ+V2exKkpE0UhSCPRT4vaN0JQbYEw0jmNTg+4y0mRlGyBu/iNIzsmmF28
YMkIgq+tXo0p0ef5MNugcQYtlq7olI4UV3/OZMCoqlYaYtd6tpSJHcU/Dq4j454PMWlUAWGnuZOG
HbDnVRLwUHhx6Mw5xDBdS8FPzFRivt+8MXHIAj8NDz8fNlTLNRwO6mhSStEc4HkbFnyZjQIRKYfU
SvWowS90xfT7U6OFKs9pjuWc1DOEtV3wtW+d1ZlKThx0I8tA/bbrYAnrQCZayQjUmm1iGaNSLXp1
jd0ess5/LeAgm97uVvfm3SXw4BvkHrOwBui1mNVeaVfMtCuT5DdyDS/HyNwKq07dLMXe1xtC8d8j
RvExe6C/Ra97x11uEXewoNl6/3Fj32T9zpNQyHU8GyzD4J7Zig9NBLzY//GPcaV/u8uz9dU6YXll
NGdnTgsT6rUU8zJ8E83V1uLRc5kfqeSwmmi/1RlKf3IqD0MP95MePwxAyZzPBdXR/NiHBg9cIiyr
6i7A2MnJNrhUmg9DGQaYp14xnyclPrI5PN7Ya5h/5/b6/Oe4m3WIS46j6qZ4RUspl6OmNKZbjqMj
0TI6/ZfMJBpJso+CTpcTFYqRxQvg5JfybSQVd0SZ7OzY+Lvmr62bmt8p0cKUB83QqippsZN7m4ab
jcKNQLmqibb7w40AcAwqPj1VO9G0+VxoscfYV+WeV/vnCYy2ssLX/xT4g1I2vJ2kpM0AMfyojSNw
yMXxAWios74KmYBFK3ihObn5IIPvYsubCMW5wNg/b5cVZ2IbZT24upqea4MYldJZ1/74B/gpsxyc
QLKxImG/21UW4TI2JFuOA5p2v6CLCPiZQsYmK0/65oPKopwEfDJCIm8/c6A+kqqDoQ29MJkN14X1
yCiQ8d59qV2NzyE90f0tJ5iecakkKeoY3CwZ7sYjikjBa/f3xzKJsl8T9oALtD/9yf7rnGBZ3EXv
u/h0y73/tudFicnQNhjd09Y3K09ZBNhLdiIaVR//+xR+KJB+UYlD0gZi4uyq+hFRQiM/IDEyhjWs
BY3SlLJLJj7qrkdmKjNaz2RxaeU3+at+YzqJC0F5gcoPypPlC4m+1NIuHlmi5TSFJJEqcZPrfgL+
y/RzjO7uVul6khx4ZmA5SZe07W7VjFDDJoV7jDybwM8mqDgmlWmjdAU77DwoiKSi4cDdPByagMe1
eF7v8XaM+dIvar+mgG8VPjnxkZ5lOVz5z1vWZknK48k642wZLuS2T1PPknowqEG6yfsKg4El2RbD
4GLPXd596nTNZoSvhrc2TYr73HaYEZDj8ZMQ6FURrfFlrxXrco56nQ8SbveVcRyAQAltnSX33fyD
x2LXM5IiijMW74VjKE3Qk/OOgcCH+l1deuzELOu5EI9v71yYBAy7Po5I/2nnoXDGCYSkJ5+EHNsF
pbuVgH7gDoEk6b+vyYJv99P22Cc0aK3mqqsGMlrq/k0xLKj5Y+FdEnL+56dnDVEAxWrmKfvjp3YS
ewwUcFUDRF44VTtR6Y2acH4j4hEEQFFzQLCdbJzfjN4jC/3F93gAm8SUK98Mp6BDADyjOVUzupH2
kKq6n8z5Wv/04pqT9b+4buJbsHU558gioASNv1iNMEt5d3ptEya0AYxL5TYDRD5mirX0yOIRsNtO
qwRgEPpuVLVIO4sMJj4oWQ9DSTRkhjXFekx3RP3Gq14aCGMFU0ucvfM3eSYgJTS8hC9VjkupWgtv
YUUwHnDaxTB3KbzEW80S4gFeWea/yTP8QR9l1ho5EtksnQxvkWfgUMmcz6d/96CIUoYebUCkY+PS
amuK5T5h2y1vDMWdO8HEUKVbL2/MeFj/kBXSZEx2CQpxCEC40nToO5jTmy7ulQyeCosEk7wfvIui
/1GYwPMVAoZjfewdOop0xIhAGN57IJOQqgpCwynh4yFMES8+lWxVGJ3fmiafJutvvAKGPasElACv
KQLyLTINYXEh3AORFnJUxfXCW65lKnpoD79hkf74XlE4A7eg5GRlkSjj+v8QGpo3QJRVY83rijeN
Fg4eg9SMzlgWE8RpPmfmW7EmrQRypBdDpPtBgVZG9ZvnLhRl3pflMGbZT42aBFEJxlnLo5I049pG
vERXKDtuXGIaiLiz4VnIcbiTybzml12P5dA+IkI93PCnCVk2uEtz6SQi6Jz5u3K7/Fzsc/oQCVZn
0BRNt3sc/qJbSbFs8TyLhcyxtwZRV1Zt95FQGoabM9KNmIWHq+vvyqu1CJmQ+CGukqx3f0z9L8DZ
YbtMmyJPpIp3h5CvO64ltZrOF5GFeP6XQY8kqIWsIYffEvQwkh0VJB0/RZUBxIZKZaTLqQvUYWEf
boDCy44SMEIRTv6BnE2oSQ/X3nRAghG+dMtOobD5qDJKefBdLUCo1fDHEi2NySghxhADon9Vl/VM
ttGddBmsTuSYHd8GBH+Sble7IGAORPGpTWENxTu9LZUgCe3enlXHeXk7V0zTakbcnSy0sciicHSY
VJVa+mwDhlMPzZkGxJXDtKPbGRkdnAlbDNapuyCTrNBycVJ2qOJ14u9gXYUN+ED5F7WJkQrsapLy
x1ENQTGHcD2S7AoOCFQRMCark+Qi1vd4+iTsqGmtDwvvfXGeTugSf07Y2Bo7mioK6H2KbrRf/Dtt
s9mCkSArWSuE3IN1WRqJTqqm626xZrSvNQ0vj9WeXCDP+Un2df5v7hTLG0wXP1KXZQQFDwgCuxl9
DuFBtjPw1/Ji1r71S4pdO/223JM26yXHf2Gamc4jrthlm45dxI5tV1NZfCYtXXrzST1UIJ4OF5sG
WlqC153ECMiyC53cEpky/IlW5c/w7AnLEMlfPrdJanIw0fKL622Ww9+5TJl5+cq4XeXSmwvu7u3U
6mQLMZf2wrm8ScxLYxID4Hf0sx+ifKU4jTikfu0lTw2IJcktG99RUVofJaeVK0Y9hlNpm8mE76U+
NTF6/4ejR8QPpd77v+j6sQlEwn5I/HmGyT5X6r04ei1P0xYgLyZ5upjcXVuNTgAruOG48co7xUgy
DrvOwLg4EEe00H8m4CgonopK9dIWUClRqR+o9rf0W3dGKpnP9biuic/kx8i6tP1zsfoQhEMV1zIJ
ChyBJdUFQ96VqqpDHJZ0St/xPRU44V9Cc1PI4gIifzGOpuEV7LvTYp9tzcyByr8Ll31UfTSrOS+S
LtLHxddh7b1iO8o8rCWO09Vpuy90fxLPbQgKf43lBRfq4sk13JSJIRFQGes5PYAXIivrE3O0eHDL
fa8ZxihnJR6g+ekl11S2xkWEaUX9dF0/JFf/ddfvXObexevUHSURb9YwjnjZGigNctpixCA3JGUc
+hAAhPfz6IFDUZipLRKOOzLX40JMitZQ2xHCZSzMyxeoDkNvIyg2OYz+fqqb3fSMWH4YLkoPSM/c
jhS3BZMp3oMbuwvzfB8aiHt7554I1Dd5e8+r4zUsxGnvU5jpCXS9QlArJBzO+DSeKyQllv6kvWrQ
toBKf+0qc3wy5Pbvam25FvA9tA2Cecb7Xch9M9fn7AxgDHlajwhPcV4Hvms3QyuY6ADg4H06QwtU
7/nl9M37QoGJKd9R0fC9WiYRmRPnB7d0sjFMPbf96sC0c5XXtoy2jlI/gJBckVjUAluDxY+WTg7I
PqsoPJUBEjcwZQrtDDWShJmoGXRDMPKTCmWWk1fknwdPLqqqPpOjG6cDa2Kq0HE57kBRIwXzgguW
+QUXecHtLSscY/gsO+f4JOAGYsQqKaYMIoYahqMGAwcR45PaAR7xhZoaWPe2n3T+V61Nw/9e3HnM
ynaEwjTK1bK/1pXTSd1GgMYpPLNtG6ccMPb/W6+0U2M92188P2Dv/uiqohCFb6oCoA1k0Wkm8xgu
RILSlQmgmvlDIhmCnNDA/XoFh4liUotPrmQV32neD/sMsEi55IytTr7799sg9yiR0o391l/JGP08
QXlbY6kkWrdxAck23cpnqdrhaCe9m5ZLxvNnHeMi8ly0dGyUQSWJqtRZrYngAizdq+VN9eSGaDll
kyuCX3Jdoy2yq/DP++C1Jyac2cd7PLs5Fr0e8AgEV4oo4tTHYI/viBkhgKPs/70eEK34UGaxn1Zn
zBzcXf+pKCuppzGpi4bQvyWXRROj6JLCx50+Puq7MFdNLFnmccdDdV+m5gnQTjaxKQvOdVaszDYx
8lyI+JWoG8MNiHI/vFGyTwHT0/U8LdZGNR+6h3Tu1fhhucC+BLjXYMa7JkfFf6BYDIVcANheSP0j
p3as1DrcArLl77C1LnbLOZHhDP8kowYgWvdTDvbIJ9bZjM5A1rj9EEMP9l07EWexSGJwnq67DnQ1
kDLWIgbeDN8OqXy0IJysu+OwlfWkgyZ2skuJd/OM7xGCMQ47sKNtKNvASKRWbIGpAZCHtlP4ggs3
la5sC2l/p5cZTys/+M4z+bQdAK9qaTT3l4t17cmB8UVTFGfLE0OYtmnxRqsbahWKRj9gX15iPLyK
pkdbuQo/jGcm9JCvNtd2d3wo/V1Hg59jXgAQN9ZCFn9CDgzOg2Ml2Y2cKW8c1thd+VKfQIRtjx6+
Nu71oQzAMCY6tR3CpfTdW8lhzqDaB2N08I5PMxNXsGJHVasMJ346Tm2ICuN6KxydGRg5sgVlRqST
HEok4zVEAgi05U9f1yNLFkDYWplYNzv9gcZYjoCcs73balJAPCczrpRZmqm5SQPoIA+/g3n37xyS
/XLm6jnLk3bi2AKk3WGgD1M76H73m7dioUjSuhEBpNv39OnV7hwPAkNir5oJ2i5jEppGLl1lksWJ
vNtifJSKXrVj9UfH1LgQ/oNWNc8vSIbZfTFuR5yEqQJtjyL/+sDYJ5RiKp9+lthJKwgxKCgdDYGn
JE2d0+2KmGU7kv5NazbSyo3Mt1Ss2w/AXSvgHN7XqSZpYXoRyJ2JE1DXe8rmPPFVZUbmkfgEMzeg
y8S53L5Pw7cpLfp6t71J5coIO4tFRxrp3yR6sqiwZw5YktwkqtS9nTC/b8n2P35v+MMXJZI0kz40
ppvosoMcVeJ8CpkzNL4KFhqb8sgLI8GFuVznSzZhbZOI6l8UU8SHurEpRInmwhPQgGW/Z5Pag9gd
Sxo4uZdy/grYEvSvqO3UP0IlMe5DQtVEct4vURU0isQUJuiqE/hMFT03y36xPouXxvIxfpv3Fe0J
Q3g2Oo8PRjp1FX8VHvCLmF79pK489J1MR5mWED4CyqRAHW39C9LeD0Rz+8btELllU9z6SEv/hdjk
SAakSlDqF55IL9nXayCPsYWt60fivoVPvAJPxmRPAw8/EEf3POgQzfOhO0OieRE/Rm7idFYqHKZa
i0+evIEtBOYVvbZZedr8dAIlCMjgyYQ7i6149zSJQ+XRmxJ7e/QjRU2l+YB69HM1dL2qh3nFOWKj
VgSyz49JBeXqgCdieuwEZ45OD7cw8oGXqXChC8IhjFgB/9zL8qCNqNijTSvztpfuNX1ov2bV13Dg
ilJx2hJnx5XF6KJ8Ix7aL3LfJIWzlPHKGUJuZr5I+0nBQpKa4ElGrZkoQgug1rRu7/SOPKaYcn6q
KZv2m/CpEFdwOAAqjOo48TOu+1NTS7Iqyd8IMLeNJ4N4jjzfN7vpKXdFQhD3Ty/esnVE/MEt9q5z
WJQn5YlWQoVP2ZKE7xsGxWhoN9jfsUGlIzPoNpYVXkAGAH3ThDJB/WkTuN+xNCmiHcexYTxGpvBA
TZR7CE8JpSm7rQIMLYjxG4wdlt2CT4NufeijrLFyNMln4D/gZc0oOTW8kuyoHoaoNjrwRJBnQFp9
mLvy/mwCW0jIdG+92TNVlMSU77zq7TjpDU37tcEP1kUiGUNXX5QkMXYzkEsOoM3hbN3m7ES9xLXh
j+IqBlWDvaLOZURhevdYVDLmqeHkFwFyW47L3kDS3TeN/CydKYfJx6SYpkcUC2pfLJCxrA2KcMLO
LwIYrjsN5Isha1BGuY1o+a0qobdakndzUZjmp56eUSyKGWXQmBuVROCIeDAAs/EoSYeGVHdwcx7m
dKDOM1AkxmN9RFsDz8v73s2BFQ9ER21px8NurB8GPfl26WukGY9646MxpBYZB/PFp8lfqq4BjgtQ
2xGCmUfkB4GvcBH8vn1W8/QI6aAodpbVpL6wtQRKwjvBL33DEQDZN7oAMsV2agHtc1hB2ot+DZ4x
+z1ORVPZ7HjTnyQr6oKDrUv/8qs+howYjkWh680IIVDYuUI0yhBF1hO0RqGp4Iu0nJWRnaB6lK19
rGzq/hhiHBc5sESuTIITTngnuNOO1rY1j+R5VX5TBTgFgj6rPZZfvv9+3tBxpqmk8FU716csCM9I
q2Nu8nZIaeOexrVx2le9caso5ekDd7rRwoGbKRGb9Pg0iMaPXQJzovnLMjwOej/NN4aJwGgdi7oM
vFjhBmaZwaqABaPJxBeqGtZo3YDQ25U20/9lRMGVd0s+Ik9LcpkZYpKXdwi2RNaVfNeQ94B1NOzT
J/rj30gNHLe9g+v6AUbyiGmohb3MiH1Lc5h7PWIz8+YWukYOGpHW81EibbEm6i6kcjHtziioQLRe
uf4kHACGy9wGCMNbgfH+ZQasSPBFKL6wzOY7FVEGPFnSZYUP5vuuNLIK7XmOX5hvhKKpNitk8fr6
YN+5I6oIZGkEghY0r/hglexexrmry0qdbeoEoeHBVZwKO8xsTPw7ugi1D5PETROIUnK3bwvAZSir
0FU5zw88W7paKW5w8x6uqqh5god+bzfyfpnkGZ1MEP+7btA6WxVY9aoHAQixFe7ocJz15kFBsH20
+8Bxh6QI01+IaxN61rcOlUmadwnhENbEYMA6sOy7LTUKmVmUDDYzTHVMOT8zMHmUeHNUnVBwpaqT
BREgbRPEjRTEXb50MoZ5yvM0x7BeCTQI/+/XlU1Mm3voxVwjrOIWZXMG1BUnAnsKGgZove4J/0z8
PhtpJmUWxM0GKr/jSKCuqP5V8KjqdltdFT0Ae9IClulYlKIrXiida8Qb9rk2BnRZNOFCx1W/pNb2
hS8pzIHYVOnsKZTti3r9k/TMYh+vENhmkjnpseLTKQS70roChXbAwc1ua6YGcz5PWZdIinXMU/Mq
7al1JTvMGcoDhC/2Kfj2+eSYhm5+S1ZG8IatKnv24nIAjdMN6poaaqfyeQf1GBohTXmqd7uRJnv4
A8xSzE+X5Gg5S10/NvLEEDxgzdX6jUXSBS11tccDa0g2UICjCCY98/LwSYM+d/KWW3Cd14Inuna6
ve6CPidyptUYelCT7anixECiD3QUxOO1EP6m+lDaHbHKcPwImIbkmD/KxHI2TKf+x8WyMflJckax
JjOiEymQGZa7h4c8Hz4v4udzurYdoT+DT1w98ZoPtd7sNIoLCnPbyLDOeeVYQtj1Qw5y/W4ECuml
NgD7ZjLOKAP2+0NaNbd7Ubn3UQX692K0OV5jhnf5K/CdEwPpAg3squowm1tfBe+NR3XMWmC4wS6g
bYT9m66RRD4LBU+Zm56ykIs+O+psJ9JPAwkwvnrkseYjidPjkb23lrIRGoZjq3XZaKtdoDS1xyzg
D0CecLJFOw4vKvH4AKZfv8OvWE1+7WiVD3UwN1CezCjrYJSqSzYLXAats6YYRpoCuhYCRDqa69tn
eJLD1USa2lIwDRu1XIqdJheSuuMIrvS01J4fFwXl/zMV8KWfo7cUIKExLRB0LtB54FVL8HbrDtac
zsKyLKhVNxtkax5WHxdDZ6woFZKzH2qIgVRl1ZgKuxTztl/qFtTyqhScKYYRSNGTmLesk3O12gr/
MN0pQIOBOwjYc1XEtpAgl0sLR2MOCnfpGxcE6MBDYsNfcS5lgbifEYgLy1CxwO7D7rivF8i2cFoN
XP9QZICnGt4Q3FLTLVCL/nfmzkpTNYYGUuku93p9Ff5VZBn9KlyKVuQbRtN1FWGv9TSfgm9jjP00
PXpbRNBLqzplwDeOQUbTOFKBwlrZzai1USREEHQlcKs2zJXOzWoIL2wWUl/EW1i4WCnAbxfJldol
Pb1Fv/l9DS6ER/K3Hsp3zX6/fM2gxpEYyb5f/HywLjDJWpO3foWbJYSxhjEa9v32HRJKeLnjd46A
szRQ5mr4/dlbSUEhHYm99qb1v9s43UKltUHOi8BgroZiCp/fP4Q10Bk1NrFTjJ9YygzhkuaVEepV
UN5ncdxxtvj2LT1l5wAkZbmyHQ7cZPvrpUcRe4SFi85a+11wxEy+bjks5tZyg9Y7o5BL16FKJnLt
0ymnXjV2UyD/1z6rEcDUchyzB5qYSP30+i/53qeuO88/GJhZ90GF+L47r+aJwQjBr6uNhkGJZiEX
PFYSPmbSji7T9Y1CtIEAQSKbIoSe3kAcYCtlosRHww7FTM38RydzCHlKzawnvJjH08rEF1lLoq8D
/+WjeWTtXqAY9nQxWs8Efrn+45NUt2tvvbqtHylBCI77Lj5Z67odZyt92iFW3+EqIV1Ih2q8O6yV
IIM3zkfphHeBh2IRv0mcmbGs0ew3TAW0Wp5S8T1GcAuSKcySzPtO7wK0/DNUzHLYIncdKAknQeTK
a/ikFKs1Sxk9WeT29iUpQfKqba+wT2O+YJmsSt+2z1kzO/PXUk2SL+V+Jlf/OJAyTIYjYZBU68bf
l+KeUai/b5vexkyNPbwibuVXNAzXHBPA0ddy1kvuMYFjniTFfZ5vKpDFRmNtN/Kzk1vu1aw4Y/2D
Jx68+uL/mZu3pccnHsHE69nl8UOgPOZy/0uyYT7WDeRBRQTnaw4A91mT7MmZpNb/thrH/0ppzy8s
urUGAywimzC+qTxzB/zTJOwSV8E5W2+3iKuZ358+6oUinE7OCP/HAfOJA9VTSein71Z8559sG1WE
msTEgaTaQn0+bAMR3z6QNrqKUsT4FeXLP1+lYw5nhjgPRNBAeUSc242YKaOxeJetdWF4TlIAF2SS
VMJoYzZa75J4GZg+OansszeMOPe3bVrko9Arisx9VTyh0Vo+qILMCizsZ8YZ7wdP94chcrH4SOBz
BaTW6zv+3pbas0VMO39+Qnwd8/adSKITjHgKgZO6itzN6W4iuCbvbFJSUgSovnbpp/6y8SmRf4Br
h0Sqv1r3CnUYsbBg/sdMRwfuUpRH23Ukmkfr6DfpfnGe/U3E9Q2/A6CeiRC9LYHl6OkNWIpE2m+q
j0qBoLi8QIwXSbHIDVQ/xJQJgd94VIb79njp1AsYmWQyBex8eCJ2DnAMWZN0uFe6rB4ocivT7cLV
GvhEBIaSMguRdT6RSIi4sVU4CnsDFMCCIOc/EruJn4notU77FC13YqlJVcP40qKWZg3G2zqYo1+8
rEULxfSDkAQEJgpALQI2PxNXmA3JObDNClWtL6UBY8gCrUlkKA6clXcxqvC+mc7ttFSWx13qbRwj
Z6z/nIlusZr/0P7mw04d/lQ7VSd6/lSt5ijGMTlkCRrOMBke0joXW5kWn57UZwYItXsrwJpt6mkH
XBZ/L90D/vdb5pnDNiyFRckf8oXG/la1YM/UACLCkFeBNSYhjON7jKB7AxwMU27KHhr5kYo3WOFh
WOJ7TtCGQM0wueHn7QDa9FBrqi1+Ety5QYuTCd8ArNQkH5C7FYXOhkXzpSK8kko3+9nZOPNrl9sC
HGWa+Ynollw7LffDD4fuewc5iBNSy8tsFpHF8otviNbMHsY1WwABk2udNUMb/lPDmf/dydMNaE47
Ox+WkAce4iHQ208yJpN4GdR6zVNctKvkZGks7fHyZUDVPe6nvQprYsJMp0Lj9I2lU+qjUqMeTVNE
dWaDsGkTxeEMXGdCC8hmZ8l3Pa6lTD8sDKIldlNOr/f9s/EoC/hFzolHof/uPc8ptXMHkWcz8W3H
bzTqfOFI7ROTI3jmmZRDT4QFOl40iBnlKwsYZGCRjWy14zmlgu2CfZwrNffvcsjyrHosUV1kA6lh
UGTZHRpuc9q9wCBrSpBlLYHJJZYVHff44M/fFFYfU2R/vegYH/CzB65yCTUuhhPe5ATvzOYf3Kii
ywZdSSLcxusT5ujN4Edr356W4Paixcm1fFLvh7NpXlUZ/oeQxtwZTDDySwDD2yrNF4Cz8k8C0OvE
yomzWy/4GSCt9wBhWOFeWJvLEsJadKu3GaKenh7wpED48yqVuz4SMmN8nUn48THd7uKACyQhVfqV
azOOs8PHkbfy6eq2zdc60XYIRwyrsWbkRrRHI90eyuTb9oRtIhC2iBx5CvcyN44ChgkfydWVGin5
Ljm387lJbeeRQD/rn703we4oZmjBto4w7qv03eMJ/DIqc/flZ5FmxF6dr/Kf/AlprAulhBSwAHJd
tm3+j8+Zy73p+HlU6G1V98xpb6tmlOMGyLUA1iuCfhsSTRu8QG4Mp3pUaAYEZN6iLePXYrQ36YH9
EOmObFI4xMndednEbqWdP39irXRN04rVUR6enpQNS8NAck+c28NObwc6qugazIFmwDtRXXBMN6SH
CG66e06s/4etKZ3XPr+r3gXntdQ3ewEThEx6XbSCOrJH60YaCzcbvdYjUNdm3wPj8JrOyr4u8M+h
sibZIqG1NolGYluiLe7vM5LKEhF++6ywwYUFQIwiwo1qq7OfYFYNYvo0KqdBWYQa/LcyZmFt0bsR
5QgvFGCQlSN7AMVoYvOq0wZnPiPLzB0MKwKnBECSGbur4+4rlosHtDvwFlzreKGxgevsjSesLqoP
h4F7QbjesA2z8bezXZj4PuvG1QCGX+yjfQKDVmoksL3FmhwCPJFJCfNpBBk1N6g/7JbH5U+Ti30u
UFI38OHkt5Cu79tDLfqPESkpCAvdqVcYbCehZtD00puuhh5jFFDPDykK4O+X4LQXUbZMvM0TmYoB
MXHiT6puWxhZklhSPQGtczto427pYMHVzYGCLa4n5vY/DOps8l3TKg/K+SYIiwNExcXczqAZDet8
DsPqXLyLVRc8b+/eRhWDY5hYS5NZ39MkwEdVV2w5W3yXDOI+rN4645vnI0Ktdsn/Iu5q6MBeNyrZ
P18fqrOIHddfE1TS1Y9jNUo7b+AvJJ+tn9viIJ/Xq1MAO1gGn8BuiLLsuZw+j4XXyF23VHyD6gKk
IXjJDAH1Upvi/MGYXcMrZTIsAqb9RzPyiOpy0uM5R/VFWxOC/cnmk+iTeNYbuHvO1hNmv41+Qy0l
/Q0IJe70e3o8qq9ZHkk01lBUU7l+v8RrgGUwmE3MQfpvrYW4HNUAtTCQF6Szgcw94u8KBVybWQw7
whrBP1z+l4nWvdaVF7sLllOy1dSthO+4XT2eoy0CSw7KLNELSR+jd3MlwArF9fgbqbM7ourCosFx
0dIZsY14eQr8lHAOi38MrrBlOrTbT91I/UGwwI0+OI11U+6PqGMzTmyp6d/XZUQX6zSxWLGjGpUj
ZCXjaUJRSgZRJzAT4OcUAntzGhKvzX9VzW69bwLbSngi5dZfWEFkwmRMp28Ywg0ItOuNj2dTeUaO
stZHmcbiOOibznO91tMorqNvwdkwotqir1/ND6UvmClL+Qc74PCKWzlYGxQ2NOD7tQWngAscz7y8
rYe7zjTaUqs/ZWAPXs2v1k2qNVjMCieHl+VauuweCATCd7C1K6GeihoXS1CGdeIINTcIHjh6+Dre
RaWTpKXoEOLzSHjMWS72+xS19U7xgvUYBrdhvgjmXknMfjS/Y4wf9ZgrfL4g3/zfYsDVCxHs5IE/
906Z1ijVRsa2ea/rBU6R+V1nNogaA9/dsEdrBvb8znUNSQqs+aIxgOXeAUMqymKtZCjfiHi/D5Ee
5IzDEJb6tjJcBBmsl0KJB1huIfOd6Ln//wW2AGw0ZQvyTbRVJFU9hZq57qKBqRSfm0T2VCkPWIxf
1TUcFbS+RNHTxW7ukUo65TxSPI9dELmLPrzn9ZO0vEl8xGjKLBlKtRRTLy0ZAKTnSibaCFJQkD7i
CSxH1zTBPBZVKznRxzdftrjiwpe5JU3G5m1+xGs7NPQUYW9pEZQai60RgiYlvG0S6Wunw0ue7C4l
u/b+yA5CDT7bj8iqVb6uefEYdzw6u2uy7Oz6ZJ95pde+1mjMUebOrmTVbHZ5yzloKZYIivV30ngJ
VUhwLXDSrmEyIyAlKMVcoILTcdxd3F4jCqVNNdtFzXDWfsekGuwPmf0vdne0/arKuYr4OVHGDaVi
lom4bg8mpIVJCe9WaDKxRKW6HS5a0vSr592RGmK/YneURCq4zFO9i7qBdtNyMOMRB542hbyy2QTL
QGTHHsR2O8DeA6a5zUg9sxa/KQXwZonL3OuwCnbDWyfilBM0rJxBsQj2IAXE1cjPgpenebeur2bg
CZKnXWJcpk4kKy5ps0GdmfxKBKyMg6oHMGRN5zgOpGgcbHYXlj24fPlOHbTfXxgfufHpSGTcJpfH
Gbgny5CurZgCLFANQ9CeW3CN1BrMJaeGPRqaWgE/7emWe3CKX/6/4+yY+Q7r2jM8qyc3jmMXLFYO
mBW06Ks1Bpm16sowCUDoro7gpFot+TDV25dmp0h5u5uhkH8AhD08FWstRzEo/SR2JhDbtUUVsbrr
iY3WAAUsBPfOJEuALpebtcSnNMwywdSL+5nhqleiEdu9Bx1ocO90ITXFFqZkti1eikMI22/kin3l
O2ePtpGrzusQTgstT9veUx4ygKBdpbYcbjSmkORoHwooPKG7OUSuwu/j1U/jEmsNXvrcOF5mcmpm
Ld+xqOT2s0TFrAJR4i7o9C5mdih6Q4zQ0OJCn/x5jsZ3G/uDPB7xNEfms/Ndc2C8/9qFJjh1XI8D
MQ83yPjNrRCqt+7zQKwwp920+TgiHo9cjlYTNfiEI0O7s9rS1Jj49WOhZqqSmwUXLnS5CVW9eci/
uw5u7lVaO2eRCEm4A/DO/26xtuNUjAioqIb/bc0YXS+FPOP4qfS1Hh5xNj/dgpsyFCZlSSpFOtPY
AIPHvtAAlmQk4kCC//y82X4v9zHHRpefV08Aj8i5ddYvMQJ+KO6TtC+w75FrzSM701h6WF4YM3Tk
WAewXPACeH8pdrtv5mi22va3oB4fqmUkmLIMbzmAJDp4zktUE2E40yTY1VIU+FXk0aky+uM5LspW
t5lF+vnX9Br8OF+lx8oYdwIpUnGPAOAhJN3t8E1OjyfUg6b3rXjMBShJYehgUmoUFknJRwrpxOW2
yvOU9v7Xew1MyljkK3Ft3zIaQW+Sgl5dGakKI3jECWymsXT6Yn8o5RHZx1pkgEaJUP0gfpSK6ys9
Ypiow9RU03hkB0TbK4VJr/bSyIHuhlGAZM+M3CbavR6KhAQT2QxzLmm8nDZdDdfWN6XFjETLTdoE
4jcqYjIWGWdXsLtTOo2s0MVfSDk0QEbuxxLnGxNQN+5PlFX3K3bK5xaZp8nSI+MrgDrc9rdHQdBy
jzoN+i9dT3dIEnJ0rm1NGLeRkjQGMc31BJnuYW+5Ca1DxKlV7lRJIKt/DRD2lq2wF8sN6h2z5jyc
KMUCSAh8/9K9d9TMIsMhll+6iczfWOrr6uY4t+hsO4FuZCr++bwtCBlhkm0v94KFIh7u/iNHXhAD
cA+3hWZaiD11WnT5O0t2oYE3qbhGqOJ8vSQC879hFQb7petN+U2dckVZdaD07SeGBK9SfTZW4CUR
KABEtChruS+VNYGDIQVskOd+m3yHqJJn80a+j0kH526aFj47mvPUjiEK68TbYaslIPhz+8k7lr0j
OSD96wr4Dm9Jae8Ni319SqhnS6qGeKGfFyRL6HBP/d6fxGqynvQjFF6byUHBKvIqfKtch2cC+6Pk
O5lzsIb7skD1v9RhxLaT6WWXfYf7f5+G9SDtkaPXeBvRCPhuqsYAk9AquisQL9kGMGOiebaHl0MS
BEPzNIbxTt9jvBte6MkS4U3FsAfWphYUvew0YtAzbjNywsbmTgpZJ6vWloD27tz9h0WlQsYXKcC5
16O2RZLtq1rFScIND1FJBz3H1TLefaMlYuux5rqgy/hy5G3duQSV9XuJjl3wiJK+RzFC2os3tfxe
99Jlb77KGloezciwrOnyh0Ih4prpwI+l/6AnpK3WVixmpALVCohwQRhYFkKBJKbjjESN/7bZ3ZMi
wtN2UAEE+6chme1VoXhaJsXls1O2aM6EuLhaxWUIsOBV0A/J/tmrlvGoOTiTjUxMLIXSy8a4H5lG
4jUckNAexrD+VvR3BDsGQISwW1wIEAvawdvGtkrv3KsSDUJ3M+9ATgDvwWj4xmWGBoYNvrVG+RSk
hcVZTU3rrHuAmK/IFQM5ibk0OHqN3/9J93znIEzKTzAV8hjJC0pVY6WR1ZiXWeo5ahQAcYXP7hZH
IJK4MCUFBpYRO0BxvcJOpPjC16de+jZZMWjLdMNTqaRj0cv3D/6S6q69RNTyFf5kbr3oaTwCJUoD
JJ7VY3vaKuKzyWCIbckd4swcbW3qg41txlp6vPGf+VrWqoa19P8+z0uU+gISCc7HBmDrW3b4ZXVC
xOFi95WpSpNygTLrHscyDEwNkDkLNX7ZKd14Uaj80XRupm+kQ0s19wl65nfsvTcqF7pErJK8AbwW
TVSoxHVh/81Jix9O8Oysnd8ET/4DLYWxaCZyrtAGt4ybmU7ekwgibjwR2mgHIVC7pl0tgf2G/LCK
+w+xzvP5hm2BYpI6iK8TR6So45epSLHtUpoKp9tsmZcK3MuRVbVFRqV/Hz67IrgtBZT+vKMqiixk
TZjDHuugPjZ+5cfehtbxygbTKCSSF4fbE0sXMoYazBihL8/WTsXtoWrb5mUmxqnKLlryypVZBQqm
U8u1EU+HVhPC+np60Tvsaa+4Q/n5VcbDgo5aHGNHWwo7Mw8v+4agtCQDID8J9LZqW0/qZXtmiwBg
KQmTwyIFG5EyhLQSOfmwzvthsHP77beGniyu0XGSQoqQlWuO+mb4sVqaX/nH+rX7HxfnV/kpOvMG
xCkF5QsVi2EGIt2ZvIuBDfxR6yXeoR3jnHa9XBsMoPNrlf0fniypzxcTX5nM5pOkOsjfgQF5j+2C
xTMMnkvegHUiQMcpNM2N8X0b6/mQfYJ9k7qwKIcEPYPmofIQTHQZO2kpenbRm5pK1CIQ9FubE/W/
0cneVF3KOHVB2fiTY3jTv7/XGkI4dKmaOU49+QruQHDXhTpkfRDlbsJx1jahAIfhJm8Rn/PiR6uc
Y0wRUO9nUcM9gbgHP8f6EMDCIDP0VIU6CTDLVgN85BZ0ziYj5Z4ZrY6ALRzhbLjzDoyMrSlM/UUq
s3kYequG9lKtTKqijBjjoEwtuNwVwySYhJCBXXXUjJz8K0diCWAKZGw+uZwHGSh7tp3u6H0I8H2s
qycasM+QeERj6EBFRKpUKRa4S/2llRRQ7TQFYswDFpMv//Y2nq1GazHKJylDn67gczE5GhzGM5+o
ZMNwqgwGJ+8D7MCXVaMHqDH6Y00OOpSJHr7TuMk8E0sYHKDLBU3z8eZMd9dBtWlcQn1YRPCjII1u
LeQgIxv+PSU+WI9mN+cgpU4m9ATUuPw9K00zMwQJBglUb8fhG+GwSm8iwXl6ZWgrCKp6l2uliGja
RHZJt4vtCy+FGAOb5eUCMngQyJPN8zj/yTbYrTqUOvxVtJqEy4VwGib1LqDIvtKEfnH13rnPOOC7
/cRgCOT4IsvNybdGVxNlhEkwZqcix5ZWxNqP0fCPalUlD48l5b+d7oHumomL8kHnFD/pdwqJyTJa
dFAGHZs6HHYtDzqXfNWnZQrqvdQ/Y1jdO3MW8Pfz46q7E91YX6IJ1TCbv2NJa6bLe+XyF7VKs4X6
+qQhWbDTFSkPPwfEOCyollVudmxw+THqWc7yH/TWrQJ5qPiPIRY9hTXd/p58rqaRnJrBXfRsbeoe
dCKVOEx8z1a3ZKwgQcscFpmRRecafZPdSCSnXnfowZtXUW3biwfxYUmstwElZWmnI9QDj5dwjlGU
cNx/dLvciYU8ZwaIGKKbD1ZgcLQr0ivshhxAoYORM807L+2HIXL4I6Uuqqh/piWyfh+oIygp4p9L
wRqYo6uYkW3oEGRV36BaiLdDLdqwrITOY1eV6Q25MrMg49ynijMf58dPier0C6BjHw9HUKnYlGq0
VBBEPlft/OFCXH/ChHHpDvrQgAzWBityBH3UXw/QyL4qZMQCfydb6zXEhg+uCfVmleae/F4n9TVk
QKRarfdX0R/wbpCk0robNfRfg3jVJU9gQq4NfbfMJcTYTn/nK/P5aX0EPatx6EqEnk61keiFRZGr
OFnohOHMPCBfcm0ChmoQHDMDh9UvbjF6uqMmln5MApH1ybHyXgj9/0ANFBWnSIsdLjpCoD3tYLkv
bOkhH/o74GAxgyeDd7gso62njhXhNoZlBDD/uepFFH8BarqL5nsbJbXSD8aa/WjFN7AzAa62xcW/
TnOQCnMQ81C42F9/9TwSUJV+VbzJH+k59RDJnUuGkvn0r35NH9hpXUN46VPQSOPNRTbEWbEEz+cY
wn3IK0oQxR6fvJUfctMvz4f0TVYo7mXzrwDc3s8njBvv+Fs2DhhBi72PUik+7v0b1Pj2f5JXoPZF
SHeIvV9pV4Q52tZdv3ewNpNhTSghRFIXAgGTk7nIq2jvqWkmA1q1EioFAnrNQB8x7fiU3VCI/Quj
Cd6GJBCdZSUULbzO9F53hi/vEmBM49yC9wZKum+QY+JxxdhpYyFWBIMFlSmqQmI659tygNFrjiE7
QhpQc9VzPualjtlOJMJeul5XPUz5Ie/xKAkBPrKuWyEoYc7rKa8fS5IUOLOxqEcWLsm5WwrzO6Fr
h6Zx683AiCSbMbNQ9iks72beY7Ohn3mw7d0YsGd/jsR62us9OOGZXzhhdymBi9jN2GQjRm29kzrR
VTbi4clm/ERy+eC26b5xIHdXfqA0GTgY4smNK9Jxlsb2PPIFvhO/fkdibXT8jRoync9j7jccBwgf
Mwnuw4UTWQR7xfd3LH1tgpTxEZtib7VZj/Mr/uaHo8HQZZhwxLs/uj7hgqT/j/oh1+SmfObCwhrQ
irFnFOxSimfrfbPCPREDG2z0ojnuq7qrDqeqJ532lqUTLKrs9BfipPDsRUWn22qvB4fo6/jsEjaa
LpkGze8ge4ttMOG+hr7PIOvN30OW568JcYDaHyui9vSk8lbW9YNHb+XC+xsnl9Yvk9k5g5AInA4Y
Og2xdVsft5sQ3Ef/egpFyRvBXZHZ/R6zDuM77F+yB+jD84hAhiiKthPOv/6z0OfOF4hiWXu1/xlq
g23BAl2AM84JQnSFo77TgWA+TMhIds7ImkNY3YljGDVqaDW6OJEokrwrkeB+a9iM+vkH75BAu0ZX
0bhBWVhs1yNyo7JWXdzoZlXngZ/wi7+6o1CHeoaR0W4QoWI8rIkpFcUIwzuDosQo0cGvwDtOT7PP
NF5d8/9jF4PLKI3kqH8BRcqkhQpkqLJQdeuX1lMkZV3nNMqv+Aksz5Z98wvhaz070M1WMqzpkRk8
9OG/kLox7za8kdVsiTKQZLZGRU7fCRDQelOhFrHOhIJgonIVWaJT9KLIqc1Ry0CcZ1LjsibnX4NE
D2t5dggmXw5GRNSAdJqqHXclahjEhVnq3wd42rLT1KJF9hiyzUy7wYokgfydypctthBsZKqOKedS
6FokA6fmPv28ZDd5FvE9TFKd59Mu1mw0c79p1s8HyzrS/boEjxdQkA4ROmt2kIHpak8pEjp1zMhI
ZStzZIj7Qd2xiNQqZRK8Mt8XUHLMe9BT/aMqN/qTKAS1atqCbX0G+P4PGlr+eSQqHB9OnyORkbDu
nDrmxsA1G2ErelnhhoHmpSmdSD5bNucA7dQDruhEmtITrKDmSRE9IfNuMzaarJQytZAXIQcMMTdE
bCU6MY/i2wX+fDjo3PtDRpuR7Aa3wQh+MOBimEqLsWXbqLcLl4GbFCLy/aKFRtq88vRxr8bwUMWZ
+J6qhBhjVp15jfwc9AIVGp3yZwytokDT09BZ47X0GM/DZhrBNm+mNqDuSSCzGYHfXB9f7+XUKYLR
H53pNGP2wXulTMtVLbkRFX1kC2B5DZTVpg1IEPLXUg7BVpgiJH+lLmuYK6v5LgCc8PEQ4J7p7LY6
fyODufloT7G3ct/Niqsu3x4BozOkQ0UO/iuYq+2z/apGN2G5bc9PLzi7vPtf406fPpmkEAXvXn22
YEdhQENZmBYR79yMUXZ57PNKaV4HYpqSbbuMryr9nfBqW/0zD7h1BOKwZKuP9eDO0t2YgGyKv0Bm
Kg4RNQx7wKQCdmUVC1bIUY/w2SrCV3Y4iROkrX7Jm347lS4TA6Y0k35Eg3eqNQdRteRTmThrWY5Q
EHJuBVnjU4/q0WTG46l8Fv7runFgr+VysBVZ+hHDh67aOqLGtaOM0ahQ9WP0RvJu5g+fHXBGz4if
yv3K8HZEr+R+PzoVIu23iLC8M4bxoXwjh0mjUyeJOmeNhJqs1GIOtSKsJdmOjOi3Q4AD0EH5e6Wz
Y1gQ3eiUAlPInUCJT7cNOKgvc07Yy8GnwOnBCCp4PczKRdr126xmX+M0udLf8KuQUI7UAcoT9h/w
YzesQpX6qkeN1jH+G82KKQ3s91AkAJP2CcqGMTHqXP+K3Xv9wFna3E5Afg36Vf/9JIP61JKlGD3D
W81sPDuRYPIcnpChgPHk8uXujySoUxn233Rp+8q4jNuhuDGNblbFnstWI8PUiC6z0zLD3kuPQhgc
GshPaRT/jGJNNNfG+BU7PEJN2MXxwSZO+6nFn7WVtTL23ra41cbNEALQPIH6LGFf6ptJfV5AL/Ig
mLuKwCBp2s7hg43TC9GMU23kVaNBtqS1EbMv6b1A/8gOC5UEG4T+hmGpNm77EK3m7W3wWAD+opyq
3ybaN0cydGyQSCXj/DKxs8cn2LYlKMkULrEWsqRMGiZ0XiOdsyH5qaK5bzTJ6RTogw+CU8MhoGyQ
Xe2BhUtnmoTgzuhAbmpfppyIdtd/6AVItISbQM/7TNN3FbLPh6ZXp/z20tqlLFwg8rCTioaGikZT
aUw/UVUMPiRQ2Xz0k+pm0cnebk1Jpnv+DnukhGlz9hpzb7G/qsz512US1R6O1KZXSL6rGz7glc8M
rO4l79Av5oOXcR17ZeG/w+jL06ZK6QpjvMZv/agbBKk9x9H1Ikh8SDU9TNPy5JFpNVGD3Sb8OOLc
07hOIBBPATEYoIStGMiv4ufXGWGTPi6Kxovwe5eapdiTiyVDoDFc96ogFhSn9ff726Sm1Au/801o
cqJ6SptJmw78GzBA9rWGQTEFhVZgAqhCrb14o0DhJI8UG8XEGSeJRe9Mu2czXlE9LibURD/uRnh3
o2oIqmR1vUBemCOSCDn22Al7FoTwFfoiynfr4XxoXihlUerXjSqYJBbBXah+C+VDbRqfvz+BgEAH
Yr5DdwoeP0KIwiw4oY91UynZdq6XKYtpujnP2w7bwX31NQR3c6MCrPvGY8ibgSGmtwSI4StDhmKZ
AI5aP8cUVuMzwcPjoGPRr9wbm2S0areT/RqMPGsq4Fa8TJabRMdptUEHczKlEe7mOuPKVHL+TaZU
QhWWzsBW2wJkS2wFm+yM378szm4RBpj9xT91WskFOCtfGI6tPpq4kiwJJspDzNN2hXKsX9GO7UQc
0qe2BIbofsHTGGCyZ29gZQVxMsQ3TsiHHPoE/6UGfrki7WQiusRA4sVCnbn47nfS5VvKEUXCe67a
7Q347zPgkOLANc7ZDfQu+2bgz54vTJLxHBcutEErdC9bWoUz6YVFvMFIlVVz1tQJggJRJ7+xFh2d
scBz2sPiZWpDL4GdiZROnH1SGULYZeq3v2gLhtaKItkiZlXgtcMWVioBckFRMVtYVXq+HKcADE9T
ICocIQ1+ajDdjLAdJys0WJVPjosVgAqrFhKF4Hj/ooqjVexLKQc75oEfe64wQhasb8KZXmsRuVWW
Ex0t6c3Nu4ZD7s9XF1/zC8DbMDkucxBYUgaJ9hL0VyhxstD13rWY38gYN4fVLuL+x/tJ2JhY+vw3
IVZdMf3JSxXOYOKpow3bJBpctraFXmy38JgsJ4swwikZ+ikNJRyZIZPSCBHEHM7l61ubQmMOBQjw
AQZe3yIbCX4HBMSRjj4nwlKQ2TuAeL6MszWxsDurIhyTmXPxkCA5PkfmgQqVI1VdxdWqaZ30BxaG
D0Y5jcAR8U60Z+kQeEZEfoCWHo6ar2RPEkTrt9rcJNwMTMbQ+VdEuY/mqoKIDahkeQy6ycWpcVk9
yBmew8nEJc8dzXYvZH/XtXY58a93VJGVhNYFCMPgCFv3LJytT1RQBpIMdl/mQJhE+A0Tm9v340zY
XLo2294kl2YL2+CV9rvwxJ9XwR2X2iAHl8Z4qUS0hPSNCqOV96LOEkFlrqlMhsU0YD6MecgWkR0q
0lDuUsC8tCgxowRSPCY8GKuK3ZypXh1P3uI5MzwRlNmHh2JzO3P9R6Sten3rPX+ol5SXfD0dG+ya
t2buREyKsKwG0uapJVcfV/F/xiXaYcmuRz3PIuysQTEfKiA87Zl448KcQtIHPD/OOx5i65xyT56L
EW2YPiNSdWDqZMLJOc5ud0nwkZwfwhr0rZeJXq3Tiy23YwbzP0X/H3KB5orGelKulec0dzB0zpow
y+L75v0b41pvpDjXEFPHpVD7wq6MTxVU++Jvqdn5gRdFoILzs4/Y7fCXpEdckjvJJ0ebP9wg+JfI
DuFiS/zqpAh9SMQOVBZcTB5gQgzs2mp8rgt/qnNym9ulrz0Rqwz/jpEol+Qvi8MVw5ggvA3UDeMv
quXmE+pntDPQcJU8GD9OsMaS5630aU+IdICzYT06niVbUdszAm3VXtoeukK+y/tEx/TeU+DVo06l
PKONo4fAhEWDZGAMRE5YPVc5dllERoEGVhsYqumd7aLi8hdS+jX7TwkAZ+ybmlO4DTUqcQr7doU8
+0E+8et/if1EQNC0iQQ26vMREiZil1urJ+64GRHtApMlqihsQDMRc6IJoKMBM0zi/02Y32t7GviI
3tnUzkbemrFSKnxfAl13jQBkAHc7qmRaaXMe9YAZPsreDL9WqbzTdOY3kKt0P548ExYS6IjrK7rh
SCflNTOtF7UH7V52c36I8G7SrTRIFyjM+jVyucfx6j8PHt3wLxesybuYZlnUiQ+Zm21vDmVKtd28
eaJ0QSOV1hAWzYPPIDLPjHRZSSgFsAf/xi1QAkJ+iitgX3FVaZQ48q/KMkieTuGhmrkk8JMV4Oop
7rDBI898Ud4W3XcjUHmxQ1BLvJfVMjpod3kEQP3MVpSzUqW5ahwHsELcMvmnwQqx9EXNBeOTupbK
t3/DbYA/KQNwJ5F5ycVAPObY+HUf4e1LVhSPJX4yB2qMF15MdwriPFvs2JLlX694DR3myZ2uAhUm
dHKVAWGzqqNKknJdXxJh7W1KDxRCbURkEZFrYf6cFdlWEKxLBKd5qxo54Fxlb+Cu3+jzdMiX9yU5
y47IeS78Au1jBbJJT9morHF7rdroA1HTqmNyW/JtFlVvN4oiafPXoEFlvCdhNMsIYcSdK0hkgjRz
TQRmXMr2WvBV6TlequHuJM+F/UEHIzg+9NAlols39/Vtehc/8vg/fscL30kI2+rhuUoJSp4ypWy1
/YbievekQz2UQLENQ0s7jFhbGyQSsFGD+MyXBT0N9Oqw90FJ9q1y1nxs4K2M1Zl4tdOenJpXBHYq
ikLiLC4bZlERbFoosiqcofGdN4PvBWoJBztyBjIuaV03jw+diz4immdzq37RnhNV4PNVK8PUG8OQ
pnq2VMcju7ITYqAJ0rTGlfpqT/jHL6ACKsKdx7JTXUixnOTU+s+e7EiuSamaNfWDIcL5wJJ44724
ty+E9RIrPkwkwBit9T9RRJYYzRl3gYsOV81Kx3N8qd53AASI+MxGidXZhxAZoX/b+NRCRsDBkvQ8
1CtcweMvmKt5PEfKK0oPlwrCnHt+buzBcPb0BpywZ7g8tOQnmnLjGFYE2Oi0UC2Nckfy7GEphW5j
V9ZXbUlQlth39UyVo8MQ5lGOcftIU3frh73A7+/4U5Kntvt1ciSZH+QB4zqfXj/uw9Zbq5/bjCsT
dQLW9eHihfvsMKYV2zOmuO+Tu6AXLabrGpaduWyLt/Nl+nw6PPcrLGTmbZ6jWROSGn77TQGML0c2
pT5vjDam1cqPsYDsLOKekJsOTXScN4IUfMGtxGdT+HEybknH9V27HmBH1l2unw+88mUHBVB6W5Gb
pQ2I6YigtmS6Hd99kxTFc4srZ/StDInW0WnK9h6iP/uGU3p8aRyWOrq+DerYSMMAQbE9rLrwSRkv
zwci8D8QkUbPxtQO081+w4cdTTbscNPA24i/f/UT6HzZA/NR1glSj9BBc60XJYSL97c/ywfFjrkO
1Of4VGLfys5CYWtm9+PwuiCC8VZ3GNT+8KzVrgKpdXXgBGv1DrF7zX+uq8N0cotbgqf2fI1Kmaru
J4bWcVm7rn50ynsrgei82jHYsBAqz0bFMAjc51o/mB2La5El8iZGa1mT08qaMO5uh6Y9aoXGxz9V
obKPQDbl5yBIzhB63O8dEYV++zXS/rYKnB5AoaX3q/MfbJAQLZF6yxX8dBz9QRQKU7Ilu+8/e7vx
79CaT7UCWymLfbyoT4B0+Rl4nHaNBNzqEQ5eV+9hyP6zs3Mti9iKDL+JvPmlzGSIg6bN03QWKWKB
vglTB4TxTm4bekHQL7ZO384RJQv3mIBrl6qB1iqDW8fvOFIzYwcmVBRkZa10PapcfbPZu7KS2ka0
X/cGxrrrFMiiTR26O/W8sL2jRCmaIlzbZj523qWrlTn+fXNzA/sQ6/9lAsAvovi1pfcc5T0REUQj
eZcpStehKf9DjaAAV8DlM34MFC5sbERawfhpncVXZdG9ZGKWPb9GdFnEh/2/R1/GAwnRbyiH8xvj
fG2UxvhElxUQXqTohxC3lfKy7Kh1y13qEUtdek+WT4JkZA+fn3aNXfxRSS72BlzrW4u2hX8+i8cy
oiWjZu370wPD/xcI7IW3a/bAimmgx/PksXZ0Q3Jc+Wf12tXzjaiJjJAeRZ4fSRSBJPBF59nDSDB0
oWpfaQ7rECadVuiaCdVKnGRWH16kAPYRhEgBknwUtd2+YIbaanQIiQl4q/xnuMEd1jbPdbyeWEjg
Zl7yFOALnA2QPKGhZTHRk5kKM72khvz8T9m7J8OkOciFOxL/kJZqoZt2t0g/7YGNwGhdDqjorRNS
/5DM27szZK+OOgZOOGm6eUHs6ZCf+nuCb55V3oRU27t1jN4VWXmVL5i+EGjzBHXRH0QshBbrIAYD
GGu3xRE9Pl6uo02Nzu0NYvkD4rf7Ts2ykkZiR5cDOIVnEfkcI2KhAPRJ8nuppwUaUPR4uhlDBAGT
nbSRk68D/UY2gFKtDTUU14QdssfhByDCx588R3EORj7EDzJosCdaWxwWsvJ0R58Gd4g0G0QAMoyG
PRajCTRo4t1gIw030m1TMl/PN5BabfUspEiOHh+kfHILEUgvmofOshahBQI/8MgoIxODOqmAVgHe
ufxcl0MwCRm3ildq/DjxsqfHkOlvY1XmhuhaY63cV/HzxUL91dFAB6phpRc3jRt14ix1p1SLNAmq
Mo48J0vebFs+RTu+e5Ie5hy0FgG+VZkuzSORGUVUNCo7uXIT3DiwEv8/Ag3ocAPt0aD3tqpavNNG
MH9CzAeod45Fpdi5BsLXah3/K4mAfCU3m+wNj3X8PwftdbdYE92lecBlYFaRJb+2DkrUjwNV+6PI
z53fz2uPauPGqQcg2hXiMPchCs+/kX3ooo5tlSLoUGoPn3t6SpK2RnCwmFF9Ng2kKvXA0NYjo6Mq
qiqeiE+EOtqIfqkbhiGJGiWmDZ7dzWRJY+4vwfPYU5scsn7qYvVOolEolPCpWdz9EINvl2SkwuQa
dw3ozDcufF8l0GsvOHyFQDGKIFnsOxS6Lvxrdqy8bpxk9gqyD3gRGew3FKCRps5X33TXNwFQhYI3
mUbBx2Bm9OoIl31S57pR17lj+xaPKjpGmImRlnwxr9S2yb737Uj0qo4/KwJO1GoqWGymBap6f5wk
FXB22mjwo0iFF9FLngEDC490hkesOA9oeeXTaBW3Ze2SYH2xto4P4M5DuqU6Fqk8Tp2hU+2ECK7a
nIoULOUk06nlKz/1kjrQdfrYPr17fAoATVLYd5cBFQWVw7AnPQ/vfqG6lo1VWTtdyjq7fs2p+rIn
w49J3VbX+S/x3w6TxL9xeMiuzY5beJl1chJ1hGNOi4ZcFzG7enPhMzZVPINJ3X1Xbt5TsA4YvBXe
w4QEXhaIHZPXtyXVG2mT2It9reP9fVS/3uSQ3Rjulg//73ZNXVMNYOtAOCQg93Ib+ij+jBOnd8b9
ttO8FimfAFvAwfXhRkdsKy8a3wo599MyjOjzF1uUBuQ6OQpb6XEAOFVxBrxJTjK7nlnmoFKMAgGv
dxinRZRWwPkQuFwWpyUJ9Kt4/DZMehAMFaoqfsw1q5a0ZUCi4SKtTfDxpR6d23pja+LxPc0brQT5
7lJBnpl0UQpdoVizhGG4rbRpgs1dASeehZLsMFj7ihnRv36wMW2RFoJ9+WaN93pc1CW+OOrGuZr2
gKi5fhACqNSror1uQsuIO9tKaX2iSCNc5/zZuF5wfv1pYkG6zuyw4aGwH+In8LfojJH58vNhaPBh
2caZwKhJQo266hjFnfni++tnkWgKP27TZRTJovsSYH9gzGxWAsCRGDoju69lAFKLkuptGhUbl8v/
ghUpz5DP/04MTLA9zRSsLhhZe8KeJvEHD6LLGRHvIjYjrmwTU7NWV32bMPVv68PsCEbBszxIYqw8
Jv1RneLH4QG4TIMJUz2FLPp+AiyA8oHNReNk9Pa9nvAX3rR6yXHeB1QCi/WmXHDR5dHaaiw7btb7
cRKHZmRF5fyZOuLTPu61GtUGFaVOihypL3abhuAIZq966PPV7RI5NRM1bOeYbe7zsw9Hj86NiiiW
P8uEknqaQQr7tJhIzEqKvf35RJEzbRi4IcrgTYLgBjn752cjQiQSsTkWhdCk6SyjsrqIJ5KNH3pf
a+q/9M4qC4MsplBN6Y7OdAyQMyimigmZICKh4C4a0F1a+KxEajEkUhDLYdyVyQCTN61iFJRi6Fux
0dQnjGi2nwZJG62GkNmk29Q0dz2qX2H18+deT/fsomZ/Unt7KpWM+ZpI3OubXNK0UacC0I5XD4TG
sYlI3FjohwfTYtGRQWHn0RGL/8giMOr+7o4CFEz0tfKe56/ctx47s/EdNgUY1pAEIMB8Zml9RVSN
hR975IsaVe6278UlIct7Ft/AG+4jxGsZnqhTVBu4jVcme1zpZpTe7X+FmHrxvjbLzpOq6VyCt3h2
8V2CrArcm/uMYm0puBoHLYxKqy0PQ6s91cU0nSU4bWZg6wE7nLewD1jNJvRmhLb8EeAJpKDnv66D
1CKUTVvqdXyskm62aF/I8KqB7EhqQ9VSlYKVHe6/r0sfHaPPlh5vCcviu2W7YPwVSwkbTpl2gixr
cE77k/uVH+R0Ye0DBKhF9q1anRu0CLfBeDJX9InyJgWchK8tOFpS/tRz5Y9cSrxLEzNOwx23Oc/d
PKfDfkMx0rHIuBwYXmxAAj1QW7zPug6Dhm5BGeQoFIbGnntJPU5Vgogn4AgE7/J4cJLXIyUogsi/
Wq/AZcIc/S7DTf5CRH85Ajj7BDPqgVY5jZb3GqbQ0ySMG3/wNi1EDMOJlxqPDkfZVtoULDrl96Vj
n7vtZQno5/p/sq2R8unFlWkboN/HFuakK2NRhDYm4oIVLJhULjjTfjk4/69/XmHzi8rfoKzol3rb
DOh+ziMOpTXvIPk7GFRuSt7XlH0QZG16NxUpWNjYu6nlaeA3h74qbVJAoDOysp9NM1yP142FQjJw
uFUoaavHjnCpWcXy1rX51qqVtHATwO28h7pBKwC0VWyQofybJo7WAUKDD/PCigkikl/YFDdk3xdp
KARIPEhiPEqCWSrNzCGy7kvO6e6K/HNL7Bud/LpQw76kljMTVGtebbvcrCMDIdzeKwRZPY9CFCzq
a0zEqH2VpnFDIkBgAy2Pjm9hgTNqZ8odM49CA2xMKNB1cEfmSMELjd5u/KgLZIzeGcYQwiqj/A3E
y+VAxb6bpf+2h8sSS/QtCCyY7iX768jTM7N40T5HE/HJt1pO5RQrifnThFCrJmD/AUqvZyooqktd
gUXpO10hjVtOcPu4LdN2yVAJQxJsKHBWN6Kp9Ns1/aAToNPylaXhA0ND7UTrHYB7oEngiqFgl/Ir
/xITb2tFbZp+mFWMdQu/9BxO4HuVEazs1pn8cXUrFKhYf6SkSIYA/N41RRpux3kkaWPY9MLcnD1O
WehX96RuNla/c1HHFk0gycqAx4t5H4V8z7/KcXexET6BmC7EuGUXLS/Kjz8njX05Nh+GXm4nGyoU
rrGaRT/+72RnoG1T8imXciHtHrvaUndRi5PfWKuPI6owsnfNrM8hh+RzisJWvv8lzKR5J5xbZ8ob
jDy2BOLVon7h+XTMYQBsPArkafB7HFDCoyqxRIs7E09kGOCSYzXM29uIqWXZvpSfEWTdwx8JKl5Z
nXR+RqaQlcuAVFStH1ZJjBJRNGvch4fWldVjznVA+UCDWO5CTzYgrn1zoSPrSJo/97oSH0symtRk
aB45ol/C0+JjnoZPX4EbdYFZ1l8ddFsMnHAaTDACmtBk6mjf9iZq0s/HYjPDAKvnC/rRHwj8wyYV
zvH8qwiP94/P6VzbN/r1WTWxXsJABbLsRhOaSWXfatoZavSAkKZM2yIG/cDGyJFyfwtj3zbKJsZt
ZZtSd7WfgvjCCPdAJ2UQKh8iNQcQH1O8GXS4IcrnlcrFHDENpMGwso9XYfe6kJU+2zUYAj5qmd4X
QyPDOpl8GxLiWx3OzF+GBFxJ6g6q4HbDrDD22xlcGVeH9Gn1uj7WbOKhuG22CKWnRfZfewbd7YGc
PNSTEbf77vbc+imZZSiP8AG6at2Zz3ug3YOxrFNEGrsRTCbnrIFXvePrNfGAKEu4yqmyWbsINvmS
vwHp3AgB7poOBLJY7sV9Sxxq35W4aVLqOZwAOGbc7G5UaMfTOeYkMxM0qFVQX/bOzFTtlJXwMFvq
MdqhCAqmf2/eIjLZBDD1K0O/YMgnsGB5/fPHHK9fApFFB/k/RUOxR1BpyuoG/ikgydPRvC11ylmL
lTnIy+eoqab8kW/saJHun8RFjse13izG536a9hIQEtjtxRe/YPvoNc60VWykMBTX0WIw6HKLm5jq
1hxifJRbZSNDkiJqZMMiRNQniRF0Y/YUu+mhqyXnexAzCmgi55FYp8Y06VtVdQQAitk43PH3ATdZ
pK60gN5hUrvmhwbLdRiRnGE/KfBFdPF5xBI7sFq5eU0tOvP+yaS7zqU7jUA56PbdlF3cEZqPndt5
uBGPwIBgLZAXfSrDOIIWnr8vFwZUoSjuIaSyXVjyOs3aTwHw8HzYDHDTSJmY2D7VveUkRUJFx3P5
bhShFkRW5Gx1Ib5yDcOGu44n/CCdoX1Lx32ZQCQwAtE2XwcunLWPyXx46/WDkkrYO04WznyeJIlf
CGdDU4vJv0fMe2cWLXNYwBjry6YCqKHOZQV9AxKLjCL2h9DdEINCViYLWElGogIu71vekyNTyZ6M
seE9H14azaDfDBLmQuInFgf+MfuIF1D+glfdEMzkV37nBXcD160OLMyBOh/zy1lmlxGViuwM5IJb
GYmKB+B0rGB1e7WQtJlA3qXNY9veD0pjdcScWACiop2RhbhjtbqlAex0R2tW65dmPw1B2dRF55r8
FQ4k4NJjr2ngblG4IdDdCg7gR0rWxCy7audZJql/bx8S2Rfe/s6ktt3+IGBiurueqYzxb3XwDPWh
V5ayG2Foo01+xymTebuuCMDhPgDupkKAP0PW76oI1S93h7xM8zFLmmI2QPO6Ix9kLgAcDe3xiB7U
yk+1TYNCN8iMTCrhzN/KXmFD/O1VoyM9dLT3XPZo6AAz+Nkg9vjGY2wF966fsdPOrc5c0E0zhKpK
ZtiBFSqxRqQOxlNzZdtUFNtkV24BmVPm0YCexabfb6AehwF1dGf127SzveqZA7Oy55TdpdzTDY1G
RVClrtzr/0cITVMAqKvntvUn8vJUopZL19qrPiHU/eSItlC8MzYgK5rvi1wGzWnjLzuW+auwzcN6
BRSzI1oLm2dnRNI7vcOpn++ZaKP4fpdMc99sTWQutzDB2ZL0uv5ExcSbkxsj8/mIzWCj2SPlXRqQ
KdOOO6o7PCSHq9ycauOcnNJ7S4f5WkP+tzAoWWLUd0xqHwLAHxbvmOzF89/2GaVnKbSFTV3YYcCD
pcSl64aKdwBIphGdduT0kyr+NR++5kYoyN3F3XutrQrUDyZN0O0wGra5QU7wp8XRPZnzztqCJE3i
MO2S94oS6TeDw7/X3N8BZLxd/UgcsdPLL2k8Nc3oMX0ZpJmEKP2u6cl4TYF7DKQeZAcuUa6cuab0
rqsrYRjwem+dEkaYwASR9zwsHeEbYtOWf7TL6oMq1Wkj5Prqm/ilWTwZvESodswNAoZ9IrSLuBJ/
rNajiz2m0ulL44s9Hl97VP3jixGIGLYebSOGvCHm1WPLt2CvRMm9NwLeO9xuGtLacP9DF0+Fq1GT
+HMHmP8I2jJSNILMEV+IishtR5pAFUpH36BF1/PdMjRvb6HuNZKM+1Vy4HAeLn0XMC7uUeKDfY8I
cYWP8NM5ydVkb0/Nu+ObCFlyl+pC04kSg6M7cgY5PeCkT4qsPLHp09nT/pdNAz6BSVlDtwJPYZHU
L8cga2FnBGkyek5P1Ty1rKMkkCS/81R3UsLPCgtlqVjk1G3mRZWlrCHYCXcDnti5RgDL/Q87Me/r
WS9GMkA8Nq6zBpjdCn4EcGYOh/pk4KU3X11mYKDaxk+9xcgFsVH/umYXbSVOFN/3M57QZ/xuF2bB
2n4ohObE6tl7/yrgjHP0pl9stt3/WzhPVXicZhw01uDb/N5U9J9k+oX8YyoGDhWUHsvFSv6opjL4
JOFvkiFO08BF2LmcFPAfGjYUMGi+EMf2EUNV9i8gRVYtGSh697XP3s9K1mVsoeYD2Z/wQUUtYqUe
Fbmr9ik2qQ7XIymlt0Z2vTJZsDSQv2LCvkcOLx2X98WjHquIZtuvBTzhEsoObyxD1Dc6Kw5uZ2xy
1aICy8LGh2ijsLwl8/UgT7NPxRUCI4HHPz/I9S06zxzwDx27T7bahlXPY0ThhLAB1NHIC7bKF7bi
WQHpkEkISdwwJzDt1tzRi4Gj9OvNetruyZ6P9oMPDvLKZ3/SeeWe1d/Z8zT31MDetgxuoL2kfCn+
3YEGfmsxPnrMihCNpopPHzJxawZ0Ydq6tJOTQeuAt8lzDjFS0eORQEeMw/Xyhdf/TB/dQffFFsZq
XPK7A+x4kem8G7GS56sRi2CgYfnYGXDF3es8Dlcnxf+VostlFAUSjFWgpvohikTTNV+mOlRdgzDz
PtcArDH4qrsryEVWhUb2CpqWq/n3En2rvKLlaDS1inRTaR5LtcNYMIOGAluXj60UfAmn2NEwqGzO
jfITCfj8pCslGHZVf1/U5QcZwX+xxJEW/GLM+18M+pYlGQHu34aHessTwg5tD5AjFZ1eVDhra0nU
gehssbt2Sdz6hxblVG1r0uw5fMDf/6R/qGUQWyxQK4jFNb2oCw+FNlpWV8p3rIbQB6ILwMcEUhaB
YomGPAh4jMha4K7mlWEAnITDDnAXy6px9bMIxzarGQlProx6GSutivXXZIxgdp1Z+77BqNSNgCkW
KF7ussJdO65QWJlIZJldva4T3VHkZdpHLTK7Dmtv9we1qTwEBqXz10q6c8CpwcRjLaDL7CAgkwGw
k3yPCwW38QtMafX8KnukNynX+E35DPtgJfA+mpNpbkirGz8Yes4Pgq53ESOZzBb71DtybG64n5cu
vhKqmusvTY1s4KVkmVyYf+8/qYGIDDV9sG72RianQ4SaPBKQQ/t8gHll+JWBbAnrM2g2NRN1Luqh
Juozu6srMNg76bbLbFyEwReAZyDQNXjfOp2Ac6juBAyVKhNdcJWXY/Ry7qSQ6mc7dlKEcQz6RyUt
mhvlNJ8yKZ8mvk5MZKPZ+ZaGjbqWmcTM2LI60whNKzoNY1EyZ9UcMHK4eEPvKTkzK01w2IzQvp6m
MBd6wyRi2J7x463LhZl7byO+gFOy+pJBwDdU1FuZETaBs8ZTDlQWEm6zmkZ/lva+bRw3NaIzB6K8
DuOXpKfNItU1KLoDhaYV29DQ8uNcEMSNU5RvVSzftSRorpB/fTAsMxc83glye5Yqy902IU0jDBnq
a4G1S8RHQg+Wmxq9HwbXt+N5xb1lm5ZY8FIQ2YIsHhQeqeMMiZEsikXcyzRL7zMD+Fuxd5CtzWOr
83L9cdSZByTBkOZmnDdEcQgoq1qa5AKw2LTXVwprWe4qf0BWeQRx43JyF0pewqOFGZo6yb/fA5tn
0SDc1F/6ILTu8ypCWTZVpxL2sKoZ5zl+gDcI0yyKiSzc1PDbcs20HvE86e9lIbw+KPPgxgkCjWrW
LfSz+bsZbpIbcVaRrMjxl8vLCtbrJJq1jIzw0Kb5xWR7GuMZpbzji4s8ZxZEXhvyVEn3VGNx2as5
SeKlTnb/6UapGMZiViZ9fCXPBYxi+K/OghqgDISw1X1DBxsOPth+4ikjnl21WQiSmSqXZjGleBjs
/WA+J5SAozW8blhv9UPlpMDoSN5N55IrcYgpELU3c5ul17o+sD81WsAyE8RcG7qLW4VqZq/uYydO
tx6vS65rqDtxJPposG0vyKF+CPS75NHJ1Q6YvslSq7qE5IXlsDW4q8J6ejWwwPoayHskJ7fEWweC
y4EQZ1sQjZT1L/XsGIVWvACNzR/z0+Y4qx1xWNH7Ub6hWhOWBxF5w//q2wrh/imNL6lCAKQQ1iny
SQ16USXZzF4bAMXRdD6/BNd+bGJnWtJKto63jEzIppM34gBFWk52fHGmJZoqmtTSMwnFSuP+78ay
WcahgOBQTjKE5ip/pAwecyZXoOHOQ3cbgz/dLwgafI3ulc+nweTJjnySHqU9Bp/ZBJSyG86y/vgr
yNQubd4APgAycT9OHsil1NqjGuKgJRRihfUKd5BshThm+E/xGeg6Olr1v/aMWb7z1esXFpu9Nuq+
84Ve3SzSNkpFRNWYjzhmcCmYH2LRGMoWNUGx/izxWpOVsWXGMpGxh2kmRvgAvzX2O7MmUagnHoen
S+cGI9FdRyP+/4AGt5cQ7v26Nk9pi8bTkMnpynQWv4yIoxlKiREPYOOyRFN+9F8GgJaYu8hahSxx
KWjIhkIJjIe8pK1ndhu0wrO/d9e2zlh4b2gOIuRTWszgNvwajxKu/hJ1vhiIwRmwn7YvB3ksXj02
Tfsg1yxmBKv47gjoIEKSTcxb6wb12Yv+1C4ExsUo9gTVzpEgUHznG/6H35J88z6qwBN40znKbPmJ
zw/KTamVLSNbXuwV3JSQbPAPIdMmrJrdBRX/KTqLUyN/hnAw+9szHMA9sLSC5PynkQ8FEMhs4OgP
A0h2mG0Lhr0XNXTVX0HJMI0QO0bQnjSaA34egzJtnEhM/Q8oVNb1y8bnW6goAuuJFHbfb80Fdjvl
v4QWXiFiBZWj27VQicYXNG6wplkpdd5RvrE2E9CcLkTTzNuuVJl1S1yFmDvkVSiEVG8E4/LclWKs
7rRSXTusa+XgLFasDs116eB43x1eWz3QVcwgRc7TLQBougOT4ht5Y1C+/uG2KDdWG+fTAsbeBVPe
M7aehFcbiv6PAK22QPJluwkrJbmFX4l9nfdWz12bt7nMm7gm1W9DYZUGAeoJZ58MhaPOPTa5IY1L
8QIwAOyGpO+vQhXHfzt+jx+JV3nZJJJJxPJJO/tHxI4Z7mTAtlSYnEvnj7WUa3kxFHJbZ1AP6phP
Y0jAoad5y2YpeImiROe6vGWonBSs8oqvJ6kA/cNP9c8IBf5Z58g0HEogkHUCVW+qoRvaDYBmOuEt
SZ8khc5+cQVwrlw8UzySJbyzHh+fno0thmrSJS/7Mt1ZNno+/OtyyBhAJhPwjXsKgGwI7dTfTc4h
ibTiveaD1A7kK7uT7OjBI4O/Y0C0iLG8x8bYLVx3XpoyB8hoH1N21dD0/vCt7y3DYaaybbj5M9DC
iItknnRaWnAlZJ8H9kzc+n0Rw2DuRH7SdFhwblD3M7OZJYPcXfNn2uljSgYyozgrF/UhfDd9X00l
LKGqQWcsAZj+pv2iJTAFLePGRzjpTszhKfTQ/t6L9H+gilAPrcRxx7v/fs1ZzrDrK92L1X9BYD4r
5vxG67vHAOMWlPKwZA6TURUVcV4BpVxDqBbIqQ5vRV+NNFyZu+IOJq2LFG0pcRYQXUNrtBYwOjCw
0prJQN5H79IuAvFO/dJkSFOxaARmGOojy5NZb97/SoLU05FYb+pqZiUgXE+G/r+pX3Pp8rEDHlV2
PAuG54Xhz6JFFrjE1mzREK9nzYNqn+UJlcGYerHBDsw6BkpMkTDQva8tck1mE4yHwJq1Gc7gwr1X
FssvBsqFpWu/2hmzwIe7yC+GcZ3lFm2DsjOmdPNt1i7pfww3PHfLkD1yVyeS9P8Q9xi6BegSlO4B
07tQOnMlAfjthO4dPzZlrJsd5lYqKJsOMZGrLp3hvMlu5rwYAZdBQZvh1M90sBcw+As4ZCUSs9Nf
aPtakfjaSkoWDULWWqFi6jO9WwlypCXiB6ZRndKkGbdXPjKDCKstwInTu0QJI9ut69jQzm4E8KC2
SyDWfsqATIP3Jt9TcpTCB9hAJSF6qRwedIjK070ROr6aD7QJfa2YRInvCGnGZe7iPLi8A+hM6wtb
SVomeSgIY6F1DEAHqATyedx9BCIGRLZTTBJZfgD3bJ+368Rr0XsQXDoo3aA5ayOX/UDfModYLl1D
pzq3b8kb98MaG9YbJwEj8zxYdu93rdh0dbhweDK7Oz4YcR1K00vQx4ZV66oHwovdPBozP/NyI7yd
gsyb0EJd1c718s8Lwl2ZXrI0wjdTpZ1dlAb6BDAI4F/IK0KZ8lYgq6XYpQp8CfI0NquuA3aRPmjC
vU2y6g2PSmgUWkiJ/3H0tJiTeLsXi5dJqe4mkdK1l7Bit7om3awAssoLgmoRfx6IF1Fgt9bGSdGc
6iDuG7KbqJbu4kF/Uxzm/GPiRP/iQyrONaXFQryOuc8ITZepGuEc3LiG5RWnB6BIBEH7SjvXbgQi
q9xSny8yZDfM4Ki57+2S9gnAFtXMj2BXBNFXjJiY822LQ4eaqaycKf38DMlgpFBtSU3NQlcwVOng
mfr9rcNIbFOgxaY8ANRZWskw1lrkWnm/KUq7ezAHVpS5LdMLpTN3c0SvYfYozqPh+SRtt9/oeXSe
a0hl+9Hq0RKyXHKj0krmYDCAPG0vVj1P0euCxPSK9rGX20mrN0/chPLE0IMo5XBLV29jBrXhAD9l
yw9JQpsIb+S1wa5mqxBqe2jHdlwV1I/NQiXrOxQoOV02IVdaYlyZ1Q3QaSGHfiNbV/Gfr81wL/C+
SXT8kyoK93Dq5fkwKdsKcZxSEB8pBwvdTaie1jgRP2qL+Cr7jzjBOytR/BIlyJp9DBBgLM0ZuWen
egQLj/7Cd180iEtmdo7Y720AIkweCOIiF37On313857FIddO4ENtd+VWSY5muBzC0qeP1xXH+1ey
JnqZNlPYd68SAkA2PdXFwn5xiFXejag3oXtKAZDwd0rgFWxfsqBMU+BgbPstpaGn1vNf33njiZBF
ZgY1OTwYKOmofntVCLzqKQLpXmBrMsccxa/nUvTHOHECtNqFJNqXUW16lLo5LZMYQqEea0Z+lFEf
HOtcqKgDfxOI+T/WeHgU2VCbRikNF9cFpHcUOLdc9rMekxxTBuuljHGtWRT3pjBsdcn1LRSHBI6H
v89DOND29edW0fJ7Zvv9m73poU7Yxj+eC0eFdkkybd2TOe5CLdhG+mXkpD4KoySBEWKibRyj3JMF
3gVq/FW4NKF7OgEFBXzOdI0lGK+EVtMsaw3W2FCursHQHfGDa4Lq3eMZMriD4S4EVO3LQ566wQPp
cTbu8LaCS1jDYSv5LayaoFNmqK9rrLIfTzWWjUXVBa6H900g/HXb7T8XoVcDT3CvRBer1AZGdpa9
AKqqlCEq6da/9+1ZrpDpNkY2sOmAWqAhlNEhTMOmJM1e1vzZOfGM/vmalc2/OHpKPWBuXMIEXqXt
v3ePKDYt1Msrtlkrni14fZjQ9nhZhTsjAWmKLC8STSrIweZmdtSFx9P21AdTk1I0uDqdyh53dspL
iwi8uTJZ4OE3qZkyLny0CUZLulFt1+RDl+vNVBxMV3oeZiblybC9rkKs5B/oemdcGl7pt4VpNGov
NCwZvMpWV+BtnE3eMfdjSh9lSuQXyHFxvjF69Da/qny2WzMQOT68xmDjJwqNyS+5SHNADs+/SEh0
2GgfLWWIa3aOovf/hqx8zXw0fjpCmVBSXp59WPc3fDXi0MzJL/cOKKpRIOBdvZzTuv+SSxCcyWAC
L2COy+HgXfE38hRqv2cc8QD6/ENIme6eQS44xUeZpRX8xZutOdv6IMuQtBcJWhT4PqyAdGaZzBD5
uUmd8S0cG8gfb405+BW29YXZC7KPlsMCXa91m2SokO6fjHAoHMFqCbEA6ysL4Mxqk3YPW4JAOqnb
1XCQorA5RAtcO8M9U97yuEdHIYESAUvFzY/kRXiGqo5oZMT2XKUl+FjNGQKH4cpnRBR++nsQKJuT
CQHKtX11BBMB1t1uEDVIK8g13N+181ZXfIgxKy1p8FOrV+zDVfkpM7ozDXox/FXZa45ObEattsRy
kuou0ialLWC3i+Y/dGAmDXcW/QFecwIWX6O9hgXsTzttnLiiUEIhdrzUYyIjcDhB1q0DrdhuxSwA
0LLr4MnhFP3h8WGSteSOzixvNWUcXd/k2pW4h4oLMGqLtg7jKM+ZQOoaeBeu1+GIu9nYjHOrdCli
nP9CkWJGQHscHWWa/J5+0oyPADfxHevCfhxbczE4sQi1Du6PJOdRfW3C2m7QIaNAT1ZApXwWBioi
UdZQLAaiWl5eLyglu0VfasDW6inT6VB5fOIRFwFGa8ayOzjYsX7/0ksLk3Dx9qJ4mMF7WnXgObMk
UXsVUSxetjgQR1fKlITV2VgAOPm6elMO3606ldVk6c4vqgVaVVVzcUzs4oRTzWiOS3EIq5ugdVnz
PU8kClco6GX5VLtvQnWdh7OzTgI5cwnWJxtzVInaIv3QIyU5QgnYC0u2aouDbH5/aM+R/GDEKA9h
tzizGJ1YleDdghc3tJ4cxvWAlnYOtzyb8BgoJNiz1+/MAHhTymCE/bJAUC27CIdfQJADs8BwKxPk
fsWVeX6qZXzmznKKbiJbag7Y5hD6X6YxnRha55R0cYGLsdYZsmijyC6B25HJwKaSqwQUWYMdi78J
aiBwhZAbkbeTeE2WmX+W662xm5cVP5AsB9+uTf4rfk98uuFVgdCuqTLa//mIBf6HWfyplcgdf8rb
Nxxc6bJZGKA3eEHaMKVnMLnXPTWc/c4B7yDWykzVFW7gp2IKofs8groGiKBtNtNtosxY5jWkqsqd
gfchpeQcgIJTgwcmfi0wl3x72Vf43gI/VkzfnIsC/anzcwqo1YPcf0rWR/t7Yql1dRhHafK5Yy8R
11cFtkTm7Azx4HZXjfMoHFChiS36OsRlg/PvxPOXNzRyIizG4js3r9Z7P0d1YR3d2Vw13Sz7v7TL
CGyw4qePWmX9xGIVOlpdvDYxc/yvRQQSptrluyC9QxilAOij0vNXgDaf9ZunWgzY5jabkFrTTptA
6klcYcRyOzFS/vawJUPHUfha0G3jjsLtnYXufSgWZ/2WGPODZAkxL7QSqHgna8PK/B4Ak1kDnl24
qmiS9xjludcvsMSzzn//pM+eG/EPbL7HBpfByk0NRcR+HKHgaHB2+/Ab1N02aJho7WVDoABJuwPN
nHUNwkx+kitHMVBneIkI/OihJzZwhSnnWANBOH8a84cVchDcliaLMp56TGPOmpw8lOBGtl1E8rqo
oS4HN2xtUSCQsJw15jQn7g7n21im31ZyhN/DjN+CmKuLz4iV8QbxlG5q2CsovXSuz0UiG7Y5wb5k
1yf4DT9mBs0c34s5icr7IGt0Zkbs/cxIgXN9aknhYWbkhjLzD280CkXUgSaVz9Gned2idt7Tw4J4
zUcNIx69O9Dw1VEQwOmwwqcuN9pHGK63GFMloB+IR8TBXIivIRxajomJBuuGef702QtaZdHXu/Aw
+jZg+vc8q5w/qtQnc+yyE3Sk9sXIc6caewtunHZ01Hoykgx1WHJPh5eFbw8vIITKw4STsFUGSGL0
7odoWrpXRNjuwfQI4eeXYtn1cGZ7bV8lgXL0icgD8iTqQzS3xnC7qXyrsH+Egkyzhbu0QBJ3hWKW
W6ocODhJpy/Hujo7KaRAjpKHCqpWb6ZjfwdQasmJL1Dq84h9i5y9ZQeS/KEE+RfA6m2moBjlWAu4
TLIRsua7Rwl528fYts93yqokq3YELfm0qLa14IAN/OrElnlGgS3uXZC438ce/DGElPQcSvKNJHjK
o4Fp0K57Rf2SS9OaU0+uiW/h1CGo4iJDfWPO9pVeY3Xtti2hR82UmE0cn6t6eOdCMCbHjCzMRQOR
zioX2XM7NOz0Bh3YWzHYqk+3L8v15S1iZMcXZe9sLzfNqvb3FVq6n+UFBNzOc1ODWMZQGnMRaEC5
wlXLNSrGNnzfyLehNog41sOX2OSimD65b46NdPaIWRJIrfCi+3W/doS7JCeP45pv23jLtDhVqC5d
vc0KSHdfrZCPAlesqp5alaXFXrku3Sh4CW0h92Clda/nFCgS1WDUu8m8y6BQ186VBM0q72yRDsoB
dmud6NUl9Dugb2Q2qsxWyOm1omWk1ZtRLQuU7NL4TtWA8zz4mTiN+5wQDh2hVu36LroShxk9EALo
mvL1LZbJGQBE/+KAkmaDCpoldZkJ8K6BOQVJxcsZTBifSwUbiQi19Kif9b5eKNDsXqKt/ZufviqE
TNOnZBeevom/1k4pwSu8RYl7T60JQBkCyu3RV30LLalijV6z/ejX/B7yjtXFIBwe/7rjRk4nell8
tI6MvuVRYWuQWtue31JAJb35qG5LqAJdGhBsMWRorHyKlAAU97+PM+EMkZHDHho7w5f/+dDtBVvd
iYs1qcDGSIa1di5GevPWHAu0mS7Dp8T/t8w34d7Q7NYrpKO4jJF1vLl+qXvzQG+l24Rcwy/xr3+s
lUVZsmbRznhJE+lMTyXeyPMNMOZ56r8BnkiB1tYc8z5g7l8pk61nYJs8ctVIBr2PPwlJNMst5JWL
wtr2KpWIYpa/DpX8D8pA6jO35IUPD30Sfwyn2Lj0I7R4W9oHHPHMxFQuz4lAc5rJThFiZkwMUlQb
KDIkG09me867F8pgL9XNtVJtTm9nMILsEBYUUp1w7r0mIxqXZKQynk/5DrJC/erko8qtp14WLh88
AwRwv6jNNvtnlHbYAN3al+erB3nAgFsJVnMKxQ5+oVefR5OM+frm17TjS/cuBlXznvmcgU7ZLx97
TpYKz0/k95E79AtfxH9m33CWUM/jAztAhV7tbN/l/jlKd8dxsBWIAxQRUDNgdnTKb5Xt0eU5No1i
lMWO34GAXB2zJJlmZarlTPVd4db4Da7y4Zq9Wtj4sK+nM6zQr0K8X/ftQWn9u4qFnbHnw3fNDYSQ
v9QK3w+evaJjvq31mI9Dcx0sR57dvw4QpeEXFfQN30I5GNXO/Qf9fvUhEY7JX4lnkxAFQEIqA5N6
0esBD3M5BzG5qnETz1lPpBNuAiPZ2KQu+1mxcNKT6H/H+SdjXDfn8qrj5dO5WgYAng6+fK/jErGy
4TM0BFzOXhi5vaZzehrooenvrk7GkXAP3grNLr8UzYVe4taQuhVz/eprbeZ5vzyJVNok1Wl/GPys
GIe6Ygkgp22XypLEaOfWV87FxXPHL/5dcewgFIVo8YKFhOGV6++Armsen/qh7exCm2gl8olVZR3B
P68XOdmV6uueJVyFDo8sm7adIC18IV6rckg1LSNBwbLqJCeDOUm2EJBsWWCPoMKkr6lgdZbj6L5D
Upb8fEJaVqZzcAyKXUUu9CFcLieX0hYewpaRbs1IrD/TeDjz3olN23sQLUYAp5fCzKv8vwdaV3fU
0dr6v4AgYtymp/Jw4q1qcBRCAFJvUaM4LBFgukqo8srK0WAuUWMB6l9UaZgC8pXDwqdgtZhZl4ub
ObxAQkwr7MlpJ1ustb826mSpcSYTtkWPgcS9ctg70KvWOsph+U/NocY+U9FuhP4uiUMHB6Y0BjGk
p2A47MlX2MZrJUCA1aPGx1JFvK9KFXJSOn3aIp27gOH32HCPnWzIDlP3v+Q0xRt2eYXIbo5GAlpT
QHzNOtgc+UkW0zlFoDM/1OjvRkR8kgDLkg/PK7Wvelt6BjP4X/J/K0EmoWTM0rChq6s2fgb9opuQ
+Ay7yeDk+KWCoQ6TIfQWgRrgXd4E5wtNqobPLcTiiUiiaXF4sYcICgEt2TShgC3m4VVPGeRt88zO
rVp1+v4j9tqg+h0OuJ3Ncaw2FFUpySAa7BN0L2cCzt4zSh2Avl/3aXa9bqaxuRJzLAu/q7YNrmuM
YMyBfalwRuDhiLF4D3qMBPOn/NYB6op6E/TE8pTM4oyfGbjmDAHjvsqteLpBLZ8JD53lPzjiEmTW
4ND0JopIhPkgI5mpRCYTrhzGjV3Db/6I+3r+s22QH+7h8ylz13h9zfWAfSNuw8GGnlMzQUHHaRlr
m+BlVk1/1wWWRLvFDUBsR0arZY9fMEPDhvA7QFjiXxBGuuBqeU43azokXwwEPDJjhOWt5kuH1IC1
L1l3LtYDXwzZtLWzB4uO5jPZx3PROVSXbPBCyIbTLWkUsiwcjkrIAI7/0/Elv6WVjLn1vy9URuXX
KZHyFsUFh217w7T1lGmjHuK0N1Iv9i17vl8PdDeK8DHwFRK4KQzEZS7Op6AQQemrfejb3yip2Q3N
WCOMuH1Xa8oUJ7xi/89fluWKRt+7RtacNUNO2Mz4xG94Q9/wlC0b4PTElSAuxjN3+e4jo4A+J6QP
5LK5leR3HLxEut5ANrGNVeHb9/AKbzkdkMBNHTGKHHjsqib9nOQXOaEAeDU2lJNMa/+vc4Vi8wWr
B1ag5oefu1+F8ZH3mw+ZAM0FHXnTDCLfGTbU2cQKjIJnM27etWhZ/8Iycr8gqKEx+Atl3E2GDrpi
b3flVw+g6Li5utpTJpQ+RDhVmrqp2tWshjs+6IDdSMIGyC94FUsl1vJac8ErcJEtszqdlWnSeMYO
shuHnhXh/ePwmSSYxJuAzJQ4VRSl9VYj+F+tXVOyK+eZbquoqiRh936/Nf6WvpUf3kvo/DUSKDw4
SZ6yheaY73sRLmXDj6u3u1ZM0gsinHkztdXdcvCpAmr44txCwsNSMhTuP7Fr57+ljGiO2+g5qPch
RxDBHWpnQ2lKvUgIQ02ur2RAgsz7Q+xpylPkD7BW15GH2tTEjJ05c6pjisFfMhaLhCuh1J6+KyHR
hp/luYn+U+x94C1b6y/PiDjvHbnt11VXMbSPx1O5czQZhz0JEeoyN9Onhk6k4KcJA63Hu4HoriIp
iB7fuGY7SPRdxUulqqg6IqNdq0ABwItbBpkCITvD51RfMwyXLmLHbV6YTmE2IBAW33cR/VGOzFJf
TGWMc7w0fEyR9BfJIblAZlRft81by/4HgC2U3fV8+r4l3p/loIyJSXEw1bFkFPSwJNWdzqI/gNqG
igs8LSM49eKlWwcVN5ysKVcikOwoag7LwLQDlzjFjnZEFqh3hf/8TEjmp3xjEgBwbx1eJXfmZbhN
atcvlGa4n+DyShNiG3ls+jXOZZDdfdPbwn4YLvWayAWwLZAx44KkbJdXzTTx+oQdyuQ70/O8XFgR
BstBhwT9RShAYtaKCiqiRGenPhTP+T601evWklzF7IzGswd1+sq2M5ULhb5glN3xCGveJlZ97vrQ
U2UGlBf3/hyr3wTc2yHUYAC1ZmxS2UhtyIOTtRfLAVD0CFzYSx5WgXBoiyFZG9hMUDcHgAMliMyt
vi0ycL7iPONVcOGb2/nz44LFf96LwE4wSqfzTAUVU927MRqappk6f9Xuxeh1Xkh01wlAQLUI6a2s
MI0DrQxYAHK9oGgTI8MFdHqXkeuszRs1fFetfWmVnrUwes3Qvd7XC4lEjdHqCuQEm1fuskr2rLmv
EegwbeqthPHs94Cemv+8go/d1ulUXfYbMG6n40KA4W4itDOHjyb3Q3njwgQZpTtqGmKcTmJg7WQb
wB98P2qJ4CGhsOb8VOZstDh5Qk41hB18XU7y9KH6tDRvhQT1wDwSrvdLylYpi6J0C3ltxbG91QTT
YrG8NxBAKAtJcZI52wV+XlrC+ENxngVioqLFVgrJxdvgSCCjpJJ88MP8nXkzQNgT6XmFYgONdxyS
pa2CrdRugKLKAyGls5fpvwSGGw9CGQXGtUcsw9H3DHdIzqbYiYZSS62U6eQNt8XQgX6EARyJ073A
WBvX3lI2hYSNptY8nMU5z6KR8yJdLTcrghn7n0JMQTZwL0QDoVKIJaA2bBq/IF+bw6ZP6MflOfF7
6zQ6mqpZxguFJsDyeLZ+puNiENiKDWEN7xoHfH3zcFpAedDZ22/+n+rFajAceUz7vY0aYCeih2mO
sBSo65akh5Q1n9URp+yyNATWT8vf+2r3A7XenBhVco6BasOWGwbWBPwJTQRHL7MSVBq4U+38rk0g
pTmHTDGDjUmaXtjmO1WH3FjtzVsZC1ZkyWNNplGeIV4IA1S/awLdQhlzOGq6EBMV85V+ZdddBtd5
5/XbrvSCrs5Yuhnoz62a/jzFDn7R2A16dLwj4N/ALngeI2xMLYuaAEDqo5kPuDoVtJkiECINPhLm
FhOxTPqGcQOX02BHzByXfW8BATOT0N47NZ2goOQwG5nhisUBdGbyCwH0F/ut5UTEJpcMiEw2EIbz
q3TQTm/3aBRX8b+hJvUlA9h94qR9/JgNY0EX0UriaX31W7+OAe21MPlsEwUJZDi48G2Z2xiK0BVI
Q4adIddE5yAqVVHYvCAIIJEqTbXyXcdK7YNt681DxZKYZ1xZNVHkbaevhEFXu6A4ZXHaIZQJZAoy
8cGj/RROWM3TnaLu0fjaLC3ZtsPHhkZQbFjAFrRuNun9ogSVbwwI88UL1B7ROFqUWWCPcfIQcu32
FigsXdXWMvs87pd3MHWI+/JrUVHn+iLh/4LhDfVEfsplVEOlU/1vCZSP+fk6w5QjSYV2sAhlfV+y
fIbnsmzHAzKS9PCCUpK3i8mc5tHGoEEctKAI4TaM41PHh9kxiPBnCoQDZSD37wMNWHDRJk2CraDD
VKOa/OV6clVYAnyE9yUHnwivNsZG+VsZVkGPDAC1iiit68K5zXo1E48r4FEw3aaNTm1myQFs1WwN
yOF3XgqNDWU1xwqQt/iWDpl4UDwsIMvbLxV0IzpEFJJlDNG7IRJ8haCPrdu7BXeEXRC5o+zKhW5t
qStAAPcfy7tdm+AXO9y+ZgtxTbVJQ1lgao2TKmcnUe5YQXQYsFTNrtobpmT+kj7QPAIJu8ss5l/c
GTXcJW1MvLJW8LMXpirL+16iLb5uSnx1SpXWmRRJxG85rtL1UHuyddjxrNwmhjklKrAA5P5Obcdi
QprStlDL3lz/z4NQT+gQSUKTy5/1sktwr4GZDesZx2FB4Tckt+1sqLDrzPjxa0O95LcvClGl8Mfp
QCrnqLjuHgU0sGIgifyTuX5BjFnuirsUWJ79EmKMteydw4t5+OaeweNW5q7GdCcwGu/YMsHIFysB
vEz434jvRTXZHfVP9pyjOAmz1+dcaILcAgLce0gFrFtjeOl88Go/EFrmbeJMqDPU/U3335WTApDs
IbInEP+8TDHfSTmJCKYAcbPc+bQdo9kcZaAmr893CdwO5ugUje+QqGEF2IUYcfEQV7B9oApOH1dt
jq6fI7jHMpgpF+GmZF1mj/iiSMOkfBMz5qi0yQMpUYlLteULK5lUJh0RC1UVoAuAwt1b+9OCD7G/
H6W1g7Jvji2Zcl/3HwPqGbAbFCqPTIQQ1Dkf16OZeIuthrBSaudQcuiWXNz5qCPCElLWjTO4t9I5
/5/wwMWUC+LEQRw0gOj5DE5/JGXE99qcx1erLuSa9T3g7WNcz5zV1AxF71Ig8+PydZrNfVE6GMOd
CqMoUCYsBTKY261onkbEzjGv0yM1njLyWTzPflgQlp+hV2vz1sICHNDNH2l1xTjNMHhOcwh29f8S
7FtIauNMqmQY4swbcNykhrC4+ZfqjqNgj3zY68jpMP613Sli8f1YEbYT1PsBe7uU7s1XSVw3EPw0
nVdVMRgn/xoHCVCou07uUR35OkvfKGWqV8+BfsxeFbzwJ0kKQaXeoQPODmtXvStsr8Lsw03ry5YM
yV7rEUPkah3zBpmIQ60DO1YoTBcZKthRpUKeeW2xqT+EqMJwbKgDU4nQy4N/3odE9VAFvN2631ta
kOJaeLmV+OufnAA8jBSdzRDfmKHhawhZe6TK8tbyRXe1fRrf653wBwns5/6sq1uQdouecF68/n15
aJDgdz/KsywLudLvlM6UWbw4FqfT3VASPvMAHTlDcr1MV1eEGrvZDg38NJDwYpPK3hAykSAtCpg7
USCVHlpotYW26LqozSiwpbfTlDsVBHcqTRhMnRKQ0mS7pV1mmOoS7GcO33H2SRs0tSAcowzU1OEs
+BtregDFyhVmdfimu8ltsywDOgvvB873PxMn0S4TxMZPSd3BvdK6xr74ODRTpGCe1bl3OgOMjNGi
RkKhS880u0BN8Q73Ge7Nl5RwEPAi9h1vO4ryFV55GYnaoOk4yF/kz8J8v3WFGIESgigy6snQ9LN6
m3nrpZEqkqUoLXPfRK5u9vtSlrtcsPCWjJLQlbCk3xMmJJxuQdbQT8o3vIWNULBCxNrqKq6mOVoD
cZJTEt5ed3MBdT0WGkSV6e0yXisaMxBdINSY/OkE2YqCt3eizOKlccZGOLBFYCUbRgG6N65U/GGw
RLFB4rOCcrY5IIK3+K00O+qCYk6wDa4InnLxoJ10EZvEIX4vdh3wu4nfxQ/CB3eLYWtGkRTdR0JY
XPR3hP/vVAU/XixBnhrsVeSfXSU4D5Yh62LXR7uPCgROcHz7cj4CQN+Fs44qePY95zfFpbsD0+TX
xwO2iTXDMoBlYJodhfSlORPZteHRr7XSAAZ9RH5aTE9F/ehmK69wtoGNFrijN+bBmrMrVyHmnZnN
0Iu2ZcoPnqhT/VDcTeoNKVy+MPCDEqGn8fRIskTuZ1z+4tbUfmjPNm254HDYZHWWx4iXQd8l4mXi
YZEpR6xfMpdrKEFIxhlBm9rk82qF5kXpMfwPmXhir5t3uaabqDYG598tcMWxu6y2ubPQMP+B7cvI
lVtChuWf1NlGmmEKv2xZlZafhV4Luw5tjqIRUfo4mduB+p+EoQu3XDl0B1TRbPBlrd7AypqKd08M
wQ8idU4o1tmDtTnVu922OjbJhgAEgOjqrkncmK80/GcnssLUwel02yT/UBPha4uNNLHN81L2UlIn
5GsAAAo6zunWQ3vk0pgTzm20MiLAvRQwMu19x7g5XcP2qi3f5e1ReKSizQLLST7yAijM9uBJqzy6
7n77dKzlQIuLTZ4q7jSRcIxfSH0TojddJ4jHp3UMbrPY/O8qYZjkctzAuYkaLMwRpeVNSpZR49ww
za+tpjkSoDC+Q7JCB5D5I5EqCDxAqduatGomNahJs7e2zQCp6QIyZG0YzKIdIrqOHXlG+4KHUWGl
YeASpunL7GOIdfHiC0CHY7/fk3TdKowW/Y0WMrsIenwGynv/8UONEm1kWtLqefn0TVPXW2r92BSj
1IMd8uxf3EpsIFa4AhGSnuFFUQzWRp2WuKQFVlPPg4miB1zqA4gT2MJg3NOEbu60E50VpcqI1ngw
1eHOizfeRqj3G5XHKN8zpmCfUK3kbAjvzBWcnfbI49iMSFGxtEOP/uagQGQq2Iek/CdIhGnJtJPE
gHxY5cnUAFmjxPIZXF7j/Hc+wDL7FT/0enOWnkgrMLFDEN+8LfHt8PbA5BNiwUBcOeNGmmOpRF4b
/Ho4NmPI0KW88yAzbQTKx3CmD8l5gPax9+1LuCSPVONlyLEKIojkrQtsjCbSTr33gbv74ZikleGf
SW2c73rzEwzIaNqU4VmBSlyYWcKVlJdhAMpDEZK2MqtEeOU5MipG79fzzXFddn7ZSZTIPUNcDlNS
jBYnm+iqGZAPo1z/1x0yrbDZHMTkJWjr0YGyEpXKMj01AJKaRX0ksvDaGz7NmevkgotNCI/qyHh+
Fr7LzkPEzEMM0p4+tLpd3XTLjfLi4VCml62yPeIHbZ6BGaCQnkW0bQ8FGYCZzSOEuSjOsfbrW95/
LOO6nW/9wUwWyrK3LWjzo58SkNnqdHD0JM8elA53OagK9xlf6PR5Y32LrZrQ6a1gwn/AjjrST3xZ
4V/4taqWfI5bwOr05o8VqupY2ntVVrWEl1HlOb9tn8d9KDFRjXbRSx/QCYB7OASHtbu5ZLU93ZOa
1F2+ICAHJCUxYcEO7WqDZQ47RipYSAX+yigW53QvNWFoKUX9r64wyKMfyJ1aOdwjsD0QppF79eJY
k+AGLrZdqQASU8H57BVhKV3/1DSoaJAY/tKROznDHMUz8eBCtbUWL+P3M3tRfj/Xj+LiRPfMOusK
3/FvEXrMzvD61jd6VXQUskV4CeSlmXU24S3+ETyq7I4N0nhmFiVphxvhhsH8PPWxOdAS2FCedydg
XO/dJ6EN6Qz5FGbElQ63zpdxbgkDESczGF5gYOC9Q2a2pRweP7xD1sv5zfgsnI3hFaGvJ6W4rgE5
unUJrcRGUSztSqd9/LzTYgt9+NDX///qXVwjFGWaXaVVfrDiTmGEdwZMnoGBVc6/46wCfDnb+TwL
7HlEWi66PL4Bx3PNJUDdchn1X3y0lwWtfBBkS7s1EHHhgrBaLcJ732p//NLVGfrQxSNM/uXHK3qw
ISaBGla7/EeYX5Gxmx2epdhGGRugsCwegTKML86Ez9NZva3xBu5swgA3uf8NReYGRgkhQ2WaJo+o
RoKqaIcJCs4xkZD/gF5rfY5n3m6FjMj9qNWJIK/wtOcJ/kePq0r5Jsn9nuauls03l4l8x1jgIjVn
J+9S3qm8TZw4LsUPhmi1g/tb37QO6Tz08VvZZsj0jp2gDvdFLrRbPgOyM9My0DEaSYAMikskcqW9
2lExFy7LQO4iitmyjcN3CqAQQv0k468UtPE2fnxqnLrgitPUZ1uWm1tiymd5uZJbLk0O1855nlnX
iqPE6SlNw3Ri6YusSakZGYc6Jl7RMAvHIMSP/jiJNyX+O6KFq6Z7xku1RIqemLB5DPLTkr6p51Yg
Be9whYJekcbTSCie133vguD5rnJ0z3bnxw5VqkwAImbtXF0pMX9x36pHWBT2kN7dUfXXdgACzxpL
qegh6A+vVrzp/XJlAXPbrF0XL1TF+G/ybAsRD7tfTlDa7cxsgkCVKGkH2ol8usoywXZ3LNTs5ULf
OVdV3VGvMdDk9OR/oCDQxkHiYmFqXSM94IfC3+kUvXcf9PulfbaYqyoJ4sz7Kt2JbUpnOf/bi07s
LFChOVqOYuok9dxtuLfsIMWFJ42ZX8Ets0QNBujVdVbMZTRuurto7XFVt8ouje3RGKQWlJT7pyT8
sFUOoaJk5dGxH//TkQ6E1/1J/mYv8BdooGIQRb05qbY91cN/ER9J/yDMonZVtwm6yQoyMZwEqpih
ULmYkTlH1tV7fTDADabjJKmmRjF/co0E5v3ztrIIoKOGJP5Eu6MxF621XzuxeBF4p20oKIzhFgzA
WTsrm8WaxCt7Pi6lHx7DAeeArJG2hwfgNYLL69bp3i0Xph4akXF4Aw6jj0GjLGzITM+R5xiObfrm
LbQWJ60otSs5LX0efc8H55FGXJTRZRfN2MWl2KwadwqrfPVRcKkSkgCYAKCSQqAxhRBc5Tzd/MUF
jJt8oqbWsM3IqIrd76NxgWfBa/hkN8Peeo5U3USJhjoJ79tfxQw3w02jFFGUCcI9vcxoDC1hezb/
wTawKn9QBM63StGcW8XaElnAXN1pEeaXMyRbDfjkJOVfKLMVE217RGnBVrBeBbPjhJsGkj0DJCln
naR9TpXmJHWwduIpl5Mm9Ms1Ri1gcgGDw/OrsNrBJtZRUVgCxTMFvjKe7Hx8/XGl7u8wZ4NauSEr
XLbUo6MBTuCDWPz3Fuvb4UxvUEWC/B9YWJAPziy7P6D9MAouJGI2/VZGBOQ1mVIKVclECD847fS4
qQhr+JfDaNtMXwTtmvE/ogIEZmyOah3GZurrh71YJVWueyr93hykckr1SKDB01WaT9qbkl+QmRmd
qrRTc231hzs6JGY/f2Zzs98Gd8xLRlqhkRPtWRdGLxK8+uKEc5HeRFCSPz4S7fPWga8Y3KSLq0bS
cUtC4Lu6EuioaPGNFtbixc52RgAWbp7P6xuiLBkzCBtF8Pl/ruUizEeaLqZHOUKOO3IYTCZrHkIl
/c6Y+Gxy5mKqozA+sI3GBqEYvF8B7wdzJxkioIpvUi7Q6tOCVNIi+f+iFWn31HBYxsCj/HCw6kJ5
5yTEb2QXUczgi4+CwoPPDVtqzxii9Equ1eRkOPxO+GEAzB4S6/fBXhzY6Q3ija5TBENqYz+h0ZYt
9VnlQiO9XrAAVYr+mNTiLa6zM9zdm4KlBiEH9WngBxxMaqMZFW3O2Q5ZVneYX3sUyrD4BIMFDNtw
W768/Hz9BSBHbjdw3XDOBapjH3w0ImpI48aPoTLIZW+tqJkfluvHLcQnMjmc/KatABBgIWOFDis9
sjho9OwJicKrS3YYW3UNTt8EfaoeSjZ0k1DYey/8e9m2/0EdPpw+aUdS1Yk0SFUnnGn/WhjATBiU
NWz1MY4v33eNCl3AILAb5gA08y5pIfhLY2c2ze/Cln1nu3h8Red+q3FIE1C/EOUARKDJr7Kg6qHg
w5BQnV5UZxNq4N3Z/Zd3gOn/mLesS8EmkAGMDZQCLYM6hVTnVjJr3dcC9p+7iJQ/RFRA33NFZrly
n4HRrPdCzzHeShnms9e8BpgHpwrZ/K9y7NmCOe0V2OEJ+xlc2YoZFhw+sOcELmrcawvmkL0UCgR2
r2AtT+cB2B1ehgeqzrgPMInPIefJG8PbSmzQNw0z49cOVtNLAuteTxPrJfc8QpOSS39VxE+2uC2X
wF+TIpA3nsv3gN0KFS0FpPkv2MZH0kW/UwEpXz3WpIwUc+BWA/KUdiIthXYaIbcJPI9zjJdO/N1g
vRVwVbANRTOx7VuYPd8M4BMr70l7v0KyVbgxrvSVbcgiw/YQFsGp7qQ2QcczhAJCsFliaheyPFPC
geGDvzc4ACJafTCFzlyOyvHdAANl7Jzux1iEndoa3EGB5qIt4tfnP3+VPfbQN2CqRW5rYmCTc0Mz
gcIMT7OA5AL1dUUvX5YcWEtcpqovEuF3VfB2p/ekD+Uj4sSBsVFNtCdzBNkWqUr3oFIH8/5rDsD1
U7E4anQ3Z2eGj/XYmvIeMP+uLAv4YfMEM7LHw8+3QfHuc/KrGc9jgOZjoO6GqiAOQ+Lk7Ap+lwye
C7sGDZOd6jePIDniIpaULJUVbNRFYww9c3FXHOWbYwAtFyYlGewCqmSyzRM336Y5eizGAkZoCOru
dsgMQ6mjqtIQnnOqNdVCudVFlc5KPHAidXQMTWAUk6kyo91h9DVWoQQXnXrhYzHODqvUAsMs0aHy
Kc7/XOqdy1kfGPvOF6zgzAtS7ECbfgoA18jfCaHolz2rkN8Vt//SMeE45sUMpMXZWFMfMjzxfr9S
N21kTdEQBbqNNkNUssccYqAflJVToOxR0Mq8KnIeiBosqYmgfIOL+MlOi3rgJL2J9yRWg2F277Ec
J2+dsN+Be9VURmnnYVrUnr1vUesI04GYuTSVNa3dRCudHuydAYA2jQr1znU9gbYq1BUu8p0Njzia
9vs2/Txjlx2VoG4fEZ6rF2jX3AV3s1Zqae4+70qgn/TfpWr6lFxv/tR/QcL16WyIbqKF+PqH3h8z
4eIBqvHUbqEP23qqQ7ce+aFs7EDh5UBwdserPCqfU2H5H/WWp+qCgq7uOgKnwmzbtXbAeJWyjx4g
O/lTruEK7W4vFJ8LR22UcOqfcT9OqFXK2hOiVCMS3MDb3Osm8sCbry2ZnsdiwGcVhmsLNuCZlQ1D
YRYdYkepaew3pkyFwCm6EUuj99x5//+qQTHj0iplKCaJgz0/r1ra1QeYHm6wXQR6LkRmIAZEj+XO
FNBdxbVV+VaNS64oJ5h4KH3+ZnwfIUMbMdG+WpksX2Tk6wO4C9e05taB/1aRwpWz4i3FLb30vRF0
peyaWIMiLQR0SFtfyoJ53sdhMddWOM1JTkUx1C0lfd1+rk8EwDPTDRcVsCCmUHuRjPNWbImXDsaF
T4otTlyc9bp788uCbswFHyFvbgWw+CeDGTAisQ5E0j91hwiDOJmtM9M3EnPjHd9c5+IhydbE9qcO
AEDMNABgdXuJR3MydHan4JZTrfe64AnDgVYJtzq4w0Ccdu1E/U3H8RL3Kf91d6XS4f8nzzf3DWmz
xeW8mz/u1LtOG0BsmUsWeTAbsEPEDf+y0Pu36ejrhGXSGQena5ru1Yn5UKG+gGWCTL/NisQ416bY
aapWTmnScwF4Igg/h30SqvkEO887pM8ornPiKLPAfBHxiMl5pTVmSgh1mB3AybBJ+j40cSOZT6XF
vXtOuFIeWzdpNXjKPwVItVF5Kv4lYvWjhKxwMfyCl99eWarmGEBXC2TyQrBBL/rLJO8fQJwJRmVx
iKHIcK67iN94owDAUk7w6zVzPTmC6b+u7SL1Vnl1wUkai27/u87/13pmQvuKQaKxABmtZ+pH7T1r
WKkXnxwFDXCvZlET7rst8mKaGvdd9hRdXcVrrvZ0TidBFmbfrESED8kjwKhvKRP1kmdIEgxjUAjQ
YeOVfbMheM4JG+VTD1KR/JSCVGcVTdopVT6VFhrqKfjKFHtkF+D/wuC6g+CvS+kjWAV1S2raVChP
UIPR60xzmac2JqKAHqNQ3UJ4zQohdW/2rlEJUCYxaemnaq8MvQ9ufFa2MDnWRmA7NDdWqya1b/7h
owAbDn8iCqdlEapTCcgsh2JrwN56zPHdOzdZlRKAYe1YhWSNgwEWdvqsFEFB6crMULaUL2nQ4wup
juVkewuNUpuDmw7OvZNfja/iesm6aHnLLN77hHlUFFe7tf7t8dp5mGyN88/K0wfH9+2M8t1NrOW5
02RZ1bnSud4vQyzbtZwZNBJtJitdySN+MDqw68hSb7iDwHEbZX8aifO1NgzyDGm+a5lDEAnSCGIY
RJiq/2wRmctWqYYOnM/3AFnWG1lmOSIaPTU1ytJywuBUDWj5zHl/z4GM0XPuJJp1Y28sGyyTIxsI
7xGpFV12CjHzPvgdtzb+LePzDUBeiy/CB00oPrLihlxPsEaRPTUlxVZE7V6/cbJKSUaU3xLYPjK0
QXCN3TaR4PPbjqhRNubl+TrWXkgIp61nP+BsjjvtMs5viWYi7v1WiVuR6kD53cuTOOPG3My5arGi
ovZwaNRLS1uFdpBMcHPCGL/kDLh7fxMJehpbgwAylnywbNZWdg6KPz1kPy6MgkqgHa82gvunMmJ7
l7EZwQkJk8W/xQV752R8cO5CaiL/zRNMr77UlLFr10RGQXMMalvdJsBMEfifCXfEcDX0cvmi7wMv
p/PSoTNxI/ipOJXvtqUsR6SZmapi0mOD+DLRqmhP33p/jGVZV+MwMHPixwHyq2SqaZPAfBdo3arG
NWMRD5cfq1DB7HVYD5gmM/JuSi5CGIn6zqMaRrjDNfTZ1FMT1evclZYTFzH042eb66p+li+exXyk
0QZwuBS84XO8JGDTGJ35chdOWphZ3XBxQWIJ0lG2Ak07SaWjyA5PLL8RFTqAcLJdV99B3UEEKzrW
q2zCfGsBNHMEQ6tuq/O0Umi5co77U93bjk3EZNlRsu9MLz9oInpiRwXcxRUVYd9tYbJXOI58XQ8I
S+4hNYBtyy4W/TGho86Bpoy1HuVuVy/DyOT8Ypw3VVWB7EBuNjnkxqC898XcQoMKhH7B5WOp5NWo
QrYmAjVClMgtahJ91I2uqkr4F3eYO4n08lD1jx1hczTonSCC41gPDVe7rtk8fvJkdOy3UUSoPVVO
me+ClYEiYS1f6rMdMrRNKkoA1MXCzeIsnNdGIfykYD6TRO48+H9JqQqMVnFXvW/xder6matW0ITP
wqXFMbgLQrC8SEZvQ6xIUrLOT50MUeSx7S3vUUZPBACvIxuyz36ZcvW0eDX14QjxmcLSWCkpflTb
0/4rwyKh041fBHa1fjMsDrqUBZ5MpjlqYBsq/0a6xBzywSAmOlk92a+suAW8bnr/RoxnqaO0mA3I
iIGhOWmmHztITal6wjYb+ZsUWcoudKmQgihnEnMmFiR5jnMuvSnm42JkyYlD12dk2jcGndj0dT4Z
h1oIx1jtDtL+CU9LRj+vJcKEPKF3X7L/YIwTqmYa10DIL4/NXeHfk0XG6AsUj3Picw4U3HmrRGDG
SEP+OWgjpwvlh+8oF0/fy3BmpqcoI9anOxliIJC3w6m6y1nT4XY6456akI/tVDR/7kKAAam3FPaR
LjkvKOHFNcYDKq++EriueGAjtJDD52Gf0ucoBnxdGEWfVEZrvcX269Fw2Atv0BNXVlfazC0SweMn
Gs6Lq3LtGZ0US6cxEJzldcuDRz6n8kfknC0J/XKIoQCbMD/aoTYDkqHyItMqOXkmFrLhYjkbgh4R
7GJnOlI3X7tXVFyBna8B103aSvv7PogcuYcAfrefWR1awbBz/OLwC5TYMsQHcSAw69/4M+Nj4kAG
xt3EXnBG+sZUJfjQZ201/hipM2bFKB+a8IMPYyWqTj81z9ovCZkzw4RCWhls7iLjowPQqDRvkpIv
ZJZjUSmt5vGk1kL64vije7PbnN+UplC9YCMKipQm+CofP1n2GoUteY7ksv70obyAaFAtulWEs4tv
jE4MoIcClSeUEl5PJo6+SCIUT5Gu2dEBZIa7jjms7i5eCaF39bxcTy3YAVW9TjCFjqx/fOZuV1sk
jJb3dXvxZPs63M9r73n6SvWroVHVVvhe328TB7L6V8D4KC4qoSSy/5LJhPOIOttCAP/fsMIWd82Q
q2b/JIdheI7AbmgYJe2KFa6BYcn2Q+hCFakfvHLYjEeXRCMbLYxvjFEfb6f/yobvt/MKMTJL291A
wOMkOPM/M6grRztnNTEZJ6QpnkL5td+N0/dDUx1mPrzN5cyhIdQ70c9Ob9Nu8N7LrZI+PIYNXFY6
CqL7ayDyf1BPePMddbcqTqe1kCrRqs+fc28qApvAktHvZyvsyJZSuY3n4xwHdNkjeFxQEIBP1wja
hujFYdyj24e9SGOryWv/ZUKTGpfIJ1MiZoCNhbm1GyNU/mpoBfiFC27EhLfrn2eTL9NRDEhRNni5
xLfrmqjfO9HzKaaMIJpNbbjV7S0dVMiQg5s9c44IiuQiWu6q8QR8Zk9hmHVS7VgkGclVlTKwFE26
B4mVKUcy/rhrY+MpqTAobCxFO74lTPUC4fSpLFiM6jyqdhXS20GMqar08AyYIjeD6O1Njk1BT15A
NLN0K1HhmK10DFo0jrNFXTOo5CZMJ/jQ1+iI8o/FwxUpOwmOnA/TZ57p1Qu+SpfCHLkqNRpTmgmV
hEseekZna1DeiGT23KPuKiT7Gnf7/1GKUftmaDkqvR4RvRrQB8bIu13lsY4o5vMvdDKrhmGv/2Ma
DUI/Ufak0ezQb6Z4kqAevuItFubxj4OjUbp0xXJdy7W+MeQWhn6neYlFdHy+6jaLPkfLdvIPuGho
KGFos3ZxSj3sAIgNtZj5SBkhSTJkuFlEBU9WfLWv3zDDbMcARZPUUeDu2mZsXg3g3jCtiNyLgSKr
UgBRsa5B+bjYeK0MOUbg7LZk1FuKKFaBdIPHkPKEEMaDZkGVVz+rc85T/Q79SJc7QMKRUQKR+ZqD
MpqfrMzT8IMiHsu0FcW/LEayLtw+nGzl21YdlUarmQTFAy3wA3s3pq3Q4zoweDZdcIY4GfGm4xqp
tXboS5MQzM90y1Bx7w8wfl6+hefEuvHkUkMoH811bPQ5npcwq9Iz7iIBBzjK/pBVaqWn1L49Q92g
/tEvnMZtlLjZfbHD7gHFd53pm2tYpXMKYidNEYRBW8RPPumOeMYLY1DQVs9CHcFAqQBltIiTPs2V
5oWX3sJR8jE8e5pWkPE3A9JulK5QpnvRm9f1QekrRnhS8zXkALDM2Enx6dGTBRD/Mh7KHjNoJJ2K
682yJTkR9f8t9YVpahv+lVd1naJ5yNjPQ9teAqZHVACvIl3+1FNuiVOZcK0I3pSDR6tvZGiC6g9g
GNgaMd+nB+B174eFA5drpE5zw1uJjdU0ntILJBBk/FBjI3uOhAc7she8+sBSjTc8vaM0dEg0cgdk
sKfwsofbBIE+qQUmOlaWJToveona9uffKWwR7Bhl8MKERdOs71cNmLJtQSqBDrF36Y3/vHbxjTDh
MRe7Jgd93yA3ujaCDZ4/EcJyChj4/djKKVt2tv2UrZPv9t8ycf72P4g4S8yfKEfwVU/nHt92O44J
+K6fFm3iEj7Kfy87bixaXLU+g7QYk/6hMppBxsYmVYq7NNY4cDNtgRgLGBKqBca75wo/JNfJzBXu
+u5cNkZPrYQMyHWWelXeX5bzTM8iOsal7DrM6AjityZM/Kg4DQ9Lu+g+4S9cwOpqgkxmbhWQjlSH
pD3Yq59p+Hf0FhAD4/VVvg8lka4scQqQ1Inr7Sym5oUO3Nj3cZwt6Fbqfn77gnGvNd/0Ljb4QkT9
8Ag0gU5TQuTVmJNTauhQgFYS99NDAe5MzCIoLUFAJyVLawftVFRyOu0Xe9dyQyxDM42bTuPPR86b
I/PIXb3TOiWSE4otZUNvYoTAJ953iZFsaXrl3bOIyU6BeIkY/O6Uem4egYFWkBoARCD4+Wfs791u
KR4iG4EkS0vrayCRLVwQLhzg+d/56s6jdY8GNJpRy0q2TvciWwCpcJwXySLiaRiZ76M/GVjjScrR
iPWpDUOHO1rp+ywcb3A1oo3cSVbPE159eO8t1wGpLOOg2Cv+r1KjXIBh5sdJd+BZJe0osiUyBNpr
uc2mzEPkDKGejVlbDHzOdYP4m6hWSX5Rv0tJ6RofpbiVMo5Rx4CsVragdVIW7j4PIk4VXPOccjgF
cZeAUBK9GqR4tZ36VFkfINX42KiKxDHQcO+ZXkcVPvHcru/fF7L3oHEUjnStT9Z09H5twiy7jPzu
tnT99Am8QF8JVvrLwWw1PT6U1c7vdE3Iz9hsof4Q2F4Hdg2k2nGNoGNfZcZttDhgqHla2hvDrGK8
hr5LXgKMMtJ67Ofy8HywM0u5GLFuUhUflNS7X1ZekC1DaSFB8RZK73krDrNOIFQmfXFXbANkZy0E
va4ri08BpGUkGceFXafnX4P0kDFNQ6paaQx/vugO69iMII29MyrYfCePKk6z5nkKdaapqIZSL97P
sbnbRNahxBTJqNLxJa1RcswHHW+lggLMlYpOfFtMW5qErAIc6qhzFt8TC2YAuMMSZHTQrweMyV61
8TQNas6ZqiyWXAm1IB/W7s7ViMtzZjxN3KNDTgM94isgV1OzyY/ALWBFgKibFkVHP9O0dUmtP4z3
1SC8NpHwiPmViBLOwZIqxzwqX0MZZp6lcCASqu4OC2+fRhX/wIq+CGCwB4onrADvE9NWuSy0N1sB
70JX5PFgHvNhrHvOVftvwLcRDkBhqoXyk9pJUwnoiwIuWFjJ2gsAYFX5YdcKSID5jXldvijeV6Hs
iC+l7bfRHA2vfywgL9Y3WmtUbGxQVQi3t/M1D6fsmput+5NOE4U320bpxnsSHQvdQ3HA/o3Rq9US
ax5W+4vf3YGMQ1P4x2T/FHzPC+/iUtjq8GgSQjF5YsnDPFaRrFKANzLv/zULzY8jPjxGrf4yVyc+
2aKts/UwmcOQGOk3LWk2l4UL7SoLkYG1DhgZoy/Gju5uRraFHfqCD6Dzo8dpYExhSdcgA8hqW3cR
D0VgS+u8fN7ixWJqbSWAIIemXigk3yPgzRFJmNe6KzMasFikU0CYm1Zcsrz3CcWFTWNit9jLk/cZ
Sf5R7NIKKfStqciSSqwCDMAuD1H5s09mFkX4EBbZI0qoDkDMHNgUB5bdPiqnBhozrNLEpT5p8lfX
AIfNDHrLx9cijHveoIj5fcp733S5S8hWblG6TR4zscbyNN/T2DsW+0Tey7mkn7VqdtXrZNZN4okc
0QPszyPdyMsN8+iaBdp4q46EZqOafJxa5S7qGw6UeYIxBdMObEV3cz/cVYFXefILc3TowAFKrprY
Dl7DMa6NSnvpEXqBLZjK4Jb68Mh1guFg4MWL3NF7LylTybntk2FKeIeuIZxutjf0CtEpYnpo9bc3
9MO+3YOBaVduN5Ld5XwT7I8EAm/OSwcw3D2KVjvf93969Bi1dFfy9ObRk+k2Bvvh9kRKuDZzwbN5
YGDjE0IldU47TtjXJPXGLGcHyUHaZTLi6iQgzXwnmwiiXXZoxVHHdUUCQ9uoWZ7WqiTwHZfzCsTR
TIKqezxsqbyuAdI3mlGd1YQjZD5ro9BdwJs04R3QxB0/s4BRvZvS+BCzPXWYLaoEUwDDWFpGoec/
xp+qaXty3cNskn+XBMuUnFUuvXhJHzLZmJHLBub2jUp85vP4oSPSV2a9rQYaodPDjzyc14MI2Eg0
8OjQ7R6A5flDDY/hnzGKprScjKFR52OWGQtztE8EhiQXnWEGxYoAIY7EKCzSxpy4PP1B0H31B7Md
c/JGjWwdCAlYfQ+IQ+I8g7oJwpvt/PerTlzD/uqFGMNA+Q7gF6mXVQJI6oV9LHVW2zFyWEYIiVXo
TEV+Whf+ZZggRJzDZQ2I++tbOL4nNpa49lssjVb52dZ+Gvpsi5UKy93icBzvVtZO5YfeIqjB2Iua
TeguExUauh1sYUxFBM5+WPt/QB7NQ0K/tYXdcCH2NH6Mt6qZXLZ3D62oNTJs/4xXVhrHhz5NExMY
a8g1CnyfR+B8qw9DDIKK8QoxCwM8aNDHWOUwWSdaesH+I2zoWPYqALmGNph8tjNeUouErpKj3qq1
+CgZ1s10r5J/2XkMM9Ht1FnfscIL4uk+lpWWcFzJd/66wf7UmpOzfnYyWvD6xfx2hLgg0c6Y9+0p
WJFkMI/vRzTpMTxfxANA/YhkD+DWh/cpAj9VVS2Es+LjNBuCtcxMa1QKt9zFN6ywLRXx3AO54UH/
HpAVYosBATPdDE8GmGBeBYIJqQBf/ObsmyMGpOdws9BKOqzMdbESLsTFDwQDSnIh/f/ixMxH+R8F
D1JVxTQJnfUXwsJrv9lsSr8dEjTkXoGUXHZrradyKK57Pvb2e1bwriz1FRkdKa64JpmVUmeCBMiR
iC7eRrKCHTxOpr8V3gHzzVP5KWzKtr/5i24Qkrfqn1E909FC54tKp8GYk4vl2dH9S+QMa3xrcHge
ekOBA1ZobDfApcehf4Al5X8A0A9tveuV65tUS5s5wSrInomK3s+rX3bq+ecf/tBFG9uQ3mWEi1iJ
VCTw1ZHQgZ4Td25zau64D2nf9Tr4lg7CyOW1tagG0nG3+RszMH+rlNU7M5gKVL0cqZ5THCouR/wS
Ia0jAGhjDAvrkVzn6eYSAjh6CTZLEb3A3haVlBmhLBKD8RSZ1aVqrXOUPTGjcwMDg0kyKFivF+UM
nrw0CgQtEaTLOcE7+BEdlY7JE1vGJ+uEGmd68Pof2W0G1nKg6P8rD3ZsovG1Hq56inYw4rx/YJ2+
QxWwjrHZjj8AELoAbaxPIpov3jT0hYK3EVgMLB+5pPobIAskG5nXjpxT0eLEybCic4++I22tBOcO
gPCMm4NZkjpt5tvJXbH26U9/I0Q7UEk9ytYuVFnhUB/WSXewAfLcSMWbuMuhZ02vWdA4hhziUahT
yPLWg4jQXn6dVdLMXxVmktVQMvdMP7aEv3vYehk6RxmQN1VeS2e7OZho2hKYzN5+ajgqsOEBR3Re
YqK6XgESdkGXQSs+edRQOp/9E6phkqcbjmrOwrwc3r2jXMlerts6jBjEBfkbEBeo1WtMIGoadLjm
B0XXbPowiCyNogsqrVtsO0zFs46IE4ZW+8Z7KFgQh8FG52z6dfbpDApeD9TV58ywFiLpolDbQwUa
3ihdOIvlMVLbpr1Yd9hRYT2vzeqqvbsYQ/tINM7hzZ5HbXbd6yshhJSKysNjOSMwJ6aFPUrWelK3
xqQnPPyU98/7U+kXzLqkfTBHugG6GOHHUUZwfWEMfdV+S1NeJGoT0fKUJeY8Ozzx8kuJSHOMCGh+
pN7r57OX+mxS+8TCpMpf3vcKwhN/PncTVQRHcA0oB+9soeMrvVqK8A7tJOJihnxAvy5wNuqj0w+8
zc4pLy2mT++NhcyWH4rbh5HCSunxiyfNgWMxDU7mAvkn8Kh+/xRnQJd6MMMq6kZBCsb3KhCHBuBq
AQeKCM3QZ+FkRfhAyPA6b2MhXa+Q9SIG1l+9fN24QHashn6Qh+Sk8abDwahpVmw/IVGMETi2RdH1
hRwO21GjL8UNGiBJ49YwjsjyyhtdGnZTg/EBcV9M/LHoRvDaTQUJPEIwRZuvmRuEtsA/QwdzqNmk
KcLWrEXWzCxX9LNmGnOh84fTMtTgTy+HciUpEWYMu1BrCLqTcywctiWKA1sj632/6RaraakAew9Z
KC9YKLo83Tbuf/WebX0FF2YLN0dpdb8n9xV7i6S3Zfqab0BczJCUbvwy4OVkWyImTQ95zx94vGgo
2X2o6V9whKf19kyzpQ2DtSTBixV51CPncpCPPww2vSXSrk8Wtofm03r4R4dQIQBFt0+qpT7lcv8d
FR5cfi+mu3gaTZ8y9NxNxsQTjBVtN71mm9RqWXvLMnfXmEtBg+zceNcjx/sHtL4bPo8mSmG7bNAt
wnV19PtQ1J/OpxIQ3WL2zH+gNAqLwfCvY8/LWSMCO9++K/JtnVr75OsahAejvtKiF+b2zKDF09RH
NMsDhk0TKaAJ9BZqnZdSo9sas0o+7fG7tqZyjOWZb1AEcH7AHurJJKzVZFRNUhWD7G3ImO/mU9w8
Lg7fDZnTwdzHxJZiKMQ+HBGo80wxmR4gTTfuvrQnxsp0UaDY3hSZo9lrEAaH32GGYA4yZmoyQUr8
eTifPPFKRdryFO5kQuLq8LDw+vpIO7Q2+4dcY5JG1Xd8Vu0jEqt6hDjFvd+MkvncrYlM5C/gzjPK
tREoVgnd6CXIKnPV7y4Xzt5VTZ2lP8xEnXuWyTO3rLb21CZQPAfulskR9B4wSm6GZr0TCTyV4l2E
CgPXYCxyZxYP483JXfo4wqH9xxP0Lv/pCg3qcbrSixYQ/s90KTna5/vKCjUhfne8U/NINAFwhY3w
jVTiNyeF3XFBDli/aVnpFB+4p3WyEVi4NTXXh7U5AlMFHVXyTbVuoqAuW7564aqPdZMkQM7r0SBY
xqicAnWhPrS7FSgTqHqNxewzMAwVwfQghBn4lL7XACIPOWKVp6cl4x93c3MOHVpGOacCh1xpWWRQ
9VkMPvPdOTwKI6QpNpx7TqFjYXdwHi4hBG3d5TiDqXd2xCSHEflroHBn3+tI2qcbHQjYNgf5QD1Q
5Mhlhjam+PmrABBzpOB/KJsETuyMjaY2ZhWYeZOU4F64CjsB53/teOMwHu/PXbJ3LEP0rRrMYCLC
y4o6VkpSbMAcIqMbtvB2MyUfag3TkLDLidMYkQOetG91N65D2msXV+tX+gLXUdLJuWircYoTw2jH
FQf8FXhjFortAiA+o+Usyve4r7p2LQYbVQpqQywXfMZFJB0cT9XLYZTK44JgINgwsBkLv4UWya7m
3qTRHOawx2ATSGBORoo8fdCDqZJjjif3rkcuYjd9ydmbCtLgdLwL99RCWHK75KR6NpKGKAxc8fJT
Kmm5qUtQ+BWrRDq5GIFsPrUPxQzBm0DGP4NQffrXCES/flQIwQClCgqswaihVybAQQZkizxTA031
JcQ93G7d/u/2uECteqKYU/E6doeVVgHBZ8ih6xYaDsAKu7hvh0f2lYbsdtnIaQIECO17pJkmM2Bf
mvBH2U5FJa4E5/YNE551WjfKBKdKPcKhU5RR8QjRR7gvqzJvCziEd3uanTcKFJOQMBvDtE+cnR0v
T4xCPnJ1BfNcdjroKjC90j3ZZqH3o8Mg/GVENbMYT0CeMsochuichAQUWMgjiCv9jxlf4J1qeIca
44RM2jdeoTcwZ8neJdoYN1nWUkJi7y4Zn24XsYKZ7jI6SFr9cIdw9vJIlEPaJZhGNAu+WZmNa5q0
zOcIuBkBwYU7zr0jOdITrC40dD0w9EuT86H/g9bFX/TIvd50WgkEgkgkKAW59cADlG8dnfXwj1WH
qzH46IIy23Ve9PfsVK1HjjB6IGdxFUhJbeVPjNEgDVLKVrkuiereqJmcUDS4oy7JTRjyIcFipU9y
4qTO0XPm2MvybWzjCwDrttP14xqKb69SfaCgJtNryBjnkS6nnVGTM25ppfKd1lCAWTKiAhQ+83tf
IZCgmpr6YHKT/ge9mb/0S+xJwZq6NmwhSCj1f0vv5fBQ7TFoV3pFtlONZq9KvZZW1cYmLSzZV3Oh
H4gisfA8n6VDQM0G5edScTtJgrZwkLE7ZyPJKMI9ZkWm0F+EzX4lB2MyYtHFqW7wz+Kijhk4Nr82
WCugZ0/rKUC1fK8tFUIMoGRgRJna52g8plwC07WA38sQU696InCjt/MIX7hwJQFcdTii0M8L9CfA
CRbMFhMb0LD757VZhGqTbRH/+xivrQmsjGWIjtNsodYAzhYtmNP0YVfOduOGmsAVg1DMlEaoyD3H
4OiWJj8MbU9zfttswwM6NtQsbsKF32udaubWq9JKyDq6LuwSr1fvbdOXrvCPvds6rfI+XZ6zP9yh
g06cY39Ddwsa+vZdwSEmkUfZJG4KEC5qQYz2yjKU69YjbqBLunVT6t2PHEvS3KetPTHmshPOChML
NQoEwheLeeNe4LO8wZIlyPnmdybGD6zyGEo+YmPVO7VnCi6VxJ/48M3iheVMqxUvChq9jgm1Okob
By2RtbfnzwDS+/XSgBXE9J0FBRsBY0fK0ofjcFo4A/Q+IgXX93E93VvlLbhVWv6F0m9cERzjTRJz
kO+BV4tvRYIyFyhcj0V16prT+vPVzoTFTdrR0P2mjX/TztvCURCsXKToHHkPkniwz6xFPkkmHX4s
d280Baa9fKfJ9I+fjWBXLtJ62HnJw83SU3zeYDLPUDerbVcrJryS8TNw4dEY7RXD78j8tENeILZo
yB3tMCfu4vivGmwiWKa56XIAAff5uTuSOMQaQvjYrjCZFIN98ZsdgpGXKdR4aocqoLAp98nVbzy8
iQ8d9OIHn1B/mGzhHv2V3v3xRsHNoW+XN/lt8Rqn1zL2k7PLUJFPFIecelYU3cmMnFdoib9JfiRX
yKJEHeSULrOFyCdcLWbdlfYo85RHwgYJ2fV+b3tn7NJZFUzdeDr6HtX68W1b0+zZJkfmPNGiFdOi
6juZHgbLhIz2UStcx3HKzvNw6HH7ttRKr4fThOXIm77NgQkEfGo5Txk4kAm7CQr3JeRuufC3YuWr
wYj0g3FIsAuFJfzH3KiB78Ss/7CHfnbXArzEj/o7/3Rork/ba1bdtwHdMaYTncmYBk4bcvBud4/3
Xuf7sDZuz1sTC7gtvqneuWStm8Zrz3k6I4UCrvUYplfki5mbBfWvJYe6z9D3G9sKnyDiX1bjiJNz
aw24LgG4owqp+l/U9345cR0gpgU71WYtgl76SIIB2mJx9FAuCyFx7jxf7KS7pQ6We6AL3fYjRyF0
wzWgAS+QvRPhbc4mG568dNrJdc1ZM+en0knfpxT6UzVOxgmnDmacHQcZjKT2j53RIb14ol5fmQ1W
gO5ehZkQuTH0vM3DdvBT9870s/CiziOtxVKh78tSF2DWFRWlHCsMy+GRskbfrL46KiYuuM5Mvz5A
B0Vq/QljkxGCXBEqTvnvx/8RdGFVvl3mXcrEDxlR00KlMrwoHnp/+g9jlVnGTeg8fH+8Y2vgPjJm
aYM/dd1CJHmudxEBzWRD4C1okY1V89lJ6MW1qavDOAHoLiaL9CT3zC/vw50vQgATza05FjMZDoL0
iwoN0HVvy8bOXx/p7RtHelMVKcmVGjDZPb43ofrjOs/uz9JRckMZqXqR4oMXg37SKZfXTs+eEiM9
XCw8Q0RncPr1LV5+dC01H4YBlcB1aRh0M3ujSESASdhZifQKCrvjUfbKt8lqIKDJavShLmFHrDT7
IInyiQ9n2y4y0z4UnEhvZV6QsyIU45UKe+/ULvt3hRUcZNlq4S1iO9zswvk8sar5wTzqjK1XLLbf
nTsUn6xeIRrS9LR6cRpPy+cT5xIF8ns5Z4jSxOVNsoqSSBH7dbyZm4nM/b/nyr9nm/C6rSsO2hRk
pptUcy83iTBBUP/ePU4iRh5bsjb5op6D7ZTlOYsafSGHxv7niRN31YfwOCfjJPeG33XIqi+xcAiM
ui4XpDuTUrW5lqymp8Hq99AfemBI9a5W6no1Sygmg2oEFLY2tr7Dz3YiFSf2JCS2vqGG6SQqUtWP
eHGRG/aLhdh36ksiXcRFSvucAUhAGrhEzt+CkPDq90SZonfHDIR5MCBSSSl69Z4lbJv3rS8JAImh
5seFc1Fgj6OOQFvrWwKfRo9f0xjalLLhW00whPrskqii+Wq6Xdh/iWympOpsxUum7M8u4k/1c/ST
NEC4EfdZpKJUjKCv5av8z0clyEDtTMuLSYFBIc6/q5HMVSbGqfOc/fZ/7B7cwncK4JFKPxQ9cdQ3
be+I26NCSsBhB2+RcweAqFEBkjqW4N4owkMfFqrKOrpdkm78uwwnASeYQCSRuOQWQvQyceO/oq66
4NykndMoknsSY+9Q/pQL7+WKOFsf0P6rYbvquEiHc7ekgKnCoQnXcKP6pU0Cc8IrZpLarffD4cfu
dLkciYRN5PY4SnuSAqBN5QahjI332L/XPyqKvtwnem3liL/HC8EVFlM9guDS3gA9PJkAzIFeZJvK
6bT64Px8UHCvbWgX8pQOxRkvJTFE5zuGp49m2HydkzIvJEeBM1oIlsAxpfwV9bulq3qQ7YAzq0rB
RZYf/ciIsr6nMsFqsg5TMgiBWPBBTbwfH9nVqT7bOrLqaOMQ4gNkTwQTsnRZRkOetmCWtF/dtBBo
GMhakHzamCMBLsgRUY110rQcjmmiMlw/2S5LKtU+wyaqzKrnZJqkXN/mIlNMVisJF8wAGKALryyp
uwCeDFnsYtnLJXc4PP9ZpdpizkJTWNk/vSNW7z6XmtWGCOtari6ElT3HB2J6oGMrBSlPPGwpOrBq
nEnBTEoXy6V1uTSI+tfCcGzpSBGxhcsYkwYvcFOpYY8ONTtxo6ddJhJHaRvUmeSSgBwOWkRXFjyh
qvNawSxjToGQ9Mp199EUt9jO1TToCJ+iTO4nzQZFZrnKxM2qw+1uIgYfJYvOFpjBnRbdMiE7teTt
3Oici2Wa0xYMiyIQ/xljrhKZy05hZSRCToUn/Q6ko7W/13BxSFkchx3ugp3SLTn6ZcFkFjv6jSnq
ks0++lss9/7nkTkODIgdTJYPsX2QL6INK4bv/jUmljd5K368nAHsDOREcUhUH4umPZLv9uJd2e2z
L/OqrrJYBIjryz+SG0++NXcCyUFg/DLyoN0imh+t4xFGk/n1GSj3e55sCTnTs5m/A6kg5rMx5wd1
8W0pU8PVKi0Q2Im8+ufPnUQYCT6kAtP8dbTBvvxJ1EfT5Vo3nbfpE1r0iFJyYPuUu0HhAUQKmKeI
cwlFWTFRvGCW3qiUB5ueDcTL0kGBFvQ3qIpeWtGSvxIXAj/WuMJmQcGNC4OKREXbEwfSWGbIG0+2
W2I2mj95ZzGUp4ID3fxhyEZtk3RPH/2KLxomCJFJ1SnlWsL+0HrTUJQA+zSDdmaBICi9CTLbtxlx
WfXkP1MzA03rJ4fLpfq3M6lMCghYtZ5/ePNxFGt85yXTVf1kmhkoq2XI08PtX8Ml/fOOBiyMWJUy
drFbN8m3hFpcD2oAHLKyyt6Qks7rmCIDSn3TVzIhMFmJEN81Vl25ziHP190JZPND7sHMboN8NMs2
dDl1y6ypoKWbitUf1Oc8uO7uSX7rmZ8YM7uROxd52lJ+RCT5SexFTY9xvci6IFcXIIhI98Sn7CMw
6pExM5BseP2SOLBN5NHp41gMi+JvgxhFj4Im+YDlWQJStpCcai9bxFcefARr9+CQ4A+iVZeOL5Yy
5H26lc6sTP6dOSFNd1Wfk5KpcmfZW79wSzq/WUGt2O8Yoe2+GU03BEjSZ1ov69GtY9gETZPtmC6Z
BvnlZ8tC8sc8QDeAN+nmz7zqHJk0Q/GNul+rv9bLUqfP/FtYy6E4KiWG5NCwPga6UiscCMFvOJ7R
zeKRCiXNPgcng3U+FCNCcwTS0ElXkW8wFCUz2Yw1JTSUvkFjyaaLcQDAqrr3YmeLX/6MeVkxNCbF
ReMvAVHCUHiQUfQf4gG25NbO/lr9KN5KXngxK/tIKnig9SjmDeL6knlPtfznFSHt4eoUnoovxOVX
nbU8ylrODwN3HlsR5GEVrIOCBZFYTNgLPqxe6hH9dlmcc9cwhQsbHSdHIx4pB3UAREfAvKsp4qz0
Ba905RQRtc9plD6jGGoT8HUj6ayLJeA8J0xOJr034oPn+b2FRo90xxHOGZ+LWQh7wksRZKCYFxMy
QEQ5ryG4V1ZNtsNZH3m2ODjR/YDQqdIzQ2q+m/cPjupLuy0i1UtweHSmJcJL3Q33NhsF9GrKTtup
rU+qrK83D5q9+RxfIZbfdDNZz0tk+c0FGGQnaNAibiTUxMnykr6xqrKDX9PIpHFjfwaaFoQ7aTeZ
qtsJLStpBQBXOxN67gk197Ii3sFpXlOxmoz5tObQaLMTFtTNr0Oj78oZ48ldSPRhuVUUWvV1rxHi
1iOVo2RA3b95qmueK7nElwLt1fJq5Wg30VX5oi7gJxCzCWtmECIvSLHdoI80Jx1vhzHHZoOvThfm
ui6Z6JOkqz1P1BrLBSIkN6rIiYycCAR6f+zNQ11iLzjoa7SDaFYH0mVv8kp2GQu9ABqus3R9syTl
6kblPaafLCoPcLxPEDHM9EYH8fGb+6NrqdKPxOJsLr79WginWXk4JF7Oa5Ae14Lzgv7n8aUpomVo
vMtAt2tLr08S5tq5ErMV9RIgx1Kb4Qg43hrgWzzV4k5QtkmKnOpGCnJfMbteVXeL3klxksYNMaEJ
0MdOpu2H235MvlCJVbtK1EkY/Tz6tPlvAnQ48jWHbeouwNjXSsJqN9VKppYqYuyifqD85eCsGz73
7bR2fI6xiKMjrh1kyRe6GCYigLD8giALru3GIE4Wyf0vO4H/EHz3KRhyNaYdizjFEso3B/TagrkT
jTG3QmppXuEI+m43hc/w1tny8oQ20HYSXPKQEK3SYntP/qAdum9p5bkhoRloZE5CyOb32XfK5U0x
HqsKvb3PZr/Opi95rNqb2Kn9VW2xQMdH/l6fdcUDYPRHFy8bANGcVZMcvETZLdBCl0+XYlm6UbP8
FV1PT0HIA7etAq+ZtqXdjvMJXuTYp93KWdAuEQomQZ0o05b6VWWnsl/QOUFgYTlOgUVm1PmUgp3Y
LPzunFLQs8Tj0J51Ve0OEtjHz76OZy+AAKPvSN2VjREV/wjPUgh7XI6CdYI5HkLYFzuIQMpXM79c
veC/NJr4edYBNzQ0lOrq2gRrsAoe8qimfKnJSmjc/OA1XDiJoqYXXwEZDLs90UUh9nqFrXDl3Pfa
6wvyjlzBYACAY9ukNtHXW0u7CYaUtucFZ1DjiM8Qa+JrMLYuKMh4AC6Na8fUNvvPi4IVHBv+3NfZ
+uLi85lZIbqY3Q+KZZhKFaRo88lzYC37073ppgAaIJHsRCQcAJOxVIlKUqEaKS2drfEpe+nUkw20
cqc1P2CsBELmNbDbG1saBYajDRrtrB1m9DBNmLnZ/BEsEN9BIHns8Umu7qrU2M8PaLuC5+wS4o4I
RzO7noaurARGbmU+JekC+Usad8iFEXCeDZLgRutglRRo/CYyhB2BLy36qMcndeon9J8FX7kT9aer
9ypddUUYJE9NPr5GpJQjFx38od0PrAZX2aIjFVj4RCNdOZS0vViTkTOe70RMqff4HtgRffpVOrnD
Yk+RxbFvb5vScCQvCQ4rgDWdPrleLk1vd5bFVDOle835hP5RwfHDJi8E2DHQyWbNsBAM9zIMwEXt
L4EKLl6nUh5ao2Q2pKxLPtGgwa0zF7XyGvGVeeo/Sx3GFYJCSl345ljiw/6fttK9FFb4R3J9JyHJ
2DyBXhLziGxpQupTNtBvNO/USIaLXuBNZfuG69ugutGa9GKMxbQOzpsw2OaDQM2HgEAviyPToLrS
a1aQfUroGg9/rw2Lp18R3cdNhH/FmQ/WCAAog0M2GOnHVkXYiqWupSI8GL3GA2ebdTELAGdcJ/HT
lILY/zE78nKVT0MTfRIbwSjZT1SCl3kXzgHSb1Yz10qvTkZjiOfdb0VKLzLKl15s/FwZAgibkUQB
EUAydk6hMftaSaVOPbLLjkmoDcr2dhMantpKi00KsIskxVgDag0m/TtKGJyvbR1dOUciqB9wlMsj
ab/yUglRg7yyFi1rmDNaTExKevFNs5L0cdYyLFL+wd3achNRYesIurM+e6RUDx3RzxlzfHDVO345
xgIz+ui8YtpFH95Zh4TY/PNRh5i1He5cUIzI9vNps3YszDRyBYJDk7mpW9DcKvSjulkj+A8895kB
XuYzc9SKOYAv4V31zIEiRBwCt94FC8vhZZmo0QACOlMbZnL472u7Z33SkA/zaXIvwvLgflXMTtKA
iB+DDJI7dmMlhBYYXyyu1kC3iJ73pun3wZDFeNHt7diCJKqaZZIC0ryo0JEpNcNMB+OqpuYcxPGZ
berfR6bfDetdTcJ4nLhdraQD/rijoSMalS5QpQdtbk/antQNsL47+cVBsPuVxq1J/jPXxVEmXdKi
RYO4/m8CFS87mEi1mbTm0Hfa8eiokcaZwkA8JVIV1dGvQORSR/C0XaHBd9Gb2tMxqZ1/9LXhtylq
816wVqIWuYN1Sr/FMoDq0T5at9eSqN1xyoHzqmbah56pP5oZKURwvsYSF21REseZxGAZhHoApcfo
Ftl8lcE3F2AjcgdNcdBohFb14wh3TaCbY1beVroUR0jQPXNizc4b+Uwg90KFwPw6JUteht41ZalM
yrB19O3pO/2/KlR86uX736eiCz5pq7ktsKvmSsynSuxQVapLuC8RG7/DNrO4ZSEF667p2JLYXzxh
HvdllcKM7/rQ070oEBh4lJky8c7UIYK8nmpdSSaM4tZjlid4Z29IL+bLf2Jc1lsI4cyCKDk2GvLL
bo9VJgLFR2rw/QwNJLzd5Q0p2u1GkE13j1bBVzRS57f0mlrS1a8TQmAgdF8Jgt2wgHtwqFdMJA9X
EEz15t6f2dHDw3kHOojzfXydXzzPf4+X2NifQCgas5X1+WgbiA4ze/1MsGZWBUTz9XkUNsblJlQ6
mfUT3rpxoYouMFFWlJfpQeY1MWTNYqFFGzTPad/RW9Nmu4fCO6k9/1GfZ8yXCgnz1R7tob8Tulkh
tKlqO3SRL8piJ8bgQUbbSOrQnNaLSEdz4+MlC4XMsNolMxkMxkVSHGEDONuG2a9eo2GGPt0sowkU
pJYcg5jqGIN9lPX7cvajM+V8XZzyWSbLw39GDTo6sduhQCyD0p+4EqrRf+ZgvpUuYhw9uORHYRfc
EgTik6mIHlmbU87HRrNwfgnJbkuXa68aee161Q0p9dsMGG3e6j3ssrplAfPNu4lJvYFwNVTg73sA
JbatS2vVKeYeJTfeQPtbZnyeV+eI0MTdbJ/qRnONo696pjq0FKO47O9Sg1lbs0ncglL0BRTXCHoE
ZZx1MdRD+ImRR54v1ehFkWFE7rtUB7QLm4rBqEnuTnk1ZODLAB3iiFIeqMU/KHjQD0tkNL2rAGV4
1VZpP7exSwbMV8aLy11nPtykb9XyxVkEGVPw5ybU2gt+c/5J9OAbZvHudxu6bYs162bp5kFQvd/6
GZq7xpw4JVxPpGI7c1FddFZtmUqRcvFXYF11Yu3ck5KMWuRdc8Am0WeCNbhYSbKvX07fDnI1gbw2
oCtmu2bssOj1IzqCXpy9wTGFZgjRJdXtfaAXXuQC8qo31/PwI10f+VTLKv14DpTdUoIiIT43aoNK
x4ncL37rMrNUtitg8E9sSssuVMlb+th0+TRSwp+Jutg2/qTpJChYrqmZxYyDyw6bwQMak7w4Koft
0vTLwvd1bm7+dnWAfUxLs9UrZv1tNzl5xPsO0nmx1St4UDN3YThCE7TFlMn/hpxKrQXBx5KPhcP1
WqI7YdbhYyH/U+8hn7E/G3fOkfP6YgqquWpp4q6Vbw3Z69ScMu5pPD9Ld60aEfKV28Lv4lk5rYGB
0BZWU3J8iP/9zELfD9NnMcOuFYJyAH+OBVF9Z8WHGFHYTVm/DfpB2T4/K/ROPJnO+nGKUFa/4Z3j
eHyNWh7ub1rWqzT98lHp1YDunpk1rdQrqm1UuDX0bQ7uJ3HbRp++U7unfE1iQjaGVbDWJHSTRcij
la+q5Zdi0OX7HkLKcLg88YKL5KZEQ3jTEiHJ0Tup0j8FONDKotMKEMCNg8agyXt+5p4XopbWvQ/V
cEbiffWsxK5/SqXKQwrWTf5Hns73jVJSeJYVAAJtEteC7CwcuUonn0IEjabXiZATgC6qq+j0By+r
qCI1ods7VnWvtqEfFtJV2YPq/DsxNePCKywp+/qsM4mlt1uJkLklMymQbLqoqMb8PvQ7LsHXghYc
ZG9XDcjeymx+XS8u1m/UDWJyW459VunOZZO7e/HQTviJw1DDBGXK8viHjhv0H406X2fKnLIBLmd0
dYFB3btNDtVWr2FqdB9I0dO50YK6RfW/IBllDQ+E+KEMgTvoZuTjEeX+x2fiRGS1CrrElkoSSHW6
yJU+eGPAj/0sg47lIjWoNEcOO4ms11uOWJFLy2aaFJophtw9/OZ1A2Ueqc5GaY5YUkjaoXmD/0vc
YY8hcrcbrqp9u3Cmk2JjANsZiy7/MAwwjB1qfSXk0KAuz398mi/mIQqtHDKYKjJ4YNvDxWXodjeA
Eq2eyrnWwU6/TydTdVnL1yhe7DY80pBjjRsybhtN2AI3sthJjqABmj3iXx68lCT7GwG4Ux4bDYTO
D94tIpD/w5vqAKetxlX1MjanblddCM4XsSx0UP+1q5yvOl7kdhWuk2yLqkwKyIyIa125AKbCiwBb
ZnjhHOfIp5xHv+s2OdCEfQTP0Xoc2ch8xYYHGiucwKpcw8h4v6B6Sh3Ims/kSoBJk4hoKkYiiTv3
wG/vnTkSZN8KnomrWckWvp67pxn+pHk169bZXNoPIj1CY/UMlkV0Qi8TZ4kPMvj9ZHcDvCLQi5YW
idnbIrMoiYUD0teNezaXVjPZWHDoGsrax+PpmjfYylCn3mBqROadz5FEKO685fPKJZd9V0pvpFt0
S+8CFMVhZugE286ecw4ZQSzPyt8KX8aknoHjWEb8Grz4EW6tFvMLs/VpVaP0LZoqQV4BJKIcFpbD
x+gR6LBVscQWB1paadpEhYsQedPJCnqlEdqUFhGToi5yhndyjvLLmf/xM0SvaomABJotSkGqtX5j
w7lDfCsKIVaj266QAjkLSi+KTLq1CCDlr7GDN7T7Ewd9fEKI5xS90vqTISwAAyeFrAmo43UBDF5d
hIjViLf+ug1C0LiFgOGa/Jmsm/ZyJNYZq3pWjqFUU7F6gr211KYrCVXP4c+Y7yyNKSCEUV8JCRQw
FaZ8NVE6bVwAvLdquArqNnaBhP7y5LDmpJHSe1QHJL1ABp/3xT0eRzfxBqntqXEsvtcsANwIgUUS
s56kT2lYWmqtugS+nTvRwUvDP7drTwRrTz8Fj9uMp/Zq6+sjAJ702/vDBXupTDF47mExJLToDxn0
G8fsSh2ZXihj8h3yzQI7Rxbw14R8JbV2cC1hcKzvtaO6QZ2VK1tgQGtdK8AWp0PHLhnCNAejD1Gv
z0pMrs55qvFvXD9pCNPw1K2Q0Yx8jLMWJvZLzWKbqeb7XU4pG7iTf0HzwVfOXjM2l65C+nVALsI0
7PLkJ6KLtz2kM9ovWBPrxddrPHyQPPMHip29cQxnIKWWZ2w0GE9qyaxNreXzreTrltggkay7X2we
1txGk5jhlLlk3NtYHfXKOb6gWGnmBUZ/nFtpglkpHCPRKkNSbymX9YafB4kmiDRNyX1fJp7ji4ON
uxZUxk+B39WKD50wrreA13r/grkKp7jB/e3Z+lpeIlnEQlh9HQPAxrHIznr06CZ5eN/B/i00pj1V
OT1ZSZGR8AgIh0AEnzVrWdi5h1j4jJC+RGgymSdBREonIjZ3s18RvRtdD+WeJdGspt1eRs1bS0qO
lTvNILNFty/rCIPnEG7PzX25ricJdEtTM/e+0jfwzVVh8eycTBlijVI8C3aKxOAUgejw8DVn6dgU
iqvzbIMExQmbASZT564H8z6aWoSzVCcV51Xwfb0bgy2dXAwzTe5TUVd3VlnBgR7EBCTed/RrDQyu
iuR8nUmm49Ww5dRpD/YI1Oy5zisDmlompdeKhD/IY0qxrVIBwQHormIfxWF8Qrtmxr+mTCXXNcPu
htyYYodqU6C0lql0UFkzZoznmB9CdLzhsKPb0uy90dMN8AAXAZmuEhzf38y6QjYxTuZ8XR+Uw/6w
sOfCS0+/bdgn6fyYpULVxL1svjNgZB6QujtbniA/oFqUQ+eyCwCMop9duJNPfsZ4DmRxrZLcF1We
ZZ5IWGh0Ync1dg0FQR5g1t2Jss2pj3d0NXIULrtLt2cKtEmtArGqMEHx8ba2vQQpph85RUCfvjav
spYwljm/sI7VXeXcRMKOogzAlYp8Ah//MnZcQd8d83K8Hims3TxNbEXQRic/xswZKYVENp5hc2Pe
VUlWCJel7mkVySt1YBWV9gqeq/ORgGnao42xEKViRy/pJYW2PHfl4J1Q0T+ZIkqHHfbodCU/LG6J
uUsebhXma8ko+cPhdP2Y8ceJie+RsI6/+nys08NAmxGTPr0kKUZiu9Rt2ncbNKb/JTePiktMoe0o
YHccxtcjQtwsyW9QknpLkJPRstZ+TxrdKH3nJkMwFnjY7/5ucKVmISfN3L1MvV5Ja/QCnH7SOZm3
Swq4SSXkm0ksbHyobqGkMiwYBHuUk6RL1ddPDX50rhnh/F+jU5E/JXc+onp2knla79smLKUcqNSI
aqxzbfnlc1wXIV8+l+Jsul8Q5UVoqoJF6OoRwzhPdNweyLKMKPqFlMogkTQX+RZIFZiOajJ2LZIO
7oWTSnPm0nIU2huZwjfpQtqh1vNks3zGMtDajKYAtlAgFg9iPxFDoJAhgzd2moKjI3Kc4CDmgIZJ
CJdb/bEGB2Uv5XshLU8i6HVByNz7VO10TnPV/MjuFDLHDKRR2Uy9WVlVx8AC8uux3g9EyhSdLpIz
j+PouPWZETKH7fbjgsYBzcozzDhkl4zFOv3SAZUMk7u0bCb+tOqr2T3EDf7bdNmGmKtrripMCXaw
IZ0/UblEOanEg7kV3gfPOi/BZm+IE6AG9DLREmfJtt/Vz3n3mcg6Y5x/UxxOOUZRfxfzdFL4Lqfj
yqpDKv4j9CW6dj/0Rt2fMPms5OtVOObcZ/5pOkAGjFjqL3qGDL8GKY89jwoe7QRXQj9XD1fHF4Gd
13V69SvYywZGv16Hntsp7ZHVzeKLtTN0Nyf4Lt+Cve0S6M6I9k5H0KZ5P1ZpT8394rpOEauwltmg
ABhSyUYAmhHrMA7jkPKGZcy+dVxuwajdP3eRVxIAl7T7ZFJPY6CQVGXigWeV+LqeQct+yo4UO3yF
5G0TH/Tjq0Au1YPA5RY4LYwPga/22WgnENfT/HkD9sai8PWsfq4fmNBceFY/srco++KBwegcD0z1
I8aJmw5Ucc5hytqL1b4Fq7Lm8lFxGOMIa/KqjHkbP7Me/fK7T/0oa0UkuQQ/Hjbdr4NaGTO/SVEp
4F229vlOzyJGU/wqT6NbsZv5M+3RGCDzkGKd8r2VpZAGCiduEa7lHkefM5v5YFqSMmzVE/NKH0wY
5Gkv8K44HU+9rVG9KaHomfdotuXz2TnzbDJ4n+OTIEF8pZ8zhn1e3s5hTOA4+NCUXQ3ljXo3cZp7
abBwtRyEgNlcpDGyA7lBxEqfO44E4U/GGxAmCVjgNl7HfiGIbNnz1cVSRUmMlWJK959LQxPludW1
b+5OZctFawkd9uYCjVWni0R4Rs3D6jfEKBbIekg0weXWg/bj7NOH/sByjB1864CIBXUzDkKD9KDG
Scc/HwY4PAJvI1sbldXwasl+hYN8LZUunbASnj3JpoaBrDy72L5hu87vX/7M/phbBUUIjJCS26x7
R/uJFuCMHQaNCQRKutPkdUVxQCl0wj7T9Wr3uwt+pdsmS/AeAeCgJ+YZLM4cl4OJaHinC9Jqe8ED
OILmspyM9UAuMh/IyFl+6HHyBo3wgCT0z84sFzuCa54KPk2Z4NfvE0TSkylCK5eDLZCx0tgqPwAz
pooxvhLlJiQK76aDBubgBIKJCqL5gjgeQau3tmfH8HRMIm+Jt/Jqumj6Hz+pS6mDR3Oa+bo5ifSH
Pv7hsR6uPcKisfpwGLkRjvVOvp0h9FfMfxDcQIAyzBOSWrqxAr9qwI1xai6bZDbUtjwXpzne8JtU
JhT3UZ5IwOPXciJEmkmshVHN0NfOWCSipTIHXy0vwHvkhn8ZOxDexHYuVnMEsmTrHaDOP1CMWWlR
rg+o8sQ0pAwhkmZh0sHrN1yLeLxUMoMSE6bCLPyKmMHaxvb9QwaDoMUsAR9kneX+NARD7lbGt1cC
dFvsceDZ8l7JgbqTX5g631XyKTJwzj/SgqNPVxFGM66DbJ4wczpj9WekPibTRT6vsgDphUW3VDWj
HBh+oL6DLeEBy+ppjrH/pY1U8VtULzw2Budd3k6zUmaaXD+NGnUUBQ0BA9xG8kPEC3UzG5/xhGtQ
Y259MZlfYUi3X41e6pgMknTa4+AkpljfdLv5QW48PQvrjAuwAzookNRq+eclDk2J26TAGDKXeoZy
WpczWqXduk1dW/O8lMEum0xvkvL5VX3rraiH/Vv/eUk3Zt1qIK7hhLJKIHQX5VrwjK9P01g008/y
k6fSYGenaMCeLIntgmVS1ZbNBRISEGSqTsSwikIoncTGgTvEHWLKd94p+thLAFHnwSOVZ/pvIn5Y
K9WhJifIRwgkgZQGlIM5gQ1S632rzq7Fj+wEEICYalbQrDzJ/O6IZ8NHUjR2JWvC0nMu0TfOfgYC
524MGkPJ5AD50gHdK2C5oLSe15CEsgZEkS3piqmvjcKd0OIgUKA3xB8vW8FacCCZjPvWEa+vO3Ov
oa3juMc5wmOdU/igq6jr9QEBXUSjmAR9lZuwC/vwVM7EseRa53A8K+RnF0D043ObcigNkKB3MoPY
0oFgkGkaqfTzB/2WH4DwdD5ci7B8DQxEgvxigF4F1mWPPur5J+fiW46VcM2V32X/cX9bcbsMSwV2
4ob2aEEDsGgADvcWbwlxjmJMdt6FZ1+QY/QB0Lw5hzdK4LbT6vOC5ShxdBV6TVQO8LRjdc8p0Pam
TbaXHc4DgwxjOvF9m+g3CkDHkpB4AtZMBpqhff5SyAdHquKqOG/PlFvMgfvU8Eb2oVUHRFIpEjjM
D5fWoFihEtK64dsB5BTpxarxMVOVAaYwM1xHTihR16BJgDZsWq6igBPwNGGEqA5TAAml2tDDQzeL
SKLiUosZ0RuiU/mQGDQOZ3jekU44tcVcMeOTZWAACmOEH8iRvez1urI0l/zDXhKkISIWuZCdvLFs
5ftz8jSi+3RB1lI7Ak7XuCbLhzwOBS2tEnuV3Kev+gClgvhb18XwZMbbBi59klOjEIsocJtoY6+T
VCVYw0m/D1UThriiLegYzv1yVvazYB/SL883B+l25nq+JNgCvIO+qYCF4IZr0xrmXxTCBAigvWkr
0EkkiBFrfUrDyBW105U0t0GgJKiD1DrEhtPSLc7cwXRrvoF2oBZxUXEjTnLy7pH9R+PqVa6Q2VWh
0wlygZ6Jcfgs+iR5/e2ePpLUwlxyQb3Fw6ktghQClYeDZhn+Y5PgBgc38yzDLcRyK1dCa2seXDM5
yGwP7Ymvsg93AGIpCrENYs6g63FWZmz7tdnaMGhD7eISJuO2jYsz3n+y3uWuvyHDBNP1PyUBJhRV
INvDmkv3owi2mWVemeCkADQ72KlWeugTNJwWqQkx0AgwplKsKpj/TLqpa/f9HJJri/TBPlPbsrKN
s/HcfgP+QkD0qFLRSHkHbjJPQldmo38WGSwHwl0P4NvRZu1RjxTcDf7hKr7dE1dZUWpKKs+VpiJA
LpIIfwDIQwnVka5Wtbi+g/sIMiMW7owcmU9uaz3sI9Dijc4d7DrEC598qbt+H1xrbmmVZI25nzTK
PxY3nu6Bjhl67xghPXCs8c8uQrzI60Uu46+99hycHrmB3jKq54+Wnw4ZuA5WcLADbz+KpOW4aHd+
ns+gYQXf08aKh7DSeqsRwR+YqjZQ5jfkOv1d3zPMfnL/GvMWNc8Mpc0BRiNHZ465gxsj5FsrtCnv
3mtRiX2hcCks01Uym+PHjUAGfmwMWEp9vCmq4TJdAQEqsOB2/DVuD6NcS7iDHkg3yf2oxgiPafmw
tNxKNr70f7XHj7jgVgcFjjmY8dSZPwVWKcYTwk0LRwErvrBDQLtI3cZ6ykOVr8tELz+adGKsFnR1
8Wz1rD0nvbeUIoljoaziEkfUyU7jDQnxXHus3qx3BLhuVHgFyIzUSChC9ln7FbdndOpzr7p7FRYV
ggxlxrzUyHiz/9fvU5wOKd+1KfY+1i8QvV8A4zocEwu7JCHpreGIMwY8gRWQOkhTOvAKZeuMZi3l
VdOy1EhSZiHt2x6jy0JaBLrp6HJ2jexje3SFsfDZ3S0oAnlEQZ5+/Y5oxHxl69loG11mihIjH31j
TywIufXOwMhRvknD/3CJBos2fZrbT3uj4XEvKH3pKyjzQpxyFVs2n56qQpAX/fmIc5gJYJw/eh7y
uugvLo1uGh0I7+sK2cmISJ9/Sce5Und54gD2Sk6HUKB3TA0tfKYKiNCloQ1mSBq8QoIN72bbfqbM
JKxIY8T/4Q7Gp+3+8xuGBIjgaDjwV2mjxeRJSz16HMyXO1QCIbmnWVb4sVyHGR371ZlPqSaShIE9
lgIEYxH25JNlJLC9tLJqQSQ4d3mJnrhg/HeXZXPykyzLVXWu+q+yLROO1aUVjrlxxvzX/Rxp0T1v
2CjnKoTpUmgJg7SYwiUdkd6SBfP1M5XKb5z/vWQxFzPTMZ8iNCc4ewDMJF9Y2Xp2LklfXcjoYXKy
WrMZ8enLTdogDnQGMxrewK94AUep/It6MPvIwDV287Q93/pQ2mvaFqccv5qgov+ve7hiKeKNUVlh
I/EMuysjNzSroPWUoBj1gmbGNBtmColGOCFkTnOrPflukVXOKKHww3enFKAdpLNcNrlw4W02xbVn
LuhI1IeiLCbxi089FbDM6TPUNObYBX6yyD7KKivwVIiyUa/8C76/02qZpk2nxyVCuLOZ+VWgpheS
F+I5GV5e8HgzM0uW3nzg7XbceRVG+nYDBcnUpDBiIfsRYqXO/BxNbmO1Gob5mB1tN5ATh+U0R+/I
2Ea86E/fVDQhlkNp//yR7YswG8i9aKRV9Ejq6GGP2dCMDI1J3/4mXPwRJprYJtDhlRAGGwhniQCA
X2rtyB7thL6HyMOxR5fqq50aVcJrV0dnU5yKA8V4/dVr6/42Ol9YZQI0DmRSJcqG2SZtsZLe7lps
K0ia5zb4CWXdi6nmONBYorMwSa9cQm4jQ5wZnAW444wszpX1wyIcp0H9xjCQM5h2qTSZB5Y6trjp
v7VDXf1YmveYOcn7XJbhdLtppM/JQ6L5QtFWD7lwHsbE3knEFlY8Ca6g3uPREXAgfg74gWS4bzHm
WEWuTxer01UXJGYDV9s1sXwkg60ndzMMPxsBWT1ccOEvXFJZsP81qyGqNXKfnM49hvhhRlDVlm+Y
SRBKB1Rww3HYrw==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity fpAdd is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  data_a :  in std_logic_vector(31 downto 0);
  data_b :  in std_logic_vector(31 downto 0);
  result :  out std_logic_vector(31 downto 0));
end fpAdd;
architecture beh of fpAdd is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \(FP_Add_Sub)/(fpAdd)\
port(
  clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  rstn: in std_logic;
  data_a : in std_logic_vector(31 downto 0);
  data_b : in std_logic_vector(31 downto 0);
  result : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
FP_Add_Sub_inst: \(FP_Add_Sub)/(fpAdd)\
port map(
  clk => clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  rstn => rstn,
  data_a(31 downto 0) => data_a(31 downto 0),
  data_b(31 downto 0) => data_b(31 downto 0),
  result(31 downto 0) => result(31 downto 0));
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Wed Feb 14 08:44:55 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/Integer_Division/data/integer_division_wrap.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/Integer_Division/data/integer_division.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
fbDV08QTAHfrkuad3fu8YHTxW95tUMQhdVQWg7Lk0bWz+eV0+FQgs7kDCzm3DECMTpUNsYE+VUOt
KQVl2yBwsMJxOF+NUMeLUm4sFB8XPsGxS0eMyQEAH6SWOnBuM7h8xbIfy/qmB9X1ppQB1gui1Jn7
P1NFizLNhriDYueiXuZvwo2MacmOMMqLDhJLVoMvLJ4+2RDIrJpob/81st6gmlKB1fWsTyTE7XvT
KLAx8P8TqMzbKnJKl2yTpY4VvbqpK6qxJHzXvuQEyoEuznlKbrMmGtd4Ezh5ssA6kfbatKO7YrVv
ZQ0WWviJR9EB0H63iruh5KqLwg7tSNgi/jfueA==

`protect encoding=(enctype="base64", line_length=76, bytes=472160)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
vcuxu5xsWWzSMBlEQEX6ea3OZeWqWtMsKj+5+CrdkCjbDtOWHAchxke1qkowlSJxUZl+Pvus2ql3
SLsrUWZ5H7dTF49wKVaB/gktSUHsM73dZZZ/L/ZhzS7mRWvPWMaA8tZDCWZIAL5i1aMlc0vdjJD7
Nah1vogJSdaNNgqH7hdKYzt7n1VWw9NVq3mY/wq50kPQCZ04KoIj5XiItMr/sVoFX9U1XMnJlTdA
c174Y/FctNx45lKlghXIPGhDDGzqHKPlxyjyqswykxEhxmk3njZTVln/vz6p1TvahfAvxC2bT2rh
Hy6DRmC5DcaGCnV2v9Z1e9j3p2gCYdzzl2lJIhmRYobfIGqzxp1z/loFkIybmrxbsAVx9+L+OkNg
sUT9Q3Cj5q7naD0Jv9hSuYkBev4DBe/1jdPfwUq2uVpwsRDOXZqIph1PIDrWvYci/fTBtrcwVe5n
6fIl5lre1mrxzhzxGD1ClLLutznpx+nytQwiUV6C8wcc0G6ML1pretSREYBCae4Wg/UmRj7iURqV
X2mHmhTBK0y6nkqut4OWRX3VlrMe5LqIXmCYoWiYFU/YZN+FZXOxzxV5oA2c/Y8ZLfB55/dPmkGq
WLgfyZpRehlCnwRbpsHFOFJ6VwRfz0474dZt9RsUlnPvvni4eIm1mLmk+qci4MIiXCnCbcVxbYqg
fEG/EmofkCFPWAJHMtFxzddSkAmkR4Xyw/3EEVfXJqNRJpE2xps1sbfjBXnLoDrFaPdcJ64lLjhh
SXo27+M5Sk/gKE9G8zsEPv7SYJNjvm2JNhuD4zDwPQFhkoN9zPWXUxVZQ7jNNBkrSaQyhvhW9VoT
GACi88IU41YCSF7xzqfo4qMaBflO1OXg7co9Tyfg3Q9OsTgM3aY1adbg2d07hJA8sfXBICQn2jJZ
uQeDeT8gbw3iTemjTG6LE9K0tM9/If1j2gm1M2lKl4lPpvCjaDy67r16lflzE7KYfFCEL3cJhnr6
AUOXwT8RwG9vA4/9CYiIKuqhAKeDRRund4fq2J0wHCR1tLh+8L/xrYe0LvLBaiEu6CkY9Iq/gnwD
KWJGcTCcYkzEdp999ER/fytOjbBrPvTOpqWvVqxF7hMR6R0agJH3YBqzr/JJsLpQuNrp8VXigDMF
free5shKVh5QgIO0PIN7dJnGIcOEMFUYMaX5pQZl2fBY/OiUwxIH5q5l9jfwkxlSifEvzXGnJiCT
WOiB70rn2VGfJe0KzFwF9PtQEww5oVfxEtxxP3BJkGmxmhO8PRUX+pKNW+dC6rvNHBFGiidhhZ53
TIectQL3FL9SuhqHB5uXFQ6ZEEqtUw09g54h6VMAY2bgEgj7YiZsvYGJA2BUlOWchzBdA9ZRsfSJ
VW3hiK7Loc80sZNvniZcOhsUcAi4/sui2YfcGRed8okAHMl5h/DqhloUKP1bUJ9SkUJmdzx/eefX
y2xEdgR66YfLyRKLZt3VjXrt0iuPTJryu3LL51pQRLxUlj4aIer50j018eaMyUfaX1j/7x6W27bB
ZrcB3B94/plj4niDPfvOp6nLCia1Vh4Dyc1ySqnb0rwuTr/MPwZMfnXnAsx8VVzLkA+sgjrqYXgl
WHctyrYP60WUycjOGeHZKBAdv0O6JNyAgLjTNmnt4Ov1c2BhWW3Lt+6ruCwC+4V/fos2VlWervxp
KC0PuybUp90RNokFHOiheVkzVmbXPbVo3sSmNho2O6Z2lWhZiQ04cF0muXSsSkKi/XwSbvpV7FOI
RQ/i9c/PfiMXNMQlPV8R0319K7HH1uppE97WUfkL5VfV4cR71faBYPGTOBwxAvSGTamhSJXaVosS
ZQeQag/HcPkicyXUs96E0FaHLBovdiLxD3niNxtPwTD8Se2mjNbZ8Yt1K+HRWS95s2rW0gjao5Lt
x1WDQQmR5YRUJqpwaJUQLB+sm3Lxneu1k/GFWX4Nq+lMpreoy1GhE6Oz/4bgpt+lNriy3RkEq+wo
tJ3MA1WzCoTRBHslZDv8dQjItBnmo+GEROjJ//4t3iJ+XruNzgK4qot8CPVsUuavnSboF3kJhLBj
3jxNwivs7gykREOt1gO/uouGdKDaSAIMhbJBjvuWNPxQC39M2tQN8DtzZ4Yl+lj78K0XBWBlea+V
1SdSgD9FqaJuKYZHhhWnwOscfHHpVDCHlEDoCKDLachqPMW14RWhg26IyIuIULL66cr2yicAo+j0
GtlpA/EHBO662zkvdD3xxq3ndAv+AslIbtREtUdW/76mOwsx6hXRjVrS5I44YgaCXBM15zq0L44/
abEGcnh86hPYNL9yb9fVc8SxfIpf5rSrb3SvaFpOROPqbrpYc3Ohqe1JnIeUSQUI2ZIXsjC4sCXr
XseZmvMPGUZstGo+7qFJ9A8iBCIX/gjD4VubxsNZgegyISHRUBqhGuieJ7E3oBowZyD8oH86wNT9
PMewsFkbVDKRW9/xQg4Ykql4m+Qy0QgMFXbfmLwAgalj0cqafS6GXXzqogt589R4yQcPpRGVmQao
TfApwuwFCjbci5NJhg1TaOEixRau4aGynlmpVFIEcnqw538yruRHs1TnPqfq/oZ1oYvo7omAWrOZ
0MitwqHuxLGt+ooJ7YhvQGOv19ML0zlMQuAJOhUqJDws4skU+Osa1WJemeDn5udjJCHMO4rk9iDm
Cu1Ivrs5l1omlSuru3yLPIYxa8ti8Erq2ueE7P0MWWJuKxXXwVCJHHNR+vNOrgKI616e9vzhfRcl
wvbQpXI2IZs+KOTwYG9eEKzXNt975ueovpLlU9uVIkmcYDSasaVhk0sIqKAAKODQnLel2OX21RL/
xwO2pI+RJ5YYrawDOhE0eiPUYK54z5lhC42zm7nGDH1ZQGDKljQEZAotR9urO+fXeg1n+NkZd3Nn
a5yzTC7yQNjXnNnEuLK7gRG8vCnc6QvvDHkc3tKQVULR3Z1xN0Gh9rpifQBVp4xwm0cwhRugeBOX
oA+CpKgYrX99axseQp0qfAsT+YOsVrrYtnfYUNMRu1vW7RNqOq8phsNpnZHS2RUWaNUUax59Ma0z
i6D6m8rzFoQsIEFPG+s+byLJqZBpVRQCf2qM3Es7SdnBmFLwWDQ4NLLopl6Oofl7RtbjDXIKcLM5
uiUgRh47B+6oTXDFJh8zmw6vSSLla5RABd1qjpNNU52Wii8msx2d3lLt+9A2e2A9pPh7w8SjE2Hn
PEVxboTZY72aBfdIcsfk6xwZ+q6eQd1nkVI8wGoHc2brdkRYupGCjPSWQyyXBZcy+7JkIM0bz6aL
IU+NvKEPYJyPPG9ttG/0tKkDs4m7SuMmGFcWb4l/pbUaSsCXZGNbCVtnEjLzJ+HVrVpYeBNsu3h5
nli2tjohjKZIRxMIXn9Q4FP4RLc7FMJ5lXJEmB29WrKrzFknbu9Hh7QfL/XJLUGBIbeN2g9mhY5o
zDLu2Dv7E/9WtR5jphLj0CRYHLRI2vtgG3TiL1DIvSpXdZuIRWuxGSQejw4CdhddPM0K3JC5byH4
jpqEA2DpxstUJsT2bzQ+olg+k4jiAAkQ28rMur03gwG/cijkC9VNU+pybhR6HjnxeCWm0hcO2FsX
PThqylIJpWXVoPjV90O4DbDUGWz9J4cbshJvYjylsa3Fvn930v6mW1mM6nPEKz6DmUlS0uAvgHN2
kEALuDmxrTY56qSail2IJeIdmxOhkzMedkSR0m+tTYmCo3D+Uj3eeTyksDkKc9z1yDDcoEYr7EC0
KSXtqtNJILOUyphS8Hz68tDppmtVvfEyTMXSBSF81pB0QrhRSpgmvXJKp10h5BMIW4atkHcAELdF
YJp/+dJWOaQjgvwWEKdsmIXxvszyd0SGVa3/a97+VR6Zj1tNe9iN/sWc8SHR6L0Bn/Dd8JADLEwG
Bq8YvN0ZOpBfmOmAKNBhcEXuQpv/7LP5T3pflSmdt0lNSghd9dNkYFgnHhLcfUhb69NSHtGGsrzJ
JO4q7XVzAsTTnLGN+3WiuKkqbzle4Qmw3nk+L2tdCnROvlFWsCKMfn+1lL1a9cinzLlPoB8i2BKp
VMlDmlOiIz8p+xbwIPGh+BBt8wtB3REgw5BNfvdE/ODPwxvx0N6BuZSCdRd1aUd84v2oub4WD17Y
RwyCPN3CXkxFq2j6y9eLFqs9zMhlnU6v8Ps2+zT7p1LYBIv2XYMon0a3+Q16D4rPlTaokOlKV++h
GhKNdXqrZE1cDAFscrIw9QbkAlZi5W0PE2ayhHL7TFa5CeASjQscAR40exvxpcCgbffwSVvH0tw+
u5h7DCT0mqiBSsTt2ixHme0XJiyg8uqyIkH4LG/M39m5CCkCs1Vh27Z/PFTVYVs0j6OU62ar1K8a
iqUUpIvEklC/d7e7Cc7hiWuR0LlFjj/nZz5MhC6sKggZOrABnldUWLh7vngukfLnEzNIc4kyvGWd
pauE8hBCgfzr3Zps7kPcK9foTmBP9xt3K2Ftk9+AUdQDUcIhi2UYj5G91ZqfgFLnxyjTb3o1BQdu
kV474B5BPmO1UwpJYJmsWEopGg2D1K21q27E/doMEBKtJCmGfniCEFDHEiFys073SyBFQYm8VkY9
szTRpZpN4l69kfXS9O9MMIoZAmL0KLH0BCCj2/bYRTDQ462CQTopYzMk5uYIU9WGFVILDOr1/2lc
K1uX5IvnyGz1YKs12bJOo8ior/5svSP+TtHgxkchVnTHnSDdNqdfdz1f935hD1i1eOGkOsut4LUd
Iuap4JwhmnM7E3K+USdBvyKPJWaY0ETIlKYu1+PUfRL2PgcyrOA+M6Rn43dQ7c2dI7+CjCCHVCXa
DPzaMH5VUTHfADQ8abdppfoq/zMgNZl+LEzgywFu0CMqsEzHAOin+UTEd5EpJgI5CHkIBvZEGgON
/Anak0CPUk3IlNTsDzrQNdw6YAkP60qAwPjeaNIrrqplzz8WplI1f1l9j0tjf7TlnIJbZC5FaCgf
iLt4nvzvlx0zG/WmMxisXUvy682ShnbAg3spQcQUvTZHTO7rmYN0xIWECKTaCrXOhtY0RgUPMiRf
7CBag98PsIfrJX4sEJXrSXD2xuGZpknLKdAHVZFM0CojVWIdLIm8RrT04RbHVFFHj9ui+xFE1ofT
F/dV4gL0ktjwP9cjZfP92IPhLAznseF8sVlH0f4sS4jwCMKRb+TEhIuVEBgmI9+LrSSE061jajj0
HBZT0Fg/YKrQ7khsWvdwyZiNdn46H5ihDxTrHzRUJTqEFBNBWk5Y/sGnTVyWuMGY3tKgHCmm6AZc
a619l8J6eYubU64vdshLSEtPl5HHNJHCR5lmLMGpyZ8k1zjTjIgw5HKNSo7E57vIsmmddHflO3Zg
FyqXddX6Po1j+yJ7fUIkOSuw9d8ryV680FQ+/l5ZjqB4dTHZVBy+g4YsxASKw9laY9cjtXliEuEr
UZCU8Tto09WFiEbIJ2bd7U/45jJ89hgdfkLU9VtI9njkF9TmSyFJZ4fNTfsG3rtayQ5U2O+S7fMd
01PNQ7Ok/bOeq8hUA5tbjRSEcfH38B+KRA2RCgMi24RybzGR0IBzn57dBM2kP4k0MLMvBScA31mG
VskVtp/lN5RPdzFQNVnHwwm5tTFRsQbFTtVh3uHdpgh57Dw8Km7yMTxMPMydVAsWs/y/x1GRM9HT
DtXQZPhs+wHR79mj/TYCy7OdIVfQ/YVWmtowtK9An90NqgFTkmqPIPiRRQJ7bKV6pvnSntP1vhxW
prN8OQUhOTO8VJcQCKWQZG++JoRzUZLt+addpKH4SrdOGItYJRbK9Sn+5vyGo7I0/8NL566dov3T
g/flsBVUx7TLwo5cbPD5ukFWESCswC+IZErEtzRVmBp0pznJS7UC+o5YiURJDXi7UIXfXaowUILB
75lwcEpL+TZ/4DGKlwzBOaasJuu3cuXpaqp8u+Bo8SJGtTTq1cPtxY/EtGlBPU85+z5rJ67qufEW
Rq+2HDDFSG7dkx6qGY/URX02TLDI8GwvBhL1bP2C71PRVE8ZCz49CC5Y0kNml4as8v1+kwi7ASPH
oKMJXxBVW2QHaqo9LTZNeKEN0QaNRey7hXff2vq8Kcx/gpznDqaoSSR9nqFUTPvr6jTgfgm3Lx0M
zLtCuhnwPDDijnqUGNq+K2Dy7cAaWXFIYbFZfGd1EsADgwTJ1wIigup/6v0foVr+GLMOtaMGYpGO
rxZ02uueXSBIga829QQA6+9Fna5+dXff7QRpfbU+D6MR6ZrAT8weuDmZGd/ki5pxPvxglPMJTI+k
OOxe0stqus1ZmxIIidYd446agFqJDKUBVBxDun/n9CusDwTlVtLNQUfDzLVlCiGQanItzxDj2WAO
z1tD4DSYfbYayOy9IdRLYnEeHu/i21Rz3FW324hcwrAbbDxdxbe7o2YzB68gsk8YKkkzDpIog31Y
gKor5elq59cUfeNbGTYO6g97ncHHak3e7XhDTYZwHnVgXlECR57x3a/235O5h+lc7V8flthH+txO
DqkWw/NYgKRcVotTJFD8S5qkHcVK83s7Hgkh40romu0dJVwhlS55IeavGA7g21cXhlITHpop3Iia
cWAPub6u4bVMWrzbeageE73G055oJJiOD+9Vlh+UVie+2h94/N0GsUFBv24V35Fxj3QE8iC6cVre
P1IV2Q3PA85QQabxhGIYTmf/dle+8HMuvvt45KhvcsT7oD6UfBxR6cStoEsJOUJzBSNIK5hye8T8
GhO0ApRHzeZIKi+giz8u6nYAQWP+M4rWMoxO4vDN/5s+4x+WQvRGzvvnVlYRkPpWOMvg3CAS7IR7
EkTXjgoL2SXd/RCXrCp4YKNti4p7mkL2cfQZlx/5+ZMOzC1ifDBIQkEantq4mZgqAvJC8hm3qT/F
3CEVFAh2Oql+NtPkAqvevrF8iOl8v+a1eAXh40K7Oul38EiAsB5cPrjudhAuorOHAAR4YW0Z605w
e+8daVMqbYwS631cKC2fKararl5m7jaBfo5oxiWoWGpYvJAM10uq9j53yngbqk8H3D/L6TJV9mX5
98mssOQGLWfvx2F0LRub9kS/w+D2U21YUt+oS0J/BBrKU6RArfv/GsDvbnC3AIU5jDevapDfS2mu
qzBg67nhl+hFZIiJmql++D2qam9yqv58iDQEV18BV/hYK0YBdz8bNmjmVATpvru/5ZzOZt9w68y+
V4edl3P7+cH7H8zqhsERoEoLbOeuxxf6zHYZ5ONjqodxIUkenL4opQx+RsmsEIjuN/yx/OhRl1gQ
rCv4UAhWctG1rXN8q/FKqn7jDFrpgwNA9deMVA/pZ8wPmtcu3hIEP/raibCadlpO96DQfve3rqP3
GzdNTH6vYMMqZxQ3diQMYlzFweyFuzYdTjgL1MvNU+H7NwBA1AJ/Q2t3LS0s/7m6byAkVnFOYWQN
cncLrF2bkSRHYzR9jJ3p3XPBjaShE715h+vYK1rz5VFo4UgP2JURT38zdpMVZgbv9sNOEF6ddKpV
xCQn3th5YxviEi6QOo/576FT7QqEAl7kpeO29BIiygepVRLORFwWD7ct4kKTahWnaB14olMzFKdB
zuRNDK2d26xxgycScyF+jARIipa8AxkebLqjk4Ni7ko+UxYix71icSy3pgokdnRMM7kp96rxt12z
DYLKpLcOME7p/NJTYca17+R2fFRzMh2zc/pl6Y09EQTjdm8M0E4ZCW939tvAe/fRL53SH68FwYwH
THJcKZ+95aYvU9EzdAMAbZAoGMtX9/79j53ciZZgSClgt72yoDOqYCg9+OPim/Bsk90X2dExjJc7
WQH6xUccsVyMGKS4Bfhj7mqa6nCbmvxUitcZQ3OWX0/yUG3Hyrd2lFW4CcDvjIMhx8y3lxAsCAZk
uycydMfrFRLQ3bj5qUHgK/y4qDVjfrrfcztKWpgJKdQx2rLY9ZgMf26d/oztRVVkaWDGrt3LfGtp
1bIywwcXjGfh+v4vD9wffbc7LMaig5TfGYJAut2nFKnf9/rGpNH0bp0JW4LhldzXVWJPhTDeIacY
ypUMT5YgkBDoYGbywDLADPAKFKA6aim4ipjq3bvjS8ffnkzwX3dBvQQwVgFyRLbJ0TNJ9yxSiW9G
TDyZUtcSgi1NN3lhxBdrykQCLFRro1PUcFXQFt9DrbPAwa8JQDb6dqfM7siZmlmN1NJXZObCx1RP
sTgnYICIazgyIBgBfXqiuUtv3nyO7/V7WJpqNLUeXEGo6/B2YdRtLBm19Y+YVjkZ8XR9qR8HiYvp
tUDjUd8f46taUxYG1DniHpinGtLUiIvLEn1U6jGyBN0Dpo4SxAFfG7rR6Lk+5mZSrVB5LOrz5fYg
YnkvRq6gFGc6nvza67rvslN5C+GKt3+ynH4EU9pEq36cI7oYe/kcygH1uWJnnxA6s1fJFcWLZ3zz
A1fYF5AMBSCzc61lDIGXimXCzHuS4RGPeXIMkAdpJyDbHS08ZSgx0q3Zfps9qcFv+n1OMfBg3X3v
BSwrzPKHLPRonRw0XcDtn/GOkbpYxPqyYcJL3S0lb0F3xeAVyEiD6qUbkMAm7SOAaXx0nhMtPD6B
T69t1VjqhWUethyZW1aI5WxQIBkDC5Gjrjk27UOZMljrCtOBE9JSiqAIp1aACPrkldRarvue7ZY5
SizDfZfNlTUz3+p1WrxfOtUExF4fAMay2QT055/54lvAbG+qJCr7shZhd8J2YC15Ap3G3zWmRFiI
eOSIn7fcr5i3qhjLsyc4LSghUKUoggCZbEE2xizI0UILMagSCOZo8UqWtkvgLKWvuoHKKNnkX1OF
PGObheL0Lg30zMltzWl2aQDyVTk33qjLp3dv7vVFTwMxtyvCFITK9wBF67ElDnI9LseKvn96Y/Bc
xv5IDoKlp6/ONeF2teUYDQHVJenzqyZ2eE1fs4BKps0LRB8NBzy35A6bjkdFGFdrRzPYW11vwffG
6pXQrkABwu2N3Ukjqk/bl70BEhbAXItGt69auuzTSLal6qPnxKPylF/USnwv4mnry2q/LX5sjDkX
2a5YXldGymlo5DG+PSU6xUwJi9WVd+C4iNt7PbaA2ksKHNxWS1kMjzfMcyCHRF5d1agINXODMHAp
TbBZC51uU8JY8zirBcpSos4kNVjJBn6jkv1iMYACkmcAvaNREV4JJOtO4I5/krivLO/Kn/X4Dtq6
mosNhqxtrJzUbBk2Drensd+utxZ2W/DExPqkd9yXtWS4p4KmArPF0vGATC5WPwZdkhYQVPcI8hWE
o1gUZV4EuEoj9MEjCOAh5BefiL3wksgLBqS6fPybiDuvStOf95i4qeSb1sSxE95isR6yOA7T5B30
ictsSAY51Le47JBuIpUdh33eKb4fbK4WxIWaOh9fiyDTLPCWv1Rjvpb8i54CrJRGRxR2Jx2EO8bW
Rf+9V2NM55sF6nGs1syPjvhaDqUIiF4f8EWExdsO6lN4kz5en9kjOVmYZbp4JR8aAIaGc7cK3ZMa
8QG8L/EN+2Nxir6wpccOLuu8Hso1dynVJo/VVzDjjzcqLfXjLPuf3YCoFtC5G38F+pxhhYyjLVbM
X+67vfwJrjHWcypKL4n0oTBzM3xPB5E4cOp/lQu0ch9bcTbMt8uSKVb9K+4vcMB4N5b8H76QgRYO
wtAkjSeXMY7/4oVFasOUImXrJjupR4iFdr/HxkCHmtVuentWl/5+WRsEVo4bJZVvfDKCgT2HA8j6
jmpcvrVxzfw8wLtq1ukSJVq/OID8GASAFBDdJSL4AWCSxq6dlcIKnFL2az9Rov7qJ80nZlvEwnjv
uAb0ZBV4IokKDo96ZjeD5AatnPCh01HYI8ZTd7b/VL9ekLCAzvN9wiFp2eXU0xVRaUQCjJoEzGQh
GGRV1GtLfla1CfTV4o7VCmiIF6WwkWDYAIojVziZQ9fWWic5OlZbpz4bfBfOM/VF0u1JiIhfKw8t
ZgociGo3i7Ua2l3vnWVDvQRWGbAzzCKYGQTk3Fx90LSImIIR7IIUAY81RbCVbDw2EkxQjopY7nFq
tXk1BOHRI4RyhmpVP66oGd8TSLNN++cIR20FTC4uMkELgR1nnMlVOK1xQCxzc+Ke2XpW4KtHNiQS
GAPNO/XLYlnL7OGb2BUdFoQ0QJFQEz+WlQK3s82LC9nJwOOQ3xx4hxrrreX7XklshUsbW1o3Hnjz
uYlK/3h07h1B0WIjs9MIcOoiTMTH5OA3Y5HMZLvIdq0CtVwOMIFPFbadII46Wm4jfE6YcJmjbv6T
c+RO8XuMlbSCmCYqcRHKfobAYSm3LduYKfIsJR6WbZ3qtA1/FINpW6UtUDD1dWsS3fAJQ74jUxUU
GwnyZOqJ9vH31q8jZj/54Rg0AopTKh/P3gQ/m1yUJ3wFID+UIhXF9kVBu3wamMtufRu0HDIdUu6B
sniJcopieeY3DCzr4d8qBl1r1GOJeNVTR9OSovJqcdi2qbwhTHL0wVC0uebfzZdiVoq9a53h5PCy
k2ekL2Fqb7uh2jXlyk7A/+kw6LEkFrwlq0IKujGx4gaXusX0YFIbK9dVSviVqn7omKMF0T2B8yVO
Xjh754CjQy60uMmu6V4/at0Kc+Uxj+H1znfk8BsGBUbYLRlClkn7htGWDpgsKFy6YLPYOnZgMpYX
aB69EygHLZDx1pV3l+zV2M+MxR7JBFELqj6bvL8c3do6oRs5hz7wpAXcHwE6cv4pTiTmM8LWtHN8
Eell8glGOtdmSObIOXBP5sKxGhJjPU2bqU+2x7bGmMcM3CkYeucGxYWlCWCvPc6+Qw5PPoP60bm+
XTfDl0Mw4l1xlMGlpgAL7+xE7kQlKo0xZ9baGg+brsCvi0DRK/4opy0pI+mvD9UBQL1Put7r7Mvk
ZKAEsZ9blg7CW49xISohe3GsZUGBtXPD3luudqgkrpLIgaqRC5haXGhFolVDvDp2FzcVOKhDhh9v
tOJT2CbaIEoX3BYj7bgIOST88s/9L10IBYVlNx+9/lgwsW/vqVkBFVQwJ0KnhxWn5oZdXt8L6blo
0MAx3qQF3aMR5OynAwgKaKFtewlq2qdwQj4TaAjPqVzw9ISNS9XAD/TLY9+tpSitaRTcxN/922zw
fJYtkllL1v1E551n5zCKphqeTIR3lyyauEgIRtbbP9M+1/yMnzUu94V5CaEejCCBUh5+MmuS4FuT
vtDJtJSeYwgGhIPOF4VOJWtLpA+yw2MmuLvzOJgl/aTn2Tyrfls746esQnzbE+pWBj25kbNwb7Wj
pgkKYtJ8XCuKN8xa1Nr16xkQ7SguaQVtnxR0gN2nzI644FOnbxkIvqQoPe2r7G2kJb+lKjEj7oF6
urqF5b5DYvJstSp3GBSPq5w6p2OsPks6U3TKHYrS1xMFcojer/0j6GM2/6KLG2EjwVADZU1xjXVs
4LdnDhZzoze4FSyWUn1g4qJJJRnwvWN86YGWF68Idz5k0Tcq9p09A2sWCfLrhrnvb3dp6we689o4
ZHkYQLmre1yUQfjaVaJe9n4W7SgWC37yzEzdiRu5jf1EqseFIdxCnDj8xTif+CEoypk0IdC0H6tJ
6kXOkqU/nrgNSaN+YpObDMLUiOG0KvvFlYwnAG4z6rR4VBjLhYDtmUz2OI+NX94y566BhD1YfDfd
gFSyP7/h9ONT2BKWMd+MVBO5mpUqXE5CfVUBMdPTtX5Nio3iXNJQOkhh8zhkq4MSJHeS5XnJYYM/
u6+GOKUF10eAGH7Mo0E+UaHaSwYsxLTTY/3NKyDFPAeojGXvXYqr0eQmBENFn3LwzvUuvImkMijk
CRWWqWJiyk4WQhxpi9FhUCn2Mw6n3wI6WHC7V6aE1OLL6TY9LdOknfYrQymRGl9xElYADlCuWsO7
EU6x/oLQdi6ManPtKcBFQ0Nzrlvb+7AGHpR7sqQwPJZmLCqcBfTd35UTX3Fx5eWTamT/t4ymL3Qu
Hc/jNcEioGCvg7g8CMij1jh+R45X04/RAPMJzq45QclKaKTUEWW5MtdxdCXIBJqLfH9fD1I8F82P
bnX6WzebygnWikkQmOwHxe7JSf28i9JdwNI83l/aa4uL/kwcmZCBn9Ciq0XL9zvNgNNPJlP9NlHl
D5i/QM/XL9zIDD+wdzAr+Se6PyCWlVnZE7LKsPJsMMtQZib45KFHVE4+6nwdY4lKIDjUFZZBsMjr
QKEMPwXuBK7Kc4h8wi+IUKcoRBaHmIi5HW9iuaOjdhmU4F9IDyNOonlUJE8zT8T9hhXrIRDQO46H
CBLorN2jumoBuLKcDnVAJgvI8akUJyZsJ9JJALa1rfv1gIbfaqVTXzB4J9Eka+OIJiTRtRD1RUbU
i7FzEhQFT3/37FPp/Hf8XBuXMC3JTgtsbzP0U2n5ylqjUeOeUF1f/kKOKxz54uClyCMAJFR6exuj
e8Xa+Dsu1UGqUS66gQ+d/dvlry8RFgKDwuEtMDiCEZPvnk8IpwprHZ5K30MVDpy3QoOfSiFE0Ngb
ELjTAjIJO78GuXIfkkJb9Hae+MeSOAUS+drtXqW6jRv6Q0ws4xnk3kOA/L00O8cEZALL81GFAcQd
ntwoAbJpzCUNKr+2Tl8DD1ClCp3kHFo4JrRTYYlJdfHT2nKmETZuJFHZ2XQn273F1JbfZ7RmDFgF
zrcEsNv+nAo9FuWwYFVHSMkUcinFb3UCZCllrLB6oG7w9J8VEqOldEG6ysc0I6EcXfy+J0g4ekUv
vzM8cygYb8Z9ooemGkTyhQlxAFWuqFmqLKIf7RHeWg7AGRODtulH69+rgoICQ9+QWjb2dFdVLYVn
D/cU/DXUZry9eE/VA5xTEr2bkYATbxIqwim90P/87K/L2eRsZqeR2Mu2YlTNXjqp4Nd2gy896ZN9
sUcARIDQ/IFvTWedve72xBVjTv5wQmz8/ACeye1Cy7fuGNhuhEosWM0lm1fhSExYNH93Tp5qHnfe
oGRcKzkLdJtN5uzdP8/gcoUTmpMaGlV7loP+b4HpODEQcfdDmsruCv6UkDXRZ+PA140tFDMcGHPA
9wuhAQDFIZkq6jAFzRQ5+MSVlXqbZlCkjr4JiCJy8GdXK60Pj3urkqdK+xejFL/hR7ZrzO2in82E
9nausFTdD5jQGQ3Jcw7ZduzmyCGJQmS6hDm1MEp3MHMIMiI13F4wrZKfOp/ZJT7AnOlGw6tE1OiN
US6vGQteIHGBG948xAlsgLO+5EZHUxR5eyhrdm8MYvUKtcz1Khb0/3Rkpb1Ezte3JQCupmZpT/1y
lttZZGe+FqTFcxf+sRT1DwntbdiOpSA9j/54qi1wYd09vi1MreKgfVhUfc//o6rOiQSfZqPdRuq/
T7um0A+zZpGrZAmbhRex2It3iNcf0KFkqTE2d+aR4SmMijjwSuIeuvM2jzSsnwS/upwSN+eWOwSg
+duf3kh6jK/rcJfPwV+8DJnMs9zI1+heaLaJPzMu1XtW6DXrYMWKizRjjWRmYVBoCM1p9pyFjske
uFWm15h0/Avhux1TDjlXRejbHK2lRIqpduyRIpCw7DXa9xhpypojpumlg4HVNAsfOFAk3PrimukQ
pDx9/Y/9qiCzzmjcYiAYE7UylnBcACIe04BVnSRB5WSGvIBtnJqZu3/VYEqKR8mkujICCfJy5yTN
sUyoBZoBqGnjNWvHQQnjF0eCckyVjVZgqUVjHzBL8P7roWqdlo+eICKcUrJKElZs4/o9OsiF+oEH
xNR2ofejkGWCam6xB4ScQ9zTXA+eOTQ8tkWf55YD05pyUxhJuvYa7R6ks+TcoRGWjLbekSg/o3IP
UocKicUGfenlHAZ8J5PbaWnr/J+5a5E/U2kDAWkGm7LIaCF+dRo81Uh70g3xfiMJXh+s8NryTJj5
hUEIMRioCRwl4C3B5SkEaR2I1YwNbxQL/OWJnxjavuu9gq1O6MRSaVYR6kJlzpRL7caiX+ZWJ/yS
aFgOEzYRNe3y7t5CizSw5YbnxRUVQ0PdlgttW4gLQ/17nAlgVQqPs5mJt6jK67yX5iZSdAhWiKKp
K59KioXPsZfm0iK18Ak6bwMg3aIIn+vP5eO4ktEEtFmmkyXnOGU3pPmrVKLJTbJT7ux2in9XvTKq
Vq1/w8DokdpZYEWnWtrHaI0fUBrFH4AACLYtjmPtXGEA0HLTX2t0sKlAUw+9oA4ltVzLfgIotoKh
AJT8Lv+kbtSduLM4XVvCmFuIkQlbuXpnmmtlk3jU+ASkS4OcgW4ToFDomu+P34P926Vhc5Xmmnbz
bxuuQ/+4RmiTyC2fcLj6gV3jfr6KEKCHIBJtr26rq2O1peTbBHVtGmJs7HxllfNdQ8dKOV4Dm61T
9b0goL2nZpha+ERi8if+9WGEnIfIxPyQsZwyGDc9P5AGj6kQuqmWE965g6g8RDXHPdwCeIY6mFrQ
TETNkXp/UluYILf7E0GqQtyUW3+VxjcmkoJXejKaA8s3GwZUIE9cPz51qHSSfkjY7mJXSuYdD1dT
tI5IphJdhZXqyv8NMfx0CRtBhEnrDWxstV3fuHUfQ53oMtcb0/5fW6a3sYkfTtLE7/8m6reOk1rL
3gHV6ayGri8s/MFGHNaUHGOBtGoosNW76uTD4j1sDJjUF+rR2+KIYz2/TuKPlw9ppdYcIOCWkagV
FbM8q8qnzVSq5SOWz1KUSFFE/Ho/ksxarEiBtltr3Kuepqnx6E4Va4OhZCqrwX5H2t37WfrcvWFF
QPv2zlBk5edhOdE49kVi9pB4QP0UeX90ZwCiXnhBOtBMoYcsMBdun9zslPyR5dFx9cHWbERqZbA6
tGJVQPEtnSdVfE7S+GiPVjZfnWD4AoZGuBF0zMgZh8xmhzUi6aiNf14P1kIGgX9il3Ptho/D0vSP
G715hp1ctZc12O2oqaDThdrhdB3emk2GnjpmorExQdQzQqZ+vZsZ4baQxuCehvYcdS8zJ6XK5+bz
31QLSnw4tgKefOg5Z0H/dtiGN5IzSczESBusaNoriFfgscWtEBX7PpnfgL1Yvucw8tydzAO/xmoz
XXuKmraScZu0AougQNAw7J20PbcexfGiEzzW3W422hhq60/ZlIXV3XhfvHu9wsp6Nkby0CoypmvP
kKYEybu1mL8SHXAMj0yVEgRzRkEn8T+MyKI5Ao2KBZ+j6CBcaQe7M2whWbxCgMkXjdYsEv7SIdEK
xliScQ8Himh4mR5R7ei3sZydd8eBPLfq/EJk81aaV+C6csQfEea4EYSWnh3iEu0pqqCdui9QKoHu
eR9DwrAXsefucJ4o6fy7zsqPM+BMwaYf+VJPV5HZhMb+iaHPsx9tPVJzuaK02sXDeebB50LXDNHV
Blsd/sMjIE4POWo3/Gypdj/6b1nSJQIXX0sO01OID4z9oVneNNhNCvLfbQykukDeoDcY2VeiI7Lj
X8w7OPMoaIYM3fbd8ylorWW5Y5HY8NwERaiDm6qHgvQMzW41DD8BXtArF7KnXT1PypUopoZrysA+
6FSfspqF8bpT6TuqMhC9TFz/ni9w3Vd5aG9EBrtBQH+cDdCmeKrZXuIt1Yj8sQCgQcsFfJUmc8rv
sJfnOU3mJaRA2OXCdlZIzyi/owRkTEZ4YsVPp1MdZ+JSBIPAB9E5qdwrdiqRCXzhv+TsVkvj32fp
zUiThpEToI3LSLHDDb/HT+Kq7gI2LFlGjcc70x+xd3HJoPPbrdPjgPzd5odlTQUIbYfn6qyZ5kxg
SaHxLchqnmUl2se1FSilCjx2yF0LV0r8lwnQd7Lsq5l/dT32NQnBOEOF7mrGIH1AYjx78GW8qmlz
o+XT7AshXJpQtJwL0mRgJtHpHZgRlN5MdFBUpweTiDWI6LqR1BvnhZtzO2+a8PoNmFuxIuwAut/R
bKuFCtkzcKrDA5TpoIY1CHB2np3GBeNfbA4CUQfHplrwPG4QTED1kLvfGFEpPr+W4NzD8AJvostn
GcE9BBcPAGqargLTAyCQIGssdRC6hiSHpxYhtT1yHZxI3zyaDAfNCHU55akVJ8AX/jJRMfpC3Pz1
5f+EAmh9d1TEKvweWZiIaHQhgwbKPOgJoWCcJNVdzg5n6cQ+sBRgq3mtmJqvoUK6ATq6gqNKQEvH
rTNCIPvyUad+6EIXoWNtt2/T0sQpbvMd2JkEbyfHV4p1LD/o4I78tWqUJ/jESg8c/8HEROTelD1D
XGiqoPzvCd7OyJmFBoYU8Q1AIs+9WUn/UjqoHnMgCkZEpmyvOKtvApktPvddSWtB44jlw0gETMXo
vc+0agr+T33Rw+ljApa462HcDNIp5aCWlL9EyFoY8bJ0tQni5SBDkvJF+zFfmtgg+BL3vw1944Fh
RDHLkBOSgbetQs1zwoPfL2pxC6gcTKOd0k7iiiJ3U0kJRFT7JEBY9xF3+pyco2L6uUwiGrJQTeS0
iojtc3NvbE7lO20pbnWEdLOU952HYCoCGFfwOEOaK1O61FYSU7LoaNammm5QQShklvarPzTusDKl
zLOwTuPekUs5d1VVhIP/EVNQAvAOmVBZInCgKwU7j6ERpEw+TgHzHuheoNeoCaz2FNgLLEAR233n
DAIcxcrrrv+w9W8xzYEZvB602/R5MHXNFK7z1KwrZ9hW0fL8B0gTr6sJ6b2kg6tV9otjByhT5A49
IM7Ry0pyXM9Hj8vrGqc7RQ470yhmVYsv5kq0dKzQXzCoPVb3qEJUXzvScPlUrQm52s/5UmhLiqwW
2jcUp7bw54eUCWCmj4MRpFBC+jx0OlYc7yWwaOAJa0aIQqQ0DGP688GHGRpSw1Kx1Um2ONSL4eAs
jH4M76UhdqFvyJjfxPDIjZ3W2a64CR0yCJxkhPRhjPPaI+ibusdZBJZMzKWOCE1pwtYT/YCmfbdg
8MHfA4vv0UixZYnJl141inpCR23i+2Sv9c/wV/6UZxQfPijds1wNiOZW4UtiIFwr5ZNHpWPo+R+j
XnpkusSfmgm/30ZAXjBlyqb0W82v0Gxx6PHhkF3YuLtOqDGqBYJfGUid+CJ+o0pBK+T5XA+arxo/
dV9RtJz0b1n88petAI3f3MkMaYewISeQEXd/iDaZplz86FvBHsOqzPepiMbzKBnQfwvFXzI3K2CR
CtDHmKkwV49pjrc4GXpCij9CORzfC4Q1E+EjVdQo8ONr3fOTeQx+u0dJfIhvMbIlqa4osMUqd5eA
yFclFZY308HXhJZxo33XYg5QDnDwPYuxi8uaL//dBib/ewEMUubSQjl+mAIJxETDh/TKK1zf70QE
CM3GrC92sfL0P+Y0iZgTgKAUsbGI3M8KErwTD66YrI6JtdX0ko7bgi6e9cpX7/0H9p8vlZw7XP41
Xs9uhUQFA9oQlgpZFVVWFCQj+2ElHzDoGaHjTFzLUYHffGw9NqVcOk46/87+RcCzXBWId9MgM3H6
CFeWU+TIncasq32lVgEsvia0f4RcgzZzmcq14dWZ5bbc9bkeNFH4X4e3pzSizM5rVlkb/0JGK13G
3Zat0okSO+zi5ONeLJg7FBZ/vhovF/JDfqfgpsUxDvUwx53RP56CNLCYG20DCuJKW8KT6ywebbJZ
N7AMYxJspD66lQYK3EuF6h3elZrCeDIGs4uH+WIrphjy+dmvwVfUQZhI61TSz0sT0m6s3fgA3i0I
lux6LBsL7yxqjMbhLYaWA+f1WfbBxZF9sDAn9oO9rpCfvZqohHpyt36I8eqlZR3UdDMju2P8be6L
gFnaw/LZgbjxYs0zrQn423CgLl1w7UhSeWsCzp4Mw30LIbC70qDyU6IZwm/CrevfBjJm14BWozfo
Nj+YoKjsiPY5ef5VIrioQjjveP5wqwJVqjoqXqBt6madR/l6oJBtSGgSx9Sb/a1SIKI7KFYEWZ0z
0eYAbHQ1bX5sIzQtFvojOLIRQra8sExUX+i85b02hpBqkS7VPJA2KSpgpfJpSiJjHo2Gtv2czTtC
Zn8jtOpq6yBhHcQ971OHrZmX4cJPPDNAyfMpFLgEQY4MC8soEUoFuwIoCyRl+nATRDxUZHOQQzaJ
EYNVJa6mbdqEmKD4qqqd1J5z8/VqWweAwVc7IoZZMU0Ind/9pmPRdSmkC16suUpA/JqVWj3QdN89
3W/clJP9a1sHXp67E0ppTZWOmK/+OZy8G/gM2JyMMRDupguXRPispYbatLIBLCArlNY8ZjV+7sZ0
3BBf3sAE81vyTzQE6eAIS/bB0nfE3ETSVRNGWg4Z2E1fANvvV2yrw892wxRJR0Z5QVLQlTUOihkl
/MBbnjHWBaEYpyfztMdyVJV9Us1NNLkNyTmyx0OsUC/M6ByMhYdCGHy2+jbxPfEHg74AFVmhVuao
Iq9jUFYmv9hu0ij/KRxmhowrH/GYRl03D/pq1n2NimxH9twyDzd/HaTfUZoaXSR8bZDhMsWWJAPR
dUUPKN5g1bdW3bQgSqvvSrMRInGDUE4sRwkLR2AjQ8qsysU4RHXRPXKtVU8aoZlTxBtkDx9ZrUFv
gOFkYUEYAi4oFMulotWuKNtd/7Oy+bQxMIRSqTgI1ccnCnGxwhahJdGgFIaZabyBtHE6PdZCEUPG
OAbx/taUT6dmNiwFVRBLnBZTOAwipME5L07JQS9qcnG788GPV7BP23prNXGqgwFchZRxjynQr9mb
m2t0dPbXo6Ac9LaUgnegl4Ny67FRuTTn5uWiir24o3oAn2cbuyHGqUHa0BpvZ1Ac+BC/T3MiWNbk
i+TzgSNzlL12eDmAy6jgj5Vi1iwwbcT8f7wRlDeUfBSkiKA073miG0q+UH5VqV1Jch+8pvj5UZQC
XYOd4uNgh8/XrjFKhlxY8FncIboffJGkt7hRrvpx5v+NT6PD/2QHdMQpl3Nd5Qz1/SFplSuhbTIs
ZVi6qFuB3SOljjahfC3PUmDaZj1uewOJpY9gNqzPzsuT5kBlGvbyz22g31VXe+Xy07cuuW18PK6q
VzkD93Hv9B5d6+6LIXSWNOu08wT0w7N7fqC+acbXGDmFqImON/KWkExGIQrwRXKZ6MNnEbqMHPYI
gQJeXENVa6fqHVGVrJCpNgMt2p82kzSdwY4YOY0ATIYGzXzDPztOL5dbY/rCPqOQWCtfr8INhY/M
OrNt6tRPuOQ4M9xMQ5YrMcz0STj1yFp4EWyoR3eFRjYWpJTbUHF97n4RqbiA9hy0+hIWnoJL7gj1
8xjsQqTOytzkJIrRucG3btQO5u3N9JK6JAN5MD0ZtOA6AF/hvpzMt9ZP7b37DJqz/TDm58gMvf20
JAoqN7WzLbLw11LUZ2ykBMlYNendV9A8vu1dN9FNVbS62FvM6GomAxl0RLObl4nsgnLZIGILzWnO
oFmOMjx+KRC//UlbXfFveQY+38tf758WH5vK0xaw4o90+55mJyumo7xban6353pmk6xPraWLbun8
OFNVPGxNwFwvVnI7cJ9QDPw9Wtc69pddAIGOpn1vZ6kBuYkDQV4nLul5sSIK5HcFzo5HsELu5JS7
htlRh4OlMcc7nvKVMC7KSgJyGZJPgvCzGetbV4WgBdcolZ4NU0VEL9R0QjwOULtOM3dLQuao/Sy+
57EucYoi7MDoeoEjg7qj0heT12bKsKUvLNEwHpP50KicvWvsBFHypNgSzU4sqacFPqP98kpBsThR
vV27MfgVQd2bvNBIinYVqa9HM1u8b8Yhv/2lIzyyDCE5goAVgTvN5R6adyks6tKziKUtUG9JZEc1
h5bZVj+5FTkVbq0i3ayuUJYBbIVcELjv2KGMuBzfNdHS6etj3kBxrHOpIOLZe4+oxkfIOi/wuUXL
5AX9ttENENRBvx+k/7CRSS52vts6vvmZJdXXbDqccpCOlaEISi3x5sjs4DVqyz3Z2MBx9TgZy2E1
e1IT3zkNKnE7lPtl526u6DE35oeCUxlkEh5MvhXCHHpeTcSVZFvOYzmQQ5fdJtjvR6Rh7209j95/
+4vPrBzMa7snL0q51+XIZ9FZFloOu+o9mqdnQk70201hSARp963zN8+qEs3Wt8nPtzVcfTHl5zcs
5o6peXQ+KKx9CVqSOWj/A3QcP3xN7CPrltZDhw8fqJaVI8bzPpgxWuCd690o8KGjaB+92XJmzoeW
QxtpemwURksQFJ+vhsSVcy+nWh+LiC9jXeJkX+ISIORstBRGzpzkdh9KV2I2hg339AlgGvZVcNpS
WnmBW/plCvLmNAtxwnDazAsfC6cBqwu6VbNVgR6J6NKSboS68LsqUjkesKE3Q/Typ0HBh8Ppid5k
cYm7spwIf0fL+0VtCqA/Le6x7iNlUl3zyfaau5UwVdj6abOj44sn6ywmMV2iyH4oXQjxB/iSKo7C
a1VvqTCAhIiciqDo4qxR34M8WdhLj8yshw5mDqIT0CZ+LrHQC7z+0xHy/doVPm87pyxYX+9vLIWe
sguZc00XhSrjWwmbtiYwrlgnqBRqFYMV1hYd1IshtN8oLfqi5hOxSsTg1YeFlst330C1hwnGc1Oy
WXQavoAJPoB+V/OvECt51QRWVkAb4bAAcgFrgPnmcTVUDJ/b5yHhIPNbunl+hvUmFwB+NmewPEmb
ESqgnknMqpmIQXn2RKPtOyCUUK/REvySyvBZNGBRF8UT5FDIk5/DljeKq5YBn7dT48IySU+yZhRO
tOxwlejLR9x8kPIq0+Nwo6/uPmnePJEa64E1jFJVQMxYmsSti6bjZ+2JLVKtnwc6Qxt5vdKR2umF
LdWYT5h9qEqEGdw23UrhyCMlGcIJQX9o1UA8uSt43TzMGKo7v7hfCLEcmxTMJXvdOtKAfI6nkBFV
BwpLl63TMWtkT3e/dVuHRV2VVRpc8kbQn8FKmaUKVmQrcEMZuqnCepCxp0cGA466FHYT9uyY6Epp
67FOWPSR9NSK1sL2mJ9JXJCvzOZxEhrZqBcgJoFGWAS1ekQPvWZfflRCzAGNh24VpW3iOyqk25sC
9DvSs5gGOze2VHG4yXYsnZ7dFO+RXkNCuHy/5LSvPOdGSyA0hh20TGB5C1XyR0YZRsQ8eCK3KD1i
Q+NSeZoaFyu4CyNEvgWovn1Pg0d5c6toAp+RGOV51bSlyFXCw7uDAUUPRQf90WB0VLjLFthtYipI
8XjuKdNBMJ59KMk/EvNMayj2GMeZVOBFsPo+jakbXbepYdukOnDrpQLHPCPvHRW9XjfbxN1ECBfk
viM8GqFvyKEt8FkmLko7qTFnZ8OGnHjPM7bXj5n+QYTgDFI5FQeCUbN04SCA9UiubUvgaj0ILxfY
xbQnVKvidXDLqmrt26i4WOg/tLfl/frrW+SOfX6hhvod7FNpcZfa3weRv4BpcYNRxxYIyGqeyu2t
AAtYUxKflcLfN13XOjo0OIb/v3TadbQIwzESudGZ6mEiUne2N0EQQ2Y7iglwpawZ48OB8mkEh/UG
Tl1W8Y+i83uoTvn69S4lTzNgKUxtUXxkeFjISnOgeImsuRZGMQHyl5zVvOLjqL6U3ggdSkK789Fj
dulEYK4GDBnbK0QDY4t8tEWpDMtavIGIgMNJqgK6PnjAX9z85B2zQtXQRg3HmWuC16oLGcjjSTzx
OXglxGzYCPQlG3OX3i6Ap3GlX135kOwIQx+8Ejpdxg0h0I0Hrn8MkFprm4DO86hSFFCPWXKdIZFE
f0yVrWHJUECZTWOBOORN6A1PEIcky/EmyDUDr8Rnn5um8p1wZQmB9oD3tyVn2JFXZDc9UrkOPzIu
ex7Dl/ZV7zf6sjCkOaYVnuemAWgtGb1t4Cq6OkYzfCh2dYDSMKRBVyjdDLjO45wjWDf5Nz0Tz+qu
xdg+GxBDrS5VMORT3/53uDdT1dRgylv7pPThMSgNaFtDIqpD3KvGrVWx6fGR+3Rb4G1y5WbX31E7
UcKS7nOjdgsP7kmK8E/GxWRqOiOvtb2sElmBXmHHZfXJGrdzBt3YGEnmiuGHKa9OybRPu7C7vAN+
Apc07wRsjKrYahWAROaDrPAdVGQxNsq9ai0Zrit4beY4S1PJ3Hx4r0o1dsC9ysWvOGaJmoXIU7El
Z+kRvLRDjygMyHYTAB5VerECbw+dfKGPQPW843IGr1obzlRZZnX/UExfVPXBLC6Jv+8S02KFrUbX
CX985jZiGXcOpWD0S5cYZbEY3dEKuq6bwBp9wS6i6PfoSgEKWWQLvcTW+yXeZgbolZT8vdKhPYfU
mosggi3XD75fj1enqcZy5kBEBHCLYf7ppQS2PT+HgxD17DuCXXbtd0o26EJ4ZFsvfr3cmBTorMc6
QzQJT+rfKuwSFdxsdYJ3+8QUH/N+yWROIvRuWZjoopLRDRIB2fqv0PXbH5CQGOSSn+p32eYwgWDB
TD27Jnd/cZlLdaAa5hyVec36sZJjYnlUbPToYnpcDXLbAToF9zfS6F7h6L8eRu/7FO3hAf1CBIcd
5A8LyCsGSzDq6JWC6QpokfoEe9KSOh45R+PZeAUUAHnOLSCnodiznF8CE8BVa/MmcZm/uiQUBzH9
eL1n7VBMQBtthxk2JjBfcWouy240lM2NMC2tc7zz1eOM2Y+HS6GLUlrcM+TnjtcKKzi2uU8oDM/Z
5DRve4B1lbvu7pZ8DI4cyrpX8/Lrupg7zggY368uUUgHeM2bmo5+iFp6EWJzXa03uQXETLTGSY96
Ndk0whFqYtk+IvlgH+RhP5FBMhlQb5/CXmksoQfW9OJkh7Jd2ZHq45TbImt2wjKnyFJVFMa3TXHl
hNIdpcrYX7CFw1rd0kwXKlsM/UBa2VAwHg77eu40Y6G1WSZEgjRTThQCZGdbwQQE5Mt+4ED7AGXt
Y6OapsLhJKVtzsQ0vp0M3dWVkveV2JoUzDZGzA6717wdXCGv1clcPdvuyZbilrj7oDtNUgMBCljl
0NOV17AIiIr//G6ASTh3f3xQHP+DFtsQL6YNn7UOZkbUBxPUt0B7QHVs9avo3G7cw4E138dIO2Oi
liqIHeBUffq3uHg0dMaNuCYRpkVwHdjWn5vmFQ4zhaJoPjR07U+R+w4VwrxhVMLm/KTdDslJQEx8
An+5x99UKcnxMmlYkIZz4zJidRdnasiBKUvcOd2NjG4Iu4LMztq+mrl/bseQFHt6devpQZk9wslI
PiBL8Jfgllz/0CKiSV3pkMUxj16IH6mcY687NUPyDiNtxpHL93BbXehZkLjjAsYUJRGszoaJmerU
W1vEbp8J61XDIp9mMK2PIyuVBteu8d4AS/5HHVM70cnRuG90PqznNh60oUi8NVq0ufs99vmT/1gA
oyNk+VD7xdOFtQEhdejZkNou7ZI0DQqhtjLKtFktHGFOFEE7Br7eSSlVtMtzmlK/G4/x34bhHFBk
rnkRmNAJjaKAexMSPJIWn9sCrO6vuOiO3SgIrutJRPKx7Zhzz8On+FerttOit3DLoInUEzbiqkPS
rKVrQBKRWWA1M3WIvQdAIeso788Vc1qARD/aLyqjGQPncgpRZv8GH/k7yS443uyE+AZo5gDXpEBl
hD464x/YSb4Iw9sLC2/iGDXJHWt1p9ZpLHr8I56p5rNk24SNotDLfQ+E1BaVIVbwqIoHm5QRRX+d
nFww20HRsWILRfN2mytfEoV0BaPlxmd6q97y+vxXI5O+HekOwd4Qf7smekgReGpufyqDLJKn4LxK
x23W+Nhr4E7Ovb8HjEcVV3qHe9EJuEeEJ/cCICpQ53POuErYIJQFCRHAVoG2238e8hsDJN1u0kU6
UgCoOvcGSUQBI9kwnls0XXtgwaNvzdk6wIc42eYPy/vmzSke+gOmloAmwisRL0Slabjl6SEwO1dp
81Br7r14RlMuA//uXmYVlDoKX7s60xBuymv3HdEXZRVz8AwU7/u989z76lBj0J5uSGvFHGQ9sjO9
EjpHdR2gE9PcJMdj9rqXa9uo1hzI1e5TxNx0Fn8/ZW4mZuTxZnjXxW58Yd3JplwKHH4d4RVpaiWu
T6SKNPF/GFjd0ZQIzXb4pngNDg5x+Anpw3En+KgtdhYh/dN6AG/ooMeMrRtxOlCbHkYdpx3bfZz1
n7gDdvZlQP5LIVJG9Ht9mL+PRNTPsNCvEgAylGQDPPDTwb/klz2ZsrWxwPlOUlRs4+Lk778AgjZU
G4w8vfE+/ZqHZ+xbiYGefXvPuih56lRkBCoyyjrFPfiNMdpJ418Xp6n8GY5lb6jGNy7QI8mk3Vau
FD82Wg55fMuWr3l2RlDMI9pG5i67hqAoGjz3qwA1BMJPD4EchYIbHicM9O2KwSnG0hCULpD9xBLN
9ahdBxtotdB9cOxZQpnX6QRnzCV3nFNLgIgxQo01oju/mLQYByVjimAKhzsFLMjVICZxNiPbwEvU
TLwq8uMfAaDt/etmbe1H5ZZJMwTeisu27V74TV6hWGfPiOnyCJ1x5YE736zE/kNHYsw4gIUCYSIJ
BhEa1yIcteQT8a4x3JfYGRzW+uywb+9gYtqRtwXiCoEBGYFpu0xNkQYc3DvWOq76YVqVLTSJadaw
jgbDcGLQAYGamEcYWw0k9itOwKXd0dmfLbqYMMk03oEWTBfi6CPOMkiVLC36itvYJlxy55BvmmMB
YaAcMxoTPFjER9man4oPB76bbBnVZmDUssUL1sdJMpRIwWvMx3mgwhjt/g94ES7nZSn7txIToOso
FOdGfVXCG6gOpNj5qzJhKEDpfkdpGF6GbEDclI5We7qgZ/WKWXJEjj/k07zmsR7jFuzDuSZlZ6X2
XfTKy9OjAR2q7k66pOeGk/woYyo9Qf06BD/2Q7MCKBobTDqBNiSXV5yNxe3lEfm21u+AOvy88GWa
Y0JPhYwP6a6D3ZR6RtbyPvXlUJIIL/Wq8rnyBu9D9WL26NhH6l5I2cHOZNJ9x9QJWb3Q5UxDNLpA
FFdmY5oMFQnBdapp/SvB6spQgEo6yg5PBl65CF5LTxS3M97/T2OVEufwzvw4ZnVRDvlh12fxnZPb
LzbjIiz98KVf2+3t0lNlVZCROH8H1UtN6LoarwPRfuAouwWnEaGKPFDiKpfwHtjhran3ySGMbkXY
CSZ07aff90fKO523j68xmdFV/WlwSo7kOA/ALUPQj8s1XUW1fl6GaHnZAA6+Q/s5dD8fbC5gxjlG
m3MVaOzgQqohvNieU/++oAWWNSvSPDxIp3XTJc1vaaBtK1a2cXa/7CPBDPwuRIMbRFLHHhzDdxUM
X0/hz/2xYOIbeYC9MEeObo1kCxViH2Pr5psStd4XoFh/3fN7TD91wAHSdf+1RNIfCw4kRdujroi+
EsuV9IOtYFm/8iw4aqoS6+ScMoz+TolOoVUemO0COymSB+keOZX04SBUuQZ0Ry31h/tm4MajQWdC
KyxTzFPMJ4kKGLk/Ys4EhaVPwC50662PG6IxUQ0s3CFs/qcherooQtZcuAk5nNcypoR/1JS7E5hK
+OnPAT1VPwbvMONAYsq6564/5leWDRi82sO1J16umT/kwCQwM0kOpEUMtISAZdPHKAi5sFQ3jYPt
1ChfWv7O/EOB7dlZ9zDMwruczpStodUue5KqWCEiqWpCOjgG7ALSUn7MHUMgWKr9c5+4MLhZ95pd
bpaMUlHhE3+nEzazTLVjbTwmVx5dBqJ8n1Wvdo1Z2at6C3ED6Mdb6qgWMtSnhF0U8RTk+Vxihs2p
ewl55yO8Boi3IhF6eht6NVKkaWPpuQtvhuU0lJy/Hx79CLVoN5CX4AEfg1n3L9o5KgzGGs3T/UwP
nAIkGDnzbmVbL8frz8ZtSjUSp+9XSg0jlH8wJjNoUgIlFgumhFCquxcPD/YWw0wuRyshHe9hZiG2
HA3+jzJf05IGatxUnddAWM2fOJlBVa0Ijc5jgPcbhrCnIdKTaUQwEwNhOAIgkb42Bv+n9ZKq4emV
7Hbh2DsQqhcRdY2g5YVZmoee5ahXl3Xwqf8HRBOuL4BkbMPthC0kFpUPxjsz996Rjb1hrxWoYv9i
yez5Ccb1pztLHQl9yPXH3LToKZexEpoavl5a92NhzsIzRFX5TpqxkfU2CYtlfrc56st+EGltxDbk
Zs1C3hb9rOuTiu6E3T8bFez8nuUJvWyu5CCvQPTlhrrbEYdzNnos+pTakiItwNAESNKRStdAsW4L
5Lk8pgxVrURs0xkRCXugOUtTKlBBrOK/kt/KOBSdHJa8ym2i+UnNzngT1uAu4CJAXca8I3GQlQIa
Mrf7j9xevQQAXtE7XxCudYCTHR+1J49jOMcasJCM3nJ8msIkZDVRvhPFvwDPB4ocCYlH8BbCNWj9
Ndn1YGy8O+wHl0YNZUVZ6ONtwRxjjJG1K7f96F+eUKM2bn/7pik8KU42Y5qbSOqOxv9DJ8AzKWgN
ub4wMQAZKcFQuQvlo7EUvnMGYzErDbqrE4b3df5SLedRV6PbpcF0FwySW7TLZJKdVy7XKgNRdUDL
3a96QwC6UdCnSUWY4WYHj745GlFI4ZTuHaxk0O9AlMbJCSUfrnpddY+qgO8UDQEJyzgo48GWy6EM
cZkk71X+lT0flj7CcGeHDO1sVBoYV8vQqK4b5Z1Hz5YdpqxOg4AOqeDXAUIOqFyYxaiiquPHG8Mw
fWzTn5NcWeQfiMpZPXL9X3TuMFQRSkh3BnSNeiNwIvjjNtGz0f19uz/Ue/hxVdzJdTwIP7B7YIec
nw80CtiuCtHTU8HM720Zk5LxpfRIKnqmn1WkedJ/lp4pek7cLajKprwqVb3KONjPbD1TnUIG6u4K
7LvqdNq40p4gr6NjRzkj6Xst/+4jg25GHWa3QYYQsMWst6Mw+U9l6uI2AiPnH+3Ja+KyJG28xEy2
ZhwsKER5p83MtIIbwRkiIp0tIgptEDj0zMj7zL1qCQIRLaDuQ8zS65SzsY0C2Qif0Y2Whej2256Z
5ZdDuQUjoA9yO1/1gGnMLvE685C/FCBQxwPxeFqh5UaoR2mMYiD2ErGTMs60Xu/cmHmX4u+yWo2X
YMGKNVO5JIbDvNUGF8ZBk+OHprVXIJUxJv/57GpAJAsS+LXRvqHC/Xr5Lax+Gafj4xMlFG9Yb8dJ
mPeBaPeR7nNCqUjtGqdRMu7wkrev3XAqyoSbuFbQSB/FhtOeemzZ7/tCTwloiqGMgrPnNSTft5f/
dJY3avRu5TYbEd42MpEnvhTaQuY2zwqewexUfbB4iDApHjl1v5sSH8Ja/xH5hX14kSdnN38s2SXp
t5GHmGRYHH+aD2g6YbIaBIRx5QwnvFTz8WS0y3nsAv7BU27ncf2iVfFD+H25uxlW09koAyLy2VEQ
ty8qRZgijCLE9iCEe1Re1w7mtHzP9iH67vZA5BwO4GBipRSBtSM5IU4yS1mv9fDAuK1P3XXYC1B/
b+7tggKYJYhiBXIb6gzR8J9QmKFGjg+tQsGho9McYNddMHBGu1okl56SXlwG90cQ8Zv5I8u4QV92
b3opcNXIsL5/+fY4ecUwBALeK0D7eCjaphE9Eav3JpWg/XcstFBTqXE3fiEQUSViV8lnxHYZjVl8
Px4s6ISIcqJNwG/iW8qdCGHQW3NaJd14VFR/FCPeLnSssgW5B59/C5n4ZWXqnYVZIpNAo4L2K9uQ
Ku/WAu2YsT0tVzva5Fl0GdEJiSrCBL7oX1jqyv+2SWV5Vsuj3/kCPyB8hVkVvJEcXtZUMs3uCPg8
/2rY9IWgqyXnyY0vZQKTZbHdynqK+q/nMjlubyBvB8qXgFRByD4yAy3wr8YcPeO5MC/KFIgeELnX
cWJGb/7mSAc8kDeGscDsJxO58a1/f4JXm+uTVowmxslZpyQlnPY6FZdVOn/AFQDWv4VbMdmzoVAg
g4pCRjM+uemwYlypt9rXbQXjRzamu5IQ97u5SKvHcYy4CqaM5Oj+BLOE4jvHCTBpwwa4IRJdTT2/
IkxrZbOL5EdtixwQ0KjIGXmAr9xEgxqfYikZbm4gaRXvT8W4nrryQG3aODtzMZ35eRb6BflS9ASf
trcKVWc3bXjenY0ce30+M7sPmkrHgbpEQWMmhKF9tTGIQxci8B3KhxPsFlC+m8P7ONadJomcsDH1
blCvABhabol86MZ9eAFtUh0a+1xS0+QbJMWy0xJ3sZG0Odyt0e1mWown1SQ94SJ9km/n0RLNddE3
cz7hYNCz4IrLWdoPdoMjlU9mN5rWn8GFUNbTZ5e73VbdyXbJFHrMcLsqa6NebHMdHQzxHSTYIa+G
uKOFsaeSxtFlhcM5DfVTmp5YpbHi4KsEMC5cEwx/D0Ht3ibZiZrLpvUoYu4BWZLPN37zxWeHY52f
JWcE54TCdKFmZyYWLDZHoLg3eSOS1aIoGjoNKn/2+2dNUKvxQkfG4Qu5mOQRYUv+0VGHtcSd94Ra
bWcPKa1bITZ/d6/e3Hdfr9f+qG0xSrdM1BUkrIQz5BOdCJMVdKcpxf4JPQUoPJ+DCGIlrpnDIoZ3
Mbl2nkqtZAqrefMkrwSK/QRHeRxw8M/oxKVO52difBSv8QK30fkccfevz5FU7e20pKFdWo0OqamK
CHTP6AX8xTbK168GOowRk8a+gmInOJ1OcNNvyNzqF1Vg3FGdIZqQs8QRunonzmdsDuMZZhfDSTkI
+9vUW1Zt/EVoxL6AQv6C1S8YiW1C8y2amufcYklW015noBMNN2TU5mnips4uBCeXsGOZj+9r6FMV
LUXEW2myChAeBzNEQXmgehAntne/EnLGsUGUHD2iAE8+yLIFg+bZN+lqZv9PLp5rXKGzajZi9X+9
Mi7XJUVW6CjVSPl1Sy/lSPFOMfG/zGuMTBkNsa5YR2JSVxcE+gVFXkdHZs43q9XmRcPnOyjjfXqW
uksuu/C+gAgM80ss3Lwnj6fjF4OtU7BKODAT358/J4XPYXlxhTrmIKSGPReNTh+YNH4W9rPy/mOk
0LaW2PjTfeh1BGxB/Vq4x4gPt4uQ5aXvfhcJ+HBY+i/5pPoVd4/DKgNIXJXEfgs4Od0yUCyU5bDc
DsL0nG9WZ0TOwZqpcoTGWYSbuAh2ELsnAOR2EDPQnvNFsuxjZR/CS9bRqGkUu7/JEQXtM2lkmtzC
8NhtjjWD7Ubott8zpYarkrWD5YC6MOpLAHfFHoKkXIlX2RbypApddM/g6WPrzYF/lTB/PLMkgS3X
W4dM8rfLnhPxixFRBTMTABBp9iuOxV2QlTSCHWJQ0B4D6RXk3TqhYMZeA3TIm3RY3mubbWw/hEDF
CIXX62TtfTP8s1h8CspXcfMu1UoHj28bMgOmT9851k3Cqgmnwj6Vc+ruvMs54EV1pwGVwRZJVMqU
AdlAUY950aG2UiLa2aNTUQ/acnmAHMJvJPpAWzGrLAoBw33oyIqq9wJxMDKChqfYSdlbf6L4fw+/
cZEk71Ij/HQQFyAI2GIMbapaSe2Z3WgJifnX/HygjgO2H7ma0OXWagSgHct99+cAeNCrgq0j90jp
Q5k4rhClqe82JX9RFf20vau8bg7PgnhXwgyrNyiM9Do4Di8Yt6dU2d1zXtC6Aqm70uol28pTnbV3
w1AH4DE7VDAkMm66sa01/AqTzhBtPF8v2ZYw4nHczpCnIMsas043kNKRQmbKl6Ks+PK6gkAZzKIs
rHJEtyRhkOrnps22GQciyzgG+IxLtTc917FVKGqd+0UYwxEM3Kt/v1BCr0QLB19rgxcINzebJ4MK
fQfRqU7uayA8tYoXV9E1fPygT9t/FBDSVDf9zDizqliNf04XlUF3j95qmSbMQw+1V08wWJxZwvZF
DBm+4He9cgliKrtSWPNo08ShuwPQhhwt0qITTzjSo06/YpcaHheJGi+7wOZ4Ksfv0O2uUUG80jyG
Xkx9Aj5lPgSjgURW6iUA2EFpw0k0MxGi6TlVPAw1UeQHkFNG+jlu4b58FHr7iwUuUbkB2l7Fqk0d
1mgtl103UNCbS8+8fFreSQ23GMtBBayMNgIVPBNuIQ9zdIXZky4vYlO3AP1rT1Y/47SWe9jf/3h+
2FfyYc3ceks0LLga2Zj6gHuL3TsSlIjm/65Ex4loI4QyUMR3tJ1z88i05KFo9wLS9IvRGutRGGGB
E69RlpnLqhOx8QiHT+RDMCnain3lsdynOxVMSUCCn0TjMklUvWLhMgVF2VjSYj0AY75wIuuBZJSk
mu3YRTe2ElFBdiNFPOg1L4AhJE2SJJUPwE7HVZzytdnrAWtjL+Mo8Jdd+DWlCdqKejzlvqNDQG7W
XP+9+UxaPCasw3FbBWE+SefecvOJlRBnLF4s5njBtYj8A4A7N1JS4DBf70qJw7Bc9NxHCfXw4DK8
RaF7qoNRD74Tyx6oTgr+VQM+mPgwl8pWIQAFKoslglBodt7GL4nOnJu05WB4u7Xri+Hb0mYg9IES
MmxESWueXuxqk3KfevcnXzgRwFJWqngjIs+7X88Q4OssKgna5YKJv9OiGQJoVXFNM47scZpl2AxP
OB76XCuRDCEIQOA/xQA7Y2j4V/x6aIAMMAZmtxwsIfFk9d45mdcioqZgRrf4BKVG+gbZjm53xW+o
BtCvzDiYSu8Yf7p3ebpEzSVJkxYIVK4h3HmLNcH7hENfXah7K2u2ZEUh5e0JFvCYjb0/K9Gjm6sL
NzcDxL21OPlIqcD2g02GM2g2CyiOa+1s1NtG7WzEMYEN99n8gvL/cbTU2PeT0+gKX9mzeF26cqlf
EV6DgIDsnYdzFxzhaTf15X5GVeSqZfADUWtVPNmfzrlxXwo6xcuIfk3oDG+znMAU0MUNzrkI9Ivb
Fu+miHtKRQL1RmOsp22U47tIHExA8HnwQ6sSMEcea9PtpxK39YFPZdCS1GHY3GJj/8EqP7nBQuOc
389Q8sUMeTmE3bkk0XgfQIpuY4Wt7H+SQjZZuLDjJJOexGB9YAlp/LfscHXh48BkswG2dcW3X/Cr
4UAa6mM1TN2l7nUsp+uBv5JG8d0/jQrAAXhDKo21S0fhBUMwSn+RJozroCBP476Adz4zT+D2M5nQ
+ko5TstddBFg6kpQp7ORalnPh5KVTYE9BOD1HXk3u/FZyPEtVj1vhicuYEdE3pfroOm/K0ugKt5Y
oOjNtsSGTudxGUi56Cb6oCPX2Pqzy9NM/9YEJfTkjDfbn84HELwe6T9buGapNH0XOmgQJWG+ekC7
YvMfAVVTN7OSs6w2ASXCTouJWSNbkUbpc8G/14D/lyluxfMrA9uAgJ/l/XP919h26x6yihTyqcgD
YpsXikr39QD4n2e5PWW+983Ov/vUTYfou8nhIEihYZ9c6aB8m2smcQ9fkqyA58+bgMUQWthn3j2l
092QczH0XsLd2ePWZbJk8/pKOb46ykk+kAZJW1UCNiRHP42Q3ZwGE9l3k7lLO8Vm8mrm2dzCgVz+
81H2SgidWKMCdsLvJayCy9oenF5auda2v3X9aTd9RxMOP7JxJLQpM7zDMfU4CiBJ5EICrIVvBtSf
awuJ1bRTSlGPoQl9VdoLrK29QHNPsiVbN14v548qkYayXNGgtm6IHZQpLLKj/9j++G08ANNOGzFq
Jodg43niFE55lUTXWYe2aRPoC/kbtLQ395bAnnPR3vNK0EdQhUUF/fT9eNQR/OtSYFT6xYvav+jU
4q8KwHwQSepjoDnySpPzUA/IFvxTeo/wkBdFxG65n8fw8FqqlaRBK3leRELYPnJetRosT7Yi/2Qy
lbosmBJzzC51M7rGshGLmFpiU1EykvBBvhOZJ0MdyvbKxFn8AWQfne0qy6AnyiOpJdR0k/RBmYEg
cAwb1AtqxgKOpCsaiGkXxq8XKVE0sdzyUq4It/SeiSzWm5yCAmlRyJaLf721yKrNbImv2UI2jWPm
96sN4ZiRKxo1qWmx8BauMIRPdwy46izA1PaQBJwNv7AA3dp26dUZQJ+9rWEYWENu287qFxSzSTDs
QokT/BUY+BqbSPL+zwUrFJcIQW/3n73Ee2i2l+4KnQgKu5zbCJt74Vqs5BFHFsuRtSJM7ByUkH5T
WyDEQ7IrO+HpWJIGVIo76mpBBBKbhL+SIwr32X1jdl8z8lyRqd9FM3wtsU4/9AXCOjx3DwXyLA25
0BRrM2fDhKTnzGKDJSOAz2o0k1MkeD70C226WgoxUBT1qM9AlDOyAliRMn8Wu6ZdgcXFiao3KiE+
DpTylDO5PQUaggUfwFL8b//x96DvDNoJ3U8i4HZPhC/ayiJJTTrrrjgUyy59U2PKbIuRFF0F+lRE
P7SkU1XUzr2YFiCFLABbQcyPMcsovbPPpz3AEGrZx1TurN7ityJr4so/+bQD2OV+ZwXPRb5O5G5/
Vd0mNi/4GM2pOToJ33fbyFWZx+gEzrXR/xwizas4P2EZD3aoPuy9+t7XlJiIDc48hwoBju85Vsnd
VlicuxkgrlG0x7+rlPYGD7oZ3i/zoRAfy/QDi7GG+gtlZIK6exSTpJi4OC+wwv6/4SeC2sGpjXms
S1a8rALCdkXEwiwwPOyOFf4gdlv7Z32OmYXHfCxSd8Wp+1Zetmqh3J6KTp/htu/P2o+xjlw+mZL9
Ckq7/bBh8cZegSxviETnZcEVGYyFvrn8nMJIsRLZlQOXDVhKcAYHQVvha7t0Vv8pGVetD6AsXJtH
QfY7qJouvLwLe6oYw+Q8arn63L7WBYNUmCa1rVhvycftRgpY69f2oaOJMu3dnr+SywyDjRe6QAaV
vErYOZpKe99bWv6t8GPquo1VIA2r1R7EYjT+KKtmqHAJimN0wHlG0wPPlfALPga8KAtvl0xDLVRD
YPkeeu+iFHCv6fObd4j1d5ZpPb1bwP/8fJA8cfhB2S3T1/UsNqLIdLutaYvEbUsZ8gTtXVsRIZ3B
7qD9GeeRThq0xsz2X2oK0fILbsXugiqnmsumIia5MuAgNsHJAiD4ZaYtn6KMpH0xuY11SLIOIWnN
VuGzBBuSQVh7J5MqL3RwFMIyjoQzOjijAlPxD391Xv34+Kk9pKwm6Ns2uFMBKBQRFM0w/1yNzQZT
ED8K2wfS0OcW8TT8f4wm4xrPA2LP+OSUL/ckUstfubsQ4+w4jn6UIjAYYiy/zMlffHbzXUGgFeIg
nJBNLj9b214uUJPpF4jk93lRe+joq+b9S+5MAH4JpuP97pMoujFwBR4fHrnKhdOtoKZlzhh8nOLO
JLtn6SuTkouJvv2kLrxj0S6HgLor/9l62uNLLEWRb77R3q4EUP4QM12KkFQEYJmcc+SOycIJKdqu
UMBLNRDFoKue4uJdfO2FUpftPMiyIUQJSNaNhdX7Q/0Rk/7RWBQnOA+jgi7G+q2BzEIV3UILVYoq
cpJqdDvOuSzzCT72t/ZtVwk+1EIexNyW5QE4quARIOJgGtX5es6QUdmxVAsGiZak6922YTRghUjz
FN6MYyQCvTvKGPz+Wgn/kwInI7ZZkRP+/ln012JWqXiO6aC2kh87lak9pkXVuIktbw+7e28371I3
gFg3FyL4u32v7uNX5T5Hz0TqzepKJJaeTV5N/+ToNtDXkaaupZaGP8XsgcXd/UvEC/oGY1AgG1bp
HXaY8zVJMSyQh7PvLztgaOrzFxStY+DKxKG7/o51reEKdvYTzhEy/1wYw203x8QDxbv4mI4C8yZm
b4qISKDBrqmKUi4G2qIMi87yypqieXUY5eXcAqsvBefsUr20QCzckb2gv9AnS8I7Y6VyBfYSYzd9
Izs42bAKvGvqt67x3P5ROvZWpSfB4QpWmei5prII6XpEafRPGOy4iKrvs4fQhYAmwg/8RaaObUoS
W/8LaFiRLygHaH0XYFQ3uY9HnSVJQ5JKxYAr1dTdDcUjKG2SqSsebLc8lFgey60cUCE7Y+MV2RYC
w/shJxR4h8SpL8xrrrV2/qU+sV77djfYgHDQZxvtgedE9cpSVmyyYW49YSViQq1lGN4SoPiIfSAX
R7aO+OnhV43NGpLV4s9fIDWlMz8iIvpDLJvAfWBksz8z/IRAa1+oGYmpZI8T7wIKrHpS0Dy33vzx
4WeoBgz72z/Y20fvlNkzNr+K81ISXRZU4nQ0TgMWvyMTPEVyA4Be7qL6HoD1jnpYhS5rM4g+YFNz
GM+NvmzrLY9rgpkoe/cDexVf5m+RUMXwWWIp/Zb26uorw4h1HgAvcP3UGswD4ew3HE/+VSN8kNR0
RHpggVb8Ig3MhomrCUxqnNbvsmRKnzmcP2jIwjgezJezqTnSXZXEP+YzseZ/OAe+AhhrrKJuC+g0
qcjTY3FqVFomlI7xE7vwqo9OcBTS0xu331p1P0gxTFwXie+dRxyKxRfNDMs9luFLQSkxG3E9uxnW
WSA9kOKyEe74o3B/EIzMftSSpUw5twmuy8YO4rcO53dK5KvncDaeKyFvng/vAwgUUva69JjgIEJi
7CcW4yrv/NeML+e7Uhm9yRQoixPMrJV+w9edOWZV0vFH9NKH2TZwDcJp74ukpMA16vQHIbnZ287S
dm9FJPOfKRlM1bofJ6Ugf2wOQohcGPyMQdnx87HJnDupxUnc7Gym1MrA8gRSeyQgwj171T5k5jjQ
uFP1SW9S/SKbVga/e+AFkZgvdOAE3zRyMTUyWOAMI+uqVjSPwPK2BuxdVRp+BlgSwNX7A2PON5Bn
xmWyIUR+bE4TbmBVcJAEaWqCzvtPIyvRWQZnzyO5oUwhkFL8WwflUp0KhK0IOBLauygWfFCHcUoO
p8AyfL9WFbcVxFNQtIpEpsQ8DmIVCHwrtHwWaIsrZz2N8bl3IgVksDF1IiYBExogqBYiYwliNpDM
fh7lolsrW5/M+w+SpR+OFBiGjwqs+vd3duhP6XSjeP9gz4kkwbiztjxfAvn62GJN4I26A7gkutND
7sGdf4Z4K7xyneNa1C5hZ8LnN3ctuD7Xo8JIHMoSwybtcPwbyhf5yv8rJD9wyDXsTI73+YEKIVDY
KwR9nXnJ+3szRyFKIoA7GA6MRGoCxuCW3f9FZuUFeIZyyYE5F6+FID7Zfd78aYdnoFw0CZYJuRuh
2NnY/zbi9VHk98huMOiaSbJsBgFkJMtqWRtSG4ZGVUJQy88N8ezAYpYBJE1FUOFQdn3DzizXRfmf
TPJLjMPWgn2KlGFeeN0qW2Di92NSJzfbKYePdMUGDYHTM7ZGclLI5pnyHCnNoirB9wBq6HzZrjSk
lclJ4Cpq3AnSo65bPpzMDp8/mJljIu6LbwHXx0Vw+KHewNVWlPGMce5bW03PeRtjVvBmSdT1EQxk
7WvMXZ67Xo2FdIJT3nyQJoCl2p4srH6dMttAWw7hLgOWPyhNQQvl88+AVh0xoJ36KjY0hNDjFUPo
VoUM34FfiQDq3hgIdDyX/LpOUBcn9TTWM5GHwNovOasbfUZ6jvSe2XIHzcAxPxYd9TuTrZLpztZh
o1yShkCx4uyx3eQ3ZF/cV6UwUSeTfihUQEOSXsO2f/U91w3mBI+yXREvS7gDg/083DDTEdjaOAff
XHN7aAOY+hqYNGgFWQjBJF3AxTfH1aMhXxA4OwCEXQtJtC7kRt1Rpe2nV9A73Hdelx9Gfe7LcFym
saIjNIS+db70NeoTSEzxj2ZBo4zAd23zgruo8GF2WE2uZQXvzqR8fXmHPunAWiCV2zilpZT2cTjm
s5kYcM16uLdjirE+xvg6O8E8xZKB981Kbty5u7AFyBsrqCbN5M0ygiLqssxRibyro3QRDdpZqQLI
8AIeEEKY0480T7aZauj3nE+9SBXofPFIMrR3Gean6Suknb1GJ8GeVvyLu7CCUQ+O5JXwRut3ijcy
xd9sClqQt1N71LuHDk0c5pNENGoilDmn/3UYXGJoaatSwDLK4NehQDHc3MUs8R3y7euMSJxdDTy2
HaQYUGyhuJDX9/qF9pP9I1HVGXeoCwRXMIw1n7V5RrOkutOPjhdqqmTb06njeMj1Va5VIC7V3bI6
I9hnyw7BZ8pBTQ71YgmfMRHh9w49USzSLijBo4NpUD4iuZ0gqMiGlqpTcSu01/YKNmGhi5Hlw9ad
0HexW1vyTEtDOKjRXuAZpYp91EJpYj72Kx6aTQk3HApkNi7Ll89E3b85N86a2f514lTgQs6YB1+i
3Hj2gMpnxi4WdhRm6n803Q976WyaM2dxNifh7RR8BJTMlyGOLjVDSxqQ5ep7EwF8OeQl1Y7PPCae
d/VZAHRRUiiw4f+3Teo9yLONh4UXxEs4fN+UT0E641H9GbYadDj+c6kHkIUcmo23LLf2bCneYpBU
rqoEsxd34OATGZpk34oAqElymttMeC8Zz536NnKW8S6drGZhHdODbVTHdFEJlZHLqEmUkPfDls3u
xUlcI/tt83AjcHC+72cCbzpH43T+KHp5f0uV9cE3lzUEpUDeFDU9Fa5VEkbXuUDGwqQ3vmd9UIf6
uovRzvlPitGXEhO7e4lHsTlQM1ZnbreCntJa8AmsowcM7PoUniM6IK4vWgTpU/eL3i9pQeIOf5ns
MPbK6kbdi3hdy8YJ/wLVs1AcO3SBVJzxgWbfl4Pva21cHLJTnGLVp0j4RHiXbFDU427QLJ+H+gpY
A4mG9HsTEopDCFQOaZmwMoVJ678BJ7amnu7CVtE9Fzhi5ExZeERq49DfS6DhZ5ZK9cbyTdIBzc83
cK2MujJfatJ5zU084cxbhLuQPzepiEsHP05j4YJxVr6mMF7K+YWMXcZGyZwIhd61FS/0ghdinMUn
BYsewQx149c7M5Cc58o/5QtxQ8CQ4lKBl3ufgmXaiwLDhouRrT2kU+Mg2Ql6NIntG5lsYetvPW6x
O/BCAzbocRcSiSK+l/b5SIs7fTVU4MgHvGDc02z1LYz0jl5FvzjHTTjj/xtgx/Pg1aT7mY0m1XwU
swDkQZbKVfm2TfyYBsChv0nSfcLEEXKfPBGQeLIwJn2s7j5pTxF10Ps+43Zqa/vFKVxCVcNCQbCu
65v0mK1f6TEoVK1Yr6ZacbVWNeOKDSOyagdM7nT6m6G2Octtu1kbQ4QpapVwW+dBmVuhqPl6gIJ2
aZCe1+5zxQJmOXGqMhTQBJX4TSrrOPO+2ZvuQYHeBqnr9khh2+8/EdbXwj65BAe31bgmYGs9tGUi
lXnVK3taiGXl/QSchDTlVmTxRJ7UiH6hshuUdldn8K3SztKs07+2QPRFJAWUg3qO+yEIqJ9e9lmq
YCPSlzKUszyMwZE7v+wjpZs1PlIA/CTGUGvEunnNGL4zKiNtYjBnlGOK6f4IWXzOVGy8gooSvgf6
LTIReXY4Pyq9cjsmthKtq5OxgWkWG7NvEVgE+ZqkLVJmH4svAMKfO6dMxWdltmwHtqwIac89ZwOi
F6dxrERKvNJ/QKQ5VFj1VaMiiR1nb9q8+vXkINLaooFvzseMV+xDXg/Y2qwyBpxg1kcenfpCmDCd
wa8QYoePTAcp4ZVZaj46360QcifEHOQ6SLZin2lAivqmLuonIy0s/ZPK7BWV7r++NolkXay/1sk9
vKwZC6zngVPWkaqdILNvUYtxzsWIp8nNRvEd1293HfwqFQDyUZn0mMDvSjGNlOmHyQnzR1tyxtRk
W92WsFkw3aO71ghV5VSyQ3YThLwy/MmRveHZty+WeshdkYLvGJdKzllNFOBSFOMII/eJeucDXFiJ
sMlFZKdSavCxdmmmp8nDsgxPSuiX4gt2hsEVqXoMGoI4HGDC5/AODK+Gl8KtaK4Oj1RFgZZ8MjvA
eNNNAAACjc6cULIldOYE7eNY/qv5CHexdQ5vcC5L39U3NMTBCg3cUXzL7xZUVoqWrh1gKA2Q8bdb
r6DzdSRBuoVYoRx63hQgiF5knq5GTvEuDAp3q097Lv6mdn5YiScLAgZo4pWDyLLcM4TLVDB6dm64
HTFsGsd+AO/r7BzP8pdLTBImfftDtu+xksG2mOBj8USfuyHd+qHeWTCUP1iIHCXv1SM59fTcjhSr
ay978HJ0el+J/7gWwC+2rrURuqNYmOCiDlAsBOW1RcEd8pYM9SUHZY8z8Y96XAo0jct9YMKiPtzv
NoTDMoKVXwTIeFfF6T0zJv2aYS1w3m/CgwHHEhzc3HqpVDVXDryDGZ/PJ4QnRDLTwbIk2ZiYjRP0
IVqXBrxitxlq5Swmj9KO9gwnuZmVRI76hvCq3OJQ1s9SWnfX5ua3P1v5Ag4VbzGDWrLJeRNYdmIY
SG55RanZ3gqrpM7YftKabdnTEkud8HDm+bkUWjrJBQ4efJ1yUNL3du/a2qKRUgbuEW6jpiyEMEHT
RBEdeLsfDTjCb3Hec/+qmKc0liR+KEIBxdlL++4UrsavdvxEc6IW4NktYsfdGOfuTjgsl9Tm9AvL
ZDWPMfIFroPCRPf3jmEFJKNrIPnf++8A6akmwL06GQvBCSFgmKZfdwDGO1TO7OlHGU5G7lR4iJ0I
vP9vevRJO9UMUv6iwpZZQiE4CdBLWBnCekf6VM1KBpHzGpmxS2A+3zRNWdnECco/dmmIdPsL7JVW
klQn3b/OoTTIT+jW69IGsi5O1uU2vSYWTdOMWGrHxsOOaDN2pJfg3IMpLewXjhI8o4KPf2RVHZ+N
kGD3aRUfzEjiGNZ8q7yTRjtSrT/huZrt/SSEO82QyI0SmQbA0JTZUQN/kbN9XzaNarW9KthvdHiP
1zEZUnIVCrd5qd8VFWOg0fHnazGyFEPHfQsAlOqu7zPNGxvs9+dB8bxT+okj6TnHMz1dzVyRvdbi
YGeU2FLavlpA20snTmRh2RXXmaKnAn7sZ3tS2nK9OsfKmQgSdwxr0HJmRoSCiH1p4TqFGFyL+vgK
YcbSjkhft15JFaGg6xsUBJ0Wkkythhi09xv0XNly8SDniz7zpTqEBfLmTvKfguH5t9WIP4E9QRaJ
Nh2Jpj/GEMfNh8vkOvMREcgAw914fmR1jCYKSNGI7uwoAhs58UehAuhHvIXzMJxqXIvyjWuAZPM4
qK9pLhd2nnpHptE17NdJGXjapKI3YxrX6ON15qHPsJNfAcTH0PkVz0y7lT0v3Vi4S8bzyVWO/Twu
Ftwhkxr+FHv6fVfxttqU3Pl2ZCktLWRwwXApzwoIGBOHmRiNLYgBSXyeukpRrkgebKXousYg9y/2
ZZe0E8bdy8PcuHnhg5mMKfJE4lALdcGvXOSIbT/zk1FH8HIWKhDqw6ftWKASIeKk6PuyC7MgdigD
4MfO3ciWsEiKYjQE/EqygeWhAiw8fCth0HBggQ9CGpY2BH73W8GgiyrRjCzyvDTnQQyO1FZ9a/nn
DNFuzYmgWJ8atE9AJH6V61ECmgfUWuhO0DqBlG+8ZiDxNDAq/4GVfei22FaFuWkuPOkv/WhiMfih
t+NIJ50aOZJfdIsVKavFiAGj84e+l+Yfhu+Wauaf95q77A+tLrhxsbZxQTwo30PDyiD3LC9xJtPQ
1NmJ+i4hK/6wjOAVc6Oi6uEVNg6EnqrVii9O16uoaCNHJKPxaP/jrREpGcqyr3ovLDuLtuHRGXBk
0syIkCaafznj6/g35uQIBSikNSsWll6uQ3/AVjZsYvrdAprM0HQefLdBFQ4szMgZRcdY/tbXaWNn
yg3FgzGv1p4h9wii3TRUWiP6VZt8/64G3IKhUE2Rv99+TX99bV1rFQuESbVRm0M0V0OZ2hhmdlXW
qBkhVJydweHt/T5oO4zWuKe3bcxE0X5rVo8l4emgNb64EnY5Jsz04guHTNY+vBSyK5T1uRQC0yLm
bZ83m1qErIKVB/Z+4vyqKy+59VYtrhzAaRiDvf6NI7pCJslqfPksfoEvpypz+1xCUdQI/XxIla97
nLAyfpkX6xIaHZXbWV8l0FGhGZwQKPP0IIno8dlSs06Y4lGJgT7eq8X7Is3k+7nROTZlPwMJgXuJ
HrIZ/gjR36uZAD1tgmmM30Lt11VGFe6iokr0DvQwaNfa6R8HRDrR35HQiEPBj78Bcr2GU4ZVBfgb
FxzqGU6Oc19Zlvhnrk0O9hfEQIDqy2QanFfbdzSSER88gI6IT0z87nvaIBpO09Y1HNq0gKMgHyLW
Am8666/DxHJlLAVk+MT352emTPTAfJnaxgOOo69EE4ZtdGqwZNWfH7hgan9EFdluWSDV8uj233/b
t2DgQ+7D4HXw2jcYRC8aUDWu3bysFZffcDEyYr56HCbzV7yMbZR7Fcks69KEK6BEqWMPhuNmVJQT
dpiPEJGq+Ul6jUb2gVIfh6kjxGy1EMxiFgc8mDgHbKXHUim+8bpgceWLRGzMb4PiNUpZJ2rNCBvi
U3IK04noZIxLVXA4BRdxFoO/1BoQAevHMVgTgjV1ZfA8c/uC+aJgpW+oFi+4lpNqrIFRJ503b9MK
TMoKQ18VIv80ZjBsR5+PpgqY5+KRsPhi7s1wGL0JN7QWPEzmzb16MOTbTQHmMtQSx3lq6DkKwrev
698nIqfx0ht6dImTydExgIHl2r6JIJrxzW1PCDegNSjAHSAlQKf5HsbUhlDD9GW8PjphuEvyh578
lyzAmZvduRXLZYYyyqVUt1YvIWzDq0+65hFBWF8qNqQJN+iXgOdHmvXB93SRpCetaYvUm86rdnOe
c5eKPr9V+TVTo6qkJWaeQiTbQlh5JITq5mxAl8OSc4j+qhhppQRobAvil9nVcFpD6e6/qccZfUZj
QS75ZZ5VR7YsMyd+STSXnej8ARXJ7/THeaLBTAd9/jbi47R1Qc/x/5EDl1c1rdNm9rfMji331Fxw
FuNEmu2AoGuUwN1xUxEZ9PrOEBXf9v7l/Orb6tpSNSf0/Cz8DtH+LKMycZqszBjcS7ZOTyKGariD
wT2yE+cfATy74ekFKPBDiJrzLR8eOm7y9EZdSJyQW7RiG+gcTPaWtccJCOtzIU+yMKL86DQ35pEA
dPKq6DzF6fU/SHnXJH0ULIdshHNqQZ0aeq52//2/vYk0DR1phnzPs+5bV2FoyeLX7XayAJboK3eI
WpJoKECdfxMj3v4lPRq9oQluwbfLRI45XS07jjXWeH3QZnFCGtcQ1JUjKX572tKuxrCccUN39o8V
wkcOhhmilnbwwKAOT2/XuiMOtbidqOXRF25w5YZ0povm2V1gvXuT80FGphHgzzYac4fyZpvwve9k
/4WyHF8zfewuolrSpGHy6me8HPDQGptDDvLIXGG9t6HX8wqLFx9tFZK5StFptczS9yBOGCr/BHRN
yMbrUH6DMJy914YJeZ3nroP8XdHfk1sdcPeShxmMnIUlKU/GQlDwms6xn/9T4aU8angLUBwXNFRP
jCX86MW4sfQTxCTDPFhmPRNtMWFfGJmu4jbYVi2Moux0lvVRfEM1m0Eyt88PuBsxT2yar0sNTxr2
+JTUDx9rdeIgoxvHWufk0KN2ZomafITPaRwLmO+SgA1ojGmY+RVvC34obwVE6iG/d6hwjP5K8FUM
1So+lBFeu6pbm3QQ47xgDtA/dQHOfLjm9aKiStqaGyhfZr8FvHuxhpzEN96WlpPNVcLkGsmJjRHo
sSWk9sE2jwuQytpaRJE3WcSuH7DKxqELhf1KBuIWD7gLYSI5L9Nh0KQRPpqsZAmVW+eYTAAgFbb+
ZR6sW1mlwNiFDqDHmkKPCqJWPuRlZVnfPpEvP/KAC6FMSGUXAH7flJYksjl48T8ju5/Uan4tWQBG
5NWMGsLNwgnTMC1PWtCGpVtfh0I9LlgrQsNikywXj70qgSSD45D0bl4/rJhBQ6uWSBjNHpZe7Zjw
Xoc6A7EPUYokqOJJTfuRCjnQMpuJ6GRPrQ/BtS9P30uY4YjlUNcRViwfAdpyLTg0l6vl57h88rR2
W7wugm0MnW6jCnkbISPcr1VF94WlMotEjYWbPnF8lnXg8koNPujV4dntnw08CwVkxSAfDjQrQUG/
qV2q36eIHRgA5tS4svrfsftemUnhxqfezQwuQxkP1uJUHY4K/qxvOSnodVx6085uJ5ceB/NgbxwX
nYbphR4dW6fQ3FKnouTXZZBtbyU3B1Y5wD/gplUkyPwCiFrYxm1ZFNesLYm8dqs7KJ8SeLsV5EZf
eWW6hIga3IgsGWFjUO/igZcRBLFuddEJb0p18uSzFK5RDgx5qun3nNiP7ddl/7Oc+xULKDC/hoBZ
9YoJeuTE563rfk0tVuQzg9a9sJFVhWOMzZ2v3zF5ATAe20J88/LBIvjdom2qayK175YUjp/ibLE/
ETUafaLh8kRrmOq+eASTAF07/GJY+pNZgYc92ldMbPUl9hzLtoLMGSzCsjmSscds85/6nMk+k6MQ
t1xz/iVWzYrA9/7O2FL5xrWUYr8gZwSbfCB0nASnBi29sQLyCQ8tXlIwpTPkleLLaFdYdfZ4fduF
di7JIyOef0SmcbLV+DoCjoQQJVuSHMyCyqvnM66dPDf2mBHgD3WCXpS4S5+m0UqAJwkcmlN3ab3a
pOsICclUCFhIDGuc0qV51kLtZlQvxQt85uM5CFeqo7nqcJ1TQ+uGE5DVdbaXLTfV7Iazi6B4Wm16
w/z0zgrjceCZRYrWdq/DJSUQbkY5FP5Zt8Uyx9vnpKaamtiIMf7qZoc4aNKTwdVFJwnk3LloW8Hf
ysNlS6zEx2fJmG+Z4n3+nETEAXD4Zdh1AoQs/Fhu86l6gmhjNaCY6JxMaYKcVB0UrR0/P59EqxRD
3adKY+8kZXya2BeoTlorC986nokssuL/vKM/QG3FDoPSjm8NZynsOIBrIcOGoBJKt3TG1KDkXRDU
oGvjRcoQSlAn/4FeYH20SrQVtgbeTjmLH55o0d86eyyEh9quryKzBd795l0Uw7+QmxIiAswAQCs6
Ml0B6NlTdsJDIfBkfhFi6rlOVUBV6xv7aKfNCJbS+hgyUSE+0tni1nkRBWRrL/F5v8JZHXIA8xUx
4XZW7Ow5TFh4YalM6ZOpjZMUc6/j4Uj8uWmdAfHgzN2C04HK3Yx1Ipz6dZMhILipWk4IxdL8ghT0
EyIdsLwpeXYXyyB4qHa1aXPk+GBkmSOfuoWM12f5ya2wb9CMvbMhMdaQyB3sAcVCwm/jaCHCeiny
VnRDVyljI0dpVgvmvi0nD7d2N1EiktfBkKRX9/iVQ2Qz5l23C6/YA4qjf8+Ngk5kjF7Acn7+RonQ
tYW5FTy7GtriW++fqCA3CPzK7fqFMbPYJAQaDWOMNW8BzJXSNv+bV/PFqIxo0AnOoGUm6nvvTiQv
j9ozkB/8/+Ll6+Hsmr/lqE8c7TNa7H893HNw8E+U9u4915CF3livIxPgguWWv36oCxVnAqGfkQL/
/+phYYwLBMzd52Sc2c/A25PvoG7QrsVGB3KsF8v8NQQPHoHPm936twRy/XoXnsP//Dq6xfAsSiMh
NEzL3AI6HurD3WPpTtA3xlC/Sd9VnSq6p4ILX5JsKVmW3Jk6+U36oKRgPpuvZTJ35sBVdACmfZVO
Js1Gnk5+w82Lo0uTcv/RAzLBwx7AQ96Ekow54TJv2o7FyQngmxhMqeId4SbiXjz1KoTfDhReNt7r
qtTwF92aeGD0T7+A1q1TqcgQ7Q+e7bVtM9EgKYusXTHbschBX+AqRxxzUfif6Ud+Z1HpnpkMLiNt
ru/Cga9vsgkcyoPW/UNfwSkxbFsIxyt+OGSL8YcLZpz57jv5w5QA/AQiY6VtGmswNYC0BRYe4h8l
iYnBU0WWDzIOK/IQAeVtYOwxIXXEcQb315DngUhdW4Z38p5HCkFEFIgWSChHTYGLpH+tdzSA/2jA
Oueb1fULJFBpo2zZIBP3aAqBvleEWP4xhoT7Z+Vy7pTwC6QDmuYC0hk3IHuWWccT4eVV9dVWO01G
F3IzpPWdH9YrK6whv4mi/AzpxxyEee4t9xt+u9qaxESf/FPmmNjsewaP7EOb/8HQTtPQT3ENM5JJ
myLz2IoA49FatqeJSnvLlmV9JDRAEd7GK82737h1gFr4sw9KEtwfosxSarmfI6t44tpxka1XB0J8
eb5mvyTydtrzQDsMNs50x97qN3+lBR0SVkxVbNuQQyZjIApwrqCkYUOg189UwgROGFKaNg6OPw4s
PGZOLC5Tty/2uYYhCsi8ZXUMdhf0IyArVTVMcoFyIY4Q2N8DxxqT+RW65e5hdO7PKHZi/QFWj7JN
SwyNpZN/ED3DqUeKcVg9rJaTLgz4YxRJ/rGb7tCiHCkbv9QtQn9A81fCESb7ioJZ4kReLwx/4OgY
RUbk0UbBZOawr5iWojaNIHv29WwCceIJApZ2o4vutYMytBhTNot4cc21AIpbzHFGb0S9kO6d0dEd
jgoSO1j6kwg5pLZyEwYWQm5aYu4iBef4lwu5q+/GDJZn5pPkjNS6/fZQaazHGrCxQWt/UidRDywl
UJc/GejpmMRBZ47otU6cogOk351wKwMguvTXEUP+a/w42eSp953ob86QZ/BzLXxH0Z+3Y+TOUAI3
ltBAIu3LCVbPIzU4iZbR67IiFQXyD91F/nyy6/w8CkqH/2WNnhFG7uhSgBEY7ISexqnsPFFdIEDV
uKty+OVl547+O5DUwKwt5i77iak1sQWL7wn+Ci/2a2H58w/Zb+YNvzm2XuDa/I/rhzYEC4CitgTj
hSpSiEtYgl2gUcaNr06m6XXPhHvRwEgGZUXyZaVu1lnZNefhvNO1s4t2OTEBroYjWPE9AVoZ8C5I
4W0+JCmB2NSRVetxDVbTJs+IDsJwsQb4xjGWcRyPOrzfyb7BLmYAnpfDqtneZwRP2sYST5RWbqbX
Bq8RL6WlvxZJArdOnJQk4defO4fmL3SBE5yRQJB+3fW2LuvFDljrCkV8kdA2bNBt9YvF/lIkRG3Z
KeCq4zAgcpvLk//hoY4TOpXRa7QpGLqs0+HJmVsP9boFEiNI1YCbkwEiU7+ofXq3XiirnDQDnuym
Bl+vBnRDp/ILuORwR3BslrlodhpgPrq70ZFr0ZwRG/zRZf9XRSIDJSft0zcQjdNp4pu/nCMr+wCY
s55NIxbbLfT2M7ivDCTmANyhWk5jz0wjMr6yYrDSFLii1AAGntuy80F0hpPJSUOeO3DTvw88DNZ+
SxSgf+iL06BJD0LukPDei9o5+y+GjPptoV90YXT879YNxtm2sNAJ9nIKrPc6iq2ATaSMQuQq6dC2
7rk5inABrWx5uQErkSpKyHPjgjmzOXvQEYxj3AjlOJzKaGPiuawxTin1duDgjJaaOZYmK5ws7BQf
y65Lzqaqsg76j4Bw03YKuOPyKrd59bm1lP96klFEYmIoL9Lre8a+FHDVsDj1K1mY6vKdMBENxvx4
F0TCPK4n65x2OdIdljiGbRmqRw9Dc/SHa7iLy7RfpXB5B0/KqM3lQARMFvYu9AHDme+FgTp+gTGD
QWB0CZc9ljSZqyfBjBJB1ukaVRNsYwIBJdBTFy+tobHAXayOyEm4S0cMNpKQ6ZuwtZM79iOTZjVs
0SyBGl85mlhr0uAwmfIYYYMyspTxNgFJn0J/MBsGSQM98tnwRkFwXRPxqbaQ6JK+psTIWvE5Zs0L
k9We29KuH46U79iabbkWb/L89dECU6bcE0rKjLfaVLnrEwc+mBMNDe87H57tOl11HZTSpSAszMDm
Bu1MB1cRTW49R2tVSqyH05PyOLW5I6FuV3uy9zmBZC7jMNPgQ7AHvt1Yr4gvwF8IKNzC9+rGX4La
wlyfc0fFblRluHiIC68ACXwPIFZjoRlR17TDl6BlW1H92tdY80kBDQ8GuZFTZRkE7XfPFA2ZtdPQ
DuCeGfDBZN7+sYmLnqf/EI0/fYn8GHOZC7Z4xJ6VHLpZkzKpcTkxaDsPWt+LmryqRZgEg7EtGp3t
J0mRcgLP1PmXbwXUtC30BJL2KF1OgmAJx2QF3m+vFuGa/XQdmzxrOJ5TRSdauGM/JtmRI6Q2fPzg
r/xPpSvOvAoJe4fv5fiR4m8J1SW7mRDu6Vt1NdR3gMIGwwZ+DEtyFRG9hgSkwbPTAc1gJfRvR3jR
Ch7wzc/bYcBjnyrWLl04kKcOWwmZUe23xLaZFohEUPtwSbTgZ06ZmNbvd8IZqC1+DCc9FF7Jagzz
wpMQyBzS7/ymfxFmkUZV25gfmn9VKv4AmemqWwel2f8GOBvIgcG9MwBtw7Ey3Kazcm90xRglUwji
yjr9OrvgXQFK7oOAu+02fiGf0MjkrMYRAt4KJx/UcQtljD5AnJOXekhta9RP3RmbTbrzlsxFPO9h
/6Hz/yIn6kcZe1WF+8uQd+pUUiUVqlz7F9dKekaAj3KmQddp9Z8OibCt+4+CIzX1E8rbswOQY2pJ
w/p/WBYgTgQmBApXsYDb2Vlwnxd3ynLEpk/6nqXM8cdI6jZXBRE1vaENE2ehF6C4E4DdeEFKiJsB
42SXfvYnbMkzhpm3AbUfmz3a0Z+kyMY+iL8T/nMIifpmZ1bG1O/ggVf4RSK03IXSAeia0pMJxLva
jS9KoaUwGVaAyZvwQ2Lq1xCmtsidmCkZ4w/zJjdbOyGvWUAXsnz5b960TIEKMxCx3fKHqmuTCkXh
3ofmed/0AbZiT5H76J/kkSakr0RV6sRb3TkxnI8bZxpT6z1NE7oncsDND/WFDx4zCFKkw+OoGenx
zDmJJ4myKJrJOxDcjvg0GNtGv1B86j0phpTF/t405Xkny65cyKaMXWrRz9wOqLAvCS65MgthHP/+
RPPujV5m0JoxcDswrmOP2dPZZEdSm2gTpSzfcQ2XL1RFe1olRiUfH2L/n/66/tRefBsWKrS85QR5
Em8N8eoqIEpgOctGdzX7AwnJToeLsnCCKqJ/rv7PYuMMZaLB6YbCsOozgOiReiIV7U2jMV7DEMcT
7MHRi+cBnzDvSuo/m4SLYivtzZ9wEKUdfMwmSlZcTAEZkBm+g/XtzOcukp+aOmWmJ53G1I3pXYDO
hewtfDNcWQ7iaT+O2YF4lNLFyIwgy8edVaAOl2cJVbZk9woOtnhC9IX0/zQ8Uf6meI0Lhfloixkg
1VPIK0kTRiDDtLIc97qD1rmFtu0Pyd843cuqN+V/CLsdRNLN1ATmRVo5NFtEvlxtq/Y+NaY70RTj
gyA49+7PRFtwPrfuXZuJA+NOSmV58/nj5n7m/nvQZZoV9XiDnD4c1z2UU8ryXU766tdHS0ZeSl0y
Z0YC8pjqlw6/Z7MWwKHkOue7fM+mfQl99XpsSu6Rvya6VRUgDiolKM9m2E81MXRUkUTOBA1qRfQq
EOINDt5ZW9yhqNO9JUutBBO/sn/pIGuDsfAg1cru+gVsyuL6jR0KLSFWFGFEjgooZIElFepyJO46
KCi7CbH7q6kWYDr+5S7zM5BoecPbvHJY2ddZ+aGCCJDHWfimgYki9mtxqBD4e2RE/TY+Tx9Alnpe
LTn8q/IC0l8m1sXTiFXm0vhuIMZ3Dnsocs3abKbUgdC1UYxyJj9uxPatrFLCeRDbYKrLv2uRAOsB
dEC83jGlSEZeBML0PM6Kipv0UyXNOO+9dtyJtp48ME4uO9oz5iD0ZOwn0Ioo6jJRTHIMH+sg1uXJ
czf6BJyLGjzGsvhjCVE0pER9OXu3UOdkIVp8pIn0S6IezxS0h1lawtyunxv7jn/F5slB/0/IXMUz
894KxiId1goP2QEFxF48rdUvWAtk2VqzQH1UI89E7+UquwGPNYv3CNvm1sL0PkOtba8gTZEqOGPS
pifSQkOKB/8dGP6SP5sLCkvylOUbKMOS5Lliwe0h+Uah7EYDldZVhNOnAitGZFxk/i16ePjGZRQC
fsIj/f8wB3qd8H1/yBYAojCQDlsD1MCo0XVa84uWmucHWQLQQquVxrSx83vR2dRHua0DxKC3EGtQ
rntEG9sUKZ8J2iB5iznpFhz6+hmhqs133H5f1zGvYbXzhWpHwySGAF8Ym/PnX5Y6wijtWS5e2t1N
hPSL+YLj/gbJ1Q8XuddTne8bVZnBjvvwS/hhcN5hi7whvh2n4nUkhmG1uRHM64BTIMLxLtp0E16L
dVEEb0g7/jQ4R+yYwEkJb4yWkg0GY0BjR4w3m73pjWJRKZeidLeZXDo1vaxNnSp1t59c4KMTjJc0
QDaQqAiieLEVfLnMcDYHlh2rdhPLmhShCD3aYDHjJdgL6CseTN95WXH/rsc84284QFtqn0yrftNc
nqI3E141C41MqtqLD+I48RH+xggOWrCnFy7h63JWQk4wdNXLqVz/4a4ByBeF2g2O+TlFjkvnVwJa
c8dBzrYWdVO3J/B+FuJpNqEQZ+HxUpz8y+qSUv91dwLAmtPcGflTub4jpRzqZdwYldgymc5YKxXh
t26HaqqZd3GBGZG1CSI9UGDrvoJ7T/fg21DiLIv2zMUSXRO1+Z217X0bfrlqsC/zvRiMEI+IFXLn
iGnE5yaJlCJ25qB0ULPMdwDqxWHsVM0fW1bG99GAz4bss5wXb++EaC+sQ/W3JANHpCrixu+FCzrv
51C2mqU+j2znZzITmQ1UHCPsAQcTzkekGI2YAZY5x20rH1Mz7ZiehAunYEWAaz3tRbppcLuwqB7j
1zYGvQkA3E5mKbA/3DdvpZuOLW9KjTKueOiTbfvBMSYS9YhtqbKq3Cc+JK66u2wx8iQJBWkwE+Uv
3wf765mURiObF81sQTAMB9736kY+dTseI7TBn++sIKhq3N0Ty5fBCnUqkVog+BVRn9uqnkUEss5W
vqo3McO9Icns3VzV1bk35X/IMQNjpPqwHHC7tdU+nk5MaefuUPoMEbcVjpEy89AzhvsjtEj45BuM
gWiizTY1wX8eAfmtbjJXW+ypMKt/1T6zAQBuZgCorUqPPpsp0QYzArj5odQAktA6WJOCP+HkkSXh
Wuuxcb4P5oB89XptmlFI6xRmaGBr2QQWcXjGOVL7aVgEeNhCSkp30ueLUGHtbtgbXLPgy/XO2TeH
/0QBQO7mxkOlRQI+qy2KdeLSE4w4QbIpOT9eUelQGXhqfbD8CZmHlftOP8LhzF28AsQlUUFhKpSM
nq99psvvuTp/260bmglQsDxaNDOBW7J0ztZaVh939k/AD2XD3PuKNMhVgUbdqz768MWJVmJcjazf
ggEUFXkT5v1JCzCFhkR/8590bHCqxAhv5ja6bZWQYSfHD+wAZ+FnwEcWrl1uhLIfVu+kGHHLJBrR
Lot5DpbunS+SNxe7kDIDfWGkj7/lNgq6vm9aAyzvyM6npbb+8/tIJ9iRvbCJmzcnxu9mwkZ+KFzJ
X90dC51/bbq4uS4q748tKXnz4GLnGJg4aNnITfGz8CuQllBmZG/WDhCAbZ9wyMGshZ22RLxtAS8h
h5gKrJZum3rLwmEUpLK9VquKhVLNMBQIS1gUAhmsqWy6DMf4oRO7GsroF09+JNuS8JpMr8J2cM+u
16iBvir5QR3sPMeeNu5+aF+/nNu5pEUa8H5Vw6IqwO7I/hclrxu4cpYah7Ol3gXCm6XL0T/ER3qn
3kI69ht3R1McmXIJoVJgNtJxFK3NWHlqCxrwjZkPY+HEo8Kjoxpdv2E3po3G+Hs5fwcHf6oRAIEG
e+BLJJAA5UAj3oHJO0qvEDkG+yjHnWzvJs/iBX3UXwdgqqnq7tsV/8m1dze+D5iCvpofl/lEGTzi
HCApnNh4B1UPeXK/HlhS/lS7uy1KQ38KVqnCKKqG/qX6iOSfbmT61mV4NCsbvs/y2DKaYev1cuRA
9DdpV1JDuDzw8jR505UzAsOiiX3x1GhdOLEDAQf0kIqiSnQ3TN7NPkiTLUEqkkNz5mIAh3idgyRi
LRDi08JMW6pNXKKACHRUnFsKpAqvZE3DXkvbFYl/o43Tzes26z+boBYYVG8hYnP3rEr1u4CRPhnT
YgLQ6g0e67ZE+84cz97SS60z5FDKVUD15Qtmi8DkgG4bc0wJn6VeRXg17f8Qzgz5kdb6Fcwgst6m
rrybCeqZ0S9Pc/lzvOsLkDKOjY64/c/PgVRr5haMtaVLap6UQwsRcriZkE45W/6thIwqm4sXdbx5
VAIw95Xl8n17WHGk6UJu/x+qklk5HhBS5UhtwtHba3fxrL69MgcuYPoTbdfRJeBquLyZm2IhaiO9
imbAABoV59LcYAMlhg6smtgx7Iah+qnY1hEP4KV6vZC5FW4X3IoCmWIaVmEBJXACSPKJNXep4mYk
pPQ8GMiaJ+NFy5HRPKjVFB4u8M32eKgmOrteYccQwPa4lKsYKo7jGTiemwoVtLOI3OswY74QQWBe
q3IwhWjMJAvMfOQ76hN6gaWDeOW7QyUFmtQfv52Abe9Ks3bfN1wk/T80IaPOJ5RHONYAkq2YPFx4
MyfQUgS80RsNhSAnat5FDeRncLOTMMmRA2q8fIcKqDS5qnePDjhpr8ItkLzOuIqqDjD+v5/bqEXU
Uw8RetXV9aucY/gKWTPmtjOSIMOPp3ruPvxyyBIyIUw5225qMzOCiIRsAcvRAM8HS7u0O2v5MldC
Mt9GGvfiNtP/kFuEcUJXf9tFDiCsLeqIM71nYw1cPmuxmyYW82dV/60QCQvUzzd+Dvnv+hVGQMAF
TG+i8p+pnXzSY9OgDaTQ12jSQ9OG1uGO+2huhGJRSEvTHHFDKxpKvML4cSRbTku4Wxq4Y7a78OLt
ta/PmTQZcMZm9CdmQJ0IHyEGdjzofGpXCZLvMHeCCXpuCyuIegL0swxezI4dE7qDQRSYHjUCQHvl
IuIUh/dTuYtWWKUBn4T34XOdM9Ezy88pKrPHKcRxPuZhmCILP5GRBwaF+t+nlv3MRK7mC91Twu9W
2Q9WiP73agdi0F4ZtdDpUl4eQayYwmHrsjEZFEnkScBfP0EZiwP7mT1zW1zaWw73FPoFqmHgmLPS
fMtGfOdbN2PV35YicSz9/Tzny8OEuRQMaFKBUmHfGqFSb9/yNLveVkoYu8rOU4X1WvkEPxsoJ24j
1pcQX9kl/VnfgFbbkitBpltSYQ6DX5k1b3q7LsXg9P199Ff3fYmFqawJ196wfe4/8oe2kjfBJPPv
1DEU4GUax9IcTw1x9yBnfdaTz/g9fikAQ4LUpQMzhE+jNv5TbkZt+pPo31IG8s2GP/xCpOfxlkBL
qEFWHqvTHB++ksRoF7Xt3yaIs7f46z87CINLZNGs9VQnM8AKO7vAuuXKwb4+qBvZ1vVo2yBwQweQ
EZT2hf+a7YjiT9oi4pauxF35D4moVEFpYnU1Qdt6NXDbgmsJ5PCeE+6Datxpf8KLL0Tg2p/hSg0Z
UjqPvsTtPCpad8T8XHj8UZuY1SBlxOXZC5cQknMYEBA+gzLJmUAqJbl5vKYTNIjFIl3uAJ4iWSdz
+HxuXXu4GwJyuIl55yGy/x3dBCX8/vTwe3Rn4yfz7OuuRdKtUWS7O+7Rg7QMxGNF9bxW0UvEZheB
uN33PG2O+CNs68B1aHPGa6wpMuzMQFVzSRGpMB/V5DbTZNprJ2z3E8IBlpIsQergJVNWSLHo1mF2
iH+6cN558F+dQhwkoKDMUyBElumbFRBli2txHmt7kshpgpp9c8lNSC5YFbQY44ufn5V/SGRgHn1o
X8YoNEjmOn3VM4AZCeWD48qdFJypiso+gCmfeRLcX93VO6ZA/KQaQq7jd/s2r3tpWxh0grb//KfT
tYYdW83/iUrfpjUfzwh5kVB5au6g8sGoQyHknoho8jW8p1tes8i9V4uLpO4uaQUHuM5AwAjcc0iS
CfeXzPsidDcZUULwXKEUx89r6VI7QwGpMf3WNLcvZ+Pjq+rr6CHcCEVQa8dZ2f3H+IosLgXWUEsN
v/iphm3FpksaZCQSc36iZwCxg/kgJIX+XH1wo4i9f4UjGs7LD4NuhtAhg6wvQYHfwnnm9et9Q2mI
dl4BSoJ0lkSQWa+IaUdKAjS7PZKpIdXp73yXaKHcOwE8G/kOub9HP5wXfkV+FLhfHGxsjAqKdhAT
Zq9f76fc/3Ed7lQsqaVik2ZfyQmIY7yJr2aIcjx1aSzclKDMJmHhhcWVXGGqwQmue8sArIF8ThTp
WG8+S/TxoONIJINvAu4G0Cn84BhZNkriVfOFyYrEVG8OwK3+w5379jeAZObl90aH2QOsdmV5ka5i
zzR/3VMJKfvOQVrBD67RHlFX7XMWZ5GrUNJyvySDZ9dnY+djwKl1dCENMt3gPldQtNxBvD77EEa0
i8GhULaOgHWe6Ke6E6HUaLG4W3frp5CeBOfAJ47OMIQ3nbR7ErsFKDKV1WRE9MpRPR5DLMdMvmzS
IQvJ9lHTvZfhRCdRbmJoiUF6AxL0MIoGLLoOGOosUhPjY7fj7HFVNJdeGZG0qtj0Lh/ao4bdsExz
CkbzYOLIz23nA+gkJ7N1QnGUhv3dERyB7EItEN3HAHD2u/T/XYYEIAmrXqfsv8T39WDlmVcAiUkH
GQ2utVtYVCOyezxEq187nzZCngQlcNC3nmRT/fdGTm22+KBKmB8vwDaPxZliEMZjOAo08YHVkFi9
vpxp1eOtp2fZtQAVMflFGnoaxXp/TKkznt9al0HbAwxtnb3RLk0CggM9j3McZY/kLnJpIYV+yLBQ
vY/bbGI8/sAt6Is0AAE2sIU4TdihiFBfzbnmxjOp0erhd4YTWIXrpYAqDNdnQCr0uEhk/gdW6xf5
1a+Re4yBI4Khv2xEq0AqR0edbAlhrE3yFEZoRVuJgQ19yFLvWGvZo118nzbe1KM/FYSHpd/bj+2X
sMP+AOXcCKJ+l+N9KxeMHjxND57DaAfpdqNuRyhYjiwxfKI5rBaFPSbqUU9W9tP9M0d3TlEw+SG7
NGjZ++GRCcXYlhpdg6y0AQxF0QUKblhxki/HsDaD9ovr2e/ZBZWpW4D/Akrw2LroT2UvLGCxiav0
4qx6Nx1vyIcijyoGqaTmfbe7n6R8258zvf5WQfhc0v2f/nlb3zharOCf3DrHEZzJacS6J+hwKj/z
JSQiwId7YGEutMKFnUevFJW/uyBH0M86WEcgDKnQcAn4yKcmJUoemmm7kQI32sPuuoS08YDTqxQC
ZytP+7Mcz6qFzb/7rOCKruvmCIvcV62eRi2BPrp7lfctrqhJqadV2g/fbFA0quvZdQIzYOqug+xZ
elatc3/8vGBncvxJWB0w+xyabNKnJcB3bg/FBheUe3/DJLqDDg9jX0O3Qw3ouUfY27+uVZIFtGyo
yyoIpsDpZNxmLr1idjzA2P0gtObGHLTNnIjj9SFCWypPfjBmpbKTnn8cN7am67mUbV1jMbOUwr3O
rcxjSUCgLrP04o8MEusVfvsUtA2byGhozFmG/Uqj+vxSoQltdCtrPgZfSQmyOZKnPCjj61XzJX4M
daHRaX//CWX7oQ7eYxCgV36hNfxznjFWvGgGjjl0Uc1k0gJuxzyt1sJzPw8u1sFbaeyFggzcvFIu
klvjj1jj1AeZHTepQk2wqGfV6Pdzdf1+txt/SqGMQvMVPaxrX3VqBKrKRlJvQuQNE3poJIDBpplG
CalOkAkyXsycvlCvLqNJ8AvNEkNG1uipVSAOSZ+IIRkBKbBFMFJldJo9ywHRGGYiCEJ8lGBm5rjK
N2xMy3QjQJAvdkUurvsfe3f1ZgFitGDgEbihe4t9N+uGI0SITKT1OsA3FNwQN2frqwUyOAd73hWQ
mqmNJe2lPs2wM46CZAughmNYEZ0c6d6GzboUEGpTV+TAm0K4Cb9RoMDI9AMR9c2SKWB8in9jFcgY
3WZoxGcX3v54loWC0qKfR0lLbFLVS3rYiEjUBl4Z4thvS6Mwd9XwfnH46GmXLCyVX44o9/EOj1Ej
YQRWPOfGzrqLknArE1d/2bxBBZyMwwjM04C8OiePzkjp87g03vEvS4XVDz8N4M0nmdz173u7DHqF
cSMqzkzHhqqU1PqUOijuta4pjnB/l5jalnoJxyBj8vU7zhCwda3oQz+jnYkMp7Huz1GPuWDE/JCL
/euJgKCSVUcBBneLfCMM3XUeH+/nbbZJYxDfaklZ9KGvr/q7zsbXxRuJ2YYk/cxOFnsI3o33ANeG
eEXHHpQhnCcC/rdh4Pmjfzl2cmjyjFQEadGyr2AHk8c9Vfxlv45uA13AN9oyVLvgFxvy/J7dgeBi
w9RhVQwNJ4EP1FxtHjHrdCghVLjDHgEWowajbOqyBcRXSZukhDZpOfNqFsTgqYuN/Acy39c2Y6bV
dMBI1jcY85SVac1iKjMkVodcaMtUOGpbhk/HUpCWBUOesa/Hy76OVcI/TBJdn32wzR1AMdlenTbM
UXll2rYflpXqkQ7oDs6E5hhQbYgbxAs0+6hK323FHJ97B25rPfenRoCMgyyggpywRZoTD07/X+0m
GSbhEAOhjXPRwWDONiv+AxjberoNidg7PxOP7B1RkK7WUfVwBFydqc1+C+VxeAHZesYwkW+bunOH
pQfnSDj4KMcCvum7PF0IUzR/18fyI4E3QPe+a3D36cHb/OywYfmPq4IC4eM+SgrjqbaGYAe4cy0x
747IMWrfAfkjiFPJFkdl/S3e9AQKFJTM0msogMgdUB6ChciEMEg0BRW2FT83C9QHPg23mMSh6+OE
7/eyKCeJtrchiPY2HXr9K5dCrpJzFbaMVWYU8dZ5jJJWowWJBnQ1aYuv77ooyUwt2VKqP0ewZsZw
e0nGdQCHaYCexVXyOZ3iJWYypYqvIKbWlYN5NcX0WIHE6uo7KrJ2jGytBRRSlXZ6RUnNdoN7ex+1
vNqy9vHA0snz8oc3l8CdfWFvB5zd3M1K8VaNRbSYORB+UG2rlLiLipSkwHjhYiZ8ED1CgfBL/tPk
w3/k84RbKt2IO/udokR20giyBXXzUGWVgblLWrgcn0MjRX6rnd3vtKx2bvbyYR+6Q47QODHpXY4V
TAEtaneGxcFVqUP50/wNYl5rMY0RnZbt2VTtR4VkMrKGgUNwZdGyCJFD/K6y6KUi0K9/Plot3Rgj
gAUFG8j7+c5myvYPKJ5ygjFl+bap/N6vpXeRdtLXEMub8p1QBC2+qEGjn0LKNGvJ5OPd4ICTb9HJ
vbOa/oEnt3RFl3WmXrNFKaisEo3F44t3uKz32Fg2M6PEavjOwGPlaKdlpJ7MvdcdTdN0MPsk1C2H
blJi6LqVHmUngVaxB1I709kM6Jl2JAvJlIIIpQwrpIw5ZY/7/BHraAIqk92ohr1wegsmL/hUNA7T
yDaAp2JOj+KwPygWsOuORrjtdmzqfcYo6qtTC13WrOenI11kDcaMhecS9iFQf8dzvIamdfYdpduP
iZjCrKHgTzqdGSkBra5rHJyzEB9g3W99xPziJvED8pVJrPGNvoVgBxfCGzfYmq50yF0yjqltecrF
zntodlsiVych49tBULvORGxAZLENPIdQBhtdejt/4rnFlFdvWBdF+lOo5XIoHMnakdT0o6JgtCZh
IJ7E57ELF6nRTjHNbQ9kkjgJQcnLo1+S/63YEnJB2zAf+HmaoBuTPPKrisSZ+Qg/gtWNCQWtWM1W
DqO0iSbptYH1r/4frrKEXZgcuv4z3oznr1lgdLu+b0OqzBdguBlo4GMlTq/e8kegGeraynT/SECp
p0Jy2bxhx2p4RjG3TF0M7sBI+9Z9kvLISJPdL9JprrUr+BnUCNoz/uxrQTcYg91/WvYfrkvmzNiV
AwI1B1flIeWwb+tXdvZlNKVuH3GD3a+pZ4cksuS0oBSfPfKvk92RFArbP8+9rAW0soTIxdkv2wHW
mLGaSu+5TMMSAK/TQMTfVG43KE9cqvROZAvkZZ0T83S+eWBbW06E8rDkVGWYxdyB5cX8xVPoNo8k
m93ViSsZ0fE5+n5SOOXR4dZ92CWSVQ7cdPO49VJfjdVuRsazPDiAYqlq53usYmiKOEkUlCY8B1dR
++TrafwdcM8nCi7FpaQXC32zGlAtP8VkCtNFjAQ5669Py0WnyPqAuguoGjV+7Sm9zEaHQqPwnYNR
vVKDGTI+10kqUMeYiudKYVujphVxWsr44H2YCZx9jI9Fg7/H9sGQmgIjsmT8S1mE8a4QvLimKTKr
U7KrsCgt8LbnRYM3/xalHIEqpF0KJ2PG/LVv16+D0xjWJ5eGGicqdHFW+yAMRPa0ilNT3Poqnbl2
irciQAODv3Iu+fqtq6yeQlXSb1wKtrR7QW8I8dfBlz2ehoxo8HDoOe8Cz91WaG1lFx5qP+ISIhA+
gpYgL9nnl1/6aerm3vIhPLbktGK7PXzeZONMIrjPjde8/j83KcYjkSeV5b8ddlbeXaJizdtfCiYT
tZWOHlgxbCQM8ScpTB+ffO1HdGptdwQiu2V4dCF8tWTxHHyq9H8q5qlDVrSTt4Fyojdiw3pgeEw2
sBY4iRgz6kjyWzsDqzyeDAds6g1bGCIc5mHgYUAlydBm8X67y8BVJENX3/dW/AAywfBqvxjuTd7b
Z1FYPB61xCdkvoEC2osVLqxX1J0BQN/W0/NevM2OUvUNoBMEXzcta2Kvvh0zIEPqnL7QRNQbyWGz
wA6I0b2TGI8/ZZqeFlWvYxNAyO9xFHAy3bX5OEv/aHI0LKuvLwSD61n7pAgg24ze1eIDuZEbpAkB
G6ta0HKnnZMS3CdmQtgw96hzGc9ZG730JcLaBICDLY2DVZ1bSUzolFTYciOwLX39Argpce9TTAAp
rKa1Bovr/QzNjHJkAyCrNUzTmiTqevc72cQzou4cS7ut2zQV2IW+Ug0GIQ7J2BjY7ddNB6N8mLy7
AQuMi6HIDc5Bsediq9YYWxc5v6spDB5g0mRe1AjSeNy7q3qgZ+ajrznf7lebqI8d0lZPH1zfvQZv
mRFo85ig5QdrIpb2VGi3iR8AuDVAyf5eX4xmiXWELk0MQWVL1NJxOD72n9V6Tsa2XVom0FMP/1ej
wideW8Bpe6jnzIOaNvUsykI2QhZqfjjewQNLDEG2MmhOLh19WmhrFyRKrHAmH5auTFkR18hKw7kM
RtAfFOgq2REcLzmo4R1RPTPHCddAsDcvWzXVg7vJ72v8unqoqru+EwMe/ptsYIogluk92kYH/jdq
twmCQTlkirHT8imDmBOsIrgqHnN0tg6HMEuUlerwfbeTr/qo9oa1szA5I3tRK0mozc/b3RIGLBCa
W5lQuDxixbHnJItrE2ERemBBpqMBnXjks+KU8xEe6BS/Uaa/JbpX8uu1yImgjGaTfWrLJHS7ixK+
VCzT8eOHPCa1Xhh3ch0TSrf9cYNpGgRDbc5U7kEmc8MM/+PNw9b1CFxhu++6rT2/LwmBz6WgUwx1
J22xJhHgxHDeHZtsM2wkyS2cPx2bNo2uX94+MyD230sHlLlZQErSp0a3IMesuZmVQYPaZjo6DJZa
djCEnjN/gge9Em6F4K+gnO/Dj1rQWH0By5J0+8dg4D6PAB3UM1Gh2CU9icm+hntuSyIA/EL0I5oC
OORtmeyQbFUSPeDWknB6ljGZwgF5fCJBg5eIvm2HiGB93F0PFF1+ddLw6LVNkNvxSAt7zz8sioCc
DB1d47nAB2R8EItb9sDALBp2Wl1CDgHCYFuEohcOMafOmYNm2udMU3tjtcb/fsHOPUm0YRnbI26C
j3mYsZ4ukenOJR8c7jR6ZSNnoi7UKyR4AM4R0+NHrXW3+A/0SFaGJklR35+LjWaEEn/NWVqt8ug9
e4lD0nfQ2oUmpNiRr8w8r7Aw5b4fRJb+dlyASezQig+HBRtFSoG4Gn//ZHzfMo+zjkDXJv3DQuXB
us+bEh9Fc4aKuPFHT05wGsm7fJ0cx/rJ1rBu9SKswt3JXXpunS/BJ+TZ743+JZipZkcM0VPIeB7c
0kvmaqk03PwTOqWvrFvcEVGXB9ode3PPnlcwY/w0fA4ZjL6bO7P+CSyoyUIcUtTxY9ux2fNba7g2
hLwyh6TWfaElB+pbI/tUvTDgyZVjzoBcZe+JVcTW7EcI5GvmlnVeiwgqaWH2sOwE7TbR8YKymaqu
m4VLpDT+htOTOK5LLVFfpHa+XEDg4WoG9re9NUeP5qBfg/K64t2WpboVAZfauIziwk9teTNUXmB0
HbyfTgnJ13EeUE0zAJI0+mLOd71ZdBF38HDoz+aoeBW9QuGcqWRK2eDH0yucaspmZPWJnMnqZ+aR
vto+t/tNPWZLa1YyuNlB4H+tyI4pyZOk9pT0EKpSmUoaZGWP0dlhXKH4Ymn7Tqe9Ci64D0G/XUpx
WE0Yct3B33osLQkt9gMgQNwIw7VeCwoCzoL11rJvCIlVwtsVqRJZ1LXwalYzIDmESX/SjNSsAmKR
pMlL9fB+GFA4kaISNlvcbYSAYON5//StcN8XHnGb3pn3X8AM2WQcGSLewGtK+1By/1bOgGFme205
v6QR4Hl+L5O4FT+Xo+HyFaitzxXt72kk7vS1vBmrkbyT2hO6ZpIYauHmYfYjvM7GsApX3nrjjnbM
scBpBEIqEqS28foMpP6cxDMfWlNEkwevhcEGbyY7VsTKhwMQrZHD3YwkFkDc0MOJaVg1GU2m5VdE
1LKp2XfzbfaYCcxKnTRe0SOBnHlubO7hzk/ddDAItMq4gyDHt2+efFSCudVtgkAOQFpBMGARD7nl
bNfVF+9Y7rjiyp496qkO47A0MS6dQ9zZoT4USH7f2IdjuAVmVMZxUI4Sj+BOLDBPrmNm3M82oRJW
01Up0qCBoPVsq/ylta6YOXPiyY9ssyaKP99cKWfKSg0Jo9B9icDF84ZT6XY937nNe624dfGY2kyz
QeeNQV3eHnmBLkVl/hE51IFwM5b8MQuL+Gihe5VkZ97QRb5OKpGlrUPE1TTbVItqzOBv4h0UdjVo
lxvYtNQWJjI7vebQc8kvfcBcxWo9Ru2z2KkvdddXMEy2n+QbwyQIZn4XQgqq5/fNPMBjbGYcNwz/
5o37JJxoVb4KYQXUvu+k3EGgIL6AkmD/kph2SUuja2hjDv6bzbGW237AxLschPkPdu9xyyDx7kjV
hcI+y13PEriTEqxIJGVxQ7pnd+R6/O9qUL1KX2BYDWvR/Ar5vuxx7lEZiQEZUrIFGmjQOetDSNVp
rs7kox5EAeim8GDlF85D5jsZJR7t7Xex2YmdvzC3QXKKUtPCKA+21q+V0yaIIuiBYMv5yCzJfeD/
Ht7lUMxQhTYBuQejP5ufeD3l5mmYUUmBsqMjZhSz1Vpx/61yrUB+V/n6VT5ix2cV8gL4BurgF/IG
heXQe6GKqJiTUIcmdfZSCu2P9q2ac3C47hk3RmjVQBBAr+Dx/oghEMzhuCsEPGy2kF20DE5sTQyN
QxOqru/DdquaG1saHUaVKHLZJTAgHJZkikQ2/4CremUyseacz6k+08PrGZTiGIqP3TzyA9AmLzb6
5eC/xQnWtyiG81tboT6cTHU+RliW0NUAkGXLbL21aNfpLOn5UBhFYCQgmU6DgDdn4UzdK8KLZxnB
y6ll54yn6S5FSBEi0bgAfdm0v7lUrEBqkkqa1sB7vMT33aq0HkZWEW6Yq9PLp5yN5vL7KrvXURfR
TmOLtBbwEfjpWjohI0zEVRCvq1QxIsVZ8piBesHOkhMLNBOoggsJdrfCTTJuh6+MCuz//DddU1vw
bvqtbak4yXD2Mc9a+MKrVrk9oQqvKFz8tEHXRupeYH28lQ27FIE/X1rtLtZrps+Hhsabi2GFYHWH
qG/tX+ErRcaeBu00Z0TG9fWzLww13rLqv0DIWuOAIR09jLRg2nq/8UaKv8egdbpv9GA2DISTV8df
7rbUaOaElittb34fAsWlO0qyh2Vzvyg1ICERwrLa2DRxmx0JSuJhTWKtZbylKqul4DfKerfc0ORf
z91B9ul1LTG80MB7yib81H6NlwEBq7hgnGxragIE62RNLsQVnbD4f1KyyRgElfkNYOZqYKCpzFbU
WR/gJT52X90hybPRQxgQflvqeq8YmAPCP5HmltljU1C8Tblax5NYEr2WIGGxbH+/OFTgKCU6I/mI
O0e6tOBDLcAFtdUPIWRbBH8QA/j3vrEqoKmge5+TP8tNEr4tpmaH+RuuDtsPTYVi8x0m4R5/uloh
4/VQghEBlfFE9gj//qmbwCq3PaoVG51m0i00fpBrCLLl+jEcJZxZHRLz7GsJFTbGlTUWyOiVflpX
VxRh/xVAJv9iq0pUZM4gEo02MpzzBwp+Hn6aFTvy4rxs3Kfeu5uRQyIkNDupSs7HnbGdSLELfrhS
33X0FM2JQ4JafEThUKn3c6/fZDhiZAyydp3s80teiIPHqGbbYMDrXcXnT22k61joDdiYYj/t3iw5
QHsbSqwzxNd0lZOdVo87sga5c/sOjReAzZa4EGBZ1j1xpH/JzmGqcAPp3Bgo0SwI9mBmX5LFAYcN
cRJgoMZ6IM9r5PdjIsJAncyXctNIV8g0Mp31bSbcO28XAc3m9596rmWqEA4Lri3KPJ59VzwysfR2
/fEKk04vu+fXKi/jGTKZ8AO7aZ06fZNASPS+8x21s840gWkIrg0DPeMnrCmU9CDb/fu3tCtugukX
hJh26T3BBErr9jfxQAtbfLNDo6XdwA6d+0NFg05Qfu25qcVD0828AzQtocc4VfkBG0409PqAge8j
suI/U87pOGYrYN5snGLufeu+znAWU0RrFKwbem+aRPi0RRB+tftH3lusgdufGiIF884Twgw0G+pi
O8QW/quJjzM+Fcews4SoJIBF4ml1uGifTT6nozkEDlnL4HDpF7jKYWtSF1khlQh+PXQxWJS65AwS
0+2KRqLSq+1kxqJSrAQLR3Lr8Ky+8ZjUdZtKGcvnwM48OOxgJKHRjcOfuryAjLQXdFD/MEb136lu
IvW8H+NnCMH2I8NDY94/SYbgtf7MubEM9KKmxWym+ATy62oeAM18tR3lm7WW9jNVyIbPCjbyDyqT
qwJZpczJVIqbWo8Kv6jDwYOvXT9L9NSX5oPi2W0+LsHqrSo2Maj3wI0HONLfASRM3eAcFWnHPOYm
iUH9GfTWQMFj8yrhUDV4PcDjRc1Ye6T1M4iS/pHIowygn0TSAC2bPoGcB3uY8hbJAGp+Bjkt4uC0
Spt00fbXCCykD4b/jIN0SnOIUHxQU9sLoIWHh+HDdtZBjaZqY2r1HWISuDr0bDqs4N49JRT+sLR4
NcvBXnYT0AwdNhUpJYDyYdlgOKLih73Q/Qu3hOHj4yRaebu4mICU4fXMMAYtBBDKhVSNfADeZEpG
Ymspslil+93AYQuf+BKPCiy65pfIhAda4ykedeXffaTb0RJMbJuK6Gv+VFS35esP0WzZwaR3NBRY
ppzrOMfIKBg5jbnVa9oI7vtE8omqi7bIS1bnCgI3O9by4hagGiP+bzyJ5aKrbnh9bRX3aXPaUIRr
B6GIcSiW9d4Zv2anjOh2R2CAcQHxqer4tMJeneF1HiOQ/LPYrOqfbJCZZ01Zp6T3QOZoOEdsSDA/
+4rc562zJnFCDvyjbps7lDU1eQ8wCGt1vCUe02ARvjENsB4+mMtifWDlqKIZDY0a+gxc7vIwSFyT
87AYsO5VVqg/iHrcfi9C3UstcqpTK72xxvnuFhxOIzS9tJ30HW9f0H01a89PeDovAML618Go4CpI
wFNlR9ZHOQH7npdo6TjNL3vsBe/UdTk9R5reon1I24XviYeJyoWAeyOWXt0cR9OzpqlVcQHFDY//
dLsRUg4rK0Q5xnQ4W5fX4Ti3wmRExaokukR6DAa29uv9YZcTOLGJHHt7qn1DL4cKJlNn69kTtwyi
CJiALLb5jJh5Cn4DW9yNSFnMdnjjQZB7ZFoPRXEljI/cDX2pIR3maF09MqmYDn82roSmWNWJ7uE+
hHrrUc47uvPHxvgmQITuvw07waVJBEd2vkV+rlKhqyF8eDrkhWisWYP3nlURzrze0juB0kjaunIZ
6umM8zOyi5Baoi0HezGe73awfWcAU0aCo60GqnUlMP9r2YFHtbLjCUyiSWUDS36a2X2aHosq3TJV
0a+2pFpYaTXEcOItdlEGe3oQo3P7tppjjEEcaAUj/KbiiW6AogeyLFZvcjxH6baUMbj5QjFG5Ron
w7UZoC0K4ocx9WMHNBEjeowFwNfjEKDhOB42wOlhz2ZMExR3UDQ21gg6UqB5CUB2TiicKDFfokug
FsL0ZkAuiYMot1YP35hei7mN0tqUm7xPzjnVugoH9TVD2IsOs6DBJ2p2aL6MyxHpVDlzjzGCmEb0
IojbCdUmUVTpb6mVDGA09G52DkRD3OzS3CfSZaljIj8d2DP8LP/1J7BxByLxah//B+yBe5FYk4PX
K88AGxz8UKz+1lV5ZjcObcfxR8y2G0zBHWU1GgIKBTgps0l1+XyDZJZCZX5WU2Oj2zckWHG/IZbf
ShMUURTDYdoF47yk8s6z3cGIMMptefAJfNlQJGneIZX+vl6lM3aeHvAyJ8DZZ9/R6cbRlxQVhO6B
q8LjxTVv0NRgA4CRSIV7wJclauw/8GjrcphqHe2C1vqH1T64BdP+KS2rwCyYGUQFenM/t0Piafab
IFXKsZLvSpAlH2x7pkJuRJcJUWDGxEYRZhIFDrAJgySTvueUXeMVhZq0V0LxG4TdoORxLppaBjY3
/zBCYuDf7R766OUAyhBNQgzXrFzC1C4vVjI+B8XPRVYPNaukSGRKQQ/3TGmSImv0ynKF0CfTNOoY
m3IrkwunK+weYa77e9+6WUBmoCrhoptMQYUTF9FDhJTTXmLnqZj1B52sQjE4XksVeJ6Nl83ukKsY
0hpfGq5s54K96AjDgAc2zo/moksAqn9yd4CSwxj76graLSLErrmVtfYExTQwROjvPmzHWUu0Y6J6
nJkGpTw/OebnGJI5P8hqNUznCFh+2R8Y6KpGs//VZDQJPGB6Mb5Dsl9czls4fjFTpW7Wvuf05JVp
vtNlUrMYZfU1BIu120Dz3F6Hd7cPl8L6uq3/tNHsNt6g39W/uFpHkyM02oinybTBGmY8sF1VzhGx
x61+IxCv9qrlCxYfLr9RS9M0yzst3ahVDXmwk9t91Z5m04p7pqiyMRfcemwGZj4mdAzsNRrvv8e4
ekrV2pFE2sO2znv0xlttQSKFaFxF6/2ULcNx4u14Ay219sw4iWn1GRWNXZCP7nwDLQjKtSM711k+
XDvErx5ajNi1/i0vw+q+NZqZD3jbOoLOmOA13gzwDwvWEGcgQIGCXeAds7/BUPtfrcLIpd914DGw
6eW51EFweAbok7FP174EEbo2F9NULJttHn+EQvSdta5KV0uYAOy+6y5tue5ZUOaPE6qigh/1W5lU
erjRjCytYvVTmUEbbHENazNXnoNYENtENYrYrXe8in2A7OtmkYDost42nnrMWhtfqROqgrwkmJAG
JgkJeCcQew/FZOQvsl1lPunoYWB8Qu9oIY1h1aWAJaHw9gQcoheuOifdxwi+ACGYdFzf8NdQdYGS
+xr0AB0Ert03l80IWLo4iUv7oP17ThQWguqtJ34gzTJNsUM1p3R+Ph8OoWpdYXDh3u70EuetATHk
3IgmvuLNNSbg8p5RmM7JarT7IJN2UHEaKET570BGsBYICfk+CCy2E44ibjAFd32Ifu5k74ZlT3va
FmjUx4Qt7PPCjyG0elbO8hhFa2pqJ6DsIX51wojD4nASK0yKjqgtg5EQIfo3C7yYOUsoMYUD8frh
unL8OF6mmwMCztAAAkhXLrqnUnYf+9C2RLb3QsY6pRUn8ZdU3zu8z8Pqci2iNNtZnA5M5oElExta
6Nsxh59qm8FEU5kCv70aZUjb9Jla7UJr+D6F9K+voH/bMTOXmMh28p9CfpH2z9RJXGEPPPGoZnHW
bolceX3o4HEhp4Bwdgb7453etqMfy9KQTy5LLt8UGn4iIEc1a7bmGf8zfTgBAxu57t07NK50K9BL
KV+2EzP4wn4NbhtGf2EVwT2mr1KBLseUE/EA3iiTAovMe/SEyKDs1tpug7R0Lf+MMWxxSExUj9vk
FShya/Hp+3xN1CK0zg7m5o+20mS8UN5ycPyQ+QtbMjd55rF/cwBXIB1Q6lqFk3zl4xElyv3OTR/S
D7QKGMA5uyEivQIDqBvQxXE11Mi6hC+BLposiz/hzvZ+wgD+sRFZCP4+oUf/eB6fLC0PIQk+3I7N
PBQ2E2p4LIc89tPAg04TYp2Vu4kkDJPCzu798eK0Ds9iCi1P7BpPqWOcqix/JFvaTMipuH46AMay
oXMgwK15x16oEQYN2J8djr6luegmoL8irOFhjEJMi0Jk8bB2m93vkycVNxgSWaExDA+kmuiJhYV5
475+f6TgN1mIxSGkS393sHMDu64wgwt9ioNvUqCneF/xs9Vlho157qm9G9WZnotalDKuNabjC4ig
CPG6i3BssgRj2ZD2jSJdq0oTODCtLISAFZyowj66RTT8+YEINGfIs2UkUdN8FUQkB7LZ5RWNQ0+J
yyqk2xFxn2xmuh3Doa+P21g5WP1S52q0sCwdj5hoR9PizFjpD19IRCjbtTJfF/NcA3HpsxzpWW9i
sENVsgX5z47JyIvNbuFSP7NItr76Iw3qr8RiyLbh/GK53ECYC2Y30iYBJISgOUfqyuOntG4Z8zrF
tGdetJSrMR/Li1e54YILD52iLhGTtiC2rTPXsVjeu3iWuu3VA7U0wZ5WAQLDSgE92DUmwiiJPvlX
FtxIiCGE2sQchGXutaSkRxsdLvRaJgHUnhodHlFiIygp77X7HvmTJZ9IeHN7+SJ93jp5wInwBCEL
6xPgTWM3B1Dv2MYk+riTYJUy0PlA5muccxVdo5zudASoR8KQJB3CPrWzMa8Q4vnBtfOvXOprxoih
e3QuUM8AHrLSC5l3hBoCDTL7A1wOcr+piN+JQJlFbIk5EcGr+RU5TOsK9buznNPfzrpUnq0hpMM1
k8gPtpYCsgsYRL17HU0cHJ35X5ieyKFbWMLBs1eL3BpRbWVsI+xkjBII+tLeIq0f8R48TBf7v2CY
Oe9XEgbOT98bJ17LRkkKppJ5iGycAXfa0G1pjSNQn+6Fq6uLcPd4AWnlKspTrFCviL/F8g8STnOS
y4R4E2lW5l7T4Tv2uoeDxwgC5FByKX8xaj/SmjreP1HXat+zg1/UevbMOIBD5bId5iLG/se4x/PY
pikquiIYprRIExOOLAL34WaZlTrrSRJybK1ozxvxdvyxnTT55i24OE8BRu+odLbAWPMFfFjoRRCx
3dTr5+z9oujNzZEhCphBLHTdlkLA7zqGIxMarxjRQy9enlrRMk6L7g/6c2LuYP1N727WIIXBFKTa
A5EAQiEcdA6lzjTvhy0nWKxkqWOEe89h1VwPMzbA9WZfV79b94/Yjsv+goi7J04sQkUSxG+pgKnQ
8QDp/tVS7jbiOLWok4skNfCq1f/kFp45fKu30ym72qZY5HnqAq6BTj4sTWaHSBgfoVqZPbe0aphj
UGEoiHhF0o2gFdrACYgc820a7Utb/L8mEcoB9JL/BHaYvXh6ngAUkMMKvLJC+5Z9w9UQd5p1nVOB
nDiP+St6KCkZDrfR/tsaEJh9MUGGmcqKTTLnprLKLjqHg8nKkig3WVjvPWfXoF2CQj87wN9RebNg
aHhPa2Gli6zHwANm0sDMSA0lG97qBmgxcT0wC1HP+hPftuecCw2iU9+3D8Ke/XHnlSHQgDVIAlZJ
RudQseHz+DnYC0jeCjmEVAn/iQioGmlDVyw2P+ZdY5DGHISP5J9GS0Ysb93ONTY9fOskfSuittvC
0U+Vzp34X6sBFJyZE9/i/rjqF4XL8Q+/nA/Bdhi8h/PaSVc4yIqk+Zk2JMm4tx/sHtkzSMjaNlD8
h6eexhzqIJKvUw6B+X0RYBsAGC6Lho6ZWcRfnuaHZ9lHoZ7LEgiOcrQ/kjF/IkpfW4t3cNawhCjT
NxLnt4+HtnhXDR5yHbhsiRARNMD+NGsEm45U7TENaD4sUkzmymeAr5xy4DIFnDOYNgiIcIgTGe3l
/FOSFv2dIOTjZ3HM7ytV2agBNETrMR9I6RcrNFAy+LYaIyVHR57TADzVrcw8FAT1Hd0N4sJCgGKj
2LKmHckue/8M61tY9k3FqIdC3p00TAXlzYW04KeBfcIVnPlfrNVUPN8eDlYkwcZecUciSV9M4rDC
K2X22fWRjx4uReIB3JDAxz18GHqzdkKv1ozUaNJJKaUjt8tPrR+AzZ5IR06Rffos+CPEFHGWqmrD
jo5X/P4EFPTf0uSr+djwHIjXEElA6MxQ639LCDxjnsHdkowptRPYrJ3e1kaYG3qW+/t0Ehle8pz+
GdiRFfM/1LsYb/1wZrl5MsgEvDrSJ9S/ZGy5PWeCEpRHbLhRLDSUV4ngYuNv+QH/rpEbrddrmHzJ
76HZFj5iOjaUr2uLc6STh/SZGFMxGAhe9Rq/1/qEuaWb4c/tYTfvm51fq2kYsfYmoVd4kBrfTfpu
2Y2lpcuDQ80j44UX0s/cAoq1Zi/mPdztq3HeF4h7Pj/VYT12EPnQefc7fD4BTMya3GZKHEg3Lmtn
F23oSW0FJC1ZenB6Pj442kUfGVE7OP4cn21TLgb7LV5WQrPsVzUf3f/RwsYC1IbUcsI+tbjLCrOG
MGqMkUJt0ccqHPftP78B5ec2QLYDGS6b6YOnk89WwHX+vZdQequM4OACfa/VtHyNkph2zgtXeX2q
AdwLZilbhTk76kYizslrq3apOPlb/82ayoqlhRLyYpC8WGLoS34uoj2hPFu1e/Auw7sHOVu+arK7
+qSrnpFKvg/gZI63cYZ88/eqtutKfrBvu7LQaWqOjfCDgiLz8+16dOVIPaUEvaKE04Q2OcaxI9pv
enQ/WthjRZ7RDtYkWWmDos7kEAq3xv/b3KCZuimyQo1s293sbq6yk+iyKpUqPY7lll4cmYKq1D6V
3aoOv4uMbPJ5w76nBgDDDnlkvMOrPph7sSl2been3o1Zu5b/AeEuipsDbzQMk23QtcX6aobkKdaW
Smh4PZGHsC/uhH7BX31L52K/P6/jXUdo4A7KcQHQQ2fgDPJfiXiCLSCw+YVDhmILJc2LEFQa2LQE
rhirXFwys5yrS2BDla7iDDoNjBouQpw+X34/f64mVsgv2OikcHIUjhn32QbIERWBoxs3p/rzBh3I
rNPpy96Mu632U6kLVIuTuAjjAw2vGusSO1mbCVXKpkj0o7hdJxvRCJaGZxbOziKcuVbJzl5y+co4
GSDtz7BRND0RnSMy+dP5FyyIFkGNuz53zzQW5xqSts7WBm69JBFXikCardviuGpeWak7EGmCoqBr
L+TZaDIR4e67t4iyvRU8L0AJVnzaY+PbkBYOWU+9eE55XFkJI/ONQCrdDHiyHevTpH+wcKBTgCl8
frEjuVd3BUHbseU3ZquH2noeQMJCtZuBaT0bcK3ur/slxpwzjZK5cI1qFcRgxaKvWIiikQfKgfHJ
VqEQP5sQivbbR9aPAg990wJgz6/S3Q55E6U3b6FZbBg+XtUsEMiwUQ4lv+onVBA+mL+QeK5K52ky
VIlFrPUeDGRcpbo+V9VymM/+bPB61juwCONT26NSuqlMuR98ewXzm9tnzIr7QEG+qIfmeJJZCtnU
zBrRLRa80mLI3yt364QOBMIfwk6d5EpzT4xnDHx3vpcTIXmBPeSUsYDi8beyKUVJTiQHCBJI39dj
/DIm59GvpOtkWzlZWBhHug6SHd1JxiEwqWBAHDvyYuAsHSVg/6eV71DVeLKPm1+MevlYfZBFlNLd
VDkTr2HbICXG+VkWsul1jQgCaNvnYY5xf6wFyFVjlI8mWbhEG9LiiRp8DzGS0ERZMn0HUZ/sdoBk
DVO8J2o4UB/tiXfQHep2JqF/WIKUhv2PbybwLy/FkbRBxKGUEsU0kz/GowOsjwE7qTULZXyTzdvm
6JCPxxT0Afb86FvseX2kkqMbPijsa6nEyVaSMbCTaTkRQGZsCjxDRYExe7FmpYPPnFiVw7f5k396
Ww/eQZmq4UHdnJbSQytVJr5f6qZstlJ7hvtQ71rsJT/pc227H67EPEPg05gIm+5335R1osp+eK30
HNTAqSpahJv7QQtOt9KKpYkEvAuj1rGe7T8SNO37znYNEoipV5f/+XzZaMd+0bp5sPVk9UnBseLb
IevGSJAQqxWQ6ndP2qWuHZEorgjFr4QdNwZHUCkQGq60fTOFU0eR4GTb4Ovushf0pJIN9zPbsMGo
+FeIQkrHknj52ha1pRSTOfqOT9uiqtZvohOSaFnxICd7se47Lvw9+x9Q/9FpHdx542ElmFDtsI26
AW3LZKLfK8beQrfj8WNWzN1pBjhptg2y5VRX5TRbV6Zw3fDdlFOMK6BvEiOkqsTL0yEn6cwkpLPD
U6VjbYYPASJW+IkPK7nRtbpziyIdileSCap3aSzqs94KWKHQLkwMMBzB0hog1RDWHjHMYrY9KjBZ
gTXsEDTjMweQ5jdLYMU47RBKNYJ27/hvVZSqFne6tls8YVCv7HbnhuCbHUZbLZohgXqp4mU4Qo4P
sq/Ax2IGeOfl/4MS8evXc2fTuGp6eyirUANDEMdtdLH2eTlWPKLC16cEni/9yFQd+ZZQo+4FgbAo
sePX7eusLWTdTtvIfkPoc5QM9m9rF8LI+AILxF1eKz6eu9xGOWZZNMMeW5hiGtsHAQ1k4Hi01H0F
OGjKANmMWC99FQy0g1WYWCrpksOdQtglTgudau/h9rHIsIqFR2UrgdVv+qMgLBBsNexZoZCiXu+q
gUn9mjOeJHydyBKrTljBfDCrBP6RTVHCyzikyfEJrYu2yYZQMcJ9vpfyIK8HdhdBC3sh9Ex2mW4C
neArizjBR8v7tDPJ7Ke6zlqfC8uSahp0VcoCtXHhojHVT6Xc0RN7oAoYSuIU9A3wvWXh7mw4NTua
v+CLiraKtYC/rnn2VSe6/VUyEV/EilXl23VTBubfeYgaYu/Ll0xuo6wjT++IvPMWAMQMGADkKZ/p
wIj7UPyfbNJKO1hGsNATbuFIoAqlSbNIU1XE+HIKYIHA2Esbxonl1S1jf4KqrqVEAkwpcKsx3Fqd
xeZ5e3q87Rd06pdnexVRdudZy4KQmL+IN2lDqsiazuBIfskBo42Xk0oXUQ5SqaEm0LkKMEBDJmcv
GnZSjSdjfmt8SdFbtd1x+6XixfFuiOZqS85EneZmknptZDK7XZVtfbO4SCzvLQx5/gjXBSzsWErd
f1+E4CtYUx8rxHL7WquURJb0gFyf9zY8DQcuY2EoQPN1KCDnpToq9r+GuNSzgZKr3AMcvIjsJ6zA
PnhBveLNIYYTUg4fpYZqZ1Z3ItT6w58xOcSofZtq2vc045zG3RNawu6SvHElN+QE8hcStdZVdrsq
ZXQtMVigKpPKMrB8BLhpTfZPe+f+6XRAIL8R8JCUQxgReZznIxcB3FMU8krFa2HjnxA4MhKLbFYx
uS7mDXh9NCKV7iCaLrDWGvBBwsgPogokeYpmLRwmUgiMKxBMOabYKUO/QEFuXsWSy7Z65uH8KKcG
5mWr4GsQxct/mGw6QvMUyGo7Bj80hnwHmg/2uSLxjJN3kofOg0/2eOCoyC5JAz5+MdQrG8sKsWty
BxIj/f7cFQQgpUmw0/jBtganoKsnYD07wWNg26iDshJR4WOSWzuZSVu32foX0H3wrdUgbnSZ8esD
PolEKoPuYw8L2R+Bw3KMpTtBF642XV/walXrb7rWasLn4D6I4d+E25GnnIHBm+Eg2Ws/lOrLKRgS
4rsWlGnq006Fiihi2b2Nqi47q2w1G62KwfOQxqK4V2xJvZ5CYdedsdSMmtMntHclziVR3qqzW3Ld
hryXAsBHJgYZAw9BbANxFgh8CJ6Vw4tBC+OjGGENUL7eoiSiV+PZQopOZkGDCGDeAiNN3Ak8nvyR
H5Ys91gkqJ52zTIinZz2hIrBXWt6iHCvb6U3Gnl3QgKGFYO0HewdJ3PU7eyYYnwX8s8h/FNsbyZM
voHhQCvQ3cSeYJoGRrIDf0xKu+mtqGUknd1u7TkYZxmd6qZjPNcxTqc5M4DrotfggTiyGQyvWScZ
/pIe0Hr8PRnNpIZh/5SvQvJ+M/XOuyXUbWhod4pII2nWX7TlkOLngdB8wwQdQg1M4QyzL9qcYSYA
tSeFSmWZIw9qVRNLxCemIBe+kWDbHML7rj4SgWUenoDj26iszbxucpgCwKpvEt8g43MtJmrHfnzF
gDPwE5ezsO+0nOJqzgmR1NX81lmDT38E4t5HKsq/+6BoWgeokctO8l/BNhCIe5MbzLKdm0XirzPM
m4K7BGtDj+iE86CbrQb06ubLo9vclqaiOz+iK3Jw+kAnfVfleS4XkApqkLHBKoJU74CAqhqALUpz
5oQIeojMo2Y+3e5subevNFx29rc5bcJUBz5Q8jPK2jxcQu9v0YCNPQylE5LLqFBiAgAa3HL+4q2U
CkafglzfXIv44+q42BD7c2X5i1bMpcHlGFh6fxfSsLFeMafstk4X7PzQ6KPDupFkvMgx8yaAqyvP
rfiMcE/dGf6dzQ4gVRUaUQCV7cEIBXW+xym9lNImZv80hq/U3cOTqDqz9Nl2I+4OyXd4f7wQC0a1
rwq0RMTLu0ky7Vv2CtCafVdhpVHDcb1Vim8AKUc0sL68mT37oqwnr4S5RzWW+LZ+561TgLeDwlx5
7431RJxnLKKtqTXKItgVSxGKNcH8xKMv399IZkXJeKsrADtYTLEEYaZxUozTNQN1uSCwgPmXuU1b
RhBZoVyqbN5NiIMEjnrpE7rHgUuMs9l9xT8qiTIVxiao32omqvJ/PlWQgfwhFItg4orGEBdemsmE
pm8tfe384scNeIJb41EWSj7PBpsi21GOImk/p/JgCLJiBZXZgLl5UrfzfOd3xtdSfXd5+ghmJyen
EtKm8ccOfWQfd7hVmt0vIJDWIkk3LesMr5aQjz3pueWsuDQkXNPw63QZOFd0gV4DE2t6u3+JQAlo
RaooqjjQoR06GtHqN9wcZRJJ4Rk0IfFRnjHqcPc50tDZAvPutaoMAnelSMXu10iaEpUhb2vOkAHE
SnFNALNWX+rDRCLaK3IVnE1e/3Yl6uILBZpqREfPnrnJObLkk8Y4rIa58aUF4HPuYSSvJQ/nVGCv
YzHi+yZuOcXCYr1XFJNwi0mLiXBrQHFkvXSAMIu+vi4K1M0TldcrIGx6RIDWQpil/FIZUQO73Nim
DMGV7gCCvyQ5EWrfNU6hXcmYEfjmV8xZM6CVmBhFmbdNf+2ClbIfN+jgULT1pHQQCBB/dZ0gUAW0
eNc/2BUvpdinMoOg2tdFKOjR1K0wzirAvqZDRbw+OPc6zi69DfLDCx495pAmDtuknCN5W54FP1Pw
c++xix2RvBk4J+42pv1kpugeRlWoJy8TJqRgrLld0pu2vwkovYd9JbMq9gCcALuZWKm+zhN9zl9G
oF9I9AML/k/V3r0vcmi1u7Fw5rfK10x2juLlUosSO2MVyptyUPPcrVqTvMhPOmLIQ5lQGXe4P/wF
lKg6cL1YYEYJ4W5/MWUiuY4JOyNhjvHPQT/btEQBxZua6Ex+FYAMfxyp+Srm1UNAMbgQ/Gututcf
MmIDo5URhNilcKtPh7hNpHpqA2rIy7ePhUK7qb9xjc/wwLbXxsgg9evNg2RIifFOyU8ydUXjPgUL
yGIlJ9QVLv/aaOUn4PyZ8ebxErggu0ACZ5UzarrZ03D6RQLrgryHXbX9fexd2DSt28VCcI4Qvc0I
UdIEMIbJaM3d1cWOjafa1GWWir6Ruk3mc5uinN0GptZndEnF7KuhaHy2+huzB2U8BrwgurqNXKsg
XFjAUsUN4D9jWhzrlJNo2BfIg4jEktmpmt5bqc4YR75N3YPzm3442i38Flm/PV3z7JgwgEVQwR/c
eKrXf39GPHADP1l+wLOFWJBJCvkxcRBrc9qtzxgb4nISM5CQyfQlZmCZyEO2VxBO+ddCbxlYx3N7
K1pNhlwi5uQAPAc7Q2xYC03/mPQ0e7+eEbjf/J7ojBf6c2FsOz5lJwDXplNyeyvcHKryRj1WUik0
vOXEA71lnnGOx/E3z0leQkQEWKlzKlk/9bngI8eJRQHj/sTiEpZt904Mh7avbFM881H0t5gvIADu
UHBD0uqLMCNZRx3VJIbxduIQOjg2ca+PYfR3vaX8LZS4MhBG+yeZmo50PIe0ubhjnWPdNaC9VTrA
901VS11qPXIVdMhMiAXCOi0QBrctd6xak80ewIi5VRTkgi0vs5selW9ffxLYCeRZab9nSc9ddJOj
M0z2iIIYMYoSnKEwHNHavjtkKhPE0ytsAOXRKSUmg0/9bPveacqFWK1RoEIHysZAGlV7xrjGSlTS
xjaH5dsOGjJrA6Y/n2gn9itL5rrtXjlG2i0M9mwZyMgsKJwI/tJLmhHjciXDg8MtJMw8IsbIvAop
tVimnXK80bsVEDNICNOyCDK64idRrruQxKh6gt6TBnIF1cfq3OZtR8MvLZ67AOpAoTdF8/l9fjDU
f9nCG/v4/g2rKJJkrhYD87Kt2zeX34RODkj2XLdyLnvOMpzSoUuq+u2hdR3SRMKWvVVRXRuIkRaH
EK8/smlrsFu1YrcogmV13ij+yPx7zA+4YzPSe3imbu5GUrVhyo/eNTg8YMfprpcmgrJhI7SmRFls
e2BewNCH31nzY/xdvEh53zqLrttefimJIfzzEsoNw2eE0gmJbAZCHiKgN2Amq6XY7E76pGUMh0j1
3bLgf189x931Nt4fQudC6XQf935ODOgbkIHxG2GB4jACCOWD4o0qhBbX+8zUI72hLS3lTVs52up+
NS+mVU0Ff8CtYd/gEQz5MCW6sCofE7p5Bk/CTF0XyU+1mtUhgDir3q1wfn69GEVXLJ/mBie7UFHq
nGZtp0j/WycsMYUkH/pA5AvZm1QwVfdBHF/Z0Eljj4PiAb9WIgXW9Z/oDrpobkfmH9PJfh4mH7Ey
EaQMG6FIjUutlKhfKh/oVaw43enu6I0uJGXY8u6sj0gJQ3YekIfJ9C3LzDsg0dAJHzjyNiuhQMir
WmcQNjyxYhyKOir6wYpkwidcHkAkDI5lL9hbqtddzJfChMyA5rEcU+hxj8axNqh5Q/EphuITd2gX
FbKqO48e4NCjojEG7kcihM0MQMZfABQwCkFvcs4lvBhvc+sNKhb5BXx/ID26nsTnOF6iUAdSxDt+
T1xHAmiKFKwMib4B0lVZ8LEIHACUCJQGiI+TgqmzXpO8ciAC+RNCVNgOK80imkUv3PvWMYsIuBYI
N+vjlloj23EgrxrhznmKSdjOL/7DqfhKHXqFKq+LZWWtjqPUXRVAmyXjaUxjglDzpeFAAp0cO33N
of4yBkS9OrVsH6+f1HxxxnRYV9EsZTKp69TIWxgSnmPo9Rjf+EFRVwpd029GhDnHypQFarDlfXKP
O86Mb3ctUVSYRqO7WihxGRiOPOqTHnUv20CriawesMvRo+hQOHLPHaJhUfOJ76zwa+5k+9/JNkv+
E4cjFdjsMAbeHryXRZZwuFBZVKiw7FNHFJpDZ4oMduk3WBRAOJzQHCLkACojAK0v9WcfZoFvu/Sc
zy3HdfUabG4FM1JB/MmnUJiY3lsQRL4X/lhCzm9ubZY80F/dYb7uq+YKoXr1wusUgPCM+IDYSM15
NcuusW73grd+VMduJ+HU1DyyOOrUl9K/VIdJ2DkAcrMUGDUChhYBUsZ5nK6Abl6Vkx6mETQyr2C7
RT11EbGRmsYJ95cL/TXIu+SBb7t7ltnZxHgg9LcsL5qL2hDI/sSIvPVIJfkR3yAdnJGvDau6brrh
McKANOxOj8nw/IUm0jwd22/QvfrBfDQ5HQ2D6gnc8AJbRcjatDTHtXqsRT97CYJ2183zbqNHTiCd
T66jkE9Yfaq4tzIJrhSmOsCHiRXg1ydc+4HqyEFfnXYbIY+uOvME7DZZO9BDXK7E1D8h9RslSEpG
zXElL/05WTAELPIcAuJs3JhuA1QnJzgJHKyWKF7g68Of4viaKnSlsoeLtaybOXfsn6dCQdNMzg1w
yXepPhLVGcbMfAXWp2MXZQhSbT6cJ0mw35e2JIUA4W4lA/YY9+ePfujjbmhx8/Mg6VE1F3cNQW2l
REkEVZ/lE5xhPlMIhkUmJ2qR+OvZVP3w8H+S/eSVgvz6uIGazhs+x+eFSjTe4UU75A9dcOpw/eR8
smVnIxO+ROmagerCDu3U1yh/b1ysygtgVOQ3AXciVIvox46WuUXQRfBAeaJbOBICjmqIzli5vFUl
vpSoFsT2ucqpdQnOC/IafJuQAOUppw5zVJItseFPuK4PUDOQGJFToIgVrxT54iNF57l6x87jh8uM
FTcvXMV5r0TlRQ3RbdpTKbIesIAnmcnjjt4kvBzCrhAph5HvWuPz7/Y72m5zYzaQZf/MkkD0zuRb
NLNApKxUM2eAzPRtV30XR6MAmVVk7T2GLZssqgymlf+ibkOr/DrOpsrHNfR4ObinJZ9y2UsUrTEU
ucxr47TNMwx6nOUvDG7PTJXDCxJFrf8RWVrS66SjzWvH2nLqCjBIHUjcxYagCYo83vJjPCY630/X
TK5xe8oFsyCsJ44bj1QBhljnYmbIESuREsR0bTBZG/xoPPdTq5nTHRbxtJOSuQVxHRGNyvoE0q1E
8r59sqqej5I8LVV4jZaM/rw04ItKWa39lFKKoxS9QjJysYwaG5w+yA/rluZYEL0QSRR6SC1QA103
DFVpaPXE8CpHF+/q7dVAOCy2JXxf/xiEWM5+Pxoq5Tp68rKUUGUj0LGQ95jpl6Xieho5UBDsYSn/
9XiLVjs5xjnnA8r+Ft2cOR381xU5FwarMTgq8zBJJjaCu07bPo7mBpwwE0ySi6RcKCGMzOmU0pB0
99MjndEK9EBuHnzHNYXbGcOc0D/2dV1n5GdPPKXZvRyaaK+c+XsDZVqtoC8Nhj9+zX9tgynS/9VQ
vF60WyhxZ/3HGOSyBSO2/lWjNhrGHQJ93zUMRefLKH1uNqmgJXVxfQw5ViJAOgNxjdW77ak31fyY
4lLZohGhU3xRIr/GUA+OeaUk+3u/XbEuscLttfNcOyEOQhyzvSrvds1c8H1AZDXE6yAZO6EEaBH0
Ekf29fot4WS6dg9tPpK/BZYj/UrnxmJeAaK/rA8teYEpdh2km7m5ITRMWAifFZJk4xu4Shk5A1rP
Yz01uQC7jE/Uj+mO3WSNVnZJEtt8tJbqOAnyUywcsnooE3WDud1puKeACJtOBpLVrXgXTNrwaRr2
756Dcx7dCyXU0Is33VQGLTZt9bvN1qihlvOqdub6Dz0rSmC8zRqJui6+Poc2HxZfNPXwERwnHGgF
tH5Avvc4rZlr8k27N+tnIhLraWoiy6INR5sqWkKe1O5XU+zPEncI5wgCIYhPs0MHNEQpJQiyqGVH
w5OQHR6spKKb1tvF6GFNCILNbsGs2FKa1Ny3CKqnTlYTx9Mtyxd8ahISK+7ngkajOn3g4U1LTfvI
ortpnkNcLXPdL/xTFGAIA8AL5oqJq/RWcJEG+UndflOU7DYZXbq/VxO0t5O3neoYFO5/zkuQ7sAj
OURhiTcdRV35X0uzfxuPOBn7Hmtx1aLI1lMJx+rzWZsUa5ml0ezga79eS/I/a/+Bxg7B3wQtU3IL
tqOPS2m/jj2udmM87Sdghd4A+vrmTSEe+bqQZQPHAPttX4VEMpf6X/ryXG0xLIzG7v1AYdN6yZSi
AqoKfpPuekPTWvuJMSOGsSotuFiEkvdUzSpve8RA17+0lSSB/nMeznygNYNkyr+7c0gXoocHVpY7
+nuYX/ndcc2g9aE/atrgk2kAf0UGdSu4weVd68rz60pDjym2YG+WAOiA4y5ROyo+vhL3avbRA8+4
GAk2wROde3E+fUrKM3boD5GWv84qLVXtEfv7QXYT11rM+qB/PesaV8eONf10mkSoDxnHM2vEpB1l
sbFalVzoY7wRZBcWNC8xtEk7oFolTLJfIIUu4mUe/qbv70frsb+JM82ssFUzJhsuBFMadb7MHBVy
qjf2LdEQ+kqyxPx5kYDtF9rm4kCJrJHFSODL4yZmUb47Z8ITfQCKoNiHyTkrvYPSXaoiv4YWdHpO
I2BphpbOAMwyBiJhPET0Q69r6qTIv/OaYucNhmxjMoWqRJA/xT+YxCN07vWwBGb+39rv8RFgkKwZ
/2jyZeopAoR5PfA5PX3tY5KNnglOs3w/OfV4+8kd2H+uc3msuVc2D5HFMWHgM37HjxrZpde7wfDF
U9HLCK9+m7mFuJL3Opw0AivSi7+nhKIHwWGuZTj8KAhILhBzTnC+d2PwwhAsYbob0jDd6tDs6Op/
G9iQGIKw4dCuK+QW34Fj/lXAwgt0W8OCD91D/Dr4cUufLeRBzGG/3K/9ue/LwKyQVTYsxOH3r4Wx
OSHap0ypnCZHi3wXXM6nmxPZ0WTe1rrNN88zw421uhvjyrhyFDpA2sowUrtLOXAmYSTbZRfEgn6b
n0f5Kh8kTfLHNEuiM8TWZU5Gs0IxbNKxE0tzH8GWRkiU5HhRM/BWWtvgTUhmmXAQxRLl8VZ2XjA/
otSJ86eWZCNvkSnPd98gP7DAWelYrwbb2XmaO9OaMAVtfkkRFUmMZGCra0k43eeoEzLNgkUv5i+h
hMkLkQz4ejc278PqQVqFsI28iln3S8xybcpg/9zblxLgUv/1y+PKPWAji8YBB3H1DkTt+6BrDJSs
zH1sstCsQWZBQFNBPyncuBimjy+6CbwXZhh26qbGvo5ttls6NyBn3HCMBzvL4FtcZ6Ir4Ddd2/2X
QAgpwO2VMK6CGmJKElGhZ1Wy/DehlyNP52J95dsjVeOJE7pIgX61jk/Qmro8R1BhjgbW1g7axEva
Y5uUsjrOZs8nVYdqTIf96he5zg2+g/LxfKR/V3qx9ly1oXGzWDboFZEtcaBMCeZVmwkW+OWKk7IB
zGiEnSkv3qw+R+p5D23JQaX3uXZ2gYQsBAifAoGb3sI6vn7VdAN3AnnfUmruoy5Cx8oCpB5xnADZ
sLMMxGojZeaKReBeXeQctYN4gZVJK7jI1MDqj8+vSmZYWrcEHkt0t6quEvoezntJEEKzmIHy5uac
37UixgGOWg07SuBGFj9iFDkDmWL8bsNDHPOaQoEP/dmwf92H1JvPuJNJfRFwKjYEPHKnKKGK5GNm
u1sPAf9x6or1FQC4KDMUnI/IcmgUI1fGO2oXCQUtne6xlrPYkG1NV6fWIG+dSkYCbbfgdO2WD9ew
hJDPl+8mOp2O1Ahgguwz9d/2J3SejCfP1L5/he1t9j9w23Qy/JnlQxRMsIoK0SND2uMgKJ6PRpEm
KLaibvQrS14teVlRmN7S2Ibet9lMnTnYW+d/VkqsROhxk0zMuX2KI5++2vYfRdNKWXCJ5rn25jmR
nPs13JO6KBv35BHGHqGJDBrYuvdCKyzxSiN0cjJFvNBX6JKaFUCGhkNEnYYq2MFTzmTzWWuO82aF
np+pkRLnShF/825TVX1xXRC5nls5GM4wTuvgUyJd2bGTURQK/yQ62wJs4ZVTF5dpjCzYeLO8OGxP
k5MFxRV8pQb+UzVUfaqPHRmzL1ZmlmwYRRjSkdsOjeHnN+rbCXLAYGjKC/h1qkPng6kUQeMwZKa9
QH7LYUcN884A9XFQDnHoqYlGA5aEtTeZpJu2zfPNejjsAt4iZhenvMQb9pOYJqWxqXMkU0c9jh2k
nu23ph9KKcYUC4kAISb2cixZgL+mac0RJSo3Db+09K1elA6iHGqAe6Q83DDOzb7w7ATWXONIFWK8
HBKE2KgGMYr87X9kJo0RPFVJjRE+Mau1kaATDV1sext9eZHeYv9t7XDmlr6bAXts/fV0uhJzJQg/
ZyOgnknEKhcTYiRr2z6pp4NoE476UaNmria97uvi34Ea5teT5aZ389gswrnY8aD/J6d61n3bndx9
aY42eo4xuJCNE9FIrDHEoqUgI4m5BobTCbTW0xdKG8tY6N+K3SJJKH/7PQSSs0maRrooFY1tLRpn
hJo42qFE7LbYAbos/+sCmmI3VbD4OKrsXSQwE5lQbGAbiKi7OItePOupsqtcN1gGwHjDckCRkc4Q
IN6LxPGWCx9KSNY4HNSnb6aYVgUdl7zm7MzdwZSO7TeI/NDEieXKtBzlAAOclU/fpRCDkCrOE7Cf
kdYi1IB8bpVGa6TOGDCDTa0qYeirOfPwW2QyVxVfMv1FSyoTa3cv3aMPFGXmKRVmIDOuZsWfArpx
VfNZM3EwvSlw447/w6NWyXwBl45jvPUYKR5R01X/YsT1LS5dmOCKsVF8qFKGHbiygSOIBGYXNWdE
hrTSQGXwgaq41/pUAjdi9sJy6FwrQOOFPAS1nkysN4BOXXSziS/BSYB2StMeAaIK3WDci1vgcs9P
3X5611ygd0biIKlFn50Tvp1VieYE1yvupJwstsmwo8j1t++/Bqr2Jpf8XvWMMF0ajh9dx3pcPo/9
oIFpFSVkSyfuw4H0FOlmwla8A08P0cXuLIh/L6+NRv5T3Apx7wJh5j6dl9NGo3PhBvM/3LLpJYas
4PTAh4nKfKOu2jFsiDdPYTBpi8Zf15aFOGrYl6sbH7viqj3spcJavX/lzYnrfmaaHeqFZT8J4PLw
NBbfs2EsYGfxOeDZSFpjvF/94WDIiXmj/41V5QjdTUHZr3wF4TZa9Jm0ai8euN9kf+gXQe3YmxnA
shWC3azCTJB7qH5gG2yMNb9+yoWQZ8M4hKcfqkbQeEfW1NX4Ax5sIg1e3UV3DwFGr2zDhMFjgfEL
fh/HhNpuKbgOSRch1i4yF84CgwrZW1ZqVV5qW6YzRL++1FrtHNOHSBekIhhXJtGaIXwsbV+kPEJI
01UhGfWLoegrExPwfVe4dv4FMdh3LWViSOTlVEUnwwpOxyfm1LMprhczZe+ZZf1D0crOLi0MsmIP
AxxHo3cTDbJJla+cPPK2q0+zNuUu6p5B4ptSVKPWlztnGB9Fwm73Yy3Cbn7Qd47945PKnxB5aUUf
HJZzbrdBDacj65+Aer9/HiCpP1medtPCyRZ+3NvChrk7MQLKi53WbT5/mmfs5qdrx9059MypD90N
pKoCpoi/P27tNP1QaFRDVlEPhw0AMc1QF3A+KRjU+088UAs5Gge+mDhn0+aXgZX0TijqgD8JXB65
9cz8JGeffBT0YNDquFM6FMdt0IZNPrqQzcEendnNSwXOoo1LV1oCJKnujKV//Um2uU3X7HpbvGWI
f8OIBnoQJLZG8w1QGupLAPIj9K4ZO/gOLrHyzaSpUhUqPq6nAMvfhHkbZ2p2vuTO25R0Ofg6RLyI
wN6mKI0X1QpRDv6I3nlR/k/lXbxBEAdmltVpvl5Pg3DyGbu1L/+kBWVWD00ySWS23FLDEzDFJOMW
UysRpNStZiBuid3DfPBfTenfPI49L0tR0qECORyRHA0/qgENp7bGvTu7we5o/3NgB4cTge7wDdfv
6mSHsmQJ/ktBllX9bIDkOcAGHicIIiK11Wcp7XrcAswzbrTZq5cEMBP7hKfMsQM2tl6J0z6d0Yzr
oOF/+R6ygiF0NEw3BHVPlIdLpnAwKy90+tgBNdZw8f0GUtYoYOhQUhFLkV7VbXgA+eHKt9F/qnjW
Bw+kqhCqq16McGTOsxieewiwaP86kJnv7mhgBDudfFEKWbyjncB2KEIJSJNmcHcBZqYmMFQL+X4F
HTDzZDUaM1wXUIhLMC4MOdSTEeKGR3FZJbpbXQsWOAvCxDITz4Rt2D8Uqd6nKDzVRC4GcK8tRM9P
kg0LkpzpB2jHW5Zo9/E6DD5lE+uWzSRbtlZd2DjKFvKZdmTak9XhHDZr1A5UbE0q8JyQMg31MrZ4
300FhNO/dCS8Ge+9klzWOCJgWEpX6gE85YG6R9+rBTad1hUoGdKCvx4gkV5fsdRpiCs0G7mVvFDk
J9L+9TZKrRQ/cA1rJpGDZj5fUH21fG66RokH/ZDpFRdig90zU1VTKhj6g1B92H/lNnBz78KuBhsm
lrdeMhnYATyWwRfUk6OpC42KxoYYtVwLbb321f9+hCwW/virhR9dAmD+YHVAGWpsM/LoOI85Ma/l
nH4KiDF8ssg4XA6N4UyDwjmH2NO6HUUHhHx0yu3UaNwakslUcGnbKg0eGU7H+YM2pa7t+Z8czd0K
DwAZt5c6YLhY9VV0uXn1CRpIuHwcOyHZnhQ4r1T+VerrKiusQ1lQwlk1wgt+i9pkoHhxO2A677I+
IL3hqqn63ocuesq0Sd/h0F4pKPG9o2tHLLoIWQdkQTNtM8FLgNBeL5vmonP70UAGzVBIxy2EeDfS
Nt0hm/fnBkhJV/N95z80XQxgpF12M5xIxzLtbLgYHsJPMsd7wR7AIgka/iCq9+I1JluN+niGDlQ8
FBv44btNe6R1Mpu+zgbKQPFSJspFb0MzEzFKBtzkzlWm7SVmaD4OOc9Qm/M6IeRxSystq+eConhS
yBTHojNofh7VvEROspowLV9YNKFHzfnLpDDG8xR5DVvkRBdBAOgaK80VoW1ihVavhfp9A3AX3hbA
R/tg99R5ITDNwT68r6Bpj3gNvUhjOh1P3hTe8ut2/K/mxMxtssrlC/7wJdo7EEJG0UOUSCuzLvSP
pyLRCsim4JlUayPQF1OjEQ5lknynpDf/+ozd6nQ8xFEuNZApbtHHXpy59yc6TNdGHxw/sVsObCTe
uvK7y60aqQuHV0nGbd/KBEBjLPIbvSwyB0TYPqdQBuwWgTChOZgT/rWAJ3y2g0Ttts9mIIYPqGWa
Fe0uRH1mUa36Oa1X3oDawopRjgKpxveEAQkn2y6T8Hu30wuUBhCV7RlGtmPu0YIMs+aqgyAmAf1G
ip6LnVyClQ6JUpGxsujUoNnQl0ivu03Wls8T/ZssGhAmlheWNLL3S5YJK+g8rvYDZvpCrNP+aO5q
q3jPbJRycL1144srsGAcFXl4KDOrjvc53KlqHJE9BeCRBhGAY+Onhdc46V2gKsNUvCRAphqF+TG6
1ba6J8YpDEapBp9irjAoHlvrzddz3Yp//oHMMOT2ZRGijBEr3YGfPa3hCYWOubi9wT1+yyCRhf1e
LkYZ0rNKjakUWZoPWLVhEOBBl9XWvoy30H67HcE2qYsK0gJvv2Dk0baHgxswwLUUCfRFut885k9r
oQz6JtKD2775Eu3nsxqSfD83Dz5QcaJ2xIwMVuuukSDk8eWCx2QyN4iBuVhFZjRN9XpxfYQTjATM
8/sLRUrCd1kDRZAGndHHinoYcexebO1+tX/wjdPQy7ukIRNavcFGnY4Rt9Qiz1reGrqAbygODpXT
QNbJAmVbMYwLvdJQreR9gtypPPj1VtThexsLTzdAaHRMfZ9sWL9Ainmb8D6U38RzgVx7TgCVvdGt
SBEWwyQdV08cIPxrRROAa91UCnScSdns1CVwSHnh1XRCAOps57Dqmsjhet3IO+Zh+dU+YTvhX/sR
buFJX4iVu3rdkUMWyMrmiuy0OWUx2mhShfk7ubHFU7DPVYbVlE/jhU50ynf+vjJVxUlF8uHShfsP
vE++KABflvhc68AlUH39Uh7Iut14ibAI/ux0lSPlEuwhqThEo1Jtz8cCKqMxeGRs1eQYSpaQ7o8J
6mqWWKmOihvoX+xoL5tHLOQ6tLFDSeBl/oEdmJW3etw85WDne9gXeRGYiz7t06FiWtausxNRw2Sr
ouD/EgpIGaiMgXr3xP5u6OVe7ZIMHlHdKYIwVt5y8H44YddzI3m7Xan4pO0QXrC+kBCLI1TyTXcw
qDcHNeM8HM0ySCa6P71L/d51hg+YL1cVTO9/BKbwxrYiRfvAYaWiHo2zrGYP/cyTBPNu8z6xJUH7
6ZqMhRtVo4bcQ7fqA2wiYMZLDtlIGdQoWeINT1gugSHPS5ulsSasRgADe++696qIWDpBzfgesaPA
NQkwtnD2IVycLZAuGVF7+lPfcCWo90FDxxAOqY3PIcW5K4WEGNSJFJ4K6bWLLR3TZubG4t1pacw5
Mx+oGPQjYsJTpW68L9+sOarpLI6A9Azyf54OHMXL8WfpWaHDiZJX/0cbzVLwPisD5Al1z1CJx+6I
p3m3yRWe5HE+7XigUvrm5zfd5r+HVngciIXu+mR20pRjvMKP0ruiwbr3r8/sFQYiQB+GsG3RMDcL
usxXb3LorRYiBn08WpNDJrmlkT7CWkQfIX2HrD6kNdcYYnv6eVWY4NR1IO4zqO9DgKLH+qrGdJ+m
dVF+tjLpT5lpyV1RxZq8ccvL1XfEpJBonszJBept1Chh6wtqzE9sLcBveEceX5PSyvGqtoujW+Rv
/ZFjz+0UgXc1Yh4BVfOvtxubrXFBz/vJzEPJJfdGDn/ENZjzHtfCt9eZXHyAJ1/4qOYegK8D4aY9
LuQjw3uIK6C61NuiYR9WgNbr/ohK5cYeuFE1IHWwcINFf2pAEjmh86EL6EFkF6YCyRTvJCPJzith
ioxAeBZ5mNcQ8x1JcP0QJRPIeoTMpKqX4mi442FPMoxricIA+HvON+OcLJ+xW5dU9TJ1kk/J66QB
t2qzW/KifZqO96hn8PXEV9Oxwhmo8pOVScvh/8o4Dm4ZVDgwH2/j0q4Wxdb1Fju6wLlYwypl3Crg
VXwPVIe7Zko1Qzs94QFo9UZHZcgRnmP14BbL43jm0Q16pxxhi6bP0IushxP4fU6UgsfNaymMgNY+
qNsQxH3ZuhZ6lMeL/lWS+L9oqZKftcAQrCdezDy86a/4kdjAFZsAQRZd4LkvxqiqHmQUgk0PgX3c
UaL8q+U0StVieT6Fq1psc3P5+kawHSKfuPG31Nbcfa2tmEDzpD8VHvDTqU01fjzeW2j/x69Vq84z
1L2T2n+v26PqtdBTlTSpW1yvU+V0YtK0we5ItxXB6v5dT07HC5IkA/1vUdnE9+lm2BCmhx0DQmG5
vjrbNI/4zSaW8qeiZeXBSwOxSM/zjWNrwY79HsmCdhjGJPia8Tg1ekKVYrjHH8or/wifRCKkYMeb
BWQM1MFBy4WBLGdIaVugB6rERARkwJ6TJzOsXS3k1cd9y8LuHdyDBCETtAgJaZrW+7n3APh0sASB
eIEVKZrSdjbV8SkUwthZqjj3417utaHmka5wnmQUDlEulwBV68ilZpCkTBB2CgNWWbWUv2jF2DA6
QT7m7+eWQVsUVqv7k11bougoyRzZJXN6oSKiEeRpAW3M840B8yVtMG2cgkGgVF8Kk4XOupnrl/mK
JawMpIvLKhiH4Zux+itgXWm5+sZbBbffdgWZDAho0KcaITNFzVQ2ttIW1wE8CM5lSWpqnWqmkNJu
pPyIWv1JJS9EFkOHjV7StLhy5UHVIab9sNyz+QLPtGCnPFbd3MknXBLOkw3tjOTUBoJTvC4PZnAC
oPRF1kYCCa++8+NaxvInMpr23aYGVZ/xW1KTR4YbYCprXiSlZAjDflLAG73iNYpefpAzsK2SjvSn
Udhpw2JCZaM0JQhALo88RWgwvUjW6dAZl9PHLKxzSF2Ht51BiUXEKl3d8tK8PR/Y/RmTtFiuXJ11
8KYdvZXy62Jling1+X9wIvdw8ZY0jNK9keve8+dGHADXm+S4lOk+w8fee0k3/25Utd3sX7M15ApO
+rTJ0sGde7hmM7m2VWo8TZ62grvPOPBTHMSBNqLaujtDVPpiSmZbIsoyl9xcDI2HfzlrRZvL0Z13
jOPxayLbcCTpOgqJu6cEgfp1/5VrY8TEXNQv+riKpaM+jOrOQTX4QBL4EIXNTuO40dJb6XIVmPCJ
0r22TONetYih8+DFNfx4eu8L+W2fki4B9jPubTwRZC+cS4EBomd65t++yXh/aiqroyabteO82pmX
Ioy7LaH0MS7/iPO3qXdtUIIj2eKo2wmN/PDweF/I9V63Cas7ckj9RO0wj+xLb4oGaV4N8LAn+VER
7ZFYLDLcebUt5cIh0+27qwe3ub9WsT1GaxEini30vFkNchc2UaHfthYAlPzMa0OdLU1fu+EHXWIP
uRRhHZsLyGvxKTGrFxQEGpviGQIMe6KK4wd693UQ6q5IgGE+uKzfCVeYfN0NHrK+mHpMRxwr3lOh
yw7cE62B8qR/5G1uZLbgbfRxYSreuK+9NsQge6vHrX9AufJO7jwhyEsHVmpgFwpcAbc0rDff6mB5
IiTyecaA1fsDwCWe/LmhKavhj+sDzeUcjz5EnCJy/fcwGT6+uK3hgdI6/R+dcanv/aWVWUVXJxpk
Xqj64xfOrPTdLyZMwO1DzG91xCTUn1JUO/JoS/Hcv30pENK9NGIIERHPQdpyTc0EEY0KWEQKI1Ot
VYzCOIgdPSB0Y0XbMqhToslUtTuUloHxyZKWB0pAZg5Sk7tAlLi9sivKG5w4/jxrAT2p77bLlBEE
v4sLunopnIYY2KO5PIpEoqLh7m3V2p/GZltLQRnf5MBoxQ2J01MWedFV+J9IhKjyRgxH+KjtBp87
vKxkPHKHwX+85wtTKwsDIaBmmgO5XKeHBYRo8poQ6TT5xMRaxpqcL6GtXU0AyFMNOSSDyFsAMTBM
fG5tLifhIZrsYkC5+tNuIgBYZ3QU0eW2jnsdqS/WFwJHzb7kaHdFhtlOCxZJ/wijs+xhUNrMKwAv
+iuCnX0DQgVyiHyy84otLLTlwxwTeFRsfbVKg9NNiqUYM4c/YG8wz7pZOuxcPRtRm91kkHPlMvVu
KK8RX4mjxPT1Ojz7j+AiJ2av8Yqpkqwyx5HAbh4Pj68ep6uWqxlXCMTo4XUxjGlu232iBaIfDLZK
I1M9E0flwWEvL8VZnlZw3HOXD/Z/jKu38mFxvsVsYE6GkFy5u9DcRqtd1IR93adph6y8Gx3u/VZn
l8586GrbECCUGo/gghA7Q7z5GpwVDfzYdgGzcr5MkpSXmacczqgQNH1RC06oUTrv3Sw9z1IVQ4If
LPY6PmoyulDtcAP+sJ2N2wZ+2tPBTXaJ11a+aC7Yl8pmoKzsxA+niy5/PLJakUWiOI3ZlBjIgs5k
zwXWsArZmN6IsFLYF21iRd9JSW9sMz4wzeCntY43AMOk4omNfWJxAQSXWjFW25lwqGrFJDgNsd1c
hn4Ns1BXJmdhk/KaGdzBzevtxazRPUtcit7ks5Qf8qRwfvlpqNI7gwsWhyaZXliEJCDt7paFgWt7
PQ6pYtaWByKnFQGRqnMq0QBPFETVGMqwgMtbqf/PvBxRWWCbgFEc9sj+nAOX2+rwEU9+AH22Rba3
j5En7TGWA6xxqigvvWPTM48wc7qT2RfcqimuJ/dUogZyMAsUkdJM9Ic8hAsrNRPF66mbvcUSG1W3
S+hl9or7SNO100oPHoHpUwH1r/4a9qnFLXk71wUYK/0zS2zqwWI+QcPAIYDwPWVLRvF/nQWl6viM
4uYEHDlHqrogmzK8UFR4tEEOc6MSf2sPF4kSbttMAicDj6rZfptNfbRrH24EgPVx7U4uW07c80jJ
GjCh0j+4WQnilLCzy12MmZy/phavbJSYDwbRh8uW8eoasIFH8fQyEI6xPhBIhPFRjx8FcUGGRSxm
/TIS8MDBIrKEXbVQqeEPoIMaVtginLnC9qcxP8LcbcFKQuXYKCfNt7qtKHyctQc7Eh8/lG6tNwjk
mXjAYqcSnHJOaplHmgsXdfRuNK6RjqHmhtMJEiQ28s2tkTiLk9KuampPLnMSk21FOYpSvVSdPcsf
961CKBaf6nz0vwVP7Oo+MRhwNK+ikQVDmuvOOPnvsGCIBdp7cjSDwuYNY3n1004WUyOeu8bHEf8J
QFEsUNFbu3r/9BMEkUtWhQAUuncTyfl0o3cKNG2vBiFxGOAWYCeImn8r77BvshktL7XJZhi2SngT
JrnHBPgAOh2oN4Sf0AUps9oqUECcQRlYivfq9cjRWWjZMOg+Pyc4UdeLH6ZVaT6naO2Zlb8EWtpO
7o2Xj9JWzSj0Hy/XkOPHO7QgAT8xxdCK+S0TwI1xQXnp3dyfu8C+RWPblKmq6yd2R+QrFpx0t+tp
TJzPjsLnJftHyHedCN9yHjC0xtpMNEO9J6odIISE1Cb45wTwWbW4CkH7QH1yYGMK+ODnJJV4I7Lz
jWzk7So8u3ep8cOKFHsCVDW2NhnXl0uXsuw4N85u519+fjlnOLf5KHIIbjjpDcWkAOom8CoLJJ5g
gwnnG1SnqWh2pDgyVXXFczOu2XyUeUV+pjJkWJVC2kQLR+L6Et3HSX372gcn+xAecJWYL1dr+HSO
k1t+0tBYJoOc3ADQhQfYclhun3pc3goqSUFU6nloIh4geWmoh7PEY6hIDw+ZW6ckVjPRhNmG7ycV
4l6Fdra3dvswDqBu5j3ARTN9WlaKBlxI1V7c5JLtLoXGgUVYUt8v9dGpcIbHWMuxTzKpKgodwReZ
06BeY8wo9DdROheGanquWOI8GL0+U3VICcSrnG4CnFbQDHAnyZ2ox06R5JgzVkYff9ZZfgzRHYpI
8NbvchjcnHzXBq+IsnYsG/OvvaYsJvPR51FvIPNTtXfglEIxoMsV7Eh5tgIHsnyLhpf+lu5pm37j
dZk1z2wrIqOacloRbNF1g25DgAmOZiQKclSY0nmQACWgM0KZw6mswioxwEtu6hcPXDwJvJccmQVf
GkbO0ACdq6hiPvzpGWw+8Vd+beyD7CRDL50kPCga1uELXoNLGJ8E/o8VpBBbhUJVr8Gj7FFX/WKy
D0vEhR3BsofRl5jwuRqu785XXDYXVKhjlkfII9EuIBcc4CF6HxQ+hkqfu6mulbV4TpB/uc1NdyL5
/gGU5FSdeXxPey+slW9liKEbruEQ3SfeD0V0O7GaHPAKdawxeSJHneHJE2IvFS174zMscfQLGISr
eVnDm97F4k8KYgTCh7tPwDJUciafhzw3qbliUZFe6MMv0VgE/xAQAzTYW/XxEJ7eZWCoa1dLOgJ9
agx69CAIq60+gqYw0yd6qTkxhe+i3td9uTvgtFbrmmflYpUPpPmLLshyODh+naiSMvFIk6sO5mwN
zz+7r0FeXGx8/EgbqUQ7MSfm/LGlZbBSOdeKpAyqhSYA6KQK5g0lE/MfDJXVDjnTCgmVr8dXrgFY
C6r+mwh9qCXNCx1lVHpMqQohKhUGvHNC+naQMr2/myV0LwOwzCWn7P9slOUcOWRQAn01OO587k/K
Oy3+aZx7QLDIkRto6ry+QZ6miYdbQkTYMIVt9LqbA99mAvZ7jetbpMX2lf6/zC9RyzDm4G18R5Eb
SrvyYIOpltwC3Q7cJINvGNMNXy6w5gKvdAx+8CtRIEua8aQtLamsYJde54mjKE9rEBIv49LOAdR9
2vcOpyfMwg6U+NzjqxM//nQEqSJDfqzHXvoFZqFj/WA2psep/MGkGtp2bynf189fV0pd441idQ9p
udD03c5ta2pHHsi26wBQf/V0o395H+C9E0iTPgZK+CkguvibySswb6mhJoiKPjllfwIerVIjWfxk
WXrL0Se+Mh2mO6knTptUJ915W7sARzJ4VkysOpgJuH3Rn9ZAUyqXEZfcg57EH6DjxQdxkSW5LQX5
IkFvUI50fi8wWJ7NY8l+VbhOtO07GEV85qmjQhbu2YvqA15ZjcqngOzEgPtByoBcNdP3IETjUFSi
vI6q7yuSKnAhGFl16HcYTuUug1oV9lLjF/KpuVpRztVNAeLh7c9+Bf3vuNsj5nS6uxzynsn9CgiY
GIJmukFXnzLNn5BpDMSPad5cQyow4Ww9WgpFn0xfLgFu06Voanx6UFhB/Lsnm7y6tMd490nOFE1L
NIPFWZGqRIxtOkyiilSJ3ACVifRnwk7F/hl7IEowPY+HUr3SW5If8q3sGXS54WRR+JSE2Uf53zG+
newJYnfVUCXHftLQy07bpwaDor8d7okaxWKmiCY+0ti7a3TIwEeh4FfX5p4rV0vVLiB1d3Kqz4eW
PGwOH+G7960c6s+qbQix/g9pG/ySj09nPrKwF+GhGSh4z31qtgPH9ezX6OjtopQtR2ttEasv9sF2
ef6AgoWBOWUprEYD8z+pQx4WtaRQOsLG+1HCtRBRr0HCOcm8j7ViwPchGvHqZFpDFjkYaaA5+1yn
6nUbxdegFzAR1HPxTU+Vxiru4xoWZXlt9bCfkJsB7tgnfHF+C+AVWEpq5oWeayoJjUy5sZhccLXb
6UrPFLQuWZvsdPPHUJuY6k3DtRwABSVjEwwFt7Oi5wRrcuu2VX1xMZ2zNBGF3/SbBR66IwU7o3IL
6Uq7bPRlE1EuaMFZgSDcErQZFKhJWY46fcpOPH2Z79+q/NcHEmO3u/bP31OUaNxZm6H6AJDyAd2N
q111bhgPrJiBirHzzbG3TEFclOsGePNKfmag7fSddsqlGUGWtek4kghnQlnFGeV24hS1tBG5o/P/
natrww+zaLYpegq0tkyh5RjhV7+KIQvBzdgPAhG4HQIW3Ebv5oYphAkoGQtZOJ5ewtqPPUOJKYn+
0xtK8UZpfkoM9TyQK/Fh9mnSXqaugQoFJDRrDknai3va/6jk3D46EB6ULESVpn7vKyOcs0ICFJE1
H/xVoQD0HjcUz/BuCpk1Vs1UbVYtlDzXvvbxYtTOTJQ6Upd0MwdM/kxtBpnjjMBudYhL5QMLZzlN
ONLDcSaRPBNLhGwbkjIKeN3W9RRcHvpHo3BkKZfjOlKbKoKNLUFCk3lW6JGVKYKDUvBihjjNtcov
XCC833/4vSx39i+9if3PrcxyZL4IzivpjZJgJlaub2WoQw8sHkDDkijurImQJIwXLfz+3cHblOz2
r6oRgLrSIvudnoO9/VA6ysCQ811wb16tIqeC49/2Gc+s9ZGbrC1rH3VLDhJTFMtmXaMFuJzA1KKk
d8mhkajvAe78bpGPMkP+PWjqOf11o2N4XKza4FH/fnuAixamtIldhQ+ZM35vV3ahv39rpHqmyAaH
z43dosESS6UYNU8EIfIJRQ8ZrxMMGt9XDlnVx/WYUySWaa8/c4jhG2VDc0+pqq4wCKBDj9gJyIlh
ILyy81CfR6UixKxR5Xr7fJPLGITfQWdzHdfRZv3mKB5aB1l0za3z1U/HZdMyGeZa+RcothUesETQ
FYzRqnX5I/74b9u2uwDPNBjmiXoqF/eOThq8uf6EBLd0kc/FTOgR/Y6whSWpiSckPhOm2jObylfu
0FcciScJ/HJ0voQc3jhX2cf+UeeUEmDkX/dYBptMYnCNkvS1dlXGmawVF/A6TrGGtq3BKlUa3IaP
WRrpXWHslr4bOOwO7uIiX5mw4Ex/EbjwYj7ZY5sG5apK+a0J9ZvKnA7zaRTsddpgz+x0JVy99YeD
eJTJqnRRLpBlhG58EWSu73iKmhfqFjWvB8Vf3JiDZJUk7aO5uE2sf7VV75vGbykBQZab8WMQQl3h
OTG5tY+uoT50CN85bAZ+k3NHAd/2CHH7eDo1Ty5fc+viFQMkHREu8FTGUefl4Ej3rWgZvv/cQGEc
J4ND9ppDaBGFozlqct5KNYHWofHWSQy/1+aP9lc0z4wv8LphzT7zflCM2xzOOvuXgoBF3L0h5/9h
csre4oU5IbA9QzqNLa/Dv7DVgoPRFRk9lGtciAqhUtSKASVZUT6D9Uvixf1v5InUnOPKWaGP0uVE
dwA1j0b4D0A62MgCCcoDCutpFzd1yJGpeMJH75YI5ZNav0BlbQJmL5Jt4qPtDFWSVQ7j+Na+UT76
7kXyfR8w6M4eGobn/5aNUUBpyq5kBaWyDMFhmdFCg6HR/kHM/rSyb82AUgZV60l/ngaEBrjdslrF
hqv9q0MKVFhQwtGFyMyFDcUEOc3JsYSlXDFhSbgFZ3RVXEp95Nzo4Pay5hCmyjJBSGzrq0MkYrYV
XJsoQvV2AzcVuQl3rz/NYHXSmcdWzu+6xM4MUudjYfH1+ICORagrEqUAX8RfZyCf0rIEJ30oRjcM
GVSS91FdKUnQoEpbn0exd2rUIsfMHWoH7ejEg/dROQP/Y0gkf2jI08aLqI7R6GeYkbkT/3sLDNHt
0/WsdwhJTEDAyawL4BmxNK1csEk/iEvqEyInDnbQgvqjmrJKuocpZ9/nIJ9ciYBe2yTb1yZ/7j+M
xrAEtutv1620P1wmikwAUKCrsXHF4ssB3gnR6ipgXiRaWFaVXhaDWs1OTJq0LtwPVbie+4LAPC4r
YDhEhGFAgVjJvuo5xj+wjsyISQIbwoY5P7s8gvrptQSKMFoLaDKhsP/pHt2yjlJBqOrZraPYuDoX
w8xcuOKTl51zD+L8Oip3Y1CxaxF3KrQwkIpVFG2hJnN/PmwZElb5yCAmt/cYCcXYxSMojEkoHemp
FF6B+1vJ5PRpCwDEfRy9gcVFMRRH8NV7Ml/3jIXWZHPcMFlGLKz7mvEdvCdVwwyZb9F/rDiiAl7z
xYkkh3FF65Z6IjskV/g0pdrPA6rD0HqHroAujPfYsm9y3rCL5Bw+X9ogeh65nLWCHPczbRs0tu4S
DUXPwacMsrshTZ+5RoZb+W6G1WtyCMJcfF+OCRX3lLb/emvHq8Ypnx0xEI/FwbGeOza5PlDdTaFq
VuFRxZ1Ah6RWsyKefM5jdQZFk8FF2aOpkSUnjtRoFtPsd2z2jNwd3T1wzNCQvbonxDfAMjtwkgIR
yyhExLM8LCOaDgODVPSJF2uE3so/SCYbpjauMQ2mZqrNNut736R9k0e0vZzgsc0BdCJCcLa5rpT2
T1LeFKNckY7bYpx/bH1Ytt0f1mll33g7HJbLCK89whloDer+iEAaFVWr7Phl8Ms3CpS/Qsm0JY/F
lTQGwNGZR+ePF4Li1fiDVbUw1J14BoNFzZurDJgWM6z2l8Da2xX3rrhT+R6w6G/3c0E6nwKPDCdq
FS0upjoXTM1NaSoZQSC1chTqwO47cyhx4pxIMeCrxrbHZvBM3aCwLyVZ2JJh3X4GRJkhg9Scwy1y
R/+ZD0NUcWX8aMlFDsnfAiVBKJGCzuZux8sFWAjQBFZwDI+kJeRY7GwFB9Pl0wtuTjTHC+ZnD42p
F3AtZH19YfrI2kRPfR4/+tIBkCMAkeS5FVHSjjhr90CL+KZ+PEoRwB7zNM6nxzDxxqtN2zivHg2w
KM8HkZMY/Fav4rYR0jLmc6N7EgMV4+UeDVzvceIpITxheVxecjOHlcaP2Zv89MLKHbDB0KL3/o5H
c+6md7miAxxmEo4j0RXFx7b7Skwvn7Nq4Cr0WOxyBSnDjAyl+soLwqMJk95mHQClYzWD89xyBsLl
AADv5R0fEsAABScRpbp7DjneTvzToeuk1LYKGu63i4If51vGlKR1sIwUPHBvdD/m9Wyuk/4mYCNT
yRjrm506DHn450Vqg7T/waTbp+TVW2YVhLjafK3MfZcF5D63A42d0q3U6fzP92Qz3nkSPVUbm4wE
Rv6Mphu5zuvg1JLHlhNuDfXGYwRql2dszJDamiwnwArToLMXoM0CzIlSTPn5gmJik87IGuuJcE2h
Gz90MCOmV+EaxuN5b+z/qvzDhcdrXoWVjJeORCLwvzTWEajMABwFnqwYdHMMKLzLyOW0ELJ+SGsl
I1dEoWDSHDxNe8r+g1bKEcWeI4AVxQ4huMONUBM56JYkY+G0hixVw0gVCNSfD2RnyTqty0kw1T63
k/CF1E/axGj25j0rTz99IyoSHKAut9gSmdrTYZWxdlfdDEY16to1VRzmKSKgL7hKtJ3MncLOUyRA
0aVRfjGNXkF9H4+/bqeV9LXnKTxKVACLQf+8G5ppkOLJnEoTjR0aiqvOBkkbm0oe8XUp+WHjRcG2
8/fJRMvKp3Pd9wWz9J8a9hbPhbRQ5qVR0R2bbdKBiRpiaObNpJhfhhVNr0KVDPs3TeEHIxThSLTl
h87xyVGb7d+wZPIDKWfQFB0qMddv0K2pkGd+L2i3eNQsnO58C+r8uL1j5i79L7hcrGejY9X4Wffl
l+H2opVnVDcJyAUL2dq1Ht4DI3biYgiF6gygTfMbF/c9sTWVXhf/nGdM3R7c5vQuhFDiY0Mj60oD
5gXI5S2ZVvy9VaqLD6Q7ptIhqqMvlYB3ISFFY+xZOafc8tOFLVMUSyBFaie3xYHTk72n+mlSARb/
pDMN8YqMb/dlRsRfmTA/EF29T9FWZp+ntFALUENMRJR2JAbZBF5P7eoDZVBc4T6LMhqOrcXN4vU3
jFS2Tob2JWmuqgzffSppcVqEwRT9LLoFZ0dX+JPNa5dI/SAUCy1QrrExhOcBnjqTdAauc12mIjwe
ynjrDa6RvhZO+MNnEujz0wKyklV5H+ZzPK4mJNBoeBDH7yIJ3O34U0Lf7ZJwguCuPNGKkhMhpO1Z
ThklIVGIn/pzHmSPVhpJSi8X72s124JtfRDlaqgIfRwvV9phf5hwys/5hbJYs1vQQTAGGUneqIVt
J9N1cpUo66mOE8a1os/NFUDp3njqBHYE6e4MYIFp5PLdh6HbtyNBmf6PXT0S9sCZ2a115Q9AyXiW
EgIhyrsieXmB2T1SFibgQeC5pE50cwpR54Lb6azgTM8k7oMYNIPYzr7ChO14zc+TxX/UDT6W8+cY
+SWWvmngNkpWrDzUlzKY3ncpqk9IrFJiXE6nJNzSNdcxnJBxVz97j6QuxYwkhLrS82zjDfSUxBcT
4hTnlnWfF8JLJLXweSkxWZWjeMKmIwKkfuQdh/hKEhS54BeNqzskJMjMUbPWlV3L4Cek0atYcCXQ
kfGdZBCV7rZCQMFaGqiPSvPQnSHpvdwYVZAaAXi0PtxGFiI/K+0laEVrWqVL9KuOTnYkTats1jbI
I7RFq0lmCp8+vJnWHKFyJoB8Cc7dZP8N67Oh4jT7eCeKpZ+DhpqimNKPmad/vdcdTmQs1grIB6rp
PUh1CRonWHV0JXqrAbiMBbEQDYz9aGPq+8SwSfbktHyZawlezfmQCiIJSoRzuaBNtuh2Pq4OWTYv
12S8RXtHYlTWtcJSnls3SoIw5KTUUJwOFFlvvYPP20IyWGhby4IV4WFtv4VvAaadT/d2aYsQcmvP
7UPbmHIUVCa97n2Vk8wHjMy9tFJoRTUN0BZ0SGhEIYb5MoIae9niypx3A46hSHTv+PXl2Z9CALaA
avt8WqgCRzHUsqMdFgu/jMJGKqisFR8nQNnXJdK/LEACP4KQRmxU8s/RiIAnlfpN3PV69JSqaiq2
O1jHKSTXQ50oUblcPwRsnQUBx1mB/s+klwI83aWExjaFOix5ex9eDr9W0HgrZd5ysCXGCLzHacD+
9MqIe+PHjPCuA7lf+OdSySNM9UQwEb8FwO/Jmzu4Nq1T0JUn+R2ADkwg0Ih+TzMdxemx1PXM60u0
gBHcb8gMGWsludkQCzF6PKV9tzvWWuCKUtN9vNplo97bwE5Cq+yVi653vHDP5SM13UcoHwnmZhCa
3M3G+fAkQpliMrKswvxt00CLrwTAtz9B5zuHpbXzo6v3SvdtelfynLWruQyOLClMmkkG3yogZt1E
Zg1QTSvFtn1mo51a5iFqALzK8dh/x3Oy9lqV05W3Js7M829tjB+0Y8kAhS2aPHWNktJLzZw80n2u
bDriUYN/F50SExRf179W3/c72RflFqT2yp+iYD1fqYcTO8MAY35RsdkKuMyRc2ZAUG91sweFTEzT
6PBjUtYlJY2DWK6hb18Vec1aWbu8plIiojDV21cTnbqIWi0N6xqDFRUbwQOQUe2lB81WFqqnWKnz
GBa5XdT5cU71wPyjdDQXA3A3hM2Bkw93HwCefUJpIc9QgkJukj1tjyiX67TOA0YP8jR4pOsEcehO
DVDK5qImxVnS4QNfcpoVrToGpopkl/hJ92uXUFQI72qqU7/fz/PXAc5j83I6pH0NkqLjCRo9QpbG
QKYFx9v0278tdk9+gdkwLwste02T+Ku4NfHUMRskpv6SaUmMgLwukh7TEhHRIx6KOvVb1BFF1DLX
OM87tsY+Sx9Qu5qBEpEM0Uyf/FKnASw2oGplXwZN32tO34C4CT1QLOcV2EQ7KcVUsaZFnHKF/Q8z
4kb8VPjbB3K4hAEbyids2lEeGbbA8M423vGj5E3H44OmFCp9nm6BoGPnfXMObmJmOx3s761bW/Mx
uLZkb+Pmlm14odeDUYVWIOiPFM+0xi/YM2pFBT/zNIimb0uwUaOF4SiNejhQJoH2UsAanPMVnGyY
xjqmtH7UA/ABVNDgyKvOsm4d50JGuQA9QeRH2w7CTrJrvbPhauBMapRRGQo88cHwy9ty05PNSKCY
RQGCLDYZHm2/PT9ibZWvn8i8GhvA/ywIEYk0Geq6neGUV2speTSDIdnt8AJ8c9lyBCHHDmtFeEWi
8gEe1sz+x+PnSq2wECvl20B36OvrSVu8AusgUumvb0M8BrItYaI/sN/6+CLbCQFSK3Fk7MzsT6c5
0HOLm/8c+V3acd0b5FtD+IBojap9CQ6sJwv1GPIa37xzl4VbDbUh0CP2oUDwhVcA9q81Ijbp19Uc
kz7f2LwCJ6U63glShldP92b1QQ+gVA8VzlltQEteN025Z2UeDjoDVgEnAGEvmU/iW+PZ1vgLGIzE
dAEma6SjUAHTbsoRsK8fo+S12Q4Gk3Or18oLZYxrcUr9TUVAgmxsxorn3gls2CMR7sJBbPFWEOU+
99OoGQbIUMMMj7+58/yA+dm+8gef379VLHqmTCk+e7D3SC07Y37cUw+IN9yN1LJOnhYE64Ct2G/5
vAorWqsZg/qrmmIy5hTDuQaVgsMfs7iEm26kDglJRLdUiQvrilYVssUNqI9CAZpQfnkPzsSAU2HB
bz0oxsCv4Q+tkBEoe3VbPU+sBTLXMWOLIQIl48PuSnALHm1RzUdRIifDoBGNNdgAK9m87MXo01zK
eL+HKlW5VukQc80532wC2MMQsqUb7qREjZOzcm/WzmsbIZBjZXxm809bwTAb/5gUoU3rxQ2SEhot
HevFRk6NvTLJueAblvx0R4npqRGf6/WZQPnTcK0kz80hJy10eAfcHhEr03dmXR/W0a8oY1tbyoea
vfBTNkmTRoCCjjkGZn/BBN6DxEClH7owfL7S70e8JhOOaOJJfMb7tLvRqRxN70sor7w/MeT+E/Qb
+wGP3qNCK+iX0QRdln0AmqaOghx5XGcoc/2tw/wRfTTR6ajJM46bPNTwShXX63cyoCaCeY4pm7jw
aAKRuSAIr8i2pcFneOhndFiWd5vXQNoN9DoMhYUP1BdsBE8Ii9JqECnZKp0yymN12+qNFflBVXsQ
3dv1mWoqn0v8opjyigvWmm8wkI+fVHAxod/6Dwyy9BD//nNqp5WlsHJt6NQcupHbCz63Ph6AikIn
QaHY/CI47TRMD2x20R4svLnUzgvK3MMbyTQo6+fusl/CvQ3iGWCC23q8QYDRwQBgRI1GUMS6DuXn
RTH1cRMqvoRzVBmxPMuoflxzw49/E6WWVjNV4J3wdBg6D4Aozrsph9dJBvO5PdB+hWxcPszigf2q
YCe02nnxMD/zzzy4iNgT+SWvqBe6vIVYbVYupcS8mbdXaDtx0wbqMoeI55iVPdenXl9IE7jFryHW
zM30VCXRzc1LzT+Nh8sPFvp3CtzqmGyzYHUH+nIjd79jO9StRUEEIqZF9nzzHXlZLi/JG2J7YyqC
RQ6SXVMAX6c1eZPCUqxeDpt6sKGaTBviI9+iY3RkLrHV27NPf49y5kVtDdiPxvLZ/njL+wJrtxkb
LpgFVIGWOLrWyqFeFhg6bbe2zSOuzKSBX87iBfzQc8koJ/zO47KgSSMCNG+E83/5UDwh00TqVwX1
hCz21eKoJ0EAqoK8XoR9Cxj8nhhRz+kHaNq6pHFQXt73C+QvlhAQnLUA8gjTuQM2T/neVzWQQWRh
Wn0dhcb+pyqrf5xTjyQLtMzB7z9IrnZHxde05BGIu0mP5BT9tY6VwrzsaGJxUxlWoCXncEo11yQx
Bb+rJbQ9aR8FfqtyK/8GbBS5PQb/KEZ8WQjjxJrHbziBKyxpkcGZ6vqigec/caj5fj7GLUAdzuBb
a1bZwt2YRCr8Ysc/npZ/NbYpkMRa4bH3jtA0oh0Ab42y8TvpzPbDvCAtuzZk3DdcASJ7nU9OUKh9
HoNPVRjE7wLyaIpcxhlin3v9gXIeRcOP/CvDSbedWGWa89uvQIiqVMsx+U5cxh39ra1BdOwTswRA
fJ+sZRGT8sACO5N313XwC1IWqPhkOZ/PDv1x80gx3s4ZbEtzalipu4J1k7zdqQ1t72fkHJf7N/aL
WuWJV2Dy2NQXZ2ODKzqc3aDJiJTBfm+7J/rNcfUtZN+WIkjQTollb1G4H0XKqz2pGSDHVmF/+isO
La1qmFsCnT7/zrK9FAhpzksRl1Xfs4sAVqZxcTqmhYWy5oQ6VxSOaTi+Iq6ng3uLvUAXwK3bkdsr
sJ1orBeokGceh1oOVcDK/cVkiY+gGi8j5/rd7Bpif6kNHPV9puy49sN+jwE1DzT6kiCfZV6DAojF
gvb/mJsenNeuvDryeH4gNc84Z4NjJh5bZdKyTTiwxf82bKceig7fuCfWsgPOu0PjLkInYbUue2Go
URtBnyFWqu3iP4ZgWQ4bkE1+Hze6cnscUfXSk23BTNLBVCLn4GQiiKqt7gGPMR8Q+XQxLYUskYC5
GAIVynsnaKpqAkojbmLHA4FwkYoP/A60AXOpGD/x6LC3hxgSLyUMJhh/KBacEYwdB15D9W9UaB8u
P4jcKTkUxFdkg5HYvz/SpAC/he67NdKQo7u9BUqUB5LQCzSVcovcrmRCebm/q+f+urdR0YLJkFQQ
lSonFZFmhDxIkhkek1SLnXMRhIUvtZohzsWEfsfiMU9LRQzgwSU8Pq6Jwl2DOPIDY5neoVobFHiG
WYVad1DK/8tGMqupzL3NNHnNa2GsyypwbeYB7cv0rRDlA7ecgMg9Q6JFjlJKzQ9oJkP4+zuXrpSG
giuF8TNCCVAw09EZtTFKPenDIWUvvLWE1gyrr15EMG+5bSbAjv8owKyZR1FG6kfv/iTqeyEmQeyV
f+FimL6kEu+12rG69AKukFeocUKncJcqk4dZO0strSqcgBMqeOZ7hVioPfdBOtJwYeyeTgjppr3K
VI/qQWIXOpeHM7UZG3SiyAjH6F6q8LWvjcT2U9v/UxQ46fk7Sys7Vu5NhIHhrBzgneALlr15o4PR
tmT4SQM8obw8Z7vgl8J/xXhGN+lmOyTq7QzRNg0FNy/pBN1MnA6pJxBNNcg8ly+rOaSImsFQskvY
DJP7a/YPjkwP11dbEf+1RQrI4e8yTH236nhNBDnvVGzuTGVFFDpkJN4GnjOtKoJgEvkRzCgU3Yws
X123Xnvu425ybynPpHMp1zr1/xPE1EPF+9ybdPC5WBiDwfeMAYgRj9iFwEVzUs5T/iZnysBUq6gV
TmjPRaOHsN/0869z6kAmC3CJfQNCggK+nDGSoNlqJnlvTytjCS/XxDgA9qFYsew+Ksiz8imNfSBT
95NNTcjS2i+Fa+fFFOvxM9ss+KAQzAO3j9JVrvVBfWA+dahSYDeWR7b6G9LPkhY8cnMUzlUmGsET
Tn7RJ/PvJe2VtZ0Mv4Dask1zh1KxhL/M/UoAwhsz2gOL487jGDKKa8MhHP4YE2cj88xssuYT/sdi
4NVi9oxaE40j49BI+HYTonYStsVs0Zr4MQAmhbV0FrYS10RWHMmRyfeJJYVP3p7pV5KPhTLQrPdm
Rg0RIrmuf+y0Af0QT31BHEFQW/T79wLDPHbmT4IQAuYrPoXzTdAd3NconmulJNEKaLYnnZil1KvY
HWwwj3dwx2peXVroj3Dad+XbXp/PSXnYD4fLSFxEK+88YKPf3bJVDHt7/fCNmV+2o1DmS65MIXCC
qxMnOTVKcyb0tamY11lYfAEHWLKBoPZL7fewZwZLPhm37Zd5JiHlQKuCBq/tCSXV8jh0lRuQe9Qy
/PDP2JJ8RuDQNvHSaIZTZbJVkpCct8OO4kipkr9d6Q4saw6pJ/py68qcp51etn3pgaKfJBMMmUqr
tPtGYgflKx43eoXrrgyvzE2L6yoi7cVBzMEntX/ZR3AdTsCY5Ea6ImPq9VaB1i/wkcjhRRAEWZOf
msdpVRh3JeJD6ZhINnqygwbnyYNS2YE180uK2TuxXMdlmoRYi5rRvrCKt/Qdn/eyJZRaeGOKFMj3
oUrkJOhIf2ICOM5y5FhA0QYq8ycUzj3U4UibQH6wW54iIfT5MEtCCP3UQRDJIypODJ+ZohrlWUBo
mAiQSgiQ9O0UZSITXfzHKgcdM41eD78rV2NuEmqA6Q9q66L2Y26qsKtGhHtp0OXBtSURNSni+IN8
HygjULoYwCFDpjCedIFKjR17Pc3Pu/SgrHDrsabANuxTt0e2NK1TeYGNdAKp6Tc1on2tmhKEJaHM
gtUKeJ06mmw8+hxaroONl7pijp78trFa3F7qQf3ysMnV/6Vg6gGEEJEWPIRd6VLEzhfcaDvBUgiE
DdzQfDbiEz61cJfgKR0mFJPp1nUxRexEJfs69sOeZJ5aKNaCZFGPFy6zTu2GRD18l68ySruSUo8t
3XFOUNye3T7zZQhi8+3Wt/Hut0hLNO3OCxiIKwGMgaVr+6h2XM3ntQ6Av3XFCIN36SCrF/k/jB52
n3jwOJt232Pioa+zPaSTaKZSDtUH6WtB8aM/AUB8A4lt1ZzdjkP6g+qTGVi3veS2GFL5TnYOvQ30
gnyx7xHbe5RjNJqeEn1q8uX4SE6TANkxYJ6PLMK1zfF34Ddg5hErUrb8e2IH0aUXphx8Tn+rFIcL
yaVrN1+bXTSXCbmsE8/3nw0zeptmhGN+V0Xt0XJHrOUpolF+IlTA+uKsX6ZWnbcyKqK2OA03aInH
TwC9G1PM35q7NCzDhRUBYqIm5j5JQLj0EsBAlOWLz1zGbCWiOLuhBKzBNyFC4sxt9UHPdz5KAGcA
4fsgmOcWT4LIy51REklqG7EemahpUlxf3fEyUXkTSDbkj5Ec4twzeYnYewoGF+XWdKVyeLSrXfHi
f0Wfj30rv4xogsiBZp34vedSlrlluwpPh5Z/FaYYjWoKqxv+5jIsU8rQ9U2OvDFuN2jwVAiiYVJL
hUzqpbMY0GUXFaexNZFr3Ah2E+XuBl14hyrJ15/PUrC8tIqah06kHwXu1Ox9Y+8BVQrTXlsQlQXR
kk6um7CUbSuzzfnlPQiQGCB929omgZrSahFfkpTWIAMQL1nes1zR5Ezt7MyZKPV8ILMk2IQDYtE4
t3jnc7AcqXm/P+PHKCQ+O8ccTJOmVkpSBIwftAtAaIl+QiTSdHcKrUZU9bJXBCVVcydzE2kfCenG
J9rbs8AdecadJhVUIBThtu7kbc3nY3qVQ2gFmZwXRr2CLcqtK8NQIUA/scM7nALee8QQDX7gxvah
fKMajhz2Est5qwbbQhsrkprDbqslL21Jd2eLxwOl3USvokvX39jhY7wqZ8hIt5cQffMw296t75Bm
oGdmovbDFVHnJ9cY88eSBJl6z2c6aW++uBd3LI2zrCnOGHSV27NvIzcr3pf1rTkxzwNhxrNGmRcP
y3NvTBJnhRHOTgz0EjiPU2cyERQ+gS/zBOgjLVPnZSn6MAibl3FeLBwThnNEXjIKvL6sFpEgTbFL
GaqmSxRuuM567cmHvi/FpCJ3+9BQIQnHxfAEJTEKMvK1XfGF2+AfTQpRc7unawFTH/en+6/2duP3
DOPfZu34D9K9D3LFzRn/ilq9R1i7bJY/6/Vsob/DeAssC2mzh121Aj7eYScsJZ1nYGnqVZ7X73uI
TALNnbRPiwR4ngDAIEkGdyVXBhRHruhB8uA1uwqz6jtvpgZ09Dg/qjnnWkb51nMI6SeQwwYOdcTV
J9KDrXWm0JKufJIO2BAfTEfLUNXtAauqXoPcZkd5yQpxEeJEtKObCShWbPHKeAVSqPsYo/bd3oZ9
GlpAbBAt2YBagbceKW1ZbwtZNjogM5qffRLUDibFQzAhqQA3pBj48o/e7fbihu1r01fN8CXD+Z68
Pc8LPd+7Zh34zNBYyfoJBwAsblIsT7p7n73ykZ+aZwIEtLmBe5+ks7d9akKrrmy8sEuUke6SQ02e
uK1S+v5S5yP5s3hVOGqpDRn13i9bS1x1tNpm9cXexZ+Rnt0Na3IXFfv2HAWvnxpChhbv/5ubUNV7
wYO5wLaQJHLeP3a7u+iO5WjQsZxGyMcFCrf3R/CidYr0BWTvI2G8KhZK2cOtjk/V12lJB85hyATv
rczU1MbKFV27RgEv7OE4gC5xElc38D1rqiCWv6dk+qyGUCirPJTjbXlghp6GZvgixHdEVxtjBxNv
72+JAE+rTn+rRfSIe+P6FF+fI8nPIzvrrdT1hGIpK9jqXaxpasneeCcbWLSsVlnEnAIWPs8POELL
h5gcOttZUQWwjv/iSH3DYjDMzFlZqpeCR1ozZS+pz8VGWiisX9yWeQbsIR6tgI4kO29TvkDqbtO2
bQ/evEP33faGAZIswjvFr146AoZOVfVYHhgYz1aWDumO796pbmta4cENF5OtDPFU8p6amRISJn8o
ICDe76m6e+rPC6e0maUGjrZbeZ6ZLV/8EbD/ia7I+Nxx3ZyYEqdzzQgsd1dGSrc9192NUWYtnibp
o66wofULKGY9R9VjAfzvhdtGvMQdlbDUaAsqSB46UZe0jQ51uzaG5YvMAdUW7XQKGQ/i/adywSK0
DJqshE4C6POj2zve/kvhfA0xRTktz3bL18T9ialjf2/RZ+8flFCm6rgPNGvc+SbpMrIP6rZXXKA1
ATPDlzc+GiCmuinv2uTbjBPcY4PE9HfPBTmJFg4FrOGHv8D1oiuhH49yNMpQIc+Bg200VRoSoUBO
tMqPe27fVvAX5LKDguIVynfvhd8Au13cE2+ckObsjby1aGjUjwVueQdHzj7Gp+C8Ro7/ZUERNM3J
vz5my7n0hb8uMjFN58JjR+XpkernWGnFm/OzgtU2d4DVjfx+g3VfH1SqVUAMx0AHBuuYsxjtQ54n
AlUtZ5BPb+pLaAoBPxk59wh8gecDcSJKCMEYDJ6JwYRmMjiMFNDR/bRtDV1wTsQVcZugwdA8hIzU
Mb5P7kAxDneWJTT+ogqZWTrI9WervfjVp3Cfy/kG0mbXtiL8RJG8MHJiKYa5ENnOLzkXITjj7hLw
A/SpLa6S6cRX7k6d6+QWMJhoUzFXDthjm00lUGyClzLi3SxTMO7tFVoTmDoUDvA4eL0NtSTIh1wZ
eY4zjmfImApqfanYBRuhl/Y4hHJ6ydKAaQ2r3iCtNwNdFLgT66/CxDN8dRqY7ef8YT9l0aJUA+mC
x9nL4ifYsQQ0QUnFtizyb/m7TRkhKZ1/7YsBMdQMMTryHS673bnXtqY85thwNZSrBGPq7P7+L0l2
p6DihtxEBFafg1k0DLj4UDYOyHpQ7LBdBRTvE6Dx4TYW41U05fJDu3DlvJ2Pxc2qu2sxud1kS4Z6
GL+kRgpSOsPWe4/PbVadQDNb+CNAnxSShYjLOy7CWY9T9su4HSzgbgLc5hYcEadTfmyIeGbtqjhJ
7rEDFspJ/kSw+bmh26wI7wCMn1UnVPquEzGWBHU/KBHXJFRom/Jh3a9aJGZbqfgr8HlVTcRzzcjR
ZxfUfL5YVYbeSuL+8fkCntkRm8oakfK8/WGv897Krvy16cf7+FVEKT4+yvz3zn87kJ7NtEgynmal
UrnPR+hQvn+eJCOpmxEPb2tjAGoDMo1/O4d6teYq29W2AQ1UWUmi7Sd/LbRlWpgv1vkt8RFJz4GU
s8GCqJ3W7AaGMqzPiBhxOaqa4cyAJnBZo6rkRTQtVzjR6+DE6QQofXFJp/Rv8dqpNolD2o1/AQ8b
IcYgnDzQXIcJ4nKINBWDWd3l6g+ShR3uAHpLKjJ/REEASk3HD0eKAMUcepbUBfogHoZ63wPyV8Kh
0up5uPXWBwsITrDIBG0sm/ZXYFO9f1D2Jj9Vrm5d8n1pB3FSxFUu1APz6FxfRGVJy0fGZ5YaDoU7
OoH6L4cnkDO3cdXtGqERPx1HjK29rdKXFVOXuea93JSSe0GyK/V6Wrz3FhS1MAJH7VvE3/HAx9GF
GZnl8dNWaQ1ov+IwSnX2MBLQyjM4BpIZ88m6U5ypsHg58fGasbQ2JtHZ3hO+7TtNtDiSTk1vY0cQ
VnSutRenGevKS1QytbKwn0AONDvftkoU+ubqReFYn7MUv73ATecy7BzljMICgA5XBEvXAW6bJlsi
6t3Z/K+hLfYqB0mxfVdGD1fDYZEx6Ep+9O5aXdakzUY4ZTbfU1Hi+5Tlyn2FF3oVX+D+jRezB9mp
6jg9BSH6KzR7E+MvOt+/26M+yUvnFb5ua1ZbCOUoDnaYbvMpsbqrUzxtu47J2i8v+kYSupB6z0Ie
YvDG0afbdc6TsLQM9NuST6V9k7AK5A47rnsUUrtoKlKo1Gipw9XXlPOcclY3nb1aK0Ua2hoFOEwf
Oz5hgsj5bvQG1qZoYZhXOC/bS0taF/QjJEg8yzHkJk8AJz8dlVs31FGt49adr0bPZoOPyIg4cZ5m
SDzxzIcsf30eSwZ/X2tE1KFqPNx4NULhxdNY7Zn5YeqzQjxwy9r6rjzxYKQcZssFgLuQgEo2RDeQ
PL0Vp8uSLwyMiMg7OvUS+nD6pYwPpuMVDv2NfU3glf0tbX3fdmX8SvQx5m4o7mBhxa7Y29yc7/Qz
0ERFrheVlPZ9QlqhTTjHdnmYiFm6qFS/4r8NbUiKJM5G/QacKcyFVDDheZaAKlG1PL3EqDtM1VJn
0dp7DHobRAtlhhfbGg+5nMDG7YFfonTjeVkuy0/10lZMacMxjL84mJljTplB8DB/fOwK8MWnS7Uo
/0eZWKP/j+5glVjsULVuhC1sDAjF+UQ3V0WDgUQ5XUuvp1NbVmbAd5Y+qXPLk4wRpdEKwMM+aLUH
AwQz+D5rkzqbaZai/YelWaBSyX5krtY5eBm5eYipIl92qAhN4c0Ib/QkvTU0LKzWKUfQ2YT43gt1
rXy8NCCitny2coCh+t+7GK4kfQK+Q3i6YHqwfM5ihPLNwVwOgYj+Y3oK+3hYDnSiUhkgIzOt6Yqg
3pGDiSq84rLd01KXvkbqDBscOLcTuTcS1Wf+xc+RpbPJe+pASh+9usWDBsVrvyxgFzJUKXe0xVWb
JT2yXkJnTWIl2KsS1ZqoMKSjDtw8nybegFShWghIIlruCVjeaHMA92IdcBUuDLPmotg8Gnj4gEaR
tIfVe5ceONVPaJUkkzj90BMjhH9f4D2Wzx1H5FQpa6pQ92SosSSzzTSLPmSIcAv5PwClSw/TtRXJ
bRy7RKxA4+F04s2jowe81MoL2cEj0jUUB1rqcAdyucmPND/jWdVFNCk5VfGVjRaUMtG1xQUQboqQ
YiEEgEvM9c5PGlc1loCtr7zpECTn87DLCcpHquUxtRDNnMkjwAYinhBcdq7pL5Z056PNxdYKP9TQ
9j7uephjrfclgbpj/pSy9OFzf7H99amvehAcIz0/qRF3/HGEXHjlCMrHcmtZQH7uA+4RWEwY59ZT
RLIbVVLWkZNBx2RF24rNvAMK9n1b1ueLlextwyFmcemyDgLH+2vMfPQXdcqmbWGCdHe4p/GcWLtA
TD20A/To8DVHRb/xiOysU35BAJsRsZRudcqelqZmNM3zG2YCHj3wBcRfLbo5crXFmocmqVcnC0ft
9fXQD9TusTXBTeipky6yT9ICVMzRNpZjzxYypUolMSjkPQ4g76bL84FfgzM9HLWci4hmtJ6sHKDl
YtvG9cNAdTwC2OLrmbNJp3Q6faN0EUj1g/VLSYjvL7MHY5Y0vfkmdfxzCds2ViZabD+Vb3qjjfTE
hsTHt59dC1feQqH/FFjaPNl8BnMFZn4eRWbnQZ3rn75FASoqP2Wahh0PQ796xdbEOIT1xhABAPu7
jp7I/2eAwrGoaOkY/JvRGcalulnZpaIhKZV4oQhO2OEZuAeL7URApyebNOHy97kYn+yu8ohmS9z1
DJjR4eNQt1mIahw3901/C9MiXs38Ro5v4jlDd4pmFVQfFgnyWgCeXq40wP3kqJMA02m88HzNBEkW
DpdBJ+fZ0YYEAn7GM2FhYSIeke61aXnkQVy2e+f5fmBy88hMtYiTsEN5MyQy1oEkyhnnRFCaBKai
DlUD5IshIkW26KIIM9FCk/fmWYcdbqArc4ZCrtTOPVJhQkSumuPZSd9WqsVS2elEhGa9RDTEjKtx
UdPgwaPkhYLBYCjWQaLGnC9tMF5VD0ZHD87HNbvyYkGqGamXrgnd7CO76daQZfmecrTWPpf5wZOh
uWd4GmXR36LaraCM65ggzK3hG7l7zV4VWH0MrthQbaWrl49gPX9oYKfw9NkyqfX1NmrStc4Mswmx
dGeuapOOWJdAmRZdIfgHIcxmA56JnKGY+YqpOktlOrzMCG/jz8dx/nmMqcEDfFR8jbStznwpR+rJ
KFaR2kUMOOoW+nkO38058PF2xV5JaDmBsOIj3VOnWHnNqaCOKWErugQhgTNPKJ141QkfXrSG1WRD
fai2YBv1j/G4bDfy/oEOzcp2Lp9bukDIH/7HEnwFypxrJZ7/wy6O/VOb/aXVrxVp+EmzelyUvfkF
DaY5kXL+z5W4JGrjxnEgLksQmFDI2pzmj/KAUnAFrMcQgifMhzVZRqmjpVMjdfWfssT9cbe+JC6s
V55uqM/B8VknY/Is601Iswi41NCkQ4xJYRRpaCl9fU/MvjuTXY1O8h9bpwKP1tYnfgdr23SJgeMF
BLjk5PIu2EKMWAYIuKBlej5klqWSyLBKJwTQNJEfdcVBwOB64y9eeSo6+zGCYRQHipBdHnHO6tz/
zfhHbRBXXrHvRMSwvT2nlbua+ru9UhQE8Py3BfUTmY+SNW6Y8c/i1EJBGMO6jMPvsJlDvKQ4UUK5
yqm5xK13TB+97EL98J9oIdV5HqtpTemLGDC8pAUGQRsWVbnGFeG0t0F4Tp8UwwF2kCn7NvowI0ac
vQDncW7y6eFfSceh99sUawyUdWS7QditxfmZHgZwO+TiGq7pYxIP3uiFSysZVl6Jk2wyAypiDP0T
f+vpG26HFCE0sVFO0hA8wX7npRtEBb+Z/3bGJUWvlmYUDdWW1NeLhiHfZx87vcjktKZJIIyd2TB8
ft/M9/XHPHhbBBNXkpMWdz1wnIJcycTprlVynpwRWu/jMrFW1P2vlsTnquJMbV4GG09BKAUN7Jz1
zCgZ9iL9uYctoPQ9FLN4fBRwl6jwWoarkQs1avAAuFi6sjCf69DRAk10ZaLnkqywqrfsKRRkQx7s
2D47suOi2TZTBzQEdltJHw3yWzJNF+s8wVPfmKsZLf3qiZV+HiLXdDPksYZUWg+ORhD3yFqgGLZM
DSLTGBBdKI2S40MgNdUZSKWe3GrtHhslILGURB19sMiHRLdYxfFCE24wQHAuG4yjXd+5JgAjXZiT
1+FqWULMUUmijk4mQETjTt/RcV5cWcbYLzwYhQyokVlg2pm+RWD5mSqac02VxikMojdtOnVaRE3L
BrziQWr2GzF2z6rfkGjzAZtl2K6AZ8+jA1j9C/GXXpMmT3oOd7e4lt1lw2dc21fQ0k5xgiYilAhS
QR4cHqNuZ0Bw9mZOag6lTreqUbWUymVXIOcRkM84+85Kc6ShlHdxQ0DE0Y1d5fh8qAjtkEq8oyFu
IAvPsFKlcdPZzYDeXiwv/SSsf99eu0Xnf9jfc5rp80oBwCPZvYYoiDqUk2uQnCUSQlc4nppmfqGm
ExTZmXehFx9qqHPq+E1ZyR0+m22U2wxf1jZh2vej6qkyd1UPWrwHnv52ZtIUewH5O9Kp/bGQTYaF
SRaHSKxfYtpomU6tyDmhanY4OWUogIWdIMnE6pPS9PH/AYt61qRqh5rb5rFcrVV3aUcjDUn/nADC
0kGB1J5bcpJk5jhwR3pOQEy3+Kuukw2Pn+0Q+OdTWaXj8qLqhYk1U40/TwNu8+Nv0D+8s4gzQEkj
CfUTlIZxDI6pTMrFgW7OrLUm+2aXkCM92+Hkt+7vYxvGCpphc1Mo1d9hV26MK0F5dO4sAsNcSZJr
/kBxoXWsxuPHVO3RaP3MB/ffGMktS8lTWiuee8lEHdAnsbISYycWCQfJCjlJI+7RCdn/YsUetAiD
vS63FRCAXnHaBPuOXcsln+UhJyS9l389ZM3MdP7JneiLnVKJqzQCcmQDKYmP8z9o+ygm3p+6q4Fo
esH3nf7nGfAt0LDgOs81GaRV4MoyV92GGY9D9ZJsk75Ek+Pu/yV3ErZyEexitakUw3NMjLb1O7fq
WKwDzX64VVXnDhOkCcXIEo3Nw5DKtRB47NbwVevkVXHJvbqAPgr2GRh6YukNqo6XmUQDyATcq9YU
A6hk+h37dvXb3L/WyWNexQbdkeedHXuR3YsnDN3UkOWnnAJkmhbCkH4ujvxzKYHpVLEQ+34V/P9+
03EWhQQvTL7MX7Sn0AJeQRGULgjYwxdXmB3zeqaXeX0ARKRiGXxZGVetQfSczBHQqeWcFrn2kOf5
Ip5vPXB4o3yvYPFTqk64uptHQVoRuqlL9Ct3aLWDzTQzXwpBIwsrUKlWefm9FiSg38//p4pwrIGR
WaKjcq4tqBnIl5tfR+8c43iGCVhwTLdvnQ8BhsoItMvTPFb/e22tcKE1kRvtepKIyZqhReoxEz8I
dZt5uVdldlfbztA8CkdDqpcU/NJ4Qy03Kgu1D6HwsUlzxXNogd8wPeDtHgkYwYKS2FaappY9uu+H
gGfrag05jzjlE7ZYoiJ9Je3yXhO0ohxq0uaVhwfqL7ocAfAdMZaP9J3ohSrlUPCZ4StKHmQM9K/X
UKRTBGpd9GQgbDjVlwZkzaisqFW44+L8FkLN46ituz+QGCGcfiW90TD66+07gVu4NrFk6hbJZXK1
VQ1TEyb5JKCb6jNSsTNN8/hkFVPnghlzqRiUygufxhqjohg0nO40YCkuwBOYtKL5T9OR/gxE57QP
GNWKbMa8Oj/MrV5w72ioWyf9HkRbJrd22c51s6UyiUxBKdxAG1ZlTXZ/PC7S6AZVlKQRHVwVbyV8
gQPAbeg4ZljZmiPkrz5yIBV1N1N/rF6l29p6b59+HmPCycw+UXK5WCIqFIG77vD+LrmDXUPH8AiE
IPrZsPnCxTWWW3FRCAE5W1BSuvDFWdNsSZmSSC1gc4XzblTjaRdyVC0Mp3Gw3f1CAiZH53u50bjx
atuZhz3EAE1CXgK2UAUP1sg289RvXTBliyy7A91XObIFDbuSIG/ZS9UiZzoj+9yCWLAWO4xlI3BD
caDjvIgiAyrWgFP0O1Jfr1U68dUdmi23oAoCzQSVVkWzg9r9jGFuj4/ilHj6S/DbSqkHI43oEB4K
kQJXMHFUo4rZXw9Qoljlyqe9LtIAu0RFT4BHUsg39QMkfvbO9ALLLJ7cUgrsFobAcoJrJ7JiIiaY
iU1SybWpOFvkKblYujuuFyLYR92Qpk/znxaDVTRinaPTt3/58CufDVbh72Czz1fvWl/WcEFFXCYR
S9YzrZZZ6DnZOdHGsKUfg0m3LFqAtMX89p6fHkC/32PMJ0Tjj87J2I2QiCk1+v4gDdtw6D8b9als
g7KqLZ60LnU3pZTJSQn7xUM/HLmy96AxLt+phn2qVtILRwldZhQJvR8V9ZXgzZKTrinq3HrobOeT
IpdzTL4tIeleXBwU7kUMoyJMH3ERYc8+WolfworMH9OBvyAnSJ+1L4llmQmpd8e6FxE6+U/fBXSb
0Wg/16HUmawcY7D8LYs/hmmokbyJZ+IR37aZbqZWKHU1D+YuI2SCoQetqvf9WNhp8kLEtVZtgap8
mjiqzfQ4l3LG8xWxkDbh2s5gRJmNWiI2682jPncVThw8Xkoo6ddML2ZmqEoin0FRCISROehqbk0u
ABwirvrusw4sn3mwoqY+ynwPyEvZCE5N4uK5exVxxkehk48nU6vWm5Mokf09G4rRRoYMns37Qqdc
dkuwROAk2Z0ajh4EqxX1nu9P28yoAvhV0fjnQxusf+TolI1tUYtpZHZsQV/PkTwLwk4jCCEdw3Bo
glRxtcnAEnqDl3kLo0sGiR0L8Xur3zNNTmlNrH/Gcqn0q3F3IoAPm2ywakijVazSBT7Lj3n0C2Y7
t1cw6xFi47x+Kd6h+J2I5aylbF9ODlJeDCMOtMzkyYtQQa0L7+UbmXWnlPyEg2P+DHlzk4cB9L9b
3SERU1vW7SwQChxtDeJ2Eqq7DDqT0+l1iL2+ZTbFsk3goKRpGsxThawUSceG1ouAueZCmgFS0lYT
C/jLw7fJoiWsYcny3jAwpOmWmGZhKsl5CjKCx6itMjuku4H01M77zOwKkEK3IOeTcblRQXDq4f5f
ROxxsbW8NgBBS8Own3Nrz4JlnsFZynJQ8mOkAquiAHLAp7n9R0HHCWMn/dCg3lIDTmAekyHzSSCy
7BK2DzN/OdbEOzBPOoap3B3pxDw+gVx2O1XL7BxbEUDT57zNV7k+Q1KgJYCOzIlOQG5cokwgT1Sd
zY+F/kRRKfqpM9c73HYigbGaIK4rKQvfkelhsr9+RH5stvBlAp8ur4Dx6u/cgN7TIxK5d6SmMppI
p9j8n/KgsA47s1KB46YhudnsdJaRqpJE4nVuabjWy+HmHxmtZCg7MLtRSgyo2PKo5HxX64A5hzRD
TQpHcQaWizrEFzegQKFLJ2D69T1ENCoZghZLpHc3OtZ4IWOhRoeCJJ9UjAEXC4t6o4JRp5nqydYY
eNqs1mmML1Nk7IOFdNqco+hccyXp4zZxr2bxpYzDpF0tQn88/LMZnSVEZQH+0eSyHx7qwGUu4PuT
fjw19hUaTcTcQAA8aDPvdHNFt3uw82IdmynwvRbc4pY+PxI2B3lLkhOkUYfmh0HrxRgitd0wqqEt
wKo8+CUiHshcmzA8RJDQXKilCY1HptdJq3CeE3WOe6uZuAzt4PXLQFwoVDXPp5J+ranRzCQ+QWLT
VV1AatZo2fC6CkEKFCsyOHCyCdtYtbZS8+tijATC53SmoE1+7kEdrMIn2S6laUO4Ju6b2yMTSXHW
RwSlNZcjrEy/iFX6Ymb5bhN/lpEkhxBGiLK194yEyF3297vNmGt26F18h/3eWCQVUnX673HHke0w
rmvhrl9N1FD6nw+uepqR8/UP7U7VZhYRI9JBFsnw/HA63AkpTzxBEdhqcoGAOGvP8u2lxF2k2Ehf
rVYKVWaW8EhmjZMUxjtRMywuwn2FLotd83lbQabcIgcAfXe6mRigahX3lGvFWuyrkPh78xhnyR6F
PzqH+kl85R6DwYb4TXxYlojTwox4cejAMxjkJXfhdSci+KMrpCBDFFBk91ejY9G3vuZEtkt7GWJe
zkOzEd/jxi76H+hQKOzxKcLbjuvrN9vv4PxAyErrK6r8oLTZ5TKo9VE3v5qWH6f/jLvLAUMRoMoU
es7L7vtOX1aLF2J2h/4o48J/L81EdNZo7LvD0Cd1bx0rJY36olec/0np7PuyiPGXPLsY7KI3cg1D
98+/bFea37Faxg4Kj9BjdXtEYXv9ZN9b4aTOm0mn+g4WXoV04Bfo0/oe+Lx2+9S0P1rvzbhnRgU0
WpLmclr4+uheHjtyeND8WvXjqh8kq2Df/N3UOXh9Lqudjh4l2k4yuRgQubbm6N+mtTPtzxO8rQRe
7ApexMKBx0weXqfp0VPVpDMs8FPqXwXYI7YSIMN6aWk5pE2WNXiNHbRB4VRyAEGqzQ7aAnyHtjS6
pX/OzAG5qBAC/OhCRYpplsw3d6yQ7M/36+M1XbOJw0xLU/Mq3XUKaydsCdptD0RWERFaZv+T9ifc
wOt2h1B9rhVAY1lhdF+dKJJ3bH/Wd49VdkL1XSp+PfTsAX7bP7P+dXoJMl847cVL3wtuk//0wujB
dA5bkrSYtLwLQZ/y9MApVfP+0nr/iQAlogaRSEve1qBMNFdRZsxLitqzkx1HWRtlm4mU9cnKYd/B
IxSY8fwYt/jPFuMj3d6rT4wx79UBXAl0WyxY2oHLBlLltO8dssEz1e/qLmtYHNCuRtEqFDO4xdUP
hZ8sVWjD3c6J/R1hevFR+kR0pl7AaomWJWfcdTb8CRo/7apNCFwXS0Um79+VNcNuO5/b/7Zon03l
Xa/FhO+9ilVG4RC/XoBy0eZDxrFwOwllz5jMa3VuqtfVjegtD0p7mgUl05t5vN+zDQumbfqnI0oQ
3a+wZjgPKj8E99AT7h6BpLEbVWw+s7kDSrA7hfHMhltS0+R1hPglZELtmKJbr4vLn2LmAKQWdtZd
P7LxG6WtPumvqIoXzNwxn7qabaGlpF8gDhddwwDayCtw/sUTU7FoZlUiQhDzn9di2I3GRoV9Z/Yu
F/La75prG9PqJgl/+ydSQm5o1dz0M2ljoRs8gVsLm1OVRuo+UoUcE6oPUCuP1680cXOcG10AQz2s
8lxqAKHsQDKQcV41uYc3EmF9O1ambRHa/Bi3oB4kAJYrtXnL/ZzoCqOn2OObWnndViHFCVhhUYi4
s/21XredX+8mtaFIbEQr5uMe6qjSeasWtNzkxqW+kBGChKO6WviNxyA5VWB8v4pjTs68P6ZZw98u
ixlkEU6ZtoJNZ6F0H9SWB6f4lEvw2X3hUFHN2OSPyWn3Mmp7MFEpvm6PkHbq1+ogkhDnnelFGW+q
ZYf0r5uanCC2mkKj8f2YDg9xHt8ovQLnwc/XnYQdaScJoJtyYZwFq2gwHR7JFyuSiq70yCdykIIZ
GUS2aFHgdA6Omuw+UdOnudXdJPLipwjRRlkLXscRcumklZ7FzylS7u49ZPbiE4C8Gg5uBWGvloQK
CWjnX0y9DsRMSK4fw6NGabMzizIWzzgY1SsCEGY5NflWHcgo5RsYKcVYNZXkNMzVjFxtbfToTmtQ
xsOLvCn+z+h6yzLyfWvWRAe2NU2WzMUxWOreJNRbSdtPhLA+853VJPfVQEZb4Q8gQ8VSGtFrxg4c
Lz4MYBOSx60FDpVZ1RyJlzSSq7GnVW71h2Er3KIbPbIuF0yrpSgxNN22F7lfSIY1PcXVGIXOO+o7
YgdWaBxPrGoHVFyXEwU6iZ1o+hGSCY23nt5kq62VlSTUZCNjGZ1VCqSrbYU43i1t7uBGUYGdAJ5n
x3Mcm8z9X5TxwUF6rYbLKVlbUbgG4jYOzznGl516UakbDfk5YpwmuQxp5S1f1NbCuqKIz66GpfGu
8X0YOx1LfSGpgAt10MNzHiH/6o/vgXf0HmzUJeghStpUNem3+2Mz/hdbdYHVALM4OQVqnvP8uNtc
AMaNzwxNilu7NfwED65wj0z8XZJp8SSDLurrZTV5tSs3b3UJXlaF5qswjIPI8WAfQejcJqNG2eYc
Suv6JBzsdupUnyxkMS02NBh6J0ka5mRgcUvzYV4r0EmXpGMuhGeZg095wIJj+ZpLEPui81AnO5oL
xzQgzJfx0/d9lCGecPJB46fwkxi9vLA+JYhQXgGTTqJYJb+hqbxMgpQSDnXW4G/P5BooZ6vOnyEx
tMN8uwVyHUDt7Z2lSx070ICvviB56IT+mOzIZ1D3kQ2hxB59RsmjxlzQOGhcFSBSXuNlWK+ZakYQ
Rw8e+SnNp0QtOQhSNJDXaEjSDX9aWBO9o8ft4em2JzHbF+IOMesGdkILJqxHZfY6p2JsikVJYW7k
qnJgeUydvKp4KM7RFns7peyS2lxrdA4FX4JEgQYHwtQneASIn4xGT8bXLB4FWjJA/o3dBqWTPgmd
i89kQAp0iMoqqKDr6qBB2gNtk3Jqjfooe7ItvDZ/jhUcz5wm1Qd4irgwVsjFQ/XrPtGr0WZWBYBA
GEYB4aDZmBQgtlvXyCAJ695aMKK/J/BkOKT3OoTFfYclzXxSDthq05XVX3BRDErtu0Z+rnDERtXI
ksZAjTjhmN1rkpvpqGoffhk6IOfDKLn8YlUFlYHFUaxBLwTU6YVa6rr8Mm9awVDpUzahe14rgk3B
m4SaNAYivNFyEOdT6Y+BI+2js/u9mp1D8QeZitsoFjM4XL0WGmkkotah2gSkq+b7eddcwcIK7gIE
rPoXOCiZ8B9+ZEgkSeAv+OTXwtP4ol5aFfzcs6Jxqr3xyQZO/YORCrTZ+fsIZIvuBXAPDYG0d/Xs
iPLzdsGw00iGfOK8tAVWRaVVHJPkB1vhshM9r0+Chb6XgSbnkVsnKQcr6InmsOsrYe6CTEvcBvB9
oOz6bK5e879IjIXpRjxlDBC7BUbYbBHy3qogxAvzOyBDa/XApXqxZFMKIVQVUXVQ05Bjy5/kChcE
vc0kQOS6bOSpwZupGo9zgm+audR/gdcD8Qqob1fwaYLuUx5Rv9CfLw/ahybL9h88VB4Bl9GA50lG
OuGDJyylFSHxS0ELFHychExucEIYsNuuhVPISZdl0UeDFnVOIMIcC9LYw5VsITBEApBhSe4HA5ND
xShVrFn34MPr27TF38s9i7xqNu7zS8Z9Ckc8PRFIwUVgxtDBzwSulcuLHIgFeJNxR07mLbQDABNR
iIUUq8H6/4SkpzYeNnI5fkCL8RQmmvEIVn2aJqbadxZQfYUI/rIcDIs3X0UI9ke5tML1Aij/gyGw
7Qxu/UVPBa5LybDx+R5b5dkVNkRCrvg7ELMFjv4gQUVsIaGVJ3pCvLRxJpR67gKSHdL6HgCkg5SL
JMmfyMmO81rRSARnN3FCJ0IYMuDnyCcVedNVLHRgGMJ+QKYWEs20/ZMceT8uMlmCQrCCwTVySxxs
GHjd7xVpBOKPYxlICoAmYpys3pbByXQ1JEwb3PD2JbA7arjgBJ8XaMW7zgw4l0XbDMD5VVS7/iwA
36MCSVVFZbwTY5T1Oh/Ft73MRM/0sq5inYdJngCMqqHY2za2HFI73yAl5pHb70k43mGz69tiOLx0
VsVTer0oklBTwy04fzYKMCZk/0nY9Myk39TxRkzRP/AJCqazqJvB52TazMaQ5rdRzkgq6y9yG365
38p1OyF33LKNu1WEpspTZWofJKgb+ei7Io1OsGMuA4Sl07Vc14RQj+hewPDwNddDIltTmnSA3JeN
L3k1QkPhRmlR0uJNbQ8eGH+Kh7o8pcXE71I3egcdyeBfNOQwXcCSrupH/i6BZ/VtUvcMQB3aJwjp
PZCdRSPOAkbTYgDzVGWV256V+6IlMNRB8d3e/PLJaSlM2m/oDrVxG70onCJ+P8yrNGOi2Ea7BFGK
GdAToCgPYFhAkQ4lwmqvATJ8IMBWX0vUTXzmaO9J+SjyAv4GW5hwYwXD5u+v/jrVy/LXWWBvsbp3
E4MrWV5C7ZPYd7zp4GsAQU42DC3qnQNrycrgtNi/+k1g9cZUkhPbE1eIHFCfOWTIQXvt05qKnnUi
HtYkIGh8MWAudHu1oalvafi4gn6xf6JLDnioXsAugf/daholCb8Ro3IeH+BPcqbbbzxqDTiePPLm
AiBmwBH8LC0rZKfwMYNWrhzVQMf8yoUKBvPYYsbirpZLpfJWGbjrg/IewdPH0+lBVpWdBsZPq0cK
yxLVV/y8uZkEwMgtrer/VZg3nT3HriJax5vbAw23ASbKBffCOOrXJ1n9QgIzWhXz1g5MOWYWuyha
Jlhl2p4WFn/VzTr41ncy4U3qtuLXh5yC5z4ypqngzZULwcnQY62rIGervQDw0dz+sJJOa1NQgp//
q/4InGvnWPMHJOsCHmHHZgvprKXhEi1WN39mnDY/jzpXXjsjbiD33wyiK+VuompQx5swJXuyPJFJ
zi1YE8Li1af1L5yCYAwoiW8RC52g8eGSVS71vGzz8gFVJhB2/vVV96kyRk8WYqZDQODwDQm0O13w
DXACxlZeq7hSexg0VLXnr4aTWj+8RTnEhp7ZTK0XrOUdfgmG3JSbx0V1oAkfDREL6LOCEgggrzYu
jmhutsuxlLduUwJmmpW0I3pHI2WLc0voIusOxwftxY5hp5OKKtiTTNoktTAP0S7sJBhkFd+DoTUy
MeK8CO+Wr6CRc1k9HtNO3OMwZIfeg7H0fT1yIaQuGh+LDyFqwDRK7gc7N7z6tEVOGGxZvsneVRXB
2ogrvTtelyOKKc4pUguB9YWFGY4oKe9nnAnGhS0RczoSY7H0lbPmPkXQsTGjAZKnQn8mK8RgwcY8
67e0ri1ZlxTkB1OEUkJlUtFwnUHCB1aaRC2TAeGw9uyKzzd5g4oYqxJg8TtPZgrxdnkmTFXUziB+
GBgcydvdtzPwYxYwwRN/En6Sw3/HirLKB/qnGgBqZ5uk50tcZq6LJNjODQU7SdPZLwJU6gX2gpak
UKAr0xi4Dr4JWgO3bBSptNSLdCXdIAkdwpnVclEU+6QesPseJF6jaq9at7HIZa9Kacw79scXSm5Z
B4+2bnFe/H27xYodmtQ0RVio2j3MVfD2Ss4TwPMiKn4/5yt4za0czgJzUW9SBY1rmG27XNjKjc9g
0QNkeVstEY0ZIrLMtwe4wgfGMOTxzbXcvtGkcgE8FZzWtrt1GCSU6UAF9Iuy2SiFI3e5ila4z+T0
WXokRl9b85YkEgIsIG1jZ1r8VsYBnJaSMxOZ3lQ1CFS2LDUJcZyuoyvM/E4v+jFxfhCJsI+TFEEr
SLFbXsI0cU/8AiYR2J8Babc7xSo8QAkGJeGYWNu+7gmnSD0SWHrlbwNvjQIRJ4DYNw5X/pvIC6ci
LP2ghZQ+kNjaLuIrYAWbgUHsBmEbaSoDM3CFI5sbMoAxXZHhVy7LM5I6IXkQi6S+1X3Pm+WiGDkz
zHZRYSdZYkOvEa5F4ZeSpW1/GW3ANfP1AMc7/I4Wikt+kMVJiISCCBWmnIR3n5836nVqGgZ3dCNp
qrwo0iXyQNomDRRvtVD+SUx3M3xdiCunP96O2cLDbsqkElbpzhkd7QwB5iEg/Dlv6KO/+8Sx2h6U
LS7406/g2B5uo/zhqKAGK92lWM6N9tbtcKynWIVYaPyEGagAOzSgpFQ2GdhNtCnzIG/0rnK+F6RE
CVWoQr9xhfBiJyVsBa1NwgXK2jK9AWgFJTvXrDEYWDFCIHCqDhL52lfKRFD1IE4j8eZegExKYqbQ
4rdo2zwvxQy7N8QrjwBgs386IG7vEpS2FfXDeZvFTP6Ly9X2Q9PrgbDSo10iLo6VkEuApr8Ic7FP
9Snzis9wtXgzuVizTgh7HzBietEMa7zgWMH2DURHQJ5y8EkOyTV3FU0ytVMzOgFeK0HABG4meanm
/ergfZxBZfPeoBTkxXkrxdSgShNbYhaifCqGghWO/zY9pBCYSYuJH70AYKM7oioU3gOTtplJigIa
pRPbQENre/iQkp0C6MgY2se3p5ISej2HTNsj/AbK8YeqoAbiWJENdr1CEeAkW/B1sHxVHQJ9NntE
SZn8RFQUXXez5w3W1h5XKd5SqVb9PbbQHVanHZDKYqghAwVNVUvRwEmh3GFD22EUzbF0C5QIrAvd
H8FsjDO+58c2LbYKhgMSiqX5LlfRE7QJEzDnXvyXUfq9x03pH7pCtYV6e3m3Nysk0tQE4dyJoinx
LttS8tc0U68xo011dASBgjsJuWt92Rhbc/b9UfZfpPYzQvuGMDIEzYtZxHu50tp5tnCRHKl99Q2j
L+KRZzk8ZBzkS6YWWSSfJ6FCFc4IqTTWS+fGpjpQpz0qBF8Ib3aJajH94vWmdTaDaMiT2ChGSIzW
9mbSu/zFrdTzcIId2eIMjjHsckQp8HIMU+DeLJ5/5PGVL2bMPoJdOhm471JKd5Z5E8zFCf3ntFHt
NrUc7A4GIJU5/JdLEnPGTfwcQyFKszptxp6IOZJGVXkhG8qCn4gpjH1436v6SeUivQiRgB3GwSAF
AK3PX71fMGtsAbfM4x6ffMm250hlDTK9zj10WCorXO8+/Pa46izcsGyEr7hrwzquKdCFGLt4gF1j
VaA3SzDAtJRi7ppP4Bfgn3gb7zjuMWzPq7c5GRlP2Y+LbDeWLR4U4RRBrdug4gmo2cOggFKe/rgY
MLCookUyGIwyaCowDbFS/TGHIQxuQT93T9OO/eRYzNjSltDLef3hunLuq3jyL6lOE9/HrGZeVyVm
evhPodqqyVw4rsQ43bFZ7KVR5lhPNnAVYM+I5Ix5YwxJkYKYjbONZZMFjmHMSxWuhKXE65fqiGGn
E+sKzdRu8MU919GvZSIBpz+2/uTT8AyOWDxeRgUKcafMI9DIP4IuzGgSvUjmFPDwVgbZ5CAIdZpY
11rT8L7bCOZOANZ/kQhmaaw8nqzmXWPnuHzQzT4nIBeirLvLd5Q8Nb1r4cwnsQDo9WsCzABLbQcY
fDCaVnOY43r3PXFr1bUJKSI9K8/qSh0J761/ZJfh+3N8kCefP0o6tKlRkdyA3Dg6oy377fvcmsV0
knMK41pTt5U/nr6PnAeQUqTqpDVhq5fviBghCKl8yZDQfcs6RTyvrrQgbl/415TkxA6DSndLVIpr
1OuV7MutPlC3GSCf5JIci8gSv+iYnoF+tSDIcS++eamzj8L0jnVT4OJ1fvhnMPJ1TRbkHTbYkGaj
Od4jPbCNsHo/0FKJvi0RoX/628qMLMPh6w3Z/c5gwFsW2sE90VJHcG3Cko67FzECYfoRNHKrJIZA
ouoeMcoE/rYbFZaYWC7BlYBywaMDVDYyKcw72rAuyKKzh0QsyvGNw+2zNSgpNkJwJexfzxYcsYV4
AxPgCG22DOy7srATz9Z0ifTRkMdITMcX7GjOumoU0JiK5MuuIH8caMNaWVaOyDMs8mbm4U5/DpUt
WlBdQMPWVsSTzMbKR3FGNHFeSWNOjQNQkU1Nb04Q2uw31FfeA85ODpMi9ayGgh97z/5lanJY5Hce
GVEEZZX3xW27jk1Kn5CBCj0eggDaQ2Q4Oqeam9FKTVgV7nUnt/LmyQqfGYZvbLWgdvi0V/r7FMz1
xuxSOGiuolpwj204fkJSog+nzvbXq1tLzwzUxhJEXI5VhPr7zRgMp8wTwYZu8JPsTShwebBpeU94
LXjx08v1Qqqjtbz4LhRFcZtJAzTUe1XoqWSeuDpqnJpvrQ9+tZj5Jy/y2fv1+/6WIcP73aDFbzBY
JjcSdk0GBIRM4eBMmzzmv8N0CcSxoAvPBboL3DVoPKflJTX6UlowYpt254T41XfF1tX++0s3tnE1
s/CVWjxSvkpsG4mVZetpLF6IQFQrCEOF7bO4sodHIgzQPPI97Ha4gRrv3rVY3azF+4JssyFKV51S
t5jDSbovMG+FHJRwWGRPC67O5eZOJezBps+XBd7OU4SFyQwC4ehzQ6zUolQTs661GB1261/NPlUI
cn25m9teeTn/GooqX/7M9k6d7gjyytZVkt+6IUmxLLKwLqFEGhvtuJ50wBn2xXa67NYkTkUSuQhU
N24WE49hiH2lQwtrqjZ0Mg5fQPczpSqnRW/Qys1m6/HnFRrG7veN+eTeeGr+FJTwGYgYlD3AutFO
g2dl6RhIkcSXsSh4kyEucJg8D+gCpVpfBY4NTM2Wr5TTz9eq5k19jLfoJCtK0305aO6KDU8F4Lnw
HQCM+FJDsDsyYw2qP7StpWjIDU4176pvRYhUIuFQRNwwfUPvUrJk0dUrOHafnniXextEFw7B/Zq6
HBTBSVKLiZcv2JI2qyuu9R9jh0NKxNIvwxWDrEbbyUsU8cRr8PFfZxePIWQkr7gloT2rjE8Ygv+M
T4iOOSGsEkVQvEjO4Krex51Kz69hJ1Vgo4GAx4xn0CciWBmEtj1U3A8RrIIGxIF8ypmGgiRFpqZ9
LS6h/cSv+gfvPVpH8/dIEKYmGZTFgS/E8d4u8PkgNILoAaIJoiXBjTOVL8PEkdMruqr2vOwqAD/3
B3ItE0AaiGmJmole2gm4y58TzXs9JGKLO4Yft+XsgqwznPbRmb67DpU4cWY/GWYa1TDTedrZZxxu
y++DeaO5ZBkVSnpT5/AjOnRJnGCINQu11LdjgtRlr+qAHbaSGWd/4DdpSWv6LsnvMpbkbPoYOE8o
qFt3kW3fhCLhlLTrwZvej4EyzIkuWMZKh5M23cHO7hl0Ufwv692MUQp91HA9ALkHNfRGarhaDb6G
Pkuh9GOuV3vo7pTSVNZ0w4xwXRpJSkP5Uqg2OCIpB5422Pr8xEux5GzVZ9Wi5Q9X9bmVPHd3cdeI
pRhSrHHSqpz2xi+9i2dTHqIYTmu7jivw9DCloAM60h4y4m+dT+GvYyr4H6eDb+JQivngR12kItNb
7YAuekmoJlNpLtVOuDFQWcFNwaGlXXPhlgKPOagMwwIPKoI4HVF2l6fMdhyGa4T+v6fDnOzTVcPN
I1Bq3B46ETUAV1bqjn6+5v4FTiKN1ppU2dEzeWfKphvG3r5zQou8mHCKyDHMNGRlnLzIvQkNkXS0
0vuLn+joa4jyAxelDxiCude3PRMZG3W2QsBylXcF6gKYT2pS/QEh9UsuSKvL+4bOfeOgL27PaaZ/
hWT1+rV8s1DgvRfuSov7pY+rjlQaotbecz5AyyzhBRkoa57Z434QZ14X6dr5Z3C65oGs5dVW5TUl
qnYCpwWly3E2OZZkQ6of0SSawS1nlbrpjnD64T1btktzh3cQ48qtcJOeD/FkSmPTz9Je/qV9zz49
TpCnodbmQThb0tIs91uXlXjjWpgLPeu6YPfH8GfIE5MHh8vLF5n/gImZcNoOeW92x9kEscUpCH4U
PnNa1OFiYZnUfrU9tqCC9Og7RvgH1T5akpTKObKki22WM4M9EowYbkk99XfdEpPckfcrWjkM8Wb6
sLaL72Fj4V9tMTwJEFNzc5q+RCjcva3nWhb//2sWcNMISOkjVEwRrZFRzIkDoco6JpBltwyTLse+
7YE48GrLaWc1lBXgrCjRVsTlbeyzTlYVY1XySfvFED77ng7s5QDDPyd6/4nXiqT0llzSX9FrLYnJ
OQHiUQ/KJXwQP+fBOQ/D93Um2Uh98Ca2v/eLWjLp/nA82KGOtDU3YqvfaQJS9pU7PH2Eqyk4Kdd4
d5I6SdNsTFx1xcxG64wOelHw7Agk6sllJnSgUzi8zOVgyK+VbSju3EGxxVUEBC+h/TSQN49xFRls
+DgrJ3OfgSPPI08dFjBmbJTb33z324y0gp5575hBQWoIu92ZM8CXjpK24dHMyq6BT0zWCBJPZAlw
sYnJ9qO6BIOzNmDSgBHqPgtalj3tAaOxdLy6BwTKs6qLkpGm3DcRsMCh2UiCRIlNHi837j12X4o3
hOokTE2Yaggi5YJoOxE470Bdr1F0t/0RX6hx/1j9+gwp1vnULOAcRkCvN9r5m+aBqHFj3nHElMnd
hg3wcyhwY17S/K/nNC1yc9ehUVFJyY5J0ZOWAF4Vx8FTO70H95OSHpT/AKHYqws9tfu/SCEO9wpt
VKAlX6llGbMcfXCcSR6E1voC7FajzrsBP1kuXJAS2qDP/VUL/xXGD/Haiz/qMzy1yhoTqu0JvUww
rACBkTJeuEq1w+3uJMtfFzqbG04YC3BtOq58g0+XfXOyK8+P8tPD6bJL+NN/mPYHuhV8fa9wzHO0
oPeEALvVv3/1EwLxpda7gaUX82RIXEsCokdBbd9dFYXgkreZrbnO04PwzJNoaxj2HVeK6CeDPsQa
xACtD+71/CM3zrhlkURS56fEHRmp7qH6jewoV51TAl0xru+sKL+KwuwO1TZ48dnsOv+AwpDVaqct
034mfIil4jknjLtuxHeP5zLl80VP3syvF/Dury/8JZ+mlzuXbhHwK7VBBV5xIo0sLcBVI53dsYjP
Vj/rOBwDkwzbmbY+ncbtuWVFnMcsGWwsE085mUcYdgFtFO2NyZUWfcTwZmdApQnLvgKjhHvDKtvf
/3iR/IgDbGEDD/8Jgv5y0Oc72BN4p6bY9EtfYNygP+zpcLDa+F2TsErthCjhwR+yk32DkFc9OzYA
XeGEMzLZ+7y3Flo70ddSLyBFyJQQ+mK/pfpIVQoKf8YIeTJYECv9kKt/vj6Ig4d49RUkbuN6kifW
20iYwetcSDSaI/vWmV5KNN4uOrH0XgShGq9tcfhkPU52UG9ppLqq8lsWWq0QImK8MtxgQQQUpw2K
5oRpoE6jgTN80hUAqJs+ZioqsgcUWEBi+LBnEGUyCZefOa+Zb4fyT+C1s+wuk7Cl5qNmtYQ6qc04
xBTfz8aZijgoydaAHLrICRMEnp5MgIhRN+ZrV7BJjKpUuMxguhZ9ztoJquejiktFLZiOvv/lDa60
+UftVbvhjKla2W6Dnv1utVBcTArkBj+SPNGE6PRy+9aBD5kDE7en6BDVDTlkFn+5TBlQ28UrObEv
xdaIylns+T3bVvWkuSpD77uBk+kuyOGcf0vgFJ66q+85rA+wa1nxvtBveSAl2LYO0ohGRzWmp/XC
YcIp+2NrEhBta86ZiYomBYiLDmiRx/wjFjl7loQxrHtfY2TWfmvxD+NCuwOI6XdZgXJoHTYJ3sZT
3G5mZhlE9M5OR3n24H06ode/xM4XScYP8ojzFnanvZtxV25c9lu4VgojWLKh978QVm/RB/LD0yCW
VZG1WzvTXgOA0VVFfRVrEl421mJRXzhiREaKS1LGjKxVhu6cIKClA3lYpjK8nhgZFCR7JTfKRfP/
EK2BLn8STGdoRYWlaSpB1GyhL2k02zrv/YtaB9oHNyzKE+0obln3+1xvscEuHe9pxm3RFD/kYpXX
6MAJ762oovMk5jcjUwYy6SKIBpR2kPQD0ep0lsYWVudoeSRaNjdeB/XcoA+v5oyKFhTEKcdhC+6C
RCG57ccTa0ojQ2bmQA0CZe4NslbX+kkVVGYY7w6plSnqQMKbtZTR0J6jg3e7esEs1Jendkcw3DhZ
spkGq3MplK0iu3rmNr2EglAgz9hm8tG28OmccfdkPXDAoekwetD/eul1AzogreSKjKthm2M1Ig5h
MXXROZ+JrEoh3KGrNwiGo7rYxG/RvEpSxZ69x3bYQqvAD9h56s2/JjGrBn9SWfJvDT1ydEj1+B/E
129K0CuGOf2GRV22ro7QNo2biOJWawAeNqYm82oCDnufcrtvekIconvIBS7Tum4MFe6wflmEwDzu
Zv3wEl9D0swrJIp6rNMmqi68up5qk3lMzyRFDPqLP/WQNyKamjuzdJrHzpGoQA9DPrYnAZFtwH4n
KU9Ngidivf56s9Bd17RvuljG1CK1CDMmW8n5THHUHfbdicAO1OQKKPTmQFggb1fVywleZydLuIZa
xp+Y+yTV/du36wKHTkpaHHLJsd7yt52Q0p8Y2GifwV9W5Wzr+Q/nxOVmnolX0wzjEO+Fqk21rspW
3GupO5bRSZBJxTcUjmixKPl+lviMoeyWpkUr4kC/DVkIOKStadc6b3uPKckMFkslmSMIvUOXBpjG
5MY9mCUM/+FAb0Zzcw3SA2zupjN/srkq0sSOS2hNoUDqc4VxusHKGBOozO4O/leIXwHRdZ1kQ2Y0
cM6w59p/qHBA6RxOJ8YLYg5HtD5h+j0EC4es9R1C5E5X0cS06F4+BjNeG5J6hrvjwPO3JcXMfk8B
6LchIBAqiHyFishxy0xnVZc8J8C7eWayDg2l/scpQVRzaq2iBTenGLupwIh7X4eS55hkAf8J97zx
YRkSU5KSSbBaxsqa6aGKFUNbvWz0gWWBO6qM/ZzwF2ClQly06MvAyo1CilGl370QtnBR76yfXS4b
ich/CErYH0dfPXMnybNOCMTR2uQkU8mCvII027e63epQavNJNO4TC12vZmo0Q9fMAVtekJS6/4Ap
qNZzFcXJdgCkvPrT4+J1VKakiGTRp/PN1IBfnejZGKtTDQXpQuKii6HuJOADd8DBPELhEVKhr35d
jjOY0ALeFOqkBBajsuxDESnsJABG+68ZZBQ3mx3Xj53fxJswKCZN48wRuPwFlXrpbD8J02MQbtlW
ZR30kaFactqxqWzMbQ0eE5S0yQo5soRcDKbnOOX/QeE41Pb0k+h7cAxileoXSnj6omwjfARwvYrZ
a/OzZ0QBIxTcGOU3QTD3W7MhO0mqAyXRKUIxg7YoLpV8rcdXRNmahuR7yWGYSZqr2QAqgCJc/3Xx
9i95SyZ0PZViWEcgkAzAFN/mI2FwJexmJh7QngMI+9nzREwjF5SbIkhj85gHQbk7vibCdeupbiEq
RrX8JTDbwgukEG/CJxVYfGuuKVb7bl9SFudlx09MnOtB81zx0ndzGls0Cyu8CNXvDa6kX4sjcnCO
L5mEOxaKbZ+8PeolIuZ2CDROr5friL6D38q7MfbLG52D4eo8/Setb6PngDT50sBxkPeazuYV5Tdh
m95XElL2YuEBFKufugIlxgsuqpcAj1LfrOtnj8x4g7FjB3Gcejd0QhT5ns7Vz1gdkeeuqZaQwXzw
u7icV4s3vQxSLOcjttOusdtZq7YbGeZqbSNTNu1OyPq4kuBmIhOZjGm5Wjhn2pW0ogpWF9FqZGkY
KRn1qaIXY+6Wmd4QQLu7i0bWyXp4m0cmB3X21dYMNRAcK1rbd4b3wOkaSXsigXIIoiC7z2bUimYe
4v52PCedOm7Mg9uuTWaRBzhSqYyynuHk8ZlhETFtUe8aORKOoXiP9v6VuZWjMZyUODvZY6Whf7uR
C6UkcHaWwlHKIBUIA952+XryoU4u3D7i6o21rsXhjDHSW1wZapqHKrxWMuFcF4x0ic3BiJvMMBLN
Bczl44NUiLSd2mf6zulnmgZ+xlYwXKayZZYkQHS6B07pSXEdq56xPrTa6GH+Zo4OFJH+WJ5jrOxi
HDZzTZQ4bfaMaIdQshm0trwbOEBperfWbi+U/ICjVHsFaNRaVZraEKF5jPFKvV2gw6WE++UUguoi
2GNSlnftj4VFHc2GsZKEuIbQCAMuUsZNGdU6wgjEDEQv8qUuLjve24XILaC4s2MWLzGUWbh3x04R
7W8kT+ZiVhIpfUQm+x0MHio2lFQS58YkB5y6/1mFAovpj1YG3P35IOqTjjtP1jLmYCKsiVxQ3slg
+E2y1XkaNeTT2dSIudvuqLbTtBkXpURLCf3yPu/YYzXFmDjrVUhGWsKmOy4mLbMYAdJLOxa18Xh7
hsBj1ZRPdrWR6bs6dJeBP6NwXPkUzQJQo+sVxO/CBJh5+I7kvzCsmf1I3ia8jyeqydxTjEOK8UNh
p8osEXEI0nYNXHCsCOoLhEV48192DSzxarmoP9tlzLjrgsg9g9n58GtkdWI5q0KiYzX8ApeMbO1z
iAAOubqmt0pBMxQI9a8BJUJ1PegxRMYP7QmXpuCTpjO+DYrt4bTW/vtz8mB1CLGqLIWv5K951vCv
z9LADvE/731YG2591qcZvU87keBfRSEiSO/2UsCPP7wx7xMRkLzKO0p2vRngaq0lbkZZpPBpAK15
jw6/+qvasqLf2jAGYmMkfoSXDsBoA3RP8CQLLeKIIxVwDRD6zm0X6QU1foNDYojq/wKJtfAp7IGC
tl06jDzi3sOZZiayEH6+Fo4l3tqWWZUV5wPNgarcWWA1lBz8ui2OjJN/YZR7d21DOcnhX8eFzf/x
MsL9SXsEvwZ4iXX55vFfrmUh5cbN4IxpNZndgGv8A5u5e9pxYvp48XDJsQdS2CJ2JuAbhqxNtoW2
AOcW7xURkdU3ycGoLLQcfcJHcflUiJd4/cLucZ/9qIuvHw+jxRRd5ihQ+0Ic0ECoKZvPcmiRyx5+
LwhZZi19LZ/LS4QgdlfOELmzI/KfdOLaHgAyaoTE+39i1GxZZbjATBwKI+J/em7UBYYharpzAndz
VwxGI1OJctlCJoszkNiphT1jQ8J7J+qY5vWQsmIfabnRP4EpeSmATWRqI18Pl6KuETzsmBYLYnns
aHYWWdD4/fdv6WTVXOEM5wGF+nWT/FEHh853z2WscYlgyu8VF618RKQlEhbmf7Eay4sn+2MeH+9S
xgPruOPFMvs0nuzAbFA64xi5U9dvFylMKqLDW5rh/ASWGBD3sCKH62K332aI/lqXCPUYXSPBl1Fb
+4fvkzlgbWvJJh9aJeVCWkkiOi3L7w3lPnJ7lv7YwviMEWEdw4KkkHHZwxnR4M8iyTp3gJbwJcnz
nAtDNkoyk/02i6qj0232eZz6Ui1g/OOTDcx6cI3eNoncB5FG1RoY6GAgx+s8RGW48wMOfQzHb/8x
18rJDIK2sTKjoL+RFRTD84VLhyoxaDZHYO2hYnD4CQrFX2SNXyoOw5rXUqt9aurIK0Uot1HMtj52
HO2QVvlMzrYA8UhWsaAfyUTIcoLq8PWJoer97zDelQMXhJBgPe60/wfPz5uHT4/PeZagEPShVq8U
KJYjvRdbYngUIPVw+s/o7TpdJlMIGaVsplUf0k/oYXNjakn5zXBQPMLkoD2mX1xY/lFfwEWB+HAG
+pvnPv6UbPIqxe23kVyoj/ry5loEeZt3HsPFoGpGYDDtT0bjyCcjn8X0KGl0k6zDXdiFu3LI3983
QXEScMOoFeBEsa8YloRofkMU737RZpXeyPR/DpW3LIhlpn28mEbtiGAbqntBfsRJNEDVZqyvTZ9U
9ESCQcdHkfAJgjthWbEKx7YhoLXakpZk/ze2F1mLpDqIlB1jg5AwRoL6poPNQjLZ6mnKk/CUYfME
e4amMOKoF97LC8TrF3ZAhVd4rL/K06p/kwJjOVIiJO7npCyUPJSHIelaxNB5Q0pm2EGhFZfNfSYS
pWF/toXEUyR0DcUeYSXPZ0PHKEukdc5cMFVUyQh3EM+1eNRRj4cWlAFTfHl5q/uqqMP70JwDEqCi
e0kQJuKgR+K5iG9u9vVVWsjTj1NMQmOQRIc2oKgu+9bK6lZ3jKgqZOp/q+fDT0gYciuZIR+PFEbT
AmXvhCby6gDlMc6X16Ql30SnWXSsY5g9rMSRGfNOox/I10nosXgoiKkhf1siDWtErSzUEwk5f5a1
V5O6b/1ghU6v+jTo3OAslDtTy2S6HsWpBk0bsHIMMR1qBjp0d/ou1uCYuozhUIKTKXBd5KBv3wup
OOIYyBS57i/hoZGQ8p45LT3TIBPep+DBX+wUFRcaWqNgqB5pOnPigoGW6AWh/2pDYk+qCQHq0TGp
0qnBVAZCYelBaM2EIxU+Vtdiu+VcckRce9k9mj/YO1HcRGmzZUVKjaC1o1d41Q/vJGruagNNyExE
zHdivxcW3Mf5mDpS8hk4zgCp0veU0llovjV73tKauwWJfHughZ8T2U9ZdwC6guiJxxUAP67Mr+pZ
hLpbXsS4ZnwPb4k6PMFbav/LkxdTkzG54pV2AeT34xDQMtrCIrVz4tFFhg5PbxJSN/Br4O50LK2o
WdHSGuOXLb6/7E1kpWdYP3426j8+8gqYG8iFA78zVb0cJCEkHH73nCa2HF7vCt45dkE3ZRAmVLNq
gU1JF9i9sbXfXMsGMC1pTZGjYIQ75utjjLeR8BJ3nqjq7U9+EHhheYalAqwCdT2Fr/ClpWCRWEd/
JA6wqdAsaNukw+B3tbK+DlK4NYw2UH69lgNPEQCQRG9yEGUctv6bnLW+D+Z89yXyRlD/cDHt6y2H
VXypXUGmoL53nV5YDBB7E7Gf+WKyDvd8PQue6IDto68OmkAek1vOxM2jYyeZ9N/geWwg52Z6bUOD
hXPjHwXEMlcXafmNW1v9r7FgEYjtuLj04F7hTkor6If3hxMgVgcJIq4e0sbxMkh3HGiZ0IIXyx/w
mwd6t7SHYCHrKQvDXIyYzv7GmALpfG9PyY4Qp2h3m/EUXl4qh7JzZMpBQfkMWmrwM2REW4kMBaRf
oOJHf07AAzmtuKpN4hOQgOxD1gt34MAnfR/i3pqWDYA+KtRkJT9mB3x38LUYljV+qTrtwTVfdcgE
O5p7hq1/XrIL6WDaerp34nZRvXMJcOGagsQLwMg/6dLorzlJihdecMhg8OgvAnQoLdlLMb1SAQ/T
kYm09OZH/llswt+v+hpIQ57mlTNotH1pSrGHu4vZNeavskO/GSzHnQIkTIqPNCFOWQiusAK1a4cH
wOiJ/INerpCDOkPWdgMgCndayD28VrLhwox7NWdisRLxh6jZW3cPa3JUQxA9Dp5lnEvw6TiGEAXu
r/uxQLX3OheKlhnT7nDj5RFQNyvLSc2WWmPQ079uDrBtvnyBLUHas/aToeeBPzezEcxXQStSDBKW
JMxZbA4GT0GEDMWFy7VrBM1KLYU2CzEqYX+VD1VfhAHDk9OeADbApG1zpg/2AnPk90xRbWDtvX7B
4kw23Z9/j+E0d4YsobnmVF521Kz4n0qMZdOYy1+2FlyBoTTEjG8qgxsx+qBFHh8cwcU08/e21Kd8
VerQvfNr0KV0JDBdaNQTDwGEC1rf1c9F6PU/cebNradXRO2PYSS+qSZTkRdGJCEcYl7mraetEIwT
K2zWmpBuUqajQbU/btj6rr7yOTnRLnmwStAldcjZ9pj/O6gHMVRdzSqDUjwK8UJiLSGgqp9U5scB
4Pb05Xl5b/UxkXsg7J2p06TCdNKk2YTrkzOouWMGSzbnpTaNFFRkf963adsPDs6r31ARMhpFty4y
aQWfmpez9QE+m7i9RmwrNg6kgHAcP+5L3v107nOONBmDn9iV3n/BzkXe0hXMNL9a3oAqrj2o4Wea
NIGMvgYUHJrQwS5UFZkhq8dtakI4DEPQSr/R0BmZD2Pduyy5LpgbO3jWfBvAPl82UFcyWeZpSvhx
sIKkpX7hFZAJWCFHcKjDNZxx3MKwMYukX5tD6pubD6xvniCVLdT/FgMaffXjJDr3C2XI0kmx5AGZ
nYpTrt0mlQGItFtA20nacEUSv/JjWB7t/l8o+GqBPjYwsYVyvNtd2IbQKgzygh8s53I9IQvURMAJ
ZVN1+mkqBJbYEmuga+WX4m86NAv2mySwBx0rhx+jkhueE5fK+LkKnpgCX0ZTRf2GzTEM1cXFC55i
NOz03Mik+gkhIXHQjoi9pjRhPfHbjk7e18mS5cLGeUQmLAshs+/wxrkN9Sny6h9d0zbkT90ryBph
V5Khh2JRve7C9zXBJswzHZqrPmh4qduMGtWwH3Pqr3hymEA6I9Y1kX8F2r2jPpIRhz10KJKCuTg5
FJFxJsqLOQaSNlUyUMacWVI/ZfxDX0dRe0okEg5/8joyhXnjxnq5CLjhje8n2wBC/8rn1rcb8vi1
teY60+YZClegJxqkcG67bObbPVVKn+Op/IGb+oUAE2wJ7iBEjzxY9ri/IhP6qojO4RAFvEaB0UGh
V/xRw7dbsV98gVabNSDZ5d2Au64f1bhi3FmL5Z54+LZA0Xf0ncdSXI9ymqOa55WABReYUMvm/Q8P
Rh5WmIVtxXNx6/DWaWud8y5/ugfin7EmwKN7QlJrLHaPWFuFTUGuGPx7Bj+W1ZGJEyMnESKJlYbM
myFmTu3r86/vrYuWHNdmjy8hBw8cYMH1uYDfYVfUNMNeZJWqMD4SVef+n583NesEsDujHFJXP32D
55b5yvIckV1VNJ6mTak7SfLMG05dq8BEXBuvLMhny4WKAJWUc7E/TAzlIDJOAZmB/bO8dgQ64JzU
ltZhlvN93XzziCgUhQhbm8XXnd/IuvBBpPHnwDe2YPZnOpjLP77CjeNm/H6rtzAp1WrBKJ9UO3jL
Zix22D3p0DezpLErsRveAjMW/dXTp1Hafc53+iwkuphnBrRP2nzLEqRW+991jIc1B/M2KTMyKXEy
GEL6P6HqnXVKwcTd9j0+PgzP11uM1VN6+53a5AIpjupvrjcBkqMnLbthrN1xuZ0cIvIuXSt+GFmI
FHHJrPFoUQ/LhVDgl0vb+5+zbOM424VpQUMi4CMhvf6hs80TQBqJKNPYyGywx+xvE8SSUOHD2E1j
rVczrAqwSo1Uu/DbJAGk9ZcadpZa5fpBqBtGNCgBmBrMW0PDKS+/rGMWzovuPXyZ31swJlnTJMsS
VD6ibD4BqPLOkKCsmeiZr+Ij4mVzj9jrAGPa0MZY1rvxUX3c2VUYtF/zGff5An/pPdQhjSQ8ayhs
dba6IcTSOcgAoEEYKdp189uSxG94uGSrcDtehDA/ROHWIoVPiL3q3jhB0Lf1E5t/uns7F2dpZe8o
nzKfjmem/1DTjGRClQ/Ffs26cqayJCanEsFDqVMsmYGu8CjU3saDaEyoEB4PXbYPSQ7tfcXiTOSb
gv93f0ugZeCQU1Q+KaCZGrbuiapuovv7WojGUrf+T/+A8pYXCJzeXfsLbp/ByZz4K0Vfh/Gmh3VR
5G1O8sm3BtQJeFSQjlV3hxDIQHNBnBAI6fHyWDH6KdM/iW8bSk0tCiq8dU8vSzTqKf1ZlNVVVN9g
kYIygxLul9JL8qpF0186YdPkVkElTNl4u4CWi5jnomJcEpAQCSj1gzqZJWmSfcWkBMiQNheZiC2f
PdeFT8ZKWnkXuww5HchW5XwUJCLZzIcEIi8fRgUw7w066VvrX4bZzkUHcniiF6o/KDuyxct/elE1
/W0W+JuZfpv4r3sm2u31bZ+jIUzYGfcCyvr5b+ThoW+gDQiEu2wRmujJnRZEGIqloQXJ0LbnMBPS
kYw/3+FNJv8Aq549Dvt9F4JUaASytkOW20RNEJeUyDA8LMWu6jYGOYBgUfJ4rpp6KeB8EJJB2sgn
DPTHrROTSoWD9wxUAgdsnY7qriTInduBRf+hFSMvwkIz7Mqc5ErfDdH2AWeZGYo8OpVpQYzmP3xX
q+qUGTOzInv7f9mXhsKVazZd2KjfwqCuV9SVz+OL93zrHbNrR5eapo/ozsaM4Old4sfe0HtxdL2w
LXMD3IoFUir6FQgOXxFZo/wMt8vppj3wkd0+LzlWRdhg0N7TBSa3tHO2C/8hPgKZa/lgLoU80eNU
+1+FNBc31B8PPKn8QVY3WnQdIS25o5rLoqwhMxAG3qDlKwKqqd0dDTgoPoC/4oqRnEevZa3LF/s2
mZ7eGCJz7Qg9OrIhL5fxRDp8ec/oVp1jUnsPdE1zHG4Foxq6RCPOGMWUe/SgY8jrg8m52csxt7rM
fn7JSOltMBO3HrCQfSbKVVvEXGICvXhwuBGfII7EhQRXPFnOfsH4OgZoi7cyakbGDzpV2Uwzt4CD
F90WgbAHE7TfWvWanwTWrdQNWwSTL0gZ8mEvuHWyQAWl/MGkEs5keql6zvYjhPs6Q2HUIkj6rP9g
qAZw3Bp+kGd1hmkP8XyHY+z/KNnXK/csV++KrVcGqGktWXIrlAQqpF2VJ7xXrLNy+iVvEKSP/pyy
B5/hq7vCTBxMXGdEEpyvlZ4k+UpkbXf4R9KFWaB8QXUeFpW4n/XleIwbQgSheZwamAVgwth/dx0x
TVFE1tASWl3VP7timnnR5aWadylC7jYTdF9As/CdrmXiePwEavFJ/b3o/ivsLFYjbSxL2eTaofD1
od7CQbT4D7pTD5mQrQfl0FVRj/54l9wWoh13GxR38K/omBmSwyRhDn2u3yXkzicmW47E58/Nwu4M
ObRmCyoN5xQ4zpLIqf7ayehcA4clEOCXWDVo1kZo0MBUf8evgTVJDbt4Rsc0RBf5+/UZsZsLkw0a
IyJr+4Ekc00Sejjeb35v8qoe+mAkrGRBdec3PUyqqBVonoBcPRMAXd2XINLQQGnJfsXaPZ6BNmRP
N+X3G4t01LWV2QgDFOi3g+zM4/jioIKoMC9ac3qGeq9FiFKPZh0aF2qU7ibvqYRqgfkzqF6ErWqn
kqlaJGWwJoCF6eZCZUoPqy1oJokfWWHyQdae2Eg3ej6miQufkgTE9r2GAr10SU4CBUzStS7/Ku9a
Zg31S+ZqVspcv8/plxxVTpU2IskmjGzQ64rjFQ6m0lCSxyovLncH0VbLR8ThtCbBT045KD58T50o
FzXwokNVo58hXKSn0ohVFk6WSDuTkLr8EzYEyq2fmyBebpKCOVTV/XSyGtl+GGYI38lw0t3XQywe
Ytm1e9sr/6iYsmLCgRRX3RAnhxtc7uQ/2+Bjvzy+pH8tl7vZfg8YshBCoH9s1SknO/EyCdKXnkvY
64/q+WYLTMaeeGPS60iV3T9G4FrNTGeursj0c62niIAYGKxKkA0yNoT4H32xbtH0VEWqP4wEoDJI
iBC9QvFKLeAlwSa7p80qbJpQNcYj4bcgAbRxKA0fSCvi4Qz5dHQA5YmwDlcqoB5HeL9hL9vCRnaM
svQ0R+NP82gCNaGfCD5LufWhHZQeAMcUgYCN5F+nmA0uPEevYkSS1NaN91ZVS1mhyiRiRePLlysf
aBieXGESG21Bv3ifU1Z6nccIH7mqvLpPsowQ7FnW5Nb+Imwdxd8LRYRi6Cfkj7Z3UkF8/j9qxmVv
CAP3PChGD/6X9CQ8FSI6ynmiKnB/WQyncgrX/KviBBuzIjzUFNKX8HgLvrvfbxWQ9Sa82/3lMAIK
p0ZXwRdp9NhUeLYekwflAkFTER1gpgRRvvSfqggaNB4RPOUvrFpwX12NPzbuew8oMV1O1dfVIoDL
NlHNISGsFq/8QNe5U7L+kBRU4sxjZxFCmb6NqlsiLsBaSdhqazav500tweaefszLfiFfWJ+Tcvxu
ZFm9JB4uApvupFXdv+8719QvbW/V3y3qDEnLO5qlTWbigtxj2smcQUsGFD+NRJ2ODcQ+d+ZzfrkP
biUNV4mVCEBonyOK8pqwZQsDkvuLULEvr1b7hajKlmU5Esou68M2OfV6XQjHeo+e6+tAc3BVpdnw
FFMPaLSfiSMBFnFkDtv0NSVQ69pk8jzn3aPNQKzzprXXhl7pTko2yvMfmsGip6ANZCLJatlXTw6o
KibyX7mext+Rqg0n+wc/C+XwttPTIg5Zg4kbMCWk8SrJh+NeooNIpM0UVNeoYQe/IcG2qA3Z+Eh7
hOCv5UPftiR9LEjBmbWrlHaNT7kIekCayaskdhvP3TR627kxPikL35Uk/zcEOwYLZjzRvaBqiH1D
8rY/5xIb3YG5BWFtha5KHRF2UsGGXLO6kZW0Kjconfz1t5mMGRH3twte2w3Udk5A4mm+TSeuBELV
Tyhk2KOOtnHr8NN1/PlS2tnQbUifH+6Q3emXb4GyAMJvI/bREMnXJsAii2qejmuz/B30+IDGjAds
vgu8bjWTxNXXWjanL0Uf60D/TyrMPdPQkGABO/EsCbD2Stl0usNhgQCiko2KskALnV9IYxfhCXFw
4Ane4ZwhCxuELTYMG62r2OR+Bw6wNwZb3CVG8IHJwSnNg6WdXVQuYR5a9PuhLn4wZLeH5tHee/oK
YIGA0+G5g9T3OZtMM8Shannb+um1sN1Xb36trMujwDkIu9vtLVd1ZI7xVE6pkV7OTsbjuBl3sx0Y
fpCmEL8iV7JLBEubhe8xef2GoYzVM10PxnapWDoOP3SS9YlVarb3YJyKzUWn5/F2idFwuEL/9hKa
Y9EnGNZexkU6Kmz5bKUS8L6G9RBGw40z2Quie54+oKpqU2xhcLttq0NZ8O4YwLqv6nCw3Ap5njR/
bNexoNid4B9fnFzEJvJVV9sd7J+/6TLP4CujyyemeJYwBe0dpF81reHHoNXg+8pwMGe0DTC9v6gA
rS/irES+g6pYCw99YFpr0BCstn1zf+a66iyYlAgQUWMnnIRj5nFZ9o6+beeFaAfOhp8d//RNG7Gq
Gopu9e1Uphu4R9ZsazuK85AbKDP3TfvaWjKLgJ8C5Kl5A4uR0pqxpXzGuCEhJyDJ1D/4B60NAebV
o8ovmExahd5hIAIU7m7r1mf0FvIDPlw2qQ28u5kNnggrDoIuTfkxxnVHwvT0HESG7PyBJLRmqOJ4
T3tsdVD9gPH65bVAYruvlVfCdacqqNZx0Lk/wLGEEC1ULnoyNekP7mzlJO1qHpLezBGIi9m6rNrO
F9mEofgGmBuD7a20gQOYOAhjeeePbIhvEbDkUzvyA+dOlWpG1xIwqUEjNgYOKwwNPanugux28lt8
Oz+R6jB4bAH14tlw5Afd5oe6XpIiExCacL3QR1rfftRQkZs8C+HI+1KAFSEzKUWI6hnltVNX/QNH
WeYKFQNi39xUkuXeJTfEhyd5rEAL1t4FTAcY8rUxnD99vkxvfU0kfhMKAcDo7bf93WYSWg31LDjh
015UrUNdlz4GAbVaYFNsekPVbddv1OV35rZC79gR/q0pnrAcI3owB0KzsMN8wfhxEHaYqZ1Zlueh
OkzmOoRDoFCkyoi+uCSEqcG4UxKzHdOiZ2gZKuU4qYoFcUJz/oZ+8yPau9ECo71YzX1v7yHL5OwE
3k97/gKrm/1M9n9ccMWdaWLbq6z6s9mS1KAW1ia9hOuT1rrKGkNFjUOQSWEj8EYal8kIoSg8boOb
TtuLjg/QuJiM5MIoeBCTCg4CepiQ/5b/XXXNJ3+tuj6tNpPhdICXDcpXQ0igsmilHs05NcMGzlNa
Ih6Uvp76OyRC2+qQ6v8moRPVScxCebv0pbpBdQ9FaAo5yN49fbR2VxFySxLBlF2Z+fYWCrR8PTK3
4XttiuGELcipRI00mnIp0n68FI3fqAqCQHwKzW+7tZY2m3ga2u5kmrKDjyYyPy0DOVFKvnFpRFV+
bM/eHbNsrp0mIQn8/WlmBMR23GJxtfYbYn4ZAVmniNQ8yZ3KQFeTmmsMVH4UE5tfU40wjrlVZqtS
LUZ0IvjKlFJsCRs/MWujU8mqCArFp3uSY8eenHIeux5o4IrBofzIURAME9JYwB1a87RBej70HwdO
c0s2leZhCftVrDexID8SISm8srwuKoaMNHyO4GnhSqLLLj9HXFr68yTQDRcEPnP6D3e4O74MlzQA
gmwgzcnlU2j9iZOcw5L+NxhfeZyfltpFTAMV2LbsRtbcSCJYTL6Gs360bsAl52EAYxEYBWLlV1sb
4yhW0KvJvqfCApbNqtcmYdAfc4ClSTEMC56E0naBUVv0MTZKUqnl6tlA2PY7/ofM2i0CAwblCRvu
Shup4cldm3Tm27Kv+t6YBh3h5Go0O0wUJt0Ud83hrqkvtYlArY1TgWHk9hgZOFatzfGGzJLVthdS
/oeLWqqaY9jy+BaURAOn3zeYPaMNjgo+PcyZj02yAPdkFnIkFQUrND3vzi4xbykxRpyVTjIt1bT0
6pUVgOQiLPm8ONXZINDbTvyo4uIjs63PS2scVCns8+cMUKvgjdDPdWJEncnV4RHbkwnMBwVg20qK
rlA2oj5UbX2DKHO8v5BWWi1+SY5r64tTbbiMek1nS02eZJdTDkzs5iVMJ3L4u2Qfdi/oMWNDyyrU
iyCCwT7g7jPWalQoNk+5IsVd88fYlNKgjizRzNkegIj8dNUw47PsfxZ7oj5ORqAv0U9+cXgrBs5B
rq/Kxw1BqoiGB3Vv7IvFvbNUrCtzU+FTvbDbgVadLSCsFW5eDDZQ04TPmkTanOzk5R2iQ2xqhxq4
se7FDVfbq8ivhw+FuiGDrQdeCUcGpH7n4CaknMSkjjy2dDd77ZHhbH1gVC6ZJ7uvkLBVkpHSNZKi
23z/tKxnYcwS4QXp4YnU2oZ7kWx0g8UEfWQvg0nwmmt/5FiFvcg45afVClUuJtjHC/XU1lUpcW0Y
hDJ4UO9h9hhDH2b/YM0zkIs554HcVIaJ1lA/wvZkEzsTZtv0IBrorbU5yMWvqixjmpz2HaQdSfQx
s1ovwHIelqzr5jGa28oPrbwKqezwBSdDotWWq7f60rN1nO0hcJZ/aSMSID09HJya6C0u9ZgoMpyH
cJpDQwyiYMCl2OoaLTme+q5FgLETrWlrsU1+UvRGysT1a9ccEo01LxcWvqvhYpEodG+xhjHvzPP4
f9NWtfpNG+vRwwUHfLZJz/NAi+5rJKW5VbWLPn39Z/XPvGTzHry5sFlRK3fgSVTdvLyzV8EhPEWn
8h1Bd740exysDsg2jPcYMs5hcggLvm53+xi7XiDjDzD+AhfGhF7cHRSW8u7rhz/AB33dEbMK440R
frzKnmodwO5WKuLgO9aUnHjD/sm5Zn0ucDa7fQ7EFMtnRu6CmElWj93Q2wpP0JW8OSKBsdiSjPEL
bypEK+TOZaLkDn5FoBcaoKOw0iSxYFcUE05gvgt0lB/+SmzFKwMvgy+HOW+5mTSritocgAyQyp/y
jf3N2tg+6AM9i7INuvWq6i/O0uv26/I7B+K9fbkr9LgBP476tHaInwCVQwCMY8yEfo01Jwt1JZDU
1X1wa4YH062bKwnPaHN2WIyrIch3Cl7WUBIOQEBWNDF9ycS7J8Q+KSLsS1TUGkqnoN8Fnpr1OPjF
OUFdDKJ85CCqleAKWBUN0/f1Qte2wJDTL8KkyxLK3RpSyDiyXOXEbrz4H4kAr3EtYadxipKzt3GN
lDITUvhgoOQKghct4vpIjc5QaP8QTQQ0gsnBdRIk/x6zR8IW4DyvAsAeDYUsisOlgGWoRQQS8MuE
iouZ9Q5Y4kBjEBlq+LJ6pTXDzxWsgATB/UlDWID0atF9C88V66eno76y3jJnqqS2O3tVfhIGuoeM
hOY/iyqkaACkLKA0kVHVOip/2vtfFu20cKaMP9zgI0ncq6ffYZ/H9aWmSD6N+Q28pV66E1qgBRWS
BSooL4JVqI1SH5xjrhsEwLCKqPYLx/kF/jGIGERPzMMbbZolC5tTZ01Gx5FeVZ9p8NLjPgCiaI1S
B0F2vRzeT9kk7chVSU+jyZosGro0AI5d69nVj8rMwUZh1xSK4baHzCfgjq7RGdckjDSlfNw4jKuF
cuIaphIeA/Su5wu8xwpev047xRBiDsGAJMUUrjAJ84T62fdaKWZ3ZeBQYln8CLo1ThmQtSEloRyY
Vxhz4wAxosdPYasDQ3M4r5GaSecXXOxV7oXws4hxHb7OGN1F9rLmC6jFMalZGGtAV6lo6ZLaKESv
fPYpYcCkfcWVcGTxZkfwtURXZ2u05CrBlWces1lVPMEMLz6jw0/nAKI1arsKahUsvL5GbbSKAE0i
Pdbx3ZYwY44B0oTtIA9d/udAuUpuIz5GPkwvKETjl5X0zlu5wtuesYhkNfgSYcGFxoNnHWqNt9T1
CE8upnPOjRFSmW/n0uvy9KQfoLMTKI+P2u7LvWNUpa9RnuI40+zs9qNQQSAoZQHLdcs53hvjYTLS
sJUjRdoVbF+1tblxddcM57/AZ5QFstXNLUR4wLpf4/4lM7Zd4J8WrZ7fx1kmcxzSmS0gP8npw/82
piZ5aw6aM3pPfNwh4wTqvP+VADD3W4SOTNLoNtZMF2y0pD+Jt8rM1efi9Utsim3tnFmkJv7ucs+N
EybvTglQMxBNxydu0OQRAXhreW/0k9flsRN8YBgjgycPWeQPzKtIKh4zoGyL0dBJi5bOGeb9SYga
XyN4Oym4LOJmKtirx4KuLtjcJBdALq8uBXC2be8lvq0qAf0WeoG8BqCeSH74N+v77h/5lAHMkWCe
G3tgfAkCVEhU/jwFdRsH6ttDaC2f/hdW/qrUJSwM8P7DHXgspjRTcfx+HdE1AvsawYw6+nZ/R866
Dw0I3I3XIfMutX+U3oKEfBkeHtLCkKYSTkMZj/R5JWT4qb6EnlVF3rGXUv03ZFfFRYxc00W/Vn//
2otFrrHIV6LX8ODaZNvxndp117nIKhbU499fQFS1g+z5UJG1eURLr6oy0loPcqlZhAPWjnZi1DJa
H2sx/oI021n4tI/eZyo8HQyaDA6CDJCydyHj8OUoLiHJkUqxo5TiMTKNUz+69X8J4cXdGOzzMWI6
b3BRoWNNxYxBj7FBKltDgEiMjCmLoVG5MXfIxEZyEK47hiNYkRTfbPGBQnhSoJk6CgeCAEVwahp1
QkYzSFIXSKneEgogbHHZWm3rhAiI2sRcvYjU1aDJRwBLt6dGT5+A47nqlBzpHVvRow2NqWC8kOk5
xydLrpX8FR7ZlpGXA5CsmV32/Hwy0Dukgm53vjTA3CB4hAeS0a5ij2tXyVZPI5f1nxnEK4yEoOg5
0SMjrMSu3RYO1kRVfJ6emBVerZ4o2aJSalvfZ/XEjyB5obtDlNKCBNGDGVU37gBrBLPMdmez33fk
GFDF1vZcEWv6VO/Nq+qUNvAJ7RpHYS+kJACfd1o5GW6o5EQWyBZmUr3ncFwuxwj7O8kfIqKsRDiJ
4cSoCTvkYoDd/z/dFMSTIlcR6iD45/aMgzOenSVx59S8KrS8hJnmDFK3ouF5F7ryUyEcsRLz8uic
4lUyC18ZADRvOrCfc6Nnkp7mnsUeS5+K+ney6Qp33RH0fxjsKYT4iOEP/FmCVHxoUhDQkKlXZBmJ
xFnelZP/vEtZ+D9YNvGtsp0xo760ytZgPrkKTW1K1KAvs1jSCkGAIYinWn/qCyVOgk62ROXf3936
Aj/Efel2rjMO7kWH9j6XytzfWnn+DfZmAbNREspowCWxQ3Rs/rYA0Z/B7I4BUSQtcvSnRWUGbDpc
gymidY3fdq4CRgm7fiVntDY9TLlDQb1Z/APlGWawtfqd204H2KzptwndY3Ky8guGECX6LDwzL9ch
vU79Gw4VQcGgbYw9H4ijOp07Fq1Yoq0r9xN2IACUqKCkJICFG2Vn42KFbtEeNOYRll3nyJQvGTc2
2begizJaOAWfxd1LD+i+IRijTN49kGqsHD6OJKVeLw58v9WnuCRE/Ib7Cl+HgXL7RoSUgFDashHS
m25HWgMi+APgUNKL6JXXfe9yL3QrdV82LZfjcmmWgBi3T2MfqB8sH1ZGWi5+Qk7nd5EofFdwvNfj
XF19zGus+DHXbZdsbRkwrxM5ITNivg/uu0hvd1WtOE038cXuVZFS8DMb7GXPyw+SlEi63OF/fDK6
kBwvZrI2RCZTqhkVI/Eq1UmgauIUEU0xeKuJDIdODsanisHtvZV+mdqdCyZVYWXDdsq33Z+uHH67
q9NR3J67Gex9wmGYx/LDHze3dJ75NAxxcnup/hH/cb1Xpqu5M5AqdYeMkhhxhIkEnwWPvtJbsnO0
YlINUNViFn5ZVugJl/MbAHIJEVIEwYdniNKfQpnI0pKPkq43+eWGLDIW6j5j13a4kG/an7ScBVD3
FAnn2xLktneOVmp5Fru5W/9KelwDZWlj0XfDRq98mHaurnLBjopQWUxkkZ+hi57WfWQ7cRxb+Orm
mY2tqbajfQ6d70Za8+AhX1T8bHbE9SQ0cvwBuQsMC1CnpZdv8sliH4NkYLu3Vl4aLOKGbGIea6oj
y9h3TfHCL/NG3APsQG36qFYAumjgvAc/mcuSBWJ02wINSkni3I26EBEps4cDrO+r6q7H6eKPTq1R
M4YMiHQ1huwjSMuX0U9cgzjv+VoXvFFpbqeJUpDfxLM5W7OEcVv8jnu9Yg3062RRValR5IzXy/e4
CVZT9Rj05WYumFLcoAwthgziTChjYqqdWWeTG3dH5VqF1CXiH8bGYq8ccD4QT3iTDiYtbFbrOJMV
KdykTiBVhvghnplgmPoIl9Db7ylr2DAU9vZLWElb+RF26ZxXg2GgNNAgfcz0yDwTAWwRaGxmfbR6
fvQ9qKO9sDXiiJ8y0kX9NXQOQKTuG2huDuIMpFH80uoR26egTIYrE9XXheyB7pijDemWu16ObPmq
CcwnbnS2CKKfPK1F76S+BzuaVriayLTBMZC33HP5wGGmlDJ/0Db7XfNl6XAOX/TTF6tvyEvbejqc
stCogEiAqXcRPifYOa62RtSLlgl1nZTMpGMYdnL5hdq6GO5f29A0t8xJdoz0bFOooBKyMRdgsXEk
2oB1cQKYgYZPsIDIJZ2UgYQe3BTGUhM7/ccqwsa+5WJCYcoM2gDOTYw+AmVlXOAq1ho08J5xgBN2
1E9Ph+hJXPWziAyMZwEJrr0HehYyQkenotYechp+smLDFpUACR9ep1FUq4Xkq44CxaLButVrRNXs
UfHqFjYnpNDrD2/0uTeg32DOZJhZPnpoqt+NNf8/G96R/Kq2vMpnFLwuko6OhA0GQV1tRgqZ58TA
SszBzinj5HKdzSrVMDcLmebgN6Nm0IyVk80dFHDeYGjVO+DdYLG8cuSY4OdHQ2b4jncc/IoL5HwT
uN04s5KKkb3tF3gwcAkbvtogEUvSgLlkSBDOytWrlqGlehY5gyZsG7SwHXM5no5NZHh7px6Dsdgv
HNAQI56j+nw8azVY8mRE+fPacwNm0YTRK416Zp1dVn16D1M5vlz31Yz76pjws8oRQ7Kafjqok0c2
nGF7AffCxKULNhdRCznO5APIp8XBRAs/n8bk4qzi3TWdJoI5JkwiWuINqhsgfK4Dou/VM7x7FTOw
17sxLH/fAaMpifsiR+8Ekm4D27lmfZetH0WkkyguaPrmxBrsOX4dfPq73NZ5DGg0d2iTygE1iPEw
stBLVaYe66aDmPSi8aezwDlLvbZDRg1ac9HtCsTE9zU7X6FnMKmXLW92Zd2LnKusD8eIWYDPpr2T
PGTvE6VWnkb7b5Y5U5hGN85DBgdm7HcBN91mzdHlrpEMbiIXdmt/M5HgicdcZMkiTKzsA8ZAOF7V
sN8jvgLoyQNDTL3bzj/JO2ccCsyfQKGCeb6PVExhT5KYSO0lok01b+/Yp70HyKhzSCUVUrfvOY4p
bqAL3+eFlgzSot2rQlQMQgxWLgao9LfA17fwJH2gmRHcr4g7vt/RE4QP04HJdO4TKrnYHsLHSf5P
ZSuwjm1iJFjpBqx0n8e68eXotwmv/DSmZBdLaQdNcSMjwqAnm3LxMEf2wPP93DzFWYQSAlP9nVMv
EB8AbmbR1MM2T+DNCDZw0y6ZMFzDctCALCYTKZFUsp6enIBFMMzU7K8vOZAoRk7KlegVqmwJOSzD
MlWSVM9QIEZZ14F96hTujrTvrsmHUxZy/vwv8cXCGyZXG3pRngpwd+BBGqII2AScIVUL8sHh2+li
vkrYzkvmENo33piGE980ZFckKg8xd31fbvwjiDu21zcdrqRYHP0LrjV5jINEF4XfS4bXuOPjYArZ
Nmp7fOoR6P/lvlgoLjoaLFLy7m+3pjPh1xnH2yDiFX/bS9rC9wYynf+fxZNPy6x9Qc1e/fDNWqpr
nfRAzP8bZsdilLW1h1RVzqvXKrXjvq7paBTpvR155lcapjY50hnfOAQr5CPmNQovmBcfcLnqVgqt
SjUxeNfsNbxXPPFOs1tbc4ISt1/mjjOnkLDwkBCnC6N8cCl7oyMZf/6pLWfrryDxvqyDlcPtG1lh
x00MHOTJDlxsO17xoroHJz1Jwk+efKlf4uULTq+t5RfsS3dDspb0KZ8aGJsZy4BaMJ9i54qjGC2k
PIRcLqfFHRew63Y4Vmk9S2mLoJpUriLwOCLMVSQib7uJYQIuPYLreWYz1bj1D53MONWFtd8mX5rq
zZCQ0yZ0a4cJBVcwiGTsFkFF6XSNGMSrxkqi4vsm8t3qX4Yz0fX+DJaRIVJwXu95pVvWUclMWfqd
e9W9AdFnE620AfYBb6yxo9yyg4X0vb6fsYOZuhaSFlCCj8ww6Bu5C18LcegtzBNSY7C6KihX+Zwp
qigfbJ14PKyqJ90fwxZe3ERxj9EY8WCiw3dRS+Rh3ucywwrReSSTF+imQdnRv26D5ZHHXa2SP3Xf
hmnbW4hYcrSe1rulIcVjgfTGpTR4UmBWsgAs/MQT80zHBzrTBeGOFOWiM/LiXIWhBiM0rxi8lHye
7hvRZ4k4KHyKoF9msKcvddIR/AtzGhIn4bl82uM6+FF7wm22DRUKvlPQ+MeAKSTR1Rhtdhks+CPs
MpHwH9DsYIH53OLz3RQ3qUF+wWKz1wvT2FFVmuMf32FyAyX8pCvFBN7FopFcxfCHkeDPMExN0aQL
p91kW6t2BURFsJQ/a2D+59LB1D3l51xP2tZJlN7tt1OkENSRcGkSgbolSz/tF5a0t4aQEP9MsT2h
6fEHTiM/FrDIyfQe0NKBDntEgl6ujqFY+VXxtHLcQVYiza5zONWtc4eMNlYO1TbCtapdTmVorg5M
P+ZcYKNJb//89oc0RTLCypgSYESpaVYwzhDxCIktZmKhSaWYwD4BvJa7Z02nZXmIDJROD8fYRlEY
w6+Fy/wp8gGAW4ucol2SCnfmtNc6x2In65ZW8ho0+mSBbncNbaa61k8Ev/b0shazizu6PqkdB+At
j/worZMGa619gLa9jiCtTN+iHMfLnwm/fpzijUmqcxxrhmjZjZ+gUY5I4ukCSmU9O40K8eI4K2Ri
hlRlq7xXO8+HMh4Trnd1chqtcb9z4qPDrHTCtU9fypZ8mEAGVqNJcpFeZ2p0loeZ/hSeWyDWDDTU
qdpiIbPc2Yx1FjlojKAihWkZrUfcLnyukG0L9h619u+iF/N3lGLDg2YYNdSrwlp1OF2DFd6d9OtB
GDy+tHgVaAYc6dJZkbb9aJpU9QAaPUQLcT3JdfctBw6ADjVBcWrpB+Aw9VmWqeaskilCfOTloZc5
Bxyo2Y2S1w9pIdvFNf/GE03pRGwHkH+PkRYicBPz2JaWRItcXoa6Me7HLcswxcJCWbkYDH2Bl7ao
GQxZRKiG3Qov6U/W3Ehpi3tafQnPsiFrRLDnei1rUtbCNoszJ8mRHa8ipM5XY139XsIymvMknuVV
DNvzSVv7OQEc1O/gL6jp+upK/6gfFHcsuSYCZUGav8Z9xtiXI8FzdK8BYr/lwaV4OKKRoRnPSQVJ
6kG6qxvRx9XS1ia/pEItnm+VukdmdEePP4zcyxofUHUiBg4o1CBe7IxYZimSmo47ydOKApnrG4lP
d7Yj0gaD7v2qDEiN1TeyZAZJRfdUAhtZKnFE0dH5aZDWo+RQapywZ6Xa0aOQMv9g/1NHKtKXmW+a
/furmXbfcIoCfphHwDcjA+Le2fW8gB0WD4vtshpT/oEDms5M7zX3jDNXUCM1mztXV9w/81ereo7c
7TMLlvjX9SCo7aDtgsiHf0HYo20MNLm0BqiIYqIgjZu5SqqrGLQBeFSTeV3c/0/3JT1zwZBNBgPr
4XTWIdbXnX2cWpj7zN6nAFrDMYkejZcZNJ8AR2BIFRvJdyGosDt+h6t86zwTqd6YZyApmXifo7m8
jSGlAFIPLhuqX59QZWEGEuVhxjK9J2y6O+7uDGkeV1AONCjPx8YD/J1q1U8amGSP+1fLGAznGkYR
LHoHGZenHncsL7Htv6Xh9WEEziQqSYTxwutiM+6hSlPEVRIJgn1UkXudq7jOCQGrVJwuEJHVvlOC
NbRhJYuF0ERY2AJq2kNlgQuc186eUP8C/x+korvF/HfvMLdoEJNvSMwrSyLiQM3WoQ2P/SQvvfR1
pU+KGJxN0VnztwjCROdbxNX0TAS8P+f6MVCftcaSujleF/hw2Dkxyoi6SjBYUGffzDeo6UpCB6Jv
L0tvELPTjIsQl9wk0lMkGzHAQ5d/Q5zAdSusKPxg5Bijm9AE9fw24MKpZMLD8x3Of3Qz7N82Wwd5
MhwZN8yo+qQLe3T/nNbo3CaYYV9/punECUQN3owd7RVT9tF4YT5crA2oIOgTy4ohBU1RkX8mQ9xr
hOEv9dKQohhG3NF5Jk2B4qJNREYimk5nrutiW8NkOnb3JJfWrOlbXUHGnYjfkTihjvn4sJnsWKmw
AdOZyaXC+ilBhq1dXmv7VrZtktgDaHH4+JPNYpFFneRM3/41bBUa5UZBvigjBsFdrSN3ch8CFCQ5
NM/vBtoFB4rd25SOh7khgtpWMZdMFk65nOuxKa0seitR291m3izzxA7TvMa4KJNC0B4h7Aw55jv+
ZSSItxxvN0WZHVtQOfiSXHk4by95E9sF3qpLvNI4XhiOjaNeS6sS5MdVb1v0I/fkBn1M34D97IoJ
Y2NgwpJh4JPPFdrnjbvEJrrQJuJGd+beMXqnxGtTaj5rhgYaHXpOPQbGSO5AoqH+BrRVWow6LozK
OzKTYKnkZYlL+EtXmeQysIpfFiAT0uv+lcUTy82qiUhyNRGsn4GjE9XCE77v3tC8cSmq2H1EGFMj
DkyS215dk1bznx9yK5yZK7qP5/TycSMlEOnyqZHJsffRzStDx2IyoywwRAleMXnqTAQbY9sdcour
ItaiT6eRwXV18UyRWhGrfUV9auoYYWhzo3fI/5+cu6o96ENeNBLn5hToOsiKfbFrZ4lR90gjwagD
T8IxhdwVPYIjxBAaWxf5tFTa6M0FdFJchC+Hmv5BlwT+M1MOhx7dNki/EWFsuPk4/nR+R0/xz7G5
ejHU80tQtAglejU27VPOqnkYK/qSdV+UT6UY/HBGJ5e7kbvzBYBLkHwBcn5kvqhX//uqOQVnDeHs
oEJViek98rxsg8IUxGzNJjxJgrsDmvId/KP4WOLXcv8WsZddCmH6mUQ935/iKqRmApXaMtmu27wq
CipAEUuCW3lEMDkA2REFu5aVikinjJjHbnBXX/XtnDKPrwd5Xh7CPUKvUODOLVsjeKz3mWo92gRB
K7LMrLtgptbYg86wQ/2TiIjKw/OuxvYF4aJbSSqZEqtemF2Z2fSUk+uxp+a4xIKwStopQH6F2cKI
BjvqbB58ikcJSapfyIbD+Xx7lIzhxj3AAaDe30kI40PUUtYpWm6wNrbIE0VjTzYlFeMs9xuj6dCr
4NyyvQ4vJa2Luw00N105TYJY3YBpymZrsIBcLHTBSjWQgUJlE19vF79ubi01jGHXCLbrD+NJIy+L
iFifLWzWujRwDDH70VR2lc+TluhuztY/XiWrt9TfqKdS9no0yPN87JQO0E9G3adLDA4j0HBqZqP+
UU6MzEAAha/8yjISTP/oejKYU56DXTPSu5lsvcy1WVHlM3eESO35frKidTZf1mGIhm6VtGOQBHe2
/ny72UOPL1LD/excuarTkYR2UVLPENdll/EbJ4zwwJY+8b5dLQ4AB7+LcJ1x8sLTw1SJEfxLhfyn
1PVp8uvbgpNvm7GTT8cUCilNDa9nlIFeHhXW5GnSYPn4tNd0sLcDoPzIgHWLDqB9TUMzg9RwF3pj
6gqG8RhJS6g+TinZXklr4qAagvd/uOLMLSg/ybuQK9k5MUUvw1wB+QhawMnT4zcAOqkP89878QnN
EwQtozOPziz1UEj9zbEgZG/UoQxVyWDa0vWBIz9wvt5/MHloF+0AMzY5Ba/Olz6bSm/ilMIkbyCF
vFsX0oMKXTY6jR//KA8SABLfulne9zPWbn9zsHXztSeRBAc0YW9rVpuqM4i2f9Q+Ph9tsnQSZaiW
blQUozcJnNxZ77rVNLnMNZsXIAsATjPP+vgVImGHVmUcUBOM1WxqyZEGCeXj7oIY/OjKCYAB9Zsj
M4dws8tNotm1Tmk8L1UdnS01RZwHii7kImEl+MTTcLW30ytXDpMaNuaskK6uyggwzDTT5W5TtsiD
JRERXUYO5YyHx5CvuDWASC02Bu9P3hk/NkUvTS/+PaSa7snH5jm0SXN8UzlsdtgrkkGsPqih6JjI
zoxeW4nU/zu6H/NyJokSnKXDS9TQZr5YCG4KI5r/WYC33z3jWqoWhsr8C7+BgSiaEx21Ri1eBFsz
NhH73/DBzTbQPM0hghEKfNOuJgmsBh8OMRPgytrlipR2rs222Vdrh9Te57o51QfQwvR2k8e58P63
somAqAUr97+OJ2qv1xG2GtCM22mszTgjGNn0++5EkHRLZGFsWgL+YRvK+WmzBVqGXOqxbjPO+xhJ
JEbPckBjpcA07Ea+qKsRs1f6rhZ5wSl0//WrLQ+tCf7kgX1LuhN1DKHOLnIfs9IpC9vOdiT/7d2v
tspLxdc8TcZSVY/cbqjpn+KlM/gmPvYZhVA8MgDbKfROqI1rqCywplseKZnj4XEJDtKtJ4UmC7JY
Z5ZnTMCwnBcZXDsdamHFMJqOypHUsojroZD4B0OiYVQAlrLmZYMBttd7NK9kd6KZBWslSEq7p/EY
g5jpmluxmn/8ku7L4YH7dtwnK4SVfTFEpbKPumNdJfa1tbew93KzbY7fLA9xrd08u+GKyky72WRQ
yjPbB73DbR7IsJFz9/Viek493fJL0Skrhhs6R0O2W9Ih5mx9NedAK40PIPJtmg0Z08GbtQn6LP6G
CTV3ezo16h7yTcV2RYzp1p/EGFM4T4vjLMWxxfvcSY4B8dVAJ79uXq9Z5pTGtX9yB1mo6oU9ecpO
upK/EU+ZsHLqEnf9zIBF0mDbMie4mk6clsy642pu9PxxeHePk6NpF8Z8lqkStJp41OB49tCJTWll
bc9JsvV/JtcighRe6JUYO9zlg1OtTj0jb4dMuYMwojGzl+y7DIm22ZrFSOJ0OK87wQ64XIMc2z1m
iVXd4UkGii6AfU8ledJNuTBEiJLrAamBQvgAej3dAn31zngLfCPnFqQ+RODiwAAO5R+lc0r6vGn9
zKALs2E8zni+fjFqRJAUTFrWJHw2ZQdTctN1bIx+Q1amN48EWdiMB3xBdDfwOIWUgoaMtSUInxQz
z0ABWUuIrckhtXjl6uuRxYultc8YrR+t5dVLJmMnnvDFa9xugGVNDS2ZwIv0UX9yMUj6pEBrm35H
1hkrcwJOozdlI9BfcfbA15HdRrunJ27QjXajlu7FMXjjQbPjZ85ZiRjb3nzmH3VRK552ds4ihb4G
b0ZeyIgDDnwSjhwhN2gIEfud8tmLHx0a7JlWK8lo5WPhBThtNBjwYp6Ty0h8Kum585GAjrvCUk0m
UsNxDI7WqMANFJbGPNG9EkFo71x7xXH2kJHjYX/qLoWe4zILc4UenI448XQcl5HLhLJNiG4+6Qlo
Ycs3GJPTFqtaZgdzbGmReQ3DodnKd/dtQYRE/EqVMksV7AcYHCjshf03uxs64BbfPe8rHDCuSWHi
ThettJSFldL5Epmq6Sjqz4ZzAlJBOeasdzks/LuEW0OS9x/fy2Go8yB4QF2nYGAwmIthpElSz3Fr
9SsM6+bbjKuCuuX+4vEIoElWn2Za8o23ldJ9Y/VFHAh4Pcik0wV3c/3fCWHuKERyWOwnj0R8P8pm
pK8mSVlrxXbZYk0+ellHmkfgCPo5HbzE4JVoeu418pEKCeSz1b73Pq/WJ6MRFGi2fZEqvWi5pxa2
mLa6+4etiz5aqR0FysQMXmJtfPUCOd6Uv0fNeaLFg1wjxkqu2ohzMU4JtX/S+dQEoVXz5D2YBXuy
29m2ovcynqlS/wwVrzRKaeNBSM58VhvCh7iK9Ec6UfGMMQIh3FDLUwtZTPIno79/WP60TrON/Fit
9NN7FkE3sPRbez1TRh6HViHkuMlTLNufqqXfT5DOb68LlDZJzrnkol7bOL6fRnc9gbpv+GWc+w57
v0F9MYBoCBOFK8nLn7jq7okpY+tGYzLtKtd30Kc+TdKj7Ek//ldP2DLzv0JhP+nxFZx4lDCEU3BR
CA04sOY+Ei+yjxf5zd22gVgTBHA8thjewqQ69gGZDo5GyaXu6S8qXRa6qfj+oNvCLyGEFLxcnokm
bV0e/hO6Z4e9LA5K4CkVQOXy0V3Qvt0VbVxe5bZXMV84kIgAzt/sJFLk+1mUc+ykHZC3oBj9i2hB
xh86JwUSeeoj9SX3SyMqwIiqd+8F0RQzuiuVBrUqjX/uZ6ETT9skeUt+QbZZT3+NFKCZBuo2lufP
DRj7FE/SD5h4GSwQ1gs1aEEBQt8iolXM4KybiHQrRimNvz2iIEVacfTDHESFJzDhru3p8G2ulPIK
nRvwsk/+XoieRquoODDQFS1VMoP2E8WfnUopElwqMGUINilEMoXMnb4qouqivg1w1t1gwFEqS8bo
jwxGHx3nhmemjhZh8etK/JIzagZqMHpleJZbPRaQEevnBzRIvA8NQHOR6ORr21M699e255cbFKB6
SEGZDLRuunu6d1M7Lia0DKrIAPB6MG6xGN17bxY38AMx0NoSjG5fLQdSh1CQc8Wq++rdtfJE+oMb
A0dLI2/qwoG+urVGfec6g0gSFjVbct4v+RGZFyIQwytMyaDUoZ96ifH8QIiplWomXjXXT3u4PPRK
2XkEwjEkHGiC5okPU9eGYN3lWN2SYKDIgmLPGZJ/9u8WRenKUO7Z8t+ESp79Pz4xzhkPad77tMj6
0SURlz7cIiuuCvRCygNr8P3yhv4yt0YCY6WFFg4hz48VyPGrNWHdWv8pF8qZ0DwPA2R0J++8vScC
OIkcwguB3R0/a8DDRUhDl5nZA7Htih00nISSxtmPSFyyOMpGMJl1R9kSyCeA+fdRyppjp++nsb1Q
+6wa3ZHN9t5c40ULt4WbbtaO+h8hZqF+79L6wVt23nbEKSPjePERlwXlt0NnU5EqYusyzxuCUkZF
HCwD0g2J4Tz3naE9xJLiL4T+139HEv+upusUBvX8uzWcyzWmzwJuNqUKDkH5DG+Q8FSK3QFQReYA
JViMdXl7WtHMdOVkE5JaPzCEWYo4sk3zvTWfx0AJ0RXaYsBcNbQZsvav6jq6GEYV1sUifTpOwOGe
TTIfuXKY9VjZfZs4SdemktIoazVEH6xTPnuC84QaOcXsVcCkG8RjessuwHgbljLREuJdw9PahRKO
vjOZKAw0+52ScphBLbTvh3TYiPWq1X84Gj81Stjq2tRJcF4075XFOZP2DfiNF13PZZMoyh7AYdot
BEhXbYguB0H6BmeBcvnsj3hTJAs2XJ2DLoAU2Sk7iqBXrmk/05J3/LZGxpdDAhd2rC3e13xg8Rzx
DeRb2csJy2qaLJ0A9t45AQoXkFG/JBY5JsAqR4AYbe/HZKIn30HdAKN+wsit98TumQagnAAYxSY1
VPyfEcsxQEz+gfMASpqzJsVdVUB2OGwC1Ug1Q/HV5B5gk7IULUhT1iR5EBrwucotHJ6241q6vzd5
ABYXupCVjveShAWUYgStbRHAPYPn9PXjzerY4QhTdbJBO2AsBpx/cFhaNhAVYPLpEowdPSCuxDCV
tKQ5rbzKsodzaMBWjq973L9PM9ytZIMaP/t4TmA6udPHvQ65uS+EXrNl3C4QuBlK0znuMMYKZyvi
gTVmhnJouAnOkeff+1fH6lfyTETMjh8q47ZFcdcNKX+6sqQvy3mgT33FimhxqFYtECTJzN3Q08eP
3Z3uXx46bAD7W1U362nmxgndLMzHyXCGh+rULRrXtXT2fjMocbrPi8YU61nL48bpKKGcT9TDU5Pl
/GNmreAaCSTlslwDnX7RZ4Ltwz5aWyuOUXWqQXftbwPnUTSQrzf21DiqvBTSGiAZQWakULlhnmgm
DfsPVk2DBB7dQzVJUq1h3Z9y0OTB3WLiqMa9SyjbH5/lKQEp4H66V2m0+O7S9D7yGyhb9Sdw68G1
IxrQ2Sl6qV50NM/SjImqi/32HVhp4TZWEkLkcKHyuguVIDlnGBDej6ZaDlTIjYjVhsEO9jHAlpcj
tD4aWgPUKMYP1/uQWAjlwsrJLEU76ZVgX0ytAdAOCalIy9PyUgUddIbdtGhzKX9K6bwiwC4ST7uw
Yx0D9+grzB96vNO7BXF390NyRanyy/TWZJbi/8RDPow0e/jacNiymTqzbMUOEz/hYUYf/iFhGJ4M
zwa8Pc1VMD8bsThbVFUvInaYcN60WBTAjkMIBkixQjTbvCYFx3/0M/YyLjJL6BcS6sRptb0cy/qB
lc/roFT7OZIb6gPP0pqiwZFFr1XdWzfjvZM+lyClho9kvCJAAKIYxdwCZQ0dKfyoHtxgDNleutnZ
uSV9UjHC4J4X7OF7IYBCmCea4uA0OnRnyNediKgE9Xrd6oFiCO06pcIBRhNDbHaIsaF7Y/YZwrcf
1LAHfoBkIaAXlgSvRsj2RfTnCJO7BAhchHOeImmX10bLkmKtaBWqJLamrMCDwIiBOMQQMvQNulq7
rpuBF/gjYUVWrEr7TDads5xUOqoXiPi9wXOS4eH/eP6nsNllXGniJ1JurjFM92BMDX3FLBbeiODm
OTXRgKDtVS2KEFh/LBtSFykNUFSRkH2k/jhB51YeET2ejDs5hdedfNCAlYbIrmXLgiY8V6sIJREx
TZ66dxBpOkWTR0iIIgdYciwX2eYRJL5EDfH9CFfI/WQwLBLyLxvwRbaUMX7W0qAiinMJMqG9Byha
Fu+tMwfuF3ho+ITh9IlGE7uU3gpjK93UfHQi5ziGXa5jGAfCZpavfP/bFo4oe4jUtXF5Pbdj4kGy
gaSm6TB+9I00359uog1vlxOpKQ9LlJ9UYPf4pzhAwVEp30+tzcPwMgyzZtLuZUjWRO4nXmAo9SoT
JqRfxE/VPN51LHMUHOSZedMgfP30cuTSsIR27UqQiNpYyJmQK0sVYi1+aYce4gj+GuXKBnT2YIiG
2apu8CcN6yD8so9mg1s4pvwck30/Q2MrQg5Vd6wdkM95K8KIwnAdQGVhRfxtF28/hIFD27WMTfjc
8GRCcAI6R+KpZFSQe53gtq2eakI4EaYTUc2KQEgosSMmBlTPVKF0Aiacqmy6+hEkCgB5rrcLfhXc
GR1wigN9jnVJT0L+jLEMb4BC8rcv20hIQVlnc+p8wZtZ3W/awKUBHiTVZR9HhD+NNAZPjL3pOvxu
2pyUWpWsmlDYcewKpDYAnpmiqqZaGzzvBWXLix7gRFalQAd3xE5cnx7pyDc6qATkbCpVtuNLeTut
pOyQwOSNtw34btFrCPPvOrn+cp0REr/q2CaSzRbjng5JmXwSQIIAftCPe1HoT1cQ4rOVqxEegl0w
qPQbU5mTeVyhtaOhVW4RXszFvevw/JwNaWYzQDbqW6VDRWmD6cyymtWpBAZYYRTjpsBD3PjiOr4+
cj1tyvrymzd1o+JSTC8X8k4u+eyMp2/6Pa10EaSWpIUNIKbyyXjQuNgAzdDYhsOOTHbTo1BGdqxV
nTgJ2E+yA4+uNPDcV+vzlVUO51cH4roAp/O4w7qBLkmwkBp/tmJWOlEzKx+kKLBKXTNCcoF7q/JU
U97yPiBcAFsjEM5OofZZnnt/Z0VXS9ucTa4ZkZM/jngHkpPmDY/HGxMXm5R0W43/NWsYRiTr67cs
nlLe3287ZPAoc9ffYYL6r3TEBtguI3MVEkktqXVSZaIT7xKqOsqrQqL6Y6lyOQgJ3qHK8eeriFJO
cSQ7l1AzLlmm3Am+EgHjyeRJVcChfN0KNlW7uvwFwBVRm0M5DoVYkspp2XQCTr3QHjQPuyY0PZR0
9ClxIXjC0qbWsxr7kOyiDpmcOyszK00WYfkrQPvVE98lV8aUBvj8GX6+uafokK5g5ZYxUQgv9Tg8
eCcUWpA87fjGrY+diP5KM0Xl0FeP3gkyCIwi4ZStUGsHpXPRns05ditXCyuaTkiLabo4aidagMnH
3Al00Wc/CJziHzktdXK9wHHDCnQNZMaYLEdTx0iJ7wCI9AFqBglN5cJRaZenBS59QF+C6RyM+1gq
nj/iGY7LvsmP9YDOqlGeVu1qUxRBQiHr4EYZfO/WZ+iHOimko4KtCfpP8UfZd8mx9EpyizsPr/bQ
rMqqcSvj8QsEv9QnwEjqaL+jJXWjBzdjWssY7Fo5AAuns3iJ5Rwg82Lz6N5SdsxLZ31foHK59pH0
QtNZjdjiPHQF49xfmVvj7RWfivvY7XihIBLo2SUoipcs2BUzuwIKBCuKPq9MpZnKdJz5lT3Z3PTx
XPpmVL6monYQTCpj5gyWZiC4vG04m0snM4hoiFoh+AVc+T76dShxiV0x9s99vJvqQ81BJXN0FBhN
gBkRVWrTzc2BxsiNXwgbt4Dh4vJhtYBezmwQqWrsTSFqFQjri+1oZjEtMbOZ8ib8aXUViJy535aa
AfhI7OwicLziMdUBSNPR6aV1tI7UY4jdJfbDQo9r7VZHYee6u0A4UIRevFJVnGZkxe/oj6D3YJGa
kFzYigGSe1rl3+RoPPCh2LajdgV2nFpbvQbNf9bq6xj8wZlB24lzB8jn92Z3GyLfw5C0fNjGPPFn
10xWimqOYdgplTsQdFEYMkimi1CIK0tW1trml1WcMzMN72RYfuIpztMJDMG+ImM0h5DpYBmgDLuM
e1YnCC8geNqf74GebyuJ2BdLE8Rd0NW38DSnw6Q4VndKi6cWIncgFECkPLekg16SjTRqhwovdSkt
Srt0+Ssmuxw8zeCJaADcnXMW+KoHtdNNUgUotyklWOGV0re3nWScLOwbsf/rcrivThDKbGHiFZUp
+Q2/UUlbVkL8G90JX97Vm/w1LPoxOw6i4VuDedxnZg8WFSUjlbhS0YeV6eA7Zb0CCPsLyOfjR9iV
IUg5z8jiE660oRZe+htO6H84fuvXUwp1rYTj2EUzoamvx9R76hStEfWcxMzpQUZpvid4pONsdRVe
9YigewtCdMuEFLFZFYI4IkHigQptqzmjvVKihVFeMBQRCCt8EGiKLvIz/9YpsFh2NTp+ZkaW9PFP
ngiOhjSO1g/rAiyYfAgYYrMew/+eAThC2N/o5NKfqkzXdwfjrHZotC/bbpIhOXt37mH56xFy+yNv
VsFYe2kR7jYIR+UzLM11K0ejA/sLC8+v2zOwLaaFM97n4bQY8uqonmf/6YUcDG/Hh1ck8n1xjAe6
7rxl5JNZC1iNRtu2f6bfanjOsXRMyHJEVdLX2my6qaBPUAIzUXfLD0pjBdMbRHxI1tfF3YFDL6B5
lqw58Lk8O4UkM20/qc6HG08eKyAg5GT9r7c7AfYBjLcc5+aEeQK7J+2LNeuPT67nUzregclH1rBS
G/Ak+2WsoUY7h3dZQQ3FVzHhen+57wM9LUTRjdV4bRUx+/R2adeizuGD4tu2B68ovM8UW215FuuZ
gZCHx+0+WjUwNop5MUOg0k7hxd9rYqBoWJnuXy39aS2d5NGFkDJ6Nz9t5ACTrMaAzJSKHslEtSCp
lskcMNSq1Efsr4zsi60qWOyHuJiiQSxwkrczw50vD5J6q/QnP+OoHh6dOuBbohZURBpEabd4++JE
Uc9n04k12t3liWL5eoRpZRztnP2wZ8OUB6AMEWDjkDGj5++Iee3/yvExMtlAvB0rBhnlddyFhKVY
8YZuOaLkxaYxag4Yd9VKEVIgZuZMR0H9lTm6ffMazlnP4I443g8Rs0uLu1ngSj/zta8UrqyfC9Nr
o+RJmbEIS5/xZ7rejZqCQpqOxcQdKOOk4CkiPtcVfQYSTYsXbOydKUyRGIbZcAhIMW2+B5Pwzgs3
C7eNUaXxeVqxeGpoZ0135E+B9ESx3kflktB7rLm8CxPLcTCtD4WQ7ps7R+HB+jJ/YU/7RrPlMKG5
F4m4vzU1cYkj2RXqgOrUlg48dGR5eK2+NrZtvMFRRhK9qNapAwW2lMMd2cKBEBwdUYkT8rOLk6Gf
VTT7y7RhbiWkFcIWi6j5baJJ4bAQqmU7anQRMNo4XP+Fd3cwjef0IVRF17b8xOBHw5niDY3I+c6X
bkhLZAU9zEbzPlSe7W/ZLtfgdY6IZbVrZ4dysdtnrraASE0SHm6QNzNEjoyc01Nmmu3MOX9lfD+j
6PeJGv+/8KtLPsYhmYGw+V/4WICc7CHe65LjtogIi8cpi1h8bYfs+/zuoMcm6ZFtmmyXyyKhjoAI
Z82GIqCDXGRioRoFKb8gQXFx3P8NwrUTO3rvgQ4jTpzlfHUuH5OwJMJ8oOEUE47mlE87Ftzvmd4w
MlRKk1Y1bnfxo1fMDVPGlvYrrH0roAlme0TmNCJ9V6z3cfM0LECwTeZ0dY7e73PLj8woYQ9k+kBL
jYDuPlHHNyGQ5MPiYmeiBIFlZCUNlxqmhf/WFD5c8f/HsEfvisyllwFjKu93Hhdx/CZV9RZyqoTM
KyoidKpICAmPFzCEPYqxx3G4kHSKFsxmwqiVtKgqYFL8BNWq84FV5fhOPnigplbivK2XjtpUO2uj
M6ott6HvOx1QZiCe5EUyZh5yuA3kgamOCbako3OzkMlaCduFcScLq0wO9yIKqZ2B29H1HxvtwgGo
cx+yhHuGwRx8Etw3ke2bn3BqrQhJHALbK7Ucwa8/7r8wBSDIRm+3lZuRgaUkEir2vzWQ95Vbmagm
al+2DA8IlcI6ZSiWEtoisMb1BHBz5H07EXvqM48gi6rwBy0ANHKUK9xyu6BUZ4s0Qw7s7X0pOxxD
e6AM991UvqMxyoOgBhdgSZXAStxVHqvJQCY+4lFgCWlqFQUwIHftRP+myRD2dqXl5kERuWiy5OLy
N9Gb7kygJ/R6yWYMjFezEqExuyPEGS5vcfVU2UQkESkjXgVdrG1bC61kQb09LpgGVQmHtbKLR1BH
k8AiUiutSN8KowizsQwIdbWS2hEhG0YxLDGlVHcKOL6PBvxSDrgn1SkiYZYXzfqm5OgWEg7nTZZQ
mpePvlYXZ1IAX0AGVuKHUCzkfMZ/X2FcAJvyirudO37gYiO0+QKq5RQoLwVhCD4TNmH43uNOSk8U
tDEnfuRhbgPS9/OScIzX2chIKJFh9mu8RJEN03Vu7TdQ99OcUgnwkjOhuseI+15iKZ1tUzBBmbDc
sNQ4sihRhw8UM5Z5lmKisGTNRwjc2FkJ7M5lAelu7jOVa9mLhoRxIWyo0hVVmK+vQkb+E1fkIGpp
JZWwqZnad5KC9vTs51AzHdq5QT84xAbJyknsiQkPDXHjrH/H8HVWXuGP8ddB0jCuqFKJglKR2ocG
iudPLbqaARxcKmj/GaBKcf1EgH9Jqm56xGrawlKnbYkXzNNBQDLOCQw4KcbyxU6lYguyG+hCdliT
o9ETsoDohLSUj2z/nLdy97EBdZzfDuKxP32LhpHXHKx5bOQGsyOwPrbLzw40ocFDwSkoGfpk5g/t
gbrJkqtYVWlNHab+mMNvVYo3z/j75xXFY+bgn9VanK2jzEgdDyRXpuCfc6wAgPZTQj75pMW0YicD
Tf4tWVN3G26TRwBTsOOMORGU/uc93E+2zsAWuDgY3xMdqaS0HndaOHlVX4GTFKziZUDNMYmfUXea
BTh6Nog0MKMcMbfBW4koRbmtRa/sAog/GrKi8B+PclV2vcQulGcbTPRW6eSp1P+7QpqZ8hZyaknF
h19byISghSAr9fLSyzf/BYVFXwrA17hiJhsqPWm4+fg/WSV9QHW1Sbn5ejiVovjoqD9JSJ3Qp95J
gFoMbimGKbo7oaKl3q3WhHwGxZIUB40IDAu8op2HVY4DfDSm1hBEORmPTjDsGwU+3kNQCfTUr0Qe
Sm+yALGSfEkHD+aksAMEdivdbou6qlfq7SB1XD3UvIEfh69zr4MDtHGonHzF+Nzn5XlPX/19JLdb
D+julNFZv28DGRtlViZUGpe8hsZaCBNHau0E17dwvMLjxbUpiINaoR6EdtoxVGpXRJ47RlGJUqtc
latS9ZRio+gMq3RIoFt8WSVIqLn6rkYJ1p2HJkrGyH6gp+Rk6nYMjIb9erD/RQ3JMGxcztHylUjG
38yuOk9bewQyW609MHWB0LLFhd5mbnZWgju6ajIb4tDpRysw7j5+V9HePjI0mhYk43rpoZy3n3Z6
zZfntW4XD+AK/Zyq/vGUreXGsK0wpbZjsddXO0RPyNhilNpeU6cPfrVMOT4A0VW3b1mINlM3LyU9
inu+rYLXM8f+fV0EbAl4TaWDf+CTU+FFmqaIpgd/NuP+3Pp9WO4tzibTGX9HmmAh35PZ7Mt+MOQo
rp5ze0g55T0tGHWJnVesWzlYaYMlXbqCyl/C4E3xFL/n8KTG+mRJkg9UnwPfgUsDBpPOXFQg16Oy
cnr2zMgdt5D5YtfWvQ9tlvetGxBCCTfoJfPvI6wtUTX/0ArOUDNvpklKzj0P/WJ43AV3e70oieTs
OJZw4kXp68dzqlTUMQcioV+pwp2Yqs1Gh6xK90JlqJCiqilvoTkUbIYQo2+A5j3WnlZ0qt7JfsSt
caOcfGUCmQl07f8icFZCnkmJ0OMzQ4dVmVfI86gQNFjsXvQSIH4RkcUOa3oMUPYavS3/5gBORCMK
9MwF60uEjgO/5f+q6kDh24+e+XOJAGhtfio8KBsXiJpPYjMMEuE5m34+hG4b8gDMBth0RAHzz4dp
kfmjH6+j0XGYQn+mvq5wpUexwufR5cmCo+Bu9m80vdCcUoBAJIWG+FUak3DGFjgxCMxK9qNJRzXh
o7MrPebKKyQ/HnqYhJdGgP8fiE2vpnaxWsdRTYcI9+oWr9zNEnbny+zA0wXqaE1YRWUxOT8coSsE
Nqs4naGxqhYnF0P80jQGYroVi6J9Y6d7p+XmPbDD8U+FJ4ReLjkG4dXsmGj8SPBdQGDZqcQ6diWN
EBCO/FYxoscDHFkw4vQjN9+hN2iyD73R9nrtD7JCijs+jWGu9HzB5FEJvvssVDd+tV1ut10Ib1N9
k/HGblgWCVuHkhZE3JrVJSXBn+rjOU3ocAMiELqDv4u5qaO0xtYaf/7LjCFBxKwwnSqYybmb4shJ
bdwfklXDbHfRGyiduvYRuL/YanqPmBzqQV7Pg9LFN5i2xo3+U0pxsHaDizZ60qv7V4HHPw9xOsG1
eN0qpJbrA+CC3D8K8zQwZUJgQvb+brzZAHx9Qd0Gu0McCl23oOKanI8PYPApcsbwGjbywfPLbj3M
58di+Imxs0AhfgBASpnserGsvR8HbXxyWEQIpyDMz2t44atDGv6f4Q49bAZHx8zRTZ0iZh899ZPT
SFltwJzc+GEpqS1VwgTS5vY0hSNB+yXN0B996EtpBazK2sAcikX6yznfguTvholHmwJgWVciBG9P
aAfAgKL737alOZJSeTneywW6xjZoVzmQvQc7aNbV13QeqcysADgwM2TlPa2w4crHI2JQe+X1FkUL
RmntnFj9RPjMlsSiuqL0AvhgAPvNyxBiGfQPT/IshURy4UPnSDbs33G+e29f9JkVtRip7q1UHSEa
7JjxlYnAPUIRrlgl3BOoQuToNC/Ygk6DkPi8cIbyy6Zp5NsbXWrs295Y7uvYXfY78fz+l6j+M079
ZBzbOoRkf3RznErWVekZk72UpwvWQ4Hh9uhjS4g25s3z2qs5huPe4W7FTaoDqHHoaAb/cUm40RMD
l7SFKMKGrMaynn9rjVKholu/atmV2u4+AghNMPAkk+RLWqsbSm1wsTh3gKIrKYRDNV5gLLd5cizx
mw2fDuddRBrJ54EhnX23W8PGnNGSIwgE0XSEExWGFWgy7fFDHrXiv2h+mEQvr1Ko4tmKcauPWbI3
ibhd4doK+BU9BkksjIrt//G+uKaoEO01fwW5gnWtdrR5Q21peLsjJ3LgP+dBffnsizs3Ylx2kRt0
0ghRXBPAhXoxQyITjzOUtiDGIHGqIjqojJRzkI0U13AZAjnUfe3yd8Ux09sjBUIYh09TwKGbSAGO
D9HBMpUf4qfciH7cBSBKQ5bGFWVjID7hj3bhbDA2GQaKC+pQW7WyZ4cdGJlyjsa6lOWyUo1dXD+s
s6aHCjMUDwAjfeAg1E/WzodJlarIZhyoIKHlv4E6GhdV7u2Gyzs/p4e/rtWllFjkb58gjX5aiUV1
ATK2Op7dJY/dUsvnCvUCAjj8wHdcnE9iCEfnMXnkJGU4zNyWbtReLb23srVklpSJZM58WZSWr4RS
HoINixYTZXg+CTBqi2XUyPywRr8p6ZGVSi/1RiL+Cfb1KfUJSQ28Oh+iYfXNhoEn9pVnrCaERS6G
pG3MWTL7oe15+HE5Taaano2TZ27Mk2czFzbNoSiY+x19+5QbBx0CwOxm8HcYTSUIonvh2KnpDqPk
8TaTEUMqycQN0n5f79Vyl7E5SHJax/z3gh2kNAU6SQWNc804EMbJUbNSKuzyyCJXB7nKlBkJkGbQ
QqonNW5UpF+JC/ok+6WQG7g34fr556nLPca5iZTjKq0EF/e+xV69GcUwUx11/fBNSgByylERg9o6
pVfz21eoyqgmXsYYZHbBcquPoJYIdZamuB2g/I6GVq+iRyCV0OVjYmlsL/U5dHNifHsY+FwySM7B
z6BM4aTu6UWjnff6RZyY3NrPl9jwDmVGJZZKVvmaUYs904p9UlEqgJ9TWyscqa++WoJf8+yvf++D
rNiMDGI9teasrELEDc3D1lh9AGMzwxGrfj2LMbFOjFTkdY2NSifH8PprY6s8Pw0YS21zm9dgZ96U
P7Tuy1R4C24fshRmMCVhA/+thuy3pfz9zuRYe5FN1DeAs4v1062goeY5ZT34n5+Jpl4QGdJD0LaL
qDGb1YvdfagsOdE7L8yR4T+IxWF/kq36HnE1hW3eViD8mprLKUfTCVgiznLfK2QMAXReTdLlKHcQ
APRnVc5oF2tGpFYTzhS4uW64PFCmr8Onq3+9VGFWcqn3tNEt8+YIc9JtF3gP8kIa+R5Ul3P3/A0s
05iO1zCCnrZQ7X69KrQH9JdI0Wrhak9KyMVShESIx0JnsEhNvjB1Z8hht+LaLk2+tWcA3ozLrLpM
GpfxQM/f77crySV3PNlbvK+SFiC47iJv3kPYhk72KRfS6DP0gt3/d8wb1fJ3Tm6r6lL/tRJWAGaC
7v9trBiwHs+1U5S7zj9D76vtx5TRCH9IIHyH8he+ETp/hmLFLP6A0NP0XkT8psINkxix9B6f/RrM
ZW5L8F0zl094rtsuTSxxiU+wIYr4xiaJATKCWE4gyFwZRhfSm4Boe21F3KErg0Zv3hwFKazhLTXf
yLXntEnJ6wHevfMg36vbtJug/bsWFS27IFIHoHD0t+VuW/kdPuihMbISWN1XRGPmh+Tg0Rfhu+cA
iEdS3Yo3pp5NWZsF33OfUDCpkYQbThwhRHjsNHbN2jiHaa8pO+lKZ7pA8xx30hGtvAgufOwmgw6E
ZlTBeyNbAE/Qn3Uu+YOJycFCkg024piA7uleu3vaQDfjuq4Yv3fjG/0wW/07K2D30sz5Bkg16VV+
/LCqgkJsVEfoEnIr3oq3RmO2p7OYSUPiV79Gi3ksxKK9buV0c4fVHVRRUaGhFNiHtCgJZxMM00fh
YrRTH4PtbwkWljYs5ekOcTnod+qt47DkQqRk5PTIjyuDvKJyZH4WSB9qfbvgecwPEu4MyP69Fvzx
k6S75Brtal5nkSciosNR+yo3YnGdSZ1JNJ8VTL7Cd3LH8X5B7lp+tonM2F5puPbOVnBdwUVcyZLh
Oc/xscJiLED3oNhwIYngFjhiAt2AGtY2LtruLmGALnMpFGwhRpv3atZu2zk1ddh8wP99i0FhH/xs
S7yjLL0zOHetLA4C3BNBzrFztjg4q9ybZtr39QYoIkH+CBF+/B7vgqIablKFzNo1sSbdyZczCmo7
niKPV3UGuryhskdmz+OYGTyq0SGHFPqOwRjaiTEAZIJZnZaGvJgjrtaqliiSfJ2mopFvmg1sh4EB
5TqRtmIMgc9sjVEOMmz7BRcBqGgb1m/ICOEY6l7EtArdVRH4uUc9945annmFOZ9Hixjg3fQtb5vF
JiaOEKJPrwAg15ypVCJoTNr5HxkWRCvhsSdtxQWeRiKGQlxss01HzoHXWsf6hto1pd9fPdj7wGOp
OILHuVapA2v+78yDAVEdJuqS5Pse2I/cfMUceNl0pgRmz49Bi1BfGoKDidDtv018YkzAgzzqsECq
hqcmsr7+d8iMTFOJL2sHsm5FjL/PJXI7ddQYCiqv5OOHL6P8daAah1a1o9JUZWR4bE0soEaIFp1E
SBVpNCZULxjKRQEZav2Gn8TDU5+52hK2ghlDBSlOCDh/3q4+jmKbAmwmTka7H/WbEqVwEDm6F9JG
uwI91qMjqqcgGaBbf0PrnNcw1/zeuIX0r2taenJyFnt0H/UH3aN9hkKYzL/VeEs/ED+GTCpPfsoV
DhVCiGen3Dq+vqlH85pCfIddoGUp1NkcwIToV9eMFWxAHwD+mZD7XEqf4+EM6MkNs9TdCqFa6vsG
gYcfCrcDUgcDvNyldJJ7L/5OAlQHU48eOkQzZ6EIjfVVa0GENpiMNCPVTS8EtJWbJhD1ed8xK6Fo
OFcZunBs4mZ7iuQjuJ/i65zaUysmUiN4X3EiQIgSkL0pEix+LDFiTeMUpcUgKCWNqjl02dPuRDj+
o+k0Tjv7RRnOq7Oa376dVPoIl13bFytgs7EATgQz7ht6TxF+qAemKh07yeDDvveDZL3igm+YklOr
+0N+9tfavax5y6yrMqj+HWYoMlqtRCJgyzxfpN9Y4ryAuf9HLE7b1xEnEp0Ge2kIeEu3oDxPhnlz
3cXFTUA+dlJq1YZ/gxC2/hr+EKfdSw1NlbZWnNIKfFoQowXv/DzwGH6lUhsDJPQX0OgUEwcz7UXQ
VtbV9NwesFUraSuCn9xa6Hu6+kFVXDnIarVJmTFVx1ORk4dKWXJtPHsSrSYaDUV/fhFiHfuK3h4i
O05k33RXpzE8VwwjWQEhfYV2wFMs1YInK3XV69qbsrg8pefCp4IlveJ9L4lwQluFVrdXKlXlpGD1
ag9VKr5ViCaQ0pGHZonrsei/o4d77G4zVNFeDLwWT7bZaRjSjrUMO/D3aNEvgOgSTWnUOkPD1Hyl
Z7zyrXMR5bDg0bM55PIiJDDKAgmUlWVGAPhyJKCKzzsK90cugi3qxQojcRxHzgmUxOOr4Y7rEKIN
wcyqMqExoAIGdnWAPnWWrUQ3qDQzLQxNBX4ggq+w4z8diK9QyqA0BR14Fk2HPgxElsQn35W2yJ+c
rQ56lUMcBLStkFcE7/bgk0JOHAU8WBsY5s7CU0OGGKKb6Jw6CO/1s+CFsfitfDw5W4bx7vsQMWua
UwxLIiVZZIbymUNSWRMbjPvfrLSkXyksDRBKrUuchQ6N/6E6nweDvDCUhyMTkE9yGLB7dXhbNvVV
+jyeeWDpyjrdiiLzmPrLWC67MGsOZvne+ODR03AdtvFLGZiQmehrQKch7sTXFdtxyIDQutO87bKG
00OCGz3wvArM22hXeCfP0PXqlHCzxnV28PQYhElbi0PEJSUlN7+XDGZLibD6I+p1twH/taxl6PjL
IKjZ0hyImZTyW+iFDmhE4ig9h7ceOJxelzXT9NDcBsgxzts3Ow0PrIfqxhEqfm0L3vSpIGdT6Y8z
rli3yrbfd0LY4EAWks3kKsgeeL6xeYlqHHN+f11J5eKyuZq2TExnSd9A5V2h5cFDXpIp3rtd2aA8
nrUEoH+/ko2ibYr0dWq0gh4/TeSnGnorY++h3u3hq9otGFu2vbXzfT4YBc9Pf5kjiIy3A1XEY3YJ
273nZZB1NgEtinuQSSAMsDhQmavYfUl+N2aYnNWK6e+rEtd+KarYZPrqaoSpb5jqj4sDhB1m/959
HDMCZgxxW88lgWt4C5bRe/I0eDixNSrdIRqTow2GdSgottTsXewYxJyGPF86dMS5UH13uMHqwYjf
qYu1bFb/cZ0/KKep5xkBsrXmfhbwO2n2J0yBZ79lYtBa5O2oe3KVEKAsRnBuQP2fcs6ee5oINqDv
diPhZkE5pbSZ6eYpWumS+l/LXwZCgbmCbgHR2S803lsFqxLFHfbwGYNFWUB/g9a17luJp4aQOca1
j0XBi8LoKqn8NMuGfpcFG9ZlAnqeIQgskmzBmcqtstgIlk+dHEr3b74vwHUIxn95HRn6MQTyYnkV
Z/0htIZPhTe6QsiXADwuTW0Jfbxz5dzfVPHkHV7t8spXc6BVIcVQWpPVXnFCa+CXAiLMZB3ekBa6
JRp3S8PiTjnfJUIt3ePtTaLzGZFkLqEPZfxKOZyZ1wPavT4jhgXBi1APGA4keVPGggnElibBCvBM
wDKFKfCnlgKEnxRSuxHlBgJiBKO8XHFAYyPfK0SCiZGZvlGdiICRmKILoI4Cs4Hu1QiXkRSjHgn4
S7OABhji+U1pG3BI3/3qoi7aU3mrQHlRPiXtLXmRmfNOdBXk0sD1ag4Pfej4xC5hI7onTXHQklrL
f4GNK2VcWritWRl7oJPau9GWrO3GZrdkfqZmyZAVEwzbKxo79dnFDLPO6WH1w4HKYwu8/6jfqLin
7dyGpalYlkPX0OlrfpUarmHx2nbveAwdvIWnpe5mw+5qgYyH3iHw33aIQ5s4hfekbupHhHrBNj5N
o/nUAZ/5C0N4m8qSvRKEOGM0pjZr2G3LpWPJr4wJrma2Qmz7C+6veZHldGgf0PRc3UiBbsdffeNu
V/uL+1I0STxSEGgXuOuH/bt+BudKUK1sh7QjmhXcNA3ezwK7DBpEp+c5QIdW/YvR6SCyLBAszU+6
ecl1Og1ihkSipAnEfGVOjwka4FHJfkj+1tkEPyKDCFVNp8ijNl3u7js7sG428yL1kfUysG6XydGV
eoSfS4vKIrm/1ATENnaoyzhWyquz44tiNMVxee6sxI/IfI4BDVK8O1HiZK5vq2o3XjTGaqMJKYOh
RztekpzbQq1gMwqWEu77hj555QD40tiNXcffVITzwPvJCm3M43lnZuhGakPnCmiF038EBJK6jiRd
Add1fFDPUmRa20B+Yg/DCfZrcSOwQlUMQEdsdLaSFwmoVdRZGzm+WIyaM1rxFnyv+m4mQTKaivFn
wuy+yNdU49hfdQeHEOPAdmDlwS0kjsAnCjuAIEZiQs5SnQtOHD5boq9UCT96A3paHK+5AS9qszrC
mpRxFdPwOfDhUyNfGIJCshPdtXUOoedN/3SIm2/rbWY2sFnvMlmhJFHcdQ3O4gbtAFn3fy9Ct3Ws
M171Rb9D/5iiEoiJmKp/3fWgMd+PHRASDbryM596dTH35K7aUMDBc1Nv1zMXiUQ4mQXnmB1K0Y5C
p6MKbAckC34Nv0GkeDiQb5wzTM7EcR93GxfSKGUSloiaXFykOWMUAptP/5zqsyVKDykxjO6ohWC2
oYPKAV6jKqkgBoSvO8kyBPjtRBs4IPoW7AjXmnpk2TN5PJet33kimequa3ihu1P99nb+WeCR+dfX
5Wkk0GcOnBNQY87A204IxuxumO6hKB/piVlPsaz5xSoa1AIXihO7RS4Fwfz1RzRr89+DgU5M4aIr
PmnjTPNfS76a0Hy0IoVup9khLjCz9O5erXAmrRcZKT9Am1rNZ0legyfJP7CijEmapvFVTcU9rPWa
Zg//Fz3PJW6VQ8DBgV2moo7nMzadcy4xXL9IuAdkUdkq+IsZTh9gdYFX1qJgXvImiONqPUaW3bNA
O72fvPl0xHJ0i/vM5jrflQL66DsVCBEH2ZhV1sBpX9XqP/bOxhispfdMocTerStvdH7dxIWw+ox2
AIuZTxYewCevl/x7dC/R/8HvIjCNkM0mI6CQs+obsl3adyu3TzpoGA+svl4YaP8xQRkf/ROfzz8E
g5S09dBbIYVcx2ehBeXq8Geqn7Xr2t6Jd7z3n7lrnahG+faTF9HsEW0KDVA0yEUQnOPkxV7QYjhi
RDpnN6HBZGdZP5swYF/I82Cxw9fmksI4SKwchw1ZwTIPjNHbvI9lPhJ1+k2Wvb/h9wTddj0QswF1
nOa8yb6F89Zx6fBhwK/qhZlCJSkd4udwUb6UHe8u67UPJh/KyCV2in8JKc/nQrDUJvwqOo6znVpL
eqsjk7VR/Bd967HRDvFzrrmak/FDhrGehjhH4/44g5sh0tOHY1f3/gTHTGMaMvDQp5S4wntxl4Hu
VPbVnQKL3jLYo0Fjd+6Dbsmm2/DooLonhVEumzpY93GbSRhT9738EVeYjFCVnF8hzeToAyMvvJ+p
H18J9akf933GO25LkUEUS22vcIfRggBPwrUTxBvNihTuBYIpGcs25/kH3NhBqKhpvJOxyGBL+Jo2
vXVJlLggykJZvp54yMUos1nFav5cOZDBZl/uc7mywhyR4bxSuAThsKPinP1ufh6amD+9DrYbhRHV
cpToLB/6SKFpOyiWs6fcTiOaHyM0tf4uemu83+nImFXxVMkGUDDPOU0N9/rPAexMTkQFY74eLHpn
WhqZs9yLgim56l6OBrZ7btoh3J0ctLgi3KBZSPj2bf2d0LnMcfcvFq5QJuowBC3XaNj4xAllM/CO
lT2VuK3SSbIF4hHTepLE1DnqyN7/ww7WuSyKHM3LANwObz42pCb42/Ty0hvtIXX7/3UeGX9c4+JW
mGQznd3LcBirrLjufln3dB5XwOHofraBZeYw0OpxET1hc2qR1XXFNcLEM7ZOsLPl+twkzxdXuwI2
v4RCb/5W/qkdaWAwh5MBbFzidMgvWPsod2zrgz3QTILnPe4nSc3Cs9RREuh0enICnBjpjORsr/2k
rZOvdhzFmOGooUgXKB9a1tPx38r1aERgQsMyS10Z/jAjf2+Pj2LO5qm8QFjUQ5qYxe4CZRuNWcyI
smR2OMAR0bhzIfzf9UypK8IhdRfpAFM/ezQ/kmu9+vCG3dAC1f2nzBdsmRLf2+Q8RShMbrtDMcLZ
5Bh29hchu8vEiIfDSlVnrv5v6qDL7Jd0BjuT2b9gYLH6TouLzEaH2Fi5Wq9wap26pSiK49b5n1ne
hU3hzwrstaJwhaImOCxvUxssBrlf8ffTIqgLL+UT+/lfMrnNae17GMohKoSRoLpLhhGl0k/8G/0K
/7dNgG7gMN30F+WsQH0UTP4yseIA8ds121HU/y70gT7dZ70DSfSh3rH9m9bTQfTJw7Lt5cQVeELE
+9ZlyYByw7fm3rYmYgyJfn2gObVdEGZSj2YWhZFIiUmRtjdHlfp/ucem0TlSYhXDU1tz1B0WxWFV
QpCBnSSet9Pll1d8P8kA8bqihC8tpUQF/2lfqvD/szI2FtKEIzsiqMb3tFms9CUYnPNX18Nr9QU6
g1zj0eNd1a8uixAWDBbiUr959Iru4lIMK32/e02f7L41zcEzTCWrUwKhwo/4TwrS+Hm0u8cMXHJv
+Tpj/nHuk99tsmwvz3h9x9R+fPsQHQka89kYq27DRmpQwx6fG3aVzNvWmneKe+1MgRi7woubROBe
RsOgDnr3PLu3hGu4NxxaDTNW4oVVwlmuAexCPdX67ftOMpEZgL/EzMZiPYTZBwFw6+Dtunqbslno
cl2ph4jVexv2UaI8XaSFkddkx3wP6sZVu1YMXQw3JXJSKj/vG+zhn9eygZxY0YpDnDsjmCTduHKz
5OeKhoH8xiuZafIU5lii5CiD8XTyN3/e8Gzp9mbbMiPQPqLlAAo1saOr1OksYuisnZLmq3djw2SF
RhyXt5+6AZZUR6E1JwDpgAeoUj0qOwrJxqqoiW9prdXH61wcvF0EGyqNEAWIAifnmIpG3AMSJO+T
XGx9fZs+6NzRNdPV+Qax/WHleYFuXNfcGNzhb7nxXRWQKK/EsWYlrBRq/DL71CxHr/Ap5rUORXh/
Rp+VvifajOQ20TQLU4JjfgSSPYnmA3TzXaT9/2R90gwimAutu+p3tF2Z0fRLnmrTGBS4XCZxbDeI
jF8TeDwAKtiZIf2zr7UbNrGP/EZIweUPyJ3SrwraXWyl+aPQCjw2GLpLEOjGShVt1inlgDmQQORH
qc1gzcgDjerrrZpabisVpJW1J0OXVz8aahY6d48w2fumZtJrxIEVOFZZGsTaGesdeaXtQiKRDAok
gEW317ZtxjbFRyXY9Yrl65IfB10Gk8PDmw2J2WgY+fq40hIXLj3+Gm2jnsATvIEgazQYxdr+V9cq
idwVxiqj5ScCr/KwVKr3XMxvxnzfY4uCm0DSLUR6P7PE+w33I4rs7Bsj6TZ9UhIav6OzzdgDgANA
B+6edgOx1iubZXVjC4iL5NsCCcizVFQDrLka1Q+axFnA5LP/Yfu2ihPbmkCqTbKv6L4n51UiePIu
CVeKyIgLhAfSJo5Q/CD4sYWlO8yve+NvE5j/CXRj/C9WFKICZmOswQF7msqTlEhW+vs2ZMb5+OMN
2b7K1cwjwJszVsH9UmJS+fWAtKCFo0okEz+SL5NoFq7v1xpdLFHEYTRgrhQvSJKnPBVCCyK9shtK
dWmLLBYLJSOdW5mpIWOASgT3kFOcf1jCWt1EHh7hywEaFRuesCpufkYfCcyZs9CEzvaYdAvzeMfl
0xKW/9XNm+iWBvV4DL9Trv3HSTylNVSsWatfE8WsrQinFVJJ0BQNhKlKTJXCIfUHThvBloPHpvtI
tAL+acD8PkFbk6Q48BCYP9GJv8QYFYQYGYS4t2sFdAg755ej0desK2MyyYBu145p+BbJ7MH+yoe7
Ec2eatuJ8ZwRIb+qKyMVz9RYdgf1+mCzFCkos6FvyTVmwmElw3wvWAdCtFewFVX3cABQwE7LgAFx
GdQvaYiVvAirTnMhcoztycg2PxP+S+f8yGEvRQaV3S91QHNQJnyu0tTeBh8rJclmAi2ZqHQAdK1m
UzIAycvboZFnHB9gNZ8ggGkigSYAlLIzg+EZ23zJAeC4wB6fvOjp7CW9jNnhe75fXDRO8yAra0vg
HlTNpL36lldhHIgEbANRaRJGUz+1z7JiI5iCortlEzxfT58PkM186eNbvU5X+ScvMB0T+jy6dOxF
OtsshMoWEs/r2fKMuNCW+pO6iZtdqVevHGxajZh3h/f88SfRr3o3OCeRrmYnmNhjNRe87v+N+w80
8fYiVyHoRo+yr2zPhaqSFkLcLZ/MMw3EdCot6xDN+vrvquWUSkHjcZBlij6CKGkuYrAUi7suSYjB
RcxrZphOjyc2oICF3UI0DFtAHChz7juwOIoD6jNyoTzIC4FdcT3eBe9kNNzNzz0t2HB+WP15JzJB
zmMiGQo0js0NtYhR/Mav6BiGnxRpII2/8CG6AjmG6UEngwWR0GHjulhJ8A9nBPEpmK9uniQl1mtb
chfVkzYt1Q8wp2W2uO+1Y4goji5UbDB+fRe73RnpSyYy5SLdsuizCOgWPtM8uB8ISaPfYQ/CG2nk
P0I0Exvkz3TcAHkuZUScIb/bRHMYRmsUOcGarUxZb1WCifc2fIjIV10FhLMqgX0iFVjfseF+fh9k
kd6NpuWa9FI6/2av2DrdFktF0gFkjpKqhzdmegr/bNK6qgu2URo1FTHL30yIE693zFvIX0sLIKUP
9T5xCBBEnx2FrwwyMFo/FLVg82liNu2HZQjWIy9c2mO/DIec+r6a+vBtm6hY8FCh9Lu7zeALpHfq
slMgsShd/RgnMnjBzhdWOQHgSU7Go8lu8zQhDJPVIKcYOXa+e1a+ovR2kRKbgoUryg4zaESlhDaV
JXUl3Gj3VGFPQkFrtGhQSy/X/l2ggHLjbnJZzVADYK6vB38qHJC4jdNm6VyGdMjsES5dwGKncmm3
jkrwcSd4RO3Fr6cU4yWbV4kWSHDSLgkLwkSBtI0ArEUPUNxXkcvflsyVxDxCEXrhFEo/wpM+aNiZ
HD1wLh7R8Nc7jvzxcUg2VPgCF2L3tYJNTMOPlUYGhGRbELKtcbM+Gwxs33TlfwxX4/a9rhPd+gun
ehitBGrY1y0prnIOPXUnf65XZh//WtTcR8Kdpd+5GMifCsRo+Y/Q6SwJPhajs1N0qQBQYGGRMwk/
smr/2zGKltV/ylKPSuzDJgBS4/6JsNlyUucvaBEs0LI8+8J/wl5PquwOLnJtnuuMTLHJqZ2zn1WB
QTqx1eQhTcLDwkJXkCigCZHWK0yIS1U8cFaL6RG/koIvaPS5MjRO64OYyxe4jnc3awa3WpaDoHnv
wrAmPV6xoARL83Fo26/j1sLbyuApmt1BCp97zxy+9reurzSuTO1Yj/vPhdpIatK99lqZZnN9u7Uv
Bt28/r6k520fK51scBnSUvqh2Kmckd4E7hZ/E/WmaO92uu2oaoXJAkYuA0cVWEIMmpDR24mzXJ5R
3K7SaW7/ZNnd1Fth+PkyBWLsEtczWdiMEc4Fg1wlDtevMFxVWO9Wp36HUhbKYmGxzLREpNDrHW6/
DLsXCylVxSYbtkHNXb2k6vzuivExv9tVGLxYxMr4uHa163RuCGorI6KHGmkvuOexrWo4kK8xFYrW
VN/U9pXRtZREcqVMOGB5JRyNi72VRw/BDwS9jEDsBlTAhY7pS8GxP8yjrkfGKjcja3p0d+zKwIPf
R/9NTt3MeGd1a0+Qeyh/8F5E0qsnUIrGnGimb0s+F0PCTjcdzTYrjNtZ4cuDRPpaETXd5KgA+CTN
HAg68bM0AhQwQWgjOWK2GBBuonOZLK+VB+Z6JQKpJX1fXxht/Fub+DEA2TUFso/t8C6jv2DC+iZm
0wJvmQm0rj0lAYrHPQ1O5F4Xer2ejleHmerR3BCZ5iOduJXx1GT53qzZFoNCUz8vHi0rIHt01gCC
WBME8nDZ8gskeGUlnPuSRy3ZwcyFf4qsPqMasMce1mTM+thnKkwOddAPvR7UCKRQV/E36cni4DW+
8U2Ba0y/MqrTjQSOaZobh2NUrfn1BZyWh1NeLB9IYt0hYJNwpUAGbj9JnBhdh3ipMh1uVQ/SukKo
ux/uelt9d95+SnXSg/WrN7o+IRGIkLzb2gAg35YPtokpSkLwRD7+y/cdo+kyvAEXWRHjrrxQ6J8f
kFp3Mk4E7rG+nMpMQKdZJK9FejsPco5Be2bpICILCtvAdZzfXi0y6YA2J/wvzj+k/hEexrPSkADI
SNJWqi6rDOh2b4XYRbPAe+wWI65mdV9r04BvscjYPbd80eI3C4KL3JxjjzNe9gbxYEAqtOJohV/Q
0VfriicTWQMglMnZYhEMmfrz46RZ8XI5RCN16NxtSb56HGrcJR2duyFsuOP63RQ4UgfIiJtheDCm
kZTtlXTXv/LWgdETxyIg6xdNuryCQRz+8E2qfsUAO3Gpr36UMWiq4uAf7lDqlhGotsba4ZI5Ixew
YaOjMb9SlCe6NQ6lQj6cozlxCE+1+aSjhGGmKiR7SzGjHsXXfUqXg8DVeQvJZEOE1wIEFePbgqfB
l/sitpf1kRU3KAopwzyZzWF8On4v47biN2tl2s0mAAUzYAymlAGM1GiTCKflVJ96cUOdDNccSHuv
l443zlrSP2MKsuP7LmQPDfu/vAvmodeiLC+XgGcImiKV/XLylFq4n5bMR9PVuAydOtqdAOwY23LQ
zlIUlcPoTr/NDFXepriu5+qChDp7WgMd+8PBSJ4EilYZHSuC3jjPgudo/cZ6cbTSBbJL77fDxEBb
znaF4U81XG3D1J1eT2vSTF+pIGrWiF5jW4UQjcFOh32HYdpB4+fU7AX/oan8LvUF75MfZ9AAqYew
TLcVmPjNrtCGwdvsLFU8RCsU9B0P/Q5F7rCqy1mFgeJ53SXqVkxjK2rhqcN3diwMSZqVSJt6fOSx
B1GyGSR3jQTMh+nRfrS93phx2O7LEP3cholyoHTyV43u9WMvBE4pHIl0l8OYSgHOdFVVZj2hJzdt
6cU+Wa45goIfxK0OsLYU91VQkO60/L5bJR9kogoYXom+SVvj2lW4/igiV7W+H59JDqKoZEXc/mZd
EFfml8BjqgtFxzVDi/CS+T7Fn/Vt4ORP3iSx64+BgokAbquOsQ5kWdxFu6GH7Cvs3lqAKtTct1r6
QxxddGd40fgYBW9//s2vD5D9X6y2BG0BAPhUS7gnC1GO2y0Ek9Av67uag9//4CtoFts5clVRG9De
+wkJfQ3bP0hHp398ai2f/F6enmTavqHpewkSLhyB0VYQJ+fQQePDjbeJvl2mVbwxmrlUPg21VyYd
ylgQHKth87BUaU2OghuucjgjWTbk8y3RKzLNel497LXG7Rv04IL0Kfm8RqyACmbg+Afx/+SiK9JS
dPmcFxitNTDkciHkCnepcIfvOBJKcemzu2mqG8jHBuuirf+KWC4HpnqrYUDtfEupr6CPTtKbiApd
9TLv8uZTXjXtqSINbVzoZ1nOHZHRrbjoc6owW3E44LAG90SIvAthnj4wsRn2T/1PYxB1h2LAN9eO
ea7UqgxGidkqDAiiNhyWzu1U0xd25s1F9O7S0B0e5nvOuYvTnceQHgj535upKniNgumEZhERINQF
XQGShtVI6suQJJ/T0X5XNRMalNjWw9fp2VaFMaKDtxrmGVeL2g9jn2RWssSrk7m9K8QMFK4+nffq
Sv9Y9JTw44Y0Q7y2vE3NAmn1De14LBVVO3GmRvsUanbwqdR5J9Dyn8ydJSK8CgB4hYHHjnKzmtbF
EZEOheVuev5RKgh4HhAZIBXD2bPitC61EBiw2zx//36IcHU88ARa61c+F67cRlzqVuUCelnPHEzk
YkeTxpHuryCpBtF3BiIwpx892zRE8FycWOwZU+J8COMUFvXfq043rafw+JIHxmsPrXe5/9ROpatj
37yR017QcZRuSTvH7Dt+c8vf7pnTuOwwQ4VVe91YEm/zpjDoRSSSUmK1GBXwjgFuquJ6n1eXDGyd
FX4Ii8jmVjL9uSNupQo2nMEgArhFCQumNTWz5BGuiLyrp7XcojZvrt7FZZVQ/Z9QjMpyDsHPeH49
C1aAQhv9OrfvmImxhjMD030ueqOAJJlDNWomh/du57fE55UmSqfUxfrLAFhLYYMiUOVEEfKcICAD
nU+YchqFn2dDTWdKwNLLnvhGjvWoNOXkXK2dJjE0fjnKUG29fFALIJlYpj1evvVowwHxDEPfCvpR
vbaxY74P0TKTSEt3/2lXv12JZZKalMYI0IVyZkg+Kqdg3KPgRzECl5uXxGiO4iKa4YRs7Zr+ZjYv
3EXtMBpDC5IcXHE5iOuqvKE3rRCVMupKpP3ZkKKwJ4jo6q4opIVVkciNb3QAb+1wBr9PKbmNyexC
rzYK7xBSiwlE3a/6r6L5udcmrgfTuGZ0j3Ws2WwNkL+M/88oJ/RL3jHN5RX/zaCD/D9zDGqa439l
r0ROWcavF9IV/g6xideFPpbDqczURUll43Wb5Nfz9Ql76xzqK9spaDZWYdvib3J7N26ksHIarehZ
7POJLb0YaHQczjPgv4/fcAqn35Ghwstk/uaR0gPpb5hgy9I97tYFUBT6vXx+gkFMh93yeOG5mZqO
nUl4H7D1PFPmz1dL9YvmETmUUqtyff1/ZcHJogQ79zxIqfPhRGs6dMjz1cug62x3+5B95dc1F4VE
oDGELrgWV5gGt1ZX3ZIsCUfIfPbtW067a35yGoNunp95oI75vpn9USaAZz9QDlidX0ajZJUXC31E
KoYEOjDPwg1gSbIYqnfmpzAA0bG5dpMN8Xk5RmvoIFniDkQHtKk4WSXDawp4iRH6dffyY53d8OV2
QGTAJ6oaOLB02RSzsBjwnYf3V16HOm5KpkTKstjbLAOYW3HVy7G9NZw+n/aG8th4bFJ/bXGgtoA2
EbFQv4Cs9GNtA8wNUTo+imJx9/Ry6qcQgw4XLCbH6xEwZ9wINxQfUiiqv3NuUn272jdg9iawVyOP
6ivFPWXfM/BQPkXZJXKQekgC8xsSYU3mCKOvA80Llj7qgmMo/lK5m2k8Z8STe2wCiyIWIWKgTDxr
qhgShRWvqyUNtj/4Jakyc+I/u041J2ieigiq17yEZ/Wv7A3UAZJCCfRVG+J6fzFR4SQxM5cSub8m
yOcX8FdTo5MM4ZQ37UTffN8YqBsXNfB+nIDynkdiUO2erlUO6SEzYOpWKQgedDJclQHjL1qpFqEZ
mPPBfgrl0nCq3l0fTKkk5Ow9uPMOgo96akdsYNoAb2rFHEXqeqV2QcUTXHIUleJsD89sQFNN5oiu
hC6B/JgxP9ozcTETBELx/olgtf6qqG1ZIGDNTT7TGpHxwvybqGf4aDhwGGrkUoBYCzfgvPI7exil
T/Rv98uefX06TfMFvSSikCDYGjgVfEHZa1ZVXYr2J7QPJyI81cuUxxOfnqRDizRmVTTK78J3ajRs
aIdaVT++yXv/Hs766xYJPGyHikCeVUgKsns0aL6w+nB6ermfdEYRG7+UmFHFe+SoX4D4cktXHkuf
NcrADKjPmEvzhTd3pAMPPM59D1UGPu+SUncFkTEMpAZqsVdVrm6OVXVAVszbK7iAEI3x6BoQ2Xra
nbIfTaejhP5v7fXGuvTn4dJJFKyZANXVsX3VmyHugB2RwKo01R/9LsnRl3/awDKm+734P8Mxs6gv
6rj4IKVx1/NKDK6BB4JJENRwKiqOJTbhEFS4zjpnhYFb1PJOzqIz+z9Drfc6dGeeAqP829NB96dY
Twj2Fgwi/2cHO092VgQ31v7Ar/VpTYYE2nh5/Uip7OcG6iVdZwt1MM20PCv4erNqWzqw31OWEsq5
t3o2fnJ5IlV5p1j8bneILanfprkg12NfopiSvc8OPZEm3mtFaNbBKBceNHz79VhqWjf71XmtK8gp
jPOQ/qX7U+d6NScqWYPkA4qwS2zXkh5iUYH0zzEr7DncvWRL+lwMg/Pe1DnTZ7zW4X259IA/Bpkt
EauLv2+IoillfUul+yfFoIYcSODKB5NrrO9iMkNgjhBvIv5+yA2Q3aEp3pPDxhw+bfqYiAaEgs22
OAaopzc0qG2s/3Od3gtX/0P+TEkKFmi7iJxLVjK6yIXbA/2mANDCtpbzGyVPVqpp6OU06gBzR1Hf
+YZ+XCISXsj8hti+ect/dyA3A8HV4HFu2G/P5jHVYBcJWexGv9lvAR0EMOqbTkvwTrFXZHbx3z+O
ID/XaNebhuFPGm+LD7mzjSlLrvr5ifluOWpq6mqw50rsrREw9H6F35whqGBkJH1xQAGuqOUXatuX
3eCYajvuMkVc6zT6HA4q5Rq2orDnWLP9CL7RMHTRM1lIIZ420zjtOHajKysoZbK7KzlceLLvyn3C
ZKoQ2LmcszPjo4ktWy0boMqzZvoCwPHSj/q7I5R4+S7bDwwX3N3I3Byifjs1hkZqk4wKw/WHn2iI
WumQmkcaR6Bbf2O0W2U1jvDRki1QL8sCdyYKfm+14IbAabxBIDrRoZdMDzOWZug+R+QtD0rK0vwT
uY6wM00cIRSi0vgZkAN+vod+CBzKDFfr2YJsP8Yr+kFOScOsB+zJu8A2PxYw4Pcb4mry/cotLnZO
AJBlDY8m2i34axpu5Jcg5VdjOW9Hf0AoaD00OHul+QpUZG5T/TU7rZwxtHFe9BEHrxRf4L4TKDAi
zSjd/SJXPXBOj7vdWKT9SFpNLl/hmTmarzjN4BC1QfKKIb3MqAsdnTz4pxHE41G2GLDFYl9+6TQx
natNXXUmaY8OUTbLiDRiIxsm+KweYpXCwg+S+RNAWrj+RcKeYk6+aP2RA469RH3xG3Nb70fAb3uX
hJ4PHS5hp1ptTbLo3+FKaSUaiZ8Qxn6h8mCpy9aToxakDZ6sdCL3m2h9Y9v0uo2YWY5QHQQPQrS3
kQNMI1VPV3hiPUmzWNB+zNc/yEwkgeVx8q11X+DKy2DbqeLl7AN59Q5uz0eRQnG7Mo41CaFHz3Xc
L1y6kyht35sJXmmdInuLoj7REJLJlKG7EblX5/i6FQPduVq4MzQzlyXZelF91Up8oYkqLXnkTRy/
mtSPbcQFnVbuP3/EGmjVqd5sbeMZL2ILOatm3PDi+LmuTO+nGKiB502+t+mXI9gC4Sql2j+ucUZX
lOeVN8BqtTbQRwAGMFg1z85HeXdtcv/s6k4RY+oRukfh62+oF38Rk7Bzc7vRAMfcnGZiWmGPfcw4
L2vjX0NSOOQz7e8CitPaYM+z6lQ6tSnFkOuqMmEFcWGU4uqc4sD2YC/wCLZWKAsHl1+79WFUO6n2
vI1bTqUoYWsb57D9HI04GcpOqX1ATbc40xqYqY6sqzeUYwVC/8cvbRqoFpXmxnUCpMRPFQc6Oo5s
loc01fVpfkB/NOmeAoxR0qfFKgDT2TqbFOHQsLrOTi1KZz9QfQAYM/JrGlhHGF1FO9LAGAOMaIG9
BRMM+uLhWMQZwE9uCuHDe2yCrvq5stofJFm1YccrFIYVIgBq4JaDFdTOXucbcYiOcv6zq/+uUJqh
DAs9F94HcC97InMQOBP2iaUj1SoAcKsDYR99YlMvaZEXZH4R5cTfmPxE/iPoICvPOlx0NTOa1vQB
fEoVE6ZZyWFUpDtVIGWSmJoNxhpZdi7ofMy6hBwoKdJxe65NYVlWZEd4ogn0KEOIa3vUaTVGPAP7
2TyoJtxfuaHTtkXTfmvH2jfpnwg5OFlqrFUE9VYke6CCysKdNqLTl+vEMUO3DHZMjVU5O5Xf4X1Q
5NZVQbo+IER+/p1wpZFX5Emb8BXqWTYGOG+m8+18I+qyMelfd0FSJQ3tV5Mpyj5/csmlLITajWJ4
v448RuY/ybseLrV/6K5V/c1OiqfHWDRumnJJzZEwyAPPVwGXMU522WtF0C3DBD/y1nb92MKgsMwK
weIXv8zDefP6+od/NpwUkS6kO0iYeKrc+sB41KfJcyQtFvA06DcOGd3cJeHjS81LgJ9W7phPmNQ8
gbJT99MEvrmkAxtF4d4HtbSaURno/ebd4DHgPdPYHapfl5On4INeZjz41SGjSAIzSB5KzDdY396R
RgW8O75QuFibfTRETBwU1mnyOT1/KvebDg3ph+9KXSpRuSoqxmQNPI479ybVpa0+auAQKSdeaHj4
kuVDAGMQJPqdW2NztJ37kfz0pAMYkxwKsjxZIUY839KIw4+9XSKgrr75gBYfk3KcS9rhRswI0tVl
sEp67CttKTIUAWpqWr6yo1elkUnZUr+sYMf+MqwmvQPCpvyxoivFug7ildzyrbQE/C+E3DI6nkY+
cq8CRJiMy4i6D1Epl1SYIKTcs5wzVstPeO8g2qkwAv1Qi1TdZ8LfpoXeUrIKuWnkr6yeJ0Ml9gRG
CZMchjtVLzCOC+EfaLMPJ0QU/tdFUp7M9yXG0JRxlXXxu8OtT+Qn62WeNhY6lX0zLN3xpa/rGpY9
iBEoV2mnFndnERwK3UzKgTwrrzOD7BFRuTfDx18w7lKHTX3alpPIOqwa49kGkmf8zb+hUN8wRHxP
0SNroxbzw3PRBjD8ysqqx0TY2438xL+wSK+qYDtwyvk2Kb7zImPEQpEoMiblfIrT01zVMxPYYP3s
BZElKHxQiNecC8Ze/g1H1W9XSxrc5OM6wLxZ+XvbovUqciwCOAd7ugkkMHWalKub/kojV8KxPive
reA4G9BMxgsfKfB1ED3hQaeso0HjorIKXy56HkHSsaZDSAD5rGKdrk4GxWgcf/QVN803Pwh/eONl
Co3WKp13POmMz3JFQAS3lUUlqGnXeCHen0OPjlq7AyCVfih+Ntfedp6NVO/9SLNBBA/IGmEN8qEF
k/xwN1L+gSsFNCk1DBR7ObdwDyQRIs70/tIPXK44fhNkLDZ2xlbOR06Jg23YiZJJshnlwXjzAxLm
tCKiAL9uXSNyEjKmiXdBgPMtu5nlfVmqfb6hLjxE2j6XpFFFfsMnBceOwIenSAQV5Ktr8AcueuK6
mMvHK8GQ/zK84ig7UB3p3iyxNPTjnIym/zOAm5L/uM7g30FgDb9REgq1g6p8qtw+KqzWwWVabM/p
Ras4lTCpOnQfeAmW6fX5TdF/pup1HrBVmzJOVRYaF2iIbVV1EUf25oHWEsF/BYPdDhN3Zy3HOQVj
E45Fa9ep85yFymdXMdanXFtvkCDqtTPmSOfBDmg9CuCXpMRAYSrEj+ksxGk16iQhjcKOh4cP9Ujs
8dLfV77/IruwupjblKa7lzoZWU9c/qMxeuVeKITHnF9UvI7fqMZsHDuTGfjjKPKIbMZ5X/FrfXQL
PBo21E3lOw/EiDd23RwLBB78JRQvg249SiVMLyZpRCerWzsIcOPSZXmzuXFKVTAJhybcb2a11Cgv
WXOFM08mTojM48b3Xjyp0iQ+/R4FhlBt2piUfkxLXLpdmyUBJ4VmbF+LQ+xAhIsIsZDluiq2irDL
c5Ndar3byha23ztROFXxvthYEkg6ND1zofvCPxvTuW4SM/Mu9PxtV5bCrX1b8/OXksTfAbog6z6U
wlg8NaF+oLECOVLRdFwUhgRflZ1CMwc3M6xFOZxKOMHDLYA/IWpBt/flKSaauXQMx9S/38+FiVq2
4/HhOuFFtHzcbMSb9WoCyYqW5vCDbPvE1mrKX03rOgtgxwreqFRYAyPDV7trOkMpS7nLBdik53V7
fFiRkMt8p3GgtJ3oUrs1lO2Xn+U+fdRLgAXHRZZga2lKD7xHKb8vHRc6XUoJe/kCocG9nydQ+tZS
4DfEeWKAnfoj+Fa7fqNRxCtiq9+p3mDm8MwDnLFH9DlPcvZv0nnqtc9uC8KOVV3/xiGeedXPOaoX
LI7HpF8rg8XSdsLJiVShQn3YjCTge/cCu0DRiG4DfuuAbE29gcsCsPhcXn5y2zTZwYq0lKVHX6ec
aC3U/PhHQc+R3U+onJ5ZgpRbqEbUR0nkAAvPddSmjiaO2sUx1fQql0tKHYbcKh7Di2uGL3C6FJuo
pSdQJs03Itbbvw2kQLkVo/cjUpjJ4Uo4/qpT8frw3aG5EyOmYHV022NkL02IBZJbdsq4WCxwF5YC
TCorciD4cKIfxThOjrZOLIgPFy0Y6umSCxo6YmATC95c6d9Bj2uAw3MhF8N4KFbr7sG/eK5gtsYC
j1JcSuLnTJwinyZUR+YjhLexTQr0S8Dci3fImeiI+mfx2BcPPfu4cA8jw5qSpldrknWbfmGUil7n
kLV9wLyqDsCc/7/LWFFbzo8rj4pWO7AkK+tIRsYJY2mjOtWm7hPtd7G/ZT4zF4Z8D+Fx1wnAQbBF
X2ouU4pnMzGJKro9yMdHE5NUitpstO6UoPhczHux43gS3IRuZTOyTtgyU65ckrxPC1N7oMZcJ/vT
JtALPHdIpKKKKWYYnhYzEe8pwYfaFYg+N/rzAdvu0psZ7e1W0Y+l6RFg0C3wzAggcOxrZ2tBXULu
3rTO/3V6UK43e/zfig3+ivYQa/InY+Kq77negrFJgbHxGteuMapIqcOVlUsdQJXfLXn7FTBdB2HB
Yb6AzItunbclCqmPsIG+gs6tJXxO4pPLZXbZJUncHQMYxV/suGTTebxUQXFcQpDk7kofQuuxLwe3
N1gJj/TeSQo2LlGRzqKgRdwq9ZnzpcOAsjATB7N/rntw6jFa839qjpjtgEcLtegCtBf8AmSbJvE/
Zj52E1K3vV/RyAoW9ZHIz0z/++EOxnrxRkekDJzEkg5RLXGoiUZF4XyuwmEhy4FsvxpggP0f/bzL
2N6XdLh3DHGQpaKXd796HIHguMi6rO8YYXZ9Q+ZCE7H9RiS5mNfK0wzNUzupVfaah1/Yj1aQ2tU0
jQjKrZV7Q1ByVEOERpHOulFl6aV/mN1AK5aBajwxAwActgQtvv7FqjCWpTamvPu1ZhsbwD6IrW5G
+upA7aqfjLB7q7YflSN4CujpPXs+8hNGmMf6xFNH6pJQjzm5JN+FoQLbUtDXshXXM5jMFaWr5PSD
EMOa6/XXGS3V7hfq/GhOBjsVl/9MNY/AAviiEPSsKDzH+kf8kDCqcNi4WM1RX353HoBunxRszVkv
2dtR/P8lEbop9Hrdc6OefRKBuWSi7oV4rIEmk/P/VyUseoCV6Vt68H9uKYbyawCl/h/5SKJG5Vhk
ZSJh8DlUmnRq5YGuC8kfobCb32u1K8ujlQy5i+oC1qVnZA7nU0sSSLfGpVzPPfuShe0HIM55OKAm
RLdQBhIuglnVvx/kq/8ZdHDEbQ6MFKqbwl/m8QIhloUeTi/7c4YSK6mezvcm+j9gtwdYI7V+3++7
N8rITRFCI/EkYiUXTEy1/MgG/RGJbQOUpoggDBio2Dd3I7pk7HCNIDS3uNO9Yo9/lnlAsNOhehJZ
NkONPTrjtwZfb4wbkaXyUcVsdgJEj3lTrVZ6LVkA2GTpI5bXkTHWYwieEAqhJBh2gP4BeFGLDM7O
MbBbN7dwExbwZgwfijy+dVKyYCT1jG0nbgPkq/puEkjaBwBcgNoSg6VdgxKZMmXZ/LV7KUWPWxQB
unijtQHEpRbozsJEjflQ1PUh8avyGFdrdQra2KlB8NQmfC4OGjUmskLjGQLhpKemJ5j0m61nxnxA
IyZzWzB8xR9UfDXbESFF/3aeepyqu1IhdHRYwId7FwEIwsQIXTa9xkUizB7KknpMs1G7qnov03U/
KC9t48cRIckuJ7IC5JwQM4E2Kb1Zvi5x3xJrA5hduvDV4oEv1l61kv5NscYhQZHgkqP8WAqF/wh7
XAqxze7X/Dp2BrQnr6VK8Yb/bbWTkoi6MK4ILnkMkK2gYnil79AKWhn1uselqwuuS2kquRU59p4G
hI2BIcllDEerGl+RV7RgdW8jgox1KklBOEu/jd7tt8yR2cobjihh72A6nZ/ff8psDT1T2kpOBcSc
STxUJ/e3eb4V4Xd6yVw+4i86NGE0okx/7Aagc1FvZnkUhVWVUF3F5A8T2Bus6M1tUcJ2sT7/zAxU
GNhRKWr+iOgjRuo+NM0+Lbo78INBXTmqRWV4m5g9CxSHAcPyMcJBUDZAsc9O8G7GhiNJWjDUEIKw
nVrgM14MvMPlivU5LnYdR6azQiXzTnduSaa5JFkSvRyTY9QiaTI7a8lpQ4gyMcQwyXJ8bDtoQmY5
pLXgOgly1hsj1Vz1e1pb41wEofwdoFhUs03I/GSljkAGs1gPEnE82nxZG6OcrVGptBLOPQc149/c
DiTjvvWRwqYEUIkHunxi7Nkhm/gzLQLObqFBPo+QzsKQSn3cO21xVeBXSWAuSBFCZvD9316rxNgC
FvUx7S5ufPHS7CZ9f8+e0NVhoUl2nCtFWRlPBQlD/GLk73lNKVtYAqGMOO5lvXEZgUf51AzadOnB
w+/9p8F957ejEHXYUGCcEKQt0mexro2TY385na6steN8b7pN8Vmly1vQxmRYJgWcZw0uRxZJhGqr
57BtGbeAitviHqlnuxzggNARgQ/nT4lsxFY0fOsLh8ps65nSknUl22USo4/EzbbCSH4TxZD4DhC5
gW5T7xvLRY93FOEq9yFUg6QTExQ5R3Gsp6Tmbg4WoVXc4wNcKoNzO6X+Elf+L8x+xXtQ0ZqUMUTh
EWsiqD+YHPs4V1OzVafXypr8oAOKRRR0M+0ExDbUDwg8XIWzMhHHTYCcPv8u3RIplFyczGgEbPrz
Zfk8kCUa3ft8P8D9FfMrgag7JNASl1CnSOk/13pijGK09h3fs9YypQfhwPfSa2P4a/+7eof48qgU
ut2qtpvfQmnmiVBfz/dovejaADRX56uiNPRFS6639AzrXWDwSZVc4rKHOJioFwyJNO57PfFe3sQQ
9WxFvOh3prydoT1IK0pyadU4Kukfwrevm/JQyZkAC7MlHtQrLDTKS4Skh5z8lV4r4RW3G7zVc436
IQFT/RkoGzr2EDp1R1gz7k+mlV9wfSxjTZj8rukhrxlTTB4nXQll7JNa9vjZ2Y2a/9HnDNuvT8is
tK4HosKID/U/r3Rbgi8VMN9YxQHO83bFbn+YPkIuTqyR89Scppy8x2iHyUU/xJL6rkkUK2/2Eflw
QvldBqf65b/xv67c9DQZ2efqAqVbGj2Iwq4NRvX1VG/uO2Vv5K37BOoDXUrm+fdRYl/NjqMGCmWW
JwmmwD1rsRcJs2acEY3q3My2SZIRiysblK6nnH//PgeTtw0g54wAM7EFnLaoTcjXBOcTRF8+g/+1
R4rjmvDZ9aX5Fo3hyQInhPlo6bffOHmngfyzHvRqca9tj20xnQbuOOvUmdYvhrw+EVSoyPPHRH27
ZTYERBrTWjNHo4lfbIErTgVF5GDmat2zVQr+ENN9xil+e5nXJSoaIk8rttqMeEW+X8wRyoPbgefr
u26iOOZaYqIJ/7iWc5GSDh8DNamP7PN5Ff2+S59HMWG/zDklKHroKDy1OCjwDHu2oLWfHMw9cld3
6i6sIBm1ni5lS+R5b0aPGBjpVQqOA9g5jiiygkP7SdAIhSO6Ze9QWgK7JhOglBjKsDDopk8g3amV
giw1Ml6129X0LNd8gs442JnJvQ/jCgiSaOOwH8hLzcRGpO5Vqnxt00avuNsHfqH/MrkZBHSmq1uo
gKhh5h0jJ0vQop6CCWkDRej+iafx/iyB6JAajVXc/x9rSIoUZAtQsjdlHXwmSlx9X4mDphV5qgi0
ObPOij3BAZxrJ9zE0wE8RuO/2GNucqkJ1jazVfTAjDxEJDjgeUfRyndh0GrscUAX8TPbIV47lX9r
62flu3ezO8AfVvPW3j+q4P3G+k4S6Tf/KJrCjCIHTcI0Z+mUH5Yu8wZ4QCxlhUDM7EdIugV27WUi
EFJED7xjxxBllBu54bHXdD4OfVx1nH3smLMQsmHcheH/OtD8qsJBMq+Zz9NMSc1b4ehO0fVSZo2q
JxqXZpNL9GTuC2L+K0swCBe91FQ28bGyRa7sGNtf3go8J0H9IZz5yh69GjItYDmVFFbKxGZsW5lj
qr9gg+IsfJLj92qGjqjL/YJUb3/HYZhV/Pqy53C8G54UIjp5Tuo8ZyIYBhz1P8kbY4mC1Qh5IL74
GBk1hiYKVomzwynCWDAz3f7ALa8bzJu89uzZ7P4kxASrwfQGyYzF0I+BSuVydNgQ+XdhAZghfMEP
Gt+jCG7seeyEosqmVOfsMcXFdW0n73JAS6BjihReKoIAoxkRli+/TTkrczGLk3yL/hMrP4NXLGFq
3QwycaugwnQ3gqLJJmk1FJhrqe/6A3/A+xU8uJQY35rcBfLyySlhKITwZ/F8igQ0vt78dblxcSYj
bQKp3AsD48VQbbXbULen0SQqSzcWIT3Sk0HuDkra9g765cthgqVdBJRZofROtVtyzCxIZpIOzn9f
AUx+sP7gMAL0fKjX9davxddpxYfry5y8pDxsuTxHJuqL/3dXt+EWIGWD+lMGeAvj9wp7AizSYAeT
LVO2B3HwBVKKl48c1FBN/MrqQUoSMONdbYeGxM9pqxd5oUOo6h4dGFdZ4+RqDDFpD9YjvUfHWWlL
8UqHVNQzbn0ADCGWtUUP6ysggafYtrNWkqckZsNSzaK4K3+6uMUNwz3e3EFVd9lySpwN1OFrK4Bb
FOkkSVFuKyL9rnQkfKqUJpoRqpn1G1ONJOR62B8gktSva9SKloSFJmmAvbwZbHpMP04BlDeV9a7g
xFvKFU4GAbN//+5m8jm9q21z5rcFoVeUvM/L5fWutb8mdIokbD6Qn5rDwrfJygTu+krPyEtVRr3q
5NJx3vxE/QpVn12wUZ1mDeB0Q3YyDxi/HkYbtRNSG9UvAPtLuwwhAWlYahCdtyJkNmwetv0Mt88Y
TudfiRD83LDXemT1TNkAQ4cOTOpolvYIx9N7RXUlJ4eO8aZHhlAfbWDLzA+Fp/untX567cpLISgV
e3M5aav6Ji5Q2byLH7A27ls+JdteTptiumRiWk32ACUcyJz/8A0NyZjcstoBYmC7c7Ux7uS+yM4H
DtE/c+gzn2u0FYSfpF4DBDepKM4xymgD65ymnWd3DAjym4aJ7qSfxShqGnUl6DB9gUSMagca1Fvj
r/5dyx2+wlq46hZeQWZuULrsDGvNp3vnTXxa/gN0llDcVE8XDX3AC4qOYPkl8P+d293jwXhJyJr0
ApACozWXdDw5WVTzxik646cEHLnEmFaErU5IFGTSC8XxdbjLvQR8ymoqsFlnaUkFgb1xn8QlrtFv
COLyaMDF0h9w65ghZLxCjkusTJkII7/c9UNh7sb1+fCjbRIFfNA4J3dkJf5S1ipjErtIfLv4JTwF
EoQ/dQyDIH1vQVoxYRuXo8pUA125Z96BL3yrQ4fT5b3Fa0uPQUhCHps0eik+0S4Co+Ucr0Uol/IK
3tgZ6smOmEKnuCS14ZXCdVB1f3qfDHi/ktJEg+vn8JPI3vOOKFkv2JVo3zqn8OgVcxOPy84vVMyC
kOk2SOUBvyL5CxWjEuy068rlkhVnzXpDWAsuxNZrFqapo/Vbue8BJa3vg2Yp7Wo0QW2wJY2RWb5U
aOAYEVTDwLc9GGOoVF8UZfwWdZ0lMw9VfaERMjCrdWVSoagUMU+ALqzUJn0Uwf7b2ss//PPgg0s4
mZv5f/8PwS82LyqfRuYACGzVwPj6XlDBiOO3Ab4uuFNpuJuqK7C4WjggxoWt8j9+UREXw5CT8ywI
Gy1yYQYDIXznf/mJghNVMzNQR2CcPr9jKF8dgyU8YzkP3jNFCRL4sx3ap8N0sEKLj0spkPMTL73H
VmdZjyd2bcBmgfxrlMOzcYjGMkV/dQfBoJTbJ9TlJEMG5Jq0bpvCowbrj4FvN66VpfgvfxowBytG
Jg6Qi9E7ypGYwXGY5EekV10TtcQ0+sm4qA2UmkWwNKgNe5D3YTRwcEd07L7/8ruNxhKKzOahLyAw
5qUiHTYh7TMFXbtNvuV6rahvb09PVFXm1RFwTa2JNz5LqzBkg1k9Mpo8ixBpt1ixrj7aZXet2AyW
R9XVZofbuo25EjKMfxQR7G52sDKRx30U+Arcl51m0E9H3jG++Ol837OQFNmAcw6Xr6voUQJ3nMn8
ZKgbdDddbrHYSj9m597HpyZZ6+uLynl5dtr2N2hjbOpvYrBeRWKdJnPE/RNrogPiCC8I2epWCjRt
ZqaKJD2yIsARY7UI66WUBJ3Z860/CiBlCe4OkdammhuMcOJ5kd06MEdpAKKd/po4b6B2bb/d+gKA
pAjiKJqAj3MBXaHbInDe3Iq6tok9n8ciDf923wq5UjzyOY03edRjhqF+skz3ysCAMvgWiikK5RUv
TBiZ//6kJgU8pp0/NVRmaf2Lcj0sVvOM1RLSR3kIonKVCBeWOMxEHh/8U1xzBVZQwvqxOYOFyydE
weKKMmqIMv1UBud39VioJCDyAHL1Qdzm9GrWPPnnGk6k3Qruq4P5o04A2Y6fbrDmHY2tKQzEvEKA
k1Ok7o1hy2/zl5mdZ2NGniXU7gxmRpoOeXO2l4KmpQD8zQeBXMkVCbfz7ZOaJCueL4yPrmWNnU0D
mBnhqeZbwiJggf6Umjvl4r7ZB8rX5f0ttIZCJBHn25U8RihuMOxUCutYqfzn4fOaSOSaa+BWcmEW
tWXMZUdKTaonMH2TIgr4ffXEED8DVSBkSZJ8tmR0lxpp+PKbiSrIlnWQkvItxDC1yqkIE3oKEQC+
ezAw/STQJuuvYFwZKxcB6XQjuK4EYyTwiB7By2szi7dhnElnsPUnjiDYtFlMRe2C9kXxIZ2JFKjG
j0h/zqSroT5aTBpEMA9wSWsghkpwnsR9kJX8y0e3GFB78mRkFopOGKb8uumm6hnSxZ5lKPo0yLs8
47zk3ijp6VtrqsjXaYAf3uvbsvlD680P1haqeW0nKVQJniJEF+0xMWOXf3V0kiLlxCHdVyJ82r+/
iRD92hELe1ydkxMXCKo1boKDSiqUiPXGWaHKwQm1C8aUDF9hUIVsul/37Eck9n+2PtA407YhRqg/
8gbrKsrTgmQPp22X8VFsdoVQX28rYugqcxcPRmcj3rAe15lGkiRKzhUUMXH1iUgMjUE7SLCvjCFr
TeBKPYpYRdmkEyGWC1ONfDNBe0pTBfeyONnsLqBxMmyQYVZ7yIo85gQO0hflQwy33ABTTXRRX7qO
7HDvjsbmuAcZoIRbrRZuTLWZY6Q9DGBOqMRzliGy1NqW9aqOLuW7Zf3iTPhNLalytjtg8A7eTeGa
f4Nx2gUpglt8cIYi/GxLHsYZJOCXepbJMQjzkdcSsheBCXUF/L9YhP5QN+nvcXI5T0ifIriVLn28
k0S7ZcA6pKIkE5uKMrtUNaOV8rz7ob4Sq7RLzTIhaSz65qR2pfByHd4jy259bUyH2+ZG2eqGQ9Hz
2/u+2iPfk7syJzeUClq1ZasTCBzrrY3qG/aK/Z+d2g62P4lU+20CfEKsl7N7qmpWvXjZDczGz6k+
l2NDVYijctn/9BcJ7naRwKvn2cCOT39h8FxbYWXp2SvtZoYrILaN7m1CfyFrWrcwPQqxFR3PdlKq
M5VAFkVN/qus8pdKR0+TMqr1Ny/fkbOgyXYbM8JNWfEiMSFG/9YrUFVCtMY9Sl5Oq3VC/08Ka047
o3ZOjK3jI6PcmFTbmNob4uJPaOHmc7IAOv5ynO2XdXeln0BQkpNBOvDyNpJKsoRamjqGuDQZTYMk
Nf7KfekiBTVkJKIFybtdRcrVcGXaod6t5aE3uXfaV30q79MRnkjKBrY5X10qdUJN/QEado5w7WK7
9Klv+yzo4ycXsVP8kM9FmhcKG8M1oKySZ96TeIKqpV/zteZhUIK3Xi4LaITwK+KUvBmGAbtLvco9
cO1BYFAw45trMHEMjl0GHjsGH0J5vxcfzrlAEsLpNaPja5sxXg2RlZ/J9gheDk50t+4NdEppGwz3
nwfjF1enHOn2gNlPKho6m5jERw7kmVUBBUqfWOxwba5M/idzJsZeJnOetM+IE8WX4HIzaJpzV8I5
h+VDUB1cqCfaJ3PKNdyofE1trTFM7gk13QZo+bwQQDcq+wVAZy8OJrRi0uc4ANG8qlDAGFrGsYyK
NF5c7DQVNC+KTEwO8DtCIpeB4zHZGBVevQZ71wY8wm7A1bv50xUAkzrLMRzxHijKkTWPpTy0q78m
mbGBrA/brrV+Zjw/Foc8hzBcRS7eYDNeHu7c9DobjxUXzdKQOyCYsY6aKILmHSP26ohUkVU4zhaj
7V7XTKAZYBl/lt0rt4DBdjFQDbXAY6W7o12meWNz7MCplURMBm+0wtze/NBAmEGxx9rn2sEaHrl5
W2U05dz18jDA7JlrNqCb7Yw2x3kn1IaPSYJQ3UZ5UxR0tkRz2hCdZCTJ8IlVlIrcuwrspeIcOGKl
ywQ98khwi80h5VF34g5MGnIBiIXcReuqdfHl2Sm5CZhXI8BJKlbFtfKsQ0I2y/X/nJTESrwSA/yG
C62c+SQ2a1YVnugtlnmh8ffgY+8L6nHaty9/cm4rYYBXU9mGBccE5+oNCPE7VGK3pzUpAp12Qejy
5krHcMrrMx0MdDejFcWbyn0dqzOXBpCPsG182NL5InPMxTILdLxEDRipG7lM8wTWAMSUgnAzGdPd
0ZEHt1dnLh2ZZsIFTKAZT5SU4LrvdHE7LObrHtD/vaE0dxr4NPcflbuTOcbPGQF/PEEPRBv2UY/q
0N0ppTbqoW0egRkN+ufwkFvf31eEHrA2xrDbPP91QUTETW9y41ZdGkDTrR352VFmxo6ngo3MxXmH
N5wMzrTtQlwEwh+hH3gI2PZrVJhMhkR8uUKaHJ9Sx0qw7j62LWzHkEMB9IKTxttkn+RrZdC+kt9d
Ofe9o8KJNPhUi7Gt2yp6figvi2l3GXLmfAsAj2CWA3Y9wzNuJEbUDjaNSOmyMQpFhePJtoqg9SlW
Sm04Qf8uTOJ+sb3DF4gJc2kUaUtBRCclVQUL0xEPb4FqC6aF+EUmKbVbILNlHPqRbZ80kC9+PzrU
Ttg+o0EhRfVJ2VYMfOURx6nBo2PcbrqHn7PHpn8gmJxtgVNANmwsNGsDKHXVEqvhrRt4y1WRcahA
HYwY9Fb6hpSc/EMhp2E/mZjV5fj+d1MHkMCqykaZzKmIB7JemFrXzKKUNaCd6E1p686G6NrUlfWB
tyu/uZYJAr4aRxBdRcq1IhfwfMqgAlDR7i5l5uUC9vG41z9G5Nt5p46vTWBRu/i97As6pR8U3Svm
BaAbpAOyAyRyfa2anzTfFDS8RmR55QmhViMu6XVCXWUYoM/anugvoB9quyFWW4f131FnCoaiKztZ
eAqD3eJQfUyh/DOelRKZek8ac7CeEfO8VIg7WZibcoeBC6nRSm771x0AiCLuwq+jJ1FWcZlJLahp
ETc73VX2kQmoU5fQDJK/jDdIDOR3WdDoBJmqNVitWEjNvBwvC4OC7YgJK+H1G7eH5ILFgBd5b2m0
SxlXGKs+vd8tZB/6Sq81jQJDQ6uDJS757y5UhPWlfpHtVV3fvZi13B5+IXZ642SkjGHdKIdWgz2h
qA6EiQ1VZLvBqCbtw+NJJSkNCWWtvHA2YV+8EE2ZWV2QSQeoidhU78cujxz7SLPL/H6ChkH8GjIw
hERTjMkS3/5IsnlfSQF7CjlYP54QmcwOjMqk3HjmnWAG88ToC2D44X4vLWDoHrCGoAbebpWnmmHd
zbRqeiN2BqQYNOuwvdkGn5WlGnUJJg25CMvju8Qc7vrkiyoVeY/GKhpfZGfN3zJbkbgQ3h5Fj0Up
Wj4VnZqVPKf7GZoRQTGx2OvRWA2opjx+aOmWV9rOBwwlqDvLcKgVYNUfpLSCpxzgweHXc9WFOouB
Ge4/MjF5QECt2Tk7pzkGRH96AxjOWazqFIRr1wT+xJ0wJ3qO9SfPvBQCxUWhHWg6D//DJij5E5EE
YlVAhBUHjlw2jvBHxDE5YhZXUi9cWYcB2EdroC/LYqyUJiTA+cr3pBN6ClVUc9J7WmFY4GMaZeCq
RKvr+qxtZH9EyU6Eb5+9f3ApPrPbRffd45ex/A1ay0I0lcZ6bim7c89sVbiQa1U2WYq7DUgeDrVW
WKaqaSHhEcUYcFidbb4/UksAD4i51XIPRps+qdz7Yj4QrBDlou4AeyRoGM/P0mNFcT7ZGuusgTdz
0BmVZosETfJod/9ps2q846HaA+n4h1+UK+1PFbrKRRymjd9u2UEbu2Wtbg1BwRx4TPVwchf3exwk
iRGzsIwAV+uHMFaJTwLQzUb3V0D0kVgCgczLeuj4xtFy8QwZaPWxcJFa7h6gGN/yiAJfQgAgJ1Ob
77jWTFCEDKyIxCdgb0Z4eCTSRnWRpsSu7ac1H6AQJQUqDpnSCROGxC0IfXTyJNR+2L/URlR4cKi7
b8pSw8fMICkQWFaCGK+IwrDIwRF+lVeU3Wvos7pLxQRMQrGIwOjiNXx3SufT29gvH9Esj2N83gQS
ujnEIGZhEOpqgeo0rh9rIVPE8Iq05Rf96x44UZF8eLsdeF5BZPFn4oep8rO/kB4M9dkZyEEaO/kp
X4Lt/mwPzdUTF5ui5QauJUG4SXbZA/Th8acwxsSHMS0xm04Idmn3qaII5pIaUsUAMp6wyImCggo1
nov7OIeu00l3g83TilX6iTHSdcjsYOc4A6afIejeGadsG3nTQUSf0/gU7YXgKoGfGH3YkmV+n7wW
WUtfaZEgIbgaFNG/v072YV3+nPuthEucmizHZvAqiaOeBhVJtWmTshH9X0bgXjTRaqkzh53lG3zI
Z+d2TpCaKAdHzVULQORK0iaDPrzgfFVLWzXn4OM3KomOWjqmke5EPkwDhhOUmm+9HPCMRKqDZhw+
b2ruUip3SJKoGbz07TD+ItvpPcjDLXc69baRaG1M7KtZ1ZDumCjzMl0x+0ZexBPq2g5JzZV6B9ZV
tvMuPT8hQT68OklLtXQnjqITdqxPbofa/sPcGXdsYtwDacJVTudMAplRndrgS/mrSc//eBjqtMW2
4KlqGKi1QBhYXJQ4sCBKJrDq+i6TtuBYs89p3yCdy5mC3R62/FEvizS/E/M0oaZYzMz/lUYkfUna
FLwNFCW8QuXHez6k4TFu8bql8wY+nN3QhLqbUlvW5eseoxMKMLIKwWHlmxDqJZsqMCryCsTCJz5m
EMMYQ6y8g/cHUFHVzqVHtLZMZ1i/e6QkJ3EpiD98jQwX3g2G3q5raGhqmELrYixlZcStOzVW44Jk
iBhJa4KCq4Q5X7xfyiRIawWax6YGzNlENjyGE2hKJSFe9D+K0HK1RAvqAqYihBxAT74DosMonQAp
GaX6QhfIrz34kvyRoP/iPcXK0rrdJuArDLpXGK1VV4jOohO/WMDv7Yi5M5Gh/YnEaHjH2LaaQDS2
lIAjtRZmkg6gc8/ttG5kBQRD6XBX/EkU7ZgklCm07qmQDwJX/6hEiRqWY2IOm0ERBddgno5Z8ptR
kaQnuZEHFWHOcDUKcO9wxViQsZkyR2ALUEET+3JqN/7tYSU714TbgFYMwz8yqVQlEoDv4nHNnYFz
Rhllm2lWgSwcOH/DVajPKdDjxb557BwPtlqcpQl6CPxj6WPBgLyjOfdTEd/r64wlxptH/+D3rF8p
BTxYwfWHkklUPSPOFRm1hvd8ZV3DjttgpOb/MjNtITpLJ1XtUhnCWG/k/cfuzruj8J+x+e4gmgcl
rs9ZTARrhkZm7Ppb2x2yBbkYXF1gJ/ZIt+bcR2x2UT3efZCJNPiGHMhcg7ZMYF+eLDXA7aS66YPm
dTscJHSDxY0NSU4M+QQ6xGkuM2A2v8wZGOdod7IVUKqqfWO88JWkM1YGD5CwVKjTbQHaeoWrORXN
NcVyaBzHacpqbX6Q0ZzDW1XiGwr9Fw1aZWJWn5cKBeqFwGlfKQRzBKmVoOpXnd/14dWGoNQGK3I8
Od8nsy8AcuyncXqMw0l3ujNjDpyqGraqHbmwdTImc0p8ImOXlsRCvbMQoLPAA4t0tqYfjeqqONrx
3AVQfENyk6Na3XwJ2wVazBPlD6gaqmj6wR36cp3Pg0sE/QrJDCfl/SQmxVXMRxRPWAwijPBfjRbT
lC3+yRIN/+xnS8KwvlVHwkQjGR2bx/vwKpJ56R6ipP5rSZ9vH1ubwzlHvkq6mA/HYgawphk9h19p
vLFZ2WuHmX/0VLFQ8Y2AWJi3bAd+OSt1d4RVV6/3W1tMTXikpWBm5dUZBolETPS/dFGUJgsTto26
emmFclA5I3Lt4Q1pzoSvAHtdwAWhcKHfgfUkYTEhzAiwm+RxdxEch2C65Wfq63hITp+TzLjVFB0o
R3MHeWbfiOgs4c4vlqpmZro401PdueJj8Lf82zPEZRja09cOrDI9Y2VyBt0aFFxMeJWT3N9zd972
6TS/geE1oODcIXEOHhooMWihHrfP5Vpa8uZPXF2N2qlboZu+MNrU3YoaEyD8vqlqSMKsoqulO+Zp
+liRaEXl/Z8CTlOgmCvHY2P4rjVVDnfmDhQRc1AOuqKPTPolr+7a5oayvVFtyo3xUEjT9vxDjE0r
sijKaOfcUTos8/uiOBHoGA9Fxq7RLmuBR12Sz2yIy8uFQ/IvZ+9r3mRIQTO78CVw7I6UaAodU/zv
HUhGSTHaQU6YEwm8b/07F6lPCI30eh1ITZZX4u9vZwfp1voOQT00kCfOVuhjCZl9zqRKTmNnsXPy
DAhAWvCShMaRbrRCl0Kg3rB9pFWMZArSftHMm/3VRQVfyaGy2/a+jVXLLw+ud9fAKJ1DOTmLb0V5
fIKMO2llG8baJr250orkUEMFnfpi3N6lGyd/wK9ba3RoZwANBIQpTJeBlH5cukMXgBZCPqKDmbI9
KPikXMRRk3DJzDiZ+dISjsdh89sMuOtonaqqmIXdWUKBzu/AyfG7+0DXUpA3eBHtggJ6RLsHrRdG
2o5W8ceZ7XELruZ1wzPwc+wYwGDd9H5HsPwauN4kAerA3N2WXYlP+PlgFGfOtwwdkBUMXmBzOwaO
eVBbG5RrP7nhhXVmTYkBsdkCi7PdojZU/bukqXoAKvE7as5jWjsVWaxFfmpwNlUN3ti2C6QA+mrh
TOvW1CZouESrLDHb4zFWOYssDW2x7ZjxXD4Yst99B75KNOqz+snmas/t8upIh3vjcRCbMO0H35s0
v4E+FSiGPaHGY7qMVk5F/4gauZg4hvNNrAPx1QXn8liegBCNAxaEFphqGC5pFP6Hq5v7szNTATdp
6Q12wyyQ1ypxStHT0Bv77rr2CxKGGVufrsOwlNT1qiZbO66v8UfzPbNAFujv0Xvf4F36YBXVm6oK
TzCGhsOIWqsEUwU1nQxvCxkDbNrfaGu7cpsQ3P+rDIB/d7xrwBLWhAufixCukOUCejJ7eIEMBTdi
cP2ITIYKjLVG/KgQrvGN7tCXb1262Z7VQPz5RY/UNr+Ltz4aYSCZHyOVBMw0WdhmITi1dM9e3Zbj
i8y1GBLLQF3FQO6qtyldHQ+PKxXYxYOD6x+z43nLBmuqs7t3MMwJKKps9RT23SFrP73Mpk/krOY1
m+4yNeqJRcnhcxy6loxfL0Mza3s+E/8/Rzpr/UM8DKhWzPCfluCGwoqgEmOTN9Fc0oYHbSfw78Dy
0Fup9NYx/mUjduAz+/9RCFjDB6lhKpNd58SDEWQb/DYqFid1BuBbrpqBltJUCMgOIoxAaXcWr2hF
VGek/b4lYis2bXdq6YQy4W050exH8w9rXC/MrphcR9LY8MeEx7lE1xKMUFZ4fsVpjA06UdvUI95p
QEWMB9MEOBF9bCgK6FSAtYFUMWu6j0a1e86o0mrgm0QxYMl4luig2BZZ3yWzNs8YM3m1yFoF4x09
5OQ45g7Z7RPUcfrIN5IIHnY9j1yCJKWc7dEahDiHdnDYcithcDzLDqpOJWGrXmLX4tTgrgntAjM6
abC8pFqI8T9kju9fO3mjlyR9+iSbzYoBcccnjwhkyGlzzX58g/MD2gFBJFkhYVnqNQDjyitJmWPc
VKUR5I6NUeuRNA20RTOPm7DYpQnkdrs4myXx4hFT0ju9Wwk7ySoT8SRyMvwB0/C+DYe9ppQUlTGZ
C4Bu44hGBdw9VWPW9A4G3W5sYPOwfqAJvGA4YbHcxQWjsCEjFX3lMhrGgjSeoMEEFe1wl9LNc/KP
53jW3lEdzIz8l+SqhvKhwPZdT3lxsBbY5UNgtzeQzu328DJ65ac3Zj2zKRw8Pdid0tNI6osJxXmo
GK7P3p5I11Jjw+hXIV2gcnjt9pOIHs4pdy42KzAOfDfuj2jsbR7R55MAHLNdvj8QZRPNPd7FKPmh
SK3TD1RwDYTHOLgu7V2mYxzhq7UAc5fSrzrenQslPhDR9mmpU/vr9pMoVZp3pPD0Onqo3IIhKK0R
tbAHn0RQ5xlw0igXl55sievfyau/H38ejKpLaXWc60gA4EGmnNdv5tccrFAzHRGuu/pyvXdeu1I1
eWYZNr6bJrC5vPRRAB+Pu6klEAbBW3mqJO12Ox9hmdzIgSgIz6Dj3UJGb2t5aPmlTp5hc8tsO1Eq
EEDoaEGW17C3PqwGzF7HBo6+m/ebrEvUaQBcHn3FDBtbNQ9wYRnBOSGVGrnliY7Udbf4G9fvTUrG
7WRIQZXZ4XJjmzU9PQn52Q7bpZq0ml9vwWExZlaorBJijzJADXoEGEDSrPqrYqSuHpqLHoFkAAC6
QjxRX37OPW44vbvY5lB2T7oKsvjRMiumnxicpNlgaKZCIZ6dghVedm11E8O37U4UVvKyYS7WY+tC
2m+156yr1Pqn42k8j0o5n4WfMRk7LkxCOA/fIRvTLZibBxEHP12JBt4mjQQQewSrRTDUngVbxls0
PER7CLA0b9IURsaD0zZD/UyLyrLC+24YYBgqinn3rSCmUkBzuyx/WBT4UJl2rKDjbibSPmYpDDgv
+VPXzFF14e7qHpSRvKqGoGqyn1F2xq3A5Ct6KcUkG98BlV2nFdxmpSWmkvjPJKt+2PlF61PlbqKJ
uokfXTYeSS68m1v1P/C2DZAJ5rkBlOMVKpIutOgcgSJ9D2Mm6LtutHoq9SNuXQdt6aDYji00a/0s
8UWPOhQsgK54JZ7bRFa5QfWYmNODG4K1VFjEifD7YPEnc1eIr9t3jYORMUy0a3qLQH/ezrwnZVMR
8Qn8RgmT83UJ5t/5ic94QEpxLJegS3bFP0OaGKnb/k2E33JScnQBRaKJOPoXvKmGouViUU7bkC29
LhFC2aNwr1CKLq4XasSiqjEDAa+sKxWfzkDBfFB5AITnJDvb9yeTBS1e438d7VRByD8rqIFGVugc
jAjGAivr4czE3YU7BLW2rgLOkxR4EVyI4o6iA+iePniZt7XG81Car7AhE95VbUrDcR4XeTZIhGXM
cVxIf0gUvSkuVFaBFa40YAIPco5jIYUSXoGH958zeABo+jsOlo0PmTGJ9ZTVOeMthwnJT9IMVOXp
Cc1m6YSZyP1xKRKUsYTvLSp5SHKi5lp0UueAn3f/PmnK3ewUj2YATEvymEbuea6Th08JFsQSwImP
KVtvz6eiuJ3bdzQ1gT9hVjX/nltgWyivFccJQ96kdYOsq4vwjxJ2F9fzt8+q/oWeIt7J82n6Fdo7
It70r3oFTWXINmfyEnoon6N4ox7JouvwiafcXNYhN1NmT2SCzIj/Njy7JXUyWJiyYWYEuLjtn907
M/k4D+109Hy5H7cc2oj4ojJWeUefbIX51KznBRs5r93j+ZcPbnr+6EJJ60gkhdbf3LdHAuAfH5XI
rEfYhRJfabr180RDII2MYliP97Py0bkbCJMH2yLnHNirY6K+zVW8pUf7QcePleUnRbminbGZ17/V
yTmGdgNdy2366EQ3yEYXuUoBk0HMnLG1cGqOz5jIwnkJP7KPwLCt/KQ7/rZuSk4442icwx7tb/Tp
+y92YUsX3PG8Rjc3WpbZ6RtZqVh114LhslWs0T2Z86qnJGGygiQl8P6LIyjRNNqTKEx4mMzrP3q0
EaIJZsJPAUFQai7noftjH10CaEQL4erEFeatKPiJLjiDgPZhaJAA8pz+iUIMKnL+grUzMpf5KdA8
F360OD5o+Rd6P5DLmsbPWgkXTw2s9/1YJVUfVmkxqjJQsEa1LqMfY4lCjXpD/zJoS5bF/XtmwONK
+XlOVW6TSTnHYLAN2kksERy8rEKHpwCzwQYLaz8LZQAjSTduQtxb20Ac447DFVC7Ront2yhXxvP7
+wxoIc8mbZ9Y/V0ajbfDgVgH6Uc3hYycd3yTM4CvB7xeBdMWkRHb2ye3f7LSfWp9CQ2+Li5AEvie
QUqY7lxzH4msV+iare8xid4U5f5LUCFiQnAaXZNYicyMne5Iqx7jI8gBKo3fLE9Z3wfP92+jZI2H
yO8yp6kSB5sT745vQwWQY61ED9RlO4mQTaNfXHcpbw+7j2ApLa+Lofjh5/tVWMktfKh0o9E8mRu5
a9SubQEiyIcJfKOgPn/Nea7eZpLKP0SLMcvMjJ9KOfgSX6DsMCisF1+iDI8eXFDWc8Jo1suWOcJp
AvIHQFwi/HpF3F8DBDrdyTYh3lfd2esVMyXGRu1UJ34//j9FvrlwWiVKM92ZMwElF/G7BhqyZXCa
zlvlP4/M6nEXlijhd8V453SAxXS+uRjtlk+3nwvwyx67gMK4k+GUm7fbAEkHL6Wb8EbpI+1JulRo
gGw5vGRFt7OqzOl4AYS87ZmhmivEw99VhpOgEMvtNDPbiTW5FHn091e4L1PzEC7U7uz7PDa57DNy
GG0hA1NzwvwcwSwAeGOtuAr/QQQ1Gno3KLZEwm8qfGCQxPhE+hS4pPutpoq/JEZDHF6ib6v2rpYD
b93RzKbjUJ4M16UTgcfORSSmBPSRzO+RwM9aMl0AVjolrvv2w/rnfjrqDparnNKPaf3kzoaBo2f9
N7i2PlRqvLvnvyeWodk9/hhgRphrShotNXzn9WGNsTwCpQn5JDgq30DHEtERN3PO8eGmawgQDNnM
sO4/t5DKh7t8XcrQ0wlgpsGZYzcLJhzOJr7T0wR95MBFjr6+hwET58pUC7KeCIMx0TbosrLi0Y7i
S9RL8VqysFyGnnrnX6/Tnmu7e+LwTObuvvbRoEDS/Qan/+RcuKbZRX4spmtqls1MDbNTN60WnZaI
QLRWOkvivzryCO2OnYNvYXuIQyCJXPBOK5tKkgFNINKZc4telJr+MW5B0UIt2aJEWlDDfVOAJXcp
E3bB+BNlP82xasn/uppZK/6MJ9S8jOwK+B3oU199n+OclgbdOS8bWG2sAMI5flMLcvnBGeqQ+BZf
QPErbPLpjsLb74VK/nBtBb3ooVWCdjvyGzcJ4p0tI1g2wagHiq47vzXhU2yvPjY+Z+hFhJibOolo
73Z7yKnPInnx8hAEE0ayGvL8V+PVV7UBUtQhxH4JLWkH07IMzpHpGo3yPFQOZZGpq0jDYSDHcBGp
8R//2SKxEpnKSDpnIi08lBBefltHh6zX6FZo6pKns36xaIT25EfdK3KzQQG/uA8VxkecdGDJRzk6
+upq59tnR1AMakvs0BHe6+quzhRfXOUdFhtdAwL91nfsXljRZWfYV4Cjcy5AuPeI2KY/6YXxPbAh
VYihz60zLa82cNWVilzt3c516XWeFcCu6LhDV8pnSUXBjIe4k6LcstbumASFOlHmZw4BlXjIdIrR
AnQfiEFq+HwEMxchFdIAiUgKdgFCP+xfcJkzzeE9aSZFpTrBEnka0g6yuq4gGEqxPBlzcex4CGIU
RefLozMvPGzTEzCLbRG5Bg79crzTB1R2Fh8ntexqitTP8AmZfTS9HwOdTCHED0UWdKB6zkA1tqTo
8qnNuJwrhSKTSojit/IeYTWl040JX71Bp2QB8l75LuxNLsilLCgRhv0sXt0AVwjEDkPv0iJ3xsFk
m0KCIRiRTm4G9bqpWlHFm0n3OfIevRLVN3wAJ9+jumIaoDtJAgEBlAkg4Af0AID/EEA+29trrBFN
ZF4Luu2lh3taO4+jXdfDow7KJfuU6dcU2P+K1Lk9bxp/APKyoI60FpmhsvPQeJCo2Rk0QjUR1bk3
kFTpWY6EkbY9n+PthidskHvX8ys9aYMKMNUbOLgZkHFziwP1ru4MYs31VOtM/W/lM1AK7U3FIEcP
82/ftNqBb/ObFxoNimlwzfOc5G9mHT58gJWtyAqb9c5MRB028OgI8e/AXiqUTM9R9pWidlunQnv7
1zQAKRfpYcqD9yJaBdFU+4PJELK1bgcZey+UcWELTyjNi5Syoj6h2pj2jMskuXMK9BhqwueXLyBU
bcP0DiqpjnaQRsBZGibvFIjwNZpXkNbyd6VUuHfmzVQocC5WBDXMYGRTYCq1SMwbrG8lZOM46YaP
cITso27kPqxWczwE9FV/nfsVhoEiaEGFdxkG0sf55OTuoJQWa9wJ0x1fAY0ANAh1J6wgA/a1nXhg
6tmF9EaISx2r/M8p5NjJHD9bUApxlfSYdzM9fjciZmAM15lwcJQJVz6r+uJj1qysW+mAUU2XLqNS
U7Lc6ro4R1ZtehcHKuGL/aE5V4gkH/qm7aeBMo/fKkFr7OuJfwWpKq0kjVYJk8J2XhSyuTwhSOc3
/9XOoTO8QGI2fPoQ+aD7lFHb7/SYOmF/aCdnGtWFt9BQHqc4YvTLbuXrAZurjS3STNKhc/PbXnn7
2g8d3oHneeWPJkQ4M/us4HlMnQWg5yONMgwo9slcdk26P6Ud0Zi5Q3FMKdFL4IZPCDDBUx7gOHTb
vayjcdvxIE8GmVbic1k6S+lBi+nrclLsV+mhJC5SKPzglUk+fG9dgPB8E5wqIW4AYXkR5d4GJ2sX
l3jlySTwTqJyMmW5M11mAtBaGdNtYo7MLK4QZ55pF9MBuxM8HslDwb1QCsTos0LW4F3yyjll4Qfv
Awvv3ct3Z61nBY8dhbphiOoDZr0qOnsDC1Tjp/xEC0w181bVfnnxc6hvS6RROlN9/vSMUGtt9dWp
munOI6F6ebnSE0Npcbv+vxbLcHFVsufru+bIuhj0YnJsHXDH+HedaSfepJUTS3VP+IFt6Qv/KQVM
ucxffe3M+Dsy2G+lJO8Rn/PpzfDo734JWXE+YLtQ+Wl5Pn+z5YIaJ+8/5r1doKJ0Ta598aFYfUbO
BcRk2L8uPOMaki1o/UW0kvdbAmjv7pXDUwIjMN2QQ1FV/vGuLsJICZ3eU5Oer5N1Jhx+hR9/3n59
Rtw7Gb3X72MjaxGOKuua2rGdq7xQMG2DDIbyMqdlEZRrqzWXAFsO17NkUFI+uGCuVO+EGBnAEyEo
PZPetgSu8ISiknp1hEG4nC/75BlzTIgXfvgwFc0YUSKEdPyWTg1m3guc9Z7k9TC/gyfZIHHwSDsx
fw9k/4PmGoIkqsRZVawspUGEG68GclvsAiVAdwIzNuuYF1iIirl6W1NE+PUTUFom7+Ld0Co2a51J
W7GbRdcOI+NLkFJRJ7MxL+lVrVRhkRLf4lI3/A2it62njYfxzG6BHAPQBG4v9kDim+hS5UkdinGP
ShZySVg3vE08Awr1zqky9jaB1CwTel8GWWoxNjEad6ZB8Otn/JNna2wUQGwPZRwcCodg0A5HUOaX
DzmrKI/zpEfB5faz09l9Zari4/EO92rSm50APUh4UKchLMIwgiKhB76xnAriq7FUQ4YnOTWISXs3
bXJctfbmRDEmmMZ4B1zFvZ3pEarA0RvLah6rb+DVx18tDhLLHyRTI/xMXwqLHdwUkpn/1JUyMuX8
cndx7RZKuks3INkqR+7sYJEju4+iBHwnxMyCAlP7TTNrsa933h/bnsPzI3Ia2ho6nw/SBaaTzXrM
ALzjnpV3GVrc3P8AKFhaBDD/OSYjpKcPpEggkcQ+Vos+sn1loU/GKXyyGXYXZ8CL+0UtZnQFewHa
oR7S5k2GchOvDLpVxrPcDLjqN1DG8bnHaX4n2f6olfAIHWY6aFY7xJyir5Z1e8Xf4koOjttrfSO3
PEkTps+p01gzKajbUWpgL/U9P7hUM6fw2XUBb/62KsZ+ynLTVH7BK+WhxYmzCmpjGYh6YIybEYL6
uKRP99c7wHAp/UhdTlS3UVwZoJh9C1r8WiKC2ohwIeuxwxl//GJIXgyX2aNRVJp3wskS/r99/OZX
EAUGG0ueuyRbh9DI29L2qEr3y9bId9vNvFI/OyGREe9IC3ajgiXEd3CGJMEbxT7nTTHdsoXzO56N
uNEiMQBEowHWMT9qFOylsTZenHNaUgMZVOcqiejjl0AwFumooo1pR4F43IP4Mz4gbOQEXJnwVYfi
GrQHZu2NAb+uIb3a8Z3zzUj5E0qpPUW8gW73IvOLK7huGkNpL7F7F4rEZ8EXwzbewucyvAriqbid
UOjhiIst0nuWSxQOW9KdeTkQL44L9Aqcbak5BxCuL19WC2/FQAn2067qLJCr2MfC493ZkDNf76VI
cBmgXI7peEjIQYbrWefuP6wlBuNMi8sWBMcbddLQrJVOzI0/93DXwlyRbZXQwGmCy2hbHdO4GoF1
LeX/zREw3CJywmSiMThYanyMlj2CgPhvhVqCzws4M/SiZ22NnOoLWrfFw0MdjudbkNsFvLjFN9o7
xh4koAxOvZXvBkky4J3jdo1xRNddt3ZUQYVvUX3dnb+ldj3sEEmfx3kz2jYK3exE7LECcPnnUa/D
OZ9wOW2Rn9e7Y2uFSqSv8ZcnlbtksMWUiL1WpFeEJGavw05S42N5Id5kKPXXcNvgQpPAGL4/VPE+
JdZ/HrHYtQTa3CbWsKKSapoHaTeg0aCdHmSLjChe++XOyRDNFIQaspH+Ay5FzREmlAVcQaTPc/ZU
okXGgeA69LoRXclpOGhPZJLhc0DCcWBwKjshmw2+thusmYZzsTj510vywN5Qnrk4OJgBNP0Hf9oI
UvA/96GnYC9+nJxQE9Tg4aHwf9Efhl26xqr1u4rDgT3l9g5VvmfnWDMxVAntx7VCk5xgPfABlkz9
PsV8oRnISwiGpdmgwEmkWr1p7AS6sG2NVKZnR4UfLJ29FhOz9mQJkLOmPPwI+7FGmsBSIocJNwsL
GJj4x9bTM46/lbA0V17Mor91NzrJdNi459zhN7b106upA2sdJX+VRKrQEQmxV5JPUV2NagVqgpne
3S4yDjwYODvNHv+Vuo135ayrDEPBq20Gymwf3TcyrmKsAIj8PDkx9FYymyb1p+nPwESfFqV47q4Q
1HMhx3Sdhbp1rojNA8GYE+j2Ym1SlSoODhNSuvfv6GNvX1Jp8n88ILHidX3kCdURwZvBv08S+TB1
8K//DHlUiToDvsEeCmeycDnALkxToqHfXkExpHsKwQpvLEa848IAPijRPyJ6pXdi/46/RueY8jVU
ScTwzijR0U8kfMvdfYm7EDzzSmvC6W+KtzZIlLPtIM60/fabWiKE8uKEjgYcDD6dlVA782Fiawnz
0vfl6ZeYMBtIFBFej4JDxyX41IosfaXoye49T6xcULxtdYnUIQSPQex2+KVjUyaphnEurYzQMZ5P
3TXAMf9xTpZ6X50o8UZZ2p3ETpd0PgIRsz+BDBNpzXU26QK2I6QynEiBq3pKVGLlUFja4+fgwb8U
WLWoN+oD7GEIHqvhBA4NFI8op26dqRyf9Vpcd7e9M4wBn6l+xEg5WRqYjdvel1HvypUD9MuUEWAq
yuBNfmzTmey89Hahq7xq3MtDJwi10/YTnh7X8l/9ch/MegQUmyy35WMAX0mNaZJWIsC6ECW1y7jI
SgCTT6KvbXyu4x5zbjYQK7hpQseh2REGo/7MzbZ0AoZ+HVsyrTTH2DvI96ZpLrI+j/B/PHBScYHH
Nem1wN42OimLEKcJYz1k1MncPlVzjFrhVVkizIVU5NXM3HAl+qy9XzPMPf+pYdJauy2ApxLLwwhN
UZAyk3B4fWX0WleeU/JofY9KOCUCgxZu2OgRCnc/CejBqB6HW3DhpKUFfbdurupJEtjBCtQPVoaV
tw8adkw4q/KmzULX1sjKrPCn5+CfRKcuaXUoh7Jf1pvme3JkSKMDqeJAtaZ0hqF+jOACkPUh/jUw
zPu3fWgH+BBhN2JhDtAqzE/l67OsfzlWFL+o8wk5r2yGLDxupO/DrqOdeEd0qxl1ih2WimOL7vnD
sjvSPFyUyD9cWKhUykSba1S+pZ3/3I+aJ2AzDXwTtnCqNCasnDBEDZF4+tEhkxz3AzGNwGokAvrw
LhPA1glaRLXPDLTSRfHhaXWtk0aidfQpaoFWthm/V4RVP52/F5FhhZvbRth1Em6rvHYgQn2MDO2Z
w/sM7rRgwSJxcC01wtLB1NvVxjsDQrq72A0lSB8WeMt5r4Qo0wsJcbOs1QXJ/zJTAHl0zLVeHCir
MSAHM7oWSSS6wvUJfn08gPXDLDFv6kPLBzuo+Lt+nlkmz8Nr9c98gkifOcHLQm6dRaINomcGwAWm
RFwnI3av7biNsOHTCQs1a8ZtuIseheDVJuNK13bYGRzXNDn4EfR/F+BZnR62P9z8FMgwq6e5inBU
nWCp0/JvNDbB1sbWOHmm+r7FOol1JtWEQgItOa8a7ooDKetLve/grbQy6JRjKvUf3jArz1xTnizp
/EUMis9Rm9xPpVThhBur6hoMwI5hwC1ySghXKjnYUakFikVtlhnj8SZRlG+waFODkrMTCrjG6ill
unSB7BVT2EvGzPoIQmYBfLBCWldQeAKVGhk8wroULEmPKwBaQyhIlymijS6o1bI2J/+fsGu71mUF
bZTebyHczGKeRT/DoaOGBGdGd/iLzZnanG17BSo7gsVmTL3jYvfp5Uk1XrXqaHvs2dYSictOxnMz
gHJDx1vI6LGYEj2TaWVgGFk8ztxfjweVjC8E4C+WaGTsTIpln4XHU/nDj7vWX1l06MuTGmEQviDC
49HeiHfl91E5V8tMQXaRQY3va3b3RoQWHYCrtCvoG10puBRh4vSsUSZGjajpZHQj3ru8ip3I7YFI
xzFmq2h0tvIXTRRzymZyA4dsFVriTf+g9PzvSomSe27S54a2IMOgdfV3Ii7wFzJa3ejW+HNvZUwv
Y3ls6kFLiIOSzrCrdhmeOmPR+zo5c90XK2D7k0b64OZseykFFiGnc7m7c4ninEe1oN0rMZuGXsek
sknz9WDCyskNd2k/NQxKZu9tthNynlaXlcrI0f0wq/cmk0DSZsrMpqSRbJhhXTfM+nArF9z7+3To
858XvjXD5QqbzPwwQHWmNzSn039pto1jkhuBsRjUG8mR3RvufQRqjhsI0CNlLxCrxerSbPtXohsu
YTOufVxlHlkWgV4xZzLBMLs98E06ZZStawQuR5yE7pKHUxBnQXGOWqGUUlMeGIPzxBvr62PWw6m0
MRFCImudugEeIfQ5suHe+tB39/h4iRHXaY3aunFQv8OaUtmxp/Bcqhmgilr1fM/woyBEX8CIha+3
gSLN/9SKM4q4gc79uf93ueU0VuUS9O7Ps0A0x7sLmkxaAVzh3XFzt5il+xH+2Fz3OCV4lqIAecZf
Byd7m3zasiDgn/OHlE0TVWo4VFgeB7XEyFou4k25cNnxZH4kwg4DdKRkTWMkuWhrjw82uRiuZmfR
tB5zwjcgWJ5aQYw51aY/F/YGM5hqEshzpOvjE0SSombvHkkktZ/TK0BYU26/ROvGV5EQyn8OMXo2
y7f4a+szOHK3Fr1zHXtpkj4ZGlLJjWJxAm10nn/HwnjPfr1IiL7IH9AdTJjO6gL3DDKoamZ6Txrd
xjOB43JfizE/t4jLFqBe2I7aGck4d5pnjHQHq3txnNusVNNj/luqKxiv3aXdNplfHG/mcj63evbD
4Z7ZeZsUB6T9cTX9LxITZfNVgLIeN6PSyfL853BvLXCDRquYPI0ETleqAtVDQj1Iq/PtU37ei+/g
mmcMXcLTKu9tH39pHtR9I/Ov01zguwkjPB+PdmPrqQsdIpGxDmwzzG5HSGzING8mcba+0Sa6u8/G
BGcb/Cr3bDOjW+xwyr6OFKCUutCfM9HdQAXvi1Q3yijVDVYrJ8hjIrJz64JRS+IutGze5mPzAryC
pSLofsMRs5HUBw/WK1/qnD7wJwiClmiM3jXhDT2cd9+z6ZxaevhrEHY5WDEflwMP7S2LNS+oga50
peEbm0xl95laxL2fhZ4P6tuCp6EvlBrLRDyRhngJYDmFfBy0SciNdqw9pJqFI/XU4xgCGeKGwK/q
IRV0hL+Ewn0Q3GR9qphc1P3RAM/MsQTUf9GZ0t/XUANAqEhQTVvwajrwtd45I2nEy0KiLgLWe20t
dnePKUGUpRtxIUgwP2L+7k8MLAzBaHe6yrS3KABNTRNbSGutNd8QmxQkvZ6gTUyGtNCmfbmGM6jT
A82sFu9TSQZ4jJg3MHrKJ/yjG5/6Q4nZErWHOcrYH7HuCqvRolVUBTb2yKCvCbHVlhImlAgLC3LT
0RJNI0bslM+cG0T+cDv4mOx9GhjUWK7TkZiUuhiFNJhnE7Y0fQ0NvZsmwQ2XNFama9CXPbDQ225a
74NTOTcgElS0WoapzGWVWCZyMteKsADrfCDWJQ2XwpwaVppC6M6RFFbphfWRwtO8+yA3i6d3f/D7
oTmBXekusEMgpI0Ji81+/aYj4n4OTvnFOD6Cv9KZqSS/9uZUadq+8vxO/KJFUI/aom6IdA6TD8wn
LAZ1DjTokKvu0EFIJwh+g3Oy5Mu7pQIDCK/x48HA+LTAQwJnl7VC5A/IUM5y832D4HN4foP5E+tr
fHng5nIMzX5nbK7Vld7TBoTiAmTdU5bu+uc2HlbgwhI8/fWKNNMbdz6a/VHE7dCDOelCINmLgryi
vPuTOqwJXAYM4qnhN/guWlYDfCeyplPi1sNa7FKPHPkVxk4hk402ANuG4MKsjSEEstuSuW5IX42f
aBYJhx4g9gNh6vHgkNhMf2+1h3K0U5qhHEvnE16/mFxgTkn18kjWorsvYHhfOKithTTOgKkCn2bI
4ztPc7rp9Bx8/stz0GK6cAsHD1Q+woOqG7acz4tNjnbfXXucROcKcY38HcRK5nINDvm1EYK8s9JU
wkoAyqGaTD9z1PTrttEMxgNF+icmyV/Pr6WLT4UVRTnz1zCaHQswukukI2J96yBAspIxOjt6vbjj
kX8aK2nulQEaZ2JkqlAlz2L4Ewa8HR0BMVePAv8y6cCIjuqSFJfkgmaVf0pcLPMGLdVj1pkacxmc
FWRZYngldRB5Xe0iXyl0ET2YZA069sWr5hGlVyEiyXpAVgdlHhaAfIDH89Yu3Grl/QMTzvuA1D9L
oXvBlFO7K9dakYkmxngFmToNBRnSXuCmOj5LSiECZO77UZRWuYMh6UDzOEhgsZkCeYgm8hNGG17D
zrfEnX1GAbFO+dhZdz0bGyb7v8xc3NuEHoOe3/auukj9RJexy3n+mtt9fLHTs/HAJebTa2kuzWJi
yyTSZlAwycTH1U2vtdwJnvyD0nV9cZMbd2uYU2TRnVp1Nmbpno50lBOMRc04J8facLhErZ4KyqjI
XdmOgW2DO6Q/b4L/+GuU4cOS62EjReZuVgWy5UFopJPhKaKmEW9GqztymSylp6FLLKt3kMwOzRT7
Krr3aslhvdN1HRbI18ORdADV2MCXFd+Bx48qx8/IO0AK8MLPSLb50fNNs04n+rgY6bJl3RVACY41
i10kCYa0tBnZ90DlasCkGME4tDy6uRArk8LVfC7jCPC7kPkjukLrIjp2xQpeiaoZNOOxnz19vhxa
CdDE44SpPpBqPy6bRT+OP26AsOPbF8uIcWvPzXevu4eVZP9tkMPMS/QCfRVTote0j8ctP4Em6B3u
cL5hoILL789kTKj7+vy3PNezKl/FtPb8DY1f5Qr+YNkZOFDqD4QUCtoIfdZ7n5D+2sQktvxi/WEN
Pw0rSx875xk7nNav+e5UlX6raCoyRYc6waGcVeNq43cSymJanF1aUBBONXaMo2f9xcVuq7uElKjw
IXXZFniAcU1KRAPcRg1TXCcSx634EJL7FcIQQGP4dG78Senlvyf+YJZRsi0MCQlJG//V33KVqc/z
nreFSKtANDIbimuagLSgHr0B1GNkxDewIXTJnBy+RPf0RuRLIaSvBH5n9Ogqsx9tA/pHu0W/BOK1
CObIJM8mZWh33E5ZAtQXg3zDyVoprDsYScSoJyacmAtOr2pFrkEdz3t8Zx0iYBKLCs/bAQ62CxHs
BODx+rkxgVQSDhnAz0BXBYCCRpHuZPpPlPVQ2ZIYg2NdaVNcSk1K94nXWiFawfYjHUoUXzic0tbV
Wi4Lm4e1hC4uSXOF36Gqux2GOwHIBYoLSWGblGCxWg92hAG57wYjkahQXFTFQyY22ebQXppoBt9N
kTA3L4fgwHeuEJN55DqOcGOUTORSqH4dMzPTTP9lCTRKATTEXQTmQTVYs28Fy5WV0UrvqfOissuE
WLu5ccIyd3s+vhlBxBoirYMCRp6TQproLzo08lBC8Z26M3tak3oTk+vmyCj6sLQlWy9uJtOKaciJ
qKXasH+c6QAT74wHAAv+qoS8/vyRSJaUvaSjV1etmqvxpCVxh0mqYipHJ1dClvqiA5XPBSphj85E
QocozPiAcGIWlu/Sh6PkBVXtYpDlQQ/Crb+2YDoppQ3EuqjEVzyrwJFBNMEOO0uf5JiihE6ID4u/
uMMRkgb6xL5zKuJ5RuzA3xqOXHI9a/VdAe0Ml8kbW9UDTcfHQ2YFSeKDpFJpFwRpTmATuPeXintd
cM9uKnh3boGhdXzqy4OUvA5xtof1Fag5oBkRvA9hk/SsytGb6WJKT3OZqhkbOyEeGMiN7h4BfPhb
+5OVpZrtDMz78DVFaYIhD3fJW8waKTIkzR0PjXiPz/mtIuw49T5zrBWCEOEOG/THY//4wOJKuXFK
QJjqOrYJ4xqbGoBD57wN06wVLQJVQSd/QRWdUiJ3g+vsnRcyf0rxBw6qcMcUhuykmW6cxZctrKEB
6VO/tcJp+jjWvNwhrwMNgqSAkSnmbniZHKXTvhsWF/Sr57M9dMBWdEZZdUk39P4B5S3995APCC1E
oAcOWjZq8M+XOsslIJw/412jJ3lmRrzfEtI3DFQSTT5mP1b9l8htpz62zqkhui4WjzH5M4GgpBNu
NEEtsK2JrZ/yoMliAprwva5XjouX6SD01kFFFKIE1o2eq0sYec6mAdqtDVahwRmaa2j4fbWpD+hz
STVK5l2/Z0EuAA6WBiQx1F7O+vxwOyO284RPQ5Jd9FNX+iF+DtOYRDR6xcwPZSItn2usAFj1kPSr
5oryqKRZI1ZiLvh3lxdj2MkkWXY3NMjhDbtsPFiDWGEYDLVmvl3BlrJjKJwUJJMdoigfNqr5zJae
/z76Ll/nKp3Mlt7fbjQ4lMiNXV0frwjz9G/ixOfObkGDCSeyUFk200rgPY6opgCyzQQ6jCgmgD7o
YM0ZwiiFS4KDw9kGrlBL6oNNf6d4kV4w5f446uML2GCLa7LGresO849jDAuweKu9Z9GkursTYk/8
e1zghm8YZLL/i2iPEQ0iVQveHUZBk60d06uFCrdGl+n+ARN+NeAINvULF8SMU1MCCzWVqO+fEpA1
D2skB1ucDbss4aLfi9ENgqy049lydrG9I9gEvX3UIuS0og42ux+qoYnAlhANK2f8Cvyox76QvCzQ
ItG0AsFQt12bIpSTZGBtcXyALQeXI3rKsHWaUPs4+HdEnaxJuLs85E4cGdaB7nFGsXlcP4qjYf0A
xK+UnZp4qLHLAORq6QcrEW1EpOdSfrh0hcmQX/yuYLUtPBomDIzTHQal/JdUKsCC24+119d1ocdz
QBWTpNOnPWr8r/vwY9k+msa7NN63vifd5jJl5YhlBEze/tQiuyS1I2pBr/jhGBPgEysojpB3VBIg
eHtFCGyB5Bti2fm9Jl0lGneAIs8/uHkhE1e0fM/FpwpvLSk9QM1aj+NVdhvQu837OWAbmzMdtQG2
B1SIOYEjXk3SXVTCARo7cs9v6IBES7q6mX+KA5ZUeRvZo7gosFqsElpXylX7KUJZO2Qe1HFSWeNs
AhK8HN7h8aMY2sNK+zv58UYpz04a6e8/WU4o9l2emuBjTne9SeTbf7JkuUrfsjbTvbHEcAwRZzJH
ax4pwC3fcy4Uug+R436p6M58/PgEU+KD/3IQ9CPl0TqBLqmX7nuvd4l5DVrAwwpGp/SD433cFpbX
1ZTgV75KTJoam/+YWLXR0HKh+Cj7e3wY4oPUYWaStAjUqD64S8Erwp85Lbrmd8yXsZznWdVK8DVd
9x5e3JFZMYJ4RMdPMdeR0K1ZpWVYLu4PPAhemNiT5Bl055HVVvqdStjhMfuJChH1bn10mUK9O4uz
uW/gmGTGNfOjOG1HuUwM7oXx10qBkw6xDf9BQGIjnSX9vV/0BikPRYL5G2jpbZBmINBSkpfF4K4h
XHZVv9RNm4KAgNbZX8+rfEXRL+augjJymx/T6PoeyprjVHv9NoLO9xlSHknPNeW8bnfJHls7DGWd
YRKep+l/BTV+RTnc+sYPUoUjssgZbEvt/Jp6r+Xh2B43q9V/QhV6CW9nDf0SDDXcTryf2vkYuDT9
sjjOc2t0DfYC9BLXKA14DPomNF3F5ZAnOIZuy/bXAhy85kEfQCf1GGq8U4BMrHjMYAX5slgPGLG+
QI6hXtBS/k9JrCl9sNwfUdKly2kzBDmk5oRP4LDLA4OGuHA2I/yMFta/KqoQDXeo+BbXihMf4CeH
tcV3VU3+LGRsULdJKbi/F5eKUF0wmylqZ/+akuaVxN0UBnbunAc0Om4ZqO6pDnYPZ5BSLULCKjw+
sVgRtR9dR7LJA3Yl0mG3mxTr1wqe+5mpSQDucG8XvMDFZyXxhmBdSxkQiCwYFzHUOyJUYUhPOvUs
EZqxwABfNSBIJyuzez6tvYRI/ceq4ENgJk2VJSuGzjhnPFrfRZHHaZMl3a0PGuCoi134Zf43TXPr
9cus4fVwXPbI6ImZa/TQgt/jv4eeUFsPKvrI67S+nLrWt6ApC3itLSb20wy2s5TLQWcvpfnHi7wC
GiPyugb3UtSlpUVv1untDnO9TJyPglBVfqT7ewy6XS8bgodEfKSW2N/hArhfPqPwFh4WVVbuP1O+
wbbu6ZSrYA2FGf2nF7PjWrTJPV6sgbv36to4P/0gvKOmyGsxb5gWDP2FTbkKTKsW+Fj/OSbaqeRU
zecxivH0gVbHXoBmHsrDxmMpIovkRQgD9YimiM/H5NZp2C0sHsqYVq+yeqGTyg+GCqZDGkGtXmpL
q2Ncf1+nWUvbtU2ZJEErs0nUCeOBQ/GRU/vr+yxxfXYuf6DPxPYzSxcFucO8BVjJ88H4BDnfvaH6
0Uwn68hAMpOsvVYaksjWnn48fFE6dKPFcXSidFNaJZ+wWqEgaHIkMgAmgrncvcgPDtqyjqN4rnXo
RNDjIAcSG0OLdSnOoRfGEFMWW6WjRRJpOIN6icSc/rJn3mO1xNenlCrruQuGi4Uyg/Tqo/an9vCD
UKLacHeAqa5eWyZVU6EOAUjXfCWoxpvaVlEn3ojUsty9pqnNKeZfVfFfjFzgg+8pM1Lg9FsZU2Cr
wIrX0yOyPI4LcsWx7VwUZkuMdcHs5UgzabiXnqmuUWFey2qEQ2CVA3/XzFrPJayqNkq9sM7G7Eq7
75nkABKm79dQGD/no1gvzDhUAqFq6me26K0NB6ENPrkS2Da3oAbPCLVkaLL4QWWi4BuTbYK4EMou
EqTjV3cn9tUle59y6R6jdmlIQedp0EX9HjV3mfte+Qcz34NJ4hYTfgCF5TO5XofW+KLFinMmebXx
48iZlnPdf8DNfrJkGArbNx/aPq6QcKm75BsgHmw69p+dvR4Si7TjTK5XzWlKx9WdhYQLmytGVL7g
YDY0C9UMPCFxczz/KMRK0qS+D8Ufvkj5Tesge5MjKybuhikt7UoqlHnuGdYv9bUOe60o7f6ftSWk
ONfXsuuylwVjCp6dVTsgBhXd3GqVN4bk0GSRyudS+r7vcQ+zWw+7trlCkkM+WKxXw+uy1FPGYylG
UPxf80CNEzliJmvXiDqRVyRa+CmkZcZc6G7+jFpugnLOjM2Z7RjtjofWrOOPcw7ATv8p79rhNs2G
FtM5Ggglf87E8OPam/rm4dXjWr5V3MfiY5UZnXBDSmrDWYs04GjnZuTfLdaa/GyHZt2mmZ4IvS05
xHkWxRI2ik7FVT6TvNZlYX2NoEZWLrsUClkB6hN65rdPe9VHLNF3numG6TJT+f1P0b3559lm/Wmv
0hvG0/9v5aTTtntQMuqutuWsAPrxonyhPTE8AFLSBD7HnULjpJnQDXoAMMoW8eRpIYJDRJHLTGd8
eZhKKDQDACeAS41pL6GHnZZbiNPtZicoRdlmmGQMz2su0ZukvF0yfBlrY1PjhfU1Kig8PI3znNIN
ziiEquZxJ5TOBLgParWhQBCz1CsSsy9jq7eGNujLVeTNQcBuuov+52ifOOQCRSZ2UZvO5LEguQr/
+2FIOTeN9JMiqCzdHkmW07NhlfPKH5T42NyFVL42dr/XYWheoKqlxaP6gILKqtCjfu7E80eiZYX7
B738gGgeY25kKsee3jg2zxPmPBF6RHNXQ4rGtuuhB2HT7ccWkAEUrJk/Cw7q+SgE+4v+kPtzInNO
HteZ9GnVioN9SGrqQRIf1QB5cmmxLe0aaS7B9elcLqY/2m4t9aY93cOWMc6AbLBh+PRtPExC6nTP
vEwytJlKcoh36A8kIiDZajZMbkZCCmTr+yHjhvwzmczigkqWshJ4t/cRoYgTB0b3z5LPr0AdxHyj
SBCAESAZhMH4q4xadCwbLpEhL1pOOQOna5bu+ViGzSiRk2ZyBeeR9uLU6LMdPu6Y7GOIRstgAQhP
phkbkkmVHxAKccIO1H54qJHwoETVDZeXjJmGNmb1EjIZ+kN3w9riV+5cctEsWU7AgKo00pGBz7Zr
msXDmtMrj/f6p1O4nioNEY1dUfxv5GyzCDCdcyQJyhuRze57mAf3pqoOJrue52gTDYVKYpbtsM0D
kFEEatozFAcS+GTOJ6xzKQF29iakbH6hpnn6MRcvR+8FvbNB9k7sV3C9linachP2iHSW2Mc06sJ9
T37cGtG6s+RC9XsabjSTJ/PPvSvdM0NGYIsMZQLHZdWELb3+DH0tARjHmhl2LoPxmndzkcbfyTS1
TnpE3bICqAlLcKOvr3S2OBE8VE2KVqyzEi9Kdq2rQLMCwFgIQWv313CIQbJaL/UjA85I0YFtoARu
JXCxc3BGhvd4J8j/nEpxzecgIbMvAq8EsDEY6hw3KaaUnJiHGbJL71kSNah9EkXI51JOtTlcWUa6
A0v+mIrhbdSMuRQhaz7XaYEvpLjTy5gDE3+lELBnzitSW67d7oSEIduwIz7DZetmtnUF6XdGv7Gi
IvsCPCGSU1duG79uL0VeN5tSJP+A3swtITzj++CtFO5bJ24X2SgCvP8m5F/B7wITAPqFML9TCkCd
PaOtv8JOXcLs8z8MXxnDUiK3AjYJrHU/6scalc0NBozwwG3XE9eNi5hsKYgrTWtuZa0i4gHJLw7Y
hFWS7d/8ZDBAL0RqrwZGbVr7Vp8uVYfn9lvJ8hLK4Wn1C1d7oj0BjfIma4asch4PBFwRukjoB1CM
2s4irX936TCVWOXkpsHOnBmgmeS3ZUGxVcEd567RtPYLsWlnQWdeH6QAQrQB1DN84tiP94az0/g8
Uwcf9it/SgJp2HnbzTiVsP5TjVNqsF7MP9GxHD8dctX4ur9jHclht/hWhIrNcgsGvcIVDB+BVu7i
7Wx1PxJvyXw8QZUpmh3VY8ociMZ78jllulMkVdBO26HSFrKf3icGUOLxTCwguVqBVsgAdjBuVVuu
jVHtNHRWq7UdmAn3w0TGwkl7ZRSrUKS7VhdybtWG3a7o5C/4jW+208McLhWxkPAZy9+2UmWIxRln
P9WyGQLehU6mkvf11jxnEptDzMGN8t1uiOhH7fhgyKIS3VUlJ+wTXuc348hRnBWcPIZCmEaVd2Tj
KZN6/LmH8jNheIl9LxfIvkT10gDF/jhagA4kgcWcOT168gp8/jS27my76+sj/eByr30BtCPQ4GWE
WIKWrXrN3AgwRWMgDyOGmpikkyVQEp8waw4I006myXr7j4TwB7XKMiq8WL4lsD2xVfi/DD7KKeF0
uUDf7allGo+myj8WLABMC3QCpAcoFoHr0kWyVBZw3WRcjOr9csCnFzjjp0gBQE9Q4O/X2+IpxNGL
RWMdx7Xy9jtxTIlR5TLpjXQd5Z3ttuX0TEldKZsoKhF8rdYiT5bHzZmlrsnzn6OPj6wMJscbKdcn
67PQm4k5EcqmPXHzsGg+PoQ1WqrtYBNC8fZNN/Y2kBTvAE4DhSnhONXIEEoW9KYTxA1EFBVPHRrR
aHiVCs+prMTwjrp17HBQYAsiXp9TxGCg98caCi3Ty37Xd19xzp6V6se4eClwUMjyT5DRaiuvF23s
H2h+pDovcCGkkeGGH4UQ0dL6ze8WUYoQfGXY54xPlLHorSfnukdesa+ZRWyqWZ+F1ytvGynGj/bS
AqvJa9+0bkahI17trSbXY+XuX/eay/aiZgpBiHlbu1xgwVROeKNIvjJUZoSq7DqdK73hygLVdGx7
LjynDwJFKToSx3u0/E1x9dwIt9og7r8/3d/HX7zleyuZQSFTM7g5UOhX55zxKaQSBwf7JcyDYugU
LxVqyu2lQ2x2Dc2RU1PnC4PA64H6ltSs7kbvxaHxbEV7cn1ixVyr9+E18Z1rkHTdIfyFdetKIHeL
+oP9SuDG3RwTDgTZO4vuGHpr8Molq8lRQ+0V021OiCtKFgChhU5a7t6apPqQrDQEfhLgZsIiTm/w
+s/4XeaAA+4ihSq4hijg0kBEPSEjeHgWWAQN9oDrdEu4WIYQJJrAiQaUwxo2REyMte1kGMUONU0T
+bokVh7rDZjW5Pb9QvxhKq1HohfpwIH+onYfO0ony7rKc7WKJt4L/y+uYd3FSoNdIXpc18iQP+Zn
C9IgipfeuX4RZgBRBFh7RDbSXNmL3ObkKl/Yd9gmZ9BAlWLhm+h60S8me8eK1qyqeZQJvl73KATi
h5R0b5wbB792FEIR1PGWEReRCqSYi7qoIlyxC+2X3ZS55FUz2sJLGUz2JlxI1FxnwVeqpyHfl+vr
sM1Qk5/vXT9dhUwotmZrV3YIBf8BX1NwY5WuH8DXDbUmGz3rDhQkAoHzWp1ICudwwVAiTEkQlSVb
EUOxj8WYxsbOj90XNQPzDpPm2oHxKklUg4pWYkqz20tGT8zobqqvqxf1URgkStsi42jJD/k7mU9p
f8WBY+7UEPqfVfcVU6AiqHnKMO3qQPq5pYK1NSLg1b1V7pHSLpRHaLM5+YsLB/cQOzrad/ENZ25K
eJGHMg1ugIFI/EJKJBnjbdQ3byVAU0BCQYWehJ6zZMuvSf5lHao09aDu9WjJyhHboXSnEFgGeSag
YhmLoxxIJ+Ofd4JY4YPQ/Om6cCcwvqv2j4DRKG8/48a3lIWWEZtN1h8cbjf/3WYIn2jN9lUfj3Dg
RJleyBxH0DTYBfLQXBkkBP/rRX6O5GmIpQoZH7TsdkpHMAGKOjjApZYVyTaehUw58BuUhoeot6O+
/aYm9qFz2QOqPr24BbjJrWdnJwlQ/ZyKhkmHB95b/g0UGPmm7cBc9GWE44fF434j9a1kC+VFjZrH
IQKAFTbW29BaV/fsdUcxVHAOgG2NB8m7JIToJG00ACm9LV4K30Cjh8dd3zS/oDgDuuWhoTncU4oC
C2XpVNeBAwJlo8ITmTa3q1/CCvosnw01gmIWkJlvU7hS+3lvbpQGTUOqLntTeGyWFM87RC80jjKm
TvEMalYErYJ6rjARMi+Mdt6sRRX3OfqM3gv2yWP7znlhf+k6eYfoZW2igckeBZzt2SLuHJois3Qd
vSRTPAHEOGK00VrbayoOS39GNOByLuSxWhXmPembddlF89sPnhMoX1KsoPgVESF4OGzM+IMbTowr
3YqITvB+NLQqYSg6Vxvw7tqbMlxKAPjBOpL/7tcM88nqQWo256u0BAiUAcR4Q0gP9Skzih5h5KhT
hms0SF5BQ0a231R/9MuYfPSvEDW5bs/vzyh1jdHQwC/raO30S4LS0IyYOQS/mdp6BBtnx75hjsE6
z1lrizU45NGBE4NEH2RzsJxNYop0ru3ECW8v4+ZqOcQWsaVuCTrb0UFJNhWNtJL2+zV29+fQauhp
N1B/lzdPhp/lmwa6HoJR6gmsGeSELOI5PVQx0EDSJ8cCZYWjrasfM1PyYMEzFu3Pg/mI0sCjJCjd
l1Rij/1SOPkseRchBY3aWql2PmpzJ+AlgrYnp6DGpvr3YKKWKIRFQx1a/iaAGKUU3c7jjjgax2SD
Rv6q4Bx4AvJGDcWC5rAmcXw4eJsyLhhmQs+/eZTI/vtSXtI4lRUCf7bWNAiArO1cRcIYCZS9rhG+
zR/N0ZxjaBNs3ctgeRkOgRKKZvudmjX9ZctD3pPAE0hTLbkiu/IRJ5woDqh1unZJt8ptYx7NUnmK
HuZk8G4OAE6QuKTVOxAQVMk8uqsTZw29K9ntP9yebzkBrGqQR1S7IQGoKLuSRjIckGE5IQQlHJAc
nXU+M/0mqXiID/+pz27cpgoobqky+aNLWBGBXti2RxUYAwM90x6c03QNn9UfSOaV8eTIs8usjc5l
lZ9PLsGAPHr7WxLWLxc5N9ukwCSBSvJ9YloAUYr/fGoEC2lrSVkA7JOqAKQwZu9v+7vKa0CYMkdL
htVR3lSn2aDQ2yXxS0qfWDkI1BUGae4Kf99cwACMV7r5vSsBB8cWrf7rgeFmkHdUaE0tpcMEpd1Z
r4tBbdTe9/W4KxwIdDmh6p0hDE/dT681g3MOfoYx6Ee62ZznJaDTnsZ10AiU4DGhfLfhAwqV21SF
nDH13kbX65yqsUHnSJl4x+a1TcgIuFLUUImCu+D6qcAft8Ql5z3uJZDRC/phlwcWvw0vR1PPssPw
zhmIXzb4duDKeiisI+IMkPyBm/pYLfQY+wCL+zgAW2+BXt4rQEe4CSGCmy9neklsdZdHMaJBbikc
m8jTFwHb1N5UZxK+brsUR/w9FOL0ti3gJoHqx7S0fYtZ8BfJiUCZrDrapGd3LA+5YuXja/qgssy3
HQ7I2Ukd4ZgCHG9/VREbrOq8amJ6KhgsZHMPrGQsBXr8alO4/13d5S8KqLG7RYL9ygryE7s8I+Qv
x+MhMRZQV3PPDLqjfaaV6d1b7nKxOTE3tcZOvYzxsoraMVILzKiPpL2JYEwDAtHGRjqt7gfS4WQZ
sxaSCYO90eX3ZoNS84cN/7cYUY9ynkaFiuCsMXHX7nzeSAJ3yZ03F9bCWA7uYxEOsiB6MI0Pm2S9
zWwPaRJibPVGvpHx+MhwXem1e8YyZaTY+hoNXoAmIFl8wiOuoMT6wsnBBbMlKaZXfDGXrm1+I1hx
+unbKogdisNpVttIxxxkdmS1lB1D4aJ5CLIE04EfSkg/rgH3MHYuoD8i0SlynOCdF8knUacgJTsh
WuwaYRabSQnUEibkJ8//2KkfJdAMLDly5m7r5irmynDIW0yUq01z+m96W14vhsiy/XyWZV0XB6FP
JA9CVrXtHmMyzJKXsqHXMG35q/A7Bpfheb4cQ8t1rjS5iU3BNNk4i/7QnC3yA/j0OMlZsq9kibuT
SSZU5CyU83l4VzhZDX/wz2cK+vwD9/cx07vT+NqfyxQ/0g1rqwEcrYrLrBbGmmiC5WOinEK7gXAD
mymM8j3UrbSHn+aQRs/6adpaGl483iZcRYGB0wpvrg5pCCOnIhgV6Qrm+vhfjceO2dLOJtojHXr0
+8LbAfCFg1rkSZkdeu/9wxdPloVrdtAAANj4xPYC6xoRdyABFDLP2gi7tI/RvMp2heV23YBmx2uN
t+oPobP33iDUzhH5wdlSGmFtADtB6maz/1Az+XYw2HIq0jqAQ4BaWvPiJXDryMkvBJf+CsrcHKvP
9BuY7VtazkPA0xDmq03XtrSbKj2rx+xQKb45ZOAO0bNjKZ/EkcEGPjFcL7kA3PsCdkkXIEShfNwR
1q9/9jBFxBk33w4T/QV+CWJLvJzZJ+4Cs1LtHLrDomxhz6eABJnhbY5++Pr7/aqrn7wTpD8GorQM
Qj5Tn8RaMLpVuOnTRRzbPWr7yZnams7u4CrtGIGS28jQHn8vXND1aGOA+R3zuSYPrKwnWBH5NmxK
Xmrq+eI6shwaAXNBhK77RRMkrKd6Xfd1CxasfpPjAu4/0pXwoHUz54sVnbXxRYl4Q2DnRe1CgCfK
YK9r4XUQBH8nxsovY/YSK1RgSaWuLoALV+x3P2VVENL7XoKeE9xVV26JdaQkngnhgrIVUVrQMlHP
ShbonCVHdLlxwi084kd0qaHIu3c3EVydvaHPeMuJ453XtsiNIbL4KHcUbHDcWo8bb6chWKN+OQ3W
6MbUlpZ1WgJ7TSIRonULM2CvxNo9XG5fkxN8/eUa3IfLELwA6TR+0ik/dnK/EZIYeGivFQzu3krg
yu5A3ES4hrTe1CYTbdT10OE16ia6j9HyG4V/Lsc5oxp2j9ReC9qzi8ZD14WnK02Sb8EQpT5HhSvI
WdHM8n9BslOJthdOoHGaz7wpvBK+D3Q9WYIYci29jmzH9rakNWJLgjiLAVF6Wzs007oVdKaKJmbg
sKRZ+pVRnjkdRCSq5mfWZsvd9NYKSrvr/TMM9/dRZLlWY8ENRuu9h5HnulP6hvEQo5Zr/mQH8cep
tnMxTekTrGcVhdISmg+CmYTskCm8WyNbS4YqiU64rv/zS0hIvxda4ufOrx/yHTrylhRKgd+BGs6D
iufomNJJR0uC2agZdE+kz7abHTFpVkvGw+cWP2I5hZoQ+V1u8OCZm/tb2sizbUQexSE+cb0Dy9SZ
DuCfQSgASHo3p3vWcx8sGGXTfI77SH2OP93fm3LTuu09BBWnXdW1z2A/JzgDC12+7VWlFEbM0aKU
borg0JIumhuhuea1go4ELAmwAbKRcbb7ORqTCp24ciJyLK+n7TWjRraV7OXyqZw2KHJ2oF72Rfbu
r2WxaoK3vLxaFZF9alY/OvKVQQycmqGwPF3Nu2KXQx2J4nnvm1hdJFYkyWkKJphmKPC6d5NvwEoA
ytKYaz2ar6H/CCEcdWFF2i/E6pcL6yV40OlSQ7f0DGCciXf+LNrqHXXnwGLlV5gJ6jFQ22lpXfTZ
19q9rhF3PpKr/efSP+iOmqx6nk6oo7wMBDCgyG03IzKpC4pgnvZqKxtY+EpOtPrDmsWmlDuwnZVg
wdT1bERRfB0kFXg64fzvql7HbSvWZRBgwQiBUwnboDKTBIBxYV3FDh9+/8FL0IWL7R+vsOtRkdRn
WLfngAMO40abY2zJr0qN3r5IXgSFhN7/hYtYTrsvn3kSvPEFpob8Z4Xi02VzhF0IK+XzTDKmbWMC
vOHsrTCi6kpHaFc3RxyhysbnckmO8ADdxp08XrE7abOZqoa8TxrSuFc6pKbh2MWBisGBfW+JRAzw
wpWXavAM+OG4p7C4ZDgqu+pVQgiYFw8qeuup0e5n87nl16ArmuEaEsBDLE3pLkXnUI89AsJg0ENu
YF2b3CrQIBaEv17ya6JU8E64ePMhD/9Hkf9Z58tQW/I4VF8IruafLXFNKnPC9rY+fTRofvoqeCaH
I1uXYf3Ah4YLsDnOoBWeH+VlBezp7jtgVznq8je/vN3pxTl+K8aWIBbIj10ANkUd44JIe6Hv9nLY
bqPpL1yYz4vzlrfMCAV915NHXEPt/e9I7cMHObGwkzoNyQZeqVyVt2F9TjJgbi1pNCskSzAKhQ3T
lWX2mhsW5Snc5spBYgAJ92fNlzzi1/f0TlDrBq3hupGjYw7/zT85VHSLRZbhkUxlDODk8ecavU4o
Osw9BwYgK+4nkNSz1w+79Fc1ejnyhj2XLR7W27bkZO6WqL2VIHeZZ2LiYFft73z5wKoYfDgplUri
oANvrb3oSvek6A5QsIMQcZAPuUXE8qKTxygQ+E38w9E7HsDqkAIzsnZ35Ie3+T1W6l10DgRcb/hH
oNZjiflhCu3UAEpWknwksiYIERpM6GGcxwuyzdYPDBZPA8mskOxwu/hynbguuLdl40S7T2vWvdKf
9SOK+5Bpj/D6F69CeNlYyJj7xHtHagDeMY0Kxc8gzEOgY22tsGuRCRI8hvDecCeItCV1cc9j0e4y
jAOL7wYrDDsmmEcHhxZ3yrjodNzDcvjcgwVjCa47+uuQ5YKsYmPfDY9QRYHtlp2kP4W0kPSwCBZr
+hLr6HQWnSpXwtyLGIs0uD0Bp8O4yBmAge9dXfGsEK2l+tveY0prFwCh82rrBJmxeQSn3VpI1cIb
1h+umlhC2eX+OvhKptkpLV92P4vYR5EoEnYO+imDfMp9zkvTm7umcHMetRMzcv2GSLocKdjOmyql
T9rymVmnawZOYJtaBl39h/hUllZbDVcKPJ/tfZ7I5jx7j96ylMQZMG8RTW6u0gfPSFY4zbeQHC4b
BQOTAB3nEkoocnl5iP9/5Q2PNDZJpPpOBvD7YhVPVUCD5irEpVJZKVkS8je84GM0eGWSSCVepykS
v0J8fbZrc4P5t+YCGYqcEHrcV9sCf3a8malheMw7g6dO73MAoP1774dwzmUkqkNZQNVT5SWTBGHH
2D92sRK8wLNXWKf+1MaZysMsTz+duWkIgXPLPtG7dQ7+lvX1Y3cX6Bdt5RE6gjVPzRVa5sGHgKTx
EeLWfT7IWztmUuDv0315QYThItBkwjMwXoHFA0sw+sEm9vWco9WMhHuqykLxntYra4jNR7YUOLIW
TBdACGtg6JF2fBWAivS+jx/RDQg2dYeIdzw7JpiRdCHNakPufxPXPURHsumoFoBnNK9FE1q3k0Al
3MA9c+085kHymTnFF6myweheKGLO8XbKPkLaXB/0k4k+dwkPah8NPPaRAV4i0Uw5dLIkjJH1m60K
sMzCWAx2mvFsNIG3Ys6niZqGaaN+94o/AchfJduZafj1DmB9HJxogvo7LgjKr8CLvtxn4RfRcjgw
Heo/gBp5mP4bL9qZCOG808o9gCTcllg9wmwhqtF1UafguUWtkU/1I/c+57llKadgpbq7Gk2vtAmf
FJs7VRn8OLJ2C9XJex6G7Ix7J1T8aKRv2veQYQu31I+W6YFv68hMwU3ymK5qKmBFCaAu39EyS7JP
L433AQPYB/XTqoOBmLlvgEH0xq1D5Ln3OxHrnwb+VGPXB3ZJ8AHFrh6DGGOp5iJtMecxXN4TWLu8
62+2xmXy8Ub01gmCCb9+ERQ2N/ncnYMe4D3tarNREbMtgtPD3A0/CmfWyHKPDnKaEhC200Xw3Vz+
DPBwXTF7VOh53jmFUhDf/NwwlRujHHGZMljqZiZFh3eE344yCY16+qX0bieIZedH8jr6yl4L+87N
YErCVox6myYe1u9d1luk3WQzchWw83keCLzTFfk3avPzFgizVhZbfaFkfhYNwkq0uyLHUvzHdK1D
Y8iTHxoXFa9FPxrUvx+9ydHRv+6Bv71UaMnkVvaerMM6VkRnQQYQE0F9PY12WFP90oWHX3YzjyMs
KaXi3Tj/HEXGnhto/lQKky1Ot/Y2AkIGbIBuKS5/g2WLaZnadc5B1Nyxeah7JgOF8CMaLuknOOTV
4CINMiHksdKSFVGlnebR0ZAIDFSF0dfl3X+Iyi41Y7oRFMryOMNGQLEc0lfXCN4JenaPg0BqyDP3
dmJwoURzxeWFryoOE7oIhBnd7C9EK8m8UzXyhtqz0qSmycoB7KfU3guOssHgaPeAsCD94fe2+j75
K7hU8PULbpM14a/3m06+Up5zt+BdlRBi77fRsG8Qyk/A7HMcSUJTztSa8Ti3OSO/L1W1n5n+stmp
d4e9nzKGgj7W5QTwq8QSEjL96FHy1+LVK7uStMeun3cJKSaKG+nbabZwAWK8ZtzJsQLauN1qpjrX
avRR5vcghkhSO74FGH7sSc9+y/IMX2Qdb5E5JBhTGwbXrGvZYcRJlt/hKFVlQXeQuZr1/pxVgECu
HLcZ46q+D4qG2bF2qGN91q0nwK9GksbObsdPn/cbBOO2IkDa6ohhCHY6xukrgZxE+q3YUJJJHyqP
0mfdznt6IyhqNrskP/26g8fJ1bcs/3ip6QwP6O8I28wX7oTOPEriyE+Soy8KmnaZCl8EU3Ez7Khy
Nq4yBCe+MtLJgZ5vbq0IWTcXKnRhdBfHA9RsmhEooII0vAotWwMWNYN08BFuLuiKKKYq6bOd2dpx
g+5PpUGy0HMNvrWJ6LJ87B1+r1IJZ7Z5iQOhMcDTD0bDZ8/rJz5mrpdLMEmfeF/X+SwpAwTsxDYC
Zkoe+saAXbwQVTOuuYrnIbjh5SMyulsNXHtw582V+KNrKPAntr2FHIL3jgYjdNDC30wJOS4jENtQ
oApDEGJ0DmH2CrWZ2qpd/jZ3I9DvAYH/EIfqpI0YiofrACgC2yYu4nNfx8wdVbp0RqFrFeXKw7Xi
3WdcOx1IsAjQ/Y40UU2U26A8GavvURfl8ybcJ2e75NNfjsoAJzWqJB6fFLTfJFw3MXv4Bc6BMJu7
2hUlrA8sb7xU1JD4U1Aar1PF8YAlrbvYfjS0TactdireEOJ4fyx9ouOPAQqdKilut+c+N6zY/Aq4
43XFdT5mt6PzqTe6yKt/HC77PfoYImaZtGFc9rJhVdgqhaZ8pf8jvz94PNG3Gg6KNzGJ5YQK6yqD
5fy8bKMssHaiU31Dmmc3AFUqr9fqL4B16RaA+x82mp5XqtmpmvCLCJ2ONUQzGpZ6rHD4lWRofpqg
Hk6e2+aipVyyBQTlTP94tKjx/ijTWio79HI7YLQrhR5p84uKERlWZC/ZkSXJzA2flUUWFZ/KRC/t
YDavM0eaFgj8v7b42PS8SwIkQ2I22bJyB9R8HFbxH1OkutSDNRAsqBGAGjWJrIDFQIN5r8zepqpR
d9zwV3xKrobILcUaEMYtENdIWGGrtiKHTQhADw9P/8VSFCFLQsFQg9VmFwdSyjH0KBKnP9oR52Ga
yQ6FNPj8YYLeWg9pP69AoGUQ48+YJC3HTuHMQkm3Ke5S0G7uYM1H0nCoo0Xqk4QvhsPRd+uOenj7
MG3QpHPRVGmwPRcdKniNU+r5n9SJvvbq/ECfXKwMEc5XIzW2k7CDKnoPTd9uGkQuq1U+Q32FLKfr
1zG1+GsFWrYIDiTjVPjRpKtE8hSR99n2Sixx4uhu5gSjWleKsE2MCsomUzqWFMdN0VTUWDBeSzRT
b6MVu94OxIWONafzeWMye7nlO36s2NDp3lnRRBn+TdNSckOL2A1f53/rj4MmOgWO8aGqlms/hvYr
zon9p36Y8SOCsqqRbfqdny2ZhMziyj8PwKdI+bi//w0jX56U025L2tox1kP3H01z0qUvIIKhPSrC
2vVdf2IHZOc8Qb9qlii6Q2YOs064c1ykJ9i6ofwu54+ySyalkqBROZSAwJ3v9VxJpkI3JNTkFZYK
5QeLkCUrlIZqqNcmcJKEHInbYcB7cht1g1InjMsAYrWKBsuFY9rZHDH7XZfEyQ7EIvbt7cxBivNr
knTjuyoUMOaCO/jAmdu65vHBPPKUduerrkysB5+YCCtZiof7fDHq+XN0MDM20hO3h96CBejWr4Vw
i+1J0xh5Y2wmIQyfycuFcvvShWOZbIC9xtDQvDNoUU3pbJZWMZ/mbQ+Th4vfj9xBkD5KWxYPWuVf
+fwEdo2Gf+Adxpcbcb4h/f5QIFLQGFsWKM1ppb8/vJZaz36Vz2cHBfZin3btqofOjybjFvmbc2lU
MNPT8qYPLqOhMpDfapbg4hK7AQeWzUXYg7RHawmCSfQLwSYxrMNn0erIlGDQM5sQ6exWX1Rr/vGQ
BNNzJRIs/bv6aMe5xCSd5I3sDZ0vKhMIG9e02XTskmxnxrY8iBOPCFPaQMrIxSEU7MhsjnH3J60Q
FBEfkk3t2zhDYEJLh2F78XHA2Xjb2K8qlNxNZSHVX39kWFFNWLX/Ib2Ri1vhi0kvDA7xzDERnaTy
/ggOFyw+uLD4jDJmukhyh9cqBDNJs60q2Ar3krcZHAsdU7PAeR3XSfGHf/LUqRGEm6IOptg4pfM8
tk3aiMdAylKW3BaMDg5dep13gmDuOsNkSsnGussDonUFQrD0YFbSY5mx4EnSMZn2iKj7JkG86Eqc
FPTcoOSDe7VqoFQWTaIOijNTYBXZQyW6tGZWuMS2A40NicJBcA/Ip/lRDWxsgKD2AjP+tuq9XyCb
WCJZr1KYsNe+jUX+WhErz6pv5gipSPGDrlbbJZ5JH/7m/SGBMui8U3+oHVHRZr9U0BzjDOPJ5Lbp
t3VnlJo2qiO0RvmYbOkc5OR6Hl3nP31HiCY4IB13OUKGdyz+kaorGxkhAZYcjuFXGFn0O/RApkAW
E2Y8qdA4ZockWmzDSuF1sH0xpLgXLT0roW2jdMXhKLJeoR6tF/nFl/E8WrJ0NZIq0O1SuLdhK9hG
QgiKcO8GSa5HMHQgXeeyI3XV3GgCIDMCzEGFveGUJoAMqWM5pGJfUNFNbm4gJ8eQdP4m3YjYODvJ
HPdgbFuFF7AbN2Qo4chWg99yOu+7n2MJBoZrWWI+TAKkDQqgY4SK/CUUGcP2VXmuoPHk0m0i0RdH
MhGYjGr+eNFf6omP6x2IWNHej/wfmnNcKZXbc9fy5b9l83UkluYVbvNxVNOBpupq/wr8XFZz4B+Y
X+gbwigqKZFw9PubjVK1K75R8gIL2jidzY6XAiie4w6+7RYiP84Wqh3DIklmJFldYGkphH5w0VGK
Say23+K6/PThfS23cFd8pI/nFxeWJpYH4EM+J3EZAEBN7DLsbxBPM3iKIYvXSLUUJLXcRfYrd37P
73fYfSEoxUY0xZr+7oqMQ8UjVOdTKulXEmO7oZMf7Z5Nh3K8MI51U851sA97Cajdt8GwIHlUp3GH
5tsjqOpmBBxKU02Bdkbme6Cgzbe9u/AjeyrIcq7bgXyM4vO308qeS0ypDEZnZM5M8GPli7ZUYIy9
Yni0BTAJtZbJj/9LP0ods8FTLH2c1uUjLSFXl4Y4bXjZRe+83jF4g5/+pyi5NOJSQWplTD9DS27P
ny1O0SBA9JN0A92IxNtPwci4JP4WUwZJqkL4inTVmFSQs1vl/jKSwR9/dPVQG1OQoeRliAomQUNe
Vf71+iX2ixys9K6UddFSL+I1qEcYufdGfQSvkPkDzTkCnwNN5Ky8gxjHAlS9tf1lkt5tKWrT0sNR
ueKC1pDV0LdS7SikrKT+XOrGwq8cZqH7ddIQqtAb46diw7vJUHidCoTMJtMF4/Tw397CCryBJ/L2
cvRfTPluGHah9D/kC/1dGgzaM6hnrO4i8a3R7VIH2Z9n6KUn8Il0K97hRuX/1mt8HUCdvVv+AC5r
rCXnGe0kAOSCnHXaWnqOxLd4RkU+s1VVrNOgZMdc28BIGOyv0GZEVN4L/fZpKtd6Xr4Qn9HikHwC
m0RzSAHOe67AZ+RmyT3e1u0ozIJW4m86NEtXNOvDuLtXOAWHdirVE0o5ZpqutZqpAVPf2h2t4vFq
cOb+s/5e4nMfmpxtLC1GqqZreDKp7S5r9mLI7mtnDf6zNYJPPs/99D5JgyN6Npuu8+9K61I/9gfh
pz30pTirUOQ4r0WhF0xOdrbFI3HlsYCH0r8upDfr/sIlP94yZItuZzaf05O61ThPEMm++9GOCZj9
SSOaVKd2sCGd1OVtpsAzTlJU/8IvLGf041Hl6spBygsIq4G3r+mlnICrwS7rwQOHIYqek4/Hri42
wyygoowVJThn05OxYqKO6oU8VhyRxcQLhtJYqkS/iaSbEHYjQ//y6A/MqQ/QptDju7FfIsPeDi9x
UAvPb+UfcyUKFVy3zjkcGa0f8RSCZKPLV8vBSGsqs1ATZXELOeXWFyMTgDagytARQHqSjYM+fmkh
8mXIQigF887Zxdqn73lHOt9A9M1+XX1G66HWAKJHJMOdfRmHLOgqgIpxjQQAwbzDEMEbWOgt6Dej
BEsMKa+p/eNUYu7JZV0otgvFjRQ4Kxrb3LScKyz8cRoGodcSrVdakG1Z875KvDgzy1u+bYGaYG/0
Iiz5ox83WCWudaSl9Y6aSsPXKyBHEBXG4XXb38sO+dViwSxAvK0SFqBqzR64tuLe/+ntc3gA9hqo
ukSq7/L8/eHYKZObm/37x3IHCf7wyFRU4cirfradC9Ws/9iCG6aa9jY0I1sWafuddichuTKrWsOj
Lwyzu2NEJwqTGLF2vhl06YTVhAQ0AeFHeyo6XUCxBrXd/edVtE+VbATCaCDXLqnYHQdGVRtSnJuQ
ZDxcNLt54dehaIdmq+MGreCmnWkSspQGRT55vqYBEgh6pIbJm5qWBO56GE/SwEsxwSzTn3eGhpin
8UxPMi/cSoYH91L8MfibiOoe6MwyDTzIYmLxvDRcRzEG8N3uDX4WNjfSNpJ2o97lwbt/wil/Aia7
aBuB459/fNSinjF1L1EVWyXEtUJR02mTy17UU6S1+V00IMI1LN3ASJzyaOp4iftP8wUNmQH/LiiB
j1ejFgjumXzp0GBabCIJ+tWoOwd3QQ+89IfTl5rZr7quOffnAId+lg+tS2FuAoGi941fTZxUuc/i
szZ9pbH0ixocPRUVzpIcj+06DJ790HYwD5e1dikXDGVB2EirmhsErIv4XJKsn6EIgyEo4w0tymUN
OlD8jW6szkFiwmADp0/dzYl8qSC92dnz/ebMJHlTnlBHOiv2qqyegcENhmbBdC2GqJZKgBvHcMhx
0Eb76eQV84r0Qcs6D3fUFbQoY+fcB7VlOcwgm7+7Hqj817mXuG9BI8waW+1CkpccZbVeTBo5yppS
/c7VTyl3K3vEDxs+dFFbSF3lAcGfEG0jUe1JVVWBt8GEyY4x9VITsEAbN+SZ9jGuEfbRNg9fkDR4
lxTKOG5JxJ9LQtVF08rUMewDTfWLshtXDQlMOXZ7/fwXz89k0A0Ft3CRnbGTd21R9QREk2sI+ouq
UQtlO67HsecksYfZO6pZNDNKtQYQqHNurclaJaWERgxZiXVYCGYnyPBr3XKCMQw5DZhwNYv6qaSZ
uYnlRNuz302yQuJgJqx1ZG4LSLL+sn8hYGkUBRnyxZtUJMgnq3S8X01M8pH/QkwvYn//43JeyBxv
Eg+N1C1QTwLdjLNqf0WgdnOniaA28wv5h4WkMsSN1Pa6Wiv3ihvLellTEnQwW0PPonzkV0T9stR/
+0GEITIPYc5nY0O7MLgAdbPmCYDlP7D7+OiZXPuY0EhwKJ2zd293sjdneh3j4Z3Dr/MQuzEP1drq
mBL7uchICmqbMW1Ohzc3Blsvh/1qjEIJa3QX1xZlOooXoTnVgCsFyy7VHBrakwW6Vs9JH9u9ORM6
a//U3ALJn+hZYlrePzetGh8w2xi/i//wTf3fVO8wVcQohuMufRDZDzbhUAaoocqQAhj0NgOFNgcj
rFFgGnJeI+HA7KXYcbGgGYPQdYenWNFdvDOsWELPww5u9XBvzQyfL9P95/yr/bVl6jjdkDfeQ46X
i5lKOBAz7NzrX7R4K11Ns0TtZUiw5RsF7uErDCrd4QzRysPSi54K3icdAvpD0n/wl/XlLr0Z+Om3
gp4gNHBztAPN39nqRKI7iJiaZ6exWrlMrI7w+zCBqcuNIuodFXWlJVfbr3YPpUtktuvVRgB4Pwh7
eylcjCl+HFJt0E90lcdy0FBmh9FIBL/sI9RGhiYEe5CkZ3w6LTASMaO9LY2YpzdN1YB/bU/bHYIy
DrQExJsK469XwTPEPbIsVxMUUe24TUY7ZMBbWT1rAfCUBHma/O4LTpWNlHNU2XkS9OLqW79UhQDl
J1K2A3BqXz7fokh7AXHzVNr3uBpwpr2CjB3yurQtr7cb+BCIJqlGpEd+Dq+DTGSBlzIhbW3wXUBP
N4CedBeomzZ7ykE45OIVo36dhjgsgSzr/rmwxdkzsS/U/NI6V0CHFvjbVdLfbfziQV5g6l2COSS+
vl/pyt+ZHP8QJckFhGT/G70pHexgi5wwk/glBHtYK8ihbewufcxFUPFzyx8kwge/ZNmUflPXmcoZ
qsoWYsKT+8tWrUkTlPJ56jGGS44oGjsrsvM6alM9xWEo/En+B85ks13gm1apdZ4gGrcELwjpvVsk
dyqtl9ZS3y9yDglkON8Kz3Men5F5anO0X6DUlC8rgzA0SReTTNzA9KWKrXcXiG5A8Azhvxqhd2C/
FlCJmwJy+r8ShwjogRn8IGLqHiK25fauRLIgMLnvqskt2KMBdFXJEzEpegiWhs6YXGpzv0D35pKh
aleY34DmzX2o02X/CukbovqBrhIZr17ue6Y9wweyltYFYbDfN/tv+K0FfTQlaBjqIqN7wOG6z70u
D2FAGp1U0S58WOx2quPcruJxoFE6QlAFn0gbDmzCwbYEr9ChaGbI4P+VoxLKa1MJQt7PXRFDANih
KLOTXGBEvBVJJz677pzRZEsxhZD2j/S8fJTw1zn0xqST7XRUwx7d5eg1awjHv8JxJZYZlIBBI3Z7
TMp0EnMeL1g+0sX80aivI/tLtOAjU6xLsbL0BDf6jWadPGpxlh4VhwynQuDVBpYenidPTP41eA3U
m3p084FSOzpoupqLCfaQFoo+E3qZjQWOyBGuo7WH/xSXgle4DqMH7fH9VLDqyNDQ2OF4/Ql2kOuD
Ui7CgARhk+XiURCSK/eiX2wSBaT9UNKy+LE9DAAJa86TRDZMVx/OweeeTtNIXVUAQKxPv+Z369Ym
Hvqpp6sBWCC9yqzjRKrjVckeOZcHEwF8XwYvj/iSjxUmnuqb6jhIwzCiZk6XXX3iepu2+S/M7DrG
BFiFub4tDcKwd191LuqDGZeHwtVA50X6jVK51gUa3Cfb1nlIT586wQzCCvj+N46W+/ByotzLnYcE
wpaMpXCWvFABZBv2kMvMPv6VUv+Ze3UAZSl9A+ydYM40tOeJe+HRS4ytuSgZe3obRO/GDPs5T60W
KHIiSOgAmLoaxxY3BtHD4sAVWZDuzJ1BkalP1XB1D1Fz/hkKliMckaKZx6trEfJqax3PFWUTyIYz
Lw/4bA5Qqz7+rPDsUyNTJeJ2F3/dCiZIr4Wn2cTWMW6DLR17fgYmP3QXB4MfEZFrT9Ll0zPTdABd
ZQIdhVYeLuf5GFf3k3yKf5MZZWdz60gItV3eCGUijBZm+NzEj2kkeZQ5I/axkaZkKzrZvvgHT17L
XsuZqRq5az6nQ43dEiVLWmJ0eVwHor//5TEIvQex0HRNmiE8+TthLIiSOdlMMa7DlCZMhnntB1CZ
EJfbb5tKjYrAj5pvktMY/u17LpCpO7mxY1uRKgIau55f0HsnREK0DuVGR47bRChIipPl9coe8/og
/lxXkF6RYZtFlZTwyF98dsY0xjnGMcpF1Lng7nwDR2XOs00u3VlRCQJt3EF0LYAvDEx1QL2TiIkt
GQrGXZdGCqu3MNtPq065ccQq9+phXfFLSOWcXUcAx0hw8ji/yIz33wjRKQWUDHBz25x9UTG5xs4F
9dWcdi1SkQETF39/duUWqSCncFLR6UbFu33mciGk83gus0miX07E/c8v42at2byeXJAuF30sbQkz
Fi00V0kJuwxPVupVbGGlsbnMWmQamheucsqDojp2Br0CsIJBbtMs6T2jJXoXbVPjqbdedHGnDtuY
kf0F/i41nuLcApOLYxY/QZwUpI4M7/HYiYlop6j6LSGz6cF7HAlNXDPSVA1grJBAZm4aUP7/i261
weRA3lguo5527vvkaKr1Xp7QnYSTKRV1RnmJUA9lv/6dFBBNA0vYucS1FsaYb+Y+oxumIoEkj8EG
IET7A/YlSjEb6q45v++hwzMQ3uniYszuQ8GBvFcy3nx3kC/erQxPCOwFYVSS1cdaZCCBCPuX+8oT
/SMi09oTrKI39lg0La8vz3F9T7NFLat4WzePx8aamUd1awiW5RvkFbqeMTHox9a+Vlcl38L3X8J/
R7LbYeKuS9sCnhb/k+3VSTuqj6hsYvhpFZ/qkzBd/Knu0wEmT2LxkVm//fTvk6gd/kKMSh2+pm4f
Yvq4K0m8dd6RIiN2wHHNiF/4zV1TjIKexq+PHTAIaI1KzAWNGm0uG+kBIeh2jDbRha7VsVi0jZgK
5ABj4lTBsrcZ4TRlViVY6OcaRnA5Hm0qTyvabnFR/AwQ92UtpuSuQ3HddEZzucy9pdDnfQqvp9R/
Jm2Ni8iqgv1erynjLEfZi4/L/6ltpH8HVZE+gv8Vr8sqatet4uMslccCYf0vnAW840+mW2xvHLVz
brEnQKBvgMahygbrUNs/vxxA8XOd0DSIaA83DHfvk8ohNxFGqaXNAFdBBbrHRDo/gMBCvoxsAf0Y
dBITqpn7g/EY6x2my8UnY0seHiPsYtiR8L6vE47MOWH10IAFBoHg+kS0v9KC3BiIKCq+6hCCtBQ1
HB9n2mVwzRIH/yq7iQy5XPivdx02BwmNsO6ZdKOajQmj+TszYAV47L5ddIDcFCFF9oedmg2Bzzzy
R/oOuMYEBrKgW/yEp73JhKBjBuXHcqIhtfz0Ivf25m6hbuInJd3Ccmv22f90AgJNK50Hc/v8k3ZD
pWqg8OfND3IDxI2A0DNJUo9O4iiMierXVLS8lHw6AzB7NXka0mW4HMTGUnREPY/H8sLy+vP2nbCx
igUgkA4BS1BVv4nHtyMNzqtIC5B9Yk4EblLUt7sh2d8yZxyCz0ayodbrf2nHPJYYPt7VUGGF2q7j
NDbRa6YjmFbjSsScy4+3B4X6orq5U56YpWY7EJR8lqKbrlRiV63j45aMPAjmuLSFv1httam4xywm
7gmZJKN5uf51JKoMBl6DId4pCNUUJqrzeDyHXK1OvDUoaqj4/cqerQlKlg4ZrTb6T6ZUy3mt0YrR
aMSDgxfXcx22/vcqdJYavhYOyJI5MvPSoJu+wuTGqbxaXs6ywFe1r846z4GqmZee3MVHi/dg94En
bGFe+qC/e9nTfiqIpOjiSM/S4ywK0yJyfUnLrfqaFJBg43XSowjvlF38lrk1giUpUCTy5XQmZYs5
E3coCh64hxpXZUpnsDJP3zTsIDZmiB79wrrN6NMnJIqNBCfrPIrASKHkjGFMYx1nm0mzeQHgvOqA
Hhe/kRUsFudzS7AxKUG3HWh376yS4wqTchoWIk10exjas+t/35R2Ku2TpmR9f8d5BkwQ1Q8pcVMd
Qnl1cXY5/vgPg0e++nlZSegTsV0suEXjMLQAxhszC+NcZ4ziPMa4PMJhG0WuzGqWurJa1L/5RXz5
2UquKCTFPZURYDk8kEFWqosmkhJ5N2I6xeolVlMChFqoT2wnWKa/XZlD89O1dZCJMLTIwcL7d7qS
hJf3sVs07Wp3F9FozCUjbVrHGwn6ESc7M6FxM/0t2qxMtYF6wBfeOZzSmUV1vgMRPLFrm6DpFqVz
SuFEi3xhRFQ+gttaEMN8ZgJv511zVCTm3+f/qcsozFbnY86N/0mZLSGUWaUu80NmFSQxB8kAh+TH
lq6srWIcjbQwLs2d6KLxwKULFvFvZMzE20fMS9NUBQ+FSCIJltb8Xq+CQCGmWzxJfb76ndnvwTUz
oSVu0PcnZJA36i9k1ta8Jr+UJgi3ni/5w1CiR2QjKt1q7cVcO8wU0/+4rNNYQuH5Tx6dLyivSV/E
kO1l96Y3DSbjamJWhF49n5ePFFnoqzZioquRQeuKcpZdjRsFDAfoqDiEga/hBFhC6yuBslmidURl
SxJHe/cEak0kCqRDYLN3W3WsKuWf4IpPanKqZRlbRjfEbktSZcw0uWczbmJiLw1VPuP/OMH/Vqv1
XFYAKjkUUXJZQ0ZlPuqoLpNd6NRwxc/Qyl4cMo1tAL3H9XN+em+ip1hmfBhv8fGRK2g4XanVyphk
Z0KmaTNcTfA4fvZaJA4OifX9wNEJ+NYXFWDkAQPxK4ke8Fz5q42d31uBzjHVpC7BwisFG/GSHZI3
fWy1v72W0SvCW73trXDO2YU0Gwd/44O5+7vYoNg2QV4EYkWwduAHZlfN6ueG6VSBfoLrG4G83k8H
mGcj/5DJWiXnR0Poqj1BDiFK7wzweM52DRwnJw5+upssZ8wkBrASgimQetJBwEpHbmWbsIFq4cil
XvwDbwoAXmDnxoPQjw7ttotk9PtloAGCO1CKIZfHJ4HwjSwpKhOJC3ZydINLQXZ+pIAXgBwCdyTC
bSUqT5UyGd7GdIReqUxJ4VxBIVVHgF0HgzsobIhYnYsLXD3sr4ho9oFNPoQVomOQChj4dfe8AN3N
eAhCCv5LRcIMQ4r6riBsLPnr4sKWb/kc6yA9KFqIdwZhiIsDibeN8/4/S53qD97+70fHvYejTzLm
9Gai/3YRtcBb5iGbuRdRtThTTq07gA/TunV4I2DCBqMcXIU6b0ODQE6sz4u0IF2uCVREswjHd2kJ
PUPLDkX1D3ogbB3AC/eJ2o1Gqi74FghC73tfpKU1ndQbkUOsdNWyEzs3fACasSQu+j5I0wVgpJtE
qoomnzWTw7v9N2xNwgCYX+RjP1GBhbKOctCM01Xk6QIxuFQqBZq+BSNVah9VzYDmW/aydZ418r7p
z9hslR1e7MT1lw1ZBLjCGUA7DAw0a++ljmfsJvMk77bASuZ9geZ0Hacy64dU87BfP8OgbNFM/v6K
JQ3nSc8WR+RItsrKhvGrDr6p4cj+dStGq0LUq9EYdVns/WurvekoOsvc9VgWOvPBun4Z1aFiCSr8
eWsySST1P19wQQMays4VR4dDjIGLR7O+Ok2UaxwU76cklctTBUY7AdF05SXFTr3GsK2LPXQ7VlxL
lufc41J9wRB5RstNZMEcPdhhx/Zd8kUKgOpulIwc/88JVV32rlHPSFg7kJalPXfByUng0rRSU2Ym
v3w/jZhwDD2JCdouYHp7zMYupFbXre6HcTuwB1KgZmCiWOuXmOrNkK5db4rr7l+eLEmLZDkW8wh7
GOqM8W/ym+vQ/nJ7yZFlvRXdN9SqUD1nGNJAzTzp0Dwo2/Vzu/4Go5EHgj1Bsi8b6OLo+w2vOG3M
/ZE+BWIcLrq1K34edxGVnfxrZyzx15NtKcPqLj+fOHmcM2YE74+TE9uM1RxpeSmHbb/epqQmfWrR
B0POwsgH5FX4Jw609e3tV63QnXQQtr2lD5Umdt5SB0rXmS9I+N4RGPIyy7RKcLHfmRsp9RrA3eRM
P0mM0yEhBeXU78/j1wLeDVBtpJqtcia5GN1CUpE2H0GZLIIuYv1ovu12+MJY0a+ClmO48vHcMNep
qcaTWCvoEIviNiUsbxml44uY+TamfNuzflJ4epMf7GCogmudxch++5dx1gPWA7zFIrkVK8vevF8J
PRkAv6yn34DjVzSAGiZU3Q6Fqjs2LmVaV3H5uvXXwCSPp+f0HhgxvFvZM3dd4n/KZ3jWGFxti9RZ
FdFvbe+5UrNJGRzS2RVn0h9rUKFqL24L7qPP5nQMabimoTuDwL236ykGHerzdOL2Bo/A3XVvEM/9
Pyrd0T2KwGfuy3sF4fEl7HGORvauWSXGDDWMFLO2A0a1uN6KlBHcFKSQTF0XFsEhgyFGqL3UKGf+
zNe3EbbXFOZvkiTq3NkdQf2hrYsBt3ns+KBLiIIaZoqW2buuNOxYeCuFdq3lT1zjXppltnTQhmTq
JQQFoAZnVfuaChxczTHW/lOCk7yaXHxA0OshfTGmk19aTq4f8P/TzD/kHVGHjIfnK/fbJb1wm3Xl
vG0pQB07rLw+pCEYQt7tkXpZbZVkEbujngZSPAb/WYE9RAt2nfLgsZGtXNxAfWt9q+PrCitYjDif
3dvTUgbV/Ih/S+clH3XdZINf8SEhGO8IaSHGWJzrXH5+O63Iapb47XAavGQ5TNMhfyaNsbdmOYJ4
roCUpd/x0Ox9jl0k8S0ugeOn/FQxfLUpRIYcMyFVIG0RO/jSeqaLBGBIUu7pRgg/WGoUG4O1CAhj
CejvglqMIEtxwJYrykpFAebljf5c/KRe84ogvtBctLdPWyt9Up/XWEjXBIDz7HT21H6yIJ2nzwnD
25l1OZlJXUV0nXu2nT5swDqcY5wv10KcEZdElGHKLZ9Uu9bQrDmVOqyG0yavA4LtU/HN/ypr4Zyt
eNwoVk75+44oCNPW8EntoVvZ3SepY7MS/XchI8Rrq1Q2I9ON2agPlor07AzBis/KaRIb4CyFBEmx
YSC1CYn9Z2RjUvxNg7xeIozyOgf7W92QTrzA87hs9t9dr2cTMh06m3bv7GuT6fhuNmATxfH3ZM5r
3DquJARhtyN/TTs3ujajtGqYZzdWQl/CnZ6kaNzSk6s1Tc7caRtJlZ4UniFvBfTuweKtttQKjiS/
fxn2Y7mcOy6p3oQyWmCRgLacqNZ4E8KxyxTuo+pnwgeKQBxLjw42F69EkkJCmWn6dc9UnP/nitcx
3RQaGm5sKX8VWjkAS5ouh/f2xFBQnFPzUyqg2CgxaBFEQRfcsI71kR/KoCfau71os3YBcVCYXuOH
p2JnRlzeMAl6bpz1whNTO0KSw49nK6TVCRsCB1I9Dz6pFRwQUTjQ9o1QTPa2qBCvGmb+rwWan1Iy
huCJekxgVsYz/zsDFMWTQxQ7r3bhi775CYKLi7Rw9r9M+zvjiki5UTHzsRHSpSSpQ0/LwZjVdwi8
38uuxRHFvIfNkDPlY6MLdDU4g1KK0sikKOhLE6nOxXR8IsYLAQnPvqP+5vW7srssni1MEDj2wXgj
d9JbF5f7lAIkurkuYfnHWPNhG/SYt3P9P6gT5uQ8om79NNbpKLJOOQEciDiwFI2p/KZ7fE9OkbFL
IwEP+OgPHAirALwFt2abhj7MR/ZVf9W+GqosLDVRqKXURVv9lUQC4jBQa1DBNhTi9ytc9abS5FD8
Uls6HPn3HGnLrY1IBvUo2xGAoy1ghIzunJPAqPA2KAmHjIqpch5wNMIce02bwPhtzFjHzmjjU1Pq
ij1Mzbnl7quN13JdHFi7etvBU7ADhm4QqNoNqCcL0PGCpN7FavZtuO2UDLGYwYOCxE/1cwspYYr5
8vYlFLD9Ax/j235PaiSXLuyUCT6SwQwmaVRwvXkm//LBbVa4GmftQr3AQl9ns4dlG1bwmmvY9XZu
0miCcl8HGkPEUjK3yEJdrQCFMnlYxrXmK69hx/lG2sVGOf+L7R+0XxABneekojZNbVcbqsUIjn7c
fAq1ar8F632Vt/JvasXMPZ4p/Bfq7iEx2wLT12dmNDtZ0syZR3XYLe/OF5//coWjzqwQoRzXkVFv
bPZNAEiNAnV7Hh49a0xvNLWc9P/uKklWQG3xgBxDMlIanYocXZPb39bCu6vayAwEVO/zquVVgalJ
q13aWxwD1MPuPU475SMprZcFyeltKOYzMWAhC/BToIlZ5NLxeXcBGqZdCmkkEETMWOXOzrDm5v1x
twopCWKjU+s+yTOP2WKW0XzcYODpy+z+359JBTSuyZx3YDCLji04Zf0ISrIQy3bYWwGc9TmHczsc
4Rk8RzUwhuc8mEm+MTwRBo2408bGXIdFwkNWLgeTJ03rKqRCye1sR8W9KNrQ/aXtFUxACZe23DqW
73YI1keplWQWzfvaFXPyURQkM9WobwsHEM7S5nNV0P9VooX4wpvJJcXlcjzbtUtL4tDmUW8ywE3f
hqRrzGnyTjuenXnyqtNBcfhbBmIYH8pd7mgQESkwm06Wl/aI2H/KvbC3/CzNJdf+cOLJqDce4GoB
GsTinNehbdxvQpFS2sn9cGtPXA4BiaX//eU/DL5k3szIbp6/++ZW2a8qWimhgnU6h0VvIZJzmme7
txjEc4B6y4YhHQ323lYeJFNjKaZ1h8xIx4F8m3jzUfjKbChEmQqUDR6QrKuQr3D5bL0zQEBPEq2C
CiQ84Ul/goePto+SPX6SbGG1heUV5OGcZ9twg7kkmXgSQZT4DqO480l20j7J+e9APdyA8I76Buk1
K2qOgkbGCkfPRnXQniJGyhYsPgytBbP0lggicpnXUS1U81owHcnz1aAKjqxDAOYtmGLNmmHRnThK
dYtBCu9feB7Zvg9hTKznpJEz1Rl3ybWgmtM0c7MJjN7sQUPR7Baixsb+8trhSf7b3VVjmBSxh01B
3iiBEVj2eTmh3p2ZaWukEXywInh6RkN416GGbmdCQBlei/BPV5clXVWfhRGYvqhebbETmE3sewt7
qUx4rdo9SqaTKqfWxIRd3FgbxIg6Tzcq7jvq+fQzcPI+bolFIcDrngoI196YBzntOUOjOhlXHAvc
a3kHbxvpfUoQPAHWtmZ8oU0PpssIKcpZGKMLHxFGhc6rC8QuECuGbvMWGMWmJiNbsAusLM66ZWwH
itqrdl2cTXpwrZlAalNIzzkXgqRj/5A5j4DocwrlloGpnl0Y1Jk/PTFVdRevB4ZR4+8NO2/JTPFH
gHclpThtpeI/5nBazS3AXWWmzvXZx27Cbf2+0cO52btvGnsf71a2r1WF3cxZFrXsaTmDDJD4xdgH
e7PddnQ3YgyVF1jURy76ZCvMjz3KlR5fxO93KFseEgevXTDVhI95a4H1JjNlgh+4H8pJLQs5+BGr
zlix2uuj0Wcge436cKsWSv6yoqHNFdVvqBZnu8tQGnFoD/rwIaSdVbbpzAFb09/n8wmwob+Aw3BT
EIve7cpU4eduFA0td3CsJmH5K21waG63JIRsdrahH8sLb1arNIPH9flEla4lFRjIGiVCbPd7+Yyy
n7/QGrhO/vanUhcgza75QvG8GcAw+Md0RJOxAxIt2Y7c/TUr90rgzYy2AnjHyCTnBe1HLqeGrarf
i42Wjf5L7Vwh4XwfiZRaTNE1qwTqk6jF7nz/tUwZG+U2NticGYLZbCBIg0+ttQAD2amEgidemmCs
Rgo89yn/HgjbupUDE5t7mdzqvbJj74g+eJ7Ci8rkeiVCrIctJ5UkWSthczC3xN/rG0hwSlnqFtMt
0fuP7W8Avk/DVDk3k36NlLZctVSz0i60OxRpd//uI/OlgaCuxW9CvYqbmkadKg0u+lCLxJ+n9n9V
HpSXnUbhMMYtOoTWJelhR4vp3/i0FT7ulzjJ7JYEfo72CyYju5ORdmBa3E+geXVIn0IsFFtJvsTX
0FN72xEIhiKI3t+lJLCRQYmFQ0QZWJvidsCcS4yspsPGQxkx3VdASknH9aX2Ri8HM2kcEIJibV6L
l7wGBAAA4t6rxNNfSGRyjMvL6tLUUUwbBZxRlQh+YwB2xBMjbieskjGh3ILoAXs0J5qZ/ue1O/sa
pz2jy9FBjUTSvmja6pD2AtEliL4l49ZUAimf5GcR08wj5ttltKceDMqxajAQv+fh4I/BcUgzVCZP
HE/Dp1v46EdqacbnvqtILXy4em0ot9f2+Pgbp44GcTFPCFOJJgF89B9zbWRwjjEK2HgWhLJB5UGs
8NQR/HWYoyzddN0nOf5jquUz7JQvs6FoUj3pl5jRvG+H/4qVLZ1xzYNc7TmWqE41G2iprnnOABCn
JJymDTNdp2QL0yGKkp4QdDefSZpMsjgpNf72UJXKpAR+VPXaNb740OmmbKWp/TmoK+jqa25/g6LI
em9+mn53xZAmAvcVMvJuNC5bBIzStm5syEnD2nQQzOqZ5fvdPP3UPJ1mKNYOZS+PKILd/+wJITPa
IXCGpi3YGr8Vrr2zowfGgRHCXk5tnKam78d1cjM/VK7OBlSIj+CDd2AynOBP6qMec2RA8HXaVs8C
bqfeF33U7h9rkl/G3W3q8yuYi+laTItVv1/e60hYp8vRHheyUcMqVpYIE1luUk7v/QXGZN4PPjpK
+OQRCrFRirQSlnkJHz6fv9CZuvfaofUFj2h/5z8Poq9QOycg/ZHa84WDzYOeNaMfb3ZBwQ2UnfGr
mj3j51l4pFQTE+M647jlDjG5tlIGdaDDXFSzVl3NOHho/uNwY5o+eeMXSPUniOC2gQ6QxQgP/wVc
eJcP1EMIoy3Mp2ALFsEVkgh/TEY3hqMUYoM/FLqfvRuUU+eUD263nbeveQCWIigc/TD1+bUR4Eb6
7uy8Pf6IZbj2T8msdZUumJ3AAAzNh18X4QrmBD1WF4jkgJWafGmaKA89HmTzI7ul/MzZKpWbVE7k
V3/ERn9lhEG+j8ddofjclzJ6lPiNfF67kr+1TKkuwsmthOzA7QQm8VfZ2rmz5ENveyrFvtPgS527
tw9wg/xCjhpH1a2jJIBshNgzg3WU+QIbCPJfrKCaQYLbDmJaAObhK+15IanFgZgOsUqqwXx2kcEE
qffBKLOgFvr+Afr/UlVeG2TxqyylB+rh16/+Or16oGzN4ikyVy/toSw4IiHaEzjhjipdTqXh1wJY
HAi9T4i3bD262owLGWv3hGlH+n1x8sLwijfa5RtrNPMW4FO+eUP1uEoxzRa+1/c+u/8K9c+tELCF
MueY1QLKRSaSveociHscFpDjJuO6M1GCvkMyXZ3pVrRW5eKeO49xHopfHJZpTyLQPK+nQRLsiliX
LYeHH+dzpObWAx0V+91hXKn3gWR4XpqDRhbeY1Ryxo7Du5ichUxz69E9sBqyB3AEa0xdIzZr9OaO
mzKbjvq72g+huVHIh22+sn1W+g72pTnls1XiyDduu/7Bb1gnvYe59wP7bKYogv8hPizJeyRQ/o+4
83PtY+Y6+druEqvN8WblkKEFlgLTO0Er9j9wFinRZQP4T+VX2XlsqEQ4h868jT9Ni9BhXGBBeyhx
O/2lQIGMplMDubD0nDSFgEjA8KliES8EODtlVs/R2M3gVeCQexIyageWkZo6IISg/qWTHTVTd3z3
zKmJ/HpvvZDQNVI8cMg7vJoQ4bM5rIQJ2ETB7KOS2dF2XvWEV8YVZ+DjfJwogQ5e2EPiScjcfVUD
tVUSRnjtog7FL2r7iIhVhsok31TQZASkGvZH41Z5v8tppNX+4OdHnYTh3mu5ZQSioag7kRSIAJLj
l/jmkERUV0oT0mYl0QIDH3HFuhqNDwHYP+XJUhJvcW6q27eAkC1jZwPQii0gBffELNjNdPEqVPxb
+NTyLUoA1mnO6VLifK+cxQRXY6E+3bwj8dcEaQNIXPXubV/Tom8uZ3OVmxBzfwnMZQ/76jOBHcGj
oXe/rzfPrNoeqPMy5MmCB3fHH9sQUtWzorWyeneTthFCdi9UPFA7K9a5671LumwSXm3Q4r/XaOPo
k+CPm5UDQl/KoDiX1oGzJcjVoVM2i0ucfQX5d4f1w9bDZCt0GGmsRd1/IGq+bRp24rxr/2VJ+ZZb
31UUi5j+YMW8+jPH88dCnaAeFIUbhD9Z6cOHfUUtuIdubFshMe5VIZFro7ex8eAkrX8bApiYjvmO
eunZ+ochFlU6bPofbC0rZ6mh7pF8y40l6CvIqMwursnJr9jw0nDWWeqZ9jI2dXLhwca/LZZBIhSP
Ly64FkZxs0e+aI4euUjvb4CrcmPd9OK/in0y36flN8oC8W2rSAjfuPIVYmNKHXcBxmdx3Q09z/ic
v7rsX4chGNZc2EfLEiE4TzlVNHUUKA7kXIMRoVwM/jCO40hECirKdt19/rY9xNsw0yAT7oA1+qXi
sWHV2DwpGkXwh+fi2tjW+TXYG1X0d2bOBZ75IwGn4k5sjKGuvt8BSYMluiDQm500sTLBCeUVL2VJ
zwncDvEUHc/j/JRMQ6fB2x8KXjqXvyBCSoaTQSdyyvR3FgmUpPWFe/DfOJGoggaixvM8SaRNZQQX
2B0sm6rqvSRHsjRvPfpMJ1e55vjyZ0Zdf3vT9MKW0vZScSyGzTb2NxRsdAVknC+qYLGHL1jQ9QQw
RTkPXuyLnUmoo9oDyZj5rIAAG/fIL1mLoqvBFgpgkRSknrqGeJa29ojVDqsuzC7ypHuf6DGYr4uJ
2+Bikn/0ncDS7NsamNYcVVKnv7M/aqXMCiyte3eERB0PVTBGFFxzjcSrte4CSOyFU78GmKQm9DI+
kbKTiggXZrediBhFkPWLOSWTZo7b/WCrMstkpoiqgP5vjQU/N1sOBRQ0LyG1k48/4G5NcjoZIPAi
taBMSN+Aeaj2Cy96Xem6uBiYmiUQEYs1zUzfJ6p1WAstn0rnccf61VnZRHglcve+NyRfdYZiERAY
NONIlthamWdxE5e1SedBqorxljScXeDhZxx4PFes5xDJ/tAixCvW3W4ZCoCsFPtj5tp5JkUzciqg
HrMKHvfUFWIk88X6PjNEW1/RPnYJzWR+xlSmry9LZL1xdZ5JG0JNnNOZ1bhSUpzTPcvXqzguMkMb
R6PairC7LYfrIAQ6mjBnlFfUJz8KdqBnso04fdiNUDE/QQhUTN14Vd89SqWZibrQYrEbW17ZEAMy
Xb3td1RewCVsgg+tPZbrwI12vTtd48fcFyTElNuY4yejZO9+04pBfolmxovnV2A175+4+6SwboXt
s4jC+0IOu3EQhN4kC+tAib6yYDFIBmeBmifYX24dn1sFhTjE+Xb5M4pUDPuk80f29qcMiw0aTYui
Lq1vzglrEcaukvbKUOPxNcFh+TLEUj3kVR5Su8Yr2pAwk5Z8IChsklTfdZKwF/jh3t1TjGH2uxs/
eZwtem58F/FprvssWKCnizROoNlPPObCXVkxz6PqQIGf7J3bhgE+udVdEZhrSzUR6G07JUQIYQYL
+yUrhcPtgvh1ixsp9wt1pZ7dqStH7fceqk6SIT5ejwUmWED3qe6IuQZRqK09pCVAhBc4ZAtk7BzP
roGvm8CpXKAh23fl4AVD3y7j1aeWjnIiIOObuOr/rviwykYZ9FaL0Aaod2iZO1S+eRWGCjKmvQ1C
EsreAO0LB/lGTbtpuJhbWCydXws8GNknTkKYfWRXKOcghejzaCCLMEG0CRBxFMsWKtaHfnQCvKAw
VMity3cuaBWudujCoWE6RBrJPRpKexugCXzMqgP+xbhZ3hj8FglcilB79U8YGx3qB1+Fu2TRtVgk
5Ncmwyzy93FmD0Tt2MP4sNr0dAGerU84c9mekn7aFbONlHtgAauNYvYhRYKoOzQ4blZvVsOwQ3af
K9o+hNaqcbells3uldFDZMKDhzhhbhEqodfcmJjjg+jplD9zIa3tK2pPghDXgm5c1i6Y0SsgsMym
A2cEXEyiNmktStj0x9RIMkmApeRUQdsEl54watfcPZf+EgDVWr8R4DgRX3eA3Da93OJNZN4TnKN/
nnvpDbjCYINuIISbCrU/TB35N7Brbs8HxeufYuyOd8uZ7faF5YA+cKAMz1OXlyucGRq5EnLS9k91
eNzEaeuvs0YhvqPvOIcdE4BBYcfQhYQCx6HpVkbKLz5m0IEE4mpku+GQYXibBvy/H1A8rKyUmhoo
hJcjc5iC7TZPKZ+btZgMZ2kMhMUgQCK/JZV0AIZa23uqm1Cy4gY5jpeAnEw9Z/MWrtfhWZXXRCeb
dg32oezMjeg0PaLyErVQ+mNM/OU3FOHBb1iUdkfKFn2uFKqESL7Lf+2uZbzFDnbOnG+Ci7UGak+s
RMTXgCGeTRAx6QJxC5g/XoRkjYtm7VpNDsWHxn84mN0S1XSXAj3rVOor6FDfzHp4vf9duDceVz2Q
tav/3MzgWPitcdnBQo9B8l24yGyNhPpzkIMgaAk9v1X1VbPoQ7PJRUxmttLMvt1fK8PrDA9sBwlw
mUWmq8CSSpeNagjaaFm3E0XwjxqBB/KaIlXuWS3hCE6lRHjJQKYIHeykmXNpsOPG5TMrAztvDDIb
TqJMf4grhoADBXkpNTLRwDIC8BH044fDIK3AfFESk1rsKjNCktnEexAdl1Rkk07Z2/KlbgMVnsp7
woxnAzGgLOe1BnRNJM5/i1XQUNB3U0VvV+7ObvhvQEeDHvtJB4hpRewzQX1z8rlNvvIj3Q2g2kmF
9Vh9bFln+QeBPCGiAzdphfS76mjBzoThBYuP7FtYwdPycYsdCc/rvFcrzz1DGw696MYoTVrdNgi0
ZFFkLL7Ghglh8RluuYDfXcxvafEyTLs2t6dbZnZplPy9jzeMmT0MORr+f404y/hVRE9CjnrvAhHB
MhHnuWYaEaSt1fV/+vQHWhjcnHY6arVDbL/pkMJKfnxlL7vNFhPOWYCTZ9+jQNwYoAWb93OLpISe
4JtFGLPvwWj8x7ph8p/akr6jSfW8or7fZOMQ410x/Uqb/IM3lkyjNVz6Jg8vTG2T6zgQPbzRKpC9
/6P0bag+hIuuibYTSt6R3FMVqBCDDY1HSpiWJZVQjguyawGSTArxc4f9BlQyhsSx3zwKCVcghB6X
UbT+tgTKYGS+H+dxRPVhY0iZo8cmUhKo85Hi0uqA0WXOPXZAuOfw8XBlPRK8kXmR/lYGp8KXzs+b
gUR8xR/uUJXfipEDTL4W3HxArx5K8f9y4fLbaX2OweVuX2eXFzGNhvTRDXzgU8+f08SGoW/wsSn7
yKEQJipjUvt6UQ2NxgZpmT1pw5tT7DE5ldXpmqzH3GQdeRTkfk/XAGSZbeRjHlOuD688J2ALFF0d
wNH9p6Mzg2bGxK1+CuwbKBb2TfEuzgcM1DesZ5gpyZQxBWYOksASFsQXdJFHr3B9PHq0AnNKoHnq
i0CK0Wxqx8oRyQRtCZp3ndv9KtJyf1l9TiflLUAixwzNgsX5j/UgzpDC2PyI1ilXHv99k7f9zEkV
6PxEWW2vh9dgCyJkaRYh8akO3ATKj9MEmKd4hV5WBUOg0ZUQL8fU1Kr5HbB9N5N5Xyntcmm5UXtw
Mz0m5nt+V2oAHCqxGxSue9X2MtRD/5wEkfNwJKE7Z1TJxDiuBLVqbYhsy/tfZuQDo7Qm53K0RUNQ
2Ajlck9OjW15dV5he3DvfuH871S0Icjf11EUCHprk5Eb44QWUdK/ZgKeG0xgMuCTTSlo7ffy9E0p
eDjybVFrTaqo1JnRKvNZuov/mZ1sI+fHDPmPInNheArYQnN373jioaXbAr079ex//k9RnOTBVARJ
u8vVjps9CdBXwa3ZaxIwdKKCQLj/quVu1nrtnzwwe4p6bEhb/N74P4K3XsPRDvrGm0GiWXG+m5cz
BdHdNQ0pSmRTBmhDUUM7g0OMEkV68DvPXQ7PenwtelwaKBs3Sd8yozNwAhQalSQ28FtuqdPzlXeH
9Jvdl+X4hnM/nYzYfuBmUj2ppg7EFwDwp2fz9N4M9Dtr96Ky8QOA3ziKzvvZxfOemeWyMIbiQdca
R1b8c0npUKBK2Ik3o1A39LoROXf5OhYPL2prAVMF7QxkqEmKrNaK+0uPnE6LOzGoLHsysLPXFrSY
ve3iNTzACqi2JsgQzFOQ4qt1g/e6DceRIIypzCI3+CqLks8iH5AndDFfvDcatAJxlRlH7nBNKVt7
2mDXcNc77oI4n9NlFAWGfAwONNRiIqMTa2xHYuEGUB+zqRhd29ntHBvNPug2xDEWeK5KExmTWWUK
v99dvIlk7+98j71+LrAMuBE34l/0vUW2Fk11Y4ezLFINB6izdJJSXIpsh2eqEnWhIFVxCWlxXruS
7epG8MK4JkyOkfTggX+WDyheZKzRwDV9EiT0H6ce1DfdbOcDt5oGhL3EX8IUdjLe5BSp2pxjbyNl
ygOe1aZSQbgEIhqum1KW4UkGx4Uh/hU+gUHYDh2/P9a5ozzzwod2fyP0bNWdE+B7w0xLvhVvtyCM
svkiSpTGJptAjoTwC3ezfvFNCyYz2GjjxUU392blaH2yc6/pOvfYG7MmMaDY7NHk4jjlOAhUYYDl
fM5wmQNxfdINH7alfh4PyHFw8BfG3f0qG+j8kv8CXWKc/T/6aKMjh7McjJaAoEk8zpRJ5XWRzsLD
ngvaKWa5u6rhUgd6nlCQ0TRcSYBY6MNcseIPl8PXnpkVOsJj1wyJgqiVhIAcX1BgAJeCI2v9xokO
PKuAq4dADsj5mvKdXDoVpEOmQW/FzQ+KaZkZFZjFCrtnvcSbHrzLChGPThYi9nEpcXR7cI+mMe2i
KM01H6Cf8/kWeyRFhmZgGRJEG/kDyGG1xPWVfvmcZ19oc7gMFarTRWmcF9hS0FYmezKVXTmZi2VU
Gm7fT8wiW0//pZRMF+T2Cr85+ye7jmY+9pSMYr4QiYJedCaLN22JpwGy+Zv+Ds5KHbeQ3ankYp/E
3S7kBwkuJd/a/2fFL8hKtShi0JlrGYvnUjiaHfo3kVLLg1rxcUUQ4+t2X9TtxYlzJqppWB7k7j6Z
wou9Ni8owEGvychu79Hs6pybNtYtaBwNK63gRmQQlZmdlUp5Jf+MUEn4jwNCLb9bpwO2/GK8f8FN
TjTILlmbNhXEG+HNS9mGjPKG/TOxc1XbYAW+iMr8WcXpqcADZTgnsCWiwXWNf1H8H7KAftT2CpZ/
rUmwywJtxFjgE8G/f6jSA1xDtDdC0f7OH9jNJLhnTOIfUSf+X2MjcvnS03K2RtpNT8CNvxFXt1i7
GTe++Y6Txv62qXeyUZNRAFAIl3BvyPui70MFE+Vqg5VYOPqpS6H+sfYU3wDBmCi03felbwUPDttv
/2Sky9Q2uSUGZy1glo17L5m86+c8oO4VpqoOQTDjCbLVfZBbc6a5FnZJxGU+C5pmOJbfxQbTdcon
nrPAg0iTTJzbL37z+T62loFkTHXk4M6f7Fzj1MnGLLPnLzKqLr+6v9my5fxf8noAiD0IkpDMo4L3
NSB7L6+tC1AIazTUgPVntByUJWfwiLSRpNuyr2H9m2cc/kwmNyYTS/UfymnhiEb/ikasMg+MyciH
14KTpXaztKKaMjPrD6YV65/0vGTpHPoiWJxuTPifC7t3z0mrLVFQPCLibJ80RESpeW+FNIx8twSl
b0EBtXJlwJq2VQf7/sWHrQ4K/ZiTunKSiKsPa0bxYf2NFAq/rHCcDyMzWewI+snGOErHcZdqYBpu
cQz20ivv9m+yjlf6Bc03bzxkQ1tKzTuJlj8mk8Pnn13MbskXJc2BTKa1vgN6WuLo8wL0F3OjyCuh
fca/ggLqk7MBKsgE/VqnFGYYmL20HXg5HTnL1E1g045r9uwCbwz7yMaW9/LIyxJR841lKWHwqb8J
m7bIGrdU2IcmNFjxQ8E6ugEp6At3ZCBy44UG6q2TGYiVSn/TPWR8tE+V27V8+F7giKQ+wNmgjfjh
NaSVPg4J6B8pl8mbt/Nj6OENfUxqiL8uFxURyIqAAxUbYeGCRWq8RakRurTR40bz0TdNXvQ9aUF7
xDVruKY2uyzckS0vnzcfXyFvcbib4cel1BR/HD2dJf0vmhU0KEB7USGdLoOHUwjW/CIDg68OkFAy
Oe7fagJWQwYM2iWjTudbmBYbuEfJf4EUUXGWV4fEUYoAd42/HA5b1V7lJThrN+a1kQBJl7aHtl2J
0Zd/mJLekeq/kYLbiGehk/PtXuxnDL5n8DOhsGxybPTYSmQidsmav8g3Zhqsw6xedE49saf/kR48
S40mpnOsxJHQyZB7W/tcAx89zZ/R79+A/EwZhva30oYGZ5znGoATll+djOqIoKlGq21jqeCgSWv2
1/tMxWKvOiykALAlMUgNchNUMXDHKYHgK5SecDrWWsl/En4C6l3r4F/PbszBdO5EnGzuIJht3LXl
DsDh7VVtgH2kHV0qEo9s+mmBdiHRa/DbMQjyh6THtKgr/8XL62q+zBWATquiNlx2hg1bTvNLtvpr
+9xhB/uEijWqBv8jL9rTzJebtO1rRJeDRj5MJJjo1aR4eIRNhx5zmf5hDo2WLN+/p5WNt3vH6AU3
4ctitZ4nun57E+2W/zOV3gXF12o4AvDj4S+u+jByjQFwKLIaP0GBACMjSVMeNDzfFs5tviVBOscX
m52bPwYKGPLJ6JDQ0eWctIIBUzfoIhzFn+7P+iPWtbvEvs5+pgN4AjPSQMeTS7npHzeQE+I6shSl
viMc12QDEeiDyZ22POfmKcLv4vZJii3UVQ7NQNaqyvJCkdHnO+ONI761ORp4fk+5VRNlfiYf+muB
gxrtTNNuw52eXafJUDSPv5WrWEcjZzW3TjmRGVdtMqJUpqgXg6D8UQl9CZgfHH7ZGk0KwqTDTKbw
A/68+d3TiyyppsZUlYluGnhfojf4ZGgsz/3W8V4XtwhXRk5rlHFBdBIC4PLt4leon2bXOZmJUqUs
RgqsRvZBDLbdumMuyDkUs9gH3gXP75SGd2crcG6LpunkskBE8i+g3ya++9PZoZslWqQ4ZGclDm+v
L1XVlhziPxCG55gig4nheleEdLRYVw/VPwnUCUr1wkUKf5Lw12OjsAv5DUnCez+QwNZnWVnCCYLG
Cu55RqVLoNwXO2+dRunuBjVhl8hRbNe3FMGTJlKZN7iCQvKZpsdMJJdubNNZkFHgd92HHs5NrXgx
7xBBzcn5Ceuh6vcFS2i1LbgzQh1fVP3eYH/NxUFtMzGYUkyY3XolETlXvcpHB9cEWHpHLBEJxm2v
6/wdskSt1ZCKu3f61vEl9sUjWGxlu4Jcj3PY2ku77qLiB36CWKpk4qkaZdqYh4vZKf3CE2Y3paVt
JWCtTKNQ7ZxZtBpUZjmU4r5WraXz2CLTkTLbv+gYTd3j3cEncqfrUoltYMD+pScG5DOfk3ARbUIJ
VG4d8s3NH/lp8AaFA1wOwK8vV82Q7lG1b+GqDFrWhr7oY2th//wrP2qfPvkDxp+ZqD9I1lNhO+eh
FFG7okuk/k7QKCpe+Lhn09sjV/xAmoZiCJzosvk7PCS7rS542d4zoYof8v40AzzQS43qOT7fCzOK
SsXnpuRURdWbIefcA01ublcK3UrNlPa4oFK/kF7RoLIB5PPFEUX0hpnfPXo4K2yu7+2jPqVNjgtp
0fd5QqiN3x1Y16Ut35Qrt5/9bbo/mHLpxlXdr+FqU194xJ7Z5lN8nFqzJfoQzikrnrqqYVntyYnE
/mJ6qAsi5MqJ/qgzVc3xWyr1TRKV+8+fTkxGIzcTpHH9b8w38h4FWpylNGsUIgGIL8ICidxVf3tQ
laUkE+LZ3csxoGHwc3QCZO01TKOnG5usLJg65/PUtuV1X4TdJFPTwquwi7doDidAsmgPSOtrS2aC
0JqrBwhq+DtE1Tj9lCOJSLk7a6bcy+hY1BThNC4hrUusDLF+hx3brEuNjJ/TPk9ALs3s/DXRpkWa
REh6xf+IAQELjwY6N6vJXd2TQHrje77u7DsyaJWrWdF5uqLgB+1dlCsA1ZKxnmFQsRlCz7fEylyp
uBVUwG86w3i2TfP4TALJcHhceP6X0rUdjSIBaHGB+5bAJus/N2vmgrkSMyUWLKdPAvDC9AgQJuDm
xxukMbOKrcTHHcblxRwPAwn4E+0zMF/yEpmEGVa2N/lWaLN1P9SkJ6JpPPNNf3Pg6jQLjvdm2vve
xlfboxomZvo3KVzPt7GMY4NBKBx497ZFVL3ffovIsnB0e4dW4e1OttpDiUhluT6fndcHIEuiU5cn
/c3nvlxuuqb91ofC2ifXAP7Ul0FALgBuwGiXFsuEn1z9JUzDv5y9R1Clu8P2pUtlwuMfn+IXtsSU
NNVCiQZtIpwPULUJ9PIMFj57KhrN9yLPzgnK0LVIzarbRSNHUQh6wPrPdCxFHGG8NJ/AuuKp479L
gq6zUqFxCDE6uMUmz9TIVV/4mYBHO8wcxtllgd0FwgxSmMIqr/fsvFqOSLQsiWkzrmFK5cT5ZLiu
UtPOGywDaqFe3QRoYpqLnilUBkgpr19ceoyFJSN01uQQMPgV3CRuQdX+fXd2VfIo97FFYtU1HKpP
wTbtOMLVQhdU9JmTUVLtFNHT0PWbhr1wc9y5+rRD+or7OSWk2fdUofqIfJjgYeFJiQuBFMH1vb1P
otRGU3BItugOdwKxKi63rro1Wip6+uQgnMmXSDOwhCNI0yRHlQ2nUodfGevWlTvnP2x8hkSE9jA8
gd1cfq1QQrFt8UKlbv/gE5/IgCtd8bpyDBv9q72afUM1khSKSOQAsEeKx9q8MhGivXakfon78GHr
PtZb/7YXcC6sUeiFgdbGx/UGn5GXrbskdrI7+qCKJjzLd8nRsU8pcipBwmrRGVIZoOWk8+bV6MU/
vVv6mIu//xO31gR9PYm5r3/pQhYsHVxuZm65X0CcaBrb7V7GM78WtKbj8LcPMiXv2zzI4Q9ZgjnN
oncKPMI8qOW+V2R8SfsHP6tWIJYQbtctDay0pBkMixArkFY5NGgJVSnwjQOMpYambFj/ajVhP7rV
t0uD6cWYNTBdWdobYjmY1qRRWzpAgzT9qiDn8k0OWtMmhKfEa/p5aVHfHWRKeu4YkV24URnxrr1d
f/ZPTQHK4q+++b02PcjlwZPKTpAxmZULH/nAHapb5xrg4/sm1Dj5OdIaAP3sI3LsVFnC7exI1W5z
iMh3Z6GmC7GmbvhArt6b3NxhEjtGifSFN/bFMrq5UFVQ767q0yaYIjsWgUgDGRNX/X8G0lbJMm0M
mecn5mgCEMenOw0dbg+RafiMX1Ail4Z5mmpz+/P6oyp+PP3nmujVpH71IX+EcszixpQweO78T2Lw
LvtZZsWO7GUWEvD9IgNiZQO4BD5880UzKaW73Ao5u/gIUnoYt+CDk5DvlxQ1uSQZRDaqRGFN4uPN
ayuKLurmoyAHM3/m2m9Vru5GKIkWcvkJauqe1yee9pt3UBLykDQXu0CVO9VpHyts4lhwaA455Pbh
QJyk5a3QkoBTLuqBB8AiwVEyhycR7LR6ClPZfs1ZcrPiH2IqE/tRkFZeNotVZMKa8YORXYJrIRGj
15eGJ2BMa7mLAh4456o5FyfzNVFuZ/ia7Ml80YWuYqerQrilLbW9u3TRBrwUoL/N/k54xGZHlebA
x0MK1PEXzisf3+iv/xyhaJVb3jBswTKJh/fJIbKttYYToVhy10B8WI/pVkrgI0DngjR0lrhp13Ni
1n2rNuWpYBbbyEYwSl8zm1KrfO1zXAJj58aufCiyzApdvSAWlLUU1Gqn1S/tFDiQv5FcYyW2zcRw
Pca1B66gJlHsF1eOXk1IOkw2y6cy4eCOvTjgFjcaB/6RxCmRw72e/YU5DsALdk1Lg41CxO2njqu1
wPqfYW5vwMNQcoCwwLINtpFi/L2rWmvDg5/EiLIOG8C2Nl7lieaW4D0rHhXcTnUt7gyRgk6sJbrO
/Nq9PKBUnZewwTssNEQW4s5LGR+SQWXJU8ntIRJTw6xqJBK+GHjyLSNHz/74WCUQDYKgFPjP1Qfg
V+gaedHIZSKiLEDKX/W3LgVCisQkHhAl7oFCh7xmBcISiR0ur8E6s85jiizxCFNdBPifbP+R8LqH
0Bx5GePfbU4Jmh7KVQSgmRsrNDX6dmSMAWZukUMoEhJpQaSQA49uyW7YKu23lrAwJnOoonO6gO49
yrbuzRWouHvS7T19Z3cX99pS8eEst/wRJITaZ3bQY22g9xlYpSGueI8kGm8NDNIr/1UdR36qxZPp
Gw7WISOzoLINY61tiO5of5buIT6WcyAMQFSDgRGG6Cv0zj7p+U1zFKU3xzC9JMbjZHACUKqCTDuK
LnymVVRLp20PnHhxXT5onUiUNw094ocHlsItjbFvHZp6WNK+sGZTEy8Uo2tnj5uatZGyhp6GKt8r
5WIL+AhTzE/npWF81wXoxFuc6neAXCUutsY9gmOy7a4C3OF0Np4+4xK70acAYe7cGo5kTtxMAj6P
8f2yqqK1BCiUEEWjA3ewRj4GkPxz3Xrh+Hmmo9ZZCxr986j3J3O8065TyhxDZml73jm78VbOMUiZ
zoQrYhe4nEFG2KFU7ctnpnzOsFOyd1HtwGjByPRjxuYVLSqhq6pw4tM8DKs4ypsSdDxWEYr3cDQG
H9MSjiaNbe3Paz+NI7acEfihmLb3PlgMXidZHJxp9nO1nc4TxbfDH4zmbg89DOLU2M715kXTtWTP
MWGTWFMLWJ9eGwwJm11Klw+7TgqxRKj1xx1ztnkVr7tyVs9Xc/aE2aUB8AHIX5ioiOqO64O9cRnJ
nytIs4hSm6CGVYUROt9MUDdP8D2tC+1SQrjVldFwgZTidGxIArAbuCtd5gqU+L2TtlPH9q5Vhijl
FYNMoec0uQ8W51z4B3BO7SJru4rD0afS3n2zKDdw5d+RJ8w2yRjRpsNEz9h7pgfg3GsTCeOA+dDC
LV9UDRI/bwcrY50lGDlKjULHrbshBrljNArzwe82yxL8Z+de01MrWG1kh+Qal+VWvkSxilGVJdso
S8F3kE3dGGI9o3gdE919pjY5vVdWSOgsvpRdq4thlNnUAxokenFO1uktdUuRZOoRA4+eWzkVxi1u
l/WkP6UdJU2XRdRD3WJdsPn22EGDtGfwsrakH8lqFM105n5IWJa/xB+z/bfnQJymhrDjGQqyrgka
Y3VPC4vSRzOOvxgyO5iOz2QdcG65xA19uhpkQUmOvfTOqSIoJrUD7VmohlqJbVvDBBc5/soOUgvo
aKrcSQMXanx4lViWh4J9RhvwPc6ILsVdDpbrimowoV7OVGgc2xjM9xEVbG9OFeouOJWXFH2YvYli
7URQuq2VH746k0S3OQvHBlTqknoGTy7u/lquzgbA5kPy6uIXm+3xAP8d+PXCvyMVWmBy1HaRUFcb
5O8j/yfOLFeNd6fNgtg7ZQj2q/hgnyNhwDAGtJBuABEyaYr1/H1fOX8QAuYSWz2O8dKAoV4bF3vK
trPpXIjc11IFWrm7IUpgUQbwMJQg3K4EGnejtv+rjmA42kPDwR2amP2Hwu5Efg2EOJ+fJTAeYN54
aLBgKYdmCuluovQy6l0AdsrL6SsfvIaIh5sqByAkKWyHlw+jNQtoSqen8uDtXxa1JpKNOab4XWZ/
teiV6CmFzYQqJdRSjr0Pp+ubQCgDrdnBa9eU9CF2ZvMXtEJ62tJQ0+ES5h5fa6iQVrHU/IM1Yb2C
i8URStzD8Oq3ybJ/g/zcEXWUlSl7uBUyVT3UBgFVZHnYfh+l/cxZEKy47WATzCc7LRMQgc0kbrBL
OLI3uBvH4PkEoMD3Oo3uZnOrBse5vD0e8SgxUyIX/LDv4nR0qEUXeteDpzBl92vglkYuj6lvd3XY
F1Eds3mo6Axcke2yQYbg9n3FcfMe9Ai269xzosJUJZUk8cym94ZDJxXNUfGW6K544+OhGP9f66Fw
Qzo9waodQQTZDAIBgZ7+SIWtCnKyd9aHYrw5JBBHkp0mORY+e49DRpSD7iFRNHGnhm668dqgpBLc
Hq2sOdkRbqA1ODlPPjVbCDZv0xB/JuvcONeX+/gB1/NTNzOREqSR9HXsywIoxa+0FPDMNK0W2fN7
EiYpE1ZfF/5BROMUzJ6vghmqva3ceHwrcdqwAREji9gqTwJ3Cqvrkj5dzr2cP6IL3C8rluwsBFyt
Q/+n2B3Atp/ddfOgCi2x4mzJJzBwuI9PuRurPMyQmLhRUD+WbL2K+gMr7nU9rR/9eLj5OlgJGtL2
D82OOlBZjWpH4c1y781zubWha6ifmGrVAor0t0QSOgh/EkJdvuy3kAkMHm0sx0OP2F7hSx9UMrFC
d7yhCwy+SJT3YAsjZsRZQ7XHxZ4rdIMP9eFfYtx2nyh1OxqUALWztMW39LiTI0MbOp6e8/nbylUg
dTCfKG3+oDlIULKCipXd6oA6c1EtVi1r2+GEDk8Lc7LsxbF0N9/NPXJiWsp5nOo5YGt+NnZAcUxp
FNxdeM6LREMu22GlrRnDxW9OD6XhywTW12s+SNyEXPJx2XljL6WupNKJ/fYH32JAN5N8esAt9fLK
PrNh/p8dh/rKnwgMkTYae4kShwgt4Try9DfeudJbmAa5TbQ4gRpOgwcc16k0vJ1LjOPHihPepGRf
IXB/jaxKT0TIEWWD4JcJcGsilexnF6uefqrVOgGVMcrBV6v4nffm9hlTvaR/2uzn1iPdLCC5LmiW
FDUAKFMJaZK0ZKCCdbWMDuii49pkYe/LIDd6Ni1Fx5rGrf3BUmb0Q3VVadtREUjtRRn9FY2icpHE
ZtAt9hXI1cW1Uq8uYC0FRgHUVOzS0yMOm2Sm4qAiTsmYQyPeH4lYcIwMR5kyIPM8fYqIJfcnmj2t
HCIn6oumjF18s67jsMJweHmtBoW3DIK/zDcGWgX/bARjuZFDqxdLa56Z55NDdMJv/tkpyaAlp8SF
W4n8d+OsE3gj+N1m3a2NTOihJ2uiKXCI76aFYA5ULYR1jx+UqOmb8g8Irmu5keoGCsaBlTmPGHAU
Z4XxorwefB2S+hyuhErw3dOQj4QEa25/iKX22oZWFuYBf+Plu235cgzeNQpincfAQn4fTTvfoknH
OuHlwGVmRDXuyPwkW4oC2S6HoovwgvvS2KuT3Su+SCou3laqvY9WEfcI6IQ+riB1x8pTXgX7q91w
/WvK+qPHoCfsn1Db075XvHDIVSOph11sHMmfTwpDYUW81ggNpsjwO7EsJN2xNMsO4740NJo03Ood
vAoYLfJd4iIhQtVgSjvlYHVG5rTSFvZ80NoEPYdIsoc0Olxykz6HZdrNIY6JHzUq8pSzgMZZSLTs
fYyTQVIOudpXaVhhrE3BkkcQ2o+EpQyLK7uzIOZCnVPa9PCd1kTd6pD0KmZpnTBS/ye2UaxeyxgE
SPChBv72O0jCPPWwloFC1226bXHFSeNdHCVPJBG8WWl71hbxNzPCPCUbgre9nDgvP0BBaiKPvxHK
SDUaYWDXFMGzIcb7845Sw2m+n6si0G8hRlpVCBBCvk8LBjPuWfmcIA2BgBF5t2OVL/n2MPc/m56O
RVhN0lCgXfSuVlq5PpES2Gzcho1L82VUfRvJO06nWgD/KUQO8I7SwbrzZTMGYBkIoV4dF5EzNyBn
nSQ+jHUDvBpz+PZup7/0rCFxn4dYKNvryoYlrtSHQSlxPWoy/gD3z5x8yJ5Wfznrwue/SH2jYUKy
e4fWb81QUTmtB8RLIpCEILzxuuM9CdAj8MH5DfEz1VxeMqN4Q2V9dxLYUhDrGW+2PJ4Ic3zKR59/
lNKctDALWhecTmeS3JFfTIJj9xahcEf9Aq7y70imccGH+Q2VEDzLroUPlcQNDRLhV8k8ufaMzRrI
AcDoDtWqD9SZnq1cFE4Go2vIMMhZnZCS+mWGdGKH8WT4fAGdj+76FjF+rGh5DQouNT9d4P15ezzI
RpQCSIey4bpXSLH3MQ7HrvvaTyGPXRBDt5ATmEM5wH+wgSffnMktHcq3XyFWnkyKn/celQ/bhVTx
r/+QqG3ssROQMXTlb6xcz65/jFOdxwdAK4VBmGFMGJfuwlwN3CqrjdwSYdb5dKWNhqX8QCnOrtWS
47E291jzvRyvfBcndymRo9mYA3hnPI+JpGbPbaw7CnZd1qfjflKQeKABOwLRXzuwWK0QQgPR3keN
a1gSm+u/uesNClvlmHOaDj9zAJ3Gm1SNGcHc4uNpPuiNpjjvOAZUp/GUs4TxF2q2gR9Z/p2nedg6
45uq1BEEbZwVW8C4kGWaG1XJTZZcJI6Xx0QNMkx/qAq7WED9gEi8rpjs3gWT3iFLkRBVr8v9BSn6
X/FkEGghCo+1DmDrk4n4iFYivUEfcMP7E2tAis7n5BuzpTPueTj2s3TzDzdRK6Fik/eLbLo0vz7P
OpEidv4lBl+r2v5b+xoOi20kmdNixLIC/cnF4kKIE5JAewRsJ8J/2DN3oGX3HSYrinW/1jmYN0BD
ABti0QRtXH/BYjrT5ifxJARSamQD4F25SwsFdNrmbkHkV8EGC+52+6edlgn/o3XAn46nM9P49CIy
FFwBxZ2Tk/8C46heUNDjvKZ9nSnWEE87oxFJRpk2ZnSZ7+17Fvfp33yP4g7IOH1BZJYJKGgLEdQS
coow9OgRM1TQyKS9FtCOyqM6bOWvf1Q44COfeILdNHFLZ+n6NW29t4PvPdzJdM9tGkb0wlFA7/JQ
0a46uxgqGxQaldlGeVwoUxEeOu7jzXGB/72NjdFfVq1+oIupc1QdFff/DEwMFQuUNenyX3wDuxxS
dDPhwP2tX+TI/LPRsm0PCaG1mfGtdnqx/f/KIF0y0m+ze9KJ8XPYDMETJFWiGhy0s0FkTEBOveCA
zGApWTgozkd2yl0AtXQQ21NR/Ah5XSaYKs2OKSzxw4eP74c1v+ganvbom6s6ctoWtjnYyaZ5PCsi
w2Dd3gYJwppuLno1y5Jb3o2F+UPaVp1D6o4AFDgvt9xLekDZUFXQ7Axona9kDaJM5sLWMCEHcRaX
O1ud4XtY30kZi6JKJtLvy+8shua2AJeGfvoAiocs4HDTaz83af1X1H+TqE6KgB4+2GLRYDJIAgzp
zfAF9vcQCoa7SqmcUv33vZ6JPMnEUefjJDI/7+yP2DfQffBMrW68Ehw7klHsKdh0NKsojLnC8OBf
KyCKZuiV9J21FyKtLapT3p8BO5apC6XYpD9t04PhKwVla2YlKMj0yLNXaWt4BMoA/6an/S1q/EY3
vBnuGCZOamQk886UaVmnNAkd2NH+HQjDqTDDdSgquHIeSfUYYalaiKJEt+BwsGYlWqXlHDdXYWbE
IOuOz4/QiXNdX0LXgd2vQGM3ywglefJyWEwhe5cIxBy9b46vMIb1h27hz52dYJtFpVYlCCf+NL5l
seRI9cmVT058RJrdHcmw86GWcH/lPyuEXQsJQE7Kj7ORUYnZ5SodjQWowwLTM0z2mcy+ctGvtSy8
NiXdkJFav63ul3I6ND4Vc3cE/Nouf8xXNZSp/LbMW0AJkHVtnO44Sa9ipcpn2PYvq8rKobYtYnpY
avGrtJVZ5xw95ZFFjy/YtSOjGNwZV5POnM4Ik1xI5pZnKrHuYSZ1ehimvosJgwZwy76HovVxxlmt
B5GnXtsHulFgh2+n2cReNDEiH7E+0zPPQBPQOtJvIQ58ohIuB6j+srAPU7ghqT3c/knw2GDCyU6r
T9cP8ZS/k2iaflI4ueTVF1j9P7LYcFnZLzBIYeyTSL4sz2V6ZtVV6AMytVlMqVHUA49Tviqh8Ikq
eN9BM8vhD9P43LQWo9/PME4pgWwEB1x3oFrC1GJ/F8TMbhh31jT+D0yM8J07vCDR+lrJen1oTaKb
Ns51Xi3VKQgU8RxNaAPWEiBG9l+KuLbED9WmLpQRyx7EA2emmUsWnyaCL6zD4uZed1cm7zoD1Y3y
Sra6sxLnGGnpYja1ae/49R0HkscUaN7DQfkVDD2zX/qHohBPduvmFzT3tocjtEWOvWkwLSfQhQDb
+4zNAFy6AIZpG7YAkZvVoxlx3XGKoEQeBIwjhs/vlRLYwYLbTJnhY6WWjq8HmF/Pp0SwW3kL3Olu
QddLal9sQNhW0xDpNPq70WTML0U7qsZfBbPsS8sCDLZikosCY/0HVYSoYL45rUWSzM1XF8bPb42w
0F18EmkUG8afsPPoZRo0IbmNpwfTgeEF7voC4fo9LM/xfe/pA+AoHX9xWIe6z8YIaXQq9rUk62GD
YV1zLY0BT4dZtBSkNde6IZh4hdXlJsRJ26GFoVwDXj5b5lt1P4cyTYWnF0/fvx8zLXasD6v13K2b
w+2Ta6i1mK3dOufDtosDfwoo5gJQWFED8cER0ckaDdl3z+2dW7qMS4FhGhD5U1IWVaph1JdhzC4o
hZ6OvzSe5oQ7ZgyQE3/DtiOPIOxgPx4W1Xbt0753qJP2f3a/W2+nu97HZNyJY+iddCCOSSspwV47
BnKjZey0llYFSN2q1skjdPPbHlazdawZPxh/Bl5O128AkmV3wylNtuhSgWDeLzeeYzNKo5fEO/rV
ITN1U5ye/Oe9hEgH+UVygTxLuCq7bG3dGzSWv6Mu7XaQ3Gk6Wo/Vnkt6ss5b0d22sb8/Cb16JHzH
4RUkf6clRwefJrziH4Xh3qchCCRIEl0PKlCUlmAoSnUT1knkWF12qsUZSMBIO4k/Tqs3PeF/5aOM
b3sn/5r8ds7VEvD7RyJf93FRSgJFeIPMj8PVFIjzGPMZv61lUhXXCYaufLZSTPoe4dFsvRF1joTp
xRS1pcvV0ZxEgrP74Lr8lrbzm2rnpJ4X2YbdhUu0oBI2rMLJcKSLVWQGkBj2eKu+920qb0ZMN/6Q
QwVN3nU7JbkQ02n+HGVbNujpRH+T9ZdWOKZUVYQvI40/IPR30J+iwZGmZF+E1jX6OPuIsw2A9GYF
mC6//EZYxU2RD6oyjoVZbn9UV79OcR0AcUEpd2ZqP7niY+i9Al8w8Z77WxDlVcxI4A49scHbNWuw
vCT4txX41H9FAnHdIEEqNQWxtMu6wx5h39JthN7evzFtpXEu972ZGGbo8e5NEm+qHc03v7rbdlGW
E3fZVkI0UWIofRFY5+jOoyb1B9AbFiBc5iM7mB3dJ6VOvrGSvnMcK9nlLOUEqV1RDqUGB9+endae
qPISlh/QnpOyxPlSZUJdyikaUdFF/fvE46GVR9u4zDK45ZPs657i7/HH7LbSXeE/y7fXqa2l3FId
30l0Kq8DdmkiWKkfz6DNOz+3IiPIYPYyYUQ8xmnrRvzycf0RSacyAehouWPX0O3Hj01L01DBOGy6
2oXqrAPDloHwdmf1s01Chjw1IYpFFJ6/l43E5ucNnGiQaY9fb0SCewZDCwmDMf/kp0gswln7RFyh
9h1SDTuOUid8DlZnO8UJXyFiIzAyGDK2Z6kElhVOzJ2GVC9LQVRKqs9wLUG9/65VPWsxSXdx9v40
SLzoGzsJNWYj0E1nKUW52I9C/gDq8UjEIX6Krq5EFWACRFUHw+K7b1PuFgjrV1L/jWYKcIjzVK/H
YOdywOHIHqRCWsXT3k9k7uGaBFbrhM4iiZ7bxpwWbtc4dou+9TEDGBz2G0tzeZXLbxruJJmZxcFV
TmEYAx6YaXf/fuE9o2i+VMmiYVzonRm6P2DmgYuHzYi6Al3ttm8L3SqOWNlDCSg+9TLhORnJ78Vs
gTedbeN3p1NxR9ZXlZeYHpxKC5996o10ROQ35FD7nfk6EdsSlTBBGwPKtHW7Nu1NNpvyUEYqrszA
aPnE4EYHTlV3+HiROtNBb07Uhktyi8MSaxLUAUAiUtxrYyCbFaA+IJQAmEOpAwOiZ8YHj5uCimvr
4YYiOSRp0i8ATgTadeUx3kf/1z0T2cMeCEK7NZzAj6mlfTi09Cu37W72srczo8Ncowup4Y6O4MQP
yo6jJdBUhyJliLGeyZ14rma3z+xa6EqMDeDOr4gjRKCoyG+Yfk005BGiO0Ll74beGIf2licsXvJs
0jyONzTRi9Mg7YlsxEPyLLNJs18mXbXmrJs0PiTTBMtsnjudDu9m+IT1FtvWayO6GnjSVxv7Uu3T
xPT1I22REIXsU715PcqUuNqweRnL/qgRLAyx51LwBBa952zJaiatphVwp2qxnoL3Ea2O32R0Q9RW
Z+RtV4Flq8b55btBgFTb97Gn/+DKJ07XicHp33QhnaIpLtqztSF2ELh0sGDTA5ZQSCWXlV0I6exc
1dD2J0kOSkqLXniO8UMrWOcmxKFhROkbn707ebf282zVfWNVCGYa035Qg3FpnNmxlykMawiIPrNn
DxTozbyVl5OR9vul+iimQAVSJDLOeb/VsqjpMVUjNf8KSVjl25KSIJMpSzTRmva3wZDv+FiP33sT
aXHd2XPkE2VnYjtQccisQHOgh1g2eXCBLWTaiPgwgasj6i9mq+QifbcGc9xyFrmGLdhJOU23x4Gv
/GGCLYTXYXMyQIOO6AFJabTjmiVpd+NHlz9xeWkFCu7d7jcv11cf1MJgXMZQR1iUi+fVKTkHIcUQ
5m4jwQf86jFWLL5W1xmmv3zumISVuUGUZZb93vKJdlsuoKvFsf2tuQDfGYBT3h3TafNLhikmODrp
WUFt6/LsQ7K0vRjHy57BidMYh+bS3M8lLI3+TmKEJrz3CFgnBjlC8utmLvmvigNL9mp5ypLQyD9c
8Yuh0j8n774LYFSp2OaNl8Y+6uyDjCxwtHJLW6oM1+i5+j4c3Yt4x5JDmiQ51NEg/Gnl7j8uvRRK
b8Z2T6B3ioD5jyontLdcg3csJhiQsGg9uau3700aZns3kb2BaOfqs5w6IPVhtBECC6U9NeoIhfY8
xEMjFl8Y67J9aJ2iooYM0CjI2hC7/Cmcy4v0hF8ZaJW3HFoOcQPUQWHGD1J6jy2K4bf6r3jRUOiO
lN/dBtEuz9Rfy8oZqPECtjULMEej60LHsXCQOvb0TZkTzICvguB8ZIJkTrVX5oRottlHNHejpNGz
T4+FQNb8P1dDmlbzRZZK99a67bp0ICMohUOYzQjrE2vKQgucSwfc1A+JVnP4HLoahdWzfs97aPH0
EZUkoEflIswLdZ+IGWwMY6IR+nKQaNS98MlGdCc6KB4ycRtWZdo4iirkZIvPoBgNpLdX83s/pirh
ufeAq/fFuvIkq7NyKlx8baZOQps7c+gA63g3gViAkgLMPFIiwhoZWheV8fA1sRbqKqDhobRoGwwU
ziZqhgswq5gzD6Zu1lj/yIoQUQPMBkJaE2SbSimi0d0vJ1YYFEthCQxeh4dJyqZo0AFYGawFTHg4
T+buWnmzfgL6wzt5sMcgCnMw6AXcnh8zWqhnBqRBj7jVwNm/cnO0e9BsFNEHMmH0XgZqEfufF20h
855sPfilfoHyZn6i5/GhErqH3mMLZr2kEvZTn6YZDhJGr5osH9xOTfIvtaGYP/zSFweT/8h3w66+
ce5qgiUHmfcn6TdgjoaHzksNjLSLqvG5fF7IPyIBYCnEK2XH7p3uJ15bAu33EfIlVLG/g+/4MMRA
WgxXgCEuVDh/Lu0E/D50OUQySKa0fIvA+G+012v8nuEgz/mWkPVFBQGJ+pvwOiPLo1d5SUQ3v4Yi
qTP0XPIwCQ0t5gLOnrwh08dRkN1NGuitApLhk3+lyoY4662uYhe9X+S3/FsnWfnKLmIU9ugD5aNu
FWEjNO/YCmr12n5YCYFJCSV5VDjI/rBIXAnru0rvDfBeCDXyMfYtsncRQsnBlo8f+KXAkW+zvXSl
Fq4Ks89DQmx4xjz15+kqo0YjBUuon2P3p23JACeoUhIYZBGiC7HOU4WqauEmlsO5xxvHrnQp2CWn
1/c62LY2TFBtQ6xbdtijevkm4IN6iItqIKwBrSEhLuziwNvxJEdZalUPi69TfjjxpFmI9ZqW9odw
5T2xayWVZTLFNA7dFZtzcpYQgkIUfBNz3UVZQOrURcJAe0cAVOGMTde6EXszr+vcvLDOS4/L/vXy
SK651qAD1KuP5OqH6h9VnSZfDOVRBgnrFnsH5DVfQzNahStDd1CGQWTDo4/e9fM79ipCAB2cNykV
ZXw8I0Pyf09lMsoznDyZIRpYVPbuwhOI46N+BP/4Ztilgk5bGGFtCstWS/nlWozhb4nDwPKrbpsc
FUidFjvtcXNNTgFo7GPac8qrD6L9I9jXJgQaZWp9SSqs0VFCDrMN2qK9QbZF+ozXjCgUp39Og66V
9xkP+Kjhw5fg+lwKuXrkgSkSiPEl/yU/cLkBI7osCdbxFTzqHLB202XKS3O0LOxIUJ/MaApPPKtw
CM0AD9rWU2pPWiDxhGe2G9xsMp52By1ler9JzFkNUXb8I1aAsxjfhvNGXVv4IJeqzctCkD+GArRP
dul1ofGf0ExkmP9DMbrgRFOHqZ1CrCVjSkvZc/kOThWS35Hbl2aGV43VBJ+93C/Wl+H1C2NGnLSu
1NwfDH+LmYwXs4FQToItTtcLxH/XLucuzbsmRRZcZ8x4/VYmnImysftrxdsLc4H35MHuedI+kv0C
gLIBxUHbrpCHGgaIKYSPz8FuxXKh8gp4Kl27TGPXeT3L8cGL2CcdxYod+HGq2cMnRzzLF9wQyomi
wo7Hs1q2rLKRO8yJGzggqPF120k8+4WnWYxseKL/P/2+F3hSKWDqQhbCcFwxMuruFvXogR9ORf6t
aFS9MliG6Zv9mbk8MSUp6TYBOCAIC3AL3YcS6FEJLENUCbt8DZZ9pvlRUIKEAvqeUhWU147Kc2Tx
ZzE2gQJWEygIvyftePPa3KwzGHn83WA7Q6/Z1eC5IWNM1asah4HwO/0dnE4IgBAAqcogfJE2/DW2
3gT5Jr8uXT0/mnPYBCiVZqciy9WU0UHgWqJAL2VhdjEDhGjNJ94NUvw7Udgu2gRCJqJojjyF5mkX
RuAhtnPebE90hj9vnpYpJ8arCv+5SCqR0Upoy/H0rxNqm+WZBSCEQX35uCq7XMlxC/wyWtuVJSOw
l6vdPdOE6a1QRHYnvAE/Ann34UMlJM/lm0BeS0PqN0mVd+9rf68i9KVDQc3mXN8UWvW8g/IzU6xR
iT04U7Ua0q6koLMr+38jHwjFW9LLX4XWod2/0ZMYE0Ssj+QGaCLilXmVT7L5Gwpz+BAU9QzGqyJR
+YtycOyKDf8OQHUqTertS42iJWf4YDdH2xb0zomqDUJmhGTVopBTKTvZkO9nxcdtAzhn7N9phYKR
4tqhz1jJmxJ4O+c7kq5w+ifnEJgZUyO0tFdW8VCiMl6RtukoPAJBrXsutBRZauLfNOYdxnpIDgML
tJdd6r52c26eHq15+CAWdJ5NjYn5g5vW1uExoPTt1jNoMGpC3UYpOfNvDQF1e0j3Kl/aYTKixe5s
KMzDFquUy9W4EjRuQGF5KVByDadiJMTdOj5VEnnO9s/z8WxCOR61uWI0Pd8FnWtTBcBpbK89mw5W
1fKT2WVrIj1VtvWJuKxQiGQPFjy0iFDfrimjd2XfBlqPmSp+qaxJsd7SBj4AUo4VXMERhjDlGaBO
GVMIBvoBg8F73H+s+QqzK8JaTShXlZBiNLz32lN3+Ro+WqiC/54T8uHBC13TWq/RcDegxcuJAquV
FLJ7h3K3l7Lhnhb1Qno9QJOE61/NgYwD3kGbieO/G0EWOpWx9paOYgbEc7M6WTAlDocP5zKYp7yZ
fp7Fz+KR3NXsZmW0cDaO11pFNWVV7zCbATgLqo9YAqgH5gVFIHSq5JCnqnRU/aEiPmZqk7nCIbg2
fNuA/IL9EUgU8H3FTz0xunYklebwXCyYkqcCG6aZQpzI/KbAztuhrfy4C0LUCiPqkJK6WYlMcO15
lyIXDuqMNSbBsOwLlpBTpMSNcMEm7FtX0ed09KnZUwgdy8u0xS8zjRyGkiNwrBfaYcqmNto5Ce4N
iVoYndjikVsmdg2GupnlaEyNk5c0kxPYI/Ay7hJLY7a00j7LuniDdmXXUvxPixBEG85aUFoS9XjV
C1/XpZSuN78frLoqXoq/Ngv1OBJf/lqP638E7bizDdgGYzzBxAVrTxfhgDdJ6typKGlBtJee/asS
yXlahA7E8JZ2J7ZvqCby6jnLqMhOL8CI0bZz4gIYozEEgjgi3Ufxl2m10h1H1DAFTBzFiu0mx2Nn
X2f8EtAT2bDFHQ4uZoVJI4jTH4yF9aL6lSPzWD5FJW7wudutiGBc2Fmm9Z7pR1eURBQmPm9fmude
yr/XkuSql/Ku8ZkKoHlLwKqOZtTQWsQ7ztUgms+3X2j0X/YLxORHXbqwvNBZVRNA5QJn3cQENCDx
cYi7+wd+8jiyajGQ3TkkYSSp7D7MfxbkWyY6JvzjjeozKtLMHirL11snQ+YGky+6B0/wC6z63BTJ
amQQPuiDViRejGFEuAMvCONRyF3aDtPbytPTDNebF+uqYl8BwaB6w2YaZtKPaxEUyhAiaFd4KN41
MobNSHB2CxVJvNpeKkysDC55BCC8fbaaR3fFdf2MdrnaRuvhJjqO9TArGuE8Tj+OWlHgoaua/ora
CE7GGMeHU1HMOmFsgnBtxhF7DjA/jJ3juU8yHioA2O+VHJYXVWQa5Y3dAG3mareEpaggNiNqQ+wQ
/R+3bdyV2rKStCFIItFyAptnV+ZlGKsk6jYY8RInOOf1/r0xQOhbwqwRhN6ig3tNvT517DDyab9M
JJH//Sbyf6sjZtfkvr+CTRW8PGgvDJaRJHliB9EWpoNzYZeKGou3Z+10UYQ4I1smCvH6PURnf4Le
B922KeD7LKTEFLTizQgIt7ku4yCsvnWXedznw8z90nKp3RIME17udACFDWN72+c2LM5Tl/fFzD5v
kpNrbR6oUkAHz0Kh6duSnDbvX2d6QUSOz8Yzu4aJv5Dt+WDi3X2Z6e89a/ifsMkCvD1y8tcLZ8on
OSwsCOkP4VCaCatljn+rt7mPRt4yn6dm93nGw9h4pf/sWIhRWGgcBmrs/XzItOaPj7qIC/GRfAK/
t3uGm2o+vNmde+kb3daaR0su1MNE29RBEiMRzEI/Nah3CfcSFRXeiisWBAZmgThnYoeUSP7LIIUF
2eoooIrzWM/v+5+uYztgFzIbQmqxE8rMpD5DjGgNaEGOptQmDY/LzAWZmA7JXwd5/u65U7c7hPlW
Eii7vI6TXL8i49ak5uG58S0yhDL6aXKvHNgPO8/VJ9OrZAAxbLwF+YGZu8+7Wa19mD4B+eXCoRtf
bm+NB8vUWUr1PrCi4kn20S+WJgh9ebAfafYdMMbG8EvRim5qomHVe2GMQUxezMLAHmACO2nhoKyK
+qa72OTfu/zLKc72rgfrYz3AYOt95h7ILySYx3GOOAhyUw4g4d3GZUa2KkjpjrMPILYNCXjunfj+
RqgExT5TgderuycR6WA70edfHaU//02mcJSGxtw3pHKptBMTRoFoXCP33ahnmlzdjAT1EJ881G9M
CzhZIxhaHNe+W1rA5dFDeMJ98zlCemHnbJ5DcjPacpel3DoqN3271S86E/Clv/fW6CfyZ57OgkQv
L6uK/L1Vein89feGTaBt19IM2ouFkhQ4boXJwHhEIfyv+fBwAlgDbEajbJHlxompnq/SPy5P/vQB
6rUm0Ioc3FV7jFgzAeCs9xSvEgoh+wFeo+bIQiEYXr2cqkwJyzsQ+r88WvQIQTGB5W8BZiZoMzuR
88vpcHcw/cAhODh5W8JDvoChYPSUV2faKuMV5zga0abxQCNDXKMw2vT201PjkOU6JIB70Sw3cD85
4jR7+929aXRRO/fsVgTalrbu+TKKA4CGJAbtoHX8uOMIa+RkBRh1dzRlCVnkHBqXFRiMAIisMFGp
cgrT0GZhe6RwJxkeKxJ511DejYQGYe/0d1uetPoDSPj1qYLzOQPu0hkLu7HGMhMoFW0LIdYBrmgH
YShbu/bBsUhTixiM2eHERgNOS0i3zEHKAa6YNGlofgJXLt4q09OwiCOuxCmpckz77Ir6+ey7kQab
yPM4xK0IcN/JyGgNGWnBYZ55OZ7m8qUwd51/XqxqnHQprGu7q2kh9XUI9IxzFBCtyDoPLD1kgoOj
jfp0qg6hOQqJXIOSyzeILumZOuIYQaCPlirVk4blkrffr065SpXUH2aeWZRm+ieLafoki1qu87EV
EDe7Bu95wMiKxnTr5NXQ7DAVxIzK9hgJyEgzA70GuXEnjBiRG7VUUyU/Awt2l3RgoRvxZLcFbocp
iKhQY8Cs/ykA6as6MK1fF8bxTmcHGgwDJX/SrrzccyTRAR7GBkvHHYct3A8t5XJzUo4uBNjKuEio
icgM28xW8sclnw0xJPVZzAegZW5j8Lnn4MSs6y5FUNzliDO1vTRzCMz0gZP94Mbx71guY/+8mWda
PMCy9Tp+z1LIi8sSiC4xwh4f8A0m3vm2pJpr/8tE2xAgZyCa0Nn/LCXNtuwguQuMxm5fhG0/HHFG
iVUfvuRHsd7LmM9YR5FFKXGcDGkVZFKLM0yYznuWMie9SfTrOD3Yrqt8CG0PXm4kIx1jUSYYywjf
XJf/ycyzMrMWW+KPV1JevZDvd5owqtMw43oVqHW2x8W2CNAH9UdXDd2MKt3KP9Ra9YNNCPBxt7Zs
9zCEKs2rMqS5j7AlHLd6y8nizK6qGoP2Gs3dsx/wc9UB0urOv0JsbJnwhfaeDDBngdiKnpZfrtXF
ZfPQF5hfMm7rboqFz/QUbOPXpVHlhaUP8AAjLqb1Eco9ho00lWae3xRsPmPQqB5cajgZEqWhTCLt
l4cm65nsaw2Fbt8qX8z5GBCYyu27C1ezoU+yHfrfUNV5FpRFyTzqGCtocsB7gt5i7X3ZfQVTOdYW
4Cr5Eoz9wmr/dn27Z9QH2KqSXxeomLVkj6yVNe05dgG0JxqX7zlb3RJU1Fhau6M8Fwo3r7qujtB8
DC3hRl9jerU1a7+s6KarDm5NgizfGlkOxXW2ooOTvvDmBDBsBJVDAksHe6XaVF4YPnwNBTzvhsaQ
efuG6e0wBq6E/ueyTKjjKS5GyiIc03oMOwj4sskGa5X/TlMbX8oMexHjANTU+opSrM6GtiA47/8f
Wqc2qJvXXzTw5Aan6jxJg2LPlvig+0plDQWIKitaN7uqPs1YfhnrNk10mxKXx4NN8juq1kVw4nAz
2KH8c4vQEOZzFTUQvWQJcXm60rPh4kUOQJZV3hvksBUtJXw1TB+Sq1nZebkiSajSNuc/APaX61HA
UWI/RW0qG7LYA+pBhI1OnfXCN/Dsawhjj/fXOX4BDR75gB783JFQYvx1ID1e/mC5f/OJY8t2Npd1
YlMwcicd34LpaO3AEidD6BnKFBT9J16BkPPRLiuEv+oC6qqcD1h3DjvMMvxHCTBC1Eb3xu2CSvSt
Wg0tjk2ycAFtgLrTFBA2Mb+X+u7AfDkeW7zVpVBrj95GrSgGz4rYbqaEXCqjwD3d/b6pmTfaO9WI
qavomWsS1nxLIOB9pmv9BZ9Vij5ecNNqL1RfG20BMUpbya8dH/aUsBmnplckOCQUJ8sD9rOEvBLD
q6y46O/N9mbvlZCrPexZHULWBALX5An2NRVLh4v47Vg/XEaLNLD0EVsb90I3NfJn5Oo2fegtv4Xs
xOPkhpo063ZFFhr6+M5eFKNP1gunEcNALnexaEsr+9JX24uu+Qp5/yM4MYOravZzArEznQvG/wZW
CGFxMOxh8lXcfEC3PRWgASbo4TpUaFWuSErBJb4DwKHCdoi+zrThTKii63l9OJtiCg13d2rGs6vm
kGzBZ5v7QJHLV07WALR7TjQ6k8IakNLuh9ogQup4aw0omj1SN/QJ8IQcY3iAIVT3OeAMw9cJtUue
jkUAjO2ypu7Ls72PDZWYmeCq5WwZG1qN0o6zzNaIpKR3e6CV+i9hX18TiIpDRh+pQAOsrg/8n08G
9b6Y8fPifTpM35dHm9Flu6i0cD29LCZbWOV5wTzFPJr3Xr72IIjwa5jiSI9I2/8P8OS+peNU0lgW
ArWtLdWced4sHALFC+ngg/X4zobDhbnnsQU1wjCjj11Hm5fn8DRVL5PJ8Hyi0fcwBXT6ivO4GfKF
S6veIlF8dh4GUToH5zvi9/Z8BQFT9sps1ANzGA4cuY6i8QlVOjoKGwRt1dh61NZD73aRyXLMSG0r
aKGHWYlbt0SiEzzl14lb8T1QRpcSc4U8zvlTEyjOgfuklWmAtdIAqjFXWuV2VaaUMxhVHFBsNiDO
3W/t9LFtciWh+OGJB5Vy9m3bpWkHqUmuU3vxvrKrm4cwgb2+4ahBJ1WGhA3oUevo6ze0oduioIRv
TfB3KYYK/3v5O1ZrXUYwcmd5HXPIi/vCuP5UvJLpkDqjDnGx9Cc7qbW0mXqdvaXywdnmCA+mcIoN
1bPcqvny1B2Mohk8cg54lPG4/zAyEf+k/xLHVi9sLotxMecVvnSD/TTo+z4Ssm0jb8R6j3UTiQz6
Sgn6Ox5lD6waG8DF7Jq0XSgtIyQWYXei2//VQ0hqLGkJ3wWPPmk27ZsefpYL40+RP+lFOJkosnBO
lbQE4ijbffHn5l04lL3a/V8OJDE4Z6PHMg24cARh4/HXE7rM+c0dzVHXazuCtNN9OfplU24wBr1L
VUNY17O1m2L/RxD9Fhm2agT/8Bb+DM2O0qrxKF8OKXE4FUmfkVBk5m6ZDntcDaTJ1hFUkq2u6gCm
qOcju4USQPhORByYyTU9raayHH0+J4UfwfU64FmaFbgWSbOJbhSNqlYy3OME/n6LJ7tKLhKKfzwB
QnbAkK+ER3nJ57jle+0NQR4Fyja/ZPls9SXWnIgh1CExA4AbpMPEMGvq+YgQpDwx3lJuBydD8uW7
Oo5HOdhRE9aTHu12VNzPKDDq00mhdPaXqRgkySlpQEqsmAkhfinjD+hgpcGgxnfvdRW0aa2+69UB
BSVvmLd8Pw/odgMTgUZNXMOP+R7ep8TNxRGHq/KxvJdfa24ktlBHjZ22l0icUaioZP6lCG+DdljS
uNVKl39bitgOcIJhgbpZVwqMHcPB7/m6M84RnNUttiSFV64J/HkIbnpgTKtoVlAEf35hSUGpYEod
SFebygCQ5paBeMmASDZsQHD2XZR2FcIs4qnESk8yVKAkNkTaf4+pfMPR74P1MWz8HwTo444a+VHS
NQ3enwRvDxQCpEkVAIQwWY8xkTR2JVu8ozPWrIiy//l5bNL10Y4sF8DLljOPVwiCntogLBEHZ77u
p93/gTcB9sa5Z2aXKMAy3QTWHf+T3vgyrVphv0qLaeYaUIjYTdJpT+5uIcmEOUyh33UXYOIfbWwI
6tiQ9ieaTVRlM6XthEzu9SU/BbdTBje5IUaQ6wFZhB7vbx5rNlZuWq8cTf24P+g15rQXhsRhfpA8
YRm+b09yV9ZNBxsXEbwoCK+VzKGQEVLgxlsxWK3rKN8zuJy1YEvHizLSZu5teJP6iAlQFkuo5lgs
uUDPfiHrk/4X+dsfKH3Y3VlHqRGVrBI3o1MTOWKaGpC6VyBHIrMECKW4fnuAEeZuIj74t9zWy5sv
c4oqfv29HOnINzycjkEknt7TQaYZFJE0KWH2s/ra+KWbgcnXS1y06oZHWCyvrgFFsPS32xo4Fgqa
Ko9RVtJ8axz73K+nKV0UmPV87nc6iXNBEb3KdSQUWhKojwC0KA0sBd295aTUNjXmrBzVRP2u6asZ
zFBuuMy1kbZ0pcleBow8lRwE1VMxTRZ6N/UZ97CLoCfMOZyuA5A1uuZuJbkdFyIhwRw9Ve+B6NpC
xIuVIBEoUiNt3KknI5K2no47A+O0JGdRD3kLAkrLzTrso606450P6iZyAUjuvrzDAKDg9YZDfElG
hooITnpOnwD3fkg4u6sSiZn7h/ONUXUI+WmO6da3wLKD7UJlSzwEPf6pu4XQzQCyJLTzvqS57vI+
FFiX0gjwibYsvU+O5WMzWbVg4AflL5V4FZ1jK2NYRc6RxvKCnwPFXYjwWfW7AbZE6gqN+aDNyCp2
vOaOIzpfWKGQACcmaRhHdODAgQ2MVctyKMabboaEr+oJERuNf9YgQIqBp149ebdG3M/kewd7/F5n
UhsKzWJCYO0bmTwRw6r+qImmx2ufHbkFwsQb6+vL36lFp2WbcadtjsTS+fD/RBXyDyDXcATDwK9y
hSRE8BfXMuGI6vb3XRNTZpcQVFukBsgUPzdZe3iyDjZKH+nMbfHIJmRgQGwA+zpXWBJctGeZxgQc
Ft2/txKrMFK+PP1he1ZCEIvqUb/50v7ZmGytW+ym9VyM7XH7YfBi1UX4KkErdR6YuEQdYfjI2qMX
9ve8k3ozZEaRv91sD9R+KSYhVcQS70Fo488+z7A/nJei3FYajfm5qwXnH9h2UV/kZTINbtb4SP4x
SlvmMDFwcSag+yGqYoX66yz8Wa1A9uRdtLfl7fL2Q6Plv3IXE40LHIwjRbCqNMUruFneoLsVhud9
898wLZHZqEwnlAI/6uM9tTIxB9W6+Idl6Fo9TZ80AGYA6abiUYuq3a0WtAX8Kh1PHVrTwQpRRwhC
+bqc36OSKD5TxJ83m1vZlxy2QFs2Z12Z0keH9Yqh+QbDMf2CAqLp6AIrCZNM1HnB5ajLwCxp9xNi
KfL+4lnEojq1kG9NOF3P4d+KPNfZtxewu0H1RsEHG72m2A1KeSCLzfQG32A7EJFfgi+QJ2Gqh6fX
+jZPgIhzc5UQn65WsTGHln1KkgqxjKlwZRend0PmKTfuaplDB7uGmtQjsfB2OozTqE6GPc38HaBU
exceLYsSvV4IGWfna2g3qwAPD71TS8J6BJBfqs83TIiV0aQOfy90N+uoWDAo0crDX0OcJqTuqRMb
KgIe0F2QukKwPs9hVOlQvOQkV9aLdVvcTiQ5AfQMqUZ/zpAhYSVOehjsAUP0kMJT/GWtdJhszCtu
AcbzFsL8R5EWOtuwFjGNFI5sQRz1kW3nMfKGel3JigNyTeK95WCyy4W7KRfe8vmVU3EfSvYjRSHK
7eHXlRJgZ30BnbldKKAkSQXRX7C+mbN6aBTFCQ8kYqJhCChFi5wPzAS1DcKZ/XDfDNwLFIydKe9J
QQSFDVlhRv/b+G3eTPH9izXboz9cLaEDyJLNtuGZ9V/HEe2lDtgGcJDGFWyxFZmSoyD3u+BxXtF1
1o+hMud81G6vWFHPKUtWhN/Kf4WpHLiWf6dwCcfqJwlRzmPwGbvYENQTnaBhlulsRm3ANIWDYOV9
4jFu3FvyBfazK07XOUpfunJRjX7qe6W8N0eqeRoG4hDDU3sN38Uex0YaU0jsh8E5sOF3AZMh83yr
ndSvB193mWCzgEMIATzUzOahPhKMI+UZXe9uzeDDBy3MF0sN5A2tTVg7vZHo4/EQYt8MofsjbUmO
txjeYEpihCr8XMgyhfX8n1aKXdNx/evFP198BKvsU52jls4N0RouIlN0SMncFPhvKZ1vbeheE9gv
ulAkZqDc19IGQNQ1tqGBf5oJs5RWkR6fIE/FxNSa5xi4k4v7N4FmShKhL0AXgQzUEbgk2+QFmkuZ
lYp6LtUOK35BAg+BjypkM29pkAzoe0NZhdtt7TP6Phbvfb5iwqzKeXuoHCUNBFdTsRh7ywyHwCE8
Q9759YTXA/mNrr/51fSgmL7vjYYseI4qbiGeSRDiAda1wMvw2FxkPMgWGgNbfwH3HXz/XwkDtmHt
aEgBqOLndvgXoxZ+1H+lBxS2o7QfTP6Bn0lU5RTMt0FG1dvc0bAAy6mOvvSJteJ8SpRulIwUtS/w
cJoTRPuTtrnUdfsxPoytxRA7VI/UIjMEmYrNM0fcLNnDrmX8W5lDoYbjwyt3fP4ChAZLaWpLz0tK
I0bDGPHb/H2g1EU6Q6qyLfYD8LwaXhjAwPPpk6LtsY3mbYqfRjdwk6/2n6+gwFmeLYJOJOjF5Bga
qxg1v2VZRtlYs6o5o2SwDP9IJ3ZhFkpcxZ2lPtbwRWgRdENlaMcrYo6tAV1CFeRnreS/Ymri2EL9
RLKLVxECK5YsyDKzXyF/Ms5QoUQ3kLyXFuAfVSkuqlRrpGpqrQ0rOafPfFbe+M3atnq9vdhPqSIi
zH6ZjOP0C3TrkLIP2C/7kkpT7k/71FTmCuIJa0VhppRisoDiOS+b9kWWZWCBCZ73hy4iBvwr7AE6
wnHtxO7Dqb2s9NltizU6S0SoSzgkPaOpK9f6fvq3Af096NeT4p3w//fB8tUbhqvEvR1mMsMFpjNb
MSqssh4s+p/jOGzI1DYT3O/gGsVYfP6pclw5oIKkuuooZa84InPYHzrIVE7YlWcNW94GQU5TndS+
BKVZkF+MrlZinDfc/CsrDBQ/T8IonlfwubT/AuO5iRCb+u8UrolwZ+r+Al6Qw14wZO0/Vlog2zQ4
Bytok8DK8XyBcVjb3Y1RwonbjKqLBg3D1Yb5prDb2o1A6OxnXwSijYiqEDjlsUUYu+xUwt4lGpMh
14TH0o5YDven12vHT/t1G40YM5LWbByYrDdjFahzjcZRg80ch3mgq6FIlgvL1pOnZ+tfCzxvFfYE
lnWww2IxH53zP1SAepbF7VzYA8kMzb15be84zu3yq5hvNFjl451+4MeZdRz3uc+DDwYig4roP79W
qnAOkTdSXTLLvP8q0zOXWA8pDgQxmdqnRt6an8uS9a3b4WXzSm3JRXWTHDibQyrUWvkh0ip4k7xc
eDo9UB5rY1x+1OBlht/Tt1x2Ds94lQYUBDYILJRNBOSo70t2v1FB3a5GEXLyK6dwxgozlV36bdRB
2Pm/awoVL2PwiUG+8iLuDOqpGycWG5L7XL0K192dM826Gn7gxG2qeOuE44OOX8YVeGqRQ1MLcEY9
xHWeBLAjEKc+kbn3fFtOU8bTAWc3p9yEcMx0At/SQtxIzmHF4YiSW5kWmBUvBeyiAJCXDmYAnkfa
5nVZ+rR2F7Kl4fwPE4IN/WXTDZQ7YQJSkGZ5sef7DUIIloevOr9zVz6axx2mqSuIgjLDxTcYcBxh
7HSHfMgFqkgli7rzBQHhPjmrjcbSBSFq1JUHKrXSTYc/xVg4fU5aPs/EN+fNI8ZLQdLdC7aw+7R3
Xyqb8nG1TN/J+HVqgvLUL6neQi9vmGwmHkKUktglccSPrDfygqlvgcpfgrjV4nxjxcHaRPGT5BUF
yndUQVGY/btcAAaav9q1aev3zDd3g/uAb1qn3vk5ZoKqQ15neFIwUVsR3zDsQSSj7kc9HnkMzD9h
bfw8D2kVEqjpv+YvFs3KWCAYK1BeXReCsmkYjcnzwxugSF9yRioZkPZliX+0bjh/DDU0Gztcpf5O
F49tvggjZ1oXSxVVoKnt3/oUfboU5rYyGBYOmQVL/G8ue6tPymPXRmUM/k1KsfK6fk9vHIi9MYW3
su0rjLB9uhme7HQ+sFDMHBqnXwD8LDedRv/WxZG6y1Aor8eJPjNfg0B98XUYSB7mU5cQSIftolxO
cmzhJFopYHHLDqp6H+Xmn6vTj83q7zhdCHpJ8mDkk7IlHAMSs1jMjGWFo3mrWIdPcfLMpKZT0LlZ
H43OACxg5MPh5wTaZM7hpdyGRrEiQpbqaNgIeyl6BzlP7q9zek7vrVr7MfkFI1TbvtXQqM5ImUSn
h7pMFCRq+Y7C3F5XaduLpZ75M5HzxzZvZMXEJ/ic3YDGE6YurP52P5G59c7s3EyYd/nH7QbxyeDA
KPk+k9rgesm6wup2EJbLG/zlouNB3IQZrrLXMjPITKmHfczztvlqN3d2JRlrFLvWCozzdl/2B9w+
QsYDGmVCx4KiZTfZfmeQf/gcmdoVrddi6GV2Gv94MwyaYAhksr2ag4XGTT4QA7LQIZbK6XZCeGPr
04rX7kCgeac/GjSjVotRo1oABfETQmUefCphHjQTYLqvGRKDLDCQS9GcC/tTJXfAN8pBtu80Jwjv
CkC3N2IlEWq+CnTDG5Vs+pyQXl5gAm2bEGSTRmBz5O4N5wQfsRHpT/GuZ0Eju4FTEA3c1mktBs5+
ZqkKXHg2GGMuDLQFsUNpEgkIHXNTh97HIQHuro3INjWBLjTw1QCf1BejiSDaA832qocEGjPHI4C3
rX2rNZCjxzfmU1xhzS2AsYqp9Gt+SFMnUmf8LK+ASmeLvS9eOF4EYBfGOf95ACNxX3pquvjCLaSU
OsTfhOIJFK0USEKi6tFAnkhHeNKrD1b3waLCwUGa5kRK5LTzweMkdg94Vtb0q3o5Flm1wo4pzDYn
8YTiql5PyDqwaEUQbcSns+ItjllG0pUwCbPpZDuwnJPCguz2OhCQbaTK721CInLwscsYqD/+I50g
82o3b3UQgPYMIC75vYaDYNjkO9zASF48soLXsn4f/Nc358w55CHezMz2u+JaDnxazxpcJKvt9oM+
xqle2mJx9ydMwM9lfFSPPGma9YGzAPeAraSs4I9veon8HuugJ80MF4BgZ6fmG64WmkUVNUlAbzDS
gX67xPpF98vAmKFr5DnO0QwBdLQOglWHZBX5Tcow7PE0p4BO19G5NCWi1KR/Hrc5Pnu00nRD5//h
emmaDzj5B2IQA9s8uP1mSDvdq11wexX1sGavupq2Nuyw5Ci1IqE9OYrAfhc3viTwg9JnTbEWE/2L
pKuVATm8MxTSr2zyQFzr4P1Ri2dIWtcNQcn+RSbeTcvbdkg9UDGlzS0MTZMjGqIR8RAPT3VimShW
5gs7qfBB/zmgS4p1SIvVEpGqxneIcUoLaGD+Yzmt7/iCTTx3tTFXhwLBq4vArlzJM2RsRQdIeHbi
hJ87iveMv9Mz/sINUyVdWMC0ioNSpUdroktAzD8wIgdY7hOERxvLchdu3FojUHmYSleOBHNG8APu
XJuhW7Fc+12FmbN8I5Agxno5aflfcW0q3LbHGEV+SRhJOkSvEouMIB7eiiQ82HkGSHvxBXWcIc55
wyyuBJOqXoZEdaPNBA97KsXdVxgoWXKaOZ9sh2yBnq1NNvknJIZuTMwgkJhheIgJhbh07rkztjkk
PIXpR2ICpzZdFCuZca79ZrW7xMNo2UaQGdB6REgcckayOwRRW//c3O7LJzeK9M3xRjqrF7lUimWs
SPZyJqndeW65WMUiPR44N7kkFG6xlbyPH5FxR5f3hcTlB7QmAHEarye57Kt8dqUJQyRHu1WmLdxB
u83qU+pc1H7a6Fckis0q/+yFtHUNv5nsNYF2I9IK0eMLQpksNdYqYHGi5aQje24dHTKrXpRDvNYw
CW18uOwg9bMT+ysfJsyfop+xXG3cgVepuQ92/wQjIyi6sJ9na5Uah3Ehvwq2eoDEGOjxnQDtB047
EK8yVAeFFWtfqv3K6Opwg8gQ/+S300IZ+QZLGG+0SbxNn+6PvXjVXAFlDMgv0Qnzg/2ONkfZ5EOA
uPEwP81S1RxyPVytEcdNtWIUXJ5fIeHeiFHUNkJMbixPSkLXeeDbIKIGjiNvS6hdKAxik7I325Pu
/baDlWGh+oTZ7121q7wwNP7qt3iWiC0/U9+sVOHgKrEqbjAdTjRufzr5oxiVxZNxiO4tS7+rFvRR
+ULh2wUTyq2Li0UzXzMg3y+gQIDRt+XdYYXU7BBJ82pevfNcxC1YGhQ+F/nezMkp/K1f0svI6Avn
GW1NdTFqfAi7sH2PVAiNnRmyr2lv3p83KYwKWKKzxulLzehw7v/FQJEgtwHqHKvKP3OuRV2Df1ZL
ViTqJGHZJFgGuUY8qO9g0HqeDSVUTg6Xj60dx/DicYTQHIBBNvK7I5rdl9Seijb8BZZyRzGXCodD
SAq97BWyzmfw+o2g5pVs0a0HVelU7n3Wmez8eWmkBMydbBvBsAg/SFdmuqxDQKE9XLPYOgCQtslq
XsTEWye5b8+Yku2XyzqkVFZQZDmN+5F569xmVAaR9nFseIVxqOTBQsLijCssB+VGQdo6Rq7jDSh3
1+WPeId15sK6ZWUWHV4XQbZwbFtdArNn+SRgn7suobBDRrJ8CobuiXrzj2VlBE6puvwRD31ZIBzG
7nG5d+ytlA57pav/ZQ6bKyHQj9wAifexroAqSKz1ZP/0uGMIhUbAoMZJflFxKxZ4UeuNqQS6zqCq
W9LD3/NHFApMRJitC9HEZaR0e0GVRQkHLwuaKb+vic7EKZggwRyD3RcDxGeSVnJjmw5UgFVJj6xa
U4RdnaJ8K9HfhUnmwSZS6VP3i29rjits9ZO7z2cHvAFw7BB72e0yNNuhdDLWtUU5u+53HzK1yvXY
femRdDh6p2qOhvTc33ly3UBWsKgsvCO6wdZlo2GVl18nQ4YiKtXtVPVXicndzRVUo3lj91dRNm6g
jE4QWzrYO2RGJt6dkZg80GSBa6fA8GLELpfDZMbEwZ89zyXPYsF6NPR/PZydQYno77YLbxVCM6D3
CMvjlcmuIMnClzhOeMwyGYx7cWizdTb8YTkz91J+hGWEjRBXJ/p3h+OmUjJPjrVYlZVbZZY1jWW4
zYea3KkouaxkpXm/D+uzlCbGIpD6iORI+bYRPbhDDw12OKr2TbXezN5U8OjSqJU0dsbk0KasvdqU
9ZnW0N6tPDsPZx0K4R7qR/nzITYJtu/MlZ7UTK+mRXlWpRHYS8pifNoc97SHDiDQz0DhmeQm/xd7
SlJEorlm9eDqZw4gP77mQSLHDsoRIrgvM3vBVE5WI2qnp8tag1yyxtaDEfet1sm3xyOY/4Lb3Gu/
wUe3XEZp2Ne3mGGeRzK2WhDHnwTiH7BzpZpVCzJWunpanMqqPpQBnYvj3VRi/HZvpD9fssZKBQ6c
1MtLg/mZOnLkWexzAi6qbQn2wrBIYVA8M639LIn2Qh6OQyXKAdUZSEtsdhBa9i4a3eNZkt8avdYp
pdHiBFPNnJIbcMOBEqz/b7+aYskE3oqB98wBk2HtCvo5oBakAGyAF/sPsRsGnN5z+AVqldGttwES
LtEkLh3T/GXZGMF5V3pNT+DBNWEkCXgxp3uLbeqIYhY37B0naw3dTed2Rp9idPFabSFykBlh3MYo
l4mh7NLxCyk4RoyteiHFaCe9rki+zb6mUamgRFPPwLo/KKUdSEUaWAVu1wyaA+MdDgM1B1Lio7Xw
W9bHs1MYpik/txj7I0CmgMnb+V11gqCCpNrxhgIr3u7WFgQEJy+hzvXXHcIg+1y/nriAfzjq+BML
6PGbCcd5AfYkhfdx7wokJjPAr6uttycFXKLmhg7nYMVGZihDqFFTQ0BeDvoo+9BRPkWLzCvMkSzM
SwzLxTeGt5Oq7LQpumA0af2cSLW8MjHDMpSxvGgWXMH+gAKRNwGMWm8fCAWwpbAWefvt8gkMYJiV
6Buq8jxQeztzMeKercYvMLQuIMHLLaKZXOJM5pGd2o1SgcZhW0lKAf3LxpJ45ZkTmEbJl4HoskDd
EWGr/9KoWkLwcCwvcM/WZlL2GuRtJQweKYbg7i3NLKMVgBt/xoRKSXI83OaN0KJaqkabrHUj3y9W
ml6/i7StDjkiwEIqNzpExDpWLHtwgNIBX6YpGYmETF/rYpL69cGbckoF+Aw75NOPFa/UlAYEvqk/
sNVzECdjmij4fy9ukZeSu/gorvW92/VmjRJtBXf7tH34eowv8Mp0KzIPi09Eff6SmnGzo69KNKCq
/56qJ3G8YOzl8RKIe1nm6uz/6rnkxkPRovmDJHypnfn57xA3/QvSUL5SeKU/A7/eI6l7ZG1/ZxMW
L3ZS3OZPP107fT4fXQo94m/chHF1qZf59Ri9fJy0n9AeFaRGOYy0TyjfvBo0HAhiGndv8wYSs1sC
z1KJmx6OFkEgwBy/hHdAUlnDbz/mSO3GOev/nqWmDDaHTF3rKEuW3ULL/jTB40IdBBwnPixqPdHx
IIdQIQNzpf9ey2J8yovp3wNYb/610+ZXdcO5OFQ699bDit7nQkxZ4NEG0+GMVsEKB9z2/awBJCD2
GZUv63OkVIZ46K1QD7qPO2fv4U89jHlM7SosK1RcTdpwFshtowBxlkxQnaO0jPIm1HSDtPtlW48O
OrlVhlKtAPll79044VvpNk9MB++OV4AFdPvdpFC5k09gi/gwur3oOgJwUBf+ffpeD2bG6jE0TML0
3t6fmjoI6jLnPven8bAWttEgMJUPtRvgAqPvKKSA6wJKHKUDE1Ac3VSYelFtJN4QeFAeH3XKUCwp
8ojXjK/6OURio8jcVsHnoh0fBJoBJzfhr/6BT37oAyhaOUePlabo2P43WHB+2tbYSti5VLude6ws
NDS+tEqKGM3JnOqMclVvq1EqFVFAmuyk1k+kiKDSVaw/8c2k9mpNsyNSI5Ik0dbH6nVxNESuUrOK
DO7kl8SNoz4W2lrmxo+md8e3IgwWnaTI4pUQMQ56U3DwTP8zRShokBpmGEpFOiWDVpeRVMY+i+Jh
CeetoP5/UVSfqmg9FIME23KCoNBxwEKHB363TzucnojbUqdlQyz3wwO9PpTbCOl5dmMDCREPMI+n
4Zetz+Uy3pr23ajeJ4eUzE+hTsqXlFc6g8uwEf/wxewY8OZIFn7xClzQ8K0hEt9uer8fazEBX7vR
hGsJNyb88Ws3Sa6FbB4nnqN2dtFIx4w63hDplwZCgnE00mEcFQ/MPkRroMGLLMuRRLK9TEdbWKa2
ivs/67p/QJNv95XdazuKY7lpbqsLF7GHo0tEqmY5yjQe2JPS3Wz2fQqlEQnu82fOspDB8Vi9abUY
pZGzb7DmKFREzhI8Bcj41s1rUEfiZEQnFg0VgmkVzD1bChFKNxfH7EWG4+uqE5MtJWkHPh25P9lA
R5UxlrQpH+l+0jYXGMUD7isU64p1Cc6b8VuUA9a9nHEJ31zHgxdw7n0z+4IJLpNG5Qg1QGhfKrI1
SAJ+5ME0Pr7AipHaUPX8dQcC5wh7qMa6T3UP6bLB83Z7PegNedTuia4abyETt6+wtAATe62jMvvw
Sk5KhBoSU7kRkyqJy8OlzGS13MlKnUOTjelIyum9UCRQzrV3CiX6qcSYo/WuglRbOcWNpthj+661
lbestAPUTraca9hwyzBGoQsC8LTkyT17j8mDUZN6jG7YY15I+6NqA9uCsfz4VTGec2R5n2j2jBLX
+SZuSHKq0ewMEU4JjCwEJP52tBTN9Md3ZjWWWxYqw0YHU8vRQZiodBTM5PIFX8Td/ZkfcouPP2Ns
Y+C2YWu+gL/VMUVG6LBcGAIEhhJ2j1OHyFrRAz1TeqZJtEFwXqzy1IU4RlraIzUQF7pQRSftBvwY
dZeY3GZF1NB1CRL9gODyi08PHuhBSsfdHc2dsSnV2pSCb0RQXBy67P6SFcs5/WYyY0TRjmkza0u2
22z7qpGcSdtGiacQbRqp1n4r46RNv5xpBOYuRUHzSehm49BZ00YWsxSm5YiLlzGC/9c7T+izETTv
eVt59HeEw/e71txmdTSviZbdm5J6JPdwO/uDhBq9xmxvXElhOXKqZ/Zn+3LtWQy1S977NyxJL9pI
hjsZ3dS/K0wkbCsfafHvWDod2kMtmFlPZa7x//H8n3EskadXoM4ay9f7tjVtaC0PGwJybDQ56jYb
wAdDlcFA+OIDUdG+35akrs0Ehx09Ouma2GBiLfoJWJ3iJPJo9R2iIOuwGC+NQXHrKOPU7/zZLuXY
xN6ssq8HXQy/uRvwagNHDFbejz+NyyfCb28YkX+oWnmOwFCVKZb2QIOpM1l1Jn8/NiI/0VMXOLuV
iK8NT5gdSC6krMjpLf0ourd3eFLVdkyCZ6TfgSAJHvMvJiCPXkODeyowEFxyk9I7SNzDC+5DqJ9g
JGx4ppy1zG0X2/RbmygQG7gqMdEBMd/YsMX72whYUqk92+QXHqaJpspNtvgueO/Id3CoUVKgE81I
7hhlpPUetoecdxghDpJfWeShsy9YtoBNND5lJQYiqLLBA8Nic1tBkBFaYoHXqgpbZLbqnNhiAVms
38mImOnG07CYPcpSH382zCq3dKdGIxUx7rXTuozjZ8yl6SjapzXxOe6yEPuzb7ZHI6GpiMSa2EPR
GPQ1A9uBJdfEvBrbENvPiNNE44qfxBuIOgusQ4wEvgusblkUcoCo6t5GVaJG5v7VmqRIfy5IwI8c
Y6Q5macXcLZ47mHyWjB0EDRAiSWdJ0w7u91VV/o9zjhLboh2OweklbuPg4oJx0n7EYoR/18M0YMh
ocKv5JV30Ydk8Bgf++HpXGyIsWars1AI24OJDWUySWGC62dauhHtKXXLFyZ+/CLoVJbuLc36BGBr
qtzwmAu4lU43kQRZAEBb4IOi0GxP5Kd6zCPOSRSXSSINTNC/7CRUa97qjxeoCb2IGqwInetcsyf6
IRHVNGAs5RYPN/jRccXVd5fqH5UHkFjhsR4IVlFtuHffbN3H//JuEauPhX1yZH7mFrBtlt65gi5n
/Wm+jVpSOqya0bw3jtvrQDz5StcnbK8jF5s92yE557weovohCYmIif/2/BR72MwNhTAd6QTGdrat
CyMhu3yZwCRCte8W7MVMxd9UmVKb0NdXRQoIyAkB/ZrYvYJ65hNhw7A5ZOxrNKsZobAgxmEpDIhC
iz/7QXMLmkOXVQGDMawX9sZTe1LosiUb5NcA6FTIaKxmOi2SIqQcuMSrgIBfNsAoyQVgIB7HgP5j
Ju/FTZ2MY50M2hnAnP15AxrNx+Yb/6yVMiquBdLX3K+PzI7oM7BMEp6c1JA5JVrzoedl/XaYmxKm
jeGY/XGZcARqGU8Agi/ZjF9/vciNggq4Bd7vp2/ZqhS8GOZiIikD++diKS0ELt4GU/N06MJsPdFG
XvDq8NQExtTYePKJDsl7Hykqf28AKkyWrOiaRD0DZMvz//vxzrkAyBWGZlXWtXLD8NDKV20szg6L
zNcp/IkYqA8mRWSL/hl9MnH3rFtBWPX1gMLQ7aXiHipKcCI1xYRNQDr6DqZGYLgo6Ul5qCAjTsFu
ILBCejW1KJbgOsFRU6Oc7x+oWJ9otXOsIMPl5cuKdQ5eNbRotllgUxQhxfdaKwCJVfe7AwpVnax/
9h3fM7KEEfu5D/XuOTCfBmEM/IvinCbc8YX3PB4box3HL0w32wsOqDRl6mgqUlepNsYYG94bCf4N
wIU+TxD0B8R7ldWF9KIoOUvU1ttCQJvki6WyvSCjTxfMQe+iWLzMuBc0sY0AXDY4SKHW1QW8bL53
bvpfkOzb3v2pTdPKVPWK+g0Lfm95ts3UtgVW4+/62h/c3yze66fWJX6WPDLi5DTFEeFLUPA/LUS/
49QVCLxvPiRTpIooTHm59aNOfgfiOQjsgu10vGFgGNGVLXYE+mhnqP3havw9lRrz/s5vdBFGjIHp
kSi3yGSuSqxlHVH0IalARsDmx09+QizGPry6ss+GMUif2l1XNlKvIDNjvCVHr7AFowGKimi4Iu+F
Sfv5kRgq8QGFFbVj8HiCEuRbGfsDEbmnIKlhvA4tRlkcQ3FO04O5sbxdFSfV6TOQAAoXshLLDyzU
ZHaik+Hi/nRfcZKZ5USTH23efF/ygSyHxXF79jPzpUg5rxMEMWlKJc03wIWXFFkpBMhXhNEKuthJ
D7F30FnOavrt3DtZZ5grO2kB8WYDPKfw75vriNeijs3PJ5mntigknSvnr41L1krMLfTek9Me0Olx
rTs5U2OU/ppwmgVaYieiQMD0V9lK/C5q478diluLqX/zkU5ChMZ+9qINqs1Mzz0dNfw8zfW2Dxqh
Mgy3s9ZfBIe+mdCqrdywvvI8SO81qOcqeiAhX7UIw1dPFRZUfDkRuWD1D1vxkHrBW7ATDsDiBIX9
PPHVJUAs0uYE5MwyolVWJi6D1SGY6O+488tJ+VDgmoAjjcLnXbyu1JSiP7hib1EkL8qH5wqgAeND
YwDY8yh8S65ymom/m4COPm87IT9NCo33x07CF9jAvp0/1GHKO0KUWKpwFrwePMDqYLnADeg6dd77
5c9siajwsCPu/dzb+oixBn7tGqQh0hKkSviRt0zX2O7gC0wkgtXFvzhFFmzDek9Z154OHQRBjuae
DgjCqewC6UzcJQZ1bJUgb/+vjJeBQ0k387OUWUD9yT1G6M+7purbB5AkL1bP+CvcC/7Qi29KBv6G
4bHx6z65nBLz8lYp2YrUc/Kxjm44dObAEo0gRO7SfzoqRgJGOB8MAAcrcUb1pnSqC6ZGERl02nad
V84cDl+wyOoIgeAKPkBuiG84nJTGOnpI7QiXb3NfCuDRD0jEFR/Jr1BqBSv5M0fi/i4wyliDtb0H
M+Hgy444lsB9RrqXrYdG0Vy4qyjKlc4rcVcMwWNs8MNkvavSHZwidt8rordtNJMUa26Shy/1X+RN
E3Ch6inJ3rnsDVQZ/32MsCnh9CIO1inJTMPT6TE+rvpylF31XypFpqk4vrM7wBR3glbZu4UvydQO
aXUf2iPpj52flDMkiTlIQdWfUII6b+hmXxuARfS007+ALJTAf8584sK7KSo3+jMNWyChQvyT2ufs
lW0jFJDuHwYSz6JICxcRomFgDNHzGYLa+wF2BaVX+R5K2eD0674vZUYyvhhX9cEccM+QP2yhPtDF
BUdISnZYTqt6Kbn8uW+0qzDJw3wAju0wg0zz2svxV0qxT2b9nG8VqKIof2ZNW/4yk2tbgSpyyzr/
soJMmMKnNYOLSfL2t34mI/6kWWVpIoQQ6nMKwtbjllBkSW1XzcTIlThujYgcgf4Qe4sXqlh2Ah4+
cHW4johAvXhHyvu+RUeH2XnxDlnK2vW7VRCrtvGGZKOzTmNaq5V4E4cTddyh0JzY7Ux8cEJ6uZs8
rGgkIb8XQCzAjc5tdNDobPBV0QmB2IJ/wueuaAdni3zX7023GPutKap7IXsZVuHHOFHjVoa4CAXo
iQVVyQWHqa3l1bs1PHBikc1+8VjvUODSREQcFKh8qE+3BN8MMC5DRAa4na0bPBb9qWDngJ0a5FGx
8mcZxmZrK+sdwgmwRoTpSu6y2zx+ssgXmLo2UQMMH2hotMLB6CXrzKSGgmS3TIXfLLUKnpaCMcql
xJSgWkfUTf3+FyCFFUlCf46LJV4vmFvoZxyRwMfneTRoQiJ3XYGqtLBEWDHgAu2+sJqqMDi4H5hG
iD6mScnDpxJuTi+FzbN1FH5oidKhf+L8R0zC6jFMJCDvXMJpdUaRBW8gCRJhPC3lGqz9WgvdfCdo
vb4G7A4NUBGt1O5f3dtZbrcJ3ik7udSUrld6kONZaQV+VHPoZMQamarQIMmwDByc3a/7JVdPhFyh
HJ+xXfyVrOfglvIGf1CLaRN9gWKOvUDJqyWBvjDPweSSa3/csd3fobkWATXqHzeTaxa4n3FGlrGC
2txOnHGoqH7TfKHsK5WNQQ1X8Nvi2+/HSWmOqOXLT5Kqsp1VEUELoPdkyIfsIrgYRde30NEeepDb
CILwkppTnNmm3X2C4NobIx4LIkno/+pKkI5/8oQog2RkiJZIdnFUBo9yAs5dk4DTwfgsfNaxRKhr
DZ7CIVE9q46MKGqYpUHIlugkVs8VmbL0RLr4zN7xx6wNc42KTuneEwlhF10d095Vd8eLqSJOf27V
eDjtPudJ0r/qU4DPRn9LNekcHcP3xPYqUqK6s3XVO1s100vxrXwNKzsC1NgWd2jfZNX4h/OIHE9c
Tp6TQ8M2y0PM0m40lSktUT2YSt+SWgT1n5QIjL8IT6NBMe+4kQF+cG/jYGsz8PKjMO9efjAkR/Fc
qIdQ+m1xIluCWrhFPXQY2g+gOpBCS8XSVbZtk83Zdm2FskCTYon672Fkadw2nNNKWbdbuqXz2JMp
PfVnUKG5kGavdkc5SHq8eNCkNhP04dcLJHvLp5ng+2IS4VrjGsBADeOaMW3+8hMN4a4u55c2KESA
19aIDBr0S6weipoYLSxKwGUqFbDr/JzNH73GzCyM1RdHFVFoyjmqFwIzozhBX6PyzZs5SG1SPkSg
4Mop26cCgPKvqU+QVGUXeaycBGvnAjqGSve1NeZv6UxcXqNeUWISWyGu3TJ0qVPlZS4f3O4jVXDn
XJPuLTb5dJnD/VNIbDP4KRE7ojl7v+B/w7O966ju6WB73dkEqaoyT0NrI3AjlTYqElGnQvq2cj2M
ON4QDakfb4yO7/poleh1sbnAJ7PZUlW966cLQuCjXmF9xNmJ7XAhckfd4Ncp1blppB/90TVAGWaZ
+3XDQxefHneryS21GP5Z4htNXgPbX9kgLCLUPS+0GSpmx6CzKwSirlDQFrnWtvgY8KpkwOzmjHvX
MyhX51FXBwX4tTO2f+nqG9N9nWgtOwWtMo/d/nvX5yD4NbImHI1D5hQDsqcGNOf86Kygi02Zcp2D
mUiszAmaaUPi2MJcY/btmb/efnwzaiApqOSfPuAjtJi/BOzapbUwdl5zoMD+e1JDch2afCccbs8l
xzwyjQ39uXIhAGyuN/n6avDZhi2lEwZWe/JCh1FFl3F5/zgCYLmJ4pdE2B8XocrlU8p8AruMarT2
0meYDqOI+r8PHGh/tXZbTrhMR4B144khPALiNN2JCFgBtdyJc+yusO56GhS+fUKOC5gYsysfDK9y
IWjA5efDTvs5NyEnMgE6UmefVMRUNwNGAc0rmMZ1s1lkJlL7wKe3Sh2bLINy96appvyWJ6nGCWVa
WJcZdRTkNigPW7SbNHNbnoi1uL52gzoSFeMAprAhfQQ1T1Y7j98urpScxz67WuRF8sgXQkDQ6HSx
WlrF0IoIjm1cRwBk2+BcaeEOtefYMhn3G6wvbGWcbbsSlIC/bVdYX3U6ucUiFOtdFcmLQkotXLKp
XRqxwsVwJ69ERPPBiAabYZqJGjd+9oJoAoWS+yyCex6EWO5TuaOou41ZTQXQjwpO15izckvUDjzk
jNSQIyPkl9+Byy2LhmloDDjceK4HeIdvoJTU5D1bs+CYh4qNqT+jZZri9qhYiJXJQOJVqW+Rym3T
nbl0CJZHo5FabpIdfVg401KHnWl74rvGlgBqXuM7TgA2o5TliCVUpFuAQGBsrZCxJ8BsisarrwmO
/Wjwi/kZ9QEBFqlTBAVBggvNei284ugRSmJMUJofSP+r6/aqUpxPJxe7wGQEIVo9AK7xcWZjB0zc
51n24ZFJhAF//u99I+jWlSl8iAYxTrCqlcR+UHOUYQMsiSbSuoUQBmBsKuElbZ3fXvgdJaCvsiP/
AvG+vkVWuDmFLjS6KGO1DQD4GqO9Hs/XSu+vcB/esXcz+M5F93s26j+Wa+9s6+n1v9zMnFW4EZGy
z/iq86M9SVn2fwnv78AvQxkXOVmTL6z/PLIQjqCe5Xz5l9la9bnbu03b3BzUZmeUXydopmpY5lPk
KWEw5EnRCerPfc+WUEoJEpsOl+V+cpIKnufy2HoWp3LXm9eTwz3sX3aegpY3ISKsJai2pQBVebRs
mB3FefPKq17nZgw3IzUvRtZgO1GD5TOsYkz561dU/MRD6t3+aVAPbuI1i2j8Ix8SUsbpziGL5Qfv
B3ieEUsvfTzCuAMoIDOQWveNFDjSXhSD0Q66CFo4Y9xtIe2hE9GjYPLUvAkrRl6S7Ai/H0ILiOXc
o2hTZHco+Jr4/6G6GULV1Wi3Z1dZvo2TC+Ez3PeF4opFP0CtM4r+chxTsiPQmcnuuHYsV4d/qdgO
rkGUk7QkedNzOvUMz1pVQRddGwxpjckjMxMTXHg4rdFTcx/oKaCViuDa0rBcyn5Zl129YDHPrQ96
pWz81FhUNabd5d/sZhKqefAAkJE0VMIZsbH3+A4cVZtEd6NIigjcO9pppAiKhqy+2RJ0WqYPwiHT
vFBhr92SV1RKtHDCDy2C+/VUKF2zwnTkj2wbsgsEG5e69gRgRJFtwBc0ITwP5SXUNjcsYdYNGIwU
eFHsm9bwX/YOaO43lyNZ3u8hTd0knLc0zBDMV/p77s7421h6lBfriFs4xadM42YH3yS4FOR+Hl05
oUPBnsohiwessAZG9Hp23u2Mi1hFhP3bXwRRwfs8hOvbm8jmIBAKBOXcwXl21ejz/iyb4LqGDzRb
XOBoXc5DcAeU02X60hUSH50xzIAa5c9LfPHzUVbFjcjMtPZceXtrLUaIZZWV/NbfUUurHE9rY/KC
JCvPrDNazQcq+RyWbX2FZcA7T1GUKhBcoPCLUmLuQjC7fyB8ycmCknSFp7hSVm6DgAUcrHiiip3O
RA7Wd/eunNs2WC1WOLvibL7IxC6vXtUNeaAgopGpP4en/CP1J4WGsO0EbEdTKxar3oVIvsD7jOkH
FKq/4P6pulLR+oKOno35YGtkSdYtxEw3Dg4lBX37JjZ5/x/0QXK9r+v8iQ4/qVm1nvaOMafwMge+
FyJ0ZWiYwPVrbCzETgjDCRP05JmhtTVqFw2PRw+SBmgsIYSDvhogLk2swcKk+2OBEt03nja8zfCa
JbDPz44Dr1z+byn1EfuG8w6Hcsa//yPSg57Q9qqpArx7SXlTnpyYao3BB9GvYG+vMgwR4kXVsLpg
OWwvVSaBFJ6NBCO2U1UzxE4NQHSs5/i+vgXKLFiwlxMfy8vwRnQQbZmuBaUdOGuRSj+XtHPHm3IL
hPz8sU5kEPuWsLGAIn82pPLUSeaVlFupgryxPI/dx6XedblR5zEV5TBbcrA/Msz3/p/BIoCh3FQX
fXxF+Qa3wRLgFC/fDfsnFSUerBlhx5Ru/AfrfT7JVW5nro0Hwv6RGxhbUMwMaBwyWYeC1B14Qqcm
ro1TONQohez2yDwFajuGjbmv9IdC4ycb0NYSjaPOu1hwEY+J1EVU6myNvYDLpnx/1DzqwadIf7HG
YjZH8ynWK5D0vjAWarCdO/yxvBRR5Ka3sQLbCWf9Jl62QFfEPyoLtyLDiaSRO0EULMLEpRvGPT5o
Dz9jPd3/i66G9F4ht/jnFU0cpegTjKW/kjQvtdc0o8y+8Hhx5ONDLnKarHkh7LnK+HvOFbgrG7kU
GDs9uuN6ZK+iLHBD9q2qATIU9rnB7kz9gaycyo+b9CVR/K+Y7uy3E1PEmQeaXO4noKrkvDhs53n9
BSNpKugzf0JL/1uEChp0kDGZIeG/pcF1ywmcZ2paaF9rgvmy1d6awksD+c2kaKU0R1XBPPydmmmh
oBbUSlqHqMPpJs70dUYUG1fP1cgUuQwHn0Qfef1ntBqkkMlAQLqUB9Mg4QLhJ04bi5jNjzrici60
9kFtIf4n3/dxfxekpd+q8PLMjRN6XcJEqbyLWTxktQUxvm1uXT/a4isHIMDyGawgcTnHYwg05JZI
hlmyiaNDXqPQZEQAkFTBKD9060O4iUChuAvv7M9893+xwTqqHQXEx5HTwLxR8zhtEEIAa58zKkRf
xmrlXmLNpu1EWucuWMFJN4bCdQg0ujp3nQIi+b/fQZKMTJoHRaboyeB0D84YO5teGOa1y0PiMadv
ESiSSNiPg74uwIjryquXXWlAh8mGwxLB1WqdNmw46ZLvnUEd7ytmhGTIb97ZLFNUE9wDZiwB/7kR
vOir7PuSXR7Sq/bzT/sDV4DVxexv9EJhS1Ri8FFYNjKIitLrDkqYOAs4YqQqI4o/nP+3sg0CcDtu
HUph4w/aiI74TRCN9rJwom7B7ysjz0LbGgzx+OzEhu4nfOtpkjLSAbtiTYzTIrA1NCK7aRu+/Usc
6JPJoYEhP8tffRtkFa3Bw33NUq5khBt3UdCKKT6ioE5yaVsvunsVXpeSiknqPLm9j7m5VxZmUTvp
Wlv9S7S2FlpTxIacL19nn7tTN80E/jtAcs1itJ2zH2CNMPyglZQ2TEpn+sHAlN2qo8DiQsFu+djh
PzNgMvpiDCVJ/W6LL3BjgkcJqjiUmJn8x9+UWmYuW2ZvhTLnYQfOzekeHspMmJKpa6+dcv96p7Xh
6kYyog4FPycsCO94+cw66XO9UyY1Za1Ikb+UGiyMPvCQ6MyOxiwXKEX3qZ7W2Rx2nRBJHuMe779Q
HqigQA8iZt8be3otPe2QtjOgnvrSGEVSimZTMZb3q66TofpBGKyaEDzXzVm11dQOF4SEEYZWdK1b
6uIpRNlH1qpwg0hgGwybCUk7tdQ1Tce+12mGPAJ+EHUSoW2kiHT9EdfV1aIYoinYzULmokiBpks8
Eka3HWtJpkp2CdVVziBqb1GIPwOEuQEF59W64PG/i5mLFFHE6cFcKWAR1+8Th7hN6Q1wD3oqh8D5
2Ar0bsmeAge1B03ZBGE9Vr5WMAyqos5ypwe93FOUKbufFsVfKAT4o2QvPbSVoyWjrZOBP13t4ctB
JbH30DSPsQnAjMHb2YEWyCYQUgygweMbVvKeGYQEmUm/fD35XRe6tFhoHtrMuXoiZnhE09W40v8v
+B9qms2cj7TdYLo8fpXvGTGR0QieGdRa41teF5jZB8pWx3q9ckVgkAEc0cZ56Ut7TGSiu/sO3cDT
UTW5NowGvcdxKL98rR2nzquh3ux1QzXNTXfOPVuw/gkl5toLU2r+agP7F0K4Z1hbqAGWMvbj2zRn
Qug9fsuXcT8OPjKEFMECxQKJiJKpMaMfo3ljnl1MFME6URENu4qXDPau2KSOX9R9PYO/UoWSnoP+
Gty4OVX4nSzDCTKgo7GwZSpwqPhhKMMDE6Ved4wZed60sT0hzmleleAbmz98RBkBzDRMx2I6MkjZ
MPWskmc0dWmKnSOpt7tA3D2tGE6YjcvyYNkDDqQcox/GSWxP6DleMrnW7Oq2gTyyB/m222TObybs
bqcjXEjjx1PjRvb/fnqx1SWc9gd3859rOIRuPbEgCzB2ZTMmFtOCkvy61Nw0YHFH+e0H0eQmsdDK
Rz8Ch+C2d4c2ZLzPDdF4XmSU8zRR0kL1isxT39FmOxtspq8/bBE1vhxXMWv9VfR7Zta75/p52nDd
qi6saLeeyYOuO7pMkk6ufnRdpP6yTrPy40pMQ2pQ79g3c9CJd2xzyMvsBGhKQtRMTvRjhYinryle
867I88wBwZ/1RJKdlx1ZSSayD2UovN1cv0E1Q8l5Yjy/6WKWE16eriG8ubLAeCdm73ik0a9+qcYK
wPMXmEf2xMuXEiYeXoWBHKYZFmHH+pDQLmosGMQxrVhIx4FjR0BccEAmUQjZ4sQOI8Utn2hmfOab
ZLokiPlB1nNalH5PvrrLH9QnXm69+vjLm04C576ROtCZltgxFW8C1hafba3kRTnpENqi/Mj6eyQW
X89/yU+vfOJ04FhDCyFtmISMoxMsZLUlnKWYfalTUU/Ja0tMsfEiQh+XifMgMhErHXyjW8n1Nz1T
+g3Pnml8yKObhAOPm8Utz87JD2Ry7WAFT9lbOJ1jCeWxYeB6y0E8uIUY31H+s1mF9plL5cMP/dyx
N3Qu1C2S3zoFgQDPJiQEhpaiOkpFm3klO/upzMsxCgxeI1G2FVki3H+OSrY3msclmSpW9U7LJE7r
I3/AoIoZDtsXVF4lwHgS7zFMX7eEK1rn6gcpzz1FY4oHXNSWWf0aM3jtsvz+uqupZwIG2j8Tf2O+
cwhf5TPu22t0xtg7w94nMk0kbUNwnf+3/IL+Qyj3ClHXRsmTo4ys1j+DOoulQT0rI6cvm61gZEZE
1J2pAJxFNInbUzcNyVXHcEO2vVwcj7GmGXBTd1Ju1Fdfrv7tRVU6xcd0s9FgcrZrC7HNnj8nWPES
XOlttyoKbF1FJCHsquONtp36WZkAszrXwwhqBlzfQ6liOdzzWiVk3itAaAVG7NanhkW4EEmR7KBi
L8j/mpG6wyWNGz6qNbQ1bYKTmdQGV3uQBiBenVhvhWC/v2n0h02Mb6LXYihjGhtKc7bVKrKHAvPH
QK9QUqh/ZE7/XHeRMtnYJCQFAqmuNXPHXK+m5lgmbi2X0jmFYZQUpMUkxJcSAAr9EGumpfEXZyMl
E06pI5miSAASA8v9xbpmszBf3Nd1iBCoIpvOz1mW5FIUyL3a5jLfG5Yl5kwkeT8IUTtBnRMI3D/h
SXjUCFQGXOzQcw3oW5/tfx9yiMmhekCVnfdwEs/JKgpFaPWCsFytAQayxcDqn3cl5RD1dqCwwJwt
eu1Yki7H7TljnW6MO/E9xTs4EVobvtjZ+4scNF//+9QpEJfzik50pCd9UTRhIy7jSmNU1bJVFTHI
tY61FyKPZnka+0GU8qVs7FQFHeBk7E+ZqyKSDxdz9B18yPZ7hqERUF9zXwoWvTUQNjXbTRDpwK0k
uoEdAS/b6odgqlW2kBw7LVU47wIOqir6A6OlRij6N+aDGYp/TyqpCnDZKXztLNQWv0ZuwPn1rcZj
ekT5kWuXCr0JkpWvogQ3c+Juqx3Vgy4u0L3/oBOFy/q9tIfIrBAPRkoWv2pFLiYTlu9wAsmqpzZc
MWlJJyT5eTif5WEi6+4FYFTU5xAZrtQ8ahGv67QC0mREWlWpCuiHc44PPvr04BFx7n66AEKY/J4o
F2mMpHqTY78gIa98kfTLKjuwLu31g9vnGZVjh8N30ZPjU4NasTo6HGOLd01uSXl5YB6Jd4kNqWoP
RN38icDEhMmlE3tKf7qzSUaDxbSLANnuKJ9cjNA3/oADrgvyfLgDh+hR2M8mwIudFXIrSQBsJJit
6FsTy/OadkkUQyciUzPsr8+Q4sP/TY6CcKOgiMDbYHiNFRzZmucjvxhb6N3ZuXtPMnpiBea3Baus
/GCT161oU152wx9vrxgov9OsPD0CtABQUUhtONuSq6KNeZQiRRWWQZRAfstigR5Q2ldE6nYXaF7v
4f7OQcnaJfWS8qRCkz5quBC1lW4xR9HkIZN5drw5JeAOdWkDoUPqUJqygbMMQtKD8Z57+hckr24a
HkBv4VAczqFPw1LS9uZMuUaqvhZaKn+DbDfsX3kBfdgQmV0taNl0FIdd9ayOQZS0PuF7KcD1luYh
j4o0n2JUczRLwMqAwBjrxS9OjV9oHCui98YjJfkO5Ii/1iqrflfzc+HIVkrniZSkHhAhiNI+q/5s
honBdmJnztNw5igdWws7GyoxVyVsumH8b52R0gKWa5Xn3uyMmP/XCX70eLhBhSwAcEBeUDhaigQ8
L6Ti7paB2uu+S36uw735XMO/OODmcASSBq0G+8TcmoUdBxnRPsGmr4hM15nKf7EkzE6amH/cVql9
jqrTuQ2syevVdqr2SdIJlXFbihu8fcXMjxhURhecHIf4CD+ICR4UjmF642shsLsVO/PTOBjOFnYx
/21JZIbYSDCxdNT9oDtoK5K5XSH0aHSvNTD0qaMpE4WEZAjaGfHvWMHxK/l4I4Ir3sEKfTUo4No/
lllDpXjVIOmGIJwcvS4u7GMFtP+Rev7mJRpEU07C/1QINlEraj9b8gzcwTDCTdvWAzDZhtGMDPIW
HJgx8ZzOoicfxU0qf/sdLYTfNVE8mKyiFCzU6bFVgu2KBhCuIIqRwPWQ43PK0qES7pfXXtte3p13
DdoLXQth1NzwJAZR1f0H4mhPF3Q5MRMU9zqSdrrfzyawd+LSfkNQqW4QcqlbCOfxOT7pCK0WN1KN
IY6isW4vWa4Lnnqsrp9oBSoNR2ynVeta6KpzsPItAwM/JOGP14NPR56EIS1X0bZVyNR5gtFwqEAb
XF5wrTKObe1aUBx/0mk2R8EfzY4HOrKhBleZ/oHn3aprX33JGTW0KnXCnK+wz87px/hFADEEzfl1
FDXblEzKg26r8cb+ApNi3qbQDtrxmjtCsTbhsI+EbTSnOvfwXF9gF80/ALWNg1IJ+E9JLj3R6k72
XmaM8SbDnGtf3jgnkFkxMLzChP0dvHuW6hrPTk5xP75UiBRF5JbwY2GTOvH+fhjJV85XEvc3Y8Ui
Isyzf3Ny+dgYscP8so/fSG844nGJmEpnfpM58oLiIsZ44MBGuL9v0Hwsz0bzQKI0hyokRFeucPQo
IHU07UwU/w2EsgBZEjB10xkOp/AlUbgD/p81pTyjL/PSBZPMVudZRgRDt3bUtS4oAKEAzK4w5hHD
/cK4P8w9CaYq2ib9WzwNkmh3l+X6YTeubZUbjO6i4JfgROIcOM8aulRFkbKmXFeiSMhzzqrs6Go7
1B3GFjWmJ9dvBrEj5cdV0Bx7zbgO43QWsy7QPuj89MQo3XaEG/IB+V14VpMUvvrNYga04W2RF+GC
xLkRmLNXSIlYC6gcOVDD/TxXwqK2I0N+eUm4hr4a6QTEB0vlGIHxs07qPp/asEn92t0e1azIoOjn
7lM2uWnY8B57zXn9EgGrslZP/xxxaUyR59wWpuDZeUqM4edHt+QqpXy3EzGeE01RxwZAu4EAFVAU
xtMHDOWgTfU8yHE/xsmyuPlpXI6Mwp2MVzzApDuYUEYr+gghKGfIuE2x9ULvvrkpkINCKbrAMguo
9F0PdkvGx7g28LmTAX5IpBr8VlMPGNQ7v92rCrLQbFn6FRxk+HGHNTQ8zTiLYFBCGrCK8omC+yJS
xOGQKopZ4QQicdVA22uOlvDeSIHBHHapclMajJ6Wd5NJmRZG/GwU8nRifgKfRNKly5cEgzfGDy4X
vJSaAKY+OA5K3GueWMUIm0klenhCrsLfRr635vKvwF0mdXQgLyM/cvHiPGF0MsY0OY0HK7huqciz
5bl1YfAuPlHBbxgpjc5OxpYKDXsPsKLq3q1LOOKMHMs7zW4q/BeJtdjVu1zuXg/Zs/87oHqodIm8
QsrsML1ZkhwT8CFRtnkmmre2sqhbFezcCPl0YmfJCh4qItAFzdn3vgqzo4oZ0ZzAEfEy2iUnmsis
LFb1SLdTKRlc/FrXbSYRN9jH6fWszVXOOz6KDKanREgdEIv6jyCP7CZNeHla1vpp1xQld0rx4aK6
MyEnB2NyHh/7F3bQS/MIqKROIK66bZFPnEhtlgzKftuWVYLaTraeY0Ia4IY9tWTgYVi1SyG3V++b
XV9iz3678el59Gan43wKnTATRZhFnkqrnq09NV39xyDx5zZndoBTFWQg2SXOCBp+KGeEhSh0xKx5
zaT+WBVhTtFX7p8Sp4577ub298zowXLlU+kHHSXCqjfAnVuszwyLizdiURn/EeM8owMHo9vUKG30
el4bSNWhMUza7+I6rxFJ9F2SAkWSCBaCUooHvFb6031VdQUebQSuxy0adQWvnoD1HLTzjO+JmwNk
Nnz9agrOQofNztj8dWXU0fSJeTbV+dGWFTMeclUiLnqXgIIgOs60VMi/zf3y5105UMlguznM3U7z
Vs2BfOFlOj9h+ETw0GTFlYdQ4Wp4i1O3EVPQjL5iSjMhQpOFXUEdnXh4rWlE+mtgRs5BNW/Z/LHV
2kQdo9Cd95keXXuPQeXnXePs4FLXQH8zqxELtal+lFSa4X2Tf3cY6PxgKtEgbe1LTb6OrgZYgfq4
6cs5N5PKyCMmaX8fiNHHHFBZXZblgRm6ggcfBwSWlNaO4sQ6Lf4SCaQ8j99roOs24vzZmIfuQFie
b82Fl9/55PUwKM0YFoPm1v+ocj0quIwiRJRvOzBn7ajRNm15+2Ab7Pw4KOsYd/i3lvwpnIOEe/pv
cji5hUBwkXdKLf2l6sS1JLRvf6SlLC6/RT/d0ffYo0D9xOa5n41eoTw0vx31NegEOJ0nMz4uROnM
lz51amCrRKwbcDxG9I3znPB440zuO6+Or8Sa7BAf1TSx2/gH9n3Q6CNGbNyyPXXRn7WGytfqLxPY
sN6yrduc13Kikjvo1oZNJt45bpjKLoJy7ywZ01dj3+UZbagcE9TLqI1G/HYIktIb3wj6ZVARI34w
SP8o3Tj0VQHZDAu6UQoqnFscjz47ArAAhCYr+5ThaeFTsWks9Ez1zvq9nFAVfJpdPjsLtgjcTETX
hxJl9EfvHrtnQFf7f4NN5GVBpLEf9h2brj+yaO/aIMVek/jI7yV69jHnQZSCf4KQFJ5P/nauiqaH
YEofG5jtHvLZoRaWC3M+8ClWaIgtYeQKaOGnhT8/0Kuvbois3tzFbjQL7XpxtfpoHQejBp2J7JVl
G3OOILziydYd2I/ciROQZy3Hk/Bzj3psNPliBVyvVQN6RVQlZ7QZuKbJ3eFU+b7TFbwtbCM1yhT5
O0plLLW/uAk6BOq9mPLUlrrrT72/PlukJ22EfVVlmCbj9cVQtELkYd6tASV/Ch9C3O4iwM8oFKqJ
QpIsnItXb8jm9BZMJWmE4QrF5PweNmNsDkJBNpN+0D7nZWB2m3OeKfG5Co9DmSWzim31ILpfnodS
7t3Q5qB6cu+yNEgdZS8x4olXdAEhqvvZ6OTCtxcAiNsNwf6DcvlI5W849rdI8Q4+LasJnQ5PhNdB
PCW1vXOOlNVM3e+mbuE2XwFOZe8jmK6KuDWdPkGDSXMrm0sfsiEHFDYml84u0eJtA9c7Q6yC5GB3
AJnVL84C2GKLHJeTM0KJQyUVjdrMbBvW5XVoDWuiydnzXSy3nE6tWFGRIcuK47SDhYQZAdcdmkDS
tnNjiLCJAAesizcJLWLDLfWN6SaYRzfer1dTnExP68eDc0wOZ0DCvszBTm4048NEeIr1mIdLN8TQ
2n/iIDG4ApOBg0ZLUo7MLnUJjMPjLIAXMHlqd8ktTQ8RV9JyeFmIwT+ajG6sptZEumpuzJWiHSsH
Mx8ylojq7z6dX4iinr3gnQ7KwVhSgsZpAqAYeS1SYFr3FARxnaaAfXxzFE008p48VBvF6ZudbFLJ
oVHGWl9wWdZjtpclel2OIH25UiWPcl1327ZqEBL343ID7OroHh4f1Khxpd3/iI0vP5gtpYnH+uQR
3BPRYYVq7P45nV55Fty1Su3bnn04BeujgR9bMyiIk5LGdpDUetIxCRA2nTPY9b8wxlro3xEJI+8R
5wfBVrFsMTauwUkDHgAykKskOhPoviDjGcKm+PvXjXowwOpQXyeZhX/dEqdECboo1E1txrJr0jDW
CoVo82S8OvHcOVM6f7vroBBL6UqFK/GBbhAhFG5nwJ9EKlayJX74Ar19jCgy+iD2qERQW2Cd3ATv
Jyk5ZkEGtpJvstpZlOgkF16PZ1TBDt+Zk+9baHLTaP844yxFYtz6jJTjhh5CwIUZCdk3c25g2p+B
kOfWbU2xhSgFG2VOGruAWLBzwY+FUO5bexEuJqzgVtCy0XXmx1zdm6Fd+CkWZazrjtPHGnq5lOZv
8Gd9UOwUtsTHuKHVvZ6fLuXuJ1W23YBAL2bn9JPh3BSL+N6xPTNbKr2T31frjHvRdpGEfA506Hnu
i+N3WSotF6O+KtAqWDhqccVXoENHw6c9FLh3B1ZrT8CPgcyEIvA/nNtnlJ6FYAcWtIOOVD3Fo3dx
6cn5IoKkiomSV3Tx0px/KFVAXm8X6O48Xo7CmzvZMhUhnc3LQhbjAkHIWra+JOQKdBONC1Za1Jzj
xbZw7XlhYREsQz6JwT974inXWF3q5GGQc/Jr/9BTW1+jEG1w8O8MWg+r8AUESevx2iENVfFEyKa0
2jumwjq6tYRlzJv6ovkIm05cUzVLvtFRvVK50iWRMhrcVTBgVQIqd+W7t5u2OXw1M601RROlh+lh
yYMqhb/5ZHbLJ3LfdG56djmSg1+pOosj+u7kT2tEe/eAYsU/Wkg4Cs0knODlkjlE8BEVbiM+SwMc
TIMgTiBD1ECwLQMnUJ8cV+OtkoYJRpV16/4O9seR2Txxp4/cxJgaOdl0pv77AffMVJ2lmFHZ9knt
3UxRxXMuXL5zIfzio0gaJqDfFtfckFYxsyc65/Az/dsav7XNlWlucUBckPYptgJJ9S1UNjq3jlt8
UlbrvY0p5hhYRc6E5conwq5oXJZkmf2SH/FnlyHFDqpvBDdzvaZsXaOaCYn1ubBIX9Ogy3IIwpa/
hrJRRPSKGYg1uU+Txa7UuL2m+cAtDQV+0Bnu1kVdnVM42Q6uk2GbuR6TiE+J8pbq06XGU4EJpsyq
0FG6UcT2UANB/zij0CPEosn9BzDf79VQbxKpGHW6ZLJTJ7gNVz4gJouy54SU4ydFVmmO275YCTUt
nUTf7qCnKR0Q2yMHDRL/LRmiBoh5IiSFu+hRGwj5NoEk3NGVwrlXuW1EdJYuEYbEJKvk1oOhFcYz
inyvn+Q/vNWDlyzegA5bI4PgW18c/LBaBYRF4rj2/p2MmHMf0Ef02nrjm2i9H159wjSYOFpZVYL2
qthaXxX4YGKu9KKk6PhBm9qkAgoEyICQnHc+DD0sPD/6B62SSItI12X44CtjqsRSPijrC3DjaP8Y
2q7n+hMYt26tU4l5V8jr8qjBzeQOs+HI2RMYUZ4z96Kq4koLtui3edjq5xBhmw2SULY9ytoBv9Yg
M6MtcnWvESpmHZ1+CBTx0vzADiJpUC5ydZChmW22kWH3cn2OlkZmYu73aUxvaa0xZoSKcmsHRBTx
YsK0mZf148wc1VqtTLSgriJiN0aO6RmAdXM9+GL01IwV4Or5ucyG1iB3JMrVk/fkrMAt9FjiDnuz
DV8d8RfgtQjtljYYE3iZONCCq99fWRUWOru9Y9qH6FcWh/TLDdTLEXe9xDE4PUFCEX3oG+sN2T9K
ivhP4XIvWEzVeRsfgNCbXIAl423rt9yMHXoxLU3y1FsfzPopmFzD2K1UDJFlr/YA6m2Euab4a9xD
Ell/Gh1KRDP/A02zyTYAUP/ofaLWf4v8R1bUEYCHUPedrplUTLHLXiDQs2xhh1sxLIi7S88NMRJh
/mwnDdsmAywwd4hCtmNHNRG61BcnaIGG4OFoJ2fJlrKYKZCBNb9Bff6H6SfstoHjm8b8g89NQ1Bf
mEtuj5aIJ0ovsaBA985SkJeMTSNq51hoanUIXojjRE2+m8MCjJg8nDm/acBly5QJNk+BrEGP7jGx
r0dqEUpmhXPft2tz7bU5VqZLpNBM2qVMbmvxV2NLkVcLKnqbmlumB/CeGV1YsKVq2hv0kXVV8b11
rvPwe4Z+04chzzC937Z8Meii50dOVTmS2giur4lwpeqG2jhkbamQh+5K4qwrVQy64dvBqg66kkg8
2amiBQMaG27CbaXaIE9fEOFUhOMfodj+aygyUZ9QrPoNiwhTQGpjBKUoohj66G73OfqbInHbRK1i
a425N4jvtA6n9Xn/jzgYxZ/WZ5LVkLmoFqrZwut6blEh4rfE6+uAWyXHUxFIo2cC3y+MlCpem0xT
y4tuWA46C+Fo9BwgeA94CRvj+7wexCsAoH7FILvtKvG7ZFSi3uaXjRKpbV3mLAvfMiH1FUORJgNW
Q/bOeDGLiKizYfO7fCMwuI1DiD8F5Vbtc6lLQpYhJHJ8UZUJOuKgeHBnMLjQCxBe2aBE5nQNsadA
+AjzJDdG8sJb7P/TZO8vBMIq4Xx/lUTwO+ntey2bydUbZ6MlYyHqChDU5PlKuK66Vq3MN5HsyMI6
458WOlkVAsdEVBlmFwt3+nFSyFt7Q65VLndsSmZNV6wP3XS4sLRLIji4X4yXI8Fm7NuamQFUzjL7
OwxunNAI+H+LgZ3kxafrMwHO98JEQ+KMp2f6DgffDcqacMA7uC7NI8YMs4MUOcWNvkWvNwlWOviG
PwhY0rvQ0awyqvMhj68clXgB9dFr+2sJoJk7DZEjoVW1JoXoCjDhkm80hIIaEQuGXZ+0tmagiZFd
WGnYIH0fnJiwLCIfkkUaagOnwlNVFdDEJ0phOwHs9IhZ6M4Ghr24ufPYeijkcafDaySutEZSD4Ey
rCoLDe2BlVusKFFyvJLYSgfba/wiwjeiuv5dPmwuTLd4y+BqpnoH8UowK4q7FliFhpzx8qxDKGkF
4QCXmgWMYqNLIhdBPGkuOzEZ5v93TWHSTtkAb+EsqEUUqoLnmlEESrdbUsPiatKg1d8saMRPPj5z
d/oHbPZZXMCUSkm15s3ZJC0V8hYSUgltt53jWmCH75MOWdGYhsaE2PHA/41YDnprtUxa5iIEtzy9
EY5DjDRdSnXxOWEyj7rf97wbh2EnCpFjR1RW2LWI+Ydu74zV1v0EGsQEZavWsvWUG7MPgontPRcM
L6A4CW/kD07gqTZEURKHADiDOok62jlxYS1I6/ADwq7vV80Bas+0rX6ykkq6jya7+M9otGGwxeDo
mULxLCF0fJG6ToaVFXp6HbcUAp9HTRWEoKMMECDkgW1telf85MI6I0BveqFHvph0iLvAGsXZ2O8c
v2EnFuWdvn/JXG+t27wLKhyoYj9UJ9HVietzk4NqJ7uiTJuli4xyJjTGSeeMJi/XPgEJAmLSKJpL
BtW8z39aKTU4pOPwVfoIjn41fk0lN3b5q+z0ztxvj6kDPjpACr5+oY5xHd+miDd941Nksg7348ZL
GWMJZK4qFrqCcY8fFWfnfgnnaDIEBdmz3pjhhlTfByxlpqFDAE+eVUj493QknbxcoF3w0kO/ro8X
GdYB211AJzD2yByYWyqsBqDUqWNZd4zuDcnxHerYgyPv1n/AceiPcWFDZZVanYC2AwwMN1RLVzQT
wn80lcI3ahZLliwz9orRWt5/9rKjUs9eGRy2+zOPWm4Srtb1uo8xAuR/yybYKsKu6FA5xBvZDPgh
FGIyC1003bYwmTiztZW8vBKfDI48SJS4oa4AnwGH9zJc0IUyNUHuZdX58sCdxL+hrQlfeG5bEn5K
xYqP5T+mSm7LZQdqq3IEtRyXf6JQZM3qs/BlawnZkk6NgS1xGAhAkPFP39NdO3y+uZ1+IQaQcAAf
Z4K3MtJSQPIjBGyjGs61HO6u1JumYW3FABAunZAcBXboMI+comVvaTiYrqIdoZBXbtM3vfpiC/54
73cTrkbYuA8LYUu/ejNeDjLZGPAoM5p635Nj3Mf3FahyAkXfGC7MNvxTWEsw0/9AWts2QJx20cpi
95f8ekGRcn6BLI1lOm2W2QS22G/S8FO0pO58GpojHfn/JmfSfBnUNIiDjKChuL8tZDVedb7gCVdY
fg5oAtbYpt32ma3EzYXHwIsdO/jM+tCZTGLiyacErofTcogXpU/27iBu8/gWq5T9bi0A9Zc5+qLl
jPf48ewZixTIqI1W2ABW+FQyXmdY1N8LZpkeElYw1pK9qUkT6cosSOt2pRQyetH1VukLT68+BTEZ
KPeKz7iz9fbbjgx791sV8iwaKUxXR5lV9QAYeMPmIDWMeARfmB9QPPP7JJB4CkBfEDd2koIvN2ON
/5zbyvjX5beNsIX1w+lH10zu6I9Iu+IX+k941f78Xdjoj/1GHJ9D4oxr89ieaS/cBHIed3O/nZOp
LRxuUJTpyTfjxJtAMdlc69entcUyGz26pP6s78s5ToV1ezBF3GHdT4zqzZTajRNd4amWRAqKhy6Q
CSD2Gzrcxb3pDbSiE/5KThmNCX3KkHxyJ/oyEp0lPGat0TdC+pOelR/8PbUROr6tM7H2unces2C4
ZD7WTpsF3MXdte5rTOoMSdp0Isx+H+1ydlguvxxqSI0NZFlSGTOImt2x5pw78weiz7XI75q6Ure1
K21CRNhh0UHaGVEBBnbwOd7k4ipIS3pPRaHKTypPh7Col/mS5GZkM/BOBKROk3wAW8w2S292b9UC
4Zw71t8CtIcBmigEnIvUGPCOkUl2fhlxDzM8Cunuo1OAYDs/IsPsWovP//wY98LISnxlCQUbGx3k
g/llPzy5fZi3jfwpvoXMC6akfMkKTbloGd47kbQ2A9py3+nexe/Kvr5H/HoN4CX7azI/2Y2SMNGI
y0Faeab/zEiqd1oFtzJMtgCfPaJTAIfyQqY4WbvRC65mnN49/ss+kRJ2tCES2TcxjC2q0LdVUfNR
cG6sIRLRvNGDnKXUhpIDoulp/ulqJPD2/JtbaZWZr4qqJAdLvf6CgTEci48IPfV2sWgqctBix5jH
9S/bq1sl/bZumCpw1+IZvkuvqAfHIoG7igkYC1LZDLlHN1DSwc1GV9g3GEM97vnFhigwNBMDl/qS
j9lbBPfCQbrnEaaysDCdUDEwbvedlD6XkwBntQ0HcIGFW48OYsEa2e45IP0NsHoX+0795JmAlLnO
xwnQB6onNNR7fSgvXq7tFacsMWodAMbxSNjIUUW92jA1MOKH2Zt6zB/MP9qtcswhqwVGC1w0hnDW
oiEAzPoiuot7zhAQm2e9hc6Ss2PJj+AoqFn4sGvslr5jK5qSYnXGWHxJDea8vUgJwle0C2OP5L/B
79ogGyfLLGcXNRcP+/i1Gs11FCxv154BGmrKBFusGrkQqr/NfZRohc0FO4QAJN/9tqLRSAkhenh2
6RWFrcgzHKarVaEaYnmG0d7ojDdgy+nQQBiKj5/2AZtXxZOn9WdiKBlTi5RWR6CukvfWVwqfmrh/
Xf+xFtUZMy6k2SUg4kySLAAGdP8T/R1Hq6D48HbUg1kljKA8NzzK6tF+LZT97zIIv2gYc/z1P1cn
6kp80cR+KtrPSbN8Q5SARLxr19Ekdi6t3Iq4nJwXigR/nLjOSCqvZHrbNgEZWqYrT0G/Zawt/dnd
jEQcus7IFlR5y8xigf6HFIXW/42oIXe4cZ5wX0lsTXmbhAheeixgcYGH3XscuC47YdZYXUd0TcLn
xSvIMAfVqq4xkfKflU/qd3x6wq7ALFoWZVQV5Eec4eioyenm2AuBo+UwRxeKW/QKmpfCIYerQ3G+
TaYFYA12H8+Gdl9w9dOUG8hfgf2I9V2WOQqoDMaX2IeOSlX0nLPm9N3+r2hPw0RmXQnYHDfFvoH3
TYfIWFlpFXIxO/jFp0onfpn0OxqidppUf7EM8ukrnl+kC53pQ7CmLbEAu0Lh/EhuuKXj0vyI3dHX
/KlF1fpPEYjdYJP6+u1PVRZLjN9JKwmeAXT28RRk9/ULe/qRCAgTy/pC/eyPrnx27qAGOZs1qQkt
KZhMGJTdyM1Zn9+WNyMOqYhKBqLTpJk4EmHJYrVLxk4XQ9DSvL0//KY8N6qXPto2NLAmzaQFC3q3
YAuDzaSj4BfFuKOLm8Wz6Y4GomW+UsxqXoqaTXcIifmHsrEDN6/gwb4y+eCkPi0czB00e4mEkv6X
e8OB9aKzi7lRd4FBNfL1TjFuKTzFCeZRFQXk7w96uHripmaBkjrfeiKYnjIjmtDaGBro3BtBqHe3
9CYESxTgpXiScL2nQmbBVBAHBMl8NIsaLrM7NOMokrmeiaffnh6QIX7tRbpiueC4gHK86Y+zKkNT
Mx0vfIMZAVM46xOVYETVUwSDZRJrJ82ifGvstmdDcBKb6ParC1nBTrppGGR6WRiFrWmbL83Q5PFj
isl4PM/k+W/pkB0biUMC0HwnBtbQHBw9Y/kX0uYGuCwdGk8vsITi4SeT2xVKZb4DMEvAGXfbbq/q
QUJ8uFw73i6w/1sIMPlxFm1+JV2darNwxXoB0WwDRTmkj7mIIpT/ILhOdOzOcvakXPqMKKaxYrA0
qkXncjEN5wScWyapDluYoxGwlI+hgcxV1n9qDHCRjwGAnpFgD2JOa7znJ6K1BEt+pzpBaKQZaz5W
L3SFwKX8puhvcESTLDNu6V3WYOh5ngD7OWwucAbGyCi9OyTa8oa8JQ8EWWaxAGZuypmtVGKuRsEg
aMluKaM9OnE/VLwlgWtmuzEiP6oN2wJCm5rde4Z2JP3Bn38AOxFxPX53OEkD7vV+S+WBZ607cSCd
I4ggcaHpEoLILCtlFpn1jxlB5N+shKE0bhr81Ln/LWCb4koIB5pW56eOB5AHBA2gdKN7WCRxs7sl
gEkM907iOVlLaL5tBmW91AS9KqMBW4tZbmMFEWPskQr/2bCfD2W06+BGLAisqhkSGl1TafXN13Z1
g/wttPoOsUuwhbSZIw2OGCzpIqmCvh7becZ8A5upyfBPnIZg/NHcuEG2aHdtk8p0x3cDA5DcP3Qd
aZZka8/J91dNsnYJnWf2oYktLtA1zl+XUVg1Edzjg5Ht9PH2qMl6C23jL6X7Gsf9w+KMFyAvTq5N
+IfUCYwZky1VDKZdWOq84X9/Vph7EZqscXQ92lSuThJ+pTdlFeKX+azNwd5nDPPa0xWQOFRvsVaJ
TR0SDUYJk5pdAACqy8suGxs6xNXbsQ5zZ7fE/9TbOd5gtjKrNGjkiwb8tJ2ZRmkvQxdNYwOm9/4G
Eq2e+n0iwIOowJsVuyKwLQVaVWvmtAxqp6fxs7nKqm+jd+NKrTN2B0MwEfNq0s1TZDktQCejhutJ
3anvmhmzPOR7pi0M2v2hhS78AgnCWx8I9uM68oGJ1FfM6h4zvVqTbB/3qh0W2tsNxDPXgTK3RgUb
b6ZtKBMD/MP9oVeJWISIYauexpMgmW2hLZTIRCoS+K5c+z4qZ7X3/rb+E5db3JuYJFutmJpdfK9/
A2H5DtX3XTzr3HUOP0IGf6fRu3hlM/MmWM39CTi6xrVGnxK6HO7mTpp01/QI2FpWIc5g0A/6zvOO
iUxh08dveJ0eZv6x8NPpVQKqHM//8rlQSjoAQfVwZRpyM6Qeb3VUQhQtal8t5TRPat2kDDv0E0wb
uZylIanAgeqeNzrvBW1EsPzszCj3KRZX9+L8jjPhkM/Zvc+EtXvnS4By6j8lphnWMY+zmpVgmshs
o8L95Qzf5G1oPzZAoYwv5q9h+Wj71fQrjoaoZrhtxftbCzbI7pIkBPQxkeT2f2kcklabwMF3xI08
eJAde++KaQdnqSrNkRWTNtLrIG5hF2Hngw7uv2out5Omr+GNsl5x/jdTv+4hBwejqb2gobScsobW
ybHpD104ByeVRA3FmFAjB081hYJnPprN8+6IcL2dySQDWQOweLr4kxQ20U8VMK9s9XcPy46cs7JH
xaxXDkoUqFHQTFLz6bNzcKbXw0aojii5gKj02El4VceyEY/oGfRCzp2Y76qAOJ3qXcQFJpMz2c46
O+CqmB+ViRbzY+I4j8SLYKuIHGv3Cw07a6yWyTRHToWHe+FbKzoXLBSXFtacUq8q8nvC2cI2D9Tm
E+/MFigVzjnjVir19o/afOgwO7YAb2rDtM3QIwB6zCsN34/jKt1tpnQ+eFm8o8OkRgZbV2X96fkb
qHDEDaWdLOZANqSk9wAt5rSGE3tbbJ3PVBe98Blpp2y1BtxN17qCSpEY//55/ikIK5iHoxVOaStJ
uOowHQRlDCoAD8wEzaudz3gaSshlPyEwvck9jIOl6BKL2gC8CLFGT5kD8sn9VLeu7r28hPJNSs+l
/MSddeqbX+4G10EpEkwj/lf/AyRWQh3JokUL4prCVrhM9VzhTVGsq3J8MY+zGiNyNjMlwEq181jt
Gvcm05B5P3qoPdhp4QHh/kurgChx8wRHq5y3XKBJ8zRMgeNxsSnEJmDWDVyZ1UEkILEC7+lZHbi5
/XIr8vNzyTlfz0F+kwFYS0usYZJg57oOts9odL2hFd5Cgp40ozgwWFkqIGEGJrFZ8mMtNJYFK1IA
flpa4cXB8EPkfW3JsJm49mPOVYJbLBh1GHBUsqVwkj4OHuiZy4uSTTVrSUeh2jrmPCoR1K0CLsi/
PG1dp/IR0cvufSXqDqtjXt+gSPk4IDYUlsQulC2OkmTmn+lulOv4gxxyMMl3AwO/1nv6hbZQrbyM
DqSTmq+2u/zHsWwXftpldKIlHYRdeNgy+T87IXurlRf//AGjGfple1X1lqfqMUjtPUjECm5WmpQz
jw553sbpw45pbtk0C+V4pcSxHWlNk97fxKF9oR25MfgN6+j0Hv54yijwiWmPGAkRPG84mpw68vl2
i4XfFigbYOb522fiSs8bujNJSYZMH92jQxRiMXEQ0IZf1ezlDxzYhcmVUvTLDOpKBN6aIYd42MgW
0lW3AIsy3QyIMLo+W7PAeUANm0df2hIyXvZdcnW1NfTUcTRswZOpV4HL5gLeChgbwFa1p1cwPk0n
yisDj3XzzWlB8ontGBhus/v0BfXesI9SByVX5BRgpOYVqhdbmVRxsDTLz+OXa18O5jq/DR4EzIL6
NfW9eLtMO6p+iKJbz5bQN/VoZbV3qGCGa8w0HkNNoHQCvQ+M893WGXPO21T6aoWBe1tI2DBFEvlq
Dbcrai3ovfZbU/5HYfd0sGX4sInoBTyWpuujP0tQlLCQwsaigVSUUstwdQOou83dCNNSlCxa+pHa
JlF1j9S0exqMDj5nOpM3vMq0ty/4lKRULbYqDjwoqH8hrwfglkLO5sHw5lihTzD0wpwV6lp/D7NA
LgqtRkqlsrzCB4g6GJZX7NZV+ANlOyW5NruJrY6Ev3+AgVynKKJ26YGMCTHzTMvyhgVcdk2hWKhm
JoIqhcoptjgL8w4jcBPaROsk9hrNPf1ehduJKtyJst2SaxKc6cBrZOjGq5KGP41TLJSZT4LEy7Sw
3AsIxWLOVGziyJWNNisnPNzwOyA8fXfmv0ZpDC99dtNtM3C1QEZACUvtVbEabcoRr38CnlXQzEwq
/3/3WA6pbIYHC2bqVOaVhG94/UiTJOrzcJOJ/9YJCEKTDmxi9Vi4gqh7QzW5x0NZMj77+a8sbRBs
xxUOzAw1+gHSUDN54vDiGgZfZW/H9zY06A8cp5otQJg7DP+i8C22+1KqbUKmKclA1Bi0X7Ofz6qb
CxLtSg1PITal1zmjB/QTfSjkCzXBxYdbx7i9BwH59BHyQ8qroEssNSGmSm5fO6nw7vR+LNQZ6gkE
ozUmXVCXDmlKWKAVm0At7/6M+5aQzySNXcQ/jeiCQTAuKuVZx/YbTkiI68UV5bVQSS5aIuNEdriW
M/5fRpmOn7vlsoVMgCghbvyCis3vlLH8vw1UW4IfujLacnwVLr6BCc4iFhXl5BzCCLRDUuJ7OVVL
3frK9CA8EcFrKsq+LcutGEq6caIr0P484l+gONk0WpUfnmN7EFKXSFYq2x2MXNBX/P9XZ2XhDvzY
+VM0lTtmjUQeF68SkmjIklIPYB9ChUQ98aMY8m/6OhYcIVINXp8X7+TwoXivkegjGtzH5HytMHpn
n7Nq4/tkxW1cCELSCoHOMDRN68VaWCT2SzZo2i2v7Y32Hr+3dgUhIpKXjI+hv6FTN4EIElst0rAk
u5BzXs/U1128DHl0STujg6zxyMmYIqwLKKfJ/Wzp5IdkJ7q7cK8aTiZ9RsrbK+mpOME8fUBhBqaM
q51GZAmfhJZ5FezBelIKfIm340vDjLlOIxna3uqTc+OCPjhhcOLfZ2J/G65JZgqsV4OYkJlyNDsX
fH3ji8dxPgqHxPyE3TBHXM66x//1PMjwGXJxKUNxCF9gvQ6piOKH9AwOjh7s+ijtEzUrmmCeiRSx
lcjOUTLoA5ZFCXGbXWJm58QxKjZPcCuwu+XdNgiRBWlcZ1xTarPVNrcEO3mOeRQxuaS51xg9GMx8
4f8XJ4LaKbi7AjAMskKr1jikSaDB7drmC1uJqsKCXfmyaWhxQmyQQfPKLngAdpZ3hX1aUQaRv4gL
m/XNC284w38ZftxOKBOSlCVPp6R9IFTwz6ZYKy/197wX+nnvYydCbOQJJWrF67ZVFxS5oWREyNnk
c+2HCBgZo/6enyiujm5U6J+MnK+pa4ywLE7bYWp241RXOtL8/2kI2JMDEVVVUhwznLrz73vPJ3Gm
GMXsmq+lBxocUHWmrGkRjhXPtlLZAJy8XN/hAHG8ok3Z8KXjDI1wyFcpl+UAlgH2b9DcMPzW9EnZ
AscLhLT73SGttVHkAuRNjmsGoTTy1I8AVz2CubNcCPUjgv3doxLp1CfTgDKj7IMcU7Dfr7jMPDjW
FmTtRaRxCq6N2WurC2nal71kJdxpmy86rpd3HjrfKl+lULyOBUA7QoFG5jPx3fFqMWjKGRI1ueo6
ConurFCEgWG1hpZx0QLmsyWVLmKB2nK16NCdNgQ+tusiJuU3+3o3IaiBiTjdLMJDshxkZ64+lTtt
WLQ98UCGpp3b5IQW7vZRlIN0OcmeyA6gKtpNgO7flxNe4qj/GZELgGXNahmXtyxfrbVbaLueDTzL
EjmhlU0flmK4DXo6S3JL0u7W+ErFnU4Sl0t3tYT0DiLfABYkBEuBIHPgKJXzrjVuQSsLuhAiBLLD
DG/6d3e/H0tO0Y1u7IRY+hknFbtIHJLAhpgORgqDiUqiclqeFuaSG7DZnzsH4dzSxDJTv71fY2AZ
PhdyUO7JO55kYWJcw9Nparq03l1vPEaU58LNOhxRhYOOi+EDO2F+mUGvXiGR0aj/Xe6aj7pRV//V
uavo4yf76bS2bVEqicpHq5/96pLCJvoYDRMNJvdbYMfl+GhgdJVMyMbiayIInhand1gKNt97Ycxx
Mz2AG7PmLN3ieOFQxXS/MbXc76aBMPkSpsN49f4vv5BygBBJANwISVLVOO28FarvGPZ8vGZq1flC
rIWrWsMVMygKSwPoy80EhTpFt/Z1tr/7Ima1VqGJvD8SiMoUB6Wj+3J9yYZJkWn4N8Kw9sbIW2sF
lejStTRFS34De9ahDO3yv2918x2taE6chPYqw+PoP1TuXTLq3h7yY20Jfga1re5w4YeqBNOm18bi
LjICjMH4FN03Lh+IqTe/1K40j9m3C6QVJFxWH1ZrYj+3zhlcudf0p9peSYxTdc+StQoKFd6udjEQ
j8zKt5YCyLwqgwjqeo4D3At1zPPDlRWX+i397nI/IbqeZCH8kKYjbQb0eB7VxJ57vG6pW9VeOBLl
d4GZYksTzBV/Gtron4/My5YCJ7VQRySDCiQzeodeKkgBMYoYh9uirjl3z0ebwe8HeeFEFEZTm1Xi
wtEF2W/XhlaLXILN6dk/dZtmTyqCRNgjXRWN+n/UGXpmGsNau7XFvTm9+h9wCymOpdq0egcW8Hp4
Cx5G4T88bOKzg6JH/oqunRO4wTM+xj0QiMquxat+PIpFc0p8Aw1l6TFnvL1o78SdM741VSALc9zr
Ou8lNAPjmSxvl8kPDWvXkWsSyykOD4XaQ7lTP6TKU40jeANSbxZdpPV9WRcY0RZIV7GuHM6RW0uW
wvpz6q7Rfkp+4ZCgw4NhXqWceZ9G5GRh/Qqh+aWata6YNXLeyIvK6WF17vpMq9DVNXpXZ5CXcm3k
dbU15Lzk+fp6LxCj/UvhMSPugwetkL4WaOIKSxucHD7NRDO4VFlr7dyCjgUHqfHR/747gplFICdg
ostwFAF4b8KZm0yyKM/Na7AOS/cH+TNwEzp9eG8MuuBj3qerihRSNrBDSUZ5lhQ8q9b6/GNmMLx5
oKLoEwu+HOYaIO79/6Bm6Ds2aC0VKIddt6pjlc7AkdImmKIY0OgU5o+kHJkr2Y6xxrusdYZF+zWT
PlHuwUPtdFfPUDNtsgjlrLdgEgGrYcx8LsW/B0Yp+9npuoosZhiwj17xhBTWJnIjes6ykPB+N6W/
bKA8ZcdrDWArABvHLOE8Pum/cebX1xvfDSY5UIVMrZpbOyb4Vgc/KsmyL0wgVAQARd0y+7NrVXKZ
JLCdZOruIBljoF71FvjkcPIxq11lpgQRQGMBmMrzuGFbUzFcfADR3QVFr8HnarAAYTHGXIjM7XNx
FQhfJCX2ag50KC6heh/WzcRS2L/ZaBc6ivJCYC/hNHYSuPStz3m+XIcpJ1xckRiP/zeL84HjGwDb
BrgaOwjcSVXMBdsvxSEqewfW0iieYTe7mUxr6ucmPRgAR2IM8DzNpeyJQKaztfXEtWjHLA0A5D7i
E2IJCLOMFJYevUz/EcVQ63CI3YAFhzYXCE0mlkqiyAwu7mnTXkWv+UEJ828cO847Q6atTZOuoRvu
yTOr7For8t8Zgtv2L/vU3JP6a4vYudDl4idcScLtcaTRHKMwdTPc0DBeRoRZjp5aSmU6ZHI30g3e
p4wQvxn86fHIBJxaSLS3KCMZcebRTr7yC5hhavZ0rdWGdFSSK2pKgxBwbq+5rOJY9ok5uT7SGxyu
o29gz8SWBwMHzKX8YQ41rjOrOCPsPx5k6d4oUb78/XqJwjPyXXUeqJ1rdKOn1YGp14ErLbQmyfO0
26R19guKkTNRvAWWqHkJEBHUWuIi/q2xCT+Z3v28c1e0YU3Ut3hKzVHGAh2TlgcAikA8kCtB5IlG
AJJgxRHPGnUzx6QkQBMbPwKcdKIAMh2KZ6kzGKuEkc32uRYeuXcPWz8Pw4oIU6Xdm6uZJTbuiSTU
E9q8g5VSYrjkavo3u5OfOiJw82wZa6utBr5zHOfwbd1iYR5R8znIkzhkyAzeiR8XeLo7aVGJfa3e
5cpeOr+tph/uaMe13qhuGFva4786WSgJoEh2h7C5kNfRKh1zwE4NJyFs0i2KsNfeRCkhMjTy/8+H
VXPDUQO3QbBLduuIPLagnRReuTfFwdVrHA2JaV1tnpCfxntJSLdN/N0Ib/Qao1hfmJwHjUJEjpJG
EPoUwZVyATjX8sMvkgXfyrlGstKz2uZV6MOdqV00unXcd1+MDG2Cw0O3Yyp0ve/20DZaLLO6NRqR
dzAhxbLz4ua0FEELb0PUbubb84nZHSyTP4L9kCaC1EY9SS0SuQAbYi2bxdHc3poMfonLedOXAOhI
dsRB8LsbdGtQvN1tcM8Rt1icNVTNuMccZ7TGWNyFSOmlWTwuaSxKYgXM645fNhqknnNFfJMFcaFB
YDm73ynZ134IAI3axuM4fT7ystK9upOvZ24W71Vc6qVOQAeQz3yiqEYATSxkrg3v2rcYBHppgdPT
gNoSVxacm6W0okpFVopyI92yz0g3uCbtBt1wQsiPY72A9F3d+5KeX20GjXWRXw5H4cf+QT+7Ru5N
bmkmpXZeERsFMtNOHDimyTJx1Op0rDLVeeKSemq7HfQ+D7Fs4g046JSU2GjFPRUGo6+XOC/5oHZ9
Tnk93YTa1WWUAURlz+jCGUzQmnAEKP0SWGKlx0ahSZ6fQVxxK4M5pefLlxZaByDtLN1pMuPCKL3u
Q80q3J6jsa+0UgnUGCphqqsfdPk0HbaEl3mRmtfza9dqULbFlvld4n2ggfXDPv5JUS2HvsvWYFj6
G/snFhjeIkl2j+YYg+gS7voDxObWzxbl7zybXsoTneKN4n+1YEW8Z3ps2DYVPe6VSK8BKoo2Qd8T
h5+d09F9lcsNiKvuo1aVK1HnaDFA11zO6fPx6wFqQ7G4K0XPvvcKSgElxTAqmiZYyrS4eX6kWCAc
J58C4gnjbWZe6ROZwlTXccc7vp0AlAIgFBo6p/kHB1Xy3TZWa+XWgRAO9gSkC4XRSDRpH838Y6X+
8KLcdMNIrTzNWxi4G7ulDB4Dex5067lN8MIfBYkv3BvJeW9TKs6vxl8DR7ygHHaRlJLS2LM3h5dl
cODxygKl/Kxa4VsZdgjlTwrGI/SZDoHqTAq5NUqZMi3IwBRnDI9URvPLVLyFXduSUiFUDZlZSyOG
SDnRNLSLNnvUqPSyCpnDS9pl2no/O7SX2yGqTLeZuBKdjUsdA2xXPWp3t3puOW2P+6xicr0ybA48
fgDNBcrQj7d+637QfsGcubernN3QwtX7hHWO9ZRxEhcy/Bo4ebKL+x8Vks86Uf/X+yB7mcNxadeH
xAw7bguQOruM9bWNIsq/HCDUkH5HLIgwYdImkh789h6b7mhCTAwtFQb8D4UidT6mxX8BBHh1CweN
xW7r0GjviYjSFIUMYXRcx/2Le8xpSjOcElKivuT3oVio8F/7KKvlVblqSMsywP7z2ejjmxWNRPye
Q+ZtdbJnFTboaf0p6N4DVDf7n3dekAePiI0xWXgqq7MoGv0gMnOFgbeQueh8++fZQnxxPMbKCqh8
lWliZ5BZh3sgQ+u748R5DNTVF/TegvVa25BbvczBKMWnEscPYTnqIY9NBKB3KPkLHdFFI3gtK6sr
xMrY7UcdbY2BoncYfNC0WXQ8iv1+F8fjRRLkG+HGcrZY3BfJs/OSDXJG2TvFB6q/X4xps7pHNuzj
wy+PMT0MsK6qWtpEqnScg4ZNfY4NfeIxvWUZXMzLn+5lJBTrTCjYwQVAWj1UdDuc5+aIkMmpQYpm
RCCgBgFz4QjIkBLNsFoEFo+hfXae9NtS1iHaC2BuAfapZDPJ3AeimXgXxw9TyLgFSKYKZDH1RL8L
rpvzCGeE0qtT6D+IXxWRfJZjZHsGCGqIuf8C5YDXVGXhd+VLzvdeoYJqgwXBwHM6HgOSct0lsKVD
ePyBJ9+q3VlgaOOY3EZnv6dctWTY8BNMkTxK0H+HxXgmyuP20nLXXtuqoi0DYkoz2vGFWRKrYAqM
kTEHb3LA9bbfceOE/YmA3pAEmpHNQXXWCRpa2kPhz3+zTztaIDK68aodgqHOG9nuWW4aVYL5pHbA
CvJ3CxaupJOQaKqZIoj4/gVmvVHgpFRNk7PHz33hv5Uj0Wb/nx5H5A61NYEHbL7v4s3MYzgdH212
WODeGx7EBPqO/QjMBeS0PBA89Wv//7vegYfNmU9tCwKg02Pz2SVo2OFJhrxtDy6WsZ28XBAKO9Hj
rjz/Th1/IXfHykZ37dXjyHJXXl+mgpiNdL3cMxA+61BzHQCY1tueBmKo/wptp2QxCQuLxv5D+LRg
EH3KH21ivrnPTj9QqqNKzBHbrGtaWf4X7/muJEmF48chF24NAhOKJGYGnBSPJSi5yGRfUJ62Y7DH
hSeZjns6odemhVLEl1l/cKpeXZ8pjZC5/S8wxLBulFEHm85PXLxNFeRdjmGQb+OmoemGe+4IA219
gFGJ9jE7kmPPXehDbkt8qRCOV/lza/+TMhjqvJnh9oXRT+eSstV75lyRLSRmC9OR2w+DvQftLhDq
aCDCvt4URjr5+OpWt25zRlv/g1B96e8Slr1MmEYIC1oaf73nB3yTUx/HT74JkOqfa0xErRk/Qzwh
QQbi+n6JiINvBQsLn/FVBpm3YxkFzby6fRFaYmVeYU/Wh/VflEwHhggXHwVFqW4ZCSXPSp8jNCAw
nOJR3kSyM8rEu7xJqxwq0QzqaPaQlBGHRXmK+ZeK5Wsf5Y9pGayx5L8chckOIBq1gEnOAnmuTjnB
xABoHYLw+4jwBlWxpMAT7/93sYeg65YbN5/EvDDlJgwDtdGy4icSlzK4QFGvsNoAABmVhWKoDz5Y
wTq4JNV7L1ZW/Bkm2kny0e7ueeu5+g8b59aysMq58Fvk0PRKQ+g5ZGfxn1Ym3+ZjjcgiFZgx9BLz
BwwrmQxFll8EgRVhWci+D5ejkoeIlUKeFt3+r63jEm/xBFGgVjem6KOurijf9XQMqyyq5g93UHo3
a8HxoB4uHyvD21+Nv/cisjHlMAbVz3Fb/z52tZ85vH5Hu6CuRgdKnCvwAoM/8dffiKyrPqcngCUM
u2UJiDYmmKZFsIdTJQ/am44E60aE1u0w4V24bAUglp7wimMj0/aGag2WAup1pLYVi+dclG47Huxy
B634yuAPPAWLUiP6/zhl/5GUQt0dIQGxBZ6L89mYJrfnqvNW++Lb9ZVoxP3269mAImkWR4CMQUNx
aUB7DOkJMgDIH70ao0mZpiXLk9SZIDWqrMjpUGwar080Q3tJtG2z0jhE7PVgpXWGOT3m6SpuQfgS
/Dw0JcIdsLLLE7qi3Bi+Pls97BgTgFoklolLXBvn0tBbgmWlIBYIGi1WB2dBGZamQwjYI+/caBVJ
pFX1t3zLtGdXvmWO3k94F7w0Jan3uPV2tTVWOoBx54/+8GbRVb5NqHj2gwigSe4xJYw2Xm3eHkoc
cLvzNV+XSJUKueaN/3xjW0nJKBOlsbMYxGaRsxVeyZRzm+w4x2QgpJAiobJucZ06TJWlp6ib2D4d
JnzYQlU8Rp9KyyqlTfepcbSlaO6AjozjkYYJP5JNOuMLozJflseE989Ft4VYrj7qYzw7bzet3Zp4
tMWOMNqIPruA64b7RDt4LIcIgIKWvPIpFjiUaB8ZmFj2yifwbrfTJ8cpb2qYnIaRCz7zLsseotoI
RnwnmOlooWa/ybnDyEqgBkRVYRk6jQwHlAeM+vQM+gToQheY/Zw9Ux3gIsfQ+6BPkSjsktyrxM7M
7MdazUjmx7viYujyA6BwFuDWDNE7AqNUUB9i2rAVT0eWiJv5kTXViibnmNAcEqDzPJtgu2drtya+
N4mDX59ZQe4SXQAcLhXP6K+ZC8Ovc4wNGADIGOc64KcHc7DZpXL5SIhHVAGDgksFrfRmmdiweUUB
6O22p1JpNZwzFdgKbYbilaUrtnllrArSkSJez4QB7LjnTchApj8fAQDouZkiqOVQnAmPYF+WvVYp
/Bl3CtPgNDhgRgIi7OdX8fKlhQLUcKyvaQbsjJo2Wj84pg42bxGYZY99sgxKm09Ck2qJKwP0aZaL
3fwLgytBS/P1bXtPdk+NZ3agSLsgv9hx1a/c+9g1zrGRwuhnRX9lagaDyiisJFTar/ppp6SZzO76
U6GSnH5t71grCIiSKJ76SK+pevcykYhgcXhuHjuS24wJ6PAPEW6V5GMkfKxTlbF7o74qN8QXuYEL
B0t+Ald2uppxYHGzs7qxoDy4L5Tn9MCtOW1uEqWE0jbqmCzGRDB9CYrZdfAz22hatzZG9uaZ6sWb
RiHy10Ng3Huw7osKSLBd/li58Kwi31sGLR8pF4AV0L69psnwcn6T8h81OCvgLNjTUt+JjWiW4f4e
myMRv6G/bytegM2d4TT/9i/P+GdRvbSgemwx07q7Pk3HyZGx9gKWWr4MHGtXSDQNwS38BvL9LsbG
adyffWOsNyJ5ldd2xt/vvA7VrA9SEKk7usstpx0KG7yS3ZL/wHJUe94o6sz32F3KXzR4nJP3xUQb
1Xu2kJENUCSkfNkcb9cuPP2nGBVkwGcbFXuLsxsxCLN9R/dktTTVh7O8oWQwT+ZyaaOthBMMwuVk
EIGyJhHWH2UpxRZtUk2Xm7oRiTQTAZHdEEfp6fSe9nipHSxKbKN0pctnhb3tgGBipYKDS94uptZT
DqIY3sNSPTFJlu6/ZtwYl6esQflK4l6enwkEPtdiD+F308y5GvXKMr5R7R/XuVfdgD2Qo7j4zm36
0WNemeNe6cdbilDr6aTpD6UkuHWcT/G63O37IUzBH0YI3Cgt8fzEwvuqgR4F5hvAmUgjOpzTXvvJ
ISYTIqyW0jYfOx/RwIxpi+a1vrTeJVvF7ZVd7MFX/4QM+R6h3Cvrjx5owsvI1YrjQrRlA9Up0XXX
Tg3G/3EkRJNrLuj1ebaMTKhWzaQ8hHSH8shgL0mG1J2hWlvmpJ/SnBaukp9waEXAEOdWZA9gLXOW
fGO5OListZ7bFx13SpeYk2J3C5t2wrmxF/IRn0I6LWbDbTAB0FVvJ92bIAj8agT35naVaKCuE+7I
vLrmxYYd2kvbVbrB9Z9+pj69/iwEIsnxF6DR8Y5K2BUIargHWvaGm01fPLVQds4ic76AUilhup+h
/eYAZCNKDDzaZ2cchG8pvRPheSwHLm9N8RpsOa9zEEi97YHPKNs0GDtD+KVO4QjTV11e9EEY5mRh
Tb6Wu6AvVbzS0HxAiTRdG877pAYgNmMvtjGMkeFfhc5e8hmPQ5+mwKggNle+DVS/DxvkcwtVMfhS
B/Oo4cNf+Y6VRy0WJP/kgzV0UeETKeL64iCe3tEosQZJn1DgSyxccR3JEeeFq0wGnEgA/FqbTFGd
A26S0f1WY6at/x07e9nc5gChRj51P1CiZWYLn/nGL+aDWcyc6EJzE/U3xQrdLcnKgkYLfNOLtSwC
NMuSF64lqxopxnghCkCyUSxSR/BIeze7Bjq7RhSpDuwkzU1buJjHd0/YboHgZuJWGZ7ZI2tRtmrY
vaDeCeB11jXuu/IcQstvmewL3kuKTBUVY4YAwebCvZXgt8p91HEHRsIoQjAVj4NrDGA3TMejk/uY
s7kylRTcAxAKY2BygForgr04oiScqyL8p9ZM3ZZE/bdY70BTvvisvS7bwM0Y3gT+Lk0CG9kFH6x6
15YbulrsameGpGas1n+rBO75n/dvtcIQUhv86RSV3hclRSyeLGRRSXWAi7U+kHlfhrWAGNH1Q+Fy
86mI0WhlfPK0zwEw8gHuNe2lf7/En0mU/SgyHkhSSul37ZRgvxZU/6elbJ4LGGyiuOHXNelCJJpv
nZxGELigN0HZq4JZ/9aHK24dPNd7adUnYzvN7xWhsUn0xX4dC8zO2mer0C08C75deiFGwLnhgj/C
8yxj1XlTGA7zhxgt9BkvTUMzcm7S4w9SvaRhR8yq3ibmzHqPKrumWhTVNSVKIfwAG0fzBh3B8q/o
u7JY/516Sf1/bEEuqoVGuvZz5j5IDc9dC4a7VDE8vqkl7NtDW8dGnh2a9c1DuC80tZKzN3WxqpqO
Lk8psuadAG7Ekjm0Mu7k2v4C6Jod/60ZRZkV5NF3SVBXXn/YcPWgRgRz30rHwhpXrTge4bS46FzQ
X9I6u+WTd7ceskfs2poSQmYHPCUwAfFDaOYT43hF9Xm3tF1vFIIe6HNdVefUHPDXU8QZX562J4s+
erkYGiVS0t8omN7cGU+eg7GrTQwyb714mx2DJdHDcvnFLnshbjpk8DJmJkNga6By4wOxACE8gF0B
XkOIotn0hTmn3XfnQE9sDVoT5G+4aDR0AlvLAyZrb7eOzfX0TuLizg7ZUxQwJhDzQSm6DVN3sVYA
Q5PYUZ+Cwsb9fBF1KqNovzAKXWbbKJ9wyB0pQO8C2vdjoMItw/I9qli48zfTfSZPKTr7949vOlv2
p+OBchcs3d8A2+iLHS89p4wFGN8atM2aFeWuSYxVmAeAPnVmmmMPnbb3YJZzn+5+6Y6j5IAAct8E
g/uZ3q//DtfRnp8/5JAdPVXV1vxM7eTqPbKGGln4kl4kJmTP5FJnDCez1DjPqkn5Erg2AsgoWXYP
nakWhFOa2AIgw5xzGDSZZLBNyy36oRfjyRqc6V9sX6RAPFDi9PbPCRBfMwWepPpDmoX0J81DmRo7
XpLeVSZskQe2kdqcEyCeukMtfLJ+/ZNP9p+ULtvKS1bF9AKG49+35R3JUvsitmbOqHK/0HmeQY9p
kJB2v95dcJA/l58n4nXbfrrwjT28k6wnD1pR9lhTWEmDqSPLlfxLeuVmxrFJY03psmK9U2T9A204
FixBK4VwY22RH3fYkJ0YfoS8MhUicyCQ1wOGCTMik3ysOtNvuhI+x3SvRU6ADWcSGamZNcjqkpn1
Z44QFIXr5V/GwUb6C1Th4LpFVeqimwma8wcLguXmCG0nHQTuqWkdghDgiFCfaIOIA3REkbmmfu5a
Dc2tGch7skq2rCPB16Y68OPCPtnfUHGlUZanxj0vCw6PJ/W8tT/GsZ/IgB/BvChSf/9+ieg9zvp4
4rQPG3N+kWCs2IOywEUzE+XiihMOszNfbNMI0SqZmvfHCNpNOoDZJxqwmB4G1ZsqiYCBZwoPiWBd
9A1BYByPNEHgDinXAHeembXUTISqRMl/0TB06KIW1RMg9nXHPu27rGr3HzmSQ1G6R5L2IIinHbv8
7vwWwmZpeM1ILv/UlAp8SfOWWJ3jBWn4PReufCMt2AgK19KzzlTROp6WMKEvM3SBHp7Hx/IYH6w7
TlmUCe0Ro8asH13qVmXSu4urrK5r+vu3bY54Rso3zjhHWRGwGh//hTOTPPmH7QM3ckzUo687akOj
pOzqUHFOe183J6qmylo7z7SMbT9nqH56YUdVT2W0L02o4lTr1X99QgQZbAWz6ht8HBUXQObtwTqe
K09aRswzadFznrSyCqWrj1xACPZdWVXt6HkKGJVBzbdKKI/MgBXOuZXU8nH/haze4MG1wClny3L5
WsGvMunTwCQf/wymWMiUW+A5AI9ejn+U33Q3BcRY54m2WxPi+W2UQ8ZsixCQSc2hd5d27fqgv3d4
X/gEDbiRtFnT+dCJjza/fJS0eaqzNpZna2cpeEUuJ5EYUtOnMwhgHRxPXfGfm1vv9UUkVJGCPLEa
BljSGReQxTczKQznZBfrkvYix7Ozr6+SzEci+NT9GxRl/Im8e7siaixaZUnW81G01sQxpHi6BQyA
GpQoBe5OKmKcEcLu9w/3ktaBQ0J70aSwPa/6XBniAcd2zPQTL+KR0IRk+7cwN4BopfnMr9kwtc0u
gx3a3nzR41Y1lUDLnmGUQXIyYUeWuQ668ZxxUWAzm2vywFPozMsicAb9IZhmL4gA95ycHc2io+wF
/fPDJ8awyba+nHNct3uVF8btaPkmn5UWusk8+XH3GITcxpj5oOKlFdWgAY/EBiwzA+T4HtJvgMV4
CuplOzXTXV6t1frs3gPrSWdkCKDFbcdHmn475goeLzxcTvZTKLPT0jNcbA+bxCd/4RPlY1QuNyUe
HGa5nUs4K4I+ICFr3tySMi3HFjH0xIqURRGsdfWv0Tjkc6klOf5Tj22BcAAE2U2vRcH0LTWNHiFC
pCvweGE82cSPuJd/5EaV+Jh7SmZ/WDkQhi84pMmkQvpZ65DNnWBdzwAxiJQRS02W9roC5OIpWFqc
okAnZRDRSJyHO/W/rS9ac1lbABhu8ke02J5PzDjGQ4l5BxN82jltzFTyipid5FJuk+ADknEtd09v
ifAhsTjLaZ1jNBYVsMmA3Ww56vVjFtqzaRYW3TmkEDsf0n3PFEt3QaBtFO+JKsRSb4O2nTCjchFB
oGH3DtgJj04E5kQsKAfZNAbwKTsokeEpc0l7C1ErGTc8Y8NRIAwTHu4mFnQY+Y/pKZCu8l0HZP2Z
C1IH/LhhoCJOnMFqw+/H+LUasLwlj6PzyCVjSZuBaq/THTX3vbd3jL5gb/sf3/husyuNAqStW0cs
dKx9EHv9jsIBXuJlg9bhlm9W8QeQQRZZE8X/ycHUArd0IuZY+HKHNP/ml7Q88F/Jpt8ROj9AWuA/
Y5kHTp2bputuIJsEPugWhF+JTk/d9y9cGhgkwltJ+tbIfzPhJRZLTcyy2HX8W51foCGNJtFLXPUU
CkWhBBgx/aQHiaxnMF4uEWIv3wSPgjaVlOmubBEMc3dFGKI64GdVEVFqQxYv4J77ZtmdtZggsl6f
WE15pJ/i/YAChuPVl2vlFO+d15CoAFMwaZ4ALU/ITzlY1XhrnbodbdGlIZ5tW2qPNzsC7OORAtD+
6qRN4vYFrgbBkmvW3d9iXR+bmxF5KuEwmlMWbive1cDOY+p0Plnv9+tYhzlxaZx2RjTYsr6Y4GRW
1G1gCwlXUeD2oxb39y/2qMMOCBpGCyHYWdyHI199Y1ouJyGROz+x/kKcwpk3ZtAeh6FMxh1VRAwv
Yx4FK2j01o2hrKZEbtmYJe8+UbfD/3ZfKa16jbO3UUW4Gb4LbTBkJ82HGju9ZToJc/W3Yptw4Av5
ZLK+IWgwJ7W2O4iQUEdCDIPIZNjimUHVoNLQpYcgf4z9Z6NiM5wQhq/CU/w9FamC0Os7VIKJkuqr
qUp2WgC4BTei2tBVJoJ4IaSQgqt8FQqnFDTQ9b24eZjSEOS7OhVzF94FWJxbccJRkoBDwO2EbvDL
qdy+Zx+RN8OpuGBp2FfAGPM76BQaz8fZqbyjBZu9u5my/OEMf3/xviZxEsHqD5cIE/dXYDSzDQFU
xERg56VfgYvTXIvq0LfR1Nl6hi59/k+exGDgi3WTltWWOUtdOQlmDu+B14a0S+D9ayzps25FbfC/
/5qu7k6XFxwsg7xiD1Oa3vsLaEtWSlNafil5CzmHXMgiXuLfbVR1j4ZNznm4Wwnw7wvBf9J/cNMs
fqBw3n17TuvLedQaflRQ4kQm3tgTi8v7HkNR2fxqm2y+I/j8Bu0ixbrVbcnrQOGX0ZZobNPL5IV6
221hkrMtJFS81YsZJZraJYn/DOxCFFbKaBO7yFz8xV6BzNTtDLZO62AfXiEISaquzfjjixy5a7AI
YGwnvqIOMv/CW+lq5hrD6VjItDWkhoHglNo7TqNIBTLOGn94pcnmQXrONOyxFJHfQl7hw35/vcCE
PLpsOIez4U3Taj4vo9X0cVvLTUncKPlK3yzZiZOCAoN4yOxgNdD0L04HKcrsv+VAASTVZBza55YA
Tb2B3KICpWolFzx+hJU2E090l4aI4QDwXj6Xww+QIzbaoLlNMRgGVKeTSmXDjAdbkuV2SnFHAWyP
0U1gmux4XLRdgnuqKlo6EZbGjWqzFB1800pFJHdVqR2b9xkk1mKUTO29ZIYTMlenNuCu83p3EAht
p0wJB+C7Yot0pgocXMvx6oZDaEcFfYnAqGcQAMTDvCte7int3cnki0E1K2vhx3nf93XrxJuuxliz
hHFLS43c1WXjMfDYlaqbi4mtoA+shosusXw5C4i/uaPXQXu0JtXMu3PJafUTvSCw3BLZc4Y4aTKL
TXCs8xoySBe3Y2HAZZbUGEyWJCGKP5feDSr8GQqZahzDK6NYnwInAATRaKeYQLLIzV5L/1uFgd0p
7LV0B/UEgYzdwcSbWWyWO9ZZFKpzFWoy2fwBCFKHcD3ve11WlBURDf/EdRin8VF9T3Kgw+OI8CUc
1qhds5S1rzspak38038Do03Mb6HaVhXgJmeGAimkrm3R3s06A0c/478035v4pet68CLMoqeDn1Ul
JqGqDLLdpaO/SuLKqkdBvA9IQe9nA1BFjssFVEyOQDrqdXMZ43ZlqfCDGelwJKVTcNu5CWQuw10c
h3XnAx3dpGEQLoX59mSnmQUC1XEzOTZrqa64mFhhnxD3KKxc4QyCp+XUF+GIXyocjDAP/yIcKX0u
mbWqm3GLJXdWG1iZfWZvStxSvkTABlHBJBg8bCk7TQ55iuzMarDPOsLvRJp8EumjMkihwMAJ79sd
UbTaXz6B6ZR6KwuMPrizmNdjFGAS3IzEo4DHedz1evh8taq4/P+uWJNmLygpV+4P8KYOdctrgDW0
MHnwrA7uZxIVLn7v3XXIuDBt+brsesyRP3++LANFy23DUhpQBa2ypUm9PPTbEW/79QGKCtNFcsiL
eaJs3VLQ+Jc41lid/pEiJxWTFhnLD/l/T5GUqx2L8TN4Lv6W4nBy6CccTlmnL61FiPMx32UerWRr
uIn0M5mSYTd/VFURDfoi7aONcz1MgNufL5GJAOT82l12kIAmXmxJ1GTLJt6GoS1tkxoVUupi1YCi
904fAFPk1815Lx3cM8LLbx3LaELXTvCQTRBry8+6s9OQ2Dj4YcwhRmcbo+8J238192p/k+hl1Wyk
Czq3hpZS94fAd5NDo9EXWwksUzwr2y9r2DTjAwXEw72j1guMf2KtiCv/FIiPvPFaAIVpPMri44zk
ZV13DYCHPC/lWk4kEXxdnImUDeK9IHMMC9a4l5KKNZMXl4ziuEW/ab/NmHujClb+piim2juZPCAR
u9DbMjp7aeHhJZ9XAE9OPxOKx2bmLM+r9ooOVqZsRSMINBdMC/mDxu6VXqMunEHnNa0p6ywEf9OW
n1ht28FBmbJS4P5VJZdMxRcdUVRgBIQAmJdvAPRiX/A/5Il+umRtU5V9jtCg86XjzUQRHD2FViHL
kk3Mx+nCTiRq5+DJn/Y/SrV8LcTobwMODItTbGxsLMwJokrl6sXbQ11jT/kpQLlRCq9p/60vxF0v
MQ/C+oeSnIcrzNKacWvPyjgoDMzKosp+DBfviTAdIapnis2CJNdGwxf+q20ITfA3pTrMOE14ZUmJ
/1oLiBhLaNcc9EGgE++G3iHMPvpH8HUkczG8T4wEnrFtms9b3PieUOQ2jY/PdDH01s+QxgMoAxRc
FS4Idw7CF+U29//pzkzTaW5meM6zxSMPO1558BNNrrZDr5+BnEti27rmDrPgn+WbzW37GhoMHt3O
3mTAsCfegn41DHMQFg7/ggMss0x+skqVsnAijREQE9wINgoH2xETSkxhBPQfMDjCPugCJVC0FY8D
B0JZiARb/omy6knB3zqnanxXyLo+rYr12HBuKx9KpKS4MZGXe//iu9n+4zIplLYhJGeydS/TNTHP
1XPrmcyJx3afqYNow4EY7CvgdecuZCb2W1h0wqYLGoV8ZINgskc7XbT8C881kFMXFwlfa9tM4Nse
GYZS57PBTTrRghuonXyvqsmLdfVVXEvpAvNnBU7+yLRAHAVja3ET+mo9bYsKcFTWxboGGRJxTX5C
UwgSqX1CXJbhAayQftHqvCxiTlCt/mQTI7tav1c3oWYEPvV1qlES+qOvXjSklTEqwBKCAzIJ2FGn
3U8wdEeLjv1arkDYAJZ4pqRBzboQ3+FBEBUkAwG6zHM1pPspXe8flPImUxAmVVR+vJ/nqhc7Czm+
1juzFkYzyn37D01OfSwOx6KtvLqjfVE9+1v0bAnroksGzIAiKBTRBAzry+ZPxPSD8Vg7WLcf7RZc
O1ogJd2mVFgv1ZZVaC8A8GW7ID99nwp9r9t4yxKs9BETgXTRn2Nn4idxH4NTnFQDcYeeRx+ccoqz
qEigzA5GDAFptdUpadA61b0W+Rqdq5gGU/pLkZQze8oZtYsTYwE0DVjC+j52ZiUlF0/3m9NoO3un
sTP1yS7cMDtAa1giX+Ee2XcZREnPcliRSfzA79V3V83c9g39eObA+eeUhA37Xw9yRautz1r51VXN
dDok6J18rwYaG+0XKxnOzhzxORJcIIQoAU7wwAfMXGrXYzhcEzBdY1bJibjpNQdTgNIayCYbTFN/
ZXG7P6sq5ULm4tdsiXh0gfGZ0DrLsfRLgfWVqT7XtrIuBep/3QaE4sgKJeaMWBtDCIJy+6OUS4vf
KAof//4Y9isJCwrIdbHXUjMG8lObxOrQ6GZLil0yipv1VGaO5DArzKeZR0WcWnubMO+j53tfiv+d
wBIaxfkYDkyZhHViw+7AS5TwMIrSUMNYIdKQxrvbnQEfzeMAJPedV+rGK8gmkX4ozOyx40zN/Rh2
MlEcZyl/+M2pyVT8gy9tA47JSplY3GtD6NLQbCpdHmITGsZOMgaSVnaUSgQkZGw5GI0VLZCq5O/A
MkpzsVf0uIGlqATVm548sGGX87YB7FBRSuHMxIiBQLtFoQdKzFD2+EDgX42tn+G9FBD99Xyu1AQ3
ebaZ6Nhj7Zt1nXl03f2pCZy5Mzsx03O/e3ebGhzWBXzrgES75s42lbfOrcxm2/+CP/V3MR8oGEkB
RPeqJ00PBVmLXSoMH4ISmT7KNCBUMzUNOaJZRagqHOg18JpWmgxXRlyi9b0iG++vkGRN6aV56k/X
8hmMqiezaDO7aWiZQDDTVsXWQgv1214GnGsFtJvXNHiBeSgx77SaOJv84eKrESPP/m0VIOkxZWKK
yQlAIUVK4fIGwbgnrb0+8VFhGCcATiorrLID3oxXupnoxP/JU9sLDRpb6bfteWY9rLu5wRQ7yXvG
CYhj78aGoghwjTTl9kAdT+LpzaXiY31HSU9ek45S2FjjwnpUBh5V7F9+FYdCeBVYgR2ZziseUM/P
8Ivc78F+i95j8UCWRYWUqJuf9pZezFZYv1Z/RXg1aONXKORZLKbcWeKQKEiuEccW14wsq9VIp/90
MeXaf9SLFAeGmkT7yuNIaBgEIJKheK5q8AMbBxD+atta21q44bHumTOII1VM5H2lHxGPpVRO51Ly
eIVDmxXxXzu8PI1tfaZbYhimf4tCQ2SDmGAA7yiPxigfLJRUzilEv4EPE5/28g+2NF0f6n4kMbaR
iZpBm/unNCAIt1sgAAv4d8pTs1sVhPVUDjp4k/9cTseX6WhgoX2vuE5KT2eBZw9MfrDIbqIU8a93
AqSPbwOMdN2F+nmEjRwl3vdfPR91/jiu+skpPsVsE6HwUbGn9ZYprmyx+QeWHh/WZW8Z37imYXW2
Zh+onAOciOPjX6jqe1XNxz0PcpRMXkjaLhgh3PxcafxHLcw2Uh5A4RWsWdJ/+ZDV5gZqpPMlwD0G
6a3qr5QXFMUlukfdAuABkOglpwN16kSGuszMp/yAZfussCFOnUyLzlOGk1wHyDV9P9R391rjKzFy
cn/LdsiLi2KKZjt+xnzVM4inlmmoyUIXBLzvEntOEHz+/QTf6vB6m23xyrrLfHxP1+hWzzSty9zd
QS/zcwy/wacXscaUj5ga5wzmtEzZkPE0XKlpIl37yI0QTSyvAfE2mj921NRXSOwR2JupGV6XMUXK
R/MtoO1biJiRcGwh5G//bM5Dv2QGUnGNyBXUrVNIIuvkB2d4yFXqyrusP8fRShTfBpM3S891/bwM
iS0UwIFOPTwK/u1E/NG8KUy00y8I4Wu8qgVxVWB4OsAns2fR882V9uE2LR46KjsWwCz/+aAT6dsR
PZ6ShoeHDlzTKCBqoSGdDNZWMXNoXK8LU4bhDC7Ah2Zu2/9cr6mNKnPiuwuYG5JSlcJbhj+OE8Ls
6MDnNUgyrnbYz+BsYPSxUXNtb7BKqjZfuz0UaRBcK53XgupYuV04kLFZ8xT96WZgINXrMFaVxQ41
MShRB0gGWVNwT5CWqBl2e36eeOS04fwjUQEzGg7HXoNskKhStBEPMdTBu6YCC7GWoScPZNmYCKcj
whcIRCeCtDqfgcc78JhTTM2oGElek3+NT63SIncUS1cepnOrFZaGwE0S60acq/83GSA9mJLwtexp
72qu3Frepr/wX/gRRrUKZnWa6MqksTDKIW4gnw/5J5znFxdP/BoT/lH4PIhR7fAEWYuAtbN/6ioF
VPoPMtrTQz/HyNfKygrJYUMbu7gkKSV9n5x0Mep4eFOooq95m34Rth6h45t+qIjtBL+ojlQAZeiy
F2otrBHwQl6rVo627cSWQoSue2D6T7HCXAtRMeGLyN4z6asBo5makbRXHwQcPiT4mu7iJ4SjSfPU
xjVc62rBAiu3nCKXhJZJ0NXgOXAWj7VqyDEQ2UhaMmoqNa3xtN8Xnp1vGhKZfk/T9cIlMHpL2hm6
e0vfIM5wIEwWuJOJaoj+pXmixYfOWUcByEmqUDZ3qL+fGofg13XTghap1irxAFOOItSemokUHKJ9
YC6qjrU5gbsFuz1gBySzsGrcSAQdZt90KtWdvz0S8A56FnHV3hGsVfgEn87AWJ1GnMHKG9VwlTBc
26ysmgZhzlxkGUQdkdrX4WdY5S2yUEZpb0wN7mox6jhz25BCMLtiRRkE2TY9k7oCa5n3qiYYMYeJ
dcDYYKdZFwvfCxxgor+JYhOeghGJtj1E/BnaHiGAemdfM10tdpbLB+vUaSTGzXP3Q47RiJYZk6Tg
goIXyKBnAPcVpiR8XteEFRY69puJtTAkgzEm/xEcVa1NnlfjnOVmKiRrJyfEB7orQZH60aQGCOZ2
4P/BlDJZeUL5xvrZ5ae9yNwgFcV3trodHytMDmh5IiVyWJbLUZWQkZXsPN/yswMtRsBYSwxBZl0s
K/HJKTdXPcdW8STc8cVUpr7lq8GyrXTx5wBlsKDIz05RxoOghz4Lsfjh2wEu6+9HGfqvloMOvruE
a8Awn0fW5z8M0nlIdl4rIMHGh/stNi8xyAH9NhASKH5CR7IMcTGuVtQ+AxtYPLZqn4TuHFu3p8WV
wgWKORIL6vG44kN8VI0DXcRAXXMl0cLUFWjcTeQpoW6e/11GWZB6lOmGGk+NDmlxYgH/rDP926AL
JoePwFeMGL2Ph1DMTT/2UjY1eSSP5t/EZh0cFa9UR4hLnJsCeX1hS917TRDZ0Ij3JzQ/FTUwoBD4
l1ksNsSwr0Wyv2jx4xUWIsReY+KlFFBXubWebkDsw/d4enKGDoseb+jLeQXX3HvCUqU+vtbW2JYX
zr2q0uKqVGUSeZDoJhVCO0u2RTtuyMJWlfie5duxBEdMmMiNImidRaqY7a7otHkxZ/QbAW2wptmU
7pZdCmOJxwbtJjgmiX0hhgitPhA7Tfst87HRByUjgCVkufWRvOvqOcBo5pL0Savlt0GPrFMHbd3Q
NZ1Ujrfx3k6P2L5DOdV0ps8gRkqrO9z53Qi/kp5n3cyFUnryUIM4p+2bLLBozgNGlieW8WeeKbrx
vKQ7FyUx83B4iAxOMcIkm5Fvwg9rjUew1iKLTYhfYgZLSJEoS7UuNOf2eKHhdeqdFdaczfzIldJF
xRPUVfaRKoEVSQ4jKu66oHtFoH0YzxtZpkRq2C1euSMLMYZSl+4zLV+BLcrpZk+TEHTmYITBDH9o
1CzNXA2JjyYplwrdZ/khU/r1IFj+eisyPn4pH+yNCdWIuBg0phzRqRuKtFggEe+9aGc4P9DdtMXZ
qAXAZ8QTHC7rANDJpEzbZ3SFA1LQkO7vIY353DRrmh9Omp1vgIGWeLA4hznbCKRwEPtsd4lyRIzk
Nz3GLt4X37Vnk3hYATJZUiw+gWwRefCAKMbE7ow4nkWuu+sx+fOY/45ktZH70gKcwI1MSeFt6maR
OdPeLrAQLUbFTe8QVD0vj/KWiOZnqy6LhHpF/iYM8kTUvRYwQ52WLpCyskt8vYAvH8ReF7F2aSR1
WUdBNOLk+Q3o/eq99a64MmfpM+uevYGhtV+Go1EYqC/lsCuXU61VvO1RONl9cuk361mSr4003xSY
9Fh8lDmHY7qIaYCtBk+n+LViuRvaaPJdneBGCWqnkhqSvt24kdr8ctrTO3gOSKL54/T8rWOh9zsh
ubaewPgDrkCpHjTbi8ag+vu37Z/+nT1QXdvz2wcQwxmR1ftEzyYHBWeYMmIRRNW5fxloeYtriNms
FQZbj3k0UAMa8611bO12rjfFu1RUoRJ4z4nMPPnTpKWwgkh6PueacN3lwK8x15SsWJSj2cAdcTPG
McnRXoFIGBiOK4Jggr4CEXhQV1T+fDlHFwAaeY1XvGo7xU98KhyQa8UOjJGtlOPIOtKtO/RBXSe0
tnjExvfElk9P4hIva6064qTy+vSaEoVk5rBLt9UG0AeuP9PtMCjrsZEisgI9y+XADzuyhRVUdlZz
me8+ZPgwzGvjrHHVJ+wS8na/dW/4RXGwnIO4IYZNfvesjZohJj2LkNvH3qd3lMuB2J7iavN3ni07
58kzkTeRZf7NU7C74lx8uXMiup8ZO9JS8Qy0uiIQu6N0KaLmAx2nHWoEJdBgV3UbfJfqr0PP1q9M
tdX1jlPPM7R5Xe5GtL9FxSXVpgkUQLOcdRR+7ojkdEfg83JnrUFga+yUnrQnV7EE24EpH73EnBaw
Cs8q4GewevbenPAtDZsglXVVn+rGfj92/IFw+Oi5VDJC0MSxredE5513MOg8fP4P0LCqHsKqr6ge
IxlRqPmIgS/Czczyv4hKxfBkQHBgSaLZ9BgnlbKzCJvrhfiIl4EZBg7hgVDeg/D7Xeg+2+zEqi0W
5jPYZod6AYdBhq25daxsC1TCwLoJtDTDryEzbx9ik7AX8MIoImP9Of7c2fG8ABpxH84zu/HPnaap
0TWxj/YWSuCHFJp9nsE/9qkYUGsF579kQQKTn+bpvTUUakJnqykMS81pEGrqSiCFrSa58hDCDQ5W
2CJC4y4DDJ28CRWgZKkU6TUdyKH0zEKcKkxJj4dsj2LulbQoq16Ft5wKHpGmZFcy53VUHUBApbEr
ZhtTaZUmxUtnmYCoK4KFjP7/0hwgaNz7G39Jir8fql07K8mgJur02rUOPy20S4fCsMFT2VLQgcEa
YlDEwfiTFpbBR7+Q8UWzokVKc+5BXb4Rfz4c9xlGQsWGNQKwjwHawXxo1TOFSHucLdhx/amlcZaI
xHhVAquUJjW4RN33xi0Pmd7BUyKN7Hlq3wxjN71bCum6OPVW1HDwL1lRzz8GZhkSDj24dCDcjlL0
UR79FtU/bX39LcqRu48kACPqsJV2ohvMur+5oMvFQHZoqeZaNZQELNNGrLb/81gCAjh/lAJ8WQFl
HPxLM1mUIhJhCtRLyhMfUrs3n3nxEgLn/JRiSWo7p5KtYTh3VddnDnT9XFyZ2VPvLE/tAM5blw53
OqdyQxQV2crua6FKi12OcRGqA9EwfCcNCOzx6T4ZrN3/2MyOpYF02VlN2wHSCwGFd9HGpb7duyNq
kZObvXykpJM8DQhJft1bloIHaVhlrSwBDym8GboAwHWCPMbkGdAZPYaNplGqx2/dEhidW/JVW1qe
rjilfEmjvEA4YBWbHUTUzJLNkGRZ4H638XpbYD1sUj0RGYx5Fxav3ic8IkQKYE1p9ICeYAOsSMYS
Jz2f4Gx00dJ2swaXjc6Fcm9nn0iGTpQ9Rp3qkz9lvp5UYauLohuI38O/RjYh353eovcrweoSCWd0
WMcJ4XQuytYfIkFsce65iHAmnq1cUuqnEtKeaZUmiWEOid1MncVhiyddeHQ0jHfh59z+8N8Tb53+
1odbU7Kpu0HcJbKH5sveIvqhICVrvoIGy+wuPBcrY5TlmCKU4msKplnf5m9rFGiMsOLDu+lIl9B8
jzi0mjHQ2YitUXkLAkgy7pGRaWj9py3so8+vL909PWEEgJZqGYhDiLB72WGL8IC+VQfyAg9QG11Y
NkMFoadEaJcwRv0uMfPeGplJGGpSCtsTMVKpFaJ94RlCIr2R4lu2ARZcvVj/ZvdmngtKlHAwkn9p
iV7/Hm2JAoA1ifkB3F+LNuU5COK1h8L6bpqR3eOulLW68TspE7TbvAhl5YUKAniOBHIDMkFYuzj5
PY3vG4CrXdF8eiHPSbDVUFzw/KAdeJ8DbiKLsjSgQzZBvOG3i4Z84poKM6TpIGushl6pgyKO8i7A
ymTGa4HFrjpdiyQXqaTMh0Sf1S2VfIXB49AbyXvt5V16VE8XMXCXi5ySyUB0amX5SlI4+AwRsvBL
JcwXYP0qf+XQJdLKR/QNri3TdyVLieVT+rldm38hVbExw8VxuHamD/sm7wfN4zCZZUEaf4wMRKGw
B3htYmLx2GPRmtp8pjClN8Yk6BlqvlJjXsY6gxmaLdCxJu6CxHt7rDhPx4mHFqgKaZ4fTfnXzDJ9
bVVPb5y0TknL75zzZkq3yDKv7CEUAoCSoWGBjj4AyTyjTwwC2CuUYCaaZ5aqE9q5c6lmugjSPQr7
fe+aQSMP9Gf8o+hQK5gVHngSa1lhh1ix19Ry/NB57a8GOWn6vIOngBECindtcO8oTYvzX6AB9ZaV
cA4nt/D7umrtABu7pDVcu62pXhYiUU6+f9N+KU0xQniVz+g/MXlrLzOR6CDXh/RBh7m6q2BYTIDB
4C1+Dd75c9E5ONk8Ph7AOCISV0mUQr3eDpnlmT4g5sWfImzH0eQyDB5n6n1ytwddRRK0bVPYNyZK
a4IQ/f7tnatnoufTY7UoeHoxGrENLl6EB7OS4qYgQzPdyeA2c3C6D1ZIwOFh/Nrq2/45xbso8vz8
TwYhQmGg2VunbradhcFHy28KI54934mxVxCBLEU7ObE+3HkixBnCcnuYM3PEzGdpBZ69G8n6Sl1d
nM7oEdQcr/aA8VLE00OZOuRCRQch248JtEd89qFwC5ASGMrF3OLZpzOAG3LrjVShXtS6f3E/HZ1c
lJmBtYh5SodzuS2zWTMFdwDT9uEPRCdwNWVM72aAJCqDRcK4tz6e9lkvsitCGomG93EGzLZQo8HM
yJNHxVvJclQDKwHpoS1kGnznhSAQJkzStSAtJqk1Ulce4WlSimWpKPAo1R+LDfYnJT6dQZujJk3T
Nq6sUUpXy/1RDQaDWnV8oJowj3U9EL3uRu/KlZZHJbxtb2qUET8ugS25xnj37NvhcLx1yxHZYEvA
b0UPrqN+YBqgC1nmFTkmwCYtgUHkLIZ0N1QAEQW1cVssNMNRaW2qdQg3B+BmLfb+FOEimvrTxaEL
tbT6lytYN9zcnxGSr0SpoZwMj2TA5aer1vwiG5o0yV8Wc/v8mvD6vJd0mM9sZX0Ll11rLrGYCwSk
VsUao1Z0m9Q3fJyQkVXhkgj+HLqHNPBizEEWon+i9HOsOFTc2xNDpBmCu5LZ07HPDgixsr3ui1CW
R+GP58B2Tl9ZQOlfx7k6tMSe+YBxh4kPeL/Tbd+F3ugTx64FmZwc2vVateBsBAlYWaP2AnOlFFEm
+zex6v0kluXpJ1vsbJfbaXc8a64nB8a7EURKeUalhEkYe7e3MSybTPZdvaYe/1/7teJc3Nz5kAGt
LekHpLdkJUkqH2wRKytHiqGuAFvor/kKMjald1TQfgfLY3cXDJeu7vjoBsV2qVThxXIrEbSEBa8B
l2P+FlS6dxW/J1d0vNZ/ZwPSGvUguk6AkCzdxycUfgV/+2lIZUl4DN5A2vopE47uTmXKopCvdO5y
ov2jrSQIR4fYzj7ptZdcRR8BFEvr175z41M9oiClMnynGpwHbKZHRcM7o+h0p4UNvnfkS8IL5z1a
zMOoODOwlSVO21MNuu61NUT1RSRR/1d3zBc4ByGbg0tel2huTtyosJeyWGA0vecwfq+PWYO3P6ar
OdXWER4Hq2usqh0/VqdH6YgMalnQlxqk7oDia5wrd5+/eWHXB8OH3m8ebyxiAuPEB31oBRgDP3rL
/4h5fgpF52PYjuKdDJ7dSI5jHV2uOvTjgyRUTSZVQUhELa+B5kPe8r7kacWTNAGk7t1Nq9B5vmKY
2sm4Y5PVoQyZv2YgNROLbdovdLNitJuaar/EjPaQAzcD68SuEWso3xMRo6J8HkEeSTKHJrPqF/17
nWjzCOjUQtbBmKJbAmcngeq/NwY2S6H8h39EIywKuvqHCcYtnO1Mw6vyBbZNFMF/036SUlPpTeEm
mjLJsSyb/6yjh87mU0UUbFsuPXvQlrxWT3668/9HLe55A5olf9RdH8mKcqUCG9cHe0RpFyZLoLLZ
7SDwv2vS6d1LQqyHC83x3xP2wbVoiYeQ6n3mHL9fw/QwPiO6zWZee8ja31F+O9L1Gl9ZLht4QWk0
5Dh6nDHpJM6fICfV/tb1FlyoWKw6UlW/QPLwiHqIp3+RrfeB62PMnoCIdbF/UXn6XhIv5e1cE92V
Sf/h68FvfbR6AO2xnJrhMBRzAyI/1Qq6ttjbZGESX65RFFxjArz4d56pdaR/QBgBZbki1//g078K
5C3pXQAdyU4A2uRoQIVibzcbNvbJogmDYXOWE7AskQbwGqr7kFRvG1BxKdgW5HEgz7LUXWX2otT3
EmUTYcfwF5bZwN8VO9U3Itlm7RIIFqsXviNIcxTQN92+b8e3oU0+BNWkbN28YuVVcxdRcCs4zejQ
R95WYmBMwybkaczudF8/CNCCCsUNQqSNNTG1fvN1G8tIewUHRwoyqmsK/2Ofoqw51+Hkg0/TW+jg
UFg5DdTIVfodmLMCE0jSfeYrq1qc+5qc/GpfEFVmnhAnIcWbL0YSeFuxbjeq/RP43VOkQZsucRo0
YJ6rtkhRM1otdawUzpKhv4LHgk6aaLokxJPdMZiHKkOo9c055+SSKdwpFpJKjLHAmqAzwOgXQQzC
NFR6CWWMmyKz4bXeQ7oFcim/SwglFJcJ1EXatE2uyewIPmw26CfZ4D7WDRdz5y8BvEh+3llGlzpr
XTxw1XdQels2/HJqLQ50k8WIrmFeeV+477su0nGTswT2zKSZ4zlXmrbCpfh3X9dbMB15Fhea0PI1
Mvukr7Nt5a5IGykAuUS3UVVgx3mOaJZJ1zYEj2X6+DEaPGFtwqkH/jQDwLzgIg1lWtvpxxZDxiOC
BrwAjMvYIJEQ8VRGutoEGZRtv3Erhk1YO7ccRVbVuu9I87GDurmy61r3mmI/QQnYjz8ATnL4G9Ks
hMqzUXPAqrkK0QiM2a8tzuPRklaMH6wpzStL1MKY/xBrPJhglTUtlBnGy2ghaqdhG9qUaVordwXD
a9RGmbORXzFSKG1Rosv62aZ8hPmbpPmGeJe3apxlJWTUY4inq5mQ7oXNfgm0zdGLnET3FNGFmlAe
JQ+D45QbvEweKvNrbe+tiOryPGHIR/4asXLnOlh6+F3RG74NAUW1GIwQh9yd1kPiodtlaAj0UXLP
zTcNBTxmGVT+65NAixwRfsfHdqx3WHZOb0nGic0aqRwpw28CDgM+Q/8WfD2y9vds+nnh49slTeSP
weOj96dQZAP6youAMP6twqPjLcScfpNQNNBWcTxbcxgnKE0+mP0+tr1iGqSCfKxNkOVE3L30FY6a
XnRIK9E7gt3/mwP70eiLEGKkAdADuysyKWeK0I7l1SrwcS4cO6rMWpNb0+L330WG3VzlXIHIA0d2
ihAsq1FJ5FURBbGxnxFH2GLhdsmP4vvsgsSG+vIbPs1992BwaX0zrFFYL0iCJa9gFt6kxfWPUhT8
bo7UtfjR4LPs+7uWw506+qd77+h02pE9UlbRlGUxMBVSytsvyvrlF/SMC13gbpQP57gUcoz20ODF
f5qOY7rGuavKqfzJ3olE4iPz4Ywi3e2/GkCX4AN5cEzIoZztMD9rybLZvismAAalVLiBEoQ7QZxo
8FvoI5ZVKWPWRpiCn1hQGBKNBKQg94kJPrlKPkwdJUmBOuR6qsLxZ+Q9JjLBRvJnjpiAI7rVQH2S
5KVSOx1VLnqBn32AlMNEhZ8YadTeOGKO1cLGwMAU0elARIJebJhYby2l2YDMAwKk3HDyjsACi4F6
ZjstRbn0lUMxcPfe51DlTiqwnxOH6TzBILOE/4ZMa/QHsV9nWjIubkErQuVDxhtjaIcBsVetqxYN
UKzweWAZVrgCr0nh8hN2fCMr7b+2ooWPgzkxHUTYuuxvYZdMF+jsThBTb6JnAZjiEJv9zfC+lsh+
bTUCFjkL+4Fz106m3OEUB9HiT3fltOpycSVeCryd0smfdXJFm1sSsIgMFQCGR/WmAqRrBqFQCenL
y5vR5hRDTKcWvXWRlyYKc19RikEvEGVBYbeRUOijXQ7dxCGiQ7AgbiTGl5wvnCA6lkujK9pqrPJf
gdDIV7LRs0+xRZorSwBbGOWg+XWaYKMqi6ihb5/25lfB+rWBe8xuY7PKDUH6GBWFSs/3AYT2Gpkp
Kxv0vYhQsMX/LVdZq447Z0LxR79wrMK23Itfo5HemU/NgwpFWK2/UW0Qi4EZHASOzDBvI/10kwGo
lr9ryx6QkUQOyTdxgTB6xLA9sHI05EeW42Sf4hd0E6Gt3bd5uWCDYXnfzSSoUfT+h8jo3ehAkA2p
/cOTBYAYtavtRhYu20Jq2kfeNDytad7fvBDf2yLtO5mpUidGDVm9gHTamq7kbzQA3n56RwFTP+xo
K1wVTGw+hIQTtCNt/0QE9opGH5hwgkqPmCSNPTOtwY7RzeucND0zcMGHLjHJEMTvUi4wDW6emejx
UQO7MvWHUjBB1Fs80R6zf2UXfO8XIUVy6OeqcWZmjT1Rw3MFfweX9BLVkkNC4M6ryf3Jcdz4cys+
FFx/pS8d82kzK7nE8KA7TcLlyfeMsddNyPaRzFxxWguR3bFOLCSSBJ13oSwPl8gPDLDffSUHsU4V
HxLVzs4IXY6xvEpcMqxYnSYaqPs0BLXIChJV9p+5nZETIfqIXnNBPYdARB4lCRcasLOnGeIEP2QW
cRfhkRtOeM7u6dsxcD2BPkjBMq++Tw8pueAchhyY64oCytsVoaB5Vm4cCViGS/oodbQFQw3+Wkha
/Fqxkw3jdNOz+i3v6VOu5kejcD3w2Lz+bfoBeH7kRxx1OyrqyaRTmBFsDkD2uXgWq1CLt4KFSuvj
KM87ksUe6VczLp8Uxl0O5Fde+WPcJ4wAA55OjPFeO5Fcv+pOX82uttlYCAGqkWN9wK4BROddiwSo
a9EceTdu4gAuLPosKfp/434IrkY4/IKkWyGzy5peUkvYlWo91T23MlcF7Z2h3xqR8Kj53aYdBF8a
NMONGBfHaQYk4hPGatvHpvHEr1+BRnBKKueynAJCQ25OpxZD1fT8Pi34t+fJUaXNoddh3JRoKWeS
e/YaGsa5745/U2cpY80go3BvlFO4mrvYAZ9c9AAQLanHh/cefVxnvMqWpsJRt3Vv3R+oWDdGG2FP
gHsibEp1IArY2ga3hacmO0wJcgkNZLSr0uKoaq54agwU81EglBY8AMkIoheuieRiA587Doh02lPY
0vW2XOk2yU3YxgVoYOuhRO51Wo4TcplJ5PlLKJP4BhfVY3wLVtgwUFWTfiGAEVBh0KbV3BfYU8wd
een7Mgu2J2jspjjb8+0W/EL7M9pyp0QP66+s/YHGGHuDx+Xwb3XxIMPqzdKrUtEDvk9mESCErlqv
Rry9zbmPjvCQAZiqNI/MOtrq8IiBBSANdMgfvL5Eltya/+oy12kTvhj1JXag5Abdno5c6n+dKD8K
RmADuIt0aZmJosSQFfHjQOlC63ABdcC1MHPVMOMdHYcsSYXKwgg+BOqAGnIScjPro3DClS1LRkH2
tKOudXd5kmsJ3VhQdCrE/V6YPrZlOFwAvpcad3BYSLV9/dY8xyirh7ORnR80LA4MRzpA9vgCj43o
HLRZ/tnLvnu+d9qVdXJv/753DqZbiI0R5dr0uu20Cbd5puuPX1zYk5iH/FyeQit7/kteT7UE9KNF
836VNKjIktPQ05smcBzWGCx6bljwD9CF+mgM+5rfSm/6IZ19aQaXkh1NeH8xexsTlIOa+HbghTJK
mH0516nAKfEj0NqzCTpFdFNUmv3HXmleXorZDY3zJBRVh/tk431+GQBGFDZd930Vdo5TgdvbeqB8
nTuBrFXvR0K2S2lhrjJd2dhf/iU/bbNf1fhI8MVgQNP1sd3+XPnbUu5S3s+AG2bkWqlsCQY4hzIu
yUr7rj5GhdQ+ovL45pBYtyNV9/GJVEdUKSYGgeZpEeUmwINfCN3sijMydzwHFpSc+391RVc3MxFd
PDo4dhAJzJobZgHw8F0snnug+zqXFN+OnEmsCktaF9n+5gHxCd04NHjeXx9eUOLl1cz+bpilUrIa
ZfYPjeI4DEliHTSFAWRaB2s7Uv1PMhu21EexvVdcqu0Tct0Zc3+88I95eeyJXB3/kSv3jvztzcE+
ME2FrHQIsUJ7zpFkNN/uoXy/gJR+87p8x/PBr95nRNk9c05CPTfacAVJPrJBf54n/y1HUbRmgbzF
IA0JxS5VJNfGj8BuSAon4SPsI66J2EvSOcba5EJ9ZLGYFCuDhztr/J/JpdVmT++yUO2ety4DLVpA
SGVOskfQIjIy/80IOvZuQEtbMnkDb/xUwhroZD/AKwWTDJ+4n8p3WzKEpU605YnwDHKSP2MJwUZT
VXtoAMD8raYsnsharrzVQJd4aiBYaqZvyM2ddK0AldU46P8fI5ti59/nwOijrLGB8ztoeEkey5b6
y1mhj35GjYBRdf5T322WnY4cnNYkwra8QYLW26T+lXCe1TKiHO1UrBSww8WPwRKrOfkuJcRcZMeH
kFCLgGrKV+ZnsVYNdnaoX8JvkQrCzQFn1wPhLkSira/NGGPkupwKkD6GZTm77NfI6v7YruFek0y5
2cnzxMEF6AYm/clTD1I7RUr2N9Ygp6wZzrLFhoZhluseJM5IewJhFbPDgQnc1iUSpaO3f1s4jmou
KBcIqiMgC8VxOpgk4AKeJ1hpCuJgN7+N0wLZwswPi+fqg1JZ6E5wOYOWacJYlbm2T5ttf4CVbi/W
G6tIaydZTQl+Dc1LVS8ruB1Kze5bzsC/+uT+1vZr1yl7ZYi7mi0e2KrpE6gFA09LT/obeRe0Okf6
rbsDE/s0Ap2IUMS0PG4Vz2BDVqqEBQ3QZrUdqpB7aifaRxD+tgNYcD8GaS9rjwQeEyEX3pYLePyu
Cv9G8zfjSZ3IP6Qp3BWhq7u4Sc+UJ+3hV2MTPxK0z3r+485w259MF03WpnIBDUxOsHuRDbgPM2pL
Bn6f8ipDftAq2CTLjoZRGhytAmiZAW1Dn+gWSEZ+vn5Anw/ggUcXCl14nT4LYllAdyCH4rToxbg7
OxO4v2RB/5BA5r5NxBGzcE89dacLAqO0tFUp0Dw3c1OKcKzZf5bFxW48vJuhcTpSTM8u8MxcmiiR
5IbJCrCRTJ+qKRGrEVMCFfjEd2AfZTgmT3YVWG60kc1hbGIQPa2ICrebo2GhGegykrUc8JrzArRM
4sD6KdwQOf32tPcnTWsNGkhopv8CpaHumDgByaZHJbbKLKZc33C4pBuMGlEU2m9mUSUgRysDTZxS
H7C/2Qi7NCrNoShUHi8TFHcR6zJgXL4ulNmKON4c/Up0DdepLhVGAsSf2Nc/UwYMmJ/kxf+YkfmR
vH0p4Ia7boL+o5/PEhUtGGsnbp315zYcUH9j/pWMkHMepoKgsJUSgXgpsx/lKyzD/Lb71wTlGcNW
1gqBUvazJQByYcMDY9L+maw5qxTVCWYDHAFN8hbVKSnv285NoOhz3UIklUB9XQC933xCvFZZiFy3
YwqqRqp7Vh3RHNHjZ5jX99RL8HboIYVA8ghHJZoZwif1aurgidrAvV+MdleqGrsuBs2CbllJCL/A
2JNGaJBqff7pn3ga2x13byTd0icdwdYJ995ojmiJZCwdUJKSeuq4qbVPpfgvW2+lGWfqEGTcGGQW
1ezjLv8xsLGex+JttAvC7IZiDobMyr7Sk+qcU7zwUbxRfTRbFpUoHpfUAPPEwJHZBZW2bO028a8K
SA/OvfiV0W660tUlPIIlJRvxoUOaHRxImmPulegLy/oxuE1n/3NLQks7dFXSmQqQCYnh/U1vIInc
OxkLcN0PY/AEsY5hLAM78OoBar6IEK8OZYvGMZpWO7Hnu/7dQ5xR3OAy2UOI17sKvFBv+2G5nzU/
FM/AfKLMDX88ef2LCnSGJXcFmwcCTqGLwlKrtNLwANz4ZRMH6WhU24zRwqvsUcBifaMm4ozWAu+E
nNeHtsW84R0nsbjQur7Z0IKBRDzF+4HVsabtaPIS5Xy8998APJilG4C6rTngNenHIeCN/xrYmxkQ
lnmQGdHmtrk46+AYS+kH63xnbgkro6SLQf/RBjqeiaxQt6OUB/+/vzYGs25o3tTopLGQMQjjqMvx
u42KyDoL+2iOB+y9ktMEhzowfW4fKnv15qi/7cuDVlNp4Re3eLO88ixr6yqrBJutPhOj0PN858Uo
uCOPixo6DmwlUZwUs1HqifiEHOgSnco9ndPU7fz3pgOkG6tjI2VImp4GibjJHwHSf8Hsd8GEqzTO
CMME3+KbBua9qmlff7lvq9xDdC/mTDHuWaJ0XdJvVdoSx0GjYUkYJY8JTWTLYk7lnfIT3+xo2VUI
wNJ05GOA7flhGmPvVv3ztkZlSYz8J7uc1KsBKvxfz3bqLbG9C4ndh7bQBA9bgx5SGiqoKj/ZR0Yu
939Hnv+DD9Yj21G2Puh/y5aPU+R33PvMU1ayrTCTTYrmJHz5Os4rhWHUcFXaEsdPyvXPSEnEZIME
VmX6nFJc1I4RMexvNPLTFM7nFSVakQnlCeGzPtAeIp4Zh+CM4AbYvn9qEKgttMOxNgAOiaRzp06s
LNG+VMQ97UMdG959bwiFsdsWRNxdNHUiTza/uOX0CKnyLSTSay03qqcAYPSzOkVcfdZkvP7ab74T
NVYXD5KpmovPDp1D9Bqcm7ea1O145jKZasZWtxGJpJwt1z03fzzogn1M1GSjhdUyPMjcHeCTeNEM
ina8y4ABAO5lxR40+/m+hbK5v2nM50kDrgABG59mHnlhTRDh7tS1SELZqAE9ixu1TxbD+ZGrduwf
XATmoElpHty10orm6KSYxfyfnwQzL1rXpmxL6Ak1fuweIrZGseok9ia10klI43mt90AwgxIW1Cj0
so4ZXwPAw+sRfaZzwp308CsOczVqEEKkAP9/w++SGkwec7O+J3OsBt5QLZLAG5zVvobrHQUN/ECr
WO7MF3lIsQ1ja+ua1Xf1I6XcFtk2zf3kxna7FRTPeCv50MPujDV5hQlEPw/X+EBzY86UIt/nA+hc
FEA73dPGvc1Rp9pkgffCCoy2WigGQLATncn52z9FEAJccfEIY2Zy+UI45VAGN41krxeyQ18cFhvd
hukcU9Lyd60Hyby3HvA+CuEpH603PV1M7ojKg/TG/lcZ3RXNk/a5B1zq7DAX4AFbiWkEqHVRfamd
EeayADtA2/n1pOP5JFU3HZ1L6vJASHYZx85fTyoKfPksFdWhxLAbMuebkc+XvtJ/w5UbVgrMxu2k
+CwNm87/5XqfvHg5LLkJkgMq6mjyta4qaB+yc403UjU/0+s6KNo5rANUxXrTYxviyPXcYWBpur7q
AK1nOd2DCsq1TzfjNtFhzxS+jKMghNNt35XPTCMjfrba6bGaKzFVHOkiBzrQ8tbP5BryCCTIeL5u
29iVQlKwP+0sgz2s0+u1CuknEtrDE0H6G0W/q1T538Cqqioq6QV4s6vTAvZ/VtVLZDI53r6ZDq7q
Nyc/xIZywBCOFnHLEqDSvtxfk6J44xKh9vpTgLkoONOFUwVGINnmFSsrrGvKFG0lLrZdXo/wNuwG
tmOOeJvk0BEz16MnN1AdzvrxQKqWKxeQGE+KrCUqdKCuhgBTOiwap/45w4OT1g8taK4hGTge5WUJ
7a0gIa5FeITxkhPWtmi7cdNvqL+LzYkJFzUd/vLUGTEyMKWzP5TNgZ/vbZitYo+za8hl3VHDna38
4yYDpFs8uqwuDU9zVsaZgr7E4YAz6UfWXXYMeucZF+qrpZ3SZkJHYI7HdrSku5XxUWYHIQ+wnCKq
M0VamztVvkrpUXO0212GhXChUaUm6fa5kaebtCifXnqdvUmvmVqovcjB6TiqTVPZVORAMmOmJ9Jh
PtDz53QY1aWMkR58Iku9yqRiLGeInH0Pg8HhsmH1SuJsjYD0vfqFoPR8ans8ccRLsz8MMvocy4lx
8+eXl/Jsk/pu5zm/NCUBpJlyxqyd67bbd365bEw33K/RdY6E5Q/KfAyV4eMhNVIV8V4VbLuOjYVV
2xI80MO2RhLVQgpxZIPzV/QwRV7RRGfWV50QWYh5t+FGCEAFpwfdGgLXsuJuqGYwQmeicYqgwd9k
ji2h3MXB9+G4VuuLdEce73BIVsOSeGn2DKzUGXvu6Xf727zPK0yJQWxclwStLBdUlC+luJ+ood1j
BrdkVzK0Ej76JvI1DbITONsNisP0qRqoaeSr5MOH1e5Unb8jWILyQUw8kcmbnsWwFd6o7dLTfB8y
FzoZSNbXN3SA+ZeY+00q4cTSnsF1NOKQM/YIbpDf4JxjHTIcWF9GtTQs2Tb4OtWlNqA6xkORAuJJ
nGyYeMP8rnRVMPCx9x7A1DGQjk15G7ifeNz6m6WE7vBTIy6X9Ahvga1QQlMv3UuY2it6DqSLUfc9
SpX6g9cpzbMFNSEDx0kIekbdlg6HLXw2yCdF2iKMYk0W9Aop0QcpIxEYn6On1IUcWEeRla49XHGw
H1I76pDrAnTT21h+aDU5fiBwYP5SnWNTSPwKyl76/MEhrC63Zqp7YTpVwTiK31FLtTJgKTdnTyDV
5WDtX8atxrm8GGk+ifbqK3THtQtAk75tkQsehllug9yCDZkoB9EG3kPewujcS8VDZ/dbQaU9bpzt
Zlkb9bmaxOkL1nn4iPEmKoWmqfXLg2OoFlSVmPJ3dF07ZVfWAW1KBGLifj90dLMLyO4wwtSGNLla
x50jQv28sY+yuFk97xIThsBJUZouRXKKL3YzeH+MkobmltVC5ArV+aOPlZVbTR/OEDB3M5Zl8TPu
CWWsvnL56A17JuZR/0Qyqm+6BdxRX+k/ZrYT/B3g7U+8eltwL0bSWCcc0slJe+bYO+XPGJxT2aRo
toGuLMZVmkICm7h2PYlPHFvmD0AvPpPIvpjEh99TQCG9S3T42huK9EbcFriS2+5IOXJdeqk0bn1O
FO2tQEFsMutK2rBi4H4rTUsvDw5pmCHNXVmsjsU7Q6Rh9rQasjOvtaw8UCIaYd6D69o9tp6Hbbb4
g8aYCSuxISCDrK6f+b4WCXriwZKB9rJ94FjQvrcl/TgQW8kxyKSNHr+MVeZ9aKU+KbxKBw38KkwV
igPlaNeOPKDF2kNo0RiYPrHJP+CqHhi15jzzy5uVFS1M8V7wcjXGIBEOrLKxo9HjSBHDhfwfwyYM
Z0K5LPv6hj1V1ndcn/4pMmYvuV7+gdVyjP1UI1pWL0g3PBlRqotGFEtv/cVbNS/fXVyxgtkGLmcV
VEA3ND30V+R70oGEhdROeLHyrfYtw3xuG6i7Wb6LzwID0LnCaga8QjRhcMtYZoe1OHn/+r0OZ0Ko
PyA7tLGsTz5P1C/Etv3ZZ3T7rpf05gSQSC7bAoc73t9TUsMXZYd+V50R8Om8QqpX3tBLIBlPadhp
UCZVRpSLAjSfCA9Ypq3MJf3JZx5ivQ6nc8Wod3vEuVt+W1S95JS9GZmK+zuFx6Klew747rXmz7da
sdsJi3ACXLLHJSzxvVe/b/BEXkQFL33f5xB6zGEZRsBII5CDyx2zf12FG0zYyETg6CampSoXQTAN
HH41thOmR0WnV7rc8lt97aze2WGhU76pplRRunxjL1vV/dFEGO9snw94TpFKWT+F2LkBloVTtnIF
XdV7tkVrk/dLbSYvpPUAvycegle0YBCieMMQ9LHq6G+9na5l+5Qr+W6yqkYYVHqjYXC/UI08scD9
PkEN1pPrQWf2xRej1QgvgsrMmH3JrPJiFXG4h9zZMWXU9YgfcPFug6M1H6SYNbfdgXeXuylL1LKP
zgrVY/OQOFioip44HTuzkJvRh2NzvtojJE8MBI/cbZhT3iEgz51vJmDMJXkWpozP0gHMxwN45ouP
2EhJTmVOZ/GNWdojLampDuobPt6/r2fXw1MeGuXyqdypIUnpoTRW8dXs36VmiMqxCUaZy18lANfj
/g4Og3nEEFSk1Y2KkmOaqhOyghIDE8E0Prll8vztoXi+Z2Xd4txkI29yf+26Fjnd5PKjIz+FAHsm
S4NLoPgcETqbXe7rVIg7fuM1Azkb5rMdJmiZM5QGtM+jUJDuw7CAsTBTY5q3F0dfd3M8o397jHQP
/ouxJTj13pgbnoKDV+102gsCUhFZqQjDGGC57UYQEqPPBA/XJv7K6L8/XGfhxcXldyjydgd4BeOv
tmudV8elJULFnqZ+juwDKt81HI+PYY0vhQ3JdwFBC9n9v619qLu6rgooJL9CMDh/SChc4TdsLE5e
qz36RGCXTYg/7sI/A5LQEkg8xwDEgBb8XepbMyp5HJJpaUAOFGJ6TtgiwxhJeJ+Wz7YgqY7jO2dF
Nfg6WOdAz576RCWk+7NLnfs8D3/+j+Sep1nRbL5p5CpTi1Y7roknjQwNF7VeK7yu+fyHEd4x0Ra5
N+OCiB3DiamEz+pHnYBEcauJHDrXPLkyuC8a9omUWvxXb6E7+H0E/osxQf0CI9GCmOT56NSnj0kU
CRwFHw7ihCer+Bu6qcHmpzdb6BKH8mIfZpR8g7fS+UJpSwULCzwlFvHI1tkIZ+b7DArwO+GF5A7l
PzxpXNKY7BRDGCO8QnHUvpvFAhXfui3HOHCuoaexi1mFYiGd+da8Sq7sNkO98TPDlhmmkLBRi/SM
z4UDgOsjFqvgBn0hJe6H/qxR5sVHy/3rePwnQ591mDXMaiQYUZf7FH22G6xj948YrOT5d6WrC+Vn
ahSnrwiXXIPjqjb7b/8hGfMZCd8joDpqhALknJ1usr1C99yRPy+yJf3jAfGjn9aRvbg85QnCtLq7
nSGm5an1upAfCefD6k+cNvAQq+160q7CbV32gLxRXsvH6/3MQrXp0hO7REv7UKjFcQQ1deQd1yC5
39zb6POsvZZLXsW3F4EYlHCYEYhCl91EaoQbjGTQ9gQO/7jDzvqzpSMXnJ3Z46a2lRzOAdkvU6q4
om5h5shURw/JzJc530AxnhHBkUFbnri5gLFqRFEkkWjETm8NTCqnfAW8iVetRHGDxU3rrCgttvHh
cJlh/AWSwxG4Y91qyPt0Cyj3LkbjJVT63uaqhbUtqv3gQYRXfismyOhdClSQWidQX2lLNsK1zIrZ
n4hNl+MOI2wDvUmK1a/29I96khiF96P2C6i8DhgUMLKd14IYdRGaeu8ZyXBWSHxxmq1uUMIlKKpA
/2EYlHdZcHtELeLyKspE/8n2hXsJZlu40lt5Q8cMeot3gfqQNRSXPT2bsfktCY7hjNeQtsKCBzDz
GfAzkR2ug4/6ojpEA87Y/ox8FkWq1dxlgILhDrLVVn/c6Mqc/242tSpR1G68Fx6BC98xnySXD75+
9FPSzuNxIvclLo4yqwqWKK108imiKLEYFeaEbeBdxtJGb6P+ooMZIk9Yd+hpuOUhOC+YA7KpY/8h
NYt6WAZgAloRHm7/x35eUnXFvRuaLYA2uYPrtn0vtWSBMtLqHFiBnPhDnWmzuHZ5rfQAgMVq/j/D
wjs2J8ukBxm462HRGV4FAwrMVmmNK8HT68GYufZLGi2OSptSziIxWeaDc41Ez1qvi6ZkEzsaxWN6
Uq7uzcaz+6P6QxsI3tpTc9I0ozFrj2gxSir28IublfdMXG0qhzFUg1E37IW2t7hOhpV19qK8lCR4
kThvqE2AZzii99Ny2fAdoNBMLpYBbfv2tCFAcqfYqctI5WGs/iS9kys4jnJj2J4Oag3i2oC5U34Y
AoWvWdGVYXgNwm0cNOla7oxeHG5JLddIYjKGKknOcXztmVnOgpb+eXN5vASSSOEGD2JzAlqmRdSM
Px2m0YNEMK+zuadAVZ/0drB6ujLNeIymJf4L1u2SuP8B0TcJO23HVL1Tqs2ixhO5Fw/ESZsNA0nv
NR6xcRukTsKfAhVR0FCSvwvWccPI+8Kt9RXZhhpEj9rbCIBlAdu2n2xU1JXpgIODy7BCK0XUK7td
xReEc1IH8djD9QbphxDvnId4p0Qx5G0u+NgQ/0i4FgCr2tjdKXJjB08WXcs0Pu74GMSla1227kM8
kc6tSa9+eXLlkqAeJ547jGJsYKHBjqmd+/ld826PlweZDlEJBIqT2f/12NP6pF5Cg1NHThd6MSZU
CJe8JtY9uFpybjA//3tIsEcWYX5mxa92GzmPqZIHvQyZm/2eMu8w1t3IxoIQWJvO8vWBUlt2RHPS
1Vq59hJvEy/juFbLnv0t/vrc3dZzXFB4RfVNmqf3pe2C+QAtuVcCZkK96RiXw7RgMYD4MoldRKUx
6fEs+4ZGD+u0PkIfLmq2h9U53PQJ0xjjhh2zXPgkbm3WriEOFcw+JMipWcWT06Sij2EQlLZF/ZoP
L+d1jHcfS2pvQsGZZdAbJNlEGd0oCoZgMOJsmmqBIDDLFxEDlfOrs5mkb4UVw+wPmYb1XI73d3M3
3RL5JC4E7BIRkmSVniAVvN9TKd6VMoFB29I/gmKOmHQCcpieVq4cUzVBvyw2UtwYwsNmzPBdvRVO
CRHmg2KN9Ode1HN/nSPHD4peN5t6Pa7iXnWCU3I31CpNyeEGqoFjM2FrWMVC8jdhWe0FDrb3U5Gf
3nFJX/VpbR3HoDLw7NhTjH1A+iBhULucSj/T3cjd5SVE6/swmtekFyGDxob6Du0wubBlwD2AxsWl
/CGz6EDxG+Mv5+HRe9Xr7ND3sydjc2poUpEywYrFIsGcW9vxnAVZsW4hgr/BH0OCOPKiGhd0+D+Y
GZnOQTcAJF3dHUgOR+5YCNChciOuimIJ6dFZR523j2vozxikhH+AfvWKGJ5MEEJERWfgkm5tyzus
HhPoGMJrRWT63tMqLMAOg98fkZ6lD3Fi8+PFdy1dBFXVrwY+Vefct6UR6QgHRBfwNHUqZ9y/JqYC
yNGCr/bGOjEiA5M9viRZAgV8n1rt6CP6N/1rdEoMYlB9G65nE0lnnBROP5IaRVXhDN6Pjp48lyFv
7QDf5lDbXZpnQgz+JXTufayxADKNpS0791EfRdU9YfGNzhraGkim0jRB+8lf4/pa+CAfGaUijsnp
73bd4T8py8MRi64oVUZFcvMcdXNxkAQBUmGT5HMZRC5I+xGgk/w+kb7SiQVB1gPfxgW4DIzgHmKM
VQ9UXCR6G384RpWmCbC1Qsjrbdoo32X0G93FxnP6+1ZCUG86uRtd9XRdbVwAgWgY60NFW6zYxZkq
SPgyj8N/fHsp6b/fl3qmpXZwotL4PQNzvZPJNQZPJoNq736VS3uxdjDLxoXCpnJal6krRgoiDStz
rjHfVGRWSqMF2aHrydxh7QWVHCY+aBHy8zotD7cokPmKQuNeDDO8uKSDBAWtny0bUmjayd+oF2j9
KTDlRJn04W/IcVA5FODkPdBbzBAG2kzKWiK9rWQwpm3HMEuijfOeUlflZ1nMyeKmBvaX12hJ/JEt
vZrDqqUasxhyU2YnFoQbyAONcI3HcXbCmWszyneVUnLdPNbqpmZ3txY6L9Yrgi3+pMN++86rxWKE
OPHowMxMv8v8CpWs9o+qeW14qvqJQu8ScgpwTVQZvkSbzybknGe2NT5sNdRA/ycB8rtv+atLGb9n
pNG0dDA6sTORIeFm/y6fgpEiK4Yf4eGQKDPinXBgVpTB0O7+7VuVk7GrjGYPQ7B9VReEbS45sc1p
pXZkyH4D/UG/0vSaIDVpmjAWL1p1TxAh/zaAPBG2uPDZtGMgPtA9UfAL3EcJtskOLSV1u8lSYZFa
T3fsvTSie0vFaL8pwV8SZOh4RIj4VLYYY2FVbuM0M23T1VviJfx1Ta4Q+2PNaFGoENLuIaaKbYTD
N+d6KpQAXy5iHzgINZjDhXLZUxELnobb6tMvuYsNJFmHZ9HhiqsXLWTXtmtgLeMaeV2YmV6RDOdf
w9+iakgmIvZojcYr9dRvp6JJI07ZVGNbZsvyJTJIyRlJVGvoy9fRkeU8f4iaqDK+/MPH2DiWMpTd
ch+VN0GweO/eSgI36b9oeerp0CQrQXzlLMPr0+OPztWruLwBd5zs54DuresWOMYKsWE7n6f7T6f1
uLqjDoi8bSkWcTkhhsD7YUXm4AGKJReYQNXGPT74zzHD3y6M85ZsAtV1u8FI4aoE5yysq+EMnJaB
kGTAHWfRypNrdTo81rpyzl8/MCy61zJgEDn8RJHQdRN2wFhumRxhYn0iKSz7QHkzdmmJHqrhPBal
xCp9D7gHHhhG/UdzKpFH4sZ8n8TqCAAzARGWi8B8IJ2qU5WocwQS2KmFyGFJZ+ZK2jcgguRggK/j
HuEAuC7t6nTFmThRg54OFVz8tgriNGQDdsUgFn6FZbZCFIx8meUeI1zDWK64YI0XwUlcPOI/TIGz
NqDm70GErxwgdhz0dix5UXmPNAL+7MHN2jbfw7qSkZnnydVs7CoTNy3fOyJu/ut3vynAukuezaHJ
V+A0Djsfy5f6petFe1osf9t1SGFRX31WoH43Bx6fcxcVOMxHRweF0NJCdpNWQ4jbMJF8tY0r1jHC
yJrDM6n/V/baeg0ucR7guwvqlP8R+PY+CnihiVHSK30JNSxyfcR3JLjSCq6edthFvbKdybsO0N8W
zqb4hPhamoDC775M9SG3bhx27pegP9AnTITcJNCWToCSp3m0HP5JLdB7Z5zpopo2xjM2dpm2RVWU
eSrXe75z8aIOmMBCXCHvKHZxXEG6SmBnWf4qN8BlCPa1Th6gQr6Xy8/tvQ3lBEBN7deNgcLwxDUb
AfIJ9y1Im7BTeO+9jsV3WM079eBNenXx07dLi/yeT2X/MZWjOoO9aryC9pgvZi8cWW3KHC286XbB
RvoB1goh33qpN9frzUdla3h4kxgZ1vxjlTwwfZh0uTeCyDH1t4+ypHYIudGBxS3QO+zYCsFPNCN4
PYHRRfU2JIT3I84ZMLgauhfuLywghhVQFcG3KLukuDFmaznuP0Gltn7mx7d9fIXtSqXLBFsteLNb
kyWCeTVEK/SN/Iq/Q80FfVTaalUZxgRXoKNHDN6uX6I2y/ShrmEm1gO/yKovlkYL+EP01ueJhFV3
+Y6T3dr1x9g0p6zpfngDOTjYSeEcLFbTu5QgRlqz5QusUlHdVh9iB6QBpxgLcLZEBPk3KbGyY8Sm
JMNXzJmOmMhbVJm/EknwRwshItXzGeU6x6JrDc1DEGuhAZQ4XYlVmFvacez40KGODDs619tO9NXF
m4dru8dslc6gnCWCPZTJ4e74u9d7NteSvipEEXZLI0XYS4xH0mbUwnBzgsnXEOI9CmLvVhEQewuZ
imPfl/sk4nNK4xt305m+D2Yp+qYQggq2UDZAFuAObzrKp/DI3urOLHoE8A/+tleyfGUbqiGMBfD1
HgOTWWNutTqEXhWGk7UeLPHDKH8iG6yy7Rs597fpr7SmvBrFNY51wksKaclixq1PsYhNwDr1ZF1n
90XNpnwHE4PiTkLeKN6jq08L4UIokQLI0AgklRZnleg3o7fjm6ffZx2bWt0ARkCTWZoEzwjS+zys
wwXmroE/XZYHdbxg/x0M/e2vuYxdY5NmDtW7OlqH2rzujlUhbXtelW+p2fkLHUs8oVbYevtGYCPi
YRpJ1n2Mghgg4WZ1pc+NZddKL+DWEFBSjdClY8UeCZaDpNDj/Sq+WiwIsU4ypABOUns+WBf21Wn/
bC6wdXInohtVOSgTRDnbVSX+u2cIjL8Je2BknEj8ILUYuS8edFlM/uovWMvHz4oOyWiiCKhH7/Fc
A7mB3WCIu4CucF3t+WdcO6ygu5+7xRhNbPNZdYvhmIDLoeT2n18WCOLCGsovFeCE7FKyRXFkAPY7
vw7AW09CgCGLEikSYheca1GZg3R7ucggUJecdThkigPP9Q0qhIdkZUELTcJ6r1Cx6n8t+ajEnUca
WrqZ5SumUhM6Nijre2yABJ7WRK2XpycNh4aUGtylgrLDn3B0rP4r6lFXkQRRezqnoja+JDKIOs2j
ObzPXALRJlXWY65ZIyYnRcAJA+3igEsJai0DIJjKjDH3gtiweq6rjLJRVErTaQKh6U0p/oZKXiy6
jth7mqhc1vNfE4pxQUOYucIXsmHP+p9d+Jctpk0FptKEkzFAqlktXNqwfpsbxFeeUyFsBAp8ebRe
VNT7phQ6TimEBimrOoG+soA9mDw4oPanCpV8wqX1VhaduTOarH7TIDH8lf1ZODQLRJbqRaFT1G06
fUd32niz9CMBmSCsKppDCgpG196EQSegAMNu1bKibtPC+67L5SbE8u5ODi1c+HiLmdbU4qfsgrG+
fUPe9vnRneVXTDOp1xO7ufKtPYdjFtXwxrdX6AaO0Y1a2njoFWsKA2v0nPgRP4yTRdKTfK00Md8J
VirCq/5Ibiryvvi1jZORPg5Cq2r4mgAe2jG130hToLU/c8cTmcyzsoKiOuNPKVMj0BX9X7vuKIfZ
6K6uaRhrG50Zt5ZwPSKrcF67eTa+CPdBYiVfHISfhnnEOPdi0scUn6lWZFXh0OKRAcKKEGiqDNoM
d2IQKHvp+xlG982PH+0hmnmouvGaDZT34Lv7hjrSyTDeMPW1Sff1CGUxsjAJtUkYHT8jsJXZLfUJ
XCOf4pXwI9aVoIweSiqUKjpZjNI1SLXPvKtdm8KljN7hYP66QLFZI46Ko7iv6umfPVARtEXSPYG8
5ygLH6pIJQUEtetKz3IZsScIdsh2piRnzAgo2xVuRobdC3zTz6wofziLFNUiRlm5Sy4xftQXLRSd
8YODOtOsInlNntSOa6t8/GPallz7/rN5nQU8YZkQ4N8bfWBYCHIjiiXOObmN+bRfd1g8AONGqF3q
oovbsHK1tlL/0ZDesfgZIjgvMATel9wq5pzqudMqA85lAhzS9HRFcdtFeJAUyKUBnZE18SRT481z
tFXFlzYwS3GrOAeHJldcwGy6LtFfKb3DfK3aL0VS/iHaNY+V2K3jHYR+SwezYhwNUuITrLIdE+rc
DhzgqC3MWDvbBu9CgpxG4ZeAjmW+W9pdOQew+2HMQuXVgCLg25M9cjeelx+UGwlOLyPgyWHeEB96
rQxfh8gbqHBC5B3uIIJqQYb+dFaKVuEyIXeT5hk0DonqEW5vHTXbm6dQPG7ICPo6K5yOFRv/VnRA
3enLU+zgU/ENhvOX4qEmXhCoYoNDEo+AA0WeRrhcpPO9V/aSLL8oZh1G9oCX8yDJ1UvIy/ilGl5v
SvodacIa76dmywzMQRrJjAkPdoMWqe9vwda7dV75fx3WGUs50sCcHGzRSK40ARodra7Fne7Ie6Fv
+7m34KBnjbYdgCXN/E0LtbexnWYtdjXmI6A0uaOnqwnw+VjKtnTIdLv772xn4RZ9KY4gYtUPt+2l
q7eTh77YewebnTEC/z6FRN5K145lAKzROQMT2FKiYKdAhqlFn2QRT1NWixac5aQ5ruG8DXOWWFAz
ZCyOtYkR5aO2Q6Uwst96EgXqOeKXeffaivTxjsEQx18W73j6+24tBkXB/NNQxEjrGPh0NnBgVZfO
AuU3KD8wEBZv/z80gIJNVjDznFA3/Zcln337Eh473xc9KYNv+E7KWJTKWwFII5kvIYg9dprWX6YZ
p54nsftKyWp3fMNJZlJG3dCtApMUQsA5s1I7EfHHgL/52uLSLgT4U8A969fNBOZi7SDSbn//s7bo
TnlQ6RyFv/s5eE1GeeT60VsMUHlhMjMaQVXt3WiKpJdG3583+kDDqfLd7FkQpAtqXRd2qBeq2QWy
KbFExEnu4CfErNjN6Z+9DXHp9MjNRgvKomQ1rVvYU9MmIe7G/ge9qRB4fkOyHbM69QQJL3zq0LFr
K2kJMWss1dA3/BBiAe/dYF4lWDlDJM+VQKIsiIOCkOEL+EQ2Zc0yHWe/IXknA5VZ82wGKvkMrnLK
CzZHeiZcpwwAGZv2u1x85mCseuom3B47fjsHYk5JW17vMqjNnYq2n7RsCTxppHS2ScIApwOJSiwg
5HUhp+oAKS3cdv0niw57tQrZDPttkaDo/Pcr3wef0VVluk0mmnpYji6ERiTAwQFv/bx8iOs2NU1q
0A/GyTqAvlcOnC/vrdZtCzLHe36/+wSYVvVBUTjKCUzZj4c8gvRxipZGcRLRAg1Dul9R1HmvpQWZ
IBSthr2atnK3u30OJU5u08v4nkzKXlwMWs4bAxr+Y5yrGe8L2hKz0ImlWkIckIrRHV1leL40VvqH
Nhw13GqXzEIV4PVPCjcgDu7oRfB8ACftR1bavkPTQK7A77ysRc3SKU5H99xFSzCeMPpiuBWl1ozL
QTvUFfFXWgH+oIG6nXRfm9wVbmJYmb6k15X7rvnjgU6ClIflAoAdrgeQVL5O9a+S/gX79JuqwWPj
V9kbXSy/bAlcKyf4BdnSACf5Twi/jcVVtmSiEn1jFBILboqX6dWsHwrIp1rDXlCcVPWjbbLWaZMF
653U34RCnqBP5eAmDzYrIeKsuSEEDzDmKY+3qmezOAXs6G7DyQdgSFVkG9DvYMsyKbDMYvTXS361
eeYdUjXjR0NCIqG8kpGto6gwMajOMeFh0yMDz+tMVak4HXyqcd2gzS62RyhcnXDAxXtkc16F0DBO
+ndbcfdtq03HTISIxbW9agLURJRFVqaBwKg3RGTvvYnNoZHGjzapLwLsFsc2NFl9EaQJT2IAZL5M
GwE145ynS0/MCPz/T4d7/MgicJ3NvVI6/SF+y274+AY7/27/STTTjbCTaAG9vydguJdo6eyAyQn3
yTUZB7wgfajqKgZ2BXS1naAnAMjoGMlanE1RcsYPGRPSMNVkYgIB8SQsS4MPzvz7R9XauyIoiPm7
xMMfgTFNFbEPjDSN4/RzlSexnL01WNgrj6p65V5qfGyIOMNPf2lHrI6nu0HlzvnB4gq+ZqOx66RY
KNk9W1TQb+c2rhIhYDs628T9JoqxIPoXgj5UGnClM5TtTnlRNNZ2Ofa3zgv9SLW1dhasOMK6bLes
Ea69iueiOMC0wut4iEY8XtTFuLUDXuYzTZcbjS8zGtSymtKuBfRmuWjaajuLfZZSIrlPYVA/tAOT
65I5GKpWUeRmuf9pM9YzeMtc8F7K13imO1u3FZOjBToYdSk1lyo00CJwbNCilAwSf/zmaOkk3NSO
bSesPD+UAYoidkA0YHR51znzWDuNUi/ADWb0t94lr8FGWlLVnhlNhKyX7EE34SpYW90M37AyKFxm
XrQ6yY/xr1hSnuoT2wXT9wMO3x6vjZtE2rrIsHvKfMKX9DrnxIR/StKMSpv4/j04eLo3pd2lEGW4
qXs9JYkzuh5UegMLtSLbERPeD09iTNF70CzIiOoYfxRoEZbqns9Z+99CCOYLM8Lc87b7AUdSDag4
c/iO/kF4ehO357xtvLN9l00QtUoppBI0Icy7xh90V1xMrl6vJKNDneiWwaA6l/rwtXLjWcx2ZsZa
ckYRJLAX/3esecslDJSzFcySrG9wL5yaxdJtlEZVnRxP2deTesCp7Di/5rLFjPNOY80vUZ29tUbh
IFyyqDlXFmmCf7s6jlurnOq4vVdc2H826kcCGyKhh8K5c3NNptWdpqnpdXmoXQDmakO/6rGn63u4
rYJw9apUlJrbXZEogNi+sO4nlQEBKtWHTTJ8CuyiLhDZlZ7EcG1+PGJJGrdgyk9Ofg5x+PMYEItE
5v3AAqzlVCwVsBZ/fjKaBY5XbRR44nUPOSpGOA98R+EAyHErELPRgJuOUG/YPVlbq8QdUdVTzOkx
VyHSe/hEa3lXiTDaJBAYcOKVEQYzl+MEv9cHb2XhNhMJG40/pIbbJPbaruzaAJxqZzZn0um7uoYx
d+Jdlh9kDsovq3P9S2jG3Ja5DVnqnglv8Y0vL1ycroSS7ubOT5eHqIOeOBe9MLT3zZ5ZX7l0xtE4
mm1yIykp4uAcIWKBjx7UA9+DrcIgWz1K0ujANCE7yi3mhljqxYc8LLQegkgnr48820Bws5zSJTR7
2ZGLd9UfRmWQUGMpCoOKylIC6v0d1Q6HC9yE0O48XFKfK5LgFMK6slKmwNDVokNMNiZy822tRNvj
1OrJbhNmvaUvRt9MexVaP9f4HEi3HB7MrwsXFGL2zYlqiDLvotfHwNCuEGCWc31p6hAhJYSsxtEt
pIlFy755sMNGev0Oy6DXBVYs+m4qSB2HRwhl0q6qqqLNyQGZyYzIKKdl3ZBWKUfOUi+m/+Z3eVpk
WCkxo2ILIqCYki3I4DV7GLR+bFtb12ZWwuaPo/7iwCJnwteYkXqKbiivr+JZpLp3LXllErA8qNvw
+Mm8t+KRPvXxQydgaRAW1sr2afqNe3Zy1JmhqPJgwqI0/W/Ax//ha0O7q02WG2VwfiiZ2BOXmb7i
3/W2hqWTuy1On7xPf6frd+qYPq68wztBkjSaVZMS8eJNVogw4rkkt9+Yqpz6ZGQ6VDVEx3FOg9tD
gaB2Cyng1QNuQdKk+LTX4zTz9TdYthv3yMdIaRaEoATceqLQTf1Ea/Z1Lkhwvur2BC5QzICe0V2E
mhKFc2W9b1HYT43t5bcX2DvBkMs4kYAMcmGEWl0uztnYFr6hAdBU1KGSH/Fb2+Ro8l4y9p8oLSWq
3/xkMPaDBPxx/95mgp0TmNJEglazEC4OCgQJ3N/mWK5nHS0ZQh2mOHOseMW54s+6RtRyH3w4e5Li
6vQTiE2/dAHp5eD//PWdNah47JEwXrz5FjCZsdR4EPniUOtjwieeo7SGGVbUUHPi8/GeQoG4+yf6
yzYpFX5p2zz1BnDBYPhRvo/z/O67WQg7xUL+Dd/V0N04PosmQO1SMzF0ixc0NkYLlyEyWKwaxrQf
ijh5Gz4SaXDj3YtJMv6+2QMwQZku1e/bFB/inzVSDtA9sO8hFlYAMcREstHbcJ+CaoW5cQgeyb84
rmfVld0icUxImh451llr5vIfCksBHku/k9wdxlSjV176sztjoAPWmTcsI7ByRn7JUzDy77QbKfyf
5cnMiYozNbFun/0PaNJWUr0hx7YP3aBmR9QW7Or6wFbNwxH+2Ig3vaG3YEpnftv/i9BdWTdVe6rW
OmxmKxui/Xfpqj0BgJPl//kWeGAjw8lzEBDSKJUgcJchHTFnuPQxq6Xvxd1Iad5DxazRYEgMh3pl
pVaknFFfQmd3EsO0Ze5FxHL9J7ouJFlKp0WtBj9k6ypFvJxhvy5IccjsRq/RJkAHdpDkPyZfTjv4
v6shHovIYPQVEQXe+rr86K839LjlEwXTWKgSdulmKEthyh8+f10X7q0/IbjdlRjEcaUok2PkwqRN
aeQWD+/GcdHwAV6z9KJ1Y0+E/21B549471zBaojYyF/6md0kaPWPFQdI/8kL42FUTVm6EpA8VK5q
YlQ98xJkxDGWYRrCG1zTLK8zCtzzxtSFgecQDO9kcC4+Nv1zLWBmgIV/aaeAbUeANgRN8IG84XgO
4oW7cvjsGTs9nGaSy6JDkOPwbilMLXVSdTDXB5j7Lb/2x5+6h6wcZUd/ZL6W5UE+5W/5FiRbNU2C
lW6HQlGlp1oHaeDndRl7RBPqgC0H6s/EQWJEW0yG20gTzrROy82yM+uSjwbhj1wRCsoavNUqfBX5
TdWpXXZrtCtMXW7BnXBUd3Jp2Z5D+fYS9+G+ACs6yTXSnguOB5F+2KUHCKTZRzvl0cIlPKwZ03H6
UCRrX0GQ3S0o+UAy7Whm5FsVWsibZxC7rpdCcH4PGRFx0pmtNSeGWGdbbM9yEn5retnAn+xyOcEg
cbAycwyK8t6IZz9pcdJim9ACUdhSoXBSGTRkfmbM8pndJO5FYAggbkwr/OTDR8dxsIhl8zYqSbL5
4ELDmRaw/NJjCnvz8z3eG9hOZ6hD+QCGwqMDxq9d8A1exLD0wBaQNGq8iK9obLepcWqmKyXq9Qrq
iqv6lWyRuLpuZHKPKLDTkzEqxTS6E2laG7GWa7wG/5tEgwr650MWl5ny44RQ0CLaJNsw6K2hYl4q
nj54EXUNnkx05kieDb75mDlJz4FaHBTclKygQL596gxOU1n0GhZmOOeTd9gYSFrial1//LGWCsJT
gvB6hJkGx6xHA0TXm2z8ZxeqS6KUGSVqptIPepM/97WKj0BVWIp6HlksQRXhjtzG+y1nEZ5ayGty
RhFf7zh1TxUwIoi8mDKnCgTMt1hBKG6cs3CWTaqxSTggZXwX9n3otPgbYKh8WHsNHKAKcfyMK/pn
5VB59WZyGq7gWPQj6/MdV9dUvvdci38uYcGAQCMlkXkT3HVcrJIPiYVwieoi7LgkFrp5CV4suVKX
jYqPGzup54hi2IKGgcOo+CL5z7FGJRLwmqMvQsmNUQTSFg4oUYlGOlemnxJcmXXC1BDurtiiu/SE
a5hqi1qqRumrQP9UEeTjbre4zCLzWH9afkdzkSGY7It6V99RkY9uJSgQIAXOz5d2/qux89U206nt
wImCbYAuR0i7xWMe6D6NM7itbdEABu3K/TZqnnIQcVEEhYcuzmZZVwKPDjmc7qf20jiYrax/b9QC
ebP/zhsU4AJR4ImEzQnj52J5bsqTkvFdS3nku8e0+gBdc8yji7yyvsFuZ32t5J/OUl+G0N5do6Ja
zP+zjPe7Ih73KvkgpddIBD+zBmBLk1uOXNXcs1GERw4ErUSWPWEnaz6YuIaFQCRgU2rVix9D/Sd/
5FogsxylzGdumr5Jz6WzKqUJ7vpvwzpCTYRKkCTlKXgu1EHWHQ0byG8H1aLx3wgtdKPqj9t1nI/j
tbD7weAe0Kq87Se1OVGBNQijg0wNUKML43Z8go10XithXfXnp5afDzhucLjbDONXa6JcmbVhmwDh
M23pYiT+B9cu48X1pKRDuNssq9E/plAfRFEGRyPfjoVuFeoRLneCabpo5dcLWLBf+yv7G6YG9jw6
8d8pUFxY+ggXRRUWa+Wf7y49EbT2DqssR6qc2pb2QPRB2mVtlvuWEMS+NxU6lDS5/ihlsRHpvt87
6VfW5NJPXtKtHIBa1HqYAdeY0lfC6vW0ExeWbYqSb8uvYiL4EU75fKPxFhcuUEXu3LUcTPUApk0h
v3zQFoIy3lE28b077m6ibwTppUZJNKcddIALYib7aSzDatfN6V+BwdI0WBfR+NZJNYLT0hDPP7+8
/EB95TddFkykWF7Ms4ygnJnLWdg5CEmEvV1S8xycgEwMUKweDCzxxII04kqN/LYiUW1ZLi+E4IKc
M8BZeVCQ9uXHZSdr/5w+0koOV5BGPJAuo9kryGTaCreg8j29ZG33F8OAV1zmegreJ4WQbP1SO3ux
LVvjLpiX39wHB8RaZminrUsf5pm9Iz0yLuGvaRlFXzBdc6xLtX+ujd3dACdTbmXxXWa1cSYymH+T
BfvBzHPq2RJ+KOgfXUCVb2mLYAOSQEKqzKoI1hc7zF4vmO6VhPamB3aElqPVLZXx7MOGpPcUQ1tl
4rB5bztCwPMrbgMX0Yyd7uFz8BSbVpECR5EFoVXms44OC6185P4l+qE0mYUGHsHcuc/rt34G4DAf
h82FXa4RNoQhxfcM00MOPk4bKGOD0oovZ7eeun6oZaZVDhADR4IkeRM5CwMFFaTBKS+Nux780F2w
GYBIpUTGDtG3M9BkUfaywbwgl/aKmwbi+gX6q+ewlgCX6fv1NJPnQNhE5NhevQ9DXwtRqmMSaUFu
1RwEusJ3921aHKBCrBkb1mbBdlp6IWMQAf12FflkKQS9RH4F9wwTZUldxgwDIb6B19ZfzGd06dl2
e3sQMG6Rp7g1XAXxSxns/V+QZ5LUs2hbsBoM5aEiwWmjeZ36jDqMXBxZi43Io0jMzNwY6bFrPQro
hPr5QZhEhpOodUfAhbcKMd5LmELNq1zCU/fVJKABuYy80nCpAhG5kHe36eOulYxaivzd4IHTrvcK
4LjOH/LYNTWj+hzKgEfL5ImS84XUx5R7r4on6Ltm15mCDuXROjqzvDapqR4CdOiWCGjFHct7SpH9
Z0wd1w79YTWi78s7Z7zBBuq0ge++T9uI9A9LbimLinlrBh9nIUC+vsReX1Q7L89qJtjeCbpbk09y
JVJKTbw5xxnz3avVjrfPxH+bbl79uD2fOiqSZwwGwOazMwtqYeMIMkKojRWCNmb5OfDVDvakHsyA
/Onn6bLbMfHfGktRKhB2aEg8OPhyzf2REDCblTOfOLYRA01oQPnu1X5OpjBDjh8+OHrW6YajV1rG
7U71RFlPN9BpVXaZspnOxQFcbAlNRisegneQm8sivIOcaqlsIgR6wYh6wqbJgUpkYJxiJqUmPkd2
tWPd2eCz1dHJ/CZNlabZGf6aNJ40ov+mOGpZwiELYlSA2J9KBA+rirPXAvSdRybxTOjTms/iaYr9
u5ww70ENLQ65HCrAdgNiRmzmb8J0IweA2x2wXrUvLW++qOoQm7tq9uebZSDju1rOj1x/YFqHQbL6
eXJeNnlKAY9OVbP/wgK5mDi6wauq/K2oF24Waj4iPlkCzB1XaeQXGg1v2ZpfpViL/hEqaVqpyMCN
NR/tIE/RZRZlNw/nKZY9N+FmpG+M+IBmnP/0O+AKYPdZoPcP6RGf88gby1F3bofdPDyg5Usm2zvx
Lgu3GlisRYGRNtdn8VbkscjEZ/VQMGHrOQm2VapQkTwqmWNN/wC+tz8y2yfNVpHlvivq0KOfXo1l
846CiLPW3IozobsW9zWiIDbeGSJokizYETHkfssAy56F6dCY3IRkpl0HOiyLl+LtXvDzG5L+GVNT
E3uf6ij+X5+8sA+dH42DPXVpyS0COMWI9fV3yghoC3nb3VC685Z5X4I7p/7IY6crUq4Vf+LDWwAl
QLpIgz77IgQ3s/DIN3hk6IOm+JhxLkzJrBfdZudHpUpBbLe25jmGPCXevgjS10nFaVHLI9EYqLcy
Ids75rNXiJ88YJlOK7eG0jbePvwaCgbNA3tmdTRn5GfdXiGBj2AWqZVQzRVixe7ZzCqOcVxYRiH3
b50RwkHS0BCO4g5QiK1tcYfEvP+9TRxtxeJDiqFMYQXVJS/m085U/QQXPP6jdgCUmo8DukvAuOv/
RVJGyuvCH5Erzf0tiGwsXjVcgXsS6Fb3Rkh1KF8DkGBNoeIJk5HDoUUgNCvoCM5rp020TIqKpLu5
WqU5q6L4R3YYdHFrISYNqMuRew/E6q2cD+HRguIiEeuWZDFPyZCQa0tAeMLJD3sSYMTo9u7AbTmU
Qf6laZRhYsMDGBnOj7MRXS6f497/yCrxqtJrAUiwwL8iNqhxKE7WmLTnaGbiAC4pcbAIs93jLXbH
bvaQ26i5veZ3mK5q6kAFA30vHJZ4tezsZvw9ydqaPMpCbYk3uM6TdHdtBwdRPP8wSgWLANzpXYSN
h5ZEFGnVtMJNs0Fz5J692pT70jy38V330Onxsq85NEAYC6l96rsW6flLXsW7rK1ZQKOh2gjZ6MjD
hQgRGJj734HMm93w40qpjdOd6MaWqi46SbMwThNFCEnTspNx/uHfZWnRC35wetE3SNu/eGeRMmdE
HdPHj4wnacXvn4Q/mlfG5hFtNwLPlUM2YSFa6ASPiNpW7dFhMUwhFwHfPPhLBluGlElpEaXSLN9A
2Zy+nDBiiAi59ID4mUXHA7dQGG/Z+ebaj0m9tVNuHRHLWuzGYuZh4HNrfUA3nHKLjbJ9jOD/TWvL
iT5fnMDfd3nkpjqY1MNPrakGADbWqmvq1PJf7lSJsqpo2lqm0YA3jg/8gouaa2gYVsNAqVYeQQvk
vwq3yfm6VU+i9CjoyY27mmxJkbGNGY9RwaXp7IDs+BjkmYV0po8xK7mcXyq646zpEqpqK6HuxpaH
s/sSx7SUoX+LvGkb9g/Klf/OT3faAoKc127jhGdcC8CtEOUmrxKwX6ey/2VzfLXneymwxUE8EW7D
XGImqVxeZZX/4zNIrCSpgccBEluJzS2JH1teK1RjPOdX6CmOG7/Tq9zMJ+LLGjB82FUQbq8v/ZsT
ZKq6awshYrcq70p7raGuQu4r5FHvsuL9uAGmFIP7hnG4HqNim8ga+RpGYzERShRf/kM2PB/hRbq3
a17hQ8oXX6hxF5XQhP4EQf8tsBYQO059j0yB8NHqG8KVaWWaTYvK3zecFDQf8SWHP9K/v+vbUtso
CF8omSU9Hxnj7Wo0gHUTytsDMRIcTzmKN6zMGM/8/qZpcnOs33wSMXA3E+GGnL+GV+6kxu+hH/u7
+HbQ86NCvWpebPt937JqHqE68624f3yH3cs6gI79jaPJmNYl/Z/ZhLqIFmSv3ysSdsURhMbz3VKC
FqCfLXx0S0A/K7ILu+kKN+8serw5EOY42giBf4asZtejUPMmjskR2JpIMzCDi7sHkS89vdjxEsss
PnNIC1tJd7jcxSswdQT84ugSfX04KrWdyeidkuBgC8EJa9Y4aTj/DE8dF8tZ/a88gw4Zvomlps6V
ZD3/E5lxSRoDVsxAxSjENHjboKRvzx2MkfwraO9W8hY+dR7xQpK9BRyUDk7Pg/qNealrZ/cQx7Kl
2gNbqEzXbwkagKN3KqaH8Jv6PNwBY1+QHRvJo2x66JdIP5eoAMthTLMAAMWPFhFg5owIv6RJQjn7
bA89HjojlSXqzh+R3H3TEmZxipoNH4zHaIRYIDDeTIqfwZ/4DEGT9vxG0CRrcQMJHjZf2tDPxDSM
f0KsqVm9GhGCCSnd18HYWVvQoCB7Dm8/1pc6bv1p/VIW8zIM360sjruUVfoSd5PU0QvcjVx/ZMU1
bRZD0oEu25x0v6/uiIX5SbYl91yP1RsJfwJoEJOCHShAX0gPNminyldoj/o8GjprOyIwRv71K14J
vOoPuOGgWmpgmSnADTrsAfpAqzFvBRd/BYxJTbp32xCRDzXBl8uYGyLryQeSAL5OwarLascmpxbN
VjiLGPlb3Fg3DnsZlfEopCbZ1Lf1giH89FuhdNGaMtuRLFplPp+l878TkGS5C23YhZBe7TjjqAG5
fep6IkBiTwkW+B/D2WTjaBNvw1KsTVdkqXMgzLtHYN6Rf4tiSQdVo2Up9GydtR5AV3oIwzx6N5r5
yGDMi2ElJdrvM+zqXHDEs/cT8+S4yyBlgckUbijPugTU7nDHQySSaJ6ef9FmNiXpQDR2eRviclrE
OgTApcGS+0SCW6ASglwAV1ZHuhMaLXLMC/MXTlPlglJyzdbTAPbSJXDP/1DiqQqaR5TKoOdjnp1N
j/Mn/oyMW79h5E3geYRMqWOkXElu9Ny+B7sf7IVaSlhg5VtdeXNOCWd0Dpi1fdp7ZhN5rX2Y9I1D
f7TD0QT3Zu6Ri4aZl+H2Iv5qnF+3HYu1UYRPYDAe4PsPGHQvQiNI55bAbeH5VMAzKZYIe/KpxwSC
w3LSFtSHSXRRU1LlCCYv5DLEdb50g+N21xyi82ulIiTE2ilL4pXp2uyNVYXFLojw5nMRhxfGcYOl
pJnrw31vHX4DsvlNPYSlc0qXvMrp03EjddHuKITCCWCCMfpSFb8pX/YvO/3JWJYCNESqrKPNzlmi
q8OOZ5BeFbtZrp9VpsCSRBj/zY9d1JBBt5sli4NHfODicGlkN47Or4uM3Cv1lOuVhP/iOFjOl1Pk
Ln9bxumS5U6qv1HkPQV42QcXGj+sUgqAZYAExR6L+MmMV79xw4/c47KYsV/aL59yuvKga8hOskYm
xklY4q50QEKG8guAxfXEgvL0th7DtvrVD9awbewUoV6DgMyFK0JBIlfzhYdXyCJqJQnFt+BstyvK
DGkdmDxpSuDP8zd6JFOI4wY0U11kjBLBE8FFMLrByK/0fmkw8SVgH4IlJMp8l9G6l4alo1jDdOQz
0LMnkI7O2njs2MGnqVTbMA8JKaZESH0K+OL3viCxFjPRPptqq+XLLHv+15p3pp0f8/5sIV6AHYUE
vXivb62XzuC9ywVuZe65QTQ1OLPo36r/t5mwGxobt0icA+lORV0lkgPuCBUOvIAbxRYgPmnYKsPj
LL1MEHewjeEwrGED3oSA99X2F7wo8pJGXxzvjmLtvDFSBTcZXf1AFi4U6eSErfi6ObUEgKqSxIza
asF3NudH/XDgQcASo6ztoy8btLjvax47nlTlfWQwiDpSnDIspGIEeUSQVTX4Xl4wpu4kZFSkbZ8O
e350aplhycPYDZqN0bgIwm8pwC5YOKV8iosXoupnoBJ8FTDgyk+n/lzzxUD/VvstZ4PlUzQDjEyL
zZYMiFbVfvCO5c0DjOGRnAOSDu8BMvOrWhV5a3WgnVJqe69jOnekfj5vexI2SQn6xt6m32A/glfH
QSSu0BJu/kWlkpyjL8qHCBuvdlTp++gJS02TfiA0BaEeuM8IRzkQ1D3nUfJ7bPrCQ6d5xlnSmnQd
xMOQnUKVyFclGmpMZWh9C25mXIfTuREEeO6L9pF1u8JQtO0GFSC5R9LbO0wBwSeP0LyMUYSwTBfi
QaLk08ZNog1bRtj74KqgboiJusc7l98fQgcjZdomdUY+9ekIBRtYMRXxxJ5V8ZM4uyLh5wu+g0Ah
AdUmepPsHx/AZ3pk3eHiDNn5R4ZS8XMmVDmPuQN06KdPGCdHUo2/toq9qc3XWjsEM4sdDexqwCZ2
XvqEI4de5lz1f6bqVzlGMEeQ5LV7owltJa8WQXJVumckaqzh/iocxNXc4b+qACsTL1GQbYJpsi0b
OK/3YQULRjJOuDTQuhDNHB5u+V8uYEJUMzjdqWRtMLecc9JkuvQ3fVUGXwn1nXGNE6p2mOHC1rvy
2ip6AZnDN9t0lT1w/re96cmZNxFnTnRE2MUQAqEk0bhIVI28xbha9I2xAsezZJUJFQqsSF+Ql3Wc
5C/xImiRoQ8FRhkJgHpknZN9EK7FOtyjAW95Zs0Q2DvdZgEECO6gbsctHdRbxgzqrMyMS8i0fNDo
BiN0PRr0QzNGQ1J4b+fgfyEPZJc940eXFo5toszkb4suvEBEPEaO0FYTH0/b1NLolPysdNYv3p2Y
cA9M5m4aARDnnAwudmkEP9aTgodnopCBi0AnvxhG93y9q4fvVPvW/LhxXrTi3Tjiqk71SywWYxhf
6jlxPPwGshdKo67v65Yl+onfwbIB7/IruA8xLSaSYNyWuPHByGsujLYbO1otm4rLoI4T2bILcOWU
icqGxGeGn0PCVRhYq59N30zCH9aRhbj38UGsVipjnT0vlAcfplck5YyhfZ96GlCArThoVbh4DwqI
r5rWlfDadsYzaGJUDKwdqgJmtbKpcM49I9Ho2AoxhbdXxc1+jwlARPKmhOOchIEmoue8zw6NIm5d
3IXnoFCU63iJlQ45t2HDyb1NeAGq7nN3AcjBOHQgsumc78xvqR4jjZzPR3cEeIYOskKUBSXnisQu
otOMvc2yqilURB/xnUFGRwPRysuy5IPEcUU91ON6PuzEDrb+cmdGQaepf7G8qTqWj61VQsAevU4Z
9Hvp1XWOekGzj3wJ9aIOFkn/WxEDa81kVMm9S207juacz8MjeQ0G5kxnoM22ksHzRxVJYzT4N/FU
OSiXeiZMQ8OQNWSZ2xQzzfcRSYMbF6jWdcajbyb5AZwpPoBVBgu5SY1sWIBqyBD0OQUoDDzPnF9c
iR4+Y3yBDEoRgN6S1+O9J/VLqh0h4mTS9O0vXlNqUNNmZbJC2QM0J4RozT6ZMdsr0lyQHlA4wXJD
aX6HNgfycxPEDLx0qlAADmaPkA3cPS0UydjBU1PhsJJv4Ei7eIHqComi8z/nHKNclCy/R123VKP/
uXaW9y+id/0bmGXjy/W6hc/7/GeSRsfCpJIVnmVW1M2c/GFom2GEooWu+SxsN1JEg8+M7VI/6ESt
KezPoPPqqfJMOEeV98OlW8oZmYX1nSbTr7xoIyOUaQsg3L6JHNgg754GZLAIigjTfTjQqio4A7Hz
mGXhlZq6E/Ba6mR4kjZFhW4bmAEW4S/YsOa72MvXhXN3ektpy464q4zgXdCfbRGhHfaK7qBy12vX
t5aBJRUkiCS6e+lenDkw0avK1ZW5Be4whY5yiJ/rmIhui3A/PMZvZf4gtjlYVrrb7R9KWox1PBxO
x746obm5hPVdwH6tdDaUr3jdMk0x/hR0PI/BKWMhmv1vlC4N6tjz+TgkdT0swDSHjA1SaStzF9bL
7bh6fKDT3eXxNPJEo6Bv+Ru5el540tzz0+KiTUqkvn9lPKXpBmjTSxzETT2+KDQT9CDUwWbOdar4
snBTcXC/FX71KkuB9GmAgkY7oP/iGJZL6RZPe9ZcZueZ2ziX5e7W+7mm0YJuf4K8QZ63lZOTnvpB
8zpKcVx8eQ5T9CZVo6R2AIGbkmrJ0KIBhvtrkkbDEzUqKEddNO9aZ4tWREnj9awLQFIRUpBohdIo
+ivVdgE3kwJJgMaxs3VJkQcVK95CpolGhfaz9sFhV5jeHhZdyb0pmbNS7a9V47bngqkKT1xV29/1
WxSRm1nTAQFCg2qqdjCB+ii3QH+KQltjVD6XWT3Q9VNK0Nk2zGi95+ERDdrz7lsrXr7s3GJCxp31
/szm4GkrPmBqDDKHRZ5qRerVY3AnsgsKjZuoGNhnZl1dTA6O8b1sTLu6RU+Ch3cP53wZFD4HeHzz
cdbH4y//cvCfhwMkYLUlTn3TIA8MPe+BA1EGPW37tRKhQXnyom1Agck7zZomBbhc/vyQ8hRpjE6q
Tw2zTwMzqD5B9RK0lXmmMC6nzco59bWLBZ3hIcNmQlFbJza/KgwF3HF0+oj3iERVUohjAazDJBFj
nthS8sH/GtjYkO5FsNxnbIrEkezZt8kxv5eb7zV3dew2X6dvm8QkFu+eJFIJWACt9i+wc9vXlyFQ
MY+WsJqF4SHczcIS/V4nP4mrlGksgRQRy32wNbOqvm6xAwDdTEoKr4j3IRRlb4MnmJ0AM6JxGvri
kqck4Bo/yij8F7IFOJL8xjBcQ9oxhmRB0d0vVQtNd8IbAYHpXGnH4ZWUj3NTEzMZ9sO4OaWWiFOv
FecjZpw3ne8EZA+t5EoNOLLbrj/vssAKbGGBTmFTz6IjR5y+p86lK7TrvapJBhkTChkKa30f86Lr
9xHjB+OeCyGHZ1x+9lwBiwLH+S5l4CMrfdqO4znnnVMskOorHfurVBHAoSP6cxbdYRJCBQ7IFcdy
kGHTj9xsBPnE36bqFFoD1qSJo55zvdf+Ff1J5vaKIQ2UI5xEThibhlpopNtyNn1KvsQ/Y4YbuyYX
p99a97vpp8tpgEY1YpeVHnuXxhiPKu8mHt5KifXEqRFuAwOZEXWUU00/WcJkheK8o1CECiWvD2Hu
9Rz34/dIBV+Y9Gt2+2dGw7qVRNrOXBD78uWHF1p2N0yemuk1XkEMS9wjh4E+osUz7LaNClGTfSrH
zVOC+AkWbMn1H02zQEopRJEwIHz/4zB11Lzkjt9N4XdHZAXySKwOC53I4cFFeyOeuMWfyY4v9vD9
JnmjTEVA98BkCGDntTtZdweb7z5jLE1WVWCFw0Zs8FTlWmFzr0tGPdy3Z64Hm1j2hj0c4ShtQ4Ng
QmnHezBSgxhZo+s4uyOAY62jI46SW0uUPWEE/pSJ5HsNpF2ZPz+Mzw8e1Q4wY8QzWEEGcazAm8I7
THhipW4+jaASoVZCNJRtGVS91du+EnAQ6Atl+rUXRvREt6jfSu4OFA1coibjUV1TkQsH/2ik0txJ
wIecosF2ujYXzeMyUchWjanwYO7b6/uG5MIqr5RkoQ+SjAZPGcThRUMYkLrFWd6ONnK8aHZPM5NW
5oD5krqRVVqM0T3yG3tnSUFxTyoZQmJEWWvCeAqPsiGwQKoxmIlTtpl8AVRtI8xcdQIBhvQRjB/z
GH0TIX/ABHt/6O3TanniDX6r/QA4e0bBPlxPaCWIFm+73eKYpLB2BA3p5xeT90d/8l3OYBrVTRmu
TNOeznyEo4IZf4LR7DpCIiA7EcX8C9S6UPejihc7dP0/XNytNgVcKZ+JNUH7u+PK67OHurgdusv5
6bHFy11unY9pXAhJLnogUmMw4Uv7Oi7wFKSzVgU4/d4U2RLSy82anSpeB/SRABR6F9VtRICMyJJ3
LSiBGNZU6Tnu0IdHMtHOC86L6Xv6UYr9zrg6nBryY+aFYktTpBqUMIRVeHuVbLgYKwZ32BUiN/1c
KXNLSieRuLfUTZdH/DGdTCTGUeo+CRTgTL91iCZtN9VH//IErw28gDwu3VKfnZsGKMwFcHKPRqJO
8pA5fbiVALhoJpOWyXY2Uv/kNeB4hA/OXuiYjFGNpHuXkxBY8eukyzkkKnk6iGEi2YrzqxFI3VcC
cuyZzCOA3mBWL3qaUxlQGMia2sZ5o6LirMXVXq/Xe/AuXQ3HWcZggXFRdyO8cndhMt8u+LkI2jmz
pgnq7aOervZfc0wNEotiSX7SWRNc90UFcOiUWJnJ3vhykPVhqfYVzAZP2lQZ3GNzZnRpnSeeQV8q
zevzg898Gd5iaxHAQd64oJvWhUFnNGZ7yNYPY8rMBn20KN9dKsf6xvhJKID8UH0NUw/dnGWXZ/hX
mcgvCBJuOgxVZy0PwHA+lk8YKGI7PaKEws5eCv4TOWgC16LsW40t4W5zmpiqdTQB29Lb6aM2jWQ/
praCEK+cN959sbmn6aQzm2rSBvvqv4VVXECjtSjlNMQWvM0e06c3KVNHCLp4cK60bF58yUXuTJD/
cD6Wqoq/rmFUM3gUTeuyYIoVTTxK6sKxZjoCQLbxrU2HwAQ51NFgf5QvJlphzwppeKad5UBZvBK7
UMKqqZsvi4JgpFxAZKJpw32Yka3/mjdordswh0KK3NZoomWMf9rs5h049RRoZX9WPs9HKUoD6bLP
wjONsx7bX8fe3beA2z0nMqzLfijMXIaOAceJm8/yYUPSjHK6JyeAfCfss8WGQZhTGA4ZM7E1r3v2
foo7gam3kDuXH+IOFoErxBa2rhL6e/66aKqjCj0gEKeJ/IKwzWa/2R5kJqYG9mz7C9jwVH/A1pHX
woQPu8Yp+xkkQ9YdBQbTCCEbyqOc2/tj8MQ7fFV6CulX5Yw3d5iHuXPc2WZAAsuRx2GTBiZKoBly
SP1WQ1ln2Skmm1OCDWAsKCvLKet+BoTkx9Ata2XsSP0Kfe+4vnNWHodRIt/UAFUeY8dcl315vzci
/yDJ/EpqSRP8tg+iOAtdlfsz4QhxKbE3aKBs5RJXJnkjR50qGmJKK6eW7ilOjmc9Y9mKM59ATO3d
WvLZEbW0dXCshgNDtgX8Xeqr/fryImF3Oi7XY9/Af/RkxnrxVX/LTEIlE53p4GnS6q/W1mXiji35
JrgkEsCRjORrNAsUst1OEI7Eden85B3ZnhE0rVt5pwj9zVqlA/EOiiCeQCwg/mcBRK4zR2745HHD
qyE2rAkelzERGiTngbIalRllr7Pcg78gE4lnsOD6r4CKisGFF6cEloV+VeE6T1DxzwgunM7pfQ1t
Yzzb/H/rxUdfpOW+LsQTaK8qqZ9M8ddhtmHxLZVvcVYvBnp1WbjeWW2Kqi3A3Iigkw3PmuCyczOp
FmpG0TEvs7GFbyGy2oJ1c7USeI7FQGLRlqkdebwKg/IqQsPkaNZFzqtB7y7BRx9hIuCbh/DoEA9E
fzeZYoBp3Zsuwli834cRdbvm0FkTcky3Q1cakiEdDXH+qUivnCXLVBJZGbBrBBInEJnNIFf12a5J
PpEzge9H8iOeTXO17MoYHkOY3OVBwrUwuVCoStkjWDG0tpoKHPq0Cm9hFs+/kWK5PhZqDyatblG5
PMN7nD/FSd1Y55CSNo6yUfNn6BurpCXCR7hENnS17Xz2gYMxl+kT+cJQYf26/N6rwItJkSTpiTfv
T62ebQOwxpIM7MBO2UZTq5GafzQDy/PHTlIjwEBvfx+ZLQX9103RX+/u5j6qkmPRaVxoavTg5cEI
ggdG7yB5qVSOCVKjU/TJcb7qRxNSGGHAg9EBXUi/cGvhkR54mqqfhEzE1FCMnB2nwvvvdC0Pcppy
BEfZNHfdcqLGvM1/lV3skgUfWokaB3BLzq3hwJ2zP+lWx+kX739Pm+pzOA8iVMlYSloOgqrrVPCx
N4+cKvnkhXDctQfHTORv2r7nqd4KWfCzyAouq2mpRPFB1MmTlzpDTys0NuacWelyqBtkSDDA/GOS
UKgDsEZ+XwI96EYxtyhrGI7gTIjQEbWWTtLUARIOQhrZ9kaIU2yjDoUAXfS/hY5Cs6LU8pyWqoFT
djpbHB9gGPJhmPB5bQtxSvEiiKNXcsm8FmQraHJLoMEZ9Ys79EJr60W4dG+Dq+31R8w/zbiZJmfD
XXeigsKpEgJ5ivtDrq3oV6uTjUcATqrF+nWw7KC3FYvF6DOC8TkkqULRVUwjeIwrC+l0w+jH4CNY
XNC1oq7iffQlDS9wtxqXjHEWpRoqE34OVLmwNAGtRwA5nmxux5/Oar1DtG+lNym/AAjdAMNaF3Xd
lQ4lgzYQ/54Ia6N48/RlCCl7MPEDaW1PaxiXzajRh1ioH4cGTRh/KnhyJeuT6JoC/0CYqfpqscKC
afGT6VVkzKXd8iuH0rJajyCZkh2hNJ2ZB+zIbdM4GPZJDsuzSemV1fAYRiQB6z9IeuO6Jt5bQCYb
o04tKqeOqdB4ytUPKrxr9Cw4wovtHAp4a8qpqPPP8Zm76OzqaL3+lm+LPgoxh9eLDt3odtuYzso0
ZQ3XGvrLJa7XyHeQTX56v1ZirEDeMznpCFnmOI1U8ikoucxFNa2uhogPp2eKuNqKWBmY5YsjDzjM
b3HR3+PeRUqz2txNb3Jhba2mXZipkA+67DORxQapZKYzdlOS+r+JO2UTgD7VJfPfetCKCW7rHdG0
tN2b/YLpDyD0FXx46RDWG/vig9Lu1Bpj/ZD6M3w9u6qLkvP+Z+t4eXUMT1y1OHWkaMSm/GsA3NA9
QLHiw6Dutp/pTKF0Cf9aRYnCNP4mMzh5z7Tkda2OJPNOxJ9up+udZqtrU40A3jg76u40db/h5JzR
UVexdGk57DU6U0ywbn1bqP+gZ7rMhvy5E9k/v+A9c6a6fcMegMkUiiq99BYGsgtEMdJsu793Zw4h
K1tfU+uoUxhp+856ptVGYJcB9MnX9zctdYv4/Vml3nwMd26TjVNpIfkb2spvk9VNcju7D0GqOy70
jXJ0WehYC/svdyzxMGww/0xv20o+z/oZ+FYB/0HOv0VblSVIw+JiPTwdJxd11Hg/bJqWs/JWVcBL
lMTaZz0J5dpIeMOQHn28JRf9Hyp4YDCUtIijyAv569W7OORZXnb+kV7lWilgLDCYixTQTmviT4hk
pCfB+rS7BhJDghnkgE7tlgDg2qgLq/Og4EI8gY86BVRRzxbOOKRNRdk92EnVSgCK1T4C/Q8PU0Ay
bCel67dvPu3iobJYWy58IMqJoLAr0ALbBuYqmd/RQ83dXsKGnfBMUeZT7yhZKTg6CdWqS10sZDMg
gnrP4/qpR2e3XW8RceP9Uru7mfN0Mz0ejXBHl4YvulMb5gN+RQ3cm/NoQNh5hJOXtXFh8T+e6nox
b/mRbj6EutzrD3sAUz3Kcg9yJOuqrZq70kuuMQU2dHllqTZrV02Q9LzL5wyqczuRlN9ExHK4a9ZQ
uP16EQVgvj7KZquTwJmWwk1ERbATmhxV+5e9E6nLi3YoLr/9EleKpREOHE3SXXClKfh/UyS7Ejed
A/d46f5trnui2emzUB5/9bAmY5jMcdCqtT4tOMRnhBhf/jXg+kOO9VLixTqs30GGtpRnVTClglv6
jDEGgzub8RJzSyikDZS2R2w3B+jqoA+vwpOGBt0nfGDs2f2o+gb8D6h3fMIM0K9eX0Ftdc80uN4f
b4Yv3ejX3a04u7NtqBzWQIFdjseuncKfhdFUMWbWQnyEd9D6DZ/BXhdhhgD32ke+rYqw7bbQ8ECp
xoJmVMq4IBpExTSs1gAR8O4icdpneIzsn2HAF+q+7c5PA020qZBn5haf8iyEkoe1z6MkZT0Shdg5
1w2pRYmQXrUPKicKsQTEx6b9kkY6nlGPy1z+JcXtXfWNygj9jA5wMvX0hv0SUT/fS1P6sZ2qenq3
Fvr6KTg34asmB0OO2pQF0H+xOJRIRNVnVTgpIuIwjmLKWzqoEEkWWYelq6SfpyX0OGPEQABbrOEi
VA4K4O2cEF4Fc/WAZR2pOBw09eKTlcvIQDLQVNhqG5UWfla+/LWSvzI7so52N+cVm+3OOZCjg0az
nKuHhpOUUJ+o+D9Lt1Pqz7TtqdKHIRuQLfLFVQulr6PDFNHTcsj1obEDMiSinaJEHhd1DmjSsEyF
iqgywOfSI4lnW+8+5l6TkpGI39SX1JLfQhvJxFh54LH3ZhNxm0o5IUrmkGpIlh+90O4HQDek1ZfR
TeylP7aPia0B9css5S87AO2cX6kDfDsFoyMdtUf+ZnphBN3NvkrYcMeX95mVNb5VNxyV15JszhXX
MN/3q3A61OiYfCcW0ZHIsI1M0HMq3Rs8EJWmuefcVoW8SeiDvhyNCbp6FmSKhBIVNUsUiM5jcdp1
/qvB+9PgfBKH0soXKCaOahpTyWcXNYgchoICjr0AlwpkpTecZBHWlQOc4U9n5gbXzZmRwhV2hDd9
Y6s0Jdn57Zg4DiLluyOGhWrLOyqFMenKWJLH78Xsw0yG89vies0r3/eb/RlhxnDa05G6yWecwrhn
QTMWKpL1lozrkRUsE93cfrvS2PtTUJFNk+dVAO1Q5OpUtG0aJsqIYTCiBARlRt4GlTbBiQVteWAs
g7xMUw6jdHBRP9OguiPA3j+ZbYrGmiB69QVrJ3NMgO7wPvOBQ88KntzoCILIYQkaS9yKU+6jLOnp
0qHA0Ww6Q8VJerj338+A23Srmo8iMTvMbUNBzSoIGmb1JLYD5Z1aSlOZ0HJSPspINFpyP9knbJZA
IgKCzoRWW4BBv/3pDKH3qpnz9cVRdbLeda/k6WXzfalUy9ZxFsk/1a9dqEUgi6UvLa2NuRtMZUD8
Ub4THmbBpMHqsJs7R0YOCN/OrfZdSs19kQH60farQI6DM4W62bai1ultiOIEvHGpfuNu1hRMDDxq
tvjVxz3Z2ZXbfeDbdTpeg5Qf7wLnKR3qKoufH6PA1RM2dT0VTW8jChQ6dpgnYRxIrJh6+XrFskQn
xRxwtGhAQSF7jU/4fGBCrtOe1Dibn8MeLMY1a4kH3Zesys9Q3Pp8CC+QZqrkTQjn/jG5O34Nw9/G
hWe03msTYWcTWaX49TAgdEAg3RD11bmPevwapyUHhWOQoOTDt9sUYRifVlmJJe9DGiYfZ5Bb5dh6
F9rl5Fv3gXdNKZPap1KMXLSMHDVDrk2oKLkWa7RIUFD6G9modSgBaIBfm506SZ6zgvBHljye72FQ
kI5Kk/Ym+6JoJ/kmV/E0fTMl0kkbzdDg6JS3JWQQUa93gOF0+5shSGzFYObXmgVZebdF+C0H6uB/
7/eynK5HMi2nc/Bjw31VYLhqH0XVHYDPw+1kgjX722BPJ/fidkteHbWhDxUILTl3Z5ruxUgnfbBd
jECgI84lfYNJwDS6TI1juTQbLIba3vz0NS5kVL6dXtx5xen3NkLtR28RfX2iswQL8yiihZSPfLi3
E2DZMS1Ze8bVxA7eAtlnSgLyOZKun3UZVVFQVxgqWFbkZxe+f5Bft/WSkKUQ7PffDi1RzLY9skT6
bmW3NLZZbAaxItn9lrgphV3kaBM4jc8KCnuuJLAnXweCK32n6nZJhr60RgMeR0RmNCv8T87v+rbU
iaQTmSJSaDdaYJjenxu0fsAQPQjtg14J6wM8mvHS8/0xhhnGeB0XL/g8d59xbSOxFxXUHg2GOe+2
yP6Qez/RHEixC3QhPkEzb/ZHosb1IhLsLIn2pqpuSg5QJfB7+0+J5w6u12nxLMM4ahz+SvWRvvh8
PC6H2N/375OJIC0E6kU30YQqZUV6nVdQAEOGBkd+/Qp4/VcRTk9xIGqO2UPRTUhBnQroLRMz1FEk
xlzFtNzr/XtbnDC0aA9b3WoJMyTERnmmUdlEXLKkrm5AboQnZZGeh+MEvDnMjGFnkabEVlom6weg
RfrG/npFperdDMnak5L8spw/zGWHx2VBXbjoT48+Cw056BTb5BEMhqJPbu/0QlJplI5UCi2PCyLE
NPaNJ+FYeQqktQBQHp77o8W9MfpooTVFC1xLsT+/XYBQSA3Xol/58BFKiq9eWe4eS7AIT3hwJ5y2
DpcJsp0CyatAJmmUuej2yH5+N/Vdy6a1Zf6cykVXTbiNIS0DiBWUad4CeEQEI6ChUqpLjzYI54L5
hbMdRKNLcB2cIeDwCrh8znWir2J9+Zjr+6JKY8XgBvXcGHWVAQncCbrDkiPYudvL2zJ+MpZsN+Bg
yc2DTX/3WQbVNnxyYCzKLsJ6ti9olhidSSiYMDMdikpXe7+S1ObZR4lFMdGkAMWbz6lpwA9HJf0M
WTOiLxCtMXibBDzyclLoIjVeYsOcGUGtKZbMmySGyTmxenc/jCcv+MSrsAsYJufbtRoAnBwCorMx
X0iE+twGMC7p1LHgZeHXAq2mOMt2qvG35Liol8Ooqhm9AZvXAAjhpGwrgeOQFNbyysJPFAN8g2rZ
gdFinlMUHhF86KyYRnlL1ODCyjTT+cR1rWBEzwwTEftxd6lFitd20M6wF68T/roZB0g+EVJSxDiU
lWMKIMsQoquxu0Rh/lMkuH51Wkeg+2x6dP5H88zc1Osic8RBzwlGiKDQ609gfg3eRiQhTqyZK3BC
arSEG/SQNTqQTP/w15BVQi77IAvLGtmND0/qx7821ZYvdgQfjyrdjZAaM7iuAeOGyfNDTsTI8s7Q
jM4zH+qxxg3QH9jKH0mtISr5ILf0Gj/WDlsa6iTZUuuJ65eYd7s0UWGyloyG/9PDtqc/GxidAdx9
11DOMFMY5//DA6xPABTho3pCH922PuqBryzcjFE+IvwZO4lTuYDRC22XU8+nZph2IFKQJFgNaZ1f
Cb0SBxufSkY/OvDY/81gEhIBDAGbC7V2DDJhq7ExWCEYZ5I4JAqIEn9uca1nP/egoyUSirX9IsGM
liKLTvVGSfC7bKNpopHmQXq9X0fca0BI76uCy6aLkEQpuUJWosz2TMWiO6U1TgJD1L4+kwBn6I6o
SOhxU0Dw07WaJme/l6B+8kIv+zLzzmOSpgmkt1omi050Y1zuTRxkZHRtVd/YjX8wEIGtJB38ZqNM
foK66UZLE8dn2Rs9JIkT5W0nTB0uo0mPxJGPOthmb0vYi4lt+PMio3SapH2ibL1cm8Bc33eo7HgL
Wt5ljBC+UISNlu4iLiGqBVB9br7UyEg2SEAt7yShXvvManU9OPn4ZiWm+UzBgKkZl65uP+/FO2kK
j/Fd0/R6jGWMS66cXOUwTK4JKeTdOHUx2vY59ftd6AmAChYGBrN53ot7uVxyQYco2Ei4fIuEVgJu
4djYpNLctxYAqSQyr8iwRpyvJz+tRRsC2hxq+GQebos5d//I/NV8eszXU5ecyvEyFc9Z0PxTJwa7
p0aqcEFdyzAxujv/ePhrJord7pl/Cfe3h4k9rmPPgz2MnIa8YKuM3NNGDHnxN6rNd0rQlOSO+Qoq
sgIEBVN3SAE1Nlm+2Ijx4RwfXfVyicWDJ3EihPmqI1FvjkhelLvK7f2pQTZtFDDdxnEkKe0ghShk
X/Rrw85NNkryuRcqbQ6xzOtSoF6TGjzXkjMNBj3gZC+Qx/X9EwFQ4GvYQEehzYU3WL/7nb6QCzeK
7PzDO4azgu4xGsc24joq2s6+qJ07FG/V+2m+ZuJn6bvFZG2YNLZoNhEs4EaMcd40klbas3hmHWJA
8jZQ9/2+BmlHBlUUJNH+CxZNpf5IhaUwai96Hcsb7hFGsNnBgYnvF/mafoHiqF43DPK6PXpO/BnO
U5A0sPi2WYMavDT7ZQ7Bk3q9heTrZpVzuotgafF07NwsO/2OIL62mJflbNylOy7OlyXsj8apItuT
DADRfi1zoj/5uBYUk9egy2TSFtMAEgPS0LggfTdFYT9WMirGeq6gJO2ux0voQPDUWo0j61NeV88a
WcHOcrdt5iJxCnvMy+Z2TfKkiQu+E1KNe1lH/17ApACEflaWvtXRY9X3EtRSY9wXjNUceJdcxjEz
ncz9YVMZYrqiWjKNqhl00yme/phavJOlfbuMe6chxXIxItumDR0bihz8cD+mLZTtqCyLBrEeEksm
T7hL8Zpb7gBH4Gr3aWhbhwRHLg91RhoDsCYWpAEIAhNCDNLxULH7qOFjxkF3oy/L7c1n11PpiNdW
8kQi2qmqZo8TQVsY6lOAQyL0uO35dSM+KfbQCDwZ6nWkNaNBWTpMkqgJnV75LyyUs/Ru3WUpwFQk
cr1Ax/tvVid2cllRO0Wb0ULjR53InkndaIhykFuGEGsGEsmuDgxIt7v2iayq5aBmThlgSp/Zc14L
NfavlcJ6hCPDMEQU+gslg9UCdZfR8h5r9lzYqSMrvwiC+EeHeR5snqKjh+PV8r4CoY/mcwHAM98J
Oi+XWxUVd//hi1/dJHtEX9m1LiLcZbzhtIMR6SzgcFrbrVuSiKBiIR0oHQ3QgXvHb59vRDYWGaUp
8jmdIMifiHa2yJdnIKin7v7Q2qWf5GFwPGaFfB0sXNkGbCKDoc31hflhH9B/FldSWMRq9TupcJj6
LrMozyQb1t2OLpE0S1Y19JKnhZ4P8XXhmGpQ6e0b/xOBPavVTnRu4DdU9/1Ct8aw/XbW2/5PSbMK
7AH1MszJKGdeRgn2eqXrJqzWqX0fDywg+j5j3oNRrWKaUDhuqMVqI95rPgiQBJglbIre1O8QMQJj
97yDnIsmbmZEBG0TlH8UTT4K+MK+WoCEAvHZaAGo392HtV81hL5+18gMA5WhEMYKMquKmmkZW3O2
RIxh9nn+PTb6bbbNO1SGmis/uGRr+naALRFi6OnNYtjAEHrDdVSkg2DzYjGiOIhidJrHVTbp86Hs
OcN9+EmjTvGDftmpYmZldIqBQrBzMCTp3xq8MVSaoS0P5xMoVbUBmChsfwYJltWVIN5iMML4EWlN
8Wl98DzictBWXMKz8+bQopK1P+758cto6hlGeK7aItRxDoo4gkeND0f8mTaFkM6sOSsTwB0xmeKY
+s3sa8g7JPaYYEIzjnP+5sgc+jIxv8s7A9na7zr/1AGBDT6FY91yhV1699/wB2hzQWVXIqSsC2lk
5+XKZlUxylyCAWEMVQs9la8PO5KELl/U3joZtd43A/Sa3/AwQiAWkaqxopxbituIfGinsSJp2cYR
e/lKNeLoJJ2lwMmM8q81wNMmYygZgW8zMPNJDcUOytHyBaHlZqrfaaAm86idbRIfFD9qFkty0Hdv
Ra0TzLRbykwq7oTAIbu6aJB+crHDXZZu0clFAUds8SvvnhuziEQP2023v5obU0doh5NDO3BEBUM1
Y5tx8wndNsOs5tz9Y5RgkB1g2rGVHGzA6v9feRcAMATPfvOwEDw49KvEzqGM5nmbrKXSosI8xQ7O
dQ4LkwQSQTh0MrAvZxVzFC08NYZCuSoRzItqKqkk8Qg9/8OhAmKJi0iSfWg9Kh/2zmj6eN+/Eo6x
Sr8vLOjY0DGcJtATCiEQjwncIPKVAGoGMSxuWx0cN8dxSwxFsPkxb+YY/4Q8cxm3rCwwpZmUQKOR
3SoAcCayHGmv9KgdUp3Z6WSpWR0bFBinpTdKH914pOLXNHg9QIpWQndkNFQKzeIhdnWk3s/Mgc0u
jYEIrN8SmI3JtMwW821+gKZLAfqBhMs/Fs4Tn3evO1bQs4LXkFk0ZCUf212rZ8SyNwgFdAfnDxfv
wu23qKonDVnabAIx2YZo5Pco1cTDBlQVyybor9QfulZTyuZOgttggV8uMNsQDGKi1LbB6LUDZley
YDV2bBeWUtkSQ2Y+B3EjVJeRP4ICN0z6G/qbyU3AbKz9OywhUsFjKuO2P34T1jABtfyd8TtAXqIV
bPapA/FUqaAuSatdweqY+1vnm7qhljh6p32VpTLieTMW2G4vnWZa9Jk0Hc4/VZC1JfKabuOPrBO0
TyynU/v2+n7iOnXkpo8F8c2WRRy5iLBIHSaAS43io0LS30KElpehQtA/pL68tJvtHPIPU7dtFQPG
N23cx3MhQyLqUaAzG0PmPhrg/x3wByn+G7i8bIWmrloaUUdM8/dnJGIXwFibmnDa/ZcXrBRgQB9v
1mgn+rgcWHZ9Xt4hz83Hntwb0kjLot2Sya5ED4QYY3FpZGDR8ikPVkqwiO9U3PNcwJUDbiFrRC4V
tN0v8CXiNezKn0xcJEE8VU2TbXZJyz21l/XV08x08S33KtFPUCHekc7vTwqupKojJY+2Fl87sS2G
SZzK9ctnNSBuZbC5bkEy9UjC039kDOtJ/Zl9Jmy3ZeUBXZGEkxAai+QnMuPdC+DG20IhsCXyPfMq
dyFtHKtzZHW/yR3asNkLjJQzXHuDZdFw6NXniDAfxc8gNmbE4PUaddYhhcZs9XFAj/gdJ4um20F+
42NZ3tDLxs/XSeNyhDliQpAUQy6X/vMDgu+ZrxpejRstrsCbe9eC1Ib4pFw5hAKyIUQPD7FMT67w
4k8kI4fCgcLgsMsNJR3+O0dIg2gBSLycQfgu2hJN0pXhKUgzcURBSdNmUc6rSQgVSwN+YFBnAC6j
6uHIk6ax69U585zoVssRdWsYnu3BABUvpPb0DCM410LiEY6vI5gluOXu2IjCKJuB0x16U0rcVefK
4xMiRZ/yKYRDrvUl1JZbsWOBqPrDphaSNKaKhmca8d/WoUCzkGxj6dBeXPqataj26I9kVTqte41K
Ld3t7ol2iGIHhm1f7VqqM3/AVgjL74mLowE7np0rFw2vjCdiWlLQGBKamX5u2rvSjrDGK+PhQLBC
SmjMKIm+oUwLIfQ4PMcxhm/iDcclYGX5hyo5lYq/aGnr3k9YH6T8E8EV7ASTf5ZxgMgaUZoWy2yD
vMNtNmN5qfSE0sf2tHTlg9BpSs4hy7ZaxowW4YbwJboyGSnKnBeYmzelr5Bap4hsOHvuMmcMhZt5
6VH3t6I8GmLdsvJEmr3FM4rYje4nmzQKqp0f+Y6xDqfH6ulEvYaSfiIdZVymfjDleVwGHKDcI5Rh
JHLQHe4TvNX9mZq36hw7z0cVRbGaQ4YeCVq4afbw1AjL01VUD8D19Imk9VgfqugbjeVkBlf29DV5
z3fnpblOdeW4MpTak2kkoeBmU6Exj5plYhqYDcz+bRvx4+DtPRSSddW974c2PJqm8fP1CytnXLWn
JnhJKZzYhuOSHZgIVOLuvQOsHXSmEZn2QWetkxvehXYF2zkfk/cWQZVdtTqBlP+F+MYDDJq0KUEw
hxiM+AvbrhKU4Wco3kwaNvOwVoHGFhE/KSQX1DDZqHvz/I7KSur+AOpUAogNP3rHj6Au1PRULJq1
t3W4Zp8Fk/gEgdLyMxcEN5wBQDcxGbPH4N3lPqTbc0fRcLzkHaBHu8cHgIwqr1BvcqZB0JsuSj6/
DJHL13J/TvcSF6QwJe04QAF6FnKjZaSSrqkJqTdwG6ZD/iK+QOqo1CC/zaywLLuCzBGr2KvKdwQ0
jDGI/dyYz77/KI/Yg4pIOJ7o+S2j7A8XdRUOnyzRuH1D/LBJX3Io1gkuuzBrh9BeI9Bi60sB/gbc
beBBnnSVK5cZRCVq/TNENHM63VQk0kFHK3ImK41DMaplUX34QFihwSdXA2XmgTGKSZnLGNsLXUzu
c0KLQ5yr0U0cv6p58xCL13X3Nvhx9y93ouTa+j0k124OQYT0V3PMtpNiSOtBQ5/NN4c8QCSRJGsA
nnJPcpcgIhTroLxv6OTdl7AiYfgFzEjB0j2ymVKacQ/UItPDj1H+13J8iAHvVGShZ7a12TX0crWs
rxhbZEBmp6l2wTcyCWcHJlEKwaJsHa92Sxf1ZaU/0DbZ5hrSh6rWNp+O/SV9YbG7U1fULgsozUFJ
6MxrGC/xWbkkLzae/L9Xg/C344gEkcRPGg50+kZQwLNzxYqK4AaonNzYyV39ZB7A0MCNlRsMbJgI
YR73nLhkUIwuJ2NQOd3bXCYYUSfSuGXxvGZsODT/NawmYk8NyCHQGUuqb5K1wR2E9ych5JW7zF36
13WkuJgb7ANl6c/FbJ93qg9GGTimFxvmrVO9iIcMNrnWjlTF/WcjWIaeeD6lKxzncX5IM2ye2fth
EUTM7ug8WWx3auOb7jLefO02NaWMcli7rPEbfbB3UdA7pi8TlDUtONkWSUn+CYoLl52h28xD4U9y
NcMIFype9w4seXIAkJtzjJY3wOUT5fawEXWm5B6kjF7bHKUdV7prWYLWs4fm/Uuba1edta9lgnzu
SxC09DZn9eEo7r/GwCJpnrRcqBDuOtKc8SOQu4tTVF4tZG87HUY0uxzXBXZXaOOby4bFCn1yjNAV
yYMlcGvfYOxbW3QfakY+EPA3tTX/9oY3drscDR5L+zb0y0RzCYq9RNvnJ9qlf6Lbk31vvGnWsJyx
a8ZuYNRQgr8Af3m2PPoJb3dwafehkw9MdQMSncm8Ehpe5I5dZtyIKcYCPh9YQS8YzpZzicjNloyv
2QZoKPZnX6X3YY0mz+rf+6fwf6eM7yEka1dtuLWfheUD7fGRdUiTz4ohyHyfr/iXmXMubWNxipG7
BsUBZpdb+UjviroTmbS+lgNcf55orRQKXSBj/N/oJZfgocytOWhvzo5c1//w+Odo3S7JIiTM7N0Y
JeOyxN/6j9zS26Gau3tVjANraXiSKjhNHlOgVSDhRdOjz+hOTl+wx2B0P2ObKEHuPGArZQbUhqoj
mUgrUH+4NTFatbS8t1NxO/Xo2Z22XlYRmdP5D56QiehSVo/YqBF4ni/X7IKxSSYUQmF9XsBTOt2e
YgnwzBGP/VPYOsHLgRfntUztJI1uccbd5Pt3MibzmfSiDngV185e/rppF8Ao76w108SEStzovnT0
dxz2LJgBH96f5WQDdR365DSFVdJ1bsfVE6t5V8GbQlEILRLgVUs2uu2o5rfW31bTXYcF9/9MS3B7
eOtFHE2NOniOdKPI7rh0yZOsVcuBATygygLTyFDY8OWhFymDvGc7R0rWqgG8KMjY0KU/CE6I9o9x
j/AaeuxThRoj0YHPezg6/rWCWQd2rqAvk6CGjx5e/d3lgJdHQlEzYlHVr1rLlcOe4Zz6ET8R6qCe
UIGq34brxYHdH5yxjqZfxNaVWQjVRU/owTofeEP53kTMeYD1BHaOrFAb81/4wIOZ2A6LYdq+yJ//
ZQXVBGYf+GQmwg/UtVgK+3wkaw9Qk/qpzHCk3dtYghYtSBSyv/LtuO22ZXuS8+U88SZaR026t2zA
2IdDdAAKxPVNt7rYGep/UHXACqxCQ6+NSP9GqvtjpVYOSiQUTdHN23Xsryq5cGuHikfniuwc/Mpf
ifldUNNhBzkfyIbpQbtdsJ5bZ2m5UVonVxWALTdUDR+RHnfxb7hGln84AbDHGadRaFW7GFBjBkjT
ZNa2BXgxS5E3mGlzfX42T1qkx8iOEcSFiWfk4/qn0dEeneBHsF13v9774jwkln/rnjcbVvTplv2E
IlpZhTDI1rnFFtcFbfkcM1pjDSOFyrpzqebScKmwXoNKMATzZre6TzMIWwbrB21xPkWj5tEUsLvO
I/K5CtOEqddCpgHr6mI3kD5yzaihADlh7eUzpiIqEPoKHzJx6qu3aX0DJteqqm0cI3bZdXFr1zVo
6P0Zo0gXW5h4tNmsIfZNTzNOexehpQAZH1+hMueoA8LaXdz3HD7gC8JMN8DKKpxHR6CA79NUGnIk
bGmrf3rNy1ynTC/mPMkizpzMK7Sxhq4bAFjzMbVkJgS0fjnZCeOXQrn0s+UWhxBz+GUT65RxFqFx
u+/vbOPOO6DebkDcGvnWyCQEHD6WWDpQgW36c/Lz9ffSDDYrw2BfEv29RtSzn3nPQ4ksByncZ9Ir
Ps96s0BwkHawFeVqI5g2ZS/aSth67CL8GDBT9kbUK4CCtp9tlKTJPGyypnRcLHvcouXRpxKnooD0
HrnGXl1tTjG/qdiYxK6OPQRgTZfQGLSPiPpDwZT7UgTapTmOM6PDroQ0+Ya6HwdKk6PHDF+3iWRR
5mrrg7kdEyDE40msle6ArGbmIEvuybE27ZjGdJ8pE1ygjg6A95fgxN5+FyEQqMfXn3O74g5ycECf
waArnQ/7BGdcDEu9MC8LAH7yc3MKqpS2v7/dDMF49mL46Zky//tDz6F087Zl/WPnj8oT6DAsQpbj
ek98lhLNHctUK9+j+XMM3fNGMwlzLcURwzoFq3mraOGgbayBJK9eWuU63jPqKsWdv1dUk4sd99nA
+MpWuv/IAcv9kG0lHAPIpabjQ1oupxy11ZDW3FodYthxRG6MQGya9ITrkrZKm+bERZCZjiMYqe+N
zUa7Yeb283o+DZ7Eauj6oMUgg9T5gqRgrudAoNIJ7L9HINdF2oIqZbQUkmNMQiMuIMG1KsEldZTu
KaW4pVgmXeTiQsb/pQjDSw7wRJMQHW9KOOyGB8gaxcaqW5OD5Up2R5MWZqHWe1D33jsQAVShP/df
uiD/m6RSjba/smkGvNeZeBa0XZQU6tIQV8zCj94qASPUJPGjSUUivowr2cCltd/3A460LruPxieQ
Is9N+eve39xJS5wb5FApm71rP8dxfipGCeXORhz5oaN6OyhjAxStvMbZMLvWG1uraIHzDJ5jmp9T
hWm2sB57Fp46IbXZuE4VdHs9VktiuPkkbQXO23xmpCnIWOyA4w3ANN6w9ik7DZBTgEFOBGf77rM3
baEvD0SmbwCTc5/OxNtUPJ0vJ47Ns+y0oT7dwe52C2D0hI6t4NPU/B3CwTY0ZJ7xYUmBU/V4JrIV
A6jCgInWDxTfUYwm7pHo5hjNcwDO00XIsfnDmIimhYQAxcPoQwjEw8D3dSoVWVssMiu9J0+XgiVD
5HkGMoI13jUEUZWaUBfVAHai8dYfTUzRNDPVla1Tf1kiLjuxLv38kXpGLDwFAYISDNZUvwFD3+lE
DGIcC5ya6WE18a5ZeX1sHNW5E2EHqNB2HTtw+BnawKuMIT2FR7WcrtG2opfRVcrOBoHacK5vablh
rX4H78ceyU/CjsBWSeIjdCmJVDqI0CCL7+T4V2AdR755kHMAVsz3cgXHULP2I5RR5nvY3PqdSX8V
fTintrQn6kwFRzb4f1tdspuIFmUZypkqHK5ypxhPNxCFcb+z/fOkDaO6V44KEx92qPEiOtlcqgO0
9le9o8URQACt3yHkzLzkyaLGv9aaw5tvK4dQMdoELi6mseo5dKZU/n9gGe7w5yStSlBCD5k3RUni
Ln7DAri7tv5vy7ReiRvTtkW8PZjk0hQMTBAQhAYAMmsuBItnNcFZIZE59G1OlxG2EiU6raHtZpqh
sh1JzH9U17mlKuaIceQaDR7hjktVMv3o+0yl9JbtB96Mpa/eSCbFDDP2xYBUHBtcKBOWLRPTaW/N
l6/A9UiEkZfZXSbFDR6qJXol2LenoFDGBn9atXDfH0TtoHAxgs29mN/7ZuNs0T4B769XE3qo39Ij
OSOP61EGkgdOuLSjtD+AnkfHpKcZN4Fo///ymHET2mo/AICTLWE6XVm02MvKm1FAPyv6EPzRabGu
wwDVhLVbRrGTwYWzc4BzXSJkMDBi6t41vpj8H5LqLfINWR795ZQEyndM9p62489c7LrkKMxesAzH
QTn9orVjOX7CDATxan+uAEipYaKGccAjoYRXYMXnZ81sD5xgj2G+Y82HVez3LJmGEMwswGhDkzwZ
ndlD1mChjXDHGGozrRF91+ufg5hj1r24A7+2f5V8IrBfUVEQZhKc1katGiE2naEtJ9rzrtJJzOfI
58gerSO9O3ksvBt68K8AubXQMnviKdo+cGmnZ6rBDFGAn4UitUhtyFKRzBomyhaPcgpvwvpAsPWC
pK7s3/lCqHvINMhTLLxp8TEcv5ku2TmT8PaYm9Y6pR8ckfhyqkSHtuu/2wCdu5+q8pKNjl8H+ETB
q59B4j5+xf5OxJEgWD32JSB2TOXJsSD6+4a0DbqtQmsEoXeTjqtkdBv9z9uz+Yq10CBVPPxDPGkQ
DQTRlEuwmmJLLVO5The7zX6tdZm/O7O4ATqh5TGJdRtCGd9lPzqEoPekHe9dGGp46+vDNJXH9AiE
vjUiTIVFXJZNZRA4KPqQivmf3ZOqbltoq6bQ04kSllUbrTIKMsdkA+lFVWnAgNEmZHVXIDNUkE7R
Hiaevbmb2MjQVEoeKYYOpF4Z8qxsFPHqlErxCnou8CHm804FlCvALD1DTNEu8YcMSt0sfVfzoY3q
+sfflc93Knne6ALIkZbgpKBO1qqQMNVtuscJmz8k0wGJw01R4v7bRXAcS6ckWYavQu8wt+Kr5RTq
nYNhWEH+jJVd1JYn0XLr7yHSknprkIltTwpvYBc1YJdtsnYmGqCGzZzP4eGjjRy8YrPfuYSvZYi2
FR4FSY0EwY4E4aLJgnL60LQk0LUrjEoQ5kmPMGH41u2rHeO9qH6VxCN29miW29eIwkk4hTD4ytwx
2wzfUqQVApDQD1u1JDdnej17QeMfpkQyznJbWQuEwqEewdsvEsQ0zmpPlg04/r5KopKbDn2ypaI0
K01PVTAf7W4+Z9K0aZkYWxcqRzBPemlUYhR1UdbXi8MJsArABKe1HLmRwOqI85WcyReVFsXY9pSr
4usq/632vYpnH32OeA9/104EST7MtirF7X6sSBB2C6yFrsgy+G2hT61h60ZS7bs2FOXW61YDb2V5
Qt4ynVmQMBbybq9MS/Fq7Xs7QQFGKklWXJCRMDOBgDsX2K87D2w8SwNCScqqLTbSISYpVAPlrAQb
jQu8r72SGbIhW06BMp63ma4++VLD9iRUL9vn42hptKW+FFkfoN5O1dJsfFUs+oyB6sLy7yTQorWI
eFjj+wEgPKaRmjB8vgiLSSTWJaIkQURDLjXg/f9+OTjsti3ZpEhqXbxg9nUCfDBjtW2G92CgGS5O
LwsmErdFi1sCB6EfCEbqED+bUh9KW//6HoAixmhhMJVcScFH3MT1ZDLYb2vkACvVcE+fXIvLGXwd
yeFx3G2Z12hzhWybTcjVSaqfhzSy305nO37s2KLXBLdGvgPEPwnxFIiWiHyQdmNVDScfGSP0BJUD
jM6GJjhylFB4Gx+LXTgtocXUnpwj2VNwunfVaKn+2bgJF9MptJ35hQoGq+XMRqseXL44/S3q8Faj
l7ob6iKz3tRYTjg85x9ja5V62FCeTVhKfyv0HB9t2Jczc0qtJSlgOEQ64YC10jsBysatqR/i8UEA
89y1WIK0BKnMhQWI7oiUdqlhPcuVZiBgj8jzK7ihZGbf5RUBdOROKpqfRWQ/85aJF36iA8zAW3jY
fBAnzr1/O93XfspsS6aNNv52Yq5CxSx+qJMVGXZipHnZjr7uvj60FN+SKYMSg0DBQPovZmI6Fv3N
IPBR1MB54tgVE4FobQEDvP3xYsa0he2s3HkXR0kxF+A8SwYroX6AL1/DuRzt/ktdJts/xYcNolRu
x6ZbDvW7blWu0zVvE5pAxp/SeiSlFYYlZwfcOP7tqSXIvUWXUcUCOXOmnOUdONDSNobreC7v/yJS
T1xPDImUwU/z0nBlHy/HLc44tuKkwm74y0RfERpSMvfLAvHTdHnWnH4+nn0ESWuarDfoIu23ix1o
CIzGDsL4srRGX2m2gWGEtWCCU3mjYsZqEE0Vpn1a8X8cR31B7oNcS3J74B0n4VVzNjI2ZR/wPcn9
eXVxhXQ61I6y+wOZPOCUIqLmmWQ1tUkX/Q/+4HQikVBCVgt+FNiiwUOiweIMqPMgV+D2Xw9oNOsg
v6L6RftEKH8yq/439DPb+mHhOwXLtxmXgy0oYVWgAcU/fiKXIvkmgn33OfFol5mPs9ZzR6mn+awA
TnEFWqeszpqz4zixJ01sm+mPUyfYVEIz9iSpBWrKgAmcSrkriyK6NoJgGAmCedz6ZoqxmXPu5us1
7Ut/Ay5QEkuRk0CmD0qPiZgUIAOomnu1Z1x9+GvgFU7MPgjDWBB6DdMVP9NncYDDEixfcnJH5OZV
Oi048TewM6D+nicNi3LnRSQDEPeYxSyImXZfGtktr+0ERi3ecN9ty/+6g7wDqmiCAM/vi2t+/DwU
WUnwUL62ncGvVYhtiLAb4wr84M4WD5QlLgfR4GFkuPwiwmEeIOEf+rhSDeteQhzWADErEEHQCGrV
dzarapoub1EfyC1djLYvRnKJemERrsIytwht8y+FGe6jzM6RQvCM2KraQEWUqVqKjEtJw4kGGdiy
ThH4sVMuUCQNYiwrDFXuFTtDKj4U+mvJVC+bfuAUGQSHx0V4tXDkUWZg/Hfy240xMFIUjGmZcFAT
9P8X7uX5w4ocjcmWEJa9asUOvl3kDp/YxLfq+VCFVSx9gMuPkI0R1ou8okncWyKtLN0Wo0llza/1
VIsRcFmsnHfSqYOB70KM0E3kX849kM/DdflCZKYBOuCMzJTGdYB3l9lgad9Mhd4+i8ICmeUW0bN/
zmAIhoZ9ZSACnHj3QXRWT499LZ5kDDUN8QUhyfmqkUS/+zkvRlM+QY7Ji9VXIX6jjmXpKHLpsZgT
0mUsvSpHQq7PHo5C8S4O5BSa3Zwc8wEnrt3Ps5Qvm7nwkGGBevbQ1TpDUU1S0Xx15AnCrfviIKdw
fOWuDRbx0LNglKyRPMI8RU/+JKHWbqKKDTubjWNeFYmu6g4csO1VepVGjKzg+cy4dZxZZXv2vGgN
jIE3CdZSxXjWzR4myKs7l8qXy5I6G1KBcL8Xdwmp2d36uAhdVkGFZ3G82rs0ocEFf9cLuN69Qraw
zm6d7unBut1npDVS7K30Be84eOcXPVFwAOyEkn+Yfi9SLnwTRdmcgI2THwX+8G7IbeoiJZbB/ktD
XFGHQWShQleVkuF53AY/pAGiPcxsQlblkW3OaZ+U9qnGCNXR6/oPb8R/rHyQZu2rNz+rYji9w5Zt
Xo+w+qrTY/ylKotmKQquyWj8wPLubJP+oLRsmI851bv5lTCmRJWi4PjADLHJ4TabxaudKrGccuUW
3fAJGwcZPsuNa1pYDl58RFgtBGg1bA16OJN6MuYvNhZS2J1EK2jHk3Gzw+XvV3bhXkAlbe7oxZWR
cvnRhFKUCKCg9EQ2n0SHH886xHIvPAjQeylWlzSBYll89+I5Mf0MlrE2FgjNkZPzjs8iUIw9scnh
Ly9ZgX7EQqfzdtzqn/9aVgHO7VVAYVCvANOrbykus9mSGsNfmMhb2Fp814/aAubVeHzixi4Sz0Tf
2mdVHTJIXWPdJVlVISTSmYjMyFOE7DTezU1mdFK5G0jfRGHP6zPokj2fhGDyPXL+njLnL/ymmoBe
Uo9k/ielvIDCxmI83NKnoDyjdNRadxLrkkcdAsDnjP4HzVOBosxi2T4+xdWLeHWY0ygT7MqA2kry
BD8JOQKmYm0NLpN5NhGiOP+bjJ7Sqxu66r1xm3TnQ7hBf0fqWDG8LrpJIdquB05hTg1whUT/8cmm
fKZE9ta9UQm2aCLIfUPZO2lC/F0oW+vX0gBijidtpTBdZ63FW8L88GPqe4ZchJw9hKQEPQsyAYav
Zi4Ao62c7b2LgXTUGlEtv5mKJSHVWT7NpmWzGuPGj2XdzKz6R7CAIrCE4WgFAGdEr7mkBSjqYkxR
0CegioFG5rEjKB4g0V59EdTl4CBkImQvJphPNR5+AJ0AxAW4tOVTsxFTR+1IOY7gazJxFRazNl3A
uCE5Hx9D39PpdwZYe+nb8Yx4m93WseZhkK7hy3Uf2sIRGbUVT4BOoKxnnDqXTK9u30CIsjoLZ9Kr
kjoOEBdi+S4vPaKqxSPaM5NlEnOZQX882qGSe7UoJdOD/PwQr1GYZOWmYtE/3H8Wnm7lF+X/rjQu
zmumjvw8xpNivwgRNvGfBDvGmYPccf/Gbz4iZ371lx/H0Z6i37OitPxVVWb1lpGriznOoT7XV+py
AQRzaQ2nAHvbDZmjegHsxzs2gCco5sfyEkaY39uRVg6OOnkAHQbTJDzwbiI8aAmeCs1jgV/93Tyf
zt5TcJElnS3yYiab1ppNb9nshobQMgxH8vh96RE2p5Jq1z5K/gh0jcPKR6PkIll1wjlAuDuk/8E6
WwBpKd2fQzEMZ3CWYkJBa4u8vQ6X5LUiqPgFL4rI5Te8k/MfnR8IX8XkWDNpisUmMd4Bv7zdHKxN
aONFqsllr0XEkA5B4ITJ5UWLPQFAdTqWfm1HbMSjd7os7SkyVUuiEihny4tyRPzqL7x/l/HnUTLn
1+IyZg+DBFWJ1qFO+paqciorMl32jMCnyBgnNf/DORXp5UoMsjrgJPiEZ55VkRzget6jm9X15WUs
YLMLGsunvJhGnIIZCfnhkNfSAeVru8iAFgBiEHUMLqhaOxeOSU8XXaADtwzQ5kvX/l1xyxdCNKm9
xbrEJoXCmPhjPQgNTXQgZhpvHE91VcX0NC5smQBxt/al+tYf/KGRXvNdYabLalHiUcuyvOwJqRol
/Uu1XljASk/Yg23Y5uaqckFxmrkbVNUl/uaOBYbIMo0i1k+Cn0JnWFE7s1kaKc8Jd3MO1KX/RrdM
KbIZyzmT45lxIRnYbmlHljPRpShU1aOD/tGB0stm/0JkHuKLTc3cCv0uspNFG5rSHXMG2ohrqeq0
4dc/D3s5r/ltA+KICyc8gmDZdf7T/mE8YCSKgRPQe8p9YTphuPKAqIs4plEcRCpLb51kZhlUNZ3w
75ovghYS07qv6rOB1lRfKINmFODbEiizUQ1mAe6xG5xcR6AwEuYSOYEiKvbjyC2JLVg+YGpqjNCE
R9NJhDYodZfiEJTj67JtxaU+3//mxe2LP/+GCPAAFol7jAb8+HeksUILNRyqPoMm3gt0lHkr/bVi
18jp6D1Z55ml5V1zynTW8MRwN6U9apPJ8RByFk1FXrWdYqu63TatSBAOxfSHTxE7AgJoMk05T5Cc
fjm3vtTCFaV/hEzyLWifEM4/jShBt22c3I1ZYjSuzL/23Hlc6abaxZx+1KEneKMdkwedtaH2s9Ii
sv1XlRGuWT3sKK4+EPBme9UembhvJyA6MqdvgigJ+xeV9BU0ytw4Sz5VZZrVIPtk7u4J42pRewk4
fYDvceDY40aVr34gks0IcxkNOHuU4hnEoTZyAvv574o2vdYekxV17bagdIRvM+0ueNj7FM+GUB5J
xHFUZ6FyGh0TTyB1RpKVJGj3C16FbVojb5Rz4mYEoYOS3bTilydtzX8yCAE948C7dC6mZsCtv/LA
SMX0r+c/OzZoWwo5OVqM7xnyTc1HMlq1oWulINVN+hKaC2dBgdqGu6WTTvX67YilKQmAZfQsmwGh
X/KfBLwgdI6sxaH+H8jPzPvJ49sxwUjisSBulFZMBJyQsw7XTGZQolDXrZATx+eT4oyfUJPQCj3p
J0dhw9KHhAynz/XKuAq5wPhxZp5T7s7IQAAQ7SZvQXp0tA8KHpzDqEysFAabZvZJqPesDNZAOoTY
4kpSXCQ9mCcGQip5S9aze8cKrAgO3xe9gkQO7FS/qHD5Yd3K9sFZbFxe8QxSaWmQJ+gp+OvM37t1
wcr5z51pJzO2QUSS5JBGgI4xZLATJqSrovLmkR6KGmJRsYClbZ5bdI6LOaPWcmJHzQ29MK7PNqaP
2B8IgwF3nJx1Zhb8fpTw/Y4zZ0JydBuN6yw5aOq7oqcSqMQl8cxNOM1GvEoxMd4MtvJ0XkOTN3P1
SJkH1lfgfKAEsZGt1NkZjTE2G7pYFqAv54TIrVQbU5ZQleiMovh9pvHPG+TxddCkR/vT3IqchKBG
AhGfJg0I87IZI3V3JNZ2T1LOHGUQKH6UuaChD7p62dq7V8b6nJaElHKQl50EYFFYlZm2G98U70VO
ip13Au/0wW01OfygkPH4O43KIm8qF0NTQmI38CZeuP3zr+B0Es+bthTIMyTq/jwqWiCX7BGexwQf
b7WnBcTFbkrYazj7yMxLYQNG0+S/3jttdRTLwtzJ9i5uR5CG91hrZJBuligdUhiOwb0UU/u4tVbZ
ZyV617PLasjqOuz5s3eAIPv42OIvSddnSCU5OVdvMTMzwPWHlO8g/R6FkzoTqyioMeQPhTl6GFAn
3zFfPEa/s4wAFhsTgUCDJIIoGaBuMC5DwqEl858CJ3sD8+l6YRuoD7Xtnoh1wM45gD2eXuTUW8xK
szMV7DQ4+0GlNvE/Zdv3m5BtrYT4us5QUGdemRHZ6OdliHK1Ft0KkKhx0nD4Qt6XGCq4c9u4Op5v
e9TTOMvZpt8JVulnFmCdZw6RG4QAvNCDvQheN+ASuLxyyxY1EZSiwUKLFk/KRbIJlXUcrWV9vkfL
ZUEHodQK3/QW+BdYfDdYH6BqIt2GA1ZMKbIk38K7MDbarPQxZKcE2Wr/ORp7VfysY0U+gGfBRs+h
Bcezhi+76huy/oOJvSeKBvjgFxsw8N4PtX3BxgD8EDi+wF8B02GQHmSBt5p8atI+8JV2TlDmD0kK
C4FLqW0oyBpnPsyXRLWWvbnaoLWnuymI+tIgK9jxNCRJjaOCGPOF4L2WAtCPoFOZhC9bgmdDPswA
Cb0ByWXpa4hIsfyPfRkO2kSqYklesUV8Dx3ad2oyVYPQKwPajY2Xy3T0uz5YjAurMpdNiosNcuRJ
qMyTN0eGf1ChGkGiEQ2CkiwovG58L7RiXuMjZ88g7asYmv7s+HGtJ/TBaQNuFiVSLyExSoGE1sFm
8C8bS0l9NHesiRsMJSUMHxu4GnNzL4vWWuEox+tct+iVr450RXMm3akYsFm+dxHZc5e7HrhYBM+q
MQDTaMi4z85SmCkYJxLHqLifNeFtStLdE1mNocpcHIf4dYjOnUiGTw3BUDT8hKmg53SHMllBSARP
HiB+u3Zdff90KinLuk+Tay624IAcTxzqeOaWtSjCDQLHenSflSUHdS6YzZA0VG3rX9IrWDdswxfo
ysQsXnO337/Jw6a9u7u1PY0PGa2m+3DfUedc9d6Pl4r6/NNbcKDqSJccObxmyscVkjXnodeK9eQb
mr2hmQi/QG4r8Ux1dLqUu+xPAAlz6yyeThVmi0ooxYxVAwHCvUXRHuq6nLsShQ8tGmQ2ylJTYGrn
QWz+mMTorS7yPCCHgsY7UR8Ih/OPxwJ5Yid9iOxOAaC6YF6WDNCm/UEpGtMpEfOWeWjtOWp2y/Nv
QsAzv+MCwpiaI6AJ+gO2jWFoR8ldUF4yWfQHWGRbP9AFnhhq9wmDbN1O+wNsnQ3nmJvIzP/DYGp4
1t110psiuEWXsZEfyieoYB9s2HihkVevLK2PskW73Ad9HrM2FdwY9XH5YlQWxZolgbIElUwO+RCt
Wf2pF4fEZziYxYKPb6911upbk05pMHUEkM5amDEFBKH5AL5OfhGJoI9GQgfKjhwDTXZjRaaZcEES
4pSyVeOO6rJZtVS6S8XJdckyhmBgIATH+32b8z8aYibv8IxJSYoT24vl+8F7KENQgEXuRcfUxTPD
Kblw8snW08c0fj1QBk89vrJSM67XzHHufxLLUQXZZ88Vu0kPGjN3JVmAo3qIMM349IMtsdtZcXHo
L8x4S99AGiLTL1bSDJp0HwvLQnRgn6lPiL6Av/lI/fCpdfzpQM2Vu8y3Qd0Od59H/F1hhvQ54Qyx
Y9v/qjut7ufMzbeCPd6FXaE/uFPRjM5VxTv5AJUcrcsZRxgZQbuvSuJ5UlQImuakGLq7uWXZRdns
scEn3uSod5SOvYIKOPYnbMwxX4C1bq3/NHrqBesLNEPUsc36s6HB2UB2ismvOO7oEkrY0dtIOzq3
z3uDnYsO2jg82M3S+u+gS+90AdYpHtB7g/zb4W0yBH+l7qxHDqXnpaSTGUr4RsWzafXhLstuU0bc
GASpeaOnb1VoPelT5GKxe5ydoszqVqoNh9idZRWxo2ByTYLorwNSykfnYGD4VSEI83/j/8VXdrai
Lzn0xEMe2eCuVDkU1UFWJGiSuoECdTZJsrCtsiV1mVBSArvfzm9YBNW8iBrjHry9ZEA+WTY9AFFf
QtAuVYYwoKILnjr3/NYu4yw7QdGXssXgpov6sbFoklS9ecePOMoc5rOCLhNlBD3rd4md3IlVgt7E
pQ5Lexka0O6aPibFD3I8EHSttBMLeEHFF20c3dlPM7dvK7AEuh/CTysHSpaodwzxW436imygWhw8
elr025Yw6j9s0eFgBQ5c/cePYzUwfQP+klY6wTyctruAsMr+m8+1Pgfpkh1PdxOL9kpCK3CotxgK
bQKS4HdYzqiRdP6o2tK4ne4cX9iwZn6RX8i7JO9dnr3sB5gwfKZZ3Wyxj7+jDoyLVCB0c2QHgq2p
d+CkT+DePZxs3TzxQZZQWUFFTLhPNSVX4Y2VeVTWU21tgyF+zOZpaCgN3Ld8HQxlvUXP4/fvhj53
RDDR2ZfEDlGIZB/PLG1n7Xn4wkghJ8z+zJArBv2oWdsVyPj1tKp7a1j9BzzxxyCEzY9cz2OK/0qN
qzLVWIF0vXF7Z7FjnSjV5t9UYMp3lOE7pD2Er6AFCZvmdiDDh2lIkoHKWgYjcrgUs8UV9cxtgh9E
smOt4AAU/4b7S/NYpJ6Iy3K2M+j0dCmNd8QSnycJadX6JFKtVGhCQGyjUAy0vqmUjjuiSVjpStsN
PY1PNHcPSZnHLciz3lS567l1ucQzBeqhatYcWFPFyW1MSshnONQitQNqpQbu/yEKOOoaEE5mJXM6
BI6I88ieATmnBAuZexcQ4a2oeTHzbOCl3juY59/VSgFP8yTO0Kh99JzmvBQRWmpkzPJeR7TU2bR7
p6iSLpddCVPja6/qMsm5rHsW8DJzy/qYVQGJ4HPAHES2NpWe+9NUn5XdQJSfDRUg11hUm9ivBKOR
r3QTMg7+O+rrC+MDTpu2NtTf7q/I/MEzlQq6pebC4Q+hiTPkb76F/V67M7oZfJiqCKXN9bd3D0RE
7Yy4j7wQwuy4Ep60RWqrD90ocF/O7UXBBg8vWYs7TVZ0IfyJCKuSlSVUvrJPOmcLv4h2tmQIbOUE
MlF0sdpmlkwg0up93luf5cS6lNRDdPy93XJPS8UI7j26hxltNLVOK/nQO4fjVLZzTiKQU48E3F9e
He25QDHXrrhaRId5fIZ/BrByrNdfYVpDv7P5yevvUVjO6AAgbKnZTQ0TXfmvlGVT3iQpR7LnF/Av
b8ZERanW615KQwXc5CpRd3XP+ACZCfJPJUTS1EYA2YxphJ+YKewu3AhnV3v0BiA1pI6TonOCkDoa
UTGVitlKmAL5BmffNo4553XVQ3SLtaqrkkEcyJuUGGp/HBYN7ifsGHB0gO3IuQuvPw3cfif3+tsP
xWPH78/Y5sgbLBcbfFO11BRk8Ip1H+Qo9kmCzUrKmlffvYXHV/ojMjKGySf2Jqb95/TYjVbxj82D
F0xzESZL3X/RltxmWcgwViigzSO5C0dUN3OQVRLDTcRfUYtsd9JaY608g4ArByop++xYaUu8EzAj
91rOsfx9RHT82hqJSX2YYzleFnnrYHI07AC1JYrPJRO4aATmXNtmu68WLArl5tw1NG3SNaQmncM/
ggGrBx+Vgx9jWGsq9AbrLTCrQ1HFGhJv/gJ3Ynmp6jU8ZLK42tEWHPTpkhxkHOrUbx0OS1CFlSK4
MWBHLwj71kC4m7g6IV5SXCbMAxtFJOT/mIVmLhj/asySNHRYhHeM4Rf6BCROlAjtnen0YInPL8x0
9cdt8qD3VwB66W3w/dnw4Ox/Oe2u9J3XbyCy5lSkZMhYT+GIMw6jKv5996ueoK3kvI9q3vLQlNfe
6USnERYaaM235pIXVKLvyx8oKZhaAZA533mlg+Lkr7jHUoV4HMKbj9D7Jj/jUWBI0BunrTeQcoqU
DhfkLx5uSA1pP66MT8AxOO3LPv4SSuj6WLgPyy72UFToC4CNMDVlzKqMc7Sq0oDYXUrDX+yYddOi
6cKgjJ77bGzuIISxGQ0LPWEeR2oJnjWlGBJQuAGxdS8ovlUuyy1J2KZ3C7nPHrFpfvpkFCAMXr07
TdUCEk/iSG2vRgiPPzy6tAdSq5Hsac3X8WXIfaeyhfG6Qvm1qyebKVJ6FtoxxOO70sH2M18e75Uk
ZSfS8hxJMoTYuKr+OOridEPUgjBAK91fqMeFTUW1BDmQ34QP9LiPHLHgQizsbbyeOER0PNQ3KTyG
I0vt10+O2V4Atx8PitnavgJkVLDZw8niRQ/TO76/Jw9vK3CN1gxQGeBZQO5cmEb5VocYM3xjNPVM
edNyirEUcQ/2RdygBqwoiGLVNj89EWGjPaWAr7Fh7Q3Llq0Rrad1PIvfvje4HoinevCjKplkJTHm
QphFBAmsGpOjS37RD4Qo1rhEvgyOgY3bUzdCfZ5ASmuFXZaazW96D4/RiUJwRr42d9+6E7y8lM4d
ulUqgaSt9n92zig8hVoOiX7rPeulEdc/xS7dxyPdpcKNxAizthXcSnntQseSXF7dhAFm6NvBaaO5
kTn8kHt/AO4JGVQFxWfO/1MQJMszSxBqh4lJe0jEXfdQLqYCVtdae9N+zvzsdNAlXQ/8evJZxC92
JVEHN1VbRm7dxL1OHWRscfd/7yFhncwgZaqyx9Rsll67NzlLBc7wKmw58UWGhiQVgamTxNkptF14
irCeAUEwaJaHBeI8pY1bEwKbDQQyVXhPwk2rMqxP2mQssrNwFw1KqGupdmEOsD06CRO4IeVx4KId
WNXOraqXLbmvu7al7FtDysdQtC0ejZ2Um0IqmeVFlcf9r05vWKitiikILfwO+xsu+NI2BC2Fi6Xp
yyVMvesoX9CzPfuM8kz84LrmtvSsvu9UnefafY3b6a6SNjT4U8ssXepf5rqPSDk6QMUl0TZYmWt3
QWgwkAX9TvFP7Y3WtfLSfz0OJ4W5gijZu2GZn6jf2c6O3OMUc+baASnWKilXKtNMdJoQ5VnsLvIU
PfFRSdzHhg9Ahl4iakpfcr0IHfNqYzTXZbuzNOVNqfMGg2x2tHm7oIA1E0DvpgBuqQdKWfDaDyeV
bBx98pk1EBNLO01dFvrTxRE6ugcl8vuajhXbud6GGnA9VatCv7u6Pxh7mtKxRbouA60yTyVwUNDH
5ZUUmHwqaK4Jy7Qg8urF17RQJAfLw3nh4kNE+PeAFtncLds3B+0K9/V88r10I1dYhe3I0q6NiPhn
S08sAFzmK0nuwtPBO4cdpUY1BxMIRmOOYyvkNjvAPP5olAQj5PfJzKnxEqV27xkwXHpjh3rgDxd7
CrPhvWSCnCV9wB6sMn9EcwO9ibBRENPbSYrUceFwvs2l2U4GI9mh/tojbe9m1eOmxCWbYoZ0PrPY
oNY5l/bwh955PLaa4YdSp1p+fIylkOn0xkyz4groy5kcHB/S63pImRMCXlnyU2eakBL+6jb3LwtF
r2Dm0jJSFzZuLKzZSZJvTT5Z4E5qehOl+N3iGy3oauiQQhWJoT+oJ9WTE+qqbcI4w41GkQebYriM
3zXw7UdsNdvDHSXqzZ1m/FQowPPr0sVH1qkuyQB8v4Shsys9su0Y5Or9jaTHPm3FVoiHwGOb3zGn
ryRMVIwHKqMUcSKaX3tEEdfp4fnme/LB0BRMzSYw/6aPPqJTRb9VfyAOpHzh8Wg0LtE769ErHKqX
fIKNtXUthO9puTOvLO+zwyYgg6QWdkRCg+6lC/TNdFFEDVSLW+iENfFJnA/xi24iNLZlFsshcJ0C
CHSXu4OAQw3KPHw+jOM1YopQg+ECr4PyWwSaI3btNNhopQI1MUqK2DTE1JHHNYCCv1YbfwOjIANg
gjhy2SnBCIKquvl4NAyACs2ryeDIvaMljfE5h1w7O7VM4KJLvpWguk3SBBzc6FoXVLii7P/ccgvT
VyifLsmodS2yZvogAT+ayrc2+71WYWHx/Befg2BCNSYfvRc/gWGpWRBP8NV8uCkbCt2PTCJRtw1q
vVQU8T9KuDQAEnth5Vbp/5TqmqNwXmhw0cp3xl+qSxv8YomOMJkvxkl1m8ecVJEVTS8v1KzHNUR0
HA+7+kq4tJGPMbkz87NX/T0ilqu3rb5BVj+nRSBmIsACGJPiRY0H03dMcD+iP+mlj3V1T54puhO0
X9W0PpkgUHKoks3VBp5yxBL38OO8cBsg9+lj1P60uQidf1iLDF/YeZB2lgQoh1682czzGSP8ZWnH
h3pyMUMDrJSR5Dg3p2EOr29dxrwZ/6uCAF6YfWoSMp78MirYARpk8FqwrK6EkutprHv3YTsbp97c
z2x0nAmb+eEE+Qlz7wi9322X41sQBIituhlcICRPB4hrHZ422sI2L6ggDX7XMLI7Sdsfait8D4rs
eX22ZtvPPt8sEVhCINWW6DfiyfyF5nhwN2wjbc45vtmpeuEMhydhe2Ybyys4Qw3IVoojeMZu0sHD
/xB3tbr2rradDq5sokJltp+LLYXkXPn5/aWaaIalmk+PQ0KdT66hAgzIkMimcQehu9JCJ8pK2tDA
GZMc4O/io7+rxcEnAxM1zapDjEpNYF3OzzyzKhIb5SIV3aImnq3m7n3JS8lvB+L+iXmR1oOM64YO
BVEUCKiK+zO7LvVspI31DAStOtDy70WC3496WEqPHD1Ozxu/OJR5jzJUzMA842hjTYmOt1fg4E7E
jldlOYBdAmDm0G3N5E9lO+9dml5UrF4ewBHVsRPqbAnm2EGhY9f6E1yJaazWuqyFo9WQfrSEno49
KhlWjf3x4sE0p1LXjedQ+FEYSaXk/q9DzRhE2YLJ984rrpE+DIbSJAAEnSD8CX8Ayrm/QXmqvFof
w1xgjxDD2Pz2zKdK34k5UT8rmtIogH8u/PFMCIb+Z1itNUfb9VhxzePErC5XKhG/7a8YqGxcfYoX
EEXb0EQYKI+d1KyN/jXN+P6t3u1MtYpw4/VX5YiLTjqIcCpQdTp+NtsWy4VXIIPRWuEyKCG/+0rL
RoY91B9i/W9kx5Y+6agRPvDyJ3YNVBtVrhShOUnrlbHHt8FjqWDQOJJ4R/6IXao082ZI0Ryd33By
4KOod2WSjxx/BiYLaryx4d6Nu7Qtf354upGG6M2mXRMNpi56YP8pbPcXdrFS3gTfzT+KLorjxGKk
pP1jcO4KLzOXMYuIKcWZi9raxMY0dT4ygCmX6gigfWZ5TBxQNSWvnALsVbXTLJjiV4kP4fUTw121
4QWVetUT26+VbkByrdhwlu3tpfPz/KQ9a6mY88S6rVd7fi3F2SVEUlZ155OHZYpmzbBE6sm3Szzl
qOYSrX2DfRFSnrqlBichy3oGodHtPKpph5cfLYSpDhWCQvXMTL2hndMZVwoJ8QJgip0rus7cB5AA
u4qRsRIeDJ2s2/d2zJHWC5yOTOdOSqUc24cQFp9lZxbK63uhOfG+Zm+WR8NHYRC5T5Zge4NeoPYu
6F3px/78zgVbDcqe7tAMcMHYibSH65yVhU/QuUr9hmDMXjHTOOYd3s6I+syFnzD04Ju5g/XiTPpq
upPSOF3gr99WbGVDKs6q4aYWzMA/NegC9u2OOokrIOX3q6H2P6lh16aDEwXkAU9QPHOdRljn1Svj
k8fYxfCCWf1sEHrQ3h56cRrF8YNe3kezJenK7fiFKRlnORriPGQJiWL6vUjFK2egMEP05Ev/o/s0
CnIbUoUAIpOF42bF/B8b/5tjb0Fxv5OIR6k6y2+i5p+H8gsI7v4x54ToLE4dzSTW2X+yTMTp26RD
E8mCwN0DrfWnJjybulG/nzOtdovQPNUfpVFHHb9anYtZP33g0JmtDQ+yhauDoWipxXvEMU5jtFSi
NBuguQbxNiIA6SlkcUrRSqzVIIp1syXTWKCcma0cFj6aP3seV2CqK9DkhfjbjFLBdhvRH/LXl1Pt
PPz6bBP5l4qdz8cGu3thvqxyc9il07faqjltYCVPiqhoUz9iE2+EJ5Vzr3+is8ugRgHloLLFk1pw
JytlaTekLEcT+ma/mxr9yiQ/+hObHCgeeEl3Ovbmo/2obl02dRdQywugpMSZz0xwPc4vidYuwP1O
D+CJzmCkbX7a5x8T+HtOCMfthWMqx4y2+I16TCkSKE1nxNlhsffa67ero+bVl9fSDK+DhOJokb3K
4BxLno60l68DC5giUwe2mMmU0IyLzzjwlgCRijfG4YjPnqJcxd/p1IrB7xcwX+U8pyoqcbLkz+0w
WIZxOiU5UaWPITHVP24Ss9HT5T+bXq4cZuwVOE9q9DNeuteCmnC9dtZViat8QD2CjcvPfUDciaHA
6BENcUpMfLL9v1wXd1/4cGOk0TZse7puRrYh/BAziHazGcHmtICcG4ZfCr6ket+ckJn5Jb24s9xI
HFnC8nc9VEIAGiIsADkBejzSQVkTRbpKyRvN0EReqU4hnhw1Eg98q1YMVRML83ajmkSdY97V9iGt
TWFf+onWo2GJUkwxLpAKbALY5GPwYCDwU63vnNty+5iucg9A/dWXij+ct5CJCSwnarG2W7Sb7MYa
O6YY8LlEkefJGvyFEmnyFK6vcfNcszQ8dn9LCwpfXrXaSD6HTxOkKw5nHeSx7hWE6kVe2uXUAafJ
k+4gE7UdxCdvl4Ip+PPldm/n6RyUmUH0aebI3TrcjnIFSGTwPg2cArnAaBYy5CLEu097HzQ5NVqk
w3UimxjpCFsHoGkOlYtoaJQ4LRlENf48rs9UiBDyXkplIF0UI45PmG9NykaC2C2fFCftJBRz0tRQ
cqPRnRijeAQaNB/A5pXcfk/yDWVZJN0sR3yYuK5CzNWD/4gyiTL8DjaCqiNftt4/7XfWUc8zngRp
eYVJFEERSbphOBBEcbokOuXGa1nkLCynjrEdUFPPpMm1GYPty4VA9vFm3fx3GaaR1lA9tPbuPs20
yQfzWDIVodNeDE/XylKWQzEjJbAhsK3Ur32IIwYtWRxuv+XlOs2mtEGghLiZQwPm7T8xDROWLOeZ
M+B36PNZK9AOtPkkSJyZqU8sxl03LkrZJIEW3VUB9GbZeoe8W7knB/vPAtuK5Eh2rb4IxCPanLpR
LrcJvV2lEkS6srB3XwsIetOVD02lWGxyogiutpjE53vsaxlyEn9a3eviJZ/vICftxbYVrpT6nOfD
oPc5KuHnyEywki+EyftbIR2+VgcDFXyUp9VdAejZQ4Zihyzzl+8WsCNRjf+5+O8y0jfC2yFHjdBq
heSPU+ucqR8CHIPBI29hlwkRxLAAGu0o5k5885FLWGYQZXeDaROWW75jAIMghzJtftZYrM6Vynmm
GYV/03UJfxWNaqUx3CUUMao6h7Y6iVQ/9/JFboqSVMHVCHqq1mknK7JkCihm7R4oByhMr9cJLsxe
Z1RhDJLfZzAiVjKzVpr2BQJszkXjz59L4pScVBujrg6DZI6TqMSR4+5/CfTlc3aejqr07eK95cZz
N0J+1FPgf8feae8Of9z7xXYpS9tbGPfLoyXB77f015KIj6MIHGKTxO6VNoUZNR7GTxRPprTxf3xz
YHWjzpPgdw61TvXE5NEsyt9I5FwnrjnsOsqvzLgcfxmwzoKpuLq+fjlvqVSaltHZmcSH58eOM4/q
/267uFoLLQgBeH57R5Uxa9X7PJCFWv3S3j7fkWJeHreSVwK3WzOxxgVTz5pYhVWKI+HxXmLy+2n6
hfWjcJQKuAeHmfqJsN4KnnB9ISxOtrz9SsDUH52oJ4wXXdS2dMceSbOSxhWAjOixUao4j44w7ww1
6A8vaVR1r3AgoQ2fPqf3m31S0RMQAOnURjzh3RdqLKhg6D7YBi+7TVoIHntznsGmTl2G2RmOys03
2audHALQQ7PEMZFDSYmoG2SBa/6lRCVYX9Hcq2fMjH5OaP395ydZLZPYPlNo5gS5eoDlvv2DdnJ4
Gs7TBW6WRUI50pJjgVM4RVi2MEu2n5xuMKom1Ng1qnfv+vXIiK5G8lolWRLfNnYahtqKk9TYn/oi
qysfRXl/bz6YN/UOHTWPgixxQV+FmdSJsVDa62RDlX+2lWAzuuM3FGAPykOy7CCPkcTP6PwZHoRl
FNaaGIYeFZ3qs9WE2MnanMzavuUHi8Knj1vVPX+619Lw8cMO6gEh3N5pGfY6Ab8tGbxzohnR71oJ
RorKFztdZ+SPEpES4lYUEkZzG65uZXPVSnQS6nHOnpDRvFQNKybAjohn4eMAPf7i1SCVQGKNLG5a
eh9OCY850v8OUtmcAeQp38Yp1el/eVvvZbhPSnUfkYJ6GyB/vT98LIHdPhvuQJ94jXlLloV4+oUL
1D23mTMOWpcbe5UW262HEzE8h8ty3NohW//WidT5d5rTsNtlxKu46eY8CHVpYazcmU7MtePPTXq9
mKEDJxDpNqn+1A8AEg7UogPP8YwIkC/C0zWy1rk1JszPIpdh+tbwXdD6mgEdZmO/fdqqPpXb8jIu
x4ENhT/HgXIqSYwNDEICNfNRVcxVBc/wdDoSgE2G03INbzB/BK7UlWs+RkArvOxa0YScgdQDZfA+
EwpKUHp1mVDxPYY9Wxnz4CH64HncCcNYxqW4iMEF8znciplzsL6sPAOKEjoskG+GKythSr8awxcj
XBmVNkXllaGE2zM+AK+KLDezWfzEVOY3UUBHKBg9C9y7XR6sKiU1SjBJT6FrRXeH4qf4Rkk4WHO7
Wi5Bx8e1UEkikpzf3dUjrQkCfBN65Ig1wO/2nBCitpzCEhGxj5xlj48MmnQWDLUHgGojenZIjch1
URIV6n7MnVMtAw47Qmb7Y6/e4PKsWL7lKN9cMM0uCYaUXxAYh4vKfUb8F5WPsVZjsfzgHvpFhM+n
wFPGua9wnPIhfw4GFnWx8CdgUD9Ld+q1N0g0RnmzFHdKSeE1WhYefGfyJ8hkOBU0VqZWE82CG+Te
2vFVzInapuqJNNhQsL51uU6dvXJGrTBHCW8PztqoDewv9Ft+h9fnfpXvKGGSp+qzZGV3fhd4FL/D
xGmUc2vQEHepyPJ/0B+fAWCksUEHmpbNZ4+6BxWOKDb1uS9Yn6JHZOYvGEKRGG+HDqNagG02F3KZ
3vXOXPVeWyZ9DtDw34V7uuKSWm9FAqEDCrtAiu1MN6VVbmouyah2U9VYgbgmsuhj7vjgS39lfEeM
IerHhdJnz8TVlQT7DmLV0JAMUfZQ2LOm7n32JtvpKUIdYUfWiSRjpV1EsDID1AxnWzenGTgS3JMu
ba7MQe1z9yTC5EUc8jQV9KVmprxAXsKUDsmUH0fpQz0btHd/9QobpTUKhWNcXceBlAL8ZKdb7rhA
cobpzjVJH9TxgL5ytxoIO5/4cuWTOkzffTDnMmXEbExUmIVSP/huxgujLtFPGDq47P/YE0cc5FKC
PpAa+QpK2e7t6z8xfivFJ1SE5068OY9PoUOBYUjLoo9n0EOdyvJEDZms7qnQV9pefyj7E91MX20X
QHqapt01sIO+pULRHNWwNkC0XADdgxV2bdyjzGN3drk+7YiLj3N0cMpYlQ98FgV7m6Uq/8I6vTKn
aOJtFKTNklWSu2VOg1Z2k5V1RxJdVrLGis2XB2ajzRhI+VeDRdjcJy8sq4LWmirWE/48Qgm3YHu8
Q/nqHZeKPiMHvd3ZnFClmzn2aS0w6R+TFTp9c3HIJ6F6UQcmMQGFu7cVSqgFRf3Qg79Tpnx8zdt4
OEKzOqe9cz4cmueDdvS88t4iutJ4YmWi63fQ0+yCh1ge1+9X4XHUV6PMIPx7X0PeTtsdKVlCeRJV
DyFfNj10d4u9qKvYqXqGiuJztSndTf9j7Df4IaSQL3Dd2FHm/eA/A7EAGmVTbjBUOMSK1KoPNOTB
zEgLo2uFbBDUE5hUt/ok2KhLfRHAbZyFE7WD3C1z7LkCTfS3ukFFMYvoPIipgv7uRfiDQKMeocFj
Tfp2j6OCW906SLEoIKE5nez4NY6MLE55Ue71Z8y2xB+kRImhCVxJKqOM50/25a1giOrZIZzixefm
FecjKm7IyjFuA44nd6Kg+Q3dkdbMcKL5sdLszpY6ubOYKm+1sWXq69D7yCTBEfkxzTrIU7iZ10l6
nNZQt9INSuTIBNQsnVr846yJ7s7UrsqDhcLWI5Z3aVD1fGsi5tbTPMGBjmFR9/B/Tp22EKxGoggT
DVB+H8wn3LzXPGsYbb4siAOLPh5d5BBr3GzmcveNdnktABKqrTnrLCEXoJrFh3vxBFGBn/K5WgZW
GG58huvgW0lahUBu91POxmIwwVhbC8Oh6sJNGtfENJ+HCwIDqoMt053ng7WUVq3jagqBy2tPbHH0
Kl3Ll3Snj3xew3X4qHRopRD3aj4/EVUvWDj6zrMYZjUcEasFQLZ0uukvhJ9uUUOhhl1ftjbUlDlF
DhtZNbfKuHNhxp7oGCSjBVTzD6KnyqB0QaCmoRnr5qSQtRK9GH4qaiqXlohzhTgGFA5vjm5cM2DH
taDlbk4CTUXZM1J44PyjuGA8mfhyy6Irr+ZG4Id5VkBEJcqCyTQ968VSRyKbk0qV7ABMr+84erOf
KbpgfK+b8FnyXtV4yXjwUTJa+e18ICeR5lFheShf+Yoq8DZ+IZFIjBOQSRxs0c3wmGYNF8YBqzpD
jY6uiuptZZACQae97A3w4gYdkrNqSBjkhgLml8HCsswEn9SiG7Pk540V8UWUqX4T0G9XHoGUiHbz
EE/9nLAUDVrnXYwvEf/37vRD8ecUYRwXHvTwXK0cr19jXySjlZj8uqdQk2YvHXcKHJkw763GtaLL
HgeaYFSuYSF7g6ZJ/7jOXluXMORCB6uvbjMWvKdC2jyF7YZFEmieMY16d1PZMJ58GTM4iyMU/Nhi
qUre2H7Zif6PI5BTILufA1W2AehzVt8Hzkaa3FM7l3EiOS6Qw0NXiYtkOSHI7bFqQzNt65YBLbJS
7AoZdtRkQ/JeAElc9IT7GaUlYpCYSIY0CkuXPtkWULbuxNObTrcN8EDGVl5vESktT43vkSRBGwX1
WdY8l1HtrLNFxCKy3zHAzaQwrn2AxoVvRmx9fyAf0KNZM7JfYWymoQkY5kJ4q83JVIBWMfDJr4Rb
Gj3JcJHO2RCLbG9mfX+KopRsq9SO6WH8xMeUl/lPy/DFdZ2Iw+zRp3zXdO2SMoNFGkMpuHNFLg+B
lvL+4WTWKLra+1QMJFg9Paa5T7yHy1rHMdp5a5CoNZwNuOGpDu8PZRocEK6g4uRYIjEGPrGTLD7y
PHinffKZBX0xACH3HBfIqjqEpLKJtQorbgbsUztw+htMXSLcWOmDAHrFXcboxDswDA4Hr2ecTkkF
ANrbxp94xrhdVZ6tbXaysTSsyXJmL6Rq+ssRPiJruCM8RGyWtpox7Xahruyh/ihfh+aTlAZgeBKe
l2I2gqwebg9DDprho0gEHNZBWxYvMBkYdJB76h2OdJ7mRALjvzEOhVIIuAG/Sc6V9vK/UnXx0WWe
nybLMY2Z2jEnteeSIZz9hmyEEVKUVvFGD8FfXatS9E+JBK0I2fjY3oLHVBe7+aar4WRapmTOQQM7
RmbAbiHcp+V3ItbBcBEcvhUrJkWrbzTFYTk0kWp7wjpjzg4PgaD+f032HtNoqjD9sTYZtbcfiSuk
l87/JvDqx1FILqmfaVKQk/Ha04igT+52LCI5e/PUnpA6hePuLejOpmBl5J/yYME4UDQgEiTxAidB
ANzKpf3iU5EmTNx7qBIS5facBJ1TtAv6h5Rtow17ZTjA7i6p/Uba4DYCBHCFKRVbT7jakiHgHiYl
WkJFy31Wt9h5Mb0Hq87nWOsLaY1FTmIqtBEfYQPiPX6Br1cVbikTzA5stgWfJK5XNm8PI0bk5N2x
9uj+qRUUqIeK+5rrrPVsqij2c31JPtYDPgzFVeZcizWIy4oNVAf++Nci+9ao9yEFj9YNj6QeJwiA
NWuJY/OxShWiAuXKa6h1jCNJ70jaCFNe70voqVKOeNf0477NIk3tA8x/xblQsbSGu69P5PB+5Vty
HSAsPsTuGF40t13MUHKha7Nr+iPw10esIrR5itfXXywQbujdTHzZTiHBN/iIMr6Y+vhgqbFYDwF2
j92w2HUOit8ZWV3+o1flaKUC4r4ooVNVKAYI1iwc3IqRA7iatVfpVMLQ/XLnIf/WugafJxDFAb5W
KT7lAxj47pTzi9wKSGBbSEfjt3NaV9Fv/2jn8PgLriIHv1IRoLOJu4AdRrFGoz1OKsdgSF4GqLqw
qUqpN3CfGVFjIU1WIGiXhjined0mCWSttfUysxfmEI/lMPGTBdLBDXTHwsgD9Tif42IJDm5DW5l0
0y8F9o1R0PzD1ma4QFQ4RY3CSIW8cC+dFVJKDqzr0awB2Q7sMNWlzQ3no7XaNnhKIDNpdGxf+ywy
wwvvNVZES2IpgLvLIrBz37RwB4I3OtMmSU3txJY8a5lDD6CyPIiEsB9U69ROB2z1HhKFgdUM81IG
cRQ/FhzwRIrFlm+QtNAh4p3vTPnAM2Q3+uOWc9xqP3KpHYpQEoJl1JkVVk8p7fYGpoY9YEyWS5h8
OF1S6MNASNKtnJkLBh7QjMf3dzSeV88uGBNsdTxklPiBBYQLcCitg74rnu0PdCSfwQtB3Qgx6qpr
PgZ2UdGNMrhYm1/210YGo+CzWm5E2mijqzrmJU9UAZt5NdGS+ugG+9CANjKgMgP1qeOU9tmBQgkz
uzkNf6brRoVvd/28qN5NBktW12FIsqFYd7ypdX3D5Fl3qUs26f/IRVfSx70n4Mv5PdK0V5JxFnwu
37v8wwKl3AeNBCKA4i4O8L0CFEoDF1ZDAnfn03aS7S2oYn5W9msBTy1Ts3wtLQFir/yUJtM/ygtr
TU2mZvFV/w67slxgSad0Pv2l66H1Ha0OIwCIXwXib/cwWVWHRlgGijGjCmAAOQdVPZRc9rgNzH/7
U5drtCLY+dMfAe045kS3qicfjZvVAf0mgvqaaZ2gwR9A6fUXIdmFszQVW7qxQgK3ON8qVkWiUUEd
VVJD37RLul/zHDysXUl6Lp2SCu5Xkt2B+xNvnyEp0xLbKdqn3ZEMmtk56255/ihW67Yc95B8K2Ge
jJdKuNfAKAv0EDPABnNaDPPhBN50RbyVjNl5ffB9y9aeoAAJ9y+Z6jfwSwWSs/f37YGhWRqKJ0SM
1yndThWkMoc8CLr8QhImMgRylLFGWJzR47QX3Y+ZkxZ8AsXyS9S7jSpU8k20WwJoLZFOwD46zSOk
BAlqQ19qrprN9c7Z9zZpXo/7FQp6cZnGD4+QvFmyZBBJ9EDM4xq7FtbJt0reXcR4aZSfyKX8M0W0
Mesag66vUQQfEqRUxKfPUrVWEbYN6RcrA/zPkOrsiTih37qvdOwLzQ6vSmXdJ0kZgzZWx5YDpaRX
HALuMed6ysHPvyMUF1F7NPY8HFREBl2/HvZYevVccndMPS6nQaHmyf4oQgkw97W7MdjS7QgEfhE5
n/rvR2nuWGSFU9Nf7tMLEg8+wsS7xAhwjpUx5mRe1nhLC8OkGYL3aCaXvCfw9ArwDus9o4ncvyJe
uzwMU1ACh71tb0qoVy1txdbZDtmuqinNqE7pn6+J8Gfr7W8EyOMIXLmGS69oLzLkV5gYrqfvcn7G
sWstT8vgiRPFvYeW+ikw1rcpCcjumHP6EhRFo2+p79G8oJApS1ehCt/k/ubBqHbo8nYfehNLY80h
YMlViNXFcxcBnOvgxxVfUoI3+C3qPqcg6BdokNqaScdcrQNG+42Q38G717ojcM03K/1rdUBvUmEZ
GlAbfZbQkwoXYFC/P8DIIDnGmVoJKFbMO9+uJvvyyLBFJWp33ZLAgWq9qMcHTKVinHwvmcfoVq5I
KVabZaLEe2z+JkND6dKLUF8BUY8Qdxt4VTGpM7C7SDHSiZTrinKxOjj7LXIY/1zfP1mW4V7UcwGE
xpKMvDgonkutgfKtOU9qegkqu6EGH/3xmtpIGvWtJuKiZQO9BTSgTws10G9Znj/my0Raaqve49Vh
/zZvpiVdxpeJlM0iI+GRDgthtQGOcl0H98yAFCGfyrMgGkpOSxnJgS3NPTJkDxHJfvsXblghbJUw
yaD/ueraM7a09odnZyWlu25ZEpJ6H2IiS81I28D3hyTgTaCzSD7LgkOHo/QdOp/LniB5dRByq1BV
Plnjm98c6hVE95KTherRFLrBZyLvsbIQT518bUzzpRG7ZAXKOkBq48ouFfhE1ulB8uA7ebEWOgIk
oHnoG7m3LeAaXeevMz7iHxxj3tW0W7gSsQ75K+ThqGP0ictRW6RTIJHx09J3M6IQW4muHwDY6SK4
7i/5uBXL63uAANbEwQSrKmMEaqjPdOZR31mG0vbNCgMGxzMnBczKS2RomBs8855TOKj16fgKxDSE
FM6fAagfJ1hw5JrjSOsMLg7OvlU8OTimx2jePP0LJEsv4bWVYVjyaW96mG0Qrl3AyyKcF3GWx+K7
VA9Ig4W5dG+JPxeb8eUKXs0GzXh1ZJmeFKRzKWb9oPfChHlI2sPMB+n5T3icQlaYaijw+aGNye9T
4J7pTaqhmrTYoL109ffERpNICSEzQEnz7yYFjb/JsViV89PRyAU6VZBMWXNEuPSAPo48CZ9yWfuJ
wLdMNICleiHajkd2jXOZTqoo7o95j6dP48+mtFUi2nZPQyM2+EO4MnfhS7DcdES1TIZQgE53FxPf
YtuLPiyqDfSvAFNfpExDtCp8zqGl1t3Ti8cUYq6KNuUVxVc+UmaTvpwZzVfijL4AccEB8EVvo6B+
ap/0rGwoVy6sd0js3GrONyqi7ntD03eddOt/l5jMdEE8ssRGxivwAGEqabdSNl7Bp7L3jctVKXu8
UP+06O3RoYjCz7p+sc1YH/xFBTaFnqcWdcYEbIMDNBdeWVAOR2FSyyh7+ePl0Nd+vzfTSxo+0iDY
4nXzu6QmUF2PRqzmjFuuNSMrPRPcwZNbmSoNWRnFAJwOJLzBr8SmKqvcxlEhz0a8G0qKT3p+htY9
BVusv9bEzmHt8CmHi9ZaDI8eKf3i8NnWRNYBjPeeWzZyHSinzfjkh1FGQsS19Rr0XGzseftCh3zM
zEc3Gmu5I/Hz4kS3kbYeVvLpqUwdgn4Y4o+540hEQMdBKKzbDzpkjRUcwucOoa6kHpcJb2nECJwV
v4M7xfKSJ8MrUmozUYGu9r8RzUyuRgfGotNAmUC0vQhtDaZ7ggMwJHiqyzGKN8PE+eFzsOjwPXM+
RvIrLjFhYyMO2aoeQd5xlGZ7t1+wbN/cqux+F5gmkTxYKve05NIjURgvhad/JmiZuJneG+QT4vnb
B1xLpT+aI8Hzrz1KpPgcPQQ+D+WYskvdlhzOQETLQB7vyj3ye8TToECODkGJEBXbkP2fVqof/IUm
baFERvNXorBjKq6mOWjT9vv/S7ajKqmmdeLrTKfB4akCbixVbLhu9N3p2Sw/YDClFy7cWiHG48p8
icUEuS/6llFK8JCK0sv6jeJAcqEilzuubS6Q9g1TcurLHccsaTSB+Uk0ox3PAYaI3w/UccgU0STE
sfXMXzo8ZhuToDH9//2lXDhnSJ6FlJYyaGmcQty5OpkzWSjk0ZV884wltQhelfetdZrkMi94NkN9
6XtffTz8YaDeMXrSVp2m+Aj8UPU1hgK5HQBqYhlI5KWlyk+GX1fL4vPiSJA2Nq8QNnnFIzYnn6mk
p6rt4K1rpbNg2EA0cKtlragSq/wAXcBge3bzTdXa6a0KdQIWwss1Ibr5pTBGZqQcNF1A32Ql8EBc
ysg849C13o+eZFI3tJNZN9xPz2HLm7gQZroVWFqMIO1OBcZ2KNRKduazYmfWZ+LE0i5VJVr/S+ZC
8zD1ImaqFG4i4uggKHFp9V0Hpi/qbeFt2KhQFuPZ5NazjDmQUfbvaJQLsoFw7HwpY9Z30zEt2KCZ
s+PAfkO7LnuLLbbEf4RdMzgvPl6lOJxJCDAhFNWb9YRIqZrjiQGVRZBH03De5P4zIzvz7XIF/+Ct
oEKCI7RRA3yhx6/yi+FK463WEig6tsvngxr1hbc/rLN7QHvPrQyqLHKirEJ6LJreqIbe8HcY/Bs/
nYh4C13w3eMFmjZQmgGeHoWqPoTXpZnGgADSQhuxySh1nhNsumLRfpgMaqZYOcw+Zo7x4+aRXCuv
wtysuTKYDWCaQTcaxzdYpKLFjmdyep2cJHGy3Nd2hMKaNnfWRPqd3ndrd+NeO9zcWCYIcJ7Cz9uf
/SglDje1bnFaf2eOYPXdiAofmckuko/q6Tk8StoZt2bzKOdEBkZ5R+RBFXhhfE0oXdnFeuR6ZzGw
VYQKF2VGjPSK3MPd/U473oFnBtsmZ1OWcciIth8I4+tGYjHlzSWT8q6dCOR1MS4ws/6mwQNQk6B+
l0vvSo199S4Gyl3cENxIBgtGVMXIjkQTK205y+ULQkaihrKJAXwNO+n8vaGhLrPSH+pJtR8zeU4v
Vrz6ecs4TeKv4Vme13XmP0TYTnvNUkqbXrHXnEjfOYT1kwEF0Ewamwi0h0Hd2ol7xb6U0bAOr1J2
OawrA992EjEXS+3zxhvwRulaGr4r8WcHWyT/fO7tqrGpj2+DmUPhvmGC5Bfkoo+bsnLRs6h5mBlH
Y/NkeRXJi9rBvZFiAowP9qYBYz5qKMhxm3P1pzhsXccTl5b2lDOkleCLPLj9Jy0gG15i4S1kl8BU
3EW+qEuzltWCLta1jAPTVSo13rqaPkxu8HC8ezMXJvJGbIp4GPcNJw5PMtazlhMA0Je2t07rK0oN
6HTejkFfphwltILGEJeBb489paYr7BT/wF4ubRS2EMDk4i3nl9dN9QTHjfN3ybqIIjT7BQuz3fmd
+tR2D60by4F9AgpXYbVrE2Y9sYwRSNFTBu5tzsXj3Wbw3GAQT2dSiOYYq07kszx2ooLzIuNKOc6n
rXwgBdf1SxDcz4Kwdx2AiduEEN/QY5Wws2wyVQOqNSTXKZW0z5KewVrMn7of9j88hMINz90fR+O7
LrwZo6EXEbYP4JX0cN0EY3qGUn9qjvzoiV/SbURPyyqj48D0c6YHpB9vMUyUTKOoVOOL/lKaNAwX
I3kEn6Haq7PmxH7vGjv7JaN8jdqgNxySTcJLKIb1x3dnLW+XNiFE3Y4feQTUF6ARxwZ7anZRzg9Y
gecfkPShcCfn9fGG6vEwklnpAU/pWOkBOdDED0Sn94qzXHG9dWVvm2ENqBOYGSipe/B45RCCYa34
2AEEKphQYhtJ2m9XQs3gQ76WOIzcRMNLg1h8n/+O6nHhe3R1fx5FOgmCP3oo3HYoiwYZ1DTUyzGW
XJrae6HMF8sLj/YgbpKC6VUvVO/2TNzW4Q+TBHoqTlgaX4CYHZdqHiX8qW41BdWQ1BY8pB/duhqZ
iLn8lYoHSUeHMNsS0GqlZEtTQBbxOPQCcPA2xdf6KTEj53XdEtlxt6q/tBE5ofsssbJx7KmrD07o
3Z/CyMHeDhcrLDtiuK7KDaJwLWewQGgqZM4qzZlTkQ11PU9hiEo/GHlqOV1cmyveR1nzvSZjb4/U
p5J4pXhmvTZtG1+p9sUlSFSXNdCi3LhIShNoMWtELvA8l5VefAJoPdhsp3Oc9VXqczcqh8OiLieO
0FRphDZMkENbrc7Dk+r/udgyA1OjUsLwMbAbU0ALHlIPZaJmx++Gyjlteb1txHmfqTfkrTecqtVg
g7/1+mk6zE+H38bWvRuTKQZoIsyHBfkgL22AjYx95DVTXOnJc6wndrR2/8+IMS5qTAq2pD5wTJO2
XRi1CaYyQwKpLmjLGLUJLtCCXOuZyMn7QaVw9F8PGXkANtkqKmnljsdLtlaJuNF/ILDuzkvHJADq
AR4XQ+RHhY1QTLsvORiVrSnF9jPph+rdEHOKTqGQ0MzibOpzOFJqGsIMhakxLvf3da/3MyrYLQGp
7BwYa0VzIS//kX9pvPKnWIy+0NbA8D2+hZVAk9xaqo6aMOCWN53uP749xNGr3CsmbefzhHQWQe3J
kxXEBDFziP5C72brZ12atxIqmOl8YeG0nFxol43r2ylZ+t+9aE1g9nUy8YvJugkntt5l0wfshvun
IL9ftiVqPpDTJeSAHDpjcuXIfJHJZRB09cHjTsktUByUOFlXIyDxG/1GROyvIohciBGdLc7LNblj
fISirEy4Lbnbw3Wsa+4BoMOakNcXAIUc3P4X1T0yu9bX3Tb8ES8z9mMEvKMaT2zwJOYokwhb17Gn
iPGrG1MxesexFuwaFmHaq7HWtTZB+cKF9LpkkLfSrRxmO+WCrOavQ57JNtjUyeMfylheEFr9Holz
VeWH0psNUqChjmEKIhNVM51sZIApvqFNPNYFV5jabc0zwv2xoRCgkxUPNZ5nEeAttDKgxlHYlCtR
xezDwhp6NT/E+KY/xXHu87R9L7k78IcffWCe2vAGPrzRaByI/3hfV52tLzneEAdSmtgVwma0UhM4
7jfP03FK0jesnO0PGC77NTNaT3OQyr0FXdHUfVDG9jzobDt8v0VlTOtTmI9aqiwWqLQatNUL6WqV
ehVwakhaRNJD2fXO/1jfB6mFPAmxH8/VIhoUe959zfK2nkkjr2v8G3PdvC2M4eJ4TbZFuXi4c5Zj
dd1uBEpoNx87vw0NycQhqZLn0k3in4XdCuKvLNZ5tqvGEYpZJ9zryFuWEdpjTkl9IcA3UZ91Puix
rEyAT+Iud0lK6YwybOeg5dwRoTu18K/FRhjiMDXUyNfrPaAuQB0nrMqHtYogfnNxffacDfT36dK8
QciWm8YyZ62MqoBF2msYvcmIesel5lnscqYQNt+M9EjnfT4OIVGcGf+SsPXY9E5ppCx6q3RN594B
ASAd8FtcruU1tNjJ2DEp5KgG72/GIh8aLpStY2KkVVc4t31UKvIADf1i2BUzNpbn1HxL2zZ1xgMW
ko0mJUR5zFpnm3Vk1pEuGt3ou8W3McUiWNcgzQ00evL4C1v9F2NlI3+TB9avVx6XGuCtnTWitQ8M
rRzmoDX2VBwo3I7rmmcJVvC/8b1zzGRcOVXRM49DX/HXF44ny0qX3SwpzcWIcWU/g6bxsam7ZaUS
kUan6g6ov/ZefXgyrfBUqYt/tQmLZ8/I5nz3jcywo2KH/bI+LfIuwKvbxf+GTrgCBH96+KJjdjls
/83jWD/rsdhuUjL3S5c6tPV2ciZvBPUyzpuzJNr9vGXqNPdEC8L/8T6d/OO9khUkX9+yUMpIvj0V
tXGZT7OXQbi3CTpShziTDLE3Ac4S/hqX0VYTY9AUbZdsTsXeZxfd30xjTVS/2JDGJWWP3ZuvU8XU
fk9drlc+mksaYShKiqX2kErecC6EG1cqJIKQPm2fPZaNJX7f9IApF1+vkya6MzgY4rksukvC7W/u
W5WD9zYVmWgnfHq47jcTuF3hjd9PdenhHI34xwTBIfbtJinbcnUq34/NJfdgSBhhBMUlbaWt9QgO
/46FfHMUEjA5WRESgLy+L4m5dE9EVGg21KDNEDQM451N41Uf1Jx4DD91HTx6lNDszrbJkhbX8f6x
NvrPrbIzjMicIVT3cLk7n8LV27Z07HxwRr0stAzZyOB/65fyxdLa3Fvv6z9o76az2uGJMkbsFrzX
mxcaHzk9lc8pmEnsxcAQHSNO6e+IXJpDZjG9+88+XL+DQw4AIm1M6tCohGP97zLm8mJuj6JR9sDQ
UiK50QDWt9DMV++NcuIzM/UgMokBW9Ra2SHl7atLeUf3rxPlRZxJc71X2y/0Q+KUFafn6tqa/Y6Q
az6f2o23sQGVtNnzrP6fhLJUxC1iC9PLmJ0VhlxJVn54IL+DD1BP8StqH9CjKokLFvs/yCdqLtN9
sYJ3jCeJmaHWw3HiH2VjXepcey1mg/n7SVGPJk++lNWcxBgqrQ9WxBINOSq6gRHuiPIbjzHg2YDF
J+xP0wL8zEs+OpyFqrt/AadHaoUCoh95JFMEUS7KrME3H4RpO4twUk2NvPt/oDd/cxBUCzG6QY/5
RcFLbDSZVH1QPbp+vldRZT5M+gupfbt7ThnmnNy+RJ/vTuRHE1lOHXN6cpAsfHj/ZVKNJgfNnJXy
aak4oF2/hpuxx/Co2vmP1iHAQyBS2ap5Q5h5x24M5X1RzNu+ayWDMbckebK6JvTibu03BLaLpMrN
TRvUdxzmoDBrBrgEqMhzDYJKUq+t/xsL/Ui2NjHbjzUYeNzI+Szk7TNDfZRwj4eSl9vWWDsrEtYZ
bjuZj5c0/KhRzMgBeOyvP/QtxyZdJBg/dRc16Ij5IQZhShnvGh8dbbtoRgxPN1p7p+jdiTh8eOf6
o+MyEmOvmXp5qy0x0lgVoicG3TFGY6DUPk0QNTJ3xB4XNXnBVxik0O1DLDQEy1I1l6TiTEfX7BAp
5jPJWsrBPyfrIB5HEZmbyF2FgvdfuSWE5Ykh2Fx2JDT6ywyGgOUfTy7R8Yb+oa7unYZ8JMO+jyFI
WgXaxt23ZZ5Ys11zIyN3i92ARoSDUaaM5IbclOMFOaZxceVV2c3Td44xwwRXu8T5IO1asJizl8Pb
+GvWUfVxLSRS9/tisLL68uTla0LoXYVxx1IOqCHeJwcpZKPjwJlRphc4GVpaYxqybI98kZabr9+t
udNSGuaes9erw3+U8wsNPbVzEeRg1737L4r8o/BRVhGj+qHKIrxlpbiNFRWN0u2NWwNpk/ftUe6w
6sPecx+ZNe+xRsoxSiocpdxX05Nq7k3mzzw76lEGfsBMY61G97w3L7Ma1imtXK56y0ZYSCPvPYQG
xeZsURwV4NEvlbEc8OBiuBosBuPoSPbDzVyzUuf5CCHAOZnX9m0v0brycSRlcCpWiVywIC3Xh4IA
New3pKIGd3Bd/efJOgTUJwxlGCgeBVRhaaRepY3aqiq6RwhgNRRp+T1T7OEGNhl0PFw4KODAPKAk
i3VjkyL8tJCjn36w3267CfikId8XyvdCKQia/Ipe4w8oL97AFcs1j1jsaYN+XkQsTY+jcCnkMSGH
Ozt21nfehpBahi8rKR1t6V3nFk5/3oaEIUK+C4M80vdIofd48I974I9E8Qtw+JD0SV80TOLDbVGh
pWZvkPMecmLZE9mgO5RJVaafLxYP9dqRDqxUEmsJvW/JTB8oZ1ES6t2+UVZFq/76EdpIVYFPNuAT
xFZph2BdpRAUi18mpNi31tIX+9/foMflGhWyUGm7LWUFQRC3ItSpxzuvN/08Y2YgWfB+rnoMTxbv
So5hNIaQkncMh/zWB88sNzyJI7Sk6PMmCCOqIDH3DpMbOkVZ5Q5IJ3nDDyriHeN7WH6bxpqX236E
rgt4neBJSxrRmsz2s6OWa/sJFhtPVJnUtXacKNkuVBvgT1eEqZNkW2kqnlgcK1JyHtS9zlVFiMaS
omz+npkjyolZSI3zultQcIHhyjOs8A4OrRSLPcNRPce341a5oHDKVEWSiCUfcu+1DS7TgJl8BEZ0
c+c136Ua3rf7WQASceTTCuocAZIv3PPM+SqeXwKGyIgwsFcV2qtNiTm9FjT7vU4tpcfSlljkDj/r
g3RqevGUvU7it6yHOFeirD7azr+YWspk6CLFjKlJ9BqY/8MFHJrp+BuOyV7RbwgRDUgn9d3PLcoS
S1qhB4S2/ELMgkmdwIBA0In27N0+JjvXlxgtaehzwfpgkrOkCFW3l7K4ROH+A61UgeTgW1jZq+/9
HNK93TlZUey+PhioXRnVY0HWTzCvOZKoHQyRxPLpzWbyCXch/hks+JXGoR7eh7PLLhwSwDzItMJA
p/uKeN+boKSrV8MTK8hi9hvuSHeACWwT+wzBXYJq2hbeSag8ERamlkjMHV9cIYmoXbh+1uA6Y2fI
ULKjou88aYDOHVgZir8yULqv8WxhFWlRVGaXwyj6bGk+6tW0SeQvyeaTLpOPMYhYTu9m0MFkuXYS
1y6eHZjm4GkXSvWRJDYVgyyIrLiEopKUDrDT5tBV6PPhZjOQz6EglhVMluzNBQrB+XRItGQxOL+t
iCwdSaZqwZHy9iEyEaE7rx/uPWFZLpnA5lCa7XgmsJm0+d5oPDs5S+qRC8ehgAkqY0I8nKfPfUY6
Tu5REzTZLZUa4sj+kQTQ4BftoQnrBNii7j3Ij0DMFiFmfAdewvFK7csNjPfUuM1Mvn/beyX5t2fN
HAdM2D5hdFsBBMfhhTcJq2IQ3j/pGKsRburuZtdGdDH7z+EGcbZNsdAW9AiD13GrNgOXQgeUkcOp
4OPNmCoswHJH46JD5gK/au7zyeOskPyaZqgLd7FGSPkjWfiEHnMeaxrMIBzG96a2285dy38UDYTE
QpS2SH8c3RN8AYk7eeVDMfTU5D3yBBpuoOfyPd10elqp+Ny/CPCdeZERf+xNjTyWjnkrAIPwu5Qm
vJQL/8627A+MDDw7btoNameBmvmN+YLyDUyUpScwGcJrSrzh3ZAHtW30ET0DD+Rorebb/759r2ZX
3OOA9BC+u+Eb4mKO368KmDHkLsPvhAQlhsOKJ07v1Tz3nMyKeDRmpTbBFX+O8W0OwtX7YshgsvcV
HDEPN/ibwetVSJd0CDogW3X6h5+Q4xiqLla1RUizlCtdaZ0VXBdfJQdtBX14zbJfCsAHafJJLd3h
wVytCesVuuau7bVlSlGlyUNmvM8pF3ijkLkRcoiInaDwlQWlcGATLu/eMSRD5kNP7dmgbT952G7p
fcwRuT5+ZAXZ/G7Vch8Lsa7sl0Cs2lY+YsRvxg35f0+54tJWsZTMYrSo1XjwthRvROKfxAdXvO9q
qQrYRrRsDmn1TGmn3AayxC463ji5L54ECsYX3KTo/g+dTJyZ+LXfrUfJHBUTWCZFwsORuvnbE2VL
LijTXW9DTKBBDEvQBgydrPQyWXHitNGEq/GLwJFqOU9cpaRcD+MTBe8rpsKq6PjoLuVXEdVRdqes
KU/tedXxZtAZZ0mSHPR7C6FstgExVfH1EsYCvH0EAshS8Ul/voD+8pEFs26d4ay+9HOhbzQ+wes9
x0I/BRy4O/NkAVuaDHl6+T6tMrmJ5TAVCaYWJ2FrTN3XHNJ/92ONtYO/xpBsshh1RFrybUUPDLxX
VN2bjH/yqpofdg92nN7fIBtFoVYL5NNi3ax0Hy1zu+v/UzzHpCU6xzEDhCcS+NosuyoIDfCCLmtj
oWxEm8lJr/FyLuorFJyx4VlJYmpAjwlOYKVE32ARLy9sIXWzaRAYI35OdefGTOXWP3cDdu5ae1pq
nTu0okBtYVJJDBO2lpmsbplf4XUymec+pX421j0jdYGQBxwbC4lnBpAncP3txUreD946mApYuqlC
I6+gxGR+6u5JtyUbY4jAATNXMCwmVWjSu9aC50ao1eUtw4IcyVKu53hoj5sW3WXeACdoiqMy2q3c
ciBIRtsYq8i7G2TSCOxqs/mFxBG/5YKmHpzvIYeWxz4nw0OhYTgKlZP4RSh0XwfBUZV0qVm6knC5
6jh8IAzZLQxilVz/2poOLjMUpY+7V1ZLLxErzzpXGeYyydfKQMgS6g8Qw0vUz9soF3PY04ZS4h0n
EI3vMeAtZozAcA06kdUavU1R22QsSG9ht6oXciRuTzXN2gBo9RF3lxFtbL7SAZy+AJMxWoRTO/EW
yLMeRe8Qz72ptB20Xx/yPQP0ZBHGAnkpTngsDkasq1ErRnMTtEnd9nmPTOfZUIaptR0JWSJhZvSN
jMWtKpQlrVdFHuqmLKawNotibyzZDIImvRs7KZ+Y4Jmu0l4VNyBh5Bx+l1T4Yv+3MdO6KH5sUosr
8PIkToIA+8TcXm6Soc/34SxJWd2uLmhEJbpo5oGRLcEinHkUF36YQ/CfKv7ZnEEk79/eyPEqNEcc
6BSk6hN87CvuweNZ779m0ubJ9cp/HUsW6kG5QFXWeht3M+zVlD5MPI9VPJRjawkF8Nigb6JI3e20
sTOqOG9Yu4scLKXAPV12yzDiTYvROG13pikwx/T7q+csLcUprOwRwA/tBs3lhoT66Cay9ay+9o+G
KA9l4+u6zLv4rCJXjgP8ks5ARQ46i52ajP3vxEedEIeU6r9AE5VzmjOagwi/j0Fk2E2m58ugCoW8
nQ0va16MfJjKyJEvCiEV2tOCt6/24GeGQK61tmBe15ml2CgxwXy6QEHXAP3N8CidkLbJH2+x12Uj
1Hn7H0e+WB+E6h7QtXMqT4KJkMHUHeIbNFs3BWTa0jGXN5hcux0Nntx0GM079ZXguipWBXK/A2bK
vLw9dR2KMW7No6fvXe6+i2Xo7i0Dx5xKnBnvsPbQDTKiBhsjzGMg7wdYhIZlrny7bpO6KAD03oLo
bNrWmugcNONyOaeuYnJwXnxhjuHuKKr0s5O3AxX88EZ5HNfNRsPF5pIlpgbtxLQ0UU5CQZ6YgxSY
LdbsJBkt48trOxH8eA8/0M1peNjk0iGpXmBwnLdnNWs4jcIf6q6GF2kWcH9LWv2aMwV7mL5Cj6uk
ojyo2z7DAg6IrSgngysRuLGJm9uUzNYmG+/fasD3UdR9wKO/uo8klVgTNbeRruIsVXN/yy3t4gn1
ntxNNz1fFPFpCPp4caWHlBPpzjAWS7zD5hAT2N0l+5IxhUz0A592JcA+bAMERndMUfTP1F79A4E7
GOzXp9wQ80um+ZmB7GlMjdMGVuaO8Tah7PYLPlMr2XUU96nldx4uAlxu/3nLQt06lqRoMvIXioN6
DsZlr4c0Y6WSniW3MZC4Wba7edHJuzbfEWL4WMdeRcMOW0/wuFePDW6cZBMJvgGl/Le1g35Clldb
/Fw/+kpK6XomloOAzxkXILAxzKXmq0Q1zRR107mePio94fmkKDF1x7FYaKL+vy7+6069ZpZ+U66u
zmcLzHoG+rQlHaSBpEZWhKcHLZroTP9XtMhJRsSRjrVTc3cSxY4Oy/E5Lf6gkwb0lfvoNEui8HfO
awrlvgDfocuDEOIvYQF+imvSDncNY3LzxApS2MlJ6Fb7lGyL++g+pun16Kc/paf0FfnQDOsDTtaA
DhHCV/srT58Ub9uOFMe9dgcvZQBwRJjln1t7afTQcUeRSlCFmLvJW23PiIvl6qKC/JJG8KI/PRc0
xCcqMfkTW5Mspd0Ay+RfgrcDGyCe/F/W+1H6AWUtTmuWnIcN3XvwlvxUMBg3r3saNKr9kzxF3baV
qTBMJ4Nac5bBUCxQ5PYjVri89aTOVjyggUDi93kFPnpG+/7TyeZE0UbHlKP6zPj75g/zIL5zLW1Q
/ZbECZ9eHxe4HJA0eEx3pcJX+8T51P/Y6yIY9DQ6IVNmblleoPq7rNYlU3J1ibPHUwy2m5PTdypZ
NXcIuOSCfilE/sDjVHbzk4hWls09hFlOk5LwWKjIO0/Wa05sDG7PpgncrtnTXXVO1gMrvYjPMDYm
e1khFq0LM5ReIkpn2oMVCJD9bLcVGsbUzVP6aoGFWEJk/+NKZ75Pd7aekWhmIDL4HEJ68iy9eHd3
e9r2R9i/l0++ATzyro0/52MlvLZ/W/cb8uQgWjiYuS3cbwVpbvGRLdr3Tig1X1pBAB/x/ZW8yD2A
udqJswH2xnsaaFqAtTag/BqU5VsJISnz09wwLo8foHuCAP9NJlmlVveCFAThJU43bLdCd233ofgU
SKNBYpUhur86mHE1AwjauALB9qgrSMpzuLFAy4Z2QjjqZh0GASoizFnxg/bQIEXqE+xgOmKEroUq
jk+WbAJLLqzxWe1jmfHhMyDxR/v4ie/plTee2Ff8WXu6F2V3nHn661uo33O4dZbQueecZgX6C4mg
KvzvasEi1G3CfKlfoxnkecksckVoM87K6MoupFjScSBrPjys0WXrntzsP9c7F14hhfc4XIDJqo/m
+DWxy4RKaTBaEqlQlXRfUnhI+0tSUqJuc6zFt/hiYcgYxWotEzNlaFr32HLzaUYelLIFaNvzjBZZ
uRQdZVotYN4hHaqKaQWZOP/wal9DuqYnZ7STNFxl7FtlPtO0hJu3e0lMxrJxYPPN85atK7e3SRBG
uYlZrACtZN7qtgSyWgp395reds3wfJ31iowRWyBZay28M4mFycoYKPXOTtwyIzZ1dMSu11cY9YIe
F8p/T8b2YP8e5UVEYjXRs545HSeuOwkgfIRMQI0K3gccGX5WyQMR2uEI8DeiOE3YV9dHMAWXV/58
sDp8Brn0G7k+WYliiWKRzzxYHuufvUd/wEc57djs1IsDE9/Ex7fXteywUbOlOZOl3yHer//59ASh
0BAHWSK6ar4zfZJDFdKrkf3qX5JMdV4wLh03/T+PiuTrrTW5SdQTkfnVSmN+xVsV9p37P5qpfuJ/
YgZvWqBGrkqdVMctU3AZYckcGumb3/Zaf3dkKOERymqknQputVlezb22LDkMM3hU9+TxzNmrLxhg
woapoivQQY3XKzL272787b1R9c4w6yj6ZyaKyLGWAmkhIZIM6FJRNVEitKLM8Jr6QIRnlmVfmfdc
Xf8uvTTqtz31gGp2MathDSRRnoccZA7+v/OTKXphSWm/QlH0ofF10MpWiCpIxeAdwf7yWiLgR8Tg
cV80xGmbLhFS/EObcs9XS38IzffCR9q/K4ReNnlbOjk31Xh2bPtx96YhxTh6bDt34KcoeUhyu2gC
I2qR465ifStZWyf6BCO+5oz7Cl+aMYXTW2evvOcV66Pc7/HFTqD/FoEuAT90S4+Xx3wCCwHrsErm
WV04vpxugh6Ti8o4wMn6YkWVDQ67hvFshuXpZWd5VbA/NFKHDUTgwQR6My2cXjQVNpSOjKt9e8Fg
dkr8uslO8cKKl9wu7cinDOHXBsm0kL+b4BddZfTgFkeqzYZ7pH5l5cqigRtqR5WT6Qjqko7+2Rc1
9UD/KJBbVdoXB+6bJe1+hEE8LJcXthTERkn2cQIgTtAorvdVJBBKVCyWblPK6cJjs6CJD99fapb7
aP+r7i3D4ifHfA5xgetku/Z1/nxDq/N2BHPFlKFhFzbgQImpyMJYjI17wnG4Ttrku6fKIIxEW+c3
LaGY6aNVd7of8xYQYQbjgtQJ4522ngXAyGkMLNjJSlqFyrbBBGHsnYfIWfgzTn9ww9QhpqS/8ajD
1Um7rzHPppGURlrG6Q7pct9684ebbKzBQbsWBQPh11AQQSbm5Bp7A2HHw8KB1CWLQwaZQemjRWFy
PakNJWqlHB1xKjjTEhmLFa5rffQbqSyT+gUb0tdVGrEClXLKzSTYsEq23oJQy9Cl+5KpTYj9bVNH
ucSpO/D2OmH5DTxg3uBsUoevNhmeGgpXJRt/G1TJaPlivDsGzYVy7BXhwJocBO+sTMejNEnz3A6w
fEDB0CORRx9VkF50Rd5u0UJiWuKtDL/xiQDRzYX5jN3seEevcochWF+lgxBcXreQTle/fBTSOWdN
Hh80EhalAQGl74jdhUuf0ZVo1NQ0NfHyyp+pqIbQuLVoo4Lzag6RVhdE3PZl4EOl4AXHzMvncZXL
UgCCs9X2K5zURh4yEbyZ07HTd0wYCayA1uU8Kf85+DWckA1IWNhd11nVhLYPsVtiHFcpJn9gLqJA
k2dzx1J9SxRhgpzbI223LkbF/8igIjPlvI1Drv0mqbtAZAJwB2RPN1oDbJcQ2fRU4rj3Y4Jv+IoG
au5ws/CPiCOV/S1srqKK9DvqAqg/vNWjzoiUm1nb0NwV5A1WIcMEQRdCQW81tAtl+mFSbHo5UBQ/
SQIFDGvao0WAHJy6ZAsM6b8QvJTqLwFDjDDnsqc8uQgDdpMz9nPwsGwII5i/GVLFFPXtG0utb/Ti
6SRcEMlTlby+/eSwFcNgBh43xlHslm6K6f615JbxpQHItYcneRVMhZQuW7bRWdXaFCloRlZXJOEE
NtyqzgHmtDEBjx3RPxSxhDpb0LgLGJGMaOHfpwIGIXX973nTvPKmA8HKgyBV4FaXgxJ1qEQtb9l2
UD0EcFIgSE73/RgKtCnI6JNgH/PbvdY49u2VxZOMIvvOe9W07MZlYsM6nFEtZ+/YqCsWAAlvXG+0
mt6TO7z1Ytu5Ql1VYsEvhlqb+zmbWEcK2Q1NTZRsE0xpowwZ06Kiu4RP8AEO1ipVnhEJqmRCScPh
xfN6eWkp0V/pJr5k9XMictN88e6B4EBZ/BvTxtR6oJQ60N9paYVN3ZpBFDtnytBbmOWA1xrc+giC
vVXgRu//HbJWKmZUUypsSxzLZjJXvadzH488qgrDquCo6m7Vh23JIqdktvfX5mZQTQhysndNc2go
nKTyM/pBkzZKkvsVMKtL1hE8FrjaC6uG9T6vpjhA2yjD1V3X/lvNfaGOLuhXy4q2DDTM31mccXoj
KEEbGA4ECmNxmnq/yPBXRpLfodjk8eZj6kAA76UdThLDW9i7R9IzmaTjOC/CdDn7Jco4yfhBEZwe
tAuuX0r4WpG1/kip70rYvqQNd0RusR7EsZdz9LVzzkBHE1Cww8QF0nz1ipHqG8soc53T6cUnDh1Y
0GAnT/2ywp+QGezppuqnLqZTE01UBfrBA6CuQA2N57XdOaO3O+4uKgGr8tpbHZOMN6cuQ5gDsDR4
1VYSeqrlDtWJtNDRt85/obETU08+zpss5fj7TDjeawL7NYsi+BznsWttNN38TqnJCIOFrL0ojWHC
4GfEWXGIkITHbzpLmomV1imwK7GG+IqHyikwpBfI+IC5oNMd36HlENNg1qAxQ4RP4nWEzhQ9SX4c
m8i1DMLbvfRi4neFAGIcW/KxFs0Lh+hAyl7xumsWgiZJ4nOMf8D91b6kc8fYrOYLrUerjKv71aqH
b1hnnFmimGGv+5mFf3p6vlhtp/dR6ttFyMOxXYFHyG7IlJIlyv+XezTTfL0VxVGRsIcy/jo7Lmf3
U8PMcaNiGedhiWv5Bnvx0y9UqwfoAOKRZrkaeu9czNIollgrS8MwVwPDpP7I71M23MnPau1wDZcz
hjZ+/4NJGAsE63FQZZ1SyAMeIAowCNEMDeoPqF4cMfkRsmrNz7BIPOaVzbwyqU+oXGMkIAg3cQX1
65aLmAoCNS4Rt/+er6ScmA0uMVzXlGI8tGPOpLTX6mWlFmK28VLZjL67oCN4URW+qzZmkFNATikm
EqNN6a7URE1sgDtY5Mr5BpezZUO9WZBzInRjG6zUYYbqDHindkT3JYTrV9rMIqnEtWYcj6iiVcIB
B3GhKoH2SXyZFqngf/MDMXtRU6ewq5aK2TPliMXWqL/BN706E5gkghzDxns8QgQ2GQgBTYegn/bn
O0XrPPPZEs+kVk53e6F69cveZo7DLMLj/mmsTrvM4jTg4WwPWHmBqve7KeoPO8GuDDFGiqEPSsn6
r4HxQTwrzxAY3Yp82OLSkS+4FskNDo69V6APAHrGG71rFdNkUgBWB2Wte/1YSwrbWwQozRge+eoe
7Ii3JuKpfGm0rbRrGevF8MDQc2F3IpL4jj7qGRQc0W6sNGVVfZ83DrBCODeSkn+xxpRni8j+JPzO
sl0f4BzN6HR4BLFu9oUCXfDyWsCtRTnbDLez1g+AR+EScMJzHlHEod/x5BpDSyQIA1DoPowFUnbe
xDFCW59mr6YpR/WKFcncST1/4mrBnqfMLgT4OhXM0PloCypQqd78qxJdPB2zinrVZQ09FUyMQlOp
0KLpuGl0N+oID/KWqq+GprIQVLkzTlyv2e4V/LtQJVdRhQg83JP8egu99KaZOoi1b6V5KajEdMyX
ddJTX0Ue+/NqnDw0EjAQyZu9j3UJDooK2XHLI2TIKrHuVGPV4Jf6dBq7qFVcDkN7lLoEXqHGwUSz
/c3FuzJs+eCRMfwo2ihBa4Ovtd+9D6EGLEGyIixSiQrsOlxNYWZLMfIgp/DgfjjCVgrgO2pSCt/Q
DS87brC9p2UiwYKRd3wot/N011RajrvtjzGMRG6P9ueEgrUtFsRCxNTrkw2OQc/ERMNt3Y9OPVPb
WwaiH4lwq5xGIDPm90OVTNBrROW2MMR9zDeGf/9/bS3yJogdiVSRO5r1ZmZfRtxADp1uqwV53ks+
5FWsmVkLXh7A3/lb5F7PcjOO2pqwLA3W1pb2AzFJAGEi1R9oYWjSqzQBzCW8A+QRFR93lubXOnZQ
nRnCk+JuHSb0QfxtEp8KaKH2d0uZDDu9sdZHGFYEp13XIIyagP5LT/zYz5rn9Lw5CO0wGucvQrC8
2tmITtnIdSdBtwWEU0LCURkaJzZRFVZTwHywpRRlzCYRpqAi/A8grYJ0oybWNhME+9f77oleIMGR
jTctIJfavw0Lo2oOKKHjO22OnquXUD++gr0eXKbdXINYF9jvqnoNf6EzIzgQmn+erF+GPQ+cUDNb
LXIlwrXuTv5XEiRLZy2dHiMGKn3LN5BkJhJ6eLvVcdIVTI8REZBK9aEcHpjwsdMhrWRkXTQLLQTx
1642ltDNk+3b+5CBMbommvCPD+JeR1SY3Y1HTByqessZ3ZFKdIDq25hwNAZxiHztxCqy3sm8YTsg
ulEpXuzzf6881NOxrrLW/jigKlGLt0n9CKttLRQB0iAVjfKO7OVxzbsV4INuUDs4DRSDzfrD0jcG
eDmQdZIRzXQBztOmI4vdZ0vwd9TfAYuRwwsYsyNWB/Xy0EwULxtPuXcvR7nrpil6AMv6WR6vUcB5
ZdyAqpRIIv2nGNM+id/KpyWFWk+0UWn3/TJ7EfsKxsRsu87aTB7XjdsmqLqGLBOskXxYxqVZWMKl
6rFlPmeuk39fQwPa7p/NWFP0kkLBwkht0hIQ95r/1eZMUTJEriakI/dBi3abi0l/lKDGGRxgGpB6
nmwc/tzUw+uJeAnOCxK7G6WML3fmfo+VYBLpRggQtF1CXHotCth5WmiHIy+azWpxnCofaaXBvjkH
X5E5uROhiCuclYqDfiayQ1ZBhqcmp9nxR2x3V23TSNIFBZnmyepDcnD8MTsTbGxXyPPIZa4bBSkD
02rkA6MGGF5C+pmby+UNqwoaKOXx8YAigjQpMl2tB6xSaYHDi7fWcuRoBSis+L2q+8lu6thVLlzw
tJczoYcV8LhCdskJD/N49SHYI5vonT/p0kroOU7nkoOx0H/uSPevyvauGPqDoBQHL3DC00+ryK4j
mEOzeU8kLs3xi50/ljpxKXHr4f83KRG9g2INAryztOwhPrM8g0SJxZ4nyYTRt182xnNKd6xvry5T
3ne2BjWOIHvxjqw1fldIk0kNSq9dvF6xNNN4DNRFL5UruFge3tAz0zvClqNJBbqZzG/yvNXd2clG
OW8+0lGtlV93IxqSlpdWO4tmrM9Vs+5a1SsFMTLHj+zOi697N3o8gltljQkSk502Z+YNkm9Po/4n
WKuhrjM8M3GTsr+gHHjKCo1sVY06ALzwfC3oJl168K6RFyqvzGxVI8hcK1tYqMeZzd+1rbiQaH0t
DMCORRQXDzOnsVq0WISnid4q+BWI+iq/XxVi9oMmdkMHZjbeeEVK+OsZjTpZG7skohqaiKcNdNxP
1j7hfZHeyyRWVvqGGEwzfEV9v50uoEk7Unsys/oT6m2EgiBT4sfzGAFyS7gVtG7tq361jLEYm92/
A6fZ5PuC2kIZaavwwuV/2v+AqlrF9qljBW8t5Zl7/yk0Mo7N8cQ4WBsv3OE6gXoWpLEYX/ViLn45
VgFBDTZQ9GBxyoUibg43IoVqfElSMXIBTGy5Eh4RcEA1+3rDm1iwJJA5WsR+6yLGm2m6DOGBa6l8
Lgnjy5/EXkOs6USOplogN6GCpPd6kx8Y8oTaObvrR2PL1/fNRUOkL1hlJFLrIM0K5zNgFfDpC8wM
UWJL1DMOs+aIIERt4NM5Rvqz1uLs2uv/q2sp/iNowZXEGAf9OuD2/EeOL+BICHtwQESupjPFytQS
JbvNCXD2PdQV17nW7eOyLsWygrD7kXeXQTKEcAfJP6YdSbC242HkfstRgiUmU/ZyW4ey1KAiFs+6
IhYR7zv3oc8HArTzawm7oOQSBSrw+uEE7qgqBu97Y5FCybvdwbuM002iY4Vde16ZMW7zZI7//qVb
/6N7CJOreyC2epntPNjq+ix15CVLe9kC+5ofzisvkR+3tJ6a/tHOQSjEo7b2CDBXfEKWnAvsr6fi
kYvbxAqHtrFsVBmq4R/lm3mqn8yXA5KVTryi8pKYC2Gb7PsFF9Nf1pymR8a0VQZMMNYY4cmD4cqW
qPhKV0sJ/WUst2ng6HSgwWjRn+C2Hl5vabTcQ/UVSqSDPCfVdkAiGA/8Ry5JugOyq5y7xpWnOOLb
0VWgicpl6Qj+e0zj477uLddtSgpVFdBrxXCdxOoycsJe2KmJfHw0PN+r9yOJUXZJ/ba1gRvLFXTQ
c/76JSunpRYFka6wxz78tUQJzoRpkEaauB6r2gnYzuK+qmnK9nRqj43HcyGVsdiPt+amBxiYwdeP
649anyME3Zg//aEHgsgu010hH/lZE9jedMAyZ4l7hdf4q43zz8BVVSZK6wwx6hrDzOd55EZmuFza
//i2Q4a/oAOp68vQnyYrwplVIiDxu9NSVElVBs2Evkf+NExAhmGgW5ovlbljbMZ6P3DJCyQVJfOk
Cmpp+wVHI7G/OIRMAl/zBhe87auHiVtyYTgGC0sonE4M0pfru+z6/Faycg2WmwvwcgXp3Uq/b6Jh
3qgGCzNZ+4ahIETYCLNuZYrALU31voDCcBGsNqPAKYdMVfOlLjo9KaPsGFSsREuCjhl3jUAwcHfv
Ypkatse94egTcLdWmDNiaGgd1RZDFXByibyW9tFEQvJL10jwwxi12PGbQXhLrO5xWd4zXj06BJgR
vCryk6iUo4x6X6sugK6rvvY6M3BPpPM75kE1GSb5BWyvXGgRbHJtqdQb9uWTZflVFRvyVcXX//5m
nc0KvQJdyvMUKK2zsDKVyBSJZTP8/n1wz5cKqSow6Iby7RVkYvvifbp/6RYdNTBNqbaG0FKqErvG
pndkrifCiNmC/rozILJ6un1EwbFwVJ0J/e5GWfEfqpVYjH+EsWB+X04WF26hqrFhCUXz5NsJMLVJ
/1gwSr9t5AN8KdbN0dIjUkY+aCN7H9YxR4TLvVw40EQFN8TworJ4K0uN26N5JFQeJFefMWmKgwTx
A0IaiUQAZ9o5u6p7cHmVOGjPuzRuF7YeruuytbeFolUia8iLAxhG/LEa1nPmH5X8TfTfqnBOqQuQ
XIOEsnLcIU6bT13mWUb2tXqnh1krEy6Y+CnmEiG+nO5ey8xMA1nq0PgLtkRSFys8W/vPQAB5SReb
s6ZlcLMX5c4L1OYV364ScapjN8zvflFVrqbvhoPQD9LSueMxgLd5wQunn+/58pkjSkCvXn/RP+QW
Zm/YJidAwTMoTjwQnihT4EKV7mj2T+XHEqrg9L5IxxadccDwUD0Aa8XHHnAQg2i4xWNqdFehylwp
2Ph+Xvzb3L//+BkSfc9yfIak++b6HrriTjRXIt4DRSi4IkRMAkdoBl5Zjrjjp84U5ZONRmJEAX2i
tr8nmlWxIt1HyWB6VY5XXslUq6reThmh0zCIsxUV5WVIXz3D8+0hpo1oIEx7oMgvX7cAXqjMBsT/
GHMMvEhbqr+z5WIcm8td1UbaukeWrHXDgf0abBBGBIqdCGXpFl27WyTAtDAWl42TTCb/SqwOu3Cm
H2xlRXYMSPFmLLqxWuDkjEggWfFx5esWmg0V7xMqWPuFJZGADXs8HlGpp5x80u6MUn7VTmlgEP68
mJ0um1i8s7D7s+X5HOVLHWrsVXGWelTuHdfcUKDuvvQ3GUprPyV552f1qhV2i1SNnMoGZ4kAlzVz
J30E5ehRsOK64PqgoQ1VwpOK2FE3hPQjkLmaz6aIPYpyMNvU0x4ofxDPA8pvnXsXiLHnUW3JkKPs
XgejBVWvpRRKLfDjtQfsjFuoJ2CTYux40TD21pzJLnL83c8JTbu6i1BhCvJANljSMMBvVwGJfDAe
Kvxum3c4JcaXCKDbvfITF1xJTkoxzWUhem3CiXlNWR4MorG8dHHxFWPXH3SJ6TZSmtwf6mS/pb+t
XHV5nwPv29yDm14e+aSXikXtQA/QvOMc7BBog9B/JenKJ8WqvmQLUuaQeKxyyzy2DdZmk2txhdC+
7SH8RpuqM7THTwOOtN9sE3epCvhua7OWdp/YE1n9ifbiXeIAMn04jgou4mbEMAWtcJRcCzSKkdF8
YwQxnJTEsZ1O75Yy0tCl9DUdsi8SMcuyDJbBAUMlmS4evyOz7O50qdXcoohRA+R/D3K3qBhxLKIF
Zoh8c7tDFt9UU2ujAqL1Dl98kubrJPJeijfoXPYO6o6faIWRe0mt/0SRlYw41oAALhnbtv+6sWab
gxQghcaYR/y0GaOaED1xOOzMlFE4r/axBHSBNr0hLZRCa37SHuFHzLElUX50CWbhRAVHQnYxVvlA
nB0ZR1Hy/+Fi0PkWewUgl2iPh2/XdQgKFfuIUlDHy4kKXQT0mEf/8ewI0gqy3x48c7qIbkdMe9Rg
9OL+5SDAYpd8vVVZOC34hu7tjQqldENvRFkPJwH8gH077ZyawDKw10+l+e1/Zd8dgoSNkTjTJgHQ
WZtkqfIdevDeAYGeAn6WzNbFtxzb31S3RzUw0bY/IbfQjsGj4Cz5N1J/gC1m9AM57dYhl8By/ika
DE1MaeZg+J1lrzaBTtJIewd/awyEgr0DI/5PfsrW7LkieM/WO1EkNjrY8XBMXt5pWIp/EHnetf1B
xyEdXNf6AkHmrsATE/NvCr9vzMGN7p/PGTxJ/KYrlvtGRzVy8vpI8c5XPiaBEYM0O6xE4FvOGHwo
4re5LTnAZrRPsoJdB0Yv+raRpr9tJsVMkocpKBs21NwC8aZ71PHZHoyieHMbRXtzVb+hq8A4/USX
S3w+zcttEpIzAnFzsd6lNHLq3A4Lrjl/bbaAad6qh46FaLKyODWfXz95hChjF7I82JJ2k+hFFIfs
4Zum/OG3ZRFmKxfsgPZlI1H3t4XPWYW9JwqPtVnutZGZJq3V8kvRyIylkN6boegw5XT0VXKWLaX1
U7+IOX0ctk5BC+iRSuR2MkYWfm5xV+W2/0J0H4QHrvAhlF7sygLLCd9IaQUAJG0B5GG/AdZuimOq
rvv38l0b9j8wNSCogrfAYZb5tCn5u7EDFD0OVVyPYJu1j5Hzt/JqcejAJg2TDtyxiQv6jZxy3SZ2
rV5r58d8zykOlKMzb6CcRJ+JV7MjlvQfGg7evQM+onU7oO6cdaXUJPJvhgGRTvxLNctqkVlQH51d
YlkOAdsJ7vpCoHB6cvAIGoVAK2Nz60Fit58uC3VeXzWiFPTxpc2sgX+1kPtRkG4kxPZI7jLiPwCu
CoYK/MP14G+9w98QXswS+0D7opboUFc5LkUKXZHqs3zxiwiqDjmTv+v6jD6Ob0QyK0BGFWqaC3xE
+I7m7my3+RW2S4pussoB5PWLKbe01rjnoWl9s5C0qQyPsD/Lq+jq93nSMwGdQBvrhsPx4/9VSuhh
n3La6hlb8QeJXbaL5d9abyqPjk11cNEqR3PKs7LmbuKqmcZpJVYPWIfdVc0SHfE7eorzXSHzPtRf
LXjnsGTcqAMXdYRAf4+jaTbFhnUKx/tUyv5WzLqcq2oBxnT6TAYBm5mUPhj9PbzSh7pKupP3ir2I
7D/7TWCMC6M9+g/qKqqY3mtyDBSXuZQKsgsQD3ZszSfh6oH5FUNReLPxOfLIkf68NbL4DyYMIn92
0ZfLI7ygU83bxIAbf4QXaQ/AHGPVJbJ2V29zy0nkJOMuX7z0+stlSJWD99Wi0oKhLBNaeM1ab+1Z
8g70Aymc6FOm2EU7T4EVXrVE11OMb/OzXOVmpsJy1faV9TddoJpQeFDjOb8+HC/9omEWY1zVi7eq
3dDLSQ6RivVhqOc81VJa6JEwkey/ykZlD/2JH5NgdnEyVxG7QxkSxGx1cioXuDSq8bY5BP9aK6T6
JO5L7TSm1Nxg9PpiziT5JpL6kAVqhTAqMvMNXr94laAgt4EoB0v5lDs6kPKUGA2m/0iRy4D6+ZrL
WuaKPh2m6EMGqgfPKveEA7v3CuoVseyjVOlQXADgZ1Bz4s9rwzAG19qm4StI8WRpdUT5YR5g7QyY
EACHh0YsQIu91+eAeoAJOjbxtgPYxIk2iIE8GtQRpi9iFe33tGKpvzhxzyBTkOaCxWQH7VQA+QgV
6Ap5FPbpJ0eKE2iNBLSyccBpcyIcbt9wCXGXT3zCKuRuMO6ShXsoFmqDbIbKAtfwOphV8Hc7Lljk
6stEX52n5m8bK1msC+3UeBBOisZqmatHgjvrL1Jrhf3hE1WNMs5nU7Hssmp6HcZcAVfyL1U41EFf
iLJMWguv5f8NRowvSLDlCLJ6lbrkR3VMQRFbXWXjHpIKSQQ6kfDFSZQr/749rRzg2MyxNqzylTQa
cWaGpMqHcgJlTCSEmWacheifzG3CeQDfB3Uose/UZRqCyppc2RQA7YVu+DVopS6IOQ0kJrE/t1Eb
rPRicaRLbbqChJMrqZFA2OmgUSIfbXCQaF3CqhYaz9LE07ecxXgKQPgJcTxUpdwW9XRoY0N5NIo3
arrK4lE00CLpQkR/GbBT+MJ8TIpSUKp5n+vmQfNx1+OPNzwGNiNSH8w6FVIuuMRSGTt9lrJ1gynG
7yg7fcM3Ez/8flrE3RYQ7taP+XFj12NR54Cud1MWfAuAbNThrHnRPyVk51WiR0mQaK0gvy7FJT/k
kAj5IvX2hWLIUNqBtE92LE+2OXQDgIU7dGbBCgdOLXJSxin2ga7dsh5hkYFJJsOK9PbjEN9m2Jcj
3oedY6YcHx+r8es3mXX3dZcgWg1TfnYsXXtLSR5q4Hng0SFRfWGMseIINCirKmZRlpSYZ6QLpyRd
T8GPh+hH5L0kBpQayNiI8zC7ZsBOOttP5xAr+VEl38DZSRoisM+Sr73SundX5sVVCtuSsmYn4mKu
8phanaD4BIJpq8ir3SgSy5rG60e97CiiH7xTsYzSrxtWgrX1KdspiSxqRAbFfFpPoPL1E2Wu2pcT
V4Kwirg170cwc2pCRYFvAGMvy9p4XQrud8WsXWTW0BtiSCmK5bMTnJ/7KRfsRZRmCxYTkOZIgNkc
Xw4kcXf1JFaYkTT9aCTgnkn90OytYwCqCja9Amm1b1U/fskyPUT+bLB6IhF8WuH0tXy1czk6MYC4
9JJqzyqxpcVLr+axJ5TKgcus0oiLg5evvQ6a2v+QkUpMBZU3KxYm/nBhc4ZAahg/iWDPh/sdEZGp
5Plyq7PJ3marlyXRxFFRd3bQurwf6GDNQofKRMpJ2fQ6zdm+v98Ty7T3egsFVdi6onheq8kUVYFb
cfT/J4TrcRoIjmNR4pLT7O4bCUMOnEFzHGvIEfUyLA1hCDOM3PDRf0GFLguIn9BGwrku3fOT0Lwj
Zfq9EZqTeMIeHKmTVrJFmFRPyT0iY63ShDy0G6TjxF/dEw6j5OPujWeXf+0QiOrDE01gUYDYTTTu
ZdKHCCQ0W/l4Fw55+gBg2VKTxJJxGvw2ZR+7bcwr6cnd0DrBnOmjFRj/pj9VsTFNEIEoOIsRKMFh
Mp29L/ruZiTy7CEhXYdy1JfJVBmRFjqyylE6KkD1n0dOsM4IxU0MqQ/jmkL+LsEAqJY2TErFj+ek
7R8BVshWRNFrSnvgXu7iJ861WBVfJrMhhyk7M7BeShFSu2BekKEuv0PoabBwOba5alIUCA+nQ8kT
GTWjE7XZ+ICYACWBBP5+22NPdh+B6uqamvQkhGZF8Pqfqe6misUDmzRT2Qi8JuKOXLTqvR5XY2Dj
m6PeHuesNOB8FCibiZwZq6+kmr6wtAkvFEfUunf2/AII5Im0FXKdZ+w7jGGBizmfCTmzLnnuzJtc
dttdnZJkFhi/OQ1Hc9AiAQz3Ik8Fb696vMJGqRoeLIwTPwkNk9zU2t2b9Ze9Zpy5+ZV0Acd/nGFh
o02RxsIYxpHILRlUo/E08zak1aWywU1mdQYjqs0OrILeFubVe+hP4Zistz/mgMht636j+E4BXEBS
LGmWR7sefh9eZp907bfFkereFh17z3pXnTU7SFuKapE+DxhrTREl0DlJEtCwmtT3n5tFjO0yKyaO
gWpJT660n8NKtv0n6eg0SNaRdCwiFveCx929xK3ehtuAzGGa4PWRZzniQ6i502kE3YvaeFYOLZX4
l+UdFgLxqikB/L4N8Sm0QQ6kuGxLlGJgAmoDs68af6I3HB+2uDJmCNFWkZR0nLJiMjJvevuSUf2W
fvlLubdQW8BdPsOMEAwwy13SNj3pSUFgJQRFj40eDsn6Bkvg18Vimk5iVpfekwKYLl/EQOVM4wRq
XrDLAEf7ZUbLyLeJYENl+x8fZXkI81bBj9YUuaqXHyv/tFSktv/7ipfrb6F5OIgRAWnDQKPlvTny
93nGCEW0dvnNopoWQiCPj1nErWd5wFaUL3uMeNgNhnmRH+o1a5J6qajwT44dHWmdqdwZvH1RSBT/
FZFa2dYUxJs9Pgj0NpKhePJ6EuKtEUlFVLAr7babXzVwmLu7Q8Gu8Rd+Fu6eQT8YNaXluQVc3LiQ
8g+B3z7F1ucGSzwY3Cof1VUXN6aOPzbhptEL/sW9g/525AyPygBcCykDIXq6QFHjvOg93FQ9slOf
FnHxDsDLA/IzuJ8zZFr2MHuaIQE6ExvLdOYN5pKTncAidKNGmXUoTNLWww49DJIhyoB9dDQlA0gD
1wCcORrhqr1aSmBxkriRxdyIZxOD0eVCa3kZ5ptFqdLHqq6WLL3W0ZodweBLCM7OgJjTZEEJ018D
rnLFDtLG4YHq7dXyDq7lPLAM4Z2uis4kWK5FVEyGwbWWltWxur3xHwCNZ3gGqTRPgUrex1qKBz4N
wS7r8JkXB1QWuuE0aujJ1oTqWK/gMQEFfu6BQ5o3aPVkXvq6reAM38GahpSZggF6K88JG32a5eBt
/JJTOS4J4nFtzblpyCByqzHBYnFvKGWzFH2hH8Zez0+Qz8M5wLanEdmq6oZvVEIx1ONwRQivjoa3
Lusrt34CtSVeZ6xyNVXE5IeSINauaNpLj4lp/lLkWaPhBAhHdRI9AoEcY7TV1MNzLblBL9NVbv1O
dAUq74EV9mB7see6sOYV0awCAJQTy6K7owBkZmzuys6jCY++/FguTaBJFMb6PsMCbUKT8YeUQZ1J
QCIah1cZtzu2ZBK7NoOH7k4o/cy4usobWObLjswf98eUsZK2LZ8aBW41aXs8PaftxUTFIkQKcgIf
gXJzPH0rLUuWocEacK25pEYxee8q29yj6uFrDToCdUVX5pZfFnWgMmpx9VcoONwJ9kSxgI1zFu7Z
YBFyBKFuWjxfaeeimcSRqWdQgAkoHQagwUZQpZ9Gdj0ALaaI6Ei2q5ZozXVbNUgaMlFHVybPIBEl
w7uLsiBA6NYY3JkqfAwCc3JH872g/of/ZfBffVBbKzVZP/QXeDxPEiI0hgiZRf+eX/Tt40g1JDC8
joFeHUetA4wwnzstBhM0hwx1TAFii4XWJebY3DQJXxXetaCmKMhPkbkmxia2nxYwqPZM952xNHEL
f277JkM/H0VCYiYklGjjVXwZWCEMVUV8da5EuijMYJ7W42HB8McFqNS/Vgrks1hwUgamO1HRDgo3
PfSjmdP8742y/v5coxRocCqM7yMGHbKx2xQo1c8TIpchbVN6v5PkNsBCoas+Gg2Y/pyIalc+IN6y
EuRp+9/b0cc36sQkGrPK+H8Hf1Qn2VsYJ3f6Lm7NAAmFLrh2XZR6PcyGxhDAM3oTkRqtmpCpJ4bS
ANm9UbZcjSG/gUBzdyGpWK2TcZC6gpFup+CfTo0/yn8evvM9XXgx1ZFTzUuNNVFYjXAdd8KDxAsV
k6EFIxSuwO9QSgJwb/4gdgZU3u21CuxB1d3QXuCFy5N5ehme32Derq2p6KXy7iUZNOXf6qXrpRyu
Oqh/ab8m25Xc2v89iZg44QBZIFYipD9UOf3MPMwBMRdFhP8R+yBHHixLuFeT5QMliqhF6OHn6mXB
c5ZvhbayUurkbSOOcxTQux5r/F8ttjGolfYaBXqNsxCZITtv31e3YxysgGi6zX0nLhLm/rk2lguK
6m2NRhvvmSyqcXVTKpse39YjsP61khkBBTqJmHHyiFGXxUw6h/vi03cVkpl4aEzgMGQRq1L2g9hP
P+bDB/Q+8v5ROo+geiUp2lbO2P7Zd6ip783noRwJKeCsNKABKkG4blT5u4nn/oplgFK9jBmpeq+s
0fEpM8MChRCKfdZ2kOkQ431xLVGy0pPwmmdPQG6mx4D1wlVPpqHV5wtxVC7ixQhKnxDxc6EvIJqg
fWjrp+TPbmSvWqXsyykyRAOGHPF3uzT4Yfk5uhBAfmM+Ep3AjrUsuoUEHlL0MnC9Rs3xfzy7SFzq
UqFq2xaVTiH2X0oXsjxWRRaIotRY1rxa8qXsEpMDcsFRoLZzLIOVSp66yrJpq5nPnNuU8aPBZxi9
yC/GqxeN7acflpVmwi+kA1SWcwZsUFbtJo/G8h+/1vWCRqUcuONzkqtQ6icLiU0pSWHRFTKg2vrt
7b1FO7kxIc4ZBkHCRjW6Vc9pbkZ42KNT9S7mt++a2DZCRh4hwkeCcoZRS7loMrfligUGosjBpxnT
SxXMwOD46UAfx+ZxmreckuJh9YW7dQIPQqbNq+vWOmmPEZ5m4puC8dxSLz0+C0Ybf+CHHyrAmrHw
DlaYMSy1P/B6HNj2dC8TuQi1xhLyVO109q8IssWdZtKrvaignhKjd4ooeXh9P15MTIkuKABpvfjg
9r7bwcP++06baF3VCh/Pxb47u72ceXmszmQk66XmfIgAIr/iamCatj7Q4gh7OLOFcDflSokNDOuG
bjDOYjGYiJrq+w0GNFA4yKsfif5P1E0UhBEwqG/+ljlP/yYXI6t8Uhj3YgEBKFvJ3lzidey5UqAV
816nuOdfwQ9CfvUfwHNukuWxR9Cg/F56jF+yx4Eg9RmjDElCQ32z3Gjt/Nl7raTHaufRu9Zig3eN
xEV14Jik9Xkt0YKdy/U/XQ+e0BeEIYHzOBaprSVi7i5OtgZObJcKeEeaAUc+hVObabtQKTxmCSoB
BbkTngSXpVjhV8oUEvzjHQy2a6Po742XMYITFG60Jy+H1gSYqoota/dydgLqfzgiMe9u9p3eJFUn
4/90BnVqfEkHcDBtSxpIxAmJmJcuhveOYhH6FkPexbcHQVAQigwhKRCxApL+hJXqKhVeNyIRE635
7pTAEQ92iPLoTSy2gcq377olETuNjflb/gMq/mTUsJqA9d0m5cLHE7jliOduK9SBLodaihtib84K
vVPyPoW2YEc4Dp18lWYh7NG3sPpdeyy+dDg83to+8YJcQGh8HT+A2qDTr4FKQXwNiVqVpWnqqy44
XbsJBb10iUAOnXGnRHJZMcfu9o2brps8qQJIx5nJ2vz6ixGgkLDE871Bw+Ikhbpt2hteNbRiSnZv
kE70jtqE+IxDP/5aC/63DHDpwnpNMBoCmoCS7mZZ/pDutNsHZuqhCF1du57nV7XRpyMOK0ZjBN2+
2RwjpOQdNinOf0izmuaNYeRUUogJ6/QIM10cDoBsZPrN1JcnpAQBiJcmW1JfeIKgzcJi/qf4mjhS
QKqn01b3bWU8VxL0Ga7RZejGOUR+bgqaVIKewh1CENHAMC1uagIrrxPV8z6OC1xocJNAGlmHf8Ke
4ZhKx5gu1XUDN5WwaAx9EvCqK95+oJ52KmnHONsA1HR3rqMVpV6NsN1hsVAA5k72yKKnjv1Ts2UL
a6oqY4Zo0nVn0k5J1QvRAsEXINhJhD600Ee+oLV4CmEWWtYCU9f/sy+IV7A6qOEG6yXsP0+30lX0
U23PqJomuK/iCZeIMBwtrceb/2jqo0H/HtHxVs6qv+MYYod8jwyXsRpePt3xqUfTd8Uxiw4HdVD9
8d92BqRku7zTptv2RYoYb60MArtTQLJ/1dwWIKa0x6HReiGiiXdKtgbjCJASwZJZg13qwX8pb6Tp
Lm+0atc8mUjYq96Mth0pW/8AdTM0Z6Nyd1n0pz7hc3921vHsbYC9oAGDa5mnErq20vZDhA8LbQdj
sKSwLO8gVQMD7kHHDS76eMV+dtTvqonWFySKQUCAwICB9L9IqY16j9WFepGP+BT05fixzN7y/gzD
cZE8JpDfmFGzdy3WggbMtvaefxOoec+inCYkXgGV/jI5VOEsVab1kYk7HJ56Wq86DENTMy3a6L9A
DHBeLRi1g9ZjQZItqHfPtbquVIamab2VQwLs/qYFAjmY2Wh8MfcYvHKO06j5AeD93OYCKNjCppVk
1KzVyTlGPziGS61C72i/t5I/gCLuYGljQlHJz5TuryeME3usg3hTToTW9GEfdWNvE3B1t+4309/g
TruXlXcknYse4Fxi1WIbWWsQbiTH+gCOFqFF24Np13ye7bIERqMWjWHHd5DWjswSoZ2QPfkVX0K0
onuaTeM2ypFmC+e8D5vDLjivdC33BcwcJpUwT0ZNyChjFXTtX8K/hNgz0S42Gx74ynyIqouahtSp
znWU/roE2JYydPW4OhIVxLSfgBayHTyaymR9b5E/L17IwZr4eoAQ/rWCVbKGASA1ctYLtbEbphgq
3c6WqNih2PgoyaVZOc8fDiprkCYwxE39UR8xL8z4ukMfr+navugTj6PzEr27BJGmqqpAEkEm1xwu
4iPMXJQQCZsvoTiMjXdQbb6VMInEIwRPBKkTZg6YCAI2MrHdBTE5BpDs+KT/cdHJISPZW8B5J6aK
MeQue7w/adb387fUnYcU9tX869kW2vxTbNQMtJEnwdeMJA2zqRtqw4pdg07H5PXH7jDyL2NRMzbz
vo0JvQpFAhIOAXNOrSRPVifMgsX0U0v47YwJxqu13Tw9nDlwDA+bWA1mfqhG++iV3JS4anl4X2Ar
01jWR+FT81lucTcpwag+Z3ZwJ3Ud2k94aYmIgC9utCysa5a17yD/dwcpJHIietopADcNax7Udf9x
+TUjlEkQ24VxWplSSDCI5CrzZAEEeQYBBQzfMRyRVyhg/7fJVvyTE6VdAk2l8Nt78uV8Cir1k4Xc
/uv8bGPUBrgku91pWDf97HuPfixoi7vzuIpRJchr5yCG+/3tnD2Zi89Xa+R4PXy7hrMtOnMzIfMx
QO6TzlqX2geUbykQv/sy+OP8W87qKTbnLNnQV8sQR2quFbMvuhzrpFOnWf0US7dmrCKBqgAyI+Ti
mqvmMsTQaF3pWfE4r/zRFkrAphQ22L5ZtMBhC7giz09aIV/WEQkhdKstBuUMdkWgI8VtkWOTgDrt
fMFngDlplBG91QYE0L2JSl6/XY8JdYeYElNn6FZgGe021Hxsl2cGytjua6Ov83HAvnol6m/vmH/v
QboBvZa22hvDo9QI91yvBwSPc2PWfXiq/ka0neWuqXrhH7p8Fp2PY2mHcjCYUnMf/UJRBz99ohKz
hHM0RWx2kI2JXYZURZSZPplHNO1AZYX/lHA5lX5f54YxlNl928GI6O7/pQSOBUp5e3/j0bLWxNDC
8DwLBcG1jhhRXt4WRt7oEbolVlKyBqmnBXVQyJeuYL9R9QjR1V7tEhWz4IzlayuStaI0SQAtHMDb
f3RS1B2r82je4kP4rrgeEl1fIQCRJ/mXZGC0nkWV5Vr4gSuc1/JhovuqQmmZX2k2jKCqmpHNFFVZ
MmLQ7oNzcYv4huAIBiHDKPbvPzxXaom3Kvz+SY2sIhA2x1NNf4WeNrzugGIyLklwqmdz7T6jhbsv
Bm7AZcDZKnWv0xbi12OsurysF/t/up+IAEJinpznJDuARgs9WKfAvD99hOPlkVJsyz/hFun9eqAq
s4Ix1gjbHhpuDat5WRUCnWAae8A2hL5OdYXP3LTFbBr53VMx1dGE+Kf/zCcuzUBWuMCgfcDZbDVz
Cs2Qv+yrd4Smqn/pTrrtRaAD70xPQZo25oRE+/xFeCdZnSMeLqrwbOKBsSWkKLEe9Zm/7NUW7DhB
VEOPgo5SLDWAiHsL8Wf9JaIDPRt20whlbcSZRtvM6KLguBMhxc1gKyqDABrzLsd3Szlc5tKgsYd0
ouBz0yJPUXHOKnoK6UWNnyrUg4achYfZOiQHfCGx1dBneYUjWyHTwI7TKF6RDWdO1tjCzj/iT9Q4
A7l+1kLR+J5IemEpj2deE2l+W4EeSbvSd2wrXjFhe2OkM6gTftyl8chySiRflQj/Bx+rZsRIRG9K
F5ZAZbDtfu2bmz0bxrzni6+pB4gRMytcnQAH6taXSTQzlkpl03BmRVoGffcPhiv/hyZ4B5o/aSkJ
nsGOgRSyP5vZFgnR03PyPjhH5TEzsXtCL0W12/CDnnWwlJcCHZhOx4vDGJkNL0VdBsXFdAWyRlOb
GV3h4BF7sULqR8jy9H0geHYll0Df4GWd1h9Crw4QBSDbh/OhHR5+qxVWUfWre8SDwWI83M2+bpP5
04gPW7qJvwdZhWm1M4Bt9Ryp0NP1CnU5Y+pndkwwxmdq5R/xZwr0cxQdR0HaVfKj8j2WQS5mH01w
Dk2hgyAUfRoKJQJ1NUhZoqN0wrlIXXdgawZRwHU4DlM4P2sPd0miQL0ooQ/u/mpLXEmBRDmukX7F
2wMjaezTH+8uekxQyIyXkiqYLb1V8IJokBE8gaEnbrtYYAaY49wTiLp+iKmdD8Q8kwt3mmWhmnAB
dIHz6aJTKPjoG4K4uil6fvtP834NVq+cgbcwxjHuXFZnGOMA8yixoD+dzkYaH7kHuykwXVQfhU2Y
vbISEwDCvkIHPQgIlLV5ZcWNeSCeSyThhygCKuvraJKfGCMbT3TuU373vIPHWQfMI6aV3ZFItJN+
cp5rVg66TqR9DAJ3vDH7EyRa+aHqMl+p4qsgXhQyMkXwoEA12MSCqlFiiN3nYEpnTke/E0mitVwR
wC2X8WWeDK6DCaMxt1soyFsrgJKUJZL1kRgQ3ul43heOnsVgXB3hEqiXCSj45NhbdKEtlNnMuQz6
rNr2xo/BPWFLgxqvY9+Fd2RxeW1bf36xIxB+KLN2Sw++PXWbqre3jAlae/8acGSHCGoxb+b8QiqB
ivjibsgJSqSu9VnwGNtuQANgu3LxTegwM0kFsKjffAV5wkt3p3L9Py41cPb9euvOa/NCpqoDTK6q
XP22t4bBAN8Wmbt7GPbQanvz75NZhf7TTPDNmY9WbvNk2OfuTrLm0+JbEnrXORB1a+XM2Tu66Mp8
BMgXYjL+iVVfdiY35t2oyE8C7aPwLU8YIjhy7cx5Rr6T0EIvqfl3hMdOUaCqsi0UJQktUcrL0NbU
ik/CiusNr4BkT1fzzlc1AXdadEAn/fLFxKChL6HDxqIo78UekUGDl2DPTTSnt8xiexQbBOaSj+8E
H0sTxFQ4owz9ePHDt0RA5e3/xJkwOhNRtKTgxmBf32Kl37cFl+s6bqS2VtNT4OzV/jbmZgu0bppj
SpsEJaMGQHIo90Vgna/DNasyTfFKpKBJMzhA94QIcf6yIpOax3Eov6xVNgLIT7NrDMa9VjAzKRNi
cYajuDUM0zK7Xbp6JrLg31+l5kCyr4so3x40dZS5hAXgTgv3P+8EyAU6gGXSHCHIX3QK3Gr01TZ4
6lrradlsH54MAk8IQDDOOI0jFmmS/Ju7KaY4urftcs9UvUc+xBh9cbCIDyit7S+ry5xpWXNIrVR0
Z7sb0ihkylwveu1UFlLQaTW3T8qABSuJHm2lvIqkNBmtU88FAP/KipvxmYX1Dttd87pRIZ7cYIXZ
Jwx6t7r1nBiJs097hOp9E34fvPAdwQacAV3DVsiiFoFj8xMXxz7InEeedPOw2Qkn7n01yGL+j8He
Hf12vO4pRoH/LsUoL9gYese+khWEdkINHzGGHzQDm6XrTy+RlZ8un8GWz3hwOY0W33Td2bmKeQXj
ebuGrYZio4xgu8RB2dYdkx09CHgJNCroPjFxwbUUXe3hCyTX2amixEI6mDgJHTE9Xvwt3pG04jsr
74Oq+Emd0UrQdMj3KqnNpJg1bDO1GZrOcMg+dJKrbYKQ1yuSWSpyx6tdxGPGCRt0dz/H0LowEzbL
frAa2PbAQNgMwQqOfYNLSiMI0sWCe8s1epOy8n4OCeKovA//p8b1K0stcLb9juZ6FZBdLA9hSGWV
pyhwhI55JXuM3sbLRQmNZMrveashy6BJAmQt39wa7MZJCmpI0987NtV1ISjOvL0QVexuQUVFv+nD
ivwr4Q3JHYf3+7jdMkbEqHflAxc5BIfL8Fy5g0QV8bXEEvtO2SZLPdGUf0X/+B3wgKch22yfuHSP
2UHelj+y3SWRDVqXBFLZbmZod16hxyCwcsjU4x1c2ZH6Mzu6qHv1fF7kd1BCpnbWzx7vzxRK4ZK/
lmZOrNJWE2zUXSny6q4f1JFtI/ZTI1LjUNc8C5bTDj1m+f2OJAKNdGyqaxoHYU/JYP7jVtxCp3/Q
UKaAnB+a71zp0lsOfRxttzloTKFvTZAyl9fJrGt3e1lpVNBkGB72zE/xmVjpj9WFQ8BtwH1MyfcJ
oqmshvEPDSTBXaFlDzUQGn6iClwW7Qsbcz7eFhVWKXvdlfls5cOjwFv4W/Jv67T6oXcZFhC+eqMp
TJe2HwRLOtr5dVCKu+kPYOLF+b56t/bYlHsYzmzdTKIbhyZlJIpk21UaOtfJ5Ttzf5sCcJeohP9f
biQxLxBTj4+uGcOW4B+UXZjjj1RIazEfw0FAdfgPHVY11Lp3iSsE9fM8nhGgS5QLI8e0XZ7KJi14
JGRuval5SwImZ2MF46yXw0PnLF+L8ZyBfzDOoGtUg1hQ3nYJjNntCw7HokOXghwsyGBa+dOnROL3
zgmvCQwSvwn7XcaKtC9kQnW/NrAxGjst8ZGC9+zm3OcBGeTNPITB/C6P/qukKmdeae8QCqZOPlvT
nR6LUJ5+rEs18bs7siaoTVP+hOnQj9BI/h/53s7HzNq9yBwgmjIR2KLlMBzSHP4gv37eMzg1/TcF
nRmaeg4CfvUqTjOH247VT/USGAjK+gJ78qhbqzeb2MFBw8JttrxzI7KYjBtKaT55Rn5AfZM6yxZG
zy3QktMBuBswzAFM0aqbWjqSjZN8T2Dl48H/7pMkj62ChJXsy1zReKYYRjWNhIxbSDDnzo0GEViD
L/dz1MNDgbLlc8w2JkOcmyjbiYDkuHhFUejVIL8HLgYIHPnFrwUKbl41ci2J+x1Lbn/lZoVu1Fmh
pKqrRO6W3ZhGHWTCHuji8PElx7/H+A2whGe4xAVi5pynkGLWtYfkRgbj859ZQsY5U4e3dzxhDyWK
Kf+DZTYlAqMF9BwPYyVeZnrv95+dlPniAW03+aUGHD3ODNLHkAd/uVYKDunyb1N3RnTRcU/iI2Tc
40TgRN2dcBs3z27Vh60bT40dXajr4BphPYTh7NVeC68KBUSXt18x8+eDffF85UXOKMgvegJgo5cT
e3tgsLsg+GMQBxsXmlVyUDsvb37cSv0BWRnKzFSVwXIK1CM99gc4xylv7L3xQ7FZ1sp95cYJgs4K
MnApD+BEtBHNsiyFGYgrjbgiYJtvf6tvmYSkpAoMNm/WFBZL8RGcoN+zM36rk8PNBVnJ3S+yy7kR
Uogzy0iAA2SDfmdO4jGcZ3dgx2jeMyHiU4XJuTb007gY6WJCJjykRHLv+CP5aj+m5Ba+Ut2J8tqi
1DD9vYQeQyl1RcDkT35T+l+qbxA4+BNnttnjETXkXNWiek3BW4W6/o/ouDmQWNxFpAch82odG7gb
+N6jGHBz+lmC71Yp77FXxJRECnRR36xFIh5x/LoxV9xgMziLYjSbHuAoqxwj5GusuGW4FY13ei+j
ZZRPaNke4Q+ZGkk8fP2jw2jg29AQ18xQpqf8vjdR1abSktHP3lnmr5LKfTV/u3tNZWzcHO5DgVrC
bsxLDDby4mt0w/RfLyAxSpweLrjmaLsktaTGS++Cg8MtOAnveOo074GOgH4a7otG7VUPY2Uly+5C
lOgFyea+enY79KaA5EB1OR0NcvlE1oN7g25lsAWphh8VvGLPb+z+vaO4obkz1MoQYRNJRjgo6bQD
0haoLac/znyJQSNJl0Jpa7OXlK1aMAo2wiYkrs0W0b37fMA8QpjolpbGr0CMO0tXZKvBWiaGR+Tb
OB12rwUiycl0rzNsR/awevzmKDVodgqP57Xn+J/WgRuvFKiRlyOcY42Mg/uGSwuH3zNRGm4i4DcH
TciPFzNV27/Uu6YrROWcX/hOKIwcC1i56mrWhFCKS6sz6l97iU5HxVfrqHP5alG1cUwZqD7ofkmX
x9dqG2rsUIFcFBu6knm46TsJrVdtn3G358Ri2pXuikS1rnIa+xmV4PPJ34YRoW2cIUjxFOvNgkAF
eM3G3U4GaR5f7dMRiYwdlSCSC5lsbDEkpfmdcA43svp00RBXlphV1GUHh99YsJs2bkIgRhGtJLG/
U38v6KWc+sPWRwUs7td33x1tDYbS3zYi8Hdxv+Vw6zO/F4b8ZfwYPLS+UVLCTOIFZccJuJ+aQZMy
cN5rQxdGZRs0ow52gGy2bIgB9lQD4AHArDborsUICW0ItaIBAcq1B+xSAy8CzeDEHps1fpYZV3HG
GVp8yGK03X83p9EoyuXZclnak0+biQbtpxXPSVosRd6yAuqLu6aQD4qTloT/cRte5pLReRM5h0Y/
XhmwIuUBS7/KrkMcB8pa4QIat/P5zhOPmKtQ1QgByMMbdLvck5Coz2s31xFDrlJdQYclE9IhScYi
FiXzZzElBDudAjxl5Lx0+PVzuvYor0Y1cgd2vWAH+sRhLK+OmNM3x/MHRqffxqOTbBKet3QFyVEe
MTpgRy6aztGbrD9SpFH/I72olK9jddln+FZsVTcH7RXbLrMTi4dMCS/o7mmpaC+0pdI03zye/Wug
5LKfHql1+1s/EyFTjkpx03Bn31u+RRH+NldN1JziGmQVFvwD6VYYDvEMFARCnB8HfKUiMwKEABX3
3Zv+OEY0Oyr/SFuQVq1Y1yJzuSGB34m2q9QYrsAEGeyD70GV3R6FHUPNET1nIlr6kFMGXH6G6qLn
ceEbzaaP0HmNrl/NHpkCp8LPo0DFLWHTgEOQzKl8wgOXymW8MrBt5MAB7iH1ucSUNhPChL1Hf9iF
D4k35BqF9Br213kWexC/wPahpN6eS4acRPQDRLvNeZpnbK5faXVUz9LNe6zeUDVqOd9tHfpcgfJt
YFuWUxv+5oXHBmlzIjh0BTwROhn2/O9LtSwwFQTxb/WPptNoS9V7AQI1xVe+Ri8BzaP1MprOL650
h6moI9pe6ljQfaMSJ/vjcvW3fVtuXVdQOjgujhMq7qBSstTq5oKxzAjtZBWdm3GUzhOg0UbF94qU
cZ9oql3QWICv2QJXoSL0hoA8sQ7gZPb2B2BghhUoXsraDqhZLPNAR7RMyipfkhaKPa25LoFTIdGS
DemI0xlh1ui/QYBVhuBoX2jdjKILk9yuMUzod2Ez7iy9d89Uppgj0Pe46+qXu8xbIBJbMkynVIsZ
U/Hyxy3Rll/31i9xQ081PnjDvkkfaGprUTLwvnxXlNz2A2nRRbDozEZqKVSTnLroKLRXLYiaqJy3
ORTV7Xssfmx6Htz4JIOH++oDX2ygHWDAMKXK2cFC7a+LXab0Ptuw/2I5Z8Xa5fURpiWcVSAZYawu
0J9ki0ui8dK0nTdhq5ErvKJDchHUmenNjK2FUY0kjEoDJilx5GUUnr8MiWBPGA275MLqVwXYclV2
H/c/QL0XxVf5Slu2uiIuDZrXjZEhPdOhvTJ0JFSMm7bjE8vQieXhOFJjgd5qBnJhY0YUreaCSHuI
B+lLpKMHOX4O9HRi26gSQa5j0v49APQ6dIskBOHNxUO0oLCk4/WipT9Wewjd7JPLgM7TS8iDPeVw
MGqUWX4VWZ9Pjx7vQSKmLEGxVWJhRHchcvBoiYOoELbiqKLtrEZCuepWSyuSNQmJP2AdutjWxOHc
/6kFHoYsTyWD6UkSprjpB2A7mtXd0a3yNP6RxQem7gekRgHaUfjqK3FH/y5S0hys5vDgl7bSNXo5
jmWuee+e+93CoB91ttirb8hXQc8zzwwHsSWMb+rRazTXP4u+FdnX9lBir/yES6lxMOcYEo62x8zb
WPoBHD7g6iiexy7keYO+krMmuqLOvufvjF5NJfQyrpQ06VijTnsaC3wRLwMnvGrO4Ra39/k4Czj+
nK+w1QHeutbJJ7xAS3lC/DWIQlS7OgIP90PH6UYAm2I1ZA/+kkFuhA5MKe4xeI0UEuVDUmpA8FFN
u8+4CCVREnCgum67uX+o4rOB9OzkX4EuwcpQdltfvyUNdmvgtd3Y8KTz6j8vpjt0OiPZySpbKSSC
DeI1yYDrp4FfnQwSW9PCwAqtSW/IaveqrUOWYy9UcKC4zFNCYQnHh1yeNNBWUsUno6z/3ztLWhBK
GuYm9QbvvNX+GCsDc1FmC9qrzlSDeXN+ZgMpAWAItC9atpc3bdNkWUM9axiE8WyLv6sQ97MtLC1j
FU3T3Aj7iPugLKHEYhMnxu26Kf8JgNWYIGvHBZzHpgi8PLX17r4wn23AjpRX3MLF2z6yZHcbpFGz
7JD+wxfNiGjgLMRcGfmaCkB+pnuvhjZbYcz6ZKQw8/jSkJ6wZU/vTsHMdO7o9NIknaE/SF3boYTt
TYJVS5ueqqt5TPyQLW875MbFkXvKTSUL7XaR609koW1hxSY2e42MDPowf9X3fO8cZAeBcMs/G1yy
aVnRXtkxWIRd/oRWSMNYKzVv2OT4PXFOYAn7+Q/WHMcNbG3aJnqELEpbIOsMAlo5leRlxGLxmIpz
jDmwxbgnjMXoNHDEWvHZEck/cMGNb5mE0UuuDUfPi+cYR/HPPb9V8Jr38ZFPJg9pUfhxDyeSi/ea
1CjVLRto7QwOgXRKygtK6TjHXU2FpM9bGQi3SgGNKxuOLNRxs0H+Ph/1tFEITi9fM0pwsTQdTeTI
WX1+3xHttfbBxItV2LkxMG/S5QRsfxEppgl3E3HGxUu2nIe32mvJZTZearUBBOhA+VL7i1TEomCw
PqxWP4nDkGBW9d69Y29NerVZXN5mxBLeQxkCbxb+qG6FLstnYgOX8D139KJiu2CoucoHuFfa73YK
cMH30AQkkVfJSYDVUVqJeIim2BOIx9mz89GU6QIuXfQUR1IpxXj4dRc6HdTW00Slg4tYvrvNB7ur
h+HI8wMyd5myAsdvlzfeetp498ixG+iR5exL95PqBm4jzq0IMy4x/i061VcxZD938gId8lMxdE3s
cnN0vCngLqacWrkU8iGd8YusIax4zjA/8i2JgjYePnxv9gcz4lCBXhlJx0fI27p4wuSSpWuR3Zz1
MuPdG6Qm9Riy2a1czX+NEc2D/rUbYW07iyleRNnoSk4erUTf5e+kQRcJQ0fr7iWHXy8MQcNXZrRE
gKT5gr4MhzWZRAqZTp17bNESyiCBi53sehloVFmrnmFOpJ0N4YVO4zW0eIe5WMl3ulMvC+pd2ich
zEv7tneMZe9NXX3AMZT1Wm7+U13wIIW1vvDZLumy3sjVkS8/ibX82UqaOyQY4iSUsgEeFc8Vy28a
/aRIMkEBWajWkUzxYbOu26LrSnnRAh1hJJCjW4LdZzjwC2tENbJmublSuqWrNTGuT6HcpP+wUN5H
LG8AtnGnE2v4hdsvsCEk3mPHw+fECMwBPwi/m6o79Uy30yH0IxCbARYyMCDUiipl8r4bCEEazguT
9ZI8vg1ccKjJ5aoqiDmwdt8NP0DOWLBmbel+W4BQ42mSklXtg5IwOtn0JOap3JLyjnLUzU/Vwnxz
Jsh8GLHk6YlLgJLpzVKxl51w1ZYPd69mMKhWDJQKeJbc6nehsoPZ416ieZZhgnEpxPqQfvRpQ+7L
Kxw7te+5i97iywBh+wIzC3stwGHs8nN0EJZzroV/NSbb7u6YcBjcTVjrxy0uud9N7BH4JvJJNPpg
b4n1CzVVbcktYm+e06fS9+RMbTOSymroZzACsxXWSHJdL6Bd8cEKbCdEQJnBRssov/4sls0obcDi
EhpoxROBOPqiHNla9F/n4BnjaIKnRk5hkQaa8OSE9CTE/mKGSOHcd3k31yWX7xS1ReFmhy/dfgas
owxsTFulueOjfQ/TEty/3zH2P9VaRDSpx9LEf4XwkAVdz1vD5FGx07wArvqxKE4+Upg7DUJQHCeG
WKzv/AbsENkwMSbOFpHzGuzEbfK0Ezl9Pn7oR1XkRJkI+Xdpo23BCoM1kBV+JabLzko+JHwTRHL9
bPIpXIcQMPpmukWtQq+FAVgegNl5laFAM3n1tVvHoEMybxKP7qmcT+v/7D0D75KRSREagHwuELgn
FsfdTxKcp5BAjS/GIAQ0LyIopXGovKNWBSFLqkPQDVQFIjR3yCb5fJBTZXlGkYSK76a2vLlKK2bz
Z+CMnHTrbJ00tNXvfIHdpLugPu3cSqHl4ft3O9r/s0nAGdWbPt4kbIlUhSO+cKhFXt473PjuBqK5
cKGMm+S4nOGXOIqUDrHL7VWqrSb4fFt+8Y01MSmssh57V3x+RzxUH1NlWyhOfsCZHWaSdqsvoFWz
uH3OBSQSt2fuWLUSfaPVY/3rMMS68cvC80QGHtGQIlTBFPcqRigtK8sQSltdzzL7YM6jZt96N3Qe
lrUqoAyqn+63F/tph20I/xZ7LSQXTB3AnF/bVvC3eTGbpW2tyjhATpowqd9Zl5ww2lDsQ4XZZBrG
8CAzQINylTnOlSGgb9UTmw+ujsGwdXhzOtvLOY14QrPNVPcl+brg5OOlJbZGtVG68pn3aDYN92go
ZXGJNasAYwPm0ojAS0I8suU8WQ5sdRD5dm2Es7vvowFXGupK7v0xLfEEz2dLoy+Xpz/LmtBHa7qx
KxFijv/qn/48IMqlMDJA7YWZDkX9ClcfpcMr6LPUVwRZLKeTLlMTxjV6RodCuahmo7dGivJ5j9NK
VvCYJhoKksftvvbSb9H9yFVheZp0OP7XD4Bm3T6sr6zRynbTuo5RZ3URWWiieM7ORivxLdg25CDT
S/blpcH/6naL1+ieihirvPR8JPASkgoaxtXmHRVvNgOOkdnvnYCLSzRvSrAx9bJaUyJBQsC4X0aT
EqouWh7h7KngohT5To5gGfAVnTQQ5SwfjWfSaVP4sbSxiRud061bodkZIdpv+7rPiXjZE0Y0wdJQ
AY8Xmm/nygoZdXr5lL+NrwWmiTiEVRhT3tBWWLKsGU0LUnMcClUG9NSoyCrG2o6fmPIUkf+Zbl1w
11Wtagdd+vtNF5CPWekdQil4yJlkmf93jHN7kNryYKE5tROm4GfQ6Ee9+51qt2gBX5C5Qt2P7iVC
t79rK5IqrzyiDuDo5a4v3dQ8t1vpySrngQ52mX448Cw8SSICO4N66ORYC0VqZXnn6CY5fbFXzZBk
OAHJ+pcTndaTgFA1paDJinw8mhBXK0iZAgCIjK2iZkEjGA7R+/9gh+5yj1UnqVfXka3s9IECH8xc
KrONZYxfCR9ozpnIwyjC/jACLrlB9RmlYppxjuXsHMoJeVal/qIbS/GxDnNbnnDLp9vfP7D5bT5g
014T/jleftX2JMrW4yIxi9YBBqObhsgxCiYuaQDAuXM/OGx/3ddQqgx9CL0+9/Jss4RL9MXqKUHA
lDdXt5eaDH2OtGXd8uAXWDHfPQasMqLen9zzravambDCaJySvmrWMUAAN8PE4w7ArrLOtxi9Rezu
6FU57tcND88kW2xFbGhXgHvetQyczFniCJPh8VhQiFCDWwIBL8BkdjxNbZxyyqgTicLcBCzjT/R9
z8JOygTI+hVycAbbtHYEIFQGT8atM5gfpsn1zT8iqb75EiBY8sGux9pbrv9870gG/03W1iO/h9R5
uzlP7mmNZ7xsoEFrilFepR2Xs0GtwNrSXy5lL2CYwm0CRsbOU94/rTJV498vYtG+/0rcRnCO5Rsh
57rHaaDlYZ+idXhEpsFZ9QBPvp2AA6B3Gd53BZyEMl0HRrjYW3n3JBs342wzkNl9hDOv1lydpOTN
L6UohN4WKVusZQzYVTLh3z6A+fnJXGB4WTLGgxbfEavFjHUQW6PopM5gYdSJ73AOMEOZME15aeC4
D419EOFVrZVJriFQ8zJHgtuT94cuCAxPkvTzxaNxMQhAmBFZnZdmIsPHDPQEv5I7GhT0x2i7+KBW
quJ+slFb0M+pUMxt40G8mqhK8NlwO0EBEfzGNcQiW3qBKomulKcSWEsnBdy45gh6PjWstZJI66Cs
+u91g3+CzV+7zDr1+s+5ntYCTMpBRgiP7I84w3VgJLhZZOOSkh13CiJgu92WA0yawrCd6BXSAO1d
Ett1NuaecjofDge+rHBI1xDAX7lvdl1+elEEeQrxSx7M/cbB5NdEM5av60lzfphyhv932z+WR+dp
U18485ZkIVx9+7VLBZoeTJGhw1EYqWxkqaaeqJpHiijmFUGF87wBzSkuFYfG9RzUa36eCoIXYDWd
sDMosGr+AAXCdCfD4395ndHxPYykZkUgZ5T6dG+85VPiAs2SizXmF8VdCQeMC4VrJV54h1YN2QA6
fI6GErwliophsmkmnu8GcBiuJb5Kzof2U1zpeA+DT2KIaPyzLzQIJrliSMx+Goxhh7n9s1ao/Efe
KNF7FUACLiyYza+6nO5G8qa/xXPSn//o7+4LIXwAMKakyhNEwp3vFFJ/80kLABJG7Kn7jfgPPIOE
hIj9bV8KXAkZKu7zVgDOWWEKRV/FRcwBjhIKXqF13CfYGynH/yT9pw1bpFUK7XaN83ZVUOZL2hoB
Mc0WrETA02vnLoiMKod7G2MzK/Il8tsVAs2Nb3BdGd9A2iFje0KzO+CIiSLi7oO27YNCF6lVwb1m
yxXvjDDJD/j1wsOKC6pWSKbn7PkMAyWeWCy82aS+ikwbUgKavklxZ1IdIzi+f5JgjTGmN6gQePff
1iMnJcGmvDYTgE7o08cjiTIv0o3hR7YSElpb0j9hRI0IihfQEYJ2W/MBojP69UyCaQEsCEDvRsJg
BhncxDLabXBEgKJQ0pIWPoYQSB5OabAoSjkAarRFgY6OfWMgyX+3PWWpJkkSULh5B6yJqDgW4PP4
x/g1qrB0grGOa1COO1ijqtsnVlapybsR+3A3OP5kqjqGoHp3SZUX4XfeG3dxFzhTZcQGkKj6wm71
W3hyC2o096cJ2h+tqvKigNiwsLW86tZf+YxYlbRf+9kMJhdSGFrvG6uRSxPy7jaj08Ur6vNtfN5K
PjaG8YYXnj8f5ckvTmRSqSbZ5894vY4HZ28VM8gEFoCJFRMDCfH+sgMbODfaoBlcnctrMiTCuw0u
G2Dt00KUKRxzAXrhhW99nY6TXb44xllZ3MGmrk18hIUJ08mDl3GZWUNil2WcJa2HrtX++95NdLlk
hvwFiKC+Pgd0wSrthTqbsZT2IaqoQGCTn7WpgFF3/zhOOF1OlVfQs9Pdx0TiuWUi0aVXjiyIW3Cg
YM4/jsnP5ASpwTV0YM+aGx8pA3cTXn5Rt7pVTmJLPT/XkqY0Klf4mo6oH3n6yjsxgEspK4mBXFbo
EzVYPARqHJEOpRTnufxgO60sLBqz1//WhGKy/0RGa+EepcGJsN4x0dgEs+eXa3ETEOe/JyrFFEXA
zw2Qgq5IUFyTg5WxNW8hN4MpaTDyCt+6L15rJLI9y+/qR7CeFyx0E1c0zpKArmUVe/X6/7EDh2zs
KQDhezWNe38bi0aV2QsWjW+j1UXPL+rD5cy/OTksX1y7Q0e7Zr6LQY2hUqvlYiTLvnK+1J+ZCWGh
FVn50flfVAsa2t3hYX/FMYNciIvjdolFHqoRDWcGNtBwSQSaPVhwbDwzIfQEPLzpj/N3kVaBnePR
211Xhf4JnY3mMAxqvKyj16+ULjf+tFQz19nCPD42Ld0se7Lxh+r6WrHwVvxApq9ZJV3WmgMUISgA
2zSfNLzHQAw1Q0ucA0WljffL80PZIozznUSbTNthkzd+ZVeHM2m0LY8Iuy1QJBpXCA4UIdSAteos
yOrEqCTkAXmpQUK5cic+Qq6LF5klDL3PuGi0daOqupZwKfiqe9uobRCKMTcHrTzelkPIepteDPVV
9CMWYvITIK2TYE/mzLm5U6yrN4wHLd1sThbrY2V4YkE8u/oW/VR2Xfp8kSVSkXiStd5kWp/Phe6o
pdcWAG80VzOsuGECJuImjLRGWGoiRHrkVnm/pVM2dvCun6mbeNBBgEtAFnN8f4qS3lx0XA2cyl/f
KHwysh7biP2Lb+M4rX3wZEkQk477YG1dhV1yiwL23PmOwAxxBaWanTZE7WyTvoM90jgNDgelTpJo
ercC9uQFwSH3/cLrsuwYf1N+sv3tzcURAqydoHkLOapiJ/US+/BALhjHQOm1gx1mD1ZyNIDXGQd2
qdvLhDYa46pI1C9fOV5Ed1kPN6Po5yL67zLgy6NSB1a5cWWPJ1fNjjhVyrg9nIHlRyV3I9dtfs56
L0pFA6n4FcXWACDXHPhn2gw8hAhL8lQXt6gb9LIXdbJO2eoR0dyT4/VNmJNia/33ALP90PaQCmkg
bD/jpPoRZHKZu3VjaMzSidghEiYwfeu4VowZQabSAiSY9ZrYs93qNznXRJ0/ratgMcGtEZIrCSYr
knW+mz9p8IjfMkIQl4MjEIbQqB5bMkUn15uQpqSGlYBZw9S+Ka9UT3vDv22YGbdSDqAsOlRJ8OS3
7LOwiezgE6njQeuwobPQlr1YKqdVhXGd9WIQSd3JW40JnXcORpEIcBHpQlYCzJgJgJlGrq75J6+p
8OqjypsPtZWQA3FjN/zklPLXDuXaKta/javDKQTyw50Ow9SmhrJOD0plpUKDD/LGPNEob4eXeQbM
jZN2u8zU2/ep6RsXrZf80k/fngnFQSL7DuxwenK8AzqlGQREaaqaTm8V4qSDTmcQ4e9i0YflrkLW
tsL8aIt4W4hh532peywBZ9eLuJ9dJNw63j8fbR1f54Suss1hJieDZhsPjrbZs16GHcj2reo23F56
Mb3kYYDRQJQkos3mA71kDENMmTUsJWTo0PfwFAOdCpTISZLKaYeMi06SltS6hIFR09tCAixOlKF4
ZvM11PlV+d+hU4zXih/8k+GMeAa59AsGr7fH+CgQXWiSS/F858fdWWe+TfWwYxU8lLHteZxFJIRk
Abj/MpwvP2ZXMD9SxFKqpSgPaPhONUQAe0sG9zYAxGSIwpEKRgJQQe5FsgFJvzzrdUiIc8S79uOm
bgUcSzggcohdRLs1W4OoPxNmx75NbZAnUIe8OAAgdYragbmHLsyXTl/iHftR7/X9hcgyS3nopb5/
QH72wFh3LKityNn6GC/TiJ2bkVidSuYJQCsTH4b0p0iVAAWQ72Pmdm5m/3po0+WMxjqmN0gST3El
eFcL6yNktYhetg0Y1Vomzm2dGpC2ZIZZ6vbVSGbd9N3CTF5khvX9TjVVkYQWvC3hzim1mg3OUZIR
kgCDhHbPPTl6NV1rOg2eCw1Xed7d4/ZjQ7Fc46R2oSwD62q4wtQpXzJuPFHTKZ6s47WZOj1jFhHS
8gh4PozJNLIPSXor9x0Bi1gzDWykxK4/3boSdGhgw4qj8lN6dIbuWlX0j3tBL+NAvKfqX6L8vyZO
VGmX7CV+gIJcJctl6gOOTJ4v30Ca16DENY0/EkrOv1Tp4fQDtrGNZk5/9JGf/pbVqvLFoiGGB1Gx
5b3Tx5xhPwjsjodQ8TonDk6iY5r/k1X4Kp/4pU4KmFW5tmVKRDj1tAh310u026bsEiyXZKV0jaj9
B4P/hXvFjfdndTJOXWAzAkvdSxXbTdbTDh2js5k4V31ArsFqj+K6tTgDmzevgEWeldLMTPhyuioX
UTceVjvTHJhHRaKdeNN3p6FG2Tfpndr3RmU5pQxYnQM1/fnOMW9BW1KK4fvKDukhZwX9IeuubLuZ
3MqRgC/OW4VXFqp4/LICdvoWT2XdMDtf8soYDHvPTKHjIq7bl+YBJQcGV+MbWcrWjEYSSzGJnWO/
H6Zsy7BbhQwjtWDqSIrMNAjz5N0TuOtTuBEZkoniWIPdiESjjffHlOH28gt7+evbK96GKAJ203Fx
d4GA4VE7YAKW72LXKjhzkE3awUo1WAIbfnT1VVs4Ji+ARitLZbnHsyc3xuZGL3XmPJDlw62EgaXj
thn2eEe6G9P+XhhyewBUwICXf9b669ieAFqPycKgXGRE3P1bxAnW7Imn3VRRJ0ZtTIlzbrOxETG/
zuVwUh/IGkeWdM3sTfa81PriPUcROEI1/3Hz+/vmIJsv6YqzVAM33GzUg3Fv6RXSZLU2oSF+CdQI
tq+OAJGT/6R//MHTsmZHr5yhNc4aMIuvXaZSlWJAvTyfpz5jN/2mF2bCelf973EvkQvdyJ++sd8k
blR6eBIOQHTdS+EjP1TGFrfnXZWellbdIdWA16sv+wDUDQ5qXEXvaChPuRS9xgRrLZEFoW0k4A9Q
Rt2BZQ/b4qn6OM/f3rPmmcSh4/ZXN6oxJiEecaANi1A9jwe2bKFWFTD/NIlcWx2z7ANKwLeJwz4q
4DyWoU78kQs3FYRPN2ZyvdhInbJqfkaIebaeaREpq3cfBwpVa0q0I2EQzqXBQRwO8Ezjjf7Tv+Wv
qlj4Qdfk9BQ1GYbltHkyp7+kzGr500UR5lOPNHFG5HUuz05e22K0LCtIabHkbUIkzrmDml8S6h9a
wtuwtiVXHBqC1zi8DcWsvsRVM6kR/7dPjDKc8JT04aR1bZVCmNJpSe5i70YkG6e/VuexlMw4Hk5B
NQ4/uzM6lFEWAmW0vKh2tYSgRSfTdKgymS7JJE8xjioyKD/fNvI6SyI5BDGXhgZQJhCVG/UQhQCV
rCYUj36CP88hTiB2ASCyGesOytHpG9dzcAaUynHIyW1bulxwfhhFzCJFBGns9wpa9cSsm9W1RpQg
Y4ayTtDLTP8zlW45VICBBpUt754sgm599zQqtHqbeZWGDLuP4/eTZf3zEVUEeqbWaiFMtREWsTsY
D4BLj+Kaa55ycl7vFlEYFvkuUSNtcdj/qGZrpkvRSCAlfcp9NXCp08NccFYX8nSlWc5UvqO1cldx
+Vszuk8J0krHspG+TgjnNfQIV8DrCdraAkE8xSplXaG6TOR2vfXawC40aY76KYdPXUB731vAdzmC
yhZ3EomV3R2HnprJ6amjyjV39rYxo3NREvVARKQFYkqUeNcAr5xfp4/MFZBevfQZTRYWyPFSGyDI
ds/WgB5hvQyiNeAvT4uaG6M2t5W/XeBGM3ws6S+rDntlnAvU9FPWOtNbmjvTr6omI8WSQmhfTwgW
PD9Kmaka+6jvhb/g+CbuO3PRJXzSiVlWQHyiQkaQoecf7jqyzLRJlV2ybrZAAI50DLZ5F0NaAaZG
Xqv4zRGdbnZQyBU57NYhqoeEo9r6rcQHU2uygiXFuP3ub81OG2DGPzLOrYg/0/qlk65Gyk3boM2c
X/Bo3ocmpSuhX6FoaTKqEs1t37wYSl4u0pHY9arcvXxSRL0wOtEXefEVDX/sAUcXfScn4TKK/Szi
aer6fSTTIAlyxaocSja72AzDHiiSSpBz1/TjGAQFjR/nlDvhA5ItM8C7aP7DZJdSdRmYsmO9dCtK
wo6Nj30sXJLcY8ySWiko3cAA0jQ1LJ422+JgV8io8oAjyKTZrpZiJLkM4kcM4K9wePBbL4UjuLGg
iVvVbBH1IUdDjnCDP4Rbz0AFu+eeMeXfdK/Ma49bG8VUySeL7/F/padR6Jx9bwi1ldDj4BvOFMvD
QDo8JaxcBWW2Ei/flzsNQ/ISkBZ459pGKQYS8H056JxYa0PYxRZPASckNHg8ddd5b4a7MElhc4+1
300RyFOX0fc8N1gOOosDyJSV3XMggFAhPp00ohLNCS5Ekma4w+CZMYg31pLxXTj4KK2IfYOUriFN
6VoEe5OtPIz0/5a/Txgr4ew8LimzPI+G1FEY7RMjUe2KzQzgCr1Lh2dJ19hbAXF8b9L3KgQa2LPE
FT2NAnalRKdxzEN2ohFSxYO1ewjQd3o7OFOfMU8tH1FKpnqTKrPGoKkpSAUPNXZH9cnltIg/S93d
+P3wbij6YXxWwtRjFz2LXTdkVqJrZLJBPh/K/QOBLFBzN8INNYzq77CLwF151Ns6r+vhLaAgtHBZ
SoGoZrZLi7nYDkPE3/LAk1g7kNDE62kJwKqgW/F24sxpeGt+JZ7RuDJnFqXf0Ea3QD49C5E1iSCz
BtIS++zKpF+j41PD8o9JTpMosfEqCs0hKSUoXJOyS+EF4DzpNQCB4V2QHLN/tD8zL0YlrzD+IDFn
IN6s2NzVWHd86P15+B6el6CY5O6R+WqM1yWHMYlTWiFYQWketcWyOEUpUs/CEJi32ko7KmrMyiAw
hyWgmoYs8O1cQwpjZDw6Iqy3ZmdhyA4MK5dMAgq/vm6WLCUZ7Mve7TODoGBPhikbYsYZb2NXUWa3
OAkzR4uNVG/5VgNgG7MMP3zi3jisnCc+1bEPLunUZyAP8+7kFN254pBcPkBZYIMhijsnu++CYEg5
E9YVV8sgbd8VAGzEW1P9HV4/i05OfS/yk81CRFpcqn+DcjJ+6lJ60r1ByRiYqrbyfWNZXhfKcDdk
EplzmGLCpYIRKiNuJ80rkprqwzcMBNGLQl1jN03opvqPSjhSCffuQEjIFybyiIwFqV3MlUtZ4rnr
pEdkpwTEvNrO9kHKAX393TENXipbEQZUGDdPccyJQzaLeguus1EglW6NQgAPaMmEaC2njH2uXrAa
oTbdG3CBVLlkH6ZyyDkCYqajxJhkQyxyk9WqGwd3VtaYViW4mycXzri7h5d9QWY5wW2U5ttiNK3L
OvQV6IzIuv/XNNBjNOdNpMtLUCnQt+ms2b47NT3p47aHy24OC5hcpMV8pU+wtYdj7LoFQJvJNbUB
GhCkoBpVTvGlgR9pAITbFzUcn3K5ftsw/wpmPbssEOdeIIGaWIp/SmYPd38KdqET5W/+9MNWLI7W
mPgI3CoWIg5pR59NY41uxLMN4/+bLS/Ewd/dqDmBBbEnpL6VPb8cYxn03L9QzeuzUd8QtlyAXdo9
p5uTkBcYE94G37pTCH+d1nBTKhO7PtExDhZ/XFDpby90AzrUtb2wqJy+p4+H8Ggm2xnW5mbhC6Hp
DNXWHjqc4XnPWzie0Bl9nMjgyoHIPJKJl7YtDI39vICAdcyERrCX0D8rG3RUhw60RzKYKmDKeC/D
L74gXYmMJpRbiifCsCqqbtIZgs6PdjTKyq/ozM0P6+Te/MC/P/ylQ3gKqVbZt6EpYny8JE90HkUo
9aMciGtWAhlIdKVkhjCaW5oPLT2g4lX/Afj4zG/Wn0DSlXWYQrpMqZG8eEEGWWNZtUK3SbOrH4Dg
8xcdXl6AS7euF3hZban86DpEEKQ3dGtZCmPd1+mWVwAmLOQjOSxNgRb+HhlsCf8oJ0TlkjX4iDUh
LowAss7wunSLr/Hzd/TI2cs58XiQGEoDoCn8CToV61Rrb6Hq0S+GOScGr4VlZ+/x7/fGfPTKrH1Y
NpsCctISpcIL8Uj7ZW0CSxqt+ON+OMm3t028z+CSho95rP/3oRztR2txroR0iUT4dJKEO6kaibHn
BFwT/cLYX7pFxPCPYUCiN0/YCScjSqhWwENg652L41Oz6VkMkhq5oWblPVBrwxEIWGbQXJxfiOTg
SZ5XQC9emUhbcYJJTaOQpssYRiYcbbFjc11ah9U/+Bl+wx+aihBNIJLF8Nrt+3XcMEQj5RMy7eRv
U+Te+oZvP6bossfOgmk4vTtRCqXy1XH1rvXTrGiX5hPnlOMfnSbU4FRAdpmQA1csKJ8e35gxl1Ym
rbN1Kg4TGFdkJOZbiOEke5EMhRMwenRTrAgdVtUaUzd1SZN6/E7dfulGJRbarwhY8rTar5QN0T8V
nKJn4V3ab1dihhIaPfCsUiGrmPTd83EujQH8ouckHWsjWdDNLLncXUkZ2+uHaOVyT1IJ6Ebdz5nw
30YnaYNusU94s911gbk7MPHgj/O2MczVcETd20Sm4Pj8ktZbmQnwHw7k8l9KoOvEo3Vc0wMhehLG
46p+G2ijC2HQ0PXGz3lTdLE9zkgDlZejaSLnTuu7zLiENWgIUz1CO6mExCoJ8lQsqDbuIWG9u9sq
ifjL59Bkf/JYCal5V5049P2Ov05lgQszT4Cewu0Crk/uJVCS/f5+sD8nS2h4a3Ew39m/kySIUi/i
H2rdzCcWUFYoeSPUXac2D+f2eDWV4Ze6no+IxYWfbeEQ1/VJfdNKnwa12177P0yrtg/HCXbwhHVB
lc3rLKIRkiKiBm5IvNRCFMCoW3YYVHG9/fStoOxh1SmpRVKY1b/qwFD6GtWJfiUE06E0nMd9+cfu
jdJssdEZ1S9kSri4Og/XYY6ystGRceXTBxS+Fbba9N4CEs9JWPhXui9/ss7vGAMKKaeamgObqOdP
UVHkESfcpcXY0vaxNsVeUYGbJCee1L4WsR4dxUeUaVACAD98XrvQTxorh7w0NkD6p+LuDmddNG1o
Bqp2yPNhXp2q96ZtpqauJ6gkXlboUxO/5xBe16w49l1cBgaJqfAdn5HfjwKi7b4Cn08BbtTFj0tb
tcB7mdnVBQVXpl03+BKuVQavK/ie9AXtPpLWZU/KqN/MasaKJhXki6ZdqAZKunKOzAeC4Grb3vl+
D1HTVyMrlBwuVXym+EKo9dF65HDcPt0bq0C/zMKcllkIK3cPA5KBMkqkLTPbjt2Bjd2BC75VfunG
qpDi06DjDmVjeTdxERcT6sFhyaVe5c2/f3I+ESSV+Yz1mC0kRD3qUP/1yGgoxRDv/3Hc2Ywvf+u3
FmS+K7NkwJPOSZfMX4gWiS7QJji+Hlqx+bkcU1c22EyEtI9K7NraZ/Xpq8xhjy/DluBHYEK97B8M
45yY6QnEnSdnIATkk7E8PTMODk6+SrrDRXnb0lHQEeDZ+odx8lOoe+o2/KzGXaqnT495Oj6lvJzU
txoVIgvrN1VvvMO8AuC12zQFf63eYf/bi7VBvTUlz1kkPqzwlqX4ybrk4/Rd/LAPoiKj/clPq1Ul
Baan39uSlGX4mZ4yoaWYztkdddTbw6ItSHRcEB6hIkwecBNVgoHzUe3JptsK8NN4/D99jnILA7sY
GR7rBh0xjeEzKVfol5DlhppQV3dIdmU8cMWSj+ofsoTQsdw4zy5TtSHbmVwTBs2NBoYK47YOAbRE
PD1Gg/alXIOBAzRlyLyDQgJNstNVZG+rdt6njxA8OYZlIMtfm/bTPxT5BQf69oSvHXsLyxKEKr+p
gzt/yyKBFZUXUoZDdK4BcRQZAFtK8nunUSGmyeCICxkjF18ZsmUYm0LIiXnk70N+8IbMRjU1Yh0r
1avOMLvsZWmFSnY7lFjNXYpVnbSlgqrDTSCzksqB8NBA30126bGMcaaGzdSvBcn13EVA/psZvnoe
ir5zyMK4ZlANxNak14wj9SDwme65kJEpeWiVx49FleRag+efgQ1VxGLWJGA4rzGHltzNtSeNlNAc
bRHOsJO1cWZHHEO5GLH9pTq86gOUPXsIRct50m5q1ZI/m2JRmZEKt3ZJOzG1y2JAMAVN2nO6Xvu5
ypH2ueHPL7tt6sIH2ncYIuy1NXbvRF1n0ZrHvK0uid/vwccrPLuOp1oCsayZ8tbwTpCSZIUD+ZbM
8kAg/f8g95EjE/t0yXV9JRHfHiGruf14SnDncX+RcsuzVOoEBGNd9n1nyZ+EN3lreHNQuSFa/vS/
Id7Bf7ajZRzBLgbkHpuAI1H501poimS0STbWcyDvaGBPs7ggRKRvVyT9rXFvla/EA9Xn1ZnoDxkF
oI6+eGtZoZBxeOobeMdYmBbWOkJc1wh67Yvty78UlWvqkg5rtYzNbvbKFrgz3ZRl+pGzpyX1PBcd
CB6Z3dBzODw0CAD8KljbzFl45OZJONZBTr6teiA+UQE5gCh8lOt3lsnj5unvJMaY9Qi1MpYH83Os
Q5oIUWPAG0Vkvy9EPBqMP/qeoPae4DuqOVf7K5CtbZXdLLe5B/jpmwMkdT3VgWN3wM3QjJznkeBb
t2en7YeAeveSsvjfcBgVx2GVJDDszxCDtyv6CTk3GemAk9DJc8IgJmrcWrN13zFipPuB2/Dv3PQi
p00HPti+qftm4NMng+7MgiFiBcMKJ5zeuE5LtFSXP+sjGgm+eW4qjKBG/0V/NrsEPNe0Hygb6nwZ
CHDg7y02YYhPK49h8c7rq2nAUGfNJ8EQUj6cb9OSvunWaXkgE+VaZRQ70HbmYZa9cVBOte6LlQ9J
6p8JsRAr+Y0YCmWczCikKPqm8E9MKa7xC7Pman0D4XxI+UkqWWz35jF8qwQWt0MpOQVha7u37T4h
Aa1v46a1PP9wQLnQVB3NBVgXS8SzmK76lIGYsuERKh5UZLovRJKkVPJjbtT24Sor2ceTZqEams5G
Pc6BA9xSKQzYJcXYNaX23EXFJeX8+wfRtO8sECpqZU6US/EOlAGlTkWcnw/CtmLgnFb9uZs6JEzN
PFSe9qMvkVM0vWSchrDsX2IG8fNimpJVF2Fai7eBgQ478w4mxcqMgMVADC/xdHzhKiVAiTxD8W/c
2EbmGNFSZ6PIbxQA6SjbMKBANi7oUhgNP+AScmoIPRtFScHYXwCkoUP77gazLI4TpQhOdEnX2C2T
a+k2fWO0m0SrODpyRbAzXgd3AeFsWzfsfbcj4wtM/Fgl5on4zdkeqgTsMRzafDmarrHMpMLyP1Lm
MpRmP3tM3oMz2+BtDpJMKjDuydKBZJN4VGssbxrYQh8cZYTKfhzFmjIBGKv0md7RyUBPB0igalK2
PJwWG3CNoC8azC3zyosKSEjShMNxZaV+srBdtjheB+C4AGHGKnVeeAvBqdi+w3C1F9eiU/pHhsCk
l4boU39q3QVmZMIA9RIuDp1a+gVPKU+iX8B78k9n4oW142edDp2ogxmAI+mdn/72xacTgtQPCUm9
anHgYh8OJr0XChzgR5popkLvDW99txqY09MLfEAepIr1Wn+4QLUhwUN3st77Dafpzl+Wb9A6hf4O
rbXgocoIEtQGBFCVIvMMiFBqWzGAtYALbgonqTEXqVtfj7PtyGryv5TevD9DsNwuuFhR05zsGurO
Zv5V/cRzszaY/bw6zyC44lKcy3BKnvD3GsBPXZ0LKsBEAe4Pgk2GpRwIAeOGhAyj2vXjwRgBe/TA
Cfxb9DcMvlGveW4rBlxqMXW1uFMG1E0e9bFzkrqMipLqUXqaxmI3gEfMFZU4D83T/PnmBYNoEW6U
R4HWkcoSV8MguNh9+w4LsSAQO01FwG8H+xNK5fSHe6s6BBB/hgylUIm+7pPn2Q609S7bwGZkNXQm
HR0a8POeH/8h12LUbPLdaQwOz5qMOSMxuWgy1xlM+/w9QfQdfiK4e6JDqcV2g8qp1JtPDS5+1D9H
BfY/kz9w9Vn2I1c+JsRSVNL1+bDiVl69fItHmzDmbAUdCLuSP+3f0PrLhjTpgWjSpPlsakGHmTMw
Utoa+fgwvZEVok7+LH3l9l51AMgObuUIAxNRvYrbgjpnRZni07LrLPSe3VjVzyJqgYixZqlzddwc
w3gvlRbZ3i+fC+FQtjI7RGDwlY0LkBXZxMEVER3DRYCPw78k/slFWgjt/sBTFeLbVFxj+69CTyV+
gmqayTccqINtoBgGHZ9jI+n0qRd29ao0ETvCmrxjd37+njbMiB6hnTc5ps30UUa/RkB0s5ip+4OW
yo4DT7dBnkcGK9ThxZfEN5csarAdQMfMPCFnLVxqyJclhm6s10cPi9KoOOYYqaKcoYivGdLT/D67
LQUMbiU6Brg4ggrP42//Xdc8nI2WUrUSWLRYmgJHvGIAYcZ+i/x8FE/WDATsYuDbAP4zSNbKeWm4
fPDcRMDEgm1fHSAzRgAIDe7ueN+YMRdpxoBt8c5h0D1fx7TymeXB6BDxNgNL0XCrUGIWVMAxSQHY
HCLZk2JO0i5xeA01bd4IQ4Q1nJ+RhIJFfg2384msKmRMGzzGVeSU5t0oOwrlpLfL3IwaS02+mWoK
HEwOp1yloXIT1gVRzIuwx5TrBmGUBFraMRsgAkufP8D+nOOx0qaub0JBkHZ4jfPy2Dtvnf3Ldwae
7cGkDhx1mMXoKG5AEJj2e3K4+ZzqEZ7rIjsmMAuxiDJwpn6i1q8FSnq6JA75UZHgXiMet0F/lUxY
64pSM6nA0d5AIjaPfcUWBsfjilm8jpoQyotyVCy04z5mQZj8vBL8xkAREbtn3bvaiC32pZRYyyf9
SpdlKqC8BVOJCxKFxz6qEg2CdWOaTH2cGChq+sCIyGoYScebeotU94sx0oQtLXZuf3NiPzgczAZw
UAGCis0Jd2vZwTQx3GVNdggAJ6j1b2tyY6b8GBtq+PQsef/LZ1uSFMbCuQnU0pW+LxjxD9Y/z2Tx
fhMIZmREFPJGd903Z9Edli0RrGAKsvsIZiU92vf0GKDSPrYUCm4sClc0k9wOO0ERRP7DOpeY/OqP
IzLq/GRrC/fF9+MAFNbqV1LRBg2yNHoORODX6zmD+Jgo3tkNAx2HT9b9+W9Cmrie8kAkrkgsxCab
WDKDX2Yn/wUkLXFYa1+rAOuX6o5cM2uIkbCkcOMkb3vxsh0Ii+duDNFbRF6mH7sh0vqbD20j3TjN
91McteUiVHTrOITvORYERiLXrQ8rWSqiJCgxBd6iqSDH79i0EcBv1OOY7pzwMsjeFuY+rEGSiHdH
L4l6GGD6dwCVk+xTRqaE1fwyKxrXHhOAt1OY4XE4YSRR1h0B1nyHRMYf23lkm/yjm85GrDEhBtJ6
jaLJkDXH2apPd1nF8YNdRqFYuzso8qHxz2yCuzusJA//iLC3rby+ab+MaqxrtU4l9s8/3GYcW36L
k1qt8ia5NzSUUR/RJ8VkNUTRq/PaEXmSyAQX6CsM37ujg5WXKDZeK3gCccIZ0k6ne5MVs9PbsiBo
Wr6ex8YN+bogayeCXI0sz+eJ2FYwTqtcdClbX7l+Qc0gwepRKU03okVBuI4CfJ6i9i1sYwMDb9nY
nie3H3IDxtKtw5t1Wjzztqa07Kzeeq+2qLmH3NxTliw6lcoIXCXXdRGacwCKbH2CqM1YNepPR1dr
q7atNY/DJxUElFm/sHAJ1hQnRJXMOn5V5E+aWw30mJXFyr8EaJEfIR57dgT6gzLEramOYVW6V6/M
T4F/0g2IMW1YFYbcycTFXpquDKyfNOc+Hbvr5jt4r4rbkJ0jWI84rEhcyF19h30Wnck3siR1KMk7
ZuSFeN65ggLN5R7ht39J/Bx9WkCr56w9OXYI80M3m/eDotNIo1Dt9NBpCaEpzN/b4QWTT7aynGyz
Z1t7FEtJoSeTOYDcd/lFpAlRnbgiuVcoPpMvM+l32mgp/rumlD3JqtuL57M2BZ+cUmhzGaLJyt6H
Wfs96haGLuFq3Wx46iNG6b7c+DYO1OhdU6p7oUhip7TfZRqXnj9KEeBpa2ahDHCp9dtpM66En73P
rzS1oE+wm1YgVqXNiIFF97Q2aovcWj+A0PkrGZXoXZQo2YJQtdJRgIIET5yMGMPqhh3CtocGMzjH
VXQJ77qKoDVzzTz8vHU0cRcKgDe5lAc+fMlKlaD072gE6dCKHi1kx+CucHU8UHtq5dHpy2SooJOj
ijr75gQMOiexmx5WTk9u9BFaavee+kF59vMVVUTd5hNpppIufIiYw3zHKCWjAgE5/++gZDg1LGEH
lWdWRyFmvN5V4uLrvDytrgHiL9ZJmn2WNWImONAfaXeCklM7bWSYniuSfmS1VjDNmROfz35r4RZV
CbNs+wL649Ns7pG+MufqyAzIO2E3UcBjpZLpBM1oRnX5ULsMGiZZexUQeAlm5AIxUVjKpE24Op7b
LSDiCUGhYaYENW8Cn8GgqnWOlk1e7zXgDG7gQRcHbd3g1xEqM4du+chSuS/f/HKGRtupucbshc5i
j0aecAjcV29QkfjuufcrDGThPVpPw1r2REMmiUkwXKMO4a4j4UYk5HQdV32KE/cpSmEJx7Gfo9Kc
oVAes9Jw8dKGa/Z1rhDcYoI3FONcikip128uutebYfBlwsTtP1Y3YlEbr2/7KcssrIlD7wFHvLY2
LhVQmInIaQYvsKvNFdOdl3oX+88Ks0kTJIRSc7An5WkxKEvds2l7/voQTs8pS6xH11FMqAYdr2gI
RLzLZkTy8miuPoqYbE3MwpmfPc4RItYukZh9CA2sS8COo5TtQAiVExDnYfOoNuOZ7XqyFDI7isjM
iuTCR6SVWQIkg0v4Y5O8OpiISWjHxN4kWb5ByaCxXv0AVlGMTsDcCc8oFefu3zhtnzGos7yL3R0Z
Q60Cy+NEMC7aZZ3Mcf0zrFCzzn4uS3/+6nedCOsh/q0XMuLLljC2XusM0jg8p+Kqd++y1A9GoDJG
DxupWqVZ0Qh55apQ+Wc9XBYm+H8/ZwMWkzGfYezBcnxry4I9YFslp0eKfXJ3nvJxDwAJg/+CDxsN
+5PxHKUanWS418vHaMtW2/7b2Id9tkl3WOzZk6nv1Q6iUfAsPMgawilaeCqaeUg0o41Un8CHOxhX
aIv41QOi6w4lWx80s97qAz/VGxDN0U0hr17CV6+hF9GvytmUU2hK9+xcERNzqs26VDJdWaOXNiDV
wRmipJ6DCEcBDbG6A5hHX51H/+xa921hA2ynsLEgeRCtD4xilMqFBNDos8T6vPF7XtLVlJJ26tZ4
iQgSiOg58HPaeFp9XH5tov5Mp5UfC1ZSQ5eGv0cMJht3pbdRTiRjqSUoIUI1hFxtU61Jx09mPV+v
KWK6sfmgsFEWw+GDlSw2sbtVr/ac0znpdAICUSYimn9MGFoHcmHBRgCRv3fVhTlHZJsy740jaPFO
9ZeLF3ov30hxu5lc5LXICRNM7P1v+VIEOneFFNb7M3pPAts0N3WIl2XYFel7GOKHvhiBPI8ilYzf
/1+BuBqhkKNF09UMCTox7jcOWP0am3gNZLIsWKDE9nGVnAqgvcnCQkwVkfeSyuY85Wb0s5B4ioht
rEIsVckZ16N7NlBd2zGzytMCTKtf5AzLpfkDouWvt2macPjdL1S/3TQdcjEttCaPCfi1OXHQoDvO
83mzDIS2up2jlbcupPt7HbJkUT/V4TpyKurfNvtE5UYqtQtK2vCESp3dnzz519pRaTwJ3/HeIOOY
SwHFywT1oowfX76w28cTw7Jdb2x1sTPvq/jm0dhiVQd5ioivzqz5lBMrlRuGOrjruk1fZ8bQwEmW
YODXDFE/6Jzvl/zw5IOgbEEm8tKjpBUertEuSoQVnIeTJkqaL+qnXhx3p36Q6Z0pW20fjcExgrF9
0F+r3eLjsIhenGC4Kp7Zt+zuG5adAiY/4XHfsKcJNzPPn/ZB+KfkLNVg8PcwuEOVONVzHN0ngzx8
6ZpnIcwn7P0lSBHiRO7taEn7hS3UB0l3l7n4lftjPg9pCmlmw8x9oSKSK7kOIeZ140Gjg7XjbTaD
2pyy+JRYaB7J5TN5imhNVuBOXKkTZiYSi507ejaPO3B5CiH9QZ2YJoRgdSnXEOubbBpVSEOJWf5k
h7UMA1l6wbNq4Mlk7GLc8E1lf1+m7qXuyX5v/yk8eJ3E8bKOaMcMdZ5/QgjKxkZW9KHGqYsXjyip
qU/hD3hCUDMi6pxMQS4168I+FZ2Y/LaXF6FiZJXeACm5ZjQ4pM2keqWr6Q1On4jxg+mro0LoZHWq
cVVkHdmvSUPrEIKLUejZ45wzxocFsmcVRhk+y/QM3NdGPLf5f5gJhWQO60W4iAZJxIwa/2npnVfJ
tFWAQL3JNpfNhjlHf8XwAd0Z2xxXik/DJM0P5w1qfTfSczSp1knvxCGNMZkWeUkYuT6TZY7zDGCw
6RCJ4RKTTZ4/rkOwQJkMwWvvkV1TQcUwZlx8qXxz6EFEeFPFvu1LToxEkedCiOmDw/UdpndlMQZ+
e9BIo9CFJT4s+Elb4kELUJVrPN/VfUzJOVvm2hTtngKELRSsuty6x5EhAiedWoqkXFE75qRh1hkJ
rxtsIY+k4KtqIe/QxFcHmp1QqmZyyPvhhzNt4oH1oCY5RwmHMixI6TD1KMa0Ckrie7uIndrh3Y+N
0wQkasXrrhkLNIhh6zdR0R5dJEpix9/Yg7eGtuprtNjC8Ib8rH7agT3Rdl8nyVuBz5H2cp0KVQCQ
h2tQj18dMi5/bc00pxbuGMYVZbbWk8SUJYP28BCYOFOCdnMRhhusa8DCqv2JeVTmeljnED0dOBqq
ZFquyGMjPa4Mafl+l+71D0trbS9Ujnm/ayr+4TGlV9yqAGxn0ZaclCl5KjA8OH64KPC+j6hzSUVh
t9Ys8JjozveG/ogKM69m4I2l1quTpDRqroYY6tZRoj636m5jQ3dvLBYx6Zo+hcOlnTsE1PpoYs3W
pAypPBdAuTHiHAAkC8zKNl5n61Es8Cumfd87YMDXbFgbG6qG82HsmbRb+9wc2gkas+H6HWLxs/AN
tC97F+biO2BUJswtwJZ0Qs9uZ7Sv1Qxf6/RG5tL7+s6XAF23EMxcSnQgurzRcWXCTDa0EnG4rG/v
kr49MiRhbxWReetZ/KcuQUku6uBpDDAvjW13ZefAim5JCIzaRvibuFIWiUvWwORNa1FO1j00jVdw
6gLtkptVLadere1d1imfhXJhS3jcHqUQHv2FgTDUl8Gbpn/n/6nEsG28Gknf5HrRL9TEop8Epurb
0+yjYbK4tq1H7m2zfpzR7ajS9lQldidLSfVyAu/V6krnbYrtITyhvGc42q4a7asC7/7MFew/0d4r
0fXG03HxBNET4fC+9JY7fafUYMKBnZdCFf4qST7gSIR4CR3j0hjr6Sj6u77BSebI+RFNEUGL1iav
nKzSOI6A5e/4ozaFvs5pvpjmrTUnGukW0dvHeAHjA/w5utBG+t3byweRzuO6YiJmlTKajo2bPZAr
ZXVQcEv8VhUJbGMJfrs0V5qSrnnWlOdB4meTYqhRQMdabof6swHp5YFnn9qBRHB7IzPIp/YWNz+x
QqgYbNIEb0b+qZwI2kWg3vGcckaT8soH9e4N5IcbcqDMWOPRjDAODsDNsy9+zyZwOtk4fpCYhmCP
/moUY+TWj2VqqjXo1NmWWd3nj8FZfYhLWekAS0cp9Kg+FXcJPdE36L8mV/XlWrbNTYI7eNqftfyI
gfgE+1aALlZ8DryKcBlyyd7yABNkaqbPiZ4n+mbj9zdoJukQzlPP8SLTfgzcwsjQwBgREK9sQgy3
ts2dWyRUCbeWe0Y0zHlZ/52cIGXdnLwVTnbGajZ5ijW9lCBCmq6qExrN3VDLrxC9rba87e7ZQAsf
+MRD2SBG2KLgvIawu/fGn4nVn9bxj4QCxiXweSMWrcRQGYlE8B23Tqb4VpGxkeAbqqGxdeD6kqp5
c1g/OlR0vHgLOlL9GutDD9DtzAiM2gcZg/JAXjNfuV+61KnIWHm8GYfR8mqJVyQ0IVYxuHmj4dhI
CphTvFYOopUFWJDacXfxwkEnUl+blCCXlPjBdg1Bs1VjQw2i7TDDmOo/dXR5gUYAwtv4RI6kXXl1
n14vc8kRIoFhI3qjNv+w/95T9ErbW28pZXRmd9tN4fyrEWEZ1Ctcus4XNNbYCqQ69YjY816CKDV+
LwMIDCnO4x6gv2nLihBrcjNplD1vWLGLjFjzsIJBHSujxxibhe2xoyLvayfSYreMaeUjgOG5zQFT
GMZ24WNPr7+thH1xiUWtPBgwsJSnqFTgsuI3lcwSHyymXs8moPGZxPeHxgfw9Ohr0HU020pj2tuF
0Spsvs3gqYKcdYbs3xJBuAbmyP55bcsAEnjyDYsOuM3g/j9qcBfbS5R49BcPntWRKnmdVb2KlSO7
YuEywNuRXJ4IjZN+omD6bO3RAyPRtVqUD6LJyCYP+zRIHjmxEvVPTkbU9ULexaGlIpMr5Tin3kPa
x1pKxyGoJ8djsKT6NiXa0SwfPs24J8WyT7TCxP66/lXMowWxtDCL2iw93vBc9/8wwtL+YXNvme7i
GXJbE/kqBSLOH4iVK6DjDred5//hUNiWmySYu6GzFjegxpaIP1HuXc4010eImrLtT+rJhM5D5G61
pomd0y5BdvS39rcAnG1ldlx6SMuRml+7EMxUjRwYomMR1EDfJHw/DC5mhoqMpABCKs0HvZqJmoDi
D6OUB6Sd8NiFbW0zMM+nGUp77wTCXn1Td8IYaDQ6VAbokzDdEK4hvZ3l/1RahSN8oSxUW401yT10
ZgasDEBPnfgLLKV/cpit+ULwFvVEUsYBIdWbRX6iFmv/ItkW8hh+iGpwk2SpHSkT1s3tSxDgMtZc
DvFEQbkS8mFjRBM/DIts5L00CKogEw2nVIVzhX47FMrI3j4fj4l/94HUgeNom5r1UZMlelIVfC7a
m1nUIw4HPGA32B71N+9/oaM268uuPahxtcUNe95WQ8G0lZRabTlDVZQGxtiW29ENpdEFN1TxYu50
Ya+dsnne2yNUFtV/zl1VlIbt+SeiePRGyiua7xW86ErBbba9H8WrkMU+J5d/fa1AbZQRf//8wrh/
MG8ogo9w35ii1ohm6A8HJS8pAzYgRAS943Mlg5I0tsrFidXEmeMVWux94fGZd1YgZ+gwlMsecWkO
cCboeKpi7yHJCzfjDD3diNw6P/4pGWAEV/FwP2y7TUEgRebpwvvfSTF0Ure20wXCXWdJNh4OrA3K
EK86r6qDXokKcNPFfRJk2QFdNeVD4Edbyv2QV5XyOMN0uMzeyFbSrXmjWNM7ahQT4uvnSrdNtlKn
Mofofb73TW1aDfbF1Gc6IhqzXq9SFtaGEdL0lbxvVpkGhOv4+rpEs6UMQQKQD8k+GZhkbJ3wT789
yTB2zWKrIj+xBddlvocdKL2O1ldEpSiFLu4iHPYBp77i41n2pd8nVlQVfqUHiX31kmF7KuvWtQTQ
b2IiFQlRC/LZtNiN3DSmXyw5TLP//x8FLmvHCdHLVBgxlMD4LGdq76TwtADhSMYKVpyrNTt1/erI
67TqxFnT4UHsP8kCJUVA/rPyP0FzAW2zx7S1xnYzJX5DMtjjPHfAAQQ320aQipSOB36sPxoxh6sU
TNxdeyo75n/Ienxh9xklIXxY2MRB75RIahMdX8h/XM7rdg3XRyZSGDfxyuXK87lLnMeP3AJWofLY
uH/vsvXQqW1Dp4cxYKc7YqA5u7leHgE0khihJw5txCHyKYCl3wfIq2L2wC2hjLqx9pqh4uf3sqhY
Kj1iCkESES6WatcHgNinzsLlIk+ijO6YVq+1bc8E2rbc8WjLfi1MREInkRv/WAmX2smYiV7WRY7i
8AYKrGCUTKKdp4/iOFwmi2Gh9XWKdweHhI1bQSTivTUGbupklmJJ95WOockq0XPVheb9rp7Z/YNO
swlfHsdD3b0bOX/hIZeAG16+0shBVyJy1bCOdexXjO9ufgOnQbpq5tRiilbKM7NKXIz7vvFQ40qA
9FsQtfM6dTdBjYHABrUDNZM9UyRSsuq8IBZgxd0BPG+Z14c6+yEUj7WHVoSQOBBjiEuL0HWm4KXn
N4Yuo61MmtZ5eht1LV41ZUfCdg6/I7iMA8EClKSS/XT5V+wDOrsc0aiJ6EFSAuWEc9fiJ/t15nQn
ze5rbC22hqZG2ZW7r1NJEdIE1vmzNAVfttZidLqC1V6fd95siYQlQANQZU0ekhHTPAcNFIRVS4ZW
oYoPLb3nkj2hInMuAVgIs03CPzgDAreCPnXrAIGZdpkryzw8OJzottBfGwvwMVwkc4V+pNyc4U81
icZEf3o8YgzNYVEXjHVVN5oddtVJX9EuTmT049Ug5I9G5d/psYX2SBs0DDqVIRAp1Z6WypssDpQE
lbQTisWuxRjhQXQwB+bGJtOt0bODCZOq1A2ay/NVoheRtAUXvx2cG4jHz1qwksULEF+DKTk1urKq
ON7y7BgXJJOWpVeWA1l9aS/wQE9Ef7WeyWGLf4j3bLi3SERFu5hFyZUIzOwcEh70pawCttHsYFKw
CPE5NguxqTvjU3rl+XIi2RGWLwokLY1co5FQvaI8BFB3bLmlhrzGLYSwWLuOPNhc7wg+S/zpb7NL
g9nPqFLaYksSiDAkJLuyKCvnCTVcjtONfGIbW6OeYBg7S9PGq5IUV/YL6BWKAccwlaKrAvNXoU/q
hrge376/psfWlw2y76UyqP9Sd9Ynk53JRdZL11wdKUIxfgXxzDISLQ2AOH9gOfe28wrHTocNW5lk
HcfFkqt/aRcxhBhhLHjQaGiTcpHhBMpCjeNkVoAXS0IJI+ZZt+rUPBZBcJ6rsYyD9tCrc4JO1c1w
gTlOXzlyhtDplz4JKYAXKbHY+Ta+hW+w4KUnJkRlti48D6+IlHcLav2XeMYJ9KKPerN0Siz47PC2
FDHzdrjGJAMDlSgJK5XqIaS2QwUg4uanA8SfMEHNflzO1g7vUQmJ0gDPjDCI8prYdp1RGPgA7IF+
8fIkQiJ3WTMGqG1oiuuhKHx7HY7cMoamXlvLcyq4z2Fq+O5wP4VcdVNPgd4anUcRAnpF6XrrVk9z
e96sMgtSM/XMWUO9a/sTBR0d4b71jUEZdaj8h9vU1uegHNPAd84ENypb6I2dkev++GZXixQQajdf
K+m/r7IE9Chz8NiJ1v/IlPz45+ku3nhZrQwXTR5JL/8Ka67SAvNd20VzDEIQ5Y4vl6HXguVqBg98
0OBn+aLestrpSjlx/iGUkWt7n/X1sfJsmZPXxJbBHOPadMcHF040XMUHZvFNEMO5fJdw+HaJVSpO
dDJrsHHmUDJnDuqEoy0nJJurVi9bKsTrkAdsLpXQHSeo4ghLVAzESoeWFtM0UPgnnfAp7VDw1DER
zoGwz7aLwgXSUQYO9FgDcDuUQulmQuBkc/5IigUJM9qbW5/5YfklHJgBfJBnyPa9yjW2dEvOvi5W
dIkIpJiJpwObGierHvGCVoAYGHt8wJNjV8QfY+4gr/FSu0Run5SZ093MdmMuj9vhVxxI1tO+ghOJ
XLmz2QPo9i5LhFD6guJqjaNV5g9P3Yx2EB3eCdZtr2B/2tl4AzABY2g/wL+7/G7dvizXDNF3qzuv
Y0/ZL4vS8zJIc7ExUz9vT8nVEvPg4MIDKQyR0UvTWXzzO4yIiFof8WYFkGQhJdBKsI5XUoZjD398
fVWbZpO5cfOPp01WqUzsihv6nNRIGSSFgPsTkBDsyRcQCHx9P8OYN2r4hsiJxurF5BP+6GwKZKHF
m4MsQv0US+6T3WT3EakHYpsx67ZcKujbju2X6zHg30i72ytFxtVliWixyXYcVg3cp67Zwyf7FqiM
SCL5UWkX+JwoOjVDKx4FbJfYnC1myR+L3oFPY+xn/TdLj8WJr6CF9w6q2FErKJ6/iOIBBdc/QqSh
4EiNxFUPZo9WBahHSh3Bppvodo3rcmhrFji18h6S/T7xzmi9E6OX+ryLsMYNXIy9LD6wPmgJRTlf
nzhoXPj8eIQq2hi/qD3mz09N9pNq28rjf0SEuTjim1ldAauoT6c/p4k6XyYNLx/lQA/95+stqZr3
XG0TLmBwZjvpu7wjCfkzeRrONgz5yJwe4h+BlUmGlaPfdDwt5unve289h5bSa53osUuh2uU/+WIq
Tpmx9m48SVGpy5iS8FnPmQAzM2X5SonmRT69GHyymONPcG+EoUetOc+B2W+//Y3+ttriYtVdEhVr
cQHMKXzqnu2vVymurSpohrtPBDw8P0R7yoCM7Npuv5Xo/fAkIgXBS48mfNg4CshA4upe5lExKcW5
LD3+d6xyFQXEX+gZobH/Ee+UPIE6sT8d/ggbL3wGBDWistZO/1lMyoX239q12sLLd9oxZb9Im/4g
vxj/TgfOjFxAlpJe7WkbNfT1nFFmy8C5SzIiFshRvmMijwRAxr5VO7sweM7dqinvGGicNFUoIAWx
pZ3kWxHOheNMuwfFOLvG4jNuzl/UKD6ClG3jYw8c51RRaeb2NbF8aDmec8zRwadFeCN/+o2PnfHo
UGs6VbdSwOz0lsu+ar38Mf5GyvvjJ3Ti7EgDCDpJ6To/NxOojlBXCD9v4JBTn2mwTckfSgOEX6RB
7rzJ14IlVMUe4X35eb3eXp527uksPahWUJ25JRtsHm+O4rklg6FHcbfNlD4dgFa70ukYUr7EtoGr
Y4pGDWr+ktA/CtQpbcRsCdFi/bgaqiN7ZK7rXDIS8Y8HEPa0YmybpCjk4eLd3VkjYW0MkJPxpTW6
hdClxrifkb0yOuCEz3i39TTbXowftkY9GifJl9CTUz7bpkn9/S5Z4UhYbLxARfaKFHsyQmbeeNcg
d3PLNwXGXFzg+Cw7dmecHb8O2pWOSYp1X3ckftazHASIR2lNbV0EMcPfwOldgrD8NUL+Jhwu8JKx
/67Xdyg9Vy2Jz45CFAo7rtKA0LHt/RQjxrxuSKUc/Cus7iDhTq+q9iDMhGDuhMuCrIshQ5oD904G
1h4WZbhqpitCiqkjlxFXrzUDxkX3Qu/PxOkzJ+ONkkIApCMItldFtX0ZyqpKcLzkJWMx5S7szQm2
csrolebL1Z3wGVDQUHlhFzaF77TZPGgwo2451SRnuwswb7ASKCNwwz9XCwJcW6HaLQb7mJHlNBod
5M2cvc2CnsNqvYOptnmyTzxt+47H+vy+oshwUnz7K3apv7X2BdhRXHY95dx4ruNHoi8TlFyXQMkR
l6IWFFcebBt0iKiF+ZGD1bnvBMSBwpCkDigZRXaUkDYfPKAZe6N0G/MoBZQlj9YXcZumUesC8Tm8
7zDed5kek6GDwMiHOUaUFYH/GESgc1TPTKpkhqOhHPD7pScIKZUX3ajCIstXBBs4zIYaBuNGGP1O
5r0n44oXIItv7QAkagmFEU20BKfCv+7QFViWGWhnOhl/vXDl3s/076wER2RHjqMkdqie7ELVc9ta
Jrg3DSwTTJ5E01kINon44peS9EEwG2G9cAEirfRrKJ5m6ZzB8neZEH5mT5kJ22/7QAEzPNtK1v5E
JA5ShNCxj5VBcR4eJWDCtpvFiJYvYdAxN3cfn1QQM2qvfpl9khP2TxRGl/Tt+UxCxCx1h3rp3Tpg
lhyqSfl2q5KbDchzyaWTn/qpRpJsaRs1Hp5PnN3SxSve5/th6a4dWjWE2NiPfl4OkE6eZIlfgs+v
DmZGKpLE+sLb8iwUS9N+6AdDg+ye7towVZXIDEI5YjF1fO8qZMBEUOj6CSZBo/IMexok8dKfDikw
O/uQLsBXhgJzTz84I4+xpIn6SPjO0uDxeOaRAVyarw3oYFOIFAc8VNm7WC3IKIIdATON1MGqShbw
fEnqTaYIYi1wnVjBrN7VJbm6SgNGPt6+AdnjCsn362pfLgZeLs/q07MfYk2/eSf3MW8alvBjc6kI
PAHzhOuVat0rad/WAO3ZNcMuRtUlQ0NjzM4pZBB140ejJUvZdjmSafxwLwuhYsd0rz/CnWNWskbB
61sIwrcdFmiYHI/OGOkpvWB4OZ+jYm9SGwIrtv+pEMssv2OnDZDx20kaq/Q9fgYapj4d6CeQ27x2
S3tgFMAJPyqm8HPtQqaNh3lPHK1MRunTUer/Uv1lr4VtbLF1KxNhcPZ3U8pZ0dd1gP9KCW4sK3CR
ZOKSd5gt3w68jlo2QYw5l2eljDLGMayfRN3OAAVntV9MVEDYhobdFQcKLkR1LDKPjVzAqVNT+L/R
q5Ru+jKSZ3JxGu23a1qmOiI14aiNNRRw11Py0o4RYmiTWuar8nsOhWzyCerO2HvlblTjjsTefJ4g
l5tQeleFHSmw5s+FRVMvlIsodqYRZf0ibCGOXN9YxHimuJbQy7DvldlmOR64yUZzu+LL0wJIGvqR
O/JlCwNC5ygnTjlowk5RPCjteRSd4ro3Aoi6EnKvST2m/1kXSs1OXHYd80dOG2pDrlN5eDxmn12s
Qg1dPsraZ8vYGxIEov54jVmyXFk58cSOhhf891c9vKm45kjCgWyWlOvqUikV9d9stoLn5tM8k6ht
tgFRE9lawofp51aNwCe8DuNFAq35rSuhdfHSDsV8W1PyZqywkrGD/q4CZXfcmLv/GXTYolkUiVZx
nEO8Nu/yMwtPDPddYhXL8A0T2oRoGwOwiiChZECajc7pzEDa3IpJK9MPd0s/RhBkrPak0urmvNuJ
N5klV3nS5hbGYsGt5VsHvDdaYdk2fEflHx6O7lqsIGr7fTh9RYvYj7kLvtpYHCNVcmj9bQf/s19k
ayRVYvEla3q/AjRfEV6eyKZzMoV3W7LRvWVwh412/FefSu51RNqZuyBVGH3uE8tU3KM905b79DTI
MVy7YCMP1bqarL4bMQPorn4u0vLRE/ougR2gb8dM1+XajIZAbwumFwQZkwd39FdkQFAYwtaH1oDK
26noIeF/1GRDQK/cQdGGKHeOL+VaTbgMC0kc6L7RytSWiUy3DZu2yCn3JrY9i2rqgGWpLRliVGgq
YqJX6xVneK8rGJDCkBgcw1BVAWqkJC49pf6d3WpkRkLvuhYnMaCci9BPfRGam4zCSTZzfNc0XsnX
Rlc2rOIUuXEmn9Viy/kTDOuChaicyu5WM5BDsNgBnum+/K/lx2/57OJ8Vm7UAZLRZHUHtlnLFfI3
7LPS4+wkq6mFcIUi34E6VZoCE6Wz+wFGG1FOJqv3/qB5jE8YXbCHDwvsLDe/kG2fPHwUHmrHhuce
bbE1N3ptFelYTZSblMC+VTXEAPY1K8IEm9J22j2air2pb/iE/PZe3qZuFMgop43EbHEztCL8i2Qc
Pm8TqovCHmPbYrVpfE3j6vVQ/kv0RRXXrdc9Ls3k0IZvQB3oCOmVyFccnirTqmBMtR3LuRwaQF3t
iMS52+LNoM/hcu3+0Z8oH1tUaJvQNCvqSjF6uvsrOphCWSXu2Z51F9P5smemGhvhl5re3LpEuSfn
VWHU1iipVmdinZV/+UrPRrc5rMhN4LFZdRdo43ZxVE3dzYt5kJybxexcR9GjkkCf9CRjqwb4eUhz
dWCYS1AVRhs1tZ4yciQjiA//M5wQcwDLQUyjw9qFX9Kwmkme2Xd9ewrOuF38myMy9bOtDYfzMBSk
P4jMJFwxeVsr+D/I2PFqffcnq4DMiDg4R+p7hMvEYNi2DHpFKF7U2ivglO5OWEzRPUYKcGIyxw66
voEVW7IJ19JVJR62LSRA5Eto5wHXMAp9F52nNgwj3xt5zxJorCWWApyyi8nftNxI6GNlOp/tY6sl
cOcZ8BWLnY9os3wLFGxsgw0A4bCOGXJvDvluOpRo6YccHvZVRGkFT/dCKEUNNGCvlzFIeoxt8j40
xpACHgtkkqwX/cC5BeLoh3HOg0n/WNHiH6m5thS4VCzSWrNCq5K+hL2/2wivLWl5r6zeYqTXIM67
RtcTbuwRNfpk4oRgRrhnozVcpmZWlQyWsNi/02ZvdDjiz0PQRtaicaxIKVktx9fg2+pN8eS3xRf+
yaOk1lJOQhklTBRakQL31zxqIC6pP0YMKSFLXkN+/f6na9ibLMhVRehFGEeVA040pay0tpwTkAya
mdff3EtkWzHX3araNH7h/d+9JLxvVljSUIqmKXI5MrhutNTqxVCJQJGdHBffRtHuANlgV0QkLEqd
wjWlggEN+nRQSO+1v8W4HHV+OMMAtK3TqzhNuRdemmJcal8HsO42PWPZ8bcu9XKsdtogvSBaqAvV
USZWb5kq1TCtmDi6kVfgQ+895vKI3V3poplCcB10VzbD5fgmAVBNyCtPplA60Q0jF93V9PdU7R84
ED7mnXhvSvBRWPibty8OegnEAvO8r/iaZODnyFMN5L0ngatlsNb5yARrDgaA2SV5ufg03OfifEWE
GQSq6VsnCeJKiXtBBw+gk2ZuFzPCanLvcUTJP+nYszSDr4PNSLSnTdVBsn0C8hdigsNH1EIKhC3O
ZniG5pI6NhgpvPjxW/0uNsdP+fsYbb8hElhQKlvAxgqMIvkINPHJ/tJisLjKmMnUcS/RLsDadjAf
/Pg/hsbPti/n+OvP/ft/puKcAI8tQF1M9R9vukZB2WBOLl15mOupUvYNANuPtFQ4NpIvu2mi4q8f
yJA452c4LzcjlsGHlK5EMUaZWXGiwI4CL9szsMF9+Gi2FNx1Ls1/NXwxS5gT8aszcIs4Vboa8zAQ
PaZct9fKVSeeoqCr3AUphNhIvLQHelNnarYP8+f6pUg51sz5mMbxCo2VqzVwmzPxhngfJNTQsE1H
IfBU0cYV4qDtpP9DI3JN13EKZlU8OBMkdm1d/mx8Gm1EnWhNPpKyXJ2uwjesEFQrP/XruiQfilkI
wcJDLeJZfT+cRh4Q6pyqLBLqYO4PVeitQv3mFsC696dy7SfFqNkvjxoH+iyTBAAeIXZ61n5DDD0B
AAlRuJTkKb/Of9b2+WevWoS3IvxbNtvsV7MIsynThWsI+LMqdvejC1TJyJGk86YOBNS7jWrFgfdJ
sEJXyG9o9JZL4fcu35lwLO7kqaeMZJgclgM2J0fW4pSed3jQCEctYGqUgkMpNrhnGnKda+sRUhIP
RUJ84fMK1igdMNNSvdjHE9yguX792+GPsfzw8pJGR5HFD3wt2Jr8vo9ak9fIqovtzIZwWf/x896k
CfssdHl08Fk6VptG+gntTEGx3NkSp0fQvYNM0+Y3OnhgvZLl/pm42FL1VtWWI1a6nNzXhs4lR68o
hduAq6ZY0RW5sxZJ606fOuImNdxelRV1QauRJ/Wq6f12FxtwQk97HgKRTTXM0ZpMlQGjZtPMy+tD
PAc6mExcCGezZmGvAYvK20sBJ9wSCm1Gk9inH3RsU6hiEgpsD0sNGAL/G9iOmyl9kglW6FIOatia
LhfRNsyjyZG8HzVAHowcmbX1ZbySVKmoEvpD9DIsqVyHbr+J3qY3oDAlt50f9yR4sDOlZb84ALM7
krFPQKeBpuw/Li8wu1uV6qyLRKiz4X9fB/wNZNTzIEYjrTyrGRDYNZHvFbZm9PAcW6PbdTJAugZK
PYH3RX5hO9YYrQ8aYzgq9ZyIAb8cGdvJBqt3WOasNiQdJZc1dQ2uRiNnNfui7X+KDTJgsPmr1wl3
Z9TtE8N7SEiGFO2muzXCvM3NgfRW6ExlJFyrk7iZj1CtzqphqvM/A8Sy6mH43g06mXzr47GWQUqg
ZvlcDdIcYdL3Y5bZOQixfJEUu+4Mbb4C3nseSYIwRPXRqduOf5CN8/1rfCUeIHpx+EakTJTZfvWr
mzirfLwu+VUVPygN1xrcCw2QnsN0viyqUG0qgLvJ3oSy02T0cnCnweNBv0hp2Vzc5qCkpruuCYZi
pfiQXQhSC/yN6a0V2pqG1PEUWfgTJ4QXGwNY+RhlssR/pegpEOml9VOcJ0i/yeAbBtNK0SNakPE5
wHkINpNYmaEUJHN4izvMTstlQNLWTZ6Zvm4qWcwrN6ZZlzUwfcnRDxMbLzCkHMOOEatb0OicJNi8
IuegsxyWryR361AhOv0mVlurcoIKg2j6KLalQmKA+xDr/NqMoiNETA3XmnLqLax5dbOjr5j/fBsK
ZinvqQ6W2656fnjXPD8uuWq2OEcF3WfQBUTfNkwwXEi6g4rJ8vsKvyPYNv42TSja2n6siWN65GIb
ie8dpbzsXRt4bOrPxDXbi/R5w4A2nCbI32YFFFcAXZ2R4vODp304GwrwEWRrMHT/kS2COKKSDv9R
lVG0ATPzs/bjAqAqvooClHrsSeRzxjeGHl2/f/hLFvN+zrlq0QxXS2v+5Twgsrg408LHVWgpXmR4
l3TNqTnKUaxbXBRPcazumITqMoCRHuoGCyUOsfp5A+QvyzJpacYmCd2Zlk82VBdbDHbEcY8Dxo3E
fSAqiwise6Eh3MskvuSNU98XaTncRGU2mZuMi6GZtqw7GkgI5rLiCqeYUUxnjOAHcXEkbv5qXcFt
GHaw8wPpYFLchiCvjyw/U0cHlwwvL47Z3HseY26Wyxcb72KT5MZ4FxPyxNMTsJrGO+gaGpW/UXqo
0nKnXH3X0hD2YTQRgxGLWcSPDf4mrUi+MugeoSx48jrYXt7cgyx0LfgIiPG5n8StSJl/Me+9TpYt
ySQEdzbanZSnTuaa92l/RWScaKyeTx64x9QGs9l7b9x+ARHdvF5x1eWdqG13j6Eisr9uHJupdLoJ
D7AaOuwV41BDI09Q3qm9+Vx0VkygLLnw2U23VEFVYijtTi4gs9E99J/ZsFzEShSJHXxrcCLekCtJ
OTabMINHOP0uGcCUsvHbCaMBIyxuGRFnMkAOq9e8dC+Lr+yX4ye8J/z0ai4rZnt1fiklH01Xp7vi
ncrruz3n/Rnh3h9Tz/mK/r0kcdBp2kENaHlJjvmIPfMdDOVhxKsgXch1tk8c4DFuJ2dkQLhUbgWg
2RyYmvUFueSHaB9HEBViQB0SEhz6qjjUBWOfWaZudoYMcqvSuIrGClExl8s1T0Pe2sQ3T0cJtYkp
nfhcZe4n6KeZQSRTiyU+eccWm/z7MWcGGt2oJVvhq/29MzkxNW/yQlDbwv/kC3kw7X1zQnI0zgza
nStTd5QTgw4C5iFnmsek7idFyOOTIgfGAtLG8U8do5P9zCmF3DED+80fZhRyxlGEmvboxSSTUAS4
oDfBC5kSxQO8yiOdcLtDcdADoLX3m2a3WoZT7oLDAJQy1nDtkeGvzS9ef8V76pSGIrhMayjskOZJ
o6Vzuu6681U/nYejZk4yKJf6+KxPAEl/YLCZpbxEaK6uL34XZkyGyn2BIQI48oEqXAUzzttw5h2Y
McbO3iCFfBzz8G3iR1TK28w0EPj1ZBtU6Ow92bRy3maEAQPOKWecCE3xj42XrZ7HYylWXQ8wXJjq
+a+jCrzBJdDE70vSN3NrGxy2mMK/urLnQC8SSmzckApxdRhL2D7qghGSwDNMFoFZC6SUKD6lGshX
4jvCqpHxCcDT57U6zcouaGeze3d0ix+QqekBmMKGSTG/FZrrL5/Nu/+z72r+NcvcM8hFoM4QNLty
AbTuaV0YJPcGMXRDeZHr7Uvnfc+xRdaly4vZqicZfSrBFikeeh+H8m0Tp788gcW83u4iCFATXooX
LcknMya3yZFyhOIZI0286m50HvfLRrBcwmlOjfVCxVYL3U0E5AIGmMAT/jONRln9uW9AbgVod0aL
dDmpNwxYVDGMR9I4/iHlxpxpdkk5hQ9TRXdO5m+n4y7bwpLgHbWxs5kpkvFOcmjv9ndFonrcVw8i
nZJ2mFR4OmmmqYEjqbYpLbtA6u+tAQcDSb0lurOISx0gSf3NZgEcXApJ4117pOeqypy34zp5yrVB
dAHfQNAkU1fDuTeLn98lg040F5S4mmCEsOmvHrdW1Pwc1UVfbkhF9cMBr1SOAnl7Li7z2EBde7Ip
FZ2un5+7xOkJsbLQ0+B4Hfto3f/hb0jV+v3/ahGUVNmYITVlsZcTGChF2Xm4LGECI5xINDK0dwhK
MYPkC17h1XkDpTuAjDenRDaBffKOeuiRClOihQocKpQzOrK11rCzqpW5rE7jkTUnhOMfZtv3Cwvg
2Qdgf2iFxC26g9bd4iqfHC1ficJclrx+FxxP3fXLzRTt3d1Wyg94GH3G7g0d3v+fNbWJ8F35dz+b
l1TWK8NkSqAGMewwi6oY8buwMHdEcB+PTiL2t/aIb7TOe3xw/mRuCgdGe8Y7j+uqwWU6nQCmF1RZ
JKMDPHz3EdVpDo02EvpPZu2SdLTqU/bbb9P/cPkAF+bvRL+4DiLYpET8+MS7Fi6+6Nk/jfSUzEVx
Og2sKBSAxrC+wzBOzGniUGz4BXOhY31+MJ/KXba+8C28wGGFYX0ZYh99a5AmgLBl5USO7aM9h0zQ
yAq2ohQUEh//MMK1nsYfHx5j2vS206Uw/LjyZAeQUS0hwXIJt/HuQDTPNTYiZ2Ip2d483drjyYL3
nO47WPmbaFYA1o8fZxIKXMiLSRCj/4ER/lNiHc1MNGkfF4ofnUDxkKR3O1Zz/QVSpJyXorQY+Lch
ZGjvT8ycCgPHJvk6+Kkpfe8dxvIATr1Al8EDKbM/7TwVO6f7fUoVUio19uiiY+B5aasVL8R6+/C2
2BLf+AgRZ+rpRTOVFcNjTnSc2pTdh/Ozq3gwS6Zgg/dhx0F6S7Arsf3DiXeo3NjfnwN9XXi0/QbJ
//A2JiQ5K6R44HNxuEYeF22YRIBOmoUAG0WkRZsIUh2w1OINzlwKF+oZ5+B16s0oYLD/1fu0Uxxd
DzWd/W8Ra74sqPFWEtaD49M5yWn762LLIj8LgWI9IGiDWQW6OVWqmoTCx1oMCJdVgKpcA3DP5apS
zOjnuEIu9dIleDN0qy6VqZ7H2YgVjNH2KQlLKzHCPo/oFlotvuIUX8XkD/Izgp5M09SDMJ/F8v4J
zNLfFHfKBPAlnloB2cKxmzn9byIzNGXi5ZdmRAl/oBo/6Yh5vUc631crDC3VQk3GpUbQmpHN6hL3
3Ijc9t3Fy26ur5aNEvlBft68BakmAMDytdXuNzD/UN8xbQRo3hzoT8zUjxafJ/bRlc2VFZbFndGX
HQLU/meewIAgc3tkFBPDpoQmfrCht/dv0cK2KsbzgjV88ogpmEGR13bRi3yh1A9LmGaUAz2zYJwg
tXI9WRg0FosCgy7zYydRuxm4ncYx3uz/MlYJ+4pCVadl6XoO9W7Huv2L2F9mzMlEbN/WhzfK42gi
2eyUVRdv1ph5u4BuN7em3JWQPzToSExAdGBAELgCDOfHSxU0jueC3mvrQnOe+4JbhI3T2E5yYC4R
2djnNNA+wbmDtemb1aG2RrFs+JSiF+pUEhE2h/YkUrCBL1pkLF24Q5X/XLVn28NPtWvav7kR1j5s
H/6GjvsBsvWLAg+RBeeFRm4YFdHC9GRx+ZuMP5VtdnzNIx7GKvGkr3yeAu27JPaxk1heN8XGImls
8LtLnQ5a4izmGSJ7eUcn1spOpZq4LfzRazhlg77IGojuAmiQtA1X6B3Dde4TwdZdEINxjuCqO1Ju
xelv87Sc96srBB/cpEkDViH6PAE0rHpMPvXSIkZmrnFb4qRmdgx6KSDYcxglQ0Gpqx8nNikvts+x
YKAF4tOXEEyuwP7lVeTL6YBciPtVqnAhz8JOiL/acBdHhUgwlVbe9BssXtl+4zXm+qic5EC8cq1N
U3IxS3SfWQ7Z/gj9HFHl3a/e71Y63TopZpsc/DT7fY59SkXAhiBfaUKbr+m6Y+F85nHU9f5cw/Tn
QnwFtochrVSwAF9S6EsaZGEdA1aO5/YUCrzGlYvAhZek/OGGKhsBKpNnBOe7PtqXXa5ExUV/hCqi
HeVxVwhGB/P7Q0N+CZuTERtD8MDbSPUXyaAbNBijTLoh1n67t09q4hW/IG4+js4n83tsFuJyVOXO
jeM/oQban8kbSDx77BMJ8g0hnifxQ6QCcrMIQk4pFJNBG5OLYyHcyWlA2Zd2nCwNRWTpkR9gIHIh
fp+SYCeJqlPGNsKDVN6iezaenYo/sC9ATMlW4oEv70dTHgGbFDn7/jptw/+hC+DaQVfL5GIEsPHy
fT+gD0hqDpD+88WFsDOCPBSo6RZjCSLh4EAXZUQEYwhF7ArrGQKat4qALGSzy5B8JK1WRXX887db
+V2cddbdIAMmMH6Lun3NB8w0moPl4bpIx3FTHHANF/Iscj76tNNrGnAfeSLekI5KRV8lQumaiBBW
6E4mhBBtDaFmDUhARQ+7+iROfDj8wc1mSNB/jpMEAZDxDsmqkFx2YK2pASHt0iC6agkGmA7y5kcR
VmFJVMiWFOU9el+RZjSYGhaQ54bnYN3mVeWaF8ZCaO4Pr/uEuo/+0xl7UEE/QWr969FXLP+0WTD0
Wp29Fo70ZX9lgf1R0qfBxK4dpN28vmEEcddc0Le5J7R5+HzTlmf5GMmEu/S4J8YekoszFJrqAamf
QnE3zGPhn1FTy0mlenaRia3akta+d+n1Hq3fwB0k93rzYrcGi0pHYCDCZ5YOulD70k7I3e7fr0wp
VNO5LGh0rugc1hBynHqK0yvwKcprP8sIgyOMAV+A8xjx6t8JNdCBZc6FylIrAmoM8kxNW38cdxTN
pkM/KY6R4D5jhStv6EY63LctUc8FGEGNB0+8fPcdOHXUTVj51Le1Fnf2JfYgPcKmVs5pdVPxudhV
NpDQUnidQamXL/YRE0feW91/IPdRzWwLxpnG9xdVyRvuH0jlxDdLo/7gzxjK5UTrLPoTHApao1dy
4Xif17YKfTPnhP7OeFfB0We/h7LMdbfE69UcngI+5nj4rmgikzzbC/gl/7xGRkQwZvK/OEZfIuaY
6HP79iuK+45xhl/YxLv6q4sL7O1o4ejwpjUbQNepPaJr7PjK9DPuOq6eeRHa9XwOBs3fmYIHcUiN
1B/Dp8AmthFs5L2zZ6qLME+xNxGaKIGb4eQIb/b81q5YsO3V3miEFdsFSWiATsxwb0jrvxK2oGNv
dfiepwRLrLylSighpHCJ4qQEDEkP8l+F6rM5dgeCcysh4EAabaKXT+x/UT3d1D+h5TpVMRZt+YwU
yzRXHOFjPF+7M20mOVUELKU9Uc7IE7UVqwrSHAX4I22kq6c5HzxpRwEeDB2g/kzK9P+c4ntdnxz6
naOeizGUMZ8wf9JQpAy5v2yahfgBqTX2GBYRLyFAIQA6OA7RFnFz1JrDOX56lAawBwBd5su5SbAL
fofBa2PyJKw4/d5V39+zVQRaSUoKDt6uHPFUOvl6gJ63hhTIP1w61ZPWYcsPkg4eRJUuuE1gSgkF
vP8H8a3BzSAlMsY+sovpgx1uWXEcsO3lu5Z4CxeMKKpeaKQcleGYsH3HNUS7YJDMZ+CtkR1KeUKx
aS945k/oxAy/Ce1QXAmnovW0WoOiv/d8tNxdUeTIk+FCh4F+s2JHQNrMyfp8C6B9xGLkoSnEAde7
7wXlKJtjSYgtCwMADMvrC/FqdlSwxl1hltzu4fgVb83I+I01rwblPZrjrZk4rRQpiaCr2Ejk4kLH
bYhboN4FB8UnU7EdMgBXfV4V0ctbjVCFT52VeDM1AUpl+1SHhZXzRsXFEoVb4uv2HEa5C25lt80b
YELiRleF/csgruBDoJrHm1FkiPQakFuZu5MWmF8mCYyGQ2hNLoONg6Nq6eaiXZ2D8GcjbDcuVJc8
0i2k5L4tngB8dGDnbg8b6tk81tsLl8gO1OF2j3Kn9NTlWJnXPrS3RFS8nQwxEN7IaoBednid5e5e
YOaGXvUWxrqZxkZJWnDVOrW1sQGZqXc70DZK8AMakqL4aOHZ2VMQv6VlgLzXlXb7PtDKItobsxXt
+R9p+LbFl9CEUdMaZfBsz1G+3jw18Wi7Aiu2J/j1EZitHKW0dErDuG22jM81sezSdEqfm9Fb28B6
BPLpKElv+26+YGK4tBFTOovCjMdZWYLvD389gAvf4OQSpeVn8lc+NZDabaSdtcrg9GN2iT99fHUs
jrc+UhFOgwNqs2YpJvwSyBnREnPVOsNw65yiSszFbjzwF2zQEBgpJHb3RuTT+gXKwYZl5yj7KPQ2
oYxgowWT9d+Us5J2/ilVvJeYwUn4yCPty1Xa9OM43xZLHz4IOnvVJtPTl9dMspXEaQymG6E18DXS
SP38UytAvD8mYRJhuoCC3obgrUMPAHcqCEJXhkll38PySusvH6ifVJc6rmd2ep6KFOOVDuPzyN7D
9TBQaN/U1ZJ4nOziCo8US5vsdBfVc66qFSORgeu8k4Y6BUJrLF+UwTPh/3Tp8ahu2UGYFsEezqbS
nKxIJJlZP3p0vSQgFlMRvvNS/rFOIWPIJdNUtXpKBccjPWNJJUouWwR7O/kBc5Tfufolf1jNwPuJ
9RuEzNjdFykGqBVFKPriiFkiTkkQWAleOgZ8d/NgCazUU2r6hMcspOnANWAkn5bNsdDiuLTog+Gy
F6bywTXbDSsFZwQuHsd/UXGC16b0vq1TW/KAG4iBqGokcyew7dPyGFYGYKO74dR4wYkVxVIZ5kF+
dNZFVWX6btsu842ZTh5CbZ4/0hqp4NmORETwrF/Cz08b07vILWECJ4Xm8D6wFr21zIZHzLLiEdhi
/3wO95rLXsfu+RlqmsfBMR3sOdN9IBYD/Ai0GgOBxAICMG63+LZoHkHZprsNghMVnZFCFb0kbrW+
PjIAEdQ/aRKkrYXMObdfQ+91S7z9+nIdSxVHxG+hLyAy87I3zHX9vNjKtah5dN/yZEvZpJR2KbA9
wNlKFXTZljpIa3PB6qlKKS7LH7XF/d+baVNXw38v9ZX5MgPgD4+ArMS2TrTE6xvhPwzq64rAm6FL
mDm3ApGRN6Q4cIkrAdTcR/j8hMzmGkdgobiv9ROEf+CMaanhw02p7HCHRJAcHEcqNAIhnmM5yc0W
Y5mgTIts79JZttZNQyRExgOVUw+37+o3Dhnfn/2ZgZHQoyNoek7gEj08sV5DktFQCP+Fzt5eKtZR
NbOVuMH7vd7Z4o6nMcyYCN7UXw2oPbCLUYUV4HyMJk1Q28sB0r/Y38y/PH+58DXkmjW4G/yG/DIr
eI/9THJBksMRfrgTcU523vfHGElgnNbq82sdM4dKWiNwQT6Mdr1BKv+qyyU2sKIKvV9h9vbURon4
ig2gfZh4r8kYBgxroo+ywpDS1Kcrwbykj/d55wOawvc788iGb9ddUwj7WPIYwKm2bywsFmbirmZC
mxHWkWsXRQoxqDNFKWt6YrkS8jDqaNZZtV905gSm+RopPfpP3aRwUulcYmtQ6ajgeANSG/ItIoC9
5DCnOcelani8rCYfSVsE7Nt3+foitz5vqFEgP3/xlhCbYqgcGTxgnfSHs8N/T/sdj2Da3z1aLoa6
OBuu1hX34JUfjKCqJw82WFkzYNyONZXLXLwDPX4tpNY845qIHqb84totucn+8dFHBIWesFujLeQT
UYPMMk/IQtknx/S2HuJAII+skVt1L/EHKxfQXWyoUKlT/PrK5hzGc3cF0i3p89lDu48pD3gs8Iit
sodlraKSDIotS00JIvwxkkVXmC5zwcbr4psOANz9O0vJEymnanVLr6KuO/2Hp2mqwi/o3CpoXvYI
txPyKETBgSVrARMV/K1gWAylGN/MgnueC8cN1Tq43oo7PCIf2nGiNRqrIYqKeg94VjzfWKA9saqS
bxLR5RvIp886nM3O0Iw0W+f9B0fIFpeUao1TsWe7EBK4BIp3hD0/pYOn3cdquQFU2k0DnpJuPxNX
KXDksS8fmg3nX0AktZ28cjm4+13jw/7f9Ov69u6YyuAzobtEK2dgEQZrFQjK0/nYMApGvKWsRSd1
iKiOxh2BXXCHtjegdbXqMbreFV0PEH2bmBZ6iYiYG+FDqyz3cPYUl8OsGJ/NtqA0e7iOZgXWsU4b
cLUcR/W9qYMpI3SeU1buDjEv/1NPlp58GeUYFG1nibHlQ0ANvdKHxIhp6uDU4F+nvT7llAmNYVMb
QxFbjo9J+UlZeNQ0ApskkFdSbN/wFBGoxYFTHsiAMiN+qfi1A0+2OtvLroAJ1AWpGOAA3O3BsHli
8iQGUegF+pe7kDihtRu0gXTvdoNHvmk9oqFl8Qeu/K6YAZsiUrxVeRRptxYpQICy+eAjpACXz0lT
Dx2csIF4bzA3sLB/+JaRJFGhDKxyRjL2XuW8Loy39HAGxbNxppRAncy6T70FsAyPJTBzzhOQKCkX
6V5Zq8aNCR5zvwodyCUBWgZ7oBiLOyyNygEbqtWwyrraAW41s8//u2LiWR9R1rOd1s0Xb0XxOfE3
UxTyx8WidYpnMn1aMysluIsBKNoUxGRolJ3jphWDUAYlOtew0MNa2Z88+7xMz7mQwPP48PRmbA4M
MGxyW9gWHbJa179bakOkT1eAiBPzLvFqv/p8p0lKpDzbaE3itidtBAASsc1rEB8TfwOjtpqZJkQQ
b6NyzILhwYIZu9QI0cZqP4xIkelwNmf+PkVGzrhkJZeSi9TGwAapY1KdW6y3EGM5to8cGksrrhFp
HS0VAsbPFitoHw+q7+/6CnFREy4jSw2xzv8GEOBcK/3ZvLehWxSz5NUhaf3SC/XPtjRxbGvtX7c7
KgdlZPYx2Vs37ZjH4FW4MdRuz1JYU2JKfROFdQ7P2lApqvkOA5qQ+AhnK5OG/UOayBX2nnJn+cDI
tUDATzt3h+woyOtcd0L1N8MGgo4gopOmSrwO5IxxrdhyPgIWTU++r2NvTsPCEKlZDemCpVIRgw+a
ZjTfbM0jnJnB6vYaiRQgO+LpF9Hp/UYPI8z4LWk4A2PIxLb0pNg6WpVGMnnGRgt30kbGhebUCk5T
NyCIHyHNvVCbQM7/PLPU2AkXF3YeZfmGrMRtvyGsuGtRyo3qK330Gm0+zmEXmV46p28tSJiE7whm
flPANueqC7vZdBj1/TB/Ty4KklCtXVvwJXAUk/6BeLMRjFljNytbuWIQeNqsrnmdQvvbdPMhpopB
ReHxtZSknYV92sZUJ6WbQ+QpWat9TSwr+LkzCOK9+l+EuwHtJFCvAFfYuIOyqm3gINfmReY/hJEF
L9+VsX+LdgCqiSG1PYPHVne9pCe4vIK32CRM/VX7NtSr2l2S93Vurd4BXQKcB5hyjjoTsa2IlDIn
eBgQUYDZfwYFAKPuM9Lic3sreADJjwczyFIXizJfvjeoFTk4fB+S1d3fgKmX98Cu/lNLtHSVSPXr
TtKUzhMEUkKBFMmDIUwHY5pIg0uwgBa3rd1635h6dZJ3zywINkgcZ/+2N/BIqyRM6W8Yt9kNZ5oe
2TLs8EaP/5I1kFZ+kl6mUn83uOEWUKSSK8QzlT4DA7mMgI5yfpCqrs4Nm4BvrFXiV3mHuttI42Ij
z/ObKoi5TJBo4zshaIfZPRV+nO2i2Zm77jbrFG0w/e3q4SffveeFeJe+KbdniJeFK/zgBH8L8SzN
NJ01FmTvbZmKlDuiFG0Wvl7CUyfOJJfzq4CFRCgp+vObgG8HBPNC8hrgx32K1se6qB5GsFEahQPz
ssqHayYnMUgEtcYxQ3L88wb8IcK+YDaNOTwzHHt3H47Ceoq8HvzgGY33j7TxdmFzKaCVdCfRh1m8
Yds6EanTWHTUyadLJVOjfTkh9w0+v/LGqf7/9j0HQgu2U+7/OPHNCSHCINi8h+wdEBnaPomWdNRF
h2iIVbLL69blCbHAP70mpcNHfM8U80qK/4SP0LtM/7PDu1JVApC55wdkjKEdpSxounTMVwztr1nm
NcCMq9AydFPLjG3Td9FwX9hHoMri3nxAx7T0UAVgxmva3X/U4Y+VIDyBrfCkqN7aQWQ0mni6ZExW
sCaOIBpyItrxZdXp2jdfWaAQxoLWwgW72C1jcJie0mO2vaoC+cfOfwjP3Sa3oLqBkjJuoyxJ1bU2
3cEm/pygMIn1XClVHJI9Cp1UmcOG9fFIPwCoA6/mzfGMjyH0F/Byvrfv+wqaC/JeLvwxJdqUv6xE
YvQgWWbSUSSFHc2s/SwWN4OFo2eO5yDf8Rub4ekYQ8m+GP12HmAJhHgKQq79CuaYeNpqx76eYT//
dAqhtPL75BpplvmgAlYmKRe/tTSxM8d3jGbH8NS5VMhQFrZqdfxtTYpBEFIDLICmt3/WjZDyIDTL
76EVEBBVTvxLBQVHJlyhp/ymNc1yfA/8YJqT0VUC41dBW/skh3byFfFu90sAvvsZZsDjV8TkMlsU
5aIMi+UCUMgGvLbXWnPuk/iQeKdv/m47p5qSaEa3DkIjkIyevYI7ZFGSwFgDiczh5WcX35Rc7rYX
CfNROcOF40JFOYAk9FtZBvmJPInOHTKZfZScvZpmO/5zqQyw5AKUg/sI13fQ/rg9m1D43D4ycsgO
u0DNkb2sjhpXkw09Btf2k96VJKSGF9wntS0vFJKXNX4Zh5jZpHAMXjywVPj3sW6e6HNI7ne+IhCL
FEUZGKiO2G/iSSjmW8vLFYj3VmJ5lHaCpXhltBxVgyb8IHNXfXuoCxoQzihiqBzh0hgU0x4ugZfm
RB9dxF0BH7D9iNoADQihFdG/HvodHLB+Kkz1S9nRbKzbabVtX20dVsIVvMt1GyPAQvoQ7r0b9k/2
F7xwjOvstxkK0Kez+7lvxsCvyS4xxYEAbFTKr2CAPqRRzeb9evzGWeCOKKQiQ6W6TMqamFEVcED3
Sqpy4BHRIgLEcImTtd5WM7Z5lO4+beBB2ozt0xBXJSXWnyl6Sh7l2k3fdQADFpnLJPTGxJScbD16
R17NifdN1OWE2fDg7O2dOVSuWfg91dOBvc754AdqCTK0mxdyHvGZGwVCDGKh6VDeTPbLiQYW8jgu
dcr31Zw8Hft87CBLA00ZQW8kXAZn3KYpFJlMZkjWKh8TYTjC87DL20ggmKHi4nHIdnRXaAz9h4HA
lt+/zGV+bAp3ciFQg2uLJGPBUh8NuwTK/xgbHPA2MzPhLva5YVG0DnsZNu0aorqR8KemPYcVR2Ec
oVBQxP1DtR+gfVm3+OdwsVvj/RR5GmNoSp6sfDHtab406VNGf6z9KJPME14VJgEJHJCRXb/A1OPB
uW09VHqjkZpaTHA42DhtCRv7fiqY4K0wOwxTTsnrGIPUE3HQtIBlpU/Ucl5OALH5E80eTeemKon6
qRwHxxmBFwyz1EGUPbj9kDcgFT2KWOTODXkv93fMfWHo6Bi4YmGFz67ho6al/QcRKr+7jOQS7X45
KRYjX9W5WqIHTinNSe6XwonXaZU4H209vjL6QkmNQ7QNnLIYXg8pwtxsBGDrCO77yCPNHOijJU8J
tEH4H4zqdTlL82fJ69/kDriD7eXAc0CoA1lP64Kzutcwja+wIxf3191Zanxj6z7ZdZyNImSUKid6
Zp5psoMuRF5obWlu0dXsOiCR/Q2r4J6LLjVdku2zRAtnLQv7skhNShJQ6WchaFrKoiec3LxfA0TB
5xkjbZNBiN/z/E9OzUgOoQ69z9EML3LvgtOXugAePS2tkttfowhgKzhNnoXhL6yQYjFaMTLWJOkd
i57R+jiiAv3gtsxvT49EO9ZpQNxMFABQam9f/anU0xwSVmSGwNw98qL1kDj1e+Q9FBkDB3VB8Oyd
Nw9ojGV+WMnM0MVk3tdAglMDV0E5wWxIv38SVP27tGjcm4y+B00E7tNn+Bodtpjb5AA9UXaopkJU
pjNbgGVrwun7MJB8Oh0aEuwIaTflRX+bpN7LHekqhi/DxOoHVmOHpDLaRO/Ox1XMoeAvgtsHVJop
6ezvzGbyVRLBMYYgcINBRC78bQzE5eZV+UfBSNnW39tB3FblgeDaXgVlHF96NqdrygmkiIcYZr+N
8BpHypDgWOGzGljNvLWv1qfRuqIP81qoXyGCZThpm5Nod8CsNSmKR82qfbdunrV6EQ5CaOlyPlqR
kR/5bWI8e8VGT8DBp5emaTLN0b+JqK5wdhsr7N8BMivb2BFKw4O8H6pu3NSXkM8rySF9SYZYY2Pj
ZEjK5jPtnoCVTBFoNUt8Vv7Or+gjrTfGDasgLV6ebbW4UvLksi19Q6OsFrj3mNza6CYtHMGgkFnB
13G85AzM7g9iHtac1Bp0AMzq7XqjpT/PG9YvezIu/dwGlfGFxhShjdbpq/+HSqpjp3wwlYajFJ97
179qBhhnwURCImCKMgKYhaMVZ6sy/Jnpv0xSxQtWE1+AVqbaVql9kHY37t0Lx6lp8xw124wCmHh0
rx6gvx/1u0pzPKjfqEVvCH1U/7Usw+8JjWFG+TFFJ+d+oE5OZxX23+htaezfFRYBZSb1oqxL4qba
uvmXoxyLYuY5Ln9s1cr3aNdajYaj48pJi4kwtmdxt+WYDxrfujor8qMuctIbzYhotB7c6yGMDVqI
p2MTqTIu+D/PVNNIXwRbpTR9KY+bxdlOMpIfjNlbGREJ9vKg34nbYpr5EdAg7jmzgYA09ybLhBRV
WxI+qF4KSaRs9olJ2+tMXIyWXNcG1yyxqPw3ZQS5WTOODHjc2COK5GlEcJp9oAbU3HW33eesyonW
enOdAu7vvyTXH9di1qF8UlLY8gtIW8qSNOImP/uX53pe31tRzRPDH4v6V4xrXMbVQRvCJPKtbjGO
YaqRh903VWAlrhHCmaW4pvU0jnv0QfB//tUoNozI27BYydSpvT04wyKMx2Gj5V52Lo5cxRZJ+SmK
TvIoehvtS6hQwaX2QSLsFwweXNqTnZ5U2uaUmrxLU7RHmjEmi7MWgoTgyfsf5G5Ys850PPos0UbD
Ir0Z6a62aCsctPabdD3vNfvnd1CdIJWlIOLF837MPdLCkdpnSBZv3SVCXb7LvOpfdk8EygQX4X1R
AueC9iB2qRDphEbGAAbL+ep+wlDkRLpWRoino2EUpqMtSjchwZYN7O826w/8HOWsRW3QNjw4Utgm
n7DmQTDxSMG7XbCKWeLD1tC1lK3+Qj5aoinj4WR7tnsLosLg43k30eL+FzdMO/QXUXUzYSi+Y1jK
2w/u+YFDwtv87kxf4Mfdri3mQIZLl3k0nGCvdJRZYvjuTZpzo+/LIJNvJxN1xF+sjBLpWI4252rB
ntqBvVioGceWT04M0GgitgfN92AjmnPiaYSbh4AFeG3D6xrW/b2iDsX/TlMD3h5bwUXKIEDhYnpF
ermbckxPMYVDde+W4N1otIVCiGj2OXOP57+V1tK6PPpLXSkSNdsiFF75jOrRnokzDZALSU+7xYQN
clz1N2+DmIQvqRNHd9oMeFivLDhFgSjQsDw1n07uzEsw3XwPxkmDImCgluLcoNT6HS8XRrYeHEXm
Lqhr0Mj4APIRfz9zD8nV8hlUQ9seGh+0wwRaXNMVoZty74+9hSfZxwx7bDLA7imF2otTwOABvNVm
YjH8Y9JCJMRAlLb66tGZFCYVkcTLhFco0mS9MomfAS8p02S0PjzsfhsFFA8BICcSLH/9qPtRNHez
6YH7lAZdF7lWOJyuMSdWWoyX7ktjhgTtWX78bhB43k5yGAFrxQs34clC/oNPnlJo3JeeKWSb5lsC
rgOO73MvNBeJBDcUeX+ABdnj6+lJ5xd9Mj7g2uy5tY48nNEVCVcOcLaRAm19jO6UC8T9YpMt+VK7
50eDhbl/JOm7Ye4asusm0fpDa92Sy1C6ii54Pv434udqWkZvD1GQdT7Bw2yGh6bYPsggxnX+6oQ5
1b7y/7xSya2RkRT/BE+Lnhd+e0IWYdRJGYjm/WwOCSFR73PLm1PznzTgEe2rHjytKXtf0mhE0CC+
ck6rF9RPlESwkE7hzsYquW/R7re7UCDT4KzCSCFn8dV9V16HNR05I1fTF60CZ5PD/eHpgh0eZb06
D6z2fCXWjQddtra4cIszGdywcGmAXyYLmVldjpHkyWi8HrnemauSQtKRcOtiF4Q96oIGv+o3ngfx
r0esKutKVddu0ssvCAD/EXVNW6MI9evgsM8+NaOjUvRCcUjWXIG6NTSC/g+EGm3+NjXZL/wjCvmV
gLoFx+qP4ypGPAMTSxVSUi+Mz2xpGIFf6tzfx3l8Zs/SBuTjh33doq+93Re61t0lXATXu9dwhFfH
VCyxeACkV6ObmJ1p74xRZVg9hbQTdI/cpaKGqOk4Z2OqUGIEkTtpSA6EDE+m+x+UoT0+lBw/N1oS
Yr6rm0VW7Gjp/GUqsKdeAUz+YZy5/WCvm5vQd6WcmgzK1VzSGMjP3j76899NgWtvcCNbQGY/5uMb
3WtJSZFfypRxE3DEdkxYOmwGPWj+sSYy7ml6QOBHbP3whvamI4WV1pDhwxF2YGIMSXH8gdlRH2Vp
aQVya2BPl/GPX/9ATP30CQ/8FjACKyFXFzNG/agb+3HfQjPg0eeM+bO62kGryx3fjTVEWASy3y1D
KcdDCoY5SWYkItUh2jA6rUmLZC+2eXUfS76i4X63v4I0tGITuBpl3dNkYwIRGBFfk3CmpbzIIuPL
BSHKmhR3I8Fb+y2m676KcnlCrVX+SyskAGIcnGRhUqwkJSV9XL+mVC0l9KUkbQ7+NvrpJ+OJ19aX
L9UHobF8QGWx5RBPWhlM2yO4m6w6pDfLUlccB7zGQRFk8KZLoRyJvKL+T4AQPobtkF5Mm09AWkB3
E7aY9XQOztzYZLkvUQVyiN9Jn288Yq0hwlZyLq8TVRqkh3XJDyFTbrWR8nd8YzNPf8BVbwuhIvPI
SCUuEgGslTHmdKAQJj2I3Rmx2nl0koeFozAuPUwl0D5ZCb259HDzihiNnkUj+0ocduM8TXKe+qux
rXDA+2m7HVZecWh8YwHuwiMiVn9uirTSP+VcKMMNWBFUh8QVgi0j0GsRiyt/UoJ3kV5sYEp6p9qj
UAfRsi8YuaOhjqaXOHu/t2egnaEHGzMU13OjxmIgyBu6z66l4iOyXMOd2UEtCICsBEyGcxrnXQiv
K50idTKoHV3THJSyYntcubeVvmUk3qJOmoYznRCwECJ8sHOPMIBpYT46azWO3jFOdaPwwLRw+HFB
tVNiQffeAlYH++3LXzhQ2jUFgEXH/laHnbmk/5qIuTF1l/g14bIW/OpNi4wP7aHU7le1pWazDdTN
r1vB9U069jCHUPAbOfSOFinENa2k46XrCMGwpPB61cBs6TFabKK3ff3fn8jwuZGH+qQmqmXoHlc1
rw18trRcrEPOTFycAslXg+rDkk/jcNbqZeN7v/ibOrxXVw+62AveoasrlnnUS5iC6/RZxdtg8+nX
1rzwV1NLqiqzxK6LQousftzGHkplVGoT45+hXNiTO6VWkXnYGJuNr8Kxik+SeNrfyNhf/TpRw9bK
00T6CLm2boiKIjGrYsqB1esc8YUZ49AJd0g+OKfDEcZuPBpg0XS66TgHM90p5GP4Zw6SRdvQYCF8
X3UZxGXSfPVtjbb1YpCX6rBMcM1G5Sl8xR+BSqiI6gHiqEw4mX6/3wQy4uk+KA5a0CAEgovKjOCE
ywtMvN0LuLFgQ0rmAfbdOvtKbJsWB4B4a+5cTyUqrvcyKg5Dy9D05wUZArkd1fhf8VkH558t4z/3
+knjQ+hMqNAjxv1i4s8GIWYYQK+9RzOaYVDSiq86kMQiBItOCfhPu/avSAyYgVRFnC8jKF06pakz
F/vTmexaBJVBnLNgopIGvKUZHyUbPOrGEx6aSsXJo580Y9Mift/XKVlFWQc7UB0i5i+zWxpGJzwz
MosgHYqfrO4OiiV6th6EmWBnwULN4ghCcIXrKAwdQ+mFkQ33xsEiEELqtLwSPJt9G96dwYaIjP80
T1ICgBrYT00SKG8JvgOzABBcDuOtMvdWkHeART2VQh0tvPlmmg4/SCnDQXvIMF+HErqS+0tk7O6k
7lah+bPFvbR9IxBiGw/DOnvMs8XBdwwqMIZ+KWDJRxgOkWYRWRgmYBcQ73Iyh8J2cTqwcOfXD0tk
wPZh/KyXGaqaOs2Jp2UvJdgXhjihUwwwj4Hle5A9TvXXLaWLnBs+VrUMyFhlEBmRCt73rD2LWOPw
OmNcqe1imqIrMiWXM9H66Wqo638jLLryyRFGjW2/PgvPESn3qvlTDo9M22IIc1f9g73qypI20goy
gd7ZXqPlD1ggt893O2J5NOdBsQOtxVy+TOP6iiqNpsP75oN/t/rc4AMzkGrAG4YEmD7gpb91kiM1
GlJq+I7jf9JSdlDI3wa7N4/JvrNTUMhyr0wZmiBuaOUs0M95L2b8Heel7EHnhFLq8ldtp6H+EI/W
6WOkWpvLvYBz9YwzIPVB8zNecGSOb6fZzrwCqUOM4OKTlwF/DU4Hb6Ia/w0qGhn0FK365GVljynT
S0H/v+j1/OTHMeNzxcJtX9LIAR4oz4J1YRme99RJbtEdQiHNCQVOgqtKzKISnfmdg43ZjozGtETA
0PJ9KZ8Asg59231HF5KqZHb2oohw1KSg9lIVCHTE9i92NIS3ftVYYWpObD2DgwDaDGJUHn1yVJNr
ITjpubz6nVrtD+GTAMH2EtLdDyOCAjZumiXvhV54XtzE4PJF+JWQPnX5JPleT8DXrHfF489NMxsx
/NfmLHE+J8gkb6WDmu/WkIvxIg3EmV4yUK2p2O1oD6/niw28p4YEqT1jx3Wom5cuBdKBV3Yny4A0
caTia+Flot5LZZaYYvj7RGpoq677/yRW3OfSXFjk3QCYwr1L49gVCNSvT4pznAeSMq1h04DzZKtB
P54gpG0unwVFhKP6uYyQlNGsN4cFRrIhC1Fv4NjhFNwTQUw4jwYi5L2d81nz/Stb+sROmDfLv9Jz
oruw2nr750EMm5UkyvT2iG5DTwH906aH8ZkrpiSgGQd8C0e3Ovlh20UC3cR3OPVJzEzYVHnKxmwp
BYHaBL/Vu+fn0s+9WCRq2zpdkrTJTQ8qY9rl6E0dXqKCwea+AFIAcTpE3s5Z1304E/Z3UmGehK+l
8emAzDPyxHrri/Lh32jHWL8Vmv/IUilV74m67QKzqHflQra9gYp2bUvuiy9T5r5a2pernJ0hDZe1
wSd6BrWNOZIUdXoJF/9GiiyHars+Ikj75di/2NNr816DPsfN30ARdeS09kuIeyQjrSXv564HA3M1
phgkSFFwXBVeJB+clMeHhJGvuyaCUntB8tPJLtjV8Pp862pvBwVU+K/UXfgCiULnhiU/asoR3C9l
FpP9YrPgf8XGV+6pGgtgXF/JQbt8QXy9PpY/RdDsuWAD9lVtfrxk8jU7wlUw218z9R894ppw+n7a
em5LClK37AKG3OWQyAEkpJ0ot+NDa+fZwRjvP5a3httOqLRv56mg4rPZEEdzbyYNr/ZwbBwcRxvP
IV47uXcAB639sGnLwN+Oa7ctec/UAjrgGWM15sydg7MmmOp+JVh9PWNXNzXt6MA64/yuPp9lQ+Mk
mc+fSmPQAgRa70Qy4TkC2HO8TKKuIs0w8PHxrC9Sm0jtL9vrt1S6KORlero5yAQ8+x4ZrAs9H83r
2t/tfkMFug2S6jrDu1arRoTDiyjd20cJAy7WWtjKc4qpWC0rvdo4pOFNKFZZ4mhYbXYQ6vtUThim
Y/jS0bo9oq8taCzyFDmNDcRQkcXtVHFNQAw2VUF+8wfGdG+rC/tLZK6plsDDTa/UwVv+9bKSUVny
HEhT5OxjnKmM+ZHihMXNPzBMHp0aLdfif4ihC/0QcPX0KFKFkFMDN4SvC7/KDmrZO1zf6DlWX0RO
mOJze5UVQ0qr8ZuuyzO4H+EPyMJI/KWkoOWAtdzTygIhqt3y6SI2esnEyLabSrSl39JmUXdC9rUc
kZcZpZilr4J/kYSXXh0L4CjfD12EwtLVOzgxEFV69GNcZP8Do0eI8WWrJ0w0fvFBVmmy9faQox0R
jj/NUKdrS3SNxqWlio+dOXEIKM19Dc5/DLh2gYcBGuGt1y2BBrhT+FhmEOEyNvCGxXh02PsXnYsq
ekE2QeXJnfBpHwddDyV3tYUYUav92/9vUOydHcJfSagXrqff/4CtIFm6jLrXYSWjS3mdfRO3DyN3
bgA+Qg/ugdnG5u1TgCNvpvKPbBqFUff3A+CqEjhjAeViV6Ioxt9IPPO9MuosdarNGNIjKWqsuVnl
bQbH74KswXt86Qi6YeM/7DDqG5ALE/rVbNN64Foihsl8hptLlForVFPNzdDMe+gbzdM3Hd1wzLc9
t+XbLSF6WNKWffPPjKJIYP/VgNqDYTJutFbzhi5xypjTg3yvO6koyZ80VbZ7IHU/1mW60v9oo8om
3dizGbd9cgRZCHtj7d2QfrbRQvoXY0K0RYFjB7vIodpXusoTGm+um/2P612oTosk+uz2F0M0h5Cv
hkA+qhGE+opUsgm3oNNZcsIqGXPQKkhLFuY1+m0MkOcPhTA2pjwQIeUV+xrP/PNnBSbC5sSynEMz
tdVGKUIY5VjPi8om8n8mrtaA8tnF/XoSj+pOHL/yqrkRBnRK+hgYvOfz5JXw02SpQDQuMlGnAkzi
y0d2p/srkugZ8s+1/+k9v45lhhMUUJGrcxjnkahWcaZfELZaNsicN8HzdKbcb24qvqEbtiCLSD5P
KInYPUfWlC6WU7+cVEtIow3v2KmyN5gLnEM76/3nLy/XT69/c9aZ5dEIGR6JwyFFpkYDpbICJPzI
kvFKoSy0q0kkUE4Iyl8mMFu0+HvUaWZ8g0N9Jt+Q73rYLa4GXAajbq3YtlvONyDetGPfW8uzQQrr
eBuMUHxJKXo8p8yW9j0ZaF87sryBV26Lbiiw7AnVdJ3E82P+vzjJdv9HODMYvc7Sql3Fdh7FXCgm
rPsQ7xs1P5VO7XejEXX8eMDV++jhVZt3QmJN4m5ONoes1JVpZwRDO1bVkRV5BOojqg3xQb7/+UYm
4g8mBd1B3rax7ecvjO2xprZpd6ojGB3SyTK37D4KmiztVwJOO5T6gmL/G8HlPhIbOpSd16cyxjq5
vhYK2dDf8CegWOMAlk1BsvGLACRx2aqAq6khd54ZgCj+xlPYC7KQGjlIC30mBsmPUUouqlATUm/h
eKHlLP5t5JnzVXMotKXnlZs1oOhhUD258QD5rLG4ETyJ1ZnSdwhej/IxInjFrX1YctQ3QyLYnBGZ
nvsAUkYw+Pbshebo4h5kux52yzXEu+xwVL+42BiGMWMR8/w36BL8jTT5Ff187opJSy6XNASJWJFU
sDd1P/+2PQfNl1K3EmFlBS4lrado6xvOEZgddYY5n5KZqgWAtEUYSTgePikXouC78/TVBGS8VNCC
UlBgPkeQsAgQbOuD3B7F5Nn82ID7My1nbNRf2ZMT87jktgQSpeOafmuHQzxcal9xwJ6hdjj+CeKQ
Ik83g9zekK7yJmTgbHtpYeDnT/cgsvyUeGOfPp+Qy0qh2O/epSMrhiaCDe/opCXnU9Wy455JHQN4
4Kgtx/KG7UiE1yX5NYQG11eqpSF6owA3hzBTiJVMN9hOAhm8U7LCqAbARaEofWYQzjb3ZdeArn1i
VezLK9am/5wZbbOOoBoN6yo3CTTAQP+rRoNtjK5MBpyhdDc8mARPwjsdACqskULDii+3hTEsxkdD
gl4F4D9HY9p5iK61eIDKNLJeD+QnbbGunVguBz/NBk8IvnkWbWXP7wlwiYlNdrt0VlUrNaxIF2pS
vcioH/cs9njlOS4mkVt989kpi7qxRtca5TLNN+9s5NHS+7V+0CDM7f7W6xsHmGwa03nPEnl1rkX0
C40C/VwMBgGHJ//TrgDdSy9CYCOZ1nWz9blPJv3MtkpVUHxYUD4Vxy11SEbQkxbgZOPatlPke4l7
s15nn3WuZxQQRIUEUtZH7mGeXpkVnsIw96nf8dkz3CXzoOprn6NJ8xDcl+fZH9Jd1TF7Q5AB4HEW
I4VUFXC+pd+Zpu5rlI6OkdDyg7cXzKSBXaMoCViGUe6j6a+dQw3NlXUU/kCViPoqqTsCCdsD3ZqS
6AN9vlX67mD+XtCHxF5MxQBqsyWkJi5iJ3U4WuSUx1iby8AsKElD8T3JMReA5b/H/NW24rjCW/qq
LgaF7yqOHLDxROcciI9oIVxFArlcP0lO+zi9TMQIKu8n1oguXpTgfXKd/E89LnX69OnXELYWf3mp
MjnCngHbpbimI6pm0uzUbBZaCJkH9Wo42S6eTMxK1zad95p/kMfuhTIQ8YfkcvgJ8lN7JaP89yUZ
WUGP/U3rxufx2J3y/5YXdJAroiL61w4ON49XC3/T/SN/U+3l77NkAf9oRC6AkGmWHBQUd4YpNjBY
fx29OnB7Rkqa8TP3do6/WMIg2Dv8zZVOrDqBxyGuHRuSO71zaCFsajO1LIjljG0fgaEDyU4r0C7s
QnpbLOG2GhALdFoVtXq01KaA5qUfHnkSgjwgr5SNXgZs6ZZ/ViDU4oiFxjypNoXxF3kjiK36K0hz
SEN5Qk0y/mWviC4tghLon7P1VW5+fugNdnh8Hy21AQGsd1A/WxYj7s/y6Bk8DzMK41/S//GWxJJH
9i3TSbZP1hCB+oJq1FMLlXmQg4rFrZ4h0s5XZDjHOPgX+aiCMAO5CgwuIkBdlhGoO8ImtByVHglJ
NYVPaId1bU1yG5q8xlFPW4GVmUyKVsxtvWTom2ZpY6tN+y/wddg2kMgVDxLFfI4EKIQxlGLOW/ZV
ROdjqeAVgNhPBtwwOC3z+PXYAt2U2xr6m71hdtq7FNu6O4UtL8yFLBC5G4UmIHTycWEkXmcoKFIE
oog+qq+qTq6vTfPBhsVX1YwupeqlVBKOsnSTI2jg3JE6SABxj8oY5Cfgzv3biUWTNYP3C+IT17+q
rD8bY1lv9FoTAvQiR8A1wBTJ+SK0l0JS/BliS7MQe643e4vh1R59BEIKa75AScrJnH/wcpyoiyx5
XjpYdtsuFa3WdPfmWQjvQcmXJaanUHPf8u5A08Hiw0MqiE3xFWdQVGhXA/0stWfQzh+UYwgRGw/S
ljWYkcTUOPrJu+iy9l60m7bllzuN8zD9UaixM3F2BjQY3NW16J5Ue0Opf77KsApToxIDHqwv9Vuj
a3mW98XBvu8O2YuC6UtJ5N0lyIymTY8wfz1bLp1VMxM7O52pg0U1ld7bYyz0EmxHQO6YcucugKv6
ZwVwLvk879jFJ11gpPLLB+zeTTpxnxrHJzkHHfJkfQZ8vF5cT3apeN9lf/FZnFUgu3Y9IfL6H99A
AGd4/JwBaawJ5T4VG1e3nHDlHlcUeJBgHI6B+7oTqhDBojUwtRJMGAsEQC/QwcJkm6sMxURgcCLz
STgNJojZeDE39SMyEahsZER09v+DFkjUtU106LV+V+tRBfssBiBqXfZXkI1RNndIVzCVwY63Oa5F
/kkXriR3X+1dgOX2nDu25P/o1pn1+0ZUPqnXZtLIs1/01nqT9WCAJKkyCoKfjwNAPDKWw/LnfHkm
YRB1699nSjIlymbu2oy3Rx3v5khsNuRJd+t21ysrWtuDmpOgT8YVwEU/B9fx02JaEEX6zJlQyIgb
AFpFDRfhn3RnL2gnWxxwkmXO/0ivRs0Ob3WDkmMVTnBjkOkCrtvjztIi83h01FRVYmy3jOQ6RIJw
NZDqUAfqPklAZ04XoQUTGTX+pgC2hf/ZpxV2qzwVZNUpSg9wt0xtt9YKEzdW5OGFgy6ZWacQPyXA
G8p+xDcaQZtdYEYrMOEqItdls4d4UjaNYhefIE62acrtjG1uiBO2vsQ3V1QO8fvoDBoZ/WQ2WIUf
z91hGBposjDDWf5TUgqXeiNzSLCP0SFAWjMqYevISt7aaG6ksdz2G61SNBXbx/xlGFbw1CvBaDyC
brjxa6vRL1R/skVD2zxvUVW5b9tAW5rTzAuJ5+SUBG/XU43avVjq7ln3dFlzNiD+Hb394CrvdW4L
4LiCVFSoShHQGxXfE8pC9glmW8PnBXifgGGTefTuWZ6wuqSJ5/hcsrUTNg4QsCiePTWXyqV/Fm33
/nMBqatc8/wTXxfGgEGmUNVNqHILNAZiuBjIqQqfdzSJnXjRpZ2qnWpIiL3Xr9PFyVfsXX72kvX7
q/H75e3XvSHjVIB9shFh3NQQNosSPBTBrb6tG7UYeewKrheYcnyl6ladcKn7VfPtdjxCv0xoDac3
Qberg8gjJyGymXJ4K4XfKm2/2aeMI5xQe2gQCrQDoNwJhrU5ZLF1W4mfrPF/MRS/GLZY865djs1O
uESghokK50vZkf5aInVLZiooZ/zQIYkJWy8OJMp2vlKDXQ+m4csFleRMH44lCc1OAxfJF20HN+aL
/S277xIIaiZSW5LpLPyh16LUkatHErX/PqnQF0Jb+v4WY1xI5hgH13hrWiak95s2+5oKsRvvyEG5
Op2CGorRyTGZZx9JwfLpmBicG+w4OpgcmNwTAuyL1CIf3suz7A3DvwG61TZtOI9vPjY7o8uyAk4T
IAiIfpKLKIfgP1kT8gsw/sdR9fKoVI7UXwb/qkWed/OpwcnAz/8VxfUTGXq4t38o5vvOiePf/Hx3
Ir7nE/bxqraylqpwgmliVos6yYy+nHKTpGXxjCpPzLsEDifKQZeUIqm9iRtiDFNbC+gyympSSCtz
WSishXtRpW4aJpnHbv50PoKJzdnRsDW19n9u+BJHQGg/L5jmXSml3Yk1ulA3F+3MSRmZ+OkV1SZk
G6IMlqhlqvrQDaaA9jqbpbN9ryqFu2irleACb/RXo2+OUt3Xz/XOFuMOUC60pZJDk6tTfIM28D9o
J8152X3FsNbg6NwXjru3oYa2eFOeC8MujxMBOpW+nhh7DK6Sj1upEHpprarswAkaHIzyB9VEDRfe
4yVfYBlv896gZ9kU2pGZi4M4tmGwqXdisbFTZtj/NuF+Rf7CvrArOTxZE7F6dN0B2nHVG9WGGy4L
UzG9jbEQp0YrIBLJYcGOrYt5CdbTg9Yc5lw5HPP7978ViQEFHjrG+BuAiBsQ5C/BhQZGVVurTCY6
CfiqtOH6Bx4hPHdRV5La97piSZA5DAsuLtD3c6nhgdlZMoeZUCuw0GQ9T4h3IGbsaGHc+yZuoQNI
rhUQUqPFQLjeF5ek9gUjKetNF5wr+frb6Pi8Cqq/69z5fFQU7O2/QGXpMgvganmXScy+SqnH3cV5
4weiACl2OtYLLPo+x2267O5/1KHHFDfbycNiIvaSVe2Uhopwb4JfBVojONZ0Q85CUTzfZcTpDiW5
Z7hLUt5pQny9rMu2ckA+tnGL7pgg2+X5vYcpmaHHbNZqHMb8wysk+xzluxiMTnDw2R5OwFKzz1DX
GLUrXuf3RlFUedJ+g/s6JROZqx9WyVSyiObvNbwb3KaGYZ/O9fHDnAzLHTWKo9B8CSybYmHsWq1w
zDqRFOXy64o6mph0yDIIawNP9DyKMDq0t4LNVhE5dNmYfMmiM63NIf5IwLMlc5Eu2Nj1fsncqr50
YmF1CjnsaKP5sGK4Aq0BMJNT90yUJNc65QuETD7foQjd0QJCOxd1jl1n7U54i0HlGwV1H4No3f/p
bJwuCHpOGDK5HyuxSMiYjm30JVWf+nK3k8oeJkNXxGU1VAqZC4FIZbyar7UhD8Rq/tiwjqPhY6+D
Noj/nH+Ixd1akq1TRFJz/Rnw+LB2VkPxdwP9IaOdO4a3/+HvTFOtqLAl3Zrf5FrbDAXamAUflVG1
tImj5KuHGqVRAm0l2VE8ra942NLAZotWAx0o5Jkl3t9bzkXNqiKjMmGYaUW5ls47r7VGQST1aQ51
SyxzskYoTGpuOo8MjPTgFWp5c54eIHRwfwehV6V4lV6mYXzMDG+Xbi1nF59ZmjpA9IbZQLBNcBpI
wj2U20sRRbKtY95qbD8iElF+ZO3MCRHfWY8RG+d4H680pAxfxHNFmVnGGJ3AuyTJFf+K2T1oDuUV
RYDJJ6GiBKtTCjCS/CLY3UjkwbYIHy66GU6yHnHWvsv90hlQXXCYnni31K49X2jsYFsisCMTVH+w
looJfZmZYzuta60XOSe6P2NKM+qKAbrbUbVVr4mdXUZMUq4IJJqkSgc/WnPhv2VtodvvrVu3pqAx
gT/1c7wn0RNES/JgD1Qax7t1HIogPatEM25jJlF/t0ZeqlsVmtHgTpuSMqdjyfBWdc8Yzew899Ic
C6jRktG/Emy3zGlGFp1rnMaFsEVaTmw6i9PtUqZ0w3hVf5gIwekYsdmBo0/NOsjS9RnTxqo0tFBf
XZnULQK2F4LAVl7wea1UwatYoCLmeN4avFBf4fLm4hBa8McWRfAQXt0RHN/AfTJcfjJmjchZne3B
ttxdqNhc2lq+nr2VOxJOSPuebDknD2CHPzLzAeQPnVBN3jOht9NOTWvY+5dwCSs7Bb09cjUyAPT4
l9VDvw4lYx1o0vb4AbHbdg4UqgtDLla28DGIxjXbgHbFhlVDemq7mh+JVMfhWDxnueKepQn18vyf
ccjznuCCS7xCRDW5ojJz+c/xu7vbRabsuL60tcssvUwSevksBA1kgsv9xBxDbQUE2j8TBqXC0D5i
V31pCzS9FzCfwAqePlhLI0/noZISAIyKJqa7wHMbin2uT0XDi2k7XHC53A+gz/DkEzwxFYUe913y
+u2+Vb/TP5HgE7K6/4RA3MhBf7cJCprA9uAgNjc/JES4StuG5gMoS3HsDnbGlyk+0xjss47iVRVC
WHoe2MJlGD6vQXiU9fBJLpBw9xiX+1JoxGaQqAvsdiRVAqc6nOzZwJP9t9TSqrdoDs6kHIjnFKwN
mlMSfphYiEVg8ocTpZ2+t8RL3zH+ltSLqx5MboJGQNEQQasTg4Lm1qtHId04QdBYG9QiB4gLx/ty
Wm0vIA6nNWEZ/YqtSysHqJLfDeF3S+f0OgkMySZggwNRaXE22Dc6NA/ldvBi+EWsv9hfmj3D4Um0
gaBS9gq17jg+SI3Vm5CiLEiGo+gKR1A8z7yKFZQ6RUYMBNRYDbWQFga887+2vUGRIOKNIkmsy8V9
xMUgnXbW4FNa8Jvaej4rkVIW03xHinYg0/Lmi4FaPc38Saau+p6VfrBrxt93mIlsVvdeYBuLfDxD
aBq1IbNHLpGu3CdrG47B55OXwfKPjowX60+4X2s5qLyWX01xMT6PKZoGsZALBmeRDWUTdn2yhLH4
x9mWKw0KgRvhHgZyThAGRqs+1OYqK/rAQiFxn/d6fHoMbzO7lYhr225Qh8X8ZOMsvu0+oJeYVrGN
qmkLltK8boMZYHIXCO0naz8u3Q4/VrJuMYdK1ynzHBm4JOi/JqAsRR+DpZhwx7XDvRTWLM9Hpa7d
OG5HxUfEpwvnJE7uD7h5AKMfdIgJ0133vh6LAJnXGPkcKQEaQwT+JqoetkItPsEisbJyMcTbs8/w
3FpKZQ9DKi85lxJMKWjcy6+C1isnECzXw3mASedKPGfhbsqHO5TTtthqfqHbiLyQn8CzhtXjYAoR
MBG4XSlB7z0F8mg3CGd6uT9Rg/6Zg7adIwj/3MW2nxd3igqo+b0Y1F0cVgN3QSbu2U7cPGkO1YJk
ouVETogeOZPCQo+X2i0i4Pf4BZtsY9+O3Xmxqg77eSY+NDcnjXG0X5Q8H530TJ42fKeUKoFXfwwU
V8wSXE3hmLZYPcAhhs519ZtX5W2mVtbVZPS2O7WJePX/XS5UuUaGpkOjWt8xS5rhPthCcMPrXEFn
Sh9kdCVJUJS0HutJi8DQfKrUF1v6bbIZbCX8OtffBJuIgBDXxjPMcMsDczBga586298PCM6ostSx
iq4VEbmBVHszWQFiRM5NxtS57NH33rbMh9jPhtwOUQVorfGNnuL1l4BwrmRLlO6lpUqNTEoGdRT2
cwDjYw536Z+88xY1re+57EMBkiW8zGcCMiW68mG4ZaHIY1FCy5Yy7poJ+tQLpW1vCjq3QpVy0pmW
hLLZpVrabwqBj3flFCz85sZU2rWPTSGjIRePo056GdL1PbDBUkAYsfoE9fbzBL+XKPss8nnT7XBi
EaRXovb08vy50mXf8kSbxIwF/IB30/S+pxKFpItzBRbtRi9qMdzyYhdUyHsJXrGU0tc5pGgY/KTX
b79dYi+Wil4WSq7dt/8qshod3FeIWWRpD2xjQzuuxCOVmGyXPeTs423GaNTeZfcJ8Gbpqa0Hqf2c
/Nkgcl3McMffHLsoMngbhBCQ5opEamzyHkLvsO6Uwu8Sp6fPWtS4D3tZ3Y5rkiuC4wWGMNnSP0D0
5HgjvaoX4rDR3YzgoNwt1E6p+rW0M8buiB+9ENujJx+S6XoxSuJ5kYRxnF/x5UiUO1hI+NiRBunU
E74BMxhzkc/rm6dQMXNANAz6OGbQF0C01XCNhXwrO0ds1R9z4sBIIuF4PY82SZemVTwRdCmrKQpd
tPBCcrPsb3xu71vhYr7qISCeDWGbgP2p8shWM9ulhUy+ruks8pjDhBMTbCRd3z58Ms/9BMwNPe1d
l54do5KhOv9RcCZvOox3yEKv0xUNGCHgMfLQjK3n/MYPBNJOOidKxPH5wyiq3HJzoj4Pz49CpZU4
AVFrLGi1LWaC3IrsCwGGzOxyG/AjagElBRSRqxpc/S++lZ/k0eAiolbgjofeycKTGHx/SoujSsZ4
tRCH6eDUOvKLJ5dWdtTW8IHyssv13ZuEgn6JfhNfnrliV0m1FVtxRlfrsADuqUVtCEmO0KwsgjLb
/7UgV/m8TewoJtftACmMvvhjMhBywSpHLwoOF6FfxOxQRoFemMhoQosg+fWReCCPPNbKl+aO+RnM
zx491fH2QsOzUegoeM7uIOLMAmBQoRrZ6ZcJT86a6hrSpjqC+eg3YxgZ0+WpYdEia28hecdEVLoU
hSu6RMTCQY9w9kxsG62Th+q/LMyx/J548wLeXywlen3doPl8xZSCVGftDZVtwV7I254THVvFBWqB
u8jyouWDaZ2KrBv1+/bsj9LqHzySmfBe5kIoyoHfYJvicAHUCcGuN2vStpdIKOL8Q8A4eSjIpRpP
dYmW+103zzCTi+1k5tKBK0uySsDEJK6006V88EXLx9FOf5fX16b8zXltfvfX+w2If7oRC21Cr6cK
7VCq3otiofj2ShM0SHzMV3uMwU6xoLxNOWoRbiFNJ+NvBZibsfkOy/3bASERRRE9u9+iJHTxQ/sy
oaMotnlVx4ob2Sh11qsCj+QPqWS0L1cJoS5AseDipawaPncjtV/mFRLPuBwB7XAV6gotPSUfBVWX
A8qveL5KHVm+nZ0eMnc8zdmYWF8xC06FWUIv2oN/JCFHJx6S/RTf/bJS1dVWXKuLkXX+A94MqWBE
KtGAGRaYNq+/7HKxOrdFQLNepR5ptXctYvWhKJIHvyn5xicvjyPQBPhMAosw0KLDxa3NiwNRWRVJ
Ng4wRLZxShkAy88TzlZUdguZM+BCP4e4+j8VUOtld1sZ2cdNbHB3LG6z9xFSx3kFGBnd7hwQ3j5G
WCLmiRPlKyj+TrJv40WdENdF2bV6o3NwGUsIgbJMNBBa98116fHvDywYUqGA65lx3r6sXM65b7S4
JrZp5OYtiX+dfur3yW2PeVKIEOn2Erl4rrMyvR9SQ5a96Rsd5M7wnPI0Gt7i00kR5tM5hOACJ5sl
kHYjSbdY/fAouMNa7bGS+Np+Vrpc6agtGXEN6bdrDNQLG2cQfHY59xQEYIU0YvqwIMvA/Ch+mu5k
RFP/eTyq2rSEuMU3CN8la8qZJVCRUikO54In2fDcmAkpOxBJ8Xq9/HR8ldnMTKQ7rsST04/z0BAn
XhJXs1a9NnWi1k1F121bs0qtSr0BZQly5Tp2/8WMcTURKW/AmL4tOZVJxLJG10CpD4KygpKTD69G
c3/9xR7RkLjnp4FmKJQ8yBrMJ1Fxt0hEPZQmpyKnJJXvkHqAF4NDUsTlIAHm1SOv2pc4V/vb+YjZ
jq0nBlnCKWaO5LBJVWcEGxqeimQenEN1nhjj91ddn/JBKt+78pUsZIS9VPueUWIW/pOSqlnD7+qZ
AaFZX/Ac1fWA4Z5Kbvuuvd2wdIDZEdsqjgurGRTRZbrUudwq1MixwFqhWGalLPmFPHjU8PVa3KSf
7k6x47JsmztTwlnQEHPo43wZenm28pxgRhO6yiVkTsH4tTTtMACZj+44y3og3xUrlHHgvF+5pK8X
S7pQOPGmDCzxUV74vwGaIsBGxB4UrwdIyMCq7IBOsxU0Y45w6v6lnDd5gl+U0MoQIuwiZXgYScNn
UG9pv3rGYRNwZFvyh1CihcuW6asxsN2Ft0LJb1w38/usSbJzp7PrzYefGcQwQL+Em5SDa8SRO9/S
nb3ssAfHUuwmibGnyW8tar1R17y7uCS/dBl6CIOpgsLHuxBPoT9mz1pTos+lsdizNn8guQbP1gp7
oyG+I4zYS9WdNtng7+/hsgyLUAYb9ZNxgkY1XlV8BcSUd2r6omnbP01JbrOmIXAxexwhmSBuQS+t
8KA37PyhmuTCI6Xk9hlVxKEnVtAxYew//oWoVEgkt+G2+/l00BltaCz9TIR9kcKyDbWCU7P/wsf4
9jIgivFVhtAc3JciximqrgNE6WGYdptbNkkQtgJmSNcEp3eLNdNLXin1wdToEHYELrkOmTinCxKu
4db2XAH3xn6XDvJvbIia2BT15PChUilsi1BAwl079q2JuHjUmIiaW+yetztSpjA5qw96tYL05Sp4
cOR79/yTC8TQFgOEnT+VdhN8XF/WSReS9gPQRkHlj9DytInLMB79MDQd5FYIY3DdP2j1Bty34UMl
LCV8MJg/0c3XhkuoX4bGqgLWjSrp94bnegnjO12cqvhwAa7qUiPlQmIvFeeZHScygXJ0I3koK8qz
rBETvBgD20+4421O1YdtaEFSlDRT16IryfeT4kh4WoH3ndMRyJIMDzNGn+EoXzwfjeU9EdNpwZpW
LiPN3Cs2WxOmmprKW7KZHX4YNfOqsV2O6vkSltcZxVPN2COV/H11HFS9iGB2E6LgNhi4j4SDtL99
sJlOeTkrTkRZh66iOma+adt8iUKhR5FCAYLOcrYlasx3pD/lVBF828E4YQf6/9CIBkjlLN+/Vn+l
FGu0nCeOSbTtTv+Uc31tTGtkcNfJKg9nPl6mrb+G9TJlPhgxfEKRMQVJJ9wCrzdv1VSGTBS0TEZ9
pYkOsVffX33d7wW2BK7WO2wLKVVC2uSLFZsYEsG0kcSbrocXzC2ItfZYMzRjl0FQHQkxc6pG9VXh
z75W1PFF3OII1//2ItsuEHY3Fci+20+oGQgHGyIkc8TzfcEMB4/KPOHHim1tMSQIOe4nLFGt7dyF
s/1hZ2Jjk72laHV78+kkYcaNPofNmCkq4vEM0DDAuiopJUReQDjV4dKg5oHKnZkWTpMgV7bOS8lW
0mNG0tZqs0SFZ46SKba7JSqrW2dVw22iHEnvObfhPp4QORtJX8UWDA81pHBOCkFLSqkioPeu2ZDC
dx0mcgcLGe0/xTGJuMZdTc4n8G1WfyB/Esf8sInmOXHYhzG3Wqe4+Zl6soW/5TLx8WLqRB5HlFrn
udUpvzTPAX8P5bvlXa4aOWlkhl4tjgtGRjTcGvTILC0Cnd/KN3A7LfM/n1L7HCmrwKxrXGOda88R
r+rNUE9AY3C338XwdP0fLw10WPgqeYdnM0+oTrR6jrQNY+Hd9e35Qg89sgZUG2HrcdOEf1ytzfIu
cSgbct/Axm+O4sSfmXT3trG78R5oh6nzXiX0xV9pwRSN04HYBrwVrz4mYSXdG1iGW0yTCdgVMFXz
nhu40EY8W6cUEbiXgu05mJbPof9NeraDv3fxRYVdvTjmfsFxlW4DP0ICnGdQFX5dGATeZL74h2c0
crJbCdsXIf7cyM66JujnfHrWSgjitYA7+Ea36dT06vV1sxOaWP7aKOdyV4O8b9qy14BUD4amlH73
X9L+k8IufarCcz7bGS9nAM39vgGDZayIjRj+QjIs8igxFrI4JSXgmxcu2QM5SZQhjWh4A68Gbfpy
gVccvujp7qbrBmVpg34ag+1/dZHxvyMGYAboNLVjLguOV2GovqlYxDb6ilQHsogUsMROnjjwUmJ1
o1+z2nrJGvPFzfosUaPrhyxUNVJ8FfwJbohiwGV2lKr01RzMDZZSl2+2jtP2JUVEn3/m3iajaRZi
hCF06xLde9VwtqFZC7hzfdHqi/c/8Le8+AWC80XKD8b3RiO9LUFMnVl/ef5ukuMz7fqNzAi7KxKX
O5uUouDElMJBzOmI3GejVH9UM3TtqhyvUz/pt1VgDJOLB1dDP9i0cFb04ccz5G+LiM4Axj74TwHo
3mtCa7PPsbqHgR41arxD+gO/q4soNpkxA5/deeMCxRs09Mf4bPhFavezmVdirh4EyNBF2uW5UuOS
UMZVw73tQ8rKQ5HVK3XbTUB7guvgslq5HhMUiWTbnTYAu0No4kN7rFOCJutoKcNI+R4QnKUzzlDf
YvqNuisKTuD8PTGepowgXWjz/mBiPPxPEDu+uFNIvN35SY3UWiWfv6Oqc3+mdjzrI/fc2rwvBto4
rY1zwNHjDLBOViDxZCZsHKkz6q1vN57ovi5aFdawJWb6sn32LTwAXHVbW8kjaM8GJNi7Es86EsK+
mIbxe10dPYf/0PBfJ4xMqUKGD0g5XQfHEk8dQSviYuyUjJUu1IlgP6vvc16SltacbqZQ9K5+rcT0
AB6Mo8NqG6anBJsYtAO1fY0+UtJM96FHCrTtP7+QUfM74hKK+Kon9cTbeQ56m4mWt/RT5mUCP7Sc
ksHNF2VtQqEufCTR9Yl7bZvngXGzAH715gONfIaZmnk2c3zfN0iuBuezpabBtUAtJ/Y0B5Ggkpnn
SqVh4N3wd50E8kZIJPffD1QFAw+CK0QoyPJrRw0aV4kRw8W91VihjWmWLsrYs9fbQtY9dFEgNMn3
78rz4GJ80x98WG0giK3aJ+rMb19eNUw3i8No7n5gZeQmmCElO/tbJl7IhbGJsuUkIweJbh+G6sL7
rx3LwZSJQ42oabV2we2PHvGSfbm8ZLCxIyqbmIKhkYn3OcNTQf2a+ZQty99GPDN0yGwmn7CZyE6g
XwDV2leUmJ5whlpdXkB7xbYWjnlBKPNenot9mBoxfm/oTpeO34uiF7qOGJWxhEBLFatl5ZZK3BHI
Fzw1Nl/5zWh9kKL+4D5topaJPOKmhCXtQEa2WQFsT6NQkIztAOh1syvvmzPGM3OBEwsFTl6P22rM
Z65Lu93bR98KirdF09QfznD0gyYCGEJkCgibtqeR2fLwQ1ttAeuhE4rcarVirtMZ0On/QPNMDfCw
PluYjyeEHI565ZMeB0vWrQZ6romY8/B69QSTdAEoGbj5VP0X3RniECPQnKmFUstrAWOPDc2aO6rr
ggoe9pX/jsbNW57wSRwQW1+x2/Xje9kGLCtInQmLqFOpRLbf9rNwbEhqlqmRUwl+5VQKg+NvwGky
e6gS71XfZ9qnsmYlXKrW7KhV4J1LFKYi7uL8XZ6rdarY2h5JA1WcglbUu+NTmeLXpp1GQkaHe/MO
qByeJw97PSLFZdMZTCbRFZLtPK+W0u43tFB8lnQ9VmIEpZkaY03tI4dO6sYNpIf57jCuVoAoQoTn
MrpAvgWBvmSha9nRfm+BngzKhVKwa1JYzjZA+zw3emeT6ql7+0blcXXpVHY7qLpuAuWyWXDSFZTE
LR7OLQn4vPxwNYZ6qFse+TdgpCknVsDt5GDUqFx8bR8trlN1WYI3n32kozgaxBbP/GtcP0ifDyON
k0Tp+OxKagU4mEus6HlAGI/9/HKT+i9zn9GFhEgqMB9fBHzY8sCsHKDv/ay0NPM8yU/fASSk97CP
p9nOr99txGa8mVYbHvmXGCK2RIMAxUZlojZAaX5JFJkwuDbrfERLBzbAky41Iw2H63oAMHRe6W9u
wHiizFoVghzroBNOyRC8TUAunATjeHEI+hKjVcnPc2P51+t7tpha6rfTlMYBufui4GW5dmeWbnRR
26w0s+yAT9u0m8Ibd6dZKoY4jpSRP63ojAsg7AmeCfVY82Rw66c+cdtdCdY4iJEXPKkG0pP8lFFy
TpIq6FHWTB5tQ2YG7ZmtLM8GUy3kkgX4+2/gyqEy30oxmFnjr76IIaDFr+PEgRsU1wIWO0yqddiQ
r5aGx1mTVqi5udfPRcb2qx7vFD2fFCc9z0wpaCuPJHZmOzfbXDXZkTEuPy58RypUlcpZ3R3B34vN
7Hn+tgPcSjJ9x7u3/22unOaWCpV9rTT0cGVa6hTliUN+pLqFuJCGKaHdQkUeWJ5EsmSlTf4vos5C
883cPluREr3D1LwTM6c1QL3gSiIeQ2mydHLNL+Tfs606VxtZd4Arn11lROmGr6DIky2DbLmZqLeP
aH2m+VSA7otPBpxFj4OJgnHDA7JmcfAAe1VhyaSG+c7sCewQjVg8dfTRI7qu9L4emlSk5iftLBgF
jwKY8XHWA6kYQHaMszsqBN8vwdBwIrXYdr0HyjQPpeTGiSxQLt2KGaSljinHjIz8Jo+Q5XL/pXXI
gXAXzH3M4QVyvom2RVmCzIIbPLODvW9Iqcv2U109lofA/c504IQ4xJiKTyrCXELC5uxOihXC64Vs
BXyVB0OFjjnjfg3VWT/P1Yd22GU/eaOIfNdL/tONGXIS9lJnP5cXHunI+sVuy9aLZ6+MmSNcf1J6
ZrVUU9mMvj7oMjKG6UCWxVAItOsA+igRYdC/6OASsiWakIr+LDcN8Ag1CJr5g3bdNPLP10LyHN2s
TKBbrLM0F22vg6am2Rv4nzDwKI+IpT13DTmH6mG8CU78OHrzDt+9161M+612Mriq61rL0DYltS4F
kG2GL+vh6ZKewCvsGgUw9JWf5ZA6wlNWgJZ0apDXIW0BdrLcV9bLBuBAMng0Qptctou9mw+I2NtS
R6EdfG4hg0BYHdwE3VUbk3Rp5WVIEcq5qFWRKpqWS+gYyrVABoVmskiP0Ciz5FU0u8VJR+lj9V6C
F9ptmIhWgzIoSt4t5GljUVxf0BxtOyh9mEeqHER8HQoRzIz8b9MdAOSesJ25q2MBSqWPTkqMYIdA
xrO7GrfJFxumObFI5z+nKU8eM2oy8p1911kLxfONqGt/bmWXFIZx1kyrQgpfyqhTV30sq1sgrYKf
XmMx5IJ3vf5W97k075vrWnHHQbnozEBELJiOw1LdB+GO9lD1uG9f5LXGBLnJAxYaZvtSXkkU6cgp
8i+Q0rVhlGk0SjTM+fE7+9/5A9efUcPjHVnW2MeZqo4pHTvak+VNLCIMiNthhDjkqDQg7JEVL3Og
BLpuvZoubZzYTMpRuoUnwv8PgrTav7WNXpWuwbm632D7cZosFlm2WXA1JVglS6difBS05m6Vzmkb
1I3Lqx1ERMHZiK3KQcvg023WhRGA5xKRaGL1opZnBldTRD2p960JqAePj2+DdxUmBzKNw/XL4Vby
BZS6ETi4rbH2YpO566L6QYh439qVfZ7v5t8pOYkvQKcxf24AVmsudhjE7EXxYZbWZrqOrPbh8eBb
0qCUzMyiMAhgd9Ejm5RxOuy+RmfFuGaJY8zL9DGllV7eiF54e1pqa4I3I6wPTpI1k+iCqyPpaJ8b
i1Uuk7YcM/tUw/BudPuWM/Nx/HbJlVrJYyGh6v8BmZb3tqbHblm9GBtbONa32Mw4y/Ecl2t/+3sS
JoR85dkSqtlgbGCYAEQE5mGy2ipJ+fdMbpQmwQjZC+GQdRFEInMCSGKWKzmdDA7WX+fsLLD3ljT+
TkgbK23rdTXy/o1FC34nAjabwOvVaxsHKN8GFRcBJ3/z9wrZgIpRro2mSRdtGFiDb4pDoUFMYS3x
xiAOX9v5IjRCaCWUKAhYdRC9ykpDq+7THfR8R0CGKGJKOrpCBv5nn57QNyx6egmcEQEOc1drkgKR
/I1FDw0XWZo7+dzdS1u5RnSo7nWDIPoNqm6C8lZCRkQE3SJrInamqpRBynWVcs6n9gmN7NHs8mOc
pZMeBFnZ/GvvrlVfLUT93Lq2YOf9moRGuHLi8wg3+i/bDaXbB5WzVCpd/yGer4/g/pNcnhveSi6w
gcP8wWYnHHnvEnJ/o0YqAeDSj+nlRkN8luLM2P/ixUQQDDx1L6BB3MtSlZmAWSS2CntwyGPsGKvG
dF1oJqH2lUsKivBsWuw47APOTksPmm6AQZj8x5p0x9K+XhohL35fYhJkZvRLB3r9GM909C/HJUWs
JmlBTa0EyL9zqiZvgyrHts+3sooNYbzDSSMIniekCZ+tWNvIKFTFs7+D3dRSKcFsFAGscEtQdsCD
wHam896+0m3zgJKzvvabVLv1UiZLCvcD2RiLHBykibfjk8A6//64StBzBIT84NvGnSy+2oLpDaxw
2FbtY+ZBMHgFWdeedWAyfJx06e0oXmVjHqo6YFgyI3ZYE62U19Xcogj/O7i2+N0JeSsaoDoaQZ5b
SYDwdV0cEpgbOGAll0trVdFr1y/zRHT/J6fYm8s3cp8zx9+XRQo9xYZPTkwZ+vr2DFQYO8RL783w
2uZXVZL/dg1OQEajDz538NxP08WS2C2w8AOtiskucnPkLRB2GtyASj8JJtgbJ2VJVxu44+T7xEJa
cPFI+vedMlvGpEuH7WyGsJJw67LzSbSwnRMs0NtgScxA2UDj7+Mgomv4e52+F740NNPpoWwIeyTh
FXNXBCbfjw+2O0jZel2UwtWu+WMlx1Xgz0HnNpjOQuFDvS7+eHmKBOItKdygFIH0VmR3jJdjo//b
BxMesitgflJXPG/qYzlnRTtX+aTgPr60ZITybkFFrWR3VX1CYPqS9MTrC4/HaclrzekGocqwXhjS
hyK11Ss7U6f2OVi3hWKPkNWG3LGwXv/uz7nnY3JkQL0Mw9+lDX8/nEn4w39bhHnVm3s3EEbTpN9s
kxej9eTTKHr52mk29L9dFP53pg25wdYy8JJHT6e5GeUeoMrAiePWtLD9Jwp4AgWwX+cIyO3y9TNU
nEjFcpauQtw9kKpK67SAiwE2YlID1Hldg48FNExkLmGpA0YkWDZdhJN07aeySdMlCp2M/CQmXU7Q
R0aoC+x0KamAOCAhTs9tCwyFZMSKA7t+HT+PnDPUXWWlBYffgbWoGrScseX2r+iW6X0FrwbKK+Le
Q4BUc7Gy2alvdECpvEgCcF/rYpFM6p96Ssf+Xol7G4bkmXxqgeJc/8IJh6o+sUB2XCMVkRcjOsO1
9yJCdgXErxfx36uYO4tSBu5S+MK9WlAcXsDX2QL0pVdB9NgCo5m7xmwriKRHoogdBiioTOk0d3x4
l5aKk4rkFjDPCZrZX1UTrsIqPSooL+ccvShXbIMY6TMoAFOIjom0AOANHOrDbNxo8Lmzof1FP7H2
z6lnFrRrNu4zkVnvIpaaKqpXmZ5YqNIAxffg3nqyAURvjp5JD+cb/wf9f1V1vqeZzECRuYxXD8WA
aarCUilohMbnPEsX4xGlWkD6FgwxBUYeCi0sdjd4WDxqj7xjDR5jWC8Lus2VQMDuPa2KvWYqhenl
dktczcLvpb8KdAL7uYeBwxbleKe9295HRvNs5U6Q/vxqNx99pfwo1AzhUvjZyHT4pcX0BukVHARQ
+FaCn88kVbS9ILAq6p1q6fQq4VFV7lr1tWRVoFY+IfHdNe9AczQN1bdbPlFkcad0uCwIQ1ao3dtm
fsEQvOur7it2NLffPyP3JxrYqE/gNNwaR5qq0Jl4OjW7UByGJ73kqrck+KscF7nbW/LmMsOp617x
AYgXAON7tajfZb8QcFHVRIIBf9uEJ3nKSq4tH7+w3vDFyhjPx61TSFuN6r+FkwuHbB59lMEcT8Zy
ldBubHHYZ2JSfYdopF58x3j8wEsOAmmSy0+Vqr8v9GS9TYL+ounw/FXeyHtDlWshlh5AMZTlDE7A
A/Je2sE0Ayn3lYp4Biqyc7ktcPQXpoRolaG1GhE0oN8u29byMqSdfqCfMe5DWpEmNQ73cSZiFFEC
snQ1EU/vWnIdE0hPVMFHnAaffiDx7ieyugFBRk6pxw3XGnxA+IQcmXj1oBu44LZgEll1O7ORYRcl
3r7ZWcy08u7YjhFSvgXwIEYNTXCCPYYMv6l365o/TgTwCQqoz0pA9CELfLC9be+V6BBHC8hNg0OC
J4twIXGeX59SbR32DO1otYICgel6UzFbPDcvMLR66Jx7mPFEF8Ntvs7dU5Hociw/7KoSuEU/lFT4
0yzVsMes4+l647mm6H5UKMqwJI2GpNwbAeW8DhWKg6Ag0d3Fd1/yzpXX7xqTqW93FF4sXqtgeVla
ECTRMevFB+F++dlgS/hQM6wU/nTqoWRtfh6DDAOJMr/idmSOfJV4m6TBmNXzNRmr1wIMYoLgLh2a
chFsoZEJfpkFqKog/cpafo1OR91zlF7Ociz6Vo9b4zYCu9XlCPxM/xxkCP4iJ9kd7J6mqYJpTkRF
li2NBdXGNYHiwaa4d3iO0PdkJgxUjt13i7tD3rNuVS4bkajI+p8E35UAy6r11Ew5lJjliAfLXn0W
16zdsCZph652UpwmtX5G895/ihBxuJYa7kYCxmSV4q3dd185YOY0hhToUVeN/m12WSbDNd18JyVl
gu853f61mHEHxIXffk3TeGUebGbSiQxIfCNfPbBkz7cLhu0jMju10pI2a8UUZ1oc9a7GyB0qIZvj
g7J0e30VYtJz5IkksQgrXajY1k1LKCvI+kPjk69xm7l2age5RN8pA3W+dEr2HDqDh4NK+Dl1bTlj
Rz6nF/QAhayRcoxqEmk7StUIhPNpiuM76+EvYotHhSDFwUTVgFkJT0BMj9MHIOuXwC2EuZNG8bdN
1mdcLz2oeTm2OxPTy8uDnVDOSADZBW5JJ5WdVbKSiZ+ZAnO5y4drkYee7Gqy5Q0h/3E5h1k6Exll
geJGFsia2P/ogZb1uF2wa6sgoVeOjpBXuZePw43ocwj1EODQjLNRPK0m0U27ktWvC9+1aI8PKIDc
rr+tt8NhjqiwOj09H1AiY22/hMVW4UAzc3AC+j7AmCGQVCcpdP6Q3nKDM26fQe/NJ22g+oqOs8nT
H81BoWB+a1vNNpQ4Xm4CX3InfFY0HxzcLLOFeM5BEqVVRy7CkksjFH/BbWrO9KJ8/2q2m3b2ijYr
7BD4HMswqTY4Bn4t66eglM5P6nK8fSX0Bi+xeCRJgGYRyOmd4KHA/9p0+9kSN2Oygv6yLL0nWb57
dSzmG7arbpkw/CQjRb9gVwktOzewzyZl1HcTHX0MaGy6PYojZpTgJZ6Jeh3XQ4AqfEnCvuvutkPp
bpd+xtD/+WJYvIxZapqOPlV4A+ZlMu2qCkpKu23aC+5KaX0cKNnuuYcUNrmAkm9pnZTBAlxu+KAv
4P2tu77awISJEfDXB+c6ybTSgA6XNF+NWHVVjuG1q2qqxWldhDU+rYqCZPxtfvW0V5lYOeVxbMZJ
M1hFgWiuHPf20B5uc/Tm7s3OryT2E//iTdLE/KbXz0x86tvL16aVogFSCJ9XX4Gk8Lhsxi0hE8eO
K1o2AozczBy0/yEFHsI4mFHCLk2cp9hplNVqabzc6W7oUMNJZuh8U9nNg8ZXPRGzbs9TCgpLwLLl
RbDttHN4QuGsktzIkUVdJqs2udFHe9tQxEcqVTiBygGCuVW8575KplFwf+CJBDgUDzfnSeaJmwJd
kmkjBmP5Qhm2GnnhuX/wbnFLsbxdobc7jP1JQcDM8I6Pzvgkg+vbg3gTEW3ajXmdSynQG13wjzIF
GuULs0DsdTSzgyefyJPeEdinDvU0A7OuYrmlU6/cWIiEoZWjT3pSU71c4u5MjWUU6FaRWmXEZqXW
rJUyhfRuyelzN6Lg/9IqecgL22drfjxsEMHiRb3Ck3WEv2uvXzGAS/JJjh1idfU3TG36qnoQ/hyz
KIx8P7PxBBEN5v+RwYuGaIb9VEgQA6FF5UpH9M15Pso9JxvsVA17q3jgKtqS8LZJbNRIFXTQNbyV
SDcq7E93LuKUcUY4LCAHUU8GgG89+Cq3yPRxgVqAnDZQLeF75rDcfzAajTq5BDrUy078Xs/otXBb
ldZ/QEj6bHT/PSqoJLCNTwEVt9T5mXnMqr8g6JDD4BaCsGTjj4SZ9SkG3D419mxJsiQT9XLLbJuK
YshXf4XPEidoAQ5PuiaeUR8rTL/NPNpVEE03c7O/PA3yyoUXEJfkPNbbJXpVEIypHYZPg/dlPJ9t
ax2DhejahTjY3WpiyBe3yv6F5pceili0onJQhbOCgYA4PZtjNv9aZ03v7MkKvCHQv0F1y4b/b9k3
2QK5BkqkZhWNvZ/X5A6lcPPzEe/owmNgNZ/CXEtVnieKMfUxlbP6z5pxu4pMmwbFVBJlKyluA7G4
Tl6RiZ3mClE7EWeiCnTB39/DVwwQJA85keWkuTVB/ApdOPf40cqFjD6V+cx+eq2fYpmq/bmWyjmA
ukTqPQHdDXmAsT9+RdlbWFuj9daPY0/mCOwWbpTEYaGhMEaCOWIBYnRHzVfM4IpGcUllmzV10Mss
YeKbRDPreNcGayulM1h19nNDN8ZhoUMQJt6zLFrHugNcwqYiBjSoco/M/IJ003nmtA6u5x9FfNZr
H3oqj0x82h7vrpEu4/G/b8f/JH9aD3ocI0UXWHUvKq1Wr0HSpSQunhSFS3Kv2uDLBVhoudnwBjvO
shJbwdl4mS92tF7DHYjVVdnAmcskgK53k4tX+bO2iyXj8QpGNB1Z9KZx2KWfcbQCchX6t2t8MbmP
ZE2/dcDQsccEEPx/kq5W0++ruoDSBpWoksMLs2Xf5a7HMZ/Fh7315Yh1wxX5UH+qhPPbEzjUPPNk
1Jx1HW6fX8I3MzLGD4d15hJn+7BJy2wmgO+XsV28XbYIJn2GF0ZSfhpckLY6V9Y0jkKE8R95+1AS
DcQiKXdxyAw5hSzjxzDyNUbkYeM/Gqpx24rYt9/F+cW1WuMrJ9DFJFByEFf+OeA7bcyTdC01nzAj
JQUuyzNgJb3DBh1WlBk/Rz+skDobA0HCFD7P9ieOWNsPk8GgE9kbYLmB7xN3/IUmWV9eDdWObFGb
l9OvOOiBIi8VSLWG+MAAbDUYjSc9wnhwFqM/sJUky3xnc/dwGkdJXTBJ5M+sM0MB8sBAOjONgT14
gBf7cmFxjPiS0kOIwtb+2F2oaPhnIqqZXTIxTIn8SzfOrsS9+qSWdgYtscId+MlBpBnGPtVT04JY
HJtMXKPW50+4w2QVlusOFMYTFR3BcV4fD0DXYyMWg6Vta6X+jZLy7B9Eax7dwkNAF3CwY/ld88tM
Wg26L5G0tdxBByinw6dGmvcu2mk90sETVjk5/+UIvK4eJDQLbSi/fYJoeuETqjIpsMW/iZmEh468
QIyyfNXn7B+P4R2jZ0ESBB636M4opegnG8piKJ0PWhgwT8ulzeafKuSB0i1/jLpWnIvT5hIjY81I
t88+6J5MaGmVzmF9e0B+8f/RdWukmvyqEOwWbP/Yc+GRUUxA11XC57iYdnMIV9qLqYzI58j8kt4N
oAg75uEkP4vWetncqmshW5mUTmEz6zrwlY3t/iy5hWKL7Eru6DKEXBt8+6PYDAplkBynzOul1lwr
0yyvlqF03speRiSNuy4KhhQyifv6aNXIpqbYkT2lvjKLVZBIU1H7Jpfiuh20mUvhtvxcNSpE4KsL
SrjIyJPUx/Xrmxf91PFRhZBYCQqq3SIPy2SQkKSYwJVYiQ24jaN1Vl48PxJCYESe8Yv773hoGkl9
SqJhFrFzDH8KAmh9SbGRFPZ6hwpsB5R8xb3z7UDrczmCNWPxu/8//psIsVQz14TbzwyReJ6M+hpe
Qw5gad+gDWaWHe7ZAvha1dbur4lhYmnGdJpg8ngNVwiPlOJmGY0lYEfUF5ANZlw2ebyXUvGgCEf4
4TmXegs1oBq+Lsrj3Q0xBSL3tiUMQPCQaPHGfe+D+fZKsHfLwEY5eQhvZA0c6Y7+K1YovQmgomQB
HhwXiHulgwAKTmA79BNz5Aq94UQo4yIbEXB+xd0QRhB3T3zqEWJMOJuv3i8TjysErpQWqyrP6j51
uM5TnFqyniDSVetTDwU1HNCbYjKcGeWxeUFmWbMhBugA5ywor7/g2LNlxV3yn+ardb2cKu1raF1N
w7YSdbRU0f1vBoe5zrvJaBCGLoxmlqzl8RdNMcKmUr9bt6mqLiOIoTbjNYrbIsN6J2qeJCX3DlmM
UPugswuTmDxaHjDela3gB8sVYMmPGtz3wuwgjcM8Kcxljo0QokThPSZn9WVEhncGiJl+6HPjT2qO
tP3pcXgE00mkznjDOuY+6nLOn/h0nsSMKfwoWrS7IX7ofb1IjkjQNLnIdhdFuXIqLhMs+bVor0LD
p+DMuKnzeCn4YAOw7Sk/T1yL1nVtTemC9OCKkaL+BO7l1mZknHBJzHeh1BkM69Rel6EfeFJKO63/
JgLXgPnKNuUEOA1hG3lXRrPkZTy28UAOtkE8kaEGJ8z+E/gL872ucch2LYlq4McbXkU3w5r2Pku0
9ID1e3Btk0SRy5RYtPwbuziBkS6EGkPBr8Adz2++uCwl76WgUG9zHRxEoMFlQpfONOBECaTGzS+m
2hwee3VR3gS3WSZwDw6UdnaLSXK9geoUirnIEaprwe6y3QYywAusMOfN7dl0fTGOjIV/AW0s7GJ+
c8GoPOrK3NpBKfkTQp6doGVkaAXpy2jM4ZBmQEG/bSWwo0sNN0xRH1MOeL/JCkqjwmQBbKX+hO5t
QmHTn4Fa6DL3tx7Ufr3yd56mRL9Fhg1RNmY2OVgK9B31dwayIuzCvwQ5XbOgLWkuaNeSbW6LX0pp
kJ+C9ztqNtX/Lt/bm2Hg0qBGU9tWkx4GgMN+w6QEYOdbiQqMpieusigB7VBEGccnjqcjSlDBU5cS
KtQ5ug4qLl0eaJD3iwSflZvaLQOvwf3bxRxsNA3B/adJZQHTiqJgGTrX7Y/Io53bZWDNM2mBBT7A
Vx8w+VTi2Fe0ApcLswgL+8WWKtxw9QbcwYdEP4UwJ+52qh3QSfn0Ed9H6jsqCr+p9Hohc/WQ1VDk
/hZ04J21BVt1w++lKmWYNS6SHMAn/t7rx3gi+Zl+wM5LO7qO5LqBxDCQg1I7hXghYc/sttwjPn7t
3Ypn/3BtygmQuCjHx6nV7EZ75Tyv6X3eeVi5qQ5We6k9hv8YWzf6uqJBWnrxp9dkhSvgpV7I60DR
mgAxsJNETIu0HwdFwuNmWepsMlHEM8xZAldXSYxNevQ4EXsdD2EuLGeTdCpW4pqmpXEUh3hERRWY
OEqxH9o01A/LeHMAKFli+ARw+7DB+oo0N8wlKX5L1cLQyVC7DWO3GbSpS5aa++lSH0OSTdHvO1dS
3sv7IunSgdB5diu9+UfVoqJUgLaazqCDvzuWQQPhcK9eYaoVVheoVjtKTbw/Q0wDllk43Q976xKP
zFoiWe01ft4//1faW9DeF+s6EdLCei0l9xq1Z4vfA1K8V2Fksp1WE5xwlv+ArQv69F47y9W25MFz
hQmWVf6Tl12nvrZ4BQEQfvxuPi0RpSddj7IrHFF01sRUxMvwvRDF97pPU90WU5p6l4gDPrEt40iK
lf7pbwqe1qZEDLDOW0jomeCbRNsWB88/ORpi498MJjUYm66y5kfjALrnvHI9DVFZasZDdlv6Diyc
vjVZkN9VQ4hvtF91sq9dpLTY6gqeq5JC0XDfull7izH8ho5B/5huI+HHgwkXoRCapH/rtnoXTQkf
ZfvjKq2qzJKs3fB7SGL1Svv9bGWZrllOzliVrDhCTCoxpncB6UpnqFM3c6Zd4LZ6/MRrdUZfVvBD
W1KoAevXC0tUuwQ6FHsrwe/sZEHfY3l5b7VzmO6TvT7TxG6FEquZhVwbYydiaBpzCzmR9ppbY941
hHVkgpI/puLWAdaeRM9PPUMNDaXDPo8sG6OQsi/EFa4yYiBy//CnJVVBv2n3JEjFwyxaMiDPpXCJ
iokFiRQPC+oPVbPEwm09ti3i8rHvv5GJkwTJxdfl2z22IuTMAwKmWgOU2Me+RLCFP2QdniQ/F6S3
L4zOMj/GRnTOu4AkzNphDwqHAxvS1o62bw1CYOAjbMt2e2kTUwYhPyyhd+pXgi3ZQer2so6IlWsc
XdaJ4N4pZu+X3moMrmZU9phsjOh5WilvH7gBLREhGHCkDczonzHK33NclOn936irNPjlC1CdfDd6
d61tsO+GhnjbobzL1sqIA58cCRdvO+SzoAJgQ82Ao8n1gd51Z/QjxnKArb2ZYLSxjRjg0u9l3Twi
rvrboCwPNnv3oFXc4nKthefLoG2M6b+NWL4oY0YJ+oAwoJCPfrJ125Spu1gsthHaOLaIqbofBQPz
Q0m88pvA3oZ+8VIYPHModY3ZXeH5K65ApFor6oP6FD1NsPZO/JmSynRUsZQ26VcpMa5mHIsTDF4Z
BuTK5Rrv9UEJCKm/O7a7ZHLKTyCkeQ9p2N63drgSHzBe60fvtlFYdwxSCC2+RGb3EvLCRzJrUm0W
2EYyyShvWKZRBaUUoP671WAmMyEJn9/AqSbvmAnux/JgMH/DyVd4oTDk6I3k2JdyYFWO1Jicxc+C
3U3W/aaooUMOSHQuzhkM+NqbynsiUIaEu3mh5GtLBNUG1ULJAxH4RtRM6MXCMIsqY5lJ8SW3WV1B
6hshVf/xuT1D8LL8yw45XI0HOUsvH2VgigXIXtucSyfblxU2aUplfW17ytzi50i/pqP+w+/c8BDF
BLqlvGpzzZvx1oXizMrRANw1yidmPMYQdNEqL7ezUaJhDcLjtsTXHJMup68hQiGqxQQjiNZW5nMH
UA/N26C/nPczHdrp1fpd5WVixKEIfViPOKT3GpmknzqSZIBh+LWulES5eSIzB96d8mfqgAcAZ8R4
12f2NdEH6ZX5qlbnbvmVwY8+//Mm/nc9xRjkapP9IJ2unhK/2+1JooUtQB6jYX2tD80N/2Phaaq0
x1fM3JxxIUE/1jH5SpxqLf0JHF6z0v/dIgZth20+w7IHajrfPCoIzq9O+rlKi7N4W5RpT9Ob3kzY
qOtljcaBBbMIh3CVn6yitsSZJV+/pgaDta0xzRdLIqKNZPO/4Qe4hx9C0aMMIyaX5RVRxliQhT2o
jIb7LnRyM8ukTeHixMyWW8Ip8pIypX3vRmqQ+ZkX6ry4mpvQzXzrx/9jE79zV29B3rg7hDfhm1XD
8mCaWbeKpNbp2JmQZ+y/yJKwJcC8wQTo4p0vTDCsRR39JJYKc4EZdaH6but+RHfXVizIY26BRSN7
1+xipBG7/zcf/5uhR6cPagPLVhoXLkXHJxsiqFKHgQ1ms2oca2YsOSn4LWJSQPIu60OA3jXIB0ei
WUx6M+qeWIAVHYGShJ9YjPT8YKRfEGCSDUQHJ39M2wgAJGjQlhlWR3fo/9bZ7KY3pz0RFHw4dIu7
dkBtOb+gsD4mjRu4jccjE190RWnayhFrfD2wcz2t1m2VpfKaan5Q82fsvQ/bSURhgWrfCu5WU6SB
t4Bw9NWO/UG01whZiQckxaV9tJ9nGmc4wUwnnRsQbqBgIG+Y853Nlq2JZaMbb1nz3Sx3shbGRPg0
BLE8k+fe2U9kfmFG9INu3HZuAGzwRuDEJojKmNUd+Pb5kgftzsGuUDSrxJ99QvCEY49oDO0mgCxj
IpSvks3IICzZ2zstkUXBUlsf1DMikgAqnqAYDmIggXfxVtzmGCfn00lw4Qf8AZDq0Xir7imm2J0T
EBLMlablxy4X+rNcVmN7e6n/u/ufS6efc+Ipv0qGLPLgfIYtZ6jTjHEqCIUTlLDhJ5meMylAkIAG
VqQulnSn9ucG72LKPOlVYEj3V0CLvmWWeoMdcqfc3I/6WZy5L1SW3Utt/PIdvIEx7AyiQ6QX9kXm
eyRSBM6woGKnDs12T4QO+2XUcMoTDyNTA1dY5oMtNzWf6HKZKx5llgijdpAltNnB1NScaAXcOMD9
ufsKY1oSi6nrw+15PDBtUnZ321/Mo4TWK4cyy9bJUHIgewEikC3s4O7Cut1FfCumirNnSnAsORz8
2SSdPqDQUPIWwTZJ3JjB/3yhHJe8tjc9RxWaMlbFRHdtIRMuD/ByAeYkxjAc1vpmxfyx1003t8mR
WDxQpKR7ydtT3L74QCMox/L6RfTRU1neKfBRO0PjqUBWGFPGZRtfH4oXj6ZhZQpLua0cbNPpO60h
qrdRDbIPSz8KvJ0nKf0xyV66eufqspEwl/ipW1a3UtDZFn8XwmjKjGT/HvkYIncZa16dtEDPoQpH
UlvQYJc8A7Mm0G8wrsXJWyk5D2nzNTdxMPGaDGLKs+hqaQ5Fe5r+WxxgBXQPMWpq8v+ejhsnNrNo
SBEdrHHSHY8tgIH7Cg5DgjMaNv2ocYW7J6Ibu44ULoDNpE7DPaORE82TnsAj867pEGZmuyLE96zj
Dtw26A3B90zPnIoXF+fKCFAzRNhi0GeaFz/wz+cbzaxGHvdtmgxlcyniP8imPbVTXvq7l5KrNlOu
D1oJVprE1EZHpFYYLRrePB6mdUOqw+xCZpfWbkMG5S3khgKPHY7Icaio6uhpZ01HPTvTleTyB5+A
4bvEyMaq044Npv6yUIHpMgVsMxn6o7b95cVJwJiJ4GKnUM6l+BObF31fLrNFaP1azgql2oM3GgvM
1qmaJyJ9ukMOhR8wnHzZvxBAe7/PeM3VFa+rt3XnYHfBU2tlVV/+4rCvJ7Ae9PNYiE4dVoWnJAsK
c5xKcxWf52afaj5V4MEE88B84X7laJF22X6CnvJncR//L1C7READ71h0LBav59CcBw31HCJfRbYU
4MCUxXzmwuU/F+Ccov1J7ENc0pCtvWZD3MAKuvmhoLdLUamkQKSdnE03ayd+Iic6l8XpWMBiZMyW
y97rLfGbHqF5d0MZ5mu0bNfRYV25oQMIkEn3XL+O0R+Kki92Tr2KjfU7d+mpuduXsB9523VLYU1N
BdSGAVegzMCHRFT2vhj+4vuje81fV8y+Oo6AHmGZVIbpFgkEu5OD6gY/CM0MYYeMQLAB9Lms62f1
dmhxsLAs7lRLojFA/qu4qfg+imKyLkv4vnTq2tBrMCqfek8QfOwscch7xUf2lYtSkUPyzQm7jxEA
KSBCHAGS9BTmq7gKZsVx1UsCjWZt5eRPLym6tEOkuEnbYbChAADPAccyKJZJ+ADupCeQXHEsFRbN
ZIEVnOwZm2PlN7CoapsYfsaqDwge3GDkfbGsh5RAjUcFB4ou1L6E5cCnk/JYdw5MZj3s1dH6OfNH
1GEZjRahqEiiMAJA7viWDz165cACMFc7xJSvIk+bRiMZQm3fDeC20CekXZQdlwF1u9YrBldu91jg
foensy9UvH55AG6tyBKon+idT4Ar2/KM3Xn3yoyQXtsE8LLZXWXeu90yPO2/jP5RBvj9dOPQuDzi
fOJACqVaOYOaQ+aKdDynVkFkzUN6tUAKzxmElr/05GHPfxH5HP9XKShZ1cajVdgFEeBtvH0/9rWA
i3Hoh7NoySONIEMFQi8iycHjGHIDT4XCw/bDMgNqdsphpqKVEUWGE6Bf7qaKU4Ym3BF36KLBTNHl
EQCF61/QpngzsCsiR18ZP1kzycMcdh3oRBEh5Cht8wj/3CigQC5yF6EohcYmFtZAwnEJpASRd/x8
z38BL9VpzZ5XX2oIpnnKu0NlEOZQ0Vle6BQHjl38VrqxFurd33TCXUSOSiVRwsVLd+zdJMdML6Xz
FZ39+DQrYNjEcn1Hh4R4GYu3PIc35dVDP1ukB7+x8Rb6kTQxxfSLURi8PQHVZOGqVOhf0fUcax3z
JQ2qUqHgu5wpsktJRi4tvvaEz/UKUUqHkkA0c4MF8ux4cwUwg9ooL6/FXXKlE+TkdbXxudzA4Iq/
4+2HlPTPNlsMO+XH2VJEjCaL3UDxKsqQytJOLqX8bbHHT6PuyyOpkNkl5H+Hxm/KjR3FH/X5MI6a
OVxBVWyWTP8fHbOaI7U9/kycx5d6jNyAWSEPL3vuL8b5ZXZmIVYLafqBNPdiswIYTPcGr1wBs5fS
PxXfTwhzeCWrbiMx4A9WZDaEq6hdqzlptdHulf8joCWKdzc+oIIAOcNMYGwWmNtSk3JOIG0n9j1Y
+gweTYAYl2ROsgJNqQFTogEc6mqockCSg+xZb5LkowXTs7ti0SDjkAMTK+s25W1+o0rmDXY45Spm
Y6dLzzd19t2hglxv9w1GfNPNfambQrRefvjeeVka9PNitUY4cF9DKW9iPpz6lHNarY19uIVJA/03
aoinDRUe6gXVH15HjqCzIwYlWBDpZ6p3qVJbfau89JK1QKxuo5PW1J/fLU3TYa+0J5NIr0NFXhdk
XMdB0jHQzElH0kgMkVN49D4fxV+KhfseQzVWirGC9HCAXW1KByqzb7VouuVoDRI+bQKf4+3gQ7PS
HhmD0P4yx2ofMmkpN0U7YuyjGFUFv7pMQ0r92GnOPVFuVHGEGTx3RkHpV1jeWZTV99txb4ckvTSM
3uKmOOvTmV8WXZZCL5oSE/0kHHNUVNuqoUyr50t8HtGOn6nSyAMS99E39EaHza3M2imaIihtZFIs
DyvIXQjx9X6DgGyCsRKCF8Kql/YhoQKE/Jk8sTOOAZKWeDs4pXVfZ/Lfo9cAn3OADd30521AwqBT
FxiEptlzEECnsHQnNHgEICfL/bv9ssaFU8xVXUL1YXv4n+uAaJAdotukgn1QRXWqxBAr/NohAlcH
HO8ubpog1wBlfGkHASRvzEqI23E1ZHHieoyqJ7StgwGMvRO10Xqc8v5xcwld5PNfiJ3yg0tJv7WL
1I1H5lDufXPltPj4ZxvCPyfP4LoUmCYrqusHUR+e4LrN/zY/zuR4Sxz9TndJjMA7XbgjLZZ8ET0r
g1L2v7Dwktjk+5bknAt2oc9PX8xGUS9QI/kHNuwS0qBDY6FSRfkzx4jc9acdodBwVqcRq7XEtyNs
kVnNlLketzg+o/Hu78DciotKlLYpQCR8DcWpcZRsbY7TkeYwdVNZaZPqAw8XvpLb+g/2xB/hfJ7g
nmcnY/HCyoHDzzOdfg3YX/EgHXUEgmWzsvi2mSlBcPH+0GRP0630uj4X7fbYDfUdEBMm6lQeSAk8
azhwU+7GBLHf8OFaQml6KXYppnJt39wC4Mgf5Fkjl0FNQ3pwVHP036wvjAtJV/PS9PpjKml8Yet+
VEdcO3j86ip1JKkiu3MVUXOiUQE5/L/co63tGnEXNr8f1tp0O905aE/YSrGMM1g8xucZOkuvgy2E
0s06tl2fJEkfy5FqGJyRP5n8X1NozoUol8qe6Bw5OS8PNfrMIohbFuerXdlxJnPZfmffHDmaPiMn
lr5v8JN5P/sZ27IiiwwiyCYyamoR4PWqBSmGXXiUStIo73zZb7AL/VMslK6Hbj1v3foOoIkwbj73
j7ehweAqLJGqT74uXj0k/zv2/4xOQf5A+6zUjn9IvqHQmge9VWUNl2hDEFJ2aJKJkChFUOimWc16
WCBj4kxLmXPkbBm8OgcLjvqs2hbl85e68UJvNRZ3DOwL2/CBD0hQvwBd1MukC0bo1AeFSk60mWE/
67+pY+joTXzZ60UWTADYcCek3x2C65PDvs0VXUiwAx1lx0xV3JB0R7bOwyL72thHqGE079pVo94A
NBfj3DDgn0A395UKKIvEmlLqBB7E0v1M5hw2IVngcHktn/N+5CsN+5BDyBhR0+zzWXb48OHPg5OP
LDo+AxYHydcBd+vYKG5T29fyIzktMJlSUokLq0mEou/IvBrXmlfkTUZK8fVvDgIm6xkpQ+/6HwjI
PRMY2MkNFX9tgh3Q3Gp+so91fRBI/1PTM7fyJB9ZypfJ3mj59oukaRK7TPWfaajjRD74FECpUZP7
3oNND01CJdsvbUjUd9oqy3DIj2o6hHCVKgsxR89C5DnOsj6xptVqelqS8JUmqD7T0FuG6PfzHc1x
FBgs/Ce28WXZwDYJVIEug0NpRmIG0SoyWJZlpb1qeTv1yJxii0cO1QVlp0BAXTxu7iUtLZAcroIm
C2lWhgLq+6McvvHS/UY3RD6HIGQyRNHhiyv7P+6574B1mtX0xjBOXYKiY88dcqy6CI4V5GmYQbyQ
Zp23f+i+jcwX9UK6xmR4OIPBlOyPci8RKJVi76b7ZndweGtY5DA8XSwGpa1vtQS2IDCsN0UsDsjr
Dz5YdU9fw+X70nCiG1cfqPIcA/6UXPc+M3yyK4zlLiSkjAZysHuwGgpQF5mjsWG/LHyd5EZQT5SN
py2p8W3hqwYmsz8MjXwpGzWM7rINZ6ajYGFKKl2jM8tyDhvE2nRurlBKv3dYz1QcELJx1Lml0kpt
faSWPKUWahn4dWKhLSaDyy9HcNarJgAGWayMF8MI41uwxfdYOi1EWm4qWWOz0NtaYDJPDyxxBUsN
xgXXQ8HFvgHUv5CG5xmaP3eeFVSJ6C6CkMu92B4zFtMOhzMKEGITtQu0lanE3ubTcf6ysxe7Ip5H
GrcGsTzJkHT9jYisPWE7kKUB0jR8tnhUyGN5gaj0fUKEhQt4olVnhQvQSvjBq5ZW1cJJyX5ub0IZ
YE1FmWsMoYsx00JEaR5QM/NHSSuOEuUQUKTWnskH2qlHvcFs8a42+uDmENlu+mbplnQIpoHLyYRk
yHZlJfyC3eNLDKgcqg+Vq7HfrdJqyGQqryWSj/SapAMaHxewLkAM4Phpsno0CEp2WPIKx+it/yuR
oDTDozq77rBPHezuJCRshf1FE1xuKcX9aqy9ETZYusHDcuNei8o7SPTfxPeyF3QsHKWrQhTtStp5
pc9kWHjzK90W8L785efMxINIv7RmVGGB7orsa+lqtdfXpF9UieUehfI/M6lJPMRBVzKx4TN/BCXn
rfKdqk1PsyAMtOetz2p9fpFULddM5W90eV/xwIOmnVqefiN8cIcUBBjn892rPc2Zvj/PaUPpfF+5
dY6VEGc8jZhxJxiw3cr+4NaHOCQfYET9Q1m0IEo3SNIPFPyI6MXXV2Kph05BGbbUVkoTGNQKwsHC
rQkGNUW/o3+eJ7pm6gTuHs5SGM3q44p2hXy0NrBPwJFg2J+FAWB28vDFo+l+Qiy/yZzF2qwxEf6r
5s5N+B3uavpHe1Zgu8cASQdOwiQo4S6MKA8CKroAQEAXikfN8Gii1+ayWSL55hmmJDuMnjzkFjTp
W0TRuxttb8qcE3a663WXD1Ju3UzrVfMKb1+wHTu7s8Ww9CcN09CM+jdw4Gy+tFRzlH6MzouZD6q4
YdOObBqls4ncijOVEd7HLOsY+PSOfLyg08v3dq266zBRdceMqBN2OJL6283zPdMxXjZO6DiUADX2
vj8JJAKhRkBlTuoY1/7lvICEQI0RhD9k0JpvGepFfLQkNDaeIbFgbby6aYJYdf/Ftb1SNK6k7fKR
ZgB6ELIyyQZ9nrFFPkd1uq6UnJd+GXWDBGK92osQt8A1CVZqqRGeMV5CTgLASmM+JSCpfQeK9f02
ERRtb8rHeqj+Nf9LQUZ5h8BCNBHmCsfs7YRBo6scyTzGdrytY4qb3NpCVaOhqJw5oD6lr2qMdd5e
OmSrEABRKUT0RY7zO/GD13+DllST/BkJE235frg0ve3u4c8w5kzhc98UE8qzcoPXkAZFLAP5YV0T
arAYcEtDY06SDxxALqNSakNSBdKaO5SGCB97vVbNXOEyOkBT3B/eREEMoe6FaM9OBC6z4LlQ8Ohy
TN5sxXY1VIMGjpY7cLjAbVfMA8h5DwNfOnxwBFsinVn1lVhdTfmdtgpIxjh9eP4mrsy9G4NWVlHV
uJrYXZXjBbMI8LhM16OhQZWqvDf8FnY+7i3c7nWeagkDPYqbH1PdCZ1wwWslRMrWlD/FkCAz0HRA
sHGx3xL47A77dmam/04hXcTzBAN2p+s8aME8KrY6pRLgyMjPA5JnQY40GuU1lySrN6KIPaNBflNs
QP5K4aa1a9WagMvKvtSljg+cnWVJ6UVM0bB56OB8jYaVe/4ESnINCXINXOiPB1x6zME9gUmoTllJ
YafInv7ZWU0tcjiUGsaJipW8ciof+P7ozBRQOoY2tzxs58/VLmrvEQ+OR/Nb5zoXqXVR3ctR9o1j
ScI4vH5eUoNGydUkOPG0PUWXSHsNK+JGv2XYcG4wSRA+gs2GcuP3+t47+onb8fbITExV8fl2rYH9
ZHuTKJlrrJKJbNQ3baBmEb6fKjcxRRYAZo86Jx92fb42n9m30Yr3dFGIA7RSaauhnu9lwAAwMMbR
K4TYSoxzdaFOTw91095E9t/WBVKSfh30Hg/162djKEBbGDxg3x/4o8SJR4kkbD5Q0n/x6DaWEYIv
5aOGjTa6A7Zn15pWpj7bbFOhqkhd1o8esYcniQ+HzPyZ+z5fPQFfPSnEGUQ03A7VxuuQageD6IG4
ABtoI3HyoEZESDvOMoCQ1nsK/wdkBsNVei4hO6a2HGGP8QDRixpjXs6mt27JaGg5CB5Q1BI0D5a4
VQ9TKU9HwOQaV61tN0mpGlR8ZhhIbIqSwReYtcGwLd81EUcnS19QhBg0BO/pl4DF1ycWNc28HGqX
QjIUhhFXrQmdWFLKBDAnrN73Zv9E4fqyGJpzlaEIa4cRpxVYoUMQbJk0lppU4kZnQJvuTP1rcw28
rpYGK4RJcRoZ+a1S2OKdK6EzX3TZwEgww1/GLZBS8LwhOlSxJLl2cdJ/eAosG6KYfnkPOM30ChBt
Nzxee5LpgZ0zJefCMDiFuku3XXI6hJ8rvI4xQF/I7KrhrrMouzNwWGKnzwMVM3SIRwTyMHbm9LKq
35fgrw5HGOQlB8S098tuWq3dqngOItzqJp829K7pDXhB7+ukUZncDTjLb5zRwBN2QsFJvlshkSUQ
Yx1eQOOF0OM7VIdSKFasQzKUlFZC5VZ3hNhX9OVdsSu5D7HmRxo+rxfTBUJKNvxvWqAZbkLk3OTy
IbMiHC3zzI2A16gangT6FndUmmzMpdTVuVG6Tu69NJVrwEBy+mjOSQ4aUvb78RGYjNy7UsfkALhu
XmXKAwXIC6G4ZSR/UZRMly1qBO0tgHuhbshl2dT6urnzvKgOjZAgwAlQBznPaJ8u1z3PtKgjr1u1
AL2Iu+4pOItZSTQ4FWdDjAWPCa4ezT2W3SstUfdtD4pxWhpR/CkwbBhOaJubBJYnj3Nujx0JsAt+
HY6fa8GACkd0A76CLQ+QMbRy/hYoFGYqwwjbQlM1HUhq5MY1zEQnj8Rq1A48X6wXwtHAyS07BZMz
XZK0SGFdihA4BjwwL1yCyivZvh5kLk14ao7rAYa624JvhObNu+s09KwjhwNUo2SXxxwVeAobjAFr
U+FhI/16b6mbn8K7kUNQmxMKaz9Q8w+5y121qJ0F5F9z1Spx6kr9NswWxxSzxuVhsOEUMwkx8DD6
xb+CdVuJefLXg5ZC0AAvC70m2dSSvaXjD2NBwwCaTs1nXeHkD2Y9UrnRef8sGnE4Ftdb8t0VZ/Oa
c74c7KVlA6M4CZQX361+WoJXsoOVEbeVjc6SmVrL9Iro79IXAZv7sF+WKVJ1V1Mu+ugyPLb5ipZ3
iKlIwdAdn6ETiLSQm23keQteK2CNzvKDNxWxbcBLeGV5V9XWjXArXIOUA2IzLsnCK6YWJ/Hb9AqL
qN2JqiZDQPoQXslxduhZhQS+1KfVN0wFAF0uNgNh4qkBxacv+UExUmzVC0+n60gLLK3b6ylzMNkw
/jp10G41F5PXdZeMZc5cFN+2ScQgSnXjuvQYGOqFMPfEy/epdidsnBhNr2KLnQTCdK2iJGgIqc3/
Gkkd3i4feGQCMsc91EnQjw79wkhu215JLC5fGFius4UHogLVn7ut2zPi8bRVuBcPLmeFAlW3HbeN
KvqU2997k34soJ3JZW9q2+ptYxoLdRVfMx7GatJ7kOOH7HJAwTFmMD+/KnbxqAUPAEMQyIK2i4Uu
Y3A4gtM89xrDkl9197XWxujRIIC3ce3gcQBdqq7OxzZFAgb30x/ayRiFbeN1giQKSivqk/DonGbd
1HqZrTOLoktsz0zp/F3bkTPsAr4y7+CRptMRXF2l3eJDZK//JpzP5Nmv9xLeoz0Dx3GOKCNJ3g3h
O5U3CNiN03/H9wxQj8TOr32ZfQszeUV0TCs2Gvumj1jT86h4Z6wBUn6FScmX03wSof2LrKY8R894
ZqG+YaUAWp28vulWul9PmDKpcjRmcJcozAuXllPPNnPVjhuwORzhXGsfFaK6irPEBhYR+cZz2eCI
eJF4aoM9PkuUbCQgobs4htU/d0UapkKCWiPF9HTsyvOj5zESCta481HTTsp/6tjv5QDfNxP7A0Pc
7YOaWTRZBNasELuZZd6KXg6sKGtaoYDQKHFyGd151HaUbGtxA4MRvWOd7/kMlCIT+/GvFeu5UC/y
VyLqWt4NIxU25Mdy1kq7NR983cKgLEaCcGqTIsxWH0z9c6I84YCT4XYsSaEqihgOUZA3B1B4WV3r
j3AsXuXnH69ZeyM5xrhGdBuxmRWYar/7+3iOdJ7LsQ4iHvQidBD1VwBlRvPq/eQk5cDdeFxVRnqW
0wmfsMOG4Dm55Z8x62uvmq9ESP36WBnv2C312jHJnPk5DRPYaz5SWqbTE94CxreuG4yCgkgK7cpy
cKHD/CCjYwyNJMyu1BbFsg8evSE56Mf21LwDQNwerA6TYFk3rSqrk/uJWuNI/NoQTpHwHfbWoAv1
cD+OPcaIiWUtuKTB/DnN6n44C3F9mJ8ZF5d2x/opxjFyGEZLqJ73qDywzams+vqsHqtizIbvU/6S
qqiLWl6sqasCmX5XSm4/+ivJvGCryARpaFHP+wx+PyTwHuDjtUcoMxyO8wbR6l9RAsI66O4QhK4A
AxsRHaCDQrS3CisbTlmBuGzcZPyRz7itlw/Btwpb5R5NgDhUSWkfFStlRBckifQKRv/I/BGi8Xaa
phX3WzJpQDpIkMFu8shHVsel1Pikap8ctAxBp7yZ0Unpr5cWC+Fzu0DxGsl/wtqui2GDPjtRWkBu
sYGyGEBbB7Qpt2o9n7uXM/AOdRF6ieZCin37/U3gs41jH1TcRqFjoJvmR19Awc/Z326QPGD1oY/k
6pRXm42JzoBsjqp9VIElKzcHxyhyIEaZk2HFel6Wp8qMDFOSvICHaWzTGxyq9Qop5qVvFRxj7ytp
Ba9XKQigmL13iIEkbvEXNihZYmeRFR2WKeOQns9q0e0fI3gClc+y4UXvDv4pWqT7dg/A2SI5DH9P
GPnWsZaRyvK4MX75g+VNoDAYjSj5nPylOY0aBGMz40ws+A2GLklvrcuTQukncx5pZ+vrezn2xOmx
icfeQ6LacBceCKeod0kNnJvxVlz1CgdLlMwUFIoyRzOdVW/jMNcQFZkXlEaLmO8paneHJfu+GfeU
KR/kaTLOPOclaKnpwU43IDY+yijxaKkf5G0gl7uQ4ZMQf3SaHG/lV1stUS9qu5EyZPGLpjHC+vu4
fDafnZ7kc1tQNapzmlHlvTTqHoEZt/iKYBeODlcFawZO0iXtRtIe0UeZq9nArGTfnR9VTm8t3vFJ
NRYxxbBunaUGQ1Qs9jIR6NwHYpyuGcLe+jKrzh/NrV290U6AprCCqC17Sx14XuGfwOEVGiatQxbo
X6V1Vrx/QDGNcZTdXzvOXL8L9jDK6xxXz+Er+fC3sl4C58401vbGy0h4MLs2ax1bydUxyiDBxxfm
ypxMOHEvqu+wQdMAEV63OXfpFcq9AKA9PKSDpEiyhObbUk+UjT4MY3YjlHpj6SiLsXpv4Y7VhEPz
TwmqPKDfClPZF3weXiR0kzvxgpVzGP6mI723jwd7/1ryh+6u19ouVdxOB3/UGOpy0cnW8Pejpin/
RuCtNP84kNqqkIelaN5duzlZpIlB3adtDrW/kbKdygDXRydBJnfi+pOemcG1W5/Mw04s2nyFfkbv
DiDPFYEJ7FQLTYfOkLu2wwbOhVHKhffNl8+8h9G/YK+yxKyGNtlV95I6H4C/d/XhCfYKRThjtlnp
oLW94jzgKHYGIBpCnrRbeCikv7Jn6A3mDGsLxkOrYa1o77iTDocNVfffHBGJIa1ExNagxKMVQOVl
Vo/fzUlD1DjI7GMxAQBWW56sFka9w4c+cdyNjWdeOLRR246/LFJiFOF5PQKvz8HOrZV5RcCRs6rn
jwy4DZKSEhceIyzFiQTWqJmbvJIu/hnfX3xMGS8TkkDsKX4X0//bfBuFbU6GFoo6A1vpDYaMsa2E
bDI7jOwnXh3QTonHl5pDMh5usG5aWnCXl/ivHcKYtWVKHV+55ZP66LzvYu6XnY3qYPZZwzw9rZai
Bf4mN+nl9UfAV03yJuG7m+kE3vtbgPWF0CC3QPSI/9+6cyxmadhQmos0ERQK6wCTVfTr4Qqq4ODQ
FO42vIWVbJJTH1d4SmrPoKczTExwGa8fyhOpcQm7OUuth5yheE4p5YpLMqwGgm5X94w2651u6UA3
ZyOk0/FmjJ/cdlz0P/pFnfrX4I51JWxBXy74NHnSoqxu0Ck9KM+i3tx5CCt44n6aMBUNUjAaBXuz
TPmFOagEubjpblV8ipkToSXz7S92HGzKDUMTPoT7jZUV+YwTO6nn3t0KkefKpvS/Oe5l6FRbVlsc
uIuCWPMBZHxVdVryPvtPNuhr32Qb8hriGZHNQUxaCFjMc1xtz5Wyx+gE1qbiPWl9iT0o/huSANMz
kQgZR7pbCvkg4xc/XGs8cPgaCm814bb0YYbiCXsHVqoESZUsF5ILGjRa16kuXxPlmdaoPTEA1mHZ
fT1WXS1pijwVELOlnr8NoWuT0EcrHOUfjXKLClPYIAMAy1sniV7m4sa4S61//mGy6ilYrOQpMTUX
iIlpx5G3yHEQflVnEobpA//SZ434mqCRBiHlVOpOwvao4uHNaClEtlJq+f9gLSvSLG+vvY/lr012
rJxwhHU/14nln3FgDjGztdGs/8BtEJtcdK6HXN793/RHlrHd+Q/R4yj5Cg0DhLBi6SwUYKavBWzB
HwmQmGsWgAqRTVFl0PTPY5o0ryX6ea9LeGS0Wjkbpnsq3iDuxRdARU4Z0BjjMToR43U/geRHfxwl
CEDGBrieL+0lMKsx0mW86XqDg5xbuZALwXE4ehke2wwQEcdJUXqWHXK8aEzHbRczEuaeIbPCubMV
yxYwZYOZ7wn/yVv0PEsqq/zKS8C+cO//SpImKX31/pBvG3h2LKumRWL/dkoswXD+rKsAcFEDeoky
YkZntP8BDok7wcpeaN9Wji4+klNMBNVyveLoXUDsyjVCrTQSRq+kH0Cl37aK2HWRIPC2cX2DCNwO
XrB96w2qQ/dfqTo84hAF0G4obeuKFkFcfowwXovxJz2TfaEW7aSkF7285s1AH5DWeHIAxkbIVlit
99ln/3r2MMFIoE5uOovPd1L30DEMTDr4w0t9OwkI09BB3mYSaNuJpksUtRxDogFO/b4pS4lUK7bP
sH8wYFRT813ZYr7lJjLyVnlizn95Wp754d3Magq0LkJHe+o4BZnntkOxS1EeTbqvqxguUeR+tyrn
Zalh+yZNZKX8x3ktTxFvTYTFiSdaxuRhyEYWNJ1QBsStQiUQGwTr7E1/c0xXtFucR458XFrYT24c
tAZVOVs59tsJsKxyF9gsfnoxqUNe6gCtWzPHUe64R1XRfpD+jh62nWnEz5rGM8NR5vL7hE1Q3hII
PKPr4FKz2BAtW1h4aKs9yd+ZXX7hBIy5d8L6KDDTmQHIg7eEsH/qZyo63mnQ+kpL2fP3h93PfKTN
yjLTqys41GvQ7UrUS2opVqrCS9PReE1ZTUc0fpdax4aYbCZPub/sEn4ApkaokEicQVOVFmVankR9
LEst7EYZc2xUmh63vNqPX+E43ZnzRkQE/r9g/+z8497PSyGOsclQtj5qjBaXK41jx7vI1OjKmcl1
GRny0VBDb94223KskjpVdl2z7IuQ2OLd3xFcOePxuTAZkcmVm/OV1i9h8xp2B38tjuhvfmUrTC0V
Jj0L5X9QV8yfEfPw1wp8U3yXY7F3GUmL/cKnu0PH6Zw4GhE2bg/YqdKt3K1++lq4cVIuKDYEtAiS
3C4NcYLqUOFvfdnMqBgd7QCPTHOktqCms0HQgBF94pa8Wn67Pbeah3OLr/mq/79UCmjK88NqLEBo
bB/NGEP8udnubv2iGCHEk1hYsL8+VTrMpmhiEbRq3pw3jXRzZRzpfxB2MEs8u0NabXdDIrq63VlI
5LoKnYCH1R+juvHaby+bG8y71U5a6fJz4I6A0PgIj0cEtL9Qr4x9QivP/NBSrNTFW1muZmwOFBOf
Fy8F8ApUhN1yg2JVYekiQoFIr7z6jAu9ne8MdYCo7PLBLRGQK0cv/voVJBPF7EGdCKARl6s4XVBW
OUfohVtnU9HFDudOI5yZwxjLJgR8sECI3YyCIILWfMg9maWhrlp/eRhwKiyAsAx5JQa7YsApi4W+
Pmao0L0A/owDeUnTvLwRCG4Ofse82OqA9jkU7kXY/j3zksXuXrFLBBBWtJU+glw4Pzin6l5AivEU
03cwZneTuDUAEc3wEeaF5216SamV+5kUykBxEYl9Aq2DIbvCGfLL37/Eqju0KGJ5tsDRr+MM6VPE
BsxXmwZQT+PcdcH7CyvEaLI4/hy217lzOxYSNIanZIF2R2ZjJ2P61MnjXt23s1t63RCWRVA1mW2t
zRNFXZ+oNrFaSTLvxEWAiS3JBLRjl3tBk9M5CDue8YFgImvjUDYYG/H27ZIHu9LVCXCHER80vey7
Q/+csoxU77GOn+ks4WXDpBQjBm3KTnk5+NhPRcDMDGmf2Y1ut+Wd/Pm7Smi6sf+n+1I9BB21P7Hr
xzdGWuBE75z+jzL9EiEOo3htjPicEZx5cVVHmp0GhlbPWINshEV8ECNANwRrTlBXwD4Cj04AJHuw
eg1Spb4nKUqeVsw2xV/KakvgV2FsR32sdhtRW+UwYE3qFmcapKs9vugqT6Qi3tLa1vvvDpMRmwSs
y8S+9AyVfWHUyC8t374z7vxaSkj38x3SRcBeVkeoal5qcCiBarZ+ODFM5W/EFOe4ldPv2y6Gog80
/K5ZGTxzm56X2UI/IJhw6FiPnTXLvytYTFqfHmnM2tpkQ14oTQI62Pt2Uwh7SQW2VA6IIiOHC5KW
gJ1kL3D9WuqeYQl87kBYdcSMRPkaCPHUIU3Eq8B8sTT1PqQhwDRA4mw9/buzj3zYGBvb3Vke6pnh
vBOpgS1h21WY2lAHldmxn1xuRr41yDkWvabt1rqBt8igRbLgg+vr2ysez6LKxjbYIK8tW0/HNv+V
1OSCw0exGdLHs4phGEoy3riLk45M+rsfJBLWcmK67wTSSQ3oaxPqcHUhDnZYbBJ37q3yTYHTPSVP
Y7QIjmabg8GUzsOfQxIHQBYJ1dmRt9MHjTj8bUz/yNYlqJIF2wlhThihAFF11kjS3Zf4tAyO5r6O
EubkaSb3o+5+xWp5IK06NzMLcl5BDBgsCjvkj2MRmFGSpJi9ulyX2/Gfw9YSKrnF7y77XtJeoRZS
BMVtKJOE9A09ZM+Wn5pFgnxMuAR4Et2u1PNpwA7hf7HI6a8D0HIvJwTpXVvd8z8kf0YwUsdT+Y/G
GDHbXC5SzCzmP19y10XlESJ9PIlhJLPXyVqjBU8NP5S4tc6Ij9tU48Z2W5/ThJX9n0Bj5NW8Bfbi
4BR3QiqPG9KY/Y8iTmAr8rAhvsqJhQ6ovE7UE7r66G3pwW/AYSQElfnBva19ltCj+YZPpHTK3sHL
K3O8YZ5OmPxIK4dyx8ZrkwZhrxv0iNp/gZP5k8ygt35YGxOkeLm9ChqtHgi70VLxOp3ATg4SYwti
8eSiwENC06hox+E4TX0PSyObHKMiF2O3pWSEAOA7icbZG3wbCP8kW/LJD7GcqmX+5XT2ot+fVyM2
+IJxE8DIrg27SROSta6Jo+lGXv9GJ4G7Y5EzllhrH6HZhFMjmB96VUv26Tg/x3Mb0KnG7xdHF41i
oGBhzfPxEBxhoorfiHJH7tMicWrkWjXhxOq+Ozwd2Nq80YTOd1N3BHdyI7Txg9g6YmFHRqlPFNtS
OERsi3FcjPJuRsFU3kqAAepql9VAjmen4rNnfxr3dYuUFSCJthNt8PS5f8cTRYcDLILrQfrGY1zG
9ZHTufgtwcv48ExxxB/fww9v6nKzUduwPxpy0bQbSd/QQaWof+YQMSqana33Rlm1tJudEFn4/JJd
WTUqeWWES524DSamRgJ00qGMxkcFGUMXqhdtPtsZTO1oZBO2vYXpujetu+EWz2VUtTr/Dejc9Cwi
8laSrAckbVRqL3xdY17jCqVPPM2C7Qpf/guq+JafH+xbVrdlwjiyYS6FuCy/ns06Y1mUmSHnoHlR
kucPN6N4J/kHjafHRUmwMuZ9k4X8yIWLTygt9Z4SAI5wUuUc8LG6FDVrbV+Qiukk9MyRN7rVvtnV
/lZuvwKMhevufFa9w9H1ZWlqkhjV+qNw443z3MFmp0ECHHVTAndhsbS/E9YqoQfBcalhXRvhl+6h
WhE7+WSvFGxovkgkIrUmONvdSo9JicLn9+JHG+wodOS+NIUerGXzUT505KJ2X8LKmS4eavthS7e3
QFi1rQiy3NUutU3TN7B4lWt7SJBtGqV+y2aVKdsO7u6R9z2SnTykQC/Fgx7rwUj7mDVZAlel99dG
dy/UzcjbWrxfZpGC3RExbhBlhjZ3+sgEroSqVQb+a6UMj9PcixF4keW6jEw5D736VgJpV9gbZ93s
5xoWSNZekm/DvDdRz4WeuqYMJGaO3OV6vTQrn1TDMTPCLCqI6vyPdAJpgW5hoVu10priOmDzNcNM
Pgaat6SLf0bgfFbim4nX6FlOUcBBualebhIPIInKMGR/5EQImJqLHr+S5+oM+MLHmB2ISULLxXGj
BF/UfalT4BYPQbOFsVGhHO2zuVhvOrjuiLMvUmH0ukzu/bQXxyObVdCufBMG5mBWeFJmQQYtRV8Z
P+JaQW7KLif1qvSz2eTWdFjq18DHGK7uhgJIFAok8MeHNfM6NWo7UcdMrW/HDywG4ZAc5f2OGCbt
U5TcV7CuFoCFoUhjcm0HY4hQsawle46PvZrRAdlV/vDcArWawUlhPrraOk+CZ7xqOVw3T/kOK1r4
32jrzwfdSXH7ld3ZY4O4OTNVn7HLV3F/dUsA/uw0tv059N9+MYgRboxnoCOJgKwKOPJBBF/vFcYO
o2mqEgNnRzDUOz1Jysq1KXmPQOf39P9ge8q9eaQmlEGznu3dSRhkUWtlWfHIAigjI/+qjjNjq4TP
Vb2b31okBxT4D56O/dOFr+Fe+FwT9hVFpfYh1CUybGXUlqbkZ0fL96D9RIy5bNhCfz0ob9rYkfXo
MlyzWcI3eLex1uv4wdYNHbppFEY9gUl+AK/Xa3WZCyVFz0rGh+Frl5Lild6sDkngnolMsFS5Qcso
zTMFxKj8LKYFxGzx94Hu0GkUoJfl7q3d3dwJVrKtYKdJgQNAp/RJKAfvO61OVbDviAgS7bIs2ike
BDqjUxyvCb3oKDBXb68uFxdiNeUOdMJucMlaP2aaNMKk/fMj/lNMXFiiFE6XQLbKYOWiwdCW+7Xz
NftxgQ8UxIwo+uHyNkYC5oyvdDuM17Msgfx01OeV4k+wwj4JVXm7VDnlcvlwtPKgg0usd6PcPjM4
KN+yaYa9IObigWJWHjzDygTlUK+yQqPDhv+hMOJE4ITIyNyLKs0SNnXrZzUc545UnnwVCkT8tf2k
+eKGAr9zPnTciTRAal/rRqCrXIaWWdm7zRImqTn2JSml0BC2Xp2G6HlhjO4snPSS8nNChQB6Hwcw
6zjpphY3vQNT5ZkUhbkeHkhKOFmDfHvUYmfXTJsvnGINDh4RMuP93fMEUk/odhcZrTutxU8q2/4Y
wXpqAMFumn2g6VDDDjsRJurOZmC+u3PXCTwhmrWWaVbbL65I+m5zQ1HzPmEShv5NyOlCepR2Wyca
5Gg/xEeoqRs2iWzohNYLK1eocl6N4r53SQki+ZhYjI1ZP31WEjTr48poqJP6SWZ1nGIMkqjxZOzT
eebhza1g72NiVJDmYXXHBplYr6erWxbfRtwFd1H1XsGYdVeJxCpGaDXqBg1/Sn5d9BAX5I9smwb3
5D4+7fS67W6V/YPIR5op2WljHsWtUfUMPV7XlH24rD2gEL5JO5wyM5TOiPW+hyPCmToTW7YuQHcp
BIrJj28upPgdn9GE1VPOJFSrIWFWfW/sa5Dwt0UsJSbTZ2hYt28a8PafWYWOjMXXUeqhhqLMezdD
KGA6o3w8JpjkRzwd87gPJ7x0jPROS7akkG+fWNYaaOVoTzJfSHRj1XeVXzyoO03lrJHkI6rnn++S
xKctCJDLi8UUa6Deh03F9wiV2I9dLPoQLkhiK1WWmk9BwKx2/th1vcMul+DEa8zNDWJBMj5ubftD
sT5ZzKT4GDgfKcA7YY86+sWuZPCaWe23QhajCMed/2tU5OBjkWTmaQxFpDIg7FzdrcsEaVG4KuJw
ZIu3pC/D5go9OpqyEVUsYjeqXnHVCQlhlFmRA4IClxVnxYyrthh0qfNCz3uceDlgOjbRavLVDfiB
FbY57/rLJEgCRttJ/rRA1+avH2tZW0HzRJfPoG7rqyYkbuJ4YwoN1Fr1cwWOQ7vbik4ONujHdwus
rBLQG9tS2WLTQQFttgPhWzQYh5h9tHkD8XnYZkuqNahAb/ndyTPBBWfchwGsTFvxoum5y5xTNU2r
9nWTGGLhj5O+MrjgGYIYmtyicPSUagFYfKQO/IJCzfZV5IRWOqBOtfKO9n4X4JxDUcPOVudjF6Wx
gMtAfUnu4ctFAy/zARmUyMHEd20NNnlxuaZPv9dz9VjszXSm3vTVloy0M/qXO0q7bRML34bUL+hZ
7CtH+czPXavfxP/dDZ/wXuC+wzxh8eKNvZKi8qNffio4hk32Uc8MWkeZ0ocyC0mRuSzwc2ty2eVa
FK18CaZ3T42x8gaY+LZDW5c5l22cJoV+/hPvhoDABUOrqVvJ6veRLcqeByImAx25pjH9lJOCvRXE
g0R0RtbOl5rVEvRRQSCxstBbW1dCU9JZIgIbHjNB3jhD2WgFfWXZrrXA5+4YF2RKJhjGu/JFq8VF
1R1G1oxdk3npE7G2+1/xLCC9CJBYPnYl9Tb8QTEw+JrCC/g3XBUgvO/foRbak2uNWsR/7CMFvO4M
QzRRdkQ8Zmw+htkflrETo6IlNLzxP8esQtiD3g6UOQsYpUdiDsMyVaOJy/G5m98WLAiVisLVQeoZ
EpUhLY8xKVbNpRoh197UTNcmcMlYma4R++MAfbI+phJteyuPjjstlf7DnHef4FyVJPkctkyf3kEd
KoJFyoC2/9tpTSr5nxlfP6nZ2VFJFiq+YaxpEC0/eVBfui241xQFqQeA5lAJZLa9cNXBd1pSmB81
ZhuMgyeTw+rbb8wpOoJuEVruOHckzOEWDmPKPm328wXPWmCWBOpzgvOzFJTvrgnkTh3YhorewOH6
qsdBJu8kCHX1qMdZcKi7wGrQ57qyyF3gRJOihPdUNuVAYMhN4qaQwWUEsEFO/4ylyZT/f6hZYFFt
r6L6Q7ng2ht9PhyYnd+Jxe2AvIFoQXREY6UZDf5lY/NzMrNL+r5QJon4xEnP4zoIxl2KSr6SkiSX
WwjN+LmtDyPolFomhCpwpdIg0eHDkjXSaJxwdo5YHZYB1bIOrRMjiEk3sJudcJAZb9O+HOynjOi6
tfH37IazJHWRT5oAMbK4N+7sKD9pM7hGHEHwRwqL098GKd39gYRa/3c6TiD4XIn3bqNZID7mikB/
T+hst9isyDvEDh9VrqnFA+8thtG06jgruh5XU/a6OoP/q/lEjfT/qaBaMcevReAUhHj0lMr7Jmu2
CatczbVY0rVxpO81Gycf5Iqm7LYLvzwyslOFqcjzJp5yeRu0Y3y8N1+igXAplmXtzGX49WgyCK2D
D9Hwpe5oUr5FlKKjSx1yDbdJwT2BB3VrrEgC5ul3SLaOOAFo3DVdO1l1/ocDz9r25ajhpMUnSuvu
nCBw2q+WNOjSXzAwrxAu+0K3NivX+nf1+GenpNPn9FGUNLXoNYZNYdqghEhI3mg+e88PrXPP2nva
5RnqRQXtx3FLabmwxtkgPGAf26ncey/JZnAxsjEP5D6c1UszfqxRNWzrtnvJrUaA6rq0bg/4Q//p
5N9ivVwaH784HY4oyp6AfDMVXnPsKZsAQ4tb9Rpml16JkvqshR0SOnjekHohxoDF6P6n21hkrnOD
CzOIUdSPC95LTbrRBM582Chp9XUHtcYMWrROE3bn+gVPRr45L+d9nFZWYmFK0esKmQ8AgusBiLah
CGws/dycVn1lTHiPHcTYum7D30n6L0fva8PqeyLt0LWof7sDcmhZgci2kKpm+iLnzXkJTyBglqj1
cJgguzK0OC/Hfo8AtxPaxTfz1bW2Q2OoFgh7hEfJIOVxonTWtRwNDQCLlyYnztEfPzEsT7tLri/p
RiYhqnoiHuwOJrhS978Re4ucb8qDA8/UzViqjEZ3DOzHi2BZqjzQFzeVfJxW9RWZwtZRewvHIOM1
HwQCCBvYf6lKs8cx88QlLnJbqcYXl+8G4RGd7sD3J7on87etL3JG/a1pinWiUIoAKYE+dKz9nd4T
rdXnXUlkqLY7AiGunEyGnDvdfJyThObnp3u/H0aCXGr6U+ZB9u9ItOKmAndSFy7DA//mak4cxNOA
8M9zkKh42/6WYBPHnVypfqCNG/GxiTpHuAC7rVJZFIjvDNoF9BiJkr/NMSkIVYHPzUYnQSKINIvp
8QvU5/HM/AkKi9LkiunrzsKqLHpQ9Y1N3737G+vSwBvLpFPEBuSisohAyyAf4w71isLLI3O5ffh+
dY5oDb8yntkeOn3SsVenQG3NP2wgO/O8+xZZQTau3CzJVd+T/i515HHnqTQkgfn04orlvma4PJ/m
yP1lQEacHQrZhM0QDqjX1zTS14omFqmxI2SDJnq5ptmhUSU7MHqhUQRdlR6aXCrbQRbD7MuBqQ5A
amfqj5rBIUcBct/KNBa6glrMh+flJ2KsJSLpRWZ2XCRwlkavivGHVcEbUl6SVNT7og65/0ztHEW2
bMhLDGrnRBJ2HnFX7JZvIxPsiL7YQOdGGKTtSnUs81r5XuNh1y+HUcR/LgBUyJ6zixLloNGCOL/S
DOzB1gjkTykW1ZLbE9yh993KpquWSqEtTTFTsaNtXOf0EgDY8f8xEtCgPkzzctRsCWlk30D5qGjM
xJ5egwKxcu0Mo2L23lI6FJTRJLDrLlC5P27kDzmHsRhl239OcN5jFvWGpUgbnIyd7kCsCMsW7q0c
l1EPKMpVTqoeCAEAWsjrPzigpEQA4f8XHVO2xd6YYzMGLWLq7Nxb7IP6M9XeOW529ELr3aD5rYb/
MhzCkQsYt3DtC1fjcplShoHZmpOInnbO8uXPD0btn5r/D4Ksais8SzKKaGE/1998bCbblnNDNLK+
XvUaegy2oJqet+Pv/JgqLHQuYfFMRlg1FOXXoQkoxbLzmGtbaGPfUb6WPQfai3vs7sgkcjpiO/AY
a2fpwRdgYNvpIyybphmVDZla19+tysW2vrMIS+TnnV3bbRRxXMbEKAw2DJ0eDOP7nbKBDwiWz/kW
6cKMmteY7G587ehXeCg94lxXegBZcArhyyakIc2yd4s3J1ezUSKGZG+V3xQHMrlNMWbQaWJRIafl
KBz8ZXEMnWjcYSMpG8PGWGYBDPwkphweYYZv4/Gnaf3Xsb9WfvDXZXFMJQMMUPwIargizRU2O+aY
9Bkg0F2xdlJH4theoJImv38eTZ41+q7BtOTSQmqkROJqUDh3t+T9RB8O68LXBLzvVdIOMZ4sB85y
ESg2A8K3bDSydG3w0g3fuiH/mlPCzT83wRK5nc8S/8QwiatTqdOKYnNMxcR20MdyLLO4hW8UkzgA
OraMeWidXjYKUqmpshv2QwAp5+100XgG6ISqxuAxo1pPp1rAGfWa1bH+Qm+bF3YByXAnTVhobmkW
TgyOyr2i+olmN2OWp3Jf1uuITGEoFNp6vc9ab6hTJ6LIzQcaTJY8MQiEgaVordzZye0q/A2wjO44
/yeUJz2ZO8REWugxElNXENzfIQ8NjbfvMmZrt+zuH5E7J4PcsDkLX+6oOYa0WtyMOtDdhMAY3/UC
iQCNRhhDRZgpVZX0T4TZrcHCjHoGbw5HO0IiF0n4T223v9t1I20WpIZTy/vXwbYIo0K2AjoYingn
GiC0zkovonn8ojPUFdxuzrbKK5Z4upZw8v6dbwcnwrl0RWVfaq9TBW+I65GV5R1L4IPQ3IGlYADc
WvJj1QLWlLN5Vh0E2x8VqFcRDQ9WqDQg45wHbpqA6XSVgpWO1xIT1G+T+tI0QyN+UnQBHVTnRIGI
RHju8sqdNgAstJCMlRGNH75VcQ2xvayJBh1ZOn6/arJ2N+/anjd8Kealk2trLoTGgeMRW6MkNrJq
LgA7EjM5MaQQH220pY1s5Xu4GRkpy6a3eUT7q34Dfa72G6zH7np09ExXexaAG7oYXyUioqFnliMF
kZu/J7V4QygEJPPR+pixBi6gLq2MWaCrMiaLcCVnoaxZaeLSCGfEAcIVDzLft+D5q8NvxlaGbs9m
SFNAXu+D7jod7j+uI5HjXESR0WR5Vm9FkoBRrF6vj0Yu5rlWhk2GzK6jkhME1sAPxD9yHsxgD8uG
e3UjN07tjyZXlbWIkR8MoWYRrefsL/NunZK7DtHmIwOi0j4nL8Q6MNImAi+nAZge0eq+6//NbGAz
/r8/6ew1sg5EY34mwLqk6X53kqx4HALBeCROVeDMfLqaQlgrX5uHS49YkUmIxnrYlNXyDxSDezZ2
9u7J6wwL6T9vdwmVWfT//FOPknB5vpeBGjCPzNJutrBIM7usaXGn2slIFXhpsfxAD77mPoekZ5Pu
DuvCde9Z95ahh+zPlfMl/2ea8yInC57/JVfb8ICoalMrxOH0aw9fv2nu/ij30l+8tXcB9citrEWv
2ag5zesZkkyU3bfBCD/ByWJ7yBCzfLGKWjp3KcD+XkMufsmDNFD+SPlCutYBm2gTunqwBuMsiWlO
B9I2kEm5hdHeVMDfct0Vav3A7frQcQObrDQqnFm0bllb4RzyavuTykBcB4XoFiHecLGEMWGXXigs
V/M4i6KagYrFz1B2MDkydumtYx4rVBvx9+RzzRLxhh1LtoYUIlnX9rp2fR8wW5PFvcV1JWA4l/dz
+3Q34fnPRY8UpT1eJgo3BNJjW4APb+HCX434u9t/44vcJrQxhrSB1DcYxxBio4YRSVNVnkBeMDow
m/QGd1GGsUk2Jycyb4jlkynFPxPhqbVBZ40+Gl/KeF+AkfbowrRvSLW4cncOSgr0VPD6v+CujXne
D+1KG8RL+w6TzZ6Ff/ViZPrlMGSDLdlAzMALOec4KsB45GdxoefKNBMmHG59R6Gai5AJSqZXPsPo
K+Sn4FnVypU5Yf2cWp+IOYjeMk3hmGz8ol3YzrMpBVyUChePCtkNYK6osool/s3fXM1MpquVNjK2
T22dwYQhVj347+02IvHbijMsmTIGRniCkrTQxab74hyv2o6uMMNGpK5HzB7syWPZKtQEt8PIfueG
b3iIUfy2TsNlUOH8hDH/6q/2PmM0gCgCckTudN/8XYy4mmADwCkhW/zymNsfgr2A0ekK1bK2vMaN
XGjlBiTYGGlbMUWU613+WybgKiacDrtILQe8eOiD8SsHrWfrBqbTiGwHv5QfKbvC1gn4cja7n7V6
AoUfeG/dtvUFeAnt2wDMTHjcx1YFMczAo1KX5dSdF/QAPCKhOMVg5VYDYZ9xjRqM20QkiBZEo79D
sH7+Mu8TOlmchyttiZ8wR4q1/GVDulgSgIJzpIeGuKIN8F1ZYzJWiptVpqP5dEc+gAi8Y4KWN//l
DARIk6yhH+L13K8Fl7XDCcdNU2KkoigN0dxTLwak7otUMFB3UnNptU8idOsIkRgFgl31c2PNyqXm
GI3fVKF6Egr17FUglKx+ddUGZFR8BxU//bR37w9ouSqPbrQcbEjbbN5jYTvclsQPD6mLHS9ZC8Vr
ePvoBVXcU1tv9gyT3AXBONucjNGkiDY9Yx2sJDOav2gmCl8d5uXnjsAWPAm3oUCsKYLqVwthAOLZ
LaD6T9v4WbY6Hf6ZjXXOSaMEb3Nj0yUyxnT/D6RW2jqvUUcj4Mo80nU7C+z12wGblXSPrB1qYDp+
cQtOn6zzs21awe0R/h6h+Uhq2OovYRVyGiz75OzqBGPAquC0/WHmg4BpZBpyXQ+xRTYfD5707Uef
1ERfncCM1meHBQNRjMdoVx68bWawQyYI//zYzwjuRJCMGx3bqc2vL924wny5Dpehitt5zGqtDjBR
eMi9y44WUGmOmGuhhMKNjJCHpISwp2a2DrJ5vUw0QNvEyZ/B66X+KwUPcvGB9nKuG01M2/2TQp42
8TE5W82nYxVBbGG0LFNWw8gq4XqEOlpna1tBGL9zjEa/fmnLmbDh3vuN4XjJWcqzGlqIJLuia6ZO
NxqCWmbtWHc1d4EXfvAGS+zVjKPgQoP45W8XZAo5oZcRd/SV8D3FIlPd5vBRBddpHdtAOWNFJeKF
emzLZDf0TqrxLgCNNigZRZJlWtzeltuoJeF1252OQWqqva2LFkemtpOFirVOAAOWwHJCzwWzcMyR
hddyGicf+ibJc9DEa/Oy2n4+MkO+TNiXLD+AH4t0nkzQey53mBK2zYtfgPrPXj0L2PRfOoNztnrJ
rBzZKd66gwtl211XEfgCNkTsenpJYgcmpOZvfmPpy1Qw4MqNnbpFfMdn2NRaMKXxUjIpVEV+hPpp
Ruv/8cJT6Nb67+hH7SrKMU+Ypcu3R5OAAXfcgYwh2mw50HZiA+MvnS5QowIF/B36s0AqolM6p/bs
qAcZOHjib7JNEOIUrJa/v+oxiyC7li8gYrMNP65WsRC+A5AmtrBZr6+wOpZXUUksOkIS8JWZcrYW
R52Wwf8yJaLKs5XSNNpu8lgItYNNIdAHySU7xfcGlRVeJRYVMOFdRRz0l4dXsSu3hnhb8zWCtsxt
t4UTKqe4fYNxZ97pl6am1N56l/a/mre4FDL5/OiDWcTRy6JCitU9LKvoDTM7snEJj/6/FCKQCX3m
j4yeWzJ/PSCjHKVGeI9duqivceVcny8eDjZoiZwpSTux+ElaiS327HJoQQJPGKDVEmlkvItzZDHh
VPGlHK2baANeH2KmuZM9l+dHqBkhXi5b6J1/lfV3MtB418JXjq28Pmr6jKMyw6CdC4hfsIz9nYnU
YSVj8hEoR3t+LpC+iVPqXdAHQnH9FgPSwlkTDdT4s/Q8q7YJr1DAmUgXlELiJalTyclEhcEAlGba
3h16n6JVSKWbZi03ZhNTTXjkPEoJDYIVcL293GnGBg/gA4lyAeh3pVvX+lAe6KabjZdr8D6QZuJ9
iH7myrFoFFvZwiVFclOxEPaoK67NtyhRJfuJrapo4LRXBIsYRZQFuX6ZQLXX15rDVHGGa/zGM1ta
7/KKjceBp82Btq3mEsY9ncidUyuGb0CSWQKEKdD9DSb2HW3WvL9BU/taVoagq7Kdb9DjTawa4aRx
gSndHnecdKL7Agj4Y3DsDP+WmJvD1laKlCxiS6xyam/1zZKltmqUIlKDO3NPF9hpgDam+039Y2XR
bfetLf3UnKjv9S/qbEYoEuI4RVFujYR6rgczi1a3tGoUSvRRG+KdI0AtWjxtyybdVIg7umem7nai
jWOSVaBctNediwD+qcwnoSVa9U1WQRGXsYf5xUs6d4JCaqCv5KIiGuro3G2ORH7pe3t2L1Pfh/D0
IALVG6hAjhiEABwNDqlaiZ1fnK0ROcQvpjrLZ1jZYBfKmoUpwvmqm0h4UKCb/V2yYfmWkrz+6gG3
R5hp6pey3eHb57JEoKifpYEgF342W6M8IJaeZURFZW2QJTrIY3BqBzNNoilfBHA8abxrp7I1EgDq
u1LKQIenoRTaaKwuFpqZZ6ty01NdUzpxnGRPLngvu18jvw86I6m6a0TqbrfYQwKwJpL8V59TeyOk
KXC4rv8AHG2Bj9UkqCheUhSbZAAPzBM6WiveQhmIVTOo2VH/Tc1kYiiWxjh95/gUwjWPXZc6WPjU
NXNKZbd0dj1piAp7JoL+hc7qOXO0aH2x1SkfBh+hhqdDnQqy+qqdGxV0c5DkGEvF0BEn6wXzvfFU
ee0lypki+BC/lqh5pvNuPkiX5gPENXiqyGitgI0x/+/1F5lK6p+qUqrJd6r7K3KT1ZBLmY0ZZlNF
/JbPjvQJQxODVy01WcCC6NZtBNaAfE/BH4zMdOYDIOv0+YvXT0vFB7cUDx5tz6C/wvogaHg99TDV
nv6AeLnUGS6QosGPDFBYTffh8ORvvfi33lcrorO/unIrjFJHqsRxeij5DK0Jgn5BUXzPGz5qHs7J
pjTjlrhi8VoD2ZiIUxlw6FX0nkrKTOUC/qfBJSic+dvJCI5AjfJhcKFWspSSnC7q61RsvOUS915i
F9IZYNs5oDMrV2JhYed+jcO2EJgeWlLR+790eZ+LNqc6vlWQiaXCqUffqGpc2vAh6AhGMaSiP74w
g1Yk7Ws6bJE8ldP+3aWivT6hWPTWaVwcEd68TyDTA8uP3MUjk2Jasseb6G2HHAgru8X+fWpJEUHE
asoq5271JOp7otUJ+tFCb0O2Bf9JxgVGkGnc9lSs2ffrwfcJ8fGpjwr2nTvWZcal8VLahh0akJex
OartLY9UcyKsPtWOVtIckuCgLqQxZA6bSKco5y4r9uL/EPo6rkMaosCtahhlbaHWIlC4FIDjlnrx
2rpll/DuM8OwsBETvCtsDpz5oVI1WzOwOj6sVTSBkPEO/t+8Gz40+4VlMY7MWkQ+B/QLd9yXJlBK
NlOYlEjt4esFautTHF4qqiqGOaUt3KgWSzVlUcJcSg5nC/xO4ycJZGeYtp6rr83WW8Z6VZDTwRei
cMhg9jxec1WbSipDNhH6vEXkHOg+zMtLxJakNqlTrJU889gQVtS11eZlAmciWc44URVsCJswMk2U
BXE5EeJWLhccOJNDmtaMx1W2Wv0LlWzNe02ktSDvQRgf55VX53d6r8aCJBfTjvaX2hgkij/absDK
uDrh/J/aXpazopJbTydFcaDvXivV6pq4mLyyquSkpAqAyJhelDda22Hc1ciI0UKU3oiA9ViPYZ5f
Mg6AeSMM5lyWL+p0XhpOFlFPXTtIqHACfVxBoOgpiITJ0+8neb/p8jfQ5c9mq1F6t+wv8YVhw490
nt26X5f7KTCBMxdSPYImSpTGexZJmM3OxPycVot7mcffVdqyozh3Rav0qpnnli6JdoGK+XSGkyPI
f3sUvMUfG99Fh1XdPRdf4lB9UB3a6udIGAnHdd5OTsZFjsBCUmlN6adzkwlnLTR74Niwh6KuNENk
pbvjs/FI83ljmHD98wTOZOxkQWKXbpjPedbo4/JZVBPZTT4pnW7G11uVXixeK11BkFDn+v1pc1nt
xMm2rWaSPzxDMq9rKZhB8ADam/zU0boQf4d3c47LB35bk+EeqDJ8CKtA6v234lOZdJuBpIAZ76sU
kdNmBP4DBjcyx360rdzDD7EdvQdH3boBwNXhqvOcKHQ1DZl2BwgC2rBACn7mM4/Kp+mx5j49H3AO
/ZExy9IpkqVehYDVgKTCPHGQIbP9bjfJMBa39c93LSPAVzezctx3w8OynPzlxBE/eg1Cy4Cs6V/C
P/klqG5AjH+BtrZEqNTX8/BUaM+x7n9KiVzgZ1XlgCE2tqR5r6f7ue9xhZkP23pLbrhC6qc+X7qm
M0oZzUHKecd6XjdXXcEAwDBGqqZS+oD6maAecfrQxTCNPLgzRlipQb+LIjrWfixPuaPkQAriiVNA
8urEs+m8/gmx+Hf8hSkVQcu8I0z/eF1J9DUYQU/ehs3RAasq+bvxhB6dSC6BIWeqGAHyb17I2BEr
otuZ9J6Gl8R31MJcPXNvHQrQ8Kyvl2bDk7gl912RCu7tTWas7wYt2N2qCKsbuUSQlTaOmTmhudGN
7mMs0g2bOuk6GvYW1nRkO1k6TwII7em1f8XT05TjG+oSLaBEjy+G1kx3xp7WWbrZsvQ3xnwRFGUa
Wsk+c1Pwx8IM0+/RVKp4HsL2KCR5APJz88l6evzncCu3d9J5dkMpCdX66/jyam0lPchf7AnspxDK
VRXtVzlPjjNeQcowfLIy/s3vMcCxKfiMV1KGF24iE168oYpuiHMqJwn1O+WwDVNkL0q/lRDDgYM9
/KJfqvM84UK9M0kVht3zcIY94zoHeoEfUfsH6MffzwbutI24zWGpadrz+Hywdo1+FAU9ErJpNp1Y
TXsdzw0ZYlytq57VkMb5AUtbV7De2oivxj1+WjFBH+Xu136fNind4X4O2pj5QEsCh8ULqkSESQ/U
Fj2YvTV2SBKFaWeL/GNteqKOv7g0cNDxbFwKd/0qv/sQK9XrO74WEO+EELRK5iQ/K4/c3m1cleQz
NyoT0DuWAKMVrPt4RRtfMMPiCChDEgyzIys0hJcyD+MJ2qN1dfJ0Hz/TbUENPrRG9ub0XBSDaNuV
UgATKEZpArrwuGYdX7wz5VSLti8PTBL7e/aJCp0D5sVNe05qluk11t72yQvi8w/5AVAowHbSkPkG
kuFMn5psjnWNcyCSgVQ05VaN95auJhYgt+VQJtNFeffApF7UxyrJaiErOr7Wme19zt5gC5I5G+BB
DZDvTraR409Sts20w2zUtog8gKHQxsVVGh7uYo3FpJevS8wkAC36eDkGFc8Uzu21R68CqkEq+3Dt
hdBElei28OkxB9L4pRw5aaQoB+fAQPdaWPJtDaO0sXIM8TpCW6112y5pkIv7TIpbeMUopXhGh9kj
as174DTb6AiJtJFfR9ycL8gTzjeCHI4W+HjAvBhbhspEHUtKizPNi2cMIcMz5jSDddaqO+f3aIw6
xiV+mRll/m2IGw/rxG8jXsHfwHjByq/2p64xIFFUVNvPeDkGEC0L93M4xJ6UGpHtha4oO+ZF1NGY
F2aHGgHIb6KHD1AQ2OAtjA2NQvRERKsU9YkkmXCuYUea24po7V44AYLbyGqBJg3wMD7WLi1T6Xvi
TOToY0ZJwW8X02UUHfTGBQrzlt4s8SVCKRJLSWVvycxdKuLtb4HurdS3Zq+/XZCberj3x77ZB0/e
0w5zNTZtyNT2VH+eSRm/HE+VVUtpdpb5lAbE4fSxegJrGEv8cKJDhHn2m7INfOAFncnimgjtNsOe
vJo4OFZI46EgmO2ePIsUJLzQRsQjDZgLJzJLQOl6wvgg0U37gekDp40/I2TpSyrw9IBul7cA/Bg4
+M27lJ+8r++ac5lphDX9JrwQyMiMYwCMJG9La04b6xlefk2yRb+2Hx8WP7meUTrYCXRJzdo4b3nh
RG03FLUGk3LjeaCBAnitpq/0HB89oJN5Z0O+DFNrOc0AVaLMRKNb6LWRQx49hWHTaQD/6JxFzQgI
imr6/aqIspdJUF+UzPdTe1xJ3OHMoQzVlzMpi3Jl+rMOfxPA0cE2sBHj6jLjl/UNonBCGwLBEZGL
gu00mzBMssgDSrwv4A7lbWINKNSF9PRZmhjwjyDm6taUM80XTTEa6yHLzZNZxEzqZsxgjPaMJm9E
sx/nnIM1OdP7HEPU1SgJHalLS3c9eqk22Pg0/WZpXnzAspRaku8+Iai5CmvpTJGodtbJ7yiiHokn
UJ+bBT/nBKHsjBH4L3gzCpZkizGzijKBd1UO746qXns7so4rzJm8of6QGzw4CCcNM7MyyqTyk1hv
7zDY+fsLJjoQESjL3a4NCAMxzA0yC/iKcf4C2iTfMypwv+VCCqow6Z6asibdPlCuxwxsVwBja48k
6EMIUZHmQ82iivkOaoQZPtUVLWB3swXk2BmT6qBvybtr3ewfm8Q5eOC7OaXncmxLnuX3y0LlA2gm
afLdhOj9EbFiX7+GduwFrPze4XYlc/pm9FJywxkwVZCWLPyZg4SDR7AjBEjdS3WB1CDeBuLdEic1
1o2aw/PqGwmVkxGeD0Dopxzx1DELj4IdVjCDqNI3AMBgNZ6cqzg30T7gXZqE9MIsX86nsmrR47Tb
OJccV3fbzXNKMxk/9xGKaZ0CgHirLsjd/s0aetX4r1elzvQB3W1IHjPZJUMKPjhgNcmhEWv3XulG
zkkbQEejigUZET86HsVujCcHPDx5ELhQa/QrI2E5yeCQ9bHf+Cq9rdLuA2X76HyIGpnfz0fqiUyk
66seA3qvIKl0vfMqrYnyWOJ55595ZWRczw7ToBF7H1RQwaT8nu9rPdLx92CTUEFAMjPBZ8uP6p2P
5jcowUboHMCjDuN4cflsaUzYyle73uXENBGdhbIKUNBq7ZhUAe4QkfjcSb3x3qoYkf1ObuJ+MOBO
nP91hJGwIEHXy4jsWvHxasAfRsFhJ2CF5AxCY1ma+GcYy2hSP7ROBkxREtHzv5c6jrPdHD7dSYNz
VTrpu37+L+sC3ADXnKxa5FBAoeC299TZ0s5V9lOOTVwiUWdPzp/U/xupT57OsDL3lbQCwyzlNiTm
QrP0zzFHiaQ6yP7OI0DqA3J2mxYpiMYVXoaEif/P6aISdxFWI6kPQhi9euiq0a6vvHMJpTBvX5Yt
15Y1KVkuNmdz9i+Vz+m8uZk5QmB5z5HsVRJ4dv736nBnuIcw7h0S4+n6tf/Xn4+ZZAaPgJG8UTID
NG8Nq+5cFahjxB+gBHLVBRKowVG5P7ilHqNVtZZkwMmL/FsTiqbswDnAA8q7Tn57503/SQ8vlH/Z
vEjTRl2EktVizmd9KEZnwQqVKzUaSBI8a9AHJAYYZ2fg/SGiR5mgoDJJnXbAx6Mm25e59UjO5ayP
gwE2GsL7TAtbdxX8uw6Q6SnK3qc7glBMfAPBL0B4NrbXBCZ5nFu8R9vcncE8VjWjaQDnWiNeBtGR
2a9hnFbX07ry37V7cTHnopBt41TX4kjB2iUHiXmluTUJDgHyNUePE0ltJfADeLtsmikXbsIwq1OY
ZuhewYfC8wVn2eFu5AftPqiTxhtmx/XnofereRK4CFcn0OCPBoT7PMz+9lN2LyjJYjaK2EqB69K7
7vAZaU+ybaAKaOd1L/5Sgmn+rXSV0T85xyCkz/qiGr0ve/gsK9pChNeptKy90Xzm/CPfiscOyD+n
Kf6iqsY1BoZWBNLMQB4u23pLNDuI7ioPCWmF4UTk9PwLMxMnJ2narH68AGVq4vbWKKQeO14sCOZR
pskcRZwir0myOwNQ2palLQs/7Jmn8vD6e2vIEMENhoFAJItHvGEnyu7PumMw1a7XfZFGcZPF6EYD
VPg+smz+Mo/vZGbgs7XcL9qJqIgLXr2mWA/QXtYeSPEMJshlesWmrewjw9Fe+JUlJipV41/+s2tW
ntaqD5PjQ8jB1GsCOYV/gyE4vM0eAZXwJ0k+M2sY5bXsVpFZaEPJIA3mVJz20zWXauIoARnYlZzU
XZWff4hNN6rfp7ecy7qpKMvKwazJGpeGsQckw1MGWGhh9rh683gR0SXRP0SyXbO3YRSbVa1rOqYp
yRstpYvGWEAXChBTaOeTlmajbkDuWEFvLSukR/BWHG+FvZFy1sJgy9al0Gr0N4XsIM/cioesPDe5
yR45tn5EdWCiA05WdKxncZu14lPli0T5DEwa6lwYKrHx8D4xIJvYJbFC0LCymc5DgLDvkuFgIUhq
x3nxSUKsz3Y6muezqFTg7jm2HjOejHSlWWJ3KYOQOqGmWPb/xlW9aphx1TL7C2Pl2XptbWf7hPgk
5hiD6tsIfyVliBrCecoQpRKnxXVPEAuSdRiaLx+BP2DKtzJAfnd9qa3LTUQnCSR7CbKWZX00XLQP
YspHYg2ozXzFKyIBfntox8EQEjCuUE8eW5dtQoWVRPasLBRPViJKkSy/SHaeUt0/VoILe3jmmA+V
GKz0JiiZ1KfL9/pwrCcJ/YyaOiVzzbDcZvn69alGzHVXtp8XhaReKofy3WfOyke/eUx8gT/WrTr/
CRrdAPOIzU33qRRhZR7C7FQjKuRcOjQIpLOkswMQraAPZnim8p5ia4klad0A8bS8bsk7dz44zT2J
6aIS0jr3eMhalGkBwlHw8iP9CImEz4+z6HPUqRWeCE4JZ7lSJBbZ5TV7hYKA+SvEhf0ri3q16Rjv
qLRLV+qoLdK9Ti/s2NLf/0dA/F/t6/qvt+sZ0agEhOIAfEtAE6VQipHenDQDnQsMnkFyds+SyZ5o
ZCb0mCXzmVbdAYFecJuBHoVBNlWEr4f9uGL8J3M6tcYUfU1336tjKsjptLrYcNCi1668w0ceLVnB
7tNnjJVcs44O5aTDVLcIpl1lrdMhmSXKouQ1m9SmeXTV1D99Sbk0Mt8AlLtpFlGPsv/ruO4qDbbD
lQ237j6/fNqeteRyZ+AspqS22SW9Qqc3GI9V66BkdNOfJcOKk5fX8e1tLaIf+tuvf65vFyn4pl0c
u9GkkMJkoPKdKB3ebCCK+rY9/X6FYI3Gjpm+XbziS7ypoJDJZo4FhNXUq1m8brfCGvmkRIrjQfEM
GECmjb+UXynas7X9/7SB3b7Mc4IRE3Q0XqNpuJtQasjgH2V1Hud84G03l0P3Ys53cVtKLqc44S7P
6DTD+REZronAlCTruaeaI1X+wi1z3wzMP2olYlZeh8xbSf6i6L3nRzILeaBnJofAnM4ejs0DbmZ9
d+GFBe9yJk0zjYu3wfvR1eNguYCl29fCzJvG2gOq+M63/hr0T6MSMf2CLb0Hw22AyAmPTPz7oOwF
k5NT/X/tFUb3pIiFSReohDSCz59p3jxMhKWLzsy8mmPHki4xUUDs/b9phkThsZPpkk0PNH30+RKx
Q0SHaNrx3nph7bROFgIhJ0L9HmRevAFM2WrFcXvEjPMITG2XGoqAWltb7vHM1OFoyd7z6j2peDAQ
gbdZUB/Zst6L/K/3gz48BBZjZpbHYb8jzszsrxcab2qTXyBMK1Hvm6LPSg2QtdoE/+8aBbu2tjHl
NadgHwAos3LQTr28xDnf7FxXiUlmgYjN/sT7sadgwKDAgzDGXeBImc/9lYZAV0LSEmfxbna43o2T
mmv2ylIwlVcg82m0KLKtpHZcrQhdidpxu2tte6yIm3B0imaiClIm0lf35N97P+iaJ8/7YRXqeZV+
n8fE4WBbWCOXyXYnU4D2YjtJ+M73WKeXLpq6B0f8zaVvuU7Z4FTJKHlI1B8sAVkh32yowMsEA4mW
DQu6ssQc1qtcc9hgPaHyZG3Qt8QZ2L6x/uB/anFpqVGHPOPzqZ5W+NThKuPl4BeSKYCmun20YrFo
2b2sHy2hmlaNDCL+FKNo+6JaP3EplqpYnnBsG9S2pStdeM8DZD866FkrTqNkwUIZ8k5Tzx9U1+oC
XiRARHYK3UjYmkoB+qv8KqqbeS2Sq8rFqgbai5PUbCQPAhlOZPx0R4B2vzSky9UC/JGWg/ruClMG
AJ5PtwImRifXU7wP2d1paab57hdzPVLo/HFk2drWLvq8vf4EITFZxtEosalu9Hb/fg7z5jYSnqqK
pe68+QBnM5KhlMtrFqGTdSTA1Br1XoXaPeuvlj9/zUkEtAdiscbuc0NVoO46vo/lgCqvUM0prLv3
osTa7OGVx9DAqkgJ8riymAbt4W1UabzyK77B1Va8Ka8JiHQhdA2Q/gBPl0GPlASz4Hk637LPjQPn
1XGoaXSfxp/bLZ4KGvk8umHJljg0T/OUQKDWHmm6JwAPKDytiRYHLYmOggagN7+uRJI1XGCGxZRe
7Ktq/vQpVGGM9jEbhmiTqhRWoI/mmjS3p2VPwbcqUzSgdZ9zbbBlu60RpwJ146ho43HdVEIrhrSD
Jitv1h7BWK1xd+JZu6Jx7BT4pVgRN3V9ZhdPeDxhYMhtYm3neFbDnnkZQ0U+XgPSn7yrreEDesh2
6Z3Ay5LCK+AdmQ6uXRlFrfLYVSgqDb86t/ZP3KDNQ5+l6JFSw1oLLeKEKn7X085/S0jSB4DxT5Ed
W/a+ccvX39Y7h2JR8ae/yq+NAvuWdNkl5v+BVomMyiZ6StYRBDWJAkcw1KrdDJbWDpiW+VYqI0ls
3ABAT/D/4Q7Wckodx6UxUfRIJdEPQ34yWPAZFK8EEgsjiKN1oZh6spdN8S03HPX/pDj7AU0i7yLy
QtLWK4+J5B6mZKhxQUSZPXq9PQt7kpP8Dalh51cKIUhqnN6fwDWz9wae+vwjzefzy2B0z4nfZBtV
QAu4OLB4kC1C6qHb1DecrZeCYx3Z+qAMJ5LisVwuWs3ZUJ3V+LV2v/8k2jg2D+VBOmzKZXHdX95e
USToZnLajKZSxWjLaJtgSp3pJde5A82ouB8Li/cuGlzQGsKvSQ3kq/VBHRpMqkwgohEU0LDQkXJ4
zcOSjLjpnXFDiKNRmkhSWfxBQ19xxgpbyAh2Ry/6xDpZIlzkVTCmAuaUOhPJS/tzo+s0anyz3NIC
PXnohhSI1r8pVApSQs6uQt88l7azlxsPvN3Al1Ch25T6jKlsTYROMeVBbYmwe1tkfGbTo62FhLuU
inmRhrReJWS98rQ6ingHf4/9RZRISvYbPPIjhLpb/gugJIEVVwForXX08WZQrjHxCIITFOmZiaNc
JmKy7D1bQv22QZ2e1j3+7AnDuw4G+t6adpcxg1Fyq1YriBUd7JoLSma0nXn5b8gKyPYowogEMLT5
8rnCYAGdep9u7kJYrCt2C4HdgB7R9/4SAJpNkLA1RdkHelSayArqiP/72HUUFAle67xbjTtJqMob
hv1r8CVWY9sMIRpKi32YS3qiee4rqphkGxfC4tkTW10VF77ZLZY4jEgq3OKTR0wZG7DVWV23gI4s
8mxW1a4iNwEqsSj/DU8MEerk90CkQE+tZiqiwf8B9dxAgE1v7tcceuyXKT6E8yfA5nyq6ddk1/EV
AmH8lidHeS0DFRlS47LIj3Orop5As2ZUFafKLchr4VizDiL2Tcb9O1BRP+VApxbhNTBKdIGcxsUq
uU48MyMAGd3XgZ3w30wBDlPH2cH3hSkjHbpvHWOKbaRGf72vhcdAGbXuhRMdIItrpb5WF22Hf28t
y6wFxe+Qx2QHX3yK8LUmNP050mDaDEA4HIFFHMoiMhU5rkQd/m87cA7r6RbVyrTGp9LInZE+mjzG
Tt8YoTrNTLCd0npjLZmnbKqJIYk6op0joaJuFNEqr4BLPUjfNxeeGaAslCTElUAzqg4EKufXEjnX
iBkLudkNTWFW9vpwwq/R/BrFhZ6uUcpz+XIuC61YywpTLtmXkP+YQx7gwfCcN+z+q32PPlUMsSUv
Ppaa6rtKpIbIxpqVMriTshalgCn+ovhQiQKt7WugckhPrVZgErvvsoSHmmpTkSKz4aE0BPSMfSRs
ZF/rSctKqTbjoBcOdA+JAuQl9d0ihogYkstdhSgN+sBuDOE3K3d+trILiVaNaUUEBEG0SRTwbgLv
38aYesO9k4rGduPWG64afo9iZ9cXm+RU1tModmCsqWCSBrs5qeXE4uGwNUR0vb0Z+wb2qFuXeTsI
6iYusl764h0jbFYQwM21r1BmDUbF5peojpjcUbAZBlMiFoNB6ovg/5El434Ds4U21isiB/skhOW/
DjZp66cbcaMNuLtx3mvO+CivP3tDQOcFLloAPcLZiFLCOAKZ4YKxrqtKmIPd+607jdHhqGGnA4Vv
RobdFzXlAJ8orYElqdsrDtVK3h9qb+8qAAjwKqp01NrO82E0hY/0xMhQgrMNuzb3KMWggAlsmWBF
vUF7la90NgJAkQC8T/szWdo1ZzvxQzwXJ3+H/Dsd67pYsh2rZ25y18/sbCNkwYuxqBmR/YwCQFvt
9rroqrWgEq4vdA/8luEdOOE+XPYdYXQrlSpT/WQaohewibm5qjwVrTzV+WXmsjvii9uAFwZzureA
eUjdG7rysNvIRfyvY4VzfqbK/V+Va09wGWgt1aiYsb5231ISbaM47biILkSrufFn/t5lZZ57uw7d
X4qReltqkzMY0zr7dxsXeakC3Ql7gnOnNP01lxwJNX4LcQbmXR13mGr5BUYC1PFRLy8zjsVHAEgT
tK4zU75gUodGQUneeFBQeVBKYlcT8YR7pYknPeckFhbPtQJBSNisHUbG93Z06QAduj2ltQTAhnW2
F1209boZhD8Rm1YdTdzx3z4FxK8gafhDPUgUxGm9zUCv/R+Na/zOTfNE5d218Ln3Mlo2fgx0h1mz
rqgZNQiVUy8xp0r9IzAegLW+Jn7sSwmJ64WK6ADYwlaOOpLndo681IAQ9QPwCU01lg7fQyWUN0cU
JG5UqRrqcdM3BPdeSuBs6jWo+76CdyysxPV7nVHveCUqwmuPWK3+Syu7JtkfjpJ901V8d+j0fmD5
nK4FXJjQ+78RC1A0lGTRsKiKxJl5B9aA0SXdSLiSTQdWNn2ieXzTC/qI/4xh5BLhuCQUaqIA3F4s
5YQMxNcbD9FzcyIsdSxjzYeTcPwMev/EnEXk9DM0HQJmPZAgg476RojZ6X72qJWe8tJm5gxdK3l7
hxx+FyTyYobYLLlJaMm2Zjeb03X6061pexWQ7tTi8mcJsyH/Fn0ATSL1wG3hxcASI8GQZtZ4ERUx
0qtJ+0QFN9IX4h4YRBxwgepNkMSxU9LHqYZst5LoFtmHdGu5ot/9KCxpEHYC8/1pipZwazfP35QK
aWT+KlGjhih2tvpIEva03X6IkNXw6TC6A/v7yfo/ho6q2mjiKVhKW+/tv9d68WJNXXlX9SZbM1P7
Sor+VWPkJo6oGk9W7yz9HUnzhxO26HgZPpWjMhrVSaqW/cKBTnsEaskJ8GU9BXTFVwPH7XA2YN0i
YxVy3Du0pQ1OEH0Soc29mDhKcnSBLn335EJnSTW7e4v9YLNai3CnLh3OYhCDXCn2EaLoRRH7odh2
c3Lf75stQ8RMCJQLHcIwjH2WQoDNOu10kXrRru6CuEXbgxwsj4ZSQvaczPE4QYxo8Px/ScPZVj2L
3SFXtJgGzEYrfYTq7XcNtTMlzMJ75hV3mlqrBB8Q1mcbCBo3kVJbYGhytrXJ7TTjVYJGxbREKgrK
0+XT42UxkeBFjkvdNk+H1CLAL3zjXYQd0fM3fHOwtG4vq86zaNV65ZwsTA6hQisyyE9ZkuixApo+
xsb18dHxVpI+SC+wzCQ6sIvP74w+mrGd52noqqIur1VAHKVJhFQPhTD5e0NtkERCNesQ11qKGlvN
tEzylIpzIUv6EPRp60i2kBtBhFaVKvjDKY79tIeM4YKcatYcdGyCzJG+rUJnBN3MnwHt59Ss5LkQ
kTeOuoAsu8QSXySW1YXysakiebVVWmV4GOocQ8kP1PR/Spc6OO95u9k9dVVv4Wriya4HsRUvuUQY
FqlqeGR0MyZB73mByQWRiE/d+VK5rmbu1ZLqD0p06iPr37GQyEULBJHz0UGCdUD3Dsr7obQyF4d/
DmO3mtj3RhS9ReLp+8ay86PbNWJ8TPrHaB9jrmhQtzd7ceWD1uyyLheikBq6jjEyxjVMxMwfXAJS
bpNRU4GNEiRFg2WM+Ueo8o2kvTGwsR1cGhUjZvtdhOLngEYN3cVr40feh6xLL85iXY0fMXm7V7Op
/kVUspXleXC1qGDSFc7l5ZpOw7MUEje4OGefk73DbAju+lvmHC9jSKmxZ0jOXFYOjVQJdKr0vIap
sl54l8exENhVz4hKwINuVz1Qoq71lft00MXsNaINeGHNT3EkuZ2rPccg/52bYrBYw4toAVJtWEq+
9zR2TvA288mDC8iLzebwJ9Nu1FU77DjjXf0eDKCn/Ih2Zo8E3HvtnCn8artpQ16Poy4qSku2OiJY
v3WJVBzGqHd4u8tGLKwE4Mba3qej7ENcYroqhm60MKY9M2IfXgvla+zLM3UtMUJxF6HHiQByxEMX
tNdjyVnDmuNKC+igoPlqv/xfJpeCA/S27diIO9gVVeeQB3Arhwf/bWKr4igNKkVvh5GvV2uIOmDg
+Y0DsSgfICgCns84VUhQkjmCcZIXJLfUILFVxIzAuHA6R8XsyGCMC6M38fKDsp1yS6jydFbXVz5l
gnuIY9oNdycLfV4NtCx5usS7mWAdpPdJEbh5LwESy/heJlXxCcN16NJCdGAoJcLn4IK6i51V7Qxc
+HV4wV3uDI7S2B12O4Eh6HdHCxbZ7p3LzdRcwjrN2thAaPK/0LkHCVUHSlcu1uJgT31gd290/WQE
u+jeXWVltKMDp6yOnmXB8vqQxm8vyPIhbFX6IP1VzSfLidpidl90W9DxZJV6NSgenjCqCFBrv7zC
sEqsQi6JTiAY/2K7FvwydbK6uC6pCn6b6VKxhVpMeRIco2OFe0uQBBzGO7VJxvxru0D0ofGw/H8W
oE+H16W8TxVFHJbVPVXLRmWpWHaELjnafOAZ7C/9BzrT9gTTfmU75G6Ma0Jvw3enPc0mWQxDisCn
F+tYRbZxTM3ZC/w8OScrUYbRGaVSu07fqd6p7idptDGk+2tB6gtgmi9byICp3+Yqng2Q8KJH/QSe
nCiF0usPYaACmQFDUcCfd1mLxVmarvN6dtshvHfAvlD4lj8eea7VoZEia7tUfqPjNJiRErbheBbP
twaw2Cj/ay9rRhSsYnfQfMNgIRWTejdSb5+W4ZavwxDDglIuPBc9W4oepCdMTrtNJAWZK6omrvIO
jn3repwiLyiLYlyhbgNQmpJr/F5Odt+4by3tHjxhQsKo/CUJhfnPKZGad2gbOgZRF33G/vEkf5eq
YDtOi+XDag356SerEMhdjW7fyzriM5dYhnR4iZry/3lz2TJW2cJSEfZ9uS2o7mqqWnKnxWbQ+mAv
SLVNNGdJd8bi7Tvv1ORp0lVj/Jv48/8SqkuUzehbblt+xLd1ykpueNoCJ4SZWQjV5sXPzS/OKYkJ
vaK0kJ5XLmk3pxo+EWZSEXsRbqdeqIXbqklnEF+Owyn4IvnlKkg/b7GBTizfupC5gHe7oHlkeb3z
RCu37zrGDAD5tqhOmjRfPTQ3LEhP1QMyN9NqsfN8ZsTrGV9udMOJtsXustNE7UJYN21BNw7bTU0X
9k+7XLbf9PgH1JRfDkN48NQLKfETriSN8ANvbh9l11fjHLLxoH+xut11aEI2YR4fOyOtJJKoP0YR
f+XZMh4vU1DtZjUk8bBlaFyPzGNMVp24HQheALJVzrxo3J+YfasVMR5Nodlu6Op2oftM9Kp3YEwG
vHQmM4KM4KzC0usFJ+OjCMCOJopIe1AV9jcb+86wnwydDbxHbMHUJL4D4cKwu7r9eP85DLJnFeEC
s9Qcnzn1L2UY5rDthISda3QEbBWF8soiQ1ZZD8XBo73DH+BZbMG+WuPS8LQm0JCQRxcdRrqVZ949
Cac4C5tt2ELvNncMjZ4IarNMph55qzcwXCmYvPlO7ZxCaSapawFcXJb2wtpasbADikY/BkIKBYj8
gRyyZwahWV7ZXdjZGnwAvF6EyhYqAqC/n2SxhNtb4+WRT6Vk0h7brMnqPy2AneA3a/Rvdh2nw6Ia
7R8CpFKrUHBhtWEV6p/Dt3k68Kvd/LR4Yu9esWWjgM2oKn6YfYsU/cCfn3Ez6LAWUPTGaortJeqr
koOLN8kM+AkqbTRo+HClm2mQG+GZpfdUwo+PHy4jdY/6dtgspas5IBks5CtCvFqRBSh/c+Bmp5iB
pbvBMPyoEMVZIBpa2EfukDYLZ1GXCUrzPhl7IUNhO/otaQB6x1sAxXinEmzS7/C5jLSTJjytAfIW
AlBL0Wxgrng5vqO9E8DNjCPArYXZ6REg5Wh5IZt4vumArt+95y4TWNxR+afobo/sNshwfqzf2pL9
xYdJwcwRnbx2dRlxf/3WU63XTjZsM5Yq6mbRe0MzPvJjbAikOudQe+pMAN7tVfjRdXLf/71kAMmx
HPy+3C+sRX+9crTGscBlBdfNxwyss3qF1aE1kBSVHzFPByxcWlvMwoQl6rwVsE5n7jdMYd2fVpMD
B/cXbcQyExzGJOa6FSgxasfLaIWHrPFrXVlrNeGCtxqhP62cpTi3/012s1+/gNsJZdD5dYo+pfPe
UT5ayq4cYwwd3gNh+gRc0iyLktnFDI+EQNNJ2wg2ARe57XDq3JTw1PaYoCjvbxDZ47w9rH7gFlHP
XuVyk5nE/KZjW9ghdd1MLRhA088eLifGWmybFPiCB3KOEWlU6BLR65Dy7Chr0yXWmAT8kQSuqivK
83coX83+e43Q/uiovBT3V/qTbGXND4aYF4le0/EcAnWcdaCAE/IR+LL4Nt1Ij2KfeBAR8gAoqDRa
qRImipITsLvCRQ9KPM7LZCPuVGLWIFDzYqeYfdGt7VtKHnlXbZwaDo2tE02MhE8FseqQ2CqPiFvz
HH/fGG7+nyzl85GEDoQY9cUm1B7unOwwPF6rxrQf1aPYC6MxVhLMbgppPeUFW46NuvwwQw46sB0/
CtFCI8wPBgmi7Rrb2JD8sC6VtG6P0eeHwAskoBH/2pFFDsi143Y7J6XYRVQXKAPMKMH2ZuR4VEkB
eXlXJCUFZhINUok59/t4VtB8oRuMkr0hedrNCLxamUUSxfo4tNjNKeqEaj/ukDSFQtIZ++eZHBem
xyCVttNLNenWd11rEp4xRpudxiOyf7KxbbOvg+mCO6yAOQQ/WbT+gHsvkQJTxeiGPdWkniyHZk0u
vDdK3iXO3oCmLtLHQmNWnHziloWL+ONxWDwjFIv50fwQMq128xGez+RoU9ABcHeAlu+VD9O/eowM
55VAx7xayTBD1/LbrOWdnyJqCFUHHUkZYcOIw8OIluXSywl2Kde38HPyRv9nm34Gjvj2L37qAl2Q
IowZsI+UCdHFFSHjwKoT23YlOFwY1lEAICaOTx0/zK97unrNrEyTPLW/di6aptLiImRNRaZxmSZ7
uZz903u6zZGS1vu/1IKF4fj4UAO7sWYmnTp7In0L23edIs14gfASO4gHo2YkfbUwpaddiKaUUdis
NQEL1RXPnt1heRZ0VLynQeM76SnyqMGGpoXy4tNjC0UqymZN8wCigItHJnP7SlHVuWUQFnHWc4JR
fSKdNcVWJwLmcZFSdm4lL/ETF86iPUg5C+y14U9qw4R+cEfoyqW7z6cquqA2jk2cNbe1otP9zZt2
U5R/WPeC/8SrRptvYPhkkvh4OUw7Q0f3cjaF3ibZ8JI7Be5OUydUcJ1H0ObqLrSRcorvjNV2A7T2
bYoh+LOzORAs2AgPRBndAleoAL9zK+rMfhC3iO/Zixl+/sYx4miKflLoVIz72PNlDpwyY9X2MNKa
80kPMpR0W8hH+3vZpXj4idHej4KIWPsEct99hjSsulZTXLYqmhbZcEYdYsPc5dytvMyPDp3kgcxD
ov5FHwwqdxwpDOF9EInaQK5A8BHpQagVAW8fMbvqef7Lq//LY+KZlG8x/ohEazvbZru4lj5ViZSl
Ktx8YJ9J2SICrGnZYOD2LaLgnNHc7IzP4wdPD0Dg7mV1Lz0chjHXMxAF+5AGB8x8aothtjWVpLHO
DGtiR8z8B/Ftq1wIl7puh7it1e4i/7vAQ3NTXPUY7nO4faZwPGG8/Co0JsFSFBPG7aHO8UY9y8Xj
gG0gr7hPpAHtU0/c78zm3a2ojWFjXkMqQGGlGdiJrM7MDOlIAKbjgP2ZUK1vN9yzEdFYTG9J65xs
akckkwpNcGRumIO3Qncr+E/Xyg/kxoTIuKQCyjooco83xEOjgIFK2cW5aw72jzG2iLD1jhOea+xC
+xSnhcJWB5jGgiMRTqNLBqg0bfOoulisjkxOQPQfJG1dRe6Hyw9pDqBCWRleI4vY5sg6K9O828GT
nwavKZvh8qZJCc88PdEQUKIPkD1ZKvGnrD7Z23uFkk1eo6DzO6fi8M2RFQqNK5wn7XyHadXYDkvp
FVN/J/eySL8GsNvQUSH5AMbzVS45OVps8i2xh7VKQV+rwAytqxR1Izkq/A82AgPJQKYXEvaKQeUR
wFCc/o0g/1yI7TQGX27OgZ8uHTYOSsYGrq3DVPVWj3Cf4+bFcpmHwa7Ab+ovvpyHxusAZfpW1RO7
WMcj8DPmLJVzBHFEkouiwu92hraE9pIEGAfHwjtP+yF0pqApOK0TWiBPJ2VpTS9s8jduhpLU+ket
jp4Pc53ANSsjrtLyyqZNqkQYlwSCAQB/ZZg/dnnZ1x6UvcZc78Ma0WjzQHmPZlaEVgAadS8MpH+a
j03GEVk1Q6MWZ9u2HXxmjp1qHwmSZASlPx5igzdueTS9I65n03UQZ4KP/2xY3Tx8mBk7jk7Oxn7l
Jdaml5w4N98rz+9vTWN2dYHyGmvQ9vJRWS8MdOfAVMet0rLesfq5WFVMjpy8yOdxQs+Xubv/rprJ
CKDz9jyRnT1WcAyf8cD5b8lmcz2qKc1nHwqaGNSrJ9OUGH9EIIfSUgzi2xm4sUhaNzMcG/Ymk3ru
tO12HOXCXKYkLC6bolWrJ1R7yafG22uXaZcQ9TvkuRQtuB6XR0XMVcNXOTyi+9y0msARe6Qc7Vc2
QaWDf3WBWytlg+b8ilYbAQcktKZ6Vxq4IDead+Ot8J742oOdnSxEJrQvFwuARJPboyRCVuwRzUbs
d9zMdxbE7snlZFb9FynmN2VRb6bwQxHb+I1RG6ShjJpoEbG/bxBez7tdXYpCX2xd/qB458YZJBbW
2mnms3V7WA7l4C38DeANA7qI6l/z9W/JI6ya3ezaSwn9zdU/IDOB51imEjptVoYGTUyjzynD8H0d
TcvrMmaNvjZwA1XzH1z2xwVnKzMdxwL/7NMe59LuVkG0kbN1FTdKt4ZEi6fWBNYbhurHV0SRnvgM
NqutYWMhiEr0GFvtj0Yo7RX9ujPbfnT7NzZPoD34yOSKH5lfsWsn4IOUbGZ953fLjCj+R0WFukas
ZIHs7WnJva52Lmsq7PLqLJlzhVKcBjSdEMdY8PDNRdYTE2Jyv/N1BL5uSfBKf3WhmcjzvP7U0ttw
D3mIhummTbZYfZ4cDYklwv/OGB3mEkp2r894MFRIyLa/BH+mFg9Y95W0ZGuCu8SNmQOXDlaMD6/c
460AG/JyNv5+0ns8diD5E7LrxT42bWOBwCHsqqlIvmeVeAnyvObsbZLRwNBKj8RAyQ8Qie02tuyL
FuwvR7KuN73UvCEaMNeItvkCOhg2Uxl58DCBKLgiS1ed+q8MSG5BoICFfa23kgdl4lZJfkOWlx0p
PEfrBAxJ4FLo7sV2yN8i8CNHxXcoQcqtIvO8zHXomrAd2cDljjlypbJ39h5mtfi3esgv0slRJ+9e
C9loDz8iZfl89R9Pq0f1h1/GSvoOO3b8Cr3lOVV+8ZBUR5ZLjbyerZQahX+XCU702XAvd7IbgRF5
NjNsJaNXsyc40AV1A2Vla4YHa0txGXCa1ONat6thIznNGA6EYz+Q5bER7ba7delV9Wpf8roGm51H
dqdBBIe/fDmCYYNQdB0koB+1MvM6xqYQSQuKJCMZhGfcxpoN98XzgDbZ+8sh1v1BKO2Pr1YUeyT1
PLwdBXDoiaESR/fa40DTRoRUjis9KWUH8XB6T4qaTh9Qh7L/XzcH/UcMxEJoKjEHkD6tr7gBrORh
mrT3i9ewBOeKRUdO5V2ZMmuG3OtZ2i+TaIObqCSRA4xz9Jd5tVWOoX29x/lynRtvvS+FjFiQYNmW
8HD9FJbXS5qsn2QGlbt89O+mQu3P/lWiBEPiwkVOEfKxGCRo3dgxpNxhT4M3mdwXMI0J2b/kQWYU
T2zl6QdFn3RSP9PCh++f7+6oz594L+I6kA3VsB/OHsWQ9J09dWLjRqrL42hmfkATaQv3xXq7fiSM
NW/GpfeRnrnpZe8dHV04eJr/ZFy5WExLueuyTy3d2Meh55Ys1bk/nV9VkQBzrmjTL6AiFm8MFMBh
n/2AnBHmXEsRSLfwAZnw9F7kJ9wkNIYTxsDLonI/yJreTPyeFfL3ziNwQUSRaclTuI50TtaqXYvK
1tgChfLlqVzPWs1XuH7Gkzr9Hs88ZyzD5D68PjbV6mAOQNQLU0JVh2od52vRIG0sUxNXooUVwTvD
RoLEZ3PuuVlJLhzqmPbSFiOEJjCqItAAi0nG3YTHgRV/wvWZ6NCqdGLwPSwb8le1cBkJUalhojcb
BC7syxvXEKmF8f7vMdW74gymrvagX41pxUmYlwccbrDj1HNr8Cw+jlJvRosbF/frbirqW5ei2rsB
BqqqItf9F/u6i2GxZJB2hSmf/UksAAyuACW0UMEDzFGhXpf9h2LiUuiYJfEQ988bMG7LsPovxWmg
DDUx+Kj6Gb8S+DTS9qO9uurowRnGfuVrAG+ax4x8JiybARu9cfiYvkgre5KFy4kZLy1EOovAb1lS
YDKtrhQae1ukRRwYLt9uy8yfzka6k62dKEzeSXuAEaz58QCBWvMO9ysF+uZGzq/eb9kSbeBE1xTY
NNX+WigMwvnTssepaPcOaXtWqlLPN3y5boFjGiGwNufbI9ANafbOE/TaTkuykuIdFzxabGaUpbJE
dzhS9oIJl3xMb99W9C73jh3EGxDmQS3wkWPtayLgKfR/ZuX5GMjZMCZsXlMXP+e5lOtbi+QuijMq
QLCkDStj06nm5vxPMuweIZDC6TFVf2TULQ8LoxQNN7LrK1zjDNp8VUBPl7al3L2ix6ObsvItBgIz
5h0y0lBMYGmvwAJP683rZip/1CaI+UJRsD89dkI4duJFbFKVYBRJULy3fhRr9fWGfJT3XYn+jXnB
kRwhuvrFRexNaKb+h5Zj+6a55M4sKKJYGek5aKSkMIZz3mxmEkG8zy+MOCKNvD4rZqxt0v1iS47a
7Qed9UEMfakghjbC/zUmqvCpVrG/WoZBaMyUEr/sr8ciSm9K+p5ndr/eVLGY6K74xmO2Gny3fNrK
HqUWLTZEuq3yN0SkOv/tgpAOzSVR1GQTYOrx0iG6VCawmJsoIDcunXJMWtB8yvQLMDhsFNYuHTT4
GLW//tVJk/Jof1mUBUHZbVnFeRKJmM1fHEcnPvqusIQ/w5EyrKHi0eU8pT0pzlVj36OvVpumBTvy
FNaRjmV1ai4zknx45eQJlNNYSq1ok7opQcg59C+/1Fgd198j5u10vjGVPI281yBFR9fv1TyTLTwR
jivaGLqFUlswZxavKOOQc7B/GfKHTWCK8xs3qSRZUnSKzjWlo1XMu+RTSmGWzpiCg4zF5QIhnPml
eXS9gxZ31qpuVtVhopn8GwgOFUFayFwaQH+BO+ER+Uin6XptsJj4EAvzzPZMsxQx1WZiCZ3E2ANO
mOYqx5nTacdVbkXnQ4VkyGK30mdWVknvCAKMRql+veBeX0hYQtJBJZjUUznQGJ+/9Ehzy4zrFy3z
IP/52c1TqTAMSHzeZnlKXNgWP0tQQ81GkrXzllCuYb+umTK17TclUbMJ01PDWSVU9tjqu/vxjyjX
n5fIB9GmwYmgQP9/lpaZBL0llQdEutkusN27CCOCtb1RkaxKZucQ5qX7DSfB+qbg+WQNR8lHehCz
mZpmtlNtWBZuzLONFgo4z7INcYT/I7Bh9cLwNOy29aDh3mnueOi+vF2qe0OKv6FTjdIVUgZ6vJb5
Huchnzg15AqKdhiPZmwBxWDTO7rPPUD5ItkAAutKWsS06PhnLVcjh3fs0meSoOsSXAjAhpISmFlf
ctNz83ixqLqh8vM7B1+w9fvNgRu84Mf5Z0xfUndV2/aKYnwhDmwMQ/a0fs/mRSgdEuYd3GymiS+p
OzxBqJ4ETzxsHTsjhmJw6lH+WRgUBaLp5OnlapnA2CCLUhWfkVcf6WUIPIPcqTXcg29C3OidVnSd
niUB9/IMiXel+RrEoTKZbAcl62XYACwLUzcm/aj+dXvEDUusmHH3OmZTBwRcd5fsHoFWgUfhjwyp
mpFUmlyNe94uZU/DVBywH+yjLcYcHRj4pTmGuSZ9ugml0iDCuyw93RvLzImULUNn5/KyjDmRh/Oa
s6pFULG1TPyl1APEjPx0QsXZ3W7RWnNogDHamC5ZSIhZCYO+1DYFUx1iLaW4gr+pVNP7iU5j/R3f
SMNZikpHI8ngY/CN/EpKyKNuzWClTs++AxAI9qm3q/SWMZnazjPxR0WLXDzJWl3A1NpDx/Ek/l61
ir6QnK1W1m0eWAeQ3P9+VkuoOO7h1qTmXo348dbb5xuHCiQM7szB5rRCeOoOrbche92JxZMs700j
FuJq6O1c8y0Nf5p8DJ4L5oS4S20XK9WQ9BMfvLetxU82N7lRS24knmZb0WhDl1rT57g37+RTACsy
1WZn0JHLPoGb/dkF5uDnIeYxCWusiZ4FyYZM2thzSvmvBNyrdSBRtaPGV89wAg7PW6x766ppouct
PieS7KiNoNg0I2y5CMp+BUYPV+vLTizfwFDODBuiwaNbQGHaH4rNsBZEWzj6WJ/g5H7z5M3MFojg
yetJJHfuZlVEbIczX3+ThWXpwxGUjaH6CJEj/fYJ7xddOf2vy8oPJDFEb26XSu6G/kKRrQxNCiaL
M5S8q3/V4HYUF0y4ApynUEIyLZbLgcXq7P9Err2UwiJ40mdQTSR5j9AKfNSLJqSuU3N5cWGvWyCk
rZzZe6KVKHtx0bGGrBJjgomK5a7AOQitAJlsY6+yVnP7hajUHeUFHuFOTxzuDiYqEnz/1+Q3UiJq
3pj6Xl2686MU+mHdqr1FqYLMI5ISwFSE94ob7H+vZBToTecn9Jvr3zkDRzKZw7jBd23KTvAppyn3
LwZlWAB/Vsys/I//YXTj4bNy6zXVR+ivCOT3uzST22p8OODS35bk/l/nUXco30QGYnCTt3oZ5xLZ
o403FePcJ7eDY60DgRwkmZ1wgWUJ6P8pGtmwy3AvRF2qbEK9ucZWMwqb+v7MgZrPV+x/Ko6Fn2B4
9beQYydKcZ8Z4ijZy+SI3dJx22snfiu9dq50zJnZ5R1Du8VShMteJq5WXibsIGSOQIs7BPFijMna
BEXnjvXFLzQqlbG13VB13gqOmt+f5u0rmS4NyaKW9hjradKy7l3QW4CDZa/HYY8nBcJxMjVVpOzJ
N56jwsD7TfG2sBGxHFFya32Peuk8R9hfRpMBm51vFjYZDcWEIbpCBlNSsPENejgQznpuJZm6LK2I
wD1rZXw3NPEW4x0lNBsEyV4ugJC+7Js1daiKbwh5mG9miMiaSYnRMbtKQ1uUAodn9PR3owddedsY
zg+N0yHSatD0t+8hKepz7fJ6YeqXcPmsO7/4mucRNEBBZBNisXaARJTm1II2jf7scRY1vvyBTCd8
kmX+VgmhG5DNDSKLyNXok8ZYdFSwh8YA9WTkPea7FauRSGQMMHUPsY3jw+2QwqN+undtH41mXUd4
8XK6Ftx/lLC0nBvY1VbsUZOvnbEUWKy7R2JXE1Cc6jYy0sctK9lRwR4GT924xB3N3rvlmI7qKQNS
CdDv/NjitMdUl5mnDOhgTrR3sVyJ9tANa8X9Ucu9W6L7e1F6DXPG5T03Iy+s3/2rtHddgmUhvtKF
rSObNGr+2AeJHibdDoUjN4eAkVnV6vqA8Jxm++eY9aapPVHWt3HzDSgJBJ5Atmz0vH8q79aEoouW
4IeC1bOjVLmYA1bAOuVi4iK1vILUvXnQfwTwiVbZ0LzFJpsDzObhK1Wox/6or5aRZRbl61au9cUn
nXDIxVzcpuAA1+Pvv3qFFp2TNMG/XnwP7tJt2Er01AFTk6WOkScohihKbZekEaDl84RKCsiPXCN0
rpcgRTbVIWhD/oT0yspgUExfMuGeEYPTnERJZYIEm+Fxxqg8QGFJ1p+OuxXC2uOHd33vzUy4kxwF
+86y/bLxXiQfHSPVLQlYsiTqi/x039MGdDm4SZom9ZjMRP/+IGMKg/lXEmzgONP6CMmZiH+m3nl8
GSYd3TQ0t3sXidPEf/kMau7+U6lhvtNFmOldoQqwETp471ss4OraNC5taQd3vXh/niidthhU8lCE
kQ9/hCLjASrpw7EPLYI6gGdv1J0q3isRcfKGQUYzILeIEG/i5pnQTx/bx+VS4v8eNRs7+eLrGWvU
DcaqmD3+lSfwUthT2afuU+ez3cfTvs4hGc3/Nk1XTP/lzYo96saFmOD1aeo2YecYvy7J8IIlWtBW
zh/DGZWZeUHksrJY5P5FSAwbogptyfEsJY131g6lmkLnpIX3bH3nyP3JMOKshCjBDH8oW/tlOWGV
hn6ZeV1z8s+fv+CCLeLZBnVUf8/qXXiiMM0JVGD7TFEJKq6cysWtolydKtYzkrO+5MEDkjHOVho+
qm+huXjeqrlcY7SMcxGFzEG6kKlBVStgQDkxK94NAJuyI0wuYAbukvkVNk3K7qUPd9MO6IQWoxgz
EUoc1LuBkL8K1hNYlyjZqBdBY2OKQeYpsXhlc84sO3AJPRzO6kGowq+OHuiaBIqAHg+iHpz21YiT
4TfAVtBbx1vNn0w2HkmCg64bwVDroGRs734s2f+oy//dLmE3+YXeKurXlWWGm1V9fM/NJFmgW9+e
HkIGEVzggukAWV9WznhdlYmPflpidMmqGi9PLcQlv0sMeo71H/ivnawc/sOZsQIYATedFozcyupL
SNUST1QgxELbcEn7qHPiNmml+Bk7DjJ1dvMIstKkvYu37wnjsRH7YLgylnxrfEZiCYVt+XmgHGiY
F/IkbPAga/gFqbFaOZJHIyGI6mTXKO5BvYJiY6MnWALU24ci4LgXiPYMk9mnVY9H+Lt05OWIwLEb
EzieZKHeA/xOOJmZPae+7fXY3/VwEO7LKcXHY/nB5w05pYtGu6lnvOFeEiY3ixJKDNZmHNoSYUoI
CBbwPRfvLby3cj+mmOiYZDznEkFZWcBLFj6cIDN4JvsocxaflKHvkwAyGYs2guGtlhbNkNqosbPl
shE/jdPUwLh/Qx0sDGvH6L2nBvfdXM0XX/J83AQOqypS5s/0RUV6kEGXF0DxKo6SuhDnzcG5IpCB
wMMs1vLuTXgk/wmCKzFHXi/fKFhtgl4P3sr3QGnuanyjL5rwb9xHqOI75e5XFQeAi9cqIezCI+CC
/lyRYUD5ZgTZcbnbYPACXIxwCFNq0wYFwAbPDOFtKeV5TVeYvl7ooVFrlhthDsGc3qo11O1Uvpt8
roVvoDWosF4UyOXWUY3o+A0lDWM4G8UNm4I+DHMiWwLuPOCfjvqbrmHyBUVMI8CmUoKYpswrNX10
D5tzGad5CvfNTbAlgRz8T9uDRZCFoSr0U7h0tp/FugY7Nw9cZ2scuCO3VyoyJnSYyKP18dXeHukf
IOFPetkwf0ibSpBPo5iPCeV7dvSD+0WEgn8LlplIpRdUtgscPzo9LRq+1nVTDYafgC/s7O83CgcH
9ofM3Duwg0I/6q5itUgdiOAJ9t2JEFXPhhCMFjfXAxQ3eJSqBWGf1MXiiYxcFtaWufmUesIzc1nu
muK505Wk05sPNFfiqmc0VGF4ocjE00MJkCVwO9WzhXqqBuUTXKkl3Njk8ZN0czEi7DcjQTK0rjHU
vjqdW676ryEnrUc3WAN3eIXIagfsPaYXOFBuq8KRGcMAWiZs4xhlMzjE6G7fxvkS2X7nb3uCf1bt
vMTITbmiy5Vn+WQnD9WTN11zDW8M7mdeUf+82VjuVBZkcrd6bXJW6cKegkNh4INDSXmRIeCXTxek
HNJlUa8QnqPRgpECxItvSeRKlQuWCFR3aRBrnaOPev4S9rHaDJJvR41n3cUR6CjxAmix9T1Qdke6
b+wvY5DQ15ZixVejlR2e0ERCKQ7K1bCI59iVmWRglGOlwjzQkusRrazLozDPKvHmGGzrqF12hn9T
7cVMtnGbAw2Q4zM+4GYj3P6tJ2Opn9Yq+By3WiHYNiICV/ptixpXnG1BBtEqibnpUBEsXtcpWSrM
0b4evE0r8ntkQmQktDYXS2BPWERMHgYuWS4cW7eGhC860Fs9IcENAgNwXMwX6Nt+BBC9Yy6PcMPo
Sd8VT/F4j/VNcHZky/WwoZ04i1S7DXCDcY7REVLfUPQfO3JDKjEEHO9nSZcYKiICkM29GlfBHdQY
DZlcrdkcn/zha6YP77WGmuxxtsYAP7Of9GAyP65r8IHDcI9u7NOo5CMmObipvKzXP9yeDRBFOUR6
vAg2g4zGBe1Qi4dHps4r9hUBnL0MlHNX+XysVWPjalUczo5JiJCg6Xe3dFydq2G+8iJefuf5PAUM
sIaUkxwbKp8JMbSsbhSmnjsoPCxR0P9Jmn4jjRWiClDEykU5pCeoDJhpMf+4FTSMc+SHKEuTdC3/
UkxASl5WwHVHe8GCPKljYNQmDv/1boeWPBBtSL95DPOy9k4gxc/xmi2E+j6QoeddQXLW6F9A8Y0Q
mfg5w2HFOJnjriQgaV/R9+zRLwNMtyS59Vt51Hr9noiUVL8G45BGq8ej2OuLEku6kdNEvlyO/zYz
E5W3MCYxZQwOQF48Fujt0BTN3YDhmYaQi8lcxcEPLAuO7mBgcUvzoJkBgnA32oatRAo7gtpX6wIg
1nJAW1PU4ZsGJhI5nQouRX5q3PL3NZgnswI0dKmjyNEuDVb7oKe37hOyi3mJGFuefMVTXv3ZUjxW
EXe9SfObw3WJoOfwKzzlzwvy75wHRZ7l7xLlAZqyeJG1eO4ULxWUyQsgD9FN2l1xY6oUb1egxAjM
CocjH/Qm0bI9b2KBUyDP44GuCmfmW/blkYlgDWjoMm+MqjxerGNjCHBJkKwf+bKw7mTGCLZPD8zK
hs0kcigzTs04K/yFvJWYJxRwud99nO90AgTW5h1marqfrQygAGbH6vy3ANzWY/GrroKZyJ7N7yGu
77XzXHA6BEYOQ2t2mR5g6Q3jPEQydEoRL+fNzY0J/iAR1/o6+8sHjJJz6Sxo7sO/8g6auTr1/MLY
CG6QoMg/FQZp5pg7CY5xgPU3KiL4QGg27RkeC9Gq3gnUR/uDps3XpXjYkrPWv5NES8EUYs0lMxRO
zQQFDp9WBMxlSpcHvkeIZYIwgnbd+CONjqFE9vYJOA71wvGKXtUn2NrIJoAlXscheu/+elZPSmjv
apnZgqsZT4J4T+WTjEtHB1jHuLWvru/JL+oNBp+Xy5TK8dhWT2mlsuJS8D6wlqKsv3hUbBbwERCw
fxdmbDVKUk2YkXWFIent0DLxV9zzYV63qInT6THTKIYvtzGdqV3BiHElpu3A8u7vv6XhVLt4M7ER
9/mYNIhVCgdBOeo6npya28sEG2ft2AHbI7rUeEdJ9tvkA5FOz2pnD/FV2kbz8VzluJ5sVQ56tOIQ
ElheYNqq+3W3F6eCx6JMpqykvsz+zDLjRgQF2DQpZihhRsWlS3bwWUVT7sr6DibwOBLf++OxtnFj
Xf5iSWLUM9R/bUUrTpAyVSc2271LesYm+NNZT7ju6+tlf+jP0+5YZNEPVN+Fu1kvbNe/E5d7r2Fc
lwNSyrzAU9s0dLVB4r+Vr4V8fQ4ZlOmne4xcLubMg13g8mAIHmu/xxYJ2PZ44s1wYeYfqJWRlR1Q
mZMBYUsH3TuN9Gq9APJmw2JQ6D0xSrTvps1g4b9aUtst9ycVDgDgn/gQpPDxY5d/hTvPom0sY1Zx
v9q9IYfRGzOO+2f7/PLljUH0EPWeHzXFYkWmjxTGAghY07Y3YfYzSVolawYV3hQOR7gjJsQNG42j
DOzMo2UFpIA43xcvF9HTYk5C8T4t9YICRQlqfmxV0GESOjrlZFhejcKD+wKD4Jy3tBTzWnvVYeaE
c04lTWiQTM7nDrf1Y2Nqbu9hOVJT0FICJbJfamc6el1UqMeS2BE6k22azvq+Qw85p+ocVKFxo+IG
W2fgT6C07yfY2oyCI8PNnjNTq85EcHBm+ehkVZ0piLVV3nCD9brEeDqKfDB/qmkATm7Gw1FaFHPn
tny+mzLW9OfMAeMCfdhGXvC/cO3cW+vhqeMuIi47o+/NBzfxWX+lm/fJAFuNzou+TK34yw53/QOZ
a4PbQ/NsfKYm1vW/PCAFLC7Ey7ODU43y241cU65IVcq9wvuC8SPWIp0Bjp/4bFWsP1CZ6lwuDQ1m
rrbERDYAAaf7PaWciOVEVp8+pbbN8z2yz6uAKvH0YJMC3Y8Mp9Qmir+LKn605VSod/6Q4way5n0L
iLUNt7z+ONFUN82acQd2k6aKlXrrFF5ohA5r7cCjoFxe2+paSUklyOU/bxalrhvlE1ti57Krvpsh
P2hwkfcnp6YFuJTR/+uH/jO2g3UIHzQ5RQ59hisdmK4mtTTAXzgLGmkZnCYDwrNz82kjp0PuBbrp
kjl7w60K7EDi4ae6YS3QcJxyGe8iaN7VM+t+nglgiNVLrTRxCPffiGd9LFPLhXP+btgfQwOoRXZg
G93MSJ5n3MfpEi8dxq1nY1mnw4XKjL/DWXp5tw+Xd/2jgPITpaAxbq8FHPW8aWQfFsQchVdV1E/5
i2OoQOpx+H587l3ON/mvSyBBDPYwVzLrmhHvE3Jv4bwPS+Xh+xiFd3Ed5/w35KLZzUbB8zFjvqYo
Cae7qz6KRWh/bqh0qrRbz0TwiJ8LdkSBB1N2Y3m+hFNHbYz+2hE4Q9qwJ5DM9LR1c8m+pHn/PAcE
6bvGy40vOEoYmK/WrhSVRZpO37qCPTctli6iBArEXc7FljT1ddzg4AkQ1yF1c5U2rIJdNyj+IbIL
98m7HxgL+FGSGqy0Z/xF08nm8WeDi/L4X4Y7B5D6VDt9+y06g63ioR2orlEQ9DpUDuFAqlhe0N+o
gg/6uQqBUwrXZTrT4PYPjB+iBnGonGCHDE3Ao7D5HGyH2cbfUcaKDf9lrIrago9PeQDKIBtSIJtR
6GaU+jhs3yLf/k7c2m/a2ujgBVp/93IoPMCZ5Wfby98+0+OuqR8oWg+6HIYW7gMVd0LLtdl/Z5tx
dC5a9kahS4DeGchyZy0ME1enU2+ont78GBBmAFD+c++LFapZwH6bYX/yqRqfQQadi0OlayVWdw8A
5yz4SGcKGa0yUHK5maL0LHXndZE35fgWlU0vji9vXdRPmD2TG5wyoEseGUjeDnHDZLjK1tglL4Hx
RSubD05kV4p6ekmnXqfGeIEv0g70HFhzLk2tkwifLgQ9LF2i376ReixskR9dQHYg/xVCxIyFjINV
cyL7lOuRmjtY/fvE4AIAeKamwMYIwAf0x+sQjpKnjp5EQBqQYau2gOnMgIKnDu63j/2DE3kk5h6O
dUichKhSIuMmtBIR6UaNmlJm3WVsGkQsw0twfsZPcRWosYgTSkXhqNp61A5fdL/1fnca9Om6510f
DvpEHIEJoh8oiBdiJmQEqYQQU1Wla7CJnOcoB/dUKaADHaM6GUnph7QNo2++rZAGLwBeqVGEOM7U
5tMCaeVIpWI1R/JhwzHa4gE9Ycb7wcoRJNQx6aB+DRknfrk+VGrmZdjewkGbbda/bqk2+UXUiJau
Eu25xz9PaOiqoV9co75xPliFpxFEOaeOqxRihdn/gwgEIoebS5QvcwWl/n7kM3drqZ1mMWzqN3CL
mirQSypHjU4sx5pUr719ZkJNOaZrBO6sBDE4dEC7CaDcOo/S7ZLvpn005yetBmdREg0L9fXHR03D
xEA8foSFeAk9EAQp9Ulv3lPN4Gl1ll7Ae0IyRMR2yoTAS9Mzz/mQjn8d8NK9700HaAM7ITj5nyRf
um4t1RFzWgwIguEZwwOCsz0HB6CmQKqwu4wpfzjcVxI/fmvhwxAeRqAjQaPxW7YbJ31iv8VZGmXR
yIke/GGYMpP83JKSxRB9d8OCZ8Bca/0wRkXISpPMKlev9KulyFDuVdXezvZ9CU8sGSklVp/MhLQH
8JQihMVl0GZv6wy9j2tAN2zYo0WNsD3BLwpCxxWrrjaRTAB0VqeZqWjUts65hzGW+fPuERCbutnE
xUKEmaxjjMYEQ0JNBexBULtJmmjOeW5J0l9GQ6TSfPsmvCbdNqOdw0zSv51d7QWWzJwRRSoRhCK2
GvASXSb8Iv5u9alPFqrkEXkwKooB9BW5X4V1wM+o8CwPRG1upVP1iv0uE9YXOPByOC3fSAUJH60D
U3BR3F5okbtxnqjkyywO+xvH+udfBgza962xvkb9Fst7azJv75jyUnfbHNlFPONja7vMGiqlylVl
l7fB02l89qB8eOewtNAHJFqBbnbugXjFGwbIT4NNz4xwApgU3g+8PsmkTQkRuoJctbiG/7zC2aC0
og5iqDcuX4FHHZ1O+C2/5Ke3g51/Lfce3sbgdUs6ZPmm+/bkw1tzaZDFDF144fCbSrE7G4LRX8mK
Pq0aYqm/T662kZWnwj1HG10mARyS4CukBO5C2246++jTHw2+jPVAPqjlo6mDB9BsG3UNcisot808
9G9EAQ72N5XSb9kLNiaLfK0T7e+Z7iZrZX+GQ42/ZD2fqxV2RSv4ft6x2fwEmLKZDabOXekWHwlN
6FU6+r9QuhC6Ppi8hQMfXPlSNYEm8GOPIWNz9opyuBMmbSgD5xhsG2vaUQKWKQoTFYFD1T5eriQC
12ZXWSquKDGDS0UfNIcNr3CpxedbjvpSCcnoL5btXnki27hZZLZtqxJumGcqJ2hljxXkn4+X/2wr
Xztx3nCiPyjzbvvQXuJsv8Y7ZfytSuZYlcgd1McGX9Mk7LR9R3HHd0jRVcSyG/cirHu3Ox5GsGCe
E8vZSWfUl0XsDELOdrXuCbgzsYSzbXy/jtpmXsmuwR38n24odekO1urnO052BJWhLkfyOwemNb4/
0CZ8L1iv1/rip623KDLwSijfoHZin9tJMYPQasQq1GHAiE4qGTI3GzR/tiTpsrShaS6ZYqQwj4Oo
WeX4bQipNKDiLHQLw9HYQp5xs7TjnW2li18+ZnF4mTPfrUTQt020fXQzR3sqec+h39dKpLJpK7wd
HifC7QekONyP373sv/EMIYjRdtGInA2OV/AHhpIgvYhaq9fg64/RKpEXBim+iW/PDkrQsJgutFTG
5rSwA1Q6JG/ig13ULMDxyP3DfIqSNVCT0U7Lg6wgN5I7ZmdsQz3S8/EA3ALC4M572bvTTBoQtVAy
QwLBO3ntT+GTwI0kwVzL/PcHG4OVe+wbobbEG3NEEHrkrstnurMPSmqGYY2aUA3cBOFa1nrh+cJ4
jCjgx62EeSETcw2FE1J7ggO6C/Kq09klbzMtBkM4wnYL68rEJFu6ZIGKDy8XvYqwcEqK3GDhMw+f
+bQvt3PsxrRPp1iYTBbitoVGT15DkYUjMuNM1hOq7b9z0t44nDcYoWJI36IXBpqkqzjaKxUMzarm
7Nj49PJ+2uQCI/mt+IFEO0E7tA1XZeKeCkiICujfiYzGQLOllIrAqY0xz2GjH9EwnYQ0vk3a+LBZ
QSI6P1MOwRfswvl3sa5IYCTg2JGsoRAB1s52CAdJ2IZ77OQoN9iIT0F2WfhHuUanZoOe3jdp56/J
O9SmTE5bspaDwlwki6w2DgLK2EwjXoBzL5+dfZwVkKk1+BPFrefAdAVdrdhoK4nlsvsjrhy1TaOQ
YlOJf1ufDkX1GXlei0TNG46VGZ6CLehQkHcdq52dMjgT8JCCMGryRpQ6CH1pDfwCjVoT0JJcaN/3
qL7/b/X6LrQf0g7AnHu1diesY+NX8sWJweqfRfT4y1tVvsz/9dBd4+Z3PVvlHCr9C02QRLM511dH
OFlzvCXUIQtfFC4wORggGuAeZU3D4feggMo4aOCi+fcQu7+tCrAr+aFe5RM1USxvSYihZKBK+56e
l6O3LKGC19A0sS6VhkZ59nLJml9QO0OGhAjAxdblagmvhPKtfsImpI+mKWSG7erL1kvxv5Pl4ltw
NGDcgW6FRVwVrPDkwlYlAoqy4+q4jiHDLifVHwVuB2ViNP4LVhMHUF710ZHSreQtyLdcsTo4s07t
Ik/FEnmanK2jNwSP6jSYfXokiypRq61j7Vw2Qv0u8liPoc/3zHb1rFUwjjPpUTrg9elYnAs0v/t8
0074gaSUsx0xSFJZXA2+iSoqTCvePK/jcaNFXBzJltpYCPUmwpaoTMr7wWncncwfgOg7FTukSlMy
2cdn720O/x5d+3BV5OJdLwGKLM9N+wc+INQ7DcRHN9GF49lX9YBvu4bCiYze5kzztH2b07ypCogT
XH7BZAWAMj91qnA5UUi7WOnvsQUApcdDdrWXqM7PhTv7ClugDo8Krzd02AXk7SvFgqnKg4qLmvvJ
kodd/iEkRNCLAC7qSaSevSrPS+4fV5aPKfQ5qlISbckNZX55QGyBDzc3GgjDyBAphTdqw3sNi1RX
9MjJuxpyjZSw3JUOjJkn/zPoTnebLTBhxI+VQTW4p0leynPFxxuVAVVzZHQIh7Xd7cr3t63EcL1Q
4fb/dkYlMw1MG8xnyuzu89LVVKzZHOW+nw0+orsVoyTsAkJQsPNtBkzEiLkhZwuBQolXqyEAbS7a
OlPL1/dv9g7fCPHMbhMsdlgRb8bvkKpvewMrLVyxDURnDaqtxc50c35kvBfw3WT1Notn0cK27q/N
ww3IP69tDrJr92IrZ7cbI0KNsFuuTVT/IVmE8htzuYXvn1mEfxllwuKJV13kr6dXGphPI29GbAS7
jBhKOHcUO8tYtrDKkqMF6JMQAHQyORZONCyS2zzWslZLBQKG6+yvw4MAcE1XV3nU27QF0fd5qb3l
OM95KMNddKqWbJnTLETTdY8z9rqFw218M3kbFB6kkMz0dvZEdlY7TqhDAykXWmWB1xUYffmiPf3z
/loFzYJhHJwlD57r+q49negNwz1vqTZgA7WYYH0MvmxUw8yjdcFOX027uJzd1GqrpZfSVxi3GClb
gg1xFrpa1pSEzJne0uj9DdTErrAvcxGq2QpGdlP+DZ8ppxDeCI8vXpLTbGLhSOqCnTqe6BrVcvV3
/kWXjBH+W/2U6vZdcuomZ5o5njK/AUFbbrFhjRFaDBuRvnuLLrU4IzfildY+4PRf5znkPtXwRdmb
3uicQKiPrLcYkoJy+91LnlJHfjsCI2/d5zFG9deOwfIESR9yss3RSwhsFkDhyAfdh7nvUtGYH5Hq
5g+Fwyyt6gjttF17+wEvyp8haxGIEdxURfnKvbcjOs4KEWPK6HWciNT/vN7KbkzuoRfpfq1I3KzH
xr5vZRInlOtFm4E3+GULwQhmQXILaQ512erOb4dq5kKFHkuI7Zn83pkuYZ71ae+rrhkaNpBcHzmT
dWCEu2jFgVWN3EJzZmzTixiZ/8hltXKjo2I4WAryTKavjH6+dwIvCkbbrGy8cb8XfwUzslmGoDMI
WYVDd5y9b0JWOIJx2L8xxpkksB87w2ObLgaFFRWF54xk96x7COIhTe4XshVQacS8636QjSw1nVv7
+aK4VnAfM/jMMsytHI+JVF5lB0LXZbECUwM+O5i2okQu6oSDqNMCO4pTe1yZ9hSCIOjUypY/Sfz+
RH7eat7qy+bjF69nXMTHB0gLxXK3Suh+z9nG5FStu4b3RuLVZBsjEli+Fgr3aq7YR30nemikb75y
8jlkVw9dmnVZMsJ6gMAzDly6UTKpLaGHkJ3VyrLkgcUykiYrRiEmIrF4ynBRww4j2U/QFrxBemkG
CgWjzYSGA2dBEj6XzDuwln0KYvMAPxQsHrvXsWwKrQ8mdXnr4pjodWrzT5IIfkA2jtIBkV4HpanX
WUx7aihOKwd25+kgYkbQjMcKDtnsjWfumHyHqQaU1oA4Im/igj18PG6syeUz7YG9Eoa1KjWZ4WTn
j4olY/TSWgR+MO4J8e9hp4rHkTJCIZ4YGxwwDBokOizjIHEs4peJkbG5lW3OiddBiFpw3wdhIKJA
lnAiBLikGmX/1ugakC1A4orj+vAjqliFBdt0P2u2Ond1aeD/2AjJunrGzuBXD/COs53DHmKRijsf
UPYrwtLqvzOMLOnSisinUVmKxCcvN/7OfBmlsHYhf4aUqfxPOtZvFFU5//uoC+ZWn93O3XvS4W11
Sp7tdyF0BG9vbf0zkhbNAnA5JVLS82fk9B+rESfH6JQwVBZe27TirLgqlHZGDUXUG5XraViHFkkr
dJ2XWq7EZ7ZST3OyF52KADnmmzgagPciCKo8nTK0lekxdfhXAQ38BhCG4FV0BqDUeGJEoIFsQ75H
5V2ZVEVa3jR9tDWDLINcFZUP3ajBzw8tv8IUWHKhp+9fv7NlvceUf667IBk3jXefGgJhYHR6la2H
vqvzeOIaz3PV1ft7N6cJPPxRQANCToS3TPO6x74KD2sFe89qCnl906cFdSQwAglF2DyHsMOSSpuf
HEFMtKsbgVkQE2tNAbWZqBlZt0r306K3CWV0GSw0JGwlCUdxz2XOvG40rYsoKPr6jp8zEMhZ9RLC
p8Ge9Xs6ZcTx3WA37A8g2+hxROPafuvJ9qOja7QVAFuYhXSKAJhddkAJMW9lTFjl1gov1yRlofJ+
4NaJ5quBCTtyCS3wzIF5C6op0jeA1RAmUh4/oyZ56YZqkfeYSEV7LCan3vh7quySgqUPfBhaZcPZ
BQYGwRmo/4mYJJcw7OSTTIkdweg4OTRKaVj20or5Y0/ARpuA9Nhx1X1b05qyr96WDL0Ihwe6M8FU
C91GnvevgfFHyAjGdMG0DvuY/zXgZiUe/JKB3UalflOehDWXoCgrUl+sdw2eZ6z4eCN4/arCvIGw
fjBMxqNCX0C3/C2UsZjI6hGcHr9JmEVa9uNNMtVvXgGFAePN4GBq8nk7y7wo7oAnnyRV9q8za3ML
2tlqnp9NKULwXQXC5xY12VSLC3+lXLGtWdAgnXNFLpefl+XQjrD1SID/aLkRkppHvWZASjiEkCHX
DKfcr+WmXxVjIZhtX+P9JmaPfxS/EB7vTRGDSczDpCUnx8LzvcsmsqZWcVqUWBAof4fvBIffAiZS
LifR6Wv54gHejtqybt6m3OycVs3YCOhj2t706QA+ARhKOsvkecNVQGZ3+ip8biKPkJvkI10Zp1za
dglQRxzgJBa02vXUMjqqZ+lXugBznrBM5mDJW40C7CcbjX9oTMZgoicYRt7CsBmkveY7mRGV71Qm
KN+0ARiH3pNg+QB4odIWwzU9R7OPMqWHFcQIv4pLi5cSk26ngORe3Q/HNaa1BRvEdJ9pgdcuw7bu
nbyasvUIoKxINh2hjw+Y9U0Ku91P2jr0Otbiex7brfpERQIRrXN2C2kdOyLebKKNhsNK8G2kIFGf
3adgQlq0jJQQSKQExXZTCgy+p8I/6cW0RhrJYPrAfO9dLho3EmoKzp6gnCllSBoPeXymAwMPRqd1
T6nY177P23uflKfsbyhNJHzGOCs2Wih/omHQmdqV+wjc3xEwtIjJTncCWHIf2RCssPBFRf1ZCzno
eDDc8tsggS+mJ4k/g4+gWiOi3Uofax73c6FCLE7pHu3+O9N71ga2hBipruM8o1RJauqkELqfUD7S
8F89SRZsotFY5lca1Uv6PUqGRUALmp8Th5iltBUZxWSD7Iq/DBTp+hpVr5XyLtDb4J+9OHclgb5c
/Jl0GAaGUOJb4H1m45z4JpSGrc2YBC7Jw7pz/EFlKNZC1i1HzMeTiLrp3hZ/FCUVem3wGFEzm1gJ
ipSaoEW7c0mBCMRysVo3K/LTdA+NV4oOvxohPSJ0t9Tn4pc8y0uyAS0hwTyHIYSs1H3bo1m/4qKh
EwyzJ7xmgqyDtSAradGiUw7yLLCDVkZ1lBLDa0oZuTPGQTufwEaWa9G//xyUlDgVPdY26QbwisXc
JjApSdkCiCUi3m78O1QLjrCyQNpj12z5gH7ecC0phfqN04xEztF4dQj7VGZkxzdR14oOrcBjd92z
dZP3k8Q8XaYWb5GYXv+DFz+9MM8vjLe9R/vzzwqq3hoeFlQdOmfwRULxobW0wK7XNbqsr/wdaeVw
qi7C0hyQGwc2Rv1zFV0RTQt/GeFU6/llNFhDFekvWgv1dyKFweYkGHYHqY12EZ8cv9byVmqEeMLc
/iEE8dqjY8m3z1D+MhTLFC6v978jCZTPCs9+b3UjvipCRT2DrTZ1OQpzdXFGity6+C4bm7dpMfIW
TYzVlnW8EVBxwY4bXXS9LQk0ENrTQyj1WwDN9QeFPTqBfM6Lv3tGP0Bu3tp/34lO6dzjqgtPC3ys
P12jYloxqSv/UhW/6LJFb1RI9unMl87RmDB7X4Ivq3u+AdH1jIaad6nG9WkoEyt4UzK0oCoEb8xu
CunKmTlgsgLhYHuJ7Wvh4VkWbWzQfqsCIYdH22dvaIrJv2GSJtpk9s2eN1ZJqjNXpiJLMm4JR31w
CBKv7DlNIbTXWMU1ln1H0VSAykL3qTuRtI8sfUCnc94pQ6aUuFS3ndE/aJ99yRKkcRMlYox7OEzp
dZbJQ90+ruDfid3Mtcitwc2DLfeOgnCVj3GdXCEUBdYB8BDMlaVs5wGE98lWjf8s+T/0JqZ942b/
VDlMtWpzqHROkmpywBUhlXpxdNQmDKqRKvykLoQFCjENvnDe8aABgjh823elhAsPgdWGdCS6egbd
ApJ63ToI7iRA+a/Dz5/ZNEUS4yv7s8wJG36U1Nue5McZ4PtmKlFTY3lAkqtBhR+3v3DX05XjnZgK
wByf1dsjf05npvUC2YggrTuwwOijCv47rRRw9v2RWWLCARNXI5G0fOL/dFo2qAu3IcfEETjPOCkE
3GGQfSkW5ghrLuRteiQFZAknDxlsroFYdv7JEeBl0lYLSXJ5bn9KczzwA6zfJyloRacWAaLmqVX2
wHcPoyi4J2xji0d6WFR8JV1ThFMz/AiJITGq+MX6EMX1qf4FXvBjE/Zh9gSBemXbfqEHZhuwXBC1
HkjixcrMmuMWKSCuUyLIDdtwm5LLmQCB/av+8oUTI6xlbD60w3Mv6FB6ZWtJQw5vDRbvRTpYCqfV
HGBtw+1w/Z/J+5T55vNe3tVBNEsrsiJL37NTzUBjOqG9o2NNNXzT56vNuw83d2dYZUcyiG2nLKN8
+5dXouR0Px+7pCfpaHiWzIjL66PsnOd3zQw1cvj5GeS7/gX4Ug8I8vwrvlvT0wj0C2ZzDGuMT9op
LvHNZfBGxtF6PJmM+1my+0UOQlYg4WvCt9p2d1yg45me03+1Nx/C5Nlbjmu3Rm1gYipnrh2y2NMA
y0FnrzaThL0YUrU4PtTrPxhFLelZdjhEVItpexiVi5Oz87Gg3zzwnIsFKJlh2YkSlVSuS193Y0QB
/nuInTEOwqVOSZZeO8JbsG+W0i+uCWpE0loQjk4NRAOFxTZU7YQ2/x1rNmh3fmVfNnZDbR+WNijf
D8LTFGzSI/SnOuWToKsayZc79sVG0CNnNS1qPACSyG44rSUJuU9Kn2LM7I1/X7TNrOiSwqBhXGhZ
0jintQrjBzS+zWRQeGZSbjdNpHC5obyn9GFXHfGh2n4vmg9/DksVQ4ZwxIi//p4JgV+JVucvASHd
VrLcxHWFnXPwOPOiCS0i8uKjinBVtFUeNIJejE/4IpYH0JXKCLJXWZoZwTQBilvxqgPm1nU70D6T
gmBW6jKLETfUEfuwnCAFyEn23h6XAZs2K2F7n4W8rbMoAwagicWZ/zuDcLcDrIQcqqJXOCBbLmFW
ovBiMXIp1jo0Du5CteIXCEKDP3/jhRiXG5UGAqmKVFda7qkGEVufhh8o8M68gxN9/CYu8rk4zuT4
sU94PScFS8mbA0oPnr+Ss8XoSg8QmGqKlzbOUG2xloDidtEK6rbwKbysDx4P/h8VeQf5DSpniWhW
7bxpv9jf5XosfyAIPsi8WroryCPiFcfgrhAgfYNsm2bqXuW5JzFc8LUUoQIReZ0rYr+cCoafttvp
qZnEELXVWVJPHxPZiZN2PcvqAoJkZdJjvC3nI1hxbZr8g0yvMlT2ZgSw85UHtWcFnCKYn0MIfHdc
GZ7MvocS4AqylqqU4O+OstiJk9ep6h81X7x88f1Lj7cG/ROqngotI6w/bBHtYqv9wZ9r5QgkHBPd
3YebZ+A937CpMg8zS4x0Sr+/57fnaQ7jHyIeSFy+RjqLctC27VqU1S7S5yKRkrjvLQep0xIZiv7a
GWuSrT/gpINseOAPD9JgUA2v86jcx9d4AGiyuwhRMxZI0OTFDPF73cqHcIGYghDVmhLWGPsxia9M
icjPr+dLMRcQyVAXgJ8FmWHodGGWffR+pPVoSKap//H2N10G5Dni7WJ9KvMhd2w+mf5GDD8sUbYm
rtq+107QEvD1Y4l3nwjCLsRqv748u6eYHFST0dgVciJvrFcFtW/8cBkxa7t8tkKoghtaSZ6xTzGp
dvfG9mb5Ocy1zpauwD6JQmWwdG4Oz+QlojzsFl88eTSAxFbbwLkDiAdNfUzq5WRd0EHkDPyUuqRu
Shl5LeN7LkeNLb7cDDY5fJ7vFt8uarMU3VxvbDYnxVQBUdchNiaLDg9PzJyZYLHtDaMN+Rne0Ht+
5CNxIIULS9gdpi9LdNUWjC8SacTSKaIuZsl8shL2BncQTDINNFAxvct1zbI/CQV6wHnDYL41j1ed
77bgT6+G7N9YogKaGztiGqwbB7Hhe5kzYCXWzOdEJ0/kEhlMdvxSEy9WQdgdvh0hDSkEcwnNW2JV
IYr3qx6zKwSHB1gHnSy/cayY1xSvJhs7/IgE47PlJnMNNG4nU0CMVHtUJb2mzRWOzOUd6yavBczc
LqkSThg3h2lXR9RTFiC2ck/fbWkLBHVgPtXMszaj4qz0rVooknatgQhbQ4hQThbesedhr1VWWZQj
xi8Ugn8DDWDhGOScz4fA4EGXd2EuMs1eVzldhfnfGILgwbQlzONAZ5n7/PYyZ9jtpoTwCVFhjw6p
aQa5MOYIv49XTO7/MIghmvO7qJsONYAV8JOrAk4jbHowW7K19nSk5rhbk9idOjxmRAz3+hQlflsy
QMKYjQrV9PRPy0tW0JHFkXC65e3ToIheLXsx3xY7rxkJGPV1jU6UHT+dJmL7E2uYPd3WPDNYs4AM
4w8/tLWzd4MzT6NFCRFGPrCivc78a04fjQ3aadCoQhokbYeZjSwokMkeLhDatgMdNaxeGX0V/7S7
lTcEJ2X8BJbAM2qFs65RTBulJT1CQPuDkynGUEeA3Qgg8B1HysxZuq4Jjxr3FScED5ov/nLaGIp/
isXeH8bfGJ5eVPp8Y6ghIRgqvry7fJmb6WicGjsUmtATuzD1YdYA6Q0T6qdx0xz4cNqYBFnN/GPv
Y2FxLpakSi1MPKQEFdn4ZpWdbeIHdWakJsK3oSE5KhQT+3XG1yyqq0056XragHvKZbExxX0ikMzr
rW2snVaVLwBQRdoIhq6zbICFsKXheni5pbtlqd4+MWFyAA3cI4h4pIIcfdR0QDCzQrbYfA9VkCqy
/s6HADC18aqIaUZRss/FybC+MEmtgCrW01C2SN4toaRb+lnSq+8luwF/zfw78x4J3mwlMrn+Qme+
9VpHM9Ux1Hq/QoFO23A0By7P78XKrZxxwDReiHZZ7+LFgTcRNOMoy2L8QW+uiieB+YAjY55lt83M
Cq5iCPnhs1adQ/toZyWyv868FwfbD1IewYGfdGqyvHmI94xLfyt9Ia0SUm2P9LKH/wY49ZDRgZLE
H/NektQn4OSudkpGQDH3w3764fwYCm+FWnEX/s2y37Yo23lGovQTqNzYPgYpaS71/jjQWhMcETax
ZW2598IVD1R+agkxDNnsEXAPmwF0X+RD7uBWjCV2gB/QcJ2oXHp0bePQ/PAcZEl3NBZiQ4KCkOdY
yKaB2sHbrgSiiVvtVzN7SjN3Q4DdSGgHCQQpc/U6ZYyIyYv0/xGzoJBZP5jaZhrjVvEY/krZsNM7
w0SDwuQAY+MtM2h+R7xwgvemgKb6kPGAFCcAzPFyhRX3redMLXgDeYIFA7a06rqDc0SNtBhk+cDN
veRraQtdMmU73AT1+csct00R6WePJGTD0TUrr85SP8XPpXdxN2DRFRYvwJATPDoTnv40KdVebNIZ
7yz5I4xkYxbZ67ldWMu74+YF9nVHiKHeZfverFQEZmAk0Llm8WKe61ALcOxdahT7XFkIZL80nnMt
5F5bkJ8MfE2R6AZ2fAiSoKF2ygl37/+gFssjoKc7s02Ibamj+DXgWG7aUecYCcfiYezLREqCgaEG
rjkX4UDMOnZWM7fU40MXd09i7H00ztrVtd9EVar3apFqmHu6pI3QtHYrkjRaS94gOaf57UvFf9/M
pi8wTxSVvsx9eQIO5/uAvEdtnFwJdDdVuxJOIoE4vdECstBIfU/6JYwCt7fGt5N5IgJbRrH98CS3
fz0jgx7NuZkKVHPCUuzSYdZD/fI/zgmhdJC7qOo2Y0utniXuib/ASIG7gVQLWu/anne4AGUavUU+
NjZPwF04OyClQ4cWo/OkRFmkhy3DRzmJJmL44afJHUn6aCHiniIwOIVruPScA3lnVhs+TYDK576Q
Wf4PltGX09MAOkPXHsLwjxhAuP0eFXhatHNeqtRsCJy49dTQ90Uoxtpdy5/dwMWDLNr5j2S1yzUX
8rjp0iID+Se+V8N3PTZ2DEf0hA8uCafMxymFTNcjROs/ugY4xzKPy4+DzZtuYMnjC783CuYcJs1Z
Ug/crkolD7a/uVRWlWDLGq1fAfcE627ZASWMHgkkaALPJ3pBWTlrVDoKC80D0y6WeAb0K32nXxap
XjL3HcDBx/cJ3N0Tpbdjps80zCPryFKaB339mnQMNziad3J5366+HKi6Fo8Pv9fPhjkLTIVO/580
/4uY/nDT1EO5NqjCo+hJFggwGU5Eg7G2ECdBFm8gqNI98IpajhnHfc1UJxxYIh3sgb/To+cinbO9
eZUyA8hSz/tx37RAgiAj/+EP+o7SI6XFp9R4G7a/zJeGeQoXe3M82+s1rYtfznNcTbKw8+TrpqJm
FaHY8LrDgQZv2SizXBDTl2UQXLcMOdARwVIY3djTyWlSz8l/gf7iIm4X0WuR3LsvkcjgjPJXC2DK
m+XsxbpS4rg0jl7q6pVuoEzd18rp2acl/B2XzvV2EZ5l3WMmTKrtBN/x8T01yESe7oA1M2ZpO8kL
LoQoXI28dyMweCiE4kiI4nXkJ1zLYxEXP/wYRwK2mnfXU6EHKgVpnUwLtjcSVXojTNtyhH14wa+1
88hWCfw1SWAMiwc49vHGxxA9o609Y/Gg7EHmU6QP87+WJfU721QBTpDJcjVnxtyTc0bQipt8UM5R
+nBs4u/8HXGbmAcGwwXM/KSQQyvncrMmL8p4B4lrQtIsSFt8KN43+YR8qE28ZL/6Qlyth+g6R2HE
Sqz06Iiem4va0zxGAMUcW5c0t9rbwlJ0Vx6Oy8d1VEfvhWppRgCHc8C8bQDP0M+dGYCOzNQiFgvR
qCqhNxaDa0/ciEKJpgJxq25cp6jNCVskIUBC59GtmBNOTkeGe1teE8CLcCrKkYCLyTz1g/HH+eBC
eWkslb3pa0O6T88QHJ2bJPzGb537LnJX9U6Geel3t+P2w8Rz9plTgKTkww+50Qps1dGEL8Ul57bA
FDUwh0uuTIWBXxwtBdIc+34UBoxbi+ZPWNDMT210LwIGjc7n6bERlQFT4kddlM0ThKvImuNLllpf
BgPtterAPXY6XjKVRUuQFaG3YRMBOk1McCgqWqAjDfGfuXsY4/4iebsKmSYu30hE/AyEMVfzBqKm
G56PnL3UWrWgOMjCCGzrsJgLh5HqHvWcuc5oy2/VS6uLwzO4VrHG9gpWOUhOpvL9GFpSxMe0tSjg
Qcx9DR4pPNhKpMEtsjN0DW89HDfhkkHKg2dZxhCAvQ9A6y0i0A9mHl70KZYKP+heGoUqULUrFVV2
h0SfhkoCoP4bcLiZoCZMBLy8iEkbmr4j3rAWr6dsAOXamy3fQC+llmuonmSd2rUjQD/uwZIIW91V
3ADIyhnEaTo2WWUWoK8Wp3jp0bDDIQ999pBWeqyZN/XO2Iya2oKG9powObZJ+SfowygivugcVmcp
2OfNWZdL0rULjSlMmUoljzNOMfoojStHNmchAQZoJO54b+kpP0Uw0+Qvapy9A9iEtPKKHew4G4qf
hMaLcN9Oqqv8bk8ALnF0QWifun2IXKzjrBIsAu2GUb876TOfBi0F7pLC71SLZzphSB8vDWHanDtV
VLyB1l2VIj1RgkkuseKhELOYULZMmpgdnu2kZpzQm2Z+7nh7NEer3WGXnj+in6ytmf9iEorExP9H
X8hRtj3l0Lww1nVs8JygOzQuSuwHRnWPQNDml62YMv41wh1rATKzAQoRPNh7bJeaBM8cNR/WWPSz
43h/FXv4wcpYQ/riBRPgk7cOhF2zUP/owE2OiiJ9T3YyDPJIFQCmKGj8RLUTea8rN5/eMzj9hdYs
2D6G+q2ZmFpkj3MnkJQks6g7IPwbnbDVK0yZfbWwwF8hqulJ0r+F7Vt58wT+SjqpeIGDHeQbAGbV
VVd/sjCbWvt3FEhqpj+yjo41yIGnEh53BZLJCJP239vKE3XXfE5zTc1GywpPHj88YQOGD+DkAl93
IOopaqbDOx1CuyIAPHPDVGtP87xM38SBOewiJcQVn6XJqXRViid2PchXDvK3NOHIs4UatP5tKvM7
ZRw+tOvizhsp8345Np5Rg6+f2M7LFuvc7+2JTEx+8Ih9Ozsqn5e52CO4ymCpda2LUXhWrHCOE6Mv
Q9EhF/eubWAU7JMYPm7jwH5ZjPHDtfGX6M3sFO5aw1lBVlezN32W3T+dqQ7y8TCVTzDsZ25f5/uT
ldegjKpcc59GcQSFY1oMh4Zc61MTDT4UojzzTB5fi/EL4lBbNnrvgt6NcIet89ohkVYvPGjpwMFP
meiHL8UzxHaN/IwGbVefVHieCHtwtsdgILK/rLhTJUOVOBv4gDs/TawE70IlFYoYOhLHo3SwFCFy
VTntTlJB1ob8Nh+dxXIBvdVxTkazNnwByeOOJhuQnAke8uAKw6KqeR4pQgR+XGcPrClpZ1thHDBB
l0kL8h7dj0EVirWpuMCjO1u1prF86P3/TxVVzyucB0HhIY9Q8noy+R8nRYcjNww+dt/MPwTufuuD
I3LjDMDpB1zK6GoBtzwg6/FSX2luIERKE4fcqDp4ro+pnsrDU/zsYTrX72zNATl6vNXu0ZPlhWge
Ww93IhyyPDcodDApieoll2aJPhaP9PAW91CVWoUeO06EE3KgdGClwSXbqlQ9IhonNMItmrY8I1pv
hHKpevw639bq25yYmOCcffT0WWYgJBWByKBKzTaTPOvOA9neWht/SnP8aENL6S/yta55KSOuRZZo
qiQertCyb+kPWBZO2uMd0LaTa8jqB0NG8+uiWwXMpA9O7o/JMtmHjqUelooj5mj89UBIcbI/TjHG
raBx5UBeahFkoU7eJW8uyNogd410nMk0nDEQPQihrLEeI+Tfd5IJM8FBj89Jiq+bNpq+tjOXJtz9
Kjb1gW6mHjv9B8HheCQaxVwJLT2EIEuwkLBkQNgoGmhyAHczG0MeoriMCguCvvQDFmiS+zERB798
kcHtZUJ2vMR+X+D3GZnLRXGTnkEG1evNWiJ3pe1QXhT/Dr646KtRDSZIHQheUv0RuXezHoWk/3aX
GdQ8dB6D7lOdOiM1yag9y3P2sTl27g5OWQKoTT2TWgzWYkwhQyuQnYOTJ8/2RQHmai0OZ0WhmW+k
DgvmiDK/cD8B678cUBcQ9eR6zev5Fg8+u4rV2MGKl0fmv4r+bqr6SYRNYR9MIeVXhd3viNGSwlyL
mjKeFi5FRvIZ1wzfiKXfaa8jFFNOuVSRwSPj86he7VhOgpbcyEY3fcR/10+eZiwsryKkJHTwxI1o
07WWa7fwZOLYb2EvF7IUc5WFNBBux+cVj9gZwVb+MqD+xjBCQBSmFP5OZWONMo3QV8y2wvMx2EfQ
wqRlvm8LsykLKhaKutunrxQYSSie8CMRVNLtu70XfLaxiTCgH38ZAeHRQK0WqkJHrbwsZ9KuLt4S
j0YGcEq9IYfWS8uzj8s32R2Kha/64eduhUoYMeUN+5OFpNCsw1HE9mpKAe4/RBLA2RXdRRMFEGIm
iSaBeFsnVT9W2WOdVvpLICBKiDmZvPDdCFF8PH4HvTDwkmNhvQfyYNQVZaqSyjfakGQMa5wUVI8x
YQq0e7pTalJmwu951f8/IrWVMTWLgVcjR2v13omkp52lrWrtPkE+1R+LsGlPz8nC5WoZs38GPW4m
VOI/n7vR7eVLuZR31YH7l000LW3GqKSKdSeldcpt348ZNjoOwdSMGdv21+FdasjW/3z4mE+7Cn/e
+DAQs4UdKJCchlES/jHI8wMwieQD8pGRstKer3OVlT5w37MPM0HbB3uXU+hLRtPkVeuHVOyYQhnp
Xa/1jdZdBJBhigz95K3JXFM025f7HAp5BTH44BFKJ/BPDuxiHaPD3QbyzL20As7XOMZlwrZxMP27
jDPvfl/BhrvasYoV5p3v8s5YxrLm8vL070TNW6Hj/sedqxM+5iHNnj4PUEiWc/4dfXXRGBFgpJ+9
faScTK8lGDEzQqrtkf42WmdF/IYqBajO6wVObmQrTmeY09gDgQft/NIZ/WLBASWGhpfv9BDfZdnc
Y8LEEfFjGJps9i8oyOySzCoQ8gxOu8WBFb8MICpe5bAC0T4nkFq530zCrif6TIJSC1Zfe0Abhtj5
HJgZKxTDZU1tgUz/oioRW/NGEmNfakzpZzuP4UYHneivIlae32AU2Ibjw07YcI6oOGOqIqSy2ra8
l02MYxEK9JrWHI+RoiSUFg9Dy9/LlI6O3oc/97lzVF/hXMY+w53GUf/VqWIwBmV6eAA67smrXbQT
ZusFQ8Yo1LlshUowJC3S113E5iqAJL7zhC6PTjCc2+Ke9t/GOjC+cv+ReXuVO3RL4crPJY30XFoJ
36rqsNKErP6+E9O4TNO2GPA9ZRAG0STFVpPB+UMX/LyywZfQMljx1RoR+kUXTenpLR8s9rX00M/R
MO9Bhob2y8T5kKdF/1Df+nOMb8bKmyEVYsKg2NdZo5lbRi7LLVhKZ1Jf4S5s3q75gxOJ9vXiMIMC
pNGtIhUY9JO8ReZ22SwNFO1X5j5RLa56lC96Lvb1Eni3A7K+lXgEUUtB6Bz3M0icEBhLG0vIlKLy
DItINy1h98ufE4JS8vQDVKHVBlifR8YrsOwHEGT6R+OKsah13L13y+2d/VkEmgvn9T2X6L75BydE
dlsGlw1YKwDqD1fTCoeea0S+nMzj1sb6k2xqu6bDIBQ2ki/XillymgYvsMUloVxNhwecXBXC9jmV
T3y1u8OZJF3aGiwkWeBoq66IELiu1+elD28QabrVwV3AyRswhXz5k2rQB9q2uwYUSb9DfWHUFqIe
LoNmq7Dnzf/Vjo2zmJhKyvKg4no2oKeAnu9s1FKbGIjOsHwoC1x5wC+NAkFk9vRpM2MA1Zrog8vG
RfMx5dvM7fnsYIZUKsXXa2lxhHIgWYbCNGTUu5E3O56FvSxPRtgFXQo36xkGjxr0PLOKGCSIoMtE
06NfpaC5Gn7YggwBXz/U58QT+XVO9dnAkYoRQ45kDDrg+Ug8dCKEHaVvlWAzNvCnsuTEdEa+8lC+
ciLxqfx5EoREmyipWSG5JLarMoKQveypW9jke8shvZytMV3NHwqibdUNfA+DT5sl6W+CvY1jK6N5
cGqHiI/Q+k6l6hUwfieSPljhRitptSeY0+rmDYhKMl+sd3pgUzjM4GWTNwI/VXx9rT9jVZCBn5ky
FcZg2syZGto9Fky8b0x39oCojOEcw8d3KLiNUFklBuFAC/IE0Hes3AF1kldO/M7+8zS5ZTycC1m7
0JCm/TQ4meTb29Cvu+3ksmu4ADUF6r61pr4fFYPqIORgTyyYlzORZ5ceEx7E+DIHnNr25HMleKit
0UUdzEqkq8kKHr5v0gjofRZ6RmcZ/j8BispR6Vb8OJCz8+u7wFNcAmDCNDlvlePdoUYeiii8GwVo
fWKhy7zSlexNHvVEbZ1/DMS2LaqfpkYMU2c4VqhKLY27r6lQFmnwzVL5Wy60nWiafICiSIkHdazZ
Pusy54h2mh8GaXv/OuM6yjDzhvC3Z8zD27F60lL738UIQj51UDk/A1R3rZyNznPgHqkHQ7fmmVSe
fWk1ct3ZtYUJT8Dowkd+Hz1EkRvMdmBIOFjIFm8q40zw8un1E1dU/NCtIl8o5BWuEw8eN7r0yRFs
Qr8neZ/B2f4737I3Hj7odwbL1CNoEyXIgeMkqPSwlyZYJE+ldpjtElbG6Xj6G4ujf64KiusR47rD
oBcOlybfTrEt6twrofSjIn90ykqQbOPejhf+rc8E1dQ2fLr9MeuFeCqt2Y/RNas5wTfh4VARC46/
X+MUq4eQ1b8FihVO0Jv3MRGNAlroTpF/ktBAnYRP+v5Q1or3C8bwu81uiVgtPkHsN+W6G+gSe17z
6G4qxcky9ZkalKyLKoKb/kb9Fi+3xBjciduMIafM3fwBZ4pucih1w37Dk6mHGxPUDmZR9RTXL+9i
sFK7s2FwfBhC1jhWc0kEiVSxVQWbaEoHasff1+ymUUo7UBRiqyfMe+bAQyc6fqhLyFYZpVhN2JBj
3p/nui/2ZokdF4jk1vcaZXUdg/fU9GMCvJJrlb0z5qfZ6znZ41xTP/iDFPsMOuK17z8gPqA2BJLQ
EFL4H97CLu6+0ouAi7+QTwUNkooWa0gmXHJju/Qe1+OSEU8L5RazGsm89faxLru2iDep4RfD8bl6
e7GRTqjMNixskeb+xVB6dwUWLFrsfUYW7dNzeCjIRJBW7xm/XgSdnjd/x4UIWNw91Oyl9M3+Q04P
DUavLcfrt1FPAEoiR8phKUkIp0tlvTDbWK53fQPLBXAE83rlcZGawBckYyCNNtuCkF16bNaPDO83
dSUx8SJ0ThhBa+j/4EdcwJ3p4k+8hQUgTcSkzrDE8w4Rp84UWwfi85IPOetXcpdzJq717+gsB8E6
b6N6984SRB8SHeEUcmv8zZE46cbpvCeoLTBFDGTGxRLznnbyhbVdkzEd5x+Mp2QOwcEYKyKn2X0U
V+WxsXrEepXrATE2Jlfl6k3U1qzZTJ4613++vjKYAsaR+Nmw/0Q0BOOGTjUwXW4unBAMcFy/P+jC
/8gUXrF6wzR/ruM3E5dVhcEcgDEYuwPxk2KBTiS7kSZAOSMtwv4NLOX3q53ANqi0NaEfAa9zRKPf
dEXeniJUXX+Is2epKmTJDTw/TaOHc95oOLBsODBR0qSRDFWqN40iqV9GFKSYLDdX4GGi9LR3Wzw3
+wV0ZhaqII2Sivsg1tieLuBn/DKsi0RT+w8POgduuWJmQqTF2xWpGmsux8plzrQMAQCSiFZ0gEHJ
q2A7mLp4LVkCkA+1xOBl43YI821jhTaF0YaRc+WKglnLBT2/hiVVS0xBGG5O+EHlMCp0ldSFX7gm
RaXqoJt68dn7q3ohtI6e/kUuzoiXwSFRYmpON9KLQFAontb81y9ju9sUmgyt7pxSiSN3qv3vVFHB
eAJVuyFlxOxdXlYKH1IBehvsrPqcyLmnTbtymeQkkDoRHQx3vYQMIpc3IFqoXCi1sgVOQbGrSD8H
Cmb6RKK1kXBF+8gOhXK7+0CjgH3Cnn+j4AVm44I/F1LU92TpxDp2GLmYVpN7kernbPOHxdZLSjJn
S9CjOdLp1HIh7GItFxoXyvarBY844mtTRuumsgUVZNv03Li+wVGgU/B6RFffvGZcplkcOuKKV9Lx
b8OPmq7I07UnmPT8/X7eZ0hzp9gmYppzVbRNYaKFSuwpQoWABApqX5VecRHw0Jq4F7oCPxv/mJPS
x8ehpPBs2UaZTjuU+GafqOQONGiRlA+ZS6Y56ebDggCo7627A/FTNn0CnT8ciPrdcy9LdchrULtH
Kq6LXOt0+SApmoq5D4ceWa3rAy1vrRNvygkFUtkmWhfsARa+w4fyjSl/nQQyxin6XThIhA7LNqZh
w9LhdCJ5itZUPDWUU6HiwfluBu3616Yzu4jF0CLcr/AMl9h8Q0/Ry/plyM77mqMX+ws1bljYpwE4
1vNAuk3M4mY8+ph5Zze9U1ohh6XCNiWiR2PJx59bYf9TKAtERV3I/B1Zhln5u63AGAopAO1UUsBC
IeoA1XvUxwpjBqgdSWmARohS9FH4xedrReEQ2OWmPyvhWhqI7uBn7gY8A7/Ruoz34j3kTIy+o6yn
/IjnrK6vlD2jafBLLGwq9NsD0AKdxCLCHFYqJABoargYkgJTz8MrPng6OsqhOqs+Beag155mQS9q
mlcbM72c47W0VucSKho4G+bpkFNmQsOEGql3muJs0MFOisE/Qj66PFiCbs1L9Qmb2oRJGlN6EmIW
aiBVyppIyxN964KA0/nMUXUTWX2sgmmtMiuV7nndSGwNrTnAktJffCm7V3M7WVvCTYLpYN6B3AZq
2THEk7IfbZd5uvchLsTAZC89y0I8GCmhhKQl6LRGy7/xI7fJaWkPB0okTM4gsvoKRzz6hGnQkAbz
EVL0ZFBjVIx0wzZwpa7S1CgxzziYx+KmLeU0nXEZTMJ5OxuX/aDVUVpQd/w9WHUJ4Ks2a+u61C2h
emjsyBUIlOgu2toFsBzOV4JoQmPL2xuE3HYt0Zs8qbMVmL8jZBV6nQvjY8RwGux0M/+8Wz5+ihx8
OJdz+ts/WRPvB6b1C4/Wqx+ZkVbH67pbj+B3BHuK4KvhItYpGoKU0O/7KNE+VBQkyM+hCgdqKo/l
LJnCwRoq3mEgZNoiEOVWhas2VXo16Vv7ONo6UBfDJHSIvXRpOhGl8irNmIciGVAaztGi6N0w7eWq
zBGFrHzNBZDCMdm70AgResxoJ7OF6/tGmuLqleU1Tpsej2rKvBxKQJbDKwBBdpJbkDd+qjyuU9Dn
JidKNQ38EvhMf9OLYtemJx6kzZJ2NBPjSBMh99QZV7nTEWKegEEZzfL+1cUlTocS74bZ24/0BjzI
Bimx0fg8CsEjPK0PKEJ+K8oWLj6xcxJuphC3fm2vMcg+UvUeEVL7KZ6yrSGruEEryGF/2HdaJ7jV
bnr6QDrZmziZC0E3kiR9OZM4C/PS1/5g30mKtyqmNbApXXAaZmWwAVFxw1l083w5YFhv9PyBxRHt
baK4+Mn+BF3GK+3Xgw49wR06COXJEVr3EzuKhOej7bFxY9Y68nzt93jHU13rm2scyRIx87LM6mp+
qy3Tk2VfPO0dMHveEr/FkjDLt6CVbJdcaUG1CXJu33LOlfVKSXGi9vRNWRQB+Gyb/dId8IVrYSUZ
uhBgAk2+hfIfF2zgVrcKkGr6IJT3manDnkALRE+uAydGR2D7MULW8aGZIRUNpt8YVX4gKf0hqSXZ
FvGRWRDo/hB6/mvw8L8eEIzrZvKfYb6wgzNvM1ZmejfBpcJImQm2arHdfaCxkn4bUP7XVxiqUqY1
3SneHZ5lD+kGjs90lM0rvsK/fTReTPg31K7l/eXYOtBoLQbJmRS6BdmbOYUdggAXgNS+5vYbxw5Y
yzweG92u7zVfz9UC8W3OV4XHyNB1mWCFSGCSUGffG8iaa6gzOkkSsexTVyIvxrWmK5xYQxhd5nTy
J1jEM5XPdyK1gEmzKMS11Bp9x7y6Mp+1ZyDUq1idhrJkcZYYThbKYtsbw5474T6yH5E7WoBMxQm6
N38rQ8uz8lW1sawdBcCIuNX5n+yAWY7zy2nLtjfEuJ7/15O9ABquuz5Ps/4wnPj14zNqxoCIWSms
MlJjrVwFDEOKgvH8fk//AkLmug0AI9ukwNnHpbAYMYv8aeHVTQA5F/D/nacD39Z9jI56HEAjHe6e
kflj1ssDHpe3zQ8no1FHHmeywHp+b8zxP8LAJnNT2KNd+9OKeO81p6Oe3r0X9a8wxFKHypTyTm0P
yEpmtGGpDxtp8IL2KpA42oWscO7pfbV/KFSoMVUSxxUSHZcfyMniH32MqDsTDV6ouzcc25c4r1uf
x/x1oI/Aj9NBhCzEpFeqdN9LHk1zI7+pOy4DQ4tViAl19uY8TzAtgHQ0OFVJxM9wO1Mkqd4Sc1Rq
Dx7/dwllWVAHDO/qKHrg8iev8G8Rcy2X4R7ncTmqLtFiGYOrpBelcG1cGrMTtOSV7ArxEg7r2Hrw
LPogVkckDYjppb6GTEUDmi39ePDVkyTttevuD6YjPXZmoXpSwE+mCNI8eH6CbnLNW/6ZNB8ErgSe
ezmemud52/MGvR72ZjVoqK4sEqVA6OK85I+Swpu8OygqIbcm/EPH0eyhoBbcQ8c2lQHeDz+urkAD
QnrAPviTGpu4n0YOP6SRmIQWJVYbz9FzRJfAQiMlizagEy+VfG5iHhb9mGFgyy4ibeMiHDN/WUWF
d8IY6n1cSGINP10VBdQl/6zWKF56DPpGqWpN5nHvGyvUqUIggcEIs9hQOmjTD8Iu550R3A8xuII+
UNsLOCn5m0wtchgIfwDPMsoPdDwBMjAYS17S+sCfkp3KZ9ghn4uxbZgg82AD21fWS9zNCiri2ZKx
j00DOQ7j4jk5tWs0edGfO5SYMtJp0b3NEY7VA1hvt849U15dUnNQ8CGjxvo2KneLTsqXWVwgLp7r
Cd8IOcADPujCyBuygtRBNAhsSy3DNoZqsrIMziUkuFbNtxHYyP++8iADRJvojBLu67d0ZvotM8Vv
UeJl5QsPxANqfAfraLrL3AiEb7cRHUt7vYX/6Qn0MkDP7QfO3zxkVziJz16CuuKQJpK5avVeBfAR
THM76zdLDTsY4UV4SbO4jTSKJ4ZCn+Ys35F9TZvml2WIyopbNuD17IkczHjd75lab9v9gGKEDBmr
pUIQk1AddUZ8azTZ2ph+yXtK+NQDF7ZAwZvec1SJoPJZw84oia4Dr96xY5mhVOdSkfmd7w/YK/lr
+/F3flTeidFYUsQ7E9RYESKyBnCx5Fs8mQSFPoDljQdcGd4XO8qFneiobkH26YLcO8jmib88rHEr
e1XG/GQyKEuh9rtw8CAyANY0sdGub4stsYuIs5R+aiIIhgFAo15BuHS9izBcM8WGPQVx1rlb3Wf8
dKut9tOV596rFaWli5HKktUz5pC4X/6lIeH+6cLB1+sQ6lPtMAM1B7Vr5dhxvOCAlzJX3Pjlnh8F
6Gj0xRaXcC95qMuJMcF197x3wZfAHKmNCcx9BYN6zFCLdrVNl7P3Wy/5VvxWqkOWlFaEAFGUcd9C
wraFLFmJmhiaQdAti2rgVX8nuWkVFJXD/+w1fcreDhcZgMUI05qc6BvCX7g5Fq55t98da1B6uQTL
OQDkdQZi+autrLF9woVE9YEWZlLLY7If8arW3c7MBtMl7/I8PnIujYfs74CtoSar9Qb9Njeb/Taw
H+kclSwzHlZguRGKeYUuWsCjdThwyWdXNP4d5xySaD83rrizLbl/8Ugis4v/08BPThD0CNRNenh9
J5fQdLMEMv/hic1qFpnrvYSkSG5liRHT2Ix83DvHm0h6IVhZq3UM0Uu57cxgi5pzzv3/Z8EEjiGF
LlnJqh5qYFfSV6RtB7iZvd0YLHKXPVP9CAp7KSTiyccVwvgIL9ZlPr5jTnLbibRvQTChj093VgmF
3SYY56pDlFsA2jqKBsgKGtIwjQk/Lmkitt8/O7QDzYKoyMeHs3jcKmqzubKbnvdshRfrE7He9eot
/5Kk/FV7aFaQkYRP/u4fio7HrLmXhV5CAjZaBU06k62bbvzKKbf+PFKT2wnczXHbBWxg3aGUn0oL
V1l+9LvvenCBLv0MsIsTCt2cF9cXO4JqLiRsWxzQnA+p4naruf+rLDWzrtV+c0rJqQpcMUwOqa4T
lSAuvDaPzIAYlGGMDE528K9DMB8YXNMwy0XBE9hyPw3WYOqRQU/8fExo6mawjZOtBdal2UTMXsAx
SvFhOZ3fy2kkF8iMrV0HhwU3guFFU1lKREDlLvQF+H4BrMM50nkMHwsqw904cOtnNAOW/4//0pCs
TihN/y4UW1U62su5mV2sREozKZ8UBrvHiRT12hDdphoNsvu1Il6ZnOSpysvebYnXmcRJr6oPnBxs
t2Yewqpvq54Uwlv2elJBroZxvJk8ywsGB4or58fICb6uagIwq7aBchZMv/jN9464y14dcRCFzNyb
xqSqEndYX0EdHKuknDbLIp81ccxLsisf2uq0skZot9I/g3kiJ1MLOi2k+XzVtuUXKw4nlx7Woeo7
Jf+tkx3Azf0IYvUZ/2GvhB0378eMONMG2XXWac2rOZBim+iqetCS+bn3jutwUbxE1aBQUiez2DQp
KZbQWejzkJF1IxeEAg0ZUPRDz9p5jxg6Euii2hXue7M4493GrZxsMG3rRkrNXMHaTQzfalnaFh7A
vGkRUvKUvc/oFrnNIJVrC/4HwHbh++Q1X4SBISYi9LTkFw13oLlFmj3OzsBjpL9qBjxERKOkv+8S
0TBEZ/ZHXa4cjQLEC4GC61wEComm1LkpmKCLI9F7REbGZiS5jNOQ9cV/3RYLHJgWC/lWBZV8CgNA
o/nrUcTNYtMKhos0q1Wx5ASupxznF8ODCzczqUz30vDaEY3rMJWPGijDdq68EUxU62esMFIqjK75
fphAVZnf4Wj/CG9MXIV9Wsnkrg3Qc1UROZ5g8GbDzYsHSBLzTjQKyM/YOtuz3IU1Al44cyI86Xfu
9tDxpywHAjyxXbwmhiyKYHNKTa35R2nECVB3pjAkm+mjNRRnYK6Qwxl9BswusoVxvOXKaIqKuVLc
tNxYKNy1xNyUX6CW6uTLAQ/ritZu9BoWDcwtaOzEKOFMMIdKRj3V5wGVUoyyEf/Qg0ii3WVYDf2o
QaGDZD4bACOxBQsryss4J6/FII49uhSVamv2gJJlAo3sTU0UaMp3bZNnN+JkOi7+1rwrssCH87zr
W5BsOeX0INj3Jd21fLC90631UX/MuoaLSXjDkYo98waFCTevwI3cqQHEGbsNHti8ZVsVdvgFRJgz
01+ZRhJoqb/eWxYItKwVFqbScjWVaLHVOt4xi2TufqFTOqVbmxhoYkifKMJ32TyyfO/E1XRYAg4+
JIPfIx+9jUbZMYYPHYHfGpbGl+KqdIdjxHdFu3KP6E452jpMTPLtJWTswekl/GUle6LXr7MtsEv+
IhHJHtVySb7KgdkrYq0chW7/jAh1hEC9eWgS4Mdwdc3ftHRsQr6xcu9CTUBYG2LeA8hlWnB9QyFF
kqt6xPoq8Td/T49km0UUEpeNIpwQ0WtUtTVCU2Z9uFOhyqaRXeTmQrVfGx333zTFmz6bU1AonfNp
zhaVe4IT4F3xVLkzX4Nb1FVrZN15BXrlHCvG3kYW4PGoc7tSPhbnZfDLMiE/0gwHWkqFjt8XNQup
hkAV6fSrd2dVDWBOW51u+ld7YrDWwmhQXJO+llBqfX6E+N5y8IchqE+kaP/A22ZSfasHb+uiOonZ
yJdJOlgFIROnYBFIK/9KcBOkepc6cNmwY4ZNAsX/lAkE+RhQPNyez5/VfgZxAaAexHbGqgmAR2mb
iaOmsFO5MW5s1jlLCZL9eZZdl2+2EiKPOd/fYjXpWgipY+9kPF7UciBsGdXZYb+l197AYrnU15tx
+MgaGZGLSaK9SGX/+JfEzwV0tvUkEG4UWIHfmUebxU4x+WyM1k7NzZ7/DFBIX5pegNoOvO+qZQYs
mOMV3Jx6Hue9orooM+wsk/sBRJbJIrmV/izCMMktmTRWPiOtvZ6cUqN7H0t8ltbRU4M+PhLM7aq2
nS0g99lHgQQUaoX3oy6JYElX5nFeFB50nsJTv1JkJekk8BtA2fd3JAMt/XvTGjaqcK4cli5LQz3g
1eDJ67nTBQBabgg6RaVud2Foxxk2DjLJ3BIh0x3Q/aRxLt3BELAvHOpwOkmDyDnvkgs7A6avdeL5
ZniprciLxPyy90YTHi570DsRS4gU+06oYW1ATObtWO9xqxkJp11aRxr45RyNFjJxtItX/jMxWuqd
2ShWpRlM2CYd+P/lfDP9E+rM4XqKZbHMh0YrTcenH7pia1yNvSdTKVGf5WhL6bJYREFAHXNuzTDQ
S8WkvU0iegztFDX8WsBzHbQWB6Wrf0kYDPa6jtrdaSJPTD818Cv/AM+/yREifj0ZqV1GMcCd9xr3
jWS5bcohDwmvS59rUTWyuyYqjUHFWwp4e9BMRnRdIaGU3mqYda+qs8nvsJ1VTn03p7J7GIJWniRO
vf7LY0CLTEEwLQhxGuVO3/iSruYY3ufkOXXC0oxbYoi+gmgJKYvaP33MTmm+yB5LjB11rjtP0zrc
Qe4c8CIyCQeT0JW5+oZy7yswdKw+UW8KsLLtA1Csa3xC47j1zAxJq05AFpxzdj4PWE0ePmN21NnE
lW3rcej/AwANwLa/MsAP0GiLTgXh7HJcL+JniEIQKBfP+SFAfa52ZdBGoUBemKKCxizZbP260V6j
BrJCh3bG3N0ffcOzT14QiNYUsJhpSTQr5iKA7iIQipzPR9I9u4Pfa31pgJFc8uD1uIA/XcZCI9Xk
8hYPEXigMCkc7cmi6w/A9mxm3t8wZe2IUl+tB5PXhVCRTl/MEpvA0khCiWsZqmQKQy8yR/KuRTl2
fjXQuPNxcF/TxT4jmxXNh8sUGR9qAoNXwEfFNCLkpNcFyrdabHvoO5lyLn3W1IClnekSWy6oEYMM
nWmFBLexUmUOp3ooVm0XeEtWAWxS8MtyiFKv0pLbGQ2kJOTXsukhBrdSUUQ/+aS8FJOWCZr5SK5X
LPfFbpfw1hvcyMkvzHTG4gVOWPweakfHZRTU88tLVENkc1r+jEssL5xptaYGlbQY7nEkkYQYdnXe
3rJeWeCRQMS/zRv1jvgAJE4PDTDBDl18VJ+AZ7UXuk92vW6Lp2tkicCENK3eFib8onZUjEX/luft
IzGYsK7YM8D8tegn8SLMNKu+5Z4JZ8YpH43QBvexrzsAdGRDU9LroX7hQsPxh/FTXNTCQUcsRc2g
A7/S42Xfyqm6EjzXpFeQQh4+aUc2aFkvMQMcYriVZL6V3xW8M9gczfsHwa8wyetlZKRsu99I75lf
5U7Mdne/rD2UOWQqTGzLUurRIUd+g3ZpaAYGh8CkdL1SYQlrFnTcOveMe15U/f+5lwPe4aG2KoYl
1UDbCUEg8d6SThGKRA2hOREr22jB9lQKAcBH3cVRGUEs9f0mdoFw82m/wi9YhBhfEWBT+XwWPDs6
Eus3tfPQzelEHsxOi/cWbrg33iQfHHiX/bs+JeRu0fsOuSfwcB0cNpI8WHdeP4bTP83gUbI0ROMa
8vx+eECSULdgO140xFdj0x/CbIjYo8w1HphJ+6u7P0iaoL4CU2dfwj/ISZHLIyxKP3NPG//RDFdr
IVUoHiycraoV8udN1SLtIce0IS+cKeN7j2vzjSg0nPbIGzg7g9BI17TnanKAP0pVRAyrW6BGew/N
mZ+Syu7/uXERBV9XdPgfahaCPCQ69LwFRNdp+j+cyH+BQvisSF/A5RiolN+baT4E3cDAyspMmhWJ
+X+7oXKpCF3P74myI5yhuxdFy6i6e5tqnaEewo+s6k4R6+jPHlTIKhCMmo6GjHed2YEvQIra1xD9
7bNPuNRZC493B/Lj83gtekwiftTbp+59TU/W63CyDQw9+dhG5vnsMzk0vSLTymrbuzoiG0jg6ihZ
ZhUWJhl+uHOqeWpFFY75yULR7c1muvV4gmqo5SG/PiNBHEtei+ZsUFxHg3+w66au3zvYnK3lCyv8
EbdvYe1H7jdttCsFykOOBSnxwX4nB/gxk9PRVS3XnfG/3ph7OB2Kkp3ZpIo8Eb5Br/fJnkw0YWEL
CIFQ6xJiTS57M4TQ96yL/HCTMu4fKTAzVwwC/AighVfjaM8AqNM2c7SS4GSY2j0j0cFTmBvv3+1Y
l2LM0+R/eBej8RtQr2m3hLHs3QMGAmHOWQVuOM/evIUwlLktfoWDQ2u/eOBPgGqmBSqLhySkG8Sj
v4P78WmLq9/TfBoJWFQUo6bcLo7UqlQm2BvGGgIT64RR75SA1Ab5qTG+IjJke+03ETdyTvfJP+Ka
sy5aGdEG8jR1GmUZdHSHgrg+WOqN8gjW8iXGX4GKpF++EmeMW79wnk0buEhVZw27AKsSNuTDrIeG
rUsFNa58pTGXKQ3L66LsFAdE2bt6wD4w3PR72UEBBGYZuU0SJCLZVqAasD3Gf/gg/s1sJzFn6np7
NV3KVB7ztcKwCXqcRYWhmLkptQ0fg8C1toAJwGIawgMz6tz15sgAxwJX1thTDdSphxrqYg+c3aMW
K3QxMlK6WxvmE5RogdnoaEPePioeRgrnYWAQzAFIZgl11Pf2K2y0GDAxkZp54qPy7PhNt0WkzUJP
ga9fsP/QrobYRJlzWVkVornOE80M0REXHAOQ4frMexKehV93zJzp4CCDh/+JH+lSa7ueonMqNBp6
a/RjtknAQbmz8BCicHNS54lsKkIc+Jw+YmSHMVKLp/tQV7oC5EXRinu5k9M8mGDzK5QK5HvpvoVk
SScDsYCI9noNBy+j9BbIMPGTyhTyhXxNpgNHRCsEMxU9GlFU1YagHX1+VF3X8PXox4S9XmXWxMyJ
ZBTvaDsTMuLsOVXjr1nAfVERsobo8AlM5weu70zOB8CNDSyLxxKJsbHCWQQtgA0UThAIHI+LDd3S
Mx2Lca5sEXgMiMsuuj/MWzHg++Xecrrjr22EGUwrJlRKCrp8DGfr22Far5EEzWNqqekOwIYF/bPi
fjGsVXHWhIhfMlLGCrFTLRrYd5GAWVx2iN2dWOMsg1MyvU+8WJc7siP1+CgcEooHGwruIPuYRPp5
e2DgXxiV+t/XaLE+yK/eY6gH9LM2wEiqoyyEnXOcRcl46+b6Xm74sQiCBfG8Hq4NvPXh+mFhE2cT
opEA5SMn9uxJtnzuNYGKa+MI1jRUYkeMU7/rNNeu0jG7jKsVTvEZ+HYGpIlY87nhmtKhcdLIH6Uj
Em1IX430FenAk41iT8xr6+TCvSiyqrjOcmaEV5NbyTJNdLCgo80Lw/F0JdbCrKG1oJeKC7KlrtoK
eIEKfORP0YfIhYB5JCJRwuE+1+8H+gogb099OsQrdYduVwO8SVjt3DIf6qM1NPOb/6RW0OO5I14p
V8Lf85M4WTWIYjflD9s2nFlM1DhkN1xm+od6IiIVNAbWCdD6rgouJelkth9aIrVld5mx4beRlVOY
h2dHrr2W+WTGFcfvfuzYcyer6AOFfj/6B0RYB/oqDvllnglbrxdK9BE3+xQiUt9kF3XcMVlUnJB2
+vpsiaF7OASKvYh0M5KpWZTFnwsIqZN0BqZnf4/RlY4xVdQp44LGMD4fRdsklAFqVK81wkt6Q0pX
kwNXoFBki9mS0ZGMNPtum8mpLLQZIesn+KU7WJ6I9rat8NM8Nvahu+6+rEZLHeiGbqpDOYT4alFH
JHlcAZGU6varBNBgX7awMuNDkacLtm20c/gmvrcE8JtRqRw+GbPQgCONslF9x9Pu2FTEainkbHX8
fDqL1bz8z04nGMxECoi9NDKlrVnWbxCY7psnRvW9NVViuso/GnmYtWycdcF/NGEfnu90OcnkZ9Dg
ThzJa1BxXvxWHtaySlI1MMZGNXyQXaEXHM/gPzBO+R1dW4QEe2p80kSjhlOKBLeHYYMRBTT/m6yM
Uk8v/hjxxN8qWeiXAK9RLakHM9O9zQWtUbwOB+l/RZUkJQ0KRUYRM+/DG/axNRwY0RYDkdIR/56g
x6/VbfDZbWM//fzgUaLiqjR5DInDsS1KKldRtudk/FHZvKMZ79X/tHUizbRrodVuLYxCnRV2KKlK
ixLSivjyLV5Km4xrPoGJFeQYQzfI0v1+NM+rNNNfKhHd32BwHQy/EKKNnUIcq0hMNr9EFzx6qm8f
i8MP+HK5e9gstAC/Y/ab5yj337UWy7rVzAWCYfWbJtUce9EYxpK4UXdTs11EQR+wsmZ/1CZeMJeM
9YhxyRT68uAmeNoRYZHXy2ZPeDa/XztE3XkhXVqeop5umdyxyvRNPrgsv4BWTVV9aAXEixN0ekoE
/lENZdEpAF31purdAmE/pY/K+fLTBA5Y0t1G+U35meUW4d32alwdbLP1ApliOqHNDKdVV952Xp/i
6YAlV6n3HGGzTa1r3xuFtZTiaPAEBUlwEc+WMI95fnQefKdowb92Sq70VfwZUyZyRt1krCyN9HOi
p/24YsOeDgarAp5Fc0UqDh07W6srNfbP3Tfip/5jZ3ZqzD8Xs97C34UGK9RA59kw7jJ7xPLPwFFE
qd+m5KVZsDbV8AdYWRLo9amfxhtG5m2wGt9UAVBRLnNytalDMm2lbRQjnXVk1FiIpP4s7eaaEY4z
Dzca4BjcowUV26kHaEG24mwg3TMfhOSMMatYhEn9gr6fu9mKkmJFNMuEKOy9VuIPst0o6jiF8TBm
FFmwraSn2glUikDSPZHaFUjOtVQzDyeZd2a330XuniNL5lHTFSJr3dJB6873PGpoDBssgngnzBW8
SBcyMOtEgjR+EZdmScaqE8d1yWaNGwzCDAfIauI7yf7Jh6FBvWiZdZbLsVqEX2gzxKvvqMVxR4dW
JpX4Ks7FINbF9YicxRxVmRnVsr/Js3R5C7H/ZFZ4VXl3gAseu6o9xKGInX6SpD2IEbnGFHKFed0q
KM50VWWcRt/FRCbEbLNiB45QRhAlK3Fx6R131gX5vngwjpr2131Qkrsx93PpXPsusB+8h/0llZW5
eNI0SPa7sTozZwMFSRR+x+CnmFrtHEAuC7PgyhwbhglfxMESgqlBE0CPbBweCFfbbomPpZruZV/I
Pw01vUrrNwE12HyfDDcWWsBJnte4VDA+utEJ+y7o+7ot0Ejn/uspf8cBWuzuRqZ/hSvkii5PDTGa
4ODTeBiRZi+pGQrKU2Rz1l/HWqGE5pKZt1oxfJFNl996BM69iNYySega+TojBuECXfplLLlD9v09
CwC2UUKuyICT/C/+5hGDUPhDsfqbOOhlF/O0yYepQ8WwfxW5as47xAY0VCzliFYU82yAwTLg7Efj
mob3f0uq2jsvbsHEH+zS2OZMQzs9jc2TwwqKuullwh0L0/Obxk1wxmDmId1INCjY3bBXz8czBRVG
I2caF/Vr/wQXQ+rMpnupQyymxUYjnN02cXeFTyqMdVLL0nBL0Tat24MmEqPtQrQzGq47UbU1zmh7
Uwv71F/Tc7mP36MInFxk2NEvnQMRNNg7cprK2EhyBBdjBrBQFIsN1VN2zmEqTIWkUlhINoiFtPUx
3XYx1yKUhcA8gKKfFWDp3H9Ax/1D8hX44T6PAHi0Qo+5Umjynp2PslcA8oLBaR44yXufAeM5wzkz
agCVo1MGVKrp16aZNtpb6tuF/7Kfh/t9RoqXi7A+ZZ3qTHRwcp4fnqmNXV1oE5lmIyz0RFPEbVT1
8hPFUv5uqgKr0Lj15nfGQBidjyOyITdyoyCuzEQO8uY7P78M3zkLbw7CAR7Xre6b2l15R5vDgkfd
nOsOla/Dsll3U9tg93/JMM8UztDVD9L2Cs+yabsER9KNeI2v16P/Kr//5ge9vn8vBXOBaDfF1oM0
NoHO2kvpvsUTB53lLWCZnygxjdQzN27B8U2W0eo6SBiOVa6IBFbhH8h6kTg6MDv9H/+oX2g0PVMV
/u8WiQShzcknXpyiEg3S16lQBam/s3qv82TLOPgcQjz4gdRWYHL/MbDuS43LjP00pjFEwL6PBS3E
W4Z9Nwq2T4fv1cWtVrAOYia2uRvpr8XcfAAKva3u6R1beK6X4IGKVPOEeuPyGl9xtKCNcpkaUdX9
/Kn0l/ODR/juyZ76wNmYFytYF45QHO3bV5w/1A78aoS0bhpZSZ4Gv/puKteDrcOntfz2ihJCrUoi
nM7PqTeqSTdBR9BprAAAmmmLFITlpIELlvhT0yX8rB7DAw8iX33oixWGWfHvRleWB9nEYDwR7GpN
kjgPjzaQMzYu0AVg0I3/jmvmq1zGmTErefIUaF9oV47E5fiiGKvexaFdEC1XmfzaqCyYEmAkry5l
ZV//Zm5PCGabLEXTMhILcaBbssqvCiv710PH+Mou1KvLI3J7CpfrMYtzTY1/uJeJ4hOFt6LXPTtw
qg7r/9zezFsYVtao3JrSNXIWo1PkAerxr26ub8ghDxyQumWzM7yUw2Ovu3STpWeljISX/VNZ1PMD
DPtk4syDXrExZTCTgOHGkLXScxLw9AM7Ur2U1GlKwpXe6PPvI+eifWlLWqZyo/JAy8/2iizT0LG7
jLJWG9yvQ5EFcCaiTDNJqhu5ztiWgZRFob8zct8qUy50TLxCMB8Dvnejk9sECW9mLDEUZwr1zHGg
RSCJf/AQKImpR7EqGuTvD0CAPT/3quSc+cca/9RPh1VvQ0sasSZe/X6T13RMSHUtinNDcO6n3d3W
WJNF7D0tey4wgB2nQ1a58oLH/6FcZBn4p5WDiMHC9u0RGYxeG4ETTqMVU27ahEqFcSZvSDjdLT5I
vhNXPpCgBCu/tDb8iLVKhdFseNQxA2sBkeoGXeqRguI5Wb3keDd5kd70hcqwjGbJ/ANg4JuN0Vhi
dp4BlBrwvd+nX4cAeDdNYrk6mTxtOfUKelyu8WkDU2I/lwzZnfnxAiPuKZqP1166nLkavcoXvplE
oBOWt0eGsOoT1VIy6iOHQIe+PMljtwy4EOvBSsha5S7AmY7kNOdaZLg2klkN77teYG707aPtqE5z
EKdwKk7ZAiZPjDnT1gl3rB3EpQXOJNp0lu0oJtajprK12Am8iAgDIdc+ZDsuRFrvg62iLCvoqL+v
RQuf64+3OdK7gjyR+r6tBOiv/YKXuCmCDvOuHfc17+8Uq3Eq0R+IPSxfJxoGvyRtp8MCxkOOVn3f
N3hXrPBTeWs2vfLbJwDu90vLwuAIQS6j0sdY9c3GFIbt9Bar1lNeAflEUH1knFDox6ZoxybA51yy
tq8Q44t0vfUEgNXrgMocy0WSiDLDwom7OolX8iTaOlXd9rHAlGRcl6EBTGazuAjM07Xbmyh1hoct
6AX/4tazLXP8+O9ABOrbRuoq9XfEo28anVaHdZgXvJH6tw+KQ2A/Zy6D+7oXGaxmimiWCgRPMT0c
y84pWBv6ZxbupLRxqpPs55HLZDvXJCE9oMgy2+qi1uyeUGSdV90KeAPc7h3KN6hOgBCihx5gWVGz
QkjDO/3Z6Ax+f1+0pWVRakMAUsIr0ZYfBiGdl6rQIEiqBh2JpgfBt1cMWWAALZEE7C256skI47T9
sujrMbNXrdgMVersTSRlkGlV+bNAJbMbKWp2AmOQsNeawFUjkc2rk/22D/AxU4Bu8WhUs0yNEpWj
SaNAsHFvDSbduy/RNC8oRkx3lruV75bIejoAlQpk7XG/7XWBogxGHguhB7qHWgQBawIWY4QLFLW1
24x9wafW3pqndQXVjLDvnsNq1+8EVrf2QCiUsgXeUfZ5dbrath7lanFeleYhFAp4SdMTok1kgcyt
NJP9eI8kSEPpp0InuwTxBxV0aAzHT3WYMEZmexTf9gff/INRwQJXqCPxGg2/bVoZxTvq0NU84cPE
RpXzZGILvF50dvjb1fJVsO1nxv5JpSPWskSmSDjLeEOfWgnwug01lyGi7TMxZH9XAt2zA7wSoC1G
RzHWzktY3RfcWRwX7I2Y0N2H6J0QQxx3k7CgC2NhhmJmp4g0GUweqRp9UnJuj42fIuc70AMOcFL+
NqAjmZHPlXAd1ewEteQfJVxzCxNVEkEJt3M3LuFon1gZTs5yFvqjNq2Fas9+5gbj+XuHo4YI2MFa
FwCc4wN28W5TUn9+cresfomXBL88tMjRPcOfGN7+AF1kn/siFo2uHa2/VHRKvU+rLJnu9l/j/+iB
lvIU5wIHnFtbsEDTzE0NWTm7GToU21x8fBq6e77bdhNO00sxXsLYPs2wj4LYz3pAZOuxmAQ7I6zC
URBwFjYJ6eCmSlufzT5wpHpCadpV2ZjgPRdFiJUlZV1W2qcVsbgD18UyVgX3MxrA+MpCE94M6jE4
9OK/FLve5K8bQ/N82iXUsSjk1rdQ4evim8YLN21U/Eiaxrvk5vVEp6+fs7xj++j2MAzrgRWupnRE
KhsnUevDQWEImMaCFdK9v1abiu5pm6UGd+RwNravTQAEmIjQMmGE7eeVHCLWsJIoEWqxVvlAUOh+
BCXKvaN3u4hMsAV65sgw9jBH0oZsxXWnzmuYnXT/p3iSr2u+ehkHMRiri6UA0C3ov2Z43nOKLcy6
6iyD5EouZsdptfgkLechBuRW46q+D7lUHB6rJbsr1ZkKGHLk0lwcG5MQU9/jWhsoeMh7gqRFV0fT
tbi4KxO8sXi3o78i7Etu6Kmq7tIeI7TOgl2+B3fV6N5V6B6FTAASeHbaiy/ZuDkY3ESAsaQYb9nZ
etb4YhdgWiaMV0vxjXgivYrjUUaWatlLOozJeMZdzLHKP3+sE0EW0JLNeBIBwvxJJ4mnDWnV1N+I
/hX/6Faz58HsFQFQCNmpioAb0hfKkthFeatjXVhnCTU38tbbnE2UDSesY7QeUZxK9T6aiIyhRiNp
FABikeGuJEK1fJo3bALPHTZJBwTvzKHIZHGxXdBtcFDjJF+JEi+10tW95f5o2jSugv+gRAkF31Sj
VN3u+vGEohgIO1KwQmL99nrZjeB/yKIz/x1D6JqoEU3RyVpRP6FVEEArZhiu5VBVUtLAp6lex3At
0opAjvOcvAQkU/12oCz5onl3njIdj0j562W326vHSAgUEQF/X5IQrTCW7l+GDtZ6/CU+8UHlM3XU
QH2U7m6SX9uou9nfjeDYhpnis/HAhF4TYRDCJfqaqnreehEpuuoP1GjwLhbhdTt0K/OAR/IOr2ei
zw66CnGa7wdMGOdjrmVlUMlENQ+gBSVIbpvbnoBiOVTsFlKZSLhjchuXtWQcF1p9m6cikfmi7KiE
kqftNCCkCDPdzCaaqE9ec/LRZX8dEwG5tmR8uFO/tHc3tPJTMVqSAmN4WmJAAAiVgw/HWblq3Dig
FliYDgu34TQlAulyA4GnTZ1cJvPijNia2qwOLwnwRE/fZh35qZAREltDhjGqomIk0xujiZYKnG8h
yR3nR6YLYg3KCqebJkxb955Vths22jcEIq37cEyt6fNBBy+82ToaPv1ciaLFhdZzz2SQwdzcYtIu
XXUzoZI/pmz9GslJ4HpsiuhPlO4CV86jJB42ArkTjdgqgmAAMYfoRgNaHAshP/9ij8gbXqEPRdKI
pqLCxyOoehqYVQ5MsYd1CHDqt2lGDUz0V9TdYhv5DHVs6jpIEB4Tr2wBPQ1FFHiD30HHZEHQFa9z
mkllOlkHIrstsoMmbMWInll1xJOvXFWRAcF7p8na/RhVI00UL6pQq2OSZcCRz0lSxH5A8eZUeK/6
Fa2WRb6ROmrFasonK1UXieLvEMxI6IRQeT47hUAZQlOuqbYTGOKdp4iHqKfo9stZHbpzFwWQ6JOd
LduPPw6aTG2BA+5ee8MwIVsckjdN05rUGGo+vVl/p2b650AXcm7Z7OhZIClJpwqtzm0oIp+eUlt9
j3Ly4FbKBABcyksnvdmdwnPLS7Y9YNceelrVnF70u6KEvaPCcF9KeIt5xgicjmgOd9I9j9HKQgIP
MOLqdHTOtA7nkvq4rodRtfDBJwWiztDdrXALt0a9u5CDlOho5tuiuFASKsdrCwdHywMsW6hQ3zzk
HLlhKqtHf16GwH/5d4+GeerT9UpQ1PZN0blWxZrgaMjWT3j8Te87N/weESy5+D0GImZUvEvzZ2DT
VvQZo+fTQXJWsTdckamWjSXx+Om7sh/E/Snn959Dn0/Ani61D4SVVjoEVIVXUrTSSMFCDH+uyiS9
39jLncuPRAiq6FSTlrVgof6qW0iGVA/1JG7ljJjeldh4EBViCmcIT+pJcF2JO3QvkaNRX6v7f8JE
E0YGdRgo5HRAmoPSCh7uWEoXXOTy6WN+haBIn66Hw388IR8hiYjIMXqyopXe7sx6tOKIOfCakIHu
OWM4tW+gz5WY2i0edLRih2zpQlwmxpQN7479RbjxQWMa6lxnOgo3uO5VA035dAi3ya/U7LeAIe5/
wkQuJxW4tMFT7d+dHEugYBUiHhPmWXcwW+Utzwh9A/DB92/FEtbtTzAZWI063XTxjT7xfTQJzSjV
v9UZSkkoywjZI8VUVeKFzP8dy93fN6/AnZlqXKNY7wcWADtMJoAA0lAJGF0rj35GwKVQmQeUOvR9
msZ8dOX15rMOv/X8ZTkfM1ABdJcUd/O1OkgWFbEZDHrZ6M6aXAe+KqK6f29KpIpofuH7pDx7t4yb
wwxyDAF+xDNPjXdi2qm5SJxm36sVXEmNKdH9UVe7lOGYSdmscNAHdvD7Qqzzzlx4UCHP6cCNRAr8
cfv+aEGVkHhzHeSm2j6tseE4n2B7UpK1OsLBxiubcCi7K17/eCBSOdNenmkf1RJOPGK1+wLrVRvr
rt8kHTqBuhW+vKgvT3AlBaEXoWeeTu0lzvGm4TsAsoIsxDYB1Z1f/mQeIHEsqVjgpYQQvnu6/x3z
vZ6c84ve1rkX/rieMvHYMmMR7GPFdoyxEPN35NqCdX51XUSLa03NlMGGwuMu5uFgoNHk/bhd5UAD
eLVAGSZYy5RG1ABM7CfpzNerp/yVa4Zo834N7yNsZ5pYCqDT2TL/sMZgz5opImQBMGThsAh+ke3u
HL+UOMWkn8b0z8VdOCd7dbkHzJy5bU9wO01SW86uKcViM/UeSlzKd9Cy6ZtaaQofZ5CK/NW8sxdm
zRczH0OCK5guduQHvDTWZJTDS1WStOzhwtVGH7jWIfuBNMbQrduZnEEckEFQNF6yiWQ61KIx8fN2
leT/FGwSENghg0fj0G5wZ5Np5CRZteDqrLpVl83biistwa0GwoQFYJDxYWP42K688uUVSRlBUMl4
GjKF/4nrxWckYuNbjYtgOnhm0TfYDx5IjwB/4PZYIriGoIyIRbTZtEovkx5eC25cO7Fe6hW3ozYA
G8naZBPEXPfhv+veIFOcEE22Eptqtc0uAoBOTBWl85EcWhBwzt9jdNajk3VvakZRQ6fZkghiP3SL
LtlCfGJGNYnxT9B0qNmaptRVsEycay3UPl67zRevK5cWz4SnsyYnyqp/KkfboxuRpiFjnFOkiSFK
Gw8mh0r9CVXsr6w9AOpMeuAj3We7hUNUunupZ6WueWVXidV35XYtr4dzugStP1JLrhgsvXoUdp5V
g9Y32kxKvMjI5tQGCJKlfA5nG97l3I4i2bmfRlfUsyrFdEBbMcbhAKNxROz+Cmk7mLZS4Ta459ls
b4bYnImLTBNnoL27YPF2hkBs0/PLISu1i0Yr5vx8lMSkKo2/sTAo+1RQYDzAFVOs0i2N65r/6ucz
BzcyJOUo07/p+nPh4/Oyene2u3LT/JtnvxQqe0yHstGPbkfE9tnm1WT1ZHRgNFk7+dPluwe0FKf3
iBHiIJhIF1YMVBsl9hGr2VltksYZ5Jk3ZpWtxZVvdd3pq0ezLBrkeYgBDtLqdB3of92bv3HPkOCr
3O/JSRwJNBPg0sGcqHv+TheCgC1WYEv+rPKZ2h2ivlNWw3ZiENbfMQkJiQmt78ZN0HFu8rTzuYyu
HSb2LT6eByVAygGO7S1vQwMT7z6N7jwlhOhXv/hHVPXMRW93lln+NgyzvrufJ+Eu3bsHKE9YQuhU
zZSixe40fkqqM6btcefXE0OUtxZhi09ARGt/7I2aXy+XP8G2Zn5Jjfmhf6RdQVWAyhND+vOkSH5e
wEs3VEe6iwzF272lQQiD4cS4V+kGThGKxxgauAoMoMw4Zr2Opl4WywKEi0I0osTX9wUdILbQ72JI
q1rUOwAvqzca8z2qGAsbUcZTITZWCtopvt9ghNCUAURm0hl3PDzo0DcduSsSjbcHmjAG5LVNdZgw
8XWbeSG5EBGg/kEdc/vrZlUCaU42y4sD0Eg2eFGWMIPPWc8cozNPYpTZjGDntswtYxr+Bp6HYbYR
eV32Fbtb5HklW1R7+dO+4vs17Y474NDs0VJHNhMqtz5v4KN5mYQvFAp1nOI2wjmaSitdWzlT+sfH
xw473fFDbJW85JHUkGBYwgUYOczMNafNEpicfrdmb/duKmi9QQafRn6J27UcUBQIO9gFImWC7/iN
wwo0wgAxfd/YZuIyvatZLv//I1eAoUP+pQvbpkyEAYsnapghAx2g807qS05K63x9zGRjWWmq0M7K
Wovil2Jun8CxYkSZ+ycw8WeZ0wBUQ5Djcp60xfoaRIXiRJQByC1v4g+/wjJDbDRtzl0RStgiIK+m
opz2Kqx+FYEuukQXSKXV3gTqXtZUgzVCxGBo9SXWTDzT+tAWSaSXt+7RykBw/ugs96+UYzSdlaCs
ZsfytIIGcbb8u8Tfe2l0uNGAydpHYRYyofXlLX73QDVMSxH8okEAxRpYzly5lpYrSNm/dUQx1zbG
dZnkbXsMHdFMXaOLxXYVqy0lefe3k0Dm19TNS5QVpMJL/JsctRnEcIewTj3jrIq/vSv+q8Cn43Sw
nRHGKZNgLed0VwfHFbk6E/eWgNQ0XM/eUf5KHPZ6YMEQbWR6xdDF7yCGRAqRqxY6xsrvtzYZDa+s
6Uw7nsTvRmIb7Ln2qP6MAU8CubINkWqRHM8odxDbzGr1fP2qDDfS8i0Fp+l/U3oBnPPQrN+n191h
HEk9WjwFQoARyHz48SLT8Lv+tia5ljoH1iTLe/YH1+XVSavuRn+CHOoyIN3VUPtGHvP289y1gLq0
CuNWwCX/ytGA5b3mOn+E0miEozJTTkolyFfXt7KZM7sVvDMGcDbtfqr6OjsesJ3Vk65jycNL1zb9
GJ+Y00VY8DiewNLrTxwDDjW7hisLX+rFlogii/JwpQ827Ot+YPjWmEP2C/4aowCFqABfMZ0v0uZK
woS3n9PW9G77ViscwE+JbaBLM4kG+zTLJ/UqHprAbyu2k1con1hAMFWrakWai+sr2hVXyCou1LTG
BryO5OpZR559tktZoUb5ooM5bh8TLOzNttq+mh81pl5U1wG4DxRLeuR0xiu2KCsWwPzi4qT6Fbs/
tL2QKdSirTLJAUcl9PVYt0MiYHSufakLPQHDCNphC5IJCxJ36p1GEbpPgyrMC0J9D8v9ZYxHRbGw
46vMDorR5MfMPnHpP0n1RO9DFAy7X1Z+1cefqi2YLrLvnwRY5Svnx0EEhT+Bf5vh8Jt6Khjsv896
DVQi5F62C6pk1+MXvJGkKbXs3J0FGwCPO/LRf4e6d4o5xxp06til+B+5VgMcbD6BxRpvekPJb2LU
rOtkFgLRAkgsMnbAIBM5CSUGq/QvsmS46/G2J9EoipcxG9+vCB8OUxs49wdB1nA1caLxu1n5i0un
apssYtxUCqzNTXbTnHypAgsTzQFURZyfr2VhMum3HybxprUjdntCDTsK8urCr24FHCj4uHNq8Z0p
xh5q6h4oOTzyTEZNnvUb3RGvxMg2tdZDdj27g9RsrZpkvxQ26Qa2WMT431MhMGnxIyQhnCX7OIVs
FINbM455ncsbJtn1IFGj7uaLHG1RGJQdtcg1/UFMHrdFYyk7MDzAFCbE4RlTsvaTR27pyW9g2CCs
+4aTYZspeL2BsHv7sA85qZwqM4HdNk/hMXz/1dGfi2HKBtEZowHvBsypsmtwmLcRA9kxCl+Jpksl
IOQ7l7dWGcjoU3Y3YvJVMoS9Uhd9G9PqgfxkfIDB+yBH/v4T6yESB9X02BWUhrVgUC5J7Pq8eUBD
Skpq/O05wMAjV9ByEtVfSn3JvigHLXN3atQ7byJMCXvKteqRQMA22yzPyLxlWOc/IQuoBju/VVZd
VG+TcigYeFgU4McVhnh7ifNDlfZHclWaErKhI6GHk4sqJ3fi7Vew59DBObuwL1a+wK5OoRrH+nTI
MPWD/HkwQvUUhJnUfSlYLTn+sfq1M4SQPtmFlio8Iw4GQMEr1mZt1vS7vojHNfIPQ9tbKDNE566m
Tr7RsoDxDILu6btpVb13CgIYPkB6Q4758RTOzwl0//1dcCaGM98S/6IZjSFUCV2617R/rPz+7LTN
Ps7LXWKpCh+82j6p7uv8JlsYyy+8auidZKYA9fiifVZiMx+Mo6jiGaeG5X9nYRcJE0lRgKkouPhJ
Of/H9Ut+0w81qm0dVVIyp7TxrONik4f5F+xo+DtDJziTG9NR0AWPeSWxs59lj3DVxkeHq0SI9viM
M9RCdQ/+UNdodQRPZKmmx6VE82gsZ6rG/pU0pOj95RL370XXJGXzULDh/iSHc49N+3PCLDhAyJoZ
xK4Q3pIqczk0Uj3Amad8vYYSe3dr6O0Hz+OygQ1JQ6aAm+5+ZrrKkPtHKtVwhsSiyCzDuGsIWzGh
xkkK7EeLhI5pjpvXmVWJFU7NfeIjj4scqJ4NbYYaxeHvwyFRqPQkyTx+wToFNUW6NqtuhVVf7PZV
gx4KU23vEA5Ea23tnW/Vt9JLrUCy3krvbzISDk6YJST2NyMLqPeYhAYzmY6LrU7uV3aGnrXzKg3/
3flyDVQCpj+gi9bxVZlpeAoNx4T8oSSZBcekP0rGzERLx4rb/huyRAhDdNSe4TYGSJgQnu3Vlyz1
RP6bjVTH8kdd3vqexYR4UTGxGFgJJ97VffkdOv8fybqd1Jt65Lfkb4tG2bGbxsEJev1FH3vnxUGi
GNESxcjpB9OYhcwmBhwrPddF28LarV7wt04CUqpxn2L0AdGi7yTEZavJDC9zb/ywGuKrDaQ8BwwP
ubnrDFZXY/2gcW3YUUiKr2jr9+cbHXH6bLPRm6chrUAg5lOLnW4wZVwSt+hVTNQmLoun5URQhh/q
epiyfRHz50a4C8ok+w68VQrbRYTm+5ik2giXxiWOqb7B8up44D3u1tcaixvEabAgqACxLOhnbe21
7F+N+zWEpJ7kLj/j0MFDaGOH7yFwOhu05VvozyHyE3o2bzcqse1hZgdf/rRG5/66rGCdweqQ81/h
51daPtfhDtox0Gshlzk6bxG1fEbr028W0g1lhsO1fWx7pMpSGcz3apyrGXpf77lPWEmfY7OuOH09
uDEDS7t+n8YaWifxZ9G4Qo7qPVrpy244wYo1j4MOQjNF6A4W9CYod0vxtz9lhJEHudXm/1A9Vmzv
VGJjyA85XOF5Y5wWUSHN1lmVtHu1gFvJsj9XRKGevzYU1JW/j+uwkptjqHubigBQ6Nvg1fY6/oD8
QjqGxVIBRApHtLlrci4MLCA2XLIytmza3Fq3dM7sYL1IPw+mJeAvhtp3bk5tNdas5du1HuEq1i3B
o2falEXUx4qsaDCHeZwRVJ9572liwH40hIv0J7vEhNPGuMtyxpQm/zmBrOaJaAZSyB+dcZ9LJGcy
j/XJonjFqNINPaFpRAXjjLrm2IKDC4kVXw/PELio3qJh/aO2H1c9dYKhiX6kTw0/6H/qp4JIN8GE
lEnCdh95nfoVhYOhrvWdz35kSblHc/6YyDVELkHSCTglkyZeNhk9Umd6+yycN1D6gm9+Wbxl0MZ3
czuVR2EKeMeLzByITa2Htv5Y+oYwTGvH6H5yLWmrutR8YsTMmw6CKlYysEDz4q3M+vv65vWRoaaP
KKSUDl3n+nf1XK0PTjlmeOxu/Lx3RccU6Jjr8F0if6mAY70HyllZ71PEoUblE4H4VLiCYC1m8YPT
Bv9Mav0aLTjFsfDrQKa/gTls7uQNWLJlp8Bc/1Z1PQxFlologdLFJ8gxbIHLO7w/MTEI6c92qqB9
Ec1DW8mMHxG5iD1sgHEPme9RSqAQMZktD5ZaxD0pR9QwBGEZH/fOhoqZi1JDmTMTTle/mIRj4w+e
nh+6mlgnbzefTLRst4/r7LaotoZoF72vnYQ3a8NgONijd0CRKgrqKUpNZXEFGF0hQNObJqWAimau
RacsDffgcwkRLgdf4NmgF6WiBT2CzxCSqu8OhgjUytcIv/dGgfxdP5Wi24/PKd3BgeqcM8c5qVOe
lkiib8/bCSsilFaGk+gy90Ilhyd6z1djj60fXSJTKLfUHoND35uiiIQfrK7aKNQmyksMiYRHHKl5
hhD80UmVXrf3E+UdAofpyxrBwiQ0RE3ipoeGbbKgzfuC6Rltwbh7SIBziUQYOITJCTJtNxLfmNLn
00wHvg4puauhF4gQXcPA0Ktu4moamykLe7vH33SVutTBqVOaER1tBHoyU85t705C2BF0br62LSc1
tS5c3EdiLFHeZ0dYyXSybr6746aHjNgNXu+oJJQxZQw01eSMHxc/Ctt7hYiBCHtKThbP/n1Yw5XN
6aN3bUlvK5m7piKQDP2lppFbjQA7l8FTYIXzp5DIvAVVfTNpnexbxYouu651W8eE4ZlBq56RlNRO
xfc1/w60uFwe+lH3yKFLs2jVnwtAzu4PT34P6SguNZqssSdlMxRQQ/afeN4naXwcmp46Z861nE2Q
O8vEf3/otDSSF2k67JNQZCA672SeRW48/Lu/CjOR6oVAA7q5BJO8g3uIMwkzebdJ10FbEuiYFIjN
ifd4bUhDdVxxvNN9927FW0kVE99lk2XbSxkZMbd8T8sQwUqdOjB5/UjExq9gLz4YGcirf6clwPSN
V21113dwoStUijPW1Rtq8mTG3tD3t35kBuD2ggxmI9QLppLdnQJICJMoA+caeKecBeI8LdR8a/t6
JuCnKV3hI+DeTCnvuMovibIXBAtyBpME8jT/vJdNy8I3TgLC7qs8OwCGcu8ulhz8YRsP/9BJHEcG
p+HXoA3o3Q8nIVcMC0ptI4f3aO65tHMXTZPx+2f1MNrkQSklqQfSGMYkLAQrexCDFCa97v/LeAOU
0klNvXp95lSDApWEVizYk1tyhkcjtIVc2lKf9UCVCKjKso+FRJ7Ml2r6QRn0Mjc6S84GMS9Gy/ck
gxCSdpy2frHBy0MVz7Yg18zh/a6K48wC2MmNQbkddBRMbozUanHS2VRT5WSYjeEJdvx2xFgxCdMX
Rc1juQVteAu6OwNU6xUooMSbIIQZQsu3iFBsX6oP+1De7s3ugHFUny9cvwW1RmfAvXLHOBH5wNPH
8JmvTKOKA4VwdwV7tHTOkDx2gHWTcp5DCHPNwiGTJluTJ6X7PfijcmF8l3zkvKH6JRSHXgXG8+bv
ShlZb7h9fxtQ/s5YiwsLN6aOzfiz4JtWnevx61t9DAg+A39wcYg4La9pJHcakV09Iauy/uCGFDJ2
BZowBNbsuqnD4CxBvp3xqewl7WzdE8EDnL2zoh/KaEetRmeMDX+DZEEA4BHaJEKQsAGHj85a7Hh5
k/4SBlfHRuaFcECmmk8e10z7UvrV9EExR7YE0p25iYEd+I7uYlu/DNF+1YdUMAGqjq/7W/vEKb4P
L49lcbpA/rE2Lx0njp/MjrRF4YjERPMcfXIpR6sROVody8DCutchfjsBSXt+Rop7dYxLc3ycNhq7
OwW9+j/ctJB7gjSWZjqeAY6SB0E+Xe25OBdV4nOM1JkaCbvVi3n8Gn5aAitwUNgSJ6aqAO2gnNI8
1SKhNbzXCLbZjGF2+QIwT8LWCoHvJQ/iP0tR+X4ZTTazWX0O8Vi+5/jhwt5FniIOkgsWopf1qV55
hxUF1VJxaEGu0L+Lp1AUOhwIyvm21ZCr3wUd20aBtswSZmHUbO/yJc3R/iLX4heH96KeyhgXfzpe
AVIUUlFmZmR0RCsOMNGm71uUo8w9R9lfP58/8imXPM84aXdsy/HWt+1MG6xQyRHnyOLj0XVTVs2G
z6WFQjlCdAmP7YIVmNte6Qw6XDPkvIBn+Rs4/MAG+YROEE1H/zW/Zry7R/uyALQzIAPrEw1bEX6U
5Vb2D1ZS7SNBQtZH6tGsZuWX26Pt5TxsQj2WtHiRLGURfW2fr7zF7Ewa7l+5RtFehw/E+R2vkAeM
gR+rfL/aXtsAX4FCyqKxsGQgUwFg89cv34FvMcwuEgLs+mzGVr8A+oa79owv2wVmRW9kFVnkSwy6
J+Z2KQaT00mzDnr68KPzg8VW883Hcat3KsKfM8RB7yy+nQ2pfCp9TQ5MeXRcjr/PKkLib6nWEpCD
USUu5i9VW19cEVOAU6mKcocevwJdJX+WKajrjixmwvdY1apIjUlaw1AmqfuPqn0NMsF4R/V4UYYT
+prGGMk15HxNO0LVNR6AWj0QBOooQLf+hmuDgQ/XOAg0gLIivY5M+PQbXL72Gpj4lIZ1JqdeXxi1
eVb9rhmAjMgUTiBRQWwkvoxkpPDAkVShwKWpU61/KxDaOfnb2qCSTyaVSkbBNOQY4qVNBw4ZqMNp
svcjJikfkpwOpLCcJJ3weBrGH+Y729VLdQ+Bkv4u740Vl3MistKl7DV9zGcxJc3qnZ0DVzMnYCRX
aMHrnknhkgsywcyq61MU+0a6F1agzyN3HmKnc0YzIY1n7AeV53Th2adR/ZyUnt9ArJoFPiHsYqLe
+BoCjHLhDNzLdU89jdAzkezIQ7UGjkjJrqocbOcuaA5W4ZcabpWvQRKLdJ8xK8wxhgtl6zNjRiBy
wvPlkW7VlXBxJAqXcpH6NmiF2iv9UohwZSJCdqBYx7F0+dYcx6HuajZBRPtcFaCm95MJlUFkKhV2
hXNpFaHi568qk93+qSvgEAam82fA5eJeXQhLgtkNP7R4dAQZR/LHYkWnO3tRfpvWgCM0j/j6VN09
YMRu/t01aqXVkAfI1Z9oZ/4Rw5NfebForUvD44IVezEU888Bur6gHKXcAeF4/4F2oaIW4/BD9j/U
Nf8ywx05qVX0WoQHeA9X2hEbSRhmAEtYlBxUbt/168Ept6mQ0nYpAZMGoRaFfAZEOKm5Bce9q1rn
7A2CCPdfiDzmiDmmqkIME+n2EG8hxy5C56LdFZ9AaWCNVvLlutFuAqElbGIUCf5GuMoXrElu5LWJ
/shCT5gjxGWRNxz3E8KpGnf32MYlU6o9rMqdzQWA/0qviTCIdWkdEDbQ8edavt5BKnFY0LffhUY6
WBOWrOTw9cK9nF4EJh09Ghq8Md6q/5DeFcpHHGHJshC1jd9ACzl9T/jpFhWrb5Vewvfd5lQYdWio
1k/VoC6RWncFLNFd7VavJEePJVSWsZObUa1y7EduBBz6yT+mXsNTCTQ1MzYrsDZyOa9ZPiw5ko/l
Nl1lzLzn5F8Ohm06NcQ5ViYsZqRS8FQjekEwuN7cKCBRRPZlg96UkB3tzXNNTgzHeh4cWuHWmDAD
bJmRzmBm2SXItLXsq1560ppl1xpH5QYNdruIKDDBMz9TEX2+bbCzCEGa/agRNgS4pfKSBo05qFpp
6wVhwHuMvDQ5ylC6jomsI1hiyEdK4anY/bPR1XSHsTN0rMaBMGyMWKKPc0zov3QrX+OGg31csUYw
Xq+iV43s4YJyVtEcUx8KKzZeaLBplvdrJ/XqsyHjLpQLjCgXXZ9i09tI9ZnKUgkF9YEfMwo4BwMs
dAwbTQn/yXFjWUQn7+NndsQekI1RgTWjiCbfYBnLeUfsE0eWVECNEw6/4lLSwOyvpw5CBmazGZzT
xgjheyLqVHUcicCZcXY2vu4SyDbwpXD+RyIlUhOGYIKN9kMWCuT8FRjv3vf7ykAR6jrjauxn+K7q
xIFRLSxWtBg0pUllXIwHGDmCwlQT1K0qrLr3HnpLm7gQv44OsUHmgMhdlaYXobSgkizV+AK5UMhK
47fZ+nbwkgRHnI47JoIpuRO0NDFnXqbn4j2VgUruhsxj2KnaHJweG1WLAhs8dlQo8nSfNfAo/DGl
8baiCiUrH99fQWcVtawvA/ylYbmwX1XQj0Nysj1AS7VpJSvqVvcn1MZCUMwcMM9n1hl1hlTRNgZr
PZ8wue6B3bqYxwVntrAU0SiVCpv0dKQf9xKIKejKdRaUmUvYkyMW2PbCQxteI/1LRuHvz8wR0eFX
1DO03b4gmkcsM/3bVHThV9GqERplAbo+5Ijc4ISen5KzrW4IXSCkY+EvAQernwZtcDxE9BCgTDWz
RWt6/HbRs4xrE25hQ3L4ETWjAC6k7iKhm9I/mB5ZT+/nMoJZu0k4KoB1O+p96Y+F+K51OhXRsmta
PBS+UQVUZWeV31Qkq7nxd2qUnn7+XgBSFGLx4EdmhhDZiQvGg1zqA6j8BnWPaFisv0AkJSOKew9U
WzKaLtYTN0s8SFyWsT4beukjqIE70fHdwsL5gvfEA7xSUY2x5KIkBoGS1cywqLe69apIScY4KCov
mx73rbzEOoL2c0pitF9wrHyxMPANxXqM9AcUQhm+6CVKPsfgPAywDmctzu3H/9OzI3FOQSFo60ER
MwV2kkAGP7QNxCIwAFXWZLVOLBTDwESLh0tTjsjEDmdf4w6uaEe6DXDEWLexGGk9/F+xzuA0JUm3
gLBWdQQK7TrH87DCSeon9mftWfS29VoUQN3THmvz95jdxvO/cMfvvKkbbbbavJ0Oa9T7wAYOUmBm
COT9vM19P6il24yQmTd7mzgNe5JLMzEwOPA/ex8Kf7sg1G1ELTt5ngqlmPV4nXP2l7B4PYm7+LHk
as08joeK8yYk0tdlWJbQpadE6/kYKvcmuItYk+uMrIc20cwz7OH8QHzN3h6uwX/GvIS+69ZtZlXV
tcUAj6hbUqh8Ym3GuPfObMAaB04eEqQyfO3IPZFNpUhYC/yDV63e/wRyPV3IP9JBjx51eJIMTzM0
gnUqEyQdZaXqbYQt0lzWhpYTlKWbBKjSenJbUg3PncRXP6sq7HpLoP9QGY6yzO8lQvyYuRH1lxEj
3kp5ZqEXgEo61qfXDzT9odcIOqHVnokqtp8lDaoxyuc8o/TXurr+9LDwi6kKAMs4X+d5f7sSWbpQ
YLvvd1t/O4KcisT3Z8RhWQXH/m2ijUhYqKoLgnDqOT0XP4KlHVUGgn7/1g68KuwfeH3bYnz5of3S
LnpIQ27yg+jEM92+jnDYXOm+BwvwdwU5A7vjPOIFQLIrBh1lzxrDemy/6QGT5erLW7OHnpAnKfvY
9E1kmWdDj7IsOfYOBbAF/wdtlhANSj+SKxsyaSjI4h6a1Py59QDy6Kfj4DLqARP1pYZm/U20U+7C
qj7F0NafhMZ59fXJmR7LM5bA2CrK+gO53dveIYNpeSwZLhTZuE1i9kh0wptNZtYYNl3M/UauGdLX
u9Ro2LN3wJuBKACDU5otUR24SGviGVKe41hCOzTiS6RdllFWISR2hOspJQe0VizyDbTonkmfw4lc
RXVbQvBJJrfgwD25DrzFyvayS56fDe3Ll+fyCRSb1J6FFS19oufBvA+a4DPiZrqGOT88CcOPPYPO
kvB8r68XZVu/0rKGKjgAUAxuQgq0K1RaH4cXQQal+0TW5FE/yuTw1zjGnzqgRHUv6SDYzHzPMrZ2
6xYrcfrWRezXpP27oq+4rsthExDXNP8DVFlJs2Mh2EDORCXIe0uU5Jp6jbPsVKVHO02wUfdZbc8d
iFhRATrr3DhBS2C953/mPHBFzCqLKXyn/UBYC/45C4KN2syepGBro6qtunW1unPJUpJv+PMSV2pC
YAZOpaAKp5tHYS/W9/SYBcDJr7Dk3nTn/LuxbKpdZc4EX571E8vo3ga/Uq3fOlp7bTU7P/XY7YFf
Wze+ZFKQiYCRRCAOWQNpOQd+fGnYC9PkqpJ8lkeKd/xVzTP+RlXDUJ4o8BkJL4Qh/iHIaHT/GBWN
p37DGJZdrUNyq/iw9vdmJXwotgm/iVkZT1NmUp9gZS7bILNQYVuUqA98Yp9VHH44Zj17QgLZRqQz
2eY/hRHMxFsityrDeRTFevRojsmvGn21iE5uWahbIMp207X3bMRGe+wRNdW2IM66eQSUlpc0qzIX
U2s/3HIZXgBPKFPltgnZkkO4k/Eq0m37pcPC0m7VsFvFMkps44xkBN2DdJS+4q0f5Pvim46sRVNi
J+cFwwVBn0BJcfJ0rMG5dD3bG4PAQigGTuRiN0ZvxGMdVlxjWPXWZIQ6Yp3AB/KJ4Mqkp/g90wSi
Y0+5QUS96GDN5rnRDfi5aoJvOgA1SA1Cb+QF6hPBS+PIFrzQaYuetw4HhCenxigLv0H628CZdyDH
oocNBQWDkrkAhnW3UOQ70N+06+xADpqoVoLiY5FwODIRjonyUEg3pMmMC12EqAziM8eXyXnCDUDI
I0QhxoKzk4qG8OnRDnpU39WVp0uKJdG6yVi2tIa43nRchvkO7/jkgRVoZRI57WbqH5VXUVfwI7bd
4wV7o2+5r8h6aLojQFjpOr4dco5y3qFaTvDssLtU/m1z0PXmRp/8WxoNzp65AeWX6gyH9NpnX7Ne
8Usx+h1yBr0u7/R/10z94crSpRnaBqGqqO4A/zP1/fi1NiCnmkmZYEBBqhi+N3Qu2Aj6Cfp2aX1q
3umvq32++RrcliIhvaW80SCDUWr8x2KYeIGKul7raidIwGfX/sOT8OpV+Q/tAv9MYm+vypQwqpto
kF5pQdHGM8XxhFLAw9Sn/8QSmfb3I65vJnJo1yX73yr5vetBHKIIto8HbMmY4OZTxcROKHg1RMHK
li/Un9NDsYWPqSXi6nJkHIfz4jDftWvnP8todXV2z6h8OqAxTlptxbhOXyAq7cg9K4EmIMWyft+g
3zd0wvPeeWrx60IOKIiu/n6TJ4zus80o84fh16Q+9VtZFCzzyRTmFZVj99LyYL2+b233taAatG6k
To4pSgdV1BMgMmNt0UFg9osOc93E6t7DmIRFwYMOvp1xufMEY4kU3NDn2yCbbEYYVJ7FZc8JStTx
LdiqiKSzv89HlxHy8QPWDU5w36QBQqW0jZ75U4FojuXYNgaUeBDD45DIbgKKYxD77KFZk17k4eA4
NN9NHUbu3C3kgF4AuWxCsrRDeL7NuSEHKUm1A7dqFLFEHcXskKQf1y8/XbrYglfOChCv9fLN3uza
a4s+tWeQTWMJ2jB+qtcraolUKvyEOC5DWQRlHo7cx20k75D9h5Z7W4/7ILT+H41DVlzfCdUYK9yH
pscAGNuCsiE8JHsX7nrLchVmOh6kylggInHXfJcFs39tvUwoeOuigL0z9n/2o49D/DFFDemSrAjt
6a4mFfP9mJW+GZbd0G7XMRiXeUWJN5AnTBZkYXJGrUSXQCt1m99uOPP+Qt3bsYodZXzoAmTrZigx
2k36QBsGcHRUbwUTHztIrfpBR9fneDcTTq8yPFHb1ktSJOZ9Nbi/e76C8B2DqPAQxxIAalSHDmLL
+EWnm+qkx/9Ir7YAjx7VpUjQ240gPCz5/yd01utMmvMNBgTQre6/JvqW5hQSxBA5nZBMDnzFi5Bz
zEewGgPpNpacFxSIdH4Kkc1yr1HQaRB2M1/1oYcBYSUqQGumjuLYZTz/zyVNdZ2crchC+vgNKvmD
MH87uRhrbiGOO0vzVOeZx6CUy/AriHQIeC3xHwrNCH2/rFDgnc0gD3flR8yDRmR43431L9CkBljd
XT/YjjFDnlKZwV0z4D6QUsG4/tMsbf5hLyPSMZgmK5/IKjpAe7hTCyU14XSIMMZc1aygzg0guEzo
x2SZKoGx64RqBQrJREDWww8epCTIFXIu8AE/bEOZreMdz8FNqR9r4AciZQcEntvKKMmzSv+iwkFz
boJavUkCIpwPPB9XVVsYCJxX6Le++dPCFMUoZZYxgyV6xDf2Q7PiXmzEsm98Y9rUOD+866RP8twG
LMEt0w3H0BoBe4mTot1zCKLseDoUOvWm02ITBV2d44XQXRLaxP0ElpVW8LINpCJzfZe7jez2Ur4e
VnFkvb1G1yjpnHdbJ6bOWy6sIdw1i1zwo22Y/oiVPf48kG55TVi+wT5Rhy2jxZ59bkGskGcc1Icq
LkMRCj7Rq+IHncG8d+E32gB5Q/8o6EoRhUA5/rqkYCBD7ff84h9NJl8HK0ESe4PXlQGToYPFb4qC
ol/MPL340PaPQOFJnceUrT0WmaiguDQOedCafMzIMIiVnYUKaUekSCjPRIQ83jkxdnVTtUlHySoz
pDug1V5F08duY8uFYhQjXAS+bYgX4P2SYyoV1594OF8/CwXOEdRwAAksg8lWmwmcMH8fMXONPt9e
xMmQzXpE9rfbwaCP8ZJViIZXAE7oqvTe0kxCfhk+NjmczJKUM0mmvIeZ57uaUSbfyl3C1lwG0TNA
2bSOqJpSm4uJK/zj1g7gK3w7Qejs9Weec0BiQaXZwoXuc/WP15ejEjA7oC+cRD44NATlPYNU9KZ8
9NHP7JT1YL6GTQZm3WO5ShetmJ17pNcHOjaY8RmT+6p0Nl629rtUhfIdezTUJORHD0spmC47RIaC
08HogdxbwWh/Ssgaq+/PbvQV4OzFj1Lp075WnvNfCn9h181r8DDtNLh6zRvnF6WKHMv112Hi90Wz
U+vEaLt0Y+n1NvlaPmcwQGjdY2qFTpj821UQwOqw4th+adCen2Qm/xy/LdXnBCgYJBbunsmOY43q
Sqy6odZN8S3UG3EBO/RR/F0wAC5O5svMJ40wlpN54eBdyrjtx8EjfKDtWiCTLyZiFq8+TI32wGuP
Qvt7uAa4tj3MyhsWrMbEBCEuJdE5WvjBRhkggCadldG3OCGDjbxMXVqo1iSzY58C6MDSxui+TzH/
q6qpRN1WcBnuDBVJBzvjsklknl/g4TtjYNfIFztGGF3uI8lc1jadBAKCI0nd3fXdZAqlTZkt5EAo
L+/w0JuwWNeLdE6bEQXAEJ5NtWACJRp7S75nO1PYHumXhymDT6dYfD9y6z/92jCDbzif/d7G9/NZ
83fLWedqpDlf9JEW+jI+azQmAxv++piDFRF2dfeiGxrKqzZuSzPq0C+dj+dUyCfRCC3wCVC+YsSF
cKHNGMhBFUbvvZUgroRtAxd7SW0a9KWpVTHx3IUzxj/xHrSTH1n8Spaakecn+n4VSx51MqzLLkdh
s6t8yaakSvxuCciw1qr5kqq8fwdafoXizmAv8KkEBC/Kgejt1ct0q2UPrYevX9iz9dTYj8UShLzJ
mIyvN4QwM4ZtN6RjIca/N6WIUCfR5Bgu/grItjMaXxuXv4+LRb4GikQs268i5EcJgmgL/gw166vI
8iuJhMKUDYmUG/wckHe5gQ3v5BAkHaQb88Grvevbx/l70Qe2lsdhureYDy8NW0rvr0b5qJZHpdDC
S0IAKLSfwQ34oeePk3ucy+0uGHbd76O139Hdo77rji5C9yYmSqiERJsg88tnWcXur2Lvd8SV61uy
W4nk9hmLZ2pjQu3jw/iPUC1msO8qngXDdKhqI56+BPJS59eurjHI04mVl8teCiaJJRszLkLxPfE0
LO0gebltZFfPuVVAVWvgDyoyOigTCT3ZtYrarHR28XJWPs3sEZu/zkvShhhOnXF9zeHlMgU/Qk0i
opRPKWKgDNaOZRoK6hW/ZVbSywvLtnPk+LhzYgStx9DUMMKzwoipy473ncG/qZAsE6i10emumxlt
dAxHKH/1wiVhe036bw8vaCx1J67yauzjeRr+IgdWQJ/a5w6MeIRN08+FUvXBONfCTlQ1h9o6GP0H
NoDZjmizjX1TdYghP4L2NG3k8yZ8KjRrxx0vWOh1PJIBc5MlyryiWqZvjHAzK1nXt99Dsz9s8+e2
oIJsRcRkv4vaj3qCWy1mbM4EK04v/LT8pDRg5/gf6mKE2f/EfzdVkkCKGyJ69czilNZMGKq2hDw4
ANI0bptygQv5wedjwCYpECkm5HhsZyu+YGOd6eI5ofCAF5bua2zkFzRt9astm5VknY6k/aBpmIlL
5oMmWAS3YML2R8/u8EnXa+pR4+EblyTuA5YwE0ZbPP20C8v+DQpHnSLEtHh42K5BHeHVuu/7KLA/
OtZlC3ATi4HuB7818czXP7MQxKUl4VtL4G1WMTOASHGxhIkHbPM/0Z/KQ+byOl48FNrfQ3QxwiLt
YfwVyOvq1H1RV2B30YxgbVpLoRqJnOEWlWMEWHoQBCej+hNzWpoQ9Ov71n+m4lvtTGcEtk3bqutK
pquUrXMvUoWMq86B6+ZzPi95OZMq2B13ryDxvnU1Hwavz1Z8NauqGjlezd0loc9k6XSm1npG68sD
+4Q06BvCXHRvS3puN92D5iTRO/phcKFz2LjxKfkTXugvz0FXt3BXUa17wdkPUxSRnyYXevbWz/G+
6AOLyYxyg6Njolidpb3hr9wAY25NO0EdxlfK0ic3by4gv1zdM1XU7pzxeqqWIAA5Srdp6inh/oO7
NTDgZQIgrVFKANYYU6ebeBR1Qq/vHctLOOvlDjRvkXeZ60+4QxFIocrt8+1YS1QflrpzXX0J/c9N
ydc63KmI+IXMvqzbql40NSCy+YZeV1ZIQufPXgw3Q34zDi/kz+1s6ufFYVer0/rC5EsjaMUwNFSA
Md0FmwBtz38Eb2eF1NRR6JCBnhxGzsKtMNSJQRY/zlnvG7CERmXQbgPHbMeVby+Zt1VoI8PzASmW
e4PinPLXPJzvV/61m1NRPDi/mjjhOP6jI7eWkQ634FNsGug0eDyjImShfxINwoARlffSuADJx1pY
DtqADFhcQJgxhS3gp3/8toyTsH48MNwzeILiL16fyyKQF4Bt5U1SkAaKXe7MO5gBppB8yqEmFfu5
MZPf4Adkyyr0REfV+Wyj1RmJXT2l5i7KPp5ldZVwBAmf95wYkqTgkWMMCxDKJ19vufCH3+TWMWnC
YWGTqBw87OHGIPCbAqDrCGQgB0pkd+74rZ50R4jZMrGv150sirpHEAQJWTKS09bdBopjL1mgHWVN
NBa2VG6+xx/wbli5KjR7GJ1/ir0V+VzQVExK9tF1D/yTTKPFAYzM3S8FakNIPR0I77aHjR3cdfPI
ZMsPKgT5+f7lolI/x+HqZLaIwrtxqrOtzEj8u4Sf6NoGx/ZqBAdq+Q3s2wpezUfNbhGMRyXjtNd4
4EZUJetW2fDFlSI0Y7AtebQY8Sz8tYWWXDgJ4ds2939r/2Er3mKkRtTpMgiVWfYSt0Tersqu67oX
eTi5pTZZirqWDlnFQ2GQvPKD4Q/Lzj8UjoA6XuyvpM2abniVrfdT/afaHtfgXuww3TtS6OZ2mpzC
NA1yUV8EUPj0bZh143jhvXfAlT0KuVBZKsnV6MiH9D6hNQEp4VITx0ywanosnE+FSOBFHBXBAh7j
lEIVE8L3viC3KZV/9nbaO53J+RV43woayJ41y6p2wr/Eqtbj4UlvKMKS+WIs/h2E9P3Refj9BeEH
SusdNjSRfBZYkyrug3JruMYDWbDkIDo7xgwo5FgIG7C6BX61R35cN+0+i4882SVFVhQt3u5YpjPi
YbC4ohSCEKcKGonch+eLAtPD2G2GG9uFqLxxBcPaEBwCD5FzavctoxahhlAtlPLqHblQSB1t42OU
k8gF15zyG4Ebw9cZYjS1AZfoZc9/0AyJPspj5pK8tlhAgTPq7VhCMqfXhDBVZ6Kf+yr7ULdwcsrF
1NjGQWNsGnhCB43OtgASw7fzuaRAERiVplbix6spn7d4d2j2AJZW1Amh0nSVpNq2PiJ6dYiuyp6A
ZL/4oxnvlodZaOJRvIyWYpPf1khOf2P7yhRAAy207t8CnBjgZpTnOpcV4eiVu0umxu2ScWPYt7vK
SO8roKvs/6+in6CkB6dVU/C9aoM1CU3cx0myS+l6jW9N+b2cicDJ+GV708NbuRo3VK0gmdvisSW3
L6+w8Wbqfcc0twdd3cnfwc2E0QI0CGGy27xCP4QFp62aEpm7Z0m1B/xS+7VMqjp9nHdrzBC9RMPj
2MaQBsL5BnX1+7nSeLL/PGhopsTsQX4XZLl1yuVyN6+yQGSV3986lr+qkY8bDqmo9/N73INY6rL6
8TwdOwPFCVa90Te7fpaLXGYJu5LYDxOxiyFUoKjRBhTjTcQosM/vWXwHbyam/wYpTpccL5B8bYBA
MvtNM5wFGRJpGRSc+cOCDgSbsaV0AnKSaOf8ZytMWIZBWqgc+L6MOsIh7KkmVL1cTd/hNweHhgRb
UyhbTqKYyh10Ib2wYoXuSZiV8H9ywy0ELTXYI3sfHRL5NykcOfWzOYJH8Nel385n1ye9u+SaD4IV
Z79IWRHxGkWpVj9zB4qwVJdC39OGH9nMCKd4ClbZjujh2u+WBFhcCZKqd6laQbsLU+BR/TYdFcHp
gwoAWbpBB40MAzZWK0sI6823NpoL0PV3uZ1HkQSWWsFztS27KcOJGsTr2UfuHaK/keIlJvdv+Tq+
1OPUyn6FffRCAdvcFbRWLx2CdE7LiTehD4rjgB00dF9vFsxdhnUvCOfhVtlzyVQNkgBhesThuUj0
j+E3j3oxElRY0RXKWzrcQwqDin/8YeYIVpjbyCF0u5nE5VzvFMQJKClAYAkrBrK+bRVNMmIu+zxY
31cKYvhdDlRTpnluBy86GmFZ5mAgtwS0PywJJcHQyqpXl6t6xZZ6QKg6pmGC3sIDRLL+6cSRrqSR
IzoUTvftAZJKKE8hfFU2EY5lO+yTSsCqz0dnFshzaTx7oAOVl3wf585yKqvVcSkqq/9DT9Trdp+5
RwyLTtoMUGWBLEJ6ei27t+x2Kxt/rGOlj/+NnbrK4yDoQOVkQDTTCbHg6T9o6UNhrzKwftl6dEsj
RyVSzphU47dv6yidOy4WsU3U50vn58XW1SBPLVpSsy1aLCAJqdnwaJEjDAb/apraK99lNLch/4md
lF/yaKzRYqO7kdR4LF8nlLENSVObqaryvHqBfNHFJhbJ9qWSvMboH7mzDnfWteHFO0jmox/Nx//j
xmQ4bOtsyBPzFfj88v5zeIbdpEcV3lqoipOeHiO899E5K5lln0SobwbNyKHD3S60GkrOOJqqGSGK
OBtpu4ejXKTykn6giu8IdUH6mCh8wfsRZrvlgoqpItwPOYm5sSLbQKRVbk32nBcE3LxHMbdLr9N/
5wyoMz9z6y8gcwspkFvYDUm0sFSwoWJakd/AU4PZU3sYpio0PSr33tddtY8+tU3GVUsZa0Y0w4G1
8HsZOiXOLSEvcl/9AirUcC91SEkRBU0SrIu5JlaLXbv8OhyBrwIUx4LDJEBZiQ8nGhCDMT0Fbzp0
dSko5jcpNh9RxJtz3RKjvAIjzY3QCMGRYV7UKZ+U+4CSHL77llnuRY+mvtMzF229xrAm83XvPRXK
Jq0R/vtXrMaMB1Zs31r7Q6YV4gbHcSwBgPXQsc9O5oRSCiHOuWoQkPSmUgUtuoZArP2IRuFPhyMP
SB9c1sI6NYNF1SGk4MixRJbQY0hnneMiS7xSMs7i4tPYQtU1HUmsiq6TsQWiQwCz4p5s1R/k0Xy5
68ShNdzjy8+2Mr7fwXwaBwhbdyMPTH7y3o5PelGBuQcJ812dqhGmL3wlLHoelz3qV/Q1maLXMtCq
cssot4QmFsOXKncXaA3UamHHFShA0QD6D8CKm0MBC9dWEq6vxz+NlE9eu05uSR3u260u0vmE9fms
qWF2CnROCyBocGTBm8KEUNSlBsCGi4Y8tKsQFyORlVYKFOR2Ly7TBHnDTGZQfCi1SB6tPyer1M1U
q2mBCh7Zj69r11qst9tRlcpnNN0WziRnT7kb6S8Q0DnpgctmF5BuzIsbJ1uYGTHtKOaMxe09HBkS
M0mDELSyE/Gm532bW6f2nW1CI4LcliJYCbFwGKGmWmw2QM3vCrpuQrolJIJECtQnGAs+UB/aXGYP
nfba0fj0z2XoJVcq+x/uFxVAGEF1JB/GSQjDi2IKbjzTQtNlKy6w3PVGXSquBReU3vnTmcaQy2aA
CQxyRCv901E4AVdMYikGLt8jsZrLuOxkFMcLyaPj/ueH+cEg81c7QMF48xSc2lCA2KaWnJATI7YQ
XY5RHaprZxcNwUsdbUZ2W4OByrlqi4AXpyz7nz2gz3bxPtzxDwZ+vsFfdzBIDcDP/BwoXC3s+e3Y
XaIPn3oGkX2B1GT4r5Lfu+OHWZsZEdlZqKouLDWUvMqjBqN6esLrIJfVyav+9xM8DowdknG5O5aW
78y1jNYjfRIyhDvgEaArBq9/nSrvByZ0XVKaFzSXLLJDclN8dllPYecvnuKYJhhc5LcIQh5MEwc9
2JFItkJ5FcVLyi2zGiVxS6zbHpuN2Rs4mHqTTEfNGuB2sMNelZ8BkILCB4t6CipoqQxfZJbruS2l
9GZm8mXnKtnLzrqeioTh5+AiOqd4/cS/33mSkdkCH53qIilZS6kZb6/px+p8GYntJ4RvnOM8p/5w
bkHLS4MptVc4meDkrUe2hlqhF+5ijO62ueQJpkmX2rkFgWaxLiRmNRc75edXTC+kPf30yTQ1VCJW
BxnSRFheGLmfvKlWTtgL5wyGkkGzzFjx1u5oGJjWrBxqkRB+eHnslErHEMYFsc3yecRplYY5kfoj
8cUzraNthT5S+9AiOKe5qcMc+4pwjOB7lApzRRGjNwCi78BKJ9XdvEevjRaLtak3wcJ7ntL564tQ
a9WXPQ+a1EUQPJy35gRIzyg8YDa1ZjMFkiHAyr7JTANUYDZBx2uWomq4q0UmV7yv+DjaGpj23wFe
9JOIxi8ilz4Rn2UieJQ5utErX+7difhMiCPc93Q2/0yyURIxrzakfQTZn8J1nEm6iygxb9OAcz2g
620h/c9TxWCjcCQk2ERrv7MVreZTZEAc9uJ3hO/pLsi9ytUOfUTxKrIzv2tJVma4KgDp00+NQu0n
AdJtfB1PTzMwq6WEECF0DRiJ3uhPIHB92ZbOO/aRTrF1JkHH3xD+atEQlllN2T4eeLPxMPaAqQRc
EFXIxaNWS2r3yISAyniFzN34A5Zu09Bc8kuCnQBPZdtT7k8loJSO+ZgM6mvSmgmk0mbCKFfVMEeh
3LrSUxa0yir1Mpj1DgqxhPCr47ljp1HuNOoP9aBCz40Zs2r1s9MexqIhVCycL7dOBeJUY/DEG++y
3/LodsIFekght3/AJ6pCtvdVOrSoBvH1z3idyxm1IFpBTzHQKGvPhMS+Ef0uDpsV0Ag8LJOcNOxk
oQaudk/tzrA7rB9/fyWMD8dDiWxcTiZZeS7F5BYoVzHe2lBdeg/Tb75MOlSkfEm59eAjwPwNeUKg
Bf6VwK7h8wV3e0hKBFibtRcVyNnGuPFvF9mnlcyJ2dHcR4jTpKkJBxR7QEap3JF6YJshYPfiQsKp
ft+OuEbcI03QbJRUqy8bKuJUUgPsenffwid4qyX12br0hz45pFaRHq0OWEFDk0Kuqu2SrSGUCvWa
mMU0AY5Wkvlx42Djs6j8Ca3VJiVvXssXWjrpSIHC6uppwlIdPXKmb8KdRrzPW+EoW0wUFJx+Gkj7
cXl52Br8tonEj9zelaVWh6exKAPFD/zsMTZVCzXt2VrpVzPKf8DB4a0zfX4/dxyam7w/wLBRjGuq
BnW1O50wnncBXxw+oW7ih6yZjZ+r7rT/WdSxRYl9eEsipIaMFdgZdDbQb+RSOoLrWdMvC6o6O9kB
jNyM9LYCi7ZMaLj1Ol2W9+kXaKBPg/48E1FxP2Oh4ZTlD6HG+eE7uDp+5iq6dYoE9WJVTPU0LSm2
UGAoregT6LWLah7AspJt64JUrGui/V2Ois/dw87pL7jxWZ27SePhH0UERngB9J68AWARgh3pgfw8
s2T4t58y+HslkKaGUkMjnIzPUlOgr118X6Zr3aOU3u3/IGSWSEWiM+G1MXvsqPqMgfZlYFea6yu0
Vf8VcnhGqm2vWD74QhfhVXPcr/K1g0A+V7A8B0znaFFWQT+IZ7taeMi+7zXvdIlLB5BedPnS1cTn
zzRwfYqUBOjYMJ81Lpx7bTWBdS1lDHZ3ZaQu2CAvA4HGPfQDsloA4zLyrZctg7QEOEwY3bDYX5Kw
sy7p6DV9BanQxuPu9A6qsjAgVGSVvxy1JKlbPPRmvjYC17rRmn4y2cRBGZnGvzMehYfhYj7XG2tK
QcRBh8Trghm5alu12Cs88xDSsKjbd8gcjtqhvYppWhaa0p+TjinFx35bv3moYtHi2aW5jgSzM9UD
Pi1vvNZXag6M389qjik70QjYaM9v1hl9yaa+Mxuw/HihjxLhHrpyFzDL16Oqpc4h8XR01V1S0r+O
pb35DZak+sKNwGq3JZ8EDcfq4qYJSDyNkuM9/ogXRXbcpBkqL6IqDnpaJBz2kONo7evsRhZJHNXh
VCz+3pLOtBzZ2gv/8RW03ZCju8ftjp0MP/KMoVgi86xd3NJ4P5zcKAegACw9R3MYQGp9bg12aKQx
NnXrIvF3F42Ck0joLX+38JGSpad4u2Xi8zrPCfTtUTBO5DdD248jhEXZsi4dQMZwtpodnMSEGe2w
BT5yXe73E6h52Y5pSsRsCiAUKxhS6fokTCw1B06qWEGt7QGNXRrvHvn0SI/EKAzK7gaO3IhE1PlH
n5IazVdIfgY+y/jkgtMis2PPa/RegQkWdpk78HvHz1guw3kwc/XqO/CB8HcxrzIXPP8ae6HYIHC6
DQiYFmUVG9WRCuhFfypqV39Iq9oVlTJYoMAGZDemH0JbrGF7ef04mnOTvEZq6MCGVPhd+Co66qVO
xZ4HaJsnIeW+oyww6FETQV1rppOyRKFu9/RDKQnDpYQ4BQ/aDhF1T2/5tvMYLqDq4trix6kx+i8l
ck5S0qrYmPhtRK2RL/Didyb4gBoQvtlGDFIJNb0tEwLzZZPfe8xgmgzkDgx2CPQyJeEljKzrLNZg
BwsNqGefKFr3mRLz02m+0Vkg8QauUzem3RDd3DWZP60YbvjxUijLGL4pEve8asc33WOOMag9XlBX
DbcgDrQ0W8IkJH2OdLayHhhOQ+oiOf+p4At14k87a5sxA8Lx3zl3y/6gBz08UkGXA09S9R/BHjYU
pz8nX5ajxMF03YUfJeaVaaVy6vEGLQKFQ/y4z3TzKmwDL4Gj9ZRzcadLlJ/Ck6rkGucYsJiYbx8q
4esdpXQdDiH52HCbEuIA9cKqw3d1g2tf/XUs9EFH1pWnhg9lM21ShrflPcAmCzah56Eh0ZPleTRK
UAB1EYMQr98xgtQDOyUoKR0ZbDz0osqUxsOb8IkCQClb/3d3doS8f+w9HfAc1wVSTYs5uRe5/UpK
Q0uJSU8pLQaZYSl2oEX1OXsocjC0R0a+yxASXp0qeKxIsqZCWkaXaOWcgn9sX4a2q2mL0aBjgSdE
iTkmaUtRDjqaGRQ2An+py24rYkrXdRqo0miM+6hNP6Jp9fbexQBr+NRnAJTkJtUyOq1cXCADfGEA
8njtQtgUFx1Fc/h7jExGq8QCNgtmv7AtAYwHXiVKY+cMN+jv50gWK5AM9n80UbuFFHD9E+PhZ6zX
SAuwSIKRamd6ZGqHhxg7E4IL55k6TXw9GQDOZWUT4hpJC9tcLFWJBeUegqcBpOY/mRXshxCWG3A2
YRiVrAd7kHK4vGMMScbBBHsOYbeG8hf1a9QfUnVS5Z65OVnvn3DPkHLNYhssDj3/dsrrhkOqYrFH
KQUPp7A+iKhzSYz8YG02tE0wUj+Vz5LluWeU8KBLvbeSlUIS3p40ozZXKlGGWq8ct5e8JDCdkqUv
sz8Egz4FZjm/V0cJTmRu27FvPI3dm9v6Mbogy6tCLZdNY3xbU2EPvtvNADLNgYylVCkSW78PvAX1
xGYeMzutMUo8iiJ9lFxaZvR0AsEtVHTl5ZiU0AwFHdLyslk+jeICaXBMZofCwi/xBgjLmwVrElJD
hKqS2zDRN2qQ8EY+mfBAhQPQ3V5Z4r8ZNJKJ7FSHs5ojUZcKah9IreIXX+SE263ITxEhRwLqGXAF
kG2ap+gb0yrAm42OCa0D/lKmk+GLxX72yrfbo8C5WZ+uqBhO8NbXbmG47gL19HNDURFD84qX4BuE
Qn/2xdXyA10Ug/gdkBUyyQFwPVYUjjVintUQbR+YHrw3x4dpE3jQCMOO0DqlG2XjTHUpLRejwpi3
qG5v7y0CMMKHCu/Rs2oldyka+uwy/a4I/bW3B9BMzz+6HvXeqJAhYJPNkPHJfHnnZmC7Sad5KHNk
+KZu6sYJPdIKUXb/mVrHgjmapbzuX8kLRrnvn4J5ywY1wm8Yt6FBvAQCy1rLw3cuh9QuEZpkSDoC
k+yQWZ+0eVtQCxGKYX2eZxARw6GdDff01lWaIOLDFtoO0Noh3BhqB8GcEgIXdBnHJ21lJKFfjPFr
cT2iK6Ip+6sRHr+K+lwLqXxxPqbsuN0P8NxKIW8ZzwR9SGCh7LCWtyV7R7TmdfYSeWBT4gc4wRKb
iQeup/BrQt421C0e6yh8AdImsA9PocrYs/bzU84hWwb9HfZDNr7skRYYUICEFOvpAhNcQ0AeZ9pc
7xk8jwPDrJZh5OCcfQYWRUSYXubCQI8x5jn0J+MBxmwRHg40R6JWQigyZ8jFVFM9jP7+AdBzfWdC
rxxCZU2E9Uoks1iK6Bc1vg9Ym+h66no+Qw6WaunXbcFGAQ96PiYFYAyjODlD5viGKC0lLu122fSK
Ztr2zDqpuUYNqARrYNG5ottkBUTUsZjC0BarxNo0R9ws9lV2NPY4/FOpMSOQeODUxoEl+k9xiz+I
qzJngiGiMHy3Z1FrGiy83Xk/bZm1SlPjOY81+BVTg2+ZuiwYNiTAEJgTfn3DbDgdHtXhkUcv+nx3
7nOXaRiVr1iPdvHcH3+YcWJeVwyjMaetivUOkbfgmBQBnywVBta5sbO897eqcoyx48Me8MC3PA5h
OOrtcatscx4VmBzyVII+B0OSRF5iEs9t5dMu1WZV93c3sE8lyEnX6OgSSKQsH46UyqJO3pLodmiK
l5LigoyNS9HYKQUGFVh/gH/XfJTcTKiMNcfzKLnWzw6sDqNpKnd15Owq1yc/6up01eAx67N0m7rq
1b11abRJoPiKU7pwEuJKwfy9jo5V0Wyjwp/PjW53rYkw01/va1yIPbqgRZ5SsfmBHUWzvyaqrajA
r012xPp2OISUH82QYzLPC6ocY9vamZrXe1gcsXYUR0ErmHnih/l+JfNEL08x4Y1YoTKudO3pOG1y
LoEXJAJlgsDsX1pNZ/M3bkmA5oq9M7iG4b88j7Zu76bA+dij6mJbE+6gKtWe7djpzHCqYqCK6SsM
ULAAl/5LHf8nf/+uTxZxg4rFiXY+jLOK8qr8iv5bROylkH2uLn5m3xZ8NsqnNF5DlGJShRpZauDi
aGRrAFOT3Wl5BXT+ZNs7xTNgj+cfvMymT9/cD9RALMi72gEJBodWUYMLVn2+1chmi+wkTOaaD0+i
uxQFpB9CgjEG9YUgsOTL0Dq68IsabbcCNrKP7gxfrSleGMPuq1n902s00KsA3rtOT5uHGU0bdfmT
Wf3J3JUbUKdMrKs+qNfAjQs3eUkMK9NBy8sBuA0AJ3qw4pGxjqHOao9aFsRl7ADgsuAMz5zx3asF
1zNHKmu2kOAL6qnSrWtN9jx1ag0mpIe3G97Mm3LzUPNh/JPjP8cdRR4ViTHYVNBqdavq834HhynC
Jml59IS73DcGF4mf1371KnTllYhSaxtz3MkQMHEnvVnasgDCRHqeR8wVFEpdocTWNOJci5kNZKCo
TJowsSHxK4FQKKizN9B//6lXb7zsMAcPW4PgXq0Y18gwC4BfciNu38tBVU4GlyHx99bIxah7qDsb
SOn+vbU6wUaUZLszPgAITomRxvALLhw1Yre6r2QH+uabg2P7Kypm11oL9FlmYNA5vw1bNG42xDrM
xPsK5LtGC6dJSzx2f5a0g5DqimWhrnDfSxwBATf2d2vIQFMLcffJkqnsy6PIrvMlAAn44/qgoJe8
uNuo7c+XaoHortBhWt+Sw8oMIl8gv29uNIyeTnVFPDHbCe3G1QY3+tVmuUQy1vvxKEma3rZFlycJ
0uyLL0gMq6630CtDrLwDnsH/D8DvUDngqay42OuejHnao11gjpLflm91cP2jWveQZVX5bgPPEVm3
WVUdkRB/QK9FIi34jsnS2U/KvlXBMUxoGGlf99kN0GeN2x7LgsPaH+TmMM/ketm3wfxmO6PcTJiG
W5Dx3m0RLf4luZahkT8/yICInf8QsgWoAE9LWpt7Q/e8cYhep6dcsaCfbW2t/Jq0L+VRIZPoCewV
RMHxFPtrVqj42VBCdx43vYpCziWn7gA77TEfgfjFwjUKe/iBykoqEfBdqMiZEauH5Cl71RfEaA+Q
DUGwzzXS9gC+YCOxICIaVompadSScLToa3yL9SrRahoWYCzZaVMgd3xVs2CBs33ZVgXmpk2YzNsr
Wc5mv11grgCVOKuKJ5rM6+ifJ3+9Wdw2cbXSLr06Anlu5TbaviVW7TppHkL9fh6RBhEzNCO3gEae
6pN4TTyNPBvQOOEHhF0XfopBm6whbzit7C9KXsvu6V7bcFd75uWUwYMrpE8nxcpirD5JZo1uy0o/
t2DnHvHPbGHOw2smIsBMPnXog5p2Wj/rrvXFzKF09ResWI6JIlbyp9ujwrSpFqpWh6/UoFEbGNTS
oEcqpGXiXPcfVqKXXtxtH0bADe7wd+fZyXWgQJbI/FTLKwFfLqqUX5xM1Ub0Cw/y3g8OVlyiVmiL
X7/g6VETmO6FfsgQXNrxBHpq49Qde1Jy+XxM0sCFXUCwxlM+rxCB68O4D0dUFirVtL5Z9eIEzTA7
xDZpiH5EUZGplhRXZl6quWJW9qkAQKAY5fdel4W0FO5N8fVlMgIHFHKsge0iL5y4u61kws1yFHtn
qOHbvHKDlwUjECy8obrkcEUj45oOZxUXjGTWH2miwogZMshMvurFVgkMDTUsngc/lazhymUawfeA
b9WCMvK0VSHLiuzs/5LZGWbt9XebBqMEnJTNjF5Ad7BlEd/wqcqWZqol8Wjx9ImIIHC2tZ2PudBd
u6vu1TcP2IjivpmyRbL4ShrV1G5syCxQid8EZeZ3yeMH/z49SDUclMjEz5qJun+DICHqsTtSO7O7
u4Lvv5V59W8BAYrzO4IImN5cPu51SxhphVSD6ksFyv2OJOpofVZjp2CjnDzl/M73rO1fvlr/flbw
fXlfA97Ha2TwFJgkVthZlvlJFJpL9f1DOpMG+BZOTsvG6Jo7wm3Ci/TM0DfGztulazgxhy15IjZc
dzDHR4fqV0ABrfSHw7TB5WWYhEfhW5qXtdvlfIiTmpFLA6TI7tz8l6dUn/2Qyxc3y/i5J1O98GUi
AV0PYYoqVC0FfH9Uo2WkmLb8OdbzY0xCCx1e1eyAg1Z800p9CALQtCRxKcm1+JRpvfA8EqC0FpId
sMbrZNGfnBfNb80Rqg/N8nZEBgYVGnI+6LNSjxjlyMNh2xfyjHV6GvdRoLOJjKLJtNSjgAKpQ0oB
Q/Tcf2SN2/VXQ89p/EA67/TpWEDY+WEqFMg4Q5MPyp+pzUDCjfx0FC/MrHVBJrGrmufof5N/A6ma
0RlBXABFY3J+v0hxDCe/UnXIddWtpv0ipbiDt3QOHglOTcgeLhzOHL0TUdrSOd2HPGFRo5GtKwz5
nFd+yoN0E+dlvDdBof8iZgy2EfvyDV5o0or8sHaBHnxMeCTleoE95kjkGU79CQVMWnz+VKUolEMH
mkbFbAFBz+pc8XiowSucFjaHsEcSkXQEK4Q78wdCKyE5oGr7l5n+4yAHaTUJSsnI1A/wByKC1TiN
iDVq6q+UX5v8dhaB+AMPO5cI4IrLpSCmn9oPlgnPFJB3xKFFcMyPQc3ugSNd2EEyLS+sTEuyw6QB
CjlkLLBavBIHedNEUl2apMj6GvhC4Jdp6yEpe/1QvKiPtuVQsEpipx29pp4JMxn7zKYqi+awnciy
aS4vQhdgQnUri6YfQRssX5IiiVbTP/U5E1krqOoS2U8WiZ+jAAiSTcQMYsTrw2KYX4mcGsOTxG6e
9ZoRRbHNBRK+4OgB1Ck4l9Np90hsbvXasiFNRrzvPUeFBT6zO7SLhmjgqBGD3wEYvqxYHX2HrE1c
Pt8S8cqClOYufGcHpZLtElJ3YbYn+zlIleai1nWMpj/otEcJABrnCykTLx86akUnhR2GLMquT5Qx
0P1NCXHH8dkdlSHvjqCiZO2zMZjnLP7pbDqQ4pVsTNAxk37w8N7vgds1uyGfRTsTluH8XIhQowbk
zf9Udb8oUffMScTMoRgNsvpZQUzPACa8mdiOTXqp+38dz8oF2EmLp0jNWpucMVxA6jpGSh4LZnEa
/L+lGSNz9R0E2FVjEzU9ORwIiQq17ZS7ZjHDCa/qm4euJsz1LNnJehig/0vdWoM1TM95ajnaiDGM
qup3ERBhufwFkq5BnZlcrThSIfHvJ0xPpLkC9CpQn8ABwCNGgf+5MOBNsrwZdRzY56yz7IBSC8lv
e6meE7SJXe4R2naZj+wz42kLDuPLQZePTMTJ8adI/OuFLZQGWOwo1HN7wKLGRhkhKjUghzRn34XC
1lbpGxK78dXlLCxZS1ROsRFDIEXPIq8V/Ysu8CHAzs6sH3CAUc+M/Poc6vY5k0MS3g8Xvrs7p9mg
NPx494vBWGr35SWrhUBVlJsjQelNnANGDrARWrR+GqwKNqc9QZjHNbWGO/kjOp3k03ckM4ehpBqA
kJBKaoe65zzUpZnGOK+c6dgCemhHtgPRsd1yCbeTQuJgxl0j4zAPCNF/BI6uPQYVVmiQ3kg0eQRT
XLpI3OA4nGMZPAkX/JuBGiM0mXG8HEElvRcmKTFC07RkU4rs0SHPwVA20E4DfRGEurdGpSkvlxdL
BPvJrwMGMqLi84YVdj4vAC4l+aT4x4y9eUoXNU6+oiY7jEdU2dv7fhFzrxqDIdjFcUnTweDKPgmB
HAep3g0lkVriQ8Y+qbjfxJPV2PVqT6Ypv2W3mzFOdHMMvFNcMOh8dAhgXQD8aDKDKbFka8+IhCtS
OHJcJzjXnUX2emP38x3mQFvi6usVHglIeAnbO9p4sYpEEC7TlDTJK+g+2FEggwENGS0sucIkNXtg
PxcOOBxJf16YPaxEWXm5rwKl5zGp9CzkiyjDRQ4pTGwOeA1kU+xKRjyVtY+7l7jJa31Ew+kDsLf8
wDyll9GJQFsI2YwByJ+OFhjZbb5bjBalVV899/ygFaiUZWh3aov7BJWHWXTZYLPSl+2YrfGQGpsA
XTQZNsURIpY+U4MtR7zVecKJjN+AXjxhYL/W2sz5quy3bqIwMoOkEX+tsVR7YVNhOXVaxGEIBxKC
K788uKNhlFG26w+Mb9bptCcjseW67ur9PEEHi28nIXmXUcd3HhxFOHKenOkFcpI36mlawEmM59Ia
Y3J+y517nhX1Xdf7ohreI7b4naBWrQsRavycjMQuPLPFF/yITod3oQLFAk0BrtVQe3l/2wo/m1CE
meiz2qcOs+Mh7bmmY+hh5SXO/l9wqw+Axi4jwesuvANEfkxFCjUF0MabxUWEmATPgRT5KuLdS9dG
Z4PED11sPWsdp98n8SX4+uU1VGx8FBREVIaGwI3SOacVSwGU4Qj7wcyRXywgl2S1BmvwT8V9YgTH
sP0RkBCB1DoZtM/f+QdXfbxEosxDibDeKU7PAH9/CfXUCXaz/E3y3Oc0+MRs5R4Txb28Br8sJrLq
J8e1o61flz9zJHTtRe2iwXM/RRmLFaJuX9daC3BCM2ufdiKmEqcYi6VMRLh2GTEJ/n1elgcCao+Z
Nz+tNFEliNyU2K+x01mnSysaWEEiM3+oQrOI1YVSzAwY3Zs76uD/OpHRYAE/oYMxkoBZsI2QH868
6fp08I6PQPxrxm5ZHXoUEc3LJcJwum8IgbTEoFpPg+jo6Wr6dhSf6twW0R2Pbb8nA826TKRDcnuX
/WT6x3D3DxGdXrgUvEXhAs9Y+9jVFmUhsx2YpJoyybCsGvC7k4/Ma5MltT3UhmRXWTCIEpiZG/Ff
SZPdiHbZ0pm9S07DAUhNY1fe3YNVHnJ/1bQKbRfBHPs4f9cQNMg9apMuJ9/Oe4AEgEcH4pjLta0w
42S38C2TPdElJCoJ96l/1LCn8FP0povkQ4gNuA+jRsRqMBwXTv0Tvz8NXcwlU705SYrCFxJojkQl
tOXKRpiurOFikJ3bGRvbFYfOt5sld7XdppQmVdQSkKhLpxhmATCK9PP7/O0MS1PJxqhgHL3i92nw
pM3xQhzXYmokD7BMryb4+Le4/KcfaoB+fEHu01irnfRYr6b5l96njHnf1e+4okHEYTvx9DSpcYSe
zfvpc5EXWq93VK09F5F6x1xsvPpisoZ1JKXgkF+eJrNMchH5HYS4NngY3kHg0RP+NzOY2/wvba1T
1qxBE6ZTQaoH0CFOS3YsFBZcsmXsa7zu9CVvEwLfOvl3jcv4HecOsiJkeJd3j8MZzKztL24L4UYE
4Xv+MsPZ2bgohWbnhg/GPc+Cltd+1jJ1WrCEgCgQEboiZInYkNRnksjUs6hkRU76PLon5GdV1VOK
h4HW+HGgqu6FdFjy6K+Hwt+ix26s+Ndwyw7GAZiRokUwdlNJw5E19Wn/xjQortqhFAx1ccP+gGhL
Y1rILK6pcJrgnMFKJ6rKua7KpNFSZElllTU2S6yejQ1rV/qiumNbNmTwQK8z9G/gokeuCBR4ixQz
uElPXnItvc/8b1NTUptG30ySVfd9bWlBKCAobYnKU5I1FAcZjJ/0ninl04wjBf5yMIXAdjEfm5Eg
LuUpqSMuzJ7yUSS2wYH1m6ng2Ejg6Qh/EusnHLGQMJC9vpSyc4rZVtzSukdn6mcs6Wguo7wBAOjf
/ytX9wGIuJbhuPaI9MRJ5pt1I9vIu29mZilutMnliIszD1anZ1w854OxCnienVDzJwooT5ybiW0J
6jw4FusLv3Mof9p4I1U5DydZ0VIlEc8G89otiDa2o+xGx2LDLly3ZJY52piN9CcOxcGF1reqF7PA
G39Tp2V7Pq0lMwsHFJUOxRCRo5fFZ9JsegCL6V3cE9a+qdhRsuEJHPdWTwkMRU/N1uC6HLw4mc7Q
WcvHXiJp/q5iXDCV6Xg+VbqJSNE9goW+BVOJKRCmVMx/ifbQKxq/x5UPa+k1xWsHWUcEuzfpKI7i
8EN5/PX8HUARXv+4qtUdn4N+j3I0llD+T7HzYlqGetGzeZotKZTiGp3td/zxUZalbzkeRl0SFiNX
mU+MSUXrPNEaaru0mRlyWq2Dul3LGE3unt2TPp4/u638PQKI5hEnpFqzs4A7u/QylcvhIHEH5bE3
DiJLpVksfPCBQieXbpEtUdv+7vz/fHMiLmBnCvZE9g3X7a4iLyhaPNcIPGmFAy4ttEvujpSiomrX
XY+6RpiK/UZeCteKJWOJ3RCa0lroCXeiaOoyerBdWXgJkMi/cF8OoM1+d2jRVJOEF4taG6wLUfTN
hBqnn0Y0PFwsFWm2Q6k2xvbVHMsjS+guFEQLUC+SZzNNAamwZNMxxgK8BdvM2QFakgnTPhZ0yo/U
WPe32ETcZlHTLalTxHaLorof88EJgk4xnP7a8ZIUAxbTXf2VAoCRp6WmSZkkYHG4ARnqrdvFqgOZ
aWWvPKsXKyw8TNgSw5vPRtQzh7CWzcqfTq6A/VC2xPp1hdAVnw4+5v2iHy2CQqisY07JR4FbiLVl
CTyGO+0nRG9IH8ropwEm81qMyRAdwAPCsRLzi2LWNisMPGpfddEP/FNKGVGNs+MMMXYxpllH4lXF
NHSPM9aBBiMWWhfUCdUJ9AaLVb0nBcliQYvCqXK7J5+uVmcj+Vtu1sTGy8u3WbsAnD+bxSyHUTeQ
9Lp3w1yInFTQ9XIBDVCok7H9NTZql6AwTt+99GtcDWlI8S+Ejr+h5N4lwIBiuqAdn+627kGHyMnV
1nI6lvdigANNdursiuN/gZS1386Id/GUzZFIGtOLJw4sTSHk1VGWjZXaMELeoyOQYhkdKcgsFHhV
kkP/JgraLu5C/J2PZvq75YiRaAPaSJ8ANsM9VBmGE+/yPSeSIsE7owUY5LaobppoKFVyQ34vVmI9
RbPibgaWmtX108cwDh+IQpFGKwLoGtVI0t0Zc+iglblcuweGksuJbu/33lRJBTmH29giztkdV+NX
54dQI1CXM3rwsPnFmi2IO68tXRZU83z4iazUV0asU/8FsH1xgDcujfxN/tVpnxu8HfeGTDRMc8wy
sP9L4uRS/5kJo9D8v2mjKHLmU8quqgjuRwjQ75/iH8CH7jlwF+tnrmt5UjTjyT6QHaYNNQU9Ze5k
8BiS43X+KHasxTI8WeRURjfmteGMWSneMNG7RU9xldq3ZhTnYEvxlQpIjFX/3rSXEQH8uffO8KQY
u5y85B5RvvYvEFVZI8aMtvjAdFByFH9OM0BlDkGRkCdpOcllCHRZiC+LoLYJPBaTXshhQdTgHVtN
SabFmPtfBBr7jcdf0uAUq6uK/Ygo8ehqlZJVChRCiHrx1kXODwgSf7AspjxGNKFdikJ+aykJs1On
eKIPlQaN9Sj3wsKJ0H4A2aDk6vcGk+o/Kxj4u/ETcF87xFylcQOiAH5WrW7nfX7Atcs3/t/IDLvc
w+QulSA7YMrsgS8Vi6lqXHROgYBE2IT8+CClUg44IYZch6J4RFI3tkv/21hJ1X4H6gUumY/egfaY
fNhidKuvIohgxM47zYDG2BU3lvEcmutJFbgfsYSgN7NLyMFq39Gm9ZzrYSb9NeQak7VmutRj5S0s
bT/ITkugT/c/iaxMdPA8Jh+cpxgKsTkQLt9c5QcKTs2C95MB/swf5qWGBJdxVfg1T7OnD2bGSJy9
JzdjokX88NbtrTmSIfz25F7C/6og43ExSgqdMeH4NeZvuZukVr14Pe/xxXD+/q/wJxH4SA6/oZeN
w1sLqTee8AnYzlodEVMrpCPQWHOMxBfJrp0k1WpTpyXPxc22AApnb+E6S/3XxzTXrtoreh2cYDnK
/WcBNwXXTb4VG3H1E6U8GCM/V6pUuyzPoZLrbJ2QZ26vrtR3nrqUavQPeFibNgtlMscjvfAR7f3M
lqkenx/NOMtAWz2XtYFgOeIg8QvjwLYHR6akhn2ZDwG20+axpcO9qyrNELTFJJmKHsprzUHUmwJB
vUZ8MMm8VRMyt0TdgqMt/eAFVUd3YmSVmJqS/uU2NwQsbJRgvtH6uHEBQgPLZEEurfvoWvFwT7Oa
yIL1udgQFgV6SppvjwvFaA8v512H+MtonLHF4ObTMTcjyN7riLRorMcmU33ewgOjLDc0NpA2UfxY
miBC3uonvxZ8HNyxsSGkrcJNZFW9rOFQm26WkabDq9hxBBm4LRHQ/3VIFx1S0DC/rTFqAL+wm4cd
UDeRQk45lhwClK8Qp8FKfkZx7xJm1FBPgZ8Fv+zwFOR+3fdNeMGo5TeRCGF20xN2l1/5ZwGG5Z/a
tTm4pVM9qaSlJdttinkUZ7S9oyQQuiaPoEaonIJjV/WJYai59OKMMwgBGGZuWZQFYLwrJo1DuDfX
ylQrPhtp69kHC3KSsc8etwWlDgplIlztYflVbCOmfhatAVijEXCaXM/+O+oOQ2JIyCZvi4sfjHp2
jeB6K85zVmmbP2f5jbNt5cKk/LF+jmIvsU48QfS4rv+DQ9UVk4GLij1Sl5nZcZfqJXCXf0qlhDhy
GK3ujXK+drLR4H3tNS1RqayzNVNKgGaw8f+biqQJ9ePwkZ+7ze4MuvX4MhenmpEPXlEZ9dCAN6Xx
KwPkif9u7CADSw2OGFjYdnKgEJzR7BDAT/Ao/ToRxJzHO1KMPbsG4AijY8dUAiJ0+xJrUz8MKdEm
wJH+I6RlZET7H8WB9NEEkxspXvteZl2gPdwlP8sqonwWOchvUUBUtSx+CDEb+lFYU4eMyhEMb7yW
8+gVTBXDpQF0KfO2QeIusj51iCHDmXVt2PBjeC8zpZ3gxOH8vPTlhUAQaCRrQC0x3nsjmLVf/+6k
c9PLBrsENorIxerk1qUcMih8Bd5OdhLVnUUFBR1j1rfVoge1EyrdWG3B9IiR4+83mZCzpEy8kb1g
/Y1uGjmP6Uc5EOStwp2PyWutSm9b2sI5dYDpYSj0vP8wZ+kC4v2RhD5f1UIl2MjrvebuaHdgFnaH
/BquAcoZxQ/FxIePja4vlXeoV0du6QWpjmAfNWQbYX1oMMy0cOVOV8M4fQoFbIrGsIbOunH8jEjC
GtSHw5GpcvGEjucViwD265k3bXZZuB3H7OlksQYJ0YwgotL1ZxjWN9sXSzTH/9wsTACTWSmHhzSG
W8UsDzMEJv5Wd1aCSzwS4iNhgFQsVMeiYi+9t7kcIYKldee+fSHwXPyajYAaiwYpT0yXrj/n5xXJ
pf4LSXciINb/ZCr43pEDngSyNVqpJH2NRpcslsFFFoyZKw+E4TLU/1B/GPmkrnU8b83PcIapPQ8V
JAGR+G5h59KAcjaw7WusD8427+rDFvJ745n31cIPyQvFUx9VnnZxPjDSwqTuNoBg+p4alFr5XaK0
p5R80jAKKEtrkqLA8x8T5gjy6tApczggOxx0e9GrDuvH9yROJjEUgGFF4d3XV5UN54sKFZowEM2h
8VDyKBghDFATWM9tgMF4Eav8cCJFU0D3KaUJqzjF+rHYwACuN7FAXsssakZdRRdSdl7ruLIiXUq4
lzLmWKeSpDIWVKbJLM22ExaNOGNn8KMfX/ZQgurAdDsNCqBpMZOewhbXms536EcbOg5ZhhHODLPs
bxcSy/3h6v81v1EwROIv9yw2IcQo2T/6oBNeUvaCnEYhNhY8oj6pX6NQPysWKKLi9rXjWetzlw42
059rGQcAB4yRAJ3j/BYpMrbwaFjN/wIl3lw7XRw2lnXR4fZ3NgtCh7gxaz3ayW7JjyJ90VPCvezf
MzmkZwCjSPAJzUuDJk/lKvXCWRrLWngzP8ZhUnnWQrrzKqUlnDYx5ya0KI6AI1rZlksXQ/Su5G5V
u7CXhaNP0mMZGiKQURkUgfiJ6dWJbB8GAnBDB8yzRbVfFshnHgwiCmSnaIbaCjFfiw1clG4J6m4r
pUSuZh0IYJe3f7ZnQdaBqtWB2mkfOLnh33CJrQQYe/ocfN8KmB5k7UlGR4ISN5qZzzathnFFbPVv
eXWHV62Dqzp3k3x1fKcnFXhw3wOeOYF/18qi1+VJUN1tF0VnSgbjbSMlyR9sK74U1NfEb5h/WQpZ
Pu6IYkYTXI0nVYjcs8TTEKgLuEWn3rgLuGw42FS18cniKRh0lscZ/kc842QWCuPEIAUBYxE8/TTr
iGP5VcqWkPz85xdNQc2b2YGde3YmQBxKS0bv0EEfe6ElNA5zrsTgI/6LTsWYXD4fyo6zSOA8SBvW
xRwyI4GdXNqKc4vR3U1Lcnng5j7z+zLZOAgQCrfOMbkNWyJtPfKnLq/hW8pUnO4auATslNKGSUcL
8bpyeGSMKGQUSJdRbMZEpQY9xOLT3FYG13bBphMUBryvEmr9eiCy+raoycJg8AJ1O12Bvb7MPYh1
Xi5JvjRN0S3bTia9otbK02JP8seafxAqV/kw8207NgBthHc0F56o5H46nPxBpCvLXaIXVr7rCjQb
VnnMcK3hJcX4O1N29ZzQ+MduVchWC74pyBgqM+TxjazHmw2kTzVG1ASwqIC/MBudlGK37C71BUda
LN7GlenAgaKgXh/Ck4y8UnmwFVxXRMXeaTkMapk02IieelMUQXh/sNzwcNhbfUqUJTprRL42IvCL
XX/njpZkQG1EipN7TL1ANqInGuhPli0frb+Gqf6AAA+i0VPlse+LKXKyZVoIEtOskFlbKgJyJx8X
x0Fa/zXznqk97bez6yRP8du9PEc65SjD+IqGNT8irLyifDPJMIKWdQYZqeI5uQYd0uXEwzAXRlDx
z7j2UNXpXctKGJrJJZSj/2tcYgQYLEFGMxj+w2QoTxl3g/IyZMyO8E6A1ICP4PTimbyANPm6V8yS
IorxKO/5naKVx+ycpHrKwc58el+hw+6pNLytmTz17E8aXSwfRvZi15XkH/sl9MTc9SC7cusqOp1f
QZLdLq4AaiwucfyKgDNBwLiJArDr1FFdaAzmBsaE5RT6j3Om03mrC/q2RD5WySY9XDNQNaTrclFe
Mx/PLCXetoEQALLg6sVQymeeB4tNppONfQ+l5HsQv1HEHmLqSInJIuOOGAGlTvnRtpS9eA6SsWol
cSp+xdRpC6/B9CPQGsm9B0Kr5HwJQY9cbVqb37OQzb7wV1einscWzDDRvGlky48dvU5gKs4TnvzZ
/p9Rnw4HBffloiA0sTSuAUxXLfQLtX23DARiOKDdpL/2bHMrJZJcdI4dbK6Th+yQDUCpHGNN+OeI
5AJMoiWjeH0EcK8yohvYGb0zudZbXamoZ/ZYwriQtXv86+5xrAtXyOpSxVRZveMETwnIvLCPLH/v
FslbZWgA7tXkb9gtTM6sNXypGxhtSQ1DcYkxE2wsQ9/p+SG3vOLJF/+r7tPFHkFXTMnix8VOLLjA
nb9+0/9rk0XjpBc1Nsa7s24VfYMx81UFGLM3+4Bt1hvpkwx4Q0Xi31+1VM1nFnZTsShfeytaIs+C
+/o8Ful8isXZAlEpMkhtYpWcLL07zrCz6b6Pw5YshnOEPqeLE9H7FtR+bTV6YlP9u8T4clZy/sg0
1uOcZXSq54/wgEBnsiSaDBQ78W/w2oUeJrKU2K3Nw/ujtWpA9N8x1dFckZeVRSt8JgLyR49zStUe
Wmmp2ITSvJy1WXzMpZJQKwn3GuMOoTBKKqFUcqqy5KAuOvdxf987CXaDnMyzAYJ97JP+tvRKJrZh
57++f2mSQ0zf9ybRSD8MUdKktexFJJlI1sZljP321nxDiW4ky87cugQy0D8k8yJzVuK3HRAqV2A4
dTTax58SaZyuHaEe0z6RJ178MaEk0webJ8LRPREbaSjPpRMohNlCH8wdLLV4KhoS/EsByeeFpg+I
ZxsZlgkqmKxfkvkVX1WjmG+qF/9rrZDbhHi1UJAr6g2LdQLf0C5yijcOGpJQU/QGrysNuoevj2d9
Ms7O2+qLRqN6tUPnmciMYYZt+FMG3hnj9RDWaIbZwlp1Eka9vvbKYBBHcFYL+Fr8ItlCueRQBbjt
uG0vwV+IFAQ21R2oK5z+TdPxA5bN7AoXchAUnqIL0TqqJSlS3waTfHQrGHJzd0ytI6ayKxOLAnzN
xXSlIx12i37dsCxeEP1BQ5p2mPZZIluOrazkFM004+0CGqAwFjmgyyCLQe0V5AUMV3QqkTOnn1Zi
yU9uQ4+qwM2gtzxoWvGIucejV+mNcXdxTH4FeRmv3tSUYxWtqn+dLRulDCdKC/3C8aG2W72fa9Dy
0pU3gpsH41Mvudh2QeJqE13gRPNzo6Lob1A+bHvmJYmg7XyDeE6WRryfIrCmQl5xBXnV00g6HuS6
Z73xL3wZrJGvWpJppqlfKGeHzuNbb3XFJkUV01jNsJIPRcJxylOtlcvXruyyFLQSoF++nk1Vq0ND
YybGv33BFXa8wd3lNlvqVp+DllvdqyyDSR25P4FpVXsAMhgGoroPTfPRheYpkddAbAWTrc0H/dVg
e3IVUuFAi1m8HsOY7TXtpwr7ZAwx705OM8YGyKk19xeszQtXlNZdHKNl36/BnPcsmP9fC4R6O+jI
xn+grMA8ij5sCemCwVi0t2n+2yeuljFoTCGQW+VVivg7W68hbAVlqZ4XMgnMidPbiYEXsXhAxoYh
nEy+jcwANOqb59zS6u6l4Dy8dOsoCZ9VXObPccpZVL1pEeoYEZFpzpkdgNMTzsDd1PnqXG141E5J
tMpqXEs0bmpDbxZ/d8K6B93eFrRVtbS9XRyAgs3skFVq1zcHYj4KNCb3iWA2wZn0tRuuuhe/c0yI
2IU3EvtXXAdJA4Hp1Tma7tj3ONSmTQR2ZYXTppB5LJ4vZeDEDTPKocxpiRfABccGisJUpeNJ8TUo
X0EznvAjQeI9Ns626d9ZJx7j2dmmEOkucYRmPmQFNYuvx+iFAPkvd4nTWV9gDXdSvDaFZIP1FA4F
WC49GgngEyHfWeNn4AtqIod5Mz3e+nABXT0W3t+nomleiH55Ko60ARYTFMiyO/WZM43dt2nKmgTd
kgrLG8leiQD5kEAKBxTE99d9WexB6sE0Wo54OQ5NET7TS4ZCCD7qLrOBib4XxNdjfmHJhzjWbFXg
O9oXi4tIe+NRtPTydqMYSRENKIgbx7xQ2cH4/6PQugPDG7ynHqwn2gPCgajqYdU/Sk/ghPl2yWE/
3QLtr45SpZZfuDhk9MQnwPsFOnke9OX+SEw+qPDH3l3nDS2ndfs+eGFUUfZZATGRQNQ7rx3Bm1tS
Yk3l/QQXYBYzFqWHXFQdJ5hU48Qhgtr6jUFOvoxlCqJAW62y2rwIpiJ7nEai4HCr9ZoU8TjLfuAn
+EGKZeCPSDdeiO2t9I4vWlti7U+qwpQ/UeJ5w5AkG7P5FgCnUnPzzHeE0ZnZWvCukA13CS3G3hAK
sHxAMr1m8s9odxXc+yS2y9FVMIq3bVVY/2tOFmzhqMGAdzbHqj5DeKMOZMRx091SiCPXxGwzCphi
nZaQQfM0sP7tG2wlJ9LCUnY8oHMdLdz+5p+oQUv8YCCYNvmEtGzemAsI6uex+echYY19IijhVChR
R0sUyB8y5xu7Panc2lD5oyzvJuZG49pJQfGxA9TAJLOl9tdH6mImhmY/t2eJ3MLbg79KA1zK2Mtb
CrGq4XO87JXSk6pVDM7mMj8ozsTjB63OanWK6MCgmsFSTQKdIz5OKJHma1fFDE18CnPGiDAMmh7T
bwT9/V4yOBGty15qOX3hbmBqB2ttNNum7nznx/JXkOfI/zyLE7aBf/HjfNW7ApvAr3E2wGtJQMJR
AiFEh3lh497wUeQi7n0RXx+HIgC1JY5wgylvD/UAWtOH/FXHSqF+jl+s/Gn1iMQGLHFBkWAiLo/X
FuYJVuCC0pz/0Xh7joJm/g+nNt7+u8a1HjhKq3LWUt+r277uRemNbVyb5SihHEsGZXgEi1T+ix/q
MLcVjExvinDmbnTAHaDXjIuQat44ZFphw5Mf/PdI/ECwLVDgvHA6Hyk1yVz7UhDw63sX2F5ApHhl
hnPxR1u5HML+ENitoD5KjBkHWxFNOvVw95mZJFFaXio6ZIsgia2eJjw/6SQeZBIg2qPex8Ykz9dS
gZN17lC0IEBMlbK5lnPY6w9b1ksGSqpeldAcq/IFR7QLIUs42zC6wdPV0vJ1GizVlK0a2iT3YIdZ
nehzxIbWGyhCgZaqMMF+kK/JY1fjTleh66X5aJk0pWWIysIMfAhTkfvFDV57pE4aEiaYw4Wgq0Pw
Kc0ap7gqnpgdh93jEp211BrSt9VfcZ+gauv28wp9gvvsymjNMxX/susppWWQz79wRfi4znSH+9As
jhA0r1EZhd6KdZt0+cSmkvi1PRbt8qtZ2k27myCO8BpHSf5hltROUJgEuUJ6JS4P6F8MyV9lFsVn
zqsW25Q+375gV/X8FeWnF5hPiFmQl8nJNn65lmnfkXKuGQK8dCWWLNI8IImfNZTZ0HAWk2/PQEb0
rdeAUT6upzVFzgKTQu3yKZaf8BeVykkUvwPSohhtxbjLEFjnRrHudhxIIcqrVxhtpIpN9L+JlbV5
YkBMrEZyFV30lfzQr4tUTghbUapJeuIwI4RmOO60bAJ/3OPelZMfPFYAkCusPBXMzSZW4k3mz2cL
jyvGkUDOAbWqk0CHuzHkg2uB2PX0TWKShAv+QHQPaZrzFebFJoyOC3SJHcRikN6xitDkl6pCMVpk
EixsJYtoZMuSCm069uV1YjoLAyi6SrXYUWC4SPoHE6p47EJmU604YtnlsBreZCOKhE+LaMFVg6mT
UJ8VuXEce4WIZdexNxzeQJon9ea64kVNc9rFrLS+A5JqH5/hjoIg03+1f/JuoE89dzO241FeP4Jl
1lRoJLQ0oW9VRiBOWNS3BZryVPH9JuS1vwboQ8m2uNjNc1JtV3FMO55hFWOqQwiZY0Sg8Om6fZbI
bTERczMcYTmmYIGRI9yfLm8G5+2eAC3GE64icVifpH1IqAk92blSqZhn9MT8oknGt+mYDUr/XijF
aRFqRD1UCrZ+4LneRVe3bh5cW0lnjfb9OPMzmILFeTtj8zwYWjRthvdidZQHXpGRZ669aChTnQIp
HySUU2N6ovtVcvT+zm7nHSszs5U8PUGEM4492pNJtdfdUlzNdG19qa82L13X9ZfdxVthiaCOqhB2
4n6/ILpG7PW4aGuZyOiCM6m2oTHwbLTeTBCXbmEhS7cE364zx8Nh4tbLMrPlAToNOkbnZvp6fkvK
f3Gbt9K8uYlejAJX4jca0HoQY0Uogfap4oQGJTYg4KBUBsYiaLzbR2AshbD4X3uq7noDQjn7vIb7
fY1pJPlFCEay25lmTjCh29YMNnyOpIYk1L0nYJVgFtozPDv4KXhj3vX8jurzYeQjjACPzkHLid6i
hBmDEa/Mmfxy0xxt+dejz1CGJ0LVZJYbIQBlrv2oqXifZ8yuo2dSld82qA05AHTbUMEzuq7U6S1D
YKxuvKzXPaDaW7c6sKvnjTnGN/1K1W1AxD7xVEkRZm2WfQW+Hkf27T2ta7zmcfpq0ErJ35nd8ztd
btnQbt2kOQi3LLoA8haJ8olHt1WIsODM8rqAPxoFGOU1855ZfvyIp6cTGIU0ZvuwXRkcRxa+JG2Q
1T2q0pTNB+4HPYNoQ+ArZF1fFyjHwBIQYx6Mm/TJqdHT4aaBWfyCi2QOxHJJIk6RKraT9o4LvnNZ
x/kmVulE8l69OBTMvsuaO4z8KAlPJwDi+oCjZnmMJxFYevZo77/F0h8VuZS5Y00LDzuhKuvEvec3
NcTzdp1YcRqSzsuTn7JxRkK2iG0+BeE9vml9DnXfhl2T2qpBtFn6jZBX/PDCKb5kASyD2ttyFzMQ
guRpAHtKNgQTwFLTK1qbuDB+0C/5Inr+vgnjv/Ku1R+IvbWcu5LkEZlaDpdEHbP7LBjSIgSbcuYh
hsIMK98DxbYThrarAuqZiGkR6SpwalB35AEwzX+9HTaqj2YEz7zX0jYhLPkz8UdgAXC6lv9bdIn6
yr1v9elMgX4NEcyASijfXsml7Av+2nOdRAEnqGcWU1ICrcEQ5yStiXVqro71+Lpd6bJ9GG4Mr2z4
WjJCBIRVJLo22DHnfqhS3QtpxqmAbZi3B6rg1nBVC3fTyJJ7lM/1obvIsukqgoE/Er4fzOrIRNjj
KyO4s+H4FR3b0Hwn16ge9XkVW0JKUkPA79ydRHhmi6UgFQcFnYvyKd/T9+HscLoCzMJ/YsEjRbV4
xL5IN8s+Ugvfy5dskdMqjmkAsl5fWmxWFp9FVvi0fHz5Ug9D7RGvpp9PgJ5nym7lYc6hdhIYWuvU
JQQkmabnwSHa7ApYfE0/iL63Fo4cR0ObgviQg1+RpGlfS7ndxBe5ZP4oEIjHmwlw2Bn/j9vml+PT
lY+sM8q2V6MZPQ8qWHMLhz21pCaUMhlXJYjERDjxaan4WdY89KoKi/7mcXo5JX5CQIsRmcqaH5RH
qwr1riqur+l50OKno3RlVDejvLDTi6WaLT0nDRyIpcJgk90J85VqvmvHs6bRBrltFqHFauLeoku7
JX8F6vobHZzXwizwGObQsvJIAkD+WPP1nK/NLYNVHbMC8CU4bFnbNDs8H8BswGjV0BqTi52Oaz8Z
cdAIRKCNH+bN0X77A3KfZLX3gIn5ycbXZgjumNEKXaymUFM1zT4RqSDumxuttPj34lb61SuGMilU
m3QxnWJbj1V1bI2QWij8qsqLttnMvYNPLfWl+ZlIoPezSI4T3tmo+GnTcjhuAzoklseV/KwyXPOC
wDPAe2NQf5LFffhK8GFN99Yl+VgLM5S/ZxqzABJj4Y5vwRriOj04h9O/0LvpjK6sAIRAKPeAvt18
dnP+Rmzc9j/J/wWFPUoO836Z/JD2PPvEYUOeadMWciVfkAUQc0vLo0Hb5AQenXffzKGXYKJL0GXD
DXeA6tRVTAT1fe7bnJ9MJB/ejckJWIj/rRhf5s/Y1fmapzC1BdXfMxPg/1Nwlezu9F7cbYINL20Z
+ShzEYjsG8eblcdWgiRDDpuOoLjazaTv1cArN3Gi3/6jQzZpR0OFvCnIU6Mk29IMaYCC7+2y/St5
lSPL9RbxYu+SNvmhHlgq+pzkyVgMTAkqiY6klQPfj8zE2M9aKDp7s8BmttrDPhkwtuwaUf7Pvnia
ksxPRg29tm/ZjUKecTfvWwCbVp62ToC46SfHKYX/gevybeQu9/DxLUlnq5N4JzefXIVGGVjz/4LW
PMHAEztuAHO6Kbi/f9UqxgNNNWwR5mpxWEBCy1FEKpSO7u215YmGpxmhwtfbjGye5s90HLbb+oPq
2C6x2BdWHmOu0hzdCcFzsG+0CtA8RJIust9Rirmb0BR8mVzrjK2NXuRKgiDufhozzz2QuF20Yes3
FGGfxKQu2Z3z2Cl0MyBNC/w94Fj/bkFBniag2aC8+iyyHrjXVKYWxSyTuE+k37nglzQOugc+03pW
gB5cVywNFimW3GOIIyUM24xv+BSptH7+8wnM8mDnKdbB/ZT1lhx11srClhJKbSXjgZ1dWPGFNUZ1
UAXyeH8VzZi/lDL7G5XTZq3OH8osqZzNgh6AHcfzbsDHh/4WL2OXJ4gayxpHB1Qe22LjmVz7kU/e
g+piKlvper5lNZI9CP8M6Y6+5ZJHvbmwHJ47Q1xl/lZvb8/go62YLBAfWVyA42pi1hrH8vFMIFx/
BQj8MPI51zqHsl1CYFCXC8On1fYneFjyX0eUIleCDiP1L5XwnoZMOWKX5Et3gNtghNIUiFKq2cV4
6r4STsu7b2hvdUixbQt8nj8u/WLNgfEp0XNd+8bj3Hcf7Gzc3XBebENSA2Rc23/Xz8Zuf1GH7gb2
8DJsT+RuXZcqWZNS802c+7WSOXqCYRiBrmGXGiGHAX3fLyKPin3aTm/rMZltxSgbO9V80eyEcUxZ
KxM0UY5GQ06VxcXe4/CfJdzS5ayszyM3kl4cFQpmPGA3uvI7j+TKiUDywHVca+U4E3Dwq8l7ZV/J
Y8tFVn95LfYPnBKWCx/zh41UHyzkqA/sgvgPk0uvXNbP4xdpzTguc8Ux5ZLdprJSGt7T7ehh38x5
OXIWQ8/jZgLgi/RbW8ccB7u456grqmlMyZZsWgzFv274snRkPjUPjSN9qU9eeOr+nWoYKLVCKYqS
y8J9s6PN93O/tolM0tk5fV3rFC4xGBWTkRIugxlxQ1oVwVqpQe9lQE6zxbHOKCQdGfdtG4TRASE0
c6pRVpgjDTjZrevQ2QAV/JAD1+pzmjd/SuGXHnAuPg1KPH9TrZPRQjAFrCfg5sJZjbBmsxItrZNY
slgtTFUJ+Jmf7bOp6L/4VXe+u9KVItN2oLQ0sSDuQl9oclqL75QWh8ZeTzG2X6681EKzHIulHcuD
0VIwfs2MTJITp0tu69lkokQDkYy76rHNOB6xWhAM5CrlzqJuN/IAQW4MRAj+/9rAddWsW1az6zOj
25z7+vI0IfrG6N1ZYvJlgQPwPMms9PTNZloaYoC6IlwBVU5byi2zK+5/4jlkYlgcZVHJDIyAeuh+
FA4bHM3DzpYZvQB1dpfO08tZn89F8fi1F4+mDRaYkXFnykuBqP2GKqY6SLWB/aazk6ed0g6Ez08S
1OXF4Oe2hayjUEmv5eC7qqPmgPfDMSzrWi5hVg5z26X6gfunlraCqdeZKnNDp+nymaHVO+ESt6Gr
I4BP8u8w1wmJzA+NJB4gxXcJW2K9FAzTAvtxohq37b7BRBJhc7PElIZwxhnM9OgWLrf1oEqEU0sc
i1dkK5ptVOVNBpMtA7RMzEhAShPoihhKJJVWDbNb8WpObJIqNmV8Gx/NFTPLlgY6qF3+UxcmuU2U
oNoz0n4AfFoBEEicruVZqXHDxH2yvD9I1Zsb105ocj2cQFon0qmoBJG/Dks02CefOtxkafoblBIr
Jo0I82TD3BeF6h0DcXbqYv66FYISPoiDm2SZ/vqlbygA7Xk0k/oJHkXtBCnVXPYC6FcARIX6AGfs
jVT5rGPaqGgvrlJQ9PDk9/6aVI4Qf+AGOOtxWhNX8NiLJNKmU6udOhR/lL/HSfWrceyKFTsUuHU3
sN4V2Z52r5mYqqsGEUQPGGpUhva3+zWkNOk4GMEF1nKCnz+twDeo0rjyJPcLpxIIPUODb/o8a7Ao
qc6MoSPQF01dNBE5+sx1TKYZ9Y7IC45FFKaMAdBXqTbvmjp1fbEG5JwB7OKNQdu9/QIeqUM7O9Rd
zzo5BH6+vA+08xcy7LKOzNqCxWumC65SGm5VsDntN8i4s9T03ZJwbrkKI+c+ro/EYu5ogDhQ6ksu
E1JpMf2O84cfXa79dNYS7RRgjqSjyWNXMnoYFMtcaDPwo9K9oy3JM4BFMHtO22E2QU39WQbh8wCM
q6Wb8nGBu3wQdaDHq3eNueybRTO7Hvd8Xn1siAGu7G/dvdvuWeNjXGoXzyAjXB+/AzKRztvjSDyl
39um3iuAi5j6n8nwekrCIC6OQY3BwgV7xGiBBKKc+YAJzXEC3oJzAP9f1RYjC3zR350rhrf2KFOU
eq+enlrqhECSRdeGtjD2TlCgUdzuIZ6bHV3YORN3GUnTwpoz3UfwtTkib8wY4wIzYReYBsuviWHN
rJ7VBVByr35NJv+AgJB3sMS4gLFW/IiUUNDpZ5/lYJw27MpIgTFGt1O0i7ZzouK52aQbX9+caL78
mTNLJQq781FVdbXiO0FbHQi7ntaiJUQ/1mY0np9+WXnPq5Pt+62ITlkjq9kwFwx4RvvJQElk5btg
wOyBeoXO+NPiY0+ZSeMlw4g8ZmZJLZK3MSzclW5hRZwLrVO9iARjSSbWdsKfoCxlwQJAfTL/vtwo
Gb46JauOjVupwk4V2RxC6pX5JF+x8TEg2zWb1U0oKCwI6kGcFjLhqZxIurKcKyJarE/g66DIziyF
EObYG5yCPwl097mLQREZ10TL7OB8P/+KBq3QxoQWXa11FT91rhWZQ0kTi3zXQ5Wtq31IVbuwqhOc
/XX6RaUZIvzln5gE/XVv0uasijH7cm2/AfcJG45YqVKIV4eqenTeFIuMwYWVtfph0GP0Qudq/En7
Ipna9BwdF64ETUXR5cdk/tzA2GKDbnAaJivxSWn803K91Zw/krSy8HY9chUUBgYl9S9k+WNKR+JY
KOUId4u7TjNjEMCr3nCsWKQ6418dfcSgcMg48OmT99hBwKqist9UfGirpjtPDWI28xeSrLq0Plcp
OoVA2yVAvYw2GT2HyM000qMCN3+FKPvtM/LnaOie/B7oHSBXuDsPPltvewEX1AAwjtl04lK+i8cO
O7acN5rMv5J+t1QqjIidMUW8UILJ0JZl05BB92SNhgXffGHbJSMblvEbZjJ36dqcwiITFySl5eYV
v9FEJVywzYyJjGvUOtro3Jy+q9PfJr940GnBAMl2qgmbgbCF8ycPUk1eahwr+ovArjP3J+XtB3IR
82iIXTjyzIJyCWxPJ2VHG0r47TYTcDt58R08xWXSVS+KV1dvOPD1qea4T6CS7AMZhsyQXerjws0W
LMU0XQO/IOr2UNwOOchV5OGKZcguU7/WISRTDbaFRvoJ7YN9w3/Oq6j6UtgmujLN2DlwX4+UFq+5
VlshdHTVt/yB/NTClpJegwzSTtpbhwr8DJL7F8MDAoapGecGWtqgwHZPqq14CUkxnyEs+Rymf+GL
sRErEnqndxpn+oPRI9sM1jOp1QX47ocqqOj8TZPBUc+jb0TIsSElimkFv6zfWQ62HZ8ro2N6h5I0
1RicOfZsQbfbiNnMlyQhJ0aZBNzjmXF10L+f/f3hc6UsaMXo+MjIMOTlW1CmJdrJpPchDyJqMZPY
eOi3V4SKT7hkyjhNv7mquKk8bOIBEkOTXLzcxLNdZtKDofDoMBNm+aDFC8H6pQFMctYpwCRwoYEh
65/1KwUhcXQZBvpl9b97RtcEPBbbcU4Xvzb6244IaYRb2esPfZC1AQ8wOPoY/X58cuaUiifiVFqR
47F0oYOA4XMgLLlmMSSJ4Q8BNxaOmceWp/QbrB/z9DN65oGHt0Ya2rn1Ism5DRcmf9u1fTHrKRIJ
sYDDtUX9SKAZgpJ4VohgHlRoEX3984/W38f175f9yDDGSeu85H/SzyVKnssVNCNnF63c0xp7GtZE
zF/Xoz86ZtJrPnsWelBno3LGUECIy9kHdYv4ffHN34fuDiqp/tu8J2zCkxav0nmfm3Iyp2s1MLHf
kJZ0JOssOY48HsVq2XIII+ta4Wt5BircNav+G6DKSFbVS3Uto8LNVFzYMxwF5mdoOqiRJI2wPS/i
rQJHw0feMT22VqsKQo6IIrrk4BZHx1Lv5W0XXAlrdr9ZsT6l++rC1eTKEUzalJpfgRWH64Sr7DnB
JP0EYgyiqqwXWlNFYjGB36SGGnoXHICpZLpRAGfAQeu8e7YdynwlcVUilZSEkRQfG84XdLyd0Sti
2w5PzzgYGaFP9VBa1el7rgmk58WJcG5YCWfw+6dTe0XcpLFCkLhOKwZDNukRQDDoXwreq7VRRJKM
geEBKHmqaoaVWsEQqUiUag5BYrqrpoJiqQh0U9/OarpUkcEicQE2RabYvQAGts3MsBMeMzqf0uFz
bigOtPiN6x/KF7uPfhm7jbZzDFb76EieqKlyECHEETItNr0D7yASNGlm+dg5KAezcZkcE6K8wBxr
ds1FaF+XqVLpsQeXmsdhaxUeeGGskABSYl6DiYfXbwMpn59hRvOubzXjx47XraQZvujR45qWp9Kb
kzd+UmMXNN/QAQyGmHUNAs7GK/S1PcHleYK5JoprWOIf+/4kXwgeuch3mttzuvik6ron/93Hzut0
V1Ceuny9tGIIYF4yryeYly/bXn1b+K9dCYVvaOTwXUevNz6Z69Qu3LN1JySNBZhcveB/5i3ejzKq
lHMYWHdeZ+7Fvg4SPfwv9tPvx/SPplOO4UFX517ni4K7WtHaLBDChQePsqM7c6CYQfCWDw1Lpgd0
4RBq9OVydoWUqAubTiT/Pa19UKJRiU3c3FFRu/yoPr/dHoC67vKjHd4bD7/y6kj4gjY6PD3U36np
Bo5Bx+m9rdfj/Fb9KXl8O0BKjCJazO28DByZN7kRfe3cwYc/7vCI+QuTTUB/YhxG3t7lcVOpViUX
gqCgYDWtnnkmjw/A+rUN/GH5Q1UBZ7GrPccf3Gy3UjVkz5CFf0ZAzDuOMSBl63FiXbobGxySyY3K
irRJ1czupqLf/MrYGeIFakVWwRwEvfJL+4UHyhdoSkHrAi117I7pdMgIUzJV1joxbg90faBoxPv0
VD0iTJAqjIak4HduNkWuxb6CyjQzqG7h0t6PeoGfesZQRVcp60y3s7NmrTsdVA6g5tllTtKQGqyK
hVzzeLn8Cn/ahBht5tn5ZMuSUBAfZX1gwjzRXY3Z5y36XDiz2SWpwEQ1H5dcRUHmwOssJB3dAOwe
Cy27+0AvQZGwSS1gWl68WrnV+Vckh3FbQwzY6hwPW3n77eWck05tq0UPG5/4DauDnYaJeskg4I6o
FaA6vB7VMntPvhB7LjtILrzzSlSqJvmDMV7qy02Z6ABkcncRz4bD7lcLLL3m4eEgDZqXJFpgmQ6x
Ip5wMLjfVH37JxEAKq+Tf5pFbh/ike+LjJmU6rlw3dRz5tguNV39YGBr0gxypF5ZEKMIAwb2lgr3
KGDRf8MjiWAy2uruCsJRcsi9vMCplrYcGZiRkiFB2BGYry09HGMhgsgH3/zQ3pNKox0ThfJkHile
EYFbek8UqPLxE0EqzbHEliAk0p33Pvz8HPsaPgC2G5DcZGK4VTgVdaBBBTUC79EWcsk7vbZLZguv
DxoIVK1NSuxfvGt18itjs97Kh587iSwMKnuoYK0DPiG/wwgzuMlc3PwHH094iyrLcJxM8tIIrJ79
vLyMSfPmX9xU510iHGkL9fohBloKrVIdM0cxno+A8stXuHQjRmEQhrdNsxy7DtVk3jodtQ9hFTrN
c64nHgS2Ft2sU0/oHRG9fd7yjc4FaVqTl49O1J/vOGjHnddI3sNq3ap7K+/8vjnD3Zse9co4g76h
u15Gwomdc25xFcOguCyJGiSn6wf0zHQEqhuWuseG1mGSGbiIBFJDhJypgT17LK6CsKLxKNOTkGRS
pBVczeGot69RwAFowRHyN7HmcqtqMDCUkjg0ZHJ0nY+TLe2l0BhGumDi5Lrls36lM5m2fMTLP1F/
ksIKwz7Z2FqN3EE1ZGtB27m9VJl9ozhsHZWZZ4q9vjqpOOzcG+7biP9+23UIpHmOOi+G3y4B1Cf8
Rr+ADKi3F+eQhHXkqFW/NcOJdTzxNvr5emoU7056rAB2PVo3Oi/7yQFuVtMU7Q0DjR/GL0fSnnQk
U7zzqvtTik/nEBY6sUqQvFPPUjoqCdysanNQqNsje5XK9rN79QzrXN8j1m/Zd+WV2ORLooYMc3Sm
CdufVaLE7hkehz08CuwQNYmIgnaA0fZtQJy3IHKG234cSSTZugdtwwoxhLUQ8k5f6HdTJBULAzvp
7t9uXpTeYzubnlJnDnLjycXiwiX9LnrJCAsw4ycAWKbwzobv7eK0kMVA9YYBTakiRf66Xy8iThPe
4pnhyEFV3H92v0c8IhhvQDvJk3XuSSfJiQdokagqub6IdQsgYgK7DEO3kg7knvblQrIHEC7e2GTg
viRoieEZ3bNzdtCafiO1oa8hJS+RBCpkf47HFkO6NbPbX847MbNAmlz5Em+1RdNM/roonuAO/geX
PahZd1l00bN+pdBDLPdsypj0atYMgqSKb6qaFA8UVIQD0C+WqDXwU70W3QhaT+FpU+iCqVm6qYE3
UYzKeiMkKqx74a8ol8k5RJNg69CfulRhMcmmkwjJIe06utd2aS3F8/P4CtOxtRdfpOZJgDBOTQ9M
yFTYmIBOcGY5EEfTEDlMa476Z6QxNo5PfbrLgfGwngWs/C+PfD1YJzW6yeCmNCOyjA0RN3owj/lA
77FSkwF6PZQQzG77rfBIcJm2Rg5AU53X1fc+u1CNFiOU72ZpHZt8EhjYbLb7yXJrRVDWHPfRFkG5
OMOCHcPX/5Rc6qKylyByytReYjtCVUHIdnyKDAHbFJPZXAZK1wZSMKHs9knQmA1+x6xOnHnXo04u
ID43cfXQbJXAnuUxjo/xJE/1ri5ejlnfRlW2paKyzUmP3d60ZQcPvF9vgF3wb5Y4dnq2OQzka6c9
Fn43LRe8y5Y4XhJhdniOE/fz3FCJOYHMZES4UsKvtdjiloYvj+/D9u/82TQqoXSjnX6H7Izhrzpu
XZymzaqoQe6KaTxF/kk7inSvOFSTl+z/tKEX5WCXDTDX3j8Q227NVU7+w0KPQDbIjGco19Rq8thW
f7BvRvBc4K6BCrcABLabJHCJIOenoWIAViYuAlVcW76G+tammKYQuvx7YdhI60x9kvmfQBemrhyl
gB6+MUlyB0qEqsIoRLhx8t0oBOYaC10AEyPISuuMTJOYr+xkCgu5pEWORv1qKTqg7YC1olzM1nvN
T4FWG9bgGEppRv4Tfnf/yA1AcKcGSl7fcAVf4g9K9enJiGOmO3wiIn33qMfIuBycPaS60w7bGPU0
I/a4JJPJjdZ3YMFoslbesQpG2WdRKC0ciekuRoqoCQstqPV02jzA4ZKur0nhoiilui6QVlJzxgku
hcVRthqkTqjqGvbCE2DaeHASve7mfTesR++tKuremELWKcRg/nEv1Rtbv+IXQqvsazV9ExoXgyt0
BoO8qnsZ2RTurxDnZ8PibrNTHtNGGnw3XHK+Y+5NCmeFex51Fn3uP0oB2jE94TUa9Zm7PjBvNMZr
b4AYjwNCApOAfWEdsm7O1tPcbGJQP8Lh1fGRtQ17Xo5d+n9+8mwLtIpHocdbp1GBJt7rsIO6l/3v
xoWhnNN4MZy+OOW7aAZmruYA0k/0RZJsP1AURwhv+d4x6TOxt13215z+3DQ9QlVuTkAIlXcwoMq5
dSleXi/utCtZvxnR+u4mnYOZLuFZF3fF75P01RSjHRLGOHMdqmBEMtxB2b19E61QGm9Dys4P+k2M
Aqrec0fzUg7gr2ewA1Xc6KiX/pjJf17QmQTXnvT9aUjvlgTRKpN9F17bwtOk+V4yL/puqe2lsV3q
MbzFQi0R7I7XJlqxn6b3jKhTvkM5Q2MyIkVBPQbumrJe9L8entIiV7rmiGKj7FEQRFhv1K7woGpH
v++SGAEPdiMGgJ7weVGvyoSknviUb8wVevKrVkSiwlSxgdp+hFQjTuKHstGjoTBa7SbX4mYgBHEk
Oo80UtFeMUBG8Bki7mQjft4lYT+C78LQLlvqseB1yHhXcKa1lg8AcG7xjlwfM+47JrgiDS4ZGWz9
ZlIok3vkWMn7S9IUDOdUv2+oH1wxV8nqTsVO8nHn0vqC/ISjyVy8NVl+xpbHyPXCs2lu5SakzUlE
+EWLeTWp0+SDQ9W2LTlGdSTPlI214qtmH80AsQyUxrYyaCvd2rd/B5mJL/+ojuZL9AvVWiNNOiSz
GoZgUl0nN1wvCX8c76SzgEer++DmchMo04r1v28Nlhkd2YlRfCFZac3IN1xo6QPngWBuBg+1a4/z
40mm03tlWF7MKtgDj126RuYq6nm0uUC2+2Rew4h67ec+N/1OyZbpM1rLgs52tnc5U6t3tHFqHgf3
OjARXINRCs2stO/trO+zXDqIrJTgkhGgE9FNZ0txYbsSuzHS2auXWy3eraLEA/YlO7VX7OT2IlrQ
0NxHEDYwHFrTFrvrPOv2TE/Z1WwoXyeVRxnAyYagMZJvlzITVFnUM5kKNmV+4ZJaOXOOS73yuAfz
ebO98+k/13yjBCRZfFRgZ4Z2tpWSOtlSPZhVjn6yN/IRBXR9EZirMzaqD2zz+iX2H4HmHyXvkS+K
Nzc8k3FbRCxuw8O5idVgq9wmqjINyl2xRP15xdhpcwvKwj3io6OF4i4WL8uS6jWBthjCsGnOsAsm
nCmE/36kflCPGBROvZCh2JutD83YXTW6dgNp+IZ2tjeFVwVcy/l55hieZ5B8UDjA0RCmIK6GaLcB
x0wLKO5Ps1lKC9OV0OXaW45Am5y8SioEDUxRuVQauVJGIZUqiNdji/9Hv1ViDFJm81y9rPV2P5Hz
aMD9xJyJIc7LCTn1k6uN+swsC+RZ52wyWREjY/pDoiON0KAP84joEfFoMM8mdViEb/LocTMAzQvq
gz5FfMX6SFTjEyCE0PNl4ff8G8h8tbnySJfP5Dc=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity divider32s is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  dividend :  in std_logic_vector(31 downto 0);
  divisor :  in std_logic_vector(31 downto 0);
  quotient :  out std_logic_vector(31 downto 0));
end divider32s;
architecture beh of divider32s is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~integer_division.divider32s\
port(
  clk: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  rstn: in std_logic;
  divisor : in std_logic_vector(31 downto 0);
  dividend : in std_logic_vector(31 downto 0);
  quotient : out std_logic_vector(31 downto 0));
end component;
begin
GND_s32: GND
port map (
  G => GND_0);
VCC_s32: VCC
port map (
  V => VCC_0);
GSR_58: GSR
port map (
  GSRI => VCC_0);
integer_division_inst: \~integer_division.divider32s\
port map(
  clk => clk,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  rstn => rstn,
  divisor(31 downto 0) => divisor(31 downto 0),
  dividend(31 downto 0) => dividend(31 downto 0),
  quotient(31 downto 0) => quotient(31 downto 0));
end beh;

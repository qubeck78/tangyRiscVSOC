--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Mon Feb  5 12:55:29 2024

--Source file index table:
--file0 "\C:/Users/qubec/Documents/Development/ProjektyVHDL/TangNano20K/tangyRiscVSOC/tangyRiscVSOC/src/SDRAM_controller_top_SIP/temp/SDRC_EMBEDDED/sdrc_defines.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/SDRC_EMB/data/GENERAL/SDRAM_controller_top_SIP.v"
--file2 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/SDRC_EMB/data/GENERAL/sdrc_control_fsm.v"
--file3 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/SDRC_EMB/data/GENERAL/sdrc_user_interface.v"
--file4 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/SDRC_EMB/data/GENERAL/sdrc_autorefresh.v"
--file5 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/SDRC_EMB/data/GENERAL/sdrc_top.v"
--file6 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/SDRC_EMB/data/GENERAL/top_defines.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
qUMhFJ6RlGpcdLLbPJdukN2yuFRAjBmjPvH05Cgl+jB7vhI3Hw4Hc1aPzkhiWBrCERsY+1biy1cO
Nnbkj3uwBKL25GD7VailzCIvujKoT6eoQmC71/A2CtUsRXmVxOLYaGSc4cedPWpUMi8zNwmmct0G
MIASB0CpKqNwC7Gh58IPsFa2nwJa44KFYOvcY7R/s3Y+u9m2tVpCtfo9s/2MVKaYNx0hyQifoN3i
iUMJhoZpqqsMUMOOdKgDUwL07FaVbjJ7EaXTo0yTXKcwZKPk3fr1DuCjKDGhWQs3y+fKJhZAI67j
NiIiNtiEgIcig9y9tOF2WQScHac6IB1uGq9sUg==

`protect encoding=(enctype="base64", line_length=76, bytes=162448)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
UVpB9VHH+BpECxRJa7MDCfkY30Rg6+39b/SWNMCYckaS9ppRJTizIFZpMLlAB0NqKtwwNBi8srdS
JKSKS7IoIIBO2zFmNWGWo1VsDbyktxkWzMXA+vwNAfi2Q6XvENQN6LV1tNDJC3TcYGK6lSCJkLB3
KCuqf+Pp112eW9i0OB15/evzBqeQEZlGWQQ0JwDR3hl2BfVu3KjzwDrmdKWuBOqOw6vwfyndAHln
xf9oS4cj6+xz/qLoQMgR3D59WjwsTbP3hL5DArZFCbiJch9p2mH9gkCAO+onGlxY7SZedlDlsRat
TcPBtaJj6REDY1Qjp+VV/ofkl27qrybSxxToM+IJA3P63SDJ0JXJLRL7XMGhmDnwcy4RaNA6V7xs
N5B+Y/37KDtfMDR4qHetKM21AlXtVdPA867e7QG4Uc9eRSyYKT2jjHjj+zIiyIC2ux+tMiw5kCAf
Z1qPL0LoKPN7gLnTiuvMuYJWuBoZQjLcnfKnQGPEd95eXHK3mY1tBMKGiL2TqGyEsjh/2YX0GgUK
DwwkPq1B0SjEi7njh4vQvI35YAsirrwlkYa6KsvVR+7BXFamx0z5ZDUe4n5LenPGRbCsVEV2xlwx
IBrfnccA5jtRPG6VPd/xfq5dr3ugmnmTuJiVFY/yN1CjE/LgTdb4u7YXOkQLfmw2hoOKNT5fKP5T
5rq0zmYNpuj9sBLxDXUrVLOAhSNegnc18ppV/QoOWlxsE/hx6S3mRgFqELT3EFgyrhhGDb6/rLY7
nkjIXPl/PqVskBfPVP5f3fh5x8TK+KjU8xBl4shU4pFtY2uLuJ7pF089GT0Q8EzV/gLdYztnrQBe
dnRZ7EWuyVw8TaY+7//F3GERkY9NDmlXkOhGxrC3LSFBkmOIfLyc1qkmQIY9YFWqFn2PyqXqYn/z
JepcoamenfTwKcBlE79Nc3wXuf5hAj2ajTrtJXBp2NEJ1Sz+xlEg0YOp7vW/OX+ZRnaPh+Y8jmnU
BehWAFDMylkKLYuxFTwI9cirNtFFnpEt0aKLb5H+RWdzCHxBtdv2l17AZ8DxxuzvqF1jfKCI6dVM
9+GIbBzJvRj7Nl9bBDnkDLkcDmFzcb0XDuUduwaq/1D8MnjdRWbYG1RoNeL/2qIR2b3GBtYgSGvO
3oiz5Nb6obxdVcNMiNi1ygBIpDSiDnHEJLsCp64NlOwocToCoFn8yPmobTCzkJ9z0sxRTuczUHL+
kmYbPXG8tTBDPL336uxId/HlZToXKfQab/EbP1yPce8UL6vMh5+p7qL3qjF9hKgKhW72n8HkF7Vf
tGI+cW7d/ybWSUc1J/JnFtD20zdOZ/TPJF1kPLa8UN7oxeQXve88NMbYBSBTK99VsEUfEjb0IUEc
/FRyq1u3/wP9A0YMdXdzIVKdGXrmUGrWkRL4UjB1cVh5b0+Q28zwyEEreNf8hJqQoBJCOM11sR+Y
YDlVuC2pAmbsIJFqPbQs9pzi9fVXe0ijQ4Nvhq9hFjiqDjM08llrIO2/ePMwLvaL9nFGrX7pjmtC
ij37f85OE9SN9vPwMcUkEw7SoYde92qNI60H2tpQ/008DPgSkin9O2I0J8OVYAX49beD7ij7Ntgo
IO/AaW/HI4U9MdbgMwWfgDaTSaDqXZ107shWDlgwzIvYrx0wBFZMWULtv2rjtdhludkDKzpRYhtY
5CVzUFnwdqy24JXLOXiN3G8QKQzFmdQJKSuE60jQxug7t3L1k6ZLzllpibcbR8dBuaqwQar8L87p
E+70TrRzV/vehAR36IP+w0sXkAuKPBeHqBPneeFKzZk1YJ6T6u6mNk+cypdlTwvlLCc2Bie9p5Ph
/RLo3zj/ODdRdojia/pw99Yi53+3xyyICojajUmJk8hHhWcvfrndUi1dBVIrOPIujy2+RxW0TfFG
6pCLte/eUqU7/eUlXAkYP9VqtSoxw1WeuCRv7q2OYlxqpZw5R6gAb32FWalCbD8axJqllMrbdc0l
Jm4hUyrNjJHguov6IT7weRpkXVBmqGzf9+pJgYt0jkPPGZF5OpDvwlGZ76RC+D/Nkgl/RLBIY+4+
93FgQiqNRwDcAQqXOy3AMXA3ID45lOHJDxz7rk1+AMr/ryAseuwazIpyGdbJTp3i3grVHe6NeCaf
dNEZiLai2u3zgHlFvd9ku7yiVCAKSRkj08EEs2eQ9IpU9tqGIMOx5z9uvpfbSlkqADPgLIMNIVyS
8w1K7fElY4PazbAxrsg5qL4bu1ZlccshiP5D6+rtSNleg89JOIw2aHDGvtCzuw8/MtwL7f+YicTH
NfdjmIjDH8nsED4rt/wy4Ua/QgJCwuVja/0UZLrkmLQfW9rVujzSJRtuHRLtjuI844s0Dbe1qzTL
0BgRWsZT3yPj4YUmC9eFHwu/WNH4tKa3K6kR2ZODLAAJrpOEPKreioT6D/tvS/d9exo7DLvds4dY
LN4hs/tqT3JUtAD1y5I6LMCCUp7/4V0rvDMfgbinUcwEao6JTLAE1GlqnCxAX5a/PEAK7MeJURq/
Z3ldZmE0JHyfFSUNcEWoG4lzUgq9uLuTJqWc+6kvSQ7Ayn2V03/J3+vi4YxaukQZnXpqi7yNZl7c
xqOVI9m9/LeaJjIBW6Jx20+W5j+zytSffOySkivamuhDWTq/jvEsDOX/ZaL9b0WZcwGxo8fiL7ft
OF170x98ZjVG2F5qjV2C2UnbDhygy9KTDuOd2nmJ/jtTmJwaqw8uqZQriQzK2cJBVjICohbWnPEK
wmCYBmM3O+TjmqPTmsLmzwe2vo9hk4Fzvcj2H3/R0G1Y1FiBvY9xT+NG2GURt2J+MDeYisqLTTA3
4CJAHnXVymLYv5G77iAEb9Y/j91oyzFMe2E/+6y2+Sgj/2btyXliBgQiAWyfykeV5dgFXs8cHDQG
t2JZIId1e0SrV4FSz2RAMXTSPY1GP1QCck/oHqlkNexsPO2xWvVVaKQhHdxBwwvI67AUfGX3tGjA
RdwxTzu/cxGY+ztv1yGZbryA9mIrsxx4IjqaJY+/z0XH/c6axUQl4NsPGXw/8Bt6n8unULqhBaUV
xG615EOHMOgAme3/isGZVYblPB60tg5c/uFUQv62XW+erc+tRCImkm0G0zrAlqjxKVcOGBx15PDF
rk7u7SZs0NUFYErvHDluZFQ66GQympxS48SMsdKa3f4P2Cg7LDO60uzZFjqwRkeonWq7UYZWcCQ8
mDNKkB+v2RFbnnEfI8R0qybSe0aNkJnphDKOr2X01o0L5tLXombxXfvW6tbNMxUjDOlSVkiwAIr1
sesY8zlBq6WkUUPjwYrRUpzdNouD6YfLTeNMJJQ7XSN9EryJJGVmraXr5ZS60s4wUqWQeIArVG2s
gxe75x2PlpMgnIAOprnhHHW/E1qWMIFsny6Pdpa2xVIw0Lzu7sRmJy7pdstdFlzNOnRbjl6SHGcE
dN7dMB8rhZdd3RRmYfNtorpZh2CDgaRH6o+8mN6/9eKth6z0kEBZa/Dh3UgH6leg6zNLSl3GcVTt
FjKH8ZoUL9xgeJ9c/1AEqU02k1F6lKw7u8SEwZY2P822aQ9hRyPn/VYuBeXclpa4DjJJls3YwfdZ
LALLG0JIJEfomih5D3cKyTmPLLtWek3XRPBQM/mXBBYH4emnKPjWTTN6VPRQ0AAaezpTOELLusxI
+xongv9cUf0T4RqqPRofIDaj4vW96BVaiHLdvpb1L7VxiD2vJV+rEYyi8UGDH4zEb1v2hfkOu2RR
jDy93+uACkwnmAS4lB/9NsKnBdP+ZbGztA+LLwyqaXz7cS7HqZf7F77mtToFwhti7I4Ij6Ij9xLp
0yiKnBz8/TqEik1I712YuVYwRbGg98R4CeQWnN3jGY2ZZ2TM79ZtKj+QiZ0Vr0rfegWJwjP8FqDA
nw1nWfadGGE57WIV7aY23LLZaLhXoNd6lX89xgWQd5m9URNjS+vxaxOgcReti5gowhuXLCP9YOzT
h+7SpuciJnqwzXFhKe7t8wwgC0Bu1brCYqHbz5Ksk3bKQQM9k1gVd6a1JYkKjaV1fKh5v/vIo2mQ
HJ/ZiNjWbHYWReARe0h9I2MCrAkAJ+e21A7y4NXAkyx/Sc/RzzjfNHDvipXoazpYciHS+XZCsxt3
tAzspHqmE5abqWMrEEsUOeOrREFIcZWAVZuXlU3rVYbTESqCFk660qbg2cTzM5qF7jKBviwNdr1X
++sg/qLI8Dp6ILojPPULKdFzpCFLAbPf6ht2rTKcFHIGasfO9fyhDc0e6Yx6sPuzh3f749hZGZ4w
FUACwcZGIDjB+aavS9NR+oxMiqUAHzTHggoWXIYV8d1a0R+MBEh1258uATzwKghnRdrO6P35Vc4B
3R2LQDzrZGeR0tBrY6Ovbj8C4Ti/E4tWCzDuMQArYpfQZTxYTQZt1w7FRxwgUD4/if7yGZJ82ZaT
tI7ZQtkhHXXYjioD9Pwkb5R3PHypuo4wfVK0un9JngiXjqwqcTlJHzSJbnsK+nre2pFyK19tIENu
ewfG3kFJu4TxqPnAdg5k4MxEeFXpd9/HAUpS1D7DTDyQsZrfFzBUtwTOd035iNl3cuYBlavm2k9V
mNaDq+u3XrYeE9JnbX3KLeBI+EpbaYi1y/bni0jIdaMwkmikAeven9bU01/mhBNkAziGr4A+FnnE
zOTVivlfawVa/jwpHar99MOfuusdNJCA1TVG5DroVV4EP/VN3YCwXSWX2enLLjIlisl4kmHQQzyn
hmkNTOFrpZyUlBHV8kZiW9c7CzkCWPuFLnxydZZdkYdZsbPNOzEDSo+WUVLfjSarKSfkzk0qA7df
W4V/sNADaaoUj2hO7N9HITs3SH2u65yQZr0/K9XbUEf+IvF1Ww84efCfQmc2Pj18lLQcIUCp4Une
m/v2F5k+VjXFms3pjl30HyrkI3VLg3S27Tw6iRkD5gmrQIOb9jOzF/u/FZFK3F0uvbW44nHQVLjd
+RrILxJpK43JyrcA84RC8jxRQBSrwOqH5fJ91Npw7CZAZmDC7NpCes/Zij8I6osFlw3uzRJO7dsj
JmC2prdVkPJ2TYPnhZ4HK/i+DWwMSrZYYW80GAdP6kf4Uv1/SpitwoSgmA948lr4re4WnWb/wZdJ
V8uRFRQZR12b24f6tLQII4beiBZzRMX+6fqQcJ6ua4MlRwKM356EG1Yaj0plCYc+ID5vR/YqyM7k
CeD5JjodmsuA9Lid15Tyr1i6Y7oixt2sI8zbTptq4Y67D1QKBh+kMVxn8Qr4LyFZcHhup60EV3OO
hN1emFLmBQRF8hHoDNARuEqgQ9Xwwy1WBEgOUhkg5mmxpoNVQQI3g/jgrTvHyK2KkVKSIl3jXQzt
14ry3PluJ0dBo6DchpCtmJYPrCpyoLlCuNPVDOLTFwt10l+OMc/y1kGwX+Rz8sVWzFJ6zfmGvIzq
aZyz2wUm1XOcONd1U61a0oDWLxVPz4EVMrKMpTImZjM4nPEnF9TW/Fml89DBFKPQvppnb2feEb2J
p7OYGaGMDZ6aVzwOmJjFQKHDiBwdaVbUkoCPotZi38Pwxfj1oxC9nGcHk0JAtS8bZrwxHeCAjSZk
DVIFFL673tgmOEUk4NQs3FufAYGMTmgmhpPw1nIYpyYeCxdrjnrYv0gigyykFZx4461zEW33ChZP
mKzzxgB3yeqh4blANVMaG2Szl28Y9BhCioBzZDaKX/ACYxveK68HiCfbwzafTUQQrmexZYd0jTzi
eA8a259NJyz+Ijdlt8YxWJhns8OKCgy0ACvt/tnHkSur9TJ35WWRHZk+y9oQ5vOdYHBZcAcbBn5h
3LvzjgZPQC8RvUMQUY5o0A4ll2lQf76Lgv93yAyljig1ZOXPbJjr2i+fB1dA1DlSKIT/taF05+NU
a1aYBwKHKc4BsaNXBODBnwzH/063HItAF571IRlN4A1BxYxq6GoDmc4L9ec8WXTTeebb+2IZGEsW
3vWvPmpvUj6xzAwCrAKAg5Ibk7J3Zuzpmqjha7FOv6zu+fp4hz2dqEZpyo6k8AHncCoUYO0X7PZo
ryCAhP01TdwE9w5vYY8wC4IWBgLAQOwJgrgq9AGMMQFe94kHDlE8sCV80XDA4o06RJb7SM9HOJQ3
uPxMWHVaUN2CpFQHc+nWBrXyq7HMUvHzZ0tiuuzMhAA+tZA1PvXMuT+ATO6yEzaT+Vnzx0Hjhr8K
a+FqWj8hXV4tue4+TmCjp/9Ka9MCbJic3sHunFsfO2gkPZBvZ3UkOPI3utxKwlJzgSxJt7Sd2HDr
Gf25zxBU54ww9aZYpKv5Q4u1Wn5mJv/8CB5uo3IJ3eBrJzudqHgny1C0SCx5wrH5N39mz4FiiPNS
mp6AsIxtqW19+d2gTxRlQB9dJwN0ZtU2Bx6xbzYiHNeGwzP2wcFzArXf1TxbfRe3fgSdw2HjetOE
MoMjzKL0beJoMMV70T/JMRvWYhjG3TLGmhQkiMN7z1z1mA1Jf9oZkpKjI7tecvYOj2chjTBrlMjp
AAS+QfMGFxRbhBYPLIP/L9xe3AwVNPK0KStviwiODhNS/C0X/VPBuE09JztC2tPGo9x28H2nLuHf
7s13LOzzaH2NLfWMfdaC+WXpTf5CpedA4p4TxXZXrHk34uzplKMlUuTBIYy8qZgx5kYR8st/gQgD
Zg0hKDHdEnPGfCWrxAxdCKCqGVoQ6WjuaQCLDA42Euc3cXDdXXz/8JqKGHb0wwLml5K2RJOW3Gsl
0zCX9oYm0FFPX+RHnn8Co/Zn4f8OIKWIriP4hwXRl6q4cJAtdq4aDlt9PdTlogOszPHctKIQ5eck
6wC975PKsUV90a0hsKFktWvKaJGqww6yRbOkxvxoUBd4E5oypiy5SOE6OcSby4S8BRdhd8fuNANy
gF4FeYUP7S1cUasEbIaayzDYKt3kTU3DDWYkBig0anzDWCgumgJ6UVmXfouPlcD4BBjePNu7pwOk
4Tf+DkGCzQKBy2VmlWLvea3H64Emdrj0cwHVs1EwgrGldJ1hSUYkpTAuJhLvbMx0WugmEQruPL7c
fqe0P0SXxjXQNeDxBcOWojiihnc6t6dCBD3Qd7lZcr0lbPfII2AfpDwyXMnYiMA4QYQZSAKz1Au6
D8hYoG1ExA3cYYhfZAywjlCIGFuj7pIgSxmoIelWEGe5mtDI7ro93BQHXTNfoIDvNMQ7wgB731Fm
c7b+kQ+r69KOYW1Jn56d6uy0jTIEdehynrgbbjrt/I6QXqE208KwRV67DwoYc+j7exFeJBfBVO2Y
iJI6DKroIRZoB4E1BGuZ1KGIA+Zrs2raOksv77fId5A2YTfsJNe/GsJSHb0i6UOEoR4ldtT037sY
P7nk2+3ny8ao70XZPFoAOZz+bH1Y7KVgCCTErH1tS48eFbIs6AZBp5ad1cf0adgOozjq5yzGiprI
r1OPcMzYf/7qB2T1La1yoELOJwVIrPHXu1gihUrdxEt/H776+GhBbC0DA3S0wjBVjkxXVSFYggUt
RNeHBw3s5GOOKGQNz4liRbCE6LkbkrbSzraRnTQMgRFs3eJVdK51jJfYfxV04cbOlpqZsApwwfXB
dVmGvdr/1IrGwN026sJD6cY5uSgee1DFEvgLz4F8yrUI6gWkY/lomRgdcUHiJvzAwb7AojNFXw8o
itNPzWTCuu9MJknCUCpmRGFr2FJcaGTf/ZofYr5TtExeZvCrzV4X2Ja7+KByn4cE/OWL6hgIV5dA
zr1rKotGMCOimNOgl07u2gRf8dXQWqtAz++hx1D2uMGW1D4I+pLP24AeCdpWU+w2Ibkuw6+c9YSN
z+KIaGhY3tBL2L/gMok53Z/DDWz+RYwE6N8befgGEDRrL38KUYb6YyUPZEQ+o/yu+VaLaODqMqbA
Pbsllvp5PCjOgXrlpI6UATQs/etsmuBt6SecH8EWDdBIvhqhJLYZBRGaE8GqKWV/sUP0JJbziPWt
vdcdYN2Zko4C60eJ3+1J9Xdivg/OvN0jlPJcdW6kgXszkK6TyVH7RSYA0ilC7sEso8VZqeQJCmQf
FA3nIoMAVlkYhYWDKI0dnYZJsLDAmqIB4peCoYbGT5xd7fnYgjdrh1E1rC4Jv3outhbzhr9frfja
+ZjANKgfPMg5Qwpw530MYdSnp5vQAn5exozzRgTRFujHVkYNSEbKeFj+//mr682UBUGsoeLdXe1h
Yb2fpy+Ywr8u2oWOHee0sFKyIyUeCIT/9SizZMaveNnUyKNO0KxBNGFBb6zsgIegPEXZyFG1VfFd
iFytryHOrhcZeQSNm3QF/2SH61hVN8ucaiY5tSmIkuR/ssjzUN9J+4SxfI4nX/8Pj6tFwbB8Ge06
A/Q+B43W2mDzrbWbPjxz7uS75Ed/zBX/IGxBjeZ0BhLQBEQUBFF7tKRFA96V5teoRdDMvbVyrtMs
046MVkR3L1mlpRLi3uG5ad1BbMfqs6Q4WwEGUkadIAAUI2XbbIBH/8EpEDmXeRUtaE4VED41PHKH
8jR8+q6VV2uKc3sKMsevJOCEgSEFbM0HO6KWEQqwmvlQV1Le3umpAGMK69F2BDZUA8wr3qMouq7/
mZuSDH43omf99OxFXhak8e0vAFHxw4VsUofCJBrOgucFRGTajJaqD4UwQ+0mJi/k7ONeVnjhLCf6
GEKd/SWS2TI84PLR0XXIGY8Hr3mnx8RKzSF6rcWaOANZtjdRyGdATGfVEzPu+loircHj03+dvUSf
/1G2jq3bfNeoX4cfa0g8BzDkzGeoeL46NpC6vQ+LbJWHEQiow+TuoovE5EQ5uYYC5dXzkCl1BHs0
tkMzboz8TWMIZBTYFXe/jMw5F8fa45y3HRciU4T0S1i56sE4jYzt1vK2n7tDrJzvpfUXI1uyfyU5
pLXl1Y68U+AAgvQLp9DN8Alzat0q6RoyHiEjesaC6bcK/KlfcVrWTwdWRLeY3xieWt8265xFAJBy
G7ipMFy/82LMApyO9N+a2oN2dSK8Mio4VwTDEFkG6+VwRheZUW7JdJAwK8ZZeJvOjMZZAvQbeB4B
hq5+I6p3zh53P6fQnXEwYKKLgCBMtUSCqPzCzzGQ6pnn8A9HhNfB5qGeLG05Bwwm1psLoT9FIAIz
Gz6PCy1R+9e6Mso60WmuNBddBUjfMTNyQrK5LWhsRpHshxEIrzkS0pSlnqCyzbIGavq69ZCffSKk
rtmaLz5EZ7wOz5vxqHkb7HqAxjwTq6RFx2nLOAkrfRpCXbfa2NFjV7m31Tbm/pMz33BXNC4+SxaT
+6VHJHoPmah/hmPlhfDwlwdcjI3WQ7kJ82oHvy0Mdcka/Cixzgq7VdoKiXN4nylnYuq425yt6OoV
h9E2Zbl4fUWLtANqte0GKiPIRzXw8rjfpUsjHeoS2anhLq5KDAlXE8VY9++J7SdVl4NUevrvsUVM
o3EJTahNAE2K5TZjFvGcsTrv+Rthb0qklGprgLzJUs3xMPbH2+foS40t3OuPIdJM3KIVrmlSNGTm
tKNY+XphnXaALdt1Q76y6xwMemYuDHn4xvxdWwHKS53krPATwtjU1TadkBtbFhov7rvLPzdMuBSJ
4+OAtVMWO+DYl5vFNFoVUpLQvElD/uZZB8Hklb0TzkT8xg1XP7vrDUC/dE0zBb3kxidQCG21ZEwd
dHyEARlSlNC8fUz4NRDVI6VCgoKaQYbVbu1qH/4cmFKPVLPVEu7MF74Oe44o/ldKgnRsYxYmGDU6
dkGwheywdbfwtndtmvj78i4U6BnW/Z3Z7577MGAqybDthF9w6qu0Lea+YktQDtaHUoqXPNU8tmt+
fqZAeCgWzrnlN2QRE1PCmMu7kj1b43Q1T2cxHS+TgIfgUwaSYQ+H/TMO0r2s5olfbCmU9Ba4zmG1
X70Kb+V6EA+5ghn8QTfRR/dgFvmrIWlheI9/SLUy/GXpTmZUMCYitnLZtUksqQZsfNyOyvyft6Kq
DMeGZsw4A/RhQxz/ghrX6jzaLDjraZQC2lMSkGfslko4fl/+mGQ3+Zpl8ADj16FSSBRO/u+4/XRM
LQ+V+sQ+boKSIL0ltXm0uaraVYBdnNiNAxoAnI19Ap+n13ftgdf7GdMmnKoExvfwAEyO+NnsoCRo
AVCjcKv6Uy8oDut807Z6P5brWzJsng/ggmwiDo4xH+YmT771QpCNfNLGIBDUMo0hWPEB4T0OJygH
CSxrMHh3I3NUQ/uVgfCCGwQ5p/yOYh+sFVgUZ4eFxQeNeq/MTzD5YA+37oHt1I486IuEUkhPw7wO
qvif+H/4jcyVpgjxiQ29IU5WBfGCi2COnBeoqyYfZLU3WUoAJhMf4eDPXhCaQBn2kTOswYx+TqFA
aH+usg47Ub1xv5HkPda3TY6tmqMscYYaQWNBLHZknz8E3UFmH6UTyzxsZCsnvRFJIFXBsO53Ih2E
dOSXcaaGsi3PTwHnQW/8PMkWZxwhdhfgt/kjIttAY+j4VhlDyZf44lM20aAhjM3heaJgD28Ehv4R
Jj/fb7AqCXY4rD6X2RB6nGFP6gbMxOsqhuGrzMGU72xbYS2CBLf/PhPBrbhzh//I/etm4OuyWL6w
3ik1AMGYHmctQyD6ZDX1EuZ9Ut4AIW7/RDKjIQuFmxcwU1ta3bF9zRTZVB76V/xuDCujyeXpZTPx
YBRsw8KDTEbAkwArIJ4E8rgUg8ZTZ86W+ngoytsZ7gGfKOH8ZhfX+ihOuMdgSigQcw+YBBtD17J7
JrHto4LJN8n0F6R9js/IK39ZkgvWqqqOYrejy3EGKYLenSlLYVW51ntGSlp9VFw2xKxVCRklccHO
t827JzYNxLVPEsIOyi7rih7Y7dbq29mpRODAVXnSX/IPKeher0ZusFDbiAqfwJSnFOORCJZ84hnX
hIokz/UgItlWlbiQTtgaM+uwY+EQdHhu03/lB1wgijHN25F8k1BV+kCENHiaHCT3AzjmucaTYqJf
uNDosunqjkQexMK5dilIXwiDebZz2jveMFiWOfa/CwOO5PhWcaZ3QDV6h5P2xP0XqxRauNS7RK5x
HFn3otxfLX7/OZXsvXMlBq/E6eaR5s+RjDhmOMlNKrgCTF7dJs8IPM9LpxEnyOAj2t0IZxMdybCD
6V7IVBoI2rNEOd+O4MZA2uSIj6mlNL18/LYUboV3M4KvIZqylLfdwPeaXAGTunPdDA4ihDmNmHEp
yb5MolVa2fcn15DDSiXIv/+SbA6eGpw05oEeF1R/K+Iee9jlCAq1iYBW6Phu4KZI7Idt9q47Ug9t
c6TqbhCpQc7iuznOxvA/XQKVXM3HN3zNWkTr0oorvzVguwpph2CLkSNNFsi5IDnk+oWe9QR0n18C
j72tb90V7uXPFg42A3n9SlbtvqG+k4PL0Cv4YNQ/F5nuEhoZDNE4G3mU90D+8POjlX1zxeJIVhPH
3TrUugdyFoziA8gQoB5G4dYVYUdgLjixUCc3Vgw1Yic5CuUMPgF/LHhGUBDYWrBkYq39QcOIq3ke
e+1rgAHxVIWHyfSPtbZAVABShKtWlmtxHfeVWIC2NzT6ZMeR64lk49XUkDD14J48NFNeKKgvZGZb
BLOUHnCiVqctXODoUeXXkUuWA4nGvdZ8S/MhYTeTam4+XbEytduGSndujQxmTsUnLI+BykOoVh7A
ymRr0O01pkRkSw+wCuKAxRt4HAKkA6OwWDPLC9CC8Po3YrXSejc+I8FAZuDzcpcU9DDTUDPE+hwQ
tKSoGB/9VTXEHc+1b85cIqCvFQUgDPJNnzqt8NKNAlPIgJTjCa5nvSvbZYNm+A8ZU05DyKXGAeWE
gFROt6x7fZjGDcTQGydor03zcRkZmoRwDcERC75YL3P8pULuWdOUdcKPHcqAXTmn5ro0cMsANZiC
Ru0FLyl1mRrtdFoaut2oKVGP4EsVYcXPGWuxqTwMIEipCyCJIiAtdT4ffCKbHqTi77n9K9utAf0K
k1d2WybW0gFCvHO/WpecSn+3TYdcvRXWxxUmGtBQTDi/fsSm01XLoczgklAkO6S71+Nz4s7W7dfY
6qTTHWE1D5+FTC9+Yi7gd36Yjt1ScmMM28kNmEMlaOkFaDEErCQpNNEJDcfTdr8NnRynGPKCLMds
vyywQfQEfVgpYQVFuW/UJeiQ7q5prIW4/fttLMtzymVJy9SLdR7XHw/IYEkc2YaGCf9IWP7sGlpg
7YYZ5aqMV8NTYMAfFgyifnPT1UVYx1+wX398lKpU6kVgWlWpoMPlYmSQ6BBbLVAnzg9GJ1hah4n8
u8X9hycp1UJ2UU4OxpqTP7mJMyokq5m7TYjfv5sW41jWKrtckIqvBXS2TbQVBzJcpo2QqpOeEfqb
a5bo1qLtbaTK9UNHRt1WZwcpeMO4azwP3TGH/P0fkRSTPeKgEOzgmEO9c4dXNgsc7vkMz9t3rhSz
SxGbcjjd2eJro9V8plUjcpKYMcMMv/SUsF6+BBQmGmFIexCTYK/luwGwYzcrsSl/qmpuww76cbYO
J1GU5R3s6+43fJuanAvVZB96UTlimqzw7wD1lGotqcAUe0q4g+W5yKKxOoithnOpjGdR9cCU21Pv
jvaQjhFugoKAf2OHXgzYx8NyOSgilybcdAqUiSidtk2Q1sQq5fsuqJ43piNHF+m3HM4Aw882eMZx
AZvPlL50k4oQeLSPcYkvNjMOntiShenWSspUohZhXOX5rL3MuTcFvq7lgIOe07F1ChLbpXZs2Abh
7ZT0kpIhRH7DA8EA8ZhRjmB+nhHt/prrMytch2swQja7ryoj/wkFkg8WCFLLTqfUkhegoaq9DF+l
YBJGe1CUKrSFc0GuKmL44iaIMmJcC0eby1Ld1uIf6w9Yyq55c+fP9H6shZycdUje/kJ1k/1xehjM
Dsx1lyM8BBuQybMjvt/2s4ANj92zDTjges3SDYZDH62BJu0JXdi9JYbSKkTXbBXAf3qOdPFg+7/7
WiPLAfgxEVUGXXU4CXCKiIsW/tYZXLhvSLTvVGhBb5eA4abq8SYmJWcgLE6IhGZU1G5dm64v9d5T
Q0kCt+zU5lbp//EvJ1AnuTb8Y3/3AZRLgx4r/KeMVXgqagnEl0qpzfiNtLJ4rL2h+O14qHgErJFr
/XAbScZKCFFWE47J0nRB/XB638+Bm/CihZhHabsBkVHEjhf9j5KjQl2+b6brwLzvCFlh2BiGEUX0
OHLvd9bbVO372korZJqnsjudOeWscp+5cwb7tqs/08orCQ5E+8Tl3zvSNErkXpbFgbnfFc867Ks7
nV1crVWJauAPNPLn0oJCp47KaM76E2Qay2RtUJD/XNzefmqovutk3GJlmrjX4zPPh9wkMrgWm5wA
Xu+K/kL+iro5WiLYVZbAUs/JZOiqaDVfuLdfygNLVbBRsCGoXUOUqHIYbHKqBqlNx/t9/j6ve9t7
pDvUjVWJzGv137RIvddhYo0fe9HJ7KEbwIEFsemJELHM3kmaVLK3XKQGEnx+4i6+EjsooEPXN4GY
ZWgCBrj8zbIUhXs69MyUZf4GBsxAVQL5Zw9p4FGKVINBwAaNFwInj/AQv5+tmGTTwmMxPtNPe6Jw
S/8dXDJJapKACOCB2huIwtKr5AQvaOdkxyI8iUkM+DRaqq5hgiVJuysnwTcDMZZGZ+kP9UaAXi4i
SZql5OT+YGKXILkD2inE2K/ZkJihGFMv06c4Xf5GbcCm2pTGQO0YU6G6/D4WVwTmAkCauj+0rN+s
0t+Mm02ztIGumQQsHzMtiJrAkY6iyphshqM6NGcekkJP07LfuxOgDCT27Z9ZnOJewPopLUkSymdv
hdgmChNN9zkJS4x1vU5+t7wzarQZFLmAQEDsQVgnOCIQO5ddTz2ZJM6gfpeC5SWC30/Z/nICe0sg
VRslrl1bGi7HyWLtpkPybASxUOMbVc3ieEi/VlvQ2tyMCe5ekyk8xM7mWhmeQvmYPbwtb0OANZlh
ixuMM6ZkLomLuWVMIZQFVWkYQK7FU1HzE+kmPtdkGgaIej5UW2SRUUM03n0+wa/AQ+90LTr9bpqJ
WhoLdqLD5L+knFEIdHhb04z/jjcUQQ4MHb/M/bxHcDPeMR/0UdJEIXt9lI5poo/tH/9p9Kh2gj9D
kXDDqxBg/quzL/E5RJ4vbEaoBNJyPuP8PjON8Ii0FQR6yyJX78SL58ZgVLdg8wIsP9Vu5RiEKDoD
c0VKNCuwrqkk8QGhSzFc6J0BPIQQqgBK0bVYhPrKQD6p8GGgxRHvKvp6pS8OXlZfAB0RojlwaoX2
y1etIh2LsaPRIIHMaq1nBpwKc9gbux2j5zZ1QLWsdxpsSHsjCf9Fs+qMZoXubEUQrO5NDoQ8uK3h
AdxxdeIOOV6t0R2qdg8NqWFoj7NuZbXWoIByyZPK+shTunAsITJ1wE0bE+km3daWIGgt181bCI4B
8UpV0CzZ2Z67rhCnPqloqv/wugQtMmvT7wCTHZQh7p3Ys9Pk76Z436qMHTeFKe2aD+aiWWbGB6ld
F18G2PLW78qrK1/UyHHBoExMkdZB0oOg50cbOgjXUQtT0hlWHNrVyhya98ukAPyiKAlPKsGR4dHI
zP9nFWIBbXmvocNbrw3n6K/+ES7x5OEdsRK7zNvjuf/vWDM/WY7H41sWg+lGkva0Dv07cYkUMqEN
7YU7rDqnt8Op1GuIMNmoVkxyrGvkjyaakG9MACTEwr/uj0V4UkRLhXjQlD0kjcfULifVGlmp/625
5k3gwTkuivp+5Ai4XqDMv/AaYTUzom8rP1Kyfd5H21XNs8YarR1tD735F1fYlNRPaYODkMESZ6qz
dmeXnqpGJsUgXwmd7XcIjpQnZK3c55vP+EmuguoRi8ehXDKCH+KeibrOUC5Vmxeemp8VBPUXdpSB
nDO0mvavKn2EzteObd1Fj/UVM497FN9i8wPQx/5YkSVIsHFd0xDbqWuYgPRRDisawkrO6LFEyyHc
ZZjvdIzynOuuU+KgaLG/rQanFQkxQ+mTWIErOBVeOOwwXmD1GJt4ZzmvLB0DQeCq260ruttCpqIU
MbEJ8VjDjCOmozbvVW3EdA8/CgP335zdEFXviMPw9dRQHRasTB3jgeQSKmzg3Cwf9k2y/VWacVNJ
ifw84HIg6/aHxou7yEqcxrWfctaiM7hHTUwwD5blyltjB78uQtPw5I6vi3Y6dIi+fYNa7uiPZ/7j
3gm61rtIYCLb5xeESrs3jQWsYoIT5kKQzdD/P5bcYc6V6H/6rcUp1L4439VCiCxTMR2VoJz1vpdA
9LZe9sLuhGBKAC843T0PJzYCFeZ0YJqi7UTfLMBMT0rv+jKgURm2H1/mjjH6XKxPhqZE4CB56uAS
ZfwGtOs2Kd2Alr2OF9nhLEJg709luay5nJ3stzTV1fq5SyTzxEj3LsgdUk6Wn5gik/LxNdAcngVZ
LmT2Ovm9zOibcSRpBhgksxAgXj5T5sfFYnTZu5INMfff4EltB6rwPUbDqF2g+2/I5pDy9hAsgZ77
g4nmu3/8pQzysNcOVhu1q1n8n0TpUuIKyFf1MERCjg31YaC79QSlg4iufd55KTuOtDTdyFFplz7q
msvg52OGXD/HS5nzs34aQIWZlq9Db4I8LBdfg2J710ZWzoNqsCmG5RzyMxT5F/DkUkIU/lVcm5fl
uWM5RXIEV+1RDHn6DRIuMGFQm5ahLmeRGWz1qMt8Ptme/xFRjOV9E6PQx5rRict5VKFyHxNMG3aV
YZdE9F+b/3TsqJiL3litgGTIFsx6bIRwQU+J17/bfYMOVbqCxOTLr/Xyl4UyAol/VfmZ/2XWk849
9DDzePn+Bz+lPiORrUL9bLxGU2xph7wYpF26AjbeiH80SXFQ4sJNtfTzM1MYaELKM6EMhL1YniJB
XolVJenKQFUHdj4N7A4AvfWWf0eN97qnqgxWynmArx660F3BUEViowuQlQUOqarLH0nHl6206Isp
Wh3j/O7IiDS4pCZs0fYPnusuxxeAdQ9NLPC/BuKp0DnWxu5tNEweAYNZxztkcXlPhOohjIM+uKZy
3hxui26UqT6Y/u/fMAMGeNCO+UbPG6YG8mH3Y7WFU8F7YHIqOT6nSlhHC8wHVy7Z8Isp2QewPxxj
UE6vf3FRjYd5Kpic/ctAN8Z/Kk1LdbhanDR78akSpB2yKG5/ZWVxG0c+7yxuGQH8gf4vX+dKA1kp
vsc+MMJgedN7/miuHnw3GAVkwrMmQb7cFkIxvULK1J5CqgUsZ8HHkdQhzdmdB0DS4RIaUEddj0pW
1JR33t/sq+TFlZG5TKMktp5OlWabr1NFOfdgKz/WkgOqAs+RlbkMeEhgjFfncYuPPaEyy6glkdTX
wJyugdrFuIGi7pGtvSQHBqqI8db3rDM8zLLcCfZvTM5pnl4c8xkS8XMP6eu+STskn6LItZjCB9nt
bu7b+xIzKmaWRXeafCqvGqmf1a88f/HB99qnhy1CVDqXfGDqVHGwyq/YHdgQDXUQlDHZKFeBD77t
SQyZqgZPuZsuZimZogajiRCRnyEfkvwpfdXHBKB7GMhvnoh12AE79Qyqq9cBzg9zAgb+Ov90j7L8
hd/HYPL9UQpWCOp3ymdM7lZA0l3MABAI+bnVAGeDKsqu0b/llfhCWqUGPIEh/LUwg+ehKVF5sf7h
rlTkBNihG8NTpRjaefg6OaFUNZoJ0SZGfFaRf50BOPiY4F+JkkLPxh0sP3poLz9i7TRa8R4v6ZcB
PmgVpQJla3ZAwYT+5Jwn5W5dAmyJ0CIoXtXai33Ozq0tFuRQuzUD3ohmCzCIzoy0Nih8x+GAOIXm
432qPWaSjRqulpXR+jsRqnfW12rOW196ZQWg1USbhWtXIi+v4ndMVgnnbIsYdArqAwmwRBie46r8
c/fsFKHjU9hDQZbFyoEB8mw+c4Rs3w5a3aLlNWmrkEk8OkGv3XZkqQ5s0+JkFqoZp/gKGQppssiQ
bokOo8naIgUjzm4JQl8HbXNE+2s+nKxeDgR1b9OJsfMSJVEPo74XGj6WcBOIboBI3MJDDOPc5Czu
2zUThoMhIz/DDiOB+erqtr51clQ1HTVqz4hgG2TFINOUpTKgijrwFjrx4yD8yejrYTbwTmkZQzzm
5aAFTLXu9hdMyXeUOMQRXzTc2j+1qCdmSbAEjet1Mhz1Uh3RuhYARBkIePJeDyGb4zAmLMcj0avF
HP1oOpyELRuKDR+CB3bV9860sijiM9PPEVM2s5m75TCvZvlwG5go4LeCpAkF3yQzauIceBhuFEzM
LXKj0mosS5gUkoG6LrSwy8ebD+kh6whXIfVA/M8u9De2hy7Ugo/lY2knobZgDLwNOzZZv+3qMdIT
lmcWJQbPm1CHOTFtuB/S51x8YA+Hd8qo3hL39Glg1e/UDQ8yh35w8OUtRJdwkdpHXkFxs+G1Z8DN
eHEvN89asos3OZjO1q4qECjSICIldwv+S6Y05G/emMhzkjcw8YNyZDBOOfft4IA3PsSoF9WFklwa
fuVYYJnjyXbfgNGBKNIehIS8nSBohh7ujyiuZWnEBWvRw77XTgnhkcSuodY0mZlkLjW0ugrot2lT
FD3t+Bus4wn92YlF2Z7KMWSBNqXXq1GYZaCAmEQyqddEqbhjOrwBZ4UWSbXDDowYfiqKMnZDX/Pc
G2D8//58Fujs40/RV43Vh/IIQSC7oohYiC7mnazZeb1k8RSEQ7yvsB/G6ggSelCmM6G7ikD/kCDx
RoqVizdDeM7mlmE4x2mueE7BwrFgEXjF2ALIW8UCCCa6eVAN/OmRRXxPCI4gOq6DnJ+uH1T9eze6
vL93ZiwwfXrB6EinDPyq913idiqfBBewxuV0W9mzRCikWqFhm2J3JMe/EBsqbvojU818J7xI9zm+
1ImFzYnFF3cepnCbxH3riCLwk7vyIPlCW9KfWmUNM+dFTgZElytlBqfvssI28Dfj6dwrG+iSGUsS
1dtkixxW1C3wnhNTilhzXL+gFyolN+XHgQKUfvSxiTQhLA90tqeVpiaarx/wKXayBbNiMDqOgAtJ
slJWxyXa4damHec6ggoYHT43gKIWDsCOoBI0IdQ4zbVxyHs0cOq5cS+m/ZfmRLPlkiTsmJ4qRmxK
721Snhg7HrwmteDUaOtL1olg59ib8NZJTDwlBA0ExOpXPehbVxbLjz8E6dyi65vriW+jh+dQgpPH
W4lD6JltLomWanQyYeq1a24lrbTwZB7txY509gtgQX9fS8E9OULRCYYj1mPm8NwQAGCqni87D5RT
/0BYfdC+IRDXlXeeT5YftEuGPTonpoyfjrWvkxSFOgtmSD6hqCRRoj+4WYy5kd7KOoLK2xSwWIfk
vXtaSrQWucrfUCTDXGQSrA4megam3iq3Wt1+nc1stzlZILxNKX6BJBEf5SoWmhECyQYl8nU11kCy
INzPZdSX1lQSg18hM+vr5AtkRKb8j4WYwN13CMjnP4ADAb8qhClqFhVkigKnVp53aLHCWFJ3YuoQ
3OS1aqljHceqHBHvJn9Wvl43ATGhWVCJPm9ftO5LhNgjnCkRFdCAvjbbAJaXb+3KNEYdy3vmyhiQ
Ck/fLJb6fdroIqD//om+2S7X9za8agFbwc5x7kT2McAOWAOfPvIHkaqXDsVJi0kAr8Ru2SQtH9Cj
pvSMgmoIKanxunXS8Ys0pkQq1HfDVRyvNeILztoIoU7tkZsHPtFTz8RJeg3VuwlBV+N7ZIpbtLkN
oBgLnyf4FTnxo6WCLKPMUZi5iXKVTUj6ahOLC/pzQLS2hrXnbc1H7uc5xtrPegIkR9urh4Swwy0O
jdAT2b22acFNAbdOa1l1CZ6kLhb+r7qQgMEtCuXFAOjIrVcHL2yGX4aGlYMJ2q37jhwUjqL1u0IM
IX1CCutcO4DPaItzSgc5HhAuNCp7yL+7xMYJ5NG+/5DdOxtoepuSoF/xsOPBHtn36Vyq5TcNElg/
qReKrJWCpDDHdXN0y0X3H20H0id8mCVOZJs132SvTKQWc2UqUBd0zME6pNNBB8WmhvE4mPx75yDC
CTJeE6/t9k75Vdzpu8ldINTuxuzQIcyn20P3FI3sjtxN8atabyuTAgNi8fOhfQOMlRGIXFv4GMYP
NfbOfyHb/FVzj1udgc2wqVsk84FxhRpLpoIvyngheMIBqSaD1XupApsiEyvVbBDYdwNs+CB7jmtf
e7BU4XTXQY/ZvfOj2Co4vKp5qmyTntp2Y/QVn1y+Dnk0v28UaAc8uRp/57OdCLDl8rLxd50mRGci
k36n5RUIxNhvHdU4Ilfs3lZa/ditAKR2zoORAfjxLwMmK5R0fBMUL25SrrUmP/HVT6mf0KXeJKV9
j8EaYNwbLSozplxVStIbmIjeOxeSG8yF1BOU3IX1Sxn9dkRXbQlW6QetRi9Gn20IVwIX0u24Qng8
m2seMzYQaxu+4ARMPrWsEfRBrR3ehpMpOQMzlqrXAzeuM1d1OaBvHGytlpyKYdGZwon84NBNJU5R
b6ZjrU2dzVVkc/rIVq6AM2JdBj7qSiVu4cem7v5fe2giUXF6VvYMUOOVmbUoygJc/4igWVuksaX/
u9p5+hr12bIu8YPzDx3EX9/2p2ZtJyrRxCvFVSivVJHBWPJqRZ3Hwovth2CaPFnZtaQtQifJViJB
hBCI+7aN0J+rox/Q+0efUcvqGJOiRJzolhWkj80X81ekxmCty/Bp6RP1ny8fc2ictc72hBE6Zdgp
7ww6BaFeABkeT78Rsc9X/l9QCiZ7DPVtqFAekBNnXxtlylP3fz2O1md8TxppmuOdQvbPzkV0e5Ta
A4w3Ax4nQQRuyNqnsEt+hDJSFLOBVAQFaU9acSj0pYN91rbRFkhtIHTKrJdt+4Jp8Azn0hFvA5eG
Z9JdXNsNrWZ85ohSHSy04xWa4K5qLfOsDilEXy2Kp5zQcTgcFCrb+WYC0R+fGyoSHqEZax+eljuj
XqVmZQOuaMDBE9rV/jhpVsyi4vdwBlD3g2Pq4Ne2eV1ki1B+1s3Ci5i8H+aLNaNS4orNMSblNolx
1+PWB9sfOmPvgQNaKAFYJhv3GqrY8YNUo5Jvm8Uh5PMKSCnGun9TbVfcQO3hqKQs1X5Uoejil1DC
McEFEoCycJLixgLLhMqkIh7Q9p4zKHMoQK+d9iE5sVXS2wm32l9XH3azZV6yzvG+wLqzFPpsQePL
2gg7df0lDBs9FSimuiFz/zF2BHXkNI1zKkuNcu7pS+n93wTRqXDarzWK7EAxJTR1VyTW7SJ07RkV
a51KA7zmsbqPp0d/6oiKtfQyXU6yRYjLYC3PgHBKpJzKeRictPpVfam/Bz0umJEDoN/ET7pTtz6W
iEjhn/Mh6Eq+HNjRJNdzb4IkpgJiF4po3WDs1o1Pbyoxafz2lcf7/LtH1lN245lzL1224Q+wJdeG
udquGUfzPk9F/UcXrUNJBIhXV5Cz/K7hBgtxUMHt1QkXd6bDhj2GW71ObHNMc/7UZPRME0YGDSPI
BBVYR0JKBFdLR2loo+3UP94PTmk4hxE2ns7EKQfQfZQYI6isK+A3JlZbk33exU5I2iIUn671SR6E
eBebkEh5gLlAJhFbByhIMVT3hYjkFLE9q1kUf31Yngz0xg1Q05IAMhV5wXouI5Dm2FUO8i9N++xT
NxFbRbLsFTF6r8VPpH+qNawj6YIVRK5FplsomQhUHuJYCmX9nQxNS/YUrKYsf6XCQx5KGpDkbnQl
UDjGuckUCH4YgVl6FcObfhaQXpDP4bLwWVIYEKHquRCrziXHLwEzVZA/simU86x+SeIhlY2IRf8/
n5CNjH+fI0ElQuJ5dyoy9v+45kxyg7NxHn37aOTbNrw1LsbnYmJCd3q4d318Wfj5KsGicY2TOCeS
plC+b/3Hwh+PIO2Uyj8OKU+I6VNNpVCU4sW4V2ayWmFFvPysurveZxnWAhDh+fMCzrSjaelnl501
L77p2hmSWGm2IlofFcQWPYH8dY63ItNasfRnoxYLQ0/tWsQndqPmvJ1l88mZBKP7P0O8rHOgeOKL
fe25LDypV7gxVQduOjv5NktS4j8RX+NoVRtVhIodsojTtNyOiznPd5lCJQuuk65Jns26CGU9UAX8
LFwkVA6C5VdL8mJRJ1xdy7CIyBGogId6w6gtl3B3qVGoLeoF7jDrHGiFc+ZxW81PdhCiweD4YrJ5
0wq1uDBGwxl3c4+exOcAn3aDfhjDzowuZrLKkwwauntrM5WIyrM44DBYRSwh1kRZQldHjHTdmpSa
jr88hR16BpxPBeCcbHFOhfbMUgADKzIbZy1sUwrQ7o4e3yS/2uVR3XxCyIYPHa3tf2CUQUB4A4Me
vcz0rXfGxt4Xdw9UJI9S+ei9KXF/2SudGxkfPL/7G6cuUByVgoRd+FZYUbgIX1UMmqhIpcl3dciO
bELFWMalBWdBRyRzofdJdfldPYE23rLbGQBTd0ghSiDkTdquwi3OAl6wan+QedXnk2C709x7jFOD
QaplyFD6EFOmGEVIXycFd0BuB84vW+y+yeD1pmo3idw9xipwI1UnOs6dZ6hRcNxaN4S+V89zcQjx
1PNCXB18Qc1CQRZ22gfGPqa1YB80sjntdDK9CqXqXT3ji4Updo3JYpN3DdvsHCaEdPkpi2xB2JoY
kslMri8J4OecoM3e5rY4pX5ds0UVLiSn5tSQQMVz5QMAoEX4MA3K8NIwp8e9gfhyUa65Oudy91Z8
Erbrse6MphOQTyBsECK55flNXBvaVLP/aFc5gsmlEpmyGd6XRwGViJyJ4RTJ4+mEq/zxgKcdBsVV
pAwTrNGDBaJK9sOniB+PbeNHPavih8Uo/6H9u8yIZ2NDL8So9bszU1fNQxFHUfYLa/fzjEvXxE6g
DgNUpBVBM98rVFSH0+L5c6P+PDwByQ3e0euOzH/lXaBvGL1oPehLVd81jK+zoMnYj1ARuvi4rwqL
yGsZmFI0sxxojkGGZYpFk+S3scuYzHsvbXj4G6qaDns2nb2XiGxF/R6P7dlRzly4Nn0RVzPxhDXq
l9PCFMeRSSVNn/R6345KCPOL42AOjRbVSmBpdD0gu2y0W7aVjuI8iZ48E5zhoW/5hCVE1bL1oTqs
dYBmeztCGuSeCFhx01/xatP6dNVNhJ4GumcEG3b9xHuk0+JgH5t/ntuUyPGFSW6xCgFiqMS3b0GL
qIqm0vStk8xHzHe/lMzA0H3t6GmyB/3usGriHvqwIhK/xqpsDu38ChB51V5iRMuGJdZBml87Sio3
wlB6ug8DABbrJmuJwebnvp0NVUltD8VtQMSmoUx0YzAKhkLWSWLzzbfqq9sps4nZ9m3ItF6e+ccd
oFxQwb8B0TnTZJKVzUz9aN7v+7hjBTNBgWxnx4sCQffISQX34jzSXha6V0dAK6pxz4mJ3oWnsoiV
9hv9zjTUojTMpYBY/Q2GaYVeVJMT72xPfztIRRBQElTYPgQcUeoGtKziZDRRFm0+BcUruNWN6tDu
FWtTMuRAVgQrWWJCFoYHQwAiehz/9709wnAdz5vdSWaxs4HpOn+eZFJ2AwCKHgQGs/9iVoXF0G2u
NKWdkxKIrrGNXoJcd5vxERcCufmNezDF2+wv4aTMhiMaHCA2LWkc52no9k63/ezGM+jBcvExp18l
LUzHHfDdX3OdVvzwc3haicfUC5y8tUrZoejJ2+8MWSp1nMT6CnbVtA3GWKKrgyu3cJnzfii4Gw3C
w4dziW2gwnvyxhMikgRbkOj06j+JNr/T0sMZtw6Ye1GWJ83WqgfDnlM8OAWf0m1yZRywT5otaQWd
WQ/zTza1JSuRmdiqG4ZdElJIVDdFwCZ0DnqVHE1CSotNQ2Hd3PehJ3ySlqix2gbimWxVZEHNzL5k
WEWB0pskeaaeromHQYEi7ruqOOSFGPgyOkpoo65V/5nY9cQRGrMWLzZbdB6CM0LGZr0Wc2jcJekg
2or2roTjkYrFazH3yyktRWGAuyItaJADgOvLXmVIn8JUjswqhPmM2wCi0cfdRWAbopsIajfZgAsi
kQ2h5XmQ59YHDQClfxnZciIw4lEPSbU8W0HWe2qjkoXF1AQ9fDaZ4XBTzUR83bMdPhtPAXy7PEsj
/JeSzf3ApjMixzOKh9IgLQSnFOK977fD0hZaGLNstqx/hcKCgzbysOXzIq5HRjNsZ9z/hwtOjzER
s9xMHo7OToAKL/nrSyDaf9uOKZhYGi3GJz5Sbnafqo4zL+aHpZFly0hnWInxrvkF/DnflUmnybuK
qYHVV2CqGiO7e4N2V4SHYXqvo3g6Z87GOdPWAxbElTJ32NJ8nSexGHPIJI26EYGKR7PUW8Wj02HV
94i/WdBhjUINldXdZ/atLU1cqsE8JZx4bZEJKnAMiM70/9J9z1AT2ONk1R06lvNFYX8Fai497LCR
s43ybY2ZR0eeki/ubX+9VLdjPthsGl3/EKIBaxO3CtjtjfaDIa8NNds+g5dAoOYIeghsGqsA6pyO
kIqpSIzs1Ww5WyDNas1/GHZBbwtpNWWd3pNHXtoT5uBHSr3I94y9c2JRCnU7rbAxhMYSj3Forn1r
oHVTaGKnNasNHIp7eVriDm8innfCM8i9anEF6w9oyRFSaqqC0JoGMBNZ0I9oVNI349dxcJGQzIHc
TJ0NNaKt0seC+y5dvS81cxmOw5urCCsWbGJv1cbrISIv3sHi+KZMWBnaGWVFUf/r77utaLA9v5+E
nLmf/RW5d15P4gKmm9Vw27dgjlq7nRmFGxZ7pZrq1ivSJpB1poGaRu2dNgCwVLycLHjmV1q68uiy
G7oF4+sF1QkUdXdT4zX6RoQDYaDM3jleS+lfsr46CqYacll8ZWAIGoz0fk/mkZ7gSlJI09Zypkdy
wKhi3bSNwWulKAy+NU2aFXtIIMPv4vE8304OrsPcjGOdm4nDN+ZI/PffvMccTFoF4XWD6YJPVL/b
GRW62YcBlsWpYegQ7mAT2OPEnsKIddPoQHWtTWMH/8WqxIZ8Oyc7YaOCtI/5q0Bbd8LaVDn0vgGd
WSRk9Ypsf4l1lXIWgbw2kfHEfUErY4AWcRXtlRWXgXaYKBkep5WKIxZMVqsLgu/XYpC5oa7hx5in
FnO5eaqxZ5lsXJuBHVcoWlvPBElV7SMW3J4Bcv04Lu7TKThfAXyJ7t8Ol6nppjrW1OmSjGytiiuS
JVWXaCxUQzTE93bp01cKpqNdTMloC2k6zJtUNaIAn7XRiyFD+XFw6OWZHJi+qxCgwDcBMAU7bQdF
b1x1uFrQBTYgCQwkr3I42ZALLccz/abkabMPHVr7jcowahkOSivIc5pqItQq9vHzNQRAHWDfQdX4
VA/RWXnIgebyF+GFA1RsEZ0ZLzXV9LZJS27Pizby0snB0maHS2RsUAJ1/VARdR6kN3tf2i9DIx0j
mIwDYLJRM165AqE/g8+cB5W3+JGfsbY3W7ZVjHA14vuSrdfdAubhH/f1BtssfNs4bul32SaVbUr6
p4gH8tJV8Kcbma2kcqq8Yv7vaICkeqMmGfwl4dIbgWCl4cy8rrgoNflBpxQ79rZDetvkJC3IDkHF
Ppjklic5jMhoqSA3PFQo0UDgoY6GhBvTV8zb7hZh69JvMUGAm/jkt5wxHBM6VvuWO7+s47GJUUv0
AxtvqOEhwKmlR2+8a3EP8aPfzidNnUfJ7jYB448aa5LirVQewNkIh2NhimE4HPsXdhKtLWX4/ZqP
lNyYRYRpBvLcZasdblsZo6t2PJOaRlHFeNANc8zamrmX/9MppHb1Wic5X5d7xNdx6K8O6HkhbJSf
o9jRCDds7CWTU/No2owXO0jTygWqwKYG3UqYbvVRDv8tGOc4EJIXvUzuYatw0pFOStuDPGTNK+ud
pBZwWgsW5MzOUWfRXnUxTUCqwM9+mDM/mwOFV0HdvbHZ2Ly0PKkwI7qFy/9OWAtVbUpmTI5ZFKR4
JEA+IUGpyG91uCLhSzz0ZO+rffhB2dMs8SIRsbKtd032gyQ8N7VkYEUjGIfc/ozJsUZAcJxwcmIM
XfhcaaCDvklHp7pGV/MraJtuhuSnzTFVSrIN7udMqOUCvu8/7ctHlNZqzA6cblQrvjkRNMHDB2V0
jPlvaNUIRFLakePHWzerruU4Rq4vMFm35L+5ZaTyA8zfxMbuTsyf0DO0bW24iUzDH2YEvx02tvWg
0OhU8GCxoY3+Y/49OxzOuY5qy91Sk6HESW64oqJm9Y1fIPjBPTD+rzoS7QYrevlqFlWHUsdvS6Bo
E+cKPbOtCPUN91w1YCT9OGfOZnWHNrTDAFOGUUTnbxpsW+4MYWte6svOdSYm3EWH/ne9zYR4Zxpa
yWDZk7R8UHXBFMjqEZ8T1fl1VcJ8UOgW2e510aF3vyQ85XSD1Qg9BPYT257Hm4x8oLkK7axxAdDP
sArlS0JSYiPPv7H5uHqdk62jXZBlJ7mww5IuJT2p0IdNBAChB608JI+n4xFljG2xjQzlyG1cuJji
u4tiWejiafmchZDL8CDu8DKpoY9bGIWT60KAXCh2/Gw1J2ko7LV75/X7H8qtxDDuLiVK3ZA6g+1W
GoLgjYFYHMBCWoCn69fArS+MK66Kc3x90G9UTzdBUPL4FruzUzhoyg5vRJCXIdShQ9eFCiwQZuYZ
6XDfjeI7aNPparcas79Wms0QgnP4cqNXn+JVwj+OzRv2Z/M8kuVOHt5oaRDFXqZ+ykBLpeMP6Ydx
SAbP2jE8987+hl6DANl4rsgoywCiQMsFfjDmRyedtLd6+uBXuhO8GGtieAp7pQkURs/pwo1GSqZ9
cN67v4d9aColrMYFXWwL/HETqtIhgRDhzX/OycfhcS21m9/4vI9F5L/iUEvEMlRVuMjmZtLmw/Zh
ocfccSNL1TFj8PyfvyKWlI+H+HnwPdwc4MYglFGaYjXnO5FSoL5S7YbvBS4zKpxz1I/Xp8mQOjj0
MzV7TC1Q7QrIq4sHcYy7C4b27IrrIth+M69wHo0krapDC1htAlMVrxHtMOhvfIvIOFQ44alXoSR8
VfXIg6vefzozRrPDIOKWXxDS+mUfoTH4TubmoySWpRYeklNpAenEp3MhVbcZ3j5tLbLH9waxiSm9
qhtE3TYIYOcYB0L49vNj094Tgkpr9vXzX0x+CmV0lTRZJ58DevcwXZ63k3cHnGlJf023ntA6iAdl
+jjyB24xu6vny2GgE3gK1xE+QyqATnePbyvVr2YXToMS/7Hi7yLtslH3n1jkZBRNVKpuulD5xNuN
A2vBR6ashmisodhsMXb4Of5+yIAzKbEIT5EYcCCiHTv1WTEIr2fuiqIxV7BgqsU/O3nNCirfUtvV
Q98jaLXzr0b1D8n6FTaP72eNOXqkMWi5Pl/qxTSIHjlgL7YrPxKiUtofdwnskyhatJR6Ou24IXax
XZaI9gvn2mQLyotBEF5P6D5K7DFEWGhMOgwd9NqJYmdpSkmWi6USuCNXCdGHGzcO2adI2+aCmmmA
JqQlQeLHqHTH3IBbBSBaviW45oke+glE5jfehSBEOeYlP7yJWCLwwlNvwtqzftrhMsaYEFd94SAQ
Dd7uyqc0XuL3gBv7W/ckwHhtJ88saf835n6TLhk+ALg/xni+pXbegJ4C7kbTTRFpxy0TXeeOPnrh
cBdmqYWe4KHoOwGbfZt0fholGy6XwrxesstIvvX0cej7SSDmyNRaCvyMpPyuw8HpZsFpZ2ihJJZ/
kg061JCaOzPxyfCterTORrkkCo4ZlqqOthE1SL707mG50inEd1VBYDWlsWu3Dt2UqnBBsN9G/6Wk
Czp6XCFSOwuaUv1BSPDUC0EqyNJI4TTJtI0wqKX3W2vGxKx9xXE5gT8JsKEMtCIEncVfogwDsouZ
SwQ980RmMR1m5guodM2tScabi+H/ptbKJIZwMr+GBsTxiS1w0tY202uqyWqjjwbCX9JzcMtA0pp+
+1LSl4bqCd3ah/6RCrQg1HHxNoHy7fCC/shSknjeT8QEFIjA/nKCPoVaw1OhpCF3Wz+7mlvnmNol
leoGb0e0NoSEqphRq2eAAOzaoajMcgR/lWvWt7FKHuRYdniM9eyP/SeB+nBhoqYPs1rPQWXnV9wr
72CiaQJV4dtR2KNljiD1eaiiH1xIDgboN8uWhuix7f4Ymhh6zrTjaqg5a8KVQRWPyLiNhP8S77EH
Lke40kuFDeWxzsLB9HRIzR9B1aI2YsIbk28bhRDISZR8Ks2nN7utAIfWcQwBYL3rGMZ+2J0sbGXv
f31GGOdTQCEaNdBRFyYiDHXOP8BDcEbc448pfhz0s26UGxfF7oOAG3wbBd2mAHWH5D87TJrxG5MO
gJ+A0c6sfmqbIiamfexghXOuLOEPficwG/Z6TtXwSSy6iNgp0rFYENL/QWK4jr574I2l9AAr2MZK
H+L8RjHYEYWxYQZ+YNhCHyNbtFpRv4g3vIZ+qAsUL2IqAL8O7i4lEt+cM1OCeNE+7PqR3TNcXIyT
SE6eRe47mcAxuVAQ19yQHYAr56/ShnOQlv44ZQADbaU6pB1x8hGp9in4Geybsx1uZ3kfHtdg8B0q
XG5Umj0v6DYhCTmG1LL+fognDZhMLQ8FwshDMAqFlG/f3l4lnKE5M15Uju9HOqaDvAWiICk8QFCx
PhC/DlVgw+DQ/zCexig1LReBm8Zh4EAuR0zXbUgDJzbfgn1l/Ew4ervRbylRNFmO5Miwi5C6+5g1
16TOzxehojwQctH6zFvJ4KjuddqR/pdCnAL9oP5BgDTHHcuyD7cKm+50FdDdSbELCCL6WsNWpYRk
RSDP/imMJWj0SBCA12tzZ1u4f3zzBCas7aJU/jmi2rZ5jwASXiYbRJWYZKxxRuWHFGP2VmB8AVqz
X6A0YoCpOMI9YmS8tpgs8qEHLyqIqBMZfgb9h9U9XRji6XiMkGcebXHoAaiGz43GwHyaIM6SCLib
h9btq0aIUPFs8Pvx4eInW6IZi9ymj68JRnWloqYIgCPRDHJEYEjoLErs7JK4i+RYa8nYpRlc1EYh
t9O7W5E4c+Y2lRMlXdmv5yBXxrYBxkk7gqiFxGoJNEdtse61W5INj9a2BQOCkK4/vAhP0HtX2r0W
MPpbsf06RBhJcZiTo5VrovFvveNKpOEBms9tYbsGnhztSeRJi9ZhOKM5WHIUgfllNninTSx++8Yf
DE9DSBpZbtWxlt3wFlaMob+B/q/uSjMa2NeAk4ieYUymyqoDJN5YnuuhIF+/r8lTswKONtLR0P3D
OmUBEqN6H8Uzx9TGvIt90+crQQ9hGTKqXibHbKsnJUcShkTQcecnNxactvh85Dm83Ua67kGeEQSp
q25Rt/9Wjlj+f53sjdukkj2qwy4lA2E6iw3z8E1bIuMJNni/mbFoCtas3dnD45jlqXLeKBrq5apA
/ofQeD646MAV+G1qyOqyLI+J/ZLArllR84ObCChyOWOT81UoJGwu90G9RTbY9CzrRGVQThiIDr5j
JFOD/SPP1fDgDRMQCjhk3wiOug6v3cBQKNyhkROerRJbsonZDXkv5RZ+2VyrbzWgay5CvfBGnugI
6wu8+Qi3n/hZ8eUBkMajdMfcPDT98Z6sERbMbP8TVeLgnUaQYJzuSN324hsZZcin0sgh/m2rDMpT
+HNBwW3hk/hgWyySyJ7kfngzn9y1W/PqAJ/wVt7fF3jV396y7D1vQ61wstn298FkBwAHD+83a/+t
YKkif3QNYr4dNGKvQRGX22h4i2I/N38EWVVmjCt8pM3XagglezaxghIeJGTWFgy1iI5vvPcdGNby
Nw81zhC41YLiKhgQ3Yi05KgG5XcVby0Sl/ebi5eLJS/eRKEQSOvNvZpflRKoKgjCXNnf6dCo/wbk
nBKAfMnuND3qXnmXOEB8K6t85kR+p1U2KH67SkuOhiAPG58GTaDndjk+dc3DVpBLMwQ8X6zT5ZCU
bj/IhMB32FKBnU7xduU9XocecXRAhOPS1yDR5hO8lJnpEa++yRjghNWFlvyP8NsJw6ptCJmmcBo5
YDi11iRA5WMGLb0hzGGjR6tOYn40EmFWa0GeBIxC6YZG69ArIyxvv6JRPN1FoJTKs99k0PQ/ohBP
kCsxVt69kCXhYhGmhLGs1PTMrUpE96J6dMJdtLrJdXYYMmedCaqETlb6JXVqWvRzQ4YYfPcv8yMr
awgvzkCBDM6xdizuhMu/dzl3E64J50BkBIfbNHTA0jrgF9UHJUTBS3sGxTUzCWfLEiz7TlWQAfkk
YVKyG/dH8ijm8y7nn8kRDJuZSezN6H1SqFE8SlO0u5knDB32tWvrrbmOJZ+jcWvKKGz6sJaOFqwG
2PfAGkxkIZDQTjAYGx9/XxsC2lCyiFc5KOxlnCn/KChkVrfrMch2wrzNIcChVznV5O4x+ONXdOuB
iQaz3bDkDQsereTmY11ru+7VlCkvOm4Zdxf5eq9jfPod9yV6I9Xw0TwOX6n91KCrfA7VAJHAwiU3
szMfFEj3QUp1n7Kw9sKd3N05qB0omvZ1lM2O0UBsylFs2fHkCXbAFu0GQXEL7plVywL/BaA/GvNO
gfYNeGUjVMnve7RjsEwCAAXFn6fxrAPSViRhVTYpoyjPpIWn+fG0msubSiqC4EdxCqYrbiwaS7CT
Qpi0saGlbOeiZvUV9sDKqwK3tk+FcGUdE93CkCcW6eK8fF6SkFMHhVUMZ8wDxwmqd9ynmK9YhI3o
j3uKEdmW+evWCwRgw4EYCzPVDKiLfNrBr8OfhCAn64tnOO31CNfIGiH1GS/URq6EGQKG4As5fxqc
vpkBcojSvqhwnM30loQPRfuwVcmvKuqV3nk+VJcXVWXpqvT2hrv0SAqBHNEKDGCK+XK+fV63AfWn
weSKkQ64/gis5i0wrukqA4yVA43czrs13fkvfyb1+gEPX51gEHSsr4knXNlCyzIMWz0DhZeGIACS
U9M9pfVXzewxHCyeJhLgKJuSaHuV38WNpsQE2FUiyKOJeOhYcU93VHVWL6MLa2N6XSv4p3coBb6U
sTRk40YY8QWc6SMg6H7LNB0dpHjnguz+3oaHmb9eY41Zg+sWw/xwWJAr+0v9v5xEOAfwlbeG9Atr
FIw1+W5VB83yDLYTwL1RcHfArz1UYJY1LAB5lTsCtjjkSwzDbJUHL7C18uQFHzihnmNYicMVSfnR
DKR4uX+kuXUEC5Hiq6j7yD8W7ZPKzC5ELWI1fZzNExSYSL2uRmvOzOhAkpJZxQE3NhTqMsYqdKDQ
bjsGn16OxDGJD7fqnfzl0piEvxy1qDlv0LmoTt0YjXFBbJ5iY95XVv/dGKqLmYW5SIVpPVHqo0qG
h53zYvQS3lwh4X/xFXt5HHmsEdM8btxUOwmPcvx6Sa6wclDdmg8eO3+XfmxgvLHHXtLAA9w9nnuo
L/j6rjtp+bb8VfGMal3NbveFBJwCqDMfZX+8SUaEc+88eWKEvL0mF3JQQJp0cBxfqoeD6/0lCt1P
SxkvddUGbzf71RB52hyB2lAqAK1R0hcDYp+N4E2l+9OpSdXiAMrmHhenLi1pKWfrUphNDPCdnyI7
5N0lILESAYN8p+kfHD0Aw6dxs8HiapmA0/ffceXu0T+ncyCmgIcjje3W+q6bie7j57YtSQvc7Hn/
oq2+WIsh+zxREAa1tJzurju30QWLdO3XGm6BoHEaTjznr0vUnD5ABtj+PSt7Q+etzUQNV911jXle
SmyBpbhaC1T5VDwr44l8orS9uM234rTFtQCXguP8d9eTnVMuPWgRu2NMN+uZKWUQlsAUo8mKaI6q
Q24qD/H01iwBWfIovzOWM8Rg/WEHCLf6u+UKJLpjAxLNpYJKi6XrvLP4bMdBHpDOpDNf+HaFo7YN
PR2To3bQevBPbCl+EIXC+LgsfOpTIU5a/3MT8IUc3pUh/irw31y77y+YbZagzu7pJFGvNGWKndUO
s/WdLmn2ThzM/QkGSqE9nHpCAfuWzPRPCAHzyqHTyesp2jeW0FJtv/ACSRtWenCwEQruBMUZZ8Yv
Kt9J+pTSXcsj6yJkzvxuGa31SIbzYG5XZAH6EGSzsEDpaQYoXaWdPWwnif7SrBM0pCorlHbnFQv/
VqcLiuCia2RWPLu3bwabgyFQeuBgJMhYYqFSnW58pXq9SDR+JxEQw43L+HuIIdRSoN+MDOpyvdbw
z9O8LTWhff2j/57i23FiO9/acjj9fExeFPgZbaLjrdyv3ZiCjgn9iAQ0Txy7Jh29torX1pm5oAOj
P0764BcyPNkLhwxt8bziH2zU0RT/YHA8FrC6U2p5VoYU1d+2Nw2Ji33BH+3Q0f19dOXLEy0sQq6B
xjt7101thWVpRCCwoUzkrCcCOzknRvMxFnw9yT/iepzTe4WeA9+9UovhxiuCh6TFmvg5fBopLayU
Cv3iBup2GwyIAexi2rtFVNb6zKDK/C145zPaZcQcRAG8ckYUobZPu6/+sepNwgYZBU2GzfffSZsl
w7upXr/6zn060Vyo1wtuB2aIYJqenb8oODXH+nMIKekmu3LW54cDUEZNBPDZTTlU1W39inpc5Y7H
Lp8wo2LYjQUopRK13QB+4E3NksergrJHvSWh+k7Wrb6rIExHD5hhJOWZFR+MldzRhcy16xD9S3EW
CEVANzPOCFuRRXrfOyxWuKTuzlKu+RA8Af9KfucwTWMPUE69a49H8wmVDiY0QIWPJmczdiPp9cWm
djkRMkXNc6Zyfkqs4TCgGmpqKh8/A1NTXBLLWSs7OiHgvKDmp80RZioRoVe9nfuBgH1vSyKjfRYD
03a/kypys6KorL2I4VxOoQpfVC9M3MK4vJyyPIGonCTbljJhg3IDb5Y/NwOOLJIhFFBCrCmG9NJW
/oQyWladkeHzRMYUTNym6hZZHxjV1QhoBaf3OHRNj4wBGYKpC1LvVfLPTDf/Y8DMlaTEn4QPjAvy
OeBtBhg8dUGl4WWy7URG8+v/PcHoxUHWPTpIrtVI+TtzpmdQR7ocu9+IVRykNA1fYNm8gjHjYoT+
UMH+cW0eFWiY2UkVQpuOgaHAk5NLzkzD3Um4oqKAE6y+vQ8VUPud4+yC+Im5q+ttfuVGnYJN5ktG
45Q6FAPd2PUaCXtZpHOjbCqPQTFeADiKFt6H4UoHeTKNgt5zKwLyEKwOMz2UjkogiCelKmRImpVr
Ak51cjQrY49qJAfQQP6RKEOKTtTUc3boYgsRHa97IniGWJ2H+8KqWUWhxitWa6MPRl2jGARBwPLT
NsKKlgiUqEghwadLH6aYFHH/c6ZfWiMfYQ3px+Ltc2NAfPKpZ0pWF9MVfDDvv020ueYRhyLcaglg
+eu9oLZa/RtPWdsiOP9sVLKf8Dhe5hEwQoSyBMt0Q3cB475M6OKAl6CQ7DESMKkL4c4R9OBePvpi
opMATOAmVHU1QFfWUQtFJx4rV+8SiVvXQr1oZzIghuFpiX8Fhdj4v8cNGJo+l7xBDVWrCrta0zVO
/Py+iGGUX3Roc14S6hvKixZCpcJfba0elgAb32+rt4iNf9MXQOxOWoBGJH4I0ua50pLwgl98YxuD
hE4OahPA9qC+Ysk+iiKOhnzLF7TDheLgSI94+27sjQFr8SEIyT0moQ0aL/dJoE1a3DNr6Me1k4Qm
Xa510e9OGRtytGbKtz2j9eRfDkW3rxAbd9aVDOl7KVYKsz2g1nsp2XfHiKC+AfhXYjRfyxjAGdOA
AfislYVHwwxl4PLh91NYnwS8h/Uop4hfSBWsIHgLf3npfhqdzf5ZdFbsVV11k9yeiumO7OPWlSOo
9sS1EkAdqymVjcI2K5f5UhQjuBbt+yQajsKUsMUNA2JprfYU/bvGNZ291OxArGX8NdCDo2SdtGdN
c1l2xmpdzqq//gMqXwtqGsGhXIQFggb3rNJdampDkv0gz17HAf7+tmb0m3jVJ3vA49rSD6rZIcsd
IH9l+4CHpvhHjS7cU4LJLgAncxjGTUmoqNwS+JJc+LvJ9UtpLvXg2+AATs2MSvqtoYQkmqhc/ebg
Vimqgq6yQpHbsOTkPiAmzDDwmLK+4ZQixlr9zfDSbDrT+vAYR3IDMZCMm+tM1iFSrWq1n56xy8LD
BXyV5LUQYuROcNwM/X91bw84zhE4t436/cWPHnZioLwH/K1wDu5YDlGQ4Di3ZqoPi/eT1B+CR67A
LSpuivo34ZVe0gBiag2TI3fWn1G1a+mDj95qWWnX8Djo7L8HjJJ9kyDJxjRMUNl07MqMVA1fSeH0
/fBKztUubV1C2xrHV/l/OnW0ja+id6+Elh0axeog97v1XDsbnEq1srqrdWwAsTtwiYlJS2ZxuKTJ
sijKFFF+7Matq8fpgCMWU8CH3/o1KzWi3646lBw0UTvjU1LDEmdE+1I2uQ8Z2zYhJMwO2+ZVWBkd
fl93Jiwa8zr+9ABqJZ4IM80OVMppJeIBNJ65qurxNrvdvLyeXT8WZEqSOwUcbGJfDV3ZkuIKtuLB
0TNqF73WhHwAzYBYsMg4G0TXueNGoLqgskOxc8rdPAgp2WJtEkzS1NfWY+KDnR2QSk0Y58hneBN7
8OZG+p7DhNrlAdopMusyxAzNYol+P1z3J/hjAyapdb8GYXjBhdKSNLV9uSqpKYFb+y5p7FEEJqcL
Wqjve2Mb44jOmkb2jjdW71Olkwv7CeT66n8UhrriiZDgY292Doqkyz9FyLZATNg6IHOxSDW7+Tkm
KPjQHU26N165eUruH6P+8i16BNSqzFWoJeqibl8RBSwBcT0e5ijEIBBxL/WsgV+ISJtu/LbJ66Ci
nQiiSITmJuN+Dlpl8j6iKQDuYZZRA+Eo/qrF14pDbExdXNDuReJ7UfwytxNxx6k5dxskatwJosrm
OfWnIahbTaz7X2f6Vll3WdhF8geWhvlkCgs4jH0tT5o/GTT5bOrPO6WFHhUEzwpcwXtCcj6/Xbnx
UiyRXQJyBWQWq15wnIorWe3XGGU/i/N2yA5YifOWCjCbsiDjEU9Vt2mTOjgDPMsljQCgfdgC4nm0
XIy45KseEKU3SHF1hr0xIr36UD3XsCXK0S9k/t3Vj/h1TeEkR49GKP3P/BLsjGvGdAdf3CKd7no/
zyi+Axk4Vj41wJ0u4hHT5U6wpYOp3x8ING8aNcegF1fG8jbAMGSPFXqprkV4JSJmoPkMB04OcMBu
Z6RkUkEs5PtgcGb5u9X5yQcR1r41rb9jBZQtLZmN1kzpqT4XvoTTbJ/12hB/b04jh9P55V0+Ydxv
cerSyZBBbZAdku6ABCRTJwY8Pxi95I/ScEFFUP2e0jzsRkcYL0iccidkZix4TAx1xcMP/cs2lQj4
zavTl4uvqaL+D+fnK5NRDUxbPnNvJbVLIMNJ8G8EbQUg+Y5G4H8LVCq5arwGRuKK3C9NMhQ6tOpk
Hqs9wP133hEVZRumQZ1BZGOBMysHfSX6L6JUCgap47kDNfzRojAhTlF7JeG6mjECHyXIqVsUqi4b
JAqfJVX0uNyga3kZ2vFjKD1+A6yZK52n03xh+4VYrpzKZ3BedIZ9JVW2Nxab9vL5xGM4Vqtyuo7Q
YsBT8gi+oVh8uqiFuQbSWgwPfkTO0lqH5N2B7l55FAYa5Nd5RXfEkN2v7CKIzQOBiQA5tg7WUr/x
vs9sJsuZcqolOZ/qoEcl0xMR/yhwUZ7x/3D0cQJaCbWSyvvYjZGsAsrsGmvF+6Hn0mI3n0vzKekS
a7QoxbiRWP+jBvNTNsgp7MB8Dkj7V23VCDPTjjQd4b5y5q16MZ8pahs6jHHkpXB4/JN5Mmb5d31s
9ht+HgVPKHu8c1V6RQrK7HHiOKtuKAgfvgkKsPuDJg4ePb43qg419gi5S9YNFJDlccc3ccPtwi8L
oVr9FQaJ+7TY3hAB5xThG4s1uebiGVSgbjYnrZkwus+wQRw32H543lPsp5xhMUfu3k6YVTst9CB9
vcVV3jz366Gh6xwXapB5sAs64Shtp8byLTsz6Du0hy7Pup3aaWnY71PaEg5/eOWthTJ+0OQDgoIh
UOgoIyGFnqcBmbScd8JgOnpbK7t/naSb3ZDxJ7MVYoZn3u+ush6py9RHUegxcWmixDD9y0SRFQWy
AZNDetyu89/IWgsu9GU/NbhLb0uI3rq3mzb9WUj13pyFWGAhKqJZ3La+Up0qTFCO6Vim6V3JkVbS
cU1bwwSep0F/3gd0GnErlllEngY9JP478yj0bZy1cnzXXtar9AXhLcbHTHweRaATw0O8iEOAi6QG
mEdvHozMuB37IrxLuhZOYNrbrNcBXAidZpUN7tzSxEkgxH9S32vpJ0uzHQPMRvOSuHBPpue/nX6p
/IOGdwmJTkldYgCaIarPsrPC754xfzzkxITMKVb0/foEKlWgLEs79d3DVl+ip3dphJ6JCExUVAxR
cOSgGAOnmDPMdGAUR9mrW2/AnMBJasYCC1Z5yBpneLg9RqB5ZoQMz3fHvbTz5jjflkne0lX4K1LF
QyOTmpDMHKbeajzyZamI+M7ZvN5aN2N1/WcLqQpPSkThq3RlyVzeinHqWc1uUwv/Gd2P6mpybXTh
qnsfdPdCpmKKDrmceTFaci5QXGeog0OsyrMeghCrIWZXNP3orXMYNDmdHgr27y0I6BYiB/Lw6Wtb
tSFQKuLnaZS7Ej3k9f5fuIi89n7EKQIx1rYmf2on9KuKnhD5mYdqCrTXNiU45XgL039ZEWJRzKIH
sHtwJ+QsjNinQ/vSr0JiVLGfWPuOlSCPd5dwOf7I3AOxC4Qq/4CLaiUuGdUJdU2ZTu5ZsVxuzGbn
99Og5ZR931tUwtBM57TgzRgK9qeS3nLII+yhfjVXTLEXHA6XJKetOt8I3iRW+5Xaz8StoaaZT1W2
1hbk41XjItV1Lk8qUz7uF81E5uEZfCktdiz69r8CM1/73FeOTkO9rK4aj5k4WUnGPSFGTc81RfFM
NfZDsI2+HYK0RQHL8IcDaVhGL14lW+Q/VKinXQgPo8mUwO/FTte0TvYTTB+VHPy+cNzUpII6BZkB
VKekzqZQM+nVgHF91dD5VK+9NHK9N8jlRIWbuUMldhVMrvLzjSX7R74wow4kWMrTmgHBWrCJjTGT
HTG44Ab7Zx9s7vkgf6CX4GbDgLRCnZcT73eAd5feIhNQOCb3h0HxlCuCHknCcDeTV6K0dDLDRxdk
rNAhDt1fBhe9wblFiznX2nQuzhtA/nlHMAUo9puedkxFcNyCxe5bziIqTsQcx/EBQSm7DIhLxoQA
tUPVoMVbLQZ3IJvHmpa0IFq8lwAdr29jFbrX7BwIqXNlqkTu9Sr/PZTMJ3ykd3VexAzsOMsT6drv
4quRmxDTAJBIbIPcGQOnPPL0ogCSxVcYP0QQ56ZvneD4FkQT1seClEVndjbR3GVpqpFXtCGr3Qa3
EcXr5v5J1I8a1AOna0HQcOKAWKJkGGykTMncjpCD268whBXC15iLnxkmrLyiAcCl5w4G0rhnt2F/
0ME0wzQmwieLrVV/N63ZPch20ukCzvhNOOwVPswC4rAKuPRXiAoeRvePNOf5OFV+w47xk1Lv4S7O
hhFA/lCSQZJh7PJqGT2r6OO8CzqivRFGEaalNTlygIJFq2JUmRvajE7H9gy+HZD52nDVtkEryXIA
+xXgxjwP4gt3Kl13753qXPpK2F2Eeq6+oq1gEyEzCZMktt6bVwp2tYHoJU9Pvq/8d2cm7sUHVsAX
SFaGye94fOJn1HhfpLCU5zOPn9z1Cn9LlYpdejEtBEmTeRqGqOsIzKE4YM/7ABqFtHNhVyWNLRq9
ZiYBVAQmgUlPsHvxkKqPMqmRHlkJpuggqgC1E6SRN2h4aecfFr0NhpRWPVg2xolZuOPpVG+dgPHj
3ehyFm8e3mMvXPxR0sv4PaOZ2MyglLcR+Olx3DnmZOHia5ntUmRnmTom1KiaCuHguaGDX44Wo/Tt
Ubv27Vn8KIUMJ2TBXIdkGbqkPM/zFmYEVDHYAFaraRmKFewhLEKZUyoLBwVAeYtqTvcg7eH67WyA
HAPhaxs1fp5qNrKPGP7hwf0d1skSFy4+7y4KG1lR+755iweMJ4FPp1RW9lxbqiQpeE/TrWA1jCsA
3SvRiNq5P2CQCtKpZp61sGDP8rwf3anFV2OmTZ6kyF9wvfv60ymsvJPTX8DoJiLsSUMs2je+aSkc
CwbcFRjUDVAxtPTHubb9S0wef2Q9VSk+mv4zoJI4lvG9ACYZZ8FdC1VPkNsoQjYvscUEyyXn7rj2
rPUa4JsM+lleCFdQUaluVg4JDl4VGuuvbDfebxvXodCCD22UfgCOzAceIYN96vcXU0RwKX3UnlOf
PXovWEUhcnrXVALVYhLcGBrwmMtPRvZuzFe+NkADIpfkF9oGy3/AR1RZsU9Nfn/DQiHR76cXNEqN
c0YhQozbT+bqTG2pz7I6METD4G7O9N74VjAc/VgIgWv1aSZv2d/HELAPdE7ZydUT/u1a+J2UNNVH
UB7U+FzAgdQgzmBpiOAUksdD/hl84zBdjJvzto4Pz9xJgrvzGw/zlrUoIhQRpcCE2KyWs4bsn/wJ
HHXNapyUd5z8LYMCaNMk1nbJmUPmtUEugiI3zu7kZTQmAqS5YO+UGEaJZ/x1URCWRTslHfIEwwqE
oGQEc2WMqBmQFrLs0Qw2ov5Oj6Op3ZmLaMp5vDO9qD62mcEK2v+evnEqnLznbx1Nt/QNl3OXMBjg
3q6O9oBxmrD85WtaW6v6U8b4ln1F+ZlpMEjKpd9WL3U6pZUvNZdScyoz5h9wXz1yJP9SqtHUBq2N
2NHDPDjRkZsb6r1hpM14H6KSoU43JJWp5ycI1eZtZEbyK6X7LQ2Me+mlb9PQOxKR65E6+sb2s0D+
e9lAqayccNLWdBR8NNdJSWhUGEeJl2eWsskvN5g9j+Xhq34vzfEP3IQ8ga6Ps13wdcwtPwRuOxp6
YLVidGPfvJ1w/937Q9T3HQQ7PnIdiHrE2DBOzqNCeoMTltd4DJiDgM0mcOkRYzHdSP6M62DtOIaf
ylytcQk8OVB9JSmJp8fRKZJe7h8fLmmsXLMzf1Q1bo6ssGJGzYwpmAGgY6TbAV2YBMtKOFxZfH2j
mQxYU/FeCQ7vC75qHEM7SHftxONqoneaOWlYxkYJqtSH5chEz5GCSv7mCZmcrVgnNQqeGbj9ktS/
PRFOCDs5/f8miqo2v9BwSed9Ybq5lQZVIE5K9XGoWLeXEz3aoxoh/7007YibQGk+CUlgRNk1KKnN
ZQ9FObk9s1/zHnsvxxZiDrYy9z9BHy2NPlcJ6u4YAoXjMnJ8a1t1h2RQRZIOMUFF4YedfcTG550g
mvXnErLIXc4J3mqDYMBEF89Ovs8bM203zLy++n5F4Uy5KgDC/FQlw3kZ5sxaPcpthlDRYgZlEbKl
cfewgg3Y5cNWiPkdiA/D2x5SK2H5LxkwYZaJYCW2v9ycbvKeqxTRylizEYvyATZ5r2rhl1azvJG4
t7AsM4AfWvOEMT6CavKrs6W1vszETpic2nqvspbmHXJgcydmdAHguC6HiEl85L6MjC/67/QieDRY
5UJ0JqXOvBXO2E/Xjh96rhDy8VWMYUdZ6snuYdkGFwDQwpR/+JR2y4TqvGLzxSg/Wjx/BepxIx7l
3Jf07k75Yo+Zjhz6d//9ueuvymvYCQvpoIANhZHzui29BWTBuHNAu3Gq+zKyb630CRDvwaujDoC+
npnYbgaTsYHuKkFi2IjnJn2Vqf8Ct+HyknOQvfCPwWh0kavZ6lFDiq+z29MbwYL5btKPyeGR1AoV
TV5Ofm/KDcHjIocHKLG6RU0stBEwEW/6R1IEehMHXcerOiXFUSnKRG0G8p3EQ/3OBVBD2gEvMYa/
QG9vdxDpzdAXZAv9IAJRzveeVxxi8t3019TL2th4rrY8/mTjFOytOQJnr0bmMgz8az8/QBJYh1ym
pzFGVSOBsNzxKdSCVlWZuMRO8ygM09kbTh5+q7/3KlmDAIIT+mdKLENkEAUpQ+MZGGLlKn/Lra5i
fNvlpTs0pQ3ZVyr0+sOiHzKPCkqwADksrpwmAE9YUv/ctmU2h6fDjj5navhvbltC2n+b6aQGxCcE
qY493yQpefiJfBzfzKblUj0R/9CqP6aL3/pCJnEyvu67iI8Z1LAF9MyztuFN9iVDtlfWdUOoEI7A
Ekzx7QpeZD6jAJ6aaD9tbBznyQtzs7Jn50/77xAHMlVQ72sPXf87MHRmxJMdE4vATCMrHsURIyj1
q1m+pHaAW0aDnhWnz21CWwHi98lJvKFfMxKTpaTOTREmYVfaGYJG3JOqQ4NBV5MqwmuFvgtxH6/U
ITB1VRi+29Wn9x9WH96AzgaauAiD4A5/07+He2aSsEYcpir9qfrosOdrxuuJQ5QJaPmkXHvKoEhx
eTHSns7YqmGfjajr3Doff0tjcr9lm1qFKIVm0gXXSp365MJ6DUxOWcPDADQiwuKqd5nWOeV6SBJO
qlafZQQixecPtnCLzlM03g4i0N8mx3DkEXX98gBQ8CcwAjD7w0CJFKKKa4YSYrw4r4++WVyp/qTK
a9a8pAMKU0BWbc6amKsmFaH0t0plWhrzESBwb0WFqVUxnbUYs9S84c/lp/7/K7fc6gkUr+at+NGU
r+akOBHia85fCk1SW6codj5WOC6wVTTWEtS0cmdE3RfdpTMqbuhzgC9VN2EaLuVuOqnm7lsTJ4Dn
Lb+9EexVei4Dwag3YWUANECP4XMy5xWzI43ccetI60g6CPkggcuCzKwpji2msRSvVjhSb0F8TrHg
Ce4HVX0IbDX+i3aNl0KtRa7ns1FN3jhfUTta/xYASmK+mkMAH6pUi7D9BPwCWAm9w6f3StN9NhMx
AWN5sAYWfS9cXzxd1iI6XwK3F/VTvpafpqBxzJJoCSxY2RDSEMQqHYFMZWhGaXJr33400h88AxgB
8FWsnhLfAtWSLCpX06v9+CRUaZRXPLGRPy61BgJuPH16pwslwIObGROFCb0GkHKaf9DZMM3dkRXK
M4tD9tU3GqMAlN3IkQCogrB6HhFN3dCMjTuBgyBPLd0dYbUvSAke0K2f8jw9nTlVqFedR0XuTjL4
I7H8bOEKgEwMljLiqt0QtroRrZ0Z/CVhCq1nqGzBKT78ndb0H+TG3YRg/JqoSwdOTzGhxl8s0mTu
4oQ2lmIEoLei+onSizsoTdQhYfCl1ku/VWHqjHNg8X/saSOuz6VrHFETkWDdpa6Ll9oKa8ieP6/p
TPSsBuOTfBc6pAisEXtq0mkBCaH1zPDDSnObdJotXnZnK2YAGsLCiDoDc9spduGtB2xnqq0WDojr
yp/6vwM9XiKdk4caf5DQL2dMLHAGZXaP5Xsp2zAmqAAaYzM3V/MkMNEMXRP7DQKCsRNaNrVAJVIR
pPhN1UUK3gYJ1vqMmOV3akckGIJTaz/lpSw71Nc4o9CTdPa/fPfSbqpxECXh1sB7+pj+Ndm78lYa
nHcfVqmIh/0OrGmW0xewaF1IBwzHY35Kt0fokM9KVsTXKUwmTGZUN4wIjAU6EYlH1dUwszROR3V4
NvIBjcWLC5IsCk8D2noE3EHFeNAD/y4XtD7CoUxPgvSCciZXWxIdkqusq0VeXD3J10xxfdQWsT8m
ksxZNLQClRqfliA0sn0ExOkM9nCpvgIMH3rT/LyZas/RQu6Vx8mltGa54IWIYN27VyisU/J7cs9y
E2db3Z7zYxGXNphW0IqkghSFxELxZsHnHeG+IcGwlDY8m+5JvhSyGCdL+0N9i0uDskY1kTPiDqOJ
zPaL1KMPG41wMkY8cWTNQDWhGfEUvQR+nS+kvDuYdX0Z1EIuqKCk96vnjJKmMwat+EVfeNvJX1CA
dQAWZgadMpk+X4dRaSWRjglCkVjPKq2/UdBz2Ztbi+S5LQxH0Q2rTBMljLtdjeQVpTr4gwp0OOD1
1iHwS+QY8AEfx9NwFVL5oBhxpFuBPbG7U4dxgL/Psu7Uh3E5tYGlkh8pMHS5lsGv9gQEkF6cjkl6
npvA0s0SnG93D8CKuBzuJmY9SD7Pebt7s7QOMng26tW4GavFeGafmLr/ZDGUv79wOPz6FS/jHBd+
IfKMkBB4o9uBnBiCVNgi54N8PnoWejJke9bAyPUmeAsvvjgtv9VWMQgBB8/hZQqTHXDtlNU5CeS/
PmgYx/+edKGAQTABWYv/WtQ6VXsBmwQJb+rGkDzsEPv6E2GloW/cUHW/XVkIAhOhz/HSVP8NsZWH
18dgKvchR/L7vcVCwhQfvOYh/Mqf2lVn4WF3i/k+WgzpzeAxP/tKMgb2RUktj1Yd3X+JcEs15bVM
tA1MaYUZdAVy1wkEcbzyB9AA0+2oDtlLF0EMn7502QQ6fZZoHFwIgKDXD8mMypDS73OD8OuAbZkp
+Hc9M40Nn1aF+m/fCQUAVy9HNT5F3HuoNK1ANpFWjcvmDzokcEPebU4gXMFwGgC3VGcaMB5Ssau1
muCODZovOfExv+ZzYX8/6BbhpvwhVbLlzlxDzlE49UoaIGXtYbRfw99j9GEMqkqqQ0s7RXoPbzPc
DQcJsMkR0Bmgu2OD/vFMYUuuOlv64bgjxjBzgnLPmPbAeyZ4K3wSrbnZrOdfHklYddtVoCLVOH9v
RaBqnEhZaZ6J4bHtpcdi7kzdU2RUYLIs9C1Jtx15CHLN4HPRUD+9cCSjD5GbLy0hRtUpKJt+9yrX
v0bd1JqIA3GrT7ZsXiI5a9nOEcUXqk4vZhqoCr5dzV5JvY1FGjr7y9VhnrNu6in+dCg/CqmUDmzi
2zTokh1zPJqHCUTl5tU9dQ9zSgzSqsEbxHXUy3b7xmpi99OsRvUeAuJuAGDfixo99p6uoRyX/Vyo
Hs5w9Udc69yUTKb76ur8aIRJs8+tCj/ERWfLsLJ1yehWEatNd6QxlWOhGJ9aU+CJBquIq1+LZTAy
YePKnd33xlCJE7M8jzVfOYN9cfyulmhPWKOzwRUnqIn/4z5gusGQucSglFozI8l3LUVeM0CnMPjv
XhIojQkf011Yj+3q7jpWhy9mDE4u5cfvG6sXCDztZyWTLwTbQ5HRENNH+29SLt3HsopY76c9XuRJ
acgO+7oErrjQdtSFqgIGH06hUwm5wsbSYCg5LzKXgoztuHOPRzdyOsuk/gNlj1zLDi83Z2QvC5hi
AoEOSAwa3f/7Rd6V+obdZ4epWox+r9JQ302kGuc7Oa6D6r9OxxSSOMkc0E6tTHZeuR3THWevr8F4
j/iM3ADttXfugOd8NTVU5jb6zf+JSw2+L5Hex33SvTLRoy6RBTas7LVwPc+SvX/96gGKhYYssfXH
kUGFHzmHlkZbFchZE0q/o3hdC6UvXWOouJytuxTjJD2/tZaVcCApg0+mjYLyCzc+xC5xtW7CCO7D
hC2bJeYRrmnuUKW+rHW467rxUgqakVanWfrwOXP4f1WEp45HJF1QOIJWbZantZepo9mo6rKI4U0Z
RMdyaZBqZ+Dnt+W6yxDWco6Cp4vZ3RjaeB7pamax0uOQl44MBd4neJg1olMhnsSVpfM9X/dC7WpW
CheV2DQWKG0ac6IrKxrkJGKV6j+NbQUTC5Tacm7VFvZGi/yrDt2CPdzxPsF4O+DIXATLvPJ1EV4g
Kfw3ghAGp5k2tjcoRBQIxX+dZJeY4r6xUZiQgk+G8oSfNBhmsisKEwN8NoPx7aKgxStWuZRZdU+h
V3/HnNZviAGBKToLC7P/Di1k/VYhJH4C+ZP2YoKCz2yK02MPi1H2aD6WbR4Z/YXLEOApfy55wW91
jhugRA27yVCYyGqJoTF+0hmlVqa9SL4hBhYtMh8q8zxmUKcspJT9rNH+dEM0HnK2+I+WN/lG14De
eJr9RuxQRtdyz7W7/l9A37Y4DjgPQmT8zoSq31uiHxghsVZQlBfnfOJLA8HvjHjSSumK7XJ2rUiR
q2d3O2wLosbw8BfAm4tMxDMnE3lqHKifrBlHYcFKDBKOPeoqgkk206yTYFyMukqEXbpbcOd++Z5K
36FJAQxyQVcX2u/SrJHQ12w5aMpFfAwdQUBZVmWVHQF26JQQX7FyHlx+HW+RstJCcZ7PJ/K5RK5s
gaVC8qUV59MDcYFDZNNrTIZ+L/DQK6rxcWafx3IrzwkYJ8+pURuW/fMmcdOlE/VWIEObMYMWKaqt
we88UD+EmoXNFTE2Hm1D0MgLL7obZd5vC+e7RlSf6JmbujtsezH7KNIwSCSADMhVNNYzVRVLylA8
qZOgdCUBjs30rwpLdcj6mGWJhv5MBbGtf6cVCQsAkkSnX402I+VNL0cjkhbJnPVuA6fkDRloxrnM
WDyaDEWWB25dikm9jlkWftCtj1tUtuAEMWLs0DLvY8i6Vbz+SSuyM31E00BVDkgemBfwTE9HqNPN
vqNkgtlsffhzI3Qi6kxGlllzKGtcC3R/6NujJnR0Vt2FHTULIXYXQ+GlyqBu4gLjtmQnRuV8ljRy
T+hCOJ53VcqkDoVELrfcXB5bO+qSsr4Gbc0p+V7xwJBiE96EfdSP6BJQAVWiiSM6ObDRzebyaw2C
44CplSJlJE8dbVZPhpoggRggcBJW0xRdCke/sf+Vp7DcUkyi0wMbQRT026e9+govlOIzrfpBIGJu
f0+a31SMonkXwRHhUEtf+lSxFiXmViFaK0RMkxH/voau69gDLbGPMgaSXrgzVXVvd5MVMvXiPmNs
JDXOv/2Vo6YRuJ/apyaMrYI7tfxJL9VH1gV8KH8mqUTlqATVcdSIg82waQh/6DNzOkN8VtHGswJL
TIQHjf6kGJg7JdLD/cTKfgApviqyWMYgW8AcNqnw9PInGAPjFH98oXZXt3aTJb/fkTfY0dEzu8Cq
pZ6C5ijXPcgPy1/XiY9AeFhFbz0R1vSf94eS1tYSDi+87NoCH4MuC3n8ki/hzA0il8KxsLgM4Pz0
lohO2sF2l3S/l4yWXtirKuxU/BUudL+3AamGnX0xzemJocjO2ETXedynugRNf2564YUqhvtkxFj6
zw5nz5Ua66WDate5gVw+gsi1ywcaQ0TUzcPFCVnG3JRgMXy4xm7QCpmtoaGDueQMjYsUjNRudsXX
HMaqOCHBw7/MHxgq4B8GvqJ+ozPGvLo28o5fFZMNiLwTbRZU9wg6g2AfeVPLRNIK+cV9iiolr4Ay
vjrfTV/e5UPPMoQ4OosT6I+WVTA10M0AAsQBI1HJDjZEsfIL/c6lLeXer/d+CoigMKbhmNc+2m4w
TVf+Bwr/52HKcq+XTelSY5IB0u1PkPOAGpn+7W9N7ZAvo3/8FzhSpUARctyQQkNQCh6jYm4i1Yo1
TIcOeWh4LMR1mn1LZoSKyK1b3+jZBWI6heptiLqYyrwkUURG3PBeq9GEFwix+UhoTJ1D488rr0Mq
Y+H6agbMaos+Q25An5FztZrotQFpeCKxON65Xt4TPCqtu1ZeBWFmZ9ktix6T+K63KqLoA69Wefq3
v3XN5QvTwqqgmuN+buumFEoDjuA8x82e40+qQCsSazY/i0ZgaU5QZ7L37rNzJm8s9oXTHrY66i4L
rfyHLx592nApiKBdYxGiqq+0vQPkHVxcqY3zJ72Tgs6aSyMDXPUpScSSowvKe2XvO/Y9SAzo0Tsm
cGfiO3X9dDsB8yZz4qbZonFy8yt986XlQIX5BKNj3v7w8rXM+DwTAX5TA54yK6ZXgYqn3FLw53yA
4zXnfGAB3zLR5z26Ocsgn2OSU/giErMMc1NN5RIV/rA4fuPFHWohgpwp0qNBTUqwnlCBYqhkO25x
aJmVW0EDuMYl+vFZjiEAFc9bChMtKHPKxSExczeJhd9YtGk1/euB0jMuSm+sgZ6Ds0sLaEgCTd5b
kh4UbsR2jM67CtjQPk34QGdrEQIYK+C5REZs/1MZazJBopNGOteFLXenQDb4x51YAYP0Iw9g/nG4
Vhwd7lBCzM/A1QwbDxwSZpvfo7MagPs0zZ7zEFT8X+l+8+lfAuqMAYIMrkw3ST1cfQCQQrTQL630
aBQaJNRygNi4HN3wAE2l3mpU6zld12FpX/DlHYWxBVtlJjypa9LGdhvDpIapsjWccTIV0bMoxjLb
bFZR/zTists/wER4a9muL+Fmr40kBR9oFK++nyM0PKIWdQZp/1G+A9G9ayf4gf6Z39Kta1Fa6a8Y
tjJ55qAgX7wa2ppH2COSF3hhDL6y72E6gmmYpIw217tTA2tmBcb8oUa0H7w5cbmBRipvnbS23o5B
bbsTn0l5C8S2LJ2j2KfJfFgmB0+mC+MtWpauddnbc3FBE2qVeo2Gjd+fRd2z/aM8xSJ8VvkyFsBV
b4F+AM5W3sk0wEEJ11wdb7PUoxjdmEyw4Igf+/OdQkw+/MEPLgvgwof7jN3FKhnmC5Rx38u6E1I5
kvx03TUkqjd0H7slPL+ziNIuJPB3pFzY07bmntmOWt9sZVjl8FxoNIJaAHjzP2YiuHu2quXyNpF+
Lr0kBqA5MB2nmQBhn4U0cRTJWE9m81h/ya5n1ZYeS/z8JHNgq2vA58sC5Ulov+zh9m+WgRkznZSy
M6JD9P4J8Th0bS3kbAKx9keF6zbzzgbZrLiQ0XmGANJsjqXhgvbelcMsXnKT5Pv7YZyqn4tCpj03
hU9gCwC1UsK44Kiod8hTr7VC9BKexftgBV4FSyIx7YhLHgYgAJaHki8sgMRJduCdnz+Q8t+m1Yyi
KHOH1fCFyGUqgDl6lv/bslbl3qhIvKTaUbGcyT6wuM2z6TtCucYkuhofEEHYZWHRJs3+Crcuz3V1
zJrspkdOqT0uiJE8oc34Wor4HfR2uT5iSz4mEkfyENnFBixUWuIy+TJKCjf7eQ8EK7MLqIViaQFU
/OV/z14fOzG8z+AeLp6bWuMc21uZpw2jcsfZtCFT3HGUlCiypr4fJp6oR4wXH9r2XKWFXQLHx8Yw
/wsnQmkOW3ihVyOoxWmxoHAY69ejZLeqnC1KmxLrnN8uHmlaQ+CVs7os2Dk+MTnpMyDdUT6tAqwm
XsxuDZ2OLvBBZ72Npoxyv2tWtL9IdyZb+Bd8Ai7UjH7IgTy6f5fJ2vknYLE1s2++U9hLF3KfVW6P
NixpjjVqhIOtvu9v8tP0QXgt7PlnHQpUU8pLggvKgeFwS7N/d1wWVk9ouV3Cy2rYie57bwJvE7vl
WsSZBRWqvDSvyVgrVJZwVT8htaNhoO4KETaAhX6ZJuEx729PM4vlsjRzy202jgop1M1UNWagcpkM
x6f5kmRqYPIy8tFlnmOQE+HxpAa8isyBffH+7s/ab0t1dnv6gkRL6EAwAsv4nOKKM0awUeHCjau+
zSdxcaV6+r41sZebkT4jll+2hDOLGsgxQb1uW4sIeN/DWkvuDjT9ZY2KheLkCQI0orTpWR2q+za0
4e39dLeNtdr6EtF+zoEmGxXZInE7q6fa6dgSDF5KzZ5TJt36eWNpxAboJxpEpsawIp2lrKAyb8Kz
VuQqYtZngTr8CjfJ4xpjuoKNFUNrc1zli2Hwk5TFcTADsuULY5X4o8p5l0VK2KYt/t8/U9xzqvfw
BjnrpXO04RdLHhVKO4Nes9l7q8lRgMjKaDViWia3QGC2PClGXJo4d7SIVJ6I4hzvcRLvUKKwRedu
eLA2edYaxD2iFWbp46A2/AR34Zq7TRywO5xs9jS/tvTpu8t3t6v6KPaNKqAu2YA++lRrGdNQFQ2r
UESzTba7eFgCtzPvOWorEKVeFmnGTOIW22sQgonaVJyo042IQ61kkQNN8sO+NFcZ38dd24SlzWGQ
yDTPiDHiulE/zmSETdlKhznU31jFMg6Hml8vPlL5nDYQ+XmB75Xexh1ylkTn3Dk5XU5JZRn8depk
l76+VHWjlWhEjeJnoa4rrYoeNRuO7kqFoavR6TbcaKRwpVWgk0FRC/p9igBi6xD8apKb8YNx1MPP
KaVFpIcGmxQOYcMhRIDbIPtGYsZ+HQOr4vbwD8j0vgoOUy1jOT3tS+uQLtkzG0DMKYDgAJhRN5EA
Td6UKuJV8Kshv9aY4m656MmsHV9Qmb9SHSgz/Z7mJfWULh+v+HhZCZcaDyy5qbt3CZPRDEjPsC3G
LapWcZ0+dgioj7o9WUr0qo9z/fl8d0C0eNOjSN4LEqCoM0XHIkl/CQFG8+6iFjab/JG/eMIu6KUa
ca9AssuNRUQd/vZ4kPSMHTscJXBvKcXhqa18rAYz/18WlX/NEjOd8wyMji003kPtM/AuxL+tL7fV
VBjjg5QVqVtohbKeWCoLoEYSRraFKpK3LnrIzwZv5EaOohoYW6Bkxwhs4EK4VFjmEDh+cmvBv4kg
Zke5wIaTzV05YpHFxqDt7462e5moZrxuh0KmGUbwEZRTsrmroKRJGdtlSBSGoWTw4Efuw5yqGPUk
8/7j1AfSUR8HN8gwhTHO4fRo5aZQjJeS7lZ8rTy98/R3aDZ0m+oAmH5z49+4pFZ8ijLxZ6YFN5ho
9sRQcqG7dS4VdVHX6IaY5fe1Wt6pMAQ14tLl2dvZep8htNqrxDTI6nEWhwPve9Rip28PbGrPoTXT
ozsgf+BF6YvssmCNSVbEVDC9+UvzAle6QqP2qG1iitnL2bFOqEcwxsNVvrGF0h/FX5zRqWa1Ooph
hS/4Y57cNr6YITa1MYCDUKsQhqSFivbhGghYlEX1FxR7F4qt71IQxZxD9x2oaDKoAn4oYWWA94sZ
65f7enAqtfA1hdSkBxi+PD3dTYIrXO1Y+OgjEvbYJmEJwVpsj/QgMkbjdEj3lWJhrGPnjOCbl4Tj
3NaOp9rh3lsjTYMG1oEpkPs8NWcjKBkeHQrWvmeFwUr8h2BQ+iq7uEz2Y7QOUcURvzdPSRCexHcd
k7i3OeUuKyCTVYelkHDbs0EpwtQa9uXYOflJGsLbg2PTft3lwmMIE8jZN56keLJcknWwCwCoOj1n
OvGPOyrM6nf9Ag1UUeRpCbW+dV+PT/XYKJCL2WcKk6ffUdrvf5gBFkcbEVyHHt4xBPT64DEofdl4
o7k/VYuHth2OD5DRQ/WvgqG+G7WS98XxwaLer9U9pc8W2fT+mzSgpzukpxnRHB+xuT1yflZ7Lzob
Z/cepwN4AFvyOWCH8kSp6vvXFGw5gGI7jfrsv1fsJjFgbuVM05KrIgwanOL/ES8WtGLz2/bO4VkX
AEoIIXT1/SlYjSjHjomNtgU4IGMaBF1ZQIOiaF8mgfeiRsDE/uukKBGce2facArugNJCzZ1D0N+q
9ufsVwDTQ+LgfLG+Xexgm73zDfK7DXknoFn3PpXbN5E7ck2li3p8gCVMnh7A/R/dH8bokCMgjK4E
wKxTwUbAMwwBpH5r0ugp0G7DHLW6+UMIBce7JSgDP4fXRm5dArJes1KM9lvpndEqET/8yZppKGhW
Y9S3EDM91eXZ4BGe/ZZOhbQMDRj4ogeQotWjZiwVlwgX8/i6of1n3TANLy6Jbhn8jyqJ7uTgrnFN
TQSKRQvk5S7Hqmj+TFDlPEg2/Q8E78sIabeDExY1Abo4NOtIQNwjmnQxfeQ5PEWc3Twp5KUOgYmQ
PQgYPmMGvc2ztAPXKUhDLUnRQQXVcvfO10D9oEsjvVq4INz52hkXUuz8gavt6UjEkMK8ZFM4DPur
rZC1NE+iR3lcDy4q9f1dg/Je7iBo8wXaLfdgZy5GQ4xno5eUrjHMVkWXtixNyMAmJ+IjUQWaSTqG
EWP/VwSpRVhQrzcKExllhzq0gXZ2uyyWJ8J3ZywYuf0VCLxVWaHzOLl2Z67zAkkUJuDwzr9mD+7O
O3dysOfhD3qq0+nZz/p/9K4kRgyfAZ9X8ecAoM841pxoAiG8Mbw+C8hekOkMosk2Y6VQvX2rN0Zj
iqpcG+SJKKJ3QTHB1TUJFVrphLfz0i2JkCZ90xkXgwyyRjuFSHEzvdbtVdrR5zI05zvFxezd+Fmk
Ra11HrWxAl/ltGmHm/pzqaN9GAf9OB9uN+0ZbmeXc1AEMSc/AVPIkXGnhr+w3RYGxBnKvoLFt8wa
B0j2MkCHb/5pw737EJGTYYuD0VdGa61XB5/IJrKC4boYEEMAet2VK8LlG0w2thVE0braf4PcgXke
8nGnkUeDDRO+gs5TPsyhjGM+nDFtt80yIv7Q/s80HvyImZRemgEjn5iA8gxo0/8vkqohq5KM+0Xg
2LXdmJwHiqSSjyyztgDe+pNR9HRhRvgmHtpUk3u19FDSnJoc+V4Y6j0yHwKVED4KjVpXMhqf+DQt
+zPPpmuuBGICrEod8vHPAd78ga41T3qj6Yv09d+LdLQaQM8UqTbnK+0QQaS4VXRk/N+sgxkrGhMQ
u+5ir8F9BnLruGwjUvitXtK1n8hsFOwT/Kgny/EBlPtqDNBek6tTBofnUpoQZN1UGO0XK/C4AINw
B9mr7bCaDv3OvGGnOMaXoEKhrTVaGOG41SBN+lNLF+MQM3FD133iLp8IjltP2n87mHhzDtmpiv/X
YTuoEcOJRxGS1X5+2UUJitKzsyQVWl6w1+ZRaQBCOQAHFXVRCchFN/AoZ3hpET3/eBr16avj43g8
lof0eRUNjcQHGt48jTzBfEbx5ecW6eLBzdIm0a3mL4vzXqvjoA7D4CwWO/RMKVHuR7Qmm4yCteBQ
0ephqDUnunzPqnpLf5fmxxXIFFwdk6U/MW0LkmjElH3MJhE9Pvs5wDn5uM88NN8w+ozPcZ2s23y7
uJziTe2WUY2BEN+HNY4ThGKYiD1Zu7QQB4xCaw5i4uvW2+pN0tQgVlynKoPHFCxgg0j+/kyoMUCA
JF6KNMeXM7vEadkXq+lbQzPN/i3zqmzQr7AyWlr7fq+miKdDH+pt1+DDgEVMW44igjpMgoLTJLNL
u4IjiBwQqNGHOTmM9N3UCMKmnpsUqr8ac6BFq/Z6n8tRWo1yZ2RRhE/XSIpOPQ1pMdTGr0akhPsU
yzQDELty13QDbK/D0qIfHzJfPrb0UmRY/Ra//Z1JM1U1RbqrY0hBy7YAbBoTSQ3yYBrCz8XiJosk
8wX2cHCo1swsbx6B23b/cWFRk5Z6RkMBFQqXc5OkiPeZOsI+poXHwKr3+2g7GL/pOXFl3MiLbaHD
rVUhdOuDEZtl8WshiwaK+ud8dYS6ornZII8wZVTTZIU9Zn9uWbvrWgB8MQbczwJZa4Gyeid3/omF
WVf76y/8fQCHKnQnBiOpa5eTfXLqvKxAU+bZ39GJVUgAIA2GgkFefw2q1M/J82fIe4/r6wcSqwlP
rcQIuUOQn/UrdGvVXfVmL7HspcCjyX8GRjjLBqUgFPhDDCsJ+oZ+vcr4qq7MYl8ym5bREA9Tf3Z7
UiiiIlhFu+ydl03Ogi1/k42t+JRWJSgM3PHv+RR09NlOtmewd+UVz8VimnZgeilwmVxif2ldy8is
dLPgdbbFFfE5Hi7tEZv5r5hePsCo49+lb1vWGRpxM14aDew/Nzy2nQTeJ7moHJL6f7Cx1iSuV/gE
cyuJYTw9CLXsLJm9YTa6zkWdGsQzY4GfKezDm3J/yy1rJnqT0ZQKb0OwcEDFoBwx81Nhg0zNVcEk
CUySpMmb5NG2rCWCH0x2qi3PgrNzx5kRQIXIVuh1XDEbnwTwpXN80Ei6QEZJpA0OqPio0bh9zXsc
w5QAB4o0CYLLFGkxH1SfzUJWDsH/+hzZVp8fi2yRv/IFTX2GmsYPjqWj+q17VR4SP05s5YNQNFgf
vJcWmXOFrSVHzxHk03ZQdGWjjkwC3A+MNjS939OcFTwWYnSFaVCrJPaSTfSKAtkmdnDeucrhOd6c
sSEuUqxkm4Kh20DWjkNrRFfa6spFo6VpgHEPmNLERsfRnW0coebex8CiGo5hKyGuKGFzz07XwI5I
n09ryXpYECkAeLD61qjOVKFVPz6s3GNYfollJJuyfdOnYsT8FTkLRTlzTZ5TJs/YcDAJswVPMmVZ
QFg35ECY++a5yVCcRvx5s6OMPJcqpD7sMi+OHS+nQLE+K2rdJVKmlRBVwr5qkf5scUenTpHL9yh0
XXZVvuj+6d84pmUaLRT2t95s7Ym6zOEcBBbOrjJ1DMCiXqbmKJlMTXBIAxFvvhIrSVa2kl9jBeca
qWUAGTh/ookbx0xPANuk+S99Q47DQ3RmxFcjfO6Qy5qbH7C21QKW2zLkpc/9TCO8D9rredNy41bM
MhgR/Funfzb57rKMvDbTvK0T3NW/wTXi3FdRIea+5BJPgY5+FV1yYrtsebCwWh1KJm+U9T2aF9fx
MbYDEGuiV25psmzHWsTqnau7JY0LtYkI1HB5Bi2poLx8fx1pA/dj57PUTZvX+ZpDun3T5lerz+pM
VWvo9/uU3tbllNPWi8LcsNW5Sh1DAwRpWViK8189OVs/Tsi2egmks/01JyRexpGP1/mUGIsuICNf
7TeDgRkQssfrOBx2JjaSHaBUsdQ4XyMSIy5SJsDy/q+si35SxVL45ClnD5SWtZkS3wPAzZabWKrW
Z1HJpvXgLy2p2+I3cTWhtUrVTCAiacjmbQ1PbFFUL9SsT2nGfBvfVXjkKMenE8rnR0+jHHsDoRZx
Rnt8VeveNUFuSjnroe2xDMEZR8lMvznRhldLylZRHaDyNOI0tBl3bRvWn6ofSnO/MZWieYFkSYxF
zVcT/AJRk2rhMsVEtTO2ZKPxmbzyJYkIvL+MfwGZqyDqrm/kWaUlSvjIJGZf2vRXeHb+c2hqLM3c
t/eCIAzaFK8FM7t8ALO4NaadjvpoOmvaXo6vm8tqjujNs22c7u9MYhDCU65gLZrEfclg770Id2qO
mzIcKh+LdI+Om+XiDAGejvDy3t0ZQbPoAIda5+zxo1LC8GZl5rA1ssZd0VzCG4Wm2+5fFwfEl8J1
ayqdZSJl2O7B8vhwtf7tBEiRyP4HQ5ITAyRunhAI6tFXE4uFU/OY4AgZoVmQ1+sLpwq98t8+6/Un
TjDTv4h3jflX+sCvySZvk0f8DAnzekS+qpXxRT+uqkPHqzGBh9sY5bNxIYcynJ9s7zbrP5mOGPLv
5XaHaHt8g1Wvb9fiuG4G//Q/vT4ZxZY0CObaiJLCrQ9zuV6vf9MOhtrgd5PyNhHBif/3ZZqvHSsj
nnMVlZhfAihcJWHZFSeFuvcO4B5LKAV1hbUvrXktNdtqXQdbtnzwI+LiX43AiUGkblvpCa8ec7d3
7UUhZKK9+1KVUiRFIXu2MQcvBldku0/yas0RQ6LE59kd/wVosF58AJpUWumq9HcXIhFR91XYGZwv
27iZYYCPJFdF3I4KBjr7QTjTefRTBbStRwqNKHHoma04Ssx03neVMz0ZODs9BRX6j92fsW9nXpC3
P85Z0FG1ncCAsmIhH9DubsJC2GkXwdRPe0jIqQIA/+zuA3LO7meyRXqrTTn+Xe6PZN7eLyLe6r9g
6ron92gxME5EacuD5s3UDetzGwPhbGzusW46P+sqpLzmk/BRUrDbdPW1DA69sBmUFyAo8koJWyKK
QiGEtYfrjkObnJoieaIaN3G2eQkamTtLi/B0Rz43p8+cRh1iljyCOQ46+6AXTXT8FDvQwYwOMgxv
yf85CMHxk7pYVGh9KPvRJzdNK88p7ZC1zYDQ+t0HDYaSo3flP+JiWkIWsgiAgo2B9LuCBgihTh8n
pD+Yx6j6lzJJEBmW4S37sb+TGBv9iVituZXoj6T7rUvBs/5qM1QkI8/nOyD58Ckm77GzyS4XHcmH
NRQu27sZkdZ9e/RbpCVNj1TD+cWMlA/Yf58x82tUjmbEdz3HCiN2x4BpJK86GBZfjBDa3MdT+ddj
PVC6SrP588m1BUorpP9VhKiQd/LLq0yW1cKS2PKvzwKqqI77tKyxEceMh/1O6ApMEPl7qS11I16N
4MoBD6FIQ48G+LOWRx2orsfShb51+WftGTWSLCKek9jiUW63wqoNZmiv6SSklmIiFaLEtwa62m/I
L35wf0HaI4rNoMhqgltaMGe/1g/p0MeIFr/fk6p8Ld1ypf2mNV+qqAw2qhgzbYwTkL1Gxmdfdatz
GMl83t6n4BkzWV7QJ41cJ2Pmc+JHBiYpHGobebRuPc5rpMmhI+BiEWhjrcP9MmJxqWJzEYUPYY95
CX6LtobLLwn8hu1RW8W3JiuqE3IJ6Y05/fICk8l/ZqerJSH6oMf6590+iFr1gagPjbQ85UbRb15W
GUBY4VzCWvXqSGaWpBdivJeVu4i9qp/k+vDVK6F5PGnsM+8g4uA3gIOrA+uaTUbbmXEgVYhU5hT3
9yxt5U0M/DGV4dLR9XenOgR/b/tn5+tk7fgyX6l2fdmE1sD0+03uKl9QnH7uB7W+Qkuk11/JZb2T
c+M3K/ctrLiYmtJHix8FENC9NM+KhKheaYGlBtEzzq5z65hVpD7MpEQho+hyESJkq8b5RkWEUrdo
iylamCmgqNBtWdp/fwm2GqkXRJjg2c6cgUGbkeY0MuzN4+Zx9uPuX0Zs7ZOGI62+e6PwKE3vF0p8
fJqoJFizU/g9cwdDzxdb3mAqbutWOtM58wa/tusXxNoPo9qSCrVerQ+JHQR7oG2UXR5ue/D2Dnyu
CdxIIt20XPtX9N9pGwW4OQExd2JDAhcj0CPEdAYxAfTv29yuCGSfA0jMXJFLF+Una3O9LkuEhtaB
UY12wWT1qRQh0Og8PoO8oIMxDXjDMJZBPqQTfTfq3YtP4vd/flCu8hOpJjX6V6rs5hcl9kZ/z9Fu
zJrFIDEKoH/Ju5Gx87P5QiiK33Pm70dPIDyI3q4iEaEPBlRWZU6h0uKMSWHXafP3jSg+sFS6sKB+
nFbmpgMX9ikAJigNaEgvREMZm4ihjkvQfZHKaZSIwAWKiRE5x4HZl+jI5AjDhfsjXhhm7tBXqkyl
DMrGWVGFoSAAnAguRJFTO/2S0XTkmDMX+ViKsT3y5sFUqCK8vrqNzj3F1oeKGCyBFhA74EbYDvXS
A+UBVIiw7JqdCZH+CEaz1W/nkZj1+uU3AWNzh75nqwxEsaT4AldC5esUrGtLnJMM81HMLi36m85V
H8sRyl/VNr+gCCEuEsv73bxEALkaag20NQOZjWBTzGEoSnn19291srJZnUCEY9fAyLQT+AHmKsNp
V7vbgv/VRmKHfPxQdxYhzQ5BUtgL0z/+qaqznKa3F9wI9jaFpWJJatQBapqDOwCjun+sII3MTsXC
WL7yY1GOMuLmCx/ewkHlr0X3XSI7OUNnioOGVf7upuUdscdyj5E/KbV4kbyYsjegopmlZ0jScjuq
cYLmr+p9hBqu99QgsyK40lFoUaaclcK0MQBEjdqZeMrm170/OvTAZFYaw9coJG4bNU1W5W7+CFDE
bdpLB015qizUmie6+g/37m0KTdT16H4zTkNbo0Y/8JUqGZpPlKWbfn0YH5g7M/WZCn1+P3kZ+sX4
+VL+6zIoxk5xA7PFDTMasIcXWJ20Bx9KiwJn9OtTIDvWqC5dsnG4wyN4OQKhaoxV22u5m6nunttw
MYJWF69rVNIEQ8mJm8spQc1cUg/NCvp+N+fZiM18cK2Shv6tcAgfZ2OPdcqXBqMOTWIiGTUJTiJF
f34vH3CJXQha3E1tHV+7c220Frx3LZIFX+0qZt6zeiHReuhPXAhXp5rzqpOSo03tzRrTOA9R5q8h
HzzbLkeNgmexQ8Nj9B95uQOKk+yhQzqTfc7ZCuDou1V1oNTEggt7marqe6DXY0uzCyLwPOJw5vA5
6fodj0tSTOuUGbL24YAdNPoW13q0IT8yqrcjmhqXFPLWEynWJqAzjWZnBjeeIvxlJR+9noK+KdN+
raC43aJUh8K3VpnXqwMuvgHjJttyb8svU7XVclefBUMuC71Tdp4wN7QFu41g14HQXedHobO2jp6J
euWZePaO9/R2F8R5dRqHUFx4GyI2MlbgnI1wNfSeYQe+402L38I1qWcXzefBC2mCsRDsrHEsenoE
MbbTJ0Ejzjvnjsw5xonttR+3OIHrBotw/4TwT8ELTf5KrIf5ocRRSaK2Ho4gaovtPeln47HJ+VBm
SQJjHuj3GsKojT2t84rysmnSdXcI76173PNhC5or+Dog3MiPKlJN50o4F1v3k3IX4Ev5/00gPfif
P+kpGoU8tLhrmnsFX/muDgRc4oYKXhcfnmNv8e/ec8MjhXK6jNJnXW9v8/32pI3J7rin4GGdLw69
HpU+tFninBxka63z/l1B4LJ6X/BGi2mQduCJ+4k+j+qJ6+lZn0X/ubSix8C4MJWQWzNYoTz8XHVd
pX4r5xNK+SSsIzfKbb3DpsAGMgcdz+NaV6MOoXHTmpKvwv/cpxND7uOywRE/XRbaxoonRMkZrcfU
6aDMqylxGCcm2GTW3O6EKNdxCuFtJSgpd3zsQ5fGpWGglGwPwCuAE6IZwCZCGICQTSQG9kAivD7X
2QEx/CzWARIQDh6PXLBrEYUU3Vel4EqtjTxHd5/nBtBkc3sDjclnKbQlPY5NHoH++llXdsi+5uWh
ENyjifyc7L0f2Qq/Lj2L9AJoQWe4n+dcaDgvkPC9R+PsgoitGhk5EIszyQIfWBIvyoVEYDaPG7HC
wNECBUteguVa7rO5j4fxLI1umTZzZUbcOx9vGlC8UeA0g3a2PMhVGwlqF0nK4aQ7pDJQff5LOF+S
OYD8ew74MlqVWtn+fdRII0WQVnd88MZQSMkqSBtrzP47sxvmW5Ys9qbZs9b79J7b4AQ9DzeF6up0
e016Met+tH9RZdOniUyl1QjXbnpypoFQE++PyDl2v3dQ/8Ul6VzSjCb0d6w1MJrW/1KEtw1LcWEh
TepAw+e/XVuD981AgbkWpMtGa1EmaQPx0d6Zca2F7OcpA+3KBHeJwMRCW5JrtP6QY26FIZhK2W64
e5zdUFDutL+QkBdRLmSSwkZKESoyTRQ0RkhcJBUbAWVIfxzK5SiDon7BK4AjrWTZ3vtq5NUC/c66
kAIFHHbmGaOIomrmSOvh8DeIxxFVyEaT4EwuGd63npzhsarjhEF7fAIMh5C9aIso7F+ey8xr5pw8
BU7fsvcIWCCiCQ4v4kXOtwMdeRH8Xv/XFGrdK+DWAfNFaudLyhO/VCTFwXxVsxYlEhxm6MlreJjO
GpAIut5bat0yj0+9VzdNL1jLluaR4tkSmHB35YsEL66/bqADetp6S4nCjfBL9/4uKHq96RAiTQdy
Kbpb70dLKRTmlIY7tUQGY67SyPOy5NBRh5MsB3fiV7OPCNJ2coMIB+foqtSjh3cPJfqycuGEm/wM
o3tEKWIkx6t+c+ySExtikQ8f9SF8oJjDw7lDzZApW1xVWcB5YrlR/HWhoeo1QP5AM3qvRbdwq355
yN1fez68CWoG2zs9fpOszYIGwnficU6wD87CPOyBpw+5H4pU/EVAqCz1mtc7SpsJOIqjqAgbJDH9
K1ouGOhECE4FZ1eogupUEJpVGEXqGKk/2T0vtbst7pH3P9fSTmT2A0UnRhQV8Zd8Oxt1piRua4V3
7gByLZJx+f+4+pYmVEQww16pSZRtaX4DpzoodNaP2cBebrkcaFErcZOiy8f40yGV9pj7DwBbkyh9
xleiF7wQgMVW+PDIJDYVEuRQfIIW/9UoISIVO+FmYjno+TjKa618TMI5c4w6/kofkMWFDhfHrW7N
PjXQ5RItSYgx+Uu3RCnvVVhFxNobA9fxlRqqWggbz+VFpC2JiL4D4Zbxclzzw3bdfKKTgNnHZona
3pyGjiGywOdeIkyI7Swvq/dYBavzcY/QNRLB/1GuRJAmEodw6T57PRQjPCNpgnNWYeDMKOGuyr6E
Q6L/5u9RRNoho5dvae1pVJ6QateqHcoiwGuC7sBjz6wA2M4INIZdX9GG3hy6mpPxBNcQWna4OSKb
F4ybVXoImzLJ6wDP/ZajbXR3jAvKXC55GoAZ154IF6iJEYOfKbjlX27O/DSokDv+a2mdmI4EriBi
5aBnjzzeId7Vf5KIMKgxiWwxounNygtcAkqDx80E8nAPVo0uYOKKuDJoilmzPwM1EkCa69l1YBAY
pEX9+lD1Hkue4L9hrUNO9TTznIMPsYLW3nSQBXH0op4n3lPRumezi4wRA4LNnbabVR6pNdvnrtud
2w1YVjd1gUqq764X/zPCSoCwvojvTUlAYWI9W9IKLONv2g7awbuhDiZi0VJ1Td4hQY+rRu6jkJ+y
4zZKy8DRAYanRBRykD9AxPFSxfq489COh86inGJUSx7BWgI/rrt3vljHCM4Sk/X4EgOy9JyI0fuA
GH7kXbZkJw2HSf+C4bIfSEkdq3B45ZMLVPwQcHGTSC1Q29PfNfrzAbs4OIuTndUYBYE7hpAlNGvk
LletsM4piWdWJmVU42AUFXt/SPmrqsCBINcOGkTyZYBg9eHdIEBnDjLqkm0/NzarLawVtyV8kNiO
4YC6tcyID2gz6eZPOQWjFq0j01KM0knIe0tLkR7mqt/NJg6u5pi/SS5cSbLClT7eq3Y1N23Jf90a
h0Hxw3T7nt//C1fuMP/kiWZmcYw9pxJME02OiG89LcMuMTaNgI6NmQHmNxjTbcqZCKLsMF54y5lb
vaoZ4elmSoc1EzZ/mt5A0sM0qPitFHYgPbE+C1uDldtJ68Rj/aroFnVB/nUrUqy/diZoA8hwafuQ
gPG3MmgTlNdX87bOLfBKwJ1T8KjUO0go18rsDdx8vTtlOzk9CnacmYIYzI2nG6olgR4NewuadSWZ
LciMYhmfLcnbATVTOWPrV4V1QYWArUBUL3B/Ap7Vd0ggOBvweEsjtqMrPyHH4dtTpuaqyOJuMy1p
YxChzjTucvhMPMiJjaT+x5F+eZKel572qC0K2sHerWezsgTti2cHehrDU24oo7i7bn20vOtaOhKu
4wP042SbtR5Xs1fGaILVO/eWARp6+z1FML0+/DSitXaXJHjADsawEtA+/jQjY1WNvm4xvM6Dh5SJ
FgmjeUZTKLVUVRvqYFO5+Grg6pvSTQsWJmyaaAZihGpidJKPAj5NcSb4cgeT3yaow7Hwc2PQ66p0
Eioley0/1A18CrBQzCBLIq/VQwtN6ksWsNblxMT6G6CLXPt8BueYA+ym1vhlhQbp4kGFwg5bX2AB
y7nC33M8vfqmPWZzK2+gg/Oafba5S5Jbo30XeBmp3YYITbmNAgEvhpDj31r9vygXT4Ijmq0BflBg
a5NZbt+TRkFuCDBvusRDBOeDjFfGp5QbzOjQFBf9eB0i66AVrLfL02FTpiIwhf7+2plkpoa87tGP
2RGOpWrC6mbuUIqgFr8e/1mwQEqXUNsTeAV/KuNCAmatWN2dsy+zprKXNGAErWf7yRGfWbm0c7dW
HMbjfK5fVecj9RlXgekcIFMkb5hkMux0/S+6Es1MOhpx3FaHIVmMCMe2Yv1BCBbwN2Dqs9hrtRi8
itghZ/qkI2pg+82d3hjYeoW5kVP2ODmnu/V8rzpr49UAq8SNhFhCYLOZpQDjvFZHkRQJJZuUfVmb
b8CP6jBy11JBFV0TlvQqwTLUoiGnRhwASAy9Rqpe7PNwZ8DSdArj/k0DN/NhXyg8r82hRo9hQ2lK
kSocCd6kGrWZs2EHP72eFz8DkRm7y7KYQtm729OcRg51JJhSJe3YqoLte0Q37M/bXfcJKrt7K5Mo
gKueGrHMQJ8q5ZkXKGtnMhhKeSbi4vNa673SQV03jlR03e7qPvQx6YTYvdwew/OOy7NBXN6VQlMi
dABjjEPmobDhmuwuTd8EDfstPD3vThue4ImOqAmaDriiswXIfsUnI8SmoEf1O8OFPDVRO4qTNq4M
RPBZMAXr8WqC/y0iWQwaqX05JNake7MSfMxSOQa5nCUBnKs7ywTObG45s8SR6Audzk3fCnzfeQx8
TnWpBe+2FAuWHOlGYl2PiDC7ExoX0kz9FjPqOm3KLL2ZOABZaxFas9gtn9/WlObiSMoopFJGjNmY
0/IUffkwzeuBRkVgIbkdB4iaLp/9W9LwjCRwlR8ZJS3NTCza64zs972TNmcmtEiwCzi+IXeTYMGl
nJSPPV4VDNNgdzgwQ+oF/2tAf2WpI9h42SnYoxi0Cc8dKVT9MRmLRxm0MEv2IE1to2l/FrOUMtFE
aLp2DkzVQ++8++rYCJ2Q+mVypMqPkDPvrxwnXGFJvOA7jzIHKrfRHiNEGCbNzDcbw892G0cgd8Kf
MhFGXVqyXDv3ltajS1JwJqD0UpOdeGqrEIBPvZngOYjbEsb2hAAYfCL9cBoHuoMcjWnaVDrhuV/A
8vpbn7WJY6OvCZ0uaAOTxB/66ZQFEFM9TsE+RSS4K0j2rwsaibi/uLIhg/YnbvFItb6T3LtGxKmP
KUqlft0zZw/i8+KsTdh8vfIw94+r+y0M2AC38FMMlvYcRN5J01jgBrnQNxJYuWcIHx27LR+n+ZlL
rgauje3/fyUetqDv0wqbCF0dr4uXp3HKg730y9h8KuWA3yP5ZvOvjtH6e7lLzf39+L0uwR/zc7UY
6pJV6r2IYPxF4zCDTE4Z+iod507Q3APBL8CraWecoDE8T0zMK7WF0jmG7RhrpuB6I8QHEuJW4Xs9
r7M36kfYwjaJSTitnafZgPJKM2b+WcJ8bjq72lQbmQFfWymqyfXIVLEJi34iPBHiX5tmv2Ex8m0A
9aJ/e2BPuAQpQlPu7K4i+oMEz5FLzpwHTVreVmGP1hoIbUQ+5qhtRD6wd77G8fMs2n8RRsHhaArc
lbpW3jPcXeb/PH8G9puMmBF7kvUFZEZj88VeHD/0vjvAYkcoRQdqCw3FqA3mocdGLRnBJhRd6R5+
Mm7Z8i0pNE0d1pB8vvkGhrIzQUhlZ6yUHop7SLf5zLCPcYKskSxFzlPdw0bswH+mnhJVDZ+WT1mr
+frQAd30d0dk73Z96cNylEa+i2a82Yrd60x9baSpPbXEMqqBgEmQtYrGHjOx41uyJmsu1pOJgXRp
S5xXgzdfR5stokIctPu1Ws/Bx0pbFa29ypw9vg9rODDjiQnigudgEj8Z1QHqa0DcUyASmv/D7wOZ
5XwbS8UWZssnw5vn1VPp0eKaakUGYlzHfgMJ3lJ0CZhM+phwDjvP0VQsEbNSRiN3UvCEMQ0HtXJs
F9eLtsE/P8Ca86EEirR38nmYBfn38ZzZ6gZlJ05cTKiDn3e032R+wfdp2OqUaK95dhQNtIVqPmKe
zvy1FWglLPGZMLgyJRbO1YtqEzUSC6UQNIUX7eIyji94VJUQyAhYViyvNYkklnDZHR2AeEQqPSHT
Aq/8rFiIKO3e9EVPV/hWp5hlCmcnf6m9jN1IQSJ6FBYOX/YcdYm5XpWan2CWT7bjqaJzoaXwVhRa
t1+LPriQ1PPDLtgehD8IyeaUp4Jp2CCkMYpW2hFqu+n//G/1odCLAv0uEMz9HK2WI2hFoNO6PW8w
xhw6FuU+6v2u7sDJW1163tTnghLBL3G2Kk/8ot5JUtGIhWIOBLH57XRHbmzkS0bO9GCf658+rPCg
3p2YPIF+8lp/F/4JqifAK38sAB6GiXuCjbdIComP50X6i+RhoTUmiO4JFLAP0FKxuSlyTTkVJLn3
so25fnahme3hvtQX2MMPfMvaAwTtSV+eueqWjGB7f7EsBDhU+KL1ZZ+NrqjjQiS5Kbxt89cb6tqL
qzCVXj947AOH+KtxMffjEX3B7qXSUWfDFCve498Ru6EaJ1BcKIA9xWNBUacCJ7ehCta2XFPp/wLa
Cdus1402yMD0XSqKmF87pVx3TM7aQJU7D9FnM6DzH83Ocj4DBfVWrHTw63CQfzu4ql/YPjXwh9aR
xW5z3EfIJN7DeeqYYVItWOw2uUg1uXUz/N9GXEDlHkLplqpYE3zrAw04nXxC30D4h18qmZ7uiWHe
hyjzpg3LHi/j2wWHwBTcpeZY+zVrvbQPyIC/K+ZSxpZMgun6U9uD4aaQ1Qn9FBeI/nlPvvaWBhxz
0wMQYv+X/7cstA0Iegq8oZ4GG8geSxoNQV6y9MaU0Lrxn1KSgvw1b/aMPYTWFc8ZG4lWkQV7c71h
2hTIo3RYjR2gMpFJxPYrHeX6FtMfSMItuv8N+EdDiCNEesAYV9sGr+oAv6nHXMn3UyIRcIwbD2/6
NiK5iPJ3vJDMJZe8uT1d0UK5Jy5ACnfszIfjPKcGIeIB1JNCrzY3iYC4E7i6XYI06GtQFrbJFQpn
iS/UTpyOxdMXnLMZrEda4JnjCk5sWi/AeQ44B8H+mg9HeM74qCy0OaQ4N07nvXoSvG2bFWT5vy/s
+2ukf8/IZtXy9DFSVlhXAVOhLUzrkGjyOLHdmEtd3QvJBupDYILdONZiL/EMbjE/fjcWAAJvADg8
rl13OSaHUmq1Qb/1z+0IGLO3/H85bJ5OwKKNf4gkcsDz4YzsebvtLHqQzFyD0ohXSdIDIse+tJh8
JARpjUQqFj78pcYFRc/jwdvnT3HhS5MEjKD+XtHWYnHNKbqMmF181zpsHDt36zoQvmzTUe0SpRnR
bocAbuROhNIbWXuUY/SlEZ+pjJ/tct0s1oYIIgWyVOmhWwzMylCZT5zGwI15GD0OdkafU7Z3EX4I
duOo0D1RtC1yrZTx/F4ynSjYtAti8dP2cDoJ/yezANm0quHf7devbcDcdTPy2wRrDc9q4BUHaILo
9NG4WdRX3LK+Ovxok2wBND6G/JVMw5s3vRPfmxPvDHnPTNPJ/SFez8WAP3irATfK5z10qk1H/vt9
j4kSmYMUruBT4OSL6wAQzeJF8LrjWtKAkG6ypokwswBz+cR6Eg54GHO/MEjwCmw+wOgzLkf/mu2a
to9aN/aDbu11M/D0HhOAXXwp1qtC8daSkX3KFNMqjCIYcx1hEbS9a4HNFvLLWrICoOnxzUfM0Ncr
AvmVv4NAYLzFLnf3GkVAHwzbzgxpIuZWjAkKijaGZ5mgVwiocTyDhAXofq4e8snw+ivf6kyv0l0G
9q9VeONHAwsyhp52+IJiqFpYOAIMxaV0BgJkVgZr55Ea9YVnBMfvH3HGrJjTj/PXd6UpL5+Ch2ik
CFlc88KtENwbshuMJ8mP1XOHNzRbieqhUh01ndnHsToRc5ZHanszcEMm5dEHK/GGbenleGtlyVL9
1Gth1z4lMSVOvrKaKqlSeyZVc+fFmSCMPYzfJCrHTFEJNbCOIlJQSM0Mp3RSQz4fl/hWmYEdfh9q
/DDKrRYzRu6X1NIk6H1gV0mtSE9kS9ZhOCO/FoPjzfnr6mKl4eEjSyEnUGhDjxM5bJ6qXXoCLJPj
U33INtsehzw9fOEUJxrCncal/xQxlGykQV/n0JtbEtdqv6I7Nxx9vS9Uc6xaizpFvYdeb7CUMMSI
hTpYJ9U6lB2VTnbHY7xiGpcVJCzBC4XnkS7gxTHK3xduiOE7YIGiJZAYvKg8AgyWQk171fnB/dIP
TPSc26y4TIw09pkDItc2TDWxiVlGVlV94BcO9rJOwKkBAr+8WgO8OFjf4Dnry24/aSDOpni+NhXf
nxVZYnC9meb3yJSFaxbRb5qARHqvR4O0Pjv6glKOnfTTqnuxQJrVBVXLPPX33GtjyKEsDKvl5Edh
2/VkEFJxlUX47l490/0F+6baT2fPiwj3baEZIBU4omtl26EeTO55LAsZMTP5YgLXRDQDibi+riTR
qLo1L1Z+nXoD4PBVhDpeeuGMacc3kezDdzNbZZ1l43c7FJS1McKWimtozKRguP46tArloWRzxzZ3
O93hbuu2rREV7A5Eli/GOFHPlRW6XRAuJvtKvH4s0t9tzocvBE8S2UrGlA+hNhMmCbXZxjPUeIDD
cQrYSr1D/1e1gLJ9YBXRh+vEjYg2XIa0zQuJHVTr2jOfDqukpxTtgxGuy3CD+7Rpv3T72sgrTyOV
cnuJ2A/cCZsptZx1S2IwE3tGI2XP3L4IQ8rhUy5Qg9hhKU93O6RSw8LG8jQmTDniZO3AssTO/4Dr
mHSJ3YBB7q8BCkmh3RzNTLRrJQBnw4Q2vUS2Pxls9S12rJbYFJ3LlNzSoyRo5LV02aea9JwHdrtW
EcOCTVnlpCyA9ANzTgamUQCcVBp1KPiY1IJC1AFZp7f/OHWpto0kt0W7S7gBh6Yrt4778DKYqH2m
OtHkMrXCk/p8zyoARK3eOjQGV0nz7vhKhGbwB45nCFBzR1RE7KFn7ndZq9Pw1WL+mIJmOpGVEG2w
xQNY9+uMUaq5zXEAfD2ZdYlbxQ1zEyRfTtBle9lXyQZNJWhAqe8TJu/P/o6eoe19vqz1ZVxJFfvS
ATLhrKx9OkQTaq5ykG1UtwBEjkxnLe5bFpoaOUScFSKLiq/nxHvgyAo/RqcH4YXWeQ6EaKFBWdt9
XJ5l39NVzpcfxjX0EJMQx4bY5/LQp3U+A3M6Rn70zCC3foREPgxRlSiZMHnDXWnTLb1GK0yE+9eu
4OEq0yB0tDPBmqs9J7CASd+MGvYyK3xpVLpPj2l6qIeJdUxryfWKJb3xyhu3o5qISnoDsLvdtNGn
q6RR4UHlJZzHHdMNi43tg4IfWmjjGLcUvxLhg7BtvFgyOEn67xbcnoVORxgbM5AUSW9FdJyTOGh+
JttaXLaZm83UJ8YbljNSjxIYDApu4/+niHWYdUfpdh4OcV0rA5OF7uE4oVGUDjdC5WfIzLlGYaUL
ayb+vo1ieSaNie3R0pdrVrgj9kcHJ+xASUx/3DxB6O8kHN9yBle7vcH8iqDkzhopupJFhlaQ8rK6
vsOShImxEmunCJUB7qMkfC02MrO0CcTyQ0CePPnvhls3aaVvxzjhr0JqIuGYdLPDEWiWAXxlkVqW
YnpAKePqmn33hCEKK4KxE5T85WTUFLd7349TkAP8OGgY7lUOmPM/+SmHjNGBxPTmji2TKTWWukoE
NJw8PfG7L/tomHlV6sr/IlZjv2AM3H7yCF4t0NmjtBB1iyJXSqyE/E6x8liH4QCaR4GeqsRa8Af2
IMc6GxlY0VdF7wwwu59oiaWIxg14zxMLGUz3rQ8CAIvz6pPRMRB5DBxqXLoIfyhvuXQHjhMkXFT4
9wXI/q9nuapI7iTEErFpe8bXMjccC41gATKvCEEBPDC2z6WFtTZFDFYWmpADAF/srH1k8pfJYmQt
IpfA+zg/3V9ZeUkeSBjra0SiU5FmMk/tbKeRKrGMaR8xX02ekNjVEs0JpRUeupgnNHw3eLQUo9Vg
uoTUA0mII6heYsb5CMDZVe5KJpzNyDh8qYuMLTqkRF+LAPCjwxZGht2g2heb8P/vpKZQFOar/Z1O
34EkzPeRFhiEC1WYVOyKrvLJ3vxaCZeovIUn4CMOkPV/SjtmOhDqqpKFi0SM+76gXrCmizU2Yw5U
0INP343OWsdtkvsT9dVGV3mIVty93nu+a+KxUjcAAv+WDlaS7B1bo93jr6et8CyexrApXkDJXyPo
2ehpuNI3nRmdGcoeG6uk+gm/SvQqJTBrKkC6kqGWiBBM4fnjQ8o5xuaKvSGxuvSs3mvfVokCr2az
l8M3dm1jB7vTb/FgrxkRq/obgAQasy2264Gf4H5K3C3UuPxLhP3MdiHc5iHotB6Dybs8NjXAV188
0oeKjyPoRlLb8DZJZEDAtdaxWazUu/Qx77fRGcf6XAHo37czxwShwXOazIX9SFHHrUEcUS+UliW2
DVHkmqQtnGxh25R/UiClTF6v8uJFXDN6dOoagDX16UFfAuY076nDVFdZfZmCXlQHS8jcnc5tEufR
sY3n4kovyJHIiAgG+DzGzOU7PylE+ANLolWCUeWxVnNzeU4tm896xrkz4bUMaSIxDtkp4YVde42K
I+r3MrLMV57sxQKcFrhpuNfjEK42WjuccpglsQ9k6sCbTU+bFp5oCvdiTD00qxGS47ogW86f4H0a
RVJPna4R0rffDIcz+qFq0ySWcJdGUMO0cCXraI3V7xgAowBohCd7OUZT50SgsJo690TFFmrR0Z7B
AXy8TLx39ap0DB/YG33gev7lqVSs6DzX1JHD2c+S0lASP4TJFiaol7WtwzqRc/zGE2IdPMvR9Gat
kXhs61FWMVZAN9UWY6owqOyA1oyrWHV50AuLhxEXQwB3Bwc1bf2+bdp+kGqdseogAayktjUGuc/h
xHfWGhy0zJRHkCHpOE0Hm9TAdRhrBOXeP6SEGUe5kNKLnc68op1PIWmx+F40skZJpg8B09IzY444
YIuhcripsbqWUaSKPC+bxgKD2+ue5oJuI1dLMUvgrOIROzl1BKmtgbM2STjZPvYtJL0BSPhRgYb0
bJR1Kzq/Xv/aE4DmA3IZrzlNRJpVGEDntO5CXmdeDTYX9fj0nVV0/2zU0v2l7kM0KgnrSUTY9k3R
lIgHbzoIZKCoKBj33LTjyN8dFK118SG7Yl0I3afgqGDb60C1DjDMrp/zwELq/qZFvzDkXt6gYZpr
x8Vpk3G/CFAPyhwLr39v8nligjvrPJkmZQVSQ3UiFyz/o+gfOyCQv3I81FFX6a0M3pf03daYgzuJ
OfSD/DFd5boFRmPBKTcGnuwT7YLQoZ1t/YK99vvJ/ltOMhLier1Tzwpph0bM00HDo6sQuirgpjpW
GbBnn3OwD7WlRA1NgLhrOJ6YxoHOHLoH6wJCmc84Abbl5sKJBVAHAPqmfIA1W1hAzZVSnKRTfHBj
IZ0l4pO/B03g36klppJhYkubwbWamGEqnFtt1ajMB2L0+9CUNRyrrg6pSymlup8BtKARDjcKLTIb
u+PGrix7411ZHw9RepjMLs5Hr/d0VKAoxTe3+5nrSRnDA+aCefWB/KJIAx74fm6CBnuKGSAQJ/PV
WYIAPIUP3btP52Lq0EGsvbxQPwjEsuSHWU6FroeGudGFUz7wTsN7P2HgJA4LojoCFmF6VNmInIqF
L1sCL6ZKK5H83cwDn775yUv0aAbv1EvDBoYiY3nfyWeXlrt5cN9SA3dXC0H0J52GrZMO8OuHVjEG
3rpqXp1q1zxfMvisuXlwDF26CF36Qa5Ea/Easu6xcD74OqstITO7rOqXWfTGPspj6FqSN5ixJW2W
//Ux9tManwBUnxYFjGbsfX5sdPoU+3nNHLOStUzYFdxoXxUB9C2rQuFlvGFWS0bYmhO0ZBBs2wnd
MsuNrufBNAtGD+EHgvGeSYih2a4Oo33ctn7HK45HrqT/cU+2NYPis5GcnsrLj276xkKc8/FwGSvV
gSjUVO32qJ+cvILH9J/gkGFgcCbWL+7vYHA8scQFPkA5qX+mtiy9DjmRIkYhREIh4IqGMdqxLOK2
QG1+uqKeAx1TAr2zD1VRz41InKzkvIDmdB3cB5dhRxXCDwkjGmovkoeIKM6/8RwbPo3SgcnsATV6
2tCzPcKVZuszw+Lj3z2ds/GHSpev6xoIlM2CwC8d8DSe77jwlyKoYHK7POSL4U62xbRhzr2nS7OQ
2NJ+QU752ehHepGG4tgR/m51Pdnt/kjxwoyNDNJpUD1N4Ib6LR+nOp7YMEfZzDrvsUL3x6hxDl5z
zEdowsb3Bjre4GgfrBb9U309o9dfkpKxHFvE0nBM1Ef7+ZXwVRp3vMbstosTdX13K+KRQBbnh+uM
LYqtSEQ70iZ0A8lMaxJ+/fxX3hCN3JuXiZxN/pO4O8NxM5QMtiof4FDxP1cNAlDO6j50y/aSBsuN
mCkuuUwkP8UBOLRGC/tG2X6KJTP+HzzjgkKu3a2xTzen9P/AG4FxtRyvgUuNMxztYXGaLQ+mOHFo
F6sp14Nci6r56KrCOuj6gF4ifKS+CGIjDDG92TLytphG+TcdNHXMRMA+jOyLWc1faQJKiQqe8Tib
4QMKjIEJ/+ZbpK+flg/PnorZkxLEmcUYkYlVRRZBe0iKtRSKkC7dJfp5cKiCJ0eXMSeUblsAEuPl
5TWf/FXNFfx4nHmmRn7k614spgVUv9apqRRhJoBZy5CDyYpog3SjuKL0ihM6VbmdJqIkdcjFSWkv
W7uzq+MeAUEjxwuXZ7STHV+XFionqQr4D6NDbuf1WTgvyD0WWMuumCPW+Skw/UOkJZ6h1BhYJa85
OCWgR0goDH0SEbq5Uy/crWGfNMX3inVBGCwUrgYO1rJi7PoUce+7QMYOsuczQf7VxIsO3TmTTNHU
Z51Utm+Wi34vc3FrPDB3p8op9KmVUAIAG7M/tqtOszLL5rX2IrGohfZUrGxIKxZxZujTE+slT+k6
Cb5q3Yjlp6Mi9qpFOUSPH8J1j7vSIYLGZ3+tren0MAdH4utyyYeeppig0bRe2HZmxfoNGdFL5bKm
252xrDtMDucVHAAxgsRTmKC2/KRp9NIlNPldugNLe6+nlJKZLh2rKTmDWO0KYU07OMMkGvJdqLjW
fzdyrurHnz/xphqeMsyzrJHchX/iyey9d61AXU918NfkdU9NFTeZl7Yp45i5CDqmnWVjX8P3HlPt
9cg/Bl6lFx1Mz1szex4AJ40ifuzrhLiUrm4nULgrOOvArKX7l5b41EHZfnp7aaCrvyVIFXXuwkVg
E7caY7TNZ2u+8Wgb+2+9g1PKeX6M7+kp8BeeN8YM7mOiYsZPNU+UXx9eF+FFIznLHFAlM7/PQuVt
nxv6uNJyxunHWqrM79aBBqUBmC6JmjRWddy6oAjPwpuX3DwBy7kCwqWIw61Be/HYsdgceRJ81faD
7XMvCsWAc+WOaas3Bdwbv2QpjL2ArxKY432fmvD6+7cFuBMvNTkciBPwe4PSMu+QbvoHoqMVAlGs
GwKuRzsY8a7dopKhF2PAhLKPsOw+kRLGrE6Byp572UBwdjuyZiR57nlihkMV56nZ2nBfPL3xgkNm
jUieCn5lq5ZhHgkHB67fKA2gXOufiCSeqe9t0rHhV2ERe9TyyEzpt5y1gEkJyiYY8Icat1qfB4yN
wHZ19xNk54k/T7GSR9Gr/ApiH5AgpiOpY61DBDaw3C56xNkyfLYCzcFPCu9IT5b+VvHq0vEqIOni
UUa5MWo37J/dpe/ZtsjKGXxorjtf3BVblLo7akygKIPd0uToh4x6FG0sAe4Q8eeyimdLIqVC5uMH
Q8K0gZAmcr+e2Ss1U17NnRdhXggzWw/xYK6CRVwwuJf6Nlz2JCn8X6pSAHwoPvZ1+Fgdi1WWkNDn
1xHAtgr6acxJj1bqqsO+YcdyXFK+2/vkezLfgjckPmHik+J14c+dpinVmH6VDb5qkHd4eK//lc3O
K5z9Uhr3uYMpJKkEKUtdLpdzLCG6MA5vOsyqLjIcBFtD2/LwDGuhwi13GDvT2uU7RMMPboQ06XeS
hnYgB/Ld5/9RhctCuVPcqWGaqst8sO1qeZ43hm3Yhpc1q4U/kd/gVDQvBljgiL/CU2VqO4CaSpBO
Sem6w4C7KnpfC/ZD86Y5LJJIr4mpLUXr2al27IctjGY8rFG6W/8V2JlKBj51nSfW2SG9PLTWowtR
kKmCb9U6g6q3C2/iwj9R8C/S8Z42h8BbuRfyT6sPXvI/pEUHRHk08y9zanxp6lQEER2DomfRW8Ih
c+nh/PYVSPggP2e4EM76R8wedWvI0PG1u0FPMCvGqVB42fQmkjSbXIQ+sWCB6Oy2yhyQgpIbSBdy
dr8kI/bVfn+fbdGVj8sd4247BiHAANPJL0A4DyIc7OLI3oms4yTbrGkn/cmz7Lb0RXt+chqQdZht
1sCFJQrP8vJEAK1HbsuzuMQ4J0Zc2s2IC+pB1zT9HobHq1mAc5dCRp6SaJXNHGP1bVCaP3r+5s6d
b9Vq7K4hal2uMrhCta2Sr9SwyAEIyH4y6zJw5tGYNRgai4+rhDEf/SwNxL8qIfnmsfGnhM7CHv1s
Qoh101q2pbqJPx2yk1KNrhdXXrhPTYf1Isg2MX+xqLXaRarA+T8Jr97VyhHZKe5yBsc0L1S8MX6/
1p9JzHz+Yjmwr0/cgZ0kSdcKGJXLySmOZ54qwa3HKm5ekC8XYii6D4NgEV5b/1DHtM2lLN9l2dPm
m7wK6tLuVObXtcI2QMyICi+VFH4fkHrkSMC9m7wiKXeSfbchDyvdPTM0dJNIYMOLzuPOiaoTrI5q
84i1UiZQfTLKafWUDsUZH3YR+GB7N7rvPITO4TqkSUp/WjoHaQs4JTgp1Ulkl+YJ2GJ83w7C+uPL
10PCMmD8v9yFjo0k+mJ9PJNN6dHO0KQVehoClkmo+AAbqq4V0n1kTODg1ZtLO5rzaDDF87+o5OOe
HR1x8gk3u5Ye/swA8RlZ3ggR3+bwiE3dtIqOYRdt8CDCDekI4aLk9uNmOOkmXN0JFiNE0hzp6K9l
Q+nRseplTLHETj+4PiOtsaMOgro7Zg5Xvrn9E7/DB+DxZ/DmQjR3tjwOUJCzPxh0vZWSmNpZI0Ok
rYfZak18tceEHUvpwmAcwY/MxTgco4RbNXGACFVAbabbIhlodJmK9oDU0P5j8uv0VRm/aXeZLV9U
QoPRGa1PBb5S1MsxP8t8r5r+Ct128olhyKgBCFdjDwrs6+Wb50A7TZ9o9NpNKpFohKCIALIrhCCu
6XRDHcg7euDn/dEMhmWkPykLc390/I3Ue9QQh52PUyXOMP4ZHcVmW2XhFlO3EebQIULisEnrZjZF
QBp+9ARJeM4jMS8i/ut9A3FLJsET7gsdvU2uNjmSrVlrwzs30KHmr72fSnVdrfVvNscfzia7syBq
DddAoU5q6IfX/UOs058G2cMvc/2vHksfpixXarYMWSp2RI1gabfgrzXGHAKvLrqagopnA4toWur6
zdZPMHHpamxvdTGCksZeGdpEJdXneaPZ39PdaAT0arIS51fQL1q/FOb7e8n/8kJN13VIzNe5r5lj
W6IYfjXs29evRoDoQBosYQlEYa12saq9lRjgZk6PIvVVoswXh71R9Qm/3e3x1fuHcTUZ/zLS/cNB
xidSBBzLJZxwJqfuxk/eC3mOCBknfPMEOXLbHh7FUZP47vcWqJiwDqDUyjJggRl3X3qoOrT+VLRe
t6tjGmzQVm2jFLcMKFgXNoN8cp6DeTS3JNNk5ODwptGjcbPPOnt35B+o3kNIk6Ypik3UZErFKE1V
LiWL7YnnMYOIW1+uLz1QvnG3Fjs2F87EJt9HR3m/skpj1YhybFPvlTD7jXrDgQZ8JOqjF1o40OvG
fQ7p8SdZpgaUKz75kGmbTgFmB5i9A/++3oGz/hqjguJ2Qb5Orw+5+2jC7CfkARvtLbDoY55Rfq80
bmHMubwPiAUTmdswQoOErhXRSXiCmb7xYRMWNpeic/QBHJ7HI8ZvrSBszucTglgCOmUiCB2bxi8D
m5GHbBYEjCrG67P5vnah9R9tz0cxFOvmng4mnMi3SqleL49fT8UNPZRZ+Om9iJaCuQIteTEtmMoi
LU3QrhPJLNdS6YslL3vWLbKhjOY/30A/F4wTg+HxH+9DeA8tk7wSm5k3YpNt+UjbDua1NQB5witD
ZXJForZLDO/SxMXycwTYv6W+/6Z/mQthye3Yc3aGBxiKV1Y/QiuDa93DJLxkiFNDm9KMQt8nxDNI
24wdzt4Nzkbwb6vyvbhFFTFS205n+X0XK5+8pKVzP/AT1pYgGW9xKWoiSxG7/rrhjM3f8srNpJkd
48GKaiXG7L596cQFOlPagR79qPAeHn+ol/iTthxqQrTCKMWFaM6GWitRm9+dRMbX3FW617zzwxQI
6R6fYGbGc1WWtqQF7fxg+lT8ht4K79JwpB01ORDU8s5da/Pi0+2m35AmlkSt4J/aE0uh/Age0kXj
3MmGo1HOtkSZEg3EQrsHc8v7CocWEOYyDhrgdJnDnKmaOmXEgnefNeUG3waVbuT7CAbQQ+n/7sEi
VOx/bmffy8VrPykwMEJw7kQHJJuqFt747skC24STPXwjhtg2UxiTZmN5+6d1aGqmRflagUGpqNvA
kNU5e6RPysDvghAxHQvHi+Rsp8JeM8RqOBs/SOCzTed9UHwPN+b86FY4bvBIP64R1QBRLIVUJnRw
0Vz2uKM+aBoWTa4Ta+CLH8Zi8uX3vu4hMmVsN2jjPNTI7b3kraZ9sJSBo9ad4Dc6fXk7qTAtipAN
KCj11KFRGplSyOhmFD97HVpUAtu/6Eeh2s+X3k9XZ2MrrwqyFRH6JHTAL4yBvOOmdAGUQ3vJF7gl
UZq6DuHaK0XWJZFzu6OrKGasadvXgf09BG1ogM/FS3Fa1XjCURDVnR4TinEMl/CZXBa73tXPUTZF
dKawUfnJurDh9tpdD8cOVJGD2vmRlxr94R3O1r+Cx2XA88O3OGvmzFnPEuqS+JYULYc9jEjtBRlk
V9A772qBk9jpFOjok0Z1Qzck+dZxoCEiu0j7wGAjhJnDNCjr0zQMGBo/Z219FIm+7v8g5fop1YaE
ibEG82oNJxvNEXqfHVAWCkom/I8nvQX/EfUtJyWZQr6U1OzrsBVgxKFJumTG8WB2HkOJVYu5SNed
99lW/JlWuII0XKONNIZm3DkmmY1QyUUuk59EFd5ombLRp0lJ4085F30RuaqUq9J0zshmgdJWejQN
+06hN5Fh707i+xKg42rW0wcpvxe28KBkHImnmkJ0Ch7NKqOFjmzN0nZ8/ZgSTMq2zzPuqD8iHTfy
dTo9V8e7FkQc9Qo+0EwmPeyw4ml8fEl1UM5iZaDqKURzyM4YT+lCWLlzH2BRHjGVff2tDS97ERL6
xGiNOXIeFoIdsQMwKSVRKyj5Z0DgIG+9Ki8s31PhP5aoyCq3JK0d5wpTohTG6Si7JiWZbi2pZeCA
VmPcRvyjyWhWxvhScZxByimXUdvQZdPKgU3vZNcsfgjjyaO6Evh4dBEanANMDYBGvZGeTkDjNHDj
z4y5oVgH4DeiiEyolZztlDuGco5ufAfH4bbjQDjwRJl/QcMaYqmD4J3BCMNpaWONt6Oebh+ASlgb
jB+ixuKyvqXqzF5ZIut+FIswWRtU8SmAoYbHaEp4U9HsPbSEY25P0gbsNzp+nPbRh6hrUDer8RcN
pQ3sGVs03WXWswIL+ZncdDVnlo68oATZYnJSH5S9sB8hKvHG5wcRfh496w/vrcx/E3ZWmaF7WROe
GpZSRSBceH4s4zCIaLEBG0jnJ0E22JZ9J0eMfUbxrbziR7FK8K/HIuZQgi6ggYrxkcGugud5h0L3
kvcgfEKhr3I8ytoFdhuAf1mBI02bYD63a42WJBVfj4y1Ymtq3GJtaguViKEEtqHaX18FuKdj18s8
T9sH3B0rX15Zf+bLgtKxCL1yYmt5ywtL1thdphgkM/tPkrcpAB5VHBAHWJgNe4u3StxSS2/rV2ui
A6bFD9Rc0Klbh4Vpv37GAxL2STGpRyNvKALSExnsgjoEC7kQ5je1vwfwt1Dpk9a2sa0/dnSZI+Dd
K0e7VHyGRCgJvOuvNWWqTxQRCNLyzyogU3VD6HUb32fJFA/muJTPyAtVb500OYl/Y3gGxFQgwzAE
QGT8W/Y79JHjcBGGsFgAQ3oB/hn92YZnCZ5BTBXY7bH3d8miLhfTQG8oW7o4NVw7WclsvzWtSr7A
kHF7MK+xgoPq1z1qs5Mo45e0jKWfW+yaZvGsvDKC5yfJ3+fxvnCmB4dSp5torPyL6anZq1QG/HOq
OH4D/17vPY959tGQzlcCT81zJyPofcT6FiyYNq/8bnW5d+NV5E70mOIMupBdcTz9x1/5UZ8KVGiP
rrAN9qPhKtYL2eDcFHeOiIJ3oLhz/bepXGUszB/Lk9rZ57/3h1ulp8A3G8RGokvSoO61HxD+AaMe
N1jDUdvc+DuNFj+Q9jcNRFA8sCXdCtuo2w8d7JGc5euvDTusqP0NVhLR/zmkTPu/Bja9tGOk/cUc
EhBPEWTeDt0XM5iWI1OOw8Dxh5iS65cPu8b8RjmAuzCPexhGRZQ49xugocyZZ49mKbtRI4Pl0cqJ
N+lnbGUbn4a01xVT1uNxbegS1k9dco8vAru+bZA3uSMCR1qe1MAvNvEtj3q171jyp3aR/4HoBwEN
xIz8ahUVONNaCBdVt5R0OU0T6Xhhdp+ihpCHjFOoxooLKPkxV3YfVNlm7UShLrslUzFtEbeZ/kx1
rhWI6NcaJfQTCjABIPfkIEjtKa9Fs709vIUpjHE9ks+Y9AhRXbnl2wzkeP0lTSCqxF8IGsNdbPli
9DkQFZnfBJfcUP5MKmdd5JaKjxEsjJE1Wm/eudZSbl+Q/u8X8uQ7TLx0YIvl1gs+tLrK5MeCScBx
CLVMCaM1vPpUHZXs9araIgjHMx3HRFe6E8sg/dYJmqGecOBax9dOS1zx3qpKdNy1UekxrbG+zx/Z
F0mUmXGYCychTx2/3xt6ZtJlhSaogaCD9poCQhHu7HPX6X8RpWellFLJzef6zaeA6PSFAhCa4Wo4
wQtMWM3fuA1S5Oom9V6JpMU/TXAogSZasGqOUyJUOF89JyNGXeU/yC3+T+YPKPRANPCMNGGiUBwT
4EnjrHcupHjfn962bZ4HLuc96IDRYzPGIOw+E1tds+BxIXKkeZekAA4wtTMqbtMpqaep60zwf8Cd
ODOb8umeE3/yohYzG8X+MyhBvJeabhmFDexWjpDzwLUwSRXSnSWLDCsGOqjoTdATi+zeOX84k64V
z28vzxpdye7GoTz0FsjB68+FsusA7KpB4o+07khVaP7/t5573nIC7/1IVhWrK//t/DQbDMgXfFtb
NxjHjXXdJAKm0KmXzPZPrfJIdcjJ8AzMyed7Thz/HLOl52o/LW9gFxXExC7AfnSC+8pcrGZ6hyCs
mRBJoiY6LCzX23W0S6qw/H3Csa9LMr1SGMAmKW92yttEbhIV5KwULpKGAX2tIJZuT3tHcIXN3Bp6
jIlEf9VwY8hWvPrV1yyDc3Ruke8o9HNjPtL+k8CmpjIHFBEtmR0hQvbc7Xo6dPoBfUCcoaD6MBsq
6M+EWT5Brn6hAxlZ1HOPHwasp+bfzEPITCWTiBiFP9tT8f4L5hHp5zpWdaG8Uz2c4BvHAm4/YNxg
0oAlMlqDD5YcR+udmmPZYe0TM6B8LHLoH+fdp5c7xgcd9uqu4Gpefe4OpUdTWtyo4yNV5g7eThA9
D7sCgxCsygmoNNNAH1GJjSGO3MaeYep6J1XdMdIk4cAjFOxFGD+56QW5nZh7y7JeJsOXABzq27kY
JWI1wqdlQ92z5Q3hN7c0Q7NUj8UmSdUR76Lz1ulm2vSSEmhNZWTTq9Ot8CBFcA8dz6h8WcBicDOU
3WrwEu7UoLg1N9UR6nFkIxxY/a9IcwwBR5zLZ1NqMqgjSvTYb5zpPuFey0ryKPqRYbDWOdw81aCe
TQQrQcai07OZx8QckmjGv7APK4wpmrTjTIesVDmkkdN5i7HXXC/cu+giIBvkczwlT7V+2UlbCASn
ppLbkUoZnA8MXUujGuQLeeMVkEZN7bFfUCatw5FXr7vX/Odl80SdBT12kJBZQ8KiKJCVMbIR+Wle
/1fuh5JLNohQI60lapMylPiMGg4t4IRmHIpz/7TogVOlOuqLwqK7xErlkAQubMdrwfDRR5xPIPmu
cCl8CM4ixfmHyAhtmXXNNd5pdYmWzWjo7Q75N5YkNMu+Z6Skix8nM0O5zS0lOTLcdm4Y5ZNcYWdT
IKGLmj/tHx2Xne69BjttCvn9LRQAV8n+gUxnGUDgif1QuV7mLxjxvjrYd5cNOCPsG+kxsuHThVVT
ilN5KmKSCWthUtdsDfEsfK9s8p9omA/FL/Aaow8RtAcZC4y6i5tSPCob8ToVeNJ6MIMElafosQXc
GbwaJiC/pN0iDwGl9sdsgzFesJzyXv8ZIkxdDjbTf1PIKd2g+ZbnE9lPm4uzS1aygbhmXn92wd+4
vYc4+4s4xuSEXOJmRLcfNqiZMduwyvtpzVKJjnwyq1MMGZKr0vd0cZocKar/ODuWrpD5F+6xkep2
VUGjWbuTCprffQ7TbPQjrACHKi9D2+oKat3akROrt9FfOXgSFtnrtGaRnX1FLRI/c6TR+7iwX4ZG
g0caP6KeALb6qH7AjHS9R807lFMlLKRQUFKWYP4n2Qajc+yuMOaey2/E7ZI+/XYbMopblVpQLc3C
lD4NWVDjGKlwzWSDbGlAsDhXneVyqbYKWAtrtgh+sJKa7OAlNJo0+suDMs1Helh6YMgYB4Xmx+JF
6KpRRDEkhdsZkCC/AdnmowQ3wxQOi/F2HyBtRZ8t5W9H+2C7osrgcjtmeuRWwUL6HAr3Y8M2ld8F
2CymIOhcupxHw5DgDd5k2xpIien7PMB8I1NHfrHTorFaPaWe6xYpDavVS6dqNyYNmB4K5LBcSoFG
rzkvtcqSH0kzV6nldPgheROEVaYdmSsD3McYdPL5W5A//QD34iaS4NE/JQGZjLnEU3VSt0DsYdkc
8mm9r0Uh86L46gylifEudmJ+ie/r98lsAhUZl0gyUgLmJNFVx0xxHx79o5JDDpKoGOc3sEGhEzp0
3f4dHnPw0QsDOR48AKmeLbvd2xydVjPyxhSnjmWVJX0z/u4C1lmU9js/rlCe4xITSsyFo6pZN8iu
MofQLsvmB5YTtDHnPGy28TyW/67iur3692hNK5jJ2AAlMCHq3mzr+0Ccb+ApYG+ALnXZUxAcAnIZ
sQ6FpIvVbgBrGsfrBABucCjQEcqsfRSd9SMyUfC+vjNIogUVrjGbpFA/a6SNqqrXvIJxriNcQFaY
pAlzBD8gf1i2V3OCIqIFEmeKe0qlbRZ2qgPFKZW8c47J/GyQMvauo0b2BSVK34jBz2bgRjGkLzab
9S8AHHlTV7DjYtQQj9RmAj5g6uzscEDJh3PkgxW2yvWplWMmjw8VU76mc5RQ3dBC0QuXUAPsBh11
c2dSKlfNqkQpa20EFoEtnOiViXlgmwWiUuppfpsUMKpjO7SoaCH4jueI3FS3It5wCkiojhAUPaG3
wUTLwYKrAnYFQux2obLEz4rOjjiZJNwPNBe3duMCLLWF101bmjwTOSPeFm911RrqWxX6P/Am7Pf2
Z/3cHzNMvQE/x5H3qJywB8bO3gb5Tfvt/1jU2eF+wekSp27afG4oEKs1tGM7+jw1bYePDt5wWmi2
TnUlOhIz/b1IJAJNgUKFP2tlnerEIOA5MsY9E0Cx4GLf1tZp5vd3lX44qYjLMSPBnY3cfaDGdhQj
Mi6JBGvyN9/uWjyYZaf3Uqg0Fm8VMFSs1DB/6pZHkryZkEhwdpuPlfsf6agVxotPc3EDmzjaVJYH
lhjCZMOFzAcdtNs6QXfOEUscf7+mYoTta1FRp5Kh3l97u9rBSCBZHPaDLPTFyJj9uN7Tb79DHfbm
n86AXRI/kAABhuL5SJ/E8dAXG6JcdaCl93NWNsyorSgoJsOFfViGvAW+QJsWUNuCMX9zF+p/nAA5
thU4i7igcqjna2YSzhIGFl1nGVs8eKDnzfL1N1WVrSSPPLjCniKtgXCJpIw3koCbrOqo86YYL0D8
6C+otTHiT34ZFs5AiNsnucnbGyg2TbBdVG3xoW95KCneT2mSKP1H1LExauAoOgUEoJyvOl7jEyZO
uRzloh5hNRWm9yHEBMK78m1Xg4DGcsvHWH5orIHjnl5jOsrW4QCKvjYw9wFzX0rBjIQuAjGTGgaZ
RtDGK6AQmgZmYv1+Z+Rzho/3wiCwk59DOkt4rIr7SGkz0Z8fmPOLSLeSgwSlr2af/7/TnU1Yxnu+
d1ygaQywHaTmwhG+UWrLORiiizz4ID9y/sQ/cPMhMSPVZkXZjqLX2AGN7tOp0/id90yllzA1l3gv
lCPv5bNKTHTWY5SwBj4UYgJGg+Kqplr9Jma40e1K3IbUsPgNcXkfi3vkxqUr/dTamOkmIq7KTbG+
HmbWS45CCNql7UyIpBIzEwb7uGmXRO8HXh4c0plIPFKfeISACW+sGgc1VIXlAS3kwN+CDrnATxnl
aXLNbwFUhUxVXK2ykhWUh4kqnpO/aKjTmzx2t+OOnGzg/VzgPPhNFpAM6FkCqwaenMzE+HD/BNBc
AlZ3xJ2zzp8YFQ+04cY31uYIbfhSChi7LMzJuYQb0QaAuD1gFbDlyO1IC/ysB3ehPFhgDMgimHgF
5InRp1qe+0PIiOJHkCIZT8hNm40BB+0hR0ghZVG68B+aedVSRctet8RYIQgDQRRgDOyJ8lViRh7w
yg6NiQBWGo4ZGBUvwgOVPVl4GtIJOWJIqcxqsQCuMzszz2IK8hpAiWLGOBM4TWKc0KRw4bZVxXud
KwGQEwysmJkhpzhw8MfjMXWam7MxtZHglyC2CPTWfcLWZgPepgyKLQYQSXoYzNFysL/4VP5UZXn0
39edYBz8qegLpu43Jq/K8YWzm0sPnhDa4JB9AyylrAr/sSOzR5ZWpu6F4QP86NXImEP3iROoyHyl
GY8DnFbWdV8T/YPyCM3Qb77dH696JnoxpvCVHWXJfKvpQc/1Ruz6S+pKYUETzRsL3f4zOu39oG9t
avgoS3/5+CmdO3GbodX8SSRdekY06S67hhAK+5oWcysWbILMJwME4CaRAW7Sqh67448FAUIqHrwM
S8hKyjmrF07eQLXzGY7KFq1NgNJACtF+YscGqDKPjeb8v/iFBvs1ochCWX85zP5nZCiyBUBevly3
jQEGfl93TtnAle0FEtSNU1RzOswtcAEc3iR3GOCZjYP554kABVUJur+auOI2VfhGXQnYXiHWPns2
xTyWhCOnVhRP5wcVekoQC1jxOXaGslzHo2QF/GA7KTy1kZXQrpNnTcjQchVWr7iM2z6gUKYpZLDd
Tu4pY/7chnlrkDPb2FnS7ro8Yj4N1j/YqR79yz02GXVAYOx7yVl9jdQkd7RokPemgSljQ0Ak4+Zd
MiVGaCaq5RZMCxN5Lh5YKiZJdL2RpD3rgdW3Con9lkGR0mc9K6riy3OXEX9SH9nHdB0yjce3T1Br
egTdT9ys13SDcdEUkc2jBmrblK86EIj3glab7YO6oQxuywwljKO/xHhEvZjyOH0ydzdpk5H2/1r8
heFSFIyngeXctIFKP3VvwYtQjsZD7HKmDob2IK7Tw8Y5IZgQvOowgybufFcMngFJ9H2ueRo32h6L
mjPILoml0nuZptXzIGSnDvX+AZfFYJpiHzs78PJtsXq50tLnf3ixDnaQFsQ8+03DI83Z0nbrihOL
ad9BHmwD1EwTQN+gqmlyxoXJYNfjK58r7cR9EFmPnpvErupXBquyglZgBjvJVVaLI8sTIs+FwrRN
0G+qQfMkcEBoQ7i59+Go7hOsUvf+b/EmJrfdNIDDy/kVhmR4Kg3SCKpOqhsV/EIU+hmffR67eQv2
UGCH9ea+eqz4v8eNiWNExJIR367P5HSiI6ZJiyo1rIvyqQNZni3Msp0/Xs//wAwmDnwV4qs35CST
S7Po3Ens1k2ubZ9Vsbc31YC3npndmadPeCh0NIIlPuvz4u4HUSYtbzPcBkU8T77n6120ZdERgd3/
xhVUoOC7UO04lPzL0Q4WOcFrbF4Xvm4Wt0nm0RyuFXdEsaN8+sSczkk8i67ccRGi8TRxz+ppVIvo
VtcZ2pRinK6e2DSYhCuDf7thPjDfPVZH/g6+pGXml88/cJr8DzsFTevl/1imumiNta//GXiajryp
8sKHLu91sIfER/JPxZDbG6kdk2bLVKJChNYOthzHfPIc9aek1ByizpoO6K/MD6LU+v0/NHR/glZM
7XOUYlx4hGPoAVTRO4B+0p0VMj5t7Pj+5hNJ/ESERyO4oT8KJX8S9pL/fNUtpANwrgvl+iYOn3en
i8WCC7inxxxv6e3ZvzaYmVf2GCj3M8W6lJ6aJABPEaWUnkJKLgOoxb9eosr5jMkdNsxDMpLnSmoJ
/7rongeqQG060dPM3nmcVo/xMIhYG4N4/2s4X5U62NUtaLhu78KKNKf7EO5nYr7AY3ZKhDtL++w1
qMkEGRhKnMYYUKc+I7GF+HGnCCpTj7iSwOg4kffmg4U9X/DVrmRgCsEGmtpWo+9ZQCd7J2/ytI7R
ffXJB7idUfompApodVapPLLEXoRB+OxQjzxQXrG5dVbvTIelN6rY2mJ2EKTZFuut+1g+5URWrOtj
K9BmfPsTmnG8K8G3QRdzWPUOaecsGpZxcPBAVcg2QmGNablHpM27Nql3IEj/QbZX4XZiQGjJTS/S
aiHrhmJuHxQKjO1IzQaAoqJOWDx0rESxdyihQRgIEUteD2GC5cNeE18m+nwxh1+SarUatJI+4fnr
6w7aFCW5fQWoCIh6baJLbgdBqPL5WBY851KwM/qxt/4/8xl2LWr0dMM2ncBUqShs5oaeRnPfl39E
L7Qjym7idt5gK1oT/F4x7qCq/ZU1/thJ/6tgIr6ixUwcmVfGrEsSIbsfk6y40smuLtl+6odziz9d
Umqb+hcKXCnXo2Qcz/nmN0F0alPHW4PriT19hOxjLNz/1OtfaCYpX4R8I9CnBLgPmSBkOkRv3qkX
ymkbim1iUOen8YA+l9D2HfdJreMcG4jz9WFGz6/t54pfk5MlAW8B/G2eAUG3ZJvPK3aks5uaqNbp
r5DVule7Uxx1VjgxJAxwAbGaO154Ey0LF95Vl7itWK1isxiEmJXy8G/JiPtlOoz5az7IcKFC3mOf
8DSsoCN4ytkr5x8NFnbIlNGQHCHc1fAe0S87L2F25EDHTj7VT7uq+mc+GzU/8Sp8147MEX4f7tmk
lS4fF4CYU9iNVsImVI2N+aIP29IG/vVvNbn3+zzRxA5QjKwvg7lu0QIpceO1NuMGrmkxMLnHKTh0
soWO3RxcmJd30vFPAcsoAq4hEKCitxr7LaLBSOJ1J8TBqjrOLMfQj0AACenIJfFWIj659VZ3xsvF
Qrh7LWpw2sOMWbeLCrjO1y0XQ49UJk5Xssi9XOPBKOkmhY15TusoKB5t03Wj0pmd+/UF8rsoO7JH
4KNxBN32jtnagNg8Oy6nzAk5mh6kYxPzfDaHk2saXv98zw/2bovOugNwFDU3efsJYKQzsw6S8tAh
+LqXa/mfGBgIb/kAHnIqdYfK/YpVzB16VAs/7wFmVvJL2/Ec0iBzGlj5moZqcvJgcQgru2VaQtze
XxOvni5SE5KNxKKmQlE8QMB6Ca4xhilnHN5qq7Af4B11ai9PYkUmoLJf9U3E0iCD1Wpdk0lskaGK
/wt7Of1pV1jb/TGwDCA64t3bUtPQky9QbHHuPmTVajmt9/D2C7aUkSsXkIHgVFGJ5Lrb9deopUYb
jOuHBzBhpmbNeuVHd11O5uO4cMaoe70m2HWvyRe0tNP0ADIPzQc9ES11ZpC3SSi3btd0PnN8nF2e
gnVcyaIzHKgQgK9+yvK8Pyh3ep50DtBB/gwYpofJb41YY87qnx/nFnZUPo+THlrIWwKYHsL5himn
s1ON6iaq2fZ4rIC+pTHJTAtvnjZnEY7OMxc500kCGSlyStxAOwN17hbrt8uhfqSjQM1gpD0LNFEi
TdPea14GcS4gk23ntgVjBeLZRPhEtfjIg15VqxM/usCRtja3IHaCQfYnAk//8sFEOEF2Al34ABg4
A8IwZqyMYrYb9atMGxjvtIPMMIbxC7SOvp4Snq/UcT1kmfGuPGwjezeiQnPWdUTIdNVr6Oo6s6Y+
IrgQa4v/cNxy9AHeifav7yzQBe99SOu0E8m2Rz7nelD9gNSIIT+avR9Bwr1Hzp1mhoQanASg5Yyh
pS9YphFy54fGqzdguPOFSbBy3L7rfT045gh/fK51Q3lnnxQbXWQ6HqK/Qj6Aa+G+ZQkLRnkouD7i
CTQVkKPPGUWYJrb1ALaDuzwTHf4+DDnSBBSGj4hiAMIAa6HOuCsbS+DP/0ABvhX1uwCeHn11jZaf
KuiIU2kGtn+iyq5gtw7b73N329uj+e/rug/7UIwFQzXGWnxgVpEuaIBADAZq0ocRmwfuD78olCGF
P9PY5UapmYrWQljncfek4Q1oFlsVDFXSDQJIZfLVt7B6p2o0na+66sIighsJV4wxnTQmnyduMgAR
TfVNnJupgI/A4QGiFdpCqd2ga//bR3eyOmGo/Nmr0rHB6+6yLLjIcIOGk7jHfCs0/u8DikIAPgiT
oYhZYNOaOy0bWyeUPcD3kPX1UqbMkXI3Fc28apMPK5/fqdMPonI4jqrgM/Hj51fuSNfr4xOY96px
Tc5GFnPBOM+r4eMlBjuAxKeHZa4Y98NpjZKppovofnzyMMZGqkAHc6wwMaf54UpLAAfdNyIUWpbI
8DzpTHeL8SySC8EfCKF9h55A69PPvK1Xh/cecS483M2MBZy3gHIhpAbLjIFZvjA7Rj+OaoUPKf+L
Sk5Xz8fOkDR5ZYthnrcviaNl4J7jwdYYoSchjZIQJDhGnxM+RbFpXhtbg/UT6tQgNWr0H+YzOpNB
RChsGjMYnzhn0BjQz1jirshmktbtLhqyuXRbSlLCuS2yp5K8g6MhqASoEuSNARJODfULUguJpWK2
YzJZq3wyEckXftdH5FdmBp/vph/bo62S0DFKdTLoldQhLBvaIWzMx3wvDMF8uCUGCQLq+aktSlRo
faZXri5QMt0TnvnU2UTZo0/xZWxSzIVlH00GCe3tAxSQnaE16CSGieLjNcMe3bxocBnO5hDZRj5m
Wqq7mRI0EeF5o6NEzCyco1LUSDSjLWP2STK8vTcWzPtarkri3njPxCf3MCgZSVpbZKQkQP6OFexL
yMqhDaNh0IAGaQmar+Ew4UvQGp+FpWjVPiue1I4nBoRAWBYi4d7KHLTmwJaIEb6FtWHWMmzGESZn
6UQrnS2+cHSzOUgZQ5+tTPIDGdFNwx6jn6sRojtcUNGZGM5PrZk/Akx2rakoG6WvYymcHgBdpUj1
yUewoilCIy4UJPSc7VgKFcrW1IImujUJWaB01ERpQYH+85qDjUv/55X7Em5ti0Qi9e5RcVoRNrGK
BKTrcySQfoHlN4cG568z9K73CZY/3ADvkj+43CqNT8g0GLrOAxfZxZHhr2YRe5N+4LUbP6Y8sjmG
FROHUbR7b/2e26dCYlFyU3JKv2o1cza22QibqzfZ/gfcmL050FddJQbO3oMytgcuvSIXsqldNlP8
ofZXdTHvMGOauHRm96cJKBvMl1BJFvhVB3IBIy2rvhUdZ1w99r8RmZ99G+buMGya6lbe0hsec5bC
s8lA48gHTcKpBOM8VR2/AAhHlEN/uHfmKzJ8dJV7SRinRuXMcIvDxDe6MskVDJfWzsHp+76IJceU
kmJ1WWUqlpXD8vDtE//NnL6eVMRj6nmNnV6lwdetnW3Kh1XXQT/+KvtBYx8bI/PbdA0KYEMYB8rY
TbAFrWQQSQpuRSfFXPsjD23cc7dtauOg8f/i9x4y+hiQ8OTKh0MVX//n0lOCwwaXWaqWGQwVwsHt
tFP3DV34EBPngRIBIqmTvR74w8A/Un2q7mMa/QCIouEDh+XKwAvan5ytT83TK10gTWVQsuqIRZ8D
Y3BTMHiI3rtRVXMgIBHUDsvzzdQCkyFECM1saEkn/AifbO53TaO4lapKJNcOT4ErhPfzfDNOoeC6
ILfIAQY8P16xKPaFvb1G2j26cEAraen2WcrP2s6k9DkdQnNUs3gtl/AJAJcz+jkng/5so93mDKkw
brlwYW7iXChGc070GxJKF/tb+oYYpQ4YdLQbgN1gdXkSgIEYQrt9RKKRJxZBNGe/Mm71K1gmuWTJ
+ALxyYplIGE1FVIzM00pfF3f/DXT5gHS46HmbsguTFB5+ODug+luujug0Vy5tlL0sWISsupBVOuf
hoJRk3HbGyuW1zC/RO5ESkpzm31n7QMC+5QPAMUdY5nsMXI0oj3wm8DazJYLmdDLINKIRm2k4tZ7
zwN7xoN11i4KLMkdQ4okPAvQhD6XupCrEsKD8GfUG/eUlmsrP39vzkvE/4RUrd7QOl7P8SR8yBBY
3Mc1Ud0Pwn33UrRXl6MTxqApBVmP3mF2Je4/XSIuDGO9MLHT5xekAMjxmqrldmYHbeTtV/W0JkNE
M/4W+SYqRL45pZNUE5LG8YtOe0TOJVcw12bTQv9UwSA4n35EvDMD8tysYt1QgcJL7Q+2oFQUnZJo
fv38aCefr4jOLjLeB8rjwtj6Ume/hBKC0b9VFKP6d61xiHYsVYDyDSZ27TBeq5NRyEZS+en2m/Cg
1zjm6OFN3kXhv3hCR70AfYBQdiUZgvTXuMbgxDuPkbLDPiKLh6B+r5NOWGcfwnSHKui9GiEbvHop
iiv9k4LkK22W+hezgPzqx1JtzHuTsvmHvjaW5sUSu3scCKMSWSKz3rOob3VUo+ZCKik0RAtPtQPj
mMeUbxNSjEpLcxx8hWrUZqs03Cue8tfwMncdifIeygQvfZlMhygIagi6MWGRSu6mXZOjidV9VWQ+
tY9VDAwooS+sE386v71tNzbU/sruixbTRO2MsDB8dlT6jnxKv1/che+kUIq9l33ph0+i/ugb8YK0
CYZ+/GDPWCjoQ2jrFMnUqngIMOMrrJVgmCa68TpXTstgRCj57vnlm4HRfZNG2mMXkCTid6AgRNdo
Riy/9rAhJvHim68V9b6uOas0RTMlkNSkAs8ezQfHt2p9yRg2G9LFPwjANABnyhTkn+DjKZrsqkvG
oc7O9gG5KT+3KDN6VF1xc3knDYc8QFKeC2JHcUjznJ3GqjmAZtjKR9PU/k4LxdagPRHO+5ihLi/s
5ZZPzVjEO/rXlxWPCLu6k+lg1ZEhiMoaTKcKz0wCC30lEJyR4sfUK0VUzhXjEgEslQON1q/uPYA7
2UVaslPaPZjOmXbR+CSjEEI+vQv422iga17nNE/G9/WIdYuIz6vf/uXUcbJVTmtI2VBmwKlUqYBu
AwB6WFGZwZhlkI7xWIgz0FjmtqJDP9cdpkncuGt8myWVuNvAqHKlbkKYLtxXwmnO2UrYzyVibuNB
R6DyPH/2sYIweXqQdaKUdpA0Uu66ChpkyjoKTjuKXNpTavWDmZhhXkaSW1OmAn7sQtSyZ4z5PnlL
eZobPhTf9dkqB7D+WewF16s5awIpkGgiN8Ah0pJEy4VkCda5WSluu8rq5LdHfXpU80pVZSvITKVe
hY1KvnEWQL5Ee8VD0IdrnTZKmn9i7zC54pyRjVAPuli4vIFq1NCdOZsH6LBZ+05DEv/Mg5QP2D1N
yRsfTQWwygy2uRuNfTS6FNzsXiP74puOnrzP+DuLeyTSGBl+XJzfM6KQCk10Dh6SziqZ+fCIeSps
lqJK+FmwaIkKgbyexpQkNRquahufqAKRuZf055ZxdLaNo0ANbKF3lXNxxZ+f21hPmpdxGIinJGWt
JMRYwWfVbuYsRqUlikByWiPKoh9dSAoSVUjPPQp2aMIacXsTAb0cnUXxqzTi3Gqzec9NLyrIwwqe
9hYDfeoO3BrUN0LTwlt1eV9CQqu9ui4FaRGYxsaS4O7oOxVTYc1NqANq2EC1SnGmK3JYhkxNEe5d
maExoltXDlSGxYPQVzMBDIeIKmMgnJR1obXYbRs2Xkiq7FMgYGyplNjTTV8vwOvjNypnLk/Xchnx
64K7aeOa1u5jQbt+SoFCmfY2d93soRlk6k2wiKW+pwjohwtCnsAEdW4v9hQlac7lDRLbYGH9+25H
4xIjNfoT19JUMTY72gQs9tASdBIVnoJekwaxYfYU3B/1yBfSk6UW0SR7CD+IbwsaQsbUF6AKqKVO
7JFIptEn+tmZMpyNg8yYyat/3Jet9Sy1r/yyeq2Y03ge7IEyeI8Nr6w2u1OtSkuWDUg+xebr9BnE
Z4Pqr3fmsCsxNm2/pAfI11T/xhhCo+mOdeilcJOaivJbBQZxXRz6UkLYZ7W+wl0onoF59C6N9jgb
DFAAThTm8bVcXI229vZf28VE12nnRzj64o+AJofqz/eAE34f0F+zJY8CUsnx+tZJA2I7NqGQFjKm
4QeYxHWkd2juroyOGYOY4HmOyV5CUOr7x6HBPfWIurxjm0uPIfV91wqdWHFpVtWwi3FFm6NsQ3Xo
A2dU/JoLGnCpLuxbQFoLq+UER9h/MUAp/qFuHm1xO8gVkRtc2+cxcv6En4okuyuN6VB8XgEOy++f
gibz9m7JOWHlIPfJL1CULa9CU8br+fi9EPVnc3AedPIULpxtG5RS5seEm/pmUXhoeT7O8LIBCwn6
B32kH7qL07yfD3ORN7qUuV/gsu5XUhv+p4S/8LaEkiX+GpmCmt48U3n4w31d5cMbuETQGTeJqIQ4
pINe24NXY1ZvhRAClr+20wnTEIUdLJYQ6YjDsPSSCpioTz6sUD6SgdHNZ5FbgupVfvf81mUeULUz
9a85822cTvRiFxYfpLuRbiSSLWOwyzZMmBAq1Mu1ZYtKqjiw29NcMMDpMNNN6IpLiSlZIVyhBcp3
xTws7TTKoLu0M6Ulduehhwiae3t3JcwVZl7k7NaLau6e5RMohHC3ycNRTpBJAEsd93RtWTo16ngR
/l/luMKmwtWB9fcAoK+WnyL1p7DhldBe7tKVQrijj33RKLuXJK2s7EU/dvT75bIjr0xvi+znort7
iDM4xm8z9sBhtmTbe34L1smwmwOXMYlMuzX5TXYi2w0bivgqxTlCvZV5CXO5Fukt+LSDS9/E0L0q
6+TsxkPxKq8LngY/Jd0RdiYPY9d+jOeXAr+3J3UkIzTGe7DbSuaLW5YIzYv23lN3smWS99RAWCEP
nyjS8aSLy+Uc5yuVongVi3vhMcaKWTZ+UEH1GlmtwFU+6RLH28gEYSYY+A0bltPQbm6xCjOUHliS
5iPcSCorox04tbTL8A1AkkvMwKc/mjV0YMi0f/tEmZBq4uruwdniRxc6Vs8Dry2la5NVkqYQdivE
78FO6MRKxddS038WQGuU8jI8ns//13PXvOtAfRNnZ1btydRP3Arh46rDZnrKFlyo+XbAOrpQYBPw
95tHKEzraAPQaQqJ9lYuxZm6CHKfxpcnGQuYo9j51pmRdNXk7aoG5zfCQkjJPNNjwEvuM2A35INV
RYHcLVObxKJGUB7UjvEGeZ1GYq2zzPFzC0oaPrtwMfoB4FkGbWlKSe1cwISws4Ls9Ah0d6srEXdc
Tvp3mY6gQS+m8Ad4AbQRean/SoPbQaZZVPSnT3aPd+50WUM882cr9+g5SzclL71WB4ybt08j+mEq
TJ8/irafVB7nXsRBVJp/kLwm2IfvpAEWHQl5LClg+nnr76DS6ofSamd9e1l1a/AUGKyb/us/YL0q
PQlCi51DHDIKeO2lw3bZD2W6e6/fJSMpfEGYXoYRJzAcJ2NkXnANaX4ssbixvwfLDx01BA42LIXa
XwohyE1rpv9gRaHLKHvtDSRJ9sjizR+vnOxBShbGw5wk9w9I+qk6LZ3l0nOr5SUxdnalm3BSJ7uF
IErmnQ4naU0PXr5cPS0+aIBDRFuowd/Y8IhBxwk/eCaooy2rQTeXQNWCB/sl5DQWc0Yf/qODjFad
Jood09D16Ut4heSRVya6g3/T5OMOeUX3WHH7nWAc/QXNg2F2qesQLzZIp6BIYehwb7Iv18PiCRBG
PnVPELp6s5T+HHHZfQmq31Ycjn4RXqkKEZaJHCN++vWE3R5ntjRSzywOQLf0BJAEiMbJueC9Agwh
GTorO+TcFS98TCJU55rzGXigGlr4B1gvvqe8k7P/WhQRmYWqTLuoNv5/3JP7yBgn9b0NbFVCvCv3
P16Iw6AXXwpHK597ozN5MGiyqVwZl90XtAvS2F4zEQReyPcfuoNCQtX7e38orUJxjZXuN7bzBcj2
H0irao3U6OXviR2DoZLov1jz0PQt+wkzidbHJwmpD0o4KI7ULUqOl65zR5h4kbS+6Qhq+9djiru9
jsmKp/fKfuYxhbChA9yHolxh30JX91BVvTbgUVdPXSsfyYnUUXIXy2Rd1JcBXYkOqBIaij/4nbxL
Nn70iTsWYVdA4eNibTcpyZ2Ad0GPDNpRwo74GaMo1y+aHtpNrNBi13UPWZVcDnsZJkRDBavZyJ6v
3bFDjOVy0uottqb2YHtDWWCZcjjlWSz8jZ27Ll8810GAXs6BrU2iUlt1pvGVDnIgoz2YsrkDcPp/
yxS3ua3WsrOymPZREJT3fiIvv/Se7q7Lm9Yxr0jT352URC9nO4FbFJXXXZgbHMCYao0V3kyvplf3
MFp9z+lOugNIdOy8FzSDSOvl4Jlo92ET1doBubyckkKfHRrigJvsi8xPSLQ2RtrL0Iuxpk7gvlZa
eBtdp9bLcOqxXw4du3lq7/nFeS3cMVWRdOkgnn8D4KfaCTo/kbAblPDrLtJrxmibb23XCgmoKLlm
sG4tbgLDkTb7Om5nomByYgirGFFC2ohRavcJpHVkJuK9i7zYCkL2grMPhEIzDLFJaTwqmB4WKECg
rbbQ8+xbnhaYAWFHw55mGnU20akyVIc2DBVonk8dn4QlPAOBtX7TsWRvmE+RE8mPgT9p++ZRkCQ6
r2m9yCOsO8TT8IZq4+Amqcj1Cxgke/udnRTb7dznDZ2uhgmbZYaV8Jupt+MSxf9aPTonWjzgVFvw
BC4CxHJQqBvb4/AG/m+qVpTnUeS4EB+clVbbHivRYf9HoKqvOhJmYpEUefBBjHcWbltWkUGCcukR
lm1OA+wXOlBtH94I2OmtI6PxbLI2DFuMzNNtXbisCQRGRbFhjICylsKVJfdE1BOWt54FFuVPL6db
Nlm4OvsbxH2KSwZZyYgULtaeHM2Dl98U49HMBkitrO0c7MquCsQir/JW84s7Pe0fxHA3U/RZfKY8
6o5WZOdeA2d9LOUXKmYcVRKbHIxYh5w6ZisI5BnQL1Z7z7j1niSYqQ37ZWJUDG3NxUO6WqERGA+y
YkVfovETnI7LydL4PV1qUawyerMrUic+5YaMH7wViXZuRg0f98cRgpdTbiBB6xnFUaxDr/75gWme
kYVZnE7KESbTmx46vMBCSzZyZe2wzMsxFkSJDt7FDdNi4P387221pAhFyGveiOY1vQqGDJrs9T63
GswvRCrk1nSfNONpRX3EbGkQjErytX6IvsblWrQ9JXaFV4+7XfYkSvrujzT+C7nWqlVgYplRyy1o
26QzeODbofjk9qHhl6HMHHrP0BAiThe2x6kxKnv2cFfxCFSwhwYJkPgvFHEBwh+IXJSUXYVn3E+O
Q/neh+ZV6i1uLRhJEFRSZnv9ybbm5rUytJVqrq0EaanjI9Jr7dGOJM1quxxZst7pa8yCnuPLBvqZ
mPhW48HCr6ggrOWJ+EU4kMAwi69KSXiaAB7tvyumj5+lx6G40gsyId9fFVHVQmh4CMguNWuLrj/v
JMPlslfOEOmt2FSqaEciA7aNYjn9w/gSYDfKNa1am6la/H4+Rvj0pZNiOInZOoznLSBSYzXbN0OY
nHUulOqJWNsIXInua72N52Ws0Y83mrXfsKpdvaHf/fte7yf6MQnzYOXOhn2gG4vPuZG2WZ6rNuGq
9phXZ16Xz5UnTott79cKTAI2MbgfIZw8RFBWGYW12O59csqHrOXlYCsz0IQb+wrLyTY2gp/g8Hvz
kTbtUdj28cjZ4ZOh6uoTZ9v22AHP+Q5HOPOh1FGjhFPlODGsXSZNL0uGuFjBRsWOpDCggGYQuLgh
TAqv3FMHxrawBTsCz1EHvy4SKGczTNN/2VCGKqZcEOFnKsrQeJ5x7WjmKk80rlRanKyirzlrt7sL
w5jIzaidSfyb/b+elRU4rc4aJ/eDnfo6TWp5iR5d4b+lY6mjFjeiiPv7UZe3gQoHTOGszpBVHcQ0
Ts0XlOSp+/OKljr5qdlvTQccjmuSnlin4YrVmT87TIiA9iJldDfJiHNdH6tWPtNc3zWZz/GyFh3p
bATD34Lxgs0cT0qxUiQU0eA7knPD554lil3K1GXHz+Wz7ukQfLX6klFXs54ClIa2H6ABxB6lF0vt
1MB1fXCiFWIvms07jOD9QNyG40U8qL3XIc+CenJ4hmh43Z/qoO5GMpudhH6S1yH5qAhDwMFvywIn
44eaY6Ga1wTu4c0N7xT7iYZOZmBg8F83PW8R/LutfKVvUTrLtPCtke8WQdwGyJmmplQto89tO5vq
FP2JFfj2NL7VU5XAo3t7BmgACtWEuxX4Cy7WeNoEOJoBrgbUfCz/nNUwO0oz+mO/DH2BKgiUJJ3u
E2VRT5t0Mg0a6jZTjQl1v5Zo7cR5zUXTyh8JsN1D5U3reTUGXuXOJktUNjx21Fn7Aw4gginNqx48
D4K1ij+gmj6nZZf3YqEnWR5YkmEtnk3vZmpif2j9sJDdO+tjSfBFrsrH+2916PrEkFXPhgqJ0+Eo
vFTR1aCh/VbJfxObBMdwCZygMUhtAqGzAxvlLRzYqyLuu4b5erVXmK/42c6Gn1zMjFw7PXzeu92/
2I5d9hLztFlr7icDkfRFdD5VdkcEowHaoUlYyFZ8AxkN66YHFAufDrhujf5yrERJpH8a+D8ySMDB
7SqKVudVUNhuN+leS9HrAnsocKVqxSgkP8DRZVw6PlMnMBiH4HxNwbdLvfEEot3MDWy2QsVjXgRK
UG1jXlI5Wz0muDqbupim3Z54i0VzCNpFy6oYqWhvQlZpF5QB0U2cNbKRBXKG6DGBGPU0h1ngeNAW
50TnR7vQUWfwxHlZ1/WJkxZ+21TcR02HWd01WQ/De9CkabrbQ1EsX0K9AJBZvuKnBb7H9CI45UE8
vULkoexwBFT2keepG7eueNbV6R3qSNKeXJTNdZ7PdEidlXrevFx44cQ3dxZtmhqnZ5vNu0UdVMdz
9eN9xdX3xMCFZfW7WEoL+TbcWcLmyXgIjF8tPCfm5TiGTt46ZU3NSJ/M7uiQkRzl/rqCGZyxeHIA
fn8RBSuczwRDUDAyLqA4OkD6jFijTG/PbQ42ByAQoEe8CBNjp1t9xkjA6aC/XKs+3A1fSc86FITC
e7xDHeVx5Zh5J5XzAWNRJ2CVjve8fi6xxHZyUQry9t8VXmZWb1BkaQWPZxYrK16SOoUbVuc6O1rc
LcD+cAdCpWMNLvFmXfjut4jNgbvpbpmy4KOozwt2AspsC18HM8NNfHdaNohJ4BAf/CNGSZTwB69S
vPH0imAPA9LwuaqkgOa7WNONmMEGJytChDvXPHG91E3QEe49qJP0HH4BWOJMIacRNXcigjczoEFn
N/m03Y1yRLNF8WU1/9Rqnk3gE/BqaziDqwXC77dN1v5YaoL/9VWO7SopAJimD0CMYSsDJkcXtcRc
zyxTY6WQVf/tdRvLmuMnR6Qpt6MH6+VBzCcHFYGVM0X8Casv5Y5I46QApxgMo0Y4ZKQft6GPhvp+
ps+DGIJj0ldEkP17qtNk3dxWtgs/dG3Cv6dGtWd+2Fa29PLqCNOLnmRqj9oDe+AzOWdSvxVGchBg
8VvJWTrNiwGe0ZK6pH72wl8LIZ2KpS7Umj4/TW2L+CFpa4FgVjroNGoCOQRezRy3W0WFyFRd6YcF
dD4FF9QI5lurMtrtwuylqUgA2x6Wx6gsAeJqQ1fbyGbGIQp1O2Uk6HqPLZcQ5XiqmGA/ddLGJBHH
fakICg9d0NrB5AwQ5/ElWYEu++2Gq7hKtlszmXwf1kxoK8zuAq1X03EOu79hV13teHJc7c1Mo7yy
QLLnno1lwW3xqGyiX9IwjUjYlJSkeFx2g85jf36HdWmJoxk9Fr8vyVBUfvfQde1YCEi7uqJVSmRY
XpVD4EOyNBcME0B9KMXWTt3cwNwmuqZPYb9gaKTpHg6eX2vW/dgXwH0RzUyGA4Zd3oEBx5lMqvf1
XJd4roawW36OGg5WaVjgqR1gijf62XKOWNLvz4d5lO467GfAY0m2e/FAGZXSSiDTH7P3e5mbyzH1
OgYBtTkZeDgW8jsUEq24d+LGhaCFvQm1c9iTAr5INp8AR2ps8/5tjdgquZIEhLmLtrrB8AVgR6WP
LmIff9F7SFMCL7fS1MEl4zd6CWP9eyzwDefiVhC7bhv+iLqtA2tUeCEv5+h+HNc9g+9XHJLaZd2b
7WYA7Bsw7mTX186iEpaTGSdfP3js7dePf1xfdebaEu4kM3QFdETLlMTjY9U5Z/OVvOTmG/qz+INL
ZHF/NA63TrHmjoBEVNXwCty/G0neAShAfU6FSMWkOGyMDzyoW/OMrw6hS+HZ+xgqiGRC5Msf0bCo
M4vz0Vq8FFy5MU0Xhbf2PqknTIwn6ktL6dRqPUisXSE8sLA/NQh7sNjl+ApoRHMb3/MSeHiysE7b
PMXFVBsAZDJCUkRLbFeWJAcC/lS3CaL1jo4IjuSj+AotCdNEPjrxzoM62q1vXMjgBPG+8EGo+qC5
rCfGweqKrZIByzLHCdvXTgF4VToLfXkoK1jz5GPM5CqD2YP8CmIWhpIdAcKivh3pQDtrphLEB1Ib
Zkh4bHA7ZE3eXCCTN+xP75GWxN0duk5LLosKLb62TD7AIcVfXbzkTWM+VSJktOgmn8Ngd6kJpYnS
2L/uK4HKo/5s/8x7te7U35/yrZn5EmQkwQbBz0ieiSEFAejgvGeqeYQSWfwGkuh/a1+gKkMM3OSF
qBy1vANdLv3V+grKT38/vJxf/GxA04s87UdAS4kuN7F8Uhjd3Xsu5mMzIzj2B9kE/+fqv8E61JPL
lMcnS5BeH/cBsfRhrwz8aOCc5dlmsdVKsrPyJJ2w4/Yo+kF8AgrTrsU4AdbbBVVqmadEETdLpgfa
Vq2C+ZP3EC/K8oXvcqsiqzehKHN2cO8FXqqvPmwFcS73zvPkUnQDnZJrDaUo5Q47Nu6XztwfuxU9
Z6Co3DvCRmXlvu3pvTYyaNctVRf+i+GWqZi4G/rjf5wDGpT3OObJFKT6E508oJ2otHa+3NMz9tqp
TFlhHcmumQrcaqbf/lVg0FLOdDzyt3WpxH9L8loESgckKgXsAenbvSQa9/4xEnXFeQ2/C/kE5RTO
82yUXOlabtTcwoEX3d8QJMpQzL0yaG/nxol6ZH2jBc6mxK9GtKdba/fH2gjjLF6EklP75By4eiUj
8OwqqQqw+YU8OS8Gjp0VVe+DtGldgx9SmKwA7gNzwMazbj1rE6CpgsW79uDSywSMk7KdiQ+1jaPa
dVmtgJ8GNfoLGKqthIWxRFIaqzV5cjUQ+1Q5gB9R093pDisGeEvtY1ggzaj8VOmx2zgWyrmLdDAy
cpbJXNpqQ9iKi79GYzMRpS0OV3vBLvb9GDV7EoUeAZAeQvV6phXr9gjbOAKTGA1tPrnGfYSN25zO
p9CgCVGoAUkIGLTququUY/mG2mQQu2hXj+xomJU9mhO21ui+Bom+9ltVrYqEeUwEI4K1+80GuUnC
q0yUer/+RfaqnXdU0eFh8aLgGP0u7HZuZms7z4xpMWx+m2TqbtpMFhSwi2BALIfrhZkYQHhSLoDN
gs5KoIAB4dr+1RG7GwuaCBAQmZmLtKfbNOyDDZpNqh61kCtpf8U80ZbceJNEna7OCgnNHcxxNzJH
z08ycLgYOPf5U0uHwuND+3ZP3bn9JQT42ah6sT1m7+JdSUo5sPKENehpNtzrTi+o32OY51YuV4sI
7wnQtxuFsO2sHnVbQQ70EnW+JdZw6u9QC3rWw6RX8iwzg/d+GOEBLKL30K2P3czLckCYYnuB5cSr
CRWHRGrVMCpQ15rWohjUWa9IXHkydEZ0IDACKNn8aILoXD5IFYjyDdUHvN08S/ChOJf6SFPyPf5P
I/dNYCELkXDnbhfBM40jBw/IwV+EUyDso7OHwwpRZ6C1uaimRP7PJXgtSmdtd9LE02mv2kB6CIr3
hyu867kUXEs+9N8r3JKGKWz387S9Tknfh90+fkmSMH4LcL/YHBLP3R2HmQJneLLq0/Ed2h+OeqV3
yK0sO7dIVcAA6mGri8SiZwFscTenFIiEOIh3diiwxmZ0i62mXP4vpUkSjr7kVExnNwjxnAf6buOR
BNM+/ufyH4NGJLKi1E13DhF0P6/0GtjKPHVcvRU4HVa2k7k0NmvDgk1t7y8R780T9adzPDKRBhfv
qUYzE9UlDmt0BmBcmcuHZCXAWRb+KUjlYorUNMHr2GLxGISIWKZB4XVIYRdJZ8W+dVcg4R1WBxJt
M4n/RLwk06AWFpG/oxbU37wuTH4TWQchwTiCLYBHWWF73RzdfRLqwa0wnLRwbIT38J5Ya2Tt9E/+
IPKf7Wr+qscPTGj/Px9MRSVJgM1rtVVC8pXduCNYFZ7JdTOBgt2mnScCSOxff4/KoBC6aTXAVyFT
m6LR8d51mBlkLjFHsD1i+Cc8REmbQoTYllohlCKsoUXZfpOV/KI9R+hKodej4JY5kBHPXikS+wmV
DR88x27dc6ZFy8bbXl3gtzxO8qv0OMYpcnvYfYAk/rtbQAl2SJI8MsQe5rmEJkCllaNfQYEG9mW7
cWKS9RIMPIaaFA2Nh769X9IcWhBCScozBxZ3WZ4V2q1IJ7dEhPbAzUziFjzBojeXGAwPPVlHqNqi
AGCi7X89bVRcg7bB62b7hEHrcLFur2UNgPTax0u1/OEsCrQLAjXUnMGyRxVbJAh/HFv0B8Ngw9mT
LOocSdnvpafAAotWOFOfQWRqype7FrGLbpAPoRC3JBEBEfSgMsEINNDLOS0KIDg2RLGtUdaC6210
rzGgqNuBYCN0G44NM6s4RMajOrqUbZvWvfFvUZ5BjuHrBVQxoh0R4oAf6j4sPXHfppxQ8YwDcZKN
moZfQACSmwmZX2wsIb5vShKbI/zqxLLqjtc9bFr1cHX159IZaYeu00UhPK4wETLOO84PC3HQ+lxz
UVkPoFFIC2fGENCVz3W/g+94Nl1AsA59kP3WKIjMVnoFauOzEIBsvf1k0JIAuxyXUn1Ozt6oYCZh
JKMNmCPJgYz5s0mYZS98utDV4jTr333jzy0MNsyWQ4aJSRxYiKPiJizQskafesQ801YGwkkLHbyZ
1W4/Stcp7NEXVoBzkwrbOuzdnJEe1gcsDetqWAp2D00bdppidkHRjFodYm6HnKiMXglWjsYbVBny
DicEubMp2lBuiy9jk3Ix7WNBtDJNCXad/cKgjZ9k2K8kSpv3AknizbL0TtY0LEX0pkHtCx+d7eBO
Xcdl3qNT00xKzY0qay1KnM9oH6yRVpPv+Y9IRDMnusvK8I/wFwcpVSVCPNvMySrWGYRYx2oEDzq8
w7BLwybzBT7NoPFhAa7cp4NUJ+VePdSEcYdcf7jABOZDJctL8+Icl18gLYnGmjo+xK/tvu+QqsKP
jB7BdaIlHDJlwdDRuepZTh3hMD46edx+Q9lHo9vQh18GHLBQsHNTH6FSknpbgwOHoBNH+B8TMY/8
13mBA840NYm8T7C0DB55pATZbO2ZymONzRW0+3UZz5Cs6ndFDaLjOAEeKSAhyluPHbDLPoEihdO2
wx+2nRZLj1bAKlsMuSVQ51US4m3bFszQtNXgNAQKcNG7Cem0HGJBt7+FCcLzVOkHTaKb+OLGzRqU
PESakfdDl76dsSVrkh92DhUOWLq8KoCSjS4beOIxTtXp3zrQOOGsUSLDcJNiJCbp/0lNJ4qamktI
7PkexLmIsXoWHqHjomaVLTiI68/DK5+VT4tmRP0l6XPc0b9eBGwLIS8/lIetQBgwYzBpRu7JjsMZ
hvyi44uiX7UA+mnkXyMKEePZspLg/LiMI3ff8SpE/kpoaGteZeFBd4kJadJtQuLjSObt+4Umcn6i
wvfz4jXx4ZChR8wlS1ekgiOWZK2RW2oKV3Cbgv/iQ+3fIyrV+bGL2lA0IJGQWchahAbhFscHsM5m
GXMjVoot4m8hoh5YLlObdIsro30za38CxAUwbkqbHSzsXpDNDNWTDGeNxnAa5sowDP5CtdIUMpdz
8qY+RdWpShu/s6340kZUWKcs+roaydFDWYZwc3+Bxptx4J4XJbTD8o+l2SjzsI4pSpE8XjcjDBhU
NB8hvHKeZtI6gv9Swy0nsxOWQSdd3BfZg1xuvgD/iqr+zoE+gcJiQYS74UIAU+RXsfMFT72EPjqe
RWuQagKKRukJrUfoqmvKaYmY5yLxxLw2WebP17aAms9Kibnsj/lJhcEHnD5H0+m5Lw6iAVu0LOHl
+QmBDh9c4d1Y2HfEdBCFA5Gi4d3h7B8eUXnHVwwwv53Fl7ziU4bs6b6yQKaOJthhUva4g2sXXJBg
BLTqvGLTRkYgQjybCyXZ1sHP4nE+kAtZbaiDISW/OU2Wze6uNKTKKCuTJqHTdtA5DTUZiS350Pez
QO24wHJ7YaE3ORqmOgAdHksoskl2cv/qsauXo8iTYeg/+DnKlHTDh5O4P25tnkDTtnMMHRIawIyG
oRmxLQqNB9eq5uEzBo07DPSIy9+auZlfE6HvXWkZoyLjwearmKU1KkAWpSSoDhlOGzNLqNDSfGtB
jcs7BKptpwqsKSn5+LHNNlg66DKbXiqT3yLkcFkDdbOg0A88lLkpg3eXhT1ItMVqmrgYHBtj4Kmw
/UG260eTrgPn4xNe4m7bVyoAWcUegdXpsVPgusSB62dMi1CSN7auUrZttN/Rul0JS3/UJ3FdcMjZ
k6HbDdNDiUVU7BmMqfPF9AvPC/drzuCEfJ9csYt5aBoEV69w1jVjkk/xMBzpM9gLkuKYqFo44fzO
VxdO4Wg2Kftm8Iw77ZHKFkp4RY1w8mOPr6NPZbe0lk+wYRwDP1gY0SvnUpWtZbSQ2zxTmoezcdy7
P/Unn5X/RRTmnejVUJHvk6g2RL5JeTQUH21GjhtK6SP//PPkCBHmWyVi2qPH65XdIr/E2VW4CWb8
VYRbjGi9TuN10nDrReBGDXzmgbQgzLUMFP33TwAxGlfajFJ3z0wAjyWD1OBTFjRA864QvANtzXen
Z1SjmAWXhKS0XY8WoYPNeIfg8iSwNJMBA39/sYiXnypRZJi06TY/EuhJqgSvl6Qcj28ogRuiULIJ
Wv209EGWOxnouTlmHZMG2NbTzg5anFBNWGC220aRYIhpSeDysE+OIeWtXcRK7EqHqFrgBlk9qv4c
ZhuKzjgAoAfOsRvD5myt0zMiOPK8bhqEMaWoez/6GHApaWY45JDXnCkH4BsNSo9fTFa4rHnGqNuG
Jsze6bPxpd98XLk1rg5ojtyoW16ylrOQ2Wsv3zyOeCguf9yKYmY9Q84If0Fumkvv6GT1xgjinKJH
IM0kKlUkoziWU64mNLCV9Qf2NPUfOt1dEJVAf1UZFdof6eRxLvJFQ7Ymo4y2po905GzXKpI7LccI
PVH4a3Mj6Jw62BkNUatd7jq9eHEBa1GgQNclpeOnHdG8eFJjifZYlQWdePO2AcDS6T8+zN5lWyt1
Mq5G/h3V+78g9W05AzddCMEOKEcM7Sjh8/5nCPKlVNxMO7c3wbkAOg9Dx79/khR/PCFsCgsF75ln
LMW+fi5HTtCnZ+wZL2lDDmavqW8uywhkEIKDFazNWDnuJQX8qlSQPVTIzO3TOFAvvEceicmZzLXb
mkdSuJsp41vtlCp0efQAKFXafD40i3P7KApCjYwzZMbm87Z7J7ls2ddVLIkMpkYwmDzZksz4AQm2
oM0TVJAnjV1zYeI18msPUdBY/jv0zM/PXFiWTERwymKC2sogcEVodJW5waONfTr9uf27rwQxCXed
1Q5wuJQV5B9+TtigkY+n49mhmcvx4XFDdusLFGTS5nVpWQm3MGL+zjKzuxjYLIYr7+mOwLyNYDiW
+v2ht9k+Yzjau/0sA2Vuieuq6hVN22RGHSg1Xpwzj6xl1/eNq31eDmH8YoqnyVsJqbUANU1g90lo
8cbrT3vf8RcJSwyjKQfLW4eAj3IMnacqLCYxygQA6DpGOtcBWiLwK7ERs3o6x9NXqDIGoXNb+9NH
hRKsatfkfG1HqZ3j6oqz34JG8plHwhiHM3L7ilFUE9amal44Zz7GQwaq8rkcUUpWenMVNBXBrD84
zmiUA8Zb7LWF91Kb5xqvj4SqNNbZJ2NP17OLx9fWgo/cl2fmPM1CTwXjUCYT6c6GWM3xNoPiMKxQ
wCPhUjb0stctOoLso3tkC/cGJIfGVUfom5cLPvHOnbHV2BQXr0uFlTzoRurtD0KXXwnb3zvDZNFi
tPXrhx0HyTAda6fOF02Z0jj105YR4k4KK6Xt/DpgI73lkS37UuoNaSOZlFDaEZ3cWnDqGDcGGCbo
PTvtcD3mOcluPeUac0gzUzphk8dfEgNQimrKOF1ag1w7l6RMIFhuaPZkJviEAKIqw2eJ7UX7xhEx
UOL0CP0FpkAt9fOalMWc8SPRofQrxM0AkWYFLAGhL797GYUXAw4lZrMuCu71mb8E3z0PEZzsyisO
oaqjd7Qn10CyANr+FABp2KVhTl5GsKGKWztwumC+ODzyGIwwLM5DVeTwG4db64ZKyTY422myegZS
sLD5ZiiNmLKvtnslqQsMzpevYsT7qQ+3e/vidYQckrJV433lnJF3LWtAqHpnm43lRB3SqLr1Ru/W
krcmPQvmwtc/QYOJnkKwUssQvpRA+Mj/cVI0nbtJwkZnBfgTVIReZ1dZNR/NvOT9weymXqLtgEpk
RoV+7Pb6Gh3JKP1SGA14mAVvRtmN2nA3fUyt+DlazRPWtFeJdaA4F63DhicTF/pdFpnGV2L6DLB6
0m8WJ2LdW0jGPtbkh2VwfM4i/FL0gaa8/nqTj6axm6/wAIDk/HgIBVf3NTI2Ctp1d0nZl7YBk9Zc
ZH61Z8LEaldx1ufMLWbfbAud/9RR/iCp0haqRMzbBSEgjHlAvjrjJa4L1397efY0u7EE6fud5+aM
0NMmLHusBbIfTKFEC9z6SdpuS8z/ZetC08WyGzwl0vQptR3W7cd5vEyt3ge0APbMPnj9o21q93cV
YpEsosEatjfx9VFlo3vEKMxagPfVWXZVxUXRgNV6IvkKa5q7n/hzVpL+pLEfA6NJZCrH56xpsDGn
yVeGJGzLhm7ROq3Apgo6qMYohhMInxvCJU7mUauSQZ+w1oxceinN3boOxMDz+Rtm4RV7SSuV3SLN
3+yWvKkYTWMeH9qqdUKW1JRMTzeWPvPL0WkrmOVTp2CvU3/YUqtp5soTbJr5ukIMnsUKrr8XiDiu
ALTsOCkpASgSeX9q4VZJmzgn7wuCcXT6rXud9gyKGTkYveF02XM/kAWbkWNPpoWyEB4mx0dTOakG
iTbpTukEcqSlH1hkh0Jx0dLfkUC6/dP2DvpmHtUUrAz3qW/BCtCAOvhsNMJ8LRko35B0RbQ5WBal
mhIs6/B+QkLSG9nY2XFRSFCbhNvabD8+wpQbgskesf2bNbQCoAHT7taJxOq1mLqiwTHh1FKp/fCP
wEKHqsqnDy1klvLlSw2dteoP/1rF9rJhJmLsW4mhJSyfKg1BkoUMds+utS1dVfgDq3ifRD3At7bO
8CoO84KGq+GkOVP+AEtYFEKr8QbxSMRS1TTVdNlM++gCQOYh4DEzkFTo5uOJJ7b/p9VM7i4aJtNB
fUVY8lK6SlxtufHeaDO19gSSo/aRvw20foS8f9L1zQb7r8w0uDfSvh3YvAP7bjfqlVP77/CBHuz5
NGJJAN+JM0sCgs9RbloZxUeBDJhByLP8bdQ+qL2RyoxIh6V1zq6OeaLSwT8t2vAmMJNU0r+944Ue
76P44s3JKy2K/5GBa/qvNhmOgDjpUwg4Slbnl/KSfsSaDQvqRIubtjG1LkoAGhLE1/xSeveTAG/F
KSDsvoGITNVEsRUnffZbSaN8OYQyca+NAHcfpoPdHYcwmHNGy+4w8KIZY2gHb6rgUPrQeYK2/zoa
t3LWl697wdGp+gzGuKeLGO7FcZ/DzN57omQ8VU8Zgeq00QTpmbjO+HkvgxrcqFYmSB8I4AuO/Xqo
dAOQQ3MziE2xpuNTn9BnHYVD+PyVt+u7R/2grOKHGlZ26QppFikJ29JuQ4QmmgSWLOgPrAW5Gurh
udw8BAjY7f1FIsetEmhbqu3tAf8ZUsGnmoVZsYj7+ZQcfufvrXKgAkF8YI04gASwW4e1QNO/Z5c+
24g8fiVMktTG2TrhB9fm3ceEEcHDPFwXVtuCiQhY8J6KfLzGysvBX5lOps+ahh+7Wcq/AWyXnSp+
g1KmSc51p1O02CUpsW/5NQGvxDMrXRxi8tiHmkTJ49L/x9u+4f4ID6Qik/a94f8ZxoW8b9qcWuUm
aqzpOfdT9YCI7nqFYbaVj3aonPPXRa4JI2abzOFOzzLjAGi0q+VrVqI3K+UOCP386naJ7Nr/MQqE
OaqzA3WXy/mTZIEiRyxOyaYZUsD0X/5IBGwvlEoNzhKPYAFy858DFlgiI846fkibiBPTEDja47Ms
Rzt/eYccvuxOJDBEg9QEzolee6xtJzef6YdQezrFq4U10naNUcbjuwC38DiXfaJAPGyowAYueCZP
sypI11Ydnw06vjImQ3ssM3n3vB3uYiBNN1nil8wcqQ/e297iEeKnhu7jx0w9HbpkVbVfgKnSTOI9
AeqD+tUabe03Vn1JFNePhu8Tn5VqKhniYmgPAozk0xpqKa6GGF/vdslW43uescrzXUsIyfs9/CyA
ThHvE8eQRJ3LZvp+sSj1kIby6/2Ta/FiCxOOwuz/cR6I3Gku+pIScge/GGRUjGV1U5ApyvGgRaM4
if/9X2VUY6g8yZiOxfUdt7f7ukf14Ba36qTf+qIZ4aXvi0Tt6AOJD2AoaDfK8TCY9w0So/zVEN89
MGdF2bg95Asib9wsbhCPBiiESFR2LGjiHxAWj1WmreuUnyODgqwGZDPZVS2iCyF0wiSgjPBSxo6s
jfZnyMsaywltULXBmvxUQSO3ToxXDGmm+Zxq0ZeJibbR/i+PhwzT+KPqV2JrY0ya1IGGjFaaEfH3
6yX+rS0YZ0HHost2DblIv5cwM9M0U4QXwLmlP2/frJ+msTybDM5UmjKXTKOw2/wR1qJlzPRLwlP6
YLsrBPlyun9lQJmlhJk62RikdPkGvuqeFMlP2XOOaxoVUZ70I18QmQTi9GvlqeQgCgQj6ARZhsEi
QZfCNiT19Ok0/N+uQqRbKF2graIYBw7cjB8xTEMtWjoE1pwdzuWYZp8xqwOCHzBOD7jFTKV8z6WB
jOySRy8bzCZWGLEkXHqSSapNnRe24/RPeNqBXts7QgRLWX6t0CC4ATsh5io26Pif13qcDsv+p1fQ
gB8tCoMZRbKYuL0TJAjQMxNt5ZvbQfRPdkdMprYIS00t/TVUoe/Qpn6FN5zAJ93PLHfhm87+WOJj
hD7Ken6rVyAVIn5hxdJXNjsAdRuDMNQS1uZuT6/zouTnl1en6f3wXG9DWM5VEb1ca2zgJDUpBurh
rInlwgFyBA4LcdDwal2cRx/+36On6Wdq9Jhk799kWYlrWWRmk8F129JRDDSk598asxWN6pmK6nWZ
OZznTwcJH5GNW9b1peSkEHomBRZ9BZNrfUMroInrok9M5f/DlreWKRJZDst5SxwQFxRJGoXI7S8K
5zHOMD3tPVuQYAl2QWHSfUmpVSd07oYNKZ0xDYwwARTnR51UoSdMYJCf4kQePkdRY4zzhIjZsHRE
cBe1q+uFXqmB3Fhc5ZGST9UFRxUksFbTz/xcPO24+9mbAPTRq0t3itks/ibyS4vI41Shk7NXS1aC
v+Ejo9Qg2fHpupvePyAkcVRLo4v7li+gV4Rfgag4gTVN3Fin1lnXK9tO1CfBUdXBMbiuvAtLkqy+
zyeGzW4ifME1DMJAsnsePEvXxvTdB+rbdFBO09xTptDwGgYmW+5NetzKqQTOInKtJLn4YMKZIp6S
SlplI2LdN3H1oQ25iKXyV6r3HkbpXBbyrWjf8RA5C/lJ2EDJXRcxjsTh+VjlQtu7dbIfU9FzCZ0i
nlJHgqipyNZdqtb36sXM0ooHt+Z4USvUihOJsp0BkQS6zcZ/9NJWsQCI36eY6Cx5XDcMrAaL4jzD
Rbnz4YPVLANjARG6KhTp+3N8h9WL+Ukl9ZGzmqEJzUNgrvJL9OgpafRyPZmqCi8BmlrPdhpZBx5V
YZZFiPC+0U6NvByNUCZQTh4geYtQ+wa8Sc7rNce7QcTHgFugriME2MHSZwsVEsyAVrdRIsRWXkmw
JppFaTVTEL6NeHTh86CT419bo0UDP9ztCbGs0S0KuCFILs1yqkY1j2CP2PBx9KW6ejVig+oiwU7o
cxhA9ZuzvQwqyN+jBJ8l7CEXll+7Bpji9NOTx0Ks9VmTlh/geMy8akYs5SsIUMY0BEjCBLc9PLh3
O6+hh2x8VY4QaO30u1WTf48i1lM4zJR33gPmEOHgu9qo68vrlcKWh8N6FnsHOMkjpHD6C9FG9iVC
W02POK4X4LetuuJzV77hsCHTT1vpphDa1w10xxJFcsB0JrChkhOOJjOTH1pJVHX1DdOF1gB4zy6t
jo5FIR4porsrm737LKChd8IFGO3Du9IEWERmc0z0e148n2+wHKKijXbDTlzs/2ACLxTih8rQW05b
etADQ1R1IlRLE4nEJd4XWuE61kAK13tnt0RXhATq9mOJdU0qk+HGRQrJ4ukE780+bpRt9Z9kZX6D
YzYJ19d/M0NbZKN+AUMNUVqzOAmu7kc8NXQS4fdOtG7oiUGG9YizHiqCFR/iPeUaqbbkwQl7+jmB
5rz9ibRx2yq6SvwMu8fnWwL/aq49s+tr3HTEr4camvWWKBzdUreOZIfx6cIgVbYnG831v+VuEjWU
gOQN3fy0knGl/u9JVi6Gtezxf64g0Ssh8KPKDuOjxuhZ1LSbWEcZZA54H7rdF7F6tZMVOrDZXo7y
YU+KFPCdJkSJwr3Bf9Y7ZEQIkqaipNhRvLZ5VOerONIJEFcdMQ9oMsh0oy0eZtHsHnL/owpY0qZK
Fr9s/oD42axi7XJvH0oolybYBiD31vaYov5JJ4iQK0Gq9/FJVzklXoqBSJWwl2Zc9L2cSJh8zFUT
/Xzm/uhWVNduePTr0vkpz+s62wXh/xjqb8lXozJX/+gbzq3CcjJADZyAoSXXFWdPsECC6lU4OPf1
B+j5pDIBCY1uq4+yIZd2GhM7DkBxDu7bd5lUSDM696yp1rXgiDg7ivl8DdtinTXftip1FpTg3t77
WXTdOx5lX2xLt7UE9eYdJy+1Vt6UXUMsuMA7pekzJZAl1IttiVRPkuousG9Rp5M7FcbActLXRqew
iXFZOj4cQ1u0KxJbjB++MlPOj90jITFVsDFez+CQbq3B1wBBpm7xa+hi+QPKfVKPBrYwV1aRNZmh
LLBjfDu+Y0UAUXXLdVp+KcY3Afhuy3yMNI5954hkFGcXTiyXDzrATWbL5XIlDmb3fizJC24IpbXf
dStlzDR7trfJplhjBV7XwCcJi1s/pEWqS0gK5oLWOxTGl80GM/4QfddrM0HdeMX1vu5IyEb2uF6t
Vua+sVC0t8jAzerdKteNQmtqLJOjO29yAHG9A7Dg7jEdESL9BJCgwNs7R4H4l+1ck9EtgN/e+Jjc
38rrZWqL/M41tP7CQbgn9jsi53Ac1OhuJ1rysot967cRe6W1EjHVCnvLGpGwWRSu4EOGyWhcIEXT
ilTc+T6aILQChi+O7vzkqxTHIZAQB4uVQBlPNmpLNXzCw7394dx7WVnSb1JCUNGf4i44Y7JX0X8x
FW9wTn1Bqq0uXkYNKAzrd1HsEm23Xz5NIIw9hGkUMTn4GV387RS5OTw0fq2Shi3Z9awIURW6wLPi
EKA+iV8/PWumeaJHzsS0vZdw8ZGb1pFGHr1BkMIwpE6q7sVSFT17CJt1tpwA6aYMXE0vLHNZ2J0L
FFzSVuh3wGQ5P9oityX8Dr5q/4XlsYe4n3NoWkYbS5dTeF7vYL7DizZrb2IZu5i8otC9oWNeCL8O
B++iUl7l967chYOAPGgz8G1D/4WbvT3hTP8uLIwNZ1V+Z8qL2Jv76B5Gt2Nc6I0oeL9+6r8QP7Bu
+nBn+agWujuYPJfSQSx9LPFWqHyq+asxPXtqXotAaLxcOLw+dv2NXXY8LfC7TaYvVIW1IFHCoKI9
wA1N/TGUEkk+Sewk0fH8sBatKGFwW1UPQT+qm5rPK5RLqfS6DPb8/Mb8fctJHKGwsjdS+JjQWlSo
AAtVOlhcryjjJ1yqpzpjxpMnsOkq0VlvGbdAwQPXzb1MbIwQ3sHABGFwhGdA9ljJbYKcCkFxKMjW
Vh6hFzyvfbiW4gjNsgrNhj9sPiWd/5FYzcGmDAS3WVUE4r9CUnG0moGFR8Da9uVuKEtasUJth8+2
nBpdEmPF1Hnh3W6DyquI/stZO4lHRluqPIPGA4zM2qKniEwNGF9LIStoykZjANwjRPhtasPejWcC
acQIOHYbgu7yzK01fMmaheEiz6y7CwzU2QIBpWj9woVl8QxZoDQO2gsOCaCxMLQrq0JQ0R/R1Ymt
RZg/CHrI7bK8jVkBQ1j1XOeE2yNhYRj0cEZtnUhysoaShSfRzAlAM5eALNRXgPXHfsBkugyOrQDD
YHx+u+PW059L8Vhay9WW0ZGzCAdw7FA1BCdjhFPkWNCJAsGYUmTtB1MJo+wGfyhTYNv5YEfi+P9w
6iqDTVp458j1+rSdr1qf1mXkMQFnJcnqvazpCxIfomsKiBNUcxMjMiZ2c1Ehah94joUC1LXbpRyq
K27v0JV3Cb0w+TIFFl+PdrUBZM/hFphH2EamYy0lEChc/Y5FGW1j98XdCf5sJ8OC90gPrDagmvli
E5JgSEQAF8wq2I/HLYUOQ1ZwGv+ncb/1ymw9R62b8v7MKOsiW4Y9gkOLkdWBM/5lLpKGVZXknUeV
AxYHGWHqPQkdEKgKEqZgCYo9K4F5EgIeNYXEBwb0xC/ePma01/0NyhkpapC13RcVo3rPoOXSS4JV
zkxgT7Nypad1acCA7rqURWB5RSsohANT6+XyAhs7fts2HZnWU+CECiii/b3M3XAF3xPlw40aTiEW
04jVA3vho0+9RzsFdYuncwALH8JXRNn8oVsJY3AQPNfnkNS+z74tPaft69NtFHtydq+J/JfaPLZi
+VIbg/jhjyLnfQXwImIU7KqsKdZcobVue2lHD1BNwh9j49RkIqDa5Dj/9lOX/Fk3q6lvlOf+exYE
48HE9ikxB7rZkNB+VWym7igXzsGgds6At3ZOw4eNs7J50rXpa5cMxxwop0B2pEgtCDsJWJ48lXEN
zu7UtLyuJR0oyLDKDB+7QW+VpjeZlYE6fXAcdQKZ3eRO+wzHmSevBMS7j/GQoMW3UMdJq6X6BHK8
YNe09a9XNK/uJG2GJwSMj7aSRBH8thqlH4HZZpZckUyMKOIsZhET5HWTMyEaCZOdGB1nc/yTjxae
DaizRwwIDKv5kP/yu0buThiUVu3e01tcozWfVRwXPDuaG8v/Z8zj8BGfWMcFwoYKuN0BuApNtQpe
O/0XjGNIlUeNY902l3JKquy8+mZ4jeVpTdBcExMdDpPa85FKbf/CiYqnE20IWl3W2m0eTNKKzNrv
IlpjWzf+OO0lhARw1SJFWiwEW7uuQIu6CEpHJpiDh6cLnqLZgl+6knlNneejybFd+xqgambS91KS
PKIPU0FdfcUsZU10UjezrAlz59nKS8ncp+QoGiq9CWG5I5OVVFQYpbIiHyQn59Zi5idOHka+HhiA
hQBISszqLatAzSd2BUCRaHvFOYe3R/YXaH8xI6Nmxex9BRSHqaHPIqqkHVTBV6KffVfP4VlyOYs/
49b1B+kDPoYs1dIJMCtjPmRXgRRTUw8e+xx6SjoPYq+MlmwvGE4D2tmeDZxwCSLi5Vi12+St6eOu
k07aj7Bys6Glb/b6fxPKe6bnNLIqdHBaXYUedfsyPG6NFrYqnqmEkAr6ehvQk3faq2x5+gijlECO
IBM0ELlcVj7zvDF6CEL7t/U4qMLa9bbjLZ/EVSUB5OtoE0R8aMh2XcGn+ojahYi45S5VufSHtXml
t+ZbEu+2PZPAgwGw3QL9ZBtStx6s0z6KnqEKSEGqVyfUV2n2n6uwaGZS2TqIBgaGe8p9Wf547qBz
FzDGDnvuimPy0QN2FBTn26kXggXRZ+d++9c8VYaay/RFSTIjvEo/nyVVLJ2YnlzIllbC34FgrWYU
SQ/npJr8w0hjFjR5XJI16ICE+8nQrAxDEjrkCi7bIz9OJixPS6VGp4gDzh59AW6k/dTVIy8kstlw
BCHtlzY4kNBaxYahTO1gZPdVCWXo/IyxiALY6EDC6O0XS77Uz7gKaa5VNFZ1346Re1vfAz/o8iIl
t50YIzU8H9C/fpQjOMIc79+SeDd2XlZEUbmjd87W06FoJzqZlSBtLWPfcs3WZibsy+zp+/vJFyzh
6ilW+LSl3YlBLDpx9Rt38bPtekqIqmtyFXq6KRBpDPM1sUpHH6GIVaFuf+/TS3O6dq2EbVbXGmiG
/r9BjM99ZFCxeDmLmNQEc8wTSGWT8Yx4t/t/J7fFpabiSjtlx8duNIWyd8bFLYZjQP/8M9C5Q530
7cVJWbUUgLPdszwyhPUDx4uqz8ZRFqLaa2poASzfVk9EVRK1PPtn1Nyw8p9xkzmFlSDRTVuy3BuJ
5y4JvgjBbB2BZbNSts0RLc9itpjparoMBuhTxzVb2ZIRnVc7ncStclVOT3Z8lKTLv7UVfB1mHecf
87bMku6Vm86c+hoHEtt+FfVISwo37rLZW3buc9LEe0Rh125/TIEf9IJNUR4t1zhY3XYh+/WbU9C4
SXb3VzxBnJAFS7gea0ERoEZIokFC53RL1pnsm4lIDSkUk75T54tzmumXVDO9qtJVJKFD8mjWeAxJ
iDDqMPk26ApjsL0g8aVOAyLLzQCuqLGXbLKNJMuuYPWWf6MbHVhGcwP3NPNQ8Wa2sYyts9DKiGcI
7gRJK2b+lxYUUOHT9NVourY/naAhnckaUaDSHfkkDPCrlJlyVylO5YT4cG7bjgca9dCV+G2fKP9D
G8rcxtDfAUL+2qWXEI2o//b+D3oJQbAQA9NMgh9ytaaCGDRaE3PAi4z4rj+K4O8rzs2yYvu7gZZ7
8wwwz3+16hSj74siaJ02F9eoPBq4H2x2xiDqcKgvxkrLOLqaJdq9hKBgsglBtNJ/EZcOGJFITOk+
37Hrd4OneUTBpaO9WgfkQqPgLafR+4Y7w/AZpZUGyVuMDEq1Fz/E3bze2tcJ20Ky3iGvdlUllmZg
Cnxi1gUT885G4hZ7ZaDanj8nASnpP0omfTpFkL8DOVR8OC7wcJSdQNo780iVnbbnMvj1IiDkecT1
q2h3suXhmbggiKTPgq4mLCGdXBbVxF/xPHgvmy1Tb1GhHA2+KUVffFm3dcgRreh2qNXQHRC1MX2J
T3xQ5nrC3zb52u2SELlofEQEpAJKwlE/XVXZfFyil5mLPRRMPQLk26rzQqqfCr9eG1A5K+dB9vLN
HuzyoiyqRGYaRX9iwmBghwnLbFQO1fP3Vn+bNLXv5EbrdzOlGI3dlaMuwtk3dOsDSu2hQ84uuM66
fc+NKjlRNaBoYk/rjmJS/TU9BzPcG/n+GrxXsIbu6FUwcglg8Q0Xcx60dxfrx4ZEKavDCVKF6sdT
hyUI0IESWfLwg5HMIpQe7i9B5Ihwp5aI8jQFeM6yCg8TzSIZZwjlDpsDefSxujQnyTwNez9MCYUq
K77hJeUMs7JeklaUxNTjIW2lStp7BlJR3BoC84XUNO92S9MvunxfoGiaMtC7MGCMRq5eDEIUBW7h
69oeHIukZn+huM5MWKPA9jHvbqfYQMBU06+h1i+xEcqvi2ZlqnStTNkwMmsGfKYUhkbXegZ/G+Ty
y8M+2+1OH2H5HL0UsnYnfWTroggAAsDrga7iKdON11BAkPe5huP2DLq3P1SQ3zran0N5T1JqqIIw
gXPhuCC14VZMACIsaYrOnQpu/4gwuzg5q/6knZM0Cr90mG0C499u8Fdj2gnrva++v42szz7MGb/T
ynK5PFcCqfpKMTjFWfbuaXG7drZhVaYrTIGKIkLG2E/zBauCW/P2zTqrqW0de4f1xgK5NaAa3Ro3
rbSTw6U6by1diqkjgokkgi/t4gICN09kOsUjCTUgiJfT5WUw9PoionGaSue41OoVwOAHYiuynLfZ
SPtFmu2bELz6h21LClvtdyc2M80NKeY59YbFru+eSk9gpKNA9XK31TzMeK8pv136C5B87I6kbLni
HAJDfsuC8St0gL+5HYl9pF9Czfv5XghpqHuFetL9yg9N1NghvTBb3jCCwEZQ9SvxNMpBZPHaAk78
NSWAoaau+Kkg9bOGzHasBb6sRWZTyYRoi3rEZWI+/tFWqNR80oAHX/RYpAr4Zwxk3+JyG95o0jkY
MwSXlusyQZNKHcEejMATqEB90sIUh71QGn7C4jJtlRRY2EkSgBS6exR+3FuLbdqdmH2YJm+yv8vK
h88wYJW+2V9FwVdZZhSQyEefUPQfSMs+/sQ6OJA2L+C1hx32tYAj7Jg1r3bemP/umtFcpNNrUEUV
tVN+pdaY9AA+RHULYUPwOQhO1egP9MKlnR+0kO2cQwvb18r8wHsBbnTNLwcnbLQsdSSB3ICaamE4
r9kpQjszWABOzsWjtCGiR+4jbkBr5xTM4FQwQUHSdBWRx/T61WpUtcI2c4zJSvEoYATaqY66ZXRm
kJs7w0fGratHfkNoUI50nNEgq7M34qAtbcE2X/RoQ/BKvHnluzT5AIIk5VZosvGoX3hfDZWMgHWT
nltGzAy8INp30MmgWRIi43SRzUAhAer9OlmIFfgSbWVujJr+8mMaMFyFVm1y6MxsMr+JD2EVfSPA
WAMzVjhieZ0sZ3iLZ4Uf6kQ+ZpJrB2WvyZ3MWP9244rkwg90okd690Jx8R1SLe2xXZ0QnU3C37F5
lYoPI0BZrwPDVdnxqKsfk+ToiLx2l3Mv83AjlKavmvdd4nfR/umq97L7MdJp2674BWFqD3JXvtj3
8wlcgdk55hqyGDB3zc6n6xHLh+QmN3kIjuUw1E3fgkrTSLE1iZkANNdtgMCTMO6E/OFNDTpVo3X0
wUvmlb92F+CpNkkmq9qulRCTIPjY4rU8AdeHltUoDzVJ4A/hvuUHTWuAQpft8WPpDMrZ7ni+o78B
80LA6gWfaW4SHxmr+d1zp9drPOmW30NT9K5cIt1XmCdyRTyJsAu3rYEdBMTJy/HKCSTOEmdaw1qY
J54xjn9UwF3Q6WhD52zU6f9bO54amz4sWAiKUtWNm6OOZw4a/UzkfqVSW7rEvYiM+z6bw8SlklUy
VJ7W9Xg4e/v4mBbH9rIzfx5YUiBcT0UC3/e9AM+g5zrQBBC5o/a7Ck3xLKSYPw8lYcP4oh/IKRGG
CblHQ8r5QknBGG7EqJ/2h8Iqjm9I3Q41XkLL1HMbAMRrhxXSjl7CZxd4ShoiMMeVxIVyuQFOA7BP
D/raj2xm2McRmubquOek1pieop8wm0bzHuIpHSJBMaYCxYyOTZNxJQErm5uTK1f5YwxJsA1PgKkq
rGg7e2BWI+45CqUrvU9YtpdD2sSpMHlk4tdOuXLZBxCvXxTThH0P6Y8eh6vkEW8Tu6D1hNODLPRU
3gUYb71lgdSL0PkQM9eQBCiPFB/UOn2Bh9m5EdLtipNuNfpjt2vGdHAYmtZD2wI+bGGZ8ttuxc71
hljgNGrO32AtLz1uHIbMTNbA/dK9LzGTpn4c9ikLklLD6JPhW3207numvxM81xCCRHBVmNq55BAd
6Xy6lppku+nsHc6t3L0ixBGOTsG6wx72S6pLqOAiqbvPMw89iD1ODGQ2BaVxcoMzHRtymlBLt2Ru
v0icPJNWpsMLwVo77Qf39XB8ILKiBMhb1wlVpx1D5tNvAD730zsrRRzML5gzXKnIVUVmDbmMlVv1
3HsfnJkS0MmaIKsRE4ZBVX7UgQRleoU9DDE9jgGpTj6qYv7A2x8RY4Pyp/nAEsTKJQBq7lHffXtQ
AegycbX+5aL6sctdQsK0/33SDdp/tsSAP5e/+xPg0MCYchC9LDFKdzd5Gcy+VwzKt34/f/f5KgiN
7oqreOl8o24oQ0Eg2JzBJJ7lECz9RuAB9Ymr8WtY8ZBAYe3XJM8cBfHpSw8wTQTOsBus8E+LOb2q
aTSVHzClY74iX8ma+ksOCjeeGSxq+m0UJ5zNC3mdXmoxr3ring4u4PG+lIhQNKugIgrvYzl9BhSK
qyxOUFm3zIs3OiltIHh5bWzfdFJEus9fXpisr/EXJC8muwfHtLOf+RTDRBwDJvZNWcQsI3xEDWzf
nD14YjmIYBE6yCwTUZcmcmkA0SkiARsZgevt2pjTxiJJR81RSieWBovwh+4lCXpAnqIqh/Yg7oPK
NJAVe5h2yKSphxxmdOwxR2dd898Y1r505PUdFbQaaUkJ4VUDeUsaV+NYNAiRCif9UfSjHcuaGbxq
nJoCR6zAZkDO59hOrhi99Qz4g9lRa1qPOyz3GcdjmSqMiCGFQv7sGJisdjNk5zU7dEBVyK+hfbah
87o6QwBhcZLOajipPzp3sKjZd23PczVjTo24RrcIGp7uyA8g7cOa5dUu9mV5fqDMoZvPDgKrutP/
f4cnKG7G9w1+p+dn3doKYtpbK4mw7mTWIH9Ar2r8Hq/3pawTOPhG/BIT/8xnaj73hXKc7nyeEUwq
dPzhP5w7zMOWQQKuqiAY47Xr1X6XnEvH5s6Jl7Z3Ah0w3h1x8VDN6OQ1BgZeGD0o6SO+wghn5bYU
j7PuF4PIkLKL03eDgJgGNkrxByTGBnsVyotjhA/fQdXqxvgqznFb70KA4hXBenNCNZM4sT/Kwl/N
1ET/Vf32dtJlWOpo3Q1AccCvAryVRai+mLZfjFxJUfZmzINSS50Ysm42zLvVVHrfwXv0bq/7bqCp
HoCIy+zx/0iZlBHd/qcFYS15egHjz7tO57hgBwozbjx5qgDsdun7P3yDBrvArv8Yr0I96uJBGQIA
TEry5gqix3EDBxrb/Y+tcxyuYsV5okkmpHCWRlKyUm/8dsmw9qoMHY5CS3pHvOqyOKovqYtyo7Wm
xy89ubCeD3aA5acza5U9+KXLPL/PSuYCbaZRWOt/gL7+adivIsanaedYfrN5crqkQOAZQqZh6NYO
x9p7+hl3UmRPhLaHyv7LsNb5I3db5Oq8mjPsug8CsD7w2FUcwhVe9P3h7bltdDze+08qyKB3ASkS
2xVp+Br5tR1/kftWeJ76GbLdM4O8sc/UP+wnhdEG6DUUhbZjmgjQ+MtwN7hyhmbDc50Y/5DzR3Vb
qGGZGI3v5Bi2hR9t8nZxlqrDZzakl7QYOVtSGjxcni1/usptYckXFHAPqKE55IoptYdMMJeMqik7
fylW9oUkLOfNU6OvZz/lOAZULI4eif8rdFDWa+tOxtOWkIvDhOFGePJn6YTmqQ+4RWkSpV52wzF0
b7imyenfZ7awY3YdwDr7UxnOOL4pksa1DKjQPxiXnKZ8gsAvkV6quTwO0rGTkH5WUYpFx0RrGGzj
ARQkMlAD/zRgnPcriOaenlygLFVsiRZW7wI2dV9WhqAHnt+T+V4mN7WKyy/mP+2h2h9KagoOT4qF
jmk0e4khP7pqP5L2L4KP2YAVhFK6HYAPPFv/AaS05rYVP9QY4fSWQIoUrXNowdqxI6x/617StIBz
BcG+jv8xfgIer2z9EYRjEW/ZqD51mTilR4GL3DHQSVMev65YdgY2U8P4oaEAzULY9R/yLQLatu+I
zsLJWWblo5LyDXk6DAr9GHpl26YllfEygYXUarUfQyd6Z6XU4nFAh/yIrKcVsgI5vRc4G1GMlod6
LOVffSlsMUD9V9ddbpjm2E0GIpsiqodqsHXLSCOX5Tr5joJjIjFFWubwVx7ovAwuZuAHnMCNGRsq
FRTcYns8Ijj5SMe+IggVWvpH8ypVj7sSHTC3OKERCS8lR4q9dV1jzaKBUn2tZ52Vf1sjkfggRvYG
Zh592J1xbcjhRmKiHc+vzBVsMU9umqw3fU38BK41utJpTAlL0hrFoabHVknNAJSV1xyXpZqBQjaE
eAkASK+xIVxLPbp5GFywxYw/S2pIIdBvJ/tbskjONVlwc5PRuyiewSZrJ8V6bcQwITMvoHv3qVzv
Xpn9KsFgYTM//cfl5e/teDLQ+bGoeepnf0SX2WOjFIvV7A4ldfCblNlF2QgjtDfWSYxrNjt2TBwp
UU5S23hE1C9Li5bdec7WIsnXo5Enyo2zl7eHzKGgdzRCd+zZ+St+mJmpOzIvGHEJwBx4imrOYE5k
sCnhU9KBAhZdYy5SWs/AqipU21mniztlTTwHskdKGnq4RNWfyV97Re9KrjfySqxdu6uSlV9mdxyE
/1ofB++69rENfCw+wkSg89YAml6uN1kySZl1GGFgE17hh5mmo/dcGBcYFYtM0RHnefZBCaaMZoGA
oHL4vPWxGdc2cyYTTEGOhfzGaP1v44f8atw0k5PliDGwzOZjCOX76BDmmkVtj/bE2wE/wzMIO6sZ
CBU+aal+bf/0HmURz32WLUMfYm8t73hSDwHxgbbqZa/8ByLIvYDt/6MP58t9Bfrl1dODkXJjc96P
z2rCcyPoyRtDO7eaZlx9YYTMB1oAMWAK/sJ2Nhz1FDOZBo/atYz3rr1QrcXqjxnSu/mIPu0Hny8n
nPPAoraiGDoa8MQGL52nuFR84U6qmaTdoN39hMajhQ5HnXvhaDWrMJVQo2hINPzTJX2tJvvHrW69
6pNFSmSbl7vfTPG0YfyUsbWVUGWWWPN5V57/+eQlRD0WvVzywoIvfQsM008uk7QGn9ykAuI9IoGd
CmlfClyXA51lL9DWnAFXnKFr6kyYI7PgRRhIUfyOgmd4JCllbecvloESvtci5ugrPcHoZligrF5E
SX7v7SHW+6nXliii+0So9heD3x1XC/NGGI/F4S4bAw0AGCmPo1tE0jIUl4dYIxEIyshe2RNUCxea
oGJBAStq3me59v4IEyUVUD+LiwxFmIwjvSwYs+j5mMeKiJHmhdCyplLeKHSXhSCzTZfMm0gx2I6S
H7VqFCjzin6a/YaTq3a1YscCSmA+07V8mgyoqC6PP3g5T/L7gs1rQEpP3XxMHaLF5hLnAfu3Lbf6
a5c5oAVru4CHrJ9CWJmKwTtBwV+YGdITEVj/sDMFuxYEYbBROriScWGo1iHtfyls5Qqo94RuDdFk
Ap6h8oHGDWSat/WfSyv1f+S1q9FGKBbFBvR3r+EEVKCzyPdp6iFPJCU5ReGOQCYPLjT/1s4uUp7i
amMJdAT2bDIYZd3m4yJEeIw6miV66sLpH5A4I/bZ4QNKFC3gAx7kFAuRewrBXtZ+41x8auvmezwd
+sK2PXmrQKrtn7mdYrFBWXkv0JSQ+YtaHgAIPC3ADJ/RwexBebtuw0NekPm49AmQClUtd5/n+lrv
Ro33NPvxuDnyTUb2Vv6zTdF5f/Quyt8+PEe5FtQvQYkFtAuTJgyrzlG6Bd9vRg9ZfkTYNbX2TwH+
F09U5rSdgZ6yesiuNaqoJjLsSMgbzudkyCx8CtT4Pp9aoLqPU80tVLVckBt08yCVxuPM/ormga9r
3SN8MPcIxjew9QbDK2g6DJjlsVLev9Zyr07v+RYfBicLBCHl0HxqyDaSMNH5/pKCK79Uul7wk5SX
+wR9s8Yh2tlwlSn2thg6swZpp1o8Yl074O27ZB4XCQPQJ40ZxTYrFzl2IH2WFaNBcxr6xt+ZJn4f
+KjO8WlLIfBQl/L/KZE0laRBAHqZHueDagEBbLe2AcEc8CIqkp8qw8OJW995gJ28IQ9nR2beVODJ
HeBEfrfqJ+DmyCPf7KE9SykVqxgQFnS8qMsV3P8mP+uAaGCBhfJE4DMcgC9B7WQRFRA1nskNoUgq
cyIRghr05R8Mms3I0zrpB0ypJdmh3HP8400eA9x9BCJm+kWDGXiOUK+DXyUPypMxax2hAMBIUSzm
arnGqBKIkVcS0sYu5PUrp/C43o4bPpTuWnA8uRW0tlrDThrY2go0LHIQj5kuUD/kzRRQbB49PZ7V
yiOLSVb3qBSguXP6VfRboUpw7hnVIkhE5oRe9MfNguaCZR7+1w4hLRszTUZXVotjT0CUmMLXtRKP
NoxaGfgLFA85sOgpwJapt5G8t2dC9FsVezez8QmNYXe/pXzVchbPxNwff/cSrj9HQJodyCIRPTkZ
10Kg0G85Teh4GEpe5XhEBSD0+3W2UK0sIKeKxvb5seVYqaLMtHll71u7HjHfJb7lG7JtFU2v1c+T
FP1bS7y3M7/I0ul36v2ovvxygc0X8vZec3asF1yemrRleH7eCH7gFOjW96wIoNlVxxV2765c7xDV
7gZ3GBlx/wPYrVsUBWFvpwLd1q9xbHD0vgueqz/XW6yvHwDT10MAf32EFU1MI5uza7+YrZS3pj1/
3AkQmFgp4m88DFBwjGGmJYaBskQlRu1vivwgeXTvZ58DM8AizlzKJDLcvaI3RLm3nDtRJ/1LOSDy
SNY/w2/7LRTNrLVgbseC3M/HEOOeRKXuhPfxQlneP/z2notWKlTW/ifmsnTZKsbjaYgwqs0VDbuB
HjGABdvyZ9nswqMeu96rgMw5lv33WST9HFBdEgf7yRVy6c0rK7k/+Wj8qA9ofd9KqSuXRsjfP6bn
sc4KLagr/zbK6oI/LarueKk7/MFdxV4JlPLVfmE/D0IVhoaIRJEv8Yd9hHHxmm3lrnqrAgob+ijI
oAC2X5XSFyfpzcn7an3SYSIuODaX9rD3s94Ths/3rAFvbgy3LjJTrCd6gCZfN0vaOHiU3t0C2pa+
4/BQ5X+158TP81D7pV2E1mJIlGIEY73Yz3dToRdYAO2G6MoXQZJmUs+nOKG7ABySAF21gBGNMTFd
KvGD5iqJiW9gZDghBYLtGo97zjocY6SPf+iKuFTmPP8jJ91C6J2A3dR1aDPqTmZHrCAqIjUx5UPC
iTG0UaCvz67X+YGxvSvhwLTeIeECK0RxK3/FUu0d3hDaBdOttOJKpDqhTeEm/9bhTQBetcGDzA0F
dQvIjMEDEvvF6US+fzomWYLx8f1WYckwa2uqRzqtknzTd1v1NhcmJiwdzWuafM3nFOtvpPHBi3d/
w+YjIvWnUly7mOetAx9GozixE5/3MSbqMtmgsmFImwgyUhD/kIB+BDka8rwq8dXuSRCHBsrw0ls5
26W4BmulIz/uZoAjlUp/7evjm+HZhT1XgI/YfmKUS89RMNbvXzb/Cky67hA/b3tD8ojTHj0OJkPm
L30yOHRMqsMR23QGrUMIszuq0SEucEWNpzypixAIrv4czPX9QJDOacpRnrITr5C6tuXCsNEXLQCG
+vJ98wnOXJw+I4KaHAKnDQaaOyUob3amBGVkeL50zfPQyFagnaPfwbQEE5UGn60bGGe60R79S2fK
XZ4B7AO9/ciwfYPqGAkMPBVZ/SrwMWOPvG+AvyMCG2IIRXLnvq2KjaO7xWZO4Y0BQzX8souyq3YK
XvI2b7qBFk9Q5c4TzP7jXGjlOjmBd39DsbR3ZatdJRsQWFVtJ+2XSMSKsyeQl6wA6wR6g5AiolQd
eKyp0PxiDFet9gp6pCgmWtxmshCJ2hE/6Qj2pwSMj7kKEFp89bvgrxzTdf3oVQn2uzIXxxYkfL4Y
g4uqp+XQ6Eberfw7FcGuAslaYHUOXgEHbdkayIZQID3hpljSv7tNa8y57m7sMxkPQoY5KN+KVXbI
XIgSLAkz5ESF42bDoI7oweZ4nHWGquz/xXc+Jnse/ImRYMcjWzjvPlEYN3cA+M8HnojDzMpVEisR
9GcWtdQReffVQ36VvuxFBcyEeKRPgAcGogoSbrjJIr1+Hs69PQavH1OJRb8uuEMzwsnR0osHMG7m
Zm6rK2ZPRonVPHgzCYEGiyqEtV1y9mgx1o0shePBShGeBnoUMHetJghNLTKf0ErhsAr6n/acRril
iRYTe3VOFgH9SyCpskxYz1TXsSY5v5481GD7W3W6jOzgavSL2NxXrFKogqulIQHuxoiwu7q/GSQj
+T2liJLOYs/Nj9olDCTVoKflG4vznEBP0DwfpcC7/tobN+uIDnx8HDYfDbbCsN1eF78hyJuWWNBs
yp2YTpIobJTqdtmjvb1VWY0Cotp81XqPBCXu4rOV6/ixcZh9Kpxad91gTyS22x3oCBZ3n55xp+An
pROOMt5AgPpSAi4j7HhPwA7GfmfuNjpep6Pdqn46qThTUA5zHGe6rbYjFk6p2fjs/YL1Xo1jauCF
alXFBtxGyPdcrmKZ/NkUl1yLgV6tVRcVUoZdimgem67npz7pBQsgBlHv3YlgkpUxojJc+Bw3QHD7
iL+QX140WMywErihvqXlZD3DecwDFX0htvVJ4wxsd6gi8kP7ydInjD+Xb6w72LSTAZUfaP1nUbzd
8KoXn7qgFV3Tg59NQNO4/PyLwXgGzroYNDz8Bk0mCpJJYDEZDnj4+Bp5IZDEjZzlTEW5qtlJqbD7
0/ALyInDynDfFfxV/48Slvmr2STKM6lcgJZAnSAItySQmxhwcvcaGU5AT2qcbAbHKqdaKthTjUwv
mD5OH5tOkyuolPN4RLifjqs80ke47ZWGtU6k5ZzZitydHd1x1rTF6ybCf4vSULnChYSxKmHl4gwr
95Kvlz0lTPxAm0ZttmTAhwvw8DyF7FkiBO4BbFVFZmrJI6+OZNYmNe9o8uIKywUHjOkT4i6l8zWF
fzrBFZZqntrAEKoNYuMSqETcpuU6sLdSjn4p+A8TtevbDzhLTlltqZ3e+w1TBkeJyVqvyWnauC7N
TpbFnZ5fA62J20HahCykqRjd81biubb/LA6lcI3A9gNgl5N+3cK8p71ba0rIXHj2CQ7mW3g7DfQa
HVe2UvmJDmWPpLzmAaDfQ992qeDCd4BygyTzOCoh45+4NPftB5pQbxDSHhwzHjg2pc83ud6DK7b0
/HB6jZlywEjZiP/F0h8hv1gJ7a4mrN3B01mMLmsuV6c0SmzCWlbrs6xyz4cm33fzZrn5fJjp9I+e
qDJduX+qQw+UCR24is0BgPSQFGsMBNnZUjlTIqj07Fze/P/MATv16cFLXVUafOImlHUPygETCSBp
t8i/7Q1dUsxoM594bcWqB4d87L2Bszsz+6PXzcDAnQdnux6wwVUa1Vw45flslRnC0zCVqy06LtXq
26Q8Mn94dF1Oqv99PrRiyk6wEvuxg3KSEslUxoWW6MpmpnyiEiK/3kChxmXc0QboJFzcjDPu7LYV
XY8TrzTfeGD3mCOY+5A2MUqf7vkHfb2pwLY/hKRGEmleCF2sDdKn/zyvv1C30vGbCK9k5G/ZoywG
6yjnEyCLEMUIDZ8Jjw75EW7DU+QSBKixz2E1ZsfbJjRqpLLVXacv4zHnutoMnG32vbLG+JtBgV38
CYjrXd/a6JHUlRs+E/uDEAYEb8LweOtSUtXf/q2OYfY2fNJfuLkBg5nC3Qb4gT1npe1XBvSW6CG+
K7135ajmZ87tuVLGe5CvV0ZqLnjWqFSrAHvasV2TRhrMbANxr298p3x5yt4HSS2Yabijw8/gVD7k
FeXog2Tc3ybHtF3CwDCNIeOCQCRWoT3Pzi1AW0TS5yp0mvENP9rfl7bFiHvyNf2gkbvOTDy+TwaZ
VT0MiNGkVBZatYObDlj/sDKfDVVKeuyrS8FdhdgA51SCcDLJwMNvhEpJM8DZYe+4AnnxKTCR/bZN
wzMfxFP6T5Kwq35vntpDdkd2yVYPaL23SwNusbHCMwJ6hGvYcZ7uXR/XjdoLjSd2S5voBqmj1Msz
lxdwslbl6aeYylDP14aCzeE1anK0d7qHpGdC9X7C//Q8EttkpsAuNUbj8wPCKGeGrV5qn3uQmbk3
o3FDm2idXoISa3w1qOWebCy99AmD+oWoeW8ZEeyW/qt3OIlqukhSBkYXjVs9BGmTjiwn1IYC67wq
TB6C0ZNBdgujklw8FzYjGX1dxm4sZZYNMhTsQdUQXPAD0JLM+OtqZyusL2HEpaeOzEGclVrjASy2
+uC5ZiK8utxXuxl45S5hy+WYdgXbO0SIdbWPN5APkpn0desYszHQKfi1hdSpznaKMJXTXr28NXLn
qOVFPhqHoduXG++IUcNg+6+4k2qFjP9R7hMn+TB0O7w91lhcIkBY0Xgvloci7XiqM/DwdayZGimP
awDeyjqyUnckc3Iet+SQfaCsUU9c5WWqSFfunvWL2Kyw8J7IB8qVJMvtARkizAE3oZcQuzkOcnfL
+xfK/a+olfKWqMPtaVVMcXpTCpSYS4EyxGbV9OlkMQ5xe1HmbsBu87KLWS9eXs/IIyBpvlb9U+d9
Dt4fjymX93mPCJZzBqgPCbjMHlgjgKRZMpyxi8jtc7K5xuLqlKg2+G893ElGC6gg1dmxU6a39995
KPfu1RCwhzek6lq5h30sdG0q6qiaUAkSG4AkB3oDr65cAmZNHJT1Tks3Xt5G9VugsYkWlFLoMxOv
6uZlxQsrabwanyprzt2lWFDkrXNmXv9w2D7kX6E0CFbpwK718UfhFNTEwPagbV2u2GySghu76o35
Ykx75VDSM92tloGZ63CqugOWhcfnznHTtQC77/GftmvTSArZZmOMBZg9k1K7v596RIkvtsVusqUc
9Snt4z3Ci41tdY97cpNA1FRwjF0kACFJVAmqN++ROC2v8PNTsbZL6xaqtJCqh6LpsIXHmeitXxZm
/mdR8CvyPFhkuK872YcdGkzKH4f6qayT99dwmFkonKzCgDZaVmOc5s4MwmZ3zuLHQvq0u0Tcoktz
teMZQuEdM/z/4VFMTDWeR+gEmTWQn6+1GexXdDlYbHPFDq/ST1YF+77MvyimrhKKmhinRP3i2qAR
7WDxZnJ3TDPRAhkD3jZa3Z9ypi9QDAAqLLfYMuDC3NY5gWjR/XGV2WhHTb1KfRLI2XusYXO+6DoD
ki39UjQzjp2rtVqkCYgdd9tna43YXbSjiGA5RVyAhabDQOaE1Lb/Dg58ITPKK2QoFeWFCEdfxysC
TiPwEu131BBvWlP9uLI6iNMnNRzF6vCatfq4BNoGVS+pACihyYwBdxhRCCNnu1ai5lZ1eGCgzJUC
5nAfo9LBI27nG1Vf3YWW58zV34/lOpjj0dJxiqiqF2UT3hKKqjChfSlMXnnzg7gyuDfeSQvDTHdJ
6UdaQ7jKTnmp9kohKjvmkwkkKPlQ40m2kvnxc4q+LtIdPGtsN4mTENMoaYW0QXkOLPILpnMFg/GG
qHeYJ0udx+zNHApCStJFF789pW/n+ujjYoiujzQHEUe7ZUUMYFGG4392Rfa5o37MzYQxr4NBPYTX
REz4VP5cV6VdaOdf9432Fn+Q3mGAkdltKwStZ9Xvh/OPfjrrVCb9Idsr7xkVt50PkdIx/Zb8L1d3
pq8kGPJRjl43dtB3CdrwKeKcioyFdbj0yClSGG85i+olTKus+lE9Ano340Yz+iqRSx6x4xnpWxTK
X8ThQOniRrkAVjJpv1MEet6UQ2mB+WLcxfmnjZtoVDelhHsZIJE/jSewNn7J7TJ4STeeTWbrCF62
UxPGRe+fZxhjkCXCWj+XYzS2SS8kkwOzTK7AhcgZMy53Czibej0cdRwbVhWVbtf8SZQ1rUxeRq97
kDRbuidH98NV8J/97QmSuN+VA45BwEg4AJmoWzGnM8Gg1aVgH7PrPudM2SCxuWcldQkD0A0dahrc
rTkU35LqZPiW8Yk2jsMoL4DphckH9AxO8mN2V54QuklBHD9j0n5L6nq4cRWrk3mhlZSOB8mBoBoL
ujDC0ffDC2Lr3inwnpqhykP9og3AQnPBfSZYbSeEQSisCPm87FUXvrnqLV27EPcjJ5G4mT1yVcrA
gt+E+5vqEQaIzw1abFsO6VEuEoM+JIZLCUSjgBCCe0mGIzI24fxlFxR5rah3YPti6TClLTq4+mWW
li/nRlynqpBUPydXNzpgZx2vQgk+Gwbz8bvDYycZvRmd/ztisbbAk+psTPlKK7ViVANyyOSSSEN1
L4ktVuKwMoJ1t/PIqmecgYPYijzlI9n4BnB3ViSt4GZMyNbuzIBf4hlI7Q8fb1lHJVpttS2bMjr8
22N7jxKQX9dE61m1Li1ZqkgOm7oJ6qYh/c/clYmgkPYAMLBp0jdTytwOhkhM5lg/T0Iz1NADqaft
iGJbki+AhBgolhb+ae2yixTbWgUeqQWidtK5m3Xs6gXUcw5B8uKhNyfxbbWjAVAyU1S85JdiqEIN
fq2nz9dlElus5crvqTeZBZDJhC7/xwbKQVxz3Z8qf33oYwaNlchqOgOQlN/HAs8Ncjm8/cREba1/
7tg/Ekv6eK1AQxBwKDmSWsI6cV15BKnluVvjXPi0/uZu643PkGWnf8WkM/qIFGw2n40NsiaFVB0l
1GzyNbaYFOMSspvZLvPiPumJzfzmzYhwOcQKB3LjoLqs3p2YgUgzJ8qkV2/HmgPvSjS8bE0iaihD
tSyrU8xGziHVr02Rc6wkF+Xx+IUxdpD/qrbeMeWAdzFKwpBx1ZCzhBOm36/ouU5j/QXegOCt7MrF
jY9WMicTJk58B+9dTsKTpZ/kmjP2Efk2/yJ5tVCrAkBpPA3UxXZ04n2D7qdihRbUhMcEfCafPIyB
e5/SMu09qIi5DH1Vnh4uR/ctcM2Pcb0NRANN0ckgnaOaL9enQMbqOxOpTsTHwtzIVTuHMhPxNpBJ
lP7oYesx5Uu3weMvzxFWsO1ZHFxiNVFPSxnLWoarBqrrJ0WncoJ7E+c36Q4cr+/sSiJ/8iND/r2l
vtxgsR99H4i3npxPI3bHaXPBj10yPoHsUheI2ujqR0VrWi7bWV/nSQngrqS6dC2LZ1qV/30DvZYn
FM0jijbtEFRX63Y+FlKG4hxVPuTaBImb90pXOmnoJFXpvECaWsgr8hkcStLd33u7rJ+/0x/3j1am
cPxwzJD9pPrXtgb+Nkmi10vn/B89M3MVvMAAfamN4gf72RwZpMCOODk/zpARIKjuxVD+pFs+3kXP
TDMHQWlfdTzf8p9FRMr6wgmw65hFSyO0rpc8qWX/ZhhJACEQJAQ+B/2z0eGuCtxpf0fpZhXUC+oY
IJjmw3rzz+KA+r2jOi6tjTLVnoLLvAeSS3imfwfmhXcyYxXnkcouLGtH36t4jUw20tKow54GYJC9
j3Y5m59rvQkdZj1UWIq3EqNK182iS6AuDBwZoAKSZqNjJW4Tcp/LvVX7toOvhe6VHMslorimMUIj
rsIoXVEnexGnMLkMlW6bT/pPObOlRzcl9dj7uDYNU0HVPubLi7Pcx4/x3rD6jK3P5e0cjw+PwqW6
nykESi+TawSIqldkYzCxComRpjCvpcYt1oyP55M3z5sxuS93hAhzDoOM2VJJKdGPzyTFn8FXNytE
kf2ybkBQWU8t9uIpQJ8+sllqDu+Nr6vpZcVimzprimmyC9uLQROUE293YQ9E7S83L7cczcUa9MVE
vZOs269GmypjC25iibzhqccqo76fBIvzOqAYRqzjFJ/vw8U6JEhslexq2B6Tt6ksMwVlzxQ40v4m
SzitMuOUPfe+x/0qgWnDnCe8x09UgRhlBydSkrNIO32qr3tllR3sJSJSvbeprNW9jphmJC4mpM8Z
CUjJD3XQ6I7F+qIwIv2VHmX3T8wGFIXbBAO83hK7NQ4oBigmn5rPXuw7xmSfNAAsskPYDSnc6c4N
EOrTis8H0A4EtPhcm1/y6eyZ8h3+cQtqpFtdxiq1/iPMEtVOt5iz4uDwficl9zaN8mfX0dLD7+AB
/0Laf9JUNhRs/YAO4o8Fo7IDSGWHtUvzdRXVcA4TPspnYujhmgs3imAmdR5Q1CoUzFss1NfKzTPt
T4TdMQqQbuCDkCbKq6Go1u9Oq2Tgt6NRPLPXOIhF188mH0g0FXSlls2jfyPCqC1rIlQneGXmWcu5
8AqT/XHGd7mInamOlwb40L+MX7DQzSUh5UAMknM/IgUAajEMc5iYZMmMA9pWlChYuEJw3jkMOT0A
+Fn8mqGvysLigOBnxpOdIbWQU+LyPtfwq9Gnw8FqaRz5qiAGqDCXmpl5cGC+ClSbA2dY5tArCptD
nOwymzopcLuVw/Y6BqV11tg/RDxu9fIVQsjeIokoGK/+xGb7dlBDv19lZATn8jsZNAteP5bNCWGv
++QpzmZcstgzokcU7cs9C13TT2MXAgEZzX9FbM62jE66LZ1a+8zlRXABREnYn+JSzwpLwTaff5bc
VkWT4guvFV9+xra6iq72OSfvJAEqmgQDnBOdqMK61vH1wHOHTHx5+uPV3SZma8gla1XKGorxSPHx
E+kLdEw9yxdzvI7nkc1XvV9G0//FiwTxwyzk+tji5myeJiqjD0C1KlKg4rFTrdpHvHpFmPXyuVlW
ai/Cw/c+2rMQazs6F12SKtFzD1WFmRKCAUWFaQHHLCUa9E5GRz7kersFnymD/ikd3Qcgy4hj7urU
h+CMdaAF4Su7AVc6i2xkB3XRVRnoDEsbmkT1WlwVeSpPRYvsvOBSYCAUnkm8MttcMFyewRKOdF9e
pZaEwVGF8xCruKG7RhMWwejPGtH7Fzqhv++QChnoHQqW0cJ+3JtznSDVdSlKogUQJOD+IZF8hzZq
Dhg1+iYuUSiJrGgTajaDAaEvIsWUQHRArqjixqPnoPXGh3KaZ8zWwPxH6zAWLP3B6wRZTqyCSVNG
BK87DWOJUqtM1Xx4F3rNNQpVTiJkBmt/mNQZ+gAXcl4THHnK+yfG6VSpF1VDgRmTLfxoPbzHPxJZ
c0o+fPzxTtxY4cid4x7pnwaNKyNDmzBWFPJQRuoNKBSt3fdeGJnCUrf5j1ba/b9bICRRNvdkm9ae
1MHD+w+8bWmVmrLxrTiNl53L06GEIlukC+2st/NBlSQvu4IOT8wEQeeR7M5Tw3T+UMotvQy1YS55
tDhQBKY3qMZK2muwFtmNtgRJciHk59jYO1VmphibuwHCuNVlGzP6g3Fv3EoGCUnr4F8jKDrkR1s/
Gl4HBNuobGW8aylPYMil5eu7T73zCJlV017O8Dy+W3qyTkhE/69zciZ1OV+qvqmGBRqEV9gJu0e1
ea5tF+4TMa+1zolB4vNko4YHqyGMissf69Z+ZdK8hT28BfDnrYc7UJF153amK25uII+F0LmE3hj1
ylb77Hq5uk2Hdwf8Nrz96dD2s4TrB/UFK77WYIUs121ry2col5e+ND0l9W8WEB43JoZELu0eaSrS
Sc86uQixUNBSMqEAcGBmQqG+zqRgijM0Ngb6do26k/bS8huoa/hqXjfhFPQZHe3grGud2vqO4UN9
WVILjmSVTSRETUtx+nsRqBH5l0PW8XdN7Yih9v9H4zKO/LN8KFXq8Lxj8iu5M8JLME26vrVU3TBZ
aCVT5PzfLsfnj2fz1ggXRcgGuLh94XXeoQ3ns9Yh57c4F51J4+ZVqLwHc/krZWjmx/NdVbbiRNUE
FLkgipVD0eTsqhhiGmh0yLlbtZMmu7dAnxhDZN+pRKjap4ztVnrkXmOlN0M5OEvj3HEbSmwfN7NN
3rN1F2dKLAP/mGnyugx/i0JSO8NtH07BjKaf7NMkhmNtoAeYFYQLa2lv5xIU2qdVfuO2qyi9+O0h
SF2HXJE/b4AoxTkKaQu0hulJKwB4CgVx3refaZD1/c/bDZsArR5iLmAeH7FJDrddbGUt5/kI0Gtp
72uv1Q+4nu2m+7hN2AfNYg2Hwd+vp2P7mUorH61/Xqq0n5UlFKt0yHFCjDsKtLnl8elfIlB4pXQU
g21+4bGs9gc3xTHHqUarTAXvyrx2LUxUMUWj5hMhlijQvskcMX7hN3HWqw/ZkYyGsvhs+wTN2Sjg
13nUOWYcOQRkYL/jicR/qMs1+NzLfTzhu5mDQyQz9EVFrcfK6tzu4XR5sjGXupoN66I7h8jThsvp
K3C6yqqbzcruOoOppC150iRsHgVhDrrd7RkPp+mvoXhkJBdMAlro2CHfoY/y6mxtw4ftTVqwSNXC
Aaufs9sUam7EbYyjFEZWWGShgvQG8dZeF9vlAP69BN8QpA5Nd80YhE8yg+PK+XGfo3BTdF3CEOas
GT62FhzR3VPYDfTCCmHTNDhCJIGqkUxGARL8vJmxrH8ZtJg1TlBI3Hw131Chp2nGlXbStPBJzdBZ
P2/+2F+hIweEmnCsG+OCvM4ZA2P4i42IAPcvhL6b6hzcqSFhpsvlSocIfUoinVGeNGlS2kv6GL/Q
FPWGbZ4hW/p2g6X5MyBXBnIVa+xftpvwsbQ8+oOtlufGf1YB7SsGrR6U9RUdkr5VuSS58RJ5tU7/
e2elRf11nAmqaM2ds0eWLI2lb+sLt+g/e7HdCzTMfz7m5qxWRxuaifA4U6KaNYDS2TWgkSkHHkTf
SQzqJ4sK82SbhwYGXO7+xwgP2h7w40/2ctRTLYoj49Fg5bcNliFHVRZX9K1FFcMLljETPEdaSR7Y
+B4NULXh2vjLRZaPSyliRSGAaRSSsTzDmTofNrzUQ8i7Cyw9O4a7WzpcFPeAtYOJBlv7gFXWHvqi
4PswWh+qj+rFZpAESoG4j3qlyplQcJBE+Z3fgmPykWCgHHCH3PMWXaIjCinKreHFHP4hxIa/YVGl
uN8G4ch5BFAZf9XC+0ht9hpcqMXO1Mst3Yh6cbCPs6HMG1krlmfCd4u08lJmhqXzCPwki6NsgMtF
C1iG0dUV7zpMzYVcLciB3UJA9o2CyWS4Uwv5zFsCay6Z2pauN353Lpc43kwgKcwEzQdwuvnawVMZ
cIMJT+mzSkBDGpyfV5C770uEjRSRmd3/5F4KUM7FM02thNHl5YSDf7T/vmCk1tXV36uOJRitLeBw
vZF2+/wVbArgzaSdA7/u7q/38DDC35ig7Iep74lTw+J4AONwDwqLd/uZ63nNwaRsI5gEoT4nF4Al
2OxdLbPP2DhCLlujYNKRkZwA/mMct2qugQVlVngYei/fNgzqTCW6B435ZI/5XWf/7Nnzg332sIya
ZTaNul1TLL+DugUsi7y5SKHxYZGQ26HXNGFm5whX+fiTMDD7K0SXSkGEDJwfFgiiUcq9fVv5u2jo
kqAEm2KKGlDClsJge5qqlGdClH34feUXf1lHTeUNXhaG+D+CEhVSJEHE+qLdpKkPDW0sitgyFWbE
XhOxYq0sqIiTGzAGw5qnLJCZBulycHld6Dk7mkdKHMjP6WPvHgJ9rRPW0LrH3BQRMPKTirPRXp0R
6X6I56ILeusiFY+atYdueUGlzHf6J2tk93GeBRAV+oF7zzcQcDcvW4LQc5/DsKom52fzOM0OuVoO
vr4cNG7IkbRRd0goy964I1TJSFqA9WOHQxiGz/eTU8wV3ZDYNyPUzzNcP/sgHZC2WFw2rLJnXPTO
W+gsmQXsQgHzpkpXhefDO4GSnzJLjlNjW3/jk/PQMa8y8/15BN/fmxgTK8vW7ad4iGg0xktdhEW3
amoWdBGvrNjBNw+caPsTUhBAruJGY7ictylfSx0yv1p3ZGAaRwdY9PZ9/702lm3NDoDV7qjqlJms
uC9NSRstbDg0Pc516nX4jiMkSlnGjHE1/AsAW/Hl3sjlUBhTIOpFcRt4CBrboSX3v1D8sX/3avJY
DPhSjG3rpCEwZ3pc+08tZR5MjWyAE/zV87m4WjDpfHEKkICeLomfFgBCYZeqBDnVFeL2JmvmbQZ1
WT/ZfhQ9aYM+noadlvPA9N0ZY1cinf/3YfY9bkTI+K3JZjJzeMTLXoVT3Tl66ud62aSEajfg3u/n
zL1X3g5ByIKgiyxx6s0Jt0b8E283Ui3PUjhGVGYZ+jfrCV8SEqkLVYMalXBzfdXcrf/qYj8vIhpX
4olCmq2bDbXBIkNGwsDxfl/q6/KCWfm1ZtD06FhCR1m8MMyVUbscsDCXUAgQAY1kvsi2uztSoAUh
XF0Tj0QC4tUFZMAwsCVaDQdwSzX5IjGye6VG0Hk7PEQiMI6pOtoW5+TruvNCpwwrI1fUPY/YmJNq
9LAgSXP64/zGph2iyTMnd246aLrdm+jmYWoP34v89c+/Ajr5r45ofa2Z8QPVwhQf+vFLPrzb/35b
87d+VhcwZlMME4q/110o5QaT5PGvNTwieRSUAeqFIyKb5Flz/C/C8jAw1ZyLxCV+m3L7Pxccj38n
0EkvBMHIMJebedaj608/V2ZJRXPBSEg7iS22zj61ko/lldUXJW/x1oyj7sID9QF1axb+OscYtMmW
BjLj4+MgAm0oSr9MuoGo+pHy/8x87dASCJYFAvJtE51xRRC/ofqnc2udkgQdpsGHxCq2QbLJfxcb
QENc/X5OW6bhu6SNnIkL1pM7jd6LXq8JBdr78ZJfwHwausDqngVfBM8ghogX8Y6Of3VFeIi9k7aq
y59WqROyr5vAXn0feO8Axz8X1aQP43xSJVe9oV2BVX9Rd8fcz5B98CBghsL66CwXcyoZBUy4dcKB
qr/U9oBYszyIGEuMwgPOKRWIY6EGo+Gybl8Q4fZ6yTT6V8bH9GoNTVFc4lkbt6J8rxt5lPCifMac
6Pc0dH09MbVxVr5H70Z9C2CvkEoOJh1qZCrMDZxvhkmORsNMja1KqYgM5HWqrhLs/kMN361CzsdO
UOFW4XUUi5RTSNusvN4e9hNCXg0P/meJAaELixQqm2Ale70PNRdlRpg4LlSWeD23wdaqNYzCCz6E
NePMx1LLV4TfIgGiFY0txqI2OWU/NgzpjHy1T0hq6aXOco5r5wiqd+QOhTM4uadUrGGIiMloUYjB
LlHXp+Vpm+lqUomhlFJz+buJN5G4DJE2U65S2LaaaHCcC+j9HpbQocVtrDL0l1M1xxS/Q9mkGrW9
UIAdibEBf4y+QYmy/q0d3zx+dO+13dnR8qDB3VKk4LvZc/wUhCBFl4qFHl7gzxMH8YPy1VgwqLbQ
5+dYwIE+QrabwWVtsnzpdlv1eq2lz6mIx5TI39x+lKrfs3v0zy81z0dVQ8Iy+xsZAjjgTf5hPt7W
EubXhOf68GPqpvPf94xwmj3BLDRM/jG0stFrTL5IK733rc1OL705dD9M11O4qlESqr9/O8+9oysr
lARtvYgkFaz0l/Di/Cy7LRe91ZkHErsqFEV7ses6LWK0gx8Hd0fbPiaDx1XPL6xhTjrBR8padDhw
mmBgMnOsfMIPG9MSt+qrUJBmbDHVWyYt9dy/XGj4qSt3D0C8ruo/xZnqvd6e4PqwJeR21zJhtDii
S5hDKp5vgjkuE+rKJy+K6ougoZ4Yx0S64zYtL5+c25RNbW36n3lADOWDGzB9pEGQ3rCHN1ZcCwEL
1Br3/CrlyQaWDPfUJx3W8Z+wV0RiELinPSpOIVX3CjE73Uf/S5U/fSP73IrKT5G59RYh/WFoDksq
Q4VQgdmjYwx3o19Y9HM527D0/ZvItLAHrmiKBETw5WbVojeMHk1oO+nDmGOWCya01DgMxd8edgDk
k2ptqyrvsXrsxxZzrDjwO4Og3Fyze8sM2Wy6Ue8y+uGhfh3cxOKOnmXEW8O3cV7HfDVBcWfHY/O4
bfkye+rVnSy/UKHTgRQZGO+6Yxgo0T8dUZGPTapTWbXxkp3Rjwyo/uLMNK4OThn7XlCBuFlR1IcJ
1s7HJvFkXwoQ6rZJ2EEMvBFFQJxFAOAls7/Y5HACitfI2mdOhTYrumKxAmr0eMTVVPFl453wZ56H
kGNqNgdO7shUjgkdlhCZjvkO24WL8fYGT3GnVea9/I2OAPYVQ/69z8Jd8LozBKa6b0skybEcRRTP
bRN05mjqy6FxnLfcnQ+tI2iDwWjXEqG0ZtMzU7ydwXQK0lUBmlkk9axGsXPEgaRqB65Ai+oehl0O
mAvbkdzFFUsP8+Y7B5GHgM0CYFRDFSASxUgEsK2NRQFi7pqFeGM0LuqrxQDzOWJFW2V6ej2yXA5G
/1/+FOnA7bW0n/+5cUws1O3J7svxr+2dXq06VKICVhwXaFIxDtcCEP1+yiMYv1GFGb5hqcR69Kzr
AewBhc7/GUoiuxUR1a2f7zPQWXdaIg/UOgAG3FicKhwfyAWKZ2seCm/hhbJkfsIRn9Wfvn2WoAXU
3jhhhTQdqajvPwi/rRsZdKsC0cQSrxqaStNNNgvbbsDwCzOpc+NUUll6PdvsfaQiNOqEHeN6S3Ro
AzfdW4cNnAN0aJnkenZAMpBikaYYnhcW06Jg1KLRu9jkIDAyXS8hb157hbFqFTI/hCGWBrJ+llJq
3px4kRaIffbqs53YCRiwPPPkU9qJofzQVPB/eqLWUMSIBMoHDH2GiPa5wWzMLyEFEKTNe0enUSiy
bqYEyTLfp/Mjg50aFS91gEjH/QBEpBLdEmiMmag0WzF3Pnk3KfJ1Cxq39o6WIk0cPb72TwIVbgbO
pCQxAMRcD3C+zNK5gAVeQjWZ6DRh4y+vYNuoztmiUN9Y+XUX8D9xJdOseHnjOeyrrj5Sc0tAP9So
tnNkR3MoO2zYL+FykR4IxY9J4z/NFeIaY9zV61JqfO6RklYpbtCcES0cYMSidTiz7kSLv/U3GcxB
48HjQo6rHdiruyTmTxoLRjvHMmLFKYyS1mu/BYSVOJBn4//OTZw/4ZXld9lg2iF/kbwCHGi/qc94
yyZxwQB4u83WzboA9yXphZAFFmbi8L5pG9pfuXWTClgzvGiREKbYn0eURtFn4g3xh8xpzwy+lrR7
SopRybatv7bSk9kKKuoURE59eyiIBEHJmUGODe3qzCDVsIfN/xchOiPeo6JRo8k1wEvQBN/irhk0
O5h9Czrdyi8EN5xO6WO3rjl9gr8S6PTlhv1jVzBHCoaVbWLRoxuFz+NItL5qbrwv+vJi+9uA/nZ/
TqlAPfzMDWVCdE73g5OtySyK8ydQZ6GJ6YSiHdKc0wGrPam0y13Vv7QP5uGFdjcgBL0lSLl8UvfZ
wJrVdOjofyVCryxR6Iywr7Xm6ijc/2F4kQ+YD0BWn03u6S/bQqETLpPkwMqP3BWpytveBriIZFpR
hcvbzKKm1fSdbJw1K/WACwk2Uqj7mxsVgLvCmVxR05ASI7bCJXNr+TTpEZ+18PJBWy+wPHam+VPG
83u06BU0oks3Ub7Pvd78ijLavwyWLMXv5p2FBzyr89HTGJbJJzzks292dK5mUbQHUm3qvw7CMEPQ
sx7ycpGoKK1ZmjNr5soAkmAyJ4HAhgqLmsbu7C18eMOLr4I4+oAlYqnFwEm6woE9KMBwqarqTMTF
ClP/XFeJav0X8qh8TukrDtivmp0UKxVGFILLp9g69LENtX7Uir1yJCGf0X1ljGrRNrEwqbqgNxWT
UWh0r2n1Vf+pGDjjljYVIxESoXVQZtiMM3ZhtTNiI9rWi4LoNI+ppzOxmKlOQBCLY5hoQb9cdOUr
w5Nh9lmCQNXkYREiojA0pVczJAGWbnCObEoBJ2LcNUe/agvlwzbhMG9c0JOe6EOdwvol5t7lGj58
VjFIMu4Du3hmsC7mxGIxZ/RaoZ3JKQ7w3JansMlJXawKKweTivNt/09+x1Iiyd5CFDPBeWTbdFB/
8ReBt4xAJj/N/ly+bt/CIhmYmiFSA5VnZSKKlbaU4ne5GSlj8TPRU6HH0pj6vxeyUG/j7cFxG+Qx
u8LlkHkgSKRaziYQR4uHaNUHC90GBlju3postJokOfX6XunnB4jOFh2vSGkgI9+IWgi0Q3Qx+4eZ
19hzB0BhBCihm++/Qwk6slq8TQRi/woaaDTCdknv9Vg5bXH/YQCnIzrrRMEGOy8pzNPTXHLeivG1
lhONKKqMakXttjc+RFwNJ2YCx8Mgrhdmi5J3vwBvn3IcnmHadzA/C3rkYy4jjW5VuzLpD1rKgnv4
wc2c8WCuXhhW+TwP7MWT6hxVdzNax8nFXQ8IL1Rzu9/DDDgKgNKwLm3SgPLgp8nC4/A6ECYLt+SJ
ZWInZt9HoPjDlgWaxtX3UjH0qYoAD2Fi5YIEtvdSiZuW2LCCEwv6tnwaupg//t/yqiObd7LnNafk
vpEuPUHtSCxsTiIlH4M75k2authOhzbljKK5p1E6nxAXOOKY6wPIne2i3vmOgxOTOgR7iiuYiLqv
czkPJKuXvodpYlcg4i0CneZgoJuShwju3C1+/6X3/PmRpBda3fJy7RuJI89R4IxjEKCT/g1BVS0F
7m8fNtOMccaYaO9aB7JMtNToBJ4biSen/MrAK+JUF7XyD9SOKZ8yTtCiJVoiLZob/KEQE8osCVT1
jAGE5IbfVTeKNjAR1445RsZ1nzllIp/uwYgn0+lbHt3hhp/o2cGK+kAFGaj46U1aF6Fk7JqT2t3J
3W5MA0YVcpwRmLm2LCvzmzXOGc1fyfy4O7X5Ak0GGx9djAFJBMMrtUZP5j6lgHU6WX6PNwRsWwR8
J1e4xyUXIfDebaHHAPMiUdwZRj6JNTm9dlAVzFKUkmrFQa6d7dx2vaeszMQ0hNLLQeTijZO/qNvu
MxeGz+svG5qFNw1tEt1Vm59f6HmiWkXAWdM2j2jt6kgzYwy7ZLvXv3vidyIEb5vGTXxIqi6y7Dws
MHfGvnph/SfUTBhhS8eUjcexSzrbOWruhDhy2hSvXl5jbsizkkMUb7pZ50CqQKodX5o8s+9cIXbK
QeAatpNhrhXZaZgpKiVF6gPCyMssOGukjnGQtAA+GaXFV37L/TluVoMNHbwtvxUR46wsbAOwlaKb
ur/5QbUX/sk/WUhSEUeHeXCSj+B4+qfd/y5wGbSwrtlUGZmKUu7BnDAsnJ36OWUk90Xt8T9YYve7
LRDrZjKIuVShFMO65dmPLvVbL4XKdG9Y/0oa8FWSZOS7TD1sF9dh19Ycu3nPkixPgFJbXcolm9GQ
ieIXy46iKrOzs4cFx/RiYFSENxUUGM6m0/A0GuhIBMVgIZS40fRuzENxbCSZiDil1tiwLilglSJT
RtNETEM7PKapI6+B/H5mLZ6VWjYZk9GD8ljwXPitqIkXRtpe313SRRP9MB1EC4jiW5REt4w0oPHB
2SHf3tYFyDNG6FcKaL80OatDQmxEhIOfkU4wU0Lj1FjvarliY/JQMQcvoxKrPp7euUN7kI2WZ3ig
zyjibnKzwQVQjwQvrDSF7gD1+dVkDhaF7yKXwL0PXyWArlmgPjH5cYdTmOcfpNN7uXJFunGkoIN1
Hf70IPTeCqmqJS+tWvA+wBEzahef9hUM5NN4u7T1PE7heqtmtoNZUw4uwpKuLuTr8Qrh4UN9NTrG
ehr4vOzZnLyqupOCUOCjoYAaDWwj3ksuMqFAZU+zU4eIaJRJmdabDSBTU8gzEWWVIKnpPW9pPQXm
uYZXJeoGmxHQi5mSa8gO/7zYG8SqFLD6FKf5V2Ps6sOgB7pGa+p0f4pP1pmtMO8vaCGs5icGTVUu
tlmnYb0Or1OUbO2y/glahDIc0jinG6hn8yfll24hDPLK7Jhv3SxRwdEwcRn2GsYflr5ctFfP/L2+
kMHVKcPOhzSqSiulS5C5LDcjCA/ltgHrReco0LMIQAix/SV78PYd12FlEZ2bmvG6myMcQkcd6XXT
Xhs3GN24B1f1WAIENBlNW1g3Rqt/nrjBptdm+X65bytYMPeG5VoEL3zX/x5zbAVEURFy4TaBpMMW
2b2PH19BZKxZkl0cnhLliEgWyYFG4uIqJbPnGHezqGf+i41JqG4RFBUJgfKLppzu8UAK+XXbuvxW
xIPbF8Xu4f70wcupehkCWwn/teKsLv4S4ACAjqWXEwBMGQQ35DO7JRFCbHknskZ9Zhtnl5XLe0LK
b7lsELhPdDvPF8VDr792Mn4F6Cfn1f/ha8u9WNsgaRdOX5GidanPB9ZXgHUPzswK88JxUXJY2eYO
r/luE4wPo484+aGsnkyKS37idrXKaZdCy+uqAF6RnUiBIh6lkNEJOgW6rp8ELFqM67fzIslluKm1
56eezHmqzEIrfrOOqhqm80v9E0UG/VqenmC31fmzkO4+ayCXWtePOqRkgmkK2r36HfCTFPL5HY6L
IBaJBYWpJFP91PguF/SwcZtu/JRdpgH83uzhxKCq6tlfzZ4QD6k2DUgdNex4AkxGlHMF9QbcVBNf
ljT2n2KYYXJv+A96SBZYPFWUm2JQLuKCkm33FzdwcDFZRFug9U7qrBz2ZmTeoBPydli7+PimKHy1
pWOOQFHsXiyYw/q0iurhYNnEzfuX9N5rvB0WlBCd+nRoeyrRDEcp4S8PQRzweGANquO69S3cKGmE
XKPLD36US+gyg7MF/CmmN+gDG+7lKdhtomX83Q50vLbyHGEqqnSrMnNlZwBExF8L/K1hJMSFVXQJ
o77UGNiFxGmlSEMiboO4PuL2sWttQECdP2QBTcBYOUivIFKKV/IBeXuO8HfK6rzuHaxANML72GIw
y1nf5n+m0NUrBd3J2C8qn92A/DUt2P9B6bUM8d7BaZRiCb7cKZ1c1N2zB38xbbcopyQDv7nOmSNa
qeuJWnvDw4dIrr7sFHqQuq0iDxozcqA0GIshk9E+96ObdVkgu3hIeWbA2Azy0nFppwgN/2we0Xgv
PhWUpyFXdARnzOqwXHWMPSf5ozhQnh533y96TAOuJTPt+TtPTXHVgtSWpyCHExzw1LHBl33noCq1
tY+7knuLifhgFiGSuF0IMWGrZ1ibOxScT2Z0L43VpCsa2QbfNRGq+RpixwFA6FwswNhcYtP5Pl45
aSF6+IsjJBggjZGBjnX8QWAKq610gH/jpPuwERT3jfCC7j5ITIHs9+82eNDkNMW95dYuIz4oLR3K
BfZog1ss4nN+CRrvj3Hx6AaTU+h3JpijJJ8kgN7f5CiJV7yycm87OCYO4wJBIdzE0lcZRjcaW3uH
X1bZn+Ufg98eRs5o1rxyFPCEhwm2/BKMLHVHiEEVS4ffiWDaqTJe5T7pwVG+bOKIUyvUK5OWoM/v
PNyNtx/D7ogXdaJDpDvd4bu0sOTEnVH7zuqRU8lBkOSxymBjIBvjGYNZBXFVmf8UHPVmF/lCg67W
0/G3w0ukdCF3pPfQm8vcW3O5MGX8oMORvsOs0pO1GmRQVzJIeTDWDPiYyIBIzIknT+T5yj7so4/Y
PgSK6g+ptRcziUOvPGKmOagBT+zfZMVIFfM2Al7kCMsMa631f9E1OpN9hAsoU1EZ5cqJDM2i0jhN
bnJWkv2Ls/SJUiQMILft2nLdD2ctL5gddWshu7EFVjbQ8boyAJSCSci3oero+h9d2Gqzw6ajfREJ
ss4XI/LqKnpt8R80I2x9BYXoXa/EVMuM0m7vyePbRfqejZlx5oqweM+P9zW8zD2RDV0RSGd09kCK
Fh8aGlU6kXDav0W2D0cVVMyI0S13SZ9G9xGoIrAIRO0bqXVrPwRlg7Xww4XniH6V5cZiUxFx8ChX
7WNgsu+RAFOsGhwvtqXdTNJ3bbRNOPVwpsnRN3N6k2+b64sdKcQNNnRDQJV5u7QHRX8PTVjKWO++
MUlFPuPmP8Y8JPC6Vq4YTURNTP0ePJTYAEniUuztxFPoqx3FFfYRkb6wZdpeO2swgmnTlbIWYKI0
/EO/L7snB8hJaXahHob1c65C3XjfpuPL5OnZ9VleBfFKipuSL/5b3oYFYnpb3mhkIOeZ6ZS4eQ2l
2SZdKVfUrXYycpKSiOqez9Fd2q4YYNMcCCQm3P/D4lLjPj6JJaDK90YsfeeEAS9zJGze/Dev+91/
KN6ToEPghxzdy6eMWe+6iuDD9gpYy6jMvttnOHCkP168vnseLbDT2VXIvjtx7Iq2pM7M3OY83Wis
Xoo8CcyeY+1mFg74kA3G5MQUxELwVhHcP0ocCJx4e4Z83XV9V6LtGTvNEq46Qs//89Z0boVA/ymE
cDA/pNFiOtyerarl05KI4X7AFxfaSyCRFGRC+N5B3ad4zxbkNyeyCQ4gnKqOOqf6I4DgM8r5myas
cikRbtGYMihXHTUVzxvbqxNPn7W5Ck+YRIKnoDaRoPo6VTK/yFkV0r9Zw3HjGKtmkk5m2kT7XCU6
+iLIZ7lNHQrNqvpfIp9oBNh6WLEW/40tcEB3srwfWGJTMUx81sO6uJiAqFLnvSvB/v2EFonpg0Ng
3+38STOLAJoRrBc5Pi9K/2bMzAMZKT3szPtqarrRxdLjnxxQquYAh/DHh54euzvVOfST+HltUO6O
XlfYR2g20mqfhUQ1dwCwRj1xbefuHXa/f84+8yiehQLilMjhPC+ijmhjsCB0T8zqQz5w+hAXuJiQ
oFqW0sl4rf7q+l4xQEJtobQIkyoNXnmXAHg9ylUFaVHA1Y6cnbsQ4CPK63Mk91aytoO9Y2BplpSJ
tA27G+lczUSa6kn96EWcght8LPLsXg+Md3K6LaL/njnyHseVX01zac2OABAX/ZtVcjqrJ90UTpTr
vmX22LPTMN43Q/+8wE4jl4h3LhM8eAIIfF9s8hCZYjinSoDcxOdtsVdal0+WPInh3kNUa6rPUJtd
vWjYYRmrJoHfVIx/J38s4kE2E7ld5zloM/AfS9KcURbYdN74H/rsaucoTqnUU0SOIarfWD0jg14V
ZVXCf168HaRfQjWaOPQb3dlAfLq7/DNXqEuodYQCbE5jqKSXip/CXFXtpUoRARxJrPakQDu5j9TL
2xOJjaRwFOoJF6syE6Ot3Za4HIq9gYjW4GoPhyqiFJ+712YuCAwFOJEQbWaviWRQE5lMimMnXtAo
jLMiuI+CNbpg2f4ktpmSo0bwUIbWE5lwH+W3hm8pho3Of7i7yWTGj69XM/jWTkMmZ6a+cXYR/9xE
ELc1bXGvHKxOlyc+GJTuRKAKtICQZ6qeTifTuTwYL6KrQ+3FZh+Bq0cDjAiSbG+oZ6UxvqI4TMeH
MmxLQUb2+F/+L+UdNnWNZ3/tmgQ1ENl04qnHoNMTq2FuCHc3d6FoVUUnWNBbBk9iYgJQEMPFBaIC
VjPcTV8c4vxb29Q7YPmWuKbZO87GoL+mDScS3qdQDX3rJhH3T1aRpfZ+vHc+9L062aaOP7NXTW9H
Xomqeg1PZ/OqnVj0cfTDV0TVWsAmuKza2/X9XkNd9k5UqEW0xnbN72iTYGYDjGGaFI7+UwcD+0Jw
teK9mGRMuBqoxqXwrH9NztkbMdXITN8hFBsGCCirTOz3sYLKKz384kQTed2wAkI9tHfSW9ll29RR
1msHpyKd6rQ0GHaq7BfAo4lzbMr4JvTWU6RnjPeElWR35os0ouPaF7EFaD4YLAGfiBJcFK6D/kFq
k+hSQ8rY0c5pLpr7BRGVn6hXjnV7/OCv97XhsNB8Rtg+WtAzQVkhcDHGEvw0X8mIlvsB+xldg5Oc
/b7Qqnzv+OicHG6sVCcyiNrHVppzV2BoZxZIe7+Uya5duXe9Vjz3mVANYSQs2OjRuooOKOFlcMAh
CcPilFYFz855VV+Ww6/A3d2Nxg8342jFNKGQM/lr84oS0bCEQ5vqFNxUfua5Kjt/sGgc3lUZsYUE
vhOjEFVecy12B+Xw5DE6qbX6/eKvfZhAqPchGv/xdsBEMJx/9q+kcKqi0lI3pxFArNBlWxbCd+uW
nQLUuar692UvTSpw3VEyUge3CF7RUbgWvsZDAKUKxUDLsNk/t1un33l7N4v09xVPKUsWMN8hiPTb
yGjfEbyhUa74yvnFd20ksfeTN24s4ucKoynt8F27pMiaTmTE6zJwI+8qrQ0Ky+6OKzlG9d/e5ai+
ZY5uSWufz0NTpjCREa4dL8V8zLh6UELrZK0PI9TO1sDKy9SRhNOzuIFcpF05d5G4SOYxpfJ/hnKT
msd90O7Cfg8pg71C3ZINvEuBZA5A1nRSiong9HFtbZULxwpiOYjbNBPmdrYsL0uDWzmqr0L6aHtv
eXqskMbGfDRrok5bkVjUCq5TaLgywKyT5CG3oytjaLsyD5ZQOTvKytO8AD1FyEqbCExi6BdFAH9B
xWSJJD88/cuP3UozovKRwl3o7pS1nIUD0MrF5wFSwAmQ4r01+9mSfwVSwrZrC8509APdtckPJVEk
JZsugDFLNPv1PWhF2C+FvqYJMcd1XYd+S36EH2zoeLdOHMGq+Gchvt6L7KUdm5N/WAFRZqsCmiOE
EcU8ILAoiblPtSFuFsXobrsyqikbEV/dwTcsa2Cj+GLfdKtysXtgCkScT49XmT15uEiHnWuzSoUC
rhFmUKVrdiq+s7n6hw/50CmVxVV3KTVXdTgB69MzfWwU+YAF7myV5INDp8Hib4SnSTo1JLALXqEX
3IVUUQ8BgPj98Up8rj8j1RA8ipjW+OPpyfD4z7IfotrEhlZQdqmQixxCM5lSw2JZRZodWq6+Q6MD
c+hzDQxkRrcR27BjgLTrNK8myEx1vluifiKgpxcMPpbvjuRU2DmRc/4z8k9HgPiwLWfM69SZeqTD
jQ9f+c35UFlxL9vVcXO9q7Avli5tqoJ8ecREHgIbxoiCt5ut0nVL2Ke+GbtuVtCaw9VkGx3ds1l3
6/Elt6+3sb5+uh4hCn4xNqImwvRT8FC4cKvyTNlhaxQ9Ig/Vj77yyIsIigJdRtpggOAo509vJhP2
LpfLicmcV9Vb0yAi0qF4qi75t1/cGla899iyK+Y9EfQJNKNOOGo0cujg4U1YcU7qe/Mb8vg+EJtl
IHfQlN2lROKbVqfzkcVK6jhSKDskA2d0/AYir11kmmyW4CrnIJJi/6njD4WZuhaNMMmGyDEJYJfb
ZiVoK6AZdGzNe3MY3UTqIBya3+2z6tpEYMh/VRIWYkzYpNwl4icOX2XaoAauGW/IK7GDoeeQsm6j
2ZOj1ZAc5S0Q/A9fUjiDAiBumEmBD+dfYlVaZIiwsg+Sp+NQA7NGM6GW0aBzAIQylZoYDIasMv8B
ei27q0NiazfbJo1cJjSgf+ZxBu8KoR+3YvhcCiwr91E5JP3joqGVc4qrg6HvArxjfRbNDIvc1H8v
wmTfYCZUhfXM1TEZOYR/bLUqDIeD1Z0KDYFwzyDPfRxZ7TErQCZ6dRjMZ4z/sKr02Au9E1pPSJTl
d/kCsiJ1QnDjqJ0gWxigTL0GAy0zL5aaEsiOxjzKzQ4sFEmhP1y0et4iYL6GLVnGarS4Pj3dLP9U
7AjhSq3toMh4vkNbx7BYk40J3IEBrWQoyquS8F6IqXW/8hhlkStg4o0S6j0d98w5KMA67VHxM8mn
7Mid1VRh8v+lEBcDYEXvDLEmp1xbhke76N26VHHg+JhE/qhI/B6PMUkDdklV0w3/xCgHyYPhdAjl
r8m1uPvNOX02gj0cjwy2gadH1w6oVzZVi6r5wuQG/XfumtIB9d4zulD62EhSIpjUPyfc5mFdiHwS
LtcrLIss2NDIcHmiXa5Rk29Ng5UPj1GgpdpMpdDdagrMCMxE9vnfFh7WHKOol3NNJSdiqJM7gEAi
rVdW+iEQjDOh+OwZ1wHTQ71n2f4jHnR0dY97kPnzy0/oW2YQLWIy93NJoQGcflxJhsuRV1iEQOio
jyLpMsGMeQXQ45zkuJmcE5BMIirw8ePvGIIS1TpUXBKEF0+EP0IoT80ZV13/jth7j0lIZzPRtEAA
iLrGM0ZbQPuBTYS3mdG0cabV3ccVYrTC5qlF1j2QGuCDlmBCaH62jBNkTGYTlI77Dm7TTrkr4v6e
WM8SySWCj7fkmYezYZD5TKX0XmoPciOJBVsXjRdiqiEuUeV4NsSkcx/HYGcX2XjAH+nvZjPuLmAo
uy+XVWC4PYi6rF59EvB7Gn1W7SykMsva+HbTWU0hPf0eam1JMddlaotu/sQz8eoe5peUMQwC9JDO
iBFeANa98mdgST19SxA3smIwtm/MkAZAz4PeB/0NzeuAXmuhEfj54+DW+StcwSloT/8C791uvzeR
pHJTheUs6yi7bzejhSzuEQKHCbiWRVwqyV/2GsUQsFA6tFBk8xQ8aoPMzTfTOra4q2Qy8g+5wf/s
UiD377p1BkxUIlW2DXbhS6BB2JqI238M6isK7CpjpXNZ1ry3/8Zw5VMpdbCSnNiEeaXU9OksJ42p
yz3X83GDztmsvhkBo5PdNJfQyyQJk2FYxJLg1cWgA+gk44SF0zkuHnDGewYNycUc8oCDES8fhGi1
+zYZSNvTUCu8EoKUIMRKcCtM6KkcdTCdAu1b0G1Dr08Iwx7pT6ziJxcIyvSQiOomSDf6DaS5RUEH
Z7x2seRoUj8kCMWwFgrPqUKp8IcFrrUhYwHhKtgjl+mwDw1kAf5I1MxBxaIAP2j1/5joE1zHX9LB
NfE9oooSP0bfBiHWDxchbKojHQhYaF5bJS5U4FaPfOzzYYv6n587UyaJWFMZ1NcbyoHoq8v/EDNk
G5JtF13MODrCvsJr3QcTktGkr45Fjwl4JvWjqgirbumjiW0H2Jtts04Iehr/6M21iT0vz7TaSvGt
gA9+swQH3oTW9Vz2Kx6FnZuBpVGsropVECJ7tVkgZ9+hTPCQunGP1ApeQqwejGgSKY3vG4GJfHQ5
PytTk/D66bQU85IMqHTIiuCjjW4AD1KzXqH76BHE4OUNxy9a8iWP5iVy1EYg1+5tEsrd1Mkrv9QN
10cRs2fmbrB+EtPvRqyJTEvp3RwSkGpYPOJ4cj2Z4f5hjlzt2GaSucGIw+VucmR64dqc+AQPz52Q
wifbgTTIA63HdfdqdfIwykMhmnhEKAcZe2QvUhqhKXhLszgjJZCqHWqVFAzDvu+59JlYEa0H6o31
ewYktc3gVGi1DYxQxurEuowLDBwEVTPsbRrlUL0ymH91R1ZEF1dfItYZ63DiFkXiRwgfSgduECp4
PxHxATAi0GtsDoErgIaVNUZ0pKz9OoZZReUvpjfnqMieOJLU72w1mGZIIZ5rALuXF7zgDaXnywfU
LJsqRIXN+/8oqCGyDiFjBqn5ITZjpKYTjJEwJE1Xle0MOSppeeLnXSMPRsz62fi/YIrArOH4V9RJ
xaJ9ZOOcFsnmT+P4pSoDUS87L9P37ESMtkmBkZEu3krBnPrFutEKGkQ8Kz5FRJ8LVtbKIOEhGgYP
nIFOR+Pye9jvjXiM4+S8QKhvOyChslvpUPvB/PQyBPtRU1SH19ObwAHuN4hAElibnJSQiIE+fa4A
NfYN1Qux6YwrD91rHc9a9B6YKjDHdzpf742rWV/KwpqW5iidrrNzNhbecQapxjDGC4OaO4wNvO2w
x+UJl+YF9xUqxouS6hlR01erYhJRAKj+5hFy6bjPBVjwIcDteIX4dAgbgQPt+3m6NYyUTPRSmSnG
fknkiZQGHelabvAaRlFboUtcCKbB8bY5uq7wrfJFK9b7Gofds5EGodfhhCTErC00TF7HDL9WnaU5
mrZIvsHB/UPLapFjMwbrqZOENdqyxzBtCrBFupRWpTpZwgmixTdSlg1igSh2Zz8Sq39TUMEDjSOo
7A62wHZHSk7pPlfxCp7cJ2pERsoebIv+JDfamXVaTM1mv9SNVgXmgMi7MbwfFSBppOmL7rHH95x4
oE4dbXFfjKTZr2LBO635TflBIHjH9mjF2TOwx+VEnYZF6sMQhUyNASijQ6tFiNx3Lx54b9PfCY6E
7747PokPE7MFKNpwg3csoYYPzPFXGXGHSO89YVUkW3WkvYvPFpKr4OKzvGtLRPBzlKIkEB/C//Tt
bSouSVVXFjaLBAw+RUmu8qZI9VTLLoZmHx6QPsyQ3Fsew9n089U5cZoHevsra16CXlPlg70buHmH
PwV5rT6VpoN7ufKlxm7SvNfq2hhGDM7gJOJ3j/OTAw8iS2WP+fxoKrp3CGCihOiB/up1Ev8uftdO
L8BXVRn/OSlYT0iHU+B0KmmypIdhQw5qohc51t20yOFlwIAGt4IO59aKJg3+JLehxxPHCVXV5my8
GvzJq/o5JPcezXZQXPof/nuzNBvxrSBsZ16Xrs0fEcocszKSC99x+U1j0ZAdNftSasd/oSOv2ccx
tRp0th21clafdpjVkVfcl5gdJEVgf9e55k3su8ND5kScoGvWxTnCFd1Bb+jq/gAqTaZdIAlMHUV2
PQGf3G47ptag+YYO9Fc91Roytz8N1Kubaf+UJ72Lmo7rMbzWr8rydrv65oPnNcZNLR8bPm147RD5
0w0E2tmUZD+Tg8guz713pqjV1huK5fKjJ1B0FGPhzIMCB3jrWd9AjLOvbIAQfMPrz2bt+LRgGWsD
LDLeG2vAKspaaRlLp+9PL9NoxD5zswK7GgpWykwf3MDJVKipoJSYZQAJCcBastMBsfUn6Q5y93HN
rZs/KFb7T6VcAwi5wlyXuI9Jrp9AqrymtSTWXl9sxWY/DvRpwLolt/d0XhmFnv7mhdpn7ZWEH/T+
GaV8erIvP+/d/j0sjr9BVS/wJndzmAAoh8BRyo5AsgwwARx5osZDaUo8x+oDvsx47Rhmf7WC85J6
kCUf0JIyMprkm+a3s5dpI8Qsg1ecOJT5s7U7Ewzd/sW7sieIoCSkZ7fYp9hjCR28Sdv+AhVzBseo
mgu9eh5GVuRaXDEUzYBUrn6NMDq3KxOMpxckiZpbrMAqE7hcs8lBCQXpxqIc4fyIyEoC8EARtHrq
ryTCjGPMdrqWh1iuhQDjyGK/oidWNajzEv/z5TDpy60apgf5rmBeBqyrNWF+Dm1SR6zCcIyzf8+q
9ehazw9LpnyUYFP+gI7X7i4NcND1ucrdmLWDafEYokTzMXPUbYuZNffoBrIKP+dcO8ZmPn3gKrgl
UfCyj+Lji5kiIgSIdGpXeR0jekn3gv/ld3W7z11McQzePwDuLPvzYzRJv2aVNeznGZSJvzYrEzDv
OxV+EJoXcm4I6b2/LOo0AhmMw7bc1SHBaiTnfwVjymlS9gKnNAXv+670RHdy7FweSb3dCrF5P74r
kwj1wsCyfeQ3nt71dmTj75Y8f76Wt1uW8oj6bqQ6K2r2JpUXH15FNRtE7Efe1Ne2dF8IgoMu8Llo
2nQuQYArpXl64t8Vjrm5c0TLiPuSQ46J+VRHd2JjlV8Ge6f4Ua9+WYXwEmu1jDQW/8yWaQBSFKX4
rizupe7qVW+fgf6IzY3phwFSf5ICHqn6TL7yOZxBPv5nLLNoMIab2WOB5odr3IN/kQYFnSngW1wG
gCTsMGHDVx/F6PyhQUH+G2T2nVb9XxkVAXLvEHgMwSFMguMcDEWsXH1KkksvV6dP9/cHn6rbbDBj
1cmWGGHnZewad7a/nq3O1imfX16bFH7/uuwI24Yv4QBZmFPuVv/lae2UTG9WWBb1GOAWnOrdek05
dKRJtu2EIdblJ5LUrdIZvv//DF/SlKnwUUK6F3APSyLAhk00/x+v9Hu+fjZlzZ1NEUecqckJaptI
fsc3L8xqI1/Kd/qXc10JCNU6E61VBMIye6kYa0Ywf/AmwtDrqwPDfISOpy9aTwzarte1i/EYPhYF
YcyIWkqyofkJJkvdtU04X5lbyK/T1xFEv6Ay8gf7QFqUlIbTlmI7CCM4XFsw+WPWlIkqSs6PHelV
oJHeB0ziBMV9MpsUhaIN++RJZ1hZySrlOO7hGd0GyHS4ZEY/3Seoshc5dV4mKxqcEz1A5GD2ALyl
aSlpn6uKW6vbEDuqi6Dbv5/Xss3hugHTmENK4t0PfCnwS8pEYWsbAXi82MOJ6FV1y1/bilZmxfzD
QFHud1HAGPRbNJrTn9lT2q/rnEMxy1Vza7OM+Ja3xlFJQJF1p8aGGr6HdfevWpcnyL1dJnmdiLC8
lxN7YvWEvtj9nPh75xU+ol9QmpmHS9qyjKVKFoKtF4hxIkczgonmyh0F/s93T4p0HMcxmEFjYiSN
+V6OKj9DBuQbQLHlhnhp5qgvlgRXlUyMQvXodZfaFlQj97mKwFtwl8XqKTJ6EmdENP9eEV/cYpog
T0Vh4JOAurovcgV4Aaa4hiM1Hd7KiD8Y7mHARb08rtYfFuF/EV8tbczQ5qOKQf6pK9D3rmDJFh9u
xzz2RittqIq9eQnfzw7IONPVOoBBXbXtn/R+mP19jfP5EQGQjPRCqUiScO0MiJ861BUVlgEFyKS/
1tadILi9xRjemkscP8Q+/M+lZ62tvgogS4tbl7Eaw0JBp7OPyJjH4s4NnEZwYPh4p5wrWaMzlcFM
JWWko0dNJrX4l/QqkKA/Eu/Vr8oz/vXiG5TZCb9bSrvhrkcq8huaLaFPEfLckufCk+FjvUykPLvR
DPQawxANUdzM6hcrFzSdcuDyNDttJtVTJ3i8VEj+fR56j/FVSGnA2T8sz8JpczFa2hMIBJum0pQO
sfGDbiQypE2IwEkSCe2Z56nLyxBNsCMYVTk0lzIkViS7ncNc6MVMauTrvhmVOr+Y1ikuPB6/7RKh
jpPpv9fSU5o6ESFPvgIApT71sQa9yBPtIgsXREELiVctetHsg9TQxD2Zp8Hag2V1x+nnGie4odl9
+bSM7LRYd/Hir/3wgYnyFNqemFt8V0GrASKt43xqXSWMnB3rpObcfgSYmYt4zHKNwgxpp743sIBx
E4ZIcPgVp18E5KhaO39pnbIrijEo7V6eYmgUJxe0/aqZ0xuBuRIcnHVPtWcbID/b+UeOaMyxK0KZ
XhlElUTFNpIDYi2pI/RaPhVhd3LBJjo17WCsCL41WBRimQanlUgPpSohaPf0vr/4w3DAMa39hOLs
EAtj0Ih8njBRIrMzAzbOzY44yqgq8XFWQv45aFb6Oqo1s4tHR8euVeuS0vOefoXuv+jgKBbGpRPv
urEK8Bz4OtmeXcxYNZs8MB3MyA2jaqVBH6GhQ7j1+ugUhkEh1tIptOYmgvhSJs2CbL+OK4nPfXsr
o5ihvHUuskKUXQgKPtbjJ3LGvSDwf1yg8CyrWZsZVZCin+5S80EhL16vzJoypL3pu7zr6H2mOq2L
fNIk5KtJzj04GooHPqpSIbkFCaRDOaXgY3wTTLpi85n8WVohKNu5/AvpwCq4D6FbmT/p3At2/6rB
R8LHMJsqhEfKZdNpIN4VHtTOyopjvnm6n/g60e12byUoCZCokP0sqfwULHzar2haN4GIzBZde3iA
qcfBZ0sGNaOvqHHLKai2LWUV9JVgHTLvkMFc3KA4TjfYgr97q3y5yJ7draaYlolbM/8pthQWWPa2
nyxc7udfEIm9TLof16TUNInhGeJtSQP1ipkqjYF8kcnX1cIEv/mDfphTzOnjH3X+HPA7SxYbYIh0
XKA+K1xXr0NRvR1m15oMlvheRAp84CTfbvY5KonYCRYZb0lEi7tmdwLvObZBL2T1MLUYyiHXMyCf
DXAWCZhDvNQFKSNO+1Wn+IaWtjkeca2L8CLnefVOlBe6n4Jeu3el7NF4P/L0AkDrdZBNiEb506Cp
RsSFvem3FlyblA7eu8johNyjKUuvPzaF5tTPgzNaLPLhHEbpUjyjnPlrz57d87x2RTiINYfJtNmo
Azc2RU46Yb9rZMm0mUjs2XM9lyOryYuiTkD0uFzOTAjEpJMN5WflVaorjO24+u+vh+MNYqcF9BI0
40LkZTHNB6b8rdg1h3zIYpL9n6WvcOG9G1GWY8wAY/ZCTwJWc2o3yi+piR9wB5+kBmEj//dCk0qd
EwA6RMGED2kDKQlficSwBtjdzRBZ4N3fq1irHwVIIuZd19mzlWxH+eZBIsUq7Pj63phP+AzTtrj1
V6dVjIsy/lhxqKXr4Y2yTTtEs9dc8ZHhRwYRvHVIeRLK7/NLN9hm1iFvYVEVaRTnZTNs7afHx4xR
kpyEMvJQ1jnY39JdRm1k24JYoUMU2ZCkajec+aN5NHIN6JysX6/Q8MURgCGCaNkIv1EVckScHB1t
L8bO9AaJ4RdXujfi7jUvmuTdj/R6lj27J17lC9tTa9nbE/FoSo9EtW6PsjK52fgsU2D2SJTT8zA6
yIztk+4VrN6TbsTy+OkXyUs+WYlT/2uhBId8DXOSooTkDc4E8df8+auOSDgw59tWlLFNpqcXDwtj
AegqATq3ylJLmiXV3+/08DnfM6qQHaI0BHeFXIHHTluBwFJE4Q9blWP9Mz5dJwpcGy8FQFk9d+Yy
TE2JcB6isZbT6EFBSlB0PqzEvj0DFt37Zo1lho2Fs05VdYyne7Dj7t8GvtpjztjbbiUjhwS8LCYx
kXRiYqZQBpb50YrWK8/8o2n6YGn2InSU5LUSJ+h8d+xQ+C9zqQNKzfcWAKSPh/RhS5Xl7qGEcHTD
idPKMqrsMLZhnzEQUsa8XfD2VhATdMq2oO8Ng4ok6sWEhYILZYs1jytJcZ3aXYQsZxDpdqpzWk97
bvGzY0hGYRpbp6gn8ssxuppbTOZsCK/GJIjf/f+/pJaM2sdbgBv5MCmyuMGFmYaBy0bO5E3MRr9o
53ErySnbHgGmns0rQljLe5OylGfS6+fIPU9fUSSmk8OEbuHrEvhAwocAUSv7VXxyvk8NIHwXzJDw
ol5Jg/ln7vAtqUPDfNujQeuIE/Nin6jHZlZUOQ8qVVqg4/Gx3axvVdK8fRhCO2pW7VebUw0EVN40
sUgqqwocOvXlso9tZIwpP8r0boK3NRHsmsUYQFbz+uKkvC59BwqREggTKsjdxDimAjD8R/QW7xPq
BVYR1rjYuODRtiD/KUExYjlgZ45kWP/+yhEDhyxE4pFViS5k10rn5NWk8limXiJTTJ54jBSONjdR
yy6JpNJDpHEknNb1dzlTUIMYTatTG0dpNSXSPjIj793ZF4y38mn+Hn7xzvfVzc0yDEDXU9U38M9o
QQMMOc2iVUSSHllFTux1aT+zjkryKqpezfmk4s57xV7l89MHVTc//mkH6ZtLfB/9T3V/DIoi3d/p
R8XjFtNg2M+1nJ0dNbCxd+TLauQ2bse1p+DPtgvFmpmWJgkTUMPEiJCwFV1MQsntbBTshpvH3yzg
/twKr1umi0bvuHP+nOZFUdku4/VRs8jtcYctQKQ29LJJM/UL76uHtCXp0S/6/+3WC6Sx5tghbb9O
u7dpGLl5qB4Kh4zk4QRbIOYe5LNxy4JXlPxW0Y0BPNgjFB27atLb+STVasepniPnge4h9ygcpNLs
Bo0ISgn/DpKVZKKZqYNtIXognW7S7BhG/ltn+zV+18/vKDmT7vKRo+ToNy+J3pnxvQFY5DTFzoH4
wu/HF1A8cyLO7J2+8x0WcqJ2gX3Pbme+NZwRXK/8R/AZb+7WvujEHcdfI3hgMjgCM8+P9ilEI+Ev
UjfDTWMyLpXIXPlwS1JfVLpgMOjaZeVzCHTSuouA5IZ+YRX+26Lc20kjzfeU1ZbgNrfwnPaGXR6r
EmXkYDU2IVjCJ5fqhx9mUNAwLK6rsBQmPbYS2D+rRLjz0ct/lUmfas3mVaAxy7CA/tBuDXOXOi7w
yQ4GBXY1UCL4zE9BPyE+5hzAcOgmU3XryVPrFkIKGSCX6447hfhqAjoEZQvQfjZbQDi54X092ZdC
zD8p2Sbzg+Lyu9QZIq4RC+KXWbMCXmjpTXqB9CnKIlldiTZMLBUC2xRSwaipfBJdcPEr6FfvEnSQ
jedmtmukNXCKVT61F9rtAxNuQ48/NiaXDXslG+EQI/TgXHLpUKkdESFj11fys5zzZ4t3EG+/ALY5
TmxBaJfIB/n2pyMmPKGi3rUBrV4EDTdIfCG6e3PYdJZwf34X6d9wn53+o7slaj58lJniVQxB7sKQ
bJDwAZB1tjrva/a03c7j0UeR3pOj7xzTg4RqwNzAHnV6ywuv+grB9oVl24N0PNrL0ZvNDIyQ+rBY
3vTO8pzDEZ+x2fJT+F250hajQYAlqnXPeYUtFTo+CiC1QRzqukmnGR0nlNq0gMXxZ3xa7xtQh7wo
slQHpeQAgDfEoSGndoNfATMZSYq2+fWwM0m6jq3THzvJVs0X/hHLJmQvZSAnkXluDJ/0SFt/HqcM
FND9HNWyqH/9V3kl5kp1NNcEemgcN3rl4sJtMYCQFjvvvdbs+W5qoj6D6o29fvvFZ7rR7XoJbILL
SOt7ijUbPS1tehiQhoox3ilv/K/pyOgXGEIKPe0OHEOw/ZRc2zsbU3vztsLxWgve0PXi5kwyHlJJ
LeONbgyIdbQ6nRqLUsFVxP5REcjTjmxfNrNCSgu+tHCz3IDX9BjFWP/HMxBTmoTA6Eh4yocIDbeR
ZY7STaEibM626MGByzmaH9R/qtF/596jcKBYjTdChYrJxcmqBDmpIMa1zIKcmvj+KllXcqPphRjI
Aw+fFZrTMq5XS11wBi4jm0gi7M6PMv+1ZmC9BhoiTCrF0+CcIJdFyFSWQDYkoVh7fma7CGGtLpio
6UInfiNgSxNiwg4lpbIPQx166ibKiIEZPxFDVvJmB1Ah2DlyTitIUPEVq+e5K1KjJfZYTVInQBMo
KmpKgeeT/fTeAGjgXiqkYW94n8XyXKJiR2J/wg1va5h8kTSjFikMvi83TrfsK/i0oPsypMHXmne0
dC3MajMXrz2GUGme/pd3DGBvdY8fv0uBxhPjinUgSZF2E/r3iEAHWVzsfhAAo3TY+2/JvgP4olv+
GzEl7vKj+alls+S9bKzbYJRPZXihc4RzeKRfg4c4v6CrodtBntsbQGlOzBlGU3WZmW01xLIC2HE4
qncB4Pd9HywQD9WRytOZMZ69Zz+WQi0jb5Rv0j2h9q/2IXBfPJVT0+va3J/HrCf/r511Mu5//Cq0
1hVlivLPbIGXNqQN/FgpY1Ak/BjFZ7AOyuTY/PeU5+Y19Hx/mScAwhr5epcvBXwMNH01R+15t+I6
blvyOyZhnj1vWokZRKzo+qlib8gslYMPXiHJ+d8r25lQ2uJbsR+ug8I9I2ZkYGYqBqT3VoDwTTmw
Q/p2iEQMlaZjh0jTrNkAbDULRE2UarzBb9u8JCo0NMB8QryTRNrv/OmVrLUar2a7IYXSZS6n0nga
JEnnG+0JAunQjt/rJ7C24tOPvJnEXGe7IJakbw2w/gibthHZzknSK8NKXaqRDsFN7Xvi0/S0tNHL
V44mclvh2OLfq35NRUYju9nTXuf5bk2DcotBluYfH13//w/3zspYQUgO/zOisLEDxwmXBsPCV0Xv
mAx97q2afMInzVWlFPpE3fbEAA1FSAzxJrDSWri9+rFlEQcCuBs7NIQkAs8ggRlc6v53jUfAR6WV
IQOFnzbU2hj2DyQExvpTaWRuY013vP4NZCnqdd5LCy5S50iTmf2x6EFgDlIIZExhqU7XHMLKo7OD
JYX2iik8VE17P/1fyQyi/zMt9txPpgwtH1yJYZipSBvW9U6hqtMYlwSjGcSUBZV1IZT2yZxM3D8S
HwDeeM+qQe6ugCS9GKhE5wRQJQzw7+hs81lbYmnbUdUY+L81lVSHJIy9uSvfpuh6dZc5/8ybu/w8
pR3tnq7fP/NrarvMg9/9YYkU2WWBtGn5bOLkFu7Vo8tTqdM/eR7Y1XpdaHW/5NZcTwHVr0tXmDLF
p3vkuRms+4as0dvrp2D6TtbieXNTUm02PanzWIIlOX/e4syPEvK1doWtSmMMrfvO7xo9lmqpv0AO
aucWYvH1rMiW9Q3+B/MX6WFuKvRboc3Wmk89u6WFXGpiGgAxqftRKn35dug/TWajfZfPTPBdfmhg
80JqvAcveNq9ugnxI9No2Du3jb9vXwCG8Sr6e2p0F6TlZuThdLteRVNUaG6ini+FHo3u4V6goaBz
QgYVyCjS+YGQ1bzobKVuf75pyvMZEdSW5fWyzFcR70VjDeuRQWydtBg/xNKaJVG+qfNmH0+gROjr
QYcb09ZR5SAAwH4ximcFeRXNGT+9UYX6bVTxm7MffcNddr1cuwAjkOyEIt46+nYpaB2ymyX4gGYx
x+2z2T/eGUmk05UeDeFkSFzIHKBsFo3sJDaS7WeRQ7PzcmJQoSPtYiwFn+vLXq6fXGTmBzaxBi72
SDXsvst5e36S2H+CCfR9oNSU/mfR0/y7yo2EN/xyqSZ7tXDURY4Vux3F4t/7Oici+k8mkGNDyiXo
YpgYO87bzEt98StpE0FyyULz3cewxDOQlazozQRLB8+xhWuS26wdtbPE3O83HSdnN1HcwR2+uxD4
79Y1TGkqHr2ZSqHEnAkiMDixjTo5JR2kZNZbJRwDqN06zPheA5lVf1B0OK6EZIVijYXT4JSmacpe
4KA8LpA6bNn3cLbhFvo+Vf4kUC6alfkw+Pwgd3ZNhdXglxx/sMZnmbK8VIGAFq/qtQEJLpKzSoGe
F8/TTb2JGLXq7lwfQ5UFBAr9XS+alsuNv2UQoxiVj3dkchUnBxeCBhTl5/fJeqTxqWNmMGJDNbge
R7Sl8OtZZAh7mCG27qnC1G8thXDtSNr8nOmyC9Qg+LyczcqRSE5rVA9Dy2aMW0KCdW/W++IFWDpx
TEBS0UZQcWaKEZFzZAgBAuzfwCDyVtSPGGwZlb1qYPGwbGw6AxN16wUUmm519XrZvc+CXRW3oB1x
C8wtPsdGSB9/uCm53RNQuU7TRRqPX81luAeI7zc4B6YUZqljJJ+CyAa41uAjK4uL5Lv5ogzdRvKP
+/70CqBeNkiHGkj/50w0VRZ88cIcqZz+nBSDJ5Y7mtJsHfMbT6P0LHhxhL27uV59fmBdYWxuVt5k
Vk/87EJMbtGAO1dVNUfwiOunpU7Sda6lltzeBLCqo0xHNCD+3MAzKj+hKb6a4buYMVygWVLv0Q3g
VFAfwaDroL8j5G+atM12Ajfi3OCpfIcW7u6ymU11qWonPbHD1DpTVYqWhQysS0oD1tvMUjUClmkj
una7KYqCKrk6bLv7xI8hw1oYK+c6+wgRyhu2+amm1N4UdM4yd3HUzfXLQvY6Ck6OYwIxK4nPdpBG
rOqfyrChve3UbRvtL7K9eh1qu+EawT3wDrIXJgpCNwid4RTasw3DSx8Wi1TtlL/b3yBvBsKOE9xJ
+e6JcMaBb6rzUpC6RfMqkBdqx8avkNQd/yp1+Uhe9pqg9ucHByUemPxkb/n16crYbtL4KZS2qIj9
V/ox7dPmsNAt44pGLpdUYhwObgh2sqJZ1KxrY4s1jNhPEYgWx1IXIqGs4N8cGMX3jHw5PETbY0nr
jAR9cVhoSeVNHR/k9CLMUJwNshuYJc+7q/QqWVfFPW9XcSkW0SFJUxa4+sgy7EXd858WiSb8jget
ArJm/zjUNJ/G2kVUoYeP554sOEkjhNtOHYM8uVj2pRrrBurEw3JcNr6jRV0asxigj8vNBovyVlRX
D0E8+8x3kwc/jH2r0h+N4gAOKbhG2E9xJpWDYSr9I+MlfrHC2vureXxvrIeA1YmcmLpAkWVGOrlY
mtYBok5MAc66PzO5i4DeqCCYZs5ZDOwZuxPrJmnr5fwDca4+pxHvphmf+GR0G6s2t6nwIM/qBZZe
xQHaZr5Yj6OLMLOS/Q0olJnHGZMfmKHDMoTMPT6ry5hnC3Gdknk2DBhSkAcHxjnYrmZwWVvyFtmk
XOsdoHDlhQN5on1oh/DDVUzLRsXx13iV7E6jsgmUHL9RtH1s9tvOW/xWMOfEmt2BznLLFTc8YJ4+
qvbAhfoFujPNP2rsc5595Yh+EWtlSDdacEcwVgjmRp61lWYlIdr+SF51W2+EqsEh1uGrd5rCKUKN
W6q6o9Ua3DJG9LkJEUOwD3cJ129y8x5nPoEU7cA+OoClqSo92/u1eG1gbRgD81f8ABVzgl2ei3D/
B6Yq7BN3k8caI1K+Y2NoC8d2DmBbVdzPiue8ihZXmz99nZknfNbxX9vyodCgyNeyyJAQyQ8KV+Hz
hGBqXIXm1a2p/oJf+AMqPeINj+O/L2PgcxHOeJm/1gVp+1SfG2TesqsgwNmJKtN6bljoGaH/xfok
pMa2XRc9bWLfWMAFkyDDY+o3Pdn3v1x+DX+4s3N7Y1SS23ZO9upQrsYT4JNBTl4l5s60PutOc2cE
vGMkYQP2ZoFe9VRLCGO8F2LgZkxeEkmhdaDynqtrHu6OHFPbT+I/pb6nLk7avIP2fgoqGBud/Ibu
VDhdFmcin39eFyRW4dbEvX9bg/0whJ4dUghe6YmTNoUBJEZZwu82UFqvjtXUGwbDVwymk3+x4nFl
quqP+hKncVcO9VZIBhZTBULIo1dRqwdeY2Ox6fDipmdRdkp3mZ4AgwAS11ZTjd6c+p0Xi8+Kp79y
DfXpdFnjDwhbnflESr551jE74HUUM5OBiEGNd+3chPkOMSq/lYAsEdVDmsQiXuc6Ars59ey3nB0P
QxCRCqDAqTyHvlqtr0KyHCDUO7kygJ1BX/LqjqG/Az4wMRm6WOStpsYcBUkXwTEpZRQVqOAQPNxF
v5p04C6wn54mR3b3qrziBrtztcfOEhA21lBaOI6D2XOnIL+AW/axJjpipGxQ1JqpV0CtJZUQZA6G
6CBNp37gFjkX+SDiM3uISooUsX1mxGsNRkocGsbuYy1JioQ2tlWJP+2CXEMI9JkshEAdyIilM6yg
qtN38q0k0lJnv7DlWWaGLdAFPBkeYDfOyztZhc+Ye+i0f4BD67hvZt0MDH/qgl3eHUEh3GRMTPi8
4ZVYaTRwWiTaS5E1SUkaGvmRL3iMdjHaYEY9qGpXSCbn75pWd/VUlOSs+Uc/zVOn6bS03hdVLvcn
zdn9pFqDK3KAjv9Gyy7DbpyTYmr9C8Ht44Y+s/AyLXAWDsE0PWTfntbimjEFpBsv01t7rZ/drH4h
HnguU8ehuvuqkaU9YyGhab4Lvhgx7XE6KQuMaknl9Szs9MXUdbnGYCVzbtfBqeA2xDeJYrZsUBka
gpc3tHBJjXWE8RcPW6RMd5gEQMSfXDyeuf/8GWk98+aVuiwo2S3JGrkFtL4Qh2ayuR8l5yEom09A
r9AbpDfMAquCruNv1IOBnbX3XyWnwbVL1gU278Z0tKjkX/7gqiq0EfwBJIKZwxVpt0lFKlHfOyRx
4ciCSNt1rxKiKWf9uI6Dvvcx4kkqWL484fGyQIuqi8fh8xDAvc+oNB49Tnzu9PHg7MFKYG1J4ami
gQmBCLOKJkJpDSxNw4dsZi4hdOMXIirTs6/MiAOSD7TcOSOaoPxySnTHI6qc6oh70rdNqAYUYWm0
LOOPbFTI9u9vdzjUy/GGqX5k9m+8yg8dwv2JiJPJkll0DI3KWZ7vMTB3SPn0gPXTTSU6FGBFnSWT
qo0+E4DsRNQGDf5a20PmtHQXtWe+xRUf+n2+PgR8uUacAmyz6xpeV9AJCFg9UokI0Uo0EQUqkisc
BqVpWDAj/+29ulQv3Ndahb+Hl31WRyw1zFMhLOax/ed26lanSOYgR/8fKRwfdzvBg9TpKr8NERtU
jV+ADMfRSaeBVxnMvvPcwP6QNuLugEnnRyMEOFAmfX4lBNboqu5FwFxRwyRMAFTCcfGoVp0O7BlC
7UuBFEikKGfEKMnlHqe2nsanmB6TKi8Jap9QLY5Glrbyas8GQi9o1lOFO9TmfjTvDHdGg+jbSVPi
Van5t/9wklDNuUFMtOyvFsjwmz/gXnPE7NtkOafbsnU3mOwM4MANqI8tdAQX7rjoBb6rL2eYbXfl
6WnYme66vq8E7xhneT4Y6KYX8VyB11TFI7axA8lrioGKNlzeH6DoOPWN33gnPKiJjVdLXXWEpM7l
7Eo8ZoxMB6Kn0dfPXXizIQXQWni+nsN5wuIIGvgJ/66SS+s0W9QiEnhr/d34enLE+cVxZtGFYm5a
KiEClSKGyRpmEhJushvK5DT0RO1KXM3480B8OTHh+q7EM47K43cyVyzEfm9Q+N49m7TanEwbdDI2
S7P4CbjWeU/leNKBFJiKzf0WtjmM9CaqhEowWCX7lvTvwyLGITykOGIHOy7Wh4E63r/i6S0SkEiI
6Snk9Z4BILJDq6S0LX4+ctGShpLPU8YuKknLO6gc/hL/yiofkDx8TxsJCWHwI/HagDnL8FNYn4bs
7+hN9kSn58D1oftKdzCY8TDGB0DeUCD00rLp/U5OlSXCRAT3V3UO9qUrDEV6hLtr2/MxxGA8h1ep
x9NPaNN+2GtbUFRkk1pRPg9DvJluldQBJk3ePN6VALWgYq0s0iI0W5YUlEAgdV/auY8nSJUpWJrg
pvj9G78wwGJnErbw5gKXfEsWNKoZHswld+ljggXKGdS8ajhzi6pCSWgdt3optphnEHijgDDqYEiO
tqCFr4fClBQHGeZO7xF+3xEEzxAdFRq//2Z7ygnQZ3OIKgC61OmroZPCc9BqwZ3bpqgxhuJUR9+h
ptS9QtoDGvoyWmQdoozAnHG4JdkxuKl1gSYTqzGmBRsNjBKPaWnE2JpvY7xzFkJTiGXFU8+7K98I
SxRy7q0FIc0+c3YLv9NoIukSkharJbPDCGvGj2J8RUIU0yw17nvvG/xOkwF86gbEQaUFJEJVFgB3
aeq9E7LAlIk42BLBpv0TTFQ74/KJK0hVNIVSTHvT9KdnK/aIZRklMH710KF15M+i0X8l8niaiW1f
5YIkerRVMOpkQiQDl9PCyfulmn8phFpAAFe3VuY1uXWfOoI2NxkWpVXdqPjvT0LBP0cLGFgmZUqm
GDW6MtzAs0Dzh5rRA7clprjZtlaE5bSYreHY21SGoxZeyQdyKpuGw5tAU5AkEhiy1RNc0+idL8PD
7V3IWjWBHhx1SnP659W5EvMZ3C1fq1MQqlsh6AonxulVatQjbSXs2CnhhT6Bcn+HT4qmGHk0neXx
Px0o9aqWZurWgdKHpCj1DqQAgGDQowj9nsQE5fCKBVkyHhdQZUaYpZk3hPiDdVEkpY3lYwOEVNQp
iyoh3Vi/oiM44mSL2O/3OJYNc5qcSsKP2dtvubJcycvFq2z7AubZsWVIVbvYqWxBVpXFVcwthHJX
S01tod7C3F1yoGzc77QldsNTDWTvIzTTfhKW4cdNeYDYuKXvX0iO2xgtJm7alL6Q/8T9xTkBi1D9
ZJmxoBEvAnfyVPjlrAZ9gsPCCnXSuySNCPhDoRQi4bW9suHW0JBTYpV7QB+h238zYiICikX4Fcai
y5wnz7E7Qi6WaQ7DqSAXka0BnMBEdItQMzTTWX+bgCnbk0JoP4rIfywnSv6guAZEiaSb3cCvL8rv
FhAy4uh8K1OxhxtrXGiEvsY6qOL9QrdZnfVMQd35a3HZZ3ghKhrfeaT1sABXAmkXMfC41lMlJHrP
BNAUkvoVBfMc9RoTPRb3uNJ4wYIvJBjZbFM6Pg6qzADZy4FtwHpuUaslPOickIMWh/kMaV50IO0T
BToWN4NKL4+WOWUhIvC9/tcdOhpcvD4N3nPFWlHG3Ykjr9ChSZSHNWPJ3vnh9AO/6UGbTV2zXCT2
iB1X0pRabKV2swM/q23/AD0ie3VfSnlzgXAdXGVek4x4QGGXDdJdILrg1LO4Xe/HqCRLrSnwz0LX
vIKOMGddMM+N69Le35aAgC8tcEKtaIuBA+mHnyjo6mMUK6OhriyltPDGny1nQDkLIKSQ2iIjze2G
83KaQ0u6COMBRsuLiy13tI+IAO7emmg6tVET6xVcxHuJbceygVmcmduod/E6XdSfVn27GyAJRrM7
+iUCmSO+jgp4c06zm9XTij8QKYGrDUz1IAjlC85godyp2sHB+ZuvxKhUivyo0WHJ+U0p6h/l4HrZ
YDfYkB4Kg7FkACF2c0kyGyi9Ls3mS27M5IJU5Rk+eUBLhzqEk6BV9+K47jG7CFRkU040PMGx3I0L
W8M7pWk58PC0116T9OORLpVborgTlTqgaeVnWOn5j0beINq7TZgS85DAoEJWWEjByhdFJvl+MxXe
QUh5ttddGZOaWicpALEdkFm7YmB1yfMgjQTPDau7L7x3O++EnUhs82pPQp1XKxVniv4qIe3uXWcH
EAJWZ8G+nK5fi2Tpeh8qxihJy1L6JHSSXUKKrCI8vnpCT7AGpsaacYewXVnIFezGOfAbSzRIW9gi
viO7QNHhJaVWwDMhwcOFoV6jtQNPSrdM0t05KTFjq3jtfuHZBMvo7rjF0SfeIlIA0H/ZdsNneht8
NvBHvzk6GNqqqsr9mt1RUJXAu4N0vn1L1XJicaQOZ9NOefkbXBCmXgiAOR+9qoFl3i+neXzrSbLv
U79olpouJAs5Zikw7vAngWS87rX7hu1kucj0w5CY2BG+6F/GJJeHNZuBbDJ51jqIoeb5YxOeWPUJ
nFLvPbP4z7421h/N2K4HYhzLiVN5d/LfktjPgH4cRWDesmoYkiHd39AH3vx/oww6yZgiv6p9jzz6
KaT7GVaKtnY3t9kkfG/qTANU1q4FYwRFcmsg6f2SN+BdnTSXRMXjND9BKz6nlzIFf4MZAskcFia+
FuUALicGcr4QfJTqLSlKez9f3qp14+hNJ2YoIibBpEwmi8gPt5eRuDf1xlehXnodIDwxnwwhKTxU
ghdfiCNNW7c3XkxQnAVWHbWwSVgoZP3ggsA1HzFONw4NHQXiNL3VWvTiWODhUmG6zLZWALbj5ZbM
ZROiVI5efTtBWrPzrK5sUC5Nl5nqS1OBkwv2O8Ifwiaxb8woJi0E0p5x1IW3P4AlYfkb1w9gnty2
rOwxQy6QbotaCTMw2sCHnZezslpoGZiJ5BmWH5+sFSijvkvkN9csVDK/XLdHyQPIBeTefaDvn60J
6BV4JPGbHZ2t8WzVDZBrGgPUmbtlDj92F7FzhVjDYmY23kmYMnTPzFDSq1UlLRNa64C/85cMryZ9
cQxb/+QI1Rrpt3RjLVO77CvYN7i+GjyFGi1+cX8q2531OJLIWHB51oVUWtFLBpfFiv5QmE25pMgH
2o+Vsy6ByEoD6gpBEWBUIghXlxyQ6JxYak2gwykSJH42ejYueRUFISVVGuX8xLHFavz2PRZBKsch
9wY5ztNEwRslqgQtmL9cNDiEaASyBO5kikMbCXIo3Vqj9VOEVZhwkOO6fvHsskHWhu/0CIDGYYcu
HdqklXiZL56aVWYk+3n/882cCEVy1Lwq9gEmXkJYnpGzABl7CH/fOyJhMZU9rqllvOteuLMLnWlR
7U2IRRCYu+lHRIG+Q+CkCmUG2ioMx7L2iunazdI4zfVQyjpABhru3SPRF+3f8q/jGevcaolh1OxU
q7tO9j+b/VqxIGzTzpvlM2p9B/dXGMi7bJvbtSYvz/RMofR1c4dvkpSHKR6PkwvQbkiRq8SVNd5P
LlG7Osj5OUTBDyGgh4N0Fy/3ApFooV7ZPj5Sjdn9ptjB0MpDXUxE1aBgROlQ0tKGGHo+7/XsKWkX
rVdjrIynA4MUb5LWA8mnXjsH1P7hobWwADWipvTD/nQRjbjzsM6pH/9/Cm767Ht+oL81XTA87Si1
deblul99CDfSK06VpzhEQARwuqzCfQeE7sjv8XDLW/R2p8GRBfAdCZX9Mk4QVlpUifNh397eM01q
9CHBCPZBdESztJfwpuOMYlM8wVXYhGXSEaEbJVgoIIBfvgniuaaXmYrqM/Jt/oTHSFvtu0/Q2dnv
Ro2EIZDb7Jb4YVtHSxZPN0Gb+ySfUWxfX2H4JXrTf4jj3n+6bENZYa7VPBbhz2ep/Dod13L7RBcI
KS/gw7H//4UqDvE9vBeRZL7Zkz7Uwyx+0iB3oJl4nh8+zNloSV/F8+nb5lcYUCbnzgj0xKGTprjm
zvQp0tTuPqbDcu8v1+RcfOwaI2emFOOAgDfuRTnBmWoZUh40mmrslhhVBh+hkJyc1KLT9vgDvENV
dSmZHMImaePZ3NJ+RSXApJnPHSkMFlnk9isYYKemZfCBQdFCTclctgwwhjUvPhmYTcoLejN6fhiV
GhibTxcLKSHZ6NTs17yXfDgoJTBP676GAHjIOYP7XKGx1DdlQgZ2Adb7s/1GupBcxsKe5oDwjMf6
Dcc+eYe51QMBW2OM+oX2/jiMmigLHclu3ozH8dz0gVdGOZgSYEgRqFRoJFqkkWRHQk81aopIxhvK
EyR3U9lvsNQWJ4cxZ2vS2mlNPgMLrTqCg4k3xFxLuhlDLgGtCWOb56NCDWAw3qQ3dhvzHzuClcKN
jF1XQ/yHzqrLvk7piHufkgUHp6rYx4khINI/kBOENcwR5TBEYL7Vv9qSCG4qG/kurILhc5Obc5qv
5gVPBdQ7sZTQpZ2p2Fe/3Okitb+E1Dz1p+IJARPXOsrcjBfKYxXXAJdrszFc7mHX7TLvf2v56Gov
Irl+Lk4+G22w6lt1Upn9XOD6jQ7F0H1idjZ/X1B+U10cfHflJb0qzQkT4j/QaoTwDL4R4GXGA+8j
tPz4154Yf2BLqDXC4v9HNJT8Gb4D6xWbyeIlJMZJsFAMvUMOY5vxnAEkBStcS+xxEssRnifUmPpZ
QnaA32y2rd/PO4nhhkGo2+WMwFU6/YAEJoBeEqtWza1pBAQccEeBNJEnfMFSNoQCVAtXulvDWodo
v2Dejy0xJBN7qSOfWk/tviJNIF+qJeLVPMjDMhChHMBCJIwN5lN965p1IVyWQLHnHac4CvVYJV6R
2vHgqz9eiYt4esVy+jx08/sbdxXfb97tP6EWudoRIhPW+gs1G01HXMmBF2RQqE5Zo3UJSyKISKQq
2HaIVEfW11Kqo+kRAEARyMV6HUBwmvjKE2Jwk1HNUU7aze1eWMFhfnwfCM4N+4MVNJq3fk6VQrob
3R0u23sn7KKPktG1Grn4UFc29z0mUOf6udFis0uiapCpid0wcK7N9Nsj4cTXlTPoGMJDkBIyFW/b
kMKAyJOOFPzGbjusAOkhxymSV3F4e2fnzuboD3mcQl2dmDBBiU+0mld1KM03Df4DAtw+Ui6D1t5l
SWRtXVoTUdL4qQGRTY4FVRO5lVyWVxdFE+ZyuDCS4ryctrqDFCG7czme5OWDZpLQfdo+eZ7LlvQS
GvBXhy3RPlb9SbIj6tRoE6sVHx+39emIBpXmKjdfxmJOoXORXpwNI4mCkPmF9sd7OmjhjzqmNX7K
kPpKWZx73VFlSNmHGo8MxnBzGQi0hhqogXP0MA+nriQQI9RQfQcaQb4szF2Nrag+5WWhHnVRVcVK
smysCXfSrk97rw4Wc+nn9U2lYEU7x1GywpSwOtbLd76m6XLIHOJnL5KO7bYiWJYJLf39VIgmDuoM
J3A3eKVNolSOrVXcw4Ik6xUgxpvDaxawZKAp2Qcx0t2XTtGG1RoD9ZsqzrMxoIIRmwyMrHcNrXw5
xa/axvYiOZQhTRBowomC2K9eUKm65IR5gIcjIh0yj0J3qLHxyae3jN25UUzXzWsb/GLKGg8vMADx
hsXMvagpt4/YwuLYFYT4rcBI+JNsgXYL/OYfjFDOGs+Lcvz0K//LKimoxDKfzTM3KzZSTi0wCt9U
AMyqs5YaMJ27gwzbK1/XOpPNvIksPRFqzSYskyUP+SvGlAwuFJVgoYj0r9w5HHQd/uiDMF/810+n
ONNM3G6Q4+fpTbQ8wzw/M4l5CP7sg96nEcmfmH+jWgVcmuonYXoLE+09pmCAjh9Mke78VM3rIHmT
jDT/6tRvdelsZSodqKy5Hba4CXP+VgZcaVrrCFv8UT87zyFKI14D5q/bbb6U9FY9oViUtLwEndPa
s5rxMlS8Sd5ZpJPIDsGBO+Qu5k48iptJY+9mh6XeH05ux2BKyz6/jMGjv0VRMCOYIxB56sSqX4cq
38Umvq6WqRL7oM8zOYt1OTKOUNdQZl/QR8q32Wno5KLP9LhWQedLDxmYXy06mu+5SX5NLhBz/DXT
srWBoKYXLm62gSIoDUqc/CDAAfffa6Tv9dEn+ee2KAHyvU1vtY/jITh5UjWBsml1LMwdNWMyqT+B
dHa5j2N9nh8AsBooi3e/I/gPJ9YI9bkoBDcGMF4iC3k2CxuhR1Blch+rqzT8ACeQgcG/e0nYD0Ov
G3LZcJPhrjeDGZvwaAWU1nMMMYvWopGefHFS6f1qeEhDfaFdUVJPwHOItMdDm8mgO3ctw/vmayMB
gd1+kQbVWsLu3wpJp2ntQFCtSpMPLooE6zO93WbjLCRKGSURHz+O8gqwoXBKGjauZUIIUn/cn9Pt
33fdeXX8VQ03ADVDXf4+K3k0FXY2/2ygMbUMP2zxCNqq6/R2GGZHO+EUMsRTebvV1rEpR/xky1zu
j61/RbGbfKWni4ubjVsiBtWU4WUiZNDZePLqBzW4V1r9jlIje4fMQ+bKX4BXMm/mM14k7fw+LmTy
4GWSmKNcXKOJx9RAqnkLV7W6cnu0NCaA8nHlXsLrOlS2Bz5qiJVYQAfcDhlfVserv+v1SD6BNw8/
daGb0CZsCNIubUDNKNqG/POmuG7ZTG0239p6EYPPVV6Tz9w/jRXfw4yqByuOh0SgHFQFywBZHRFD
KJ6G80Qr/Xfrx2sl5c2v4I8cKvF7gAoOdcLtOJLq4OY0bnu6WS2xbjaD6RiYKQvtUh4mVkmH0YFh
QrnOrEbKMJMWMod1d7liIZdtFh5RmB5zEW+TTO1gWbnreKv8P+Llq1b8Wx7CW5UW+xgA4hY36NSQ
J/6JWE/w7widPifVINRHs2FXxEfzkWsFKS0kno/MYWBkpfmrZV5uk8cW8LSdxZa0vqKe5BVuI18d
FUslTYCW0nr0CrDjDnSswMvTvQT8+ECQ4SylaA5ksUaIINwLKjDqP5mXnB3qlp0C55NMbmzil6Wk
JLV1bKpzR12XH3H47EdtkS+fzJoFq8rL3loNgwg1JOqSNr0cdh+cNVtwqiOkNLJIisjTdAkSvhUS
35nNJzkneqSI4O2nsxkOm5QHIjmWcfQNOemRGvhxj6HW0QywC4UN/PVDui7Jo1cbFQJUIxJih6Yz
C71OIF7+5CndkD+tPdRwAJPlYjiCOV3jCnGvwLN23iechJE7qv0588FsKrQl2IoI/7Q5L6Em/Ify
zB83dnj2nMJE7Pn9+5MV8IcwDy8E6/cQqaRyStyodgQ+nHQhE7ZibiImcSzhMAK71HhkalVx4PnF
tK8Xe7cWsjYeHG1GCUlcj/+24aXMWy/vGsVfRirVOEOv7py3Xegeckef0/rcis5aTYoO7JIK7kFA
wz3VsoWGk/f6pib2lfEviKo/qVwVcLtLGvA2CKfzhcfx4msRp2X6IGFSxldb+8VhiKNlGFN7YvMF
vAbhGBfuG9MVMS6ubEc/B4FJRMer8eo/2vtXQGD0MwFxb1Z2xxhC+U04vmuIzFGYZPGeB0K23rOi
4XquPBsQlo4VQKVLXuUK/flsNg+ipaEVbW0juP6Nuw6MlyAvipZAtl9Bfic2UQP1oHfFVvH4NYa1
0sntUwXMoVrMBI2yo/nnza+aQl15zpR/3O7KmodbS1bKrxZHB44ap7Jzil99KL4CfUYmtGRae1z/
5c/9e8M+vz1ncWKl5kVELB2cYaHYUJ+rzMQn69L0xFVeke3Ibpv2J2FvGgDHBOvT50UxkHQHnL8t
C9vi9k+qFJSn6oC7/Z/XH8g9BhiGgco6zWpp+nYl/810vTvgTpe2yms07OoXt+Rj18Z6MMXrl/Qr
moZMSh+emDfXCewXM0h5mEBjM2qtEAo0d4r1iWi52CARnPaVIYW8YoLzMJ6HgwTQIgrzwR2X2jWU
5AidXjb4XbmTjRFdqQJrkNAl1RbK+H6oSWWUHrX4gzdfyrem8oHbbGJeiQMmER6uK571Pc07+gWH
PwzL9fAzQ2LrZPgqllQLh6POmOsnw9OoQF87VinvAox36wMEKIZ1mo+33EHVm2SJoMc2U7d0kom2
avFEnjpDbrIJov6QMfgtcpcmlrZcu40eWjJ8C1GUf2FNo8nulajQgRE8RbaxVE1r+xIlauXWEkLx
yMJx0ZqO9uvc7BCU1EiHw3XcCF8uA7kO7Bt1sRP55hVb/nl5Z4BXlkqH4+g/yYPfGcCED+BMRzEg
TpHUJ+X+vNiiYq4iPLHg3Yvht+qU00zbH2lMgQB7MRz+M/UGIC85GueyJCi1PdMdFC7FFBoJNr8T
NIGnoPgDPofxaJKAj9hDvYVzOKR4OKry6oCzc4fDbh2lqjOBTFFEVb9pZFzTR5yjZYFPvJUxSWel
AFEMO9gsmDcJdQN832mS0RoEew7n8xdDoYHspx5EMR7ax/QzKFzPSs0It4uw8v6E770GvSZ9Y+ps
cWZ7mxg/c0Ybu+VWKpfNLHmus8Gtz5J1TtqfwtiGS1ZDOHSVTdC/Patlz9+9OxfIQwqNEJqsdUd7
7uEfAMLa49E/+c8KR+iI1FGe2c74sZIzQ0Me7XTFPrEAmbbLjpzpdI34w/EfhqNTONkZCyiUZhec
np/4BhimNAyddB7dupkRUhqR8u/gRzk4TtMbFJzF9wz8OnEQF0YbF/fcr8GXRxYvyhE5H0seOcK0
B1w102PaWEF6imlgvdLtWLLJ/rdF0gs2E0yheBmRq5Yr+E6pz0psi/gJoJFnpK9Te9NxZzRGyG9W
IOJ6NGDk4QtbAchmbaRb/EcdfSYAq70zt/dIwl/LCXn1d3vFV4cmuY1LLsG9cLzNIFwY0R9EmpIn
3VLdTjos6yGZWtiR8tk6iRbYXr5QZSaB1X4PzKUe083/J4AO3qX+F2QWyiW+nbAPyNdXZ+IxZhRk
gglgUPJfbItC2fnytyqRUGZODQBhvqqJsFY1xmMHjY6qzcwxziXT05RYGei+RQMiTsQ75Ywg1Nsb
eewMbj+VL7efa6LrtNUFuCL8677JgE94O5m9olWn+9t68QAtuyO8jhsTlDMhe0lGyQVwmosNyx5r
WpEBjLytjKe814YGSRhX95nmccpUMv6FVPh+gvUn20MAQvvs2fQoCtLFZarkeFvBcEHYKio9lPI5
R7wfgBvIjDhnEIdtTiESGeFy7E9k201ea11gAmEfmCZ2cQx/yp8/6VtVqlU0Sess9kzq+yxO2Cjy
Og76qGAoV3yIFFOxjF9lL8EECn0SlN9F5iqaDiYrtEET+B7U3Z+hXJEqQsf/hKK9BBfw4Gu+9qjP
2nNmwl4DGmngDnLaNJF2onTuraojAC7fzVpJMQSdRqjFu+KKwoYTh8rJdA3YF0pqkuazuiAhayVi
e5HR/0YNpTyBxaw2xx29eJYWcRvDTb7DjVPYyW9ziupKsO3C0NO+fHZKbhlXz89RQ7V+76ZnsYw7
9J7f5suAWnXbjriR7FvLbgFctLsaeJAzjIT0QiMShDwHN1/0G4IApBvww7YVRB5LtrUxEagDYth6
OUOaj6wQ7omYcoq7IiolTShD1dp3FDUDiGjJn0CvCAkzr//Vx0ypxg7oDSa1oqSLTzH2iBgJt09+
uAGY8GTodTJJ1Q0NHDiPDysUF7zaNkGWsU3lYUJUzIam98le+gGwTxMUi2XigKeaCr0NpV5SvW1G
H6WAciEtcm+oqf6+hYRNJR5KWBuCUYbE+V2Czvx2un2EryGubnwZmActy+ZB7xHgl8KlxXXMxjja
r1nHRn7D78R2qrmEJ2ngrRzuU2GhB57vz+YgUx4D3WBT9zg/9oqq7xivhABufNuCDNI/7F+oBc4/
/uyeEkyrG0eYUoFFZAn9aroTISdNcRpvZMLIGyeqly1jZx5J9B4D5kEzgM3Lwy0/aeoOnYhuomBy
LywmO0gUV8T/rCMZ2pmQlICXdTeCQYdS3xMvz4SlRGRB4pPalw50OHJO2A4F5tVq6A/QsNu4JwwA
Df8qY0cLYYvwXj/mJZSZWgWWLaqRhfNHOeT9OC/V3f+4+PXIoYIcOWXLPPIsqwflVYHFqkIb7Iz9
wKqGVMo9R7ADFKPusNojenaKq1HQ/hAzO+KopYzcitBJBY3IrebjZ4EA9RmEj1cTBFDaNTFg5QsJ
BNd0DX4SOdWkAk/KrG+zDZAwwGtgKcD4rWwzfRJZqljhzMhZqXX6X1FY1xRWfQms9kS6mX/boG/Z
OC09mMIjgUElxftG66t4Y4q6yLpZcSEbs3HtwzCx4acXQ1reWWMAwnksHIxBBVuwb0JtNXPyO3ks
wjqkaOlt70Jtk8I21ZIkLkgryktiythAMNnSbaTw73s1YP+CtO9lGEUH6TrO1NFdmmQZIoTd8x76
fiQ3A7iGn7SmtxgqtcY9buGnBEHTb1Iel8Lt8BP1ZIfe8oGSDhlfB09Yl2cK0PPe1Oy53nt+Fhxy
b41O9t/Be6EvhCQNikKCk+ZZfjcD3VTVyrnuQpK+715UuAjkVU3pF2rQ0Q8Y1ye4Pkn4H9FfuhRE
GCrDO50xpbqYvXZBiGjObBmqH+yBiUv1LQriOXH8pR6QjmU0mPfXXOxj8pR2BFUHjG7klO0BWoly
wYCLiVo9z3xibX9Wpbjupj4retOrQLA6SNMu/XfMUQ66drksxIni0+ojcEFZF/81EIkeOyOy8HsT
lXkUxeXCQV90P1f5zrFAVtJ87Cit+fegOTYHK0SuA7VuOSqFrr4h7+mjK2jwmI8Xn7ma2Q9y8Q9m
4BAvUxHH7ZFtwfkdv74JG8bXAAFtKZGwRsvyk3vcYVSbibKBU6qtxtCqTQcGBdB0T2/CDVX4ViWd
+vqdY1C1TdxpkXPTgGJ2Iznayp1fd2V5YpvI36aEE2KkxqB2WSbRPT0S9lijafB3Bf0K/1W7E1q4
+9kxekQvel5IlkSBtFeqpj8cw+am/omndZ2Q5Q1yHQjTkrHcHRAfO86Fad3XT0F6yqn2qQt0rh3l
2Iz/4XlGaD7D745/Xg8Ib6jhGnRxAHGNVeCu2X3Ero1Vbep5iBsNhNOejwnk8PCRmpyncch08IqK
KU8awFPErufmhaKWN1KL1nxYF1iHBiWeAnAvaUnMaorSiWShgm7lKUnXBi63+jRJxVKjqMeK7xgU
Fdrnrdo7QGUkp6ATeyG5+k0yO9fTqimMd70UDZOTy7j++LI0p/paYiIVzMHuRV1NsSksZWCkrhMy
V+z6HD87uP5nIsMmelefr8wlkdnnWTsoptjJjOJ8bpxkPEKr3c3hWZaWbTGjO0zC7YmGS+aYxCy1
xDZ+Cmv78dS+AXfKaH3MontifCnIIWI3rQ24j5ESXuGMhMoK4aRtSAlFCooqFqD3QBjpXCcb/2Rq
82es7I0GVxQQFfBApK3AGz0ybxvJTMJbVx/PwieXXQLeOmFdNROhsUQaYwkLcNCifxKYqb8ZXZlS
NPSHkMG9hpwG3Tf7yzniLUirBFdB9Pl1AMKC0Jv3zC/L3K88EHugo2iURXJczbQJ5q2lqWzNkfYK
iDhaPTWfUcApkCJwKgC0OWppH2q/ZIYGBUzJTpUDE0rGMVJuOx/UTAaCnalZr/K/wzheJ32rTneF
f1OzAPsBM2+AvI9QJxDM+0MKCAqQi4L6fDTfKToVKDKJaF+GWdlcELVyWIbi84Qyv6UWpUGZ7ZCV
1IuLYsi6Po4bRzwbDlR6q3CmP469YQp/l8lDunjuDQMImyJlP0JdECKA7JdYK6tjGW4GyGH5f1Jg
oUNaKt6Ls8bHPT2NyunPnpJo5eoreTbkNRdZwWR6vZVnuNKqArpGhhdsOhLzWhP31DJV9P8AGopn
L1NWc0J0ES96/5WXO6klAZAsJijNOZI15hm1cj0qAr9Eq1YNEnT+VoAHpwt97PG2Y5JhtdL8OwsC
5it0OCgBAsOEilpweDscW93sHbk6r5OTIPm23vMR+y1tH8G9yHM31L9gQwGdiMcX8ZyTWOFUbhe6
1zGG5weumD/rb1u1Bxe8oXnEEdGeLcRe3BwxrsjDFQ6917iMkRDk7yWz/U5p+4SSSc9v6jYZYwTw
4YNl64DvNE05NyJlKw9bdfPU0bSbLCILxsz/fmUBkfDHQXkZVYLQiPMsvmF8bHc8lwvItjU9/9bk
8kNHt5Z7Mo+uhJ7yA3SdTP4xongRAmIxG/Go7If8uYtkuFT89dkmKOMTkOHOrJNwPxjV+JTDFrrc
18Vqe7lHxD8027hznBwUBE4b/LLiKnNTLW93aOzj92zIgCyWcYxcVQl0zFCsDaoxjh7c+Q/6Wfp2
dHBh5QRQTDGoI5AEjz04qv80EEvqRtG8NBal3Jd+I9+lhw3B+q5WSBLlvqqNyZh+Z2R3cagfv3Yu
xUoLseYDMsvzAoD9+Weq9304LVYNxeZRPVdbr2jvZ4WWYrwWMibS+QHMLhYx5Q/j6OFbTWnh5uar
OyeZ3T3utS32BE+ZgN39TcXHE5ngjmViIVV1X7PlRzdE2+owtc2HxiP3t5joHekbovuKf7tDoxRC
WM/K2PLG5oUOPGUX/ec1+/xmOwHFeGyUPZyRO2haZ9iwWpO/r87gIkdHVsYbsreayU7X70+p4bxa
gJcQ9Pq5O8K1tCaCOAXxqLW908CyKs0LTlykuhUmZ/lE4rrnJB0zx84SqCga90QBFtdSF9oMwFOb
2lrzlpXTFcJ058t/ZzJYiJ+FTZEZMDCdQcq8CqYrCGewAhG/SCkO+xrCczo9WYAjj855b7TuSazn
U9rAtIj92SzXg9W8vlvDgVmu54AdlQff13dn+GnvtMu+0fc72LquT5f0YIB/Tv3t6inY79rJcDzC
AsD/dPwR8jAv44DnQKLeg+zUCzD6wr+08YDkDCNPiwD1PDfPK5MUEX7Uc8ZNK/9Vi6GRko8nlqtO
UQhtu0csbrZ0+hXQufoauOUQOg2SblwqZxhUB603D/7nXTXmQcAsfX71fj20FTEGBfPCillBW58v
SyamIsfdyv28pWNZi0X7qExCsccpjMkI9qRhyIn1bzqXq42B09IHBeEYkw0LG9UafQHF+MbxMCDy
tavdRcIggD7MWEc5eTRYQeKEWj9e+6Z1y8aeJMgQF9O3VK/wfT+s3UXX/fUNC12mmTLJwBmMHtCT
UvV08BEmR7gHyRaXNPxr1HDgkt01Ytrnd2H65UjPdS5vNCEgFcPtGch5FMvc4mQsiIuCYJreI3Et
j4pQVQbvfPOYgcdyzOGZKTr0B7qorjV830/IJZeX0vOCXb4oFJOZu0f8VK5LtpFSkuJKuE96as7u
Wci5AqdgzDCkqC33w2du0dbYxXueyqJXQgC78hIdrYnOgwdKZbF3NkkREwmbPrT15HCdOCUvP88d
CktFdMFLgldiB61I9QV19gK9WqwRODhoqpG3u+dRIbaPTuNH3pBfr1oYJNQ2A9YPgPxnLUGz+332
vXzqGTFuRJtjR/ngoEl7CuA28KKAeTSZLAyXGcKLz5Erd0aMOS4klSN1TdICUoRbjanJexmqIce5
0CiUdssfE6r8wFLFsmsFIScLWAOeTosSx2VuiRsPbh2q1JNSO5IjwGXPyq+1zMuf2U+EP2gUFIyd
Z9ezhMYMvP2DW0Q19CYpdg0nbH02GU4tANOton4qNtWsEnmmPdN5J8wyVbo8RH43E0JVDIuS1g7K
PQruTzydyld3N83fm9goaPS4LO0I2T7MNul6Tjxsf2ZbbEhnmsa2yNaxdMbTcaNt71a7NxYituHa
IqAQJzm5fvvXhOoPNxvH0wfjykgvndmLQ2uG+IP8ZKn3IXcX6L107nCRsVaLSG8l+pfduGqmM+GG
G7VcaMOh3xC5yqYnH2B/TIXeCgIAsdItYD7vuZBQ1VkPeaaykUKZkVHzlnRJ0y9+TuNpDqo9CGT6
aTIT9H1MhDrMlNWSTK+TIiR7BMgeFS4rHiKiIOLmR8G8LMKMgwVLFtFFrac5qrhR7pnz0HAeNyP1
3Ni3UtvEeT6RN71EVsBo0acaW2nLCsibQIMvZKAl5KY/b7MtlSyiuZxaM3hftDZqQMPc9icnoQN9
IHeWFLna1ANPV2unr78450xCFNGR7t5sPrrsRvpeP4lgKkLqJN9pp4SteDGNmFB0RrmSbDSan8Q5
bzKiXNQaTY4dpkTe5Opi8DP3Z7gw3UZMA+i4RxkZavVMDpGBdkXmxFrwJQeHlHuM0/dBCb/PALqO
zyYbPS9/MFGYqsrKUGo5S4/NxGEvP9965qdWENZJonsJlC/8as8glqUq7lJSgSjKrTB6qvVsK5b5
vzFNw6b91zaPmMgEnRiX14Ne63pCAftcv9mlnnlmlm6JlyEzulcofQvSvkVLrRy4BL5B6NFkoQtC
7gS6aGSJaQ8zlWBYmm6Kry7RrZr/Psszv5JJJWsDeaYhOKAkNGBm0Zm787JIPml1WeoO7HhhEPjk
Uy+UyXu26H6Mk9z37tTZCfh97BsRfvmQTrRUOIJxBElMC48Aqu7pkG8lG+Pk5AExwi3fNBvZRsfP
xt3D6EjGV5W7Xmy3U2YT6koxAgsjuS1mcQb3Xbz6jcQK03iUDQfX38QGfFrodK6698IK+/jXEl4z
S0h0S6+cVNVExOgjHHAgrk4SjO9ME5jPbobPMWqHHHxthMEWD55cwwN1Gzn+z2FBs4NGr/FI4bY4
FVZSIm8BJrXsljyxlKELuoUR/X1dGUI6zgyKg+Q1eTQOZfUL1klrD8AgOBhCPrOm+pdL6mwscYRT
8lqDv5MPsPqlsIclOjJa0jSoXsJD8pH8b7yVDzZOyoucHyWy6/vTH6gEvtsXmh5QfyFBdk7fWj0W
dKPbLXY6CvHHNUXf1k/JeHul/OL9PVB2AnL1Mvv5EPADzqHbtc14px8AEL007aO4Wbofeyw5VCC9
6CpCTduzbWpltEc1dIAopYsjymSMXvEim7NsOJd1S9+M/4mWkf4lWflKwV3YDhU/EOPhMyQZde0v
NzR+MPXqSwJLn2f6n7RGIfuWytlClOg8CP37EMejaXGTBJhvirb5FZ+wcpehgaDvth2hUMss6yGL
hhA0hP6TqTWiTpPKHbLGMlHfr7navLZC+YsbYOfXyL9UGsjymCGRUkk0IpZDZZI6pSKmeTfRNt8h
YWH1FmdCEX3gLeNWYdTfRTxlO2Rce4/2q7IoRCR/4oKwkfyaLV8Z1dxnWvl1Ohnsh6B7umTRnEnW
uHIVWpti2jJYWMw9WK1ScP5xaBWdPleMssOEsfX/UH7wHGRb0AN7ysObg960duZaFQyrE/zRyy3c
kGixK2+aB+TmFShOhCkiHG8utVw5F1FFDabyR1L6E1HhxHqqwNXJbZkFjDrdzRsY+LAjFRYIxfbe
7pRBvUNFxgps8dAjUbAyodYLtTndc/Bky5S4O9GEuueJcwxOu2UtsD+QRR4IokD2eaK8tqZiHcBK
Rhg1+MVsBF8TTyjWhS+QQ3n9dD5AZuINcQZJka6e/k2BvwJNLJSyHYai1+BGtmaeIt8kTtrYH/I3
pge1/nPrfqCNz86Pr+FiIK1nLyX/lO66+qgQkn8BNt5i6FoefpMx3HwXZXnC0hLVr2t352mimzMR
ipU2wi73jtO+VGi68evU0ufOoU9V9EyeUOxhjBA/lKR+e3Fjxu1SsZf5ehH0jXUWxb3L9nMhf0lE
BeR4ZMwCMmjMjSNuF/iXFaUUveCv+Hsot3wHDrxDTMSGGyzcHtJqg+paVAf7873GELSkUj0+jsws
+SJaN0QjSt1Ljrpys6+YojpBHdJURZbRXLxaQDWRUaleNNjy1Uf29ObZBs/WwQqOAqvJN00LE5y3
JupOAyUFJ/mt7fbuCDLZYzRXbnBRoKV1Ib4TZFmrkIbcGPlGonykenSMHuEiOCWGaQDW3eispN6k
gRUcx8t2gd9hikS6Nh5C3cE5nggVL8gZ0Bj9kMC5E9kbBlmHElAbS464dtCCCdawmqjF80zopyZ6
9wkvo/a7FqFfoVRy5mSc/h1GeP2eeLMLFerds2DHC3xXnQkfRsJPQ7EKD4l4g6IurzOQnSf0BYZJ
MIokHdliNihPMwPtt0cGi35VJ9nNwyTFvQvGJWaRbjRbqGappA5qPKXqFpkzHFdKOpJpT6hewkgP
qv5vY9MsCNRDIFiFozra/ZLNJjMUx+y+HOU3i2CqlpnC4u3P3SBbwrINPx72QfxGUz91/D4wUKIp
jnMAFqgH87lKsB7tzLUHI5SMpuSwEpMYQNfmYvkakm0u6+ibnVPtmfDhF7MK3wcOy5vxdq9FjQln
2varoj6OYCUEC6/qtZ49A0aavrD5DS/3K7I7cpuKoqEE2joX4NTH+5CyM+obxWOOzEOySXTqMXUH
/zk7h+1lfQDPyRBKP0If7JqgV4IDfT8kzXqFAKAhif3cNeAEymvp2vnnbfNOISTIy9H87LQnglkk
71aShFFECNFKRxJoPZ2NoveXyHyeRHMBXpqEiqQf9MpxDhRR2lRsMjWMfvR0m18V36AcFlgqHdic
1bZ/88GYTVQkjxBencNeE2Ng3s7TFu0d0VWA9/+knrNXMoOXjlcT6tzxuxJfWrs8x7yYyO1vEoZg
SiViJZFRP3kLYjCx0ntiCC09m9dgUfWIEWXrVeHUyFgEmAeIsM6wVph2BGtk8c891dlF5qZxnWc6
5Vei7c0IzUaWZLIKtITbNEjZatbl06RuN20ABrNpNoKc48ju325HWcXbcrRF7EWEjoaT2UhinV/C
dcGYRqK5kZLnkaCvjRpM/sLbAcesOSHrXToK/F4vffIsdUcGLhoGkIIVKcOL7GZVpM7qgAVgdNKZ
HLKX98qX+7HRJyfULoq0WGXVoHMjoBRrAKUKGi6b178UtxLmuXipof30INZZVNTQfRm3ziN7ruRU
YyO9TvhumbuMRCP3nDyXteCxWv9GFk4YQ+RVeuAhWVyhcbnXbBnX5k6xYyQyCbyH0QjvEjdRghqP
m4OsdUYnQM5w/txnQZ2v2AgJ/oLQZHCWfXNVyagPnbceLaq1e327ueNGazY3iMjgblAPwWLaH/hp
ovsJEXWZPPlkMaMudXGAC73QhJftO5E2l8usKLvKCHlrOnMDez1HMoMIeiqmQEvQGA4sO3KRC6/n
HT0weWuZpveZov7YXDB0ZaVtl+XdGHV9ysJMityS2o4jNxRd8vXjRB7GdScK0ohBCgEnOIY0FTt3
zoDvss6HWsPJmNlCl9l7+rdpghqw6tH6RDyOTX/ffarYxR9mcDcDHT+6jMvWzDJYicYgBga4kzBm
16V53vZ4oTnCZl1owY3ZcpyKaBRKAbHZvfJgDuQf7Z01erILjW4CjgBSnJotfWNjy4RK40CPkgue
0n/ALbI+ZUkNepc9fpCpSLFzaIbeU+hBoTRi2HVtw19pHI/GKO4tiHZmpGyUbgccfWjX06HjcRJI
R44+777MxvKVrUEHBLUpNUV7b1YxbYb00M5sEXy5PalqG4eH8hGnTGlRgJoFoygxco5jstdMX8HL
JDBy2ystLDf4H6RiaeEoEk0ANtZUVtwpYNeb0uOaaqGLEmibbdtTxIzDWuKRPWKXROk39gRSi8mh
vwcUV7acQP2o0rQ1zj9JNoBjdlPYasYirlQwXjgbX5+LHX/9sUDOaWrBYtunetCqQtYzfrQbKaXp
TKsU/OW85/EOXTF+H8SQuD5YzLPItHTTqRsn1FOFaKhcctI3A+NF2njcd8A1vaAXFtaNdfRT7FPB
8BGtV7fWtW+boL3GvjW6g9fRoAW+6yOoOggiFYlJeSi7oovMKZQkjcYXggj17hxAPPJstjtkyrL7
fWQNgaAC9kQFvXlkFT2cm8VIGu1QId23LJgSaXNgrak6vLg2kQF+klU0X+a5kPJO7VNAbQcadwUo
nYCCCElE/vNtaWVqKps9TwfgBn5uJiMGo+695CNyH1+yqyixem4IVFjvy+nrk29CIczCieP+ieFI
pJ9ZrmOuxoZUK0oR+OK1gRiANspgJjgCN6Adl5Rudi0bVbgCoSnhWS/Y0ho3ROUJS/3jd3FAQ/Vc
QyDQqxzr5URPMwmCXkC5rITofPWu5kFS50UMdqGdvz+aBEduMsMbSyUcT1Wv0903jVkhdCSOyarm
vxrqEP5tbdZFFAeqblH3stXSeiPIYYQMCj+BuTKgqhnU0nc21UKXbUW6TvmzhzQAr6SSRl6Te++E
2SWj8autLxgoB5kMQYK1nmWqCZGbLULRTN8mcs/prPchtqE43AFWdCG9rYZ4NeaBZuhuamRYSMDb
+16mpPNZb4s/lDtFWQPsDxZX/MJRvRgX4b1AAq6uxxD4648nkW+obeG96Fnv9374jRMp770yqmgh
sdlcOEOvaFNPcVr7zOUhMj2kegK3cBolNz7FYx4+WOnMCThoEoQKAFdiNQI1Ml+72RV+PyCnGz9F
VenSSJ8TAitq0UYu5ZhMtwiXXEKjpIeoZaknpAuKY1fd26aLjdEOBfxC80Jsc9ZGt2BO/y9SXh3p
UTVwNiNPKtXedSt+iKStDzct9bHULnyvf1+uU4tGEx+HM+10960suy+pBPnGPJmRstvKin7ZqZK+
hXG43EsLsS7Bk6jdFkAilQKlFBBhQo5FHVQX8QLi/I/jnBgT1yDFJUEgOfz1Khi5Fz7oBN/Ktrgw
rBjkR0zvSFuxuzE3JDqzZn7FdoTEW2k7Qj7Ae3u+mwE7Tk63lKF0HNjLPjpX1hxoJzIfgEGuTfrG
uSCWPkVB2Q3FHJaqU4MBQbsy2OkNWil1MR2in/pDgMfTqyY11JumTpv+v3Uln/uOmClYkP95DNJx
uWFgCyHSUjKnkrT7JFIH8QGe2096Gl0nS+h78baJTaGAucU9/v3uk+x2+A43pB4biYexZOt1t1PC
WnRw7QOkEg3R2M252w5aQy5F39TOSzmv0b4MdnksPCt7oer9TNAWVDXTjK+OktI9kXb951hlIHzm
NA+8vX7x1kldSB022TLwmNNob5mn/jBwAp3vortE9VraHxEYXGKbHH0GKFokm+VmYk7sOP91v48i
yiIzX8WBsEYQXgoOtOULuVBPXGQEKACj8HIHOVMl8cBBMjLMv1gllUkslUT10PnjO8kpHceE93Wk
ZqcRqzoW4MGoK1ii9uEuRoS3z7jdVyX+/6mpIAvM/YXAoDlchGo5X81R5NvVYtvuW9Ea1M0XEGgd
zbskkwRAOhHUGeRII5KEO36RzCmKOiRW6W0veaaeHYOLh0zc4go0by/EZOleMYqLDKXnfIfL93+n
MmmlZDJIdPlkDZWWGYFrAXr/Vb4waubq9DOlYjnp6UjP54OBLJEzR532+p/6HSbzUjKYxhXqwuiq
RhPR7AyZVP9e8s08lhcSPRaRWRmGE6ipyxW4iLpKeedX4/JI61pY3BN081vP183W/l4b/5MpktI2
w4QI2DvYLra5n1Nox4PbiH+Z08vXDYxg3/Uoy8F/30cAME8+wJRLo+Qeu5a5DL43gqfk1NygYa/9
Hi/KvHjmqb2PWEx51zqbHJB1AyQm1zGakbn/NSb64/+7VosHii8hvTL8A1dXG8HqComsr5ob7K6F
GR6QMh7ePqcrnWqeGXv/aMDfYXrr+jqWCmgqupWnVKH7g0X+aEgW2KTnjxRuaYqI4Yx7KT2ITBlE
sxd5BCCPI/RUekVpPoeDPRY0Ficth97cck7PVi5Kew2coUcrZ/NsKBvPJqTsx+1bN7vayxVfmhZe
qVCSKNhM7sXmNWJrplpE4MOkWP2SAjx6qChT3/nvrSUbxoAgaosOHBu+no0Ip8x2qmxTCvgi9hv5
iaC8zjyx1EdNaF6ZklJhgrDSysLEXAAUnyUad+fPByj0B9kclnGGSZYwiYx4WIU1IJQtIciJM6G9
XqjcIlGIKpSR+i+KqGqe4FUdTesjjSqneZLl6nM5HuDOMx0SDulTc9VrnrQLbFOqbTTDPV9N98y+
bdqyumgRvgmfwdgWGBiHnCBgfD5ZKhqBmCSIQDFSHr9H5LyjX10R/pd1DEofxMjS9+igTovaGs/Z
Wel1VMZxn1DWQAVKZJ0XscnD0Bv7ONv4YmyONw1kFAsy9EBGzfDSBgBMqlGF3gNxhTvi3T47dgJs
N+zG33lnzUsGlkncdYwd8cWOQY8hlQqol+5pLB3ycAu6eUFVfLijZ2XXSUQEyBdG4Dc0bT3dM+NV
kwQWdaHKvdgbQOQ0sS/8KQD2UpI8JaCqI8uMfc/CkQaioIpgAXVo3z+tn+pxza3SFYPGwyhxsWzR
VX3T2pewFdlX9xPZ5V136i2CqiTvbC7jmK1XqtJkazFTVTOY6z3rx6Hcv9WGELSISJ/5sMU8ygqO
iiQuQGz5LtU9Hq3pjsYG2B7MWxQ4xh8xNQwMNKrH0GVoA3B8dZ+c0M85zidO7xnhcqPhWXfobXnV
dR9qb90ZKFTMPhnd+l1OFrgRL2TIhxWMLeJ3cKnL/xwhIu2nTvNci35pSauklBwxYbwCEnr2N7l3
AeniJJi0Gdyi9V6cu/A6O1mITpIzQEFPcC55R3/thgteCNihd9+q4wqNWKvveX1d9gR3fXSd4FNB
1nBUCNc5lKoVxL3tZJVrLj+M/txul1rWqLOx/IyxnQRPsGBkQ4i2t3PBJVm/2Z0YM0ol4hbE0S/H
vVNZF61vK3J8Z/z5ESR09a/P7h1eGHbZImfcJ04sCtVnqRPsSNzB/2SB595YjLySgar2YvHBawgu
vpBdEeKyrFsS43RF+KXeWdn7o50iK+MOKxrecceKqZFANX0vcfjHOR5b+rE1Y/IXKNo2cn9xkIrm
GnOPptgZaRPWKVcPxVZBpmGC6kkmckEZqfclhgdbvHHIli5MfycEQVWbAUys2diVYbh9f4Cwbrlr
yR1ss7a8ankWl3TK9cwebtngcXTG8894aTw8NmMVgX2tebIaY9oFSOebYGcbXKh5UXptcCuEZMw7
Zug5F5cJKFyuRr8JB+CpUs8xumb7W+VSIU+fAZ5TbRncAwE8TwembAwkUYajXSo3MIOWKswU1p6D
IJNIM+35AEohqPfyuDhHuZB1tl+c5ButmfeNqMFN2q+7qi9ERGfFVssFf3GlhZ5OzrbLZ1d2tf3R
xrHikL53qYcBe6GvdP8Qce53QxNflrrvIMHbYQ3xRky5kOuuqqgC2r1Q1YSymQNa4VTljbSw65AQ
MPG/BkWOBHm5R7Gxe3W/cLAAvgCXCY4uCamNaszyl0Qs74HoVL0YISI7pfXbzkxyKet/MOUE2fbs
yOMFRG5KqNr+imHg5C91nINKNgLSNDzy/q0WWMxnP0wJ8kiE3m+iia0nf+K6dj7+17IAJTz2b+Cq
+HlD07qJVyVLjlXI4d5n/ra56b6CCV8Nieyeo4SwXb6e9QjNbDYczQBCHxsp1AHMLmcUeTrkOxnG
23BG8HdVwAwigM+NVZNULRjBwMJXke5jaJ0PXu6kXDZoMqJjdBESYohSkhP+LrC/xTH4j7xPI4FA
POcoD2gOOjk8cphbvcypnNc6fzQINMEZBZkMFNzC+j8p1upxEUNrgi73wHHyWpYi9LRT/hx5fYyq
qEGkX6C1zyCvmdE6JUtYr20q5PKSAqIkYA0rxk4VI80RZlixdNLxN6ddidx8G2Wr50aIMGvt8fk9
fRtMqsEBKAgVH8lwbiw3EObKzsp9oNrRwrFDBAA7IhlJn3Y3wRbbhED/fMLldWbkzUnQ2JTKEahK
g8pQeZaLA+hetGyGBNqlzLAXKwAsFb67smyW1ARabOW8XLcUON3cg2mITrLOP2+0KWGaidht/Yv6
oraHGcP3817Ewov6CVYNFqfn9sOIihIPVocQv9k7LkAgB1kXQXcsrWBMW2TnKzi0XyguEo8bvTQD
nNWHYG91UCCHAL90u22UDpKFhSEYSi+6osjc60eckw/82XkEi5csxoxabYbNlsBWpV2Lqpv56AT7
DGDnLz6PSWkld5tMX4DuvUDNYya8ZuWjciTcNnLyt7O+B0evPx+6ujo6vR3+rBn7decV29++Ye/p
uc1o6zt10Nycq/OfT5WO988i/i70wpjrVo/YKeSSpgttNg+CvkTpE+PGj7/aOCrKZihF170yoEl/
CveN3AneVXSsz/164FwvuEU5FrTHqzYaZX4Tvf52+8OKVHvONdOkU5mVJs2oBoLNRUNxzt5J/3QO
vRrQV1iou3bamRkp7hCGGNrMQOeInC8Ee7OXlhhiEUBEYhM6RZLhGACmtz7bo2AG+lGNfaRFUGwk
VIs4Z6Ad4GujpUI3sl/b6fzYiJHCl1zymJ6kYYex9+d99AB6HJpBEyrMP1IZzc2cVxw7bV2Pc30B
kMQmztjPrH5ucFlr4Jn7S26/ty0EGZ3VGqRcOz35vqIpC5he4K5lwiifhDYJ4/Qz2iYvFewOVSk9
025s4LA0QC/lY7OGg459IMI02dEGAJJFeH0EfvV7HapuhPSH79H1+fQY90nwmsiVeVL+XTtHPx+B
PQgrLW4wpd0nsYovI/PlpNAfb8qqFN2v1lDqQJ29nKDagjO2qv/uLDsKIjIXWbvbU2C/O6p1+F5D
sEt4zfkDPH501K5sKEYp7OeTjk5s8CYadARvKzLTDywLlcR8ymyg/AbCwzpOwsOVcoIAjDxuIcTZ
bRAiBh/Hy+4U3p+3MuDYu4uA1kMmgi2+LnjwLaU39BfSv+tNdALAbXtA8r2NtYYqHWgsG/z0znkB
V75cvsuZOjdQVG8rxTVVzHtXDSprNbbffoGXUuVd06CJ5jUJvUDJp8N1XrkamNSKqJWVVHgTIxuW
0DGwR8KC3UqSPCAhSR1jSCg4AiqcdTovKpF1VtX3lPbHOFouhdlpMpodRtQyaayzmjOmOn3TBaRk
Zuazb/QTRtNLHZTyFQHa2Jdxq72cQAaoK7kY6U+aROzlrLGhK1LVouqSSZRyCSBJZL84W/nh1Imo
a4dbR6XHvpWmaX7fNEmReRI9f5O7i+RzldtbqXmBpQVCTpf6hdPI9NEU/LWRxlAqn3x+q9jWvHGL
0CesB/NFpAGP996AOJ3JO4R750haUZ0QvQOVOZpINTpopUKfwQL3NDS98qGcl9XAbNPW6M2wPrnK
wq7Nuc72VpOICKfa/DNT3AysF0GbmJNBlqY8GJrg/v1p+G3OZLzVa7yApaChOyouKdckGWCgvHNk
+tpkpXeE0Ad+b3ZuIypx0FFKJsZgTZSMK5yFE/RXnkP87ZElJcrR2GRZDopl8G4DuayAngA0YA9/
nPzNiHGJQNkwdsU7BGdACmLDUDBQfNNk/oDdsrpyPBWY6YDd1RFT1agR+IIc/zRpQb3VsfXO4Gj8
NR/PP09Q8AuU+8/4M4cG/HOqXop7RygONS4Kdw8HNYdYkyxF1oO0vH4B4yYBf1B6A55S0udQ0fFt
8DpHmGannQvSLW64dbZAbdFisneAoYGhNWpJ3z79qqfYzdifCTk6ksiwlpRqN1IiAuOSPZPi9OtG
XV41/dzP0EaJ9zX1veTX20BTRYmA/ekCLeYZw2YzVCxoColnMIKzbhlgXVS5gMQqECnWApKcZH85
nD+K33GV/0s40AGmHBsWmeJ37v28BC2rpE4msR5rwlZRORbD0/G7s2Du6ME9ivHVe387PRyydCjU
W50OMWhw68TdRaUM8nnvf8FdOVBXxc3XUGOIcruxjKMgnhVG6lSaWuUfO0DRvr6CbadL1O79JQus
3EZGYxkCA42Aw3FLjVJ88/xDJTEjdACLKJJD7LWivuZHYnfk4db1kLZpS+hgWRtupUFksFCAOjmS
BAJbhRLnSmh+/p1FZewc5+Qm6OhvBrQCOkisGJcBNrGfpHYEopXC9Div6sxDAfeGCmnEg9tlW9TX
vJfddU/JKzPbbAmzzgxNCA2T9q7Kykh6vaRe5lEUBfaaKnJOge4AGiC2o8X12lrVeTyHylSKqPZP
MlOX6n+67+OMPo/epcSOWQkSt+fbcL4zkfyztFn4yztBJRM4mExRkZ1Jnv0/hohjKzGuc0mddTs3
IBPgGgJv+PwFeUH8UVyApuFDaARStNHdXY2hg+Qn5+4jE0MBAvLIAByT6WGJc7mVau4lOCuDXZ1T
rRBOwOM46+61nChYli6teNw8Y2F5MSQi9/RrgyElB4EIPVHFryTXIycb2GYxTYDNiXobuh/V/8Vc
vcRwXzAy0YaIgGiypKMABXnufd+yKb4sJsrqyPgpvAhUI8SYqFeNC1m2SCkPyGYqTcpzQdIzmpS5
cwQCf26yr5lil8jvcolmjfEB8S4s9OAmWWiNs6mtEct6gAeYkpgtR5QIiMb5PFiyPaE0TH9o4Egc
JHSmqQ4hYcRQNuMP6HcKKBj3jFTFCtVtac2FPKtPBrWYUeV3kKAedWpVLYCyrNVnz9bsyOmnCc80
oUpS3Mi7lFpcPBlXn7YJuGbACtIl4M1rGuNXigY6qSVLpJH0gt/F1gni/uUdKNXbpJyitp8wDjaY
9YO2qhhtEcMNPTmHRIon1jQqCJdAGUeC4tmvg22yek3MWbT9ptg35UOpI2INj98K+qrGOdxCLPET
Bq2c31dgItah9WrfmA3lNkfEathiGkjPjYZYFWtudCsEztynC3g97x2MeG1fWaEAaXkceHgQvmBr
GEMlRZWbgebUduhfCwUC0LcQ91xgFR9hmaq6zIb+cfNfAiLrMfy51BL7Gp3DwJb3uifxWfhhGV4Y
/IXNd7UYzS6BWeV+uMXQyfk7s/s/kPq9mWlt1A4TKdnhzWTSmZ3Df4rMFp6tn5qkKfM6Occ7ZB7t
scKWx5R5ryY/gnaDuhJrTwk2My3SJ3ReVTyh+fI96SaV/Bin/8/foMXE5d2VK8zMh5hVu6yyRzex
BFs3SYxPmnoSoVNdRFsgB/BtsYGV/B7HHN5pE8tF2IQy+EeKSjJi1orqOFEKmaBgV7ZFvKeJqRu7
qVbpVEB5UiS/ZyLaY4GxYjTqyXqscF7KffpKTrz/ALJPGfLms08h/ZddWiD/h0pWXPuvsaR1Co1T
JAQ8Qn7yX6Buhh+iT8l3bu4CWeSH0L+2LEUhKh8VCKbiyI/pyC5UzEuD2yQYnFBpORASRUvaPhYN
gDSJQHtggGXg3HIRDVkkU7qjQXd5Ij1chFVMLm46cSmCKj7O4cXDDDRFMrZ01tdgD01R3cKXsFx9
jTKjXCkUWAQ5ob7CF009t8nZtNGwInncpkhzZ2Ofx15vy65u3fMYOEv4fnsdnVUmIRRzfih5QhR0
XWrn0Eh0oOrGFB6DcvDDt3SgUPFyCSqG4rggsxmp+Q2h5MQpJc/i1blm8rBRRzj3CnICBdisjaPr
wwf8j5HqQRw8KZtr9ZGxblymB5ptGqlAKRpytslnX3rGOgO+NrSv634eSlT0Z2obz+unI6d6yBGq
2X5ZzlNsaPCTM/ZryFfSixB6dcwl3TLHrdrDCS/KFERqCi3otxuk6xOWWpkePEt0utumH02k/glT
qPIDHgDADY90FO8e1dX8S0KdhHLT1PgKhSHHQS988XxrT0pIGnT73r+iais2cK55c6bRHYG/dhI7
5z4VCBua1g5V866B0MGSzYtkI6sqBlQ/868uHw9gHgh2BPkBFKZMKfB2ghA5+OSbwB8XnfTZs0XB
V5bYfyDhVWC9SJHmiJvVLlg1bkBKz7Eafd0vyGfDIwJkzHMs5QIlvIvRw+9xZuP4gXH751zXQS+5
t2W3qvXlHeBQCucd/7z0cMxwRifGcremMVOSzdiA8To2DiEpY+wQBLjGToFqPU7THh3T631lykJp
c5HerMcMt6qXhWO4NFkYG1txQ6QqC0tPOKuvdSD9wCPDfBMQlGDKJ9QBRUmNfOQa9lgNhcmELTxv
YH+MJyx77HZ3X/+OeF2S0k2boYfBWGIrorf17nJ44gmxzKRseAfMqqs0e75G3dZyVUUi2BRwElEX
KwyvxM2aHiUVoM90LTuM3IjBQzlahKCn0nQK5v2qTfFWgO2j8lNaaevVWlmqWyd4Qc2zluIXzTdV
NP/ZGPw1e0lsiu8L3wVK7v+cIjhiuk12Cjn2iPpEDYNYQJDW6BI5ecbDbb5IWOS6lqY1WXyPxE0K
sADl9teq1H2kO8IZ0M4UFpPLo2DrzU1S3V1RVA/ENFaUWhrAnP9k7axeysRor4xuKXdFwlcz6P0n
WhqmH12CR77yP6sppVYHe6OsYNgit6fEaEuhcnZchrFkN4JGoZifyPcXBoC//nMvtG2FH0cgBctt
xUnsB6AYH4KVHhsYb55YV1rSlg0PNiQCQPyERtOqDl5GDu3tJnEoZ2Cs1NiJN/iUu4wDtk2CtgSg
TpJDfLTnftQagbi/mpcpyoBr7eebky7uuN2hN/UD7HRUcM7Bj+yYTo0f298sd8bk3aW+DmyU257X
Ms3VhVgtVOrXWvm/RR/xlQM6zkm54BawR1IRN/SA1NFBk8rPuAzjZLp4UqRprEndsLzpu8WicDh0
/cmILjYB6DB/RGo14/mqYF6GL/afuSnIYxO8QsReZvbo1ags4PN9NhzS95Q3ZhfEF2ritbhXkoQO
ko+/4DK0s4xgx8phSLWUi7lAYF0d9t+QRbbOcOiQCGE2u62ml+qByWkrf5eRQZpL8dXeWw5H2T1l
WHj3Mpb+M5wLWQLlvb926BBHIxQWKQotMGAgwa9hyeDEqj3K0Qfv6n8P305pMGbBE21bX6GWwqhS
1PIR5hc13J6hG47BMNv3wjeqXc8aZVaLRwC+bU96MvV+j+8XW6+Ll8+WmmAHetrsNMnfPo/3zyIv
2OurPgK08WeEVY8mh7l1+moYO0k4/zxfmUqneA/4WeTvkx71vKN3/E+0nxIqk4oLNkAOwaHT5f8h
1z2jTM4DkHZxL18K7K5k6SLFO+MqS5vSreNzHryNA5ftM2nrvaRnPufNuIWxiQgISBIxZA28tuRe
NNSxGJ+nXvXw9KR4dn0wGUyKrXG9zq671aoa8YdCEwb9X57b55kPS4xResyec+n8fPWATEKi+Bhz
eU9coIhJKtK7ejy+93BUMjCyEYe7tN0BK0FyErZR/FOeYhojdqdiJ5PiYcQB+ZmeA5b/r0wwzKRf
AtYPWq34LuDmWXP0oIzbzeSu1ADg3SRuQu+KEfOFTEDC/J+nZOd5jtpEvvJ/7m+mvHtczU412/Ut
o3gw7YvP6YxCr2w8hDTz59+69vmx9c24A/NbneWvZtBgk7cLuVgakvCoWyAlX+vn/7RB/9PJwCSa
4JuoFZXMX92QyOeVerHzo5+l7h1hbRQY/XwK4my+iGNspv56RPGAAYrfsA+jvTgaMThsaO1qABOt
hN6bSVAlCwmQMMQJ6lmbIbbl29Y3fqhsQmTiDHvfellLDAmJM8a6qLWh19eYuLDVT/h89EO9TMVG
1vi17AxWb7nO9MsQYXrZJLePKiT9HCHtxTW6dIJCiG7c5aZq8yP9694m4ZVuTlaYzRUTzzt/Q2uS
ArYR2FKcLmC/8SzdR5IzDZQjslLTVVKooPr3iqgQrncSK3AirVH9nWVOrGXgLS/0nLAjtGG3yDcQ
j70Exirg0OpOv8Sdnya+WMSfjUyaR58RKIw6zRs0D8Osnjl+PuT5LhDD4knAS5xWiIzFgIRbyDPS
rlv0KJ5LJ4/H2Ho+Ltc4aFPlGRqPdBETPRudV0uJsWpXldbIvkINRcJpaAOaljbYKekU1mUO7co0
ONxfB4Y1b2x0ahozJBzx6mOmRNvQVJW3t56tLiPYZF9uygJ5X9GMzU1mNzMzupj4oeyQtsxFY+dL
SSBSJ9ZInsD4lZx8B+l8v7W3S0bN4p3r3+4obXnPWzAkQB7sFkZyF6sUzRQvrXanJ1aX+OmUgX8s
IK1mWfQDh4NohS9y1GWj6ipJDIAN5TluMDWlDp8F7nfSRilyMzkxsIiwx/BULKhG5iyo023KrArr
1DoT2NUG2CdmBpdL/HdW9zkYAFftxBbtxW9Or1bnSAJHscIqO34K8LULXLItiHAC5J47DMpIbKh/
OSVM3TnC1WthsOAlm74NkS+yPF6uc2SqwOXzCyfdp6NTsckIMerLICnZxWqRtHVwYuy+bPzMV5rq
nOZeJKjFkbwHvlSX/8nR8TFobBxW2OFuDtplYZS+ZheNUnwOcj146woV/eQck54+P0P5SSPMz19X
KUxommA179lUy4giy15X4IGyi2raLdHpn+12je/0cgvLBNBJqqLIvCcGR8Zwa/IzOhOT7B6X0SU8
Qd7vDINTvFFE4d+dca8LHGPPrkqOjc+c0oXfChYCPaWe2B/MGRiaNNTw4egDH7r8OJHR0d5weCMu
k3A4uPkFA5cYihm/2YbT5DG4gFzemUYLV87CEDxZvw5QLqRpzRmazkevCktFtK23dbNSpMtX79it
3wc59WeGZIns6pFI/GhhEYS9IwBcrZZ0j/JZhjavmZNXrfYH+/a3RoGFuzzpZIlXEsYwmb2C9Ejh
oGxyHMGIbFnZkNhAbdqrYDGecg0TYq048TGcvhqWVuNfD05bqyHU95hQ1ZkyAn6y3WmJiPgkA6Ut
fJhbbuK74vQxhYyUbcvodord/wIHGLFmstTNISMAd9l5YEJTUhw4SHgtShNA4qk8FjwSc9YaD7oJ
TbsgUcHHmFto5/ioqRwnPmmXXbVNxK5+BQovY6LlWAg03l0d/fhXjsyBsgwl7jzmqrnz826RSbLY
I5YATtQAVQ190LUFPBv5uElc7ukm1yNW7tIFC3jBfM2vlSKZh0EpIzWiKJaCh6m3HkqrB9ZRryOz
4uUPifcPekoL7jEWRG0Oap1/A5f8Izui02GrTT4WChsWVtT+dgswwJeoHNJmDJOWV2VJFyTd/q7w
Uj7dhm2IfIR7aRLlb4ZS0OLPXxP0pff5SEkBx7rqCMqM9PYrve0/cxUM8xwfRRRvvVa3mY1L6Yx8
OyDqQtgLK5XFhaDKBgBXz9u49rD95BqO6ST24eHptEc2Sv/lOxvlvn30GbFKUVTmzo5jHxjkH59Q
7UBVwOATgweltPSrQTjFQCyRrnYwIJwYoFcY2MieijImtLVqEg2rTWmzxPVFJ+86OtPDYAHBpNOp
xYqsLa7NHTVVoXTWBi3+2BG9SDt7xsKabSSlJ8tcfsHvKjHOf/VYQLCevQ2xm8gd8xZdUx4Xi4pj
wRDqu0mUF1zj3wZx+uFhQPrQSXihfWWZivQCWyJqRPfE39m0fkwvYQnK8EE+nux3DePMKhgsCsSO
70mGL8PhK/xPPmPIgAxc9ea82V+ECGbaz+uKvo8nBIBNrl6nzR1uTUOSuG8HRLvwfGZmmyIRRlRl
kFZVe9X9xjPCs6fgRTq+hLqqXmuB5BrG5KH+86a5rhkuxGGo3p5/fJxCLJFbfUwTJnlmwx0ibTzv
SFkFL7qNydq6JrHEybgYxwQF3k54sXrutwuMsn4QQqZmZaMjHM1jInF90r6t+8zm5dd40ywWYAF4
y9RCoXKDDxPGQm2i4e0Os6xvhsFB8QR/DYfjA/c5nMfnr4KHQEONKgQ+SB1z23ik10atElUOe0Rx
4VBseQPA4vFI4Ur4FksV3n5v96LE1Htrdflq6APuOXLjnh8atrRivV3mqlFK5fqf0BOYRDHGfTqI
BK8gH36M5XnA2g72iPQvgVi5GrnTanNLgjF2CUOZ6z4mAf9ag2nbAjoluucqjLft3P0bD8YuzKeu
gmLo8bbsyZ8tulvgQL8fq/O8v8N0JpMRQ14YNaxJLs5eno6ZqtD+uQOHaWcAdqQw4mq8fmy2tZxJ
Dr4C9kg3O4ts7esLotFGveC5/KZgJ1rEKqEn1j14YfbMTVbBkdZR5/SpwE74PpwlydjKwln9qNHS
jmcdO7/xrEz9KLAen1y3dCEU3fW3l6NULwHu8h+bthFTMY9Yph/duHigTJVl552Es6QvdyvxDxNp
tqvgsHdbkYaDFkoM8kUkMdu/ZscYmqHVkzswwqrP5tkGGMwuM+JgdGkOZgR0CFjpAwk7hwNTRkW6
ikg0a50lDpaesiT7/Y8k6512KPGdaVI4SpfaJMF2Nwk4wlx/IyjIrBv5ItGIL0gz7Q3VXAP4tsie
UNEJAz6CEUDNyWzMd5nKYaJznzuiVxGk1TYCgI2ayuIccw12g4HchNH8j0OrJenW5VAvj0vBULJA
gr2bxbnZ7apM2oHK++bKlColwPGVlSNAT2KdRkoGQrQnU9CgxwFK64F7DFkkjY3RqaLZz3hl3ZqU
8HMztd0ajUwwe0ciK07QSh3VumNK1Boan7D9yfurBxUmU3BUVBdPZ9i0OVSAbCdzFO20jkGWekwv
nIDKGd5EgpcyWopsxt5LIJWbUezAKA57du0eOwpeQplESHBymD5kxhfwk881d1Haw3ZutZH44Aci
CLqr5LHmtid4OOy/u+4Ti6OreKaOdJ4uzjNyBOknKWEgElS/hYTkS/B2GFnBiZYhKA9M3SmfADYt
1+WNpqXX/o1MDG3HdWaOwAOLjv4L+EwsNOt/d66ZZZLqIb1iwQ4C5nhie9p1DPfWihBA3fHvYfGe
sFHi1Juh9IbwdlZTEzOtPcc2dDbFkeT2ltCsXCRJKlLzRqsjWMayVmZfRWyT/R14p7Gxv6ZKzX5p
yW19nz8NO+EOqZkUrNywNkxBGNnT6+OB0AKUpSpG8ArYKJgpXiZipQeMZqEXSu9iqBW4yLFqe+/B
gWCGaQw2fVdjq5JwK3++3UtPkZrEjzcmC92SWdgvEOA9BR1hJakMAr7xEcRHATWhvi57oF2TJrls
BP2YFoPXTZiFBArn2BwwHJMQ4phdUlZjphLGMU4D3eLOag5wo7pTE53g3KLBmkAqFIokQvByD+Bm
yOS2adGHWSFN/FdprsmftjqbLhqXrkPToZpLShi4hGesocGxBKMKGE9t3UhsOM1bdKqmrTE1r7z8
MFU7kvD3r4b57EjBK3swUZfBJzjQHg33K1WRlF31LMwQZiw6T8dTqF9EKCr0RYM+1PEvEDQRj8Mt
ZsILrCj+PNTpT8pv3TFeHqYnSHCfGli9Zz4pDD9Xx5eUSMts4BXLL2WzEU1Xuhid6YA3jVz/aHsB
6/Jo0cKzLZRen6Dk0pdWV5BucE1QfnX7LJ8x4FYqMRJ63wdLnysx7DK56YZVdwOQzJ/8+7BWlVEr
KLiEkm6K7IRm4PsIQjaXhrzVgaIDgsI91Ym7BvphPusvcq+6AXuEqDADuVnNdcig/gVd1+lNfK3e
pVQEynG70HqgSsStXO611G8eyjdH7RPL4tXYUwbr7qHvDlnfOJZV3psm9s0Bp7w/mcKAxDwzg1lA
Iebdc4NIrBYlHlw2owU94hyk2hvbXKqm/okZJBU1FaPOCj+AAGxz5ie1VJbGKegEPyTPRNjNfGu+
y3YOUTyTi/A+7CW8U5OLHB+7FRT8pSj3Afb3CzaKB6IgGVMvlle9VzN97YGdckAyxtXQftoEORb8
XZXbWTZZjKIWvslRCR5Wfr0otNLTMkqDj9gsCuw0d3yfOjVq0qenNdDMfCEFQqMJArMBW+B5oor/
vIoTK6hXZGbdly6BaM55bNHDve/feT8KZhyxQXBilaDV3G5phPmW8Ck7J5Q0K6TndHBRNuTMNIvk
juQxM/4Dc7phNh2Nf1m4W10tJr11aM867t/J1ulbx+E4BgBdO0/ld50kKUrKwbINl9vVV+GjBQ73
qXV++3mxeLEbGtEGRmEKFT21QU37NXBeOHUFlKulJygwtKWhInMx2hwY/yR4gCzsMM5vEgXFt8oR
7hxjnCFX8wfHEnjNHaeTTI0g3+ecEcJGHEma2x4WRbMcJ3Q5+/S8EkBPiRXUxT1I8kpkVR4/iQo5
egehSvEPXu+ol3z1WR2qp+lXXdWLO2+v3LZkGMUy6eObR55WyCT2hrUmyoV6lNdLYMDw8oxEbuL6
pYGFMp6hVEE8zpma5YemelUmxbfoCUe0XqK4Bif15eT4iKyOZLvbXOxFuVwaEcnSTO+G9zCY9j0R
ZIDkenCDPGxPIZJZrOlzx5uQUs6EzvRSysH5Z80vBCc9UkhauDH9ZWyq5HpWEm3EZFTqPx6q0Qkk
BKzIU38x/NRIpzZTB3wW7g7oJH7QkTQhNJ7ZSo0MRshJfMqQttsU2xaVTsAgb9geWvjP56eq3+j3
l7nFJrdQG2qNdd6O1vcdDWIeiH5B74ECQF/8ERzts+6ELebKx3ezSiP7Xti+B36iwkoSVrc1M9EX
klA7Dxy0XjnYXcxFM5cLm8NrHLkzbrvJ7bMR3MsrabhBoM2T2yw29OxxTmPHPt12vCILebuNZcf4
pUAHMgykeaHYmf/m74yk6u1F/CPJEN3dnKJ+8wxwLPtwMbdUsrSqJvMAZAnfaq5mnPhnR4tZfoXJ
DrDYcaOTzSv7jp/NW2NarnRvqCbKNEyMTOfu9iwBcVT3wKds5IsQ/M1BNXqYpp4qKau3LXUWlCLO
Cb1Cc1NwknNO0zfdK3D2P9R8NIu3Cmo9bwN2QgPulmeqDXfsjbmJSAdxjzx1qDYZy8L1061GaR76
dxK5RbvfsYspObHIZYBooIlq74t0UK5/4GxkuF5MgbQBeyp1pVXLwaenZabIfGNQnjPQ7WagWkx3
hvZ+WLPcfIXrMdVcwJ5vAskP/iUdazKPTh0pjelUBh9tva+s8uU3GkzTdLBdXOGZyD1Xfar5msJG
UkzEZlauB412SfDqyw6Np4tLXqtPHfzg4w22m/GZLAJ1vtlY/9RnjrqfCx7LC9lYvDUZTv3BpdGa
I7b9vlePiCpxA/0CyZHJeVs8e/hGE4wgDUtOam6Bv/BZGpj4Y/qdEKBMhWRMEg5iQBUp+Dpn8XKf
vMZo5LKq3ozSqYCbZnZdx29g6vNCE8hHkz4f3/mH013BpaLWqaeWsGUTuKVrsYSMhb94aiC/g/l9
J56x5mHtIIl1l6jZBA1Sj4WUNTUpqkBlKuhuld+GJLLX6+ltSn2bdCRp6NeOxVbAzQ5JwWeUGEDT
FHSAnrR3J2K1YAk5+bYhvoYNMAjlIYLQ3NVLxZuoZgfAo1AjK4Oz4170LE+iYlfFiW1LC6rn/Bgh
hiUTP0QwZds44UsX0Hr+tA5kRlfQU+Zxug7VGe4C/Q0ZVw/ENgyESHgN1glLwwJZ4nWhhcMmb8rf
i8aulC3B1yYrtMR+uEk1CdmMTf73pUhz9ztwxXnFWerC5Gu1MTTw5GQKDmLHBmyWm+RZ+3QYIw7E
NxGbaqljqZ2E0F/Nu6ZuVGmF3zN8N9aeMiy/Ot023KeiF7rHTAx2XdHEuDkqUhEBLVxQkZmMZ2Iz
pRMCFFzveHx557GnkNebemfbpgXqhquUvxT4MGfuOD1h/9rtVsVIeQCAf+xPx3eVhi18MmlMW5Q+
TMRmihD+1cPKk/65FjuWOoZo38TnZEIfCuI5R7OvBvQ0DuTb+6dnpaOg9vmbjujfIOR/cdD7IDw8
QrF35Aaa9BVn4Xhg5AqfUiabsV4gXcYT1FFfJjbFWkqOvXbUAlevyVqHSugEOCkMQtFPW2PVLjK+
YuywuYzxcAuKn8ydLAu+Bg3RI5ttfslSIHVDpVQBMQ9f/Grg7K4LrqaLxliJ2DIJZCcKtqsVDtIy
fbmYhJr2vz/O9xNGR6hZIfFwnzli3aNTnnGpJL+NLTlrUw9uoPDog92chtSl01KoB7tl4e+x69fN
mxRhsgw6krVgKBb/fZ0xboXubyH6fHom94OH8esveaPg2sbdmCVHj64RXHGAVK7+W8qof6miOuqQ
N+78FRo5qMswwpNfD6op2GpImbcDgyOhGIBVU7kjqV4vENekncsj3pShteDRDD/4LCjLXdzLvrAw
yQpCGuNRiPEeeyGeNf0neg4pEdpwXXpSO/dHnEouGvE5KcOf/tqHTY2V5VRMKjGsjkwD/U31tc1r
rSYpZ+nhYOiLMjScE6msKSfiaPQ5TdXMF9M0EL+i1OkWilwDzSd0UZaWBrM+dLguhAhDXtEJxldG
MvOCgPbABg1sffKaDR4fBfEgJJ79pDAiXWLaxP15UVNcHPh3ZOVSGXsaKEqpT3k4Fd+BhNYQneeE
E0FJcX1jTwatn4C296ZgPTK3kJyuBG0F4mlgPj3Qd767xzpVHxruMj+ImBZPXpEDv2aZn4M3ptGi
Pv6BRDbNCfZGpieJGjc8GyZ1Z9nAuy1isa9Qpiyw0l8QjUG1po2RdvlJp5f1Qd+o8sRDUdWJ/T9V
CBZykDgdrcxt6TKKo2x7EHVEV3hXBhzmOlZXe1mUUYf9lmzAS6zIXb2AsnqASMHVCCPYMFFHWGRw
VbzP9E1LwxRP9795NhQSuT3PP1wba6Tqs75P+d2sWQdLRCH2l/w8yqkZpy1rm7W5J/ySW/4eWssz
2pmqT64ViRNkT5qB7r0j34YZcK7BY0HF3XQHUESABkb94DCtAJUhf/iWKABduE22kIiKpiUOwjIR
ZE/1Km/2pDEdgCLd9xAl2BfEYq3iotQeuZU/sBFHTfwo2yNVJ+m+iruvDe3cmTsqlbnfp3h0FOIr
kj5Ng0naXP6ZtlQ7s5gcQU4BTOFs5fWfsuOxwneZDnLXuL02+J6I+ZnPmxee/YelaXA5rpdeE4Qf
5SySD2XHTaoEmgEvD9ZjL5ddP1L2PGoPLzIsw59HXclHhztz+BXwu6Yp6I/kcMqR1XVQjNfJKRNV
71kqpitcTzZop9N7jT2bWut0zaQw85gxqmPRIHHEXyFU+kQmIZjSDZn+v2BKyM2WH/rl8y4bZLtI
gW/7vSQgy6hA37pt5QZRuasuOVnBV39GbjwcQxHCwxIqQgYn2MS9I85/gexicvOoW6slVqc5mWsq
8dAZ32Zl0CVFEEk/7or7A+MeGIBtfscKqko+DN3nkmJbLkKBozFCOaHqoEQvLeWSRWx/eoq1PGQ9
ZXC0Df+qj/IaePL7LJF7s5CEe/xqdXkpdaVY9w8RzH8pyOKbmweZvGwrgsNabLY+0zZ0xO6RB9Sb
viD5RfTJ4C3kpUOSpA+s12fDN6/9olx7tlCjZTY+utDCFvfv0+2FFZNE3qcCIgVCSp7grPwCUsXZ
4Mg8n5574kZmvBGNAO3w0wDEL6Vn3OUWDF1UKeANnYerBjJuss1yNxbQZ1MUCZ3hD2hF9pzGpWll
gSL1YE4eaKk4U3aUdNdKnCt2F6EZw3sAWm2uFsRfbArZnU6etG2PQP29iL/Sn2CH8jiSUEB5lT/Q
oI1Dn27rg1dObPHvufw68IY8EoXoQDPxCv5FYtYBqpxwqx7eucHuBBeCeYzkfDSYa6vwgUpeWX8L
lA/TdBaXSx7dW6T/G+eS+nqA5nb00hPLmSs9eWhdweHQ7PLsO9ctXUrXM+Odd8bYQ5nrrYKxYfOj
i2GPmXaDYH2juHSM8UaZJ6H1guZWEJwck9s0mSTHQxXMrHtEeKQgxX9AmeBUgORNQKt7WO1/tBiz
9cT286PCGVZwRF6qYvYybodzCL2n79ebGvZ1dpXWDXrJofcuACxaRAybM611wzYsH3wR0QMXaM2l
c6jepCd3LKl9+f7BxbNlXEvm81RiiKIeKhDu07rOqCahnpJ+trbID04bIkEVU9YIxHMIZd2dNyiy
BLUJitxIE5a+6jis6z75eJ3IeV4Vq5+X7Co3lr4UUkDT8EAEl9vBoDBUuHCCY5wfZDvz6Q4Mc91t
wBUD9knKDpYHO1Psvp/ZXpzFn6FalUJhBen2YyKsHR/0+v8Eh6eAacxixQouvD7OtPKt4yu4QxO0
9yWY76XQNFaUOVG3IqMS+PdwzmlgZp6nZSILLShWVgyjM4CcXSas41ZV5hWtv2gL6vVYLaFDZFdv
qRQ3IrKyeNGvPDCNQl5iTL3cvPAepqo3WHHpP0HPpJEbzynJPwtfpbrpexSkmKvwOTMUkbe6i1RV
qudfOKnNkmvQ61p0zRUv/aBQzEWNdpQpGZIymPJi3mJTeh0Bnvj1GSSVPkJmk57ZKp7M4yAuMphH
ZHrbjtPx6IJC0s/MHAKoDA8Yf9WZ5Nvn9vVU3+jrs10Kr/rSGNBCYFbWQN6ebpLJI/TTQWOcO1aB
MiHU332jP5R6XnosSAUVEeKCrzTTQjxf19pCnLz2KXpu3mYrSpY90nrIswMgTpo/q9vgVhmjMctG
szvoLtRYennNWMGKFJz/tKtLwW6d7ZOvA7R1I+uNYZb5teEV8Z1MlvkSVa/yEOuGQkZeqldO9tYf
9azsVmOZEnTXl1WY4BOAnVzstOU+OmHI5A99+G/Uu8AA00TWr5xFOHivdVYVBAlYhNOGxaEa9Yy1
bi6tWZc/HnGISZdsufw4l0j6QUlaVIEnhQPyVn2WF3MP6tX5UaElt12InaD1cp15pEk3eu/cehmn
jKqY0TncgI7UUT2L2cVeNZbtFRBl9dGEV+Brs1F+VhmBE3z5a6ui9iBmKgq7qHcF4NLsrQADi935
T0dHQ1P17idBJAbMc7xA446dj1H4VpOVggO9eE1bEU80ksWgUVREN/jGPzXZ42mHfvSw8kMrIPB4
oAFD4Fs4j+c9kO0JFPg4u88iLJ1YkCy3IsVPBdQl71bfClHjQN1fc3RlaKb+/4pxHYxNA+NtngST
e3+gvf0YhwrPH1XoLOgTW02fIopxOmdzNBI3Z0xq/GMEZcrr2xQMy3bPVCLdWOZsaxFXrfNvvV4i
2ovqqHyD0H6BBzgr94yf85mmCkMGANVUeBtBjsRyh290vxGvBkYe/0z7N7KVPiLidDlyFw5T/4sQ
+BSDRj00PTljgLOkwRTv8N9HLRSspOHF7CVjRew/lE+OYsBKD6lCAWds3RmlJqeUe5PCPGtqDv0B
yq4IBmJmR2S6Fhfmrsyvp2BR7OPhyhZ6Q7eMM+unn+A77kIoOtDTDs14rlBy+mFd32bUH90MNl0D
6cAHO9wwfFmY3Nlbn+m5doxu17RXcGEHntZ7gVQpFc8FhjvXZOm/SnnaKIoN+jf6/J+75YwvpXlW
0xcEMbkjXZlQZpiGNrHnXocrjir+px7bbAYcRY22C1nPXv10Ae089DJcNFJVkC2S2RcVo12CsCA2
RICwyaLD7PDwX2Svqde/HoCPvRAmM19S4JD63TYiD2Oj4Mrr8eWylbiF4QgPA1in8d556sGP1Hr8
YRT9zzyEBiVlfqyjKmU6n0L4vP8+hZ/wO57x5EA/eWvNe4HiLunoTHgqqG5hSPHSVjQF0xXg77r/
z/ZDYjgZzdDvEK1IgHHkouCh+qAtU7fhCK+nGr/BR41x45hoDyCFV2QFfzyiAHLxv1mW8c3YDMxM
eSlLhO5DfgCJymMmbTw1KtDKF+rE0vBrMukDw/UvnGsTps5MTNqBYNl4/luK5ic0rqRYw/c9xgHY
u8StBqhlDFnLa//pDO7lsswmqQSm10X+/ydykS4In7nJcLqXBU1fqwtYzN+Ocf6eJqfSITfeWQok
vEYxerBhy1GD3R7x6taoCvHja3pKe/PYvIckPUL23BktkIeRHxrQHMotN2U4J1stYBAAosRjxBTz
jOUASELm4MIG78okKwoUcNP4s5Cxl1isk2NgmovaiJnHE1pKYngxogF20E3yBWmE5ok353X0mMaq
DkLaqRVWRT338HmWeWGFdEdKQySeJJvcJGlH20ZibI43ZzfzabuckwDCFKcr0tGsyHorN69fZDuf
RU1Saiod4eDKAjSfHq04gTwQozK/dvJzs/hZTP3NXlFlzt08P7vcY4I1tH9UA2uiCVjdR8WLcBEo
ROb/KqWn7pZt6raRZaRPRGYr8EH/36vfioYHHaUGBSh/AvNCZvHwBuoWekD8P+yhXPp5ujGA71/z
m/kMTLBBrIeGz7JdJzXsmLEAwIvlptIL7DN7WWBfkuBT4TCPamPSCEsrQ82i2WFle367l1IvjFjz
UvYRaxAcC7c4sZbOOSHe8sroTKTRsIUmNl7qQYgLXe+W4G7F+MpC6/h0cT9+Xy8MTSycblqrKlbz
jwMwFSyr94wjhLmhoTLcNjh20erwUa0F7b73+9nAg1klT8SIwjyRjmeJ+Z7sDfacjfhOCoaixUQj
FXP+HXYM1HhxSvqo+Dng7OzcC2tHAML07ztBXeddeOmSPFrvyUlGFPsD/ALWTuqEBnY28MKOQJQT
zV2JLZpsecOSf+isRj8kuKXZI4jRZUaAyFippcl3MhnNFgtum2L/NQA1MxkzLfB9iQZseneyWSP6
/FzjBbYQoRb23YNQPkbhDBgjNpuYnaBMPYnOB7/XidnSz0LFqoXSOKpJIto/9xxgyNmqVrccPee/
S5gWwwCN2+MEL9w2yzHYTPjg6f2jZowJDUf6nfe2zUajsIJTGEYLOVq/hwoXiv3GQupMC6a6rkeD
/XBAgLJtFHSVMG6DUfcoZOPW9QW379xOmLTl+wxW0wfGmyU78mdydSi/Y8DnlWzgoLzJvyt0Ma9h
U1QtDUqd3tihtjgucoeXqqEi4vXFqEhYdbgIQSxDe8Hvqp8G2CsEUkS0U2TfCsO+ggxVBh+Mkmwc
zio3/6C2zW54gD+eI4IcrJdtsFXKot4YAsWVYnkxrobZyeQY36kWwb0qmgXv5FWoyIPYX5rXTQA0
qBKzuHUKzijwOCrt/qLNy1dpBno564D42OoUXp7rJgGJIX/FeUrYuqIyF2x41N/pw9TpTke9crFN
aCC29mh5BpmNGx9F7uutctBoed364yW2Rn2UlwvuS8pVeQ/qTSeY1mhaLJAg0oJfrdC5DgCpK55Y
zQY7+B96GvMUzKQFId6LpyJyns7H1WoausXu7CSk1F/95bWJIP1k15v8vK8XSGy0403RXTsDg4IU
YTEsvPGuhAxCnX35u+OmLHE2ylWFqJcsDbjqYn+H0M0sQSl1ixmOy3LEZiimspGozCXUqtJt5znF
lrPN4xBtqYHi35UML2t21HE4EGwuHUBMZbnbGeAzW3xokVhVuuWiGm1HJjzyDg8t3OjUd1xk0h6K
HYo9rvgRw3BfPaxNMZ1eV841NDWxJPrTxijDLrnoQX3B62ulpbQ7i0p7FYj0bRPrkJS4/K+u/pxY
usHEAzm0Oa2oiAcce2PKDSdDmA+fImcF3S4OgCwKt1MXIjN2C1jmml/7HwNQUoSXmWS8BWgyfA9K
9XzLRlxemX6B9QutZyknJomsDaWa3bi1dkBMfWTYv6gJT/pBLJajvYzQFsWFDlPaRCKh6kcxXp0p
wWy/SD99zc/ztNQiu2RJjCAFEq00ktuXghKUbka3FRYT2q0VcYzr0glGfgIdibtIQk3POb9evjrG
xprlp2tYoh0mG2eS6rksKlO07tEkN6AqbgLuyhMssET8EMNV+Lk+pUDFW+Tw2GmzwTHhVNDUY6l+
Or8CTAAemk3FXFrnzO9FUD+vtfqR+Tvi4gZUEEyqSzwD2Xb6w671+9eEx7RDPiVvxxm+ODAvD1z4
1FpNlX9y6sRM4xbD2JJFEdZhI+hFEy2xA8ayBy1+RESkHHIsE12LZnoCca0QreDcgZxNcAmcRYpI
lbvVRjaSGGdCpeSxj7trGIaJIKb2By7jOauoc5uh6wO/fD2/XQY01ExoEhg5kXagKvabXX0MvjGm
NEcW5CULP8HTNfg4V7mCVL+5O6dDALamBeoo0jNmjIBmer1rMV5JPvyS1U9LAaeZQbF6BpCkPfv4
eLpezN68zWgLkXepWIhjyNASKG5zNlUrrD4Cg/dXsv6lcv9QYzU6nl7yHPHonk3rJLU5NifGOPHU
l/fqRamg/MyTVE57bSXoGI/WGjz37gEmVH3Oe4c5ymYY6re91DG+Ihsq7/gJqyVyDYff9luXhxQp
arNGURP7wXn0UxtODNLxQW0+NsDuEnL+cwaaXGBdH5B3NWog6sE6/aC5lP+HJ1j+qmlDDETpHEXZ
qhXl1hfrdALpSEsrextNtZ0TemfQN6MvwP5NXxCBSiRMqVN+T4kB2u3OyZK1YmhJxVhvPxYqmoGu
KwH1zHXHqItrCn+ycOs2hsMAQ6VNc2s4Y5rBJIzGkWemPucNYCrKqs+wrUd4HCnRt9YK5XKzUJd+
6nAlN8CHLXruqh88wWB0qNNq5jXL7t4Lf5lA3Abxe+aRVReN8LBWQ5YrrCUgFNQz6DDEHWpnkUNI
K19Qu1QCh3LcaES6MdDSUp9NIolS1JkPdDvZ6cJvDiI0rCoATLxRuLYvTS+NLLAcvmcI6JKSKfWO
jZa+zE5Vs/0eeNIpYYi0ASWbW7RMcu/so4BZBKS25PWgwbG/1jGZEWk4oblgnCVuOc17O20PYACn
4Ch9+awyHNy11m1SY+Jto++ue9dgkB8zn5c7vc95F2Ea/zK0mVh302VDNml/TH43YGXWWT4uont0
obTKd29MNMQ7hDF7AmSyvuN0fnreZiuoGqm0FNWWqcorAlWVby067X0q+v57JRTcjaTiWIuYXGJs
8C0o86m4mMvW8Qr9vdsJk+iPZpJufY7opSCcA20YY7Ooou5bTjteHPEXW37uzQgXhukVzgqa3SKw
PrtCdP77tgA6P7rPe5hyVrUZ27FV7N1HLjWvecMDAPRev7Ubhk/pi2HySyxBWgJ/8v19bzAKGd8X
7i/gyyF4KdoTjjZyLOX+xBlp1eJV9xFBuo6qi7qTbccRBYFRUeP4t0WLs2+aUvEcDeYhTFO83enJ
ZacGy9hPQhw3RfvA/Czzlm1pp1svr6E4uW1UVDYEbvyq74VeUKErcjFVWEqCY04PjOLT1iHf1T/K
PzqxDt19QLVEhdFBThWnFc9WoNs/KoO2dZ2zCxjT7q/BRW59gqxXpixJ6O0deIhlTMe5ecq0EC79
6CpxcHd0jETSonwL9M0736DABX8pq/q/amlQ3Oouhq/W4FVTrTZuAjrPRpnsoJttqb0ee7VLDg3A
d5jQ5d511MLzMS7F/XXqBLwKXjmdizNj7S5AjSqj1PVz9WXo9vRxzVS+moXZMSAZ03c2CON/aBXe
NGaXbj7+TpMa8fLVZKFhiG9vbWZyXzKFyW24xeV0k1EuZSkmVsSSW+7GjxsIV+nhk+OxVgJ6CRHH
rNxRNuvWy3HHZIYCokehIVAvgPTr/QwSIYF3Y78Nn+IhOQrz0r0rputm4pRD27uwEhHIirAudjvO
/UJHXjey7I8eMcclMPu7qWU3+m9WR/OyQ0cdCjMsfKtWGyCMkvVt0jHGaQGF2rMsKnyLX+6LwFID
hx93azky7C4N1ueeqg4rWKsZDMllJZJO/Vl54KLFaSsjR3r7FyIGs0CY8cRcV0SpWK8Ni8Jx7fL4
Msf1Ds7an67fRDSAEXbapi+4n21zeFD1NfHvawVR4ZLZAbk8amlO2bSSE3lZSZWX7/vYWhRSN/LY
tQ66J+W6VfwXRztmTMupqevS6k1BlpAp604v0sbSpF5D51zTBFsxP3Z8RauP7MpFzvc30Ot/hWe1
xdT0opB8n9lG+rqHGg35qz0EWyHdTMCGp5fpz1egbkaYNdekx1y1wmqzv2qVRCi9eyVU31CnDTvr
gndLlVhFbJqw9B1z0MVZMs7rxhtMTLtDDMvQeat5sI0N16OysWyak7sFbJarP+K/St2kLl1efzbo
FYKko2kgEYDb3PyIGN2A3QVfObHN+qz4DZHdsYSEMa2VjGO1jWJ93zLuPsb2bXdN418nllyvR5sR
3fLPvo0ZY5tINR9zJnYhp5PGwLaV5HhtAzmQ0BhgIFoDGyNdoi8ihsMlPBG/0uvC68sNCe8gsa1P
4P8+1/oUWjQkuEhh87xO9ekjSEIDpj/30i0i6alePb7yD2tdNlnF3MG9QU0bUVNUmDAgg1QFLq7d
rgEIW+ftZ1DgpMlT0QP47/CMOP/YAmNRdrOEWQzf94CfwL73Vx/umaonyoA+7io5Rur+42qa8j3q
o33QUUB7E6VKXpdVoi2FKKtfUQIVi441NXsR8A8X/ZTyLIVVt4UVRq51iDkWSI//lv0eS3EL9RG+
oMc7KBQAuhdBa8Q0FAq2uDDmrhmm6bF5JEmDGbwduVIzEpXtd4PJ8FeeRxnFeJ2Zqt7DsOoOi+FK
iit+c+dDo50eQexU6gZTSW4lu395nzmHDoh88l9skX1LIBqEk06IJ2oLSOU+GSj0IWXwSn32clkY
Cm85nlD7+qN+MO1svMNZWbrzQbu4FsreEY0alzX7Nn8EGwr26NvEMyjmrGSKyUPX6B3NhQB8fj7q
jDirfEnswILFNchQMbdqPPYlsnQ1F60sR4S0cqX+enrk2oE2bk5fpTChN6n4MKYLlPJAKY36SfM8
LZoFkcZfzFkanRG/vhpsqKtIcWeMP7jz4BN4kb5ZTJ9zBstufB3XlijOq0GMSvMcZdq7hMK6MKPw
2JToS6FIygu8AaKr7/SSvdBe2vsVqOw8N407FvdBWVAXlK1PdqtlNgZb1DrrSqhPtWgzWOFImK+r
d3ic5N2e+MUZjeoxVvgD9+QjQkxFQNIH9RVITWk84xP3TtS2Q+gWEg8FPnrzI/F+NoQkTbh7Q1YH
ggrrvUPWG2oDkOFT9zYThq+wGwoVh5z40TCOA7tNTb5EJJXF6ERTQN0wsrnq2AirIqz9NEj0Ncnc
bM8frCGPn8AE+Rb9GHKgiiPKkmTh3zOswpKSXDemRLSsowHHDTzmvaPREIg7lj5YPKbV33NnKK/K
1PusTRntIFZkIe+JbmWtFk6aHczmWJzwezGr48w7hgMJQbz7nIpyDoVAgNfZSqT2TyBK6gISOgzI
GNffg7ab+egUxhwaU4dDBa+LxxFR13MpZ99v9F8GwM0QAhOoBR4+LIoLL5DW8NR8rSfJwlGdFiUj
5Cfnpfjvv4GI9pkcpsqpY7vCzulKnbZgmoypsiJpRO/iWBfi7mSZ3xFR06cfU/CihSiYdD6aPfn1
zO+1ZGT34OjReU/8T4i7+iQ1fF3amXbwwLDvTvwrTFCRuPmH0QwUC9NYNiJfbs82skh7YN6CiWUa
kR8iaw/WSwsR0fQSY0sH1CIGXpcuBKD1Ry2C5sgHSlFnt0ivrTdjZA362V0LhgKGiCLlh7tONxen
EvVQuj0JqcSTy9S4hTHuIgFe7JHdbpsEzHhLPVxIQvmDZ9sB4aqjuPBQ6F76ZFEWrDzRkbmf9Cj4
C2Gi4bn0KWiKa/DXi9lJd4rn9SsINNLfnCct/frWbmAU/Ivu6A58jmFZlI1Zh2LMx39v5O2aNmA7
okzRFgq2mB96V1bprZWDxEjQk1g4szO0UmF4h3wlh7voNFgIupKvnEZs3xGp17GsYoJC6iPoD7aj
V66ujmrfBvBpMg4OMX/r3SivVRkpKzp3X91uAIzXhXWTc29aM9a/ZwJYfow2kg5N9DyoJ4nhuPSG
BcHlxHKPvjafx/VAsSPxAmyirea69p/J0TWIgl7hr/6rofA8uVqcCNDlX/vUME9jWLNPASWETNhe
K5UrjGqvmbaIFpIyEa+M6Iv+4pzh/aLzssDBt4yNekwJJTFHqOeYm2G4jYS8dWkZ4ZO7rMEhBHIg
ADKYHhAVM+LKmAzrdhdOJD5WyAVCnVz8jgDl3ZrwHwMGWUEB6b7b2auC/46Pqfwaz7hGdPtxsU5F
1UFfMqInGEBw2eR9pj7t3p2c2yBGKQlEDEYotvLGEMrwDOV0ou8JEzsFG2RB2RvnqzvH+6XwOXhd
Pc9emOjbileSqXbL1riUbpT97GBstjRgfvEBEJJD8eFlcj2ssh6lpo3oHnhjztkMGzOrCMt6dTkq
/+nh9+1JOkBzku2pi5SfWFRrMg8v7G6CA4onQacBx2A1OXypgcZWuGOuyK+yBdxK4tQl4rHHDgDg
cvsIzyddYNRcIgJq6SJowu519iiTid6legvcchDlmIF4MDdkOLuqIXPJ4LtaD60ipEJiNDGXQhLb
bS4pYzQFu7pN9zO+/MeXSi6SdefeNPL9vTN5V8J5il9KaAMGMMuKTO0/S9mPU1t7b1UNKTdIjHVT
5vVj01PkEwXXRFTffghw1Y1ZW4aXU2CVfIm0mzRk9pB+Jt0NmTdFKk8nqE4WfIDDy3PCGWKBK53G
GZAxSziVTXAjDZByR/JGInvXxKiXuqZZy+CYOfXh0wpeSjxgQDnXM6VIYTJlejDFum6fhA5IfaHr
NoqbmYZgZDuUtzqF7g+R4noOwhXH2W0Gyg+Cahk7l3wnkZTPa4Sh+UedgSBH8P3Y+AuqMpefvO4c
XhUcq9kuffGeonARIRWgiPmOCJDp/mYb3BpOGzIlTSsGaUoOwSFYKSd8CTPMQ7DVt0N8o2+6uSbM
9e0sfAZnIQO7z3dy1mjSxVyj31hT8MSlM7y6/qqtaMYds7zFst5KTVnoSW/GiLmEWVFyvTairvQX
zI0cUFTjhZ/ArRcYJIXRaaHKGaVe7gjuxURQUrZcRkfl2FUKHFFzf0pUU2qjjSwVMgs6GmdYCjKF
Qe7Pkbx7QMqn+Yq6ZtdTzJ0Pz03XNwwei7RWu3XgqtfaXigFhptztqvaAa3YFN4a5Si7wzG9uavM
MKirI9DnsizI7uTaloEq1Ja3bdq4JSeM3Y0HDOHdsVhMmfm1uxw645NKE8BtqCXpZ1OWpdPchyOb
AT4438OIkSbdS57jUQ7+99dcjablyUpaPp8sFiHdj8ZOBG8Jblh7yEYfNDSWaD2Y7EzTnJn836Q7
tN+ShuECnYnV6Qw5LxjNpD19ouA0YPjJdVdN/vFSr+jkvxf+DL0/l2Ms27rdxwkc51YarkH2Wz5w
N6FWkVj8/jhXkviK3Nvrnl0bG/kS405mB5jaqKSIUVhE9x9piWKv12skUhIWXrPOGnOCuWP1M2ng
kICKmj3p4eLrYSr/bvo/6OuolVWjHdfxE6rIf5tNoUdRw8l011SIXEapzlyMaUvFPpj5FsEMZGgG
D//hSzBDuOD9viuKfqqT6nBTSYHqsXpnCao8bv5GL1HvcRy+ZHiZzuNZ+Jl/Hzujn9KRH3b9e7El
kljeCqJGNVhKIXS3+Szn20GTO8rHb8fIHPMmwf/1iTWm2GDfb3KB4ugKd8sfzOi8HvvW8Y6hh33S
ONhcG071Q2rlaLbSggMtGrApRH07ZRuSRdM5SV8bVFHTHs40rGwwXkR2JUswBqTimmW1Syr2vdoj
i8qOHQz0Ja72bmyiwLAdDGA+HreQUnGpn6zKNu7sdX9jrjmnu6Synhab0UCEWXVJTApFBA9Op1eM
mVl2mbEDd7VI6SSG9SKmAXDj3sjsnLSSv+xF/If4SNyAarYnMcq+9MbEOwky+m9YhFxVQDNyWxew
RXm9Mr/WpvhwX0j+f9bjUi/Hp2Tb8mhi/YaGxv2fWl5k8eWLKBGmZ0PcHO1EDComOR47NyLFzB2E
nuMOFBzO7eioTCQuMqY5lL81ypkx2UvaYUQTWI4/rciaZBoJcI+y4+yw0f4SrUCJQHZno0rmzM8Y
POXmZR3WWnhbdBuUnJEpzhKsNEQ86jWC3ODTpFwwnOPp+2B31GSEybWaOeN2b0D3VTf/KdP34SnO
GsZHGZK+IPM4wLONtqo9iovxP+bfMfotmLyvD6x6z5Knuop7mbCg/nckWkt1RVqePgylLUxiio9v
avfcHoHcuzmm/rJlviiupw/POfHf3c5BDxxNziFN1MxXoNIQnD7wb9lkIg6F1L/DsyHBQtioPZ2r
U22zta7KNCY5djG2ALzNaiirJcKmktt7+jGgBeAE8baGg/0IDX47lVzXjA7AwKOkd4TLtfHd8q3i
pg85QU+hAmS2WoKeAQHoOw8s+q0Dq94k+7dMy+mLOEDS6xXBlnRlAE9w2kxhtIJ+VPhhLmJFLDez
oKGnqSOFR2ZzztJH7yRqMvz6ljPrh1NEz8vS4zVfbcF6IXNH6Fv9J6s62yCZc4KUccg1mjD9w1nn
Y2sQUr6X4DtEGmEbYiVhlvuwczHcDVNV0hrziAg+vpF5I2X2PTtBCmK3AeAvUtCDfC5F3Ps2CbSW
vnbaCAlj++3vWp/RTi2ADAYYYhyrNTWkOVf6yjp9G9+q7dhQXXx9pz/0zVLUO5L0HTAE7eeUMdfq
rLVs1JmRUw8l2uY8bBveX7BokXqdKnkB2c6rFHX3bYSa3B5QGsnFqepSyS7tAW5HdqCDMZtoROPR
523nJsnOER0UEu3vq5TLr1P5Ofr0J349tkljJU0KgDIwESHA5Iaqmz9z3OS0n0FfQ1/AtCZt/NNd
unEI/kO5h1/UsLio+HlW0L0Cwygu7F2fs24ok5zFRM6lfgqInupPmK1GwBSNbmsa6xf+w8GVF4sE
iHAB9xdA4FuFCUXXnkqlLlYyursIT6dWchfpySqyCSjpYzHrQaw7p96EvKAX3ZdgwT/Xm6C1DNmW
uHTZzrBb9y+DhRP2to7FZiIO4PYjYlg6TLck+Ub8EhwwwLKG4Wc9wwwIUyY9XqJpYJ0IdhVyjevH
xGsYPcajr1y6Iz6zVzexgG5LG+2YdL050E1XVxHh6bEilnIDKkDryPy0dAvxQnxBC2UiKsm9zQlF
L6Iu3lM/jN3J7h/qkET3DvwlNYKCfmV0kILBfFHYH3wQ/PsWA4BEdVDieypkwGm/dR3Bj0nOLlk4
FPBgsFyyWSrOnTI13Q0ANwmTwSwEQouszf3KpQofPb+3fBZp4nDDiTdKS0ApTDwB0R4H8NjZemNs
gJpVocLLOVV5+wvx7Qt07T6WSG6nZvjjtK96rHS9rtbJN5jFnGyqIDZRiBJaNY83twqyoEyUNAVu
pU4dYYYNKnXgLHVNEbtCOBjk5GOv0gvEZOXZa2CQihknHjSGclNhhpN7+Bt4PG7gb4dwZxqSAfiz
s+p+Ve2oxsWkF0sUzh+Nd5iC2lBTDXKkBtwmFeeQ5PJ2ShxLqfio6EpAxvYroEdhkFSTImyPjX/2
+snPctljFg81lsaTSkLOi+YwIp9N5cw9MEY97en1KCtDUPDi0Y5fxu1pyGAsy2boxUMebaK9YQyD
l07ne2jEPwc0MZB4KPJTYX/4NTrF7dHHn5lNC+eYaLI/NudLYJFpZ5d2PX1zd6ZbuoIaxx+dgX78
PhpgDmBRBuudzk0GQkAIuZsyo6erjKDp1O58QRLzSoK6qQ9aoKeGqy7uLZIa+AKMlzakHqOJUYA4
zPgcGfFFy4sxU5mssxZedpFlzz2WXevx8aTeRLr7hQoKQUoD1yLdPWCMqWkDic8sDt/6WWMH7IEp
ocHFKwGvNlCb97pE43af3RQ0tjwphw4HBVtsyBVAYuJ+jfo2rk7AKCHM4HkJb9Jr2dxzbv6NKvaX
4DAdxXTtMivY9I0EBiHjvFlL+bDM1fNXd9BOwoaBywf0GoTCioxVCUv0a2O4M5O9YkYYKUpWBJ5q
BG+t4zr4gAGAjdgYlEyv2WmnxfNEKHpDIOMfzeLMAza53gOBdOPHF6Difi/pZOr+vsRpN+KtVfAD
21kCQU2ArcK/0AynFB7EpBrxFdjTIT3sIXdxd0qZMxuDYg04sHHeObEh5lTm/iF4dIiR6J6m/tX3
9xEW+9EeEOCsEv0oDSRPg7oRWD1YxxCTgl5TH94g5BIIT10VQ/aE4NJvVoV1rY2kpmTAR/Llphe2
vJzOd2xa4jKvvjFUMkChbg3u82PU9Ob9ry8ijnTp01xMR7FVLZifilW22FXYsICJHldU4yLnCe+n
F0WbwRfff+90tisJhHCu5Of3kCfBFHjY+45z0O+REGt5NGQu1pidcWyHYy09eS03yMyVP1sdq8Rq
n5pCxes9d+d1qkbslkXhKD63h8jimTrCSF+0YaI9sabtT0nvfSDm08xwoZMXdl9rkARMWZ88Awk8
5QHvJsULQW11DPGSpWy0SOftbUMLiuGI+f2sZO3AZRxFz0z65ODMpa7DGuhsS8YEwtlMWS5e3t1b
lcdeH3S8OwDS6Q/QRn/yqU6J3AquNJ4K7rwV1WeyTkjVFprJRLMn/i5ZodYKKoyLSp6eJWm9sMZs
GjDsFkiW3lCEPG6g9O8oWImEUJhhVSyV87UoCrPEtm+VLuDyUbxIAFuRKrjY4WHEviUIN5mnZXP6
cMC6oLx0YLfq8F8M7aHTW0o4r2/X7evjoQtCmrH2sS6Nj0YuphRQcpEIHnPYCIj7HTAdngAZ2vsd
oVdCFNLMcd66BjdHltwnAKG49CCV0jwCzqzReruRM4aGbwqHDcAM2UznRgadBAGP2oLhIa99eUqB
34c46MmLlnaqlUEdopOVS/LQe9OZI8P4DXxoNaA2anF/iD6n1DQz9+HT+o9gzTsMNtyrA4mUwXfd
P8njxmumxqN31WGf5vRfUY47qi05eMDkFwcKj8yotQQfYdVw0fQ0kK02fsXi7jBDahWNzuL1BzOT
DNaGcbXtI524jKNgcsbJdnsk889NYCf1POLeqLxxFtisnM8UEqyCffvG3m5m6iQT6MpyIwwRbZ2r
TfUrXA4qXvpRbCaSAOlR+nMOMR3DP98+2SGPQTHCVOT8rATI6T5eG4pQnpOj2r3IR5UAsmfediDY
iOnBu+KfFoAlRI+XSrC8RfXs8C/w2Rj6WJhQ3aXQs2tCGbObOzQALXW0nRpieVZMdaSOUGDaBjOq
i1Rr3pDKnTsx+h60U9YxEh85FBn9B8nDPMf0R9H+H6ib76O5ESEz1Qdu+f7hre6HuRTvoCYVRdIP
1CZ3uuMlOe817t2Nwed4R78n8qMNQzD2q8qPPjTOyE73NMl1EHsjPE0ijX+E8p2XSUVi7aWtPcuy
zpi0n3G1eymxBokZoLP/RSYIstFaYQ5JpE4TSembrsn8VAB+ObfvmCQBXEHkgg8SSu0M8PJ8UkOV
BdOeaW9bh2V4nS7GgBqwO3RVzkZa64Wcx1EmyCcqdYkJK19eH0uk6wJAPAGIP9ejOVVcdJ2VZq84
KpFNdDgNSSeNzXaQH+ngthoowuNtKhA07ONV9UkQFOmACs1XMxeFtFH9+XzQJ2ECa01ds1wrJUvv
tOxlorI4xbJh88ptWNBRcLYvQG9Ske2QbqiRdFD85E4yEAU5qJU8Oicrq6/NsGR6RKJB1miIWMWz
kDCX0X1aSfVzH2ezIDuFuhbIWNR49CeXw83bRMZjScqATsfjxkDewUK4o/Pd51b36nXhR7Ho580V
g8gY+5c3Cwab6c2j3HOUEs9a6MBWgU6QlFE2uaR/XBbomh3sULzEGIVbE/7eOSC67LCKg+qZciM9
mYmCTe+E2U8sBRFPzVRNPUfdaNHyhHZfEBid/z03GpbS1I5fiIfhX1IksKxcvuGym6Tof76mQpML
OoVMq/D3GYOGVkQxWx22NN/6dQviAQh/J3/TCnapmUdKi09rztLb4gjvwfQD+9S799HfN9egZc0Z
sKuBFL0ggkmLma2yhEH1GgCqnVf5EyncjCVGIB/btyaYUfid8mq8Af5QE4IXxdW2dTsbGUKRCrJX
j8kqg+FeaAiDQllHzEElntGbMwGuC+ihQttCRa244S3AOhAl8aJ/L/fR8a7lglOsxBSOzI+WELfd
jus6aaQNz4hEO+s3VaB8iupjl8WJuO4+lQ+EvTqcUSlv4D5BiR7ItteZnm23adppL94xfWMZTnVJ
4sh4pN+jFe3XV4+ybm7but/BU5ISws/Lu+9LYgkEwyKgLjQtJ5a6vbAufnjj1Twi0ePhDm4GSCwd
QK320lokqQj1I3tc8puV/JJHCKa0758H9yFtSugUUJJ2e4QwxVmjxgBTkjpZyJePiOaJjYGKNaFI
AyiSQK54opirXpOZRF6RHFJkngDaUk3RGtP6dWmYW6SYV8mDYIxQq7758ARd7t5EkWz97kW/9Hvz
sGiulojJvAnykafmovxnZ7jq3uU4FNXErtNHC31Zm0TbYonoUBv18RFOET4tPda/yTUtXwVs92S7
fgnOhi5AAfeiDrkrM9ljMsoW3pzwr6mf5SY6friJaBE+g+dTKAmgUV0DBs1Dm+VLiug1iYYSxMVW
AzaFktBJrgopXI1CMMn56S1oVDB4iBzqPmh/cxpz8xlYrMunWpMi4k2EKIqwBj9FlzhTPo7PtF5h
eFNS8oekoSpewBMVb2faVM3mFhWjv8GJefIWCtZtLZFh+WeheJrCiQZy13OLVrggQe9aBxBolik+
ntrFHq96kAlGl1xrlGeITxpVrxPb2wRDuAIvddVOfiP5CcZCKGDle8/9VGT3gD/KYatKJCBJRlQN
opKaz3p3LqKMH2c4R6U5Ewvqz4s6RGue7FpjfMfFBHXPys6wli6GRh7CcuDumeQMvm2a/PCCgiex
S/2s1ehg1Y85LO1gV7RUP4z2x0yW9Fvj+E4UsqacElIo0/Xu8iwmhos3JA15Sc4XcAr8lOia0X5y
TbcvWW0UUZuiSFLzGacBkX2RAq9Wi/VnjdZQItzlzr2vkSO1eGN88ISG1dzic2MiZeUSZv0YJY3T
n3n1PE891KZT4vRAc1fmm3F0HwQfKbJZgudAFSu3PCylPgWeAQoHKcDdsQj3RWa8FtNpCK5kj8WV
AtkjciWN9BOLoGDIn10TaFEUYeDf1SWp96g3s3OZ54RvkgSdSiiz09/9AcFrlWpsBXlrTi9lK7SV
nXoZCDWSXctEFVUL3kG+/Rzu3k9Xz1M+ai6wWKWdqPfuLdYzmg4N781+0MPZzRVlJlz2sEBXbxax
+H5Bl9Ws6bLOaIPoG6l3eVz86yCXFchceCmYozyqS101dFyws3sU6Gn2XW8h0Ha4OXbr/I7w33F4
c+Ttm+RIr7Z4Xy4B5DTVy45xjE5Zx6DzNwOX/PVtGqV0K5cP2mBeKTtxD4eqOFix+s/1n34Utmbk
CAwIxLvw0E7CAD3bjcglrAbC+H9wodgjJ6Qk9IFISCYHqoN68xZi0xxouJXchpNYP7IzjFsgowmp
LFt8baqRfdFSJ81RiTC8dmIkhX3/e+jZoCcI0pC6Kn3IWiNayMgDvb1N4di1n3SYYR1eXwuyQa0T
KZbqlnJ2zi5Zqk8KAr9uvo5kWKHn+KkMs+gHNznChBfsLSHMM5JndKn+XPFDNBMzEIy6yZM4RhV9
xi0nqawmpfQEVkbnFOvtEM9K7vOOhcaWXTfxIBGvwb1CLUNt9FGl9GgNGgnz+rQl82zvHe6G0VyL
mrRDH9NRfMuo6RZ+kPzCoYTG601cVDvlGlpPKIFHSnHiMGUG+K5X/8RG3+5/1vwlNbUvbnj23WbW
X/J79Qd9hGykPg6gF7/fHx3PXQXw6Fq5YiV3ILmiUnrlG7FpWxTy7Yv/UsNS36eHoijG22aZAOsC
5/ff/7RhnzTqj8JJYg0sckQb4AwWUVa06ZagHfAEGQ5mHo0GhN08jveH3mSyr+IhaUrGmngeySEB
kCm73DJ6kQSrNYP7VIVYhgwgORFfINl4TXUV0pPixO+GQIGd8lH2bGmkp732gCNj8w3eXtUOcghR
fDJ41LgOxS49SX/zVEfS1A65LziornOvNO97c7XQEpFUW8H5YGs5UU60gty1NCE6E3+cj6pcFKVG
yCMMMxLZCGTmERDvvRiujpW78RbrIku7JgO8mLFpNSB2+iolziJQLP3NOSjOKlIL1o0J63+EUFSc
9W7ABX46tE0gEo8IHNMEgute53JR+BtZpvfiCM88vSpp/lJ7IgufxHQ8fwnghh5K3TiZoofet8Lz
BViX8mqAVyabjyYHAD0NJZ1mMhnbU6QYw4LCFFl7relgizfjlBoK+pjAbvmJUwGdT6Nj+6Cvy+9m
4HhqCEOL8S4/bEWFgLggEAQ8ckcE/K5gO6+QcTgaPFJ5UHWvqnnK8Uy/DpF3X0CSx7u1zvn9LCt0
WRRvoXeNNy0pxAxDvFQ6FOmzxDFz11MBFcEW/orkZOQM6YwkKHgQxsWTgT/kXjycbAv32gxRO0nn
H3jfJRyJZnomTX062w+q++aYwDCnVefYvH0mr+8SmKieDYlznvDLxmEtPygrbt+0TpYsZHyJnyo+
NEQg4KTtjYuLkaGR+Zxlk0M40aRePypokdWtVvlY8qX7AK/1IY/Vwh7xmbUivGtfh4QMsUlSNZTp
byFS/Aon4Ydc6hx01kegoQxz3sI9WroodmkQr6QLZ5VEam1NoniA4gTELfnlXxhvQ2yoMGSXwXQm
hgGZBujxP+nz7bJmJh1y5ncyeksG+Urp0fIPJqnflxhuWinYZzmErQhGngWbff660qk+NtgmsnNg
oDPGThZWXZY4vj3/G2PvHQPLmyRuhcc1dYGY+KkNslenN+xLm1px8zG+Yn8PhCc009zjw9+BqhSN
XO6xAQ47Nf36sU1LczErK4DL/H7N8Nck1q/+CZ8iZs08PQ1WQno7MsYyQcVBcxYkv1HSqbakRjto
xF4Y64zX1vYJYkknguIDcw3rLgqtHiIsdaeBDtat6Vw4y1VDPEk1e9bv8obTHgvcjpiNBh76T739
415iEk1Uai0uFZu/UzrYSdnhvFunpVCAVQp5RX5o2Vo67Kw15aPI2lwuChAN4u+yam05O7pjPpzk
ke9aZFAaiMQvRUHUPru0MsvBTaZZAsLLKwtxummPTH+AdDkUgJfxP2soZ9T8J/T9yxwx5W0Bw7mG
BMW3NFytS9a4Ou3PCqLMaMXeM3h2FIQ9jgmEFjxq+x+EWKnLn5enkayQ2q8F+Ny+M019UGvLgjIf
vVJOeLZqDOM6PBkKaoG+fdNJX58Oe3eG+k6V5mcRgQIy9K5ZvBvDPamx1JOoo2VsYhxGsNQELUyV
Jp8vM3Ra0qLA2zh4sJoybjKjEuVdd9mcOoLnFpQs3erukDBsuR0NyNJLDPXODpPsjE/DylY43rQ8
1pWOkjDaGvinO1L3e8kk4LNO8VoTmI7S57cXqlKw29XWMbyjlcIlkHqJmuQLZpl7vzCRrjQzPSBM
SEl1ghmbLXYPWTGWFS3M82Mcdhmk8sZQckT3emn30/hDySUQSxsYjPU90mn8BbE4FBWTdhE3U8z5
9deBY04p4lOSUafkK49krWtKwdFIqETYLzqsDQuVRRwtunlsHGtWgZ/jxgiWB41svOffZTJal+l0
FcBc/NIOYAKvmQg9Uzcj6cUy/afjTS8VyJYZMEdyaIrMNnhz/XaK/FfoAeiii3EMIWzbpAVfaP8h
8n4SBIUiOtDU1vEs503c5whGhw1Ag822tuKS89Yr9YBmHTss1ycyIRUcHyqUtNiQxkCeBMJF1ctS
cA/PpNWUo+Lag4tqOtpGNzQAuVXIM6qU+uOnwEZPKng+uu08Yws+sb9S4XF+PVJsuYv/4vFGEvio
rGNg/MGzYdTxJkE3AHrTcZmToicDVcbJG+dCZpivJ20UsudPkiXAAbaQPx5pwe3ZAVJuucshA+2L
VOrlo0or4mMglHEFeNHt/sRGc6MVEseAGcp/rLwje5A/c+Lmlzy1pTAYxUycJ1lqlCXHucTCPDW9
6cE2DwXUotKSEWgtYyetqL5mjQjPxExDkDQuVJZFqcJ+GQ3cFuJdwAb2a6CpyksppFOXj4dXANfn
fTL76BoeK/PJScWh541jdunvGtbelkBnSH2HO9ej3ncGYkoWaKsuAbNAMzvhiaCJl8q6MbfmyywI
qqrXavyLC7nG6lk9TUT2BlsbONrrDZ/atS1F139Hu+DsMDAYJNq+ClrDOyJVHyLll/Gy5T0FLrjD
oSxZgGldUTjkcVbCy0TV81XcuEXSlgEt7+IkHrB0YS7MPZzX7jMRb/2n1LYfte81qpx34mkOTPcW
WlNc5bBgF6GLwsDrJhNY3pX3UduzxG5FhstSI5Ze0PJJakXHlTsRGke7HdbzVv8qBzaZBNsLcJ45
/9/cWJa1SdoOSEBbw864QE8GPIiH+EwR+dodV3lXCpHnDe6lTheRt2EvpxHjY0TsDjYp682oVM7u
dWztHiVVh0tglWnJnAe7t6/VODpjKHxa+C+mBpRPDgewzL4qMtEesSsla6koNRP8jYo2SHvtojkf
Lsqyc/6PJe5MmIhZJYJLVy7gYnYVdLPOpC/WjTx45l9I1xaOkrS84QutO1TRkFtMA5d+zsQC9BL/
MJ/DJmezC0tJrmqDE3g7YrHms0tatYyGOf7ePi2Pki6aLUMtsGNeakcUupRguq5m5DN9YXfDQF53
T2951DVPyfVZc4qlf6KhnkmhMiVUtGcQSDhK4Jx7iOlcTZtfjnfVZ3xXwSQNecBq5b3aiTgzLUAR
2aOXQx5qA9sl9C8Rjbqod0oAywTESgfAFMQ/cDEpyQ6z8c++UNDXgYK1+ujxg1esg+TvZwOB4ebj
e75rkQDVhkl5pjIl4DQEcpD/e4sPwcOlVJQNTnCsr0SRuVEwRIo1GGPJUl67lMf9FA9o7RPcpLFb
KEjRAhhQiw+L/QHNB65VuPty5/0hWBk+/b5MZMNEX510zutOo+RQRFEvLMdOdj4gY4AMFo+I3NEX
RtUcVmTLOto0LmgosZNtEGNVGjxjysY3fUh6TFYhCPf1Arwso3iPuPM08YFpg/OrnH/CmyG/xLH6
IuftK9R8KWsTHkZuQoyDDNmWtz17sLJGVXYlzbdk+kfTJSJBUQt83jrdy+oSlTGanqcSbPg/Rb6E
EBpgvwD5wmDzWQ6IU7NsVUQuZDrLsQkaabtLd85nCByG6YgzJdvGLP+bb5/whKlQUie2EBUHNaCu
9byeSnii3X1dIktDx5Bp4mm0tjvA0tzcG9eDBguWVWgbcVEx7NtvdT8OiLMvWXlGU3vUm5+ahRZI
bptRmJZV724ooNH0inAYifZq2ifTQv4Tp8KAByueTpe1T+fHD1ulv2eo0lfRC3NoGliXX3GPgV3g
V3xyLREAHZ4C8wpygNo6oIbYwMGax+EVub8LGtV2jOtqo/ymuilZ2CCVrUS0bSxof2rz69w2ig9B
YxsJULkpUJ2oDUV/uxurC/Hovp0b9yLHu9bZyKiy//CvSXVgQSH1+/YpSaRGOP9Oul0j+3+YKTwi
e4SyU8WONFiihiXkBbsx/3mOSnA9MDqSIYMSF432zllrjUHLuX/Kg1GwUTcUX9H0gcjuKiOVqLTq
ZgmN0Rhrt0v7bmvjjG9UxRG/Gkrezo51qvA/Jc2yWg97UzG3uqgv95iM9FNnvKNWlUGSAeQCvvT+
ap06fQcgy+d4EXdIOZ5U0xIJ79Ls16IM01Fy/++Ng/MkVd8pb04oU62BFEoOZdPqQEekxc94W89H
5d7jXVm8SqI5YiwG4m8wBckPbYXfmwYgAs/vIDLOx/2cFmR59bYNTqN8z1RiOjpVeM3hjyYE61IV
3oYpHAabBVTBXdXF2dSp0oK4OLoW8IsmcSCcgUehTq3QKBH1+X9W1+f75uai1lgyrVM0MSKCJPkb
9hv9WImUrhXNWktG5Du92YBD4C8DnijYvkKro+PbL2LoJcIYzLNE8Rf1ecBRJcfCUAw8hASngzDx
jexAJWiWpR3CsoCmthtigTpKiTFZRTFb20rlwopTVxqYLH5VhK4hsrJip3krQisMW05xDAZrjve+
BiyK83y+aK0R2EZRoxsQFQNto6PAa5NJpNVoR3fC7eHR1xbzQDoPbKerc3WKAYRkO2IgHCxG20Gl
U7kvWP9P1v3MCM11W5gA3GINC3uRmZraRBnI7gUv3udPrd5kUllXfJqqfMxFMtSErFdy0nTadXQ7
TLA6u0+S6eE8C2U7ZDyAFtEkTUmhcYKogbHlEGsgx/4tgNEYUBT4m8ZVkoWCZBR/kNYzK5Qd9vuH
E0rx01tO2mH4C8M7LQELi1+W6sQ46gjTLM2o2rYW7ig3yZLTb8ex8GUkWsgVQsNnQ00rjoWxXlCd
AgcmlnSx8iMdw2UvO42L3E8BRLwYJvGaNZlUY7NWiMKWoFz2w9R4j95Bg6WfRA8lTp6VO0lsWQdC
cXa3NBZQH2vO6/ze+YG6nWHAbX1goXS8Mk7hHX9VqbHTwAe9pY0/4VgC/GnnUW6UMxzDMnj9/Pwc
lLPRK4undtoJpiS0G9j8m/PzplmjRdSaXdxy2pyq6LZ+BvRACjdt4Wiikud4ks9kQ9AQNzNewDTR
JlkskTuAtIme0PLYrt+yGFhteQ61+5amsL4oXmIFuZCI3sJ7OQOETIUGg9RYBAgNnPIag8rQIQ2h
ZY++zAOWbd5bUSrW1f3la7mpG6fizholrboht5gzV5lAsLNSMaAuLQIS+Qf6iDy7aQNSxPKJgT+Q
T8aPnshZk/SEa5BuWt9uOPEyUZSbfZM9DKLQODd8elKTE0wTJeHmFOBf2S87BmXfxLly/GL0O5Iv
HBpH82sQm8OfHvyHNzR9//BScSmB1aZGPXXyV2mik14fYOSdNuFNpOi0Z0vVN0Z/nfpxM03b2mOS
/ktfoa6nbUDB48vCjhA6U65edxhCX8uLsWuJGH6z8mNzg52YeQHYpYdN5gVJ4N4k/KxR5DljcXAm
z6FQmB65TlKpNRXZqjGnThOI1Xbb+t7h0/2ZqBt9nSiUr2egJ3aKZvc1ZE2Rp5sH4/9/jxZfZA5e
w1WcYUdD2Ts/gs1df97ZCsqfICAu5TzlWDDkd7eVnIcgJLETnmpGq8iqfTkbKDF7Kqc0s9TM6BVw
O2QAXSfmJBOGlQNgJTmJqt8hInyyZJ5L2FimpeNerGo0yaXiCIcPZPUiOx1/1QU/jjzm1Liq7r0b
xK1Gl5No70sMQ1Jz3zR4bMSwfP8KKcYJlazk4tWr2A7y/BewJLm/UeMrGSbXvPE3wgZNhhj4VwSb
ANi4UIqYoIYmCAJ5d5JXwSFaEFcXTMZ1qTbMK/XJNlIUYbimKxVyS4X2Xem7rdVbkoS1Z5tPrYy4
KlOSfE0jVdhq5nwPyIa4i5D02a7q0n+1QiHFkEC1C09QvcOx0fc9NWbEEQ8xTdmeGGIZTJFKivjc
NimKpy9LEB964sC1kPn3IhmaeGdKPfhk3ONGuPhKwTLcqHWPWKdIMNCi6mskVEdGyBS0+FqVxwkt
5YP5/XJohzJyQOt0Dd3k+Hq1dkWM+XuH/ytSmH6Et50KxypdYU6mLuiV+Tr8SF6bnYMWt7ZY+K8c
byrlyiy+3EeYK/J02zMOKgqYoe2Cn6hfGyMIReZ34rQQNrWuFsaeFF+iEnVwTN51LYGCeVHkzF3A
ft/iLLxsjpWqoDU+6E51cYQUkUogj1csAEmBVH+LDXuoTBa47S45jeR575iERWpqAdMLZtsgu9QF
vmV5ZNyHw4M4FuxEzAbi2Y/RpDscbpIGByNYhKsb8QkbpRT5R80Sf78uh3T1WXIe8m9xRPw56Oyb
a+S+GUpNO9mvYtZ5wBw5pVKZyKa9g9M014BhPkolJ7ohgaddeEU1fDlCekn3s0nw99w8s791R9ge
fwZRtJWTkJZrgENW7aFi4AyPvhYsbzmc4PbgLnpUdVFDFr1YCCIxMeNMTuaooon3A+1WG29Fu1cH
OG/lS9bFzbIHBxLt5pCj1t2KTKZhu7pBieIIGwvTmPLQnAOI3rpE8E3uMSru3vxa9PBarx/7DCeO
RF3sI38Sf8W+oECJ0OvE9VUNcqupW7NE9UCXNvvv+WJcMG+lsPMNkrrVQk9RubSPcuhclifwa46d
9H4J490Yh2FFRJg2wxiH0TZMt1ZgQIe1Dat/IWEACf/mZMebGNLImVmM0AoE3Wr9FfkRvyDBk/TS
l7ouc0IdC/LP1p2PNa1A8Wbr42y1nBHlumY+Vx5n801ckFPrHMOK9U1nQFbwDajdFsSGCNR/34uT
EupQjI6LsI7tXDD8lgo4hhVS2wkSsOwcxZ1I72C63sPjintQO9jXXUe/V1dnFW6uIOAc0Nt2W4+M
T0murq5OunNkFbMSfoRLArEpnxPoQk3nu1Z9jtbdYW9WUgvXRvB7rzWvS4xbD+05WtmpwIXxUtxM
QqQjUVfVYOv1g0NYfQimFaDJRJtIDSZ3svUjbA2/qjsAfdJ4JGuXXXiSg1gfVXF7N4NkVOjmAyC9
x16znLaXy8NsUqeDa234Dj46js1caWVraC6XcVpDMaZJS6x3lI6Eej9LdZmRfP9/l34SggeYLwXc
jjIewZ7rajUSJZ+T1uHqcOcClR8Bpg0yM+/I1sv0PfiDskVsvZ/h3cGswFyADGyugk4MZ8yzByQg
E07tcvSyIyWCcIJCH9eSBbQsomf+5NEzchpjDrZmimQIdHI/7YA50zihAw9oi/qKZ2BTUGemj+k5
JoS/oORFRckq8BlHVl5WoIM0ZTnfphhnM5VbhsKpv5IwO0G2nRwCDx0y2VG64ltyo3jkFl+Pa6Xt
8LrFbYPa5uY21rQ7FWgvnqTc4KwtrfZJu2cVvd9DZ1ZKdEUXjAzQ/QtXZGYFQXncKbQzVJWInphR
gyXtPiAl3BGyuQS2DLaDD8RnRQ73Jy01Oj1amNcFZeAMl93XQUjbluxkL6igvX1YMgA/Agw1Zjmz
9w3s7WlqH8JhJInWJcH4Ue4xPCWxL9jRc8Ibzok9Q4TtWQa1fO0bQYPOUNenX9TRzHBjvuyyygOs
bFWaGTvrKc6XbukCU8C1vdBu58XwD7DRpgylA4HZuTU/XSF0dBZCcmavt899LvK9BBwI0Lm9aeO3
GoDoI9ol4ZfjuSJ0Qo39qEZT7TRkpMdgmwJIQU+eE0rVftVl2EF+NBk37hLTP5nqHZxFt47hN9za
ECmvf0aZodr3CPIOBfJUdcCyTQayb4zKkw0gZJgXFYjpBhaegQHaT3+GfhdSAYT473KkqwFfaUoY
uiL6rPo0hah7dArGWTpeVJ7xWqukVUxYKDj7C4f6OhLny1YfEqsiw92WBH/yqp+beW2zAKz5iHZl
IkdZxzCeQIz2Ae3QtLvezjoHknywyx2CSazqSd40HxIZQ05C+36BwRla13shtyeZ2PG8gUrkqf5R
gysb2dO5pReEzR91mkwFBg3LGSvklP5fv/t3KswwvmMBkfk9LM/xK5JIVqLaFvvvz+IfeKBVOp5a
nogkJdq4bpfNkYdBWX6J+zJk19Ol+uLyAIZaC1ZShO9lV9zZ9/Rqwn8qAYMX/kWf9wy3GaPIL+B5
Ar9ZH/qhA70Y/2XgkFIVizd2PmK9XGanaIPzR+vdkGc46/nPnxYV8NRgbUVPIUCvN/MSR3DRLwg+
WcjnQCwY5udEOlCygiFqLd66Yt14xlbGTwuYIBgS/XLPMH/8FhU/NrRdJ6JB0Z9mQhzaWY79ZGO9
+Zg42WvoaTdxCybvzY6imh1waco5XIP1RXMN0N0aPRC2oJkHOyRFw6R3gSCtyRruveBI8YhdCAwU
hUvTVsRc15+8RI+NZfpXagyZYUqkd9twa24Q/NBFWq8aHW6AhQK+dsbQnoxcDhVTdmhNlOa9QQU3
eu4kmhQi5ROrHK4PLa6W9feakLNN1Uvav7QisBNnRpBJ6RyU//kpCqVO6qeE9lbeUjDBnUxCDO1G
dOor2CEy7wZ8BiC3G4FBrZKgrNc8Wenhv7E+W+hswSaamZp+41CFOL0RUvUV4DyJRLw9KxXf8Owo
MTk3YahPE8KteLlQJjgCiNzkdve1GnOMoaUdMeB3hsTtZxdSQ+qZYF0zrcp0/zcp5cD07chYYlbf
FutYFUF/8aACM4Lzrp1LtgSHP9+eL4bhfJ4ZkOtTAsJ2xQ1uch4o/yIQwLAXjBNggb/5QM0dn/Eg
wrF0cGGHMZerBzaLHQOiShR8VBii66yiDk8IABfrOXIzCaBEsEWvWSSMj85Az4IpPFULB2YQ73Zq
nvpgIIVLALxHvdcG2wSXsT5OOGF1G/12i7NOm5nRg21z802bG66tC2TEsdbzB/3CJlNa4R/eomlH
a0L6rtex31rKPmA5raC1+z1d2AQUmzGVrPxm74wGpNR4fJw9dHk+cHtSaUlP98d0YnYprXMfzY7D
CpgCzs4/qVh2Tt8iIgAxfoi6+v2M0bisJE5dXC43KVfH8f9o/yinFseDKh2uAIuZn1Hf/cAocNzj
tCslkoEXTZRZmg2dPtnVPTyVj0TZkw8N+J6mamkzpv7+K7UXdJs+wkmIxJU4+kmLaNOwd4ipV8Zu
xIf+HnyPIxV7EREy+b/5PyiyOiyINcmfBprm7MvPQ+fVt8tKVgXX/1mVFUYHtFTujCmzD+Id+37k
XjkW4Vw3u7i2BusQAjKDV53mmAvIiRK0qY9PlguZnps6HZT1xA1Ddg9gRE2TEZAeP100FagYZ1aW
vC9RgyB3SyUS+VNc6pu5/zILIyBHt4W15j0p1WqDy+CWPJpN5gK4kJKXxVYruAfc9eAr/va+muCs
vGhFNJcloof1LOOADm4o/4sjv3Vi9ZK3RULxN0DHoGBAi0TxnqHAutTcZrljyEE8kx1EiTJRmfyo
5mmfO/j8eH3eTN1t8qKzUcQsYyHqZkrucdufMAFkj/mwf39ubJryCEpCe04PRVjTchjl8dDniVqO
8GxRVOa2ZZHXteQz2fMQJi2nl7Q2Y04LPIHonAiFy6Eiro3/Is6cDocP7UIKqR2TeaBe3Q4jSNq7
RUs717rOvZQH8NuFQx2KswwWgmkhsBoiCa87HGYagUtembFn9Ft+ptoDfeYO2UTWhn8O37npAwB9
x3P+YEic7jeQ0OI36r5odMlSobHWPdjAJ+4z7iJFAmeBOXA/ZSOVWqB33udNzmmZ8z8RF0x+JY+O
jm5N70a+A90pc7iAEwyvtsdTVHupEEmItHZSWMyMfd8S0rCF0Pv37w8lvJ6x/RKsxMJpJFeC45xQ
rj924M0KSwp/pp1JOUOtxmVcFIE8tFbg1UEWTC3Qq4/VFiS30cz8CmRw8LoQUzZL9m+LG8gLGuM2
Qfz/0R+VFUb7wsRorfX4rOqvL+VcLHSdBNWpkGtmSW9nCgd2IZR6gnLbp/SmxFReFsUoeI3/CwHM
zD4GE8/GH63wwRYNpVpOjvDIMe8QV/O9fYc9AuV99r6NP+9T9XpcKZXAe8iCV/NiSzxg/bTXq2BO
h/+RqKBvZiwnCKUnvw5DeCReMkUu2OSC2HsbS4QXlsvknwVE7K75KSH0dyGlmrpJaBg4iHT037Gz
xeJVnsncah0dw55BlUFjCA+jkHhmGx08Fi7kq5Rx9dRMvgtVlalMH4HuyIHvw2Tu7zQZoJ61E6nn
9jPWV4qz/otlpbmNP8umq00hoEGTkK8ekm+vOIQ2huzeU6rVyZQwbH1BCVDjAM7AXir8JOvAgBGj
MpvBzBG30QZhwWDiv23Ru4sLKp8RUEoieTZ927sJAPXczsGezIARNb1ZEvnbNu2adhm8phsBZe9E
57tW8rm55tS+qmEEWNb655GjLktjL6QseibWd/+IS1Nq/0MzeFPwPNlMp5FxOteYLlfc5BQflm8P
SoRZBRl9jvmNuCvoSYfxDxd0fngYxFPPpSOVCQAo9OLxZykQOvgpuKLd/ooO23+BXLShumT1dqRV
kLEm2uGmV1hIjvign3ySeqU/YW0I6gSvTWuaOioFI88X5ZQvB+fFmV/BUh8/IuI8GxJ4NNw3xR/2
zWU6YFGi//Lt0XHIj9ie/l5V8rnveT+Ijl8p9g5jbpf7wlsJIDsL+7PqNYMDEnRVSt5gwf/amP6N
ydw0QPgMQXTyM+QkdZqeOe+SYeq1EcYd3l1hvvCRXfgGF8VFE4wt3kpfF05xkHoFLECSaktp9fg9
a1ML4QYEpIe126aAOzX9CTf42tRQbLpeAfPjc2AWqiBiEq+k5igKXdAi6mBRHk5U5J3UtjI68h8F
zt5ijJN923EQektM5dB7Eq35CSJzZq60hxKIY8tdSYcWHFc3FQSY7BmAErbnbrd4XqldUTLWx9Op
BttX2B7cF7mHibPN3cm4j6lHQNcIYS2B7QiYcXp42ETH6i5NydZNYqAIdUEsUrA8JGz+/J0hiXFm
HZr8BAmy9GGH0Yc+PxBD4DDJwqmWxrRAlUl3M6H3ZoHXVfYnRdPpQNiR6vLH9n/XjSnWT6rNaSch
3weNxxzeKwKyzRxUrqhRnDfLeEjHGtO2qTkBXdiDOiTKE04w8ADi/BPEi8dkeb9Q3B7BC6Vr1FQd
GTVp2iDAk+1X9fc/XbglwHjcsDl2uv531VOhDHDVezUpy6wuiEhOmd5k8fCjna/ND9j6gozkxsUf
N7JwQmAET2FRKiYCKlqvKoIfoWqMMjrJ73vhUEoXE5QiI6rPJZ1XV0hVy5GgbtATElQ2j3u8AfqJ
Krtoq11vstdDFp4TVfner7D/WkI7ZxSBmh8kkIzlrWMkfnnMTCMX5isTD2RtCl80ooxZOZC8kZoY
B99xtd9bn0DPy1mQW63/UtSmy172WAR1Ma6bump2yCpf4XMdutchHqMAfsG3Z4B8wOtAZCO54YIb
M4PVZhZXZK8qrZEwpJWJ3/mgqGt5pGQ3zk07a6w0lujF8oo8qL8gDIoKQTaNMo3h0/ZjSo1GhVqk
BP+DeRSDqHg7rRLJuamPFBBM2cwd2N3SeI7ORCpBOI+j2ryN0eazjS6RW4JeZv19tj8V3l1tAYQd
Qn1W0hAM+0eudEaq/ZjryWSe9QGhaegz1MBJFN2lLjEsZCqIVDDZDdQPS4T6L9MoBccjWBkDVVaS
FQVtBexmIgZuBHaLx/F0OxVZIy9RBpQrG2xukuDrVBB5gInNqJVKoFd7kn57E7qQdVb6Cn6lCgbG
4ylOb5kPQD4JUKxiPNkNwABiiIiWe05Q6+2hzXKXFnFT0Mdy1RjFck35Np+MkDRSjKI4CCkYTHAS
Bega/lwUtVOOPbZFvi4HveunKplXATnZAqHzV4zt6+i3oabHw/6T0g4hvsFD0zLWl+QoRZ38su3E
6cc10v3cDKQ4wMSUR6rL92NBzMN+LeEpcKWNSJ2yqt7ZrpkDt1TL4Hdp1P+p/Fu2HbrybNxWF8VG
2+/FUReFHLgKCE7xoN1TvB6bH6e7vb00Syk3IH3uofkSyLhZ3D4Ki3aQaKP32zv7exCPyDm+7ohl
7pLpoWS6SJCFeaOi3bmzif92LWyZhNt3rz9egtSKU9ESJcqlMJWlsVm7nnzAe6qxk5PN+0i69Oda
atYNDMrG4sS4M/yKdMvKs6kAxs6XNz0yd25Q5Q5xvgjtYZuu3Sn970h9nLZAbC4GWBAWH7NUQUf/
0t6BgrQCXXg3xA56xWr6NR1JC+UrbQDo9mxRtoacTLJ6lI4pp60kfzkjhO2NuHL6Z8/qkhGEbWoP
DJ93xe+cJ6PY7gxyVswRAgh8Wd4B8TS2FuNfjf1ggvIl2WtoTQuFNuDIrSEO+JFLbHfq8VTn6/j+
FGbtrQzkybTnSXAMZrSmIYAExschhsCiUdY079owxIZdZ9+KmLavTduLc8CIY5xgjX+V6Kg1E0s1
WQ77UGZUmJa7bfR53u/6tIc7yWZ+89e7F2wU7eEZhBOg8HL6tzhwFTe1BSAriusZu4YNVXXCeOsP
MwMwkN0yykiQk6l208OpbzMW29HcqQALgdTYX+5Z1vpwFQzsHqZ0GGaBX9PecbtJvz16ivHQ3HtB
DsEcRD6w180EemYwcjnrv1wfoz52SHsGN7svsl7ToqiBh+IGb88RBkUvyI/h941zI0oGWej2glqj
xTuAx0kW0K9SrZjCDdIjCJlFTbu2kkBimgqhs46X99DFldBk7oZNMqMr3PkhZE7NTjHCa2lNKBZX
2S7yyMcD9BZLLNcsiQjJkNXSnI7KhgyuAH4cInrbodltSU361aVLBlg53cm3+bmhtJ5TpjHiqFbM
tVCTFqBeo3eoWZsCvPqOvAtBm0r1nw7+zVSRmzsBUFB0duY3IKmiCR4Xyza6V2dphIPJwhb41twV
maOM34r/b3dehrCXKCgkX98d0SaS5PVGvJYP+KTrPpUCLwMlVAMzE7PT8FgT6k1Wvzr9jDwlG5ng
wHXu8jZx57hFhcGQdnv4zIM6pv33fJadUpgTB/LfCtPJAeQ8TYol0ZMOWybQ+0VZ+IXyCpJOdg/6
MamwFj2GcA0USpe84oaUp2sKn4ClNGULatDiOldsyHBaQS9pxFuQHFX/btaYrJVbHW7nMQma6iJr
M4bg/x7xaV2WHEZgzFr0/5xvgiQamXhz8fK0x8dPftzez+RUCVuh9q8c+P04s5fqaVkUEeia3NvK
/kzTj7P+F7NrFL71cthbnfyay5IqiJNYa973FV2r6xVNQdQRUCM2XY9Z1xZgPtcV4v9pItPh/3f6
ZZLZg8EBi5/H+y44e0A1jJ0dk+FGxk4KiiD+RB/7OoOq/1rXEGhheGTgStK4F89x5KfxoM8ALzyV
0yeDZ22U6/FC0wbgEkcb9wdorCThD/0qM0YQi8/l7g6znxAlR0cl3nksp2l/KRr1PeiKnzU0TQrq
u3yL8FUp5m5BGwlG0TtcsE5OWRTmcMwC1AGFDCk88peEu1s79W3UbCCyaX143TEWCrYj9Sb7LNqu
Ke2DN4RmkvVhbdzgdxOsfw31+sxcV5GwjOvb9Ebbugw7NoDL0kuENkgeA+r+JilsDX91z74QtB2A
gwzXUrm3pwtibGzK/TwgbCLXAx1q86qr82rRoCamVG4uElc+w1zy4XzqNJ/sIcTYxIw+K+tjOaGC
PEOy50T7XngO++lIVdMrygxMQgmwQ+oOaeZXscXPvnHDZ3VLlFXViCh5KM2ZcfLZ0EUGgSzyNz6A
iGiCPDJF4v0YMpGc5gqpg/3RNGmQ8rwnDNu85To9i1T7jzpgVyRksiZJLclYbN4S8F/H2V8F8VFa
EZBRX5egow+7tUgkhFfseazZ7vmlFp3ua+wSXLyh/iMh7qMKEQtoyw+PX2FzXqS8kc50+CE49qnS
QDWnwuaC4R781SpwHqm5RvafCUmOKj9fSu4UYn9UMBkp/MZKGF5tX6/+1Jf7XR/B5QQ3wJN8WV9W
1QWtBoBmx03p6DaszRWafG71Xoumuf/qqXD3kSgisoBFB7dnfD8F/ks38EqGvRbzPOuar6HabzBT
g4wj7oayUOBBhIRjm7OCDPC2jwtyf4Ok7l4X9XBP2kr+hLzu1mgp5W1QYZYnUYjdOf1AiE+EV40j
Gnyxbh9php7zT38v28lRG+rPdxTgIniY8Hh6X6zSBKA8lKYByGKd575aZwMKR1na4Mfo+CABUnqr
40QgTlWKkfEDO8OphAM6Qv04p6DGJ8z+BxT3rPkSeWvPseD5WbOHeo5au/Rxm60f/3squnnOIVlN
2CnWUEmVMHkE8XFE7U0vKg4dfX8kq0yK9vDFv5hw36dhyY6PhQG2CLU2/x6+W07m+VTBTne1A4ac
vu+wDLEZHcjMeGAu1Jt0rO06PlLnGGEsV/SGIQrrydjC4jNnaczmKJ2yzHPwyrGuoOT45mOL6XQE
LH+RRPS6Col7zQogmnW5aqgRnPHx70GIoNfciDVliaNMS8eu5Bs/Qhq41s0y1TCk838j27CkuPL9
8RJLqNYlNkUA4bpFV4zwT9E5hF1/JI5V4H3QGU9bmjL47KgeRGOuaofXCYFALy1F2J0RqxGdBRfL
55QbVjMvbIQ1AdyUOsu6wXml4eVFq4fXVSM25FBWF8nyD1IqCqtfsvfiQfSxvrkl2uqppkVZK+Ru
z/pn5+yJH1jQ8D8P9aGtRnY4yc9TjBM2tBW8gFTa3uxTGl8ODm++hWuRY624kw/DQ3/GlQgZx49U
AZBYoAyY/L18n/BPs38OrCdsIj1nlX3Tzia/Y46b4AMoLZR5nhjrL25hRVNLSuGzg/NIf9MItzLY
xP1WdQ+j4hoCBo2uLfakFSBhhjWi6hJ59eheCei/OYg3Wdjq+gtf72YWz9U2UhTyXdobMhd3w0+I
GUyt+crCnnMQERpTKlfvRItiVSxtNkU7YYpnDYgkmqp5lHUy7Blss6RjG6I1UWJWKO+Ez5PvOry/
rc96aRJvagwjnunHQr724gk9nsCVzcwrU35J0ErX/kWmcuBh8pm9UchqJ1l7GhSGwSjuJ6l+ERVN
mEIUW70gdaeq3Fid8CVjxBFk1ca1Id/dI3ufDh/LkO86xy6bw8/l2+H56R/8ciDrjKCBB+WFwtYa
whWFcULTJP0RMhSmqFoIRy+cC7WbbTezWVD0guf2QxKpvkqQGLgVOeuAFVm5EEIDYvL+K7gySN5O
leAXaUVDKsPruQMUuphJsve11FNUKYY+Py79VeJQrusjZWoqtLxLtquxe4q8mrkBOYwqlTjkHvIK
CgkF709wnxtGXqPmLfdPk6lF72ufZ9ka0oq0Lb7VuEX4jKaQqIicZrdifH3ILCajQbmCcyyp+rxr
3DYaYLgesNpP++fLlsImE4Ta2yUILyDkBRfKWr6rIKISswZzDEsFlj07pqFzuCqmZawGqEAuCyWN
j4DSwws/Q6i8PbqBYWODBBJyERY0BwGJnNpQXwEiwQDdJZAC6khcsu6EZoGB0Cp2dwHTIfd7pG6m
NwXcZUgf0SHPinPUArnAXBigrIbyMWi/dnccBACeo4/zimQaQ+5lEW4WEKHYCOcqOIr6VY/DufCZ
VqyAtD4dYl4wQhKBXgjONSNr9ohUWwOHyCZInrzrxKGIW2hvABix6n/Y4V0A9a70EhJhHs4oIlwE
9CF6Aa2Qd1i9BgBm8+QlcsE9yJ5Hu71h7aLipWceQMqB/BXD3A8tQo4vZ/dwXR4qbvN/XxCJkCXW
2sY1zasP6US9ZulRiOdRS3WS/z9orqeWw+Haa1LSDvd7dTTlA5WGckhflFubCe8/nryMhrYO+RTK
1MO60pWFKcQsMi1RvE+XTjkDPWwKkpVx5PHSKYRU5gDn7mjd/8AOvK8O3n/WKp21aaYN9heSGUm7
sUVe8q/bFfueHvADkaJ8awPNjk+4ymQvY/8M/k3g6u1EGMYFhOyew4He/acvwJwYt4sFALvabWB5
vULjUly8xYgg+f0k/CJHtMHwolpEEWoqKZ00jzGlzMt0Egjt+VGjuPqNx4WKOJ8/rCnO7QhfT9xH
BVNHL5iyFwOeT3bP81/iE+XkwFOJbMSbGiirIOCT8IW/lQDs9A2hLfXSiByTI8Pf1tW5FkZFCO9R
HdSfyIa3sxPniULcBirr8kE5a8B5Bp2lC4DO1GrzrKASzVOKr0BM1ez+4xOzOt++U7S7axbcEhxi
xAFTaYFKvyMIASEinEWri9z9HSfQym/EjI//O1qXHMBF5toK0sBNbx3XDYY3sz/CUx6wG3uJBnhs
xLwJYzCKdgParabqEtOUgfpaAG9qqj3UoNjqoA4aePEvTlvdtLlKooOQcqboRjRXIJG0ZD9jnYrW
LkPdrr9EEaiBe9x/5VRiC0OJphknzwki9iV9A3SFSDPo2sAHNC+pq0WxtEF+w650IiGrO8leP5ZS
7DRkb+4IZIPJLoB+oILJ+RTGNrB8tsoEJurS7b5ikkTTGsMDP01AG0cXFmCPI1Q1pt+l4JxDSnR2
iz2rpjW+unhEBkAePR0lgSW2gUt5t+YbAyGT6Prc/FqaECNSuxVnyrlB7UCQQh2osTd5dbeyYbIW
/OTO78jC6aiQlooS3FBj1YTNtZfoauPxRPY0KwebAnmQ9PdECXzLQh8xLAddCfqDFoDYBzDRoEbp
WGDbYt9iv1k1TnGQ1Nk4mSVPHcZnfXr2OM969Kr0pYsSILZNwF9w238jdl14CL9RQiFLfw6yN6f+
ZAD8Sovy5EwlVx/tOzqlLJAPlpAqjxUwEGUo2aLkIHGNWneUue5aW6Lb8X0+eClzOZSWeO+b7+vn
tjH3/sO8ZfbfaP1Ybdvz+8TOvw9old+Y92oISzx/fpPOvG6DzTcv2w9dZCc3hBoWA8VeyMXg4Z7u
Dl6jFN/oWIh5KR/HY6q5U/DCJxibLaHSMS2PkiBzelSiGIvEXoEbcPahT+rdY1ZpsOr5PtYDXDvj
MeXeReK9ImfkB2naS+wDwreSSg1DA893+rUNeyyy0E6Hfe9Y3GeeK7iNq5XXzOkHKQqItpo5TTE0
KBRCNmUI9Ik1p6dcBKsp1Kp0Gc2ZxFuNI8exz57aAS6zYBvEZu6xtyL+/CWxts2KAkHGLN5rgoRU
ylAMF0TitYuhwizDxLAjjzZ0YoLcN30HjYkr4Plc8eWYR5PZunVq6FSRfMDzgA66AhGlj7k8Gx+n
EdhVQyrmr8AYpP2NG2smdrkR3VgklwEo6j8GKxmIucND9qBIM7VptK1+n8RHi5F2EKhTwgrysRof
amZioEJw0lrj+Jh+vheniK50ilRXREr01nuu6vvR7ZYFZe9J5QhtGDMsOUOiIz47rvxH4DXPGmI/
ZTdMR+cjpzXlcTEB3jUMJE2rJ9TAmSXqFsGbvzvf6hDsS3p5x0agUKkIwtoB9pgZMHA0WxCPv6EQ
EpBNqwvLldPDNOJeZ3kg4F3RE9dQBuLw6CieyXMjn7v/p0NF1J9H4KAg2Pw+OtRP/b769iVgU4bP
Ty9fgCjcOA3yFoTyJ88edpzvQOwjMtWeTfj+cSLvWA0gyhu/PYwRuOVx8OUTo8xg4VFW+ovLTScm
FOqi7mcKVjiWUjWAEH5xs8KsCt7YXe2p6HDGR499VvhavAUa4Sf/njGWi1tiK4KY607+na/Iyw==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity SDRAM_controller_top_SIP is
port(
  O_sdram_clk :  out std_logic;
  O_sdram_cke :  out std_logic;
  O_sdram_cs_n :  out std_logic;
  O_sdram_cas_n :  out std_logic;
  O_sdram_ras_n :  out std_logic;
  O_sdram_wen_n :  out std_logic;
  O_sdram_dqm :  out std_logic_vector(3 downto 0);
  O_sdram_addr :  out std_logic_vector(10 downto 0);
  O_sdram_ba :  out std_logic_vector(1 downto 0);
  IO_sdram_dq :  inout std_logic_vector(31 downto 0);
  I_sdrc_rst_n :  in std_logic;
  I_sdrc_clk :  in std_logic;
  I_sdram_clk :  in std_logic;
  I_sdrc_selfrefresh :  in std_logic;
  I_sdrc_power_down :  in std_logic;
  I_sdrc_wr_n :  in std_logic;
  I_sdrc_rd_n :  in std_logic;
  I_sdrc_addr :  in std_logic_vector(20 downto 0);
  I_sdrc_data_len :  in std_logic_vector(7 downto 0);
  I_sdrc_dqm :  in std_logic_vector(3 downto 0);
  I_sdrc_data :  in std_logic_vector(31 downto 0);
  O_sdrc_data :  out std_logic_vector(31 downto 0);
  O_sdrc_init_done :  out std_logic;
  O_sdrc_busy_n :  out std_logic;
  O_sdrc_rd_valid :  out std_logic;
  O_sdrc_wrd_ack :  out std_logic);
end SDRAM_controller_top_SIP;
architecture beh of SDRAM_controller_top_SIP is
  signal VCC_0 : std_logic ;
  signal IO_sdram_dq_0 : std_logic ;
  signal IO_sdram_dq_in : std_logic_vector(31 downto 0);
  signal Ctrl_fsm_data : std_logic_vector(31 downto 0);
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
  signal NN_2 : std_logic;
  signal NN_3 : std_logic;
  signal NN_4 : std_logic;
component \~top.SDRAM_controller_top_SIP\
port(
  I_sdrc_clk: in std_logic;
  I_sdrc_selfrefresh: in std_logic;
  GND_0: in std_logic;
  I_sdrc_power_down: in std_logic;
  I_sdrc_rst_n: in std_logic;
  I_sdrc_wr_n: in std_logic;
  I_sdrc_rd_n: in std_logic;
  VCC_0: in std_logic;
  I_sdrc_data_len : in std_logic_vector(7 downto 0);
  I_sdrc_addr : in std_logic_vector(20 downto 0);
  I_sdrc_data : in std_logic_vector(31 downto 0);
  I_sdrc_dqm : in std_logic_vector(3 downto 0);
  IO_sdram_dq_in : in std_logic_vector(31 downto 0);
  O_sdram_wen_n: out std_logic;
  O_sdram_cke: out std_logic;
  O_sdram_cas_n: out std_logic;
  O_sdram_ras_n: out std_logic;
  IO_sdram_dq_0: out std_logic;
  O_sdrc_rd_valid: out std_logic;
  O_sdrc_init_done: out std_logic;
  O_sdrc_busy_n: out std_logic;
  O_sdrc_wrd_ack: out std_logic;
  O_sdram_addr : out std_logic_vector(10 downto 0);
  O_sdram_ba : out std_logic_vector(1 downto 0);
  O_sdram_dqm : out std_logic_vector(3 downto 0);
  O_sdrc_data : out std_logic_vector(31 downto 0);
  Ctrl_fsm_data : out std_logic_vector(31 downto 0));
end component;
begin
IO_sdram_dq_0_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(0),
  IO => IO_sdram_dq(0),
  I => Ctrl_fsm_data(0),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_1_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(1),
  IO => IO_sdram_dq(1),
  I => Ctrl_fsm_data(1),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_2_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(2),
  IO => IO_sdram_dq(2),
  I => Ctrl_fsm_data(2),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_3_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(3),
  IO => IO_sdram_dq(3),
  I => Ctrl_fsm_data(3),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_4_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(4),
  IO => IO_sdram_dq(4),
  I => Ctrl_fsm_data(4),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_5_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(5),
  IO => IO_sdram_dq(5),
  I => Ctrl_fsm_data(5),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_6_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(6),
  IO => IO_sdram_dq(6),
  I => Ctrl_fsm_data(6),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_7_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(7),
  IO => IO_sdram_dq(7),
  I => Ctrl_fsm_data(7),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_8_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(8),
  IO => IO_sdram_dq(8),
  I => Ctrl_fsm_data(8),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_9_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(9),
  IO => IO_sdram_dq(9),
  I => Ctrl_fsm_data(9),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_10_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(10),
  IO => IO_sdram_dq(10),
  I => Ctrl_fsm_data(10),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_11_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(11),
  IO => IO_sdram_dq(11),
  I => Ctrl_fsm_data(11),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_12_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(12),
  IO => IO_sdram_dq(12),
  I => Ctrl_fsm_data(12),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_13_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(13),
  IO => IO_sdram_dq(13),
  I => Ctrl_fsm_data(13),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_14_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(14),
  IO => IO_sdram_dq(14),
  I => Ctrl_fsm_data(14),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_15_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(15),
  IO => IO_sdram_dq(15),
  I => Ctrl_fsm_data(15),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_16_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(16),
  IO => IO_sdram_dq(16),
  I => Ctrl_fsm_data(16),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_17_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(17),
  IO => IO_sdram_dq(17),
  I => Ctrl_fsm_data(17),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_18_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(18),
  IO => IO_sdram_dq(18),
  I => Ctrl_fsm_data(18),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_19_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(19),
  IO => IO_sdram_dq(19),
  I => Ctrl_fsm_data(19),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_20_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(20),
  IO => IO_sdram_dq(20),
  I => Ctrl_fsm_data(20),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_21_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(21),
  IO => IO_sdram_dq(21),
  I => Ctrl_fsm_data(21),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_22_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(22),
  IO => IO_sdram_dq(22),
  I => Ctrl_fsm_data(22),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_23_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(23),
  IO => IO_sdram_dq(23),
  I => Ctrl_fsm_data(23),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_24_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(24),
  IO => IO_sdram_dq(24),
  I => Ctrl_fsm_data(24),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_25_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(25),
  IO => IO_sdram_dq(25),
  I => Ctrl_fsm_data(25),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_26_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(26),
  IO => IO_sdram_dq(26),
  I => Ctrl_fsm_data(26),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_27_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(27),
  IO => IO_sdram_dq(27),
  I => Ctrl_fsm_data(27),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_28_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(28),
  IO => IO_sdram_dq(28),
  I => Ctrl_fsm_data(28),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_29_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(29),
  IO => IO_sdram_dq(29),
  I => Ctrl_fsm_data(29),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_30_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(30),
  IO => IO_sdram_dq(30),
  I => Ctrl_fsm_data(30),
  OEN => IO_sdram_dq_0);
IO_sdram_dq_31_iobuf: IOBUF
port map (
  O => IO_sdram_dq_in(31),
  IO => IO_sdram_dq(31),
  I => Ctrl_fsm_data(31),
  OEN => IO_sdram_dq_0);
GND_s2: GND
port map (
  G => NN);
VCC_s2: VCC
port map (
  V => VCC_0);
GSR_3: GSR
port map (
  GSRI => VCC_0);
sdrc_top_inst: \~top.SDRAM_controller_top_SIP\
port map(
  I_sdrc_clk => I_sdrc_clk,
  I_sdrc_selfrefresh => I_sdrc_selfrefresh,
  GND_0 => NN,
  I_sdrc_power_down => I_sdrc_power_down,
  I_sdrc_rst_n => I_sdrc_rst_n,
  I_sdrc_wr_n => I_sdrc_wr_n,
  I_sdrc_rd_n => I_sdrc_rd_n,
  VCC_0 => VCC_0,
  I_sdrc_data_len(7 downto 0) => I_sdrc_data_len(7 downto 0),
  I_sdrc_addr(20 downto 0) => I_sdrc_addr(20 downto 0),
  I_sdrc_data(31 downto 0) => I_sdrc_data(31 downto 0),
  I_sdrc_dqm(3 downto 0) => I_sdrc_dqm(3 downto 0),
  IO_sdram_dq_in(31 downto 0) => IO_sdram_dq_in(31 downto 0),
  O_sdram_wen_n => O_sdram_wen_n,
  O_sdram_cke => O_sdram_cke,
  O_sdram_cas_n => O_sdram_cas_n,
  O_sdram_ras_n => O_sdram_ras_n,
  IO_sdram_dq_0 => IO_sdram_dq_0,
  O_sdrc_rd_valid => O_sdrc_rd_valid,
  O_sdrc_init_done => NN_4,
  O_sdrc_busy_n => O_sdrc_busy_n,
  O_sdrc_wrd_ack => O_sdrc_wrd_ack,
  O_sdram_addr(10 downto 0) => O_sdram_addr(10 downto 0),
  O_sdram_ba(1 downto 0) => O_sdram_ba(1 downto 0),
  O_sdram_dqm(3) => NN_3,
  O_sdram_dqm(2) => NN_2,
  O_sdram_dqm(1) => NN_1,
  O_sdram_dqm(0) => NN_0,
  O_sdrc_data(31 downto 0) => O_sdrc_data(31 downto 0),
  Ctrl_fsm_data(31 downto 0) => Ctrl_fsm_data(31 downto 0));
  O_sdram_clk <= I_sdram_clk;
  O_sdram_cs_n <= NN;
  O_sdram_dqm(0) <= NN_0;
  O_sdram_dqm(1) <= NN_1;
  O_sdram_dqm(2) <= NN_2;
  O_sdram_dqm(3) <= NN_3;
  O_sdrc_init_done <= NN_4;
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Wed Feb 14 11:06:46 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPMULT/data/FP_Mult.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FPMULT/data/FP_Mult_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
JhbjCPusrmUQ2YbR3+HbXrKQkeZE1qJD8Sg/+jNG3CIYlCxvta/Vkv5cWrC9Dj/3sfy1mfdEIVp+
xKuhK9PVJaJz5mPR9ROXk5VNXg3Etid2gNhPvpe6zSHqkwUtdLF6RTZPyva3ivENluXrJRxhG85k
I7MwA1sXSCLv5lqRJfJbWeITfDtvGBUtnMwgkPoe0k5y6m9IXITk5jnAf7o1FZpFax6f5H9GPoNH
g+QiiAxgJiXQ23tU9KBjTFI0Fx7hzGItpKy7FVo+rRIDnf0YW5SVRhI73zaRmP5/+AZLaeeCyc8x
k0petEoCDsQ2igGjto3bVA7pPuYwYrcC5BUCwA==

`protect encoding=(enctype="base64", line_length=76, bytes=220640)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
TlKc6uvaL/iz88ulY/qxRJDzswAAkQlg8cyshEJVhjQdhPOoB7WeK8MAZA2riu+Atl2VGEqTpK1F
FNi3w4C6pxx8lfRKw/5xLzG0eBZMRX3y0mm1OkrOOHlxWJRQsuNKrXm1SVFql+c9FZoYAbhCw5Z7
Oh7KJcuioCKRhfQL0CwufOIGpDZWYqEpTdmOmJJZb+FDpfSGt3cJsoNI1KR3ALzF7otyH3gv1Hk9
436qEVkVSJYDlpCFnJ5Td8vQQXbe8xRQA7TOWrH3zmXrUPFZTpyjlYHKPkUfce3HvlAEwmDxekrK
Sn+UlBKegSNK5y8obXUPkdSdT4MZhH1HyqgmTz+WLlVgdSwTICMiWearGPBGkp+ARhde/ZmPqWg6
TiCF/ItdXrC+61Lcv1gJScgLxjP+ZnYblsNe8izDcuTy0AxJ2NIXCLOJhbNqmvUGpncl1bOB1LRq
n1PODOzFQgPsfOnWTJCDjPGe2d3c4jxUDapRFNUf22Jn8dwGQpiY/stRKRW+pYMaUMR2O1JTH2ZZ
taXsGm6ldGRBnA8xsTjNAjCmrd0c5Bjyaov6/tPPOM8AqHuhlXWe/IH90D9Q92rEyjFDu68vLxxY
AvpwcwO4gF6pQqftH055UKRi8/CVEFZ9IG28VEwZ9US/7EGriCyeTEJnx4vUlp7nN+frEutk7dgS
aIONoa81dma26KU/eFWrshEbx8uySxPzc6dgnLhCVX4YZfUqagPyLOUMM7ZoMwp4M1Uo+QeuqHpE
akrXdsG6jSlZSyq3Oj29uHhcAamipbEt2VHW2suwjhkh4gi4hmYed+d1gcbW26237/i8VdKQJoK1
U+FoS9Yc6qDzvT3LLqwHQka+eKe8MlbUaOBGPMK2MqG63QS8pA3JS4wkGgwgIn0UFNwqtHZhkivr
OnYM/MVLydwGRuOiXKCI2GHWri+OMBhaokFUY1S8RowBVabNoG4bHdRvzcIK6PJfs6kJ8cVMu6xJ
QMrK5pLxU44xsttXoshXJKUoOEVlJHzZUwFjXE/cebu3hVHUYQ3uljOYYXM4XNhEwlwKxBG8Cjjc
4A8EbnVP+JrjgmAgaj46BiLYNg3haWOSfW23n8QZzfUWkO0XPEoFrbUCTHv1NxQiMJtSXfAAXL5t
z6g0nyi+vzrncRfYM20LTAEB/bXY+9hkOTuVlEht9ANLgBbLWzTnFv11AWdwyWMLjnFrRSa2Ze6G
OjaKQFxOBZwJx48Ge7uytxcoEa2tKVFcmuYHO5QAL0jfgvknFqoU7SC2BAl8nyQRcROY0DIY3Cav
f8NnMI5G9rXPBQi3kbbcgR4IgiBpo2bhOm3nKwP2qgif3wqHGYQwm/cLbHxMLcj5wUeiaysxXBIs
HRtiPslzBNhLHySFzQj2rb3y7q3hWCSthhg5mr6EZZWXH75pF0TEZvXWKobafGdIWKpp2GjDod5V
1ANtx0fuNDd/ZYErNym7WVFBm0htOXNSe+VlWsIy/BlpmSjXO+SNU+PBtY75KznUHZWfuJYkrNkh
UypL8s6NA0OFbeDpUf9G0kQzQKSFIkB84X1HXecT9Eg0rJE7oVUr/f8zjxrc0aL3xPhXK/nlz6SG
Vh5KRWXl0tprm7p/qeIVaeYHx1i7I/aoaH0V8Uyt8VF8Pk5yk4QiF6tI6vLJ+uIeLGhMMrGnMLbL
VaT/6vNaYdGeSPIs32bjvYchQx6oyKAmwOxls/xTyx2zd9bV2Z0ikyMX+RAbVFAtPZo9og+X0xnO
xaw+YwMGBYceIm9hFR3xTeZaF7dTjyf6FjpRBzGQVRENp2Z6tit75ca5xB0AxLqR8bIXeR7LfhU8
SblPoCKM5iDLPKm7Xz3MtAXU7d582/vI8XcgBsLMPpDcjcjbFZtwedHI/vo1t7m7Pc/9Of62aCE6
kyLROcEfL0Uxm0NCuDr8bH/fzqVNj2pL7vbk1IfMABr8nxwmaKT+4MUrrK5ilgVi8PEDrC8R8w7r
OJhWfyDDoSQvzsZ0A8a8/GhllwHEo00R/eBGH45oBWTNJjBHIL+mG/Oztv4bZplMBgW1V4mzb4Js
kPeIXdsPPcbDToFS8Pr7OYjRYZ5SGn6/l0fRmIVNXjSvtE7BWc6PH0WGyXOajy/imVZ+FN/D/W6T
JPHVCWKD6tdZZ0urmcz2s6UtZC1ps2Q2kEoxHFeLif1TEwL55Xnd78V1W9ge9AbXJqlWQ1phq+fE
FFBL9Y3L454sQEM9JnOXHXgn4X+XSR1XY0gosHIXYioBoF7eFMArHDqSBiRqKPryUIbjywy+oUna
HKCEYPXZH8cwtiBVuHsvqa8dVq4HMBNBxrMvY89qcZbScF56aidS8ryD+52dIl129PEVPujPr8To
KrNQoW/yno4T0eNE8TsvcRtPLOFhtRlkSyISHLUWIN8QcFh78jysPiq1lO+//qYQgW+sc5sPKiBc
rXWC2bzo08RxYialDXZ8GLj+zhBEUsswGplVv/zgc18ePT5kuJcw7mjwIMrMnyg675BmYcsegXlp
IuAbNCma3xzvehwXMP0xNK5qfN5EFEQYX0YmVt048Xjlu7IeTp+8ppobvM9YLZbqaJZsRJJWjrHv
M+0oscCeCDCvUBJXM89MkgJ6/AJNyCy778aRvUgCTfwb40p90KvaWZ9V3/O8y1T6GvQLZozC+VV9
8r90Bg4I4vzlD0FaywyxUqtjyMpHGt0bpQhVNNkInyjHUM2/PbsOUWg0JzspUq2Yff06Jxw1UXpv
upSNRpyGqIfqwBRY1D538f5Rx9B/IJVby25iWQkU2adDeIH5ZUC/3+NGh/2wjQaYJwPG4DzVcK7x
WOGAVKcYVzUAQ5z/WuuFrjSJBjz6Nnq5dpttp60QBQ01AwZIN33p3NPE95TbvQpHZt4Ow6YX8XZA
ehpOJd8sU8IGiXfYYoRuqXT0WMqPOniy6x1/8pTiThuVDon784SuunJ6nDbAmucZNNxwk+U9PZQR
RKcQfD7WPUuysJAJBVhzyz3jnxwo0NGiLn5F8BscqhE6/NkC6YyL5temcy0wSWdF6VnL1oysQqxp
gOj5WwOWFanBY1jnmYZkRowm182jM7IATcpfE6LR00Jmx1L+t+XHS8OsJdVTGE7PKIa/AGpP3oLG
bksQtfkLht8GSLEw1O6/ZhND9wSUZSKNlr5jSWe2wGmVFzDB4+rkA/xc8ymJnq0Yza1LR1btv11c
b72BRhl8zqOa66XjS55dQK7vtgSuGBeK8HKNJ27zO7g/E98wUlFTqtdLerhxDLNmSdfQRaAFmtO8
it2/dhsvWDMiYPhcZKllQhapgFqAlfn4w/fVtBWSd4LZlGfpfTld/l4zMzjAaXuKRLUpwBI34dZ+
3QnTd93cLbTVjfM/Q20XbIplJ043EhSoUILm2M4oNkIl8xPGNbgZrNVnr1Mt8BH+Ot4Q3ePUJASv
TxPt+Kx2awA85u92Ryk/zCENFRBZdwrlt+SANrf6TbqtIlfQyR1J3G56W0lNBd+0fI4wKfqiutag
c90RA3fOPRC3zHb0nySBCZf7m9VD5gPeKgjM2zSH6CaP9jDpBY25ooSOblFjS/9VDMgtFeVwDqlz
YNI37yVdwx+JTopQYsNRv1v1FlBRjiOQQt4qoCfNi1wIaHDnI2SxFGNF4W0nR1LrAZV92iEzWLYE
E0ZwOt0E1tsiV4clPYd7pFy6b9BGxIw1gWxDOCfI494h5LACH27lqJ5slnD3y3uCTOF7TtNhARFl
RMjGt2u5H1GJ2l+CvasiCOuejj52y0PMrObRB5Mdi7tBK72lXOp2ulSF4RYjAaTwXeW2EEvKJNxe
hoAiHRoCLjIEYYwIfWDZ9R3VaDgeaEVZZr5yeyCDycmWnGpZEYhlQNsnP1UsqHXnkplzPvPjUn9v
tNLa0U4rz4k+QOJ+btUq1KvSenaK4hBN4lQ18+AqECqv/IBEcKDx2Wcjh4UWptk98ytn/7AmDlWe
mgaAoxDJ1W8UDUM8kh5b1fC3m5WMKNoQubsuhGYjVEM5FuvSkmAiejNMmPrZemQjnQen9oVj2ZVs
/3J6rRHWcJMv/Izm62tNMeSLYuCP07KHiePx8HiELucV625PCutx+1Z7vMeJGwoQXvKa4HCEUURm
9LApCnuy+Dk6PS8xOgZnt5hSJeshcYZWvz/LFL7Tu4T5l9FfPWRkJv4nUAPAglK1XsQtMqALKnuN
+BrLYr042AZbK1v2wbFxR+bpI+Px/HNOBYUa8YNdrPbBjrrAGIP0ejhPlQjDR2u0tYF8JvZjOT+7
lw4d6KhH/w/n7xW18mdoWC0+NE25KW4yPQj7T2hKFzMcCHJY6WFxpSWvNl6ZHqZ2rxBg+vf2h3CC
cr5s6otQnAwPPsF10inG6YtITYhnw6jQaoZ1RFMbyzc6HBeMcO3uNwPAk34MaFM7Nl7LoKeKuh//
00HLJHOai8c1IeuySgPdtqbIKbtH63njNoifHX+dowzbRveLVCdF8ha7C4DwdEdTSv4KHgE8UbqL
1cIfzpIgk43rW0s6Fkch0GhmWvIKGE9rSD3xFWwwn/YPbFZHfmwM4br19OPlW/MLIJg/oS+q/03j
X6ZvCPrDnAJU5/R/rKBFJ2h9x0fYhcrVCHzrz1J0UJcU4vPKoRHyfTYLIgg0Bj1D2eXzRd3FInOF
W2bMPiGi8tNBbUJakCC4STOOzCTiXVfg9v5R0bwqMBSMkm1OyFacCFSlBcsnNoElCcLycNHvpLcW
zZnLMDgKJLS81yW7OPPXpsPVw4se3rfKUfpvHLETLP5xKvQ0PTIGsdu+bBBW/R/TW1IJj65vGTl2
WbXH6M4uzcTaNaGipw0bu4q4dpzOQ57a0CVkx3Q+wYZbA8IJw9tTvHSzxMQrIEc4cIdZs/oVY+MI
KXgKBNTgd7RZ7QEccsfD1Mk+M00drwwSb3TzuuZ6dHloZSFL6fR9M6I5OmeEufHV3cK07U78xKrk
dUGoOHAaey4Ah4EOWpZtvr/OBMveey0507S+UA2gAqyjjM9d95IndQc6wU6RZQjBSu990swj1ra5
0gcvK9iJuw7opGDMx7plSAOoRaCjC2i/yEtlc3lQlUYj+76zqb6gcaV226Q+DBsBM7vSVKxZA1rd
JCoaJcaIhlQnM3qrXRW6ZNhg5CWI9IKXsTAMZaUIo/y6aQi2toD/z3gYceJvwRjpX1GQ68IqsKA+
4c6f8BcjaW2hpPKOg/WjYtK9IIRfqEbN7dI9biEnQDXXjIp4gbvLA7q4LVB9i/IeyD2bMRhSqenc
jPTCw04THEHiV/Tyu9O4gqraSMQ92sJYJY48Hvj+nHcCWv6eqNFAXeVj81qngmB91tCLJyi0jUwM
n9NegBlL+ChUafnQYs0P9Nu83+zreNPi7nvo4gmEzcdO/N37J/cBZkopYA8U8Kgg377F7qAhgr4Q
/zD4eBxOv84F1wj8in/a86Y8k8mt03N90uBWvkcHdZd2mkKhRTCHNzKFQnDgi7z4LPYkRtxyKRxJ
irh1osRPJPFPwppvYMVBa6IOD4N1SsF5RL+NE2O+TOm3yrALwCScUhOsgLgW592twFeEl2A91VI0
DrUQkO+EZFRSWecJDWiZMlFgWw5aOd7EvK8O5Eco1KkIvlNrojPwxY7+hNeTJ8udrKg4UhhQTWex
xnlmGwXoUNyaIZJ9n0lxn1sg90w617KaqvQVrH2cj32rodggAKmWequUg0vLnZgItXMjTd4EvBuL
WcSYKnUQMQkzcYruhosjx6XcAQnJwFGjSt37bszfNGcnBuMPR4GogTjqcjlqLQn0bM6s3X463T0w
NTVxYtuETbKLv9QCoiu5cI60OneYTFomkoJ1ci7Wz/QX4oVgRQKMZZ0/88HEoF3nRU9BUYE225IM
k7pD859CdeMuQ0jxZpQNoGhxU+/A9Li5CaUok/EUUycLH/co0VE38ZNUqstDATUaYjf5ZdUNblCz
dJyy9Q0OJ0v26EphvP5fOHvAf6APGlakJ7ZSjdIrqp4eMr5DVKES74kUCS45LBk3OoeB5GHPDYxX
98kwow11ayzEpCbt19enQpzQSgFotsMUMQgAt0qCG+N/yqh3pzHf3p+aCbMIF3jdysLEkY62rLIY
TYawi7qjAZfYMAOvyMktx+9/YBt6l3Bf8Omq8It3k7ohfI8Y/GLNvvhELhiq3uVly15QZ4R14btK
yD8ywHGmlT4lB/Geui1lAuhK9kNY7Qf4REwkBSTwK2AUDV9fnbGB4y8VXjIoPlrO6G+zSeDzQGaT
QfyHoi8kOVvlsrpTumGxd9uKP+PVoOAEdllZPOeaJ8XOSFTfZT3cHDSITxxWiLr8H2VHcd1uB+sQ
f//JudAvY8QYU7bS33GInW+KQaOYJ+bZNv4Q6QXExj0JIWZJHVpG/VQt74KC2+uHyuoU6gJYs2sB
s/qJ0ro40q8gO4ZwwLyTb40DZTelxdV2+LzXCY8ZZDrWhk03Mbe9KtJmDE+YyWg7ks1x7s5HHb8y
1xDxXiU8qVVUvZLKe2izPNUjBTHH24MQDyAi5o4oAJ2FANcUcDrCatCucCQuN/iSXylDhTNarRhc
x3UGTCg4Ukgbj81UNveSDxQHJuzEw6EwHkwsivmLMP3ltfPxL7pevyuMZUJvniaa/qEVWrKKO1Hz
AP+IRW6zpLXoWSjY/LdiUz6OL6wkYqoINLHj5vQpkbChMqSnE/F0eQewgw28FH9Z1sQCZbaV2PeL
EU/juAy4469M3blbYvfn/MsvIT2xsjpx6ZYYRojCw+ndSI6akc/Zyesj2u9mYIPMGPSVMtkjb/Um
0arBBC/wB+ztWUOmoBnoPKJGIoKqehaJtD0NK7ILVLf4J8BTS5kc1jJgU+H1vaX7UA6PaE79MZ2g
uSboFRauXdRmTrweIJ1KGBLHIJgEySFRS4Jaa9MMTg0a/hCKZZ5uB7tcKtKQZpbpe/rM0CRBJQ4J
IV8l4ucqWi8admlpLaWzm7UApe3BhapwBTAoKXFRxs7T7DYi+wP32de++Yhg8YWqtvbUOIQDYrH7
0gzXoB2KsqcpoYL5eZowys+HO7w5tj77LGwNsp9Ppo3QBz1dHCkTmi/a3SMWMSn32wI/EVIR8iay
Ds7W6cBBYzzeuOmPcT7+AVw1EEZECGoxSBKFEeuWd4yvpLvrBY529tcq3gF3k0VXbuYC0GppeeC+
w04ifbQEqLPSfhvk6JGWyG3pC9ISGC9EAKD2A++Hv143BdFocqGLSAjKJtUYGqdlXtGmBAKh2jOB
xYYq95s4arLOLVA1kz8IatpUobMF6a/BYtgn9XNZ3657y33OhDK3ghoL6BTh9xn5g8N5FBIjEptY
5FfgRWxrB9XVi4vM7DfPvv+knMSQ+1YTxK4qevvyJWtAXAIg+cCIU/iZByufQ719y23/TdgHvM6j
V3rt9a/GzvYdjWIzuADAVMGHW9FEYxTPoOS3Ks99yFNqhxgcwr+rZdl1QZks1Ehrg5D69yF1YuTn
3uZ5cwxIUk+hNX3HsaO51hyvqUguAqv4tYlE25S+CEW5j9PUWtsOgFdpLoyjASwN/kba/lak5RGq
xP95PwwH8l2UQT0fUCbKPFSpiJpevb6Or4DvZGldkoYuuesDB0TwplDsYwUkZ2QrSHQaitc9jiaj
AheNVWbU3L9NrkDC5t7dDoh+9TLCNuB5A9TiPaDg9PMmu8N7Jxuuc+SEIOO5npvPaObB3CVZBt1U
5ovJYXirxbPx6MHllfNj69M32RnO2wppI6FeD2jKMB8j6XnrJNW5ejxTT4xFaS/jjNtO4Cslkk6N
YmmLtrdfJe4JM1zjHtX4EK8K9df62JUfoaEg244Wb0A8bYG0jHSEooL6ri2TbBTS6o0jiFs1acNO
gYJJA/4Yl+QNhZ5Bx8fF6ubks/YH3pkbTRaF3xxS+eGQPjUJwGsrda3gXwtg8xr3Mzn+MloeatF7
vSUGlgvZX9Xn3sFOxWZZWsPfzt1a42n94eUveA56oL//q/MdYL+7NnoGqZ875SBIL8tK7UKOQp8v
ELoNhqaf2KQRvxeknD+r6J753WIBW3rTKgYl1IcJaWFTjUykZxMfKKKadP3m38a3qSJKkcuG3Z/e
+k9MJviutwMqZasDcgLmvvZLn4IPejchjWkOw7IXHI/CvJvcNX2+f2O35J5VZDZxdrPMO9rn7hFR
Pih/DPKEwiU9UWgYHcBMmmY8oMDf1JyJUmSjPcaoV7WmYC5I81W9w+Ukae4bbNrC2a8WLaN91bb1
D8Y2TE/dAoFFBSDuTJd0WhrOL26qjkgCHs+o1QX78eFIzH6QNzOL6sjOt6qsIiZE2XimJ6gSBfHr
SnJxetu5MUlWPvgFrb9Z8NbkO2CeMmouPjUuUYuGWdJ7I3PD53sDjdIulppgRyPbbMmYw3qDlKP3
iuMGhciM4gvhC3LIpvZ5hFOllbbjmnmm9grhDtXdVnpa5Je3FD4nzIIsCb8N9di/QJHjLy16Onfx
Enj45NG5jXEOsJWYbQxtY1XkfnkJZbCFQly7v9KbvtldvxmQn2Wdl4R1tlUKO/zzYuR4hGtVfiYF
ADaBjkuFg1zb7zYfH/0mYNZRYhVeoJ3Ua0om74hIMtbXTSAAOQErPOVAYQH4ETG8sYhzlr9NEGnD
PzCCG/1GuUgYpui+WGOkU3UKS2DzN/lzS8C7a/gmoK1tUUpG8nOf1qltzFRaeCsaqCK5zdv3O3Gh
7pEAE4gu5evNQmDPCYaZIUz6KPJVSd6xnBYIKtufcpzpy95cmncQcfLJpR9ZRBy56xOilGsM467A
GxXp+p3Wtnw4da2Nd8ltS1+lzdsnDtGWCvb0XxdvXCjFi3vsUsB9UrHwqp334Eow9rNfloKv0kzh
4KIyLSapBlhOv75JbkikjwSECcust8f6phiD3UUVVsWfV9n7Zw2hJxUDYpFg4Os2C2mxtPgLnhIs
7OvEM8/bKNHVYrQXGM+ITNZXI79jh+ugVAYD7UnXV/qn+Rm+8jJ/Qy3tMJFNpsQRhpR82tSOauVT
KRIpe4vZ5mE7FyecWW+8rdixtPiEHbiL4z5QMXhBy3sw3SH4cS384GSK2KB2ERV9d1Z19ZFt48jk
+Wz6ezApiZWXNeXMcfIDVg3SexgCSzq+C2CIPst/rM23v+qdiUSpwvWK0aSkhQFjMvX4tethTDn+
+jgJANqec6wbUbPNqCz9yB+gGyvxs91eWki6Y4Sr8oQqun4R0qTyVkT/8h8TBFWWpXavqapfTZ41
lf9VRE3JDcWiQ+n1/hzc1sBf/TrN11SVXbX1DElgR+h1NcGdNeTHu6e/BQ/c5Fm8jWmDsLdMO5KC
3wF+UpuWhQ0PeTrgd3GaTXLWWQce985hVRMpMcBUxft1i2OZ7+++m2AS0K1aoSUdHBh6v15nStDT
BrnhOqmyFFnEwLb3WP2kXAmEWlpxxwtcixDsO78BiD1mTM+3grjKvNStTz5gCZmlMdutbYQ5bG+v
QWteWn5/+zsDT9yRT7yCjrxJSwVpBMxYzNiMGTbh5tm9kr7GvH3hOzV3SGrdg6JFp4CvB0+2L1I0
D72QneLYYOVzjUu5/DOYYkHr3X/0i37JsCKyiCpG67DeJEZRSpaqe+vxCaZfhBZFiXpPpRw798V9
Woeg5WT6Ch4YNnJcsgNUWJKt0iQ5gADio67K/DAgxrud4F7es3fJQfuMv0HlkU3XIUf5IKRusMk7
O7HzABOTzgzFLDS7TAP8c0u/PXSHyfTK0bGl1elR/rbo3oZhxDrmsnAsR9KoljlT/F/osvJu505/
ehDYmbzdZZuNHb4wse4E42snZ6I2q8BNaDUw8oEkAxAH5kr1FZTRsdYtfGp43EsLrz/uqpCYiMl9
c9J+0KxvedZRY410H2B3Gz85l+iasJni4iOW+wrt+4eZJ5bY8IeyLjyhGfwv4fqBxAAzjY1a5/jO
SNiGFc5y2TNjEcdL0hn2pWeACjqkI2Rm3+P+jWoCqvqTV+2gp6eHVq9cCU112pZljVuH6s0bVRef
0w/PYmhbCS23kiQxY6+TJkoaOE4eTWm/7ArIFyAlVORMwAgumV3PAvvhJTrgTo4oLZ+ic9gFwPFj
h9qcgNH5q+jE4MEWRCTdp2/ZjUylfdBqF5ErIMUSgbbJNf2EjCvnI7S+RYDYMqTIglK7t7CowrK3
pEbbWxU+aEZLqb+s87QS1w4uf+RDbl8YxgXamshOdU7c4P2kkIlNi6yAfj1PWAOBu/JQV51OgySK
nysNUxXJS2WWLuQtSVJfxC7Y2654jnedWuStBQq26zD3mOCqvbBKlYfOzWmjAgnUEw7ZiDfZjlts
J/kevgHVzX8GCgEnweuu579/Vinfwhqm0VwvZXOlVJuIDlx6J3LBrHjA1O0+IVQkd8f3N8MEG2cy
h1S7718Z/j8ZRnIo1JDqBT1qU02+4p9yzLkMKDRgSx3BKIZ33q5+lk4kBE0Y+biiUQ3O6okfsiUa
KSqm4SFasINgDC2bWZNfN25ppAJk53XTFfDBtM33/dQ0ptXwkogOCbngAwY3w7t69yOZrRBRBNuk
l5KxDF+mjfhp/CA2HOPsgl7yaMpzz1yit56HKj8TQ8cjLw1tw/RBZrcqvjXKE8c8yMAPhghz+Kzb
RtciJk4oqI9M4qf+9hryAeLnnN+ZiQ/DPEVNU/aOKTQB5ikpGzNnF7cWqvDT1+iU2kOzLfF9AWwy
iMJwrXjgSCwV0UVCy97dnMpUbP+GtIf0BxAwhLesY2UQBO532UvbWuvmISS4uUzBvHwe3CNdXjet
LBgGABHSxRNNyUaEZL1armWHQuu1oEr37a81ibnC/d2nr3GL6EAZ3vW9qEsKDLHk2J2mwgdUwo0u
Sb+OiUaao0okxPPO7JjsYXHE8l+X/VO9gRB59p670htq1biQZABBCcx+Zp+E61fuUeNR/He3Nzj2
cqqy9m1cHG9UDIs5w0dZSqJQRI3HOUg/6dxPlwwX7nesc/4SsHpmXJ7WcM+ECCshR55k1me+B0HT
bL2+UVQCs7MTKGagzXq/ArVpGa/GWaHsNAZqN3BAGEqO9kvvL563l2KffqfSq5Ub/YTE+9LiLqmV
Smk96Te25WO3p9dm1TrK2oMJPCXIQqQAvHYxFy7y6MyPOOCRyNTzQ3NVYrrHymUueCFjtGrSniYz
GFr6jX5cmneUSti8f+jwTi8V5D1n7+vZXAgGRK1BRMFng0KW4Fy/57qFoqpI1kSOtWhaC+BXcg7R
GI+nxoIyUGoEsgDIWV9tdZ4TcISR9rL9VLRvvShAErFoTWZ2ztLFZovLAXJyzakYn4etvR5oyC8J
zC1IsaLrkLPVLOSxegsxPByZsZULctBJW2UWueXTFd4r6nUN1woZyiwMi+xWnrbox60dYQ67o8Er
c3oWbMuFJGLGQQf5g9xlCXvOdx/N3VJ7GdE7pW1M66OrlZ1H0oMt6C6jU28PnPpBXCsv2VuLfmoq
CeT4lezA37iowFod2gURJGnT2NUmn4ulIO6UEHdAMVzbMUH0kA71JWLxVRZ/9oOscR3sSStfWAi1
Qtd8x8TRy5Q5KSZ83Gqt19nk72mh3SuE5pHXgn+eLx66aPuwcZrgxWA7+hVIaiixqpjOlsJonVKU
Okv010uxSQKyFqzmioIlg9qqqoFFtXdx5+OchjoCCyjK9AIu37xZ1uZ1ukrRsfdEDGqRn/1dOUZ+
RHV0Q5ssJfCrudiB86UGtL43ooUWG0CvghR6PLGODCqhLIXXPCEoZf2FnIkXRJg/2MF5/vksg5Op
or1mlIcDDo+YaNM8sWCqLT9lnqWe3PpfJtHci66jcSNsFSYlxIzLUHk+4bcZZBJ4mLaLum73/W8V
SP/wPotFK6QX51Z6VWjA/MdxyK6lWtER1MXyUsZR3+K7Q3BMM2hs9FUFFT5J+zUfsAJvE1DQSEtk
ki1MxxG42WGEtUSCZf6iJRCT21gX+BImPNo0EsxGcBYPjWf4XumMLGB4U7GkASvrKmPLhE9/s3OV
oamMy7EYezBgFg7g6AM1gxgOji1/2Rqal1DhUhVWm1wM569PlAFNk0pgySm36wOCyXkZ2sFNS4uS
1wdQ6CDfEuPdsvAg8kQ44gQFwMXZyABa8B7OAukfTfC9cn/Ad9anloBuMR4InSO6PMncxcp5IWcV
/zN10PFyIy4T4cBtrc6tcVtqGwI8ON1xnrKnrVj9PF4jEzXYMYcwyE9tZN8x2ZASbrCH6CeWeMRv
dTA5lTPqJY9AUwEaLioMfBwSY5CCBHHUP0iGYfQtXbQyWKqvll/iyclq+EaSZZmouxcpZK6Qq5yn
q2FJyy9xmYQrv/Wo/I10kBqR1J1TRM2qPKAW8y6bggO2/cWdTRadXwiCa6ri6wj18rHF2U/Q2Wwq
6OAbWx7zrldRjGSwkosKRksv7zr5j0hrOPwLp+1yRGQ+XXYl9JspdS1SWNSKd6MrqzuEkCEnwnmr
5XiZrXwrEcIh/4lT7J4dxT6hz1HtpV5OeH+Tw/nrRYmS5TibdY3iWaar4P9rh5DdALEoFBpWPwm5
/pmbz4L+VYDVYj0aNgSPe5ksO+42ocCo64dgfg5K1iH6Tz507pDGqPIwz2TXkfI8iLQexEAsPaTh
WbzqHNzt6P5xepk+YEhPDZ7sr4Xpdpb82Jzd3SznXOZ3DprDrT9tWa9Aa7iNsRThziIC38WVXl4Q
/HnXVN4qGJt6jmRkh7zddxO5jlVXqwZ91T7ia0/pxKKWOHNPlmssW7GIf7pE/8NDFTKPScJReEMj
/0GPOEIb3hK2Krb0m9w4GQepDOjQY0nY5vCyINHZVeApCuZZypm1gs+mTsEroDnToK2mTcSREmge
9Cml60Og65DIQSiwI5lMrb6q3eKrdcaJSyf2nIwt/FNZQ4TSjNim2vnspybulIzlafwi2hZPKuB6
QVnLf0zFUUHHeObXkBWdw6jo2RNCce6v3tn+Fb+EEsgJkZxhDHZsDXKs9zdCSGg+sEB2v2L4ajcA
yiE9vKK4F/PX3axfVrgemYkyHHws1bdWinKTVWfQKQ52VUVzPTcm2vVsBt9OdDYLspFOLcFVg8sN
I4dy5oUblBK9gQa93ttO393N3QLgfDljHfDwiUffcy0u35oU7aNSOfawabNirQoo26471iGgG+Te
4N1v4L7HHmRx03Tu0W+8At/kKWy77uvym901i1PWJxfcoEjbB4CXzaGMiZLFWXnSB5AVTj7VfAme
wqrEF+d/3WYi3hzbedMnbJqNSHRbnSERra79RcCtiN0aiilzsfyn932kaHVYMVKyjlxBBi59a+YN
lymnQiaPiiYI+FaVOOGTBWJYVSeKBNdvHAihTZ2QBw3wcQasUW4OP05TWASgYDwYm2ddMaGhuQ6U
WJyGZ9s0J5Qi3YPSsaoNDb65nfn0EN+IFgEtx3H4izMBbMwMgX8CRA6JmxluncSXGWe+/Lo2/hES
DQw9tvWI3g5Sm8ahCcROLxEANbspR2bRr+ns3gpfo8iWDDcqfapCskyQeHTp79LUa1cI17iEYifk
+MP3IbYbu7/pLDkxJCt+XF3CGuIkivaMqbsmFfN+vKLpgESS5e94KQVe3a/bnPWlH3BjPwbBGR/q
hpSqu0yYOcIiZXnGvmHna7qOqJcNUEGrUb1PRdO1IUzbTaiaMoW9LM83OZBHeRCB0x9MD2e7CBqX
VwhXYXXMuJC0ALGMOKo3SncVqgz5pm8fx7VzGkak2rfR71FnGezZ/fSXaUdBVDL3zeTtJpta+q0R
RXenxgXNCsfm/jqmK1steschK3pNsHvblEhH2AajpV0vyqUvyQikURp232auAnC6iwokZti8kNHa
H/02JGK9ndMcn5mHueauJMOWRA5ME0r4tfsj3cnkVEqQuI/+xWZ8SRCOW+JJYA0AVVteyjdmoq7N
wzmGyTflzwy8qR5lZ9xCCFoxJbzEVXH3cYU0Rxe7dfG0Cewv1728v8ohrkT+5Dtv8IIUqdTsU14L
CYWtfFH0v213dxdPwkYp6fJIib+qFtE+9cRgRgWrBe+uRZBNd1HGAl3PIYixrsn2EQVqzNlBTU9M
S1HaRVnb3F6jGYibkeUu4DmTYJnv1ELEPz6BNZzFRVZIB9FAg/JpuVKX/JQnoKuVoSA+yqC8aeQX
cDCR2NLqVQFjmuF5NQP6wgJWc1h4r3moF8fZ6YEYVr+JhQP0jZVmlkYEIfwkh7iGUc+5lZLwvI9C
vwP+mwKX3W3mtEV6KMy9Q6o5WP/veJrKx6hdP94iJsLSk+CiySYIWxo+q19eIv2BjBu0sEINplO5
3dJozJHBtgp8KLOcmwombRvElwht7GNOnrNnU8FkAeOJ7eQ8xDpTZBUhAtXN13iOwAQ7a04d9sqK
VmtG67WPkVUKU2YwsGusXc6lv8kJ5l81F4Uas3XKHJMYbKQ2Z0irq8zjTruPqn4OHFkEezsk0I4m
QN5OrTkWPSkM0AP1KwuwxBA3cWmyzsS2IMU445UKNQRYcGxjh1Zna/vH33+CQRDxOSPvdNXo/ITT
e63WpeDqVdJ4O9xFo41osqHQNcWTyHSaQPtMKkU8NaM/FuLIrzFaZyY04PVr9doSlhT71M7d+9PT
kIfsOgAtTIB0KcEED+ennBr/fHiemXWKkHCpGeRfV6yq4P1nNLaw2Ia7jsQLk4kt15A9xKFT+zzc
oUAeCcaSutySZH/RLC9dPzhIF9KjtQk6t77amb9o6AACBm42o2nUGnwSApMsfWo4zAWTAkI3T+z/
zLIIFmp97c13eEZyEF6GoinDAa4zvKHydNXZiMO/WQP+6CnziWciV+VX5/eFY10B5EKvGvZwpvrI
8mbL6r5W0dst0W0qxhMIW+r3CZB8LI60x6I6WxxLrj9efJeXSptVjoYR16F1l4rQImg0UKfbuPLx
jsyOtNxN//qabYN0E3IHd8XwR5eFpt1qU3qAuhRg43p6yzS6xmR6/yOC7NH0vfywEqznfdVvv81O
jLuq2dEYE0hh6RkUrY3qKMbmyuoTgATftTBAME7gaC5ppV0G2Zk4Wk7G5f+3+t5u4Nd+KzyFNV58
IbWj3hqlZqApet1BsTUQu38M+k/f0qDpogmbxEiEi/4G7ssqKVUGQURj/nCeV6YXpa+H8lKyhZpQ
ON7izHJqqua43DTXglWJS8bk1S7nBYQBw6cSDDcGFpuRYOpBYUxksUj01YJZWisKnxRHxlobYU9D
NPSTinsqtNNJw76mpcjNf5SA9fkSVmBCD2owBMDeub1lRW3beuaXM/Uoh/Duf+V+JTlMQbKsA3Tv
er7Avvuh1fNNeUE3saqjDej68ZuFJPbIlMPJc1302wuKAeNGnJ3mAv179mItmIKcyvhFUE7CALaM
D8o+jY/2lO++FKqkoQ8l5dsJQPstuLkv/eM7+R2HEj+mQiUCIVgjENeQrEZVMPJiqrUSxbjV95DO
0hJ6M91kaW8khhSDOYr85FuMi5J43ZTBxqfhEf8ozD2fsMMU8sK98h2Z70Kv6dzOb+VrbX9JJbO9
t+7faZ8tdbJmBDGeQ/8jYLdrXYfZewEW0xihUHDOijjUo9aVynAD3zWv+Cm5k/MXe7YYSZiRPIHX
654+T2Y3ryzmH+/YGjI4MQxwKSD8NOEbSbkKuxfIIDxBjwIrz1oQPUxtGw1DiCkHKr9cip3A8hnP
i8gIBXS2RGbp9W71Je42T9513dkJv6aKcN4t45NTecJEYENbxCDqT8mum4UBCndR4m8ne3hTsf/S
32nl5ZQvHU4GKHg4PGfZyRwMLcRIMAG+E1lubFiY54fKQ2E5OxG4qv6EUOFHawV8hBxnz06TY+Q6
XstMbrAmtrHNgwJaADS3jM2f/HSHBzT6ZCgCuMERuUM5XS7w++Y/oF2nPaNTgHtaUa+3zdvh6KMD
mgXzJvPKFWZzLMMW332wcK/woRZTnulAcqD6WPo9226iBhCmH1ZxVpAINMlwu29rGSGJn+NvCbky
jpKUaqqXc9iGz6umdw4MYSyjL1MSKRpeTqp6kY2dPt7WZlV3IRONr92lTH9qz9CTwEMxt/hZqCD/
RGAZtNZJ4zaPED7s7spfNGxgX55nON1WJpTsL29+8UjPFUcTJebgPzb4IJpjvOjPv99gPy06HKnE
eskOqTO4iNOVK1Yk2omdzHL+i81ZCcsUdbLTN517yljiiVS0HEblE5W5/E5pIv9Q5tsEtZCamMjS
FkJ73J43PGjryVoP7DXztSRdpSAl1zrZ7sci8xB+AYOzamjmZz7j6YedlBg90JCs8auDmfx/2nB5
c99MZ7Bi9ArVVtbsxIju/++bd6WoPVnRIGLLQJOJoSY/SznpRzW6WdQHbRPSwnvsQGImJ3bGgGfk
2JFoUDc0YerTjXsDvVo+PYAQJzczxyc+KdIiQ+JE2sgIcruYM63PrtUq+Wn1HrtDzzGmgEiG7ZpZ
y5gX/vLBQXI3a+MYj5fBhmRt4FaJU4fIJQS//Ilpm/f+Ah3/sImg2tJtS8zUXDmKbmRKG4zPxgHh
eOjtzEm+Z2NL1gaPIpeAkbJlx6onexnF7sNr6YSSBIg5TAjTOgEB1Xf6nOl/f2QrBEc9z1fG+0Xw
t9Po93PYxVthmc0M248gqfwH/Yc5OitLn5BTCfffvzBnRsRDZWzmf4MH8veevG3g8myluURQAp5P
ZBtbzKldCFLzkTuKeAXKn2zgiJIgVfzRzaGX88iqFS9b/7VtGGf1QXaTzhNKknkiH7LXTdUXTfXN
WBVHPU3mA3xC5aNbcZbUwW8/vMNbuI+IJlxiesLwz9m7NeFuVlS0LntYRKRi8HG/W4g1dU88ifPy
3KEB2QgvFaR8l0LpoeHK5T0qadgs9Rr0hxqb7vp3+UL+yS3m960mDYeAU7gpSmMmSPHpGSo1Nyss
2MR0K+5mbMdGokDY3Ug4sgF5D6W0dKxS07/Z0YoF3aQiBxcmT2zlXM7G2xRFO/1/NeV5uuVma3EG
MJxCTRAZi2bYnA+Prl6sTIxmyES/PxJA9DZ95wjm3A3zU7//oG99wOlLrWA3oz3Ck3iuEmrL6VU0
PdpPbxMvCQBEbx+1pW6jDiGqXO759pyEYsWeAqMQd0vmEDXXxbM9hP4bEOJxSUVASu/aID48qS2I
TTF3ouLGpKOAizf27hgrRcW8lpYWxSoFKV1+kKwXwSjayRDMAdPM6s5OXP2JYPnh20rGgIc+XEGM
SSOQD3wtrXwuSKNgffDzo3phzdkRfGXzqSGIV6yA4mafjnvbqoWDoY8FAoGKBGQ0s0pVSDor6UYC
cBR5wblVWrgBvJ1xtRLR7g/MCwTLUiBlA9PEaj6jAVqZT0HARzD0B6K14FxdvJVf90so3JmNWdmv
i/nrz+iVXp++XMbOi4/xeX/arZXHpnVKW1KeE5+eqmk7hNYFEF8rNdxeftXPzEfCD0+Rjh01vEz0
51mujIK8j2haqx/FPNXfDhP/le2teqQEgPEqfkrhxtuUzHuLKCO14IrQUukyUnpjV9b9+D9SU7bN
J6hgble1JNnUalo+g5OaS8A9OlE/QkmDJjHHuPK7g3lGCTAphPDpiwAB7SEAZqDaL0XtDbrYEISp
olax7wdK8ElHAywbhWJXuf+g25tYCvuRYWa07qRYtbURZELJ3/gjL7Ly82StdUtc3kp/ekxEboOy
A6XgRBNsP8FABaaHWQYL0/gBhAqWflfoYG7VJkxKhIGHRv7+qUAIFtsVOvj6BFLWsIZxxcve6wpP
3cnk0t1iDwLCPM1JnTA3eN8VFg3XwqDHcfCuq95hgejv3ONX/SgOxin7vbeJGbq5LMo1t7aeoabU
Lz/EuNbQRqbZ1EwbVUCfqDjJfB7t4mm8D+0KGwdCdQJM9NApM7wekr6U54K7xYeJ44JFxwZx0VUq
ONoHYsMAGAU4nHAEpvAvgNb5fVSHaR/DXEz0M2U5UBy95iRutgOXkyF5L+2wZT8KcOJWWJOGnKHW
pJJjBOxnQVpxfGodGLrvmkBN3Bsubl+3+nkN414FEH0HO8VUSGI/TwsS3ZRsRS1niyYNq+7yGy75
6aG8bIYFmzHRZdgc6JYy8Jy/xuoju+RzlzZ7LpzwMDHGXOJPLgsVQ4oMiiQEqzWAqOu9aIMXm3tF
8BpW2vQ9WAT07yEaNiArgVERXQ6uYYLs/oGR1nmwUvedBz3FGAWW7YpThz18Iy2fPJDP/hqyV5kC
3XSv8nvyxPjniKlKmz6aToP1YwIsXZyjUrIcileCeJdXnuUVgIm1b94e0zxY9QnGZ5oGIIr7UbQW
DSvF9OPMqSgm4Ql/7iYmEuotL2zU+/Ea6hh0oB/I8kBP50euRDeMAKnDmDqWLO385NQI3tUJuUkD
qwqYuHcYbsqRNInBbEdrPw3aPsmwI4pQKNwNiW8gBG2PIyHXeYYEzUe7/0WCTrGiUO3+/P5V7UWF
cFBgUghnr/ku74QHbMK4CpsW4fRMuu89M7M4I3EIrUmuXPcYzsYaUdaooMeCtZSMArd4Vh+XeypV
upU8yHiDEJKmw9H9j+WDCsl2nU1UnEENNbI6ltNM/Lg9F0nPl71no2nzgGhelXKkHXm5vj4998GZ
zK9bEqVT76OIufwrNx+Lvq5K6VShzzYY5jOrEjMHiWk8PmOoeMif8Fl5NMw0zUR58+1O7Tqxzh4j
Q8aasYQzAAjkTiR9y67pvhz0QpzsBu8hFvluMONvuho4gRwtPz3OyE5swW28pI8oxXJleNlgGwV0
+xBvkDLBl/8CrCIymbKrlUqG3aFFp2F9YraUYnNHChMTgNnwWC+sKvDC1GdFxrTRBuYSPVt/iJET
38rVic+/acXmLGhmSqe71Zcj2Ke7XTWt5nNm2LB/MWvH5lSqAZHr5QhCofm3Hn62EgEoHjI2z9dm
XTNl/ObszQ1d1gIpqHJ3vTxv0wz+0m+HL6DUecNL0KbTKBbnAYb3iKd6aNloG8jboblycJGXju3o
+8Ag5iZnMO2hZJqSFVpPjQwS6+SygfEM/821gI8j8mt4+09SL3oXD59ZeXvk18INBEOTbLWiHjp8
4pBRZoH6WE/oe5T9P3b6IQhwPzGRtXAKz3qkgwHprTWkgxI4i3LYDm2yf+O3X9N2XI1uyLqUicSD
wAfwLlXBbofAtCXUFLVLioZaSG2pItbIo8SPflOUnjIohU4Hq+wYYt1ft1xXXXgzlE5ePL0eWadm
WELQOgh5lvyiHPBdy+6pE0xSdAPDJM95Kn7bIhOxchu0Y7XNSwQoRzqf5RlIMzN9/TkTP2KKBD/w
ozwDT9KvTh6Iym1q9mKKiqfq4HM8WlcsKOwRoxiAXF+Q5VwRywfBFloyXeY8QdGZKhnM3/lE66Cb
9dBz5sVSVl7CqPKYJMOiHNgU1Hi9PgRR+FKAm1/1dU4TTGSgGWo0w5duiSrNa9r8Wsc5nf8Z2eJT
w7n8HK9SxSd3CFUDqRVL5oTJMAw9KfYH+TikcAdgj8Iqjq/duuXqIzip2qW68CSjrQFoj7msQEdu
Dl+oGReUJbsaJ9ocNRS+yYF1e4VpAGEQqsZDYxTfyaco35xcpO0ZR1A7d40AKHWImSsQ8N+9n0e3
405xWmNSedacqx0i3KW+BP5K5Y5vfNsoJfJKZu5CZ2ceiTA4UTvyZ2NI0hIqbHGWmotYW6G8dlt2
4BI5fnP10h4bt0qJaI1bC8vRFzojDw/TB+149TCLpjjQ/+WyyaXeWofED/xdSg75X/TDiY/10bm7
8wA/YvLqfPRcOlV5GYfDvVUgQ+iLG9YsUHE5YAisnzj++k6njQgDp+CJ36dJfi+jYm713Cv1A3kH
K/8sgfpdtV3Uslz4fsPsHtjwu8tIoiNPb/IrSOKDs6LFWbKU6+sVYFTvvFiI8341SxIDZrOreHdT
25tbD76H+mYlQUqPBb9+QyfqGXCrTSwUOIIgkNDCtle8g3LSwpZiER7s4hSslkEyPB5u5YOmUZm5
T/Wu9Gwc9C8W6qPsRpw1X50IwMXtDtV6vGoBLgmXtvKCx5H1o6b9tH8BOPJ3JEhR0MbAUTMA7PqA
2Xhm8/kexyo+UMABO9sRg/p6bYdBYQcef9AEVjDwgOSnFZyNe0wkAr17jZCK1cLpqgWcrB6dKHSX
rqBfHzFd3iX4A4wtVJOgtOLq1K+g2xrFHbJFR5VG/vp7gl5c5lq3A0QI0t74/NJmaLGes8vOJiO4
ED8pbjSMptCMkVe8oncNWnJxZfwYG9lu3H04zeWwauzr/c3ergl2XyCZegebmHjKKhqeduwGe2XY
X0/y99M86YAjccit4hO+21mpxLuUg0OL3t9FBxpRm0/SmVUAJdFolx76Lt2MzKBBMZqnPOuRnpcR
CHWhVenyTpRm7oloJhNMWwkxcVNkFvlGcz8hm6J4gUiqXPlO/xswT33GAMDWDpZt8RVCnIRQYtAJ
FreAW57q6n+8tWI5xmGG7Oik+sIhsJEOhwd9Yqc7yaUJHqao2GREztHsXg2Ha1pNPYdR4S9up2zl
swbOSgbK3wHsQWxh4/23G3twmrU3SsiU2hF/b4EQEX9zwuWzbnZRb964BWjJw3U69VXqjpnI1pCK
ArPwxI6X4LXSCcrPgM/m7OHpd5rtne9j7QqxWuVeGM6iFNFX9egKnd236tLEXbe94XJ5oGGm6sfU
X0nlNnTrhdubNzgjtIcj9J0x1rSMn6Xqvl0tyiYrdAmG+A0/PRyEe0Sa4R+cQoRXBF8maqJ6w0Qe
nvkwPZ3mSknQt++un1kP5ZnSLL+rI7/OejFwUzFLJCmTsSIixJLOVWMJGCO5iBl+KR20eKmNf+Dl
HG6dg+gyeN4t2AF5VJwanrvouWVZtBD7vrV2U/UwK9uWlmVmUu9fqZHaOHqa8eMLdOPKf0+Vqigb
ZrjxKOZC4Nh3X8EKqOhDzCB7zdKOnk3zI+rPpYbK3xXglxG7Amu7tMb7MEoXS/3m2a2hSK0/SnKu
WBS+IuVBzcKN24y8CqjrpZ2wOz75ftpngrEdLeNCHXjkjznviOrXjVEex4luFQoWcqacQPkiZRfS
Iu/kxFHaf4J0oDehTZjrOTv52w0tnRGCODwX0p/hSyB+KVRoRUekSHMUEjYuh4MYiT1296yU2Xap
4c78dYlS/iB6iTtlQtK2T2VRDNPi94fRhRqeIZZTMVN6dn/TSKCcyVxEMd4GPFcFG+uUAYWgIjjB
Cq0OIemIRSo8w8t9gIWILFcf6mWRxR2KQfiYbT8wO7lv9B2VM19vemAsz5RpjImMgA06stTw7vGP
BbWswxeUJExAopaBAgwHTak6B0lBmlHw1S2OJnyjvHQ1Qfe+EDXQNrBN8za8J09jyljwigm87fZ8
LrmGriro8qG3OZTcNI7A6peK0y7lOlM353XAvfIzHYzWBIOUsap0w9RIqkqYMihVyLoMRiIo+7Zk
aP0EXW8Cf7nZZJCqR3qWwJbBGMP4pTTuyIC6M7DbkjdZHEV2wjIywxWhFmmlkybBMHfmcPUm2B20
I1w1rm1y5Oa7FXPfWJf/aojsT7FFbMc/g6Xy7+1TFpy70Rj6epJf9PsokW+LG9gnKlAZUfML5iWb
qtnrF0X2Ec0ydD6QfROHZo5fZtS/H3GfbHyd+IIk8OLGJ22RfzqBQRJPyKQfn5gITV5v5khCX9Ot
3mSAvMFtBcvzm2E0+MoHC75P4QhcskMiNgbIE5VnjRjseH1/Z/dLrlI+im93Xp+/I/vnZMxH/K6T
eEK5BqMA99ayzv5r9FdKh32JtX/F8KaLWIwHq5ReCFYISHKMYG+fUJ8ua00dobveH17xaVvfcPL3
t5cNDGBdnWK0UoGk2GQIRNV5QFry05TG+atAe6rw8CiZX9rxnnY8jth/lWNqQ/EHbPBoCYc6ybmJ
GpQqTjnANbtrYZCrwr1kFBMcdR4LRavnjnkB6BVF0j3SIioZqWysydYhuR/xsseM+/8Vr4IhrCYI
xsOXzgCC3xUCJMDhStxEctTnv7PDTAP+It/3qvvpyqbqULzJrqIKxwHTYJjw920xLCpZQ5HQQRwi
o8FumQ8OEceHd9aaj6KOlfYnErJAOFHxPqb9y0xwG897G19QWJXCTndm7rQiTAsTibTUixm5xgXG
4SB3srrmFj+irQjzJL0bNVwZmNCEz8lDrRHzkQCniOKSrgkOrCFL+mUGEPmaG5bPdILDjZ42ZonZ
bVdq5rDEGQ0nobNZ37BP0/d3JtxcADkbWM/dYewwPaGrbcfUeHKkfbEvJX9lqe/JHVqZX7YoTjPY
47EMzSna4bnyPsFxZpMidZw+I3Tqh5BfmJDReby97xziDpD2tdp6tvgzqgpG4vGyxT+2QXbHNQQa
tbuJr26lppNB35+ejqhBwPXPt5Rnv6SsCIra+29YE2bSUp8udzpp+DTQt8GCg2owjmY/bI+Sdvet
LLeJhgmI3YbhYKepG8olNBDo83SJFL6sY/CCKgKZ4gGOQ0GVM1NzI1MQqfGG0yUVRhmqai9r7dlO
9kCEQZucjRCKn7Gf3KgfErvAqDRuoCw46i5lqo9LrXybz9EcVxzO3K3WbrpWpMY9lrMY1oJOcYmo
OfHU8Ppi6PvehgR5TffYi24BRGVn4DY0p1FTZFxwUAISDxsD1C4k2f7KMWX3j55JYXlbqh1S8u4I
mNjji2FotqVfjt9Uua/6wvOlLqLi7pkP02IXfCFwEu04ZE0J6sxuIL8T5hO5SS0lWQXlSHjOOppY
2O0o9gx7wfmgIKJIbMTCU4d/siVSIGT+YkO17ICy/YBulPPoabDS1KEFIxmqVvBI8uBpiSLytUxt
fkHIimnEX0qwFn/M7SoNXsDCioQFW4Xnb7URU/5X4DLRCzWub4K72CYHXS4ULVYruziy4odd1lQj
LJh1Dr1tHSPFeS1wZitm9lkSbEmYGoa6/ySeK1P0ZrjotIFQMEKd4Fi4ck/5UyCjJ28RkZZwZpWg
JlCxgm/9J6sFqyTbmzRrEET8d5K5syYPXv1MqTzMY393+UC/PwJbag0snjO+ZMHs2mUgKBPXPc83
AXjSwt3ocpRGXuaiEka2ULl/vNdy/r3LFLVpf9UdrFLzp58tVfFuCHkRhVlKUAQUVJGaJfm8inuB
gLSVJTJJZrvEVChcOeImka8UzgEDir8u/3fgWDCh3mUJVbXemuejhsHVHzuOJGrBmOTd6z1mdOa9
U/Mz9YczyuTfv+H4T1DzTxugM1Ca3aclIAhEPEoo7mZYXTc5jO6lQFyupI8ifyKTAP6xQSYXTjtm
W7HZZL5JtKvhfY6Drw62tbi9R3/L3Y0qi4xE3SC/0zYEBa52GFL8CWE0VfLKNphgaCyxYMiM4Hf/
ujWUPdfL91UUEbrC5tS0EvGznMdL3odLJ79NR8bQl078pIGBZ8gEJYU/iNEnZ/g2Ehmdo7Nkn6OI
fuCh4K9mgeM2tM7+U4JVqH382+ItS4tYhrj3gn+LFSueWit0D1z1w+53K1IIPf7hsZ3B6AZNwH0o
ODQw5hDZlmbTc8mYKuuPPcWmuxb9VwosAEs5aUVMvBlQZBM1Mb0t7aQNVeRJ/pks0a8lhWTX5qEk
i8xdz01iEbxWDnJ4ziiW28l0FINQzf4xlFgBBrsZKz6DopUhH5iMucqPJssKyx9jp2/PWqOyEHCJ
qQ9HJgC1KXlKgJCkP+12UFdPZcE2XBvwIfXnYqD8jV45Hbvoz9S31/+OteWmQDT1SoirBM6uRmsD
YtlwYnVLsQhyKIBTFNsl2P5GQg20ZUbgaF+WzARDLGvJ8355znyO8PgLmt7WV+qRNv0lj4IMrtWI
3rrqbXJLLdiiJN6aksJG87FXxwhQzs+Bf7QiPphq05ShmrxHiBnSG6aOskGcakvWwQ/4l3rnL0vw
+NzTstTpaZtjNT6x8jOkHqNuCjOYwgbNNTqcn9CmveAmaefugNDIvTbWKdRTm+wfiWaQxokBGhjI
BtE7hfQqdtlbxAzjZc6F1o4A1SjPdiiTMj46BB4NLLstdvEjjjE6gG2PzRKlW8GmeAsr/30OLlpf
TvRVx7+CdMvR61HqdumSDt7XocyT58NYCy4s+g/WbhN66W4/1lZn2VQTjVoBEMfLptG1nAmps/Us
7NcjNNxHl+cNFk2YljbgnOL5a9rymXJeBvopBMxJ/rykZyfxyZtyl4ssGtwDob4zWTDJH4Vd8rHj
JYyYZMag0r1fgU/lveRhaWWvi5aXgdTOtT+mVBvwFhBkp7v72iYGdzey74CNpRTfLnqU3iCmJewi
1jr218cw9KfgJ1N7xlV+4RC4QK5/9hRQ8VyLQGLZqGW63Ud4kmDTN8fMHIx5yxzhHhvMWlkrv1zT
QXfBLIIdgs6SxexjCjfCxj4PiCSGRCY+CdfiQiWu3DJIz9tOR7gh8VylLrfjpuyi1xiLPMpaNJF1
EouS+NN+9eM0yl0uto6R6G0EVEU4rOg1NOgoOczA4c9gSum6iMroyscYpu8KzYpt/AmqL8xnpGBc
y8cGtcsi7Sb0/q4UP10ksdteQHq6F2T9kls2Jq6kpzcnqL1dPfVZ3CoxNibegOrzb6paPAc6XoRz
qW0FVs03T/wCLBgqGzOSsb6Lxcv0sP5VcN/igl92ccdsi43piVmx/FwEkJFzIyB67ZPr4w9HYsO9
0ykcidbLRZamTRxw3mKo7MonYZko5f53Gz1YV5ey2SK15t/9P6cmBzvgHaAP5vTQ+5YYHLtxX4jz
YJRW6gV73Co4l9gFFlT4W+snRzqkXGkt5q3s+kbbTJlKtm2p5PPBAC41RX5sRgEtwVeYqNN3rwkm
+/0v+xe+sbVPPLP7l6DW/UKyZS9OvL/bTQdiBpWYejlrnkRMbcy1+Q5Zm+ZgY0UdyAIr9jaqe8pB
vnqheKvDfvz4kk/peePszAOYzwAuwEUSg+/r6lA1PMu8Uf5dZbiKyxO6VlHzOStH+UyXMPV2VwXv
fefyQ1CWolLjjWK1Yl5Aw5DMn0oKLdKzuV+AbHHwGvdeAcIxNaVDBXuhXzSkSYzpHK7ili40KJWf
NQv16LTCdDeT6/+2DpyhqjgILfM+21BSUlt2Ev9LYveDR6JSH9gg4lMxB9EUmZT1hZYDVmdRHRZO
aJcG5WD5qcvVdVWeF4LnaZb5BNl6g3k2fGqqHtcNbdTp+DT6TA3niWKq/pCEoG1+7tRQKQHprQ6N
k60+0PHsfgU4z9nNMdA0bcaSKsKnxZhNF+2QUauoP854YRrpz99hNY3tiL4uwufxemyxk3OYC6Cc
Bki44c5MN8E5+xWq8595P40sWH5Yrys0N+qhzay/JzEV94ztideQN/NgjC9PHO3pgrPekVULP5hC
KAdWpZNCuYZ+dq/FyZ33GoAKnpiw9VaEr6pQIRvlG0mKSFnkj1wsJ/fRDlv/dRSD5TDyJGYadOi9
0mK00TSb9vEDuQl/YyRCkYZyKQi1oL/HOtVwtLRW9R0o6VLiMTpsG35Fcf1Y0QEnsFM88BY2s3dK
RArLfDcaUFvSNsUsWBogrF7KgIKcaRNtL8JQn91pGLzUKv771xsgwCPjfD/gAzqwlrb+lIwkfavR
ydKT4XIfUM9JIE+sCeeMBo6mI/jjcZMYthOwigFc62LoDrpTZH/CR/KNftvxX5JVLUHFQz0FB14R
FCBNtIByAD18H/dkOc9tViS77d1s6gbL0TERuUxlmUyeH9SGJ2oswfVHzcaA6JH3LbOAR+oQAs/b
5uebQbJLI8M3KvoCBBOPh0ymX+ANafJJt+bJRVlH0j1907/4SUvFttIcunpq285AZirJzgL1NdWr
uMSnq+a1ni0QZ68wInnjFdxko7g9IuIzywZqcOKf/pp5L1ecNUt8tpRyhx/Yg49j7tHzetR//RAM
EDYpKikhF567S+S3+YrhzQKptgRks9fXA8po3ykb1M73U1lWv7rm/ixBmAhnQ0GPhs6tyzZxKPQq
+QuUoXyftCHH5NiqSbU2lazG8ADUZHEvijv/9bGRlFG4+pMePrsS6yfEL7et5edzMVZ9zVWmaJRf
i9/9NL68yHVOGu6QUO8NCpP9iZziSGtDvlB+jhAWbbaHhrIKyMKpgvHJ6Vn7tFF1SnyWFJGDNzHP
vB+zl5SPvaFw/26zapPpjgwbs4e7TEvnvTmDw0MUGOYutc4mz44g719vDzJkZdVHPB+RPzYHCsxF
j6aFFi97WHEPw0WF+BdZsHXxy7uryx+71k/G4MCzOIcaHzGDDSm8UtfsDmdkMmDB/T9Zbc1tvsXq
HMk1Gjcf6YBPr/OGWE/QzAgNE5xVtRcFi+2Ypw/3GKAwMo9ZdNbnZZPjajpS16nVSZGvSpZ+aB30
OQgrTmUtsMuOnYnRkuNpanYvzCPwg/GIzDU/rw8be7DV3eNvVE480vom1UGxtpNtL/QYwmlgcedy
Fcn6Hb+o6u6f6a+FRDUscqqr1R5qs9NI1gRpXvJVS8BTap9fHnnRjyN4kfmMYAgdl6+m5xCf0RHZ
9/sJlCGEhKPQEhkkLdebEgitHviEmRIalfq7lasFjrYIj3Jb9/DD0SFNUkYh5gUEo2tAAkA5Usrl
cVHXJtGFa5j9OWrGdnxwuu/E9IiTHrNT4AhS/VTcPZF2h8teJu1BZYZtAk5GiKUnyJGfSbTdpbV3
HCxvcwnM4LcgV7eoLpErVpjFa4as2pIsGYh1i9gE28Tf8pWJTO9PPfn7+7/V8CI7sLcwHTR3/OQk
6BJ9QWJkVVW432FlI859mA496nYXgc9BbweUAYk5WWyEBrdc9dRlbeYqcHWqbKhHwTP45T0r2orH
ZGLmy3gXI5NtjtIpehmiGDJ7D5qVFWn3zqw7WSHNxHy9yi2czprtdqNZ/e7phwBqPxewvA5RZSqK
WO7HrHIMu27G5ckwMlxCiL0aE0jWYlJ1dG+fvLZg0/xWUJCkara4azNC8JGhHuRJ1FBS+U7L7K2B
CN46RkOLQTDlc/9F71hO48nOsE325TsAFiW1tiT8sQFFZcncQA6rSiKBNk8DgpHD3i4e/Zwr7zVz
UrAPmpWpBr+YOqJd+Yl8QsmuOYRNORGgDgBfoVxhN42i0ohZlbVYqv/Ql3x9b+ur6SD6b14uo4K0
cFyJ+UtjbdNYBQvW4pZa2Xwpw4FVb01HmssmEOO0VCmO6JiRL/dEKKO9ztjv5zmxRp5doGg/BfJ5
G54kQtu+UWwfQZwxzCTr8nAs9/FdB0nUIRCS2STQKldbM3YiUDpd62rnoKHx5YXHDoUd1ZqBt8ix
dpJktlbjnQyixISZPiqLhD1xCkWDeJXFNaTbdQB3xUt1ZIhNj2gch5tWChrCEBu7caHBJKQ85GuO
l8WMN2IjO200wBnMrpcleVcO70wI68oFoJGHyj+YtHM4S4Ffy3wu7Ku3o0Xd2AsPWdqX+39j0rGn
b8YMAeiXNchwGa8FudWdStNE1GNCpXWMh3H28xO4i1j5nbuwegwf6ji2KwsgNTYxy95cwu8kScHm
clPCCuXweTf7/50EyHqifKKhEj7VehM1qUQlO1cEQsUQkJMyK/z0jF4izAqwla+Ihz/x+ZOBdMEf
O5qLEVcRnAPvpzfvmDJvb5wioncaWptcI5stqrrlevJhOmEtddVaG07jQQWJXvo85TVniU5HqMXY
EdFZjAqbALYJSRGs1mZLa7Am815bqrZktLtLXXnlYlOvAiNLpU0KiBKRjGbRzRTCc6yB6U73NCFm
R5Q3M0VHG8U/sSyzr3OKxZk7+fLdUK+6Uw8MaQtfbGq86um7Rk34QLNRzGKu72TpgeLCM8HQBWev
BBuO7DBxmuXo5vRpLatS4LY3ZNp2XvAfBU4FK3YmoRp/ybN2NwnDDnnAAquTZDOk5NhUntqkamtc
072rYNRaL6082G9xK/o01QaA0sP+3lNC3X9H/bTAgPgCS7SEV4hnG0H6gbyY9+BAWug/FFm6cgqu
QNAJuzJDO5X0jTV66Mj6GFDssfscnfduIPeWUbrNcNNfCHqzd0AULnTAWor+5Y24EA7nAYRwNTQI
RtHd7TNpXl74O+7Wab++MZTrbwN85dYiEfkcJ8jcT+dzEtVL3570eO8g9naHjfnviwIjQZAVtk6I
0IlfkO2itjLKSHO7JTK8ncqpIJYPfXUFe6Wq2Wtki4WuOSDEymF5BEe+JPPDHe2ZtwOtzQxxDShh
rWCZqIHODhPb4WYF4lqbdQdXXe/mdZM8Qiy/C8UjcpSKVslmoywFpjbp7oYKoZDZL/loLjytETVH
hPvtvsS4H35ieg9lSQLgl6v1PDUDPHmEDsCduPINaC5vqj5PYM4c8ewOzyv4HK57/7xF8pgh8zyM
6iuRs9jkQYeQ8A2mbQcwEq0S0UIa1O6H8HU0MwFTLIQ5ARjK4CJuDgD897N4uhzyp1U//KxJtsaq
iF/R2kc/6GGiiD9Q+CHBzl1T5TK5Yq8ELkBJpXQRAGR/RF7L6TBKtiPa/K3OsNBACQp4a7tigPj4
ZNJAdEC5v71/od4M6UTmtDkQFg23PX9wbfBwLgKMDE5PAke4h7/FPv6e/7sgegNRbkX34IAND4sw
NMBbtj6XgLQM0jsgiO0G5nS9wlsIZrwIyqxhS8g8pgaS6A2sKcWoL1YbZwpsLO4WBRqnkwY/QZy/
SI4BC0qp3wdiibP9sOs6O9BnTuMchRG7wUkcD0vfxokWlP6aOv5H70OaZpYXL4S/CvNonvcbs4Pw
01DHM9NOuxQLIUAD2/BMxgZGgGShpH/KcBaPHl6GvU96vEvlFzrONEMy9QttOpzHzsYzPvYi3u9P
c9HvYFL2YJdAzU9lBRbI+x+YB/8/deOqmIkOoCKsHEg0e/n/fAkDqKKYevCX0tGZGAwtOLDapl+i
vyRYpT1MtqLli/Xikiwru8SQoNnrHSPClrzql7OTjUNDYnJ8tvi2tFcZU1WmrSHDWTCph6HGaqbM
3T9tDw5+EFyzQMtwFoxaZAXyzvcPlJZyz0qyfsGZ1SLqoCPcV40qU10RSH7txNUwS8Rad0QTNk17
S0C7ki4mbrr0XDldzOdPjmkq/uqwm6zoJuwXZ+fzNvpilixgFDKtXbEZR5mqS0ME7YyHjEfl45+y
nFzPJCu4rl9Balpb8IoxfpfTU0C4xw0CqmlM6OsevDC1lpLwi/mvOGNRB+4HeB8cE08iUOg7vmCa
MxwRvfym2a7gg4AiwMbe914o3xNtvCqQxNb6cuvOD/QM5Z7iynpSUJmLmrgCaeYm4bEJPDU+4lJP
0Ro3q4OeixopoCJ+fC/scST/9N7K+zwtvcxo2NV5ArIskgUsBOuRbvBeHW6J6F4A+bpuzUOUWL1m
6owIFZA105aNnQ/ZoInVtTtyrXfRTXzvTY78xX7qbMlNTqODFq7rYV1iyWeMb0Sm2onTEbOPVilY
M3JKeOGLFeK8V4zcQXUBHlY52bv8xNargtFMBelDG5xUfhOyAQgrkdDAWpl+WuETXlihSXZzQQ0/
5hV5P3r1JvjLhFj4dKS6XH/+tzJ7A3gHkm2+4iY/65xzMNe61Fb5dPGHITcUIB+FeiaNadTjgpA8
I+lfn8Wf6FkKx6N+Ss2LqUETnsc4eUs+XPU7aLUt79C4Z2LS7SBvZPgyNbHbIYig1GXf9kPZxqnm
N17oSBotVX00hIIQrJmmDWSbaO4bDNRfmyynDhbuz3ke07ocEvM4ioct4VfArfaRGclZ+LeOxlE+
31UlLkFiPn6ETfJYmC0H+s6/lACih3yn8GzPp8pQl1X7Ku1qiISrO6DlX3UVmzXXr5bYisJCpR4S
FeM22OeOcG6kVJjtQ2AV9zD00P4mqaHMwBHLlJTPi+dISQowmE8yhvKJvgnBfrny/9jdwixp9oUh
QElp6c1s+7YWeYdXiwonJClI3W75mVLH2LGpdb8GYbLLG37JRMJMJ5fA4LKoDmJuR8zdd2zmSlsm
fZORVIsuP6azScoebZLk+aj2aXFHU1zWB/dHgSlELamrhXAXq9J/AYcvQIA2eJqN3XnGr8U0PaVz
UGFnCCnAArCTy//14j7AfRiMDJglsgA0JEBQ+sKIfKW84aIGPW6qtO9PmbKqPqjTd5lplDDM22Qk
plKtyZnSL0llSK1skpLEMnFpIR9aeR4pjQi7FxagfSs1zqtmXBRVLYbXhV5Gf+K/wOuSll3HNpPF
eSsZaO4GO5tYw0U0/Y5f1elAOuN9zrxX1l16RdC6TBcn7fsPmH7N1s2O84cYECemLA4oG2NuoRlR
6jeDbIfG60blhvssJ0ZhcOwJ4TlW5erdumSs/zr/j+i1GIAkQ8mL1+dPVldwQPximb+6PcxFlOem
LPE9jBtgDUcjnEbScuU+EgOdzA4aMy39AfMMkaaV7batt4jVylpXYEW9g2JJ0B5qz9Kja3nMYzMb
JTcMVSnSgMGlQBTZnjxf0qdNzDd6r9D0am6QZuhol/WIeCSZ4pn6hOzdBywynGVTeaVp0qVICP62
tGOgKEABFQfkd6xuGAdr9yic+IiDU5wlCLGepIByLxBFo2F7CiaJsT3VrCNITcgsVHePWcGW5rSa
m3KPtZXVvorggrR9V2dBIY7gPDaxQ+yr4j+5A8otXKIm3lbVpcBVsrKQJQ8IXRYiPodZ2xBQP2G3
CqbyDjVK467nA+CukqWu8AmaJVI0ozfHFLWn+y/2hm6KJOu6eaPYSRFvCQwEY78KlDJRqVqPKS9R
V/W29z4JSReBTEMyshNKoB8VvB4orqxm9kJiQNozp6WLhalT0g57up6dzboPDSXB52VeGMtUr99I
s24vnBrQrIO2OmJclyDg0SoIRArkKPKmHEkKK/uWX6Y6vJiaa7THURcwnL7cO4BmTK1R6u6D4qph
EaeIgCod6l97UmAsVIcbISZ3h4J3HzRNbb4FD20SZWgxuOlYlb50zxwEcuFBwsl5YiafOmAjK7sc
kN9URuFO2IgQ9L+P1fR3/wgzy8sBMz2iisIN6E/x6E1GBsyhJb5MfAGwpGPuaJ/HnsfccKq5zuC7
dUXMx5+DAcL7j3E3AeEojknu+jQFjtuo27OkCwceS12eKRpVbbtBz7s6RxovVxVdqNzhQihtXMke
5rZrll/S7rJrEqeZVnQl91QS/mq1sgYmTwF+8l1Lt8rzsQFR2cznEhUhOPaoeigacdZ2V83k9sMc
zg0jr1jxD3mVs39ghpi1jT/d7T1LKyO04kpFXn2otYXd3G9k0tkIuDM2WGqYyEasQBGOoO1/6G5r
w4EbpAiPEXAyi599jNo2fDHRuIWAiSDRhOXo7gfKwu2+gx7iU8tN6QBpkWBNVKyJPp9tZULfHg4G
8yMeXYk4b845OTP/XZtd75SFxetLVvzx7PdlrYQ+AA3mklLq7tVMEaQ82iTjk2fZlcEudH3epGH6
spBurcdE4QwtmeoGPGyIpKWl83pJMRUVsQhHpunLdYiyPxyuT9XH88Bw3ueczbGQy1Xjc5gi2DHH
hGVqkni2pFNeD5vSJY0OE7Ziw0HSd7yOTfe6SZGzA2Dl7ZSjsG7RCyPrw1Nob+ZR/NJKF0h7EGD5
2gx4S3uLbNmnWtHC53zLJklhPkqJPYBuXgJoVMvfft+CL0q385hu630AnmwSBTSIna1TJbkvk6tC
/2s6z0uk5TZ+5fTNtkyOKB4YNucsv4g70TJy6CmQ2+af0hQ1LXC/oO1IvAWoqKOhzujX5YO2Q5RN
LyQPcW02cZz73M4wYTS8ZFHoVcu9qTyEAerNYavYLl11ldN+TyUQJTkk2vCSSPBWJd06jcNxjfMw
6Gfp9TCVB4PF870t9OsmjgXRSW6Y19Homyv+AvGg3AKpDKQGJHkqh9vpFSh9flr4z+Nj3xQw4nAL
wqEHu1DqTpBFPm6NU67aXfgga137hVWiwtjAx9TATI4J6zzvj/Be+6W/naBLsqTCYzWu9ICj7pzX
gp+AlqfG1ubFsziaBg2WGFxAngYUG7KKMs0XbG0RBnoZNbstJKAAgvhuYVwm496LeuWKTbWlDApN
BIFebo0juZQZCPzg5jzeUUeqaqhMBDebaToH2d9VNxKdL/Q9FR24INAhylVPVWHBiPs60P+TOgxo
XHFcoVmUjjXwlmm57oVWyjg3Rc2/UHtYteObt4Vlh+/H1ZaajSZB30qrcPtFjVmAPOw69ruCrSyN
by1/EF10tnVBGQyMGaWQvDQEdbRNknWIIGuhKMinbRE7qdpEf7NhdBghRgbBd/STju5YJJubeK95
FL6kL4/mOHrqpgXzuwzQ2GfSEeeToaxsCL1wysuDTcjwIuN0KWtnPPsE59/59ywfLLsE4QSquyrh
qdxMfWkM4zAHnKDwy3QJmu9+hs+n0Z53y0qq75BFfEKwkiQn3/QbsVtqvVEl1/rPxSl3oFexbUpg
ORiXzZdeF9F7wBmVdONR5PqxUfZFPTavFkigWNSvrWqe9Kshq1s0J/pxuFYtUAlvb2xAf2CLKruZ
FnqiLpntv822q6wME/q4jxzfMrKZkmJwjoLAxm99af6d+yAdapSJJxq+Ads3M9fTbVwcl3nch8JK
PV5GlJJ4theM/060y0Rjly6bhtndPMip9mhbrBp8w427fXwBiQD+G3p+bKaGGVJ4oyCP/B2gbBPN
aY/VkoeR2OAjnDYuqjTjCPPS8BJyaWlTa4vxa4mhXBIERsG9Fe2lgCqOvoSzWfk3CYkP2siJLyTm
UT5cx0O9o2bjAcWFdhoYetWLiljh/i008YSfJhj99OganoUidQSS66ZNKNpc+0UUXMcpAc1B/+2S
HmukcbnDKRI/LUzQ5j2oQhDAFIup+vvmWS82oMLXl033ch+sIgePRJbJeM44XxBUhx6cRSSy+qHs
REdh+NCq55e8mxVWHvYAlgWwzhcTLRHbjxVJ7tyDhy5cNygaWosOrOekl1en4BZEpQV10eqQbvGW
iQhod215jx74FrBrPOVueLr27QVM8yMAwxucJ8UtA1UAt2eCf2a0MPb6a7lTQ3gB91tbP96n7BrT
lQfyWYxC+Tt4G0fUnQFYa7jvvwJo/rm2aB9Z+sXcxnoDcAV027CBzBjjPg/Acj7RLmuuQ89bVobb
m+mKElLtTPCrch2fvcdJqUt6O263QO83+zizTFKzjof4/f3WU2HNtWuUoi/p0zZZDSUkC19RH88Q
ddrE7BCJ9AB+NCl/l8q63qfX0PpexaDMJrmWjCrPxZ0Ks6/oWfQ8GVExl/oy4hiOUAddqTkW/mgI
BiAT85O/2V8UZPEv3QRwNmeQVWAqalH5Aiz2IXwhQAB8hEH0LZeIjUObMngJ5AfhQ7bN2jgS/UGv
7dld7jT2KMkvyg6q65D0a4dPkk+2NdoyI+CzF7PW5XNIwEeCnac2nxLJRLtdFpQA9hZoJ+Hvuy0P
O+pz4FRRd2UbCyKeoc6tgYVobWvTvzNrKp3lr1Jt3ECMLIvwy2M/BiDjbi+VU152F/e8zu8D6shF
bxWuZ31D1EcJx4Tkvayf99BJvHmqKcSQeEI/AArXFsiBniI+dOxNWeeqMjvPaaAb242FLiFLlNq1
tU6mfQhbo2m7jubRuKRsKk+wcAEP8yFjSIs6MJusMj5sTp7S8GZ0V9xWTRCOFRf1R5nkaYTBGYIf
x/E3t98ek92VAJpG1hbiGfKwVcqYNlZBJrd2HF78lJmqqXk3ZQ+MqkXLU4T2LUEQ3C0pOOR43XTL
aaafZ+eLUSJAZ31AWHQ+RtPETv9IMWjB8IrcovqVjs0TGHYoOEp9L6YiRsbyz988Dzd44uQcSByM
TP4nWqdQ8RayrDnh+eiilq1volpkSclPfqE4BvRv7NK3l0+ns/Sjl9RMUOEc/k9ovijQvsVXZMeO
Lrxzgnn1mfZGumwwx1zwDjxMauEXKTCxc2waySSz55Md2q5FVy9mjLCPO7n9bziTEx2nptCydTgf
9poG40cIBwYdYTG6auDy7FtfIeQNGtgaUHcmDrLnq4mGL4zAQk5q6jS+oRv7Z6GGR+kqZLCIMWAO
zcut0lJBIzUJnYPy1v1wwUXjj9dJAV0ZutC7FZ8GZ6Zgc5k3w/ln0ObeTp5PxTKiaGaWloOLR1aa
DwSgvDpidVb89g2htj3pfOLxjCLiJKJeScnbths3mU1gVuTUiNInR11ko+KDC++t9eR7HXO9aiH7
Rr1hP2/BDhdxfN8E1zHP9AJwGDySAn2ZeQvSC5mS6CJFfMcFIufE9aRf5Fzn4QnB/q8qshSCq78U
104wjIgTxeLUo3483igIR6ZjqWybD3mAc3BVWsPv5RgXDuF2f/wH7BJ/7Pl5iUHo1byZyy2agzS+
s/MUn/9UUa5Lu5x1eG6LxvoSfUNx8MNhW+rO9T/BvbD/b8kA6LnvqTPeD3Dq4EIJ4tzBPBog9mlE
5487qWCPemhFzdxvC3/ga6wLuLNguthG0J/iU++YdND8vAn7zmsHtC2NVoNcpU06zjQcdPCDv4+c
cL6xFA6rRlh2cC7Ib0+sSZ22K90jYjfM45AmUQliR7cjZ+LwFDEUQMpYF+dPIwe0zuYNMQtkci5R
NXzU8dE6QDeJSynUFpaw5rR0EcyoRXi3KQnYsmJnHU1OCQ6t9hwupYWGRTJj1Zu131ht+KUXX78x
kGYXNhU/CDV29tz94tjRDQzZQ8nZ66alT0vzgGIzK6a8JtmHziJ4QAyTEi8FGANn7TjpGTshjnaC
6vXuKyZgC7uLyBrs87ws44xorA/oiTWWM9YBlnMd8a7gkkFg6PTDZob/DCP7kjlZT4hnF/NXJnJ1
xTzU1W1+dIzKEMxTz7p2aIMfmrJ8Hn/B0IFPaHHl3s5G1FoqxMCRU5mSy+ipKQnFjYAAd0yE52tw
sxuENG+xCHf7PbLdwJt1FXlC4TLr7NJi9FQHYLAdyG4oiBjKNqYwvEOcczin4rROnzqXxfvLpHxQ
qFyKPCkA1ZYj1TI/F+RZMIsIiTAD5oeJ8L7zB1tt/Z0TEkoDLkGeWG0DkSX1msoHOt+gS6affBGx
1ZiPIfOY8KDrRYQu5UsZFLRiYdxyCB9FTrBBLjj8YMf6ExyUatRk+k90jFnSY7eY1vMVvVMynCj1
u9a9xuywmavO1Lmamay8duBkYGqGjKvTDGDyQ/MgPKP+RUbvctQ0kp7IEn490Cc5PVrG0m5/xXp3
+7SgIzjF+yNgW4+Zmr45ZGBgXJXEiiIISwOzJtTNmxpCmt0JvFpQO+PrJIHBBzI6x86+TTVC3TVH
l9X27saWsLyXpINvGkEAo8JmLG3h9Adsrzx8oQOoLTIOUOuF6WO9TtjYCgT9VmDrCzzLi9izPufu
mqxganyL/7mbzDKEYZg7Y6TeelftTg4GeAme1yF8GkzdtlmyWOyrFClThHIYdQT6LpRgghEyIXT8
DsL19igOM2mYhVYaPlQjYc8flYAkZzuD8W9twl/KDs3ruw/lXir2H89UXG8WIiwCvTXrkTWqzz+8
wqXN9P42QiX1RpWVitJD9aqKT7LX0srD0rSMTCV6KTpuB1l7Av+UzK9Cy1s74wReph2AMz1C/pTG
vnLwm/eMk4vKdlAC9pRCrff8L8lcFdKfUzK4B9+byKpWVfPTf+hTHlJ7YLmDGWeH5JBuuiIbKdgt
sRvPPf6vloJ9WyNhMpuhfu6pPHu2H3qKUWKDpF2OxC33h5j7vvRly0yL5XSUIRJehWmwqG+GAZpQ
/xhGcePTki/ssnSx+JGYfZdm9UCKWxjZgIIACECg3yqxs4X8tOPndIFIh1j8F4hgh3UvVQ9GV5lY
ABak3VtPDU7Rox+VoGZ4C/4BdVww+i7CVsHBW9+iQljMXarOQcbSh2xflEUQGSQncjUJSQ7lD1hd
PDll/UkKKznvCPaJ9Y9M0YEeLsS4ED5pJDAXjW3dC3zUxRguXNLL8AmbC4G7IME4lA33UOdiJWal
6iqkTxqG86w6k+USFcZbJs3zEIQAKINO8jmLOPSSQD5a3DLl4676vcAv2844LNhBGsSd9dMao6nI
oAHwGBG/LWnMfjnktgetYxSu9a16fcv9zqLcs21a3t/RaZxyymi0ef/u/pY2Rc0uhWAmPN+5RT1B
KY0EytkLSwhUqYxEregjvan7GN7UFWRzyftumOrP5RGVT4ikep/MK6QN5fvA/7vZEZ7HqwD49ZnT
nQOFNtILiAItM5R9HKHE3hiXEEHLvOO9BwQ2LuIi+yDW+7uzhlSPQz42H7yo2f1KjwvPsNcx2HtQ
RZDxYJbuJD4sL0yceYCApxEPaQc6riKFJw5MjntMCGLMS5nTDOgUVEvxEazy8OvFN73Uym1x1DpM
UXhOhPJiF5gXVBLU1YtkoYBjeCt2HVoWNXZSN71B2EhA5uhBMR771MGd9rmMmdq3uSeLQNIlmNnI
ql8pPzgKGPGtx2ePqsNL/PLZzDG5zrSBdHD9o53S8f8LdNGAz7zo9QigatiuHVZqq8rPt3OEqqM8
SK7OyEffUomeTXVBd+njfEIKuE3YtZ58xk8KB6fWW/hWCkX+CiItMEvvVmbOSlqGXUiMk1SQqcVF
cL4E+XrlBTT9mtpBT9MvtLlKc3U+DV7n1V5UXAUcSKm4CAsnWyVq3mz9n7P/AUUmcpn3WBImJlsw
c+I14osZ27mS4AcyiX9keWRh+LAR4oTaeiKQ7Rg+2e4Nza4aAeGwz43HZC9nY4xyVOCC2/UXQiwj
84780bavium1uB/ZHmx/SiFu6U6newcWDgOpaY1L+w8KXgRPKVYGnLoRoNvBg1NPVQf1Qv7vht+o
42CbSwzl+MKxSd/m7ZSTr5QOWE0XK/+JnJifOaIRMIuGZ/7mc0B7z8dvPgy9biOznaM3JLd7GZ5Q
ZJkAHsW/65b3pCv8fnuXyeyyYCVC79LhWCOQ6unj4QaW83q8AmwFG+aooyQzFNSQL6ZeCqXjKcPi
v9bDcqCTBUrbli8P3Z1n6SryNInJlmOCgw7t1h3U5H3MESLCjOIAvwoY9WkmyMXRuaWpdWdbz5/r
wTCzELxBepxJuyavWz7pe73lkBYA3v+JEqytRzIo5fGkPG4TRGnoXQfQqmoY7oc7Oj1t9GosRwXM
Oy0N5jLpFsuakOA9KCWIQSq+ahF4zkAvGDv9iAVNnbfPlWj1aKlduyvciYU07YsovfsD3H05Qdnr
wnOx525rST54MUtH3zMtJTgtK/h1zRkjmmAdG8qdk40Erol6ZwI6mcNQNda+qrjeBxtl5g2Jcu1M
C3+/fJX3bvQRxH+wXbC/JFhEl8cN/Zlx7ICPuEeiOq2uFtCUB+L8Wz1CqzC1qwoTeYbfIpjiSwgQ
JELlKU/eT0ek5temUGA5NhIWFWXlzkS78Gy1zoQp1tzK3piUpMYXDZAQM4lvtFfDK+MqCg8MZOx7
I5qBtm41vNi/IhLVghfAKsIUSd6+v5bO/9spY/4tSWDE6XREAyGChKl3T9Qd8sfb5VV0htSaKxU8
hwvJwuWZ6eQ8ZN99p5A2DhMphqPce9e0m8j1JQOSxmt1Cv+2XUJ5cv13RcM41THF3MngfGyH6d3h
DrxL5jJ/anzE3BbqePc0REzSpn3EROASISMSe7fOgOYr5C0tN7yX/osuxLIYDnGKyRV1H9soOACO
+ThhADnASW75inE+jvDXz95Wl0jGMoTL++PqS7/RqERtVdCh/KMDTI8/6RbwR6uMtt+s41uXxwpu
UEJK30icpbe5XxTi7QpSk3HqvI8KtkocHkswIj9VySF6vqixcdsyyiLOE2eChv1qIRlRXkzqaxiv
TdPM7aG8247DWazwLRronIrCgIk46fhRHozeWvKpsXW2NJ3vS9vqe1gZ5427hVqMi3pp3Lr0UnVr
BrvxZuy1sldRaqdjVjIz9D34kxtFB6BdgiM0oaA3OZyYoGRjMOJ0ECR2YV0JU2dAsEvoDNhRlpUB
eW1431bigTJ11vYD5QiopNWC/BW/eRCh9GKPYXWkhownAAQTQOPxD+O1EG8z9I4oEAOOHGf3hTmX
5MSIVBqNdc1+5J8Lt3boun8CtJaULDyRC0Gm9Jgt2Tx9qGT8diZCZU8aLW7ma7DupIHS/kkC9OZv
MBqCaY2dHsgpZDeyMbnAVYSWWGa1jd+Yweo2i/HRSD63CrFBmdnFgdiCv0L2JJEWfEzu0kHFXeg1
4joeq206fbrlSnO27OBUXW4wK4jQ4zx/vpW+gNT98OoGaIc8fPCvWnCZ2NLnpPphHoGNRWOaixYI
l9TIvXOdSoy9TZmuQX7TONB2Ep9yFj2SVL1f+Sx4feyDaDicoSqKVbqjs0eF/z4xbPZFHWI/yGuO
XS+jqrGeNvs07AxUsUtTfuMlihUisAEXaYUYwEyj4JhAOc7VVi4wqYEU9ht093PICD57w3KtGMkM
sQu1pCVsHVRFxMw3KPcWHmExg4gnhp/xar+VMN9ILYYeNIqDETolaNNq5FZaWh8IpYlPF34Pjnwd
qWBB7eYL1la84DtOACSsg/si9XoTkwvQTXKfWSkuAhYP647IKsURwwtMTZnpkyeY75Y8MqPSWmbb
1wyEIw4gehbotZrn27YHZJl7acAq4u/M31Q933msOCMXdnQQ506XcpeEfIAk2CeJiNiQZ1t9v2dd
0CentJIVnbKgGftpxwyR1FWR/0DmYkWRvdcS/mZhmNzoFY1peU9aRfe9cCn+XZTiAxRQg5HP8cTm
d5lnhEo/MLufuYZn+pQ5fWH730674ZK/L+HfLVl0udPrq62GYQKUrMsRV0jM4ckRSS32X58PR5Gq
gsf8SG/iA2HzB0S4vIflXxCHaAymwhLgZbjxvKoNkdnItrhse4VjgCDHACbM0onHypSBEr6FdGbb
wFG1gSpe1//KxHhktgCezYOMAquh+neFXM+Al5nYsMrPlK+n2Y7AKua10MwY/HcSyDFx1Eke11in
OuPOCckHSivJ5yk7Qevv11uVekLY4EzWhemqvES96NDajkhuZQ8bnMfrjnogFUSzRR9JVR4zRDRa
DAu4sCF6CF+PaGDeGXaOnJCSh4icYt9QuBvqTY1xg2fIG6MZT4hp1IViZrTEHnAYzRMBkb9FJgNR
+K9Feq4Onp3yihBPKzTQGkudleckIwDwVe2dwkBWNX/Le+pAMpePJYlgzDf44iwTBNVdx2FuUPRR
Jwh4yxDTjJ8R1DSUxn/Z8YmCvqFRqQjBtiJRdKMzGEIAVvnaUPog189vdkfX5uIW4wa5lAfsIuYY
2gsClS3evyqkQn+Srl+s3XoCPzmY0dhvPrig+Ic/I4kZXEwrEjUqj9pJY2nM1h8pgr9jolHXdHYG
EqjUycgYVN7jJthA4lxjWirkimnrMyiyV/6YDh/1kQIamvp85kHQh+yj0AI8A8CRa7twiXLhm5Il
r8Y9gtroHEQBJz2KvyV51y4rHglrk15u0UrFMaiR/iA1y2R88iqD4kvv9murNA71++MllypTTrR2
AsFGD1y1Of/sRf+gSDIdk2pDz2wWWLBKb+TZ4h8tPkmDTv6o0zcXt6cAFvxCAfv9L29+p8mIxDT/
lqM41Am11E/WqfzE4decJlwVoMAI0F2xpjrzzeKAvjB3CkevlFMvkZgKR3krlcdnhLGHWWcRdb5I
U+JQUEB5xY9aqmaXEJJruPJLZ1hT1x/g3RFzzuycvXRUsnWjtkhClXFRmxdMxmxH0NL2GhGF6H0w
A4Zl6YUxHUQZjwLF75RdQS4o21jHLCLux7enSvnD7xVE+jwbG3cZUzDESxTWmuZuE14VjIJilr/8
oVE1011HIPaLwDQcC7apzyixxYbHBNVf58jk2geNQ6I3GpsAhYBhWBjKCpqcYNDdHInnZhe7Vo6/
U7sOmG6gSj0K9SGQVT63Z0uxo9/cuZzi7O770RZbHQo4Lc/vA6lM6YOIKOZlVa83XDBjNDKnk/15
VvuQFLqQAzK8RokyLMLQBaCoLPN3xOTi9bBF8lLkw4hjOsACLLnN3NSTOHEPf1SZxG5+py4zwJOh
tJucT48jBq7l3U/Dk8Eao04f5cRbPTtgA7tWbuI5zh8TE4vV/nOnHCStrfsIhLv2t4nNpRCZHj/p
8W6q6s+r9XnSiSBnGSFOmk5tkRrRktbKTS3TGoW6Wvavk28jdrwKvEssMtw2iR/hkRU4udW9WqIc
9joKSc821wj/q4PFkZytr0UGxmD/+OJhXzJQsitgpQODfs+JGcO7XBZpGY8OstZOF5n0am8KdF4u
Y3tBpU6z20gdt6eKhTaOYT2Q2gJ5d5o//orq5ZGA0mAo7D/MNbwspRe0oEHC4KpKj7jdn9Caolig
Le07Wsr6E3huULvHWXpVjMOyT8xzsCrJBxbR9XcmdcowedBG8sZy8kL1d690e/MlNM9NZwbheoki
ve9+VSFxpBY7U9fJ4uDiGZgmJWsiRoOcJNyfFV/y5VfQd8peMf7VCC0CXLXh8yMJmq0pMMXtuiJx
VkAN9FjlUXTnK0qVB/z0oLajh1ApHZpwJAEyI54fvqTQtTSzK8++Cv/52LekIOFqcfeVgWzddGkt
OPo8Do/UMiCGYGAOCcvEIRH7opxEM7Qb8ePWjAHxks6LyBVif4sD+Yihw5mHsUt+WlecqX3KpTZt
GDOIMm9IhyonnMcaVaicLxJr/4NPDEnuFXdOR4O+9gphZI8YOltMhiOoaODLCYaaajuKQz0Jlj/f
WknDZj49mjSXP3dT9b5/kfwK6qjYL45R4pF7p729wzzVYivGrZON9NqegiXxGedUCumyXzbVW6TK
/6hcNDLFDvJdtwon5v/ZYlJLVo91T4sJmAwHkpcJe+OVsfWlZixgwUwzNbJjdLmGMJncWI+fEu0W
QsJ/7JI56yoLDvV+65SqZrumvedhq6WU61ooLqHoOq9X8sdWgP11rZfNsec/eiOyMIs22guV5TSp
vCYxzA+neth50zxPoZdcy2nnuZxrbeOTjvnh/74/pnvj9MopnEMCV6IcoglI5sMr4gnn6/mh+iZv
gd9Ada/Ch9jm6iOKXFtwTQlZElcXg9cj9XUnkg1k6Z3SwvXccDNbwkFnB8b5i/7if5zsM7Iu0FVG
/Sq36rgZxglvxckIsz9hr60DYVA9pMxw5r5C5Df0RRk0rBMl3eh6kV1ZjYC5gU86qCRTp8sIVXuC
Z6q475e9btrpkkFCkS+jpwDL1ZpYfC0eMW4yD8y0UDIlA9DhYp3fDq5t9vxFJ9KajMN9Q1VBVToB
5OvK/5a/rzomUlJhChbD0D2tyCJMm4W1L1Mnq0eXFlnV9UEMuu3MoF+tAIcXUTCdieSEthlUBnBg
TAGr8aiN3LTtn4Rx8/CjaymJpI76GhsPIGBxVi/pUnn3Khv8pPoqANakqJDnHdaRL+g/xvOT0Qbo
BEEkf9j53CN2fCjUB6HdYUSgX12WLaSdQjuNFLBqPd5we63lHUK4aosUaDXzLXw7xSqVkFR35q/T
mM45wk6XDUNntILNuZoxVw3PgIa7ULyC6WU3uLzZUhGEt3dsSrxoeaTZF5OQz+pf2x2KThELpM+h
9cyhcqcrb7vaX+cEyz4RFZECXReMpDivEFTQFS96V3JGrjgKY8SDfP2KZ6I5Zpv80QivWs+ii5Yy
e0nyYSf+0ksk1zFQmT/aL0l4JXdFQUaMdaEordU92cPPECXvVaapOj1To43tSZoEqCgr46YQe6rR
BMOtJKUna4VlumNTsF7hsf4TQPYQsrxiFYuILVQj9e8bp62aedPoCGYUtPMOpz3PSsloQmF0Kjpc
OUcx8T2fetN+FNkDlGKdi1cw9bUH7SmEOAKd3yMvD07/7E3MW0v58VPoqwLkfQ2/4bTIx7JfxB7Q
Sg4IAYSPQ1cc6yXc36b7DZzmUCy+ycBd/ke9mPo9trS+Tx9zyM1w0ft5D436eAFfIX+VMzQ1wRIH
y2f3yH5zLTmA5FxTKLLr3a3bF0MdLmnBlnTqXG98YauE4i2fA//PFIOLkMjUU6hgp7m9Qps5Hr2V
Pz6Ke6diHzhBQ92C62ObU7TMG+cbA3/YbOe8Y1TT1KLNXF5SH2AYFREsVgnDeIaUdZd2abMZlPdk
CXEZSCbRFnPTVD/nWPb0SwX8I6BlHwPSUpdinGZ5iY2cQZTBLMiQp5aUeTuYTMOJ5OpiXSYksI9j
Vy94XA4Ig+x/tsCGaagJQaLTiysZnj159YvvUgStXGk9GH88EZzn/J45w6D9qQ59wTIceII7nHSj
WNifNaZy96Td4wP+/zTntZg2VDLq3na+ZajAwWrBzfl6nEXYd9M08HWsifj59eeKdxSsvsrSE+c1
dT4l+Bsk9pyFNgIFJWk61/cYEGXlU+AjDzTD4SpzUKU/hJcd6n95Uw/NOW0uvU7Gm+09MKuE95se
1vfhBXt9gDOmI/cqWc7J3uxCMgY5eZfVkJmCRL97L00s7syXgHk3VxaJVajhpafyxqWVs1cqGrPn
jBz6nFuqhyiz1dQL2lPELHU1/zTWIV2Mww/Jjl/yzOqRx3yBH4B0uchaHFE+6SiBW9nCQNS7bClG
uZ19rf83C5i6/LPxfw2BrdirRrkTB+PK7XxWSCWmc7cM1FnUj4fL5zJs+6gdmJ1/RFutnr4aV83l
/ROrYe3n7YAcEr+G8ix96p8xPS09smqF6RsOd1Tlr/ia11Mlv9+ECNsa7Uw8NPsiW8DwH0kDxL9d
BUs9jAzvatFP49ThlCPH7pst+8ChiC5/2umgqgKC0HqUkwnG5g10RJQq7tU8kO3QpAHURQfcIvl1
9Yw9ULlc6Q9C8pp8jqcARKL+DQHsZaNhZ0avmoNbdLTBK248fIGSlhHOeAeRnZ4LCdsvC7cGCkL7
tRCIpqyreEBpfmf8xX4x+ONJBj2KdC9loPxON+x3zZ/mgo4KRg6rfS1A8JRZbDNqhHEXXN1OTEU5
AJh0IxqkgtUH1tlwAUb98k1RGbC+LfYtqE9ot5eh6zKkcK/GvHrOhW7aJU+jAUaOF0T0M/o6/Giz
213/oT/iLRuEHpXatFJeaWP+6wL649yitGFtLcaMcEqe0zBW4IFcNuZ3HnKSYKkAcCM/km7zOP3V
yvpwBPeamEZuYPHvD7pxesXnlc/bBiYfiuGujGSFhp2PWjkafdmPWTxIBk5XcCF5oO8wESzxz1RW
Sf9Ifux+r8ZDqLEUG0Vx/Ur3in9h39I6IP2s3hrlHmFW9/mY7vHUhrFrJLTKu2YrYwUedMZSdQhn
uXjxLPiJDUhbudsR5UhLSwABGA53bNpdhcyWxXrJ8hfABSXOdwTEoZZeAajwH8LD/BLlPLFt8pNj
vT1wT5nPBC/DEjWJovy27YzIM1gXEniBC4IjS3gDT8qo7l+1P8mqiGhutH38bnapt46vG2XizR3/
fbKEjbxSTzIESH0NwJdf/3HdjfTd4tivR9Yw33qb2iMrqiTELHPoHK01XXcC5eQxJq/nlaHO+hZj
Vndle1gt3WIFSYKRkSmpQUv0eQHS1sKJaE5MKhUmZ74KGrFq/fAvVAobUgOC/1Oh2nPB/KSGBdJt
3A2WQG1Q79+zuwAjJS0Gd85LLKmFs3KBSVKqX20ANorFXDwXHe5A0khJojh6lJb8SX8At9jfnUUr
MmgIh8whPdbDlqHdIC3npLiBaSZH4dQwclnAjV8Kk2E/0rcisUjie5WCUYG6cAi7zCpVIf8X9mVD
GspAArg6w4lo4grtMCyvt1BbyUQR1+7chD45tuM5dibd34BYikCgsqKabzdgSX6JJVQh5l4psx84
ypo5tzRCqYnCCWDds1/NJhSB17NyAjo3VAGVV9OrZ3nDc0pKaRPk+2d65bXontk2T46LDXvDN7qE
H+CWayO8d3m6GFgEJtnP6qVt/WqjIjk5Zh/ezZGVGvvIo7PxGRW23+Wo1bZaIhCiBpMJtnbsZwLC
qMG0iXnuBTCoq/IcCJ1PDDkziOPsWuAuEEW0P+Kk6Fm6KPkYRLM7C1uTLap6edDp2pl7+y0Oke/q
83Tl0dT+F/6F608UJ5DfQBNfgx57ooN53r7mOHSY6+G+hLhfMZ00NlAk3h02RNKrDBMAiyCrkZLs
NeXJk2R1tf/f4z5s0CeSLCPwwrCdDj8RumELCpT5UY2Tu5nBuHrc3GU/OkvPy+KljlPYqdtr7sLF
2SmmgjWKPgYbhQFjMnT/T5M1xNLy/+0hSkKLjUWSjgzZyFGcsw0gqlnoUCIQ6YKp+7M4/7Ehh1Xn
U9S8eKm6WyBM/PVo0nXZXU8jnAdgMptt+YF7bXxG/XPUicjHOZdUNRSYgfpgSocnIjNY57IZUh65
5QYYT98vw79Z4mHrLWi+2vCAGy+GVitcmGcRWsMbAnzbJo8a1WC387RA8EOwmCoCq2PadcFzpTMZ
muPEchLiPY0NMJ/8v9pKu85T+kpD+Mnq9ltobF604OXOM1uY6LdxMydUoSFZFmpVBy3F2QVphbac
1BJ8M1Xhip4PHY7pKOfKgSOOkYizeNXwj4JeF3rIco5ZT6+WPSp2crQW/yGRE43SMA3xHXJuqUUs
X3mfNKULdzU5VCLtqymvQlXKDi7+SAPVA/7PBV7jWvaBbyELsDjfvuEHNZGYwmqVBeI3kVJ+YXMl
ns+fkzO3Fjo2vkftT5PwNmkYWyjwMDVRf9RZvQiu6iOBIONoJ/lluayg5l6cT9s5CUbem0AdF0zW
rkyTTTGn+1izzNbEiTT25ybK7AFLL09e2ig4ptotY80oEE5969Ayo61UwcZMvK/pEu10lQM5rhAl
c0LuH1BrNbl1siayDJpYktPqzG2jlGK9Wonhbeb21GuSQAOwwPV2iW/yqeZJQD9gZMib5vUm/ym6
9nvo55KyoYB12K8yhsqNPSp36Y9GYnOVVr2/qAsxI4qvBTdkTKul8H47bMhuuW9v1vvahmqHT4Zu
bb9gvou81d4fz31n4dPMj2cctV9QKTvM1dV4QZ0i2VnaefZHERkWeUkOwU/lwlmyemDfjWuXyase
xPZ1W6OK2W2AjYF0ZUIUxJEURYy+gOseQCNq07knnf1ErdgH+sEl3b1cXFYRE+ntDKjl6yibSBsc
58Y6g34MNy79SEqZVzNVKt9kVEGBXkiWIwThP1tJZDarUZ9QvYGjGic9bfZahvRhilROrYyK/ovh
v19cmwMkY4xi9/kQPmoEme1aczzF+uVO/FwcAk+c7ouKRlvYgF7Th2bG7UoAv7EWEsSrglQlYvwl
eMMCS44Jeh3jjpOekTv/Uv7KWnwNRCi8YngNd9I6ssJRSZUAf8brV8quth+YOj6d9/dbwmPgqcf+
1X5M/VcMiM9sC5gyB6xsZ9uw9Oqze2xtfMOnPBU8m9VfD4molW0zHSsPEKQLJ+Tp8wsQKOABMymi
CPSmfWuBoW3srPJq3WujL8ETrg8FOjBWQjnrD6rxLW6ZnxX5sacnNXvDGRS5I7P3yLFCvo+McWY9
RtyhRuziweM19T7vdexSl/9sNxSrDkRSVJeQQKxMinW3kIk8gHkFfkfq8FXUQiR5d+l0YYZawx+s
qDnE19iAl88XGheDaPeMztXaJmjhuuuXiRZfq+zHOXKJozPHFYBxHuVu8LL4JuK+WmqDcVQ3utuk
UXfTZfRCxhfX6779Urxtqf/2qYL/SvCWB6yGjTo8b2ZHjxru06pB4szQBzII54Wzws4QruR+8rBG
xxMmXHEA8jU5ZtntsQ2Jdy+gYaCWwxWILhqrbKyz18C9xVI5jJ1O/1P4zB0m3ey929zdBvTU+0Kw
bZdVDnPgIvPJTlLjcJ4CH5wvIZh2Qcns5qAA0ZiXLxagXJ1MCXqgLfXXz2U/399ZqCzCh9Ym1lyS
imwkx4PEnwMfHbq9DoA9t9Oe7ldHNnu+BsM5/AGkYlr/PboDnd6n4zQpTXw+pgwD77FvGiFy0N7U
ZVxGzr1yyPzbcndfN7o+vEoTaL9v5AWVIDXbTwWhcxbjNCTWag1O5sl7mSQgw3RE7GtCC+QJX8TF
do1VTDapTewils6s/+9L+OmpMOwtfbJMtUY3WeUYSh6ACsFFI674bbXo8t/dmn1JdjfTustYTM5x
hsd8FcaDc+Chm5R1kZy7bUrPy9UIm5OYLelBw6rSs97segI0z/VI5LIrjcq/kFhENZoBzYgeTmix
uGZZfA/II2kPRzp6lpAf68MjK7O0Be8ZefEGW9IP8OzJ3oNL+SUyaxoy44hAJ3rvTLG8j4F6kTwU
rECBxAX+ZxAUWfFSDpMKfX3bo9vpUbujzZ9HjFy0zyye2Ofs85iLi1qHoA/HKwNEwIG4cImYN9Zd
xy6IEr04PTOv0JhRniM+j5jRB6yZReFkUuRDfij9hUlJ1v8Qq7EDGYSMgG7UfoGI6c2BWRt+Lg4L
pY3wujF+BtD5aY2gDdTgr+6YXeTr9ONSZW8bone4KsmTl9Ayyz/LWnoIYQdUx3wH3nWDjr6WsHqk
1zYr6naipZCG6Ivey6JfOgckrf5MLN1pqSxIABoYiun2HPg24gEanI9hLN7M5u25ErGFH8hb7d+P
tOpF9e5nRF9dqQ/l/iN1F4kNmWd1gFVWKrIozMNV/an+ZpOqOxLQzLll+fIQcWfvAHHVmX+PZAbC
eJE1K/J7tlyML14xrMU7M1MjeEw4c3DprDHUMAf3cdJNxLTpQWrqbZCPCQWO1GTz2/NNxLfrm0h9
gIywy9GGiukjtHvoZAWZVEglN7OtVltAhneXPOvtn0HNkPfa2XDo5X1QuzlXSxYBaCSepWan6TYV
roK/suvrFwtI1Vdv/YQLoIY6uOdoioiQQ2oGbi2wAeZpqsnGeCAdr8/UR6+1DlYKUWtGp78okol3
sRDslwIbd0I/F8h0eKFrYtQqqjJcHBOQj6RVr4Ws2OxuK/VP5igyfvBLvIHYDYSmUHd2p4aW8AFg
RXKNtRPKApPi2MS2+4Lij5hxTS8MKAgmpKZwlSEsyts6sLKPZYzdFPpFKLv5EtOjjGH6h8A8hsaZ
sHWVjXwNLtyCUAtM79Lg/fgqoQyA/C36cBYgWS0Dp2dZOapaL9VpRaafNlyR0u+AviVTKAB9DAJb
Y2Sp5m5kKM6l4tTLvj8/FRt7DjtPSkrFFS3BzOG/IkJR9xqimbeBrJoGYblDBLug5qV6EBn03V3b
Np3NPMA74KDLK//RboEJkaidD/NZnntnC6NTtEZ+SUpiDQ9Hcm5sD0lwLOy9YE3V4lhqq4NmJXWx
WafZo/ysmpdNiHOjAuJjI/F1VaBYSBTWJiASEZooKCSeF99+8qqyWN/M7XB9LxDtO8a8SzeuWZI0
wBHZu8NcfYgQdYCtFNyYS6kT0lIp3vcJbRDKvkTvB8362ABsXxDoS5ozifOJy/LudxoG3aGtja1D
Lz5Q/Cm+92lByIfATgMDLMcaiDplZ1PHLNnWPMO3H+5Fs8QSqksjvYFSuK2/qiMTD276zXxKJkkM
MJIa4Xp5uzUq2FSc65hbVP+6gW+v/uHJYzXmjEuyO1x5+DSQvgOIqKYQ3umoFd5XSuDYEKbgLd06
W/HMa7nMuIFDlBQUHyF4eGXScAKeq2Ltk34eIYn/1syWAthw+/DqYcc1aouBxzNL9tN/ZHRDj7Fd
zyWH3lpksD1Jf0MoSkeHsjrDSHo//CC7puGmjG/B8TAXhXgo5anSZi8UY+u8HEUmYwf7gqqbQLjx
vcr1nYWphh/wWQXWQngoLL6aPqHIuQjDUPUZa2BYEXMH84djVBOnvaBt243K7mVrtklGJW54BThA
4cUTRDoKsYxl8sI6gAyXfPSLu5JLe4S7g2j0DRs/NOy8HiVr8cm9iMO2cJ1T0PNKR++LvjLIQ8Lj
9nleNkbjbU/df5grrzSXKmUDeMyS1qBWFLCKkiwgjxuC8xt7OVey3IcPCfhzKxP4pwJPSq3fdINe
Lzaf4h/4qSavYky4jMpZRN6deLGjlo+QjD+zTY+jFlwHg1V66XxCP2jql79q3N2/4toySHC73buZ
thSts/iuGhq4brqVLXW0yUhRHdZZlStd0MeoqR97d1h7fDYRhtbjF4dSQvFpGD/p9n2t+r0ue84H
5hQEBO+hUOglrRvIzxAtBZfHquUSGHRwfBlhVb46wLJ21PoucNHkHu04jMfGhCfV+v1zhKpQqOcc
L8MCVITWoy5hoddLLqGdIQT1942pHb1Fv4OUw/f/wegvak1tWXaD127CaZrNru7lqYvv4sM72JFH
C4nrShwLytZmC4FOGNgko/fEN4E1nVgw9uJuQ8F00AjDzLt3Mc7rLZaPKfxTT4ClZr0+jtsI6o0s
P4Qi67lMUL7ZH58EofAhyFGH9Y8Xw4+RD+Afny1eC7mY6cymZVIQXQOrKrn4ia4p6iKcI02C2cBR
/uovUb+ltv1UhnRKRYQ0ezj0e/llHrXCOU5tDMVT9Qttvd7wBdq6YcpswJliJp5ukjwP/efygfic
EEsdDtFkpqhMsUXzyiATEhz62lizpRslVFtWvyT1vfW3ZPgZl8gPFyCz3yNZkTNZsiyY5GOfwrZR
Mj65qrbEhWKd3NuWN1XTeEASRTOh5P54yMqIi7xiKfbQenpHdK11HzaXVJCzHr0wqHvjcIvoyyct
lmyQfarRcqgXbO4jXNauvjtVZjt46iK0G4svR+2GD7ICu60bwW6D+1E8lFHxUX3BYTMB+mcjvS3F
A4gsOulqO6/Vnn4JzvwK4GXVbOomMzX2nMACXAV24P0JuHY6r1dQFiZh/oeCYhirdtl5v09EZcf1
Bx0GXTMAR6EbE199xg7iLiwrgj+YLPijPLSctqHWf3CN9bWsgOyzwhx02H75/dzD6hgXim2a9gZb
aQy939xabH8LdsplB6UOM1YFqavA4C30iADlVaeJOk8ceIaMyQfqcwaGv+tfAGL7bNNbqzomeVhO
aDXkwN84RCnlvtnALYZGpozHUcvpxj+cDX+r/SzWdURapqOyoUcKQEoMcM0pclwPZz8GKW1gFCVW
DEwBKIMERufAvhvKPNU26hrahmhhMdgGa1gjWA3T3O3c6gYoHEIbf7/xn/YpOqtuYq8t35VzFlhD
/ihvCi0DwpVd4XfxTv3lS9L9psj76Wf1ipj/bXL8yIy0jR+Nt6AyU8m4goUMKfvuR6vYeCmgsqvt
j83qUgdqAyaz5/CdS2NJ201gI2N3eZ3xXt13JXDVfpt8LA+lD6bzlsESV01yMFcmbYkHRiNe4TUr
A1vhA/8vm30DS/WOVcykV0tX+buFFYnPkkQBxWcIVfYt1UwtMSMUL6Dbj0OKsD18Vv5JUhXPqw+K
jXUNTPrOjfOUyqRA5LLAsiv1/UJGaIa1EOldqDjnwaxvhtBLnDgXUJuxkYe7w18I43i84FjkNf/R
xhYnxA+Qetz4JYOgeZXhKf5hxXiVL/ZiXoz4BxFA62NdU6vCgwpWqk9MiLYa63ArGlpKTtorPTZC
9z4WSpKx7pbcih032gGGqr6CNeGEJ5kCgJic3roDS75QoIlOX9OsED+kMT6TDVMzU2HvyKYnOWFg
kR1JHergGPUKt4JLtgequGMM00TTuWI6Eb5oBlF62hehUDFXFXuoO1P39X3uNSD+Rf/hEnFYQPrv
FJaVjQPhKX8vIUDSZwWLaUVE0VMyRaeLt0By+ul4jnljaEUbkg25xpYJOlPbrIOli+CyaNobrZ0J
dZ7ognvlGi3ysginj1lJWBe6VIdgxNmZTZyq0a/lwekhFDQusjS8JVw9DlABZZsHSS8a4at25B1O
sRk2567tQie91XoI40XJOzxmZX4Re+hlIAETht8n7omak9yiCo1WhCbJBSDJP5b47L7LhhJnYDlZ
AWiI8yRfM/iV9VKSjckl/aMBUxS3B8uqG1flvszLm6QdS1oVdXiciMkcwUziM3OgkmcArWQVUn9j
aV99Uuczzchez7JlYVtX+uXMFHEfUFt/vLDhvhNuzFUiiZ1y1E1QbKcsbbLagu6nDSvLVoxXQ+6X
Dkvi/pMSUPrtWmV9v8BgLVhC6m9S4JmTtvGdJutQdeQ6JHdLls+SzKzlY23QfeJQB2+bisrjQYxd
I5ICuzFY9ELLI1dzMD+zx3L+ANYeygxbaKbKuJJToN57N27zg0S3hg6ZPBoEPDzGCPFNtGugWArh
3uWwxFjaVYllSZOeD6kOEQke4wEIBwkGPC4cr68Y+IL1HVGThT+zcsMK4puNR9hh0BZqfLIvrGTk
A6vhFltq/A+bIAzUbSBhmu8gsAoe245CjFXzB0kb8xUtXmCkhQ1hbOnF/KcGvxNPjf+SZcQs1Ka3
jzJpC4R2AoXzte/eit/8DqOECQ9zcJrT/fLokag/OavHQaKD57zfrtVIXgcl4vbgsOnDh6snqzTb
cEu3P7z+i4IASzd+KiTgDY8tHgKJgl5F6+oDBIGIKsW1ZNyeMYCCRMNXL+mFR2CxltZZmzHH3aPT
yhCIZPX7jIh4XiYXFn5CQYkEt/z5qddw2X3Xu1JPqvtiDW98Dbv4MvvqE04CMyU1BOq0l6TxwPAT
V1m9h9X5UgXjq7Nkk56BQc+aKPYlHCklVB25o5VIw+N9TOV2eO73LDd4/viZJUC+MzBqeCWKRTdo
zsyC72G3CjzLJHHLeBs+fo6FijQTiZli6TsjpjgJQltR8ueSkcTmJI9tJc4cc1uEOO7vytMlYkvj
fD+Ji/wzErCt2xbJFUQ49xtFxhYg5w5Wod3pxrjM3gN71PdoeuanBjLc5EVSxvy9NzsNVZkmNaWE
xpU+6dVcbweePMK1gGcEqK8+e23p41tQ3oUonykW1l0XyQSEXAMRqToZaWOcVVRfTZ1fJFGWb37X
wqhM3n5TGpcc7rQWLNTnkONJtD90tN9IddiC5sSTHkmblOOD4KsN3iLORETCGGUlKww0CQfVKStt
LocpjXaMRm+6kMFjn0c0Pwfl7MF3OLilixNFvfrWMS+Pnmyd/M8yoLwEI5nCud4TU3d1lmZlXJHm
kXKHppjwKitoXYkUxO4jkm81dYhZ2Me2uzrXgexzCO/r8NeyUi7QSAadxtsddl4858hZO1daTuhO
qnAuOJ48+w2p28UtwQRBwXDFDAj+R1Sr1w8aMH199brW4ARON6REHE9jPAU5/APvVXpZ5Ehvhk65
gYPbQScQLBkNJuJzhm3MChvNlVrAjflLm7MsnMqsPXfsb3BiB3Jfjqmx1nEK4Cqqfs/WTvpzA0Dy
T10xjjk6NvxNVhiaXvYMq6b+JMvYFBZh+r/A3mgpFx7OVtTO2sQkGwFACZKVdwr7/QqXBJfZTa2W
bInHsCkN4fTlHa2wn1TG2WzbKEh4zO5zxlw9lw7nt4LiLLdTh1hyrFNrsuE2C8M3wxFsTDQYqfIx
DflFUP9W6VNPWjWS8he0Ka3CvEYPwu1AMzXl21RnJ9z8PNYxoXkCuEmAN0IjMUPu+RfzcsRAQZ8w
qD0mfWmv/Irrpz+lVPijlfiYRRR6WgRH6Un2rWTCGIlaNBt3FzWB5yaGSQ9TSxHAE7D9W3+QklAf
fSYKbainFnAZcAshQaIs74zns+7A1WnUOI+Z4AhJyIwo6yRJz0y6lTI4lwT76XbWxtdridmMJYcL
4RTL0jw+mqXNJGRei+rXbNipAD8U3dmTTc9suolaxYpedVmmavwVuwvqI5JWIlBAIPZelPTumtVo
cABkXqlbCT1k7QvifdmNrPZw7g73BhSsVmCmbhgkQQ0IUSMwkjzYKfbhbrsvZ0fTLTNqvJS4nLvN
yku+V/t6jrdFI4wTzUqcCmQmAjFy+n5HrAjngJwpWtUYKDm5hTdU+n9sN7Yw52opFEth++mxa7Fp
YiMNrHjmS5l5ldmDnQ0YwOQCVBrSamLlsrFPecoy9k2u/e9OEgfA0zEaS6rODCpeCgvxZD2Cat7P
1bngAPbKzlWCy7EMTvqBBp6fGQ+lpf6TqEvfXQRvw4H1rH1nQjFTyggqguLgUh+wlH09NVYOvHD4
9oT+XUxuuhg+cl4pYc+Mmq/BMLhVOOFblgOoUCU7Jd2HRE/9azWpH4fk18YrxceAGzTK8L8GwlPN
CMVGVKgXbLV7v9HaMF7se/k/NIARqS1i6NoG5QmpcBP5cypF+8enMIsizBG0HBrEPsUtCrumGJ2B
lPgq8dhU426y9fWAC6FKfTJexGIlCkax7Az3hqc5he82aZdos4iQ94mKGFCLgHjlMLYduAXbolzQ
7FJib3k9lt4wxIQAsbgYoRwLvxKDroIuoMQHJ0q1IJx1KBMkynLSwi+QdjjKmumOcI9bKznTyjgF
XlYcrRfvtcjtlnjJcE62FtGkE3NOn3MhXtuMmxaDZJdWzqwqrTlAWxHwxl/bo0S6Qc1PAvz90HWs
Zf2ueThEi8t9pjtCXVFrKYVkFUNgppqYTnsWDh/I+DIHRPr8KC+yiDd4vp4KVzv/YnpW1f7DGKKW
DBlNXCdx/FMu2i4+2xrLxShkpz30soFHz9kudapja/aCo4pM4RMdHKz+T2wyfbWoZvSZv2cOUlVw
a/X6D2KIq5fesvjoGHW+1mIQTh5urxzWUAPqhl4ed+CBn0AGb0I6QWp51Emt+xh/z1EQVr2ogQY/
w9QSMZUM3WgK+yzT8ZUNnw6gjnxw3Xtb8g/604jG7kFKG0K+t9WiITcR/wrriTHGFvna2jMmXWVX
1PMfhP+5DRYqHeEbV/qiooOoJyrRVBYb80K+JGtbesAguNC/f+q9WrJfOVOR4bcJimgG36EN8x2T
phUFBzZNQaXZJzmRLYZd0pwomt+cOTPoYJU18aAaMjZ7vd7UZkvOc1EArCSdhhrLRQ90PbhFMYej
cshUbe5knrKZ/Rd4/H2bcR7lKgsaXeWJW3nnBiGD1IeZw24pio+zG65vomH+kXvGru+Oit5iFJx3
hLt7StVA3BlblTYha7CksZyOt4p09ejHnVXKnWFLw2SBLBCfEedlN3h2MWV8YnlV/CL55F8ynM/8
p6Gm+25TBQPLAMMY5o+hvwixNAlokgTueyzIb8RzEWIngnS8eYk3kMA6nDwOrxTNFpKUOyK+psSA
7xoXap0mNqNyp7XRmVjBOE/KmK1ZFuGKMKIsoqZRTbrhLK+q8ZGpNgE9NFRvJD/dUerXIyZxxJYN
CWmERtWPNuGZmsVEATSAnLXVaekQhnilumkvxIb/kVcVm0JpiQDYpU0ymVqZNQRlBLNmW4hq3c1B
xLd2OR9c0V4p7ROR1Nsr9q4vZCZLEylVux1HHr3nL3KfFp9eP+7PScWoops/GlyKx96vr4PnwTjm
vHQXm6sgVXCPjt4dDiEXnI5AR4Y2DJr6ruk8lYYqfUI2QQBD6dvxkMXIloIEXMiX3btFMZq+Dj3z
/6mQ1XuRrJIu6uesmI5nLfYLrP6brtPb8KR58RttbngbCfHwH6HIbPk7SEaWIWR9rnIwfntjYiQE
CSoVRq0MB1WFP9TAWTwYoVvMpnaQmztsilGgZZma+kOlMIjYypEijThNuRR4H9GrEzw3+DsDD1Eq
WhW1f7QZwEYSleNtPc6bL0V/2rHFbSUCoMcmvKoY/d1+8SSKa3Q4Y81zvx70tlTyjMrn9niGDOdq
YKvXxf1JRjuH6goNvwfyS1ZKn6mKKP+i0nLk/GAUE4Lsd1dGVwmZlfiOH6wS8+NMegHOcn19PshF
RP3OFs78x/Nd5M1NE03/Tx86botZ3FL1pBKSBxRlfr1Prd6vlURd4ANiB1610Icum90DBjIQnvbe
9AdSZJ48yi0J7GAMy4hjlAleqK58vP4a0hEQ1n9VADjMw6Dg2qRnhD/9IAjSoghORdGeu637YbQF
1s8NKegcpAiffSstFeU4bb0lSQKlH+tEmTcmCivkzcMJIrYiWtJ4tB//ySejZoHht5OVInO4EMS6
yP6FeVbf3CP9tM5dPshKk6eDPTVhatlO/wRMT7BQvqLGw4MO/bV44fHpTuysOoQfjCttVy5EXKGB
84MKMz9TTen3Z6Jjs11WMHdHJnfRDq96xVi5I335RGDvB344qo6jw4y4gkQJQBVWnxZapcGgovTS
zT3hWVqEp2dm/2dcm1/IIlDIz8tQVdNeKeKfbYEyUIjilqLJZ+Bo1dUgelROuA40sbdnrBXiTkco
cm88eW8B7wp2MsY1J33Pq4YclrmZAbpmnfXemYTQy4Rwg+12/NzI/qHLl1Le8wB/X/HqLRxjQ4CZ
YGeGsFKgBrOsrYWM/yQ3Y1cylQfZy8SYxdJLCe84YMGb3OtfNqmsF+TqeNlztO6WFqQzv4yX8cpm
SjHofvWD0Wld3jPQ0UZBYzQymFmG++BNN1zRWP7uhWbZ138M4GKL/TyTpZbra7LEaCDY4GBaHdl+
R2mc30L1MStsVXNP8gisVS6rKvo261lRPmAEeHsl+J8g1fV31tth8qcBM9QCXCvo2OmY1rDp8cN7
58XaUtfCZQykQM/1QZjbSAapfz62MAmq5tSsNPB3cAqlhmnVHLyxRZSqwzFXj160S+0+XV4UW8yJ
ZbEuyi1x6x+uQMvFXRKL+bCds1CnNzl6BRautY0Yb4RWNsobwSnXRkcEJK2l7lxSs1dB31ph9MTO
9miEK7ViEXKAoclwoNeaq1y1j5AK4D3GM6/Q8HYq892OSS3HTFbHaJB6koGwtX7V97AATASs4Lwq
4JQMxK5RhTMVN7aZK9S1CTc+CwHHWyyjt3cvzAnOJ6W7aehvuwysuC4jIcyqL57yHvoFsFcNRDtm
NQ0wNtfUaa5mvb7o1uwjtdgi+FNSoNkeT48ikeVykAyKoDiYlUYEK481U9JrbK/4W2wbc3MASTXl
V+xoWoFelY10kVZJoOLkUQsDIUGyytvpwZIO3MR5HCU+qpydpwa1ZIhwP99KNNC2csnu3mqs/IKf
oYmxvm/dP0oANhJy0a7McVen5XfApqC9AmFK/pPe3MNbNDAggy7ujVL0WZm5y157hlAar5WZv/vr
vf5NYAsmlszLVpTcHTfZzXhN3JbjCK0nbbTBtQ+poiLdGJdZsQzzbUu0zStCb5WGyae9gF115c7V
mJdatsy7b4dmmVc+q9trpdRQaOQMMZ9yW24RRCEoMHUwIks3+VWw+2f6r2Wth9iRLUBEc6uUZ+Ty
YPtS4acS8HPhJZZRb/+2zFSpbge4Om06SAd7YI2KSk0dJOXNpMtFNG29rTWN+IgosifiTr0YXa06
DKJUlsjKpQuCLFyS25V0RLwi41KXbfKVWHz7Pu7mZY9Nlo++23xJRBfoD6ZXTy+BDbBs6qNklmu4
NBXpx1ppt0GBdOiodYmFj8X540jFGRCuEcImetxiyDSz2j8h1l6dAFmVzOJY9VfPDfH07qTB+hEj
PMbudsO5i0MCWuK+sWWeUbEOzEjll1UP00KlJOaoFUDitxH4mRt+xUIEu4aF40EJKQ6zev4233nc
QFwV/K02E6v0We+olLiWSyV16S+DImOXnKbMggaO6w+MiRXdVPB0ej+OeHG9i9mK/0CnJ4MSiXwU
sUBerewj0SZVBiB6Mj18R7N1a8XigQdYaMU1bK/BJmdRH3W1WIkN/loedAC0SHPTymC2plkyr269
0uD8/nOahNTNt/mwB4QWhNYNpw7ewYjrW+Rmy18dArBaTQuTjVGn3tAWNvGxyldUvvf1JxPIgNFC
2WPTUJIKUyMVzEBWrx99S5xL7CtooZXF5pmCcNeEhT/8677vCeoCxGmegi0WsDaLwc1zEP0mpBAk
cRoVPXAYFP3Kyp8H+Mx6xan6d76nB+IAsqwfVxbUlGkTXBvXcC3Clyc59GKEtnarT4SmCB8qkdxl
cj6rppnCQnbGAjNcRo+h0xw0R9JSU49jbRvgTQTtId7wNOeTwQOVhleRrFzFyOyehgXwagfw/DX7
OL6swW8qiwrcgrXQ12W05dBpY4ogdFgeZE/TU4dol+m4h/weYirYb0JB7j0PlwVMi4Bs2+IRdSz3
RY54gFAVdmIB8sqj+6p88c8AqnB9iveJB1vzNHt5isMsN2DEzYGAC0dDd11nuKJwnfhFvaNeWksn
RhiPOEIvuApynl2E+70YkDHNSwVqR94G9X9mnBN6KjeiYLgen7U1aUk46R/5IZkeOS0wdeMEvGA3
8RTypJ0N09yiiMc+zKEce+CXX35Gbx1TUvkT8n1WfckeZjBrHHFnGJe12S4g2BBXEJjD1YjbFkcq
yz1kZTp29IB019bNk7JgNo4xmzvLEH2duzFUOFnIZonAgyMznDbxC7ez6hhSOAby8Nox4e5R5mBL
TmPTYSYEPx+J96PhHguz2t36C6Vwl4qc0qH/mv+S+LcO4VdZm7IZNylOwU8Ml3+s2SeNdYCk0Hg3
8Sg9CbM0rqpBvKk6I7f7m/B7kadddfTtfnozv5ZB9NsrTOO4TcmKJKXHUMCK0zayAIAjFtBslevH
pCshNyajcmVIkhNZ8fRTDefqGSMGnKyqQaPCgtEehAPaCRxhNhhpIao/C3ctVeDnvFSmG1cTUNAx
hsHppYQmKEKGhcDav7SStY59qm5ZGrj4mIt8f8ky7i+kz1pgqz0gyTpIXd7yMTd8kfFwpXRLHJAG
dli0p48MkJlgKTyXbSCJV/9Uc/JHRGaEplt3yXvdUujJ//IIugz1DwR0EdG+K3Xpt1Ic5TehuuDg
vB51IifY31NH1XeSqDD5Efji1yDTKoyTZEi7g/cW7b1MqzwXJUtXQRLBG3vqIXgxkHHhaMygdPsG
5+qU5zwRE4BEDsMliJ0hg3xBlDAWsnW4Vbjfw7ej1iQEHY+NcoJ04fMti0AjXHJeR7nvYqliSaYn
Loeo+EqoTGl3K36Tpy1y8z0zt4pFMQwHBjzKMdzEx26w/bM5JmZkL1kvw76XqnOm7EI8Qwf12Rxq
dDkN8rEZu+0t3J7oFbDld+PIhJvA9+T3j+enuhnWLfiAyAe7ECGQ5ydAZe3uLQ9oh9dAq5AgQmRl
cwHu3diCTmmoug8vo5ez+V7tD/VGNMU+I5aC6I+sBElT5v/pn2xvqDt2uj68RtRxPpUG4ftOEXdY
2uXmDxNzq9LCJp8dC6I0Wy7sx4CiyMPm1TQrf/BiOEiODcln0TLJDqh+bPU2u4Yg58LHpeW7coCT
IRSaVERozPhJgdtuZzdXFvreeHdMHPhA2/gjSTVloXL+wYHgsdqGOzrRB6TDfAO/8m3Tf1jvIBOa
T0zA/mSk/Ef5vcQJ5rqLeknwFaTvUtT6hFkcAQW20UO3RSnxc8mgLRv1JKnVjyYJWHm7fMc+gE2Y
b5z+JIVy5tp1h0ht2clmfQULLx1ChMZcBiyF0Bfeabo23pK4sI1rcj/OVyxV9G9FzGW2PSAGs9Zp
WnoHtJ6U/ztmRJ0SV+04E8qS3ozmpkgJ+bSPyyFmyWRojMuP0g5AbuybWzRFNGJ+gdzyuqtax5r+
TKaHYY5xTaau9aj11A9BRvXBlYWEct5tyMlOEYC+hdWg2Xq4uaGTJk40CBbHqBDb08U2vQHSG7f3
WGDZaeVCGjQmjy2bWOLAvFrO7MfcD9NRVNDBiNTV7TeTEd7xdOcAuBmMjhhNH/4opR08zuyCrWJ9
6Z5GBYKZp/C9E2e9fkhyHgsUTNWAXDVtL9uQQF/0/rmQD76SFvmTqTz8nwSihNxTyCzYeEv5VS0e
8yYuSyy7U+N++dX3d57t4Ul4NYENrsOjUGTBuJJ3JHUVeLuuyBBzROgw6PcN6tVzRXRHQbpS+BLh
/wR3ee9+Yk3fslr1tnvz2RZBzGCodONRf1EHR2ENqqgBkvMBDgJH4/pKUoxcb7aWGCWLp4qFtcFV
h/aLbyFC45HDqmiCF7l7NJHYoYugKfBjwBvVwbxFL8MeQpLS7J/meDSVlytC3gePsI8WJF5jzKE/
GGdYILXz7n9a+VYQPAAYDzH29zwyJJGEFKRjxE8DL4vWx0zzSOkcHgaeH9bpX+8c5oBHcIP4VlMG
4QxSZEuYM0da/ULkXorIf4cn2exjeDexCtDlGd+RXSHywcYWMJUIlpjbMQO/+dc7DJp9iKJBNJyn
n7M+bhHjYfWYKBMXq54AdUfpMzKcQjd7tX2qjW+sCOgLQ+3ELuG4XlNaWuZbcsNBSGX9FS64C0Xs
YaWTFFf3uZAxB85vcYqwCIoyS0CPkH8m6yLzrJIqcGfqlkx6eRkkqltW5RSlT5WFZG0j6r+AEcg/
5md+wXw+l2IfI2q99eZWYMmJW6uOayuDg1hvgP0H97dTiB+mCH6A+1He1uHUEAO0bQ4OM2w8nbjz
cgY44fMF5/4x/X0etij8KHIEYpJc4a7ZQOi8kUyZimdE96oTfX65SsCuXMZn315gg5b764JvWY5X
dEo9Jnpf14oWbRVploGiDrsnb0B/OxTG/u8K5Hj6z3JheKKbs/iheT265t9XXrKvX4ELKGDux55Y
0twPcNYZGQV0KA8+XUk7lpUOUCI6GIoDhj6xX+DhIf8c5YpKP7QOLPSFzSI9G0sqgNZDFNFxOVDG
68duvls5Ti4aYqjXAltfrOMqOrsW8ArZ53/kxM/3LgEwDTDqhYx12skLDTJtYbLkPQ/9RalA0XHW
03K043ek1cfnfuzyiW7wOWHctt0wpH0l9Hwts7ip+jYpZJ55hyYF2TbBkLIAitIeyAATZzeP1tNi
mFv6gkjReL4/62E6pVuqkc5INLR4KS8aAtbencpvxNS9ShMIyEETKU+eyd3B90Ig5f7j7AGmO291
uOkkmeoLnTVjaRfvqrneaHbihUgYgK9KMGDPCbQNC+pPCWlGndb7SMgAh/k60VoYg6ycNXXtOEYy
jAyAAlpn0EfRzmzaMbT9omCgH1SULwsTNwrSceD2/jhh6hK463QCBNMugjXgaFLlGFFOrcKcUC3X
M559E5H84u2d88cHd/22Ek9U0TNniN8LKPjNsWcAT9n73BPWuuHW6KIblv28aIfcgkzsJJzgTmQ2
w/mGugmUjFBafSqnSjWv4yP+WTCnKddGe7Ikn+qfeulpf+62ll5uW8V53iInO7To3XzZ7pr28qqP
tAuyY2/qhsEoBGs1OPLKWIEok/5Bnbzlg93Q0MVnmGyGbKgfkfhz1E/4tcBdFsnzqifuEZyF9x0T
HAZUuID2uWCnj3GqNXIUOlowl0ENdJwM29eyL3Lc40vqpPhSOVVo1KPx8Qb05wNiSLkyKnwX5QW4
WHmUr51eqw8aypvVx7I2sTPi6fE0odxAEY3H/Bteyb1fZyl0IckJmWBAJtcqcC25IdiM4+J0+CNt
aY4zzzTop3fE6CPIyvMwKI3agUKFJOzFrTCWsnDWE2SXGNZ0RNJTFVO94mu44KTchmN9vZkrQV94
kKyhnMKfpXlJL9TqJq8uejtbmS5lXucbsqMNSI25ceE8dmEOj4tSz0RURc9IFmbkXDYNdgrtrBE9
28suCamukaaNmeQmJUu4XWYqjbwLI5Pp2NzL94MP4Ct4Gh7Sl/HSSBmKSX1mw71ZTydvd21jfg60
jk0NWlBqF9zvPJq0L0xxqGvzUyV0+fshOiwctsFrCo9TW/HPkGKApWEz6VJ5qvlbmc70rHJ+sEWP
6Agb9v8acNrJHMrvNZFGLbVX1IGXotR2fyCm2P2nVD5Mab4O02bZ0MQJLLzRk03OVwXhMv8x3ths
OamgVWxs6rxZQR1oTSJp38+KY4NJxHsHcK8fs0Kn+rJD51y1hBqIYdxsz2AtFQuAOeHmMrJJeQ7Q
8yJRB3w0PTBsmH9VFvl4TvlB7MA7B3YXbeNdhbZCzEte2OlJxN2vQ4q2tQutoy5vPaTDu9LqdGk6
exL9zq/eSs+PgmJhYSLP3vknI0TGFY17PO/KWWNSycqJIPQy3/TVKlATD1GiGQcRkRPvIc2U7L1+
b7mSWej+sLOW0vxaQr1tf+Hg9qRv5cd/Ej872efWL/dZ1SlBuETOc/J3cHIarm7QcJqSsvOPE0zQ
NTrpoyjDiyRj0mVUDBsdeJG1KoBVWkogLRVjtGStQl5ZECDFyaPziEq2lXc8g2V7GtoKyR3mtmzF
Y2gNA2//MZAJCKaI00NdkY2gHwXq3YdiigQPCydWt86mJRoUVXxAcnUray59OlW9bspyHbbF2v3R
aAicFuBLmR3T+xWGAaVzOOrw3eVZhQVD1AZrkr/y8NntHpfdmGReOt3anxKcGcEcGeYkjdMgpuiX
dKKad2E5eIRZYCO4Y0/EaA99j8pF0Lbx3nYHosZnRm6WVkvOw9CVbQx6RGIMvJ+jnYTRqCLyN0wE
WagR3gzESeWCxtUU5V74tBzyMPcpF5B9wZEziPyW5o0lSbkwIVtCSPF/Z4w8rs4bGpFKEaP0MzRO
+TgQv1Z8pnLbbVMJ1cxTTubh9esotdQkh8lhiSoMj3IFbyq2wG9DmcSEsBhlmICpu9nOyQ20tPIf
4ASI2x6VTUu7BdvIuKeGX8tJnUZSGIWwq7npqXPoo1V+id0EcoD7ci6ERgXA/BsZ3BQa9RIvQlzt
vdtrVg3AX9pGAElnMLNllL7YrKbW2QbqMeKD6MJZs3CrKdbpOrXsrgKh+zZqlJGKyCZkTacIOjqN
EKEdy9viV/sgt2B2DVwwurLOas4fU59cxm2r3cxu2r3i5rNASUV/lAWHeiJq7bJNJI6Hixj/gDWX
S82AOUrxucLrYvIgCnu3ghsEMQpwT5MzBcT1pQM3iFSMJj3QqVoWqyTWr4gInEpKFJNFPCtZgQ6r
FTKgZp/IlsuoUzchNyGbxRm9SY2fHkLI5mZf9lEZh7oa2DFxXvtjdnlHw5ahBO+ZFgadUEJq3y0r
14TJL5H6nSz75gEOZhrHua6EDe69nimk55ZSETIfgaQKqi3hwOc01ExxcLCeq7DY1gS2BXjRTGx4
30QOjp/7vaBqf4M2/h/AyExQkgRa2tOn98EE+iyCHIDsyHBl3R74lkqKir1fzLJpIjzh6XfzFI5k
CS5y4kFCXSYiQIY1HFTSJRLstpDvtyjD+pSNjrwTXhXF8Yx/eSgi2iPMs5XeEy7Yar6/4nDOijFD
arAtkblwmfbmmIjvyjtEqGGUasoAwNSaGp8NcAIqdd6vCr8MndgmdKfmju8WpeTrjSEtcI+AgYni
RMVKekwKdre8A7zpVAPYSuZAfR/9pupl/vAXFtvx4+XjBLAZVm7KDWzl3kQsP/Y8xv9irAQO0ILn
5IhI/QMLt07Uy0PeIyqxmQWU5sB3rMoJBvgQMZ8qV24sIJq9flLxxU+M+Tc/LMAQAuKInEQZn0EM
xSpRgCUpmXgkunV4j4aOOf3LgGgnX/NDDpC+rbpaVd/y0v9TXTcPtd78jLuygF1zYOvP7+5pvZhM
3GYV1W6WABSDE4RKg1YhpnB3fRyw59p2xQ5QC6UhWGASCZ7B8BtdkkRCdNSygF+OhfnA9/X1XLD7
ITkp4kLldz+37P/CDxhhHmOXZoji8YZuQsdZlaAwK0AR69tnSYf79xYqNQ3JbJ/vv5rHvFPKn48f
QKiH9SX1H1iC3FpnmyN9vF1ilwuRBJUkv+aU+oQ6CBXTXsqGmh4zQjwXMlpnlvgQJifO8n/Hbs6N
GvQ0y3Ykd84UFyq2NaFFV1rJSHTHZZjzQ1N+ABvJt6l0Tk8RualbqXb3StkxTOWAbxGvMIwYFIoS
rWrrQTYckZlcGj66ov9FAs3l8GMajaCNlrx/uR+w3ZM47cJLVXLtWwlHt1Vkukm3R8wCcpwG4Ot7
AARLLkPt+vZMeLjntm/gmqL/sIyaSsjWbYqSjA/YeI5pFKXQqjc6NxdFL8sc682j/hBP8x5T32J1
mmmPv9jrT/dRbzmeUJIzJh0Hl8eUG+ESxMzllQnFpGOWYpyn925WZvF8OepyucsmzImYNPabHhsb
D3Dw7McdKzLrOFwF/rLlbheNTPciWblKGNJ8HWVeJ8W3c4bHloaqZXqKNYE4G61PiGIpgdyqzf1z
XG0PskIYbr4FM7pIBhhditot0lYWR1kSVJwjI46pM2fH+50ZCPdSuuSJXDYiTo8UPG7uHGlA9BUI
IbUcNbduH0aindGN6UeK8NB0yYFLzmRIaPGbcLT2CnjW/b9W+Tsi+btbqJZonrvDIP7wsfyZwdWq
u/TtRpQDMTIK5IE4ESCh0uY7lpXkEd/B6cDoMnXazYrnRSuN/GD7bZrOdV5/kCn7mM9PEgKk38BP
4MCRI/6Mf214iwl9I1cW6CyA0qmUug0UNWWKbfnrGZdKQXCCN4ko9gL4OjV4/LR2Rw/B4uRpS16A
zQap5+MEhVlA3NZ9SyVt4h30QioesaqPzzg6yN1anm84NT56Ld996yODgcIsFsVrob/Z01feo6Ea
fKbpsyVcFHwKkbmxX8sL5j3QkV+oTh0GLypkM3JpGH70a4jp4/gq9z92DQaxeNzt2He9V5hR26Qp
Uj/4LQvwrHvHGsTPa9uZD0oUsb/cEdV97wOY+bGZraSa0CbHYskIiiaCNuMmB/ayuPhZ9yCMQ0Ot
PupO/ik42Df9agJXD8c/cswIN14KqT/xHE510I+1hG6gABk5Rsu6Wv8BHEle/oTnHO3ySunLS+gX
cXWQNuuHI/nVmy3bKsgP7lbunhfjnKqWVmKMzNzMJk7uDG2xpNx+4ad2oNPSstQWwdnLaH/ALaTD
38gtsQoZQPtSQFChoD0o9CmaSLIRB6dgeZhbXdSkpmmZJfzw+UjQ/HZ7gV5475C7EIovTw7phVbM
Q+5gkRmBq15KviKtyWHvQyO97JZ2ze504spBFGo6cRBHZETX9AOZcP/UUSbChyINj422Es9/sqsU
eqUKq/oKyO7wgUQsE/Ozjr0H/I5P1i6L86Zj7GMfXR1jnj8Y5jJ+3Q6QQO1sHrjRlJEAGdqasAMn
X6DCSZtoEdXx8uc0aFCLMM075rIecEHrABSH5cU7kXsGf0x83kNwlsD/Z4I2YHVlhyMK9w3lGcNh
IkOrKvSA8HgrkSNsPxhqlVINHmm9gp/V//eIjbmUiszbIWeVGD188bdsADOfCpALPjI3/g8G8BLW
RnMyPl9T4STXiF6DkZCkPmEIR9j/xINeANAT4GTc7yc06ILS+GueoHXQh+mbbwrgd33SWV46fbx/
lVyU7tmFheM2FyiloNO9fcQJd8Nj24wKimj8xQjttTah5x2J9F1qomG8fBpfQn81UmBFWVBLYDsn
sUGGP2cRAtQ1we2TgWFHGn474YhLu0Gmsu6IFyLwRZTmeqaVxrtkgAR/Tg7IDNBVlGMtzJt2XBVF
REYsnMKgWAzYXtQchCL66VSnpIaPxbj2Pl3TiEacrq4M4Tl0m66Q75Lpr9T5OKPVUojNtqh4zIlC
UME3aQey3AI8/lWHF4WTjmfH712lTUXlfpsegwlhyZbeaRa/Qr18BriAyMtphQ6FGASZ4jlhsnWm
t2yQTnN3svEeV80zm6p0iI64JwLMeNmwaoaOJdoR9z1z2iRguvuZyh6nx6OgZSbOo9CuKWvk1okk
oIqJvwDdpbfFCDytRFWbSNSXj0OEgTGd2yE0bOfhK2ZA/geabBfhnmAfe+0E9XUtb1rtlSwIQyCK
MMMxjZhqejNk/gQKEMx8hhSBP1ApGeEc4RUkg725tP/HU6vJM8VJItCgtlWjRT9viknM8kzjNS8b
C6Ag3R4jAlGA20MqCuZGtM2M33Tdl0j8Xx+JpwEitUpzZQeMF41PqioMfkOG56bsXEWTOYiWG+g1
E8wGQAv98wPiHKjpNYU/hetv0/r628yaF1M6I8xYcXElM5dH0qbzFXl392969W28VhpXpPq7SBbS
ORnkpbig+9T72xPT6cgufSEEOQcsKoOzANUZxYo57GH9o4JQadZ1APbUmpYShCjZ8RkhkGL6NErw
6ZFOt4zRiPCCbY2Nc0x3BZsOf/9zLnEaErGLWlNdWz7VigUmkanwe7cKbTh1mocbU7aBDPW50trL
O1g5+L6oyDyTZaPEur4WhZvgNBdBAR+TxMlDkgX9niNhTZn/N4ojXE4wjcDbcLf6Gdr/xXcCmfH4
dpFwe7/DuUCvmQdAoNJveTGW0BtPqyrJqZdmXrusAIq31jQR5uNPx+EPae+HWnWaJu9WU9teiCt6
GdhYnGABij/oSzANiJJA1Zv9GMJvakEEX4dZszeICJ4/xRRmceuP+LMLNs5yAILrZljuATqWd9+w
Uz6NuTZ8s8QVzm+hWRRCJh46waO+Rxtjk3aMHxF4a+bCIlRL9R/jBy6/V2psBd/3aCrJW777lcOL
/LI6cg7JWr6ny73ndNtmXrrKvEVro0S1Ao1LOKA5GWWO2YYPYRHoh+EDrIV7VIWyjZMP1Ilb54qy
+OXbXZ+ZxvUk+VG6nDgwJmpkmHkcIkloM0TMXLfu5ejMJiYR2vDl6V+/7AW1iaxpgn06gDN3B7DV
XU/oPeOlLKTMmxFofW57zgJ4dxGBQt/GFvN7UpzVff7yIdwi7XxD1FHUgSjl4WAg+j5qsc+iHJO2
bCGqeCI4D1h1aPTrsHf8nVFJR9lPBEzpdIMEM6Mqhm3a9XteV95RPLXNxYoxCBYxp/ssTH3XcLRL
XPSY5/fUWs1qEcBEsUvlQVh/0pdVmYr8NfaTjaDDHgLaxOc90v7btZZ729b7dv0bCspMMpgcXtOq
h2UL2/5pKSrnW+kB8/osr3ir/Em4JUkkBQyNWx7E1DA6m9MdVE/eRiVeFgGCyHBU65wN4pn4Ud1B
wd59nKAwHIl/a83wQRxvEais8AU92bcBwAc084mxCVn9mBH3Z49TkFxGFmb0M8yioTaIU+hg8tfM
Jt7VSz03JXrLDcMDI8GSR96LRJX57dgm/DKd1E3Q7q33lLCGy3UxK/hav3cSW/XuW/UgfptfoUXi
oBuDP2jGTr2f7/z/6cw1GgmXTtlptCVaAmsw5hZb9oXe+qeYWoKB2mrZK3kIGCq2e63kEqaRPhmw
SKRA3ucP+aJV/7UeTdVW9UenuTiz1SZSgc3wBLrfPYGlJ5K1pbML4iNTT1nm0ube+I0Kx8t/tMeB
vO7zHiI87wOsDL01+qOowgDIR/bXqEsEByGE4XjDhxLFr7D96E3hFSySfH8Q/DbkyTbEG86kW6mE
rMWX8ZM3FCqGuYOkNBKFgBUELjQmXR6k5S1KXDOjMtqeXvm01eBxAUDnlzPTSYA9W927b1lgM2M6
1/jy0YB3w7W18V2JCw+V6K/Ha590wnT7EXBpIsV9tAGGCd9MFcQABdDCdhm2VP4yFVKuLH+kk1VZ
5bb2btEkQTsIpTMZ16i2rhAlaiaAFxoB1u9lHw5MdpdAMtspHuxxAQF/8PSjqirmIM/whYYop1gy
HOwBL3PkEnyjWe9MXfLqMLX0S10gPDsFuOJXf/qtTv4tqKmLmCyB6/ULWVnT84bhEid6uUuCb+mt
VC3h1B131sHs/7onNu8afz9clGe6kVcpis8eGky8rpSdYk2BqNhPy6EIEpHrn+2znlPmkp3vf+JF
zWeixvWAHHY5KVcGsLN/bXnP0xY3V3c0MxZi9wdy3fitDNg5yoF3+SHrA8lUjLIQh3QTWrzZCMz3
x2vvgp+a3B79bHjoKZJBa27dkuVVdrI0IasJQYCol+U+VZmr+dd4dMSN1Mz4ZJwL0Dirwjiwif2w
Mx2yULuJgK6oOauC/ZE2JDQ3krnwqxcUzwlMwRR0N3E23V37wy1botoZq8Z6+BrgFUXsHwySVGAy
9gzVxBudmabHRPU7y9ulaCrFvp7fmmegxinNOBue9A3kq6KQyujHz3CrWv1HPRNuvCtoSJ65j2jd
TpjWP0Hegfm+Qlf4vfnaBLoQr9Qh45TmQ8I892BYfmQpYYVuJW+q9g8Wa3T4UIglXcJ8GqBFRuHy
YzOznPJTHcpc0GJOqffTJ/Xk+ytlKaUYIhrBBv8pcLfEfrV9HH7aQgLZjEqBvB7HPpVoi12DwyFq
kGCcqg+1E4wVGgUqoNUj80htYbjVXFoiHXMm6c7pBqwSEpWGTPVITm4iRkPhe+EV9Ze4x3TVEUxj
PelNgt+YphHFQAFKM2Dcy9KClWApov160Cf36NwhuWSN/nOW7Of2Vzr1/jItFDk0EAL8QEcOCiw4
YE34irtVzN/jPJwGWAIgmXxcSKml0Mv7netsEVxMFY60ag+1E7yxJiRKQgHaSBKD1RTv6X3Yi1gR
LTO8pRiX/TGAqbCe07Q+TRtgG5uEVPewCwAQ5aS2oYIf8okKn5eXo6n+2z3+TS5BILt1mq49uSQu
QKh8gQJZQ3dGQSh6PCwih745KZT7ye+36YkqoyrzzGgT6SW1m3bq+rz0dTAlTNTmIIYRQlGYLpHN
c3ERdDcANmx2brrPl1ZNwYYn0G6Zn6ReRHZ1HbSFHm4EC7o5sIgKf5XPR6s6in9FFauD/NljJM+/
OqQleSMLIMLwyeqMY8v4TFGxGn/7Tp2VzI36/mumh7Ec8W15SYKqpLEia+R1Z/zu3agdDY+Rr6Ab
xAjsq1w1FvlY4yFVOoMvfKgHKGepSEDNg5El9AymwD7y0lbgcBv5/uBm+2YFTzBA1H4L22XdQqgl
freflbYkOO4TRh4QpCoApZqx0fiLKgX1JXvRBLlGKSVn+Wdu+KnTrLP+8zf7FgFhABsBFp9nv/Ny
jpiZJy0sIu+8Db7D4+IQfVg9wTb4BQes6Ze0tB5FqqiK7vhuYGBUHW1wAot328sMCWo8wZeyVwpi
0C3ItNnsRi73dmuL/CMcdSITeOlcS2aWPiIPvbX3c938AVoY8luscwwSbMbQmSuyYiAlYWMuhMXC
uz6Yf7X/Ib8O5d66tg0UfOkATYVA2mSabKnjSveaXFSLUHFJ9f7vh569IpB9C2+2kYpmgd8ABWLd
ZKQIiIBpl224j71aPEGP3cmUgG/BXKNYnFDTHmIVZ913/xdCv3p7SLda6qMmRmUoIBbPtrI+Snqs
oajdfuEo3XMiFXkEJEiWVSk4D8aHuuk2HEwo+Ke6+cprrldzegzsvEMB1oIpUUXCtl83GRqlzKpg
n8IeXrsHcpWC4f7VxtfX3szi1xxFpKNQnrki9+hTZtLWwdJzy3LXrH1oZALd13HsER5QFygA/qd2
iWefmJQnUoUFIw0zEGEjxZeysF4ptfLcBpQNg4LWC/rMhqpxPl/nTp0T6WNzWws9BRPF+qRvUexO
j/hX5ZT2AjuPg11azsQP0AqwGbWNlykRJrb7CaBEioz1hRXDngHfyAj3a3zqOpZkOSgO254dphya
pNWYhIR55yCOYYGcizE6OKZY+4sQ1VxeyjazuiKP9tcrxpHxc7TYOXo+g9UDpgvdUgW6zW/4X4Vy
9YA3+WPRPB0yAC6mPKVFNtQYOA2Qxlj5lF0Dhjk+syFWBf/kMwYbOYOw9MHPOZCkTRf6HLGjpVrC
M2JbnipEiWsBfJ630S9kn/HNFJpHJhJ1Zb/gHlFOaWPftHB4R6P54BHOm9hTdzbndP9Loj0wsL1+
GY0uyFoHBCizFMeiqUcO/Ob4MJAqWBMKVW21y5+s5LB0zy3IvpDpJol95atkbSTvGFJnb5/VntLr
+4rE/enL1MSRtZgqCvuLi7m/pu5Yh2DyxvuCqQgKWdus1ZVTSAVtvOQgl5OzYX31w7e11QG03kn8
h/En/q2DivakZZ/N9wDf8FXPTTB944AbXofZ4ffEo5/PayBnVRNl6h/WpREYz4aapbFUDq9Sd7W5
QHo1i2aqnI1eoX0fZMZnG7+TYn3cOo25JfudpU4yrlnrgRzv2ApL1KW0WEtqet/x5mraoY7jN6Pi
KlbfzoH288C4BlAOoKgPc5n/Q+U5CQqArsZ0ICoNi8BHt8Riz0pUtseF/imBY8HApQW1PhGIFcHI
As0csV0Nq4icoRnPq2ZRKUN1I4j2i72/zLPtoemYc7IcGg88b/VC265Pgk8itqMfJDH8p91/7gu9
WqCSOHzUJpaf2BlWhiWQ1bWpx3LyhNU+2bnWr5BaHSFnkwzkAilq0KZ4EfMneXax75K2ExIPNzW3
olpxBqVABleg/pVy25bjzSaqbISftoxmkMOr/9ijqsRsv4W1o3eBopov490urm7zdVTcrBjTVNWq
zS6BV41t/R+GLIjZSAFv5fBDiOD0Z9GWDoqndwQG6MvDztObIEqWCztR5Q7zjjGa2OxDsO43lFMH
gEB92RfRGGjI1Ul1DxRwwM6zWNfQ1ay3HPdpbn0KL9CSxcXBCKxvJB0n138UEGZuqqVmBIyLGHfP
4ET0kz3uxyjYL5385Msgm8ovVSfWRp/JiHiBLtk2Sbiott00V0+mL/OS6jTuxwXImsGa55g/zOnw
iSGe1hD3jCR4FB8MKPSrNvO9ChTW60YviIDySqOXs8F1O/TmRSko6J1Mo8UNjDxMnKAaf8nlyosi
0kPGdHbQcjIkeBOy/6mtEv3oeCg/umLIO0j9lEnwbBazV8E2V9GK/Twtz3DYXtY44xYjCyA86lAj
LpNumXZT9xPYKujGfLoLJVtFzxEKcZBn77ProuJq/IN+6eS+igHON0Vf4p1//CvjI/qJSQ+nLFB4
jciYAW4LY9gzQhoW7gOYL3mOmloMpfknc2ZiWZtanNWx+SEFmQ7hDN0bIz7ZqfSOI2u4dVScG6mB
drtMaJn5F8pxKY5vVUKur6DHGDgToWEqXriXbqrfcQZAbw8+w1yZLDvwDELWrFI0tyq4PvcW76jc
eulakNVs4FhS0OhI7RRefGX4Oq80wdZJ8pUjBySTXBa+D5uuC3bU+WEg1P2PLr99uBfZgL/fjw45
YYy9yayLmzRAtU7eMUPZSPlKTMOHLpDgN+grP30IGgXLh+aZTFoeD9OS1k1ErmVbgmU+OdyXEHCG
L2kdUohzkkXsDU7mfNWCh8hEV/Q/NjbDXw+IIoG3J34D774POJ35p0Q68w6J5Pp6QetfDVSVkYoE
PWhMBVPyNXe650ueYG3ulfxPh3SWLwFcyybXYSMHkGf6aBBK0HxTnzZN1J+W4JB112ndVmFlctsz
ViB4ADqUNuTuLplVkSrG9RcWaOpZXaUPYYYPwBf73kwxYudSazoZjBxGToaxhu2RXP4UnXy5/TTW
eKmyILSW4YoGYHXdnWXilkrTyqceX9HzxFrBi6xWertpV4gMCAWbpSiPG7fyQK8KWoSE9CfE2PZh
WfEBGW+oz443DQmoRR0O54lZ8IMsIboW1jTybr+RH/I2dr59itzlzCLIBn6QFUSHGa7Za9a065ru
xXVcAG7dKWkU9HkAnw6k+AMNHRJH8WfvMAIxlIgOS4VicY5jx3oJjyYon77YQjjJ7h2Yr3JxUhkm
mcJyYfAMOCwg9SfaY3SpESerIZLBhXVGlosHc9zAbClVtlQ1Cv4eX3LjTEEU5AUAJOkYsNnfmrgR
VojNkjAHqEVYMFo0w/3jf9QLvrVvWXcAcWWE0OCp9PrbhklmpNME+WBitWKrJ7gvaaDs93U34cY9
nLSa0De6sABj/TqnuBb4i+9mvgXuuDsGSRVsySE28rznbh9Ux/hQb5goZhhAaddV4aRM3UME8JVP
n+PH13uvakYfgBnl2gpUgyxBeMkHZOHJpY7dB3ZnEFMEffYI2qmlsM4KoWHt1ndCqvRFdnyI9hms
8zG1xHBQbz+jUUCLtOOrpmh6hQeHG71HCZ5GVn8XSL2LSuZ0RUz/OLbYgy18vQrgE6+DoV3aDAZY
fNdgt2pvoAVOlJt6JgyWnDguUjLXt1Pv4cDh4EuVcNTgXRb/RpGWp/m1wL0GjSimmH9AiOaAz5VG
SYwgacTbXEr8UwyXPX8xO5HDqnbN2HVqZLC0+DrBZbjavURkzaJ9bxqb2/1NNZjXtX1Xhv907Sx7
CcrDAcNGiSFtWe8Td/V0K1nCIb6qWzBz4SksDLQrAJKHsa7F2gksp2JJuRX+fYACJ+XfhKnufIxi
SVyP3yX0DTrzlW8rhow3tKim++mfFaHc8STx0txZ0QDv7/X+qtkYbw9hSjl+j5nGY0Fp48pApLMW
vZt6oKjaCGCoc7b+PkT/dCluGD50grWgaBRfiaQJdHkYnWY5Z5y+begsc/D0MkQW/5vdeAxAHEuK
8E16uPObs7Hrs+WskEd6CuMrG7o2Ap8wLgGAQBLA/REaHw+kSOpDxqYNEp4gZyqKPqCvMkPMFycZ
8Xu6KJR/Dq5nyuoe+i9mGN4HYnkoWyFq9sGQS/Z/XzlCDJ7mmV9RJYrjwh9x1/YcBLbvCPkDifHs
dIH2FKa9Wl4beYeVsSTs39ipERwuYFtg7QTiSVSWAeCzggvsJj+pAwb+HmdLtyKr9GSo22I0iJ4y
iVlDTxlB4bH3a/03o9EsZJlfr3S3NA0Fhp5bYATG27Q036V4dbD2g5NR18fZ/JufTwgQu1rXt77m
AUpDhVayyQgazar8VeQIlnxc9o8EdF4wJZB/yRA1nHih+r3By/z7TPyR6Cyl49Lt7qN8e/NTOCT2
+6MoQCav+mNp33Zj0SwQlvF16uPa0s1ftkvDCS6A4htolPvaKIsdSfVLbplbfIVHBrCnymUDqIvY
ANFTMSGQiYRloO2xZBCabOVW5Sy0NW4cCZkD/aosf3XBPQ/7NaAFr5CLg45g/l2db6lgIeg15d52
tAflrLnDHsiJ2WhRQdnjGj0A7LWpVuWeWQ5KhaWZHGPjW1uwFtYLydJ22PmP7i36KyUERX9O8hD4
iikeO5hDT7CP+j3dCOEAXWFXmIZo4SoE7gK0jye9Q6IHiu3CHZmfI6yxQQ3W29nBj5m5cjv7tW/I
4moRPyrDDB5ERfGz6F2WRFKJe8otLv1hCUGcemW7OFd727XyA1brjDSo5MrVMI3yyG+J31jubPwp
/fqDSrIAgtXK7RIYVQVU3SM7WRV7rxDxrkpYs9f7zkgLeCq6Pbybokzh8dB2pcx2JlvLmeiG2Uko
cdCfbg4LI4AwgLAUXvWot1D6c9zTlZ7/bNgJi0DQlwtGVKZ5cbhPeAYK4fuXXmXdGZm2G+Xux6Z0
z8E0MaYG89dvkzGP2/vXOM5S3W+hAEkkh73JROnIVaaII/Y69zbqK59YH2lw+6YkIagA0ddbNH1X
qIyvLDi15rZxei8vLSYxDQ/YiQPr2/snJ76if+z0jYrCEM9kGhm0eII6Q4EhRuGXeTJW3WHaTna3
IllLRLG00f2pi5OyYgH8u8EAJgiA3Cxn9NOPMnnzWIqYDksxYHTIrHTQud2TbwnhUYwOwr52zkU3
rKDsDhq4ShXRkqbfuzAWF9g14cdr13vdHLlNMWuQxSHxmm83fLvBcMH3L7RJKu9BryF2DcaxXlnI
AGy1EqPivXQjFP2AhgQ7a3zyBXN9FcoMtTL+CG1WdAJOvjaCI12NHYHe9Hunf2we9GjEf9+tKoRi
OHvLtcP+LwTBNj5guiQ2Wu25OMm22BxBZf7AT3grrCr8wUprWHgBdpE/ljIQNnbijw2Ap8phQoKw
cLkKVuQl1J6gKIQdWuPwnaz3rN42/ODoip6Bu+oU6aL7ihl1UDhWBvBGUQ3sJxdmP+LlUnMenVAY
9nsfwKRvarJhphQFpHBguv40jgzZM9s1u/kJn2J88KBECkxWmn/nCCiSYozd+ieIPwcH4QvFBmN5
bpIJ0jIoivxjZ3nqG6Zus0yOrmwYgNoNpUPeEASlQSYhBBIBd2hIs7XVw1XKcayCL77zdSj18zFX
gpAZ+uK5J3cesT8qTUEQwuksLh0l75S9PLswFIJVCZf2lGShhFm1RDVN2jOwgL7yZDS5seBwK9tK
ixHu7lfaGhuo9+YgmefdXkj9i0Nez0fMhcu4RozXLhudyI4fDEpstdPGjrTNkHWIWTCFND+dU9Fx
8wiNpUpzclorLD2+uJMkEdwShgBxeED7pI8Pq8ZM44WlSxSsssjx3MeGohBaaG4nDMoMPu2I8QCP
6izgfaPGloRM7cAMApz/DuEqKW/hyghEjqEOxt3vbBOyCOthEnlsslnC6SeJkRO+Oka69fPj0H2L
6NY1j+LfkLbZZ0hk5pv7+JxfScTtQqR1a3vMXDKBnuqfxiHJHBR3ZSmGOC8BSzpZmuiXEaetFYDH
GKQzO+7f5vNdPWj8tJs+iBzWlU12p4Y0FNUe2tYicyYo0sFk8PgnnpBeqbJ5xCAlsvY5IzcpJKWO
5wCnh3ajFVuNZaEbKO7SxeHyezm8QK0kj4Qp+xpe/1+vqmag4Ln4rvZWlxD8LNkQi2oHru9Hm0Q5
ff0YzCxYzynsBZeIg9XWY1zbSQivrQRjMFNhqPgboOeNxdoBeUZeBK5+Dn0idDjRfMKV54G6Mq5P
diEb9KuQ28boHLidmJzQBpJMlSu8vBaKlE7QArzhm6rEyh84uRmIFT3ih5Z7Je1xhRSEJZ0B+9Ro
R9/V05/uApSQf2PKgo8gqrTjQNT4pEoWEBW6LNAQ8tgJ2xUKotqXNR6IaSHlW9wAniUmoxDzFMJt
wrAzQHHVM/Cbxjn9F5laDWsz5w4F1Ufv1KvpEisVbD21NHZFsdTv11n1eASkX0M20WCM9NZzctkZ
j4h4BrYFjdK3yqKdwHS1FIXNFWp4cdCe6aJN3Y7AZyPu1d8zov92BiVlVD5b6csblE5bPnWb91y4
tgXaPcY987DNQ0C4Tkzf9cfG+3BV9Ntl1YjKPH38WAiUWJEbmA8zOouoRBOmkIVe1ymYBU4/Zr2v
NDq7Xx2kRRuEinCuLllaA02pwGHw3BsZP/VcN4nK2OxYAZ8NlL6gd2Nc1+hpz8dcEgMYjufY6Y6H
NX7CpBpzSsmi8z31hXUqa5dXS0O0Ddyt+0VF9gLIhjfZgA9BUl5B1ZR7oZ1UFAr9BQk9fDwDrDv8
sgFoneBuzTZoyfHRkc17G8FltnRF006qY1zkoolB2EeUvIuNONnyolRTfmSwzlNOLBrwP6VH7dEu
YimFJKnlBZQVzE9k93apL41zULcUa0fLzMU/TlSaF1hY3lWaD2kh8JHIMQ2LHRWdhkleAviHP74l
nGPviRbZqsXFzoJOVD1nRcqecxFTczs7AVIVtZnBfnIRvbI/VnrxKgx6oEKsD6uy9B6tvWQd36oy
bTegBQCl1k1a9SY/hmOewk+r2E5oL/XyKGXfZZ51T76V8u9rNUbqhoPhtuKgIt+dNqB+br8gLhlQ
km/77s2YByYOxUogxE/9iQ8ScpBa75F7CsMKhsXpYAZd8V7wePAiVaBavon86XpDya4bB5bxT+Qc
kwL2IA3aqb77YDaEXgv8QcEcLdnQxzHLKP5a5NJvkk912lm5lkRclNOLXOCKpx1lfLjNFZlSnFnc
AcLiUOMrpeKmutqW/6rpNLreqNtxxQ6uF4f9YHEUtQn3S9rKwZciTA+2K/Cl/LnqrLxOdDHah3jm
SnxpMqvUJmb7kedsAEz/eCoNtcd8nSs7p1UhUPUyBc7Foj2JWrhAA6h93UfosVIEEM3BO3KJbuGB
ksOzICkP6VJzL8ELCTqs3ErkScS4nXVOTkdek8Y24mc1bP4/wo69V2BqVGAmdY4+sSzxZSaKPsOT
5OjxJADcJAJLUjlsyMWwGoLSjRtoeS/atOfI7rw8sIhUWOpZ+esDFaB38zjAS3t9vHqXVpaUPjzY
JKvTjODn3d3VVUMaYrJaz0oj7eEIlggtW1tHrd/PpFvBcfEqMvSLeeU+LpZDHc8G6J/4HiP4ieX4
rtpjeZ5dxqn14NvGXoPIWe8qny2wnCBlcqZNpd5qbyfUAmXDcYWhatlTa4Efj6V9uv5uGtHbtB/V
K6qxQTxtQCEThEijifFvCVuurZT2n7JAomgrtYrkmVys4yFa0i2XFgXhe/O1V/8TqNGrINvqGU/G
3+QI4ypEVLMGwWikbJPesdEqcy9VZvWij6iigYfCLHz8Ir3iGQrhcY4HaX0pivWnwRc9DJE5OzZt
L6Z8lS2ySlDShKuQRLS8URyQhRC86MV1++jg0DXCuLw3T6xdKlAh/J5dWzlzS+noAMN8jlih3dVH
3t3Lrof3ZIV93qcI2AchKTBjAejMPvTCqvx/RHsvcWQoZX4BDkhrF+vIaOLrsyXlR52nG2WYyJ9k
YdRg5YhCNlTTdR4iI37kosUoRaeEDGarDCzSmXLuGMubmcU7x8DiIIYBWkx+uRbWoS4cwwsRWx9P
c9oYOvmcoNFVoegFtiMky5y/hGxlpkYHYg0gz/FsD+YehDjIfcQ76kD8SdX2w5p5o5AlzVRr/oHs
HDnyD5kgRUbJYYVSM+C5b/b8Fvyi1ydQ2J1CE7Yf5H/Ana5dYtOXahmS6UnYQtlQl2FzsuYJz858
m/1eGB/yAxrmb+Z75EIet8MiDs4e7dnx1MzC8Ss9PMK9EKB7p+IvnrNw44rvrl1ACJ/w6s6hUCC+
sLg5vug3hrG5j8DpBBPS8Gr22z8+/byYR1kddCdA5C5Rt6vzs5F4KXsp41Sg2v8AAKMmiJmDhBah
xnGhVafLfXHLj5cl7pSjfJeUQ3h2RmRdWRCR+fF1Vc0EZM2s0LkpI4WwyZjoSdxSqqIT8nA/K9ye
OzWKgSqvSamEK5E5Aog9wbwxara9C2yydbqgb8TIP0L/G3PUOgE/cyeZMwahGKVSKCEusGtmCkb/
2yzoKCzIvBGlhjDTtTgx3S6POnEpPnOZNPOyTV8sloIbJEe/3fPSt1HevZZe6zkgbX9RKKPrhPj4
Q+E5ITd9a/HlUarVuK1Eb7tri9w26nfoQWzNDxtBNBGspkkT9OJMRe0p5FzMtBpz9VOelID9wcr9
DG6agAxz+jsE5V5++bijML3YcaVxElzVneT67kZWJCuRHoBG1goZYscCsv/jZl5KS2J6ADtujl14
rxAzOJix4CNaIrmas18BtQX0qkn+VqhveBQpXxXoD3NUyqBKOS85miXOMQmYUyIjN7iaVtrLSxoV
+4ScB8EZ349kWMSSH/xNQixjn8IBVPSmydcapFPOLCccurLoBdwRWZxyb8RxXyTwwkj6N+uC22V+
IK4YMnEgBzK/skr12B0p//e5znlX90sdaVmF6epiCwQ+RTkhEkoBNhXYTSOH9bk5BUdON9zzMXKR
Rhht/77wOOOohXHudzOP9aoQ80ABdQqePeg/wGYtafYgU38LR+sOlPQZ2w8T+dzTAllbZ5w1HDR4
jeN3Ut58rfGAqdLImmwxFEcLasiFoGU05wwKPFTl0ZRVXn7I9tTIStEFMlceAjWtzHr7mcdM99ld
IPTbirBQznuwwbKFy4m88XqSBf4Rb0pDybJAavySjfPC3r+FawJYq/wOOgffQ3+/SntoJ9N+8ViI
pS7gVFSdkyfOlY3OWE+45R1FcXl4BuNus8J4UEubPUNX5pW5u1dOV8kY/P9FUY/SA3CXaxV3VUh0
61CtgF5DtkTQkhQLyTup2/po63RpTUk7Mxn2ir9l7ZfmZmYKu9bb0rinSKzDp3hEvvAacjtKpBop
5YdioJYY5YC75wHj4Zoao8567Wl/cvBNuN5AD3w8jORQF+K1Rdd3fd7oV9VVJnKWA9MOl0k1/+ag
W36I50HCjOSptGSfCSoOpU8X+BLrdBevIl0xKThtQOFfKuigkzUjIxTykflJDNb4zcyp8Z+Yt5gO
6z6EfQ079J6TTzzObjJhN0AUJzcLTqXPmuR7SXzU0+T0E1Ic1IDjsXKY18A9ozEwHrDD2P0rAgNL
PXs02qv7AFT4TEx2Do/XOf3SlA/6EK7SzFdieeHNcJUTIUQrznVOSLOssl84f+Z9JUw8hbAWSm4E
086NBkMHVhkpTo0oh4+wBfBWZxurSW9c3TsQ0m56TPXGe4OPspAl3f5bUU+Yv5ehSf1YVIYMBBzo
5may1BcXiip6SEyTxU6qPNwqo/N3CUU8nNz72fxWkH779UzCh7h+ceXoxFY6DmGkF55xYGI5I+nL
PwR9O03YfiUTkJkV6NQhYkXJEXq6yFAxjkuHzd9DActr15pv9hKKFr2m4Te2O8OPT3C9a9FCleFL
VsGdBoVewfWFOb7rrMedIVSrOGLKXwj9pSoYFv8CSlNT8v0jHH/y5zFHhEYC5xsYdLLTy36NB7ZZ
pu07y91QxUQCKQ2a6o1y+gNTgVWt3yoISpUGRELMyguhmFQf5mkdObZon5EzsISOZV5mesrl+lkb
xnueoPE0HzL7Vl4UPbgvvMl1O79WGVq5movg0D+f20/JntI9ilr9wlfUewAnb4EzQU/LAj3G5B2H
+z99PJ53Re1nG8kIg/afOKclZbLZttJMLwK2elGyWpx2YHUwYPaWIl9iuOU3NmbyFp13R3/RegVn
z38JbaEyH7A+TYKZ+vjLyLTnOWkZpICA2RRsFYOgOEr0N9KNCu4axjNDjt2tWe1DhGiddnVPolYQ
79L0xo8hSy1eH1bT6FdgVgUco0uC0Ms/hAcwrEIrRq/jZHebnu9WAyO07ZnZiivaWwcCFF9I8+UI
NrRUS9cUyHwvgkWeKxeA3R+/p+uaOyT6aL7ht0T3fGGI5JIWqUXiOSo3genj9LTFQuze3EqlpV1a
6IjvKn1FggkpaMw3SAc1MhREiEuiQ3o7IePrxD0mp5bQXtWfg4Ga/KbHhZk5yhE7orPIKSR2r48E
X9KFKwWRJjn0SBPA0GPlcNTdT3vfWZFM3kh0MXAZVVJNtccHZbpzmnVT1uXNMicR2VpBcgCXJ/DO
BtD2CK7JKWgeUqcE9sB8kLfa/8pvf6fnMqI0nlyQgg9IT868qvuFZa0B9xqY66PctKlHcT4OyzUl
7ItCv5JO8BnOommvsLsxEdYd+92WDJ+irze/DrwvRFpdu77291PiO6rj2CcQLxxvFbvDwT7t43cD
S481dOiK4rlzBmZAkaYEy2O1FXfd3lSlcKYzHn05iCY8AwNRCbsqf0g6+E45Et5dkX6NI6Rf0LD9
oUj5JojpiuHa9Lvr8Hnw1bewLMrTF5lw3qigjkoc9tVBjsaTXD+Ci/A1sxDcOt6nKcVPZqtSU0Ln
qnKDiOkwv4BT1yIhNJGboMTyi8/GuyfJB5nHQB4zuScIexHvnxjgkrTpp/d8T3jgeo0hy/mhikOE
5Q+11jr1+SJTmQrIKeFiUfft/z0rR3EIzBrdO/8pT+yDmhjhLiQkBXwyD6sMkZ8TBxP00C7XMTti
S7Mj0mY2VHl282qUKzccyKWdgIcBK7ImiASneSAx6H5E4ANaJ+9SwHkpGPyx8lyCdYVsFbaKAw72
XwZxhYJMcgWdMiPAEz6pdcddaprRUClz+ZfQHR2lae7mFMMfVjGPLMuXP+7eNRMZ0W0owwc7tfkd
MmGrq/iOQIWgr1h9TGoh+4lHKqg6lUobMSHdPBaigm6XPMc2o5ZIaTLGxxHv0r8pez9NT6yCUOs7
HmSlGg3hdNclyF4el/a0MsvGejWjESx31gyzjwxcLHRBdjeYrZYqx3WDHRy1kPMsdK94r2GYhjjn
qsgnbUJssVp5JXijLoD1GoyljlgG72S1KxvHxAI5nZW64v/WtwwwAphZaZHVWx9fe0GwSdOqC0or
or8318HhUKeavCWRLNcMiCHXtKa1k19eztGxPwVKf8lsjuogDG04Pa/OxRzTo5Aa9hcatTJCaQuk
SfZrsKaD/LnEGdLNbXpKzWhJwG9IaX0fcfJx+MBTW7zxjuO+1L3V2zI66Wnj2WAjgGKo3NzUkQkD
zviNj6FRZg67g57fQ0NqXjrev7M5++kftVkQWCUqkqXb2Hta7zX2U6rEvbZHMS5YyPWntSZ/tcE/
LO4X+NqWPXVl2XLhBaYZXzWxO5kaINKrYXKpWuA6tnXO+dri1sVBNl5p4dPuv8siv6hMmdERKIoS
1wwLFA/uImnn2zkW4P5VKq+b3pbissLBTpaTQYnadhMCWkLDJwb4n/Zf/gYsROnWowXaMnDSUOH6
OiOtM1N5ZukLp+bWttrOlSCjD+AS/6CYgn3IpbtOaJ/lBL4x5eW2EFjLopxvq14uMAu6dJZsBYcS
mzLCOBMqCm79c3UhuOw964cmzUE833uu7zVTJC6oBTAYmhCRnj/vxwOMug7qvKw1OC0peNMcfeIN
TYVuAigYENCoh+8UtB7qO9CAGozlD0/UQ3zrgfo2y6XmgGSuXhALsnLiJjb3KIHDPpAsgyUGaWE9
333bdmDlRJurh4AomNtWJNNDN2+A+f80/yIYsIMLshet0EVZnYM60iaVjPmWP5T2Utd7XtYSJvm+
hz1xQCvYCoOOqgxnN6b+2fSgeRdcOSWxw4De8tzDRsBdhO4N+SVQe9FzaRk8AgcZr7VR/aTuwjOH
LN82JuJHg0Lh3gyxolaHMEfsALQMGVK2nkZNki2/qTes+qDTQjipBe/rRgmJFG4bo0VCv0cu0Ocv
Gf8ukohM/ehXDhOB6El1V9OVFTZRNdq7wNMcO3Wu5qrAjezQqZuUav72MAMdXPZcsOeTVn/HOgPv
TYMp53398GwCIILuombvsmdc2Zt+w6oNZouCaySGHlGz6D0MRxxq8L255032Vi5AHY7clH+xWFFp
XAyGwQ7eu4kONdbE2RXxMq1fUWd4+L/wF7vQTC0Q0yoJgQxz21BMIS1sDa1G6ylYLCixBfz6xhK9
GYoL+nMAaoFE0YXqHuIPbP7v/0ZGCSfLOx3lBHYFTIt8QbQOXFDdMsEvtHEf/CMjW3OhJpJ0I+d3
5RYTvC1MbNwNzC1pP/o+7NrEns1UJ8TfvSVpMwoXGHqNNgd670Ajmnu+z+WAAhQ7MXqZZUKC+2WY
QJCwzVVdUqwGMTVYd7wXX7V03NItmnAlSFQMlU5k+cBe624GW15UhUahST/vdqgpZihTv3w4tMyL
0BLZCrPKFgC9EfTAg3HZQiGv5CIm7RzOZ0MoXjHmBgWJFGafhAZMsVJXxN5V//PDiv/g5TJ+7CFZ
UHlW0KMLpmrAEHbDyOpVCUAGmAXlWp/qOkYcuM3VSQHO1HLxW79qk0JZDgzKcWQdYcRbLQNJvXlx
09wAx19/W7NYqD3MxuPHIYJ9IBSGfKjUzIR5SW3n6rFim/2gXlOdugUwcb9IqWABw6eQ7bWRBelX
Dnameczntq6SRynGqUp2cxV3Ali7w4xNI06EQMH2OsfZXwvLOgtHCGQyy4XQ7tv4h3sZNpOVBe9M
Z4baYhEDrWgfMBTMjw5lGZAo42xlczDrttIhAfB0cELKjZvJuh3yKRe8h/evbUP8gnzX7C8hadOD
AefRish/JK6gqvh3mmUSxlI65hTqc7p0Wz+Cd5m0/y9EdBMVgUSOcGSQv6CvHEYRQ5Uk1+Y73RNY
6hPqn/b8y/gAWiqE1hrzF+Ts1PsZEsrvBk6N1rAOuq3wsI6EnpaqB0a1Pg2ZzJHHUYoE+43itjvL
iDssP2AG+naTdcWYuIHi3mAAfxS/fRql4n4Tls7/52XKcj0Qn3ygzGGY6o+g77SQ6RDWKv4ydRkn
QJRDX+1vn0A1ZK2vXcIghyAF1xgt9KpOP3FzPn2/fiYdeWCevofM0gTex5lH0O9bXLWMDQV4m+WU
8seplEC7K30DcCwTNHGgzoBGO0z+KuUw6MbypOQCj5VZHw94vDCmrLrGfUO97pldlRy36k0noqFi
Z9ptwelXr7P42dMuOKhfznTB/HM2IyWxIKHTd/X2uYP6yZ7TACygRIECIZmoZYg5OUxxvYGo3u3u
utw/x3WUVPwEL3AQTaeLWo84XZntWgj/VMl0eFCdk6e6JhutRARRNoQhR/mjlDuGTE5zjSoFzW2U
9pJSPXagSsoWUMNMRPe/l8A6fPUgJzne4k4581hf7koavsGSGSdVCRGDl+DoJSxAZoDROXAYF4V3
VDjm//TtrePtIjoHijkyX1j5vlM6+NXswqtJrZyG2XZo1XQv5p3xkiiKBD4pqM8HIC/m30Bt+J5O
4/Bv/YVWj24/Rgdo1sQr5p5ky1c7B6ddrEhakJl7tC+Q5hkcLJdvdnCbpioBt+KChHQLFQP5oAar
mykc2FfSQkiMNhFSzjEckp+p0wkosjXDoW02mLaRmrzowBfOLPayQbpzcRmxQMaLoFzxsX0eNifS
9YlH6H3yKjcjsA41/YeB2FIJOJRro7ddhaxjkLUNoZ8nfCUPQhg2nkLoqcO+7qNJ3LyHkzAMMOW1
65YPNs4YGL0SFhmnQy/NY8MWU7oUKLEKzBVxp+K8BrEwImk3inyd4T7d1a1p+WCCOvl4ETjFr7lz
QPV24tz4wEUtzNMhAoEDzuN4t7yM/dp7lEF9czxH4Cebp+/gOhmML3rCGEklTHR4l3IiQKmtdIPn
EWbxIH13kgdadRxhpo+Sx2ZxOmGrn+IDP30o33gjz5gKn/JVCUp4V8dAMhRAmWyev+hJL/oCDTnU
dZtLBe/43+LQR/J2WrRss2OC5Roicm2B3oW8ZyWjOcFVQAw8BdXM/UpAhWkf2fppWCmK4Fk3w0g7
fk5AXcbMfesOh5QvR8Z/ofKSlNZF2ZiFZNvh0oQHH7+il9I64V9S/FkQJkGxo4yLmf+J4mgAqjfL
Y3zSsoOkhkTjGojXAEsr0+tsFmZVE9m56wM7tKvUl18JgA0Ozs9DEdsA00dVufIKkI95Zn8B6wKO
IdsIxD6Dvaw+cVHBts6NpzSG4YC7at4DZcJlABo0V9mfZ/un6C1k8dN5juSBTKPhnBg+yPO4D2LJ
9Ze7/NrklQNJUIoafghrwDeahsWkov8kzY7xC4eaYyDmcoZElzZPPIFx9jomUCVbosWhUAx4+D2C
+QXrSiYq2ZPHnU4EZ4F3y7r+ZUy8MCdRHM40sxU20wRanxl3kHHCvAW+muPI/TDax3HlJXc6v4Dc
4w9GCOrMH4KrQrdX5m4oO+dDxrwBsaIvS8U6acf7eVUx8jGS+/gO6M1Cv394b0CKtxwPbNVDN4Ul
6sN4iutwj3HHEz7v/GaBQcMBtijr8tlfV/u5jGVdoDlsBsRRGAa2sBd3Tx4ed8DYlgp0GEZpody2
bE02mYszrIYjRKXllSiLJI588cVsacDpkYdHZDWC+2I3rV+3207UUPo81a/8kZ/gW7hyf8zL23cB
ifu0CrIJISO2j3AJO5NYLOFfRzB4tbYPemifkJqQc9tH6bJmt8E8kP+BpqKUbfqBAxQPQsDq65ip
9BJyqziqjj1oBer+kqaCSQD/6hLgWGMe8AEN6turE6TXaIGi62Xnef4umVZSXcgaVRVTQ0CGJXNn
JDbL7w31iGdt8wectJH+JZ3CCyjspc5Ylc32NR9s40KFBVc11ZskzJTLsClNJaWXLyp3sNU8NuCK
w4BtFN0w3C3MjxoGWgJsSPBBhKfDQNvzW/fys0w3cEFBIC/9tYrnuR7j8bHNoXCX/TE/8XvNjQUX
W0sUUCHxpOwx9875RqV1GxAKA4/m6eIFhqhxdYePR+1j7el0si3nX/QLY1KjwmsWMsA7qCDM6uLq
CriAn6DooFEsIl0aVTCsexg5gPbSg2xXVprLKbjxPi2PlIAwmigF1QveMa6j0MEQ8KAisAYMO4+S
ZUla8X1TjLRl4gLJuDOoW98v5kHyAp4tpX18GawyF1v4qs73oVHf5PwTB7LZkPF44+BwYOGq5jiJ
XMRVZlnJC/8zFwtgidlIvLV7vM7NPRaVgVCdR15GN923A13To1OkHqWDslXAkISp3AceEBlPQpNY
pkfx4kkom+hI4kg8ZKVHvJ7MZcMcuFawKmZxRG0yvvo0E618SbP+sEpaevj0SrFo6pIWtr7V/ZYv
Fr1fBKB84u/O/d91IG+2pl9xiizIK2ZpvmQu3VMeo6F5+JqH9Cc4Qml65caiEJMH8LC+4Df9/we/
Y3qq9BvMCvoKC0az2oCO/PP+ZAzEVgtCTa64OE0wXqoK7FatDkDgU6YAEiWjya7yVNv3n0HtYBke
8ZqZbiTdFoum5JWXQ+8/LWrKIq65Xor0Xdo5HTjptHl8gdwiZ1kU+ctVTopQ3yCtERLcpxCVuaY7
8iY5wkh/Waj9L0/v+DBF/W8fSNqduFli/bdiJagPvkkpO+wSspltAu1cm+pQkLU95B4MnbfJp15M
GpXmRkVmjW+11yR+dz+Z2GLUo/94ydOf4tji0//wCUOJGYSwts3mmOgjXJHHACc1QAP1orELtzsv
GvDeQt72XDqKhGGNy/83VBmSTJD7mJmqZN7n+qFo0CBAAMp5IXm9qiHFDVJct9BmDlWxhiokbprH
IlY+20avU2dqVoFS2EyL7v1ssSynb4CcMUm8BRLJrNMqoiclxCGVGjHCmvIGW125p5bnGgos9avy
qQehFH2vZJKd2AzytUwsW7qDH9sRN4jhjLrt5gixq2QvLDgBzsUiKrQD8qnR06a9ELwkRs/1n1fx
RC5yqO7MkL1tbgZl8dANhnEI36s8bdWI+E7qW8jKFLrGWXHfuyiMolyg5OI5uttbq7vlk5OlZi6U
O25NyRCkr4sVUWeBs65d12NoHPSF4bBCOj+jEwZoPmYcpt9Ihz57b+XsSalJFSPRrtVCQUk4mETi
VrtWZBeKO7EmM5iJarD4UHeYgrIFqWdx9RSDG6bOw+vK3YwRvGP/4fPZcYv7wXiYNYWa9ILCzQTj
u5l3+lVOJKnLv/P4z86/MrHTlitVc90gA/zTZaqU0zYEVcpBkapa3XOzJGPiYXGgES+NWbybxSwL
ssgnDvwd4xEofbPPEhuNNHxswRaxOw7fcMOMyNym49j7RijIBjzwjTR2NpR8LmuG+THmeKrWIWIP
FgY7Iws46slLW0Q0lg8MmbXJFzbB3w+6BvsKVWRVJci+peUg6hkH1hIZzQq/5nk9mYTSE6N0iQ9a
pgNhUX7DIgHRY+XJWjlVTP9plnVLq8l3UJh6JyPOmsaRbzn5wgXbm8nZCi4pZSJj/BSPYAFpIfo5
1zt4i56C+CzXoT7rAh23Ki5vMqNzyu9lnoCV1cY7Hcn8pjKdgh2oMMbP9KCmItDC3QR+n3MkgUBy
Df81dREwvTF1iOnWi3TQxk4B6TMMojnw/ZeSwsBtiud+KIGPSwn4LuodA505DFIRaLfnX6SXw5N/
GRHSEqIZ8o7YdGqbm89NisIlWh3/XVrIhA8ymSe4YWPswTsUVJQLifupFs4cfeiDVLzaOv4PkkC9
22ztQyTwjA6yInYyTB5oWDbgYXCfTHEUiB7bt8VTuu8Jbw8G3FRhktM04oQujjf8fCPYR2Xi50H7
FbYV8hae9OG2OpFWK1xuZCp1l3NCJzwfpfY6iQtPFaQ5Ic3eR0+49W0ikBGzP8uSBIkZgrkeY5bZ
JBL+4tLb3KIat5W3TNKmmuouTczwji1r+MSCpIrtSi3tKazGvi0TENSs9vAGpcgqKDM8l7bI/kWt
73Yyi9hJnC7AhKrcfTEvCTZVllL7v9egWdsN0Od34BUdVig9kLG9Upaq5EUu8Ztnd0pu4wS3igy2
RIC0fuD3iZE/+H2AlZgpBZuz0dFycqGvLMHqpJX50EbTS+I60+WAg9INFnRlmuWZ67kYCxxV0WR4
tovJw/ud1Ke2mNntSmhrzt++Cdfbt2zPGiHQQowYSVB27d1KSN96AuT9RWhCWD7DGNAQUgZp0st4
7TPIqnfm9O4n/00br2eDGpLDZny07kG/xdANIQDhrx3/GlUjol8S6/Ug41ft9JiVsad3pMCMu6jM
X0BnSF7CxDT88ujL+FPxl3Mz72YeYHkRwYRm9vQ0EnOqH9oSXC9yir6T4Tqe3Xax3AQm8jSpClgV
5bLpqN3sfwnBYIUxEJso1vPVusC8Y+AUMvxIM6X6VG3RAkPKyU1sfo6M2hXmuOd5rvYqezdRWJoL
ETeVoQ9yI1TOHEmc8Ep+fFQD4J3ucIPOkU3iQa+gHgl/jmJklO/SH4GmYGLWbPoWK+mo4WGP+va1
xAz0OHkNfqr2iySHawDxzbUC+cNqwbX6f9I1taaxiKFBmMpC7OsWaz4rl9l093YxJikBYXE3OLYE
mPe5VwvBbeb7DhoK82qBEiyKuyDfmPh/lWbDSSGc+Fw56UYsRRwgcx7Dt10+xBoD1IcTNYiOBWBW
oSgQtRnuuU03aE882YHX1Zmt8i2rksYGunsPLtaQzh0+2kbKPHN2UIjgYzePeAglPodUPqoLuDw8
SlOiV5/GQyvGmPDrH8qiXB7C0Q7IFTF7FrM1ye6cadvVrAaRXwgI/21sX4KGTMA8AGM2XWOFhrPB
svXOCbWniI0yAA+V7P2b1tJ8jG7K3FvpA8JDceIbUTvt/5zPQCdSbMMq70NERhmi01qEIM6gBBuG
muCosQY3tcTsvZhhVlccs9wDTMqXN5/7vCriiUwSoPmn6cyXoYvFNWe0Y79pdEF/MgzYuJm4r5Fy
spDPisnBldOnmxusGlZZS7kU3yOrOTdDAfL0GkDIjJBldCYv3WLrbN0nTF0PV0qoDheFo2U5w5sm
E4Ca12mUY+s6rE0J+NJRt0uLR8BIMlRTLBARcVAefyYJtzFuFYMPAOvc2cHpFO/FKjnvktND5eoY
ekcB1WqpiS9iWfIGe/wTQwg4NYf6FYpsZ29yT9L+yYCdE7gjJP6nsLv2e/7lQUpAAl0S2vO1k3Pc
8ubC83w8p8SU1nlkKuL5MQKU0VMfjeTXLYhNREwueLS6ORI2wbqaGZzU8vtU44RR0H+OOVVi8ZP3
uNfkKIYw+Dt5IXN5OSJPLNetrhY/sivjLGdTx80nryOzFf8xammp1r9kriV19n6WLBSw4LjLag9S
60JMsbXsndm8LVZIjN7x0CI46HiqKk/2AZvYyHHGAEsGLwq+w54/w8fpkF3CtUsg1pz9PyyMxPDt
CQfreDsT7U9AOjs1L7HWmpVmLWKw/CpLdv20k0EkrQY5wsb/G2/0XqbJLre/NPvW5uKjnQ1NhHRC
8uPJQYRRfzh0Vdb2fELZqxbyRu6XJF5k4VWYEuU3bNEUcnuLFJMtqoZ0jA2+Ea+8tzm82YANm6a3
vgaT1CmbKQQmCV2AaA1HWqlQEK/yzE222gAkuR5Sgy3+W8si0Mdi6O84+QLlZLX2lPf5h1D9Z3lw
M+bI6kI1l6EQczVUxhxrCo0FMzi8i3MJ4S7v1HClH7tJKWOfQPBJhZM7HZRXhRN/fxvLm58i9fpa
BDdvHeGsozKNwtkj1/lvcn5c9UweTRJePUUVcLJlo3CZAKjEvB9VBSbADk7lesjf/AE7f0C/5NTA
wFQqgC5o1iLlbhM6dDgWUVW/AU9F6VOawgRVqh2BKCl05Z5NxLarNUSDLYwANNym/wEeSxIxmlac
3aRI80hE6POFWC4hPaBsgKFH0Lq6dtmlElcyqWOIgHkuXYHetUsEYl48m0PduCumqCLLPQk2fHdh
wQs3oEHUhhzOmQBRG4vRBb6sET0cvRAFRb4kCJVnPbNxAOvpWgAXFtpm3C2yXeIIWgeWNKjXtF9G
p6SSLRIIXp/M9c8oYZyWUQsjBxt0alKrZoO7OPxcDXZ/2dO/H0Uv2BvGF0TeSsP/UCwQ0xLz2XGR
FoCtnCNhISEB2ED2fm2ZWDpO8FVSX4lFuCAtMtwnxwUf7EXHf4BBGKjrnPGWrKkqgytE3fU4CvBg
7ZyEX2iUmm4c+5IJMFj8U7Ok5r9PIYg95gAUrCpc+XpnocRMpu0pHChWxyZo4W71UJQ3DtwaoMkH
o99/BTcZM8h3dLHKDJsldgnhwe1xBOSk0o+dVgRfpuliU+6oZx2y2nOaAv7bCRZd1kvbLOtK6Emn
8+JS2XGL0RmrK7HZXF5mymTMWrzEsoz/GkqESAswTY+KDH46WSzvFWWT3+uyRKJ8gqsvOr6pGUYQ
Gv7FHHLF6741DTnp/9ub4AvHwtDf9jd6bYKhtcUmcVbSIdAQnkwrdAuuBS2gCZuvrA6LWiZROzva
9+ThkCL5SSbraFG70DCJgf+GGsZ+E0+RpHqtCs2urdHbnuAhZxJueD48xTUQpKVG692ZJ0MWXtqF
MLF9fBjZWWTQdiPDKRqfB3ba1rbfJlQ0t0ZlIPglA9eEph54mUOH9XiLQ2xaCVbmDNRjNdykrIgx
kiBDdnMHz/U+VGxZ3W5SPIcGo+htajaStsoAuSBLKXsMreY3cOCtr7p3nHA4osrWLBBxfEE8+85d
dY0jBUNP1W7j9WnPLlSHopfrbmXFb9ktzeE6ecR887e/VD9mwt4nFOroSBCkL8qdRa3sk6kwaKWo
FAib/BXe68zVEFtosbTBmq0nhS1bkSzJF9blQAAwMiDWvifvcKh2wOrRsfM+DDxr4DwduR9nneRs
pI1ilUfRKkPNWFpC39OtelswIjWS18Etr80WlyVPj9UtrfJaRfj5Nqv+4KckFt8VEgUl4w6twyWJ
1SnTtd8vB4C5y97NaoNXmHTex4XOHneMaHQE6YbU9PAyPb7hsIe68U1U3YYHKllV+X6Uhrr4K2kA
j3WaPcKH460jo+Miha+tR7iC4g3EPcawi16Lhkzxt+kC9CQarDm+58UHD7vRkChD9DvaJqE9+3eR
EzHmQXlWopxJsjI6YxyWTQU/cytMmS3Ll+1HMUwqEAJxbr7QSYW7PhugZc8Wd1wOGbn7MMG+wdHt
u3MzRnpccXvQiIuDqHFXmcwZUustpx8Vri7N4Md618HmwrOSg7q3AZhiwaO7Vq1DQfE6Gw1HTXG/
ChDu+9Pa5jyjviI/eOsrw8uOpre46Gs1gV/ce/270ye33BHbYbd4UySYsHe6xt8VMz2dIU828cLF
h9nbWDFBRKn1ULwkJvgOrJXXbX/24DQTsU/yrsWNJkDkGolxR73Haw9i5tfdpX5oGkkoeY2EVHy3
Zhl0U31T9y/APBi1IFokCfdWBgfgp14QMmETFof0iyWxXiM6K+teig6Les2TjdIw85m0/J+LrlD+
l9zL32zeTEi9BRJIMBr1pdOqOlsgM+aVhrMIxfVuDaalvPfQgiA2a1WhT4u5TU/Vm0vfdlVCJOTa
TNEDlCDeCYDcgwA62010NgNlbbaCfEE4cN7AhTkpSUF97hZWcVTJKHGso7MG0ekQZg25EHvcSb9K
/OERPIEgC4luW+LAg8xWtCbYpM07VqTYyR0kZbHY0+hqE9TSbHKz+ZLu+1s+vSPnnV5w+XZzJ4nI
zNn7+0hKzWQ3+kno/JRh8mrA3X/CUBNDtCF7z2h4DwxzuT9KoLicFVePWwStCe802/tQliGVcCvG
EnW5oLiNhUZsXsJhTwE5rI13UJ2sjNxQi7ijh37d6dHEam6wanNKSarnZ3Q8mb0z5ceWPW9RkeK7
mfjRwC839pPbe3se2h4NOy9NckGfqRVxhflxbnnNilgCM0EtJ6670RHUgsz8LTFO+1ywLZXzoreS
cHd9io6vwzmFuoJsyzj87jKTa/nhe4vELgjuZwJyZbyWfcAx/Rm19jjJI1kZM7YW2PRlW4P2OKD/
zdq94GnVNhmVoba+Dukh+wuGkvle0hA5Xh9dRvQzBdLQYYHUjRzaeD1YoK5c0aJJLrmQHg54UxW+
qCVhQLaq7i20KovaRaoK+wYO6toc1Bp6sLzfRFr53tDlnaOc9UN2Svct64nRGruwR38yt1jpFGdn
IqbLiZYLvpCRX6t1lRIcnhaTAEi9ppMTUHBgDWKMJ8BoIKk6lt7ZEh6LfruCb+aQjcbEGexZQ7LJ
4bR6vfwsXnbOaZRr0lpJdqVkNimZSpP/mc/VU8AzCsm5SFa30gLg6BhW6dUN9QQDLzKL7SDoYPMf
mPkYnZxiilZFyB+RLf0YqcCaHra0F2pcx2V0wMuKEIXckfL3Wo2tcMfGa/oEKmrG3XnXuQZUQWCA
qv2T3KbPTvTCuHm5Eq0d4OQUFO3fbKbskCtf1ym6n/kSmKADvFsqbWYHSDWFXerqdfZx+F6PK9Su
IadMU6d3Yr/9QJI4p8J3lCjhvbNzNrWaTKGBD1fVOTDWyatNHecTrZ51vVB2R8DR2/mPRX/frARI
qg9RPGnOMWxkIWrFd3iSLO/xbV8GYu4GpM/4bMbi5cJLgwHzhz3pbCYkjhFdVSc0hokqC+aofEae
HKbD7doTS8YGabq6TzpjHOM7iM66qg4vDTd0W3xnrV6/wYyb4OOPfEVXHDlbA4Fg5Z+Lood/KGRF
ugyfHBCJuNzanjczG4TJSA47jGxfDpIMyy0NDf5wy/jCy3TRUWIWUZFE8rU8zNrrWMUIq/GZMTaq
Gyw1bmjVi2/gPZoOVHMTU1cVwp6q6dvEBkZbvU7kAZZ8Tilt3Zsi3SzdfRo8sW70cOuLZr4Kp7Mu
c+jK3g3UOKKPxU+KP4XpVaYVGQFHUfWsEwYJknLDE1/FaOStxvzgge7CWsn3Upc9KmE9tcKNXkbY
MFlAwsme9yTV/E5VoYGxDut50AP4PcNNizN8CkbrEnymd3se43JOV1GIN4MDPL75HznXZegBQWaH
7VGO8yspCk0vBFgkl2TO8BjDCLtxxpKpn71qOsdyhyovZki2UZ8J+4xQFHO35LtslojMZQ4SLSNs
UBMbsPB1049DSxHD5Zh0Rq+RwyQF//dkGv8YengsvM72l9T6Z1gqPNPM5oIjuRx4qPy+zIhKPsNl
6emPVGiI5QXzFY+ABYr9+Ga5PZSYCIcPlzBi2L18QlDrqJpNvp4cy+dXwrR/iubAJkMRqCXtleMP
2CUf/98n1fTx30gTpHVyfqmu7qWlPW/MjkqdtFlTKycJoMrhh6MJD/pJZLgFNqbpNdMk6jGSD933
Rz/M6x9FX4RBYrn6TgiqMtvs9fGd5EoGxhYTO6u90ezbzSxFoIbfXZ2KYWyGgmnGDi7mC+D5cAF/
L55m7XVxyGbJZXqkhunSj1/s6x35E1ic1I88ohFjakpOu+ahClohgmU8uhmwUGpaTkmssUjrmEOs
Hdccv+NKGlMJZFFeFgRLV5mUNpit3c+L1htDiaT7x07HwggSm/wCX06YCxNCNNS054CHgeVTPfHT
7kw1ronsmis2qhRPZEz/YyyznlaW9dym1cr7OeOg20Gc8wEm37nlPebIaquaiw18NIQiuXegnKKD
PTwGtVMiakfHB49NDhu10XUzYt/MVbwANz0NVGGez80yFogucaI6/kpp9S8sffhIfqHjjiuTDKSn
7IqO1jWcCJayLkw2pstoHelGb/yJjZPBXPa9q0Nj5XzgmwuJmQiShYsKTFJqPi0GQYGmwHxyJBkB
egVBpaCLJiAkjPpFdXsqRiuIc7hxGSTJYb/qA0pbVjZrwNkLKgP62McHng8FrJzzwU4+wbO6Z0Gv
qeAExz1UT6sb4Td3+hKuVPBmSOiES8kLc1taVTnNSoSep1Iv7d6NcF6ZSkWzJoJ5cznWwFrXWmeY
vJvf/lx0gmocwryqA8mmGbLiYOeXrk13ngAHMc5VDdoLI19+Ewy6uGh5V8SasEwy8NiusDW95diM
+kz6CthtiIzI67kC+wPMcmz3a4DLN5PQ/yGefJrwVgJqGgel48G8PqgeJH4cACRuJyCd6J2U8z0q
LODB1mPFItGdDoiWYGEKHznjoCzjvktsbTF8YPqZGqxvekjieUEwJaehSkiupEpuqbX1bCEPCg68
w1+wyfx7zx6U+Su8Y3hmEJO9o63fxSUm16ipSKGQyDy8YXIwDgYikw7PLzYFk+09J8ntzDLU5di7
MXoIxKtcd5pEbzYBaPrOZXvft1Amz0IPxVN89Dcp9r7zekbH37Ye3kfoUra2LDjiyh8/VAPg31wg
nw6EYRS5ki4DkpVpNOZDoHqd1bSLhUkQvfCy4DHrWrCu8ikfGp/3n1WY+i5gojoBmzt7xtqW3phX
Uofy+0k44UeN/f6f7OIfe8pLHFuypf9Hdg8iHN0YuVYm82DEsr9W88uPfGseey6naAEcPlgtnh+N
DbiV7TVbjguutmPksdi/9PJkfio3mNICqwSSEvWzZHXV02tKmhYqGQ1oU6NF7OzlOnqAwtXqh2oU
3sJjOV8SQDQhRGs/wdKJ/3izqjdbAZjouNwO5ISDI3dFQEcIVDpDIxAmiXTHDHCZAEjppYr31xAi
KMqHAP8VVkDoLO476jRG/HgtpDfTzZijnKndAAC9mIzMgC1CD0yZ8BNjarGTHqSdosvE0OWZEny/
1WUU7YbEZIomFPlmB4LKhdaLi1ha/RtU99cZ6hPQx87VhOx6k78rFfK75nZQQ4ju1ePoXAPDBsBZ
pVg4K948Zl9KqWccueSSkuwgDAmeTqLa/JrP2QCH2SzZVpOCrShh5yL43zKKJ9XU6pYjcySczvXw
EKV3DrkZNzMWlFCzaJT6IYfsr3QeDwUM4zvakJfhZnKMkgGtoHEuYo5DIFXgRnBDd6ScGSq/f2eS
n19Zt1whuBcpdJQiBtVKN9roXkT+/pX4FmHQSs4e7z2x+7gBhFqIgnqKgQ/aJLA70xRjpLYhELuq
S5YV2fxzJOLcfHNFR2liI6p0df6FPA876oz0/AxH3AxiH2VK3U2BS9xAQ21CbhqwZsISmUJFu/Bv
PNZ5W6BrjETG9cbHnqILUCyoRqfOzIUooEtt32x7jgCRWTggrhVTLvKMY22HaqU/yvxoGQf9wZKE
NRdVE2gFsY2QEFPEEHJtrT5LT5PwZK8uAZASFaU3dDycXniPGvcIKNh70VbfCXNwP/AR4s/hkrX3
XQsu7rEWH2NWEKibs+dN91eYIidFk4F1W6auRShwM1lcuHQ0LtSontnfIoLfNFKKAeMUSpq+Qrh+
J6ExCw8j1ze6ZGgpml9kbaZPitGEMURQPRJa0CYbTkDTD4LOkk7WQYHqNcLLiVQ8SS5+Lk1V3/Q+
jvG9vAI8lXjs9P9yUjGD1R/jFlpM48dN41ga9yh8DaWHLbj912SQWIfl1mm/8Vkl2Ko1uNKafm3Z
pplGFIiEaenDpJFBvUrmCZaiGB2AfDFqK/prk/D+zKO7abg5e3hECKCB0C6+UFuU03gaDqXFed74
LknYWHhRqfVIOnDZQB7CS2RAeyEL2TfFND9d+XLcrzfQ0msz/9nKSwSybgsLO/zS2azE7a+MwrI2
o0b5y7Ej3qI2wLEPsgXhkyViaUVKbdl52YbfLlpOJ1E8OmwjOOUXvqCNVyBXL1EpiAsMTSSk+lLF
2bUQX82QaeH0gTwgFKdMlq6QT1033KKpTRrqa21MmOEhmmUUDJoJ9j2fiqwPlsRVlgHZv4aqPY0S
ChfvJiw4D0yzZ/uS/D9kg1Jc40XAoNOt4NODN+tb836AueX5243A7YKFznANC8iTRcP2CjEAGYEs
WnXNTVVsyt1vDlV7tgwIA8OBP7l2+GSPLF/XqF0XPtZjLMIiGjsNwvKZMRygSPSWMUbFAEN2C1Un
MTwu75dlR4xZI0idnaF5x8eQGmipaiYQng7q48mDI5cV7U6zKG5SFH/HxDxXYsETvQEeXAnEVAWF
PtC7rwupHv09l8Oxzr/HaVDnL0NuMx/cN9/iVhly9nSI7GKR7zPbYmDONmk8y+RdbnYfE+pxgOqP
mE1VZBXu8m2UEUV+RIi6I9CBfQQjKgq53tkzd6rdlZEpwEs8me3otb+CgTqD+qGNU6QN2UMuXDac
+GiS/HbjgKDMZZc85ySSeMO/DvSwAnzQ+9DNvpBXXxVYYlxT3HE7BowIX8bXk11gfrTYOG6d/tAH
ca+gC7CGDd33IO5JL57k9IjK0ZWqcfVdagjeOppUizLr8z6ANUKuyGvvXQaVDh3iT834+i61mtq7
tY679dZus1sDNv+Z22jHwN6cIh5iBIIVjeeKSbt8pp2JsEzWAemBbjAiglzbSCb54ICVscNUECI9
VQQe/RCsrH8dxicdFlYC3FqVg6UH1IgRWqGTY+FAirRTe3na1NRWJippjHpVevNIFjGMRKWxJqIH
BQccHIFV/Zn/SueI+gnIY2d9WqWPTr3LtWMBKrXsb7F12pMbTZrRtAZ+/YxLutRQYnsap/+MRWFN
PRgpPdW3In0Zza4go0NDm6gU3wQAhL253a0J81oER6HmLOjIHENENns2QmeSbuRXeTN0WCcWKtiU
Anc2wCFNMmvlr27ZZRqe/ZVJDPdkyIMpW78vw9QldW8xkoRyrcW7CBfQ+jSBGOzHlBWQBqIQL+Kl
h0oSb27C1mcAWo/1+SEvMCzwcNDOznH62TnCejWwZ5UfYm4PeFj5vrJYuOCe9/Yrz/yemut/ixpX
T5VmGRzPjGD3huGIYaCSvkQDSvEMtU3RRNP7Mk+Vb6e0EJApuGOK9VvVDPQAu7jkkVi1uafSvVI0
3kAarZMfX6oawfDVFC4xoszQMfrhUSN+i2ggX91PF6lT54AwBP7LeyIZy8hpRo/WJBcXupuRP6Xn
+2irO6YPzp4PbLoGDEb9s9rQjCSf6O6Mi6c/983prbhSf5WKrx30nIH/N0/ZHyATRpcUJQS8zvrf
W2F/oymiyWZsWLxUJdkTYFCfD3AbVP5K6Io07cc/RqQj001n4sljJXnMGqAQih6rn5d+g04j75jY
+ZKzkdhctJdN/w1DopJMfNdM2NIYynj3NSwoXVgXFCXTMbLjhPt47WpZLjMZzRok7yXTRvdUSBoW
jU+dG0YuDDLZE6y7pckZrWb3lH4FlgoNJyAZI331N7wIjEH9hftHMozUP/JgklVK5P65Op4Wfc4n
GMJ91hWl5f/MSAdoEwQI3NyCJ0lQzwOQG+L5/t5lzHMsXvfWS62NSCxvAkMHiJqTTEugJ7izsmNw
UHznW5JW/QeEnF29CWB9sT2pxiWyrMru6OqmyzJe6SY1Z3p+nEBATRv00JsemaeE7TgX1/tF+Rv7
lGVxp/6azwB1rZyFNxSphFDQCzuX+25DuYZT3Aj2Q9mfG8gS773bSjs/4OR5e18MIAS6+TX/ITXS
zXbk8DTwSW2WRGyVwcPVDoPEeg5J6NC2CwSPj9nIVn8NS0vrg6ISpBBTOoqOS5rhvd9qj4xe6JTu
3REs8oMp1FGDbAWSFqq8vk3ZSwz3vlEnbW1K72J9oGhbAbJu0iRn88ZP3w7nlC9C0xzil4w9iq/v
XpVpFdJF0Bxh1RCEIETNhMQRwOrpzSRvJg/yr0/t95e2fByhFnER5Jty/vTAeLlWWwWEd4x17YXW
vMb0n1nA5thpXwHKgtLfbADhgQPOIFW8/2zJGV6ksM5h2sXEu7V6U1mglGOrqonx4XSbizBu4LdR
Y9Gees6gy32mx7moV0jXV/qnpm0u/BbbV4vv5bYHqG/ff+SLk40nQ9HqEIgHfDB65pLiyVa/618R
NXKdO2TUDBJzDi1nb7P6xLwLNcQwwWBHV961uxl/R29Wt/O7o/XRsAgoP2fMF8w/af1czqnvuNFG
JVZXgziRiYllDLyLxzsPjj4mg2tZiwCcakRsRsW2PrwTMMsxJBmMFb7Q+ZREANE6NsRyJoS3Ep+i
IUGw6rN1KUzp3TP1HBRecDJckD7Av4XI5o2tglgGjRPJco4OONfFrfHWlEAEbujFNi+58fLqxREZ
fVPnwUTF4nDK+qAWRWfnm2U9WC+fhxEf0dNJVJZ0WZgBgrDEIPmbh9HRmxO/gmx96HK6dvTpOdt1
l+WFV3GHXIHLYXEqwMxxpBkVkIhBQLYLjB1p8pDUQ5I184deb8jCpo4c3zB7rfLbhHDXtOySp3m/
Fe/vV6HN+iwPQapbCHQJ5UI+voJryQWoAk4E0iVXVxjynz2gLXpijsdcXX/tfntN14z2IIwS+oGI
D2eu+OFa50QYAoFg2phcZYVz7Sa/xNGxfB+TwiHi4Ep54+QFovgv0SldQDZg5YrYVsPM/XXb6ZG7
pgnEloa6fNeZ6l4sUtdZ6rh5W3/I/hn/QyABLIrGHoOfUSNnBvqZ5kBSHx2u9xGOvzgFxcmg87Wa
adGjF1J2fLeI7IitTYAeVc1wXgNJaix3qoypl7hCAEy1ztxHeguUtXx3IFtqASABhGIAn9TgM61O
naL6W/nOBxE2qPwZ9sqsRj0H/PW44F29IAC8PRIrt06mFgd2++RW+SmcGHv4lbAvMppiInVI0dG1
N3GD7hR+9QSdNBGht+Y7xPXeilOqNAWW/f69720V4Naf5auEhtnBKFOt//TYJ59dE7CiN4EsuNsI
bfaBL9sSa4Xw46ieQ7oeAkivfpKuudJpEZei5RplpqBwbj+3XaRYeS91wcHnE0jMIf/8sClGGzgn
gFvHLFWYWs9YmvmtxaFwN8IrO6fLYF0LQLKJ797aHCpScc+EAshK/5lRZv2R+bm8xf0KtogKMvz0
p3nJs8N5+Lc3JrjXE++uvhfw4h4HPrtVQsxoF5cLtOHiRp9uA6hmcEomTTECGN/gp6KWdYggF7tH
u4EQrPJqiFRgAdBnU0H4UDpzuNtraWm7LYPu94idIgAF3Xc9eBrTViNg37EWvunFXd4Kd+CUlKsx
09aI4m9b5jqPmtRSkORdT6JSoO6AJ9nUS6E+uRloj8G6CYYNP38t5iLew2a+c+leFX2oqAG9iexV
tutOygmyPHTgMzkBY6bma515Ucus3fabVp/qZV0KEJOrgTxGSifaSJdDYlxDbolbNyJCCAx42byu
v9nTP3SpRjigun2gBS2V1FPuSI8nssdcsk7ydPsMb5JlE69/q+BTj8WLRsgrNINqy6SM2n+4qPYv
u9p/LIn3CwMWiUAJ+VnnM3I0y9CBabMlRZTEeQeq/AWwRAlAvzg4AN3siZUUclLDhiqInbCaq4Ex
+x/q9EvOgW5IDTBNN7mxnvbCVBCrRWD1kq/7FDj2OOHPOmR6s7DhzL7OVjX6C13iFq/Sh1kxoZcR
s0MohIbTiPxAGUp5Wkj4xIwPOxWG0YSdKp56AWNDrGh8PTMaqSseHH8+Ru3/QPJb7mASoUsQhWed
pZM3EQKxW3RQW08njvRVMruqbU+CybxPbOO+emDg/6s7P+EaHu3uoGxMUlEEEKLD2sD5sAFkgsjE
mrRayJUMMJFkS4k8cnNZIzxjOiBSgOyvamozBWrD4HkP+mC8mJRPxA9pLkQAhLaqtI2QlsJb9zTV
rAwkwGumasXlMMo9rU7K8G6cmEVKOp5WdYmGI5s2ahqti698VhnK0M0bqgC5aMT3HtCHagrsxqkC
4VwZw01rAqGJodzGR/qEfhQKdo6S6STupINY/mjJciiA0JbECeww1Xp+ozRiPBhYESNHKs1hjtKs
fe0ME+2g+9Qwt4xodGadyw2JEpWi4O7y8lXgubOyw/NdDaBfAKOcBlWNpk3nx+K0rSNwKS22/of5
o7UdXj6b3HjNv6ClCPLjQZLAAtXB8nBbhHlU68SLl4XWea96MvlhdSoCCAum5mgo+b0mGLZjHJ+A
jrYbUTaggK+qc0eU8pJkHx15S8D0zZlnafe8Z2uP9Z7W4KTUb0x3M24qrWSSHQjKZVlJdld9I2IB
YA5ZgZkkutA8W4NXfF1RcIeL3NWyCUY4VKskt0iAWElSjL33lZvi4D7aOrJqZp8P6VaRyKefRJQp
MLvfdNtiZd9fqIWT0F1iIGvZ9x+YQ3L+nGOXBBmGr+OsP/FLlw5jKXpGWqCxPYan9HIeUmFKUSgg
WEauYX4pSZedfbsUt2NswSdBDvWNXLrG0Y18FYqrBVb81Z9FExsVoESVWHIuSyB8sYg2KCbddzdN
nG33yDBnUckGv5/5ZxwxdXq9BbXscktmZSNtFdplRlpzRTfB6dFj/3kyHizt1m2nNi8JW2XoO0Yg
hECcj+4/eS6VTrfQxd3P7hnwUYrBizoGliG/oeD2/ACY+NNCfjWyO32CVPZDnKtnX6JVyQX/ngky
KFVeqBWKSQio5EKI6yK+P32iu7aN4BlJKF6baYJmwZADo82AI1nbJ6H08ERkSG1UY2O0YgoSD8Pf
7CjlnAAVpnar4TsabrOx8JLIku9FTO7riGkXGh+O1whWQ6xJs48mmdEZs9R7Fq7zeBOWfx3S7L0K
HestL6eME2e9yRqJxaKJsWVtsdNxAHhrwKoaQ+fPgZSh5FWRa/Y6WVek7VDHrGy86oxyBdpmySgT
/VytrfQwhmUl1j4IIGljWifcJ5Xl5MU0N21LmmBO5dwHkFLqe4J7f4+rV41S2JMzP0S2dbh+ySP6
6JeeKTehv4AqiiZs0mTHlPHyZv2XA2dPlSo9Ulp/zlWq0inmzqa6xRbsNgvnotT2kPdqQ1/Fo7Wr
zHmWQQdeyv9eemGI8IEpwlbe4TQrSYJrWcO5r8+bTGcmROje0eJ0ZzQdz1eJyjI6UMAopo74X4bf
iyJlhylZ6CQ2Dj+3iGo8BFyd0vQyviGiELCOePjcLHmZiwGkFzXUiUSEmy6y2UerGtjs2aL5OZNd
vSY5r/cDiOxjXrlkkrzPTNcIiC6Aq1fxe1uwtUVPWcuDVu4qzyzYmQlFcUVh1NyUxSPYyMONbL88
LNM2mFnWJzgNWjBNplTYr0grd4yzLeVTqdaqxFw5UD/2pHEVwZBjhf3bQmqkITga2gBu6T0XvQhB
a/YebcLuIm3/ZwTzVCGwvGgs5ArVAg8Zh3gcaUnMO3WDnfWTJc3f23djtlSrCXy59fLpY3EBoa1t
s5crY65NShwoPGnzEVEfY3A8fHnlp5W8SVd0p6xVOzkZbA2PZREmAQ8ijRv1Gc/QQFkfTg/KGTgv
TJNNDqrGB3NrQZU4MGRFvRAQt0Qn/Zzz+v9z+HwjmEjaZI54sUGGOLFmVaYEO/gE98tGsv4PPjK9
SJKNHVmATMuQGfyBPpZZCy4xRXrtGeY7u/WEbCLT0R9xSGflF5Wjx5bNNWpYEF9uOIi84J9s5+pc
ikYKm9WxEt3O/4x5JRy0HMBb8cXp7iXnnc6fqikrhd0FgylVzY8GTGnHCkn6SHNV7YmybWvxnPXN
l1dV9an28HWT+ai+wu4o0OcYp3yGGH5o6cxV8txoCobPg0fct8r63IybVlINIAfoljk5sd5W1OI3
kUewKtvff2Mvyd5Vxeub3RlO3JfWKFZW21tKPHNy3fN8p72jfIMiH52W463YBY87IJO7zzomhxEb
tCkeOEGgvujSqgNEL2TMKUYJZ3fVyoh4TvWjEYz5A/UKnCoOsyc7JMqGx382/+8a+p+MkHX5600j
VW7EpwWS2jrVZOiITA+ddwDvOMmBGeW+FK7LD+Qci8gG0uek3+cQMo0TdTB3Y+jips2BGSX9tQ+b
+Ij7epp9KAhMnUwaR1zMdkBwIsgCL8FJ35h6GNX9Hw2IZYDODnWNteI/a601VDP6r+YXzrIbFUjq
35k11NfMTths/eyb1hmvVzpPZets5mnYw9BlwjidDTnWAYfhss8EpljnTqGIWpAthyVuZtILhKHo
zt8xtLL4hAOLH0QD69hEzGk0z0pmYA+YtoQ/qQB1+Q4Tis23fpS/vNi3AShJEqyPukvSwazFS441
7ueO2bDNhisuaGanSA9CvsLcGSjMD+/fwpS5RPQl4rrRSNvFzPag1YjRYNiC20UzgmtwdwT6nMj1
VH+5PBvfwS+AaLHI97CpK2h8DCEGO/lqX348SEOnZIY54umpUVjxKTx9t1X3EWk8IWLBj25OYXxC
qQsAiSfmEnMyAqP7T1oAwcXMxO3Fz1pZCR+cLTH9DSSSiFknH6Qkt/BV1fzmoDSXLJ5aT4G/8z2j
zPv5TysIJrgwt0by+6KeDQ2ec71rgcn5NVn7h3yVpii4FpjOZhHaXNiIeyagZm3+a1z4unxkGrvL
uQU3iyzMy3o8OmW/A+LKlalHD6TmISoxEoBjDyrJfcWqWmvUFLIHyrWCSMpRtksEViQy/29yAA3M
EzNKYB0+USnKpiZQDZUcaYIaZCxRVT3ORHyDUwIIwmeOaocyu/kBRUdGvAVUI9Q+U5QQv05WgxBm
/rTGxn7qhiCnTFfnVVJEgMa/JgZyOLB7evJ8XHmI1x4AVCnzXqZ/tmwkqbTynKQ5U4+zpHqEho/b
HrapGfHkl/RKtwNk+XjYvbP78zOEFctiS5x0CYu1miq2m9xj8qjGibDJ9SkvyjVeUw1FNfQmdqvT
Lb/XNYwwWXoM5YMrlv2zXkrAhjjFgeboeD6QuzR4k98fhNHZl/AWzp8bB2jFazAECkPYWhCorEtS
EegObELf1Pq14JztscmZNK2Rh3p9ZRLau6gVH6TmJpLNk7gr5CMvnAUMnp5CV3CjTqR84UEhzjUb
ZIaAkvVAvgllenRnPVe2pscs7W116gb3Vxzoe0gBv4+srvYN5Vn1/hCIXSFuLbSIeILW4VxNzN5M
bB2jIkkm3/EDGM6L0GipE/5jGJI2KCH1yUbz8IzgIsGqfqArvfs5NW8d3kFygCttgetSQf+klYfI
vqBN+xS2zkYUe9b119bRnvYjw8VblJAuqkemtBzf9wWnPo6d44XrJ4dIe7/lHCypuidaUQbY4iHo
skSAHbRsJtPiKnHDtR13gsp+BBLmohchVmrUGNbhK4MJS7oUTcQfVZ00E/EVwTDsBGMl3fiP5RgX
OufUtuYUxwwDlz8GcH7Qsi6MGHzHeWthZdWnrcYtNYyrONLzMS4lqRJlpIZ3G1rV27kioq0sQQsu
GmyWyxOeuhbp+al6XeijMOdA5kxKnYDfy5B3SArVPUDKDUkgXN18goKI6RrTXVWVq25FJRlXWO+/
2QX4rXjFlIEos+GqgwsHxfvvHsKu9jZC7bVG0gBBmsyREfwTJDll1pd/mHrh7BjrMgkLN72Fdsy3
puzYqQ1nppXRQxzTd38R9QSUs4jmNB0RAtV0ckRN158b33iz6OUEePdz19uoiRq/N7fzas/rwWC7
745ZTl8dnkZxa0/xjv8S+cX2GLiV0wHMCGJsgFvydH5Jvpm1uHDS8hX0WPts5eD/r+nfwabuKpsP
NbVS5gqkFrUsaF2NOP2WYxg1fcUNOEMOKlTDYmotL2Tjk+Vx9ny7VlTTcguXVnm6JSitH7L9bRaO
WLfnfiRrUDc+dpkaBB2vTU7CLzRFjYnPC406aFi295/fgqBhTw1ExAiGCr3AHU9q0NCRC/G2gNsR
JtWKJ3b1tz4ASXnBwS/5ybxVgULP/dWZKxpssZ9GYpygAS9mjUZAhCnDrfNguq5mcULG/CgMMn02
qDLY7t4/e1KOm9A8Ha2ULuZMZ6SAUTQBlV1xtaA7yHCCmYIqfMucFRrA6pe8XLxa2933n6mocFT3
ezpIPr2wk/2wuN+RNCDe5KIsfNpHLXMw/wNDcMf8IdJQjhh+BLNsNbSuEa/NK2uvSREJSttxyTQv
wlEYSe5cZMp0I19glnCK86LE5xWegf2MOJRoPhufgVlEdEWIGV/05rHkTIqsJupB3FM7L9UMpt4U
pdvUj4FpN3ku57k8Zjc1ds6kMLgAb6/Bcz+22k5mRwpgRJg+GiEWnnH61wEiKC4Dzl5KVE4eT54/
8HlxKJMWEJ9A5YAEWIDtUEsZwQGL9THuk7qfCDetgQ0csWWIBTJHuB0r1hAyRyWa/yDMUHT/F3TG
bJVXUMJpLO93aNLgeq5CzW79H0YC75nkrIYPSeopea7nMTnEM1OUQyb/CWj+Q64D1emgdseO1KNF
kyDLZGYWm4O56Tc3nvc2ExgIadZlBuzlizbAwQX+aRmd+EwYLSxttOPXCsaA5NuDv7YJ7/CJokJf
sRypJdTHD7PSvXGkvtAyiFBP5aI9qZ3bmgbP29bgxPcj90lJNNy5PEPTXE1hTyT1VjV5/I6d9HEz
rPdhhCSVRv5N23doB7eiHhIwWuVaJSp3ETtaDL8pmNXpdEFk4mNLVuw4tqRD+UvlFD7FDbsIwT2u
y58u67gcMorQyhVP7qIorZNazb5OT2aVOqwdx/lJj1Qbd/DKffaBJt46ps9R3h7/S/6DVtYtQjzG
HZT3PjQk+O78HgDzpWTAmG57gxXhtvs8mSGNNqZZwLw1yWkanFSiENLjC2G3R+/VmaFKTHG8ETY6
35xH0yg5sa39dRASm0PIO/RoYjXAqmsrKJrrnf77c8eqjpMxYQ/KKhYIdC0olzQe6mLSSD6EHZTR
qb/LI91otjyOtPxeyy8z1djPGFhSDOFbROv9J4II5PxdOrJpknYBUdh0u4bGFtMEgqbY9AgHnSyL
G7tuw2g9flyWm9EC5j6JrJHc8l+PCgykuwx+zzW5x3suZatfE2W7ltEfsxFhUk6PfMqMvtG7gwvg
JKnemtp30VvV0PSxc2trJaD87fkpp8mfS2t1+5XvAYg7jgIl7v2epiaQA9WhysOeXjUJF9bCxNqE
sB+LP+WHaYoq6XnKahyg1/KykvQ2lLTO2s3o/JnzDbfHNNswCMP1/+TzL3qKQGQgKuBWUaKg5Fny
oip7xqN+CM2GAXJLYIhlPmQEFLV2Jbg+AzPP//lwHzyrx4E6NfRTaoNHFKHiSZ+uGLQE4oqjF/MP
ShI6FkErLCjt53/aww6QYA0Y4ZgN4Jcbm8vsv1c5aeGhdmDRxAy+438GkxryngC031EVe0wbylU5
zXzm5RRRQDjL9RuEkMRfT8kCVTNmj/16OjMZY6XI+Wajyn02vYFs51V3cgo15Gn2NnLX6idMtZWr
3e5F6y1KC/HpfrFDy3MDz84ahmMPDlZxiXUASChSGZmczBQQ5fbOxIcGRyO5Yr7QknY1H/zCesk/
UCR3vMGLYLHNHXuIV43a5h2I02hsDCFh9W8pWTQFUe14trJj1a12hV+c4ywRODFRgOmUzQr7SM7D
nMv7BeXhdVTrANouxA3krpGmGwhREUFSTtYT+86cRQSC4j8u9czMM2OSIDMFt2Fknci1apptE6BR
B0beYEhps27PXB4OF2uo6KlVrYKjp0HePTHB9RcOy2blT+S+QiTL63SC3XUurEcKaid6Zw32sDyr
SPCgm2vrr9Dtdr2QWIdBnLwpoBIJ8bJ4OTQtf6tmpvY/TrHO2Hc72H7aj3D0kYXwZ1lZWWdnvaMm
4kFZaqFhL63FvZgoDKDYSvqLiJVaGPX58KKzbNuDmeq5OZW+Tq0WZC4igOnJqqJ7XKsQTXZY2+40
ROQS2c4bY4xdPTbmUQQjP14Q881fI2cmE9kv5QHyzaLgfcadF08V96kKKenUc5a3vdON3vl8ynoP
MTUVRNdoefMSWkuA7JR7es2EcYZ5B5yB9MiHVYeI+doS9pEXBvmrTw6KEZ2QNCu5EV5weghUdEPs
NgtaRXOpq/O+HvfI06+vj1Irqor6KzoUCYwm65aPXljNwaS57BTgvYEk8tb+25plQZJWn28UojTH
GylF2aVwF2Onakt7mUqW2uGyv/sm6ghPt4TxFVT1MPySS5OtsRAA3zYZEVh2tyeVozqOjIODSPFr
fhAjsVYrh0BT2NG3M5kfmCZPbAhh6QiCh7frDd/Jp/XR6c90Pe2xaadgiu/kM4RCin9qHjHzw09o
BEMLtPOw62iPp2WoQqr/FR00ZppSciKd4QZzyzaNmYlw/2yTSIiN3kSAxW9y+l1dbbG6wEsUu2U0
nMaMXlnPIJIEBciQiRhKGgsxbUsub3d7oZtS1g+u/s/8JrGsPqy0uJ1ngqSSypPVM3O73U4LgyRS
aVDURUuUicH4ErbyCZlNIPMxCd87D0ye4n4QO09TWP/wZtNY/Lt949tFlKJX8CCMhSLlMbviZPaX
CockBXo2Tw7hK08/HglDY/FL1xXWMrpgE3Tm8shrkcRWkTf+hPy8YUeylWbchbvtSKZfyE4tbPYd
C5zLX4vUjD5Lt+Un6JVUTEPfX7ikw1Ad7+snIlrGnFag7hAHL+UEAb3naUUdEuBtHrXs+bQj8kwQ
O6xTMchIdmVHDmHVg3MGBjtx//I1HAuWa5FdIaPhACTkrl6PmHGt+sGUR/KG/pAn78Ql9GGuwX+T
nYkmwlcQXtfuQAVc5RxlmsUeazI5T+JffGuauD+c8B75cW3Lc/I8gjx60mUAGWJ1DVGjdYuQ6o2j
uvKzNDIaURekzp60l4rJbtHXIzpe6k17WMP4cvyQ2Rs/LII/vIiTFY4OYo89vmzg51Q7r9DcpT/p
d9Y3iIkmHULPpGXQswWK7HsItZ+5VqjUE7neGwRhb+F2Uaf88AayL/sJxkJ+rGG41aPveQ7XnI+9
rUrL7bTPm9N1by/X1iIZXswG2tzvtaY+KJauJk396Rse016UFqmrmy5XP8qwpwWITtlcHkjswA4h
2VEwTQ0IoFVLWYMQh3yKK7TFr7bAGVKSoAf70som8QsVo5z5R1TIeVhia1iL7Pr1I94GaBIVBRan
anI5gqk74cIEqJ99V7stXaxJTIUfbxbqw0sQoqfLa9TIJm+tklNGLoaslH2i7E3ErPYrUdB1vY3y
i56c4LbCsE52rZoakMXZASf3jhfpnDCC3Iyn1yhLX464/WBYdmsBUdaGsAQb7yI37MByO62Z+Grt
fZIG4VF1zSJjKz1e7Y+Mqw0F0jpSfd+5Znw8JB13+1Rgod225iCRX+al93nFBuq8cUeWAtYh2xWR
CC/QMpV8Yo2tNbMM7npSkk1p10aKI+Lw8Tgf5D2T7kwLmZr/9D7oSE1TE5jD54r2U7PL3lWlxGnn
npUHxTlyECC0nUmsvJEoGJ/ZenmY0k3/aPeEa8SNyh8rqIOtwni7hFUWq3Utg6j9w0OHYOte6ILY
ViGfgvzn1ZzL00QxpbDK8aNkH2wymrgeucJ0DCsyK60o00Moj6USaffK9tiCpW9NxDmbkMI1kt1H
WK7fFgZRH8wTC8Qrf3SyGCXPCzmEBjOHy3NMBYrQvs6AteInIai1nJ8McMLhuNeGTzJl/8fOLfmo
lafarjP0fJRnvLTt/euX04GxlkRqnoBL+hq1QI4wMWYXvJzhov349F31c8UF0cBqddC7Blg3IKAv
E/sVN2BZiU/pA4MmZ3qFHuBjWRIUSHDK/EjKno1HnECZbtVQp+Wz3XPq3l2QnAS5Z2K+OooLCZyV
0cFtwVM6mKzRGs+ZMM2MmlrooKjL8xAuqrGuwa8Mz/rPM1mvUep1yXaB+amE7OH1TUsruAcrDXvl
bqpL4/7VCID9xlEln0SgZVwAMmphvS0ripxdRbJNkATV+lvAxwhcJDdRWJG8sHST/G8SUOcJADrL
3H3zFbXTCuMFFGAJK7IZF499QrnXwvLu6PzEcxEsviE8ZRJOZqAh0/mv79mR4Tk/y+l5FN8oNAEQ
cvZ4zz5XKi3eSqP4wJOD8puJn5Tzdrs6iX2DOlVGehy6PywTWlkGrHv9dBYWJL0Nzxn0+JGwLfnE
LbYoKbGNWrEqarAYetdlTPlZpfyuSxnDuouy9nkKq/iIZJB+cECDx6xc34kwwozEK6dYrp0s0AeH
9l+ZB+GkbYQWDEwi5VRKG748+fxVn42FOCS7lXU9lQ4U4LIXTaTrNY3hk2tjUEMWzt7aX8hHUuhJ
IhWcKK0o0clnuQKtkcI4yIympiB/PIanlICIppD7tt/iix+yUujdKbsXX3nhxA/BopNrcrifPC5j
pJ1o3yRhLbl251IcyQVav4h44Bi5td2/Ut1CrAXkz24K8/MTH9uV9KAHRhBaMJwbitbOdNny0dDq
ePxb4Os2sTpAJGBVa0VLhwefTlf9lPAoiVI0Mya9D5DwpF9jltVthw/B+O8t4YUXU8YZCL7xNZe8
IGmx2zjYgS/gC4J5HLMecmVUSpzInFaGmzaj9Wch5IMBiS9udPYtaAqwZv/XSerQ4xuvtHy6HZh6
i+4BbFYgATTaY1EI7pvuU5A/Lvoe3ZJ5hUZdlw6EkxRE8mjhczzSMYTmlFALnnN5rp4k+rjNVALU
A6vd2+QekKM2rAZRNpn9kDWx6nh352g5T6hPR/WrKHIjU5/J7SpsJyo49Ectwa+Nwhm9fWlmmOSb
17VDSOFVcNw3xsH0yw0ArCmybM1S1nLQ1bFo6haYROg+35BMQCMjqmqDXY+7Qd4WQcf1AovK4ntM
giz69Harudp2YtWtRDpioNbB7fkQg5BEP52avztakJEHeii0KFOciqnCUfH3M3z92NyVekGpIg+r
/+ZZNeO8DLihTvs9+2h7/RFf7SngD4HSvxS13Gt8ULGcP4snXkzTfD74uMOUcrdqY3FW7OltU8+D
2fEg1YKebQg7KbgAQRr6kzKNNbIpv1PkRs8S2LDdADKqyswBXzIX83wIEcm0SsPDacc2t4qvXpII
y/2m2Ua/XaBAtmtw1EozSlnQiSmG5ZgTZFSdekEE5nMQlBeoCExMY5ZmpFodD+O4voBpUOMdz5h0
qCIHu7Ar4oO2e31/NEPTC32KJKdAeYWDgndrUosdpjoc7Z72BfOJazwyLHKBc+bZ33qXu2zj4K39
CgxNOHIRx66CvNct5+67Zev0ZtKUkaIr3/NGUaXszLpmz5sMXP557VCO4kwmCC1KQrRU5PsVlv/R
orjcm2wpXrcazl52VKjuFFhvnPK/jxRKZOV+KL5ni03ylJI2DH/SAGsNss4+dTkRbPGUUvgw052l
1/TNg1w6amMN8VxfgnpVTAHzUr1VNlscu1sTNLV45dAZNnm8HHV2AcPtxJtTzxVXnwQ0gBhlHL53
UGg0e4h6SrL9Lcwnja+Y9JEgHVfd7oxcVt4Af1/7ytMBSP82ZFpDQm1MKISRBbe/eyCT06AiWklQ
67BLVuew480COGynT1hDS7jpjxANt5wbvzLmwixKySuengbZwXi/PQ0B5LSOIbwXZP/kvGqHMG+g
1Yqv7yQD8REJ0lRVj5vNPC5wE83rrQ/h/bgF3dy5b8sJGZDR1V1jFP505p0XM/JSoB2RmwtMPO4A
n+INZ6/HASyE8tXRirPJjNHJ4jo8h4oxt5+rRYwlWF1sQlGb9RwuTxZ8qkD+arW8rsE+DFnHfK7I
Roix2njKVXTTIkwgcbglp4xsHja1Y/wlWJBBMy4f4L8y1JVMVX9R3G8kMGMymCmhJZ3QZiReKG6B
lyGa6HIyCpQmRVbgYALkoPjMsAOW5dMTyYPynZexhSzaCnL/Wh4BGfNjqIZlnO7ic4nomE8CC8AH
dVn2X+lMNuQ/CSAOWsj/O/24ZFTYs82iZ+57N9eS4f8jiyM656RJ4I9iWa4tUeohl+2HqRAk3uRC
IKLu46nIMYEOMh2DCrv3pwgC5V3Tj8WGbkK+WOxTQDkJMQL+UbDaAjTgMhmq41UniYchAWaEymFp
hjv7rJm5efgTUBWJnqe+rBLlHvRyQhE6xwv2t9z95nXH11TCcMywD2W9G62WbFTOoP7dpTrP3p8u
ORsGhjrFFXbF0j/EMBgOCxqv2jsu52tmaIVj2HP8c0Gn6Jl/fnaTwyphDyZXG1BHmB8MgH/ABuVT
ouh7EhhgN91PqTwYPWfK9hB4lgRZqL+a2A0mnop2ia5eiM0dXKPvjJQi/hE9IgZFaV82RzaoHvxb
Er+ae1Jj46gq4dMurqWN5+Ru632nAGSP8fQzWN1dFeLggh3wlbg1b9ACtfVb0fNh03OLSydnc57L
dNSkb/eB8DymXuFGzbYnmKx5DdzzHgZWGgPG2Hg7St14XK4dwfBJVO/1OAThJu4r9fTTAY/XcMQo
EQX96fjbj/F3RAx5c4/4bFCw28mYQKnODp0/966jo8ZFiLYGTaD8g9QhsJzfe50fdNFHiwTWBzDn
7PBC7baQ3hhSQcwdXIh8CKumJ4qt8CcPCza3Cw2zEQ5lW0tqh9ygbwZLF4IS64wShxW5x2bXtv2C
pz5FHGK4uFuUibZPg/O2m/qLpKVZqz4YDJUW8NrFIhktZR5cQrZxNCNXb0+8vSoxcLF2hrSP3LUI
khpae97G5W2jMnH+gPfLkkJgARneoeKmC5UmoefQXRu1LrWUW5JS0Ti73Iiy8FSO9PdxdeSL9KQE
m/lkBK2jX/tmhEvbKsK2oVDw6jz6jnK3HhRGbqVeUWJ+CCyuICoH9cpVhukauAj6QE51e9bTY4ZK
kQKA7leMZsxzMadLOhSU2LdBcyrjEpzt4oRIfjY831ceEv9Zu8BsvCyxaZwMScf0P21g8HkqHFfb
aUS0RMVg9a/uHGfLHZzgGpuYdcLESiHccOmxr0Uu5eUe+Y5OVVtQ7VRF5RBRrIqnKxQXqJB8NZ8H
ZBRerXGNrP4iDi45j9vXyVHTmhzjy2b0oYW/5vA/zdyBr3+kdHipXxY7ZuTNvdeG5Y5a1KhuPPTX
cz9UXmQASQVNUbGkOFEvUe6RaC7pTa/YWk9eHQ7BFy7Wo2xmuy/QkvhqHDkTJFdOYHRKWm6etcCm
BTy4bXKRASDUGpBBVmIaYC3i0HnCCG9MOHbHyPGqbHtnF54g/sfKSlys2KX/s1tKTZ3AKt8hv+nT
SmVyUXsmXB8OaOJQb/V8fWeOChF/hMG2zy0XOJivCJiJYdNJe8DNlwX6acMJhIgsD+48wlOK9oJ6
OEgcsUcRJeBadJQUMp7oIzmNw/c3vLtY6EHlhXox9tPFDfqcOhkT4GoUrKuwclNaF4KG6PhHM/RW
aZeslW/pzZBzfJrismit2A6WbTWfg3LQGg+2Tzgh/2TYKYTPfB6TNfok0aMewU+xE9PaswMTbNam
BkdKWxSVQmB0nw4rHbgF4+Ftm5tfi4DH2FEuqD6fc2HKYe4zwkMgOQi3HoYwu/E+KvDWz/P/60k9
4VkxxWbRwmZQi7EK0ZlnCp7Qv7QMmkQCilZ2gK6TMTyGDe0bSUdkUKid1TqipVnC2c3jj3r9YMQ5
+lsZ6cQV+hI10ZbbroB1kEjEq49JhkCuXXZWLDcw80DVuAjPbZ+SnRzv/w5gD+RfJfpzZWICYHIj
K8XaN9ElOyeNe6q5MC/eqQJmQFJbNvWfrqklFGeQRT6kb3eSuYo5kZ31/WU45dTElKt6ceHKucjM
EiUg/5vPzToXngfqTYkHDb99L2SW3H7Gf5djrer+KFUOKhp8rFsh5w2jqp/CftEOoznQKlXhR4m3
apGioJCiy9bDiVhEUCbj+T7tJMelIxGy7tiPOfXNEShM3PJ/SlMEVOeJklsIWIBOMurHHUbX4dNO
94skwhFkBLMsGOALUOOWRdD1Xv83+RrmF6F2gt7msJEzaZ3jGMc7ZrRhXB87GvrE+Ql9v+aapOck
M38aoQ3ovqjTdRzFwfHLgdi0RwjDBXqw2wLW7jjHaw98rySXVUEv9Asr6eImvbbDGJnz4+695eDS
3AYh0JFCCKD6XBCBTk9/bhugE8BPa7vELSvzSfAxVp+jRKflc8GhBX0qHE03pVR5PZiHXf2gmr/O
PDzwe/1ekRVWpt7XUO6M3M9Ht4fyvTMx7D/108/lw8iNf/YCmjohiHmDZmtVgGBnPnBUzvQSKItf
4gSR3j4e5/7i9cRBDYjB3IOT1+bmgBl8OR4e0VmSrlqk7Qh0GuJNQKVxOPE0J4Ccq2TlRKgZ55V1
DBL4UOPBs9L0Z3Zi9cGKgFi5o8XnvyqTF3lpSsemBCfm/GR3CeQKVEY+Ta8RbnazfdeaEnNgQG+h
wR2sv0uFRxt/LmvO5vhBNV/ISFDMw7lKxzxB9ENIZWVM4pVsgsHYd1tkGaxaD+KzT+juvr/7ICwm
N9hruQVQRRq5rXobjo5wA0g2j0P/W8nClWgz7atwMlp7b8Nb7ZwF6bpDke9KZ51GkyFdMbL5hZiN
U5qfIC8xsyW/IS3/Vt8hY94vbyk13xUGAap8A81O5RSd20bN3DoQl92B+Yb0liH0cvUigdCD/Lsu
ky770WhpSU4HI3XbMFPjpAPRKfyvy1MzG7D0uZ9zsnHJfP0WuE6g4lN3HSAspjPooGBmMteIESvt
mvuDFCRLmMc5NDHzvGLmj5TMUUS/xNa4WcSjJiOp7KR/5aY5WtQpfZvVoLDcc7KLK2ttH0HI6/Hg
90zX1AiwWt9dhRmRZMWTxbs40Dvy1QXwd6J25bl6pEUWzqdWOL2JJNAoiCgMh1kx2fs890bpOF52
CRLvv7z1B3TwaeEpsWeNQRRitUQ/mwciJ7KCPiHkyv6fodiyrN6JGcbMI/O+l/S/MhI/S4gylGi3
GNDya2/3xcxZx55mLG84AGQamwWbtZrPRl2XlKcNyfhLrPunwEuGzCxAIpcLxqYykkDMDN2fJKXT
EpdpFQDzGoiPu+Prj9pIWexUHY/6bohWunqwnxnpdkc6eSni9+wAS5TDwVS8lMHiP8In9y6Mb/7e
Y4C5XRuSvSRPSiXjbHgz6U6FlollMy1TFsVKfzteikKKr3Tdt+Fzp5GxFssxBGGKI96Ja6hrdEfv
ECslU/BkzkEHYGZgd4C5c7F63GHmwVmu5TuLsPb9um+f2V6Aa7I3y46uJw1uIGbSYdKrrxEPUdx+
tJB8uWgtv8NsgCo8GHMhXrwvvOJd88ySujXqu4eSrX5ceUzrt7sYmYgfdxgX1x9IZQF066I1nsve
aPwhid2+qnafnjXvUIrgN+QNnY6TZpexG8/+epkgUrVLIIEritfVxKBne80fmGPMAZIsafdf0Sb2
eHF0f6Rvme1BZpCvRJ8Eqy/BgGrl+Wv3Wdac9VHZdSuFWGFVc/Z9iAuHii6mlBRDjokrSh+on2o0
oCTCIXdkcbk4t9UP3vbSZh6RCLcavwU+uRipAcTlil+KEXrdIyGuUKkmejSKkGGCK6KhJfY74GrI
zmZKQ6vprcQ0JfZq+TM7+JwQ26Cix97BjoTSU80bPy3DzVB7JKm2YyM/kx7ZpW2xPnYzD9BKHpfj
kTBwI80sMIQcys2HriSLofndrgDtitDfJMTjoFqfxG74b+UwrVC9VWXgO0T4waJ6mz4cQ4uVeWoj
xxr/OUJUK8EAwvIyN0OYviHxOZs7jDcST5IIctQy9xg0sAD7PFPRRNc6KI5OJM68vmi5nDwJQCUt
K8Ay2PAteCJrvcyh73sx3swVl5THZ3IQuf8WsGEZm+ri+w58vWiT1lMYZ1SPmL9Q4IH9Yc4sNIxv
ibDxEmq8AxQ8jkKvDhYIS51vXgFmDHT9XEVM9itqwOx5QYCWAHVGWEjR6Z9y0101uiSAupmkELZA
repwnIJx9xNLRhVxjJtQ1V3O/MA+tc6gJIUYkKIcaG9/sZ4EMfDZBrdEJvnv0vVJ4C8demL+bWhU
dN3C9ZNEQDOC7C3/HbzJQiN8zq05mZ5BO1OR5oWsGU3HKbP1sbIee71T50o56xueEp0GSEYV/EYK
7T7xydouNs4nccTkHFwzUsNkzKDmdi0Pe52aGg18Dk97mlTbNG8wau5L4d5XyC6A+XVt3sTjhJtg
XcbLqVR5q+zg9uvGUHobWP2fSvJZy+ye7wzpN7UmwzUxQxGLlmKxo/OJ6hXSIBCbSiAXOzfE+wHn
rZExA7vk7ZHtf+0vRUKNF4nhDcZ2Ku096S1a05Fiv6vKvO/1O8iXHNdE3aAzUlzjadu9rMJfStLo
29Q/jQY7CYcy9KJuhQN3jOjo1KOoM1u4glENx6jBuuc7q2LS2E9W3UlxReCWgvJZFa4owTacsJem
KcTmOS9BkwoajKF1ZRQS9w+adlmpS9XTtjXlRQ++4Es84lXxYGwoI3RB4hKZm7k09aMy6CIVXKpq
26eGmSTS7uP+DpoRVOapHfo3tw5ReV+C8Zui05i4SME6iYL9xrYqu48DTYkEYZhOFU47eyHuTRU9
86XWASCyqYc9cry/s/4MLtVo+GhyFoHI8WDppNMf7/bKEEo4DqIDxLr5fosx4UwbmHDjb/7SiegZ
DNh6PIM6ZNiWcH6OfSmkMHT++k2LeECpYBT413c7/qQxNia4iFh9tMDVRf0pmhhkBZuGgSOA1Yb5
dNWxEHHZZmv1QAQYitKvIHIpP/pEFv7Yo4bEkUDtPCSTNyYYUaZpM7+GdNLMmpwEJ5OD3ev3w2zn
Pcqg7h9vgEyUwDBBlOU4VtdG/1xF/hBvRXrgFDE3WP83ES9L4973IKhZ6Slx8DNci0D+jgCcnnCZ
ErJizw0mjGyM1UR8WRIN6+XNRylFmNATadJ9NSwYXpdsfxp03y857jkt3wjfx5mIBJQkNGW+Apnf
kdRVSldRV1ZxSk65FVGl8zH/5Vqo/9Icx8aj71/BKA9/B32tlYicdNhUHeox8b7o3CTUf9l0VHMY
f7SGem07kuJGtMmUm4TYeLAj1lZp+4lqpKnopQq+o04mODj4vT7oQ3QZovL1N6aR2NU0MzYzaen5
49bVqKxL1hzWAO2atHJpz6TvgsP+YTPBOIE0C4hr+msKc/yPj0NheeG/7tLpqhKLD9fUMy0K5qzJ
mcug/RVchPEyKxWh3WYXqaIpYUH0lzM+TJ50Aq9vWD2ey5moZF7wXcCp82v+JYzZzmWyDOGNvjJa
nfdC+NuVDiJKHpgCpUJYiV6Kei1PEBXIe5YSWQITtPAH42j9osoi1dS7SRkhRxmcHOIDXzn48zBc
3riobWgx8jTlRyghqEchiYDoSfp9krL5Qc/1WJ8vmmzMaEGIyRBEVFS5KYqwCUOoJO4pmqSpHSUR
8VrmwQTsKHBkhUM/BTyXIN5LyfPkXxa34MUK87lo9x42gZEMXskGtwiMJrHBC5nNhm2YiCdTg7eu
qo825hkfIWnn5vskLEq9+wd0vxHeRaoqLc6LDgMN8mwiEjttp6OjL/4u1keKsj9L7Ja6yX1fYLnh
+1zbnristMsG5MPM+YoPkkC109iulEAlvW7bb6wLEQvkiE1ZakmwjQIbQi1ejUw0vsrrGAnM0Q/7
ZRsk35L6IDOnXbscZ0V7SiIiw7kDiXyaQbFOYc2AjnJ3lLu8n5rs6D9/BpZnYU6IOdt2vajC4Thl
+S4umim2BePmR7xifbYEJBBxkZm3HXiFoV+AvGoKt76YfTtfjQNkmvzDZGR6vKZrNramNnU+gznK
GRw3dIfFAFtRORkmo9Br+RXVMVAyQmmBeYJPzA4b66yuKfNbESsh31k03QwbB0+oQSe4SsxcHlYf
w27c6Y8Z8FT0YeA8U9e3RJP5Evl2XPmjLte28h/VaLmXakLyYJV2tVB93pU5kbcuXJ5kOXJshbKw
z4rji5C9DrYd/ptn8atJBfDw0UAT3F7v4iBevcCG69ffDnEgug2ls5KEBamz1JO/Fmix6/t/zTFp
5WkG7HpeQqAgZfG2CVOcxv02Sl4Mogkv+lERdXKoNcUorPn5/Md+7wM4mAb9WbY6NE/Z/bueu+84
gkSmj/xZE6nabVRtgLm8Zjd3+OVNmKfOYTA0ZZZ19tEcwo0zTCJIj1nc0yIvoByo/lliaB0UJMsA
Nq/odhrjxYpjljz+jtHBjGCC+YXYL9TyOSuRP23sTtbgYJHFqTAo2Q7YVCycH4ZyrCWfilYJF67W
4srodxAbZPoNP5JLbkDRyIFBAkjtqwY5tlN/m2zW0GakPScGjEyC3IUqZhEs0SMfntXPnioMN416
siaxQc5lB3CP6gOo0ahvpiBVY3FMSx9QT9kRfHdEKiS/ZsYVZ00oEL05uRX+i2rGs0MvZQ4TDymt
jstA48VluskqE9Z5e2lYFyzP/+b5eH/vsTzHa51BKXk6hTax+odgq97yRF0aOt2sFUVsIy486u4o
GLTrbSfWx1XxvO3V4rcr+gbGJoLxrgkIXQEZWw0jRWAzyd24TfpXAz+p2BfuOdSMzIbrVKM/WFGL
5X5P8p97v7u1BaYPvuS65ZDznVO9S9GYAULZOhNrToXWKw4T+xh9nBX828iDBSzrGP2qa3XtaE3+
W4SSuc1Alny7+QBaBAgAPCUNXMl2JBq1YwJMclOdmmuUiuNkqNyWCToCUhjZklaafLMncG7aZ7gY
J3gcfW1BYqxYkn3lTWSobIoqfTpG8BkSgTTGE+edLBWrsUheubFp33SKEdK1p7kYMa0IC9dhMweo
QAtFsiN2GM+g3JNGfAX1dvFkWP5W/Y3LjccEsrV25GkdTo6Ckz+KD6B04aFT9Ov7M79veuxu9k2Y
nYiP2JFAWpCQFzZgMqav7Vj7QuZm11UNABE/3aShVj+gHUwmTumA551P/FmY7ulnRaJ7SbT1VlPY
pb6wpHbA8IMyTxCiir/rttW+oWaab/Gq3omedCWrajW8OAjRM5hT6zQkv1bFuMiZ6DkpnNqAdx3W
Le/ORRCMiTauprIi8pLuClLCO9+agA0GCQviKjMo2DNCQPbHUpcQ9gNylysdEDpVV43EvxVh8i1x
kjfMTmvBbmvtuym2BOWp7u+pcUkzZBGYeTkSuIsV5GRzwJLbcKjRWK4PBSlpkcX+BFILF9X3k8at
xPdAVEVna2nSxSzFjSu8d/NY2PSAinawp4unDP1QhaZTGqYpb5nWWak+oP6EI3s10MKcZpP8wAxA
C3oKr2SN0RZNCy59PnQOzcYeHqUEVyMeARlhzaNlrlLr1zr6rNPUj7HmY3+5HxPAxJ2lrPQVMWUd
IBCVZBYQ5PJqeWe+bapt+8tJXHqD0i+rcTVmc7TeHBWVVnU9DJYmYr6t1kEj2yiJpj1rmWmNQs8K
bJm9lPA9TGuWClZZQL50dWrttUa8UUHxFbsmXOdhGzuh2bH3KwtkpSGgUdnP4CReS4qPXZts87HN
U05Fnc8x80lLg4uO80rqMS0AG9C+P5nfo9ujYQa/4HvoMA2rF0GXO5QqOrBKDOGL/elNSYgHucf2
+NjXWl/zoswDRSTVyc+EIjoC02Aadu5H4QX2bg3I0olIKSHWp9FrluMNwu7+bl/OdPH3LpyejKdC
k3ppbF4upUn/CMPfIHTpEudi70OwwTX0OEIlgwqnqXLzcPeKFu4Wo2iZuZXQiI3w5OirUnET0h37
g5g6XIY9CjpK9iEbltfpKOc+TIbLlss+NWUCMa0HUNSqTxR5e/jNLkBL/czKYqBrkAGh9Dq2VnE5
tT1lNOxT8018sMUx4JGSWVnIRRI3NL1wB8N2/Zkpx/RPa+U4J+sLIIcYVdk2mGySBKHpZknWhol9
gkCofHz1gQp3Qpyvbbhv6LwrMw78tXvI5//ufAPg9YbXypu26GOBjSaHdN9sYDM9/CzJSdAWeCh9
MBX+0oH6SUeOXpdLWj1/or6Ed5bO1FZ3AuEFjz4QxNSJuynq0C+dEVN87S8ZXkA97JPxUwRajuRT
+b/6MB+W3+/sGIEuhpXx1UJBfVdeviCZIJEi+RycdDtXJJA8+ydLHAR2r687xKgDVPzDMeYQk3dF
rNNqq3nC3kA9ewYaL7SH+ut2va0FHrS8g75z+tNPYZwNQvhpVQQelTtVBMddPzCciXUun7kMPxLM
WYBDQnz2iFhKh4SVWcfS/MQV+o7rOx4bkp4jqTVzsJ1uW81PI7K2SQBJEcxA9fbTkQrnefNR36X/
MJEYpbaCArg/MduMMoVUGx9EXaTm1FigIGKIRSArwSELVXreXdkOdHG6/wZrJmmz/jIVy1B14skV
wZUZvSZSLuWAIhwjiO4UmYfrHtIVg7acNJpOo4SvtnVhuc4eu8sPAXXeIuiYIFAPsvedcLvN0Izq
YI8FITqZ8nSEAHnglnIu6u2x3LZ1c1IfcvVstFTHEhJeLw3sWLBohELNrkn2zXek0DMvxWyriD3r
DNoQbKmHOnqu4XV2GDIE16lTO8a7aWXWxf4dM5DDTmKTKUfg+vbkx/dM0QpJzOz5P+Mfvr8o2LxB
ymLV3lkEIkmGnkITDpXAtus+7aUBQucbxFd+4fFFTndocnpxs2pOAbW30P5Twik+VEzBEe0fg30v
TX1sEGgTdtHKG32bOZYjuA12UVQf69wqznnBEx3xbsg1UGYHKrQgIpxffYsQbXdubTPO+rLIsUNY
AVrQRTJPYM1vwVxXVqIxKpGzJWkjIm5dAwLogNs7at1s7xdlAHvLSlNgtas+/TeVclK1jp2U50Af
HtkTyyvulR183LjN7iMZ0kHZroyv+kFJNTxAlpOIH+FECnX0Uy6ALoSwz+cAQADKvywc/Ub78u/r
6urZKxUalV60khKMt4JGU9TXFzxx9LHbgV2ZTvDeTFSkhGpTDevwISI58Q3RcHclqub3lo4G8bQm
NrCvk3yxlcYIY33J9DUyX60iJLcF1+wYEkYVmRz6wFMjGAoaDe7ALbsenST2zSStwGx01mfgvBLm
x4FGAmVVVs8W4z/XdYtX9Agn65KW2ypj5FfbTAIlvwFk7tO41Tay6iHpmlZnKAsWjsGGqRKkxeGU
VC0DiERb7/hP7li5vuDJcVD/5x0QdkAZVMQhzDaNanFaMvVm8wc1BG/JTO6N3X9P50omXAULsMFe
zJExzfQImUSjjxa1FF+L119QreFVZb4hyeNi1fFeVTs1T25iPSTWqmml6peyJKRNOhM/3B3TGEWV
OEl05m3jjnBvyGtYJjdVI9/q1GfNkZXkqpNG/VmUvlRSl9YnYDGsXf3+EC1mSmQvs/LTRwNiZ7hC
IcC6Ajq4RfCgGFY0+hYRlq3sMpuRp02fvdlHWU/SuBw32sKAeuRKY7ypu2ZZdL45aV0UcG0rUS88
xTWunAX9tB+NWcih6xU+4QNbkTMWGjhktT2x12vMEIlP2/K8wxK5isnAVATZ04o7bFkg5vaE/aAn
Y85/mrnqT4XCYEQP6+EP1BPqCv2MpktNAkCHmtlfiHNxQGf7Xp117mCSqMdnSg3JRKw1hPfjiluR
FXwXnX0mVYeXVl6blfEadiJ+xN5Y1A3JsRnpE1hzyei56NTPVtUEiI6ROnsm+yzWoczDOwBgHd+U
UNOUbLDJu2YfEDtMzrDpiuO2OuoP8/JxND5UREr5vUm9Usla0MoyRm/HGRtG0xQ3XVAD4P6iZR3A
uH1ktioKLiws0UnuYKV/0WQT8CE4JiJMi+Qm1qxrs73AimeD7VQHqczrD8EcnThuOEYtj3y0/ZUW
hfzDZO1lS4Y2jNxY+k01wiepfNygPur+/v/+3yuK9sZ2i0q9HRNPsG11QE38txQMKwkKCQcApAqU
PLRdK6uqzhz/utZC3fHI8kzM7JPXIN8lfGqnBhTuFqIkhYSP4ww/SVp2bMTKZcvjJGKnihn+ht1w
HwFrLc96r/gYbxCLbbhVjS4lRv/RZU42NYNMLXrJB5p4iOLfdkC2vAkW1AGcZztUrS9nkRQRB8/A
Fw+sjISQV8jDpFrHB2UfJbNuK6h7UaIUIe/7v0KQhduzccLhOq7AB0BiM1E1W6bT4B58PMXCRrpC
jMSZFYiC5l7kIH89lMDSoeHnNFlULRM8f3skP70VHfP1OGcmsqLWvnXZUF7vsWh6TTswcDI14nmS
9dfmLCwmqap09Ws0KZpTj6k96o/MXbwHrJsVl278XeWRUcxqGC4UYOWahcEeoBHWopX/A7dFzL8m
X5gMXeVhfJUYzmRvoFVhqt+xj/br0yeBY4PAcV0tGqVwaKwvPhaRq6VyBl6QNyJ8VrS4ZokRx725
aRWtQe8Iaq7q7clSKwt8ZF1hX/IAfCOXPLrVyA5xMSpRk5QsCzxRf7h/VRawR3QxviFbFqfdO+Kq
n9ljuBSbkTTv6Z9yVCiECdal9iyrBAXGwuspCPPPXrWonc1LsZjz69uZr64GjmNcVCjYk6jNwHlk
AKQdi0AtTu+/qaLg3pQ4DrGOA+NTro6QBQIuRW7Uv7QQUYlNnDs4IpL2VwpalwYzKvn0DrkxD+Rh
wAhVmpbIZKy2XBlbAfGmYQOdzT6SvkdrRfz18QhMWLfqEEtkioPZwy8ArNucpEm9AiFFaivBFekl
AYhusZQrADfPZzxreiRNSchiUAw+bNKPhvj5/QpjK/pBkVflwboVoCkaMd9rM+U6eQaqAZRYq8W3
4APWSrOqIBoINnMyTZmNj4QfI75glkRD5ZZsyuGjpA8hOdjIaIHEEbMJM2UrR5rngXGYlWV/KpLf
iAZyJgOzegqilmp3Of3J8xNsQYVc8iYPBDpHmhUm4gTgDJSmq1VnN+CaQ07WKO909W3iBISuIkpJ
XsQ/7B+/5IObxbqerE7peP0khmrmMfP5J8vXYw6Sowi2Gkyf0xXqLdH3W7jPGy5FDZbar+oVybb0
yQJKhHOCt7fLDBPkyGcA+0UHbMP+jBZEp67TZJQpiomjrXKApJc8GrpiTl1RaKwi0H6ulLix2cmy
FBL+s94hx6JVbCs/Dx/6nmKRZgA2j+K5b/+kCzGwum3H398bJsdqUSywL9ZcHXLwd6136ScX7vjJ
eViJ1V4NY0dkOozJyNYLrK0/sNvva2gW5F93vsv/XLMa9bl/sC5ezW9PX7nyyDbzrDKXiN2AShP/
ZGK+zH2+h3D5uWP/Lm/XSSVqkCg/5hL1+maBfiNHzCG2OXy+zgH0vWOgkTxY9dNDG1c5r1DfQYQ/
Kl5s+L5VDbcJmvSvD7uwqsHuitzrgFbIJghp8zkb8UIs5ZHsjkhXAQsjPAK6uJ0oYd3gLl5q8aYs
ty7JrDWdL9vLpAC3LehIbV+h5QOCMp4VXHLYfD7NyqdaWzLQfRHjJ0F/kgQ/9MnWuPemRS6aLpHs
lJKkJfkHj7FFPL4O+DAJqJhoO+sgyArN4RPOu3IaPEdQLS7QJijPmB7HCJZDBKFWQp+Z0qvesa32
Q+NV3zohZV453OYfbHbYCMhaavnA5C209x857u0JPdDZVpA6T3uFkMYswHekIUQ9vY3jtzsN0ufw
FSk6vGuFjQCuLFRg8ya3cIQr9z6YqIkLGAcYWs3qqCmQCZFs1HUE55UWd9SZ/VOp/zemMPhu8RHE
YHARWv8qsSad63jvXpJbKgc84oyyK20N5cyzlqZyTqvld5BoFoujT22jaSbTypU8h/MKWaj8ComT
QRxXD1+IAU3PKiTx1pw27MQO/tZ/q4keBlHgitR1x5C37a3D+zBjiDeV2LazXHscRVFEVLLTkgHN
vvcyYhmZlf5B+BWph8NhPIGQQfd5dMwKbVQdJ7ftAWNEL4+hc1RZK+gPB27kN/qFvA3tMpvZSWRk
VNdr+dB95hT+gCkDbYX4sCdCwde2L6tOPc8Cz+Dwk7x5g1sipHZKSjFDUMgFhIV1Z35OfZIqWKKN
0ZUgZWuvoRLTZ9/XHBX/fqD1ZEMMuupYQ8llDVYbwLudc+rJlnAAIDK5YIgJlEs49O0yVAmBYbkw
I4ND7geEFNr/wniI+51JiYQ5PbAKR76WQjXtKnneBXJ1WxlwS1eBpQVQ90f0IdMBxpaHrw8EcYG/
sL2rVpgH1Cha56NuJ0pB2rjkCOCRWh8PllEyntvxGBO7N0Q3tK882RFq3FMSDoIZnuvGnTsXjyZe
3N1Cwmwb2pUH0vnXYSfO1j/ik9eEfRs+rbh3YjjVtpYjZgvJyox7oCUsEBbjW2uk45byvXxc5M68
10ZiqUqnVJS1BcrtAFILRLibkLL7TQvD2+Lr+pRoYBr6lyKqPxmKhWqO0/IMrJpoiYR5u36fvfey
J2hg10N5mEnYpV26YWQtWfkSPqloiJITs+ZCfNh0FVaum6J8buGYeIE8fWE29+qczHKYTXT3r2r/
YdjouycQ7wsfjqLLIF+opmbbSIDUBNXfQQbKhjMUtpDETUiwvx3f6y29Do63RkHfmPgbkRuvlHZc
MlEbDptAX+0UV6u+JoIMts1fkV5rKqQ+bK0Q6zxD/0UR9oK20NADt5M0u6vurwoRZMZtN797OaZk
R0gsi1BChUKtdLPmGvQwJY6Rq2dx3ComA8xvOYKtc4LFM+5Fdhm4+rn7LLHhYQex4/gg7PGW/TVf
ldL4wu3vC5ViqI+lihBD4BItZlWXAAf8BkuBR7jnRm7lhjPMs+y2yGgyZA34/fU+N2Wj8HO5oE24
nQIFBOzImLOeQp/M3N8w6Ntl8jQqkZEpp5lYZ00Bj88yYQ+IJOefSMPJWERRJ/ifU1ou1yx86ONL
pI9KNAxDR5MZUZrDAYoKW1XuTQ04BzdqzuY5Ym0VnBShmXcGith1NYpU5x3x6+XgeoLHH/1SgQDp
OPY6BN0nIqgzB5HQMAXF/2jY+YG1d61CH5VTz65P6dPZ2VL5QP3vNrbiXIYq5HBZ/BdJ9x0H9DSo
JCo1HINIcjj8EUFuYjwzW6aOpXC4J/7oHoBF70/Pe+S/zm6naeQXs5x8FND/4AZM64AEZZ7phHVi
e8vrgft6VMEG8MOpwNIiYPJVx+MDNM10GALJBmOO7to/w/LVDZczvaPoEALwDCGd6Zfn5c4uGQ6c
yGmJo3RgH0XHoXObi1LxZt4bxsv/z3AqWAKl7mM6GWQt4CGLpiamKHFokNcdOV1rgcVotm5Ui3q9
5y3yrLB/jCExNcq3Ux2y6/NhsREJ5Vu/PPzn1j/WKiORvC+U7V5U0AWDzaFJHh5UHdiv2mp1JNnd
uTZ1YvrN84ECvYtMpaV0rpavlOGIasE/BZQ7xFQjWpVceupUpcLeCbf5KH7W6tLOxr6+gymtrZsU
GJ/Q/vmSxnBabs2oZZ0QYk19HF1C7EdK9o+zwNYFfE6q9RpvagAsJAC8Azynqw/6uXDIHnLGOYYk
zaur0LNpExkLtbTsoVKLCmpguxARTpaYREppPwFhgmKhyyWj5Aub6PEP3IQEmDIAS/NLeja+UwBm
ed6e0h9iyKHwiEmKRWA3w7zVa8oWwrXCRNlUpQ68cufLIgWxaC5d28IWDIniNI67rar0fkHiYHYK
Gs1eXJy17GWaQyxvpRrcxmC5Ms7a2SpCn/hKJkPIVGDQoIhYELiUS1QkUPJJC1YxwOngNvgvRZQB
NRXM6ICZtUINNZssvNKsnFAxlOfZYw3uJxyrxoeSt2KZ+5BHKDID14bvxthbYBVDmheYFxcka5k0
8Tv3BJDcZjzWVZSUN1WFZvUwVrxebiZZuYNw0chzBDf3St2h8gmvzMu3Y2YjxD1mrPTKUSlnrDj/
o9CVlrBG7B7jbEwlf54nXXUmvZAWXlSiBa6fz83lsujQkL4qibdq8Eyh6oDFf01IOHs6UNcbVaGU
v8YDDkLVbbnTjqMW9IhIbE9AO2xNyuzoWn0sJTwXNGziali65lQAewD7YwjgfkSpWa/b9BON9n4l
v/bU2INE4cQldn5FGtA+efaT2MIdOxvX9xnVi+Iwg2ykQEmHeiU9t0sOQ8wp71kVJ9o5nNCWh5Kj
jrj2z9+YfOroHow+R+mGP0UDDGu+c/kqC7ZvwTblLOdZOyTxKT9H8hHjG2tLc3Q5bZq7G00C117w
VFzlgTsb9RreywLKD2AFSA6qZvQqItUtJ4LdVGY6CO8eWYzd93mabr82hwfXs9nruGuw61waNPVD
umIgjrYAdYXZVMoQYpMJYrbKO44SXnIO5td7MfBtkkw9b5EMQiLkQyvzkQXNeBVUtt4U9IGXG0Rw
oU2Zxw6CMgvDb0fIQ7TFTOjNXl2/GuU9cTOzN1+KSDgK0AT5QimiHQeKECIrXlmP0MVqJ09fucB4
5CLEndRtiqS61BuvFgT7jRBlW+pCiDmNl+OaXScGnvFCojw82HPE8na/T6A2SImH251gXX7SEl9o
HfQg4G1tPQHMzTmFmlSDrquLXTUbZSQa1v3NufwKdGh4cQWkd7uG3VecBrrOiXZCY4qtFdKM+fn8
NfUOrVurN6ZjPQUjEcwzfgWoxqAMy5BTTk4YAOe83WAjnGDmuv7p9auZ1ElGHAkiqR+pejH/A9Aj
5Y1t2BiCDHYT3Zhpi3p3Xlm3DM8ldx3JjISnghtQZcbdNKj/TZgJc1bWI/G8RNNT5bQTrVkCMyw+
TA4pLAeFhVsB2Et2XStMvgpAwiK8AYNB9ZZjEuvtaI4Bt0xU0avjealqJoC/GLADxo8lhj5TUsOZ
bzsZbAvDbj2SY6rruw2MIlGKWbH29F9oRT2MiXkeJzjcUnTjJ0OYUCPjVY9YESkbqcLW3K8fMp0s
IiquYxnqbxkdn5VgipgZRGcBMR0V26JX1aSPmjewitfxzBnR4X+mVmleszYe5ghdjtXXys1I9mf9
ehQuLalBdtgjpp8s59O6XSXfwQ390GFAmlqBM0zJmMs/QaONPI+Xc5Z9MfFLhbYl1PQV6YPQXrPU
lzebDj35iObyaIwuduPQ05SJWsM0RkkRSFwhp3HEQPKgBkfdxcbjO5B3Ay4OkV4jzIUY7NKYhnWd
9t9yibIT0mSOS16gLp5RPvbTpcp/riR9aohoJjQL/6+RDC7UP15G6xvmC4YMZR5+Jqc/GHFvMIw1
+YqlqofAmp9+enJ2NkZKtK85GX5j7t9IWp/FVsUWshoAzFd7/i2q245v3+WXKCOjjBeFYZXaSiZ3
HJBjhklI5IXvEXpdtoS4fSAchqbecWxXYlf4bAFQkXMzor9zeV5N59y7Yt/6+NLOe3CYj1uhpHvP
EgSLfqbrSdFDHeb0fGvrI1amQ+kdMg9EO3dQASHcmZcbxuo3hHUci7p1LmhjikfKe4gs7QQxS183
1MYVI9RqFxZdRV6ngebeOTH31qjI9rY6tSA8rCmB6G4uVJegaD6Gx1wuX2RI/u/qYRFP+4bS8Mgx
NAYmWQN+1qiQb0aiBwzCxR+Tm7itIxV7BUUp6myDGi2a4woBkMXvxrm30J3mqnwPiz368josTqKx
3QgM60H6VS1we7X1xj82hM9aoRtDZ2HTpz+jFvhhobzKStJFJISrUqKMHhPmFLRwIIYky8ZCsW6n
fMw2BlW6RLzcenUPZs1Gh+xtxPriLF0GWdRcuO2TeV99XT4TeSlxeGeS94BnBmadOsy0AaPkmBcy
wh5jpWTa6xTtlsK2iCTNZCSkvWxTXY1rFSgYaz9j70DyuYNlQ3ZmtysA7W/ntLa2wNBVdEDxd7Mj
gKiy+CZ6muv1G8rinOgZ+95MtkBgBNiEOJ6i88ynftJ+MWNQP/JSkLlmqIlAhktzVsyPydqn5/sO
i8lLaVEUlyZEuwWUORjosNG+P6Tq6+wa8xOd/ouqcow2ANtMUHApAs0sCfut2vMdYK8tf93Dc8kZ
dIHUp5rnbx9L1Pfonadw89XGL3vK0mzCtWzCluP0eQAzSywI+1dk3mFCGzyRerPpHXtx8G9yWi+0
mkq9yjLmfB7o98R3DOTq9Ir94m4jqHDjXDPx3FbdY0PK9ySffxDxYGtU+9ttJvapT4dM4zO1yhe0
ADw1bDIbMWcC6COGEjNrcNVydVv+tJE81H3vJqeQcxwthUR+wn5nIbD4xfIgacocQb7/Y78W3Qfe
10m9HcPdqGmuqw3VIluOQlE1kHOJhEzH30Yt9ItRSojeallFOKVYgTvLRbWZ0cpft/8qgsF7p7H6
pA9oexB8ulpcMmMD854fWICT5hBPeFeafw/w7+VHChemS15Zb6MDWWSJemVMSv1fTQ28lQw2WrIz
xoKMNKpHrVbAS/00PpIVCjeJukiV0Jwq0hRF7I3+O4D6AHJMjsI9K2aLMa0UwvlCetMa8egi7rXp
+Hggoq4w4DGo0UOjx/MhZWdlUvShMN0PW126xf8Zbh7r5HQ8GnTECATW6xlbjHOFRMmk1Z4GDnEa
5s3exy0MDnAo4veXm5T5lf9xDFFEIKUkscvaPiaL77hGJLN73u1n5HZrmOSd89dCRHtiNDRyY0yK
APDm8+FEtPwZH/fC0I1D/VuKKmxIa5t3uaZn8eqGV0kYpkdwi6rvsnqxrfr4/GRihFqP+19h9yN3
DmUb4bi9H7WQpsrRxMYgOZpBhOQtG1u/gHazDYeokuLnNbenH0yyrk17d7ku2b9lezjkj3qb1Do/
VJ0fxPvTfSQIs1jeUQqhWnAh64s4gOPBKdLSkKFtfuir5TFxjuc+c1d3q7/MjWbeq43EzGaz/Lss
lHH30pwq84fPIv87HV6stp0gY+Nzq/olEp6QKiVP1aoWtsQQ7p8eEaQYM2cBSv60PkQYzK6dswOR
rYz0djVpRzWvfJlhOH4aL+YCjJcRPRz8lMSO9PXGDKnG2Q+FSAQUQS/pELhtLRj5FeS9DKcID5S6
1rIIr8wmDvRDqA4HQq8RVxpP1sTiymuXWfBillwty+prty8DDFLVij/GGXdN4+9+WEYIdNtwpvbp
+ZoToTgXQKOL5QR0z98OmRnynsTvxW0DnblA6lQRqywnVb4UaDlraxBKkyI+2r2OjLOM6Gri1gSn
QHusbiD4vkN+hgvTN9eVhicSDODZgbq+bTHimeA0Fno+N2WMsOmdgdX5Y7/bUGpHRm0JEQ3RZysx
Ky2Y6H2Z84m8e5op5OlTfjjIrDDH+y+bTD0ntEBDHHBgq3V2Vv8uuZWbN0jSQHEOm0cTNNdg/sqr
v7F/++DjFoAUAC3EiQbA1x7ZnVDt5JRMqz4P/JdSZN+8SvR1xQ6flLVgblQhW88uJbQNj3X17ei2
LT0KvtVnKGZckNlTyt62Dut4D7n57SOxbYrEsCnxv39d2Z47ZRyPX9pGm+u+zDO63h6gRm8RAZWG
hhfMcWoDcXM1F26cZYCc2ZQDrnWGc7ysvGsjGtPYhmxnGVINtnOPMfog2ZsX29QsPBY9G8XVpcvT
KF75eT9dKrY72BZraWmbWp778vbjL19ozdYYTq4izBudAPs/d/UGsr378fAwfplnlwL+QCuCti8a
iC7SqZKZqKKs5DK+FNBptvuKR29Nnky8QhiSXKvaw89UvFHAPeQde1/j9iYZn+pWxyVSW0ozSGlj
yXOKInUyqiKPfXgdy59/3/SO2Q5CRQoqKnvsK38LsL02hU8unOL/jSQYCH386FD8DpMJSJT6iUTK
zgctblKnn1QFRSvxOHWJlaE1zTLwVA2xhZ25C+dGyb3V4uwc1Uc/z3uyI9SDIW+otgCaqLGeruzB
C6lX77OrO3ZakGhnDNVt7o6GyubSvO/ekBNi01T4xgGUR2NutSXqdUIk5gRYQyesiS+n6AnwSo3e
XUMNwxOpcXTjGWgd8d+zlRpp5kSEkQwzNB2pdbZ7i9q1lvJBweZzWER2y3DQVbGG4EyKttr2jy6m
+sFqrfeCeo9gMva7/KrRY4vt4snaPu+hEFxaE3iwmhze1H5H3dAk83nlBvNc5dRZr2nJCBwcGP3v
rmcVSpZsbjUbhk01czllniZAbokPbHgtsgQNd6+XLg4BcH3JzH5fN1qsxl7JY8OlSg1Cu1ykKDob
n8aK6N/g9+p6xzZA7pFN3RuvUij0AqKWqCoRHAPyuq5iYeFD93pOgLiTxlZFOONIH6j0QdVS5vAB
wdlmos4QmAA10uoVxWXhYdhyn7cYmjjPinzCzL18kTucY/9j+ilcL0+wZ64EPaTVJ7PV0fWP3tfX
FN0+AO6IYpp5HLAwE9iiy9Ic6PkGcxwUrlLoMED68ZgPk8QvmEJuXvgKQlXmLwWlHgxmvn9sUU+H
Hw9ri9nzqA4JM2Kvf64nY1fIA3HIvxo2zb87V46fFPxk21rVpSZS9CF4+EET3bEMrGw4YzD2uk23
osd+UkcN0gnFb9CxII8rfj0BedT6vevU1nAuxibOHqNNij9xWxc+CohQ5bKlqJ28SLVUu7pSHrWe
PQje1BTGqO94my5dUh+IG0zxueRKUPwEfI3QDTo/5ngktcwB2hfcCr81qJ2DoVlnrxmps0vWSoI/
EgGwIdhdDdcjQGqMiid+izKfv4eaxilY3vne9QEpMyglaN7t5so3SjsSUj/koT/H5nPieCeQ86jM
rPAwsWph5km4S8SP+7lVRvaN7aWzLCQXVA5MruDpB1ttFGJlbJfIsGN/506d8eOM+A8WfnHyZ/Bs
/20ucWgvfGEiUYyCuZpRiDSEJc91bwXNCaCH49pL5Z7BSl3T0YbTQUxsSbLUoTNFGG4q2sziGUTT
VEK2m4N42qslntngqdujIuk/TPNDoDlCQihJoLmXhlr5v2cefEWOBsitSlmxdYNdPva8zF32tW2/
wC3kRirkS9z++HZeVvUwGEGvD8a/ykG574I/B52p8f1cG/uQBAwT429whfeEJ9myXOXIqlTIqNpo
S7pBTzLO76x+9u/NAyuk6dgt6iyx2JreEVjUNY58G3Q+SjPFPewsuhfplfje2ieMFcBzsRoEC5ZS
sGNJcHsHUNCq2CmXwIo4g5sr9ztQ3S9NUmKl6xZOd7BcjmnIqJMk58Kkx9LMtVTTPudMNe2HecMA
Exi+UAGBzdzOm0jO7FrcK528fvTudLaYO5bzrKfANTqLgAwBwXK2ZLglNYkXJscmX4A9QbRl2+P2
0WjCqfILSg6K5ZnZ338RySC14bsv353k221pBRUirf0dyDhnA6yt24Z6w/NfQLbobPkYKG7X9/KT
RFV3on+5IoGxzlLKFI0eN4HEiU5v7A8wEbZO9KXfgmzUGkoZgH1zgCTTkrkQXMRcqMaVK8nGX2pI
xDiLEJB7hURlbsSE6bnFlYhOlZLttHr+oe9PgVzVvBUvLv1zvcIMTtlFKztMmxYiJ4xvKvttMvN7
ldaur5UCSj4kpbPzQEMqoqYwqxW4wkvbSFajHnc6ipC7dRvNcYZziDNx1OFUFiVDZAYMQYy4InUn
9GYSzkKG3w3TGPFN3jkO2KaXsag16dhEFuln2Vqb0hCUJL/RbGk97XmaFTXqEx8KtITg3UcR6rsK
TclnJNUvfPD1hVAONsrr2w0Y5B+oceT8dVg0Yy87HZBBelmqtx7JwhLJPx9ia3WVQ1WyoD/KKCy5
65RpwtqOFRHa+t1CzEfmhXHxI+3sIgQicE0hwtKqwk0iPOdzfVbFnkETbJO4ErMzJAFWdDgDiphb
hc4G7jZp2gC1wjO/Q4kE1iaK0oDlubLF8cTzCMim5lz3U5KFV+iTC8OUn2Z8IO2JFmxMnj39ddtU
Q5ASmAra4Ns4hZYVDtb57T1Il7HejL9IY5nPl7LCIvQVBRel6+qEBapfFOuMNTYeAvlYr6SGv1ph
1HN/y1LFuPz8hdNu1iReOBbM9TK+zichmz5ZzRjOoZg00sByRVfX+hY0p40iSdyl5K0Rmd0S0hu0
HLsO0weCS/ixfKvrxWfDt2HOOeXX0O2wIpxhpBysC6uao/yt1Bd5vMGnaXvPR0z+Bzti1DFm3zUt
XBWRWVrJOMFOKvjhKRjhwK9SfInRiu4UjPtvNBsCgMgwPdOuOdAVBL3GqVV/0CoRliO49EQ9DnIY
auhsftIF7b23mWUH/ykCQOaMPhjuyT5w3ubOQyAENzqiYH0Wn7VeQ++rPBOu0isAtAcapq40A+7U
GbCAtBx4aFoWN7/dJoKvV2Vntgs4fpFoO87V85WCeyF+GfHTHeLCqw3ACruG0HDNIb1emzYYLeYJ
jTnHahbY9dVBSACBj35rK19FDN6wYUgJHoHdlBrCMY+fLm32dULhd0ZYIMEpbgKnbPPPruSsOWXy
zqr+feEtW4JyLL29FY+pz48NHmNLJ2YzY52wLs8ToeEYwB4RkBQ/yoUm1flya0x025W8RNF6MgcP
br7XHRTVEPgpUwkOOJDPuNFM7WsCheii/Qn51No/OANkBUf7FQFetOCKvex3NssFH3qRQPJkgeTg
TVhVqzZY+45jC5JLu24N9fTwxcCjN3HdS9QuoZ8/lirKTj2aWxkWA3744EnIWjwpOTYWyVFFPUu7
3uJ4JW1nWy4aBEEfPc4nPpOVzkxFY23l+OSdvkbsUmL/Oa/ut+b3jQnI04y5DT85b7TFZs3pdZ08
KZljIBfytb5MYw9VyN+qMKeTpxUoEzA/8qzQAiUoPT7YvDo8lKBSNNQnUhUcZwoAmLfxf3ccGG8D
AQEosupWregHEEMZmnudupPDeaCXKMUsyg2rcydAgk0aVQjc9KYj7isVgrSApC3hANsgeIfVR/oe
XNjjzhgS7x3Ds/Hqpkv1A7t5ABTyZ2IfKwMXwRM8ubXDdoMuWCxCKc1PFQAmLPKBW+0F0S25wHa1
CJ9PN4KQ7jpynLMzboXfwe7KUMuixx2qV27SDYKsVDMTPOM0YeQBaJUvr3pje/v+6GppfQT1yBIJ
/+zF8kmZYofFi4hc1KefesmUAoDr4/0xfUBW2FcwPAlKbu02N1jdbKgUmNtav1NpIayncHthd40s
PIpIGjxp+vjxMJ+s+ePrRrzXjiPtpd39N53dG2ky9nt0R79eAkAX6uqUmjdvxKkFbQDw2EV/1MyT
DkYwudLf6MVjCuws1CDceHVxh4jrRbzjGUoJJ3eBksaAZWwgsVErIEBVJN+pIpeeEgaBuc5SgQKN
MQgCY8rFXQ5MR30dJowwBQKAAgrEGQRc301hSFrvzWc/Jh/nSDfOLmv8BV053q3Gk/HWIx4qp7GU
MYQKFp5FLz55CdtHTgdOq5Sr8ZVuCzmPLrmmYPRrTsXckY8zYFRaZjx9ykhF+nzNDbRlWN3tp/4e
uLgu57Hlja2vyVSREbMf/xUl7jQHLw3SUdHAM5IIA1oXlLoseDO9MNgiEuAEoIRDJdh0DKoFrR92
0eBK7DXmAMZ8d8lreOjrxzR95e2Ht9b4veD04RXdTxec4b5huXQpJkstTP8akpMohmrmSoRsZFtw
3MHeAos3HVY/pOsMQ03ZbUmSCyZULk42VGaiDUb1vlYTVWStKafzU1g8X9S23Ii/A7+PKactA6CT
VfWWOAgWl6chpz25KJy701A6RlOi8V0vQsG53AVf9wIZHEaeS4OtAnSvHPLJhFv9QjNr1IzS9rcq
3mkDN33z/wx3SQEkkyHJDbzZ9IGCbb0bTcPUHNcr8jvNMztDvy9F8/Q+8IZcjo3lNRz2J0eiZ27L
em2/X0ssdN58BhyOfJ1TEDCLjdxr5kTsMLR0h7EaE5pVAKEK9/5I194piVbx81zOv1sbx+Iy4+jr
oI6m02pB3l0EBtevGhUMnvHk28x7QYI8HUXrCDZT8DDGhBjNvEOCqgBYFm90mohSM5+G5JH52xqy
6Lg2WX4T8D1o5t5XgHXhonuqzOk8o1TVVQ5DrxhVzUM/ltL910GwIX9NQDPipK9ypvvLBk7sLXni
8Rp3t3NjaKn8bxsFAQ41NbmGCboBmt/E8q/d5kdt6+ck8hZmyDdkFlbB/FW3CooMDuelZU1KpvNa
UaQAFimtyQwBj7X6EAS4eICs91fTY57R8KkUARSLwNkgNoyAV0HecDCsgoSrnOhHbx6cIiouQqSg
CSTdaCJDWWy/unzK4ZxUvdt4mrfEukhDB/nJoj5deYQc3eXBj9cyAg6zkYOPcDIF0f0mIwM6nQEB
ynaGtvF0MaKWJkog5e5Q8A4zDbnPbPJthiwRUG9VIE+IqDhlO+zx3jmpZxlMT+3JIbx6PPAEFFut
R0O1DFFvvPq5JLvJBYzLcAWpfkh1nQ+Vu3h30bFyJZEHXSsBgSTNThWf7DllaG7rK3SXrzXgeWGM
4I5Zor1aFhOjKYdghUfCuqwd9h5NYje35lATrTs7nwrorEH4AYv7hl8RafQi9QzXOjejD+vhjOXt
8ywYczQvK9+Ew77FdlTSUQqkNYgoyY6FQozUNmqmqyLCXm2hH6dfojNRzVBZKnrWC4zUoWSxjBFb
wfbyJpZjsQiWVuwg62XccxagfyhNw8T+K9Itix8/eEDY2G+t72jPF5KaaiInvE4NF4K0ZzHT9NBs
DVWf8Bs0Y8DYq+ajFYBvuO7UuGAs+a+ebrcwumWF7GhPICVJTyl10BcR8IotHzrtKt7T3evTcK+0
3Ogb4lHAJtbdFFqPPZ2a1nt4W8HYZ9tmG1IV+miGozeoNM3TBdbaeKBI2+Nwiaby5kVpYVpa8Pyd
Lm1mvg71xRdqQrqG/msahuz9MLoxbHvS+Yj2QsC+X9pY9Y82Qa1Ztfm/ot9raFWxwSAV5P67DJGz
+BpjCEYk0yi2C8vBkEh3Tv3rfUsSsOzL4RPlzIfsjkNEA3rq34EgaE9HghxVNZFJWS1AY288lgga
wkHel4GLgw+lA4kXmONmMYHBLYYue4rypUxk9EBXOx842wDJQ9yC5wP+tPluQqzIoZXrthhOOC4G
h6OHPd8zB3w38oAzqZCOngDuLYWv3UJ34JJFPO8aYLZwH1WN2K0jxcN8dox3FO0Cnka2PWaxrAk/
GdC/+QWATLrx8nm48l50Jfl5FPoS6m7exyyeg7pJUoA3EjfzTXVBsbW/RF21GMp756KMecsqOAq4
JZE4swvD6QVJ+gKLxAHbowHc0ybA6pXG0CKlv59iChxYtuPbnO0mXfd4LVvu7nT1wgPyKO69OUk5
/ef+qY2QMUhhnCAceK4vlJsPHLW+mGE8aRqT2fqqRxTu6NosyfRGxYfiYt02lwOOy54hGteWu+F0
++bopmGo8ItmP3W8m5xmQ/BV0yFNlmr/lGBbNDnuQhUYI3MEWdJeriiluVqzp0rK24CsC1DpfUIG
TjykmMcDFyhRVcxUvdKRZW4oEIeVRXTEdIp4eHf8ajD11CQIBZQHEPNUpq3RCtjdrDtPPiK2qMlB
jFHRWvkfKlXjRWJlzVm3fofpOgKWMCvfjTvR8/FhZogIo5kbEB5F+sKUcnptNargqciu8lxRL8LN
erH6e9ZQJenh+Y4t/HdIdKYeowF+FPZjS1lipOSejaV8/rLI/A5RK1s3JPCKHLVyv2AubktI3NPH
cbDKN5QIXRt7TOMsxaf7x4W6kNZ06qIsN0eBNQsrZCBFZ8dSta1Bo5kq3Rll9z+oUKdCEoS8smhN
CDvL4PIlx3YH7fQ66SzFZfbZCKD4aon0U81tvNp1Bjmwin5BOohGvoYJJnewoOOZZ2vV3CNTp/YH
9+JyhUK8TnqNQqwP08pGl0q3ETKR6EkSK79fzuZ3d8hsOsjRL6nDkOzHYcYhrUWUOxPsBsq6aMCK
6oFnjWu7iKUiPzSGeAqZkX9piD+mp50tQE1LhQJacqqGNRHHQ8NEZLZ0ID3V6Nw6c0oBnPtVaCA6
JPx8xtARW2GWs2vU6UT4xKLQzVCeLOzHnRb7Vf97iw5z0CR93iP+O1tET86EZpsMorfqQSFRP/Zh
ZVrofQkh96lh+ol424N3ji1iK8bFx/RQuKE54birRIh2nF7WbvO8/pqFRBVnQRL2HQ9qXCmVLcxB
IlG+QPr0Y3OJ0Ae6ffvXQamQItsIEN2iZTXjgNKzTmO91JH8BhmU5eNHOfv6vBBUrV2KAJ4jnTMa
023SSoF4EWf4f6q3zEZg04llgNBX5hPQJsTiwdRCY+Fq+si1nx+68GvO0rZYdfGNXriLa7OPBSqs
X+jYpJQwo5FaOOEVmD/EIqbaey6i6Qw8S3vqjo0fIl59abb78uWcjl9rNCw22qzPl0erEp6m6eej
KSqRlYcvdaFx6D7rOxW65qwA5AcBoyGwDiPMoo81/p7btlkHeAAsn5se2EEIWm3r0rs0tZ8Wo5jd
elJtq6xjUsEOvnfHOWK4a741trLAqEB836CXIeeOblssZTVy9WH30qtLQ9UUClCpC7fFWQxRq/en
LhfUaW8Ui7KfdJWXrFMwRCZGlKHQf1PMSFmeRXzmneJCgY5jl0LltlFymqlXFPOQFIF4dBXlpdar
yChb2E8zR9X30S+Ub6ekiNQZgT6tPSl7lhHuCveuipy46XK0h19m/uJSWB3AxZt6XSQc94tCQAg4
rGLcMYEUQ9sUw1KtIc9UxrGVtj53aoqFqZnn5UfOOz/BzP2unXUXGevu2PiMWy6Jp3zG2QcBIrVd
01X/IPAG92bW+bruSEk2FF6WBjRKVk7Uf8E1WdjFQlrsXbztc9uhV6nhgi7yx+xurR0MUG1w0Np3
gSIQcs+7ukl2awZjO3cqo7YUjFUdrL5qCva6Pe8owORKizyHbWVckx19DHG6dkgljVgB4P7QZRzZ
a9SEqSr9WTaW4ByUKXOfvGHgHRFnERXs9PPAsZUfL8MEtR6d95TyryZENU8OMTY6Li09jwDARHgU
vgRVdpX+CDBaLgKdCqWKV9/959RhNlWYWpHhDON/QaPsB3rLLRo0xCzwoJ4buiRPn4cI4DvpCmPe
KfavdvdcJQOJdVSmBhPpe/e/KiguVfXya1OVD0C83sGbkGOP8mjLT9lGU3wpV1zOJ4CxScTw9sV3
S3HUoEFqnfYmoXcVyXqOenZM8ngzwgBphqIR0SVgNV1fAyycpVrglsANLuOGg55ld4zf9TjGoFhl
fNkiOU0ZQbmdMMGCpHwFbr6uo/VoTdjZ4I3idYGtz3ORDF72+cfUFWegVV6tLIrOHlck3F/RLEcL
Hf//tc3fRCyiVDgGWgnSJBDciuBydxwJ7oogU4agatOoGE96GCR05bKQkmZGinN8kupJUwy31gCc
OM8lbIqeujUKiaP8vF8egukUWoKDjw+rx5OfqzyPO+H1ZQwjPf/TetegDAkgewQV/2d41Y2mOcH8
zwSPjmrCtfKj2VnTesiIxNHLgo/UsvkG+nYiLDaVNi7EjoSTEJMnByVlVi9TmWB8tKES7rMws4hQ
k5WvIYSk6Soic2Uu8XhCC257AVwd0zthewdH4nps7rGdXecsFa3nm4IMXHv3nb7q9ooUBb6fj3Y2
IR9B6fOchR9g/Ivyz5JSpmmLdAEeGMtt2j0iQu+EyWkCVbW7ygIjtd3ukdLZNR68gaEJ7WLQrQTI
XyvEy35OwHrV5xJH7vIVvbXPt+2RUvcCGI7rbYqfJnGf7IltMo42Yo3wgzbqDTCXjJUnGuycldE3
bHEGSyWKMPOTEtkv1a4zHQ2E7NiW9XmO6rrPltNAcMX2oBQrUU0KJRS6Mqaio49PbY40CYZL4JmC
MGsBeW0QRkhmzQtRipBL93Sr9rcxzfRRhQcroqGt8IERY3dvIt3wH+tp3VxbY+gi9VjvpbqtBTzM
guWOj7jK/O7KNi2AwJ9uGp/HpXtXwzkznKQAHJoenQaY/WV2c2pYbCTNk2Vy6eKryxybMwAYAZMy
U/SvtmK/uumOskmjnTmBPVZplOPCSl1PxqLoUuQepaRlJ2YC6pcAI3mTxf8u8NYvVK8Lzpx5NMUz
gtVHiucSyptiLKKTYPwpXmhHzDH4xWyB/SwaVmCRwAmIXjwo2ZeO2MX1RbEMJDXYZbpWO9XReP7t
f48fg8+hRnSelk08Z6+AU+haxnSlSC3JAvgTcnqABjfaGwmBe7XcAcmdqXnCwQ2976eoyNnJjTKf
W2H8Co5Fm0fV5zR6pobYR8Nv/hGxuAYJi0G8RErqid/UhrGnDC96sExcLp3tnl5RQ0p2O8AUUKsV
ExYsLDkKEpWapt757PyhFizv9hlow7vqAdtq0M7DPWIbgbaywf3vifyxya1js/21MaqMJFN2r0cU
nmJdpIeL7TFQ/BVt+m9BXWVC0/EPlCJXFfinnCiUu5AuuE/yPyXj/ha0PqDQY3QschXw+JlLPFLG
evMHBK9XLMsStglNDy53u3LVjE2qn6mNf1jj/fPTOTTxHoOeQW0mskW5mPOtxeCEo1f2eVJLU+3y
hpOIzXSYqZkcjiAoqqOi7EcqcdD9aYbcCKmXv+bPNGw4dyhF9VJD5oiKQwHAoj0n11SOomDFThKT
0J76WBmV03weU+IRRnmWPsUBqcHmZUOaEKUsfj+nqhrWrWljaXQgZqIKPvV0wmpEhAg1q8qhhNmy
vKhdrb2O3QnNXHbB+xbYtubPEyVTMy8UaqMkSJ8QlR49nSrG0zVoxW8W9TMoBj2S+EgdLjgLr7sS
H1BQqduaj8OWTIkVE98Hjhbx/97VQcpT778gls7LtGdVu8uzcwTZoUcexJUz8ouoHkWhUXqbIskY
eVWfvNSjmojmtD4iLX8P17tSqiXU2l+uXPbYgwOjfqFgdAYEVE1xB41e5/Bo0ddW1VZvMClCCP+L
YQ7p+E7o+HgYrTQhiGUYOLzN1cwNgwpQh3R1ScWKKBZfTfO8yxKZehtg5kMa2vcfx246pE+p77qm
MpCkZwhayGYx07pUllwq53oK3z1JJPnhqeuObfvjoLZzK6wO3GzzKMH99ZgweBrAozDHTCYLEeDe
5TX4+a6tKsuVR72GTMRwDs4ZHlRaYG/ue9JkePF+F5Zugjxu9bhBSTq0yyb5xiJlaawP0V6J1pyd
QpL7dE0OrDSUavhVQYPhsf57OcbB1PByk2qdhXRGfX/zQgwOIcYBP7WAIqzH4xbi1XTsnX6dj0mg
ONlNQ1f6299HFvD0xLA423uj14+I8SX7tXJCYJu9cP9b/4YW4dCrOo/JLiuOu3alwZbkS/GqxlFK
TH3T0SYoq4urXZHq9nSSdj+2XxkodHfZiExj0Z9/gzD8HPapSDc7ZEoI4o9YmHX53B3N5mZimVWY
0FE87sI1PTvCIUwCHUlFvBiOfobn6xb1qk9T+AcVBhk5nbeuJAbjLN/3HyCSIe/TMCeIvEUTqflt
cUYKZu5Cyg6gdhmGuNrXJhDkxp6d6zTcVvHv+juAc1+gUvxHPv2UczAkOPYquBnSVSBg9G1qwusm
S9jPoI5bX7FX0WAOsmLbhdKh2h4EmedNWZyG4lJl8o4FYsmWLYsVB+w2pJ6B+oF1SG7yyfschEpl
89RF+Zz9Y6gCiEhBf4MOJPGewlodoholr+MQ2Uw1LjE4Bu9o3TDsrdL5QkWlauPQRa+fhgvxgjWe
OWdUDjn8e1LVrolWLkSUjejmFuhhkc6y/vWHM9994tuepn/NgJlSUGoW3R1QTCqf6bVgIIpeg0f/
a29xPRtKxx6hd8jaiWL65d6gDCj9ImGYtwmUReN+nsP1NrS+BY7HVqIK7yF4un93BW9Jq8gDZVUH
q1/UysjlLyomtPVwv01RG21ybqJl2DcDPkw/77RvBaY9M3hgpl+HDibs3tId4cFaiPeu9EH6DQik
Jo4Yi63R/WHEqoHm3aEr2kExuD49LzS830vaTDf4LNs2FbjLpNlQ9TnaCuH1xpNm5q6zPZuUcd9W
8aphIohtwwvMkdgB+wy/OtQNcFCTlk2gRlIgDfE1b6tUzW/z/83Ar/V3zG2eX04B0eN1zu4CBaMI
2BbYODerA9eQETVoAexnLmKGRfsEc01b4TOZd42uKha87lkDU4+OTao4lYF4cxMTKPuVhJTQWW51
EbhuCaPADrZwtBeLT2qnOtFT55NAfFtBaCQsLJc44VYrFeuohd3mkB55AdpGscPN+r2Rz3BjWOaL
E7sdWo8uxJZR+LvdhtPCbcxsr6LN6yEyDCCmzKKk8SJJcreLAA0IYsjhsHU5oZv68bY/xgbESoCX
6U1Mr676WSfFfEYzdmDAldZxhTdWOpnex3ZnLWw02sphvE8YxbFE3Wq/a/hBAcTU5/18XDPFhBo2
g127UPkXzOa+rVDZHRahga59dgHqMlGgobXh6eBeAu81TjJ1+jgGojq4e3v2Jox0Qn5NLIK+sJZW
opHnujWMQJZwSMCacf8XTIKPCgF3mjdLmZoo3XndB4RqOggzcVds1FHKR+Xhk/R5QVhPzTfcRkim
UyEGQa2pDqBj3rlvqBtuHrG9QoXYtRtRwshkXX038LvIuKEoiGnyVE5f+5yeLUk7zc/GPle+FK+o
fbs2U6fI+nUE59b85UMb+2mX0hg0VRLSJP1neQ+eKaB8wmukkFsdrxUA3gdeXd+McoA5ydPp4ZYm
6qMeKUxDcLJJWiRLdN9CLIsGf1nPGkM3ubR3iPstKv28wm2S8dk7yatZjtexkI+mSEzg8DXycGLr
3SkA5Wl/w0j9oAIA64yaiOY6cpDEoabKDTY8Efx4P2hR/+uidDotTVEoGcs+677poUNkucyiFiOM
xXhb1oc0HFnxST8TJwKahvnSPJTheZndiBV4DkNjbzCIlQxeeoelgoNdAhKR1WNNRvVGghCxXE6/
+caHJgWcrLffBx7IxUCXnlHsZ5YmeJjEnbybIf8vJmbqnhzmBjeBFymZt+E5o3qstCaqul0+JgZq
QTjWbIsAESD4OfjqcNQeAT/6Mztfc1MYP2Rfk+OnSLgK0SpGSpdxI8ruPYp/b4OjwFELL6f1pPtw
NBe3VFJrFELPAqvvX2EQFFeIG1XPqo5/BqyculiPNc9aGGcI/GcKHFQ0R79YanhqRb9DPbIqemO0
RSlNF7VQDaaPFD75U1l6jNW7h0OcFe7Yp4nfDNKqbxdzJMS5mHBZfm+J5LB46q1kaj0yovwLrfr4
0kSO/LDOuK8hN18SXveEaLfPtpXETKQcXJMUn/eTnlGhVgOSRVaXxVY4LmnGmNZNYQQH4eo/qKWu
3ITg3NlcirGB8sT9evSk9tehletxhGZ13IKoP5K9DcAJGlZOtSM/bsYEQfiC8dDCM6aDe2ENHYDN
+w0PX3DnYOybeGbeH1ufqLDsHk+hGsssTSNiTVsDcgLNusaBPxjEsjrjXAoeX3JucKfoHyZ4i+L1
eqblXuIqA+/6QTZSsSV9mG08QPw/xYLt/2Hl4ZOviih4AGkREm04buL+TswmiarfYhFGQBGKL7bz
SAbKAp4/Mgm1odQcRynYTSTgBey5OyKUs5XZLFhFDCJvmQC1/Vohq5ojcdp4FpHUwZNwcEintq8p
TkJqOU1tbxxAmhx5LHaMLfn4nUtErQprw8dbdNsuGOCHcqIDozy66QFVQuRHS5ws9EXweJ0Kbk0w
+XoAmgsIXHJ5WcQAbqrYSU7eemgPfTig4+YfsApJczL0mZknM+MLEhzAVGaUCpdo0WkzTFDFBmPx
Ozi2RvIPBN0R7RXHo9bU+ZnhBQLLjg/M8eQChKX8IxTuP5KOhp14jN64W0QdxiP9njq5TMxVUPBw
JR6OEEtbc2OLObXYxSaW7R2EFNCpQkjK7mas1E1FDtba6aLjVWNw8OSFoIRcibs6G7ROTJDn+Ss9
8fakmKpxrqUEPNTxkDSkDkog3iwBTjGi3EsJ6YUmwHGfAZhu4hPQrwKzncDwSOc790Qbe1wnwvk2
ulLErag92piVwcssELBFMJIdiY6WPf38sLiRYGIk3Vg/LXGUnUkF9Asy0f1jEoVu3KmTKAAowrvi
BBiEW3dOwiNoGSYy3/HN13sIfp94qDHZuo89E3OMYDCNHqobZcqQFFB5xW7esDHWah98BwP8ZGRw
o97vfnDSCpzWDXmCjw/jxW0GH0V44IVQ5dvx1AgI8Wdb2HvKh4BEdsUXj+mR4SU6virvNjnI4Efe
xqOOix6e1tgONBlT71QPqZHOrjIVUHXfuKcvts1YDtDGHzTNkWPau7q7tdD4tJTD61kCfR+36Zea
Q5hzpDhBjpu/xTFc5iciLCK4ZkAfy6eN9UHnOy4p0Yll2xqRgrq1S3wtb2mVUI2NDFkp/jf9X4p0
WCNpF9aWj698dd5yNHnyAcbQqDI2dO5VB3wOGTqfWTAS21jJ5DtQyy8gNk262wePwRxHrSHOdNuL
zqoT3cqSrdbe576w6wAnIJT73SXktnoO2O+j78YJC8MbVDRu+pJCRIXvfarrLVUr+qBrml3GnIga
76t2Cx2ZEMmRhNPQxOboAmKi5FpKexaJS1XDNLYPbhGvaNQXX1ySKGWdhT8IVNtzrFxcbQPC6g5P
5YlOI3XvVADEjXB48rGCaYisXYAUz8iZhSlxULCeynNiAOCtaQcp/A6FX5crLb+C2qPCSCxIBzkQ
gREcVrJx+9suw3P6/kyBDcEdiMz4za1HhMEFGroj1FodIw+cEfFiFPXPsrLOP5VLCjrYJzT30Zki
tGKB8G9PsR4qg8Dv11HvovhMObX6qIvwu5fQxSbTjkAijqCCaHUGPmVM0VjEgKtZrdyW7GGiqtGw
YVRQ8+Us1GcXod3wGConihCYZPRiw/WKkwCsF8PsYG5Dk9kZz7Jn0vvzKwMp8tSCfv13jveoNL8K
gL6fWeDwC6DEIHW90y4LJnWJEOYJuHyXUPf86NpaQwj7yDGnsWiEQxYejLrPalyVeR6Bh7/Qngpk
2v7YrjGa3PGZa+cRly/IrP5ntSHLGoXyOBEilKB+Kpct1w3sBLbWHPni02nQXPxIH2mHnlIjAgfF
H/EtS6q2FbydRinL73Axizg3jPrG+0OZkD5D3F7icl/6E9pq1R2T55Nk1vSR0Ah8eMaMc5pVqyae
rVDEQg0nqIip+cjj8UN8Oh1Y8hOO3cA/gaSGjdq0pX8jy1hdSYJbY84k/eNtLDnCj96b9zZujQsE
UsxlV+8IlEKnf2PmzwiZ1hvMeEvLmPx7+njCL21Wh9tNEbGCONNFWdU/IcJI/ibYxNT4zpOIe9EG
kE2Pzcn6ocjBnsZoS+ljwhg/ta5iRGGwaJSmhqt2GN0dPpoPbCcZ2mmA9DGMOzZbKmopGn+6lt5E
j3szunfdk92I/Vv2f7F6cWBaQY1WzyFVRW0c3ghBVhED0aBMz8XXXLIY78VMpZCQfVVu7hQg5MkT
nWJe6MZ9pFVoiwekqve4JwqYpiejol4VkB0uUTVpLk68osGfZPTkB9b7mLgEjDFTfi92tuE/EDFT
HEGjShcBYslYCveeTv2jryBTIdwNQ2ZtLO++xZurBdgj09lJGXL7+nmF9x9gL8Vl2/cnQ2nL3xRZ
FiF8NFFGzzEH3Gmn+7dKsKSI7oZXL+VfOXuLGDUTlUVSD2LrFivzGcd5+8wX5Pax0pEMvSIdAf2X
Eb9/lXZoIpKek5DsKKSph7WXFe8b1I999j/4reDqHCXp7TW+GyJuUYiUxkqlYLtL9LcF5pofVgyX
2FUh8IrsuKgDeTlmZh7QLr3fI+3CTEkKl7vx/rmnzc4Phhsckk7C75j+BGyKAxU3EVUh0OUFEjem
l0d2f8R3a3JsiS0OIJfP+/mbt5QO/iS61f3nFRRvuSCMIWGGauMUrQRTvh2hXaZF6B8UwMG5t12z
OKTKyMcq9nrAFlPv69wOt6QSR6ZQ9uKobpWYr5xPylGicIdLNi4U1s+ZWBwro+Iph/25Veu4uUhm
K0X+UeAFfOejdZpCy0wxpF7Pj3RY8jaUvYwVmxCLfyiWqX6zzUyxym+EoUwrq/p7LjPY2aRCPPt7
S1x9nygpjYi9jefqqYbETHl/4RtNwV2Kq0FJAWsDvy8cbcmuo7rDYTZkNuUDK8UT/rEVfXZxOpsx
mq5aNvTEyTNC9rDAsnXUktk3mqE3MZNeQhOuVNjSeI2e0RZFQpyxP/yLo8FE9f4g0G6+8atqkmSb
lCYVKsJEbtZd8HEcuqwzBiCQcapmxEJgZbJlaSmzt1jEKEILouzgIpQAg6Mh/Z+h+PT0HRlxGE3Q
1VLG4E0fKVhPFQNPNbqigcmCEYCWhJN9et0tcG+ZnDk/6c2kpOBG1DYfZd67nJ1aTB9WNTY322Bv
U0n579X7T4dcY+ghQlPCk4VvO4F3tF0Hlj/Jx7JMkc3IXjXAtFXj+HVTo3z59TxRduLqk15LvR0W
xMMvoC+MUJWUgJSXfl7DDBtU6G0nCTyzKAw/7/VwdT/fxZNBoaJ86aszgGE6HVKmgIL73eTz/Nlj
ZM4nKDXXRshgt6g8E+lEL1Nz3zaceXi5E5NaTP920nD399nQEwHRlZbQZKPtpEC/1rpo+ZiQL08y
+Y6im3hTTGz9SnaL+D7AgaDET5IN4xYU5Q/PLCzWsNvMXLzBF3DcSAAk4pB1miajor8+jMLKXpUB
40zR4nfjGa3KIULGd4xBc84iTfOJxZYGmcQtQ37Y4Jp0exLfRFxdEKVNeIj75Bue313j+078f3Ay
aC1LFbEhbLDKaWSNgoNwV77xCZmKvbzIEFQJ+eTtP8uYZXxct0E+gCpFRJi+O9Q9Bn2PE+PYmFon
Xon3dLlw8AoANheMIY7tBjhpnAGA9+GlZJbWg7nz6FHPAtif9Pl7RWMi2ERvzFhY9N4BfhMbStNz
mKrccIpDCmzsPj5Tr7GjdfVnHXPc0VgOjLG3EVCF9E+68bnGdZYez06Hck/Tg1ZJKL31Ig7ktd97
sOP+XQJTEvdx1Cj/ApMeSCEam0R0kOfkjOgpPn0nioDiEeBr+eHUdMmK6XHJ1LPd+JO6vkx6/Tlq
dhpHhQcfZ7duXeY49cp3ySoeRxdjmys7vap71WjjkasGF8aZju0lF8EbXDP9nKIMnbBSU4AprQ+n
fnWEze4rfaMSr6t8G9Tm4Rer+3h0TP5IVMY/CqBw75sok7fPduh1JWzKCISwOIBBL3a8KiqAbpna
/0wwNI1E2dLcl+NKL5UM4gFduNm+KUZ6V9r7Q74sr2ivIeGBEH8EoaB/uxw11yEI+A8aFNafL6ur
WZ3TztxuoOW+XKiZQ7aif7dR4B6hpQJ4MM/aVkM/Uow4buk5QpMnIzX/1nNSTQ8zqZSu6f/M3GHS
9e/rHsL4/Ndazm+49oUGFLJ8YGyOwWxElER2Mrp/mtrGln98ExNkSZFQS0AXxru6jLfHk0X6AuCX
9Xrp7d0T7hTQt+9UFkjnjO9CtLMkytj0sxZMooSU/PdyEoqGtPjnh3rO3Xi0x55pWUHx2yf9zADe
WgRiNXCjS4ou6PLt2d159F3ZI6hfq0lk/0bPltIJRFq8aBDIn+yNN4Q4RFROg667S94gXvRgnhTw
CcsjnTioM/9ZqRuo9k5XQeXcGBWcMADEVwKxodlh+mGk+lEESpbuPqgtNXy4QlLeQGaLoYfDEcND
2wdcAebJi3OkAk+lD4tNVlvTPO6JexWL/6QvDT7MnghO8AIzDJ4a86q5eesiYBJqznF/5algM5G6
DBOOpJUgeEJPQTazKxlpu4O9WzHWr4H6t7m9xIBjKWnEFLT4LeR5euHL3pq1XGkLl/ct0l7MZPzh
bQyGCqrSaAUMXx5ItWWYxTh8t4nv45/wWR1Ntyj4oU2ijnHwmDULsG8Dp2w8dOCQL/ScA7bFrUCm
T6pPwJW4lnn/Qzo5djb0uo2ne94w0Su+vE5Ks3iD3ThM0jz7MoilLEW5ADqfRISuifMvKGiavcsU
b4bgZEouGqqfE7jt7/0EfJuWAs6SBP0H8GmWmBMzyN1a6qxPKoM+2XYuXkeEu4A8LLeq3S/yV8ja
m/9dFx/Jtb3k52EOLmGOI+zboAJiNO9IqQqHdFI/fRmq0RL0PO+JcdXASfqwmU0NXXYs5x/3SI5+
fBpszv64ol9gmG4fQQvVI5VSnsfIdsZzvSqo/MEK0Ja0/v9YMpU+dHdltIiBxt5e1YnEy4ZFH91L
FQl8GZ3QLgISc1CHA+pboFD4XKKkxOa8VJP+ptZO0EkY6aqq7L10zGl/VGIyL4kjeudBP4RjWxXB
iobMNzTQkOhh5nmqepGpAwQHXDd80y+86zKMmD3Krqptg8E4KOozWNFttlkYafy3/qs9N1GX1Z/a
8N/T1cs4zwyFZz4MdzhDcSEZ9QxBrGfFR28SitF7Dg6/tJ9PH9PCPbhboG1OIYNCMd1kQ/AGQvho
Z6SBDzF2vSV4n8sNeMUHoJy9rPOD+xUZLVrhyhHCDe7betjeyEw/v/f3BZZEtF5/u/SDRJK2279Q
e1UFof9mdsZ/c+zCTmY2O2HGRnB7Xz6JI7CpfCrp8xwicE/iva4ogbu6duJUVMEGvJJ/affLf7Rf
OS51VNZplJXKXqbAaCYBIkJjKYDaovteqVJxE/qRpnGqfSnwdyiBXPmc2MwEb/myVFXZgh9pJSuh
9kIs4EmZVpvh4Us1Vbi3pcLuVAEOebVQiRFqqKeH00evyM1HULg3Dtsd4f7322e94pmnBvVKNVL+
eIZqHCqiRFwyD4dM4oCWL2lC3MxJzPHCIrDnTE0jVaNhXHqZDrbBQbchOfsRY44uqH3qZFKbTLKp
svFdUk4GQoAy794jsmoXr8u98CG5tVBDF/Ie483bP8EzBv+hKp5biaaS0RB1+3BdPdloVcHJ4GLx
E8B/WQo2MgX4rkyxO6cs0dO4AKa3H/j6+aOgcPuI6oqiZlSn+rktdF007uUBK0TeBq/BC150HpYN
Q9/A2r8IXVGdcTMqmFEz5TzUjo0LT3JkCFbT4W04u3o7CgBLP4iR2DmA8DDc8GgQ7FE3ryzI8KiF
tTX3Jo8drYEObOasM4LqFQ9+9VyKs9aIO8wDZvmIE2LVp+25RduL34M/KE4tjnElH2hUXIw+TwzR
AnJKTHhZPyqTQTZBvKprpKtg8bunarE2OJmkNt7CVg2WawwNfZjHmvwgirAIyLTjwZnMDxxgh8tS
XMEc48oP5e/WAfyPv0cnpQU4pUgVNaRHh2EKWqzdiPbMyhxaAUQJ0mwcUmggvNmGGAWdpkE5EY9S
Bg+ltcvcg1O7JJVKr8uwYmR4JC0LQSiMZbhonNfWK9Gy7/9RaI5G9wcReW4CE3p4BVLh39uQPUaI
qu3IYN0ExeM8AhoGgDbHAZ/gJkcs4bRc7gSlk9d8v/wum/kI03FrApk8V+7/UK0oF/jmMtlJq5Zq
Xc2SVLukomer6D4X3GdMvzsiAHnHWDf+8pWxSX2lQTWQNo6F8BShWZVv3YX9AC7KBh8W2plZWv/A
NK5NEkfHcS/r+IQATgnzGOtKrZEjNGT5vEjf6b9LIzassj3W0CVDPiEC4H+LzGMcwBTRSkwFH7lO
mU30Y4jixDT61BS0ODGBlIcXErIxS7/KGN0nzSLd7WquRCt0yUs08pUUBIeDJQp2CeqsIPQTKmA8
UdPxmeBuwo1QW1q/fhdjc8jcnnZk05py6fenB/6GFI8EkbP4Qz7TZ1t31orWfFK0PSjzv5oHu+gp
NqF3QP9DYgl14M5WfgamE92u17nBsIlKQFOalITZOYNEHKKaUE0W9x5OfObh8qBQUv6zCfWxrz9C
pkvv+2kmw6VaGls8+/pML/aNg2nQZTYUe2llPlmaDcNBJtJfcoZUDXDFgmP7OsZ54abVG2fd0Fpe
JTKEFCX3tDfhCfw343pPI6lAR9kyRXdKpEE+Ziu0A8JhfeUvelrJR9Z+Zv9OZeE3FmLswz6mxScO
EjAVdNbGmP5LiM21yAwTjec/fph8pCFDpZip+MvGMN4s/0z0jt3rXhgECb+lEo5aC8tRYilgbTMw
9ROErSVSI6USjtlTSY/sm7dOI/9XHnExI5QprybKvP1RAoRndB5laPkl8SQVAwWQ+2x+KXxeiHqz
5mKHwygDShzfOLjoC0Yb998pLX8z7ke6ul2QyBe9G90yUU8q2B5+WChnGuD5CjzStY4Q8QnMu7BK
iwqH1tLgDWl8tuKsJGvqzj6YpeAdJPtR4Tbwf23mFaun/lMqYwZi8OGD9cw6qbx0+6/Jwz4VS347
HnLyyfZxQTsjoMr1GHtgsK8NiErdi2JdeyGq3FH/HmXxKmz9LHge6qWeH4XCGQ9EH/EJvHgja2YH
iBRcqAdv+IVrNlt/4Y7/nAYZnYdlbdAdKTIhxsIJG6wL6wdzuqcGlXu7RZJlO6oZ8ymx8fvRRLCJ
zM1ZptAHlEGQn9SGgEpGKgXISkngqEN8avsfJQA6gAlArEO1NXRgeqN1f8I/bJA+ZgMDFWT/UX54
giC/J1qxSCdQtC+mIXhhjHNigjLFgOfIF/SjMxs/dFzN83ClAYHBwnlnZWaZJpMekay7hq2pqDse
WVTfrMJWzQNOm0QftzjujbKkfF7ggDiPa5E7wmmUsDocyq0VGs/gsQ480msdbPfSVvWHN8tHf1CB
V7XNRGk9pjkOjlRQAt+DB+KpISRf1lWrnY42HKq8P2Rq10rTTEeQAiM3bu6OvHRJtFPR/G/Pk/PG
00Z9Ww+lBg+8crY98mHWgK1mJaUPSWmzAttbd7aRNWllA8Gd1n+cl1CsRsWmdUA3mPVKNlh8Wa6v
E4mTb/BsCJya6ClwQlSQJbugdoMNxATnzdvnqdwvxEdetXpK9tGCmOKVoR+uo0KL2Gl46E6aKyFI
t/oSZuu39oBFYPfxdJuklG7IKpQQ1Tit8FE/4p1FAzMNqwodsCK1pYeleULKWRkT/bvyuqocAXLK
dvidGxLqQTe4bZc8yGArWOvOPGan4tx1zrMlEmkdO2A7hJwmxPhXrCnLNZoTx67jw+27fD6uvpYW
/DFm4/GnT6PUospIb7Imald1Ec5e8vqPgXOoP/JwU8u9E5MPqLxAlcaUtWaPqgiL0t/RvQvffTyl
AsdD3vXRDhJqgSeDyv4IIR21d61r9r4TpVBzfCM1XABIRfJ48hqD7JZOT8u7E5wIwB6zVkHrzpwR
I8Zt+sF/mKZu2RoAAaQFs9epb/qqn/BYay2o16MD3ay3R0Sqn97Y0S7QYUhQ8u5ERMegs35+JXLz
NmRy4CQ4vHMelyEeZbBSHIWrVcqzwG5iYMDnLYh0F340p9Mhl8AMR/mHC1Obwz+f1aNS0Dn7KHUs
DJ+qiRi6OQrIwkdxfZ5OFueIGrXy3KU7JglcimYUwudbu7HtKU8ZZH0HyWZ6ePrrww4bRhaRDEUK
5IdwSL6HXMYaaBzdM4141ikjzLUeXGX+heakwegkCdxemDlhWrs9Us3hkwpfZnCrd01TRniAUnqx
ICW8SwcBwlQOp47jZ5XygnKeMIX66WVCJaSjgFheOvxWkAPcLISRV8upZ8tGZA6+yXHAiWjaBBjn
o5/9J+4BaxRqs8l19vWv0Jh+HoHoFOABS+t8HB3psakk8wvL394/KxHRG71f1yajji7OFwwuQDtb
Bq/cs3mM0PxW70FmR0WbdQ4XiZvO8sCRhVJqk8nWyOUGYm6QZuh+qDZqH2+r33ttzmtejYOEBSka
rUoFLJyebHEuOMPjJ/SjxoyOmsrJesuqNXjUwPRjDc7FJhElxdMWOniTysHvEgBlxEBYipLTHErh
ToHpwvUDeCI0xtkbUDmcK4JqXdvzRy8deU4ceuuv6GO5XgipJpjACn14Gpcf2O3npDjptWp1Ch4g
LNBZMtn57dmVhEtzTy5UPUcd3yt91uIPUzU514tzMvF9uZtq9XMrtv9fCVoRuoOEDJxLVCRqHGrg
HndFx45QpW9v+af4hx0uFUh6nRKhSB8mHC0FhiwmUTx/i9Gi0t9+mxycrn4OO7CFAsMrVUwlwQ+5
Ulx9Ep2SlMt5mhaYDTU45w1XkyeO7T3mtSZgE1Vi6tn+3Lf9yWEiq8Ca4FsZUVM9igDVWwd0gwHf
7mlYHUXyW6LF9a+4wDX9Oh7mKGwZ+wroFcqshWAM8+3jjbKpz2EsBYwV3pcaau+/vPS683NJXUqb
HZ1enApOi5tAwTOM3M2wudhnNeOFjCsCGv/KcXGVoqnaGKra+nSzLCcCkybTilUUFJskmtfPWAqW
Ic8j78xQL6TMZF+sMNcexcL7o7wXDPWtC8PfpC7prgsW5725y8XcCe0JAlAvXRmVnDCAM4/MGouP
w/m8aWqhMTZwQtbl0B9gutVOV6B3m3hSufs/MKA3CA5Rb3ft+FxrlOnqc+QDX92736qzfOB30GXc
CDSMVAYpAJKLQ97/xhGwa8o1aSAQeUJ7XohfweDOIR/96gGiAR4tSxCr+pwA6f37PPbEBvfGLLaJ
tjHT0Bp5E7FYCztpVWRSplJkJPjJ/YITzZxvZTbVk758CMIjmrV/gvCYGWFzJ+hx4+phbcpk63DK
zp440ZjnJh2PfOUIptxhTAvrLTFoWE9ArwkjSXTHJvOKIpdm9/gM4EJVHXoya3xqrno+EIWWo3tX
+s5MY6OgN+vhE0CZzzXIwZDDmS+0bO58is872BVvac1Ge8kQnae34Sg7UHWis67Ra+XJOmaLrCAD
SVwL+3IXQ6P4E0uJuuy7gM7sbGX4qA9E9Gw4V7e3NWN4IGDgzfcHf45g0rd2QDL3lvrvQ16fjbTO
iFq/YaJRMcd5qsbFIUHYTAuVW/rCY/MFbS0Om8ga46wzg9HrRHO5uP/C3x7uV+rRxpigfx+tQMdY
r+1dJTlzqs8i37HjCXd9Z0nrCozWgJ4f+9suvodvxxx50/i3MAXF7Zw568OfkC3oAACba0VgVgza
MTa+yzyabE9RbvgcUrv+fGROn1r78EnOMYqGZxgoBP1rI6HloTHMBQAYVKKbOX47iBv8C4MJMu0B
zbllZtIvsAyke9SnsQHY64FveMtB9UHgqVvOwb7NKJ2HmGpRuOhwUZug5zaVu9JyBNGatN2kzdMR
uL8kA42KeYPmpVI78jiiP8nyr3uWufjzBGNuiDw4R7ZFGbUmayr5/27ibUtlYQE2VqjudqNFhaPz
FDgyxfRVv21BGRpGZzBZx0w9k291FbBgqg9lRZnvkRynXIls01WCI39z+Oxt7PEC6KcSPfqWXyhd
gswhF2irnIqyNrvy57XRf5wjSI+nJ7xfFLdiFuoMfWhlFobQy9GLfWZSDbP+NUi3GuqlcScy33L3
8SfIWi2LiK/9qg9cDdVkyyeqpAyxp24JzbwnncB5E6VdBte7MEpDC0G5s3Y7j+c+1sDmXnFHt5BL
GcVECVzNVpVCBL4z9M4y9Ff5H+0V35if5lZ0ig8IY9MQewlBhnasj0w9b4TlRxBdEJFrXr82J/9E
gCUVWy5trioRVuWxoJCP7Ttw3HwLR3n/6sJpWeuYjh1qeoDUEYqPot/w4ooFB0G3VEFt4DYncUj1
j97qrLE0Q5O5tHAtawB6SZr2iINFmrhXHcGzP32qqasbtPa2HQ3AEWgbTzKgf6PmtIwh74oi3iCS
7fP00CBELeEOove4lUhdx9u33X99oMYGFPYbF+mH5+3HRKHEWBcUxmmh8BFnCe0bm6HpJo6dtfoA
cV4AE7b4BplPafY6drcIOI9K5J9P+Ll9gbK384FnguQqGco8mLvZVqJKIkWKV5YDnMV5Ld7natNk
vS9wXYFQbrLYpvAu/iF0AzAofiSSFgjtcZuSQfRyz/zTFr5nXymgntWsfpzOhfhoqDFBv7rP7ioz
FKZDNmroMeQ4SvswOPHaSJgtGGqDuycF5hq4DM/DrbNz8REl+/bxEXa7F0DiJ1PFLg+oiJFLOsyf
hPGK0pUyXdkAn5Ko/8g9XiuErqkbI0KpQFLPPdfMFojbWyuxHatbTvNdDaSQf4rvTGxJpGy7hdjF
pSmCnp2JRmzRCzKMU9IocPu0l2PfYxsKxTQSgky7FYmmWuPNbuUUkFGOPoIg34DHIy0XebpgfxT3
xkm2Y6SufaskoVHUuCl2Axbll049ujcy1LUKFLQ5U+fK8QKi1VsBo0U+xJZIsamqb3ngjG+Th37Y
2smSr+7Q2nqe/qcXOVk0lI/zt1/NuZ3jN6d8J+KJ7WxTTeNW8VMSDvihS0fQCp947XAmz9imvuXA
UuH/ZXpOghqnVPLt1DmFsF6f2KL0Ql0ojE0xQN3fchW510tKm11itdHxT7Lx9QnGLFaINvTNvHBW
Ov0D4skLTZwqqH8h7eb3fmCiXjmuB6uQRA05wf9tUaMvL5gL7T5ptit1a4P7oWqi6Vmth9RXBPL6
btmJiSL7a1yhh2SvAP8Fq19OgtgRHBfHVGgbr7twtNifonAJPOksxZVxD9Ug1kXCLPBVhvocv26h
cLy29dO2PMg1QL+prL9SWdGk0ZIQeRmcyyknnr7a/ShZq1eAEJcltQb37Q6lb/FrjhiKSG22iJ2B
mm+tg1Nk3SCXxSldCJJlZ0YoN/gGgjihJkd34QuK+deHlCLUlq6H/upefmnrhworb8KuH+f4sQcg
/ZnJnBq73K/ik7xaZRfvyBKuWIbUJxdGxvufP5DqStBAZvkUv1PhyUe1B3LVF6IYth643S/F4DhN
IkHi5EMUo768hw6fz6QDJwGftQCJCHEBhh1XZ6eDwWP8j85BnsUt3zeVpl7wI69/0Za0HYCGQ2I5
CSvieCGRMA9rGDPvY7jeEkFn6hou4NS61m8+sv4d3CTQFnRjG/UmLKQ+Qyksmys9KM67QjZe977j
wO1INaIGzcOj8mwjejdjdosn9WOEYMYtYjZVSvozR1ZNMGqV9Tan91PpUOEHTnv27exENODgjvqS
WSiEQgDTu8WJuY511rr8W9qpA6E9U8+6aPatHmI6ti0upTO99kCyLbDK3wzvLY/gIAs0Nm2uWDEX
dZirUpPnhCRX6hvPZCejkqXEvJOWPqJW2kAob5SyMiNXRJ4Ffc4bBo/w5PZj0I4fcOkOEkc2vsDu
cKHcT5FNQ0vBctvQo8dBWmamT4Iug4HvwvJYQR+HZvalz+Ti4YLw0FsniHinMsLUMw1TZX1gXGWd
4gQf/oAaZp6SRHvQGI5hi26KKX67blv30rd8CP5JpOSMm31bF/Qyye7z8idk0EIPWXrVpia893Bk
XDJG8rhlj7V6UmvJHkt6etZjCfgNsahfx/ACFOFTt/vQOYvSvs1rFAlnOQtnIl+m1bunAG21ATbP
cx2rcmwfEvWDDLDMnpkmAi+DqQ5DtU9h60VfO6QT6Xz34tkhVrePEbbWqqhb7GFGNh/TuqScvKYe
loYfAV7ps591kc5jN1zrfNZlsTuxcNHLX2Z7kGRVaKaTyV7aXO3DAzpX/i6i67UnxkhHT4IOZ7WF
WUVV16gTAKZiws2Axe/8G5s6OMRWhlbS6x2qB2A06g72/Uvp2xbXIbhjCIpGopcmst7Hr86/lU9A
CuCcAjKoNaVSKoApVm6MmcdvmNCH8G+b4P1fazBwTmTOB+kPFLcFMV3FCc420gZFTsYBW96c0GH3
G7EOpvHH9b0H7z1GDNMrZtU/hSk+kFEvLE+IywrtS9MnwAmwECRDWCbEAtZA7dqr/8T1VFI6p5y5
hvlZqGG0Z9raqXFVryjwLtuhXZ6OJf87ZzcvWiS9fpJNawSMorEeFSV22Lod+8mBx0Kr3TBPm4dr
LjzIs/kYyxli3gOz1FkiYEfJqevwmFEAzyC9yagQr6LMsdqaTZv8RYl55v9hKLgMW/7xhY4eGidx
r4U65k4vRuUWtc3AuHS0RjvEMEIS7w7E8TLqnbhKMnNttia464LW345yFeGkPN+/k2kj/4ZqaJ/S
EGM206oKgnn7oTX5CT2r1fJv0DtMzK9HOD2ST36wvcXIct8H0ERZmOrVhqySRuACljPbGwHQPjBb
ABA3bDF2Tsixw+2Gyr7WTmHLZp5njujpg0FwhIsmI3igK6YkMaXjxolGCMfVG7MNcR3JT/2xQa6r
L+wY5Zq7Q+s5mtUtcpfiyRto668OdAXWSOdjSPG/izKdtTwrd6bZ/XzD852VYmZ+/V4oLpcPUu6r
Ne+x/ZRGOaPXuURZQlIaXO2hvybbn/Lv83LdeLV4RzVJXDyMJjr6Zdw9W3yeLHqjnAFSHdnvuudV
1Owrz296MJaa60LaCOHV95I1IiUsYUjs3z0b2Zxcx849EBfC+Yg2sFnLln+g94s8tOzhxDsUY+XI
KR3VWcJfxzy3viv+JX+4X2VXmrEVzLk7HzrxlGQfYKLfXFanLiXADNOuETscJ6Xpsk/5dUpFAbeJ
wslwRNPlnYfI8Ve9HfaJ/BsuUKDSkVeaPqHqt5qEmXqSQjuq9guEJltcwR7QBQNQnWFTEmgMLPOj
+qmjbg58dAZFi353MAl4ojQ9hhQ2ST3OrEB9LgQ12aNT1xT+Olf4eDtp8xSLR106zmLpkMiWxnzi
O/gkMpLPAsr95mcD87pcEe6JJxdV3vuBQkfZ4Es8fYFTtagvUBqpgw89EneXOBwkWFjvWhhVQveF
AG9K2smsduc9B8tipHA3hacRt8PV0WtP9N4qYqXTNiEfENMXC1M8fOeuji8aiqnZ2fKzVPk4grPk
BRRrPsqNfLuBhaBIsb2yDPcN+M3yzWUMtaspZ2/kT3XLexag7835WTTKxccKQTll6gcaQ/IKIgiT
JkDf4UDKoqhyeg/KY72sK7fiFvrg7WtgDdwrJNW9GTn5JlIu9znMG5L+/fOoGR0MqiYFDiBALURw
fVS3ckcd9z4XVVBmCH1wz/VHiQQe/sQACx59QKVgKWMRxbSi7Tq6IO3e/5nlAF+Yj7Qm2zccf44k
GmMiy/8r0/wX71AjyjygCiTH/uQ1+1j90SMZvzyY3tYNzbaASu+obg5uYLbWLmnjzVvcBnBBdbaU
0AX3sqqQkXdp4vw/Sh5/j0+MDak4aw25Be8JlC5L+/oUrcN1M3/sAIiV4cCh9Yw2k6U+u2DhRjhx
JvaZMrzt4rJ2W3keIs4zq7BaJpuQQbEl0nTMzdXTcP+eXrxnMF778VTVhX/Abd+EZNZfj1rJg1mq
gFgzbGRJAfvuCyPPhdKIeZGIZXMRDWKTttPoObA041LvTv3HbGKwifVhDSOr4hdV9ttaE+XMSnhd
70++TU1/VSIxAgggoK7ITdZ85EUmvt6sJQy+TqJEZGkbydW9E1o7JTeNuC1XUZ3x/5Z3LnoJBVDn
kbKsftoviabr1IXa6w3enAbdGvX0z5in70Uf/6+2TL6+PzUOT8nVmDeRmIUCND3tObzw1/87KfYx
1GUINXN/zusEDJ8cuaGDboh2+/uTlndzE3F+0aOC32G/90dPFJncrQLOGFAPOTlkippI18CTMr0t
SMySsDqyzvJhpEqDR67RWsONs4aIPARQolfXGYftd5uLXiUrd+kBtbeppjadaQlp+YcOWMAZrOW+
rBGfB262V316iJ5ORCLc4XKopuOUu+szE1qQStZzc0AOQxlDNmZB3hBajXeqVC4PtjeHBJ+uOEHL
IV8eJx447PnpSUlK49UIPkowWYyAwr1hIB6Cyc8wijIWXzy+az/cEsjJLhsasI0bAFDMK8JQMjlo
5rEYv2PKjzeRdlzDpTqbaWC2XNJ9+x1wEhbc0LKKT5MU4yYZceTlZU1blIiFhWnJ/CjZ4EHRLnlC
iiHOBcA9aTriCy6cal1FrlLWO5/sVt2eA9AZloZQ2eN8mXQGAIOOKNZVPJBz3OB/RqJZTCHvxJt4
nBhImyyOXhXdU0GrHvHdinDN+Y/AQSc9w3AR2ApiGmZrowPMB9MzRYlfjZpkfXFCEeGsA1+N1A1W
VXUxuJ+UWmBkRce708SH5Xud/F1hmOwP/a7zuMkY0S1RAxJp0SRC3t1itYlN8n2Tck/L0CtXc11B
3oJSiMIzXJvzcJhNh3yKaItGKgrqGg+D2xZUPFVJ84bn0RDjE0myj8goh5WWqiMoK4pwUKtc/vgu
yre7UgWDQGxY7VPxHH6M+k6ZixqRkwAPT9G4vP1Lj3VCLPV/L682V8XAMjidmJMMp79pAy3aquly
lPPNrVMhRTILgKkXspMbfaCcflpSOfvSX/PC+UbbWHLppppZ59VGIyuL9GJDYUHB+QF1dwc5nNxJ
8vCg3D8bgbcGpZeU77gKdV5Hl6snzYujub0em+XUEEBULHMFkTWqjs48+gcL3av28Gvm1LxHKbTV
RLGIIHC1TdRHDttT9yZRFcMl4bkbWBUIbR+AePQ4hZNmDV1pe2VZZrdfVvy8+Fd1WlRFgqvChP6d
hTqlT3833fQL8dC6Yhr3/rRdbwNw1kBr4QQUc1YlQWdvzBjpuzTGJAU2qjbKjZDmp+jMoErtKOWR
GRl2TYn9B007T99h8pa/5T5wFBcoIzq+66AojGp4S+C7BNhLCGGldT1d6Qv+nBK2HyV3bGPsySwD
0UW/A0TfHRWC9Iw/2bXwf+ebTUmvEbM+fcuqXVnFGzxPccXPgH3a+sbxmc/EUDqGFEU7wdHAcGwh
9YSrf2E7Kr1pqlX6HdRqQLVqhDV8J7nuCyJ+oacRvNwhqdxUbtPIh6sx4qFkV9qKrqWx3GOWKa2e
Ne7CfFvLzLWAbOgq+jLOW9mLb44N1tRQwdqtmgSkOBRDgPOVthmoitymSY7sxWLhljrRwgvuuES4
vs2zBIrvgXPoiv7SCNDFwfaZHwEIFIUOLOeINlwfa/9/uNa18GCathZ2mHn1zN4DVvH83+4aYDWD
MRKLhpbN4Ckn9zjP56ugxNiINe85ZccXe4dEkItQIc6d52obrqL8qgAf5Ta/Q2hPGBI2EjfeKuQf
kwQodD5i9u7xrGZq0NsCh7KLJgWpCb6YG0qWUOorRglVwO46wn9cWhvyUBD6wjAr5xWFsyR1Qk5M
6ADMVdzD3esO7zjaBX+kZEqHDVyIaOSgCSrKSUh/ovWZ4jZ/Lr34osO9pcJgoZmSIYRddUgGzEzo
wHBiUINTifX6lqx/n3eGkDdU9sEotEi2bNs1qqQPwDpruiKBDC7+WoChBNyczLdHvRsBjpbhq9gq
6vW/xqWEkDlI7So3kwCRBzsnT+B3LKdWGRcwOcW+jK5BS5baMJQa507lZro0PDqCqdGdLLRZJnqs
Uywzo6nPEibMHiRS9McMIFxPHbiVwt2b8vcwjL8Iyy44Mv4LaFK9zS+EVeZOadSPpIR5VCL9zKeQ
SEmKr+/F6geuvvgnAhntiD1HJVzZUnTNnHZYcubGGtbnNfEkCIEAWBQlC7WN7qJupyOhYpSChzDT
4jRue/XoXaPm2WARufhZNVpsi+Ih1MUY7EMIAtJ/u5eo946jpJohWpj2sVA4P2kcfbH8dySXESxg
PuRNYhm94owOmpI1UcyvmGM2KYT1gFzXIRY0EcrtOEAlXt7fLTPVRg75OIWqnnYWScwzRmYYRt88
mF/XU2iYmnwvGAFUhg48i7kqXn4+2im3b9zG96ynTPrNZLkWiyQotYB57dCKo9nDn/LygU8RS+qH
0Ojb+DYKlCOsn6FC6wsam7c2wqYFU7uuO+ruI2aJZMoKBpTViQ7yMHR0Ez1KYRYs2hCQmP6Cf3CE
ntv5EThGg39BlOzHFtynYFZnukAFsRBVZYBP7+psUkNov9B89LNkrmgA2gCONjFtPpS6Rmtuq/PL
kM0i4yJ4wkFHNbE8hy0Sj6mAWuEsjbMu+KstvuIUm0HBJo67QsxVHm0lgW0yp2OmMsJMeBJqkz6J
yKwfryXgl14tXXg6Yf0nTxiRyicLKHFoJ8HVFXywzAkwbynrlc4ec+LDRtTlRjIrsqSJ23aHYqbv
fVUKJIx1GNxZquIrL5JHyvqfW425JdNWWV7M2nl3Kj+Tkm/HECrVuzTx0yEiaUr637pU0pK0PYCn
ES911I/lE08ANLFJecQSSjwBCtGeXiBbhG1nMNpHQviK3oUw6Pfl4q1aPhJbarrIKE9EzQghB6ry
GuyaoQ33oioAWRzASfzpyvtjBL4rPoa/brYjNzNUAQ6DE/JeiiBriHT7/+G02JBS4AZMTwCvVvbI
DHxtzw1q6FEvc2MEtGnVj8Lz8d8LKZ8SryQ+BjvazszCexXSWeAWvVYn29QECvMcS53wPlo23wcg
XlAOaM7kQdzZrhVSeBlBJpTf6NJoffp4Vekco2u/DRuDOXdGo6UdtEUNzFC9whxYryLx0cJXuWCt
k0MGwzlceQ9+mQJwOIHRiqSKnw8R/8sv4y15+knbRj1ruSRmdtBx10JWyAIj09M4o6kX3m5E9bu7
KiYWHxVwxiKg4GVGrXMbtoT7vUVhjj9WGzDdSWyQ/i9oyIXXoRQbxquLP2MN5S/2eYxH76ZWnuaX
HGyI2RREYeg8QhWZdzef9c5ahDqxCE4u4TvXbsvRT3ib8tBU22fk5BFu/tCXQVww+rg49XUHWYtx
B++XtpSfY7iSOJUJhZbrhlTKrKyx2fF+V6iInefvlEdpWQNg4sRpNTxUfmdFJg8Gb8J8soGiA11J
1i931ra6MPlUPDh3BtDl6LEkZ+CsH9EsRZZsentEhfwY8KdtZaOK3bfyXndoaXbXKsGwOdfruItZ
ys+R1+Nko7dJzoTgH3RkRUMwBXEbdoNjjOvCcwBPb3Tnu2vP6M+IPUDR+HzzZZmNJPa2h/Az5Ggf
1mTycluzL0/cEsD4A+ZaQOooYPFP3FwNc0AtlRavvcpn7iPkNj9udITxTbHDQNxjJjnw6R1FKncm
Mm0A61xRh4fcnUu1YmZs6QM19g+syLErQsbwcAdYyR+9ZZY1eP0S9JI8W03XMgZzDkzFmgRWrRTq
xzRcLt+r5UMRGNyBsSi/WFJyajNRVtuVE7PaxLtEG1en+RqvS7VoGaMfdIiJQMn/PNhFqURrRrvg
sff6n6YT3yWA/B9YjjicVEheAhblmsLGd75P7CsaoYLh3KOEfPj/oGyF/qDrAx0EEqqFS7eKKgaM
q+7wWlOdpJ9pmE42QFoI1Q1e5itTH4RjIWKkL+FQVN8W0dEjJJsWNqx0GtCW4N5+FRqb02iJZsJT
hc1wWdCuozM6XiusM4Ev8ukXIaOIW6Lmthgq80nG9HWO8TLLDNW/qWf4dczAF1LddPRla9m+v4TO
cIjST/vPt13Mm9xp6cE4EYoOieXj7mtu/rwS8eftWNyt1u3mXJmN70tva3xQLlLWDm8nxdmChqns
6sD2jn3s3Xt0F6r65mUP21Sy+fGg8FsfXDwhtzejIsm2zhEOAjdVVBumzWvQdy7Ce4TqlnJJGV45
IqqU5JQByvLp9RK9wi9HuUl89si/4rUJgNQ/DtQl5YbxAH0c9F2H+ESM+Y3tpBlFTdcKjKwoICtZ
uXkUvSekpnszNSupuyfFA7iYSQ4P5Os1fZkC8NEedOnBdL/+1OMgN6n7AXDWwZp7T+YtX2Xcpu0o
8/85xbVzQ0RujFZ6nliZY+o+sYcIWcCkB7mWYvFVRGRImdyiUbVRaSHbLPsgRB8clwiil6rIZDDU
AqLhXSJ5kNY+BWy0Kp3I0OPawpbe+9n0SBXu1xj16cLFN69rjC2v+iYpEwQLZbdmVRrvQBdYYrhq
rew7IHYg67WFG1GZM0fhx8D6sQLBOOEGREdUU9Tz5V9Rn0uuZlZPoaGlF6Wh5B32veyug1zY6Zja
3Jte8WFaA7Y9XyGkhOahuFyKc4xjB39aB72iB5W8b3BzOGC/npu4KVaS/RGWVJo5MnF76bNQkI2i
Q2IUjYYlDz8hO2XsAjKApUWaBYQhjFLr5lj6nwoSz5vp8BEqLIHdDadVNDkhEPUBxXqRc6zuxxlP
O9Q9g0KZ/R7i+b+QyQ8rc3nxMeq2VvupN8rx/D4ejmVYSih/BccN4z8My+tfIH6qMkz0HkaKODh5
h2eOQac0HtmFxOnlAJALhHrWe/K4OJ04tnCR3JzCAFSAEn0JzLqX51OLHCt7LhGmd+b58553YX42
6OYq2mj+ZAoCFQQFk8ubZK5wGS37qlVflDsz06bl+yG4+1F31l04VZo/RqvTUz2npKqqneiqyf7o
jcuPFFMhL0k4/ud4AVaMP2zGHxgPGuSKIgmzqSLvRUObHSzjWyYJAiaB3MbD2qRhqDdBVRayZrsa
31cFaK2CH0Zdh6uWlRy91jkmorxK1V8t4LdRfqDUke1ckmGSnDckqfq1UO3pheEw+w0BOvrexKcQ
CWnGjo03qJj4ostlP3DKaen+t4b2qIXb6d4YkeCrXjOM1s/9ByjRU/aLyz+ebmbh02SMXPmAuJzl
9EzSqqKcd7cKgX2Fu7M2js3fu/EmST/YMEpK2N3ljB3sJwmWTCFaP9HCgA1ey2x/ShDd7V3DYihZ
O87hyZj51jBZmDn9ypqtTlvVahix3T2RC+eyY1/X59bhrO0XVgTgC4sCBu/0UnhUg7rPzmLPZTsO
dTKLp3GyxMxgDc2b/ff+Hgu4aqyqk9VtZnZ1ckF57ytcMGhc2Rtm1Uf6jy2VjasmnfUPsuClVSsq
6ipcKPOiAtCR9vH8SpDIh1kXsT6FSYkcg9IqUZfXgdhoR6pl5sZcg3k/qYlmCpFcI2e9gYlMHvfo
L1xSGTzfUuPScrcYlF6ImgBGfTz/6kdePEQMNIod6DLzWN9iTkoQJI5lQFR2zTmpIW3u4mOZlF5T
5pvlDoEnGnUV4y2lWFoHegGgNGClJzI8Gn58VgOAtV9jksQ/sV0H2lC2AATtOAO4f6BYXW3rCoJK
B0bnzmJjioT1uWkoa3H64Qri4wYrsnj93fUBAi5rgBQLHUGvXM61eLDEhowS2wz0sXdW6mHkgTeK
nvGSVWU3nPNjiWlnCe0hZLR+M/DeeeQewmlp2vHsB0ZzRq4wQ9z3GpbATMpTHS/HEOiA2OyKUMAa
dbbicHwqHJqMNAUNeWMrloa/U3wIwqz4euKUNkDdXr/c4pYdviGpQbiB5ngCqsYls0iloOH6OtQj
WR4aIjCyXHqpJ+q5Jm+BFmqM2LftCKeSdQsb+iWgFVSMWdnHvunCagaqz+uR6Gk700SRxy0wXfyW
J12vU3GuF+sXp6szdze87NISBR3lD1/fp3DlbAJ44kPI8be1pGWm4EUTNFBanBr7JeQ5Ahrz5Mu7
hfZFfZQ1KN2WGX3wIjNDTLIRPuJ4D1/MP8I6llXKhnJP/wygSmqxWr3a92cgCoC827GjTJ2ZHEpQ
obfYfNQHjbvUlsBAaUPeB+LHiGEjNZBcYcEHgpdmbnnGQvAtcbuPMnWfEvaQAd9OP01SknN++Gif
xYM7clyijDv6VGX9V/NjDOGor6MXNDwfHP96/hspWf8zIsA1ASZjSRWNDNIjThf9bTa7GpYd6gSg
huWVDowaVU7TfXee6KAHEAHho8Xx05VWmmg3FXUWbSuYJFLSZAPafdaPHVv7PWTTomaf1CCfWynn
n2ZEuO8clum5rd2sR3Fz69aqIK6YIJnQfGs+cf88TQGa6P9TbQ2hF7mK0njePX8NPu7HFMhyfQdh
QKQC4T1Ng0Di8fw8dE3TBi3Kk4cZP5PGtr+XxDI7QfpZ5UKcDJWJA+C5zCVnWiPaJmj3DwTyBsd2
EnmCC1Qk3+ihcAGav9lq29QrW2Otdy+xi+ozkbCuH0mCUXRbmwgo2G7b8ll+TBq99IpdFgjqt30t
j5XzcHWzdzwkjrUPCTaUevvBiJCRolLO2qMqIMnDps6gfYMHdjIuUqOSS4WpiRiQdtNRq/CzK7Ht
4vBrAIHwIJ7SqeVzWoWfhQy8gtIcN1TrggP1y8n7gHgKre18dBe4Rjzsy1Exga0us/YLi51T5qCV
zUJtOpeSGHrxH0KBAABlz3Yf44mpEgVeTlpihaJLUQwIehjN0/wj96+giFIib6wEN4dVKBBFWUFC
/L1N+bkwGuYJEwhz2NiKWezCYjTAIU2ZJvqI1nfM8Y5/w0W7iu8O0l0oOUrfZfPX2+dS3jIghTlE
qkiUJVJoc7JBsO6ET7LZvTj7dPhgaIrhDbi/KJfv6oqNhELp1fYJZ/eU2/MJkSYdQe6aVeVA0HoO
O/o274mZCxTGvaoqTKpnFzarGfWChn6CRahewcQu+28kwFnJ4OK5bH2+tKOhXc8DGxquRVD9B2y4
NOEo0OWn3VZlZzbHHrZVYCgGTZU9GeyD8BxCFCV9jzm36mqZrXqgUwiyf8hI+Ore5OgNUCUqcoYe
78Oef9DJHazWerm/cCrFpiwLKUOmJaR8mWnTaIZ1SeOVVCeQ0QgeDwLCVgTJqgw/nX6hI7GphpX7
TVWPr4Q/PN7WtB0D5fQHN5z/t9Y0y0sf8gpAefRSQ2YWv06Kn6uycj3v3hSL75gHglC1tsPB3jxm
1f6JHaHUpePLRs1Kd1rBc9uiW/T5TFL1iUQucUkmnSnPBPpnvr6KXptZYcl58Dtn9bCQASHiP043
ArMVx7f4dzg/FLiEerhBzqTSDmfiu04C3hXzvbVvhtZDUqfVbLxR4mzTx3dm9Y/0AtDnHIW86GCV
OoBlLnFXLm1WgskY++L/qJeQqGBzc1r4ZFqwbrdGBYi0y8lnRdq/49/ir7aStzFPKPGlZGyr4bKq
ng/zpJL9a7RqFtX7eso692DPFJftkerW1jLKvZv4xwAP2A5LGY4OZTRjZ3OOzdUyV/4hFTScxIKu
uA3LXQBWTiNquphlf6p39Pv8QVRrdMUiZDfX9p+Wh/NZIOoEMNtn0Ot5V/kwuYqhhTbY6RJ0uknK
q9ZU4BWle5LOAxF5xhOHext6+ccrTAx8+JetEtQEmXhr0o6CBEQvUt1DS54FEkJuJAYl/ybkYIIR
/YtyOm45G2EhWFyvjoLoXvdorecEUL2mYBUgyBg4s/joQ4ZkcsMxW6KmRMD0QR6dJQIWAtoCu49T
Pnaa/Ku4Q77nc0s2/Qcp8WElIDc85pVcHqxi2W4Fqn/OtwjGTDJUdISJJhNGg73ASQpImUmBAQgR
Lal9YxIops/OYhJlhAznlkXlLwQVYK0jnvrFewginSvDt881aK9O+TxCcSeyv50wTNFDnkKcdMoE
rmidcj5/NemAKyAfrpHQ5RCGVR9EJKXHOpH380EhM5kqQRPqMZJbuW4J3MWiZRVV/m2pY+kTKn9a
OA291SzdEUCOS3doghyGTtdyHXMka2cXAgb7sXZ23lrpio832hkd4h67KrAxCNK6LedOTj+9wt4K
mjW7Fdu4ZlRlbozjWvpco1LCpfqrxT1ZxnQEo2kXTdNUAScD5tx2uSrDrtyra81NuR5eBz6dTkdj
VuZgC6imVd7Qxxca5curB426ENw3X6V7M1NFFBMuUl/R8AB87ga7KfW8mSglYnxfXzWXz2k971XL
DT81tkQL6lE4CllRsKDAhsg/JT3EE0x+6IFlVHM+uFqJXLCCZhpwMcHtAOCMsfji3y9yTCkWk5Fp
BsXPsAlZDglZX55We8Hj5eQgEts1VLzPZjf315zxLAk1qybtAP3KABAjizji1tih3jQdz0+LbqRF
u/YCiH+/NldIDEbOem29ffNSMOm0fUXB8HIxjQPD+ZlZWSL5wIl5WMGwQ/l9xHWO4FViJUCKGz73
GAt/qSV2NkoYjzXT9l6sWS4dZGXXoJ9OV2KVe01fmNjfselJw9qXM3VUJQS9V90ictmRk1N+vI1x
xdineaRjC2cCfbnVeUP8KR4+H1YJW69sxgzvYFYQG0KccRyAiEjvy6hoB6DJ87PP64bmudeUgdDE
GxicjnURtBzvVQhGLnb6Hr8BCJVkTZMCKd0WyOH3elyZiuVb+aRPGeXWqCTmvypYBS6qJJkSMAgS
U4EjxtQXa8KZGZD6xwqL8H2LxE25iX8ak/Q3uVprarCftLEZo/erPDryd6Bocvg58wFbCGGl9u/V
LS2wLkCfbDcE/aWSCWc0u8ewwdGzjeZxiqPeEo4bL/e5Fq7DgiMx0/zFpaqQLX9byI2PYIbSOAzm
PkntIdpmSN+oO7Y0oiAQSPjup8ZPPN7eOMgFSMoUygf30+I4BlqK9G0yWN1gebpHwFaZOeOqbyIr
9AvONlD1bDuQ2wC4KnC3ETMWNOcnG6H9ss7g/Zf2ZSAtr+iMO7FSIllVE4jn91S8E5cZP33qJlz7
du0fEkdXNWe/k5TVG/NAg7uu2QuiEIC+qmF9ZPUx4HkYgn2Qh0T1B8u2wyOayaztM3n/LW2BtsqV
zs+n5c17ONcnqhPzsDVZMv91jEUP+Kd3HXYoIkpADpknuN7CkoI4PlYm1pgDaRAiUxtkrd+pPVg6
IDS8Ui73ZETCAkWPaGJQnAXtKmBbPbYhX5aHnsOCuf7n49vsllQu7or/ms6jTwrhljg7Osa/MiIB
LG/RqkfsCO9KUPR4qXM5GqpHkZ+iBsxU+0LPrbLgTdICWQsUT3q47icGVQ62DHxG6bKMV3weF/CT
BB4YOiHL4XKl+oAsV1B137oOM6waxYHB1j3Obpbqy5/4tdKvxd3DnsqNGt1ocDctPJh3v6WJDUZQ
jDkDVdbfWmCeL5Jj7zHaho/TP2iTngq9lRGZDB7j8XLPtxcRQjHuV8OoGiHkt/DepSzjqID+e5nm
B+iIGrlK4roKK2AIpraUHJf6YckJK722xb34vVPa7boQkTVCupgCLLd98IYMErBR8K9JtUj37HzM
BT+bKaqRXppGwXAsN007UFyj9ZKXwkn/ca/HBhZgOsnVlElwLZ5+QRZ6DV3p13iTcFUkdCCcN1Yd
iN7jwQF2TQNCbnINIGmrbZZPHOucwZL0kN11jdGMNuh6M0I+ROxzEbxtcDBx1/8eAS7xfk+XW5h4
Us9KoQQgCk/m+RYR+VeHgnoxoLEiSK1EgnBfa1zsrs/b7A94STbH0yxA1Uvijbr05Y0JZz0Mtk16
aoCuXVk2wSye8iPP46FdS8NlfJCcbyo02DkMucLsHcgiO0dih8GMiYIex1wuBU+38jt/xaQvvWDk
mYkk+LdUqkM4QL8W8x4ivnPDqW4eBd5Zdjh3QALunu8LFYmo8kIe8zP1ddAbJoyterRXaJIG6ZpQ
MGBwE9u0TNevdUiJRhnx2R3A5ADkRfsPN5fyx9sfk4oG5+mdK5Jrxao0KvACXTFO0M8FRifh8WhQ
G3kYASyY+y7bLFzf+WpdHS5DwxGYzWO8a3ikpiLKOYkDOTldvY2+3IFE3anbnli7hvmBZqPaKttg
nOhhT2J5z1z83wD9uzhIlJFXANHkn1JV73S/2M9uO96mscHNBpBLsmXBwCtgku8kzXvmw7Kzflsk
EkRtDZkSfFdvixiLcmsm1p/XJL4JI4wDR5fa2HXjtiWuCAY5RJqshewYjw8cu6zK4l06qu/OQzpO
vWUbh2Kv+Xcs5Y32t30k/FRsh5gt8mkOha+o6tB+f5FtBJ0bVUHiKwtYhsEAs9LSIamMORbD4hSL
9mxeSpSLC6OYtHcdlavo0EUalTvqi3gWQDUbGwqZN6inPCzsdu1kRV6mVqAnnJGqffVIyHWxugkC
gtmmg9+T/Kc7ehvR35Icg2szgd7rhs+5GXZQQjPMOGMD5A7wXvMLPgAwUMUCMcBTTzUZ131Uf92p
7ZTDFh/5SDPg6g5VjO5RSb4A8OAg78un1CulLxFe8zkv0+IDr2zhnL3mQYCamD0B+2eMcpp7SRvK
GsRvyA46eO7/muQWowRJLbUkQA/Hte1GNIWDld0GcAhbGO/52ZS6c2ZQUBphyKcgOaXCzTiaoP8P
Nk5BNz4Ar2GqpuF7irmt6uaZkq+l1Ct6qANK9ZY1FIVQVzyCWaH72bko0bRjUgwKjSImzq12E2p3
Q4GIYfFtwPivqLO3zMK4ol0zzxCnbQ5LSjfFu7lQ9iIinceNHDsacZ+tXfrbmqR+o1gduSMuxyDu
e46AIox+xmXAu+qZhqiwoXUlBpl55RHxfJVFD8DXi2x/TIuwDSAqX/UMH3FhDufmca5hgsOZ7CBC
+8emKu9kmwR0FxEboXoaPIB6eW6jqc8XNMfNBe1DQy3yt99Jo/SwUjkQnb6ueAPlBi2OX8T+43C+
QgYPgz2ZRWAqOT1BCBbeWhSIW+WgnV59PEML0bIUQDPSIOtHQfcS1hhm3JleZOc6judyjTxblK9M
OIUR3hf+uBe13L5h2d+uuEP+eyhLN+nCuASgmTJRDjNUGzlzYOwwj4UB6yPXOIQKPRfxBlsgDz8j
0j0HRZnbHPQTmzhvjbwV5E1f3WIrg7eH8S4cfHzXFHtXtDlN/RRjd2phtTMA+CXZPXtEWYSZcs4p
PyzO0Ty+WtVc/EnkyVVfMjFUb7uRi9oE8jRzgYnZIJlb4oAo//CUgGVPTg/glDa7nYuOS4Nr5SZm
TGfzVpHi2x7SjnNhCVHhF7AdDQvoEeSxcKvA9vM+S+Vij0xeg5BoO/gMZtB5YVpqa+yqAYloxuNe
jQ3d983NzlFKLKbsurERsmFRD+MJyarP7N1fOK2pUPhJUXFIpYeCqXR7d4uaSS83KIDHHuRQYNOg
Xp+GdgeK78QqCYPodIcKMFuMxoxmxry2FhIVCwipi9Lg7rT0niQaHkKEEfVdzU/+DfeBnjStviCs
zzErD569NzIpaQQ/4s5Ge15lu0fNQMRYTbp8aArABQviSUdR/6OAzggUOxqsh26IIXXKiNPn5g9A
42yxPlkVJZvuqWJAHe095uD/q9lQ9VEe/MMSIvrTiIJp8ZgoFo9M0p8LSThP4hlA09MvN/HHd+oQ
xfsO8jZ//OezhjczlSyu2kYAp5l6or4S1zjXgPQ+6n79VtpnHF7Hurj8ZFSTKk33f2fZjZZFwOK+
z3lwPe6uacjD3pK9uto1B9wi2XsnN07Is4TNlDOu3gXOJw4iYAUsdnXw+jzbXTt8VvMDQwc6kozY
4/rsFwd9dQ9oTGvILETMMhZVEGMZHaT7bH/POq733BUQZIcDx5QrZZdjmi+gelefLwVOgmb1Qiw8
zqUVM0Inr/8UBO1VT6hhDBwi86E7TXojHlgme4u1WDWk222DSkkyvd4U+4zwL9MqKY+ETzgJMyph
cHiUTYKcshSpd1+U7d5ZKUxzP2NkoBM0N8wjCYQVWOWBHqPFNfU9338BPbyM0MKlbiEXbn7wUbeu
RAvAmM9OV448snn6lM1H7r8RxvblDTUACmiQjLG1DYROMrR8z5uKRfj1RuCpvh1o2rlMqrW+0NOr
Wm6UReM/NHkjDCyMrNaZ6QxMF0rB0/k7LCAnROHpv2XbPO/Lf9u+QcdCQ9hWlNBhkv5j/FVdTeCa
5oeaVU4riptbEZboUoh2IRgxKEYxmlDaPTQKP0zDnk4b+R+KR8UcuUivmzdbfQ+N5zus1bXnSZFS
5e5XYWaJSrHPKw99CkVc5XTkgW6QZZ/E049en1MNhZCB3kVk+jWPaoi5NOeN83ba8fG0couBe+ZG
FdwT3O4f+1E2D30+BubVCHwRz9jXyr3SCMpif9OMhhXe9f6GdQuZSadrtqyR09YyCqKpXrIiJnVL
lACZXoUqfhdifdcEcs9JEgE5t20XvosMlLgo/dbu26DEFyXKEQkE/pCcrAwP90KojRAtckjyD6of
kr7NZvniCHfFVQQCwmmcB39PrG56y4Gvbd7p3W7/v3QCOVzJlaP+J6vDPutic5HH0pyvcwneKkRi
K0uthhj9FEEHv0VMfVZJElt6kbkYin2vxsZs26GfvHY7abIMLHwALpPADJxXuVYxcYELnjDjWARC
a8pBIBR3E2BLAGfMSNrTbGfNhHDLo3JAGpMIVP1MNqa9fBhPZdcxsiAytmEX1/3q5ACo/7+y/0Ii
huu1WSIc9fZs2l463jPKa6z0jZrLJo6Wnm6uNQL/uOyzBgalvp6h97yt55Hm3h8qKVoEIKMb/BGe
1WVIo03DMDajxyuWKF1JRb5OFbA/JLsTv0FShBisgR9iOCNzyzNjBGB1I9HzAOBH+YKWD+G5DAG2
47p2i+URGjP8RtPb3pow8QSB1C0VW4dniqtFmO3X5NXOsE65p3lxZTqF7gsBfwYDEmSZZelwffCr
/+Bb3qLX6wRnWkipH5pOQ2Euv3OSjNPvixBwJAezAUFvdVBqjTCwfglSM3soXVPmVhVVp9Ye2gew
U/jR0zAz9D959jaQjoiPVs1O6pp7w/qdvz/ou9XeJDqblUX0ItHTzsL6HEkrmO/jcVd1RW05CK0Q
0SirivC0kYBwWh+deSWkwKcLSaWNB7yli9T6BU/StHQyNtNWGNaMKSfvfQq/aBhfb9SERScFAXJS
PcUeU8LW2cU9fX0NmIMqcey77Oa/HELqMdpEgAtUVGbwEDj741lPB8nJRMXQo7hYiEu4R/pOPM8N
yzyDBvLSPLb2Pem/tcKHVn1wr7AY+eV00HwLuLiJdYMrT/VQ8VLBPM/Yxf5hMOsu1FvbfjRWxwAu
x7FSJN8BU5NnXwvig/YFw2Qxd/atM2iTpMRSK81jP2flr3S4IZ6OK64xkYSaVnFDPtvF2bmaUKzd
mcBuz6p3c5KpttrLK8W3g7bSUnTGfTLE5o7MFSLe2K1b4zD+O8BYE9Goe1xy9n6hchkwBXxeZ/7m
vDHDMeGb4gbmxAkUzo17+oGRANaiCb0LQqRgCdf5AB+zJqeNfQvt1kEtn7S559op7AH9aize+ivD
Lck8IYa8HLpXTIPZpY+lGRCziilVuAOM28bLilJZEwaY+UTfEbDgasLGWKg6Bsmwld5DmgD6TuMk
qO6ynVHf1vszmFPnDehsvkPDaqdQTSDvJsNBxyDPfd8L4MKNhDXKN4RS0rkA2cQg7BLezheJIYGz
PoA4XRO8/BRspj6Yu69CEu4L41h1nTLFCv3RUyAEAYn498qLpJalHRu+W2Q7kL7vvOlHq+lEfYE5
T4c1dTLAWCJMbptrpjBZPNl3fwxtssck7taiDcA6KNjzV2fx0UhmYGPQzEJ5kV+YZ0SOdx0JRjyo
C8LZxVhli5wyW3NmUVpPN79Rs8cuyLRv3bqR0A4TYwrlf54qGUbEt17f0bNCAPmZt5u/WUSURMTJ
eWooLJZZAHO4kcJegRP8ckvb+Dm/Oq+ok5rknUtZipsLtjFzacnXivmlezE+OdWCFHrbkAauTFGi
i6yOtBXw4vRxPa59oFWG42W2NJAIenqmjg9Tu4l+28VhMovLdDe9wzpMGbUlgv1UJPl3hMjMzVRZ
fD6llY/JtB+TMMo46Xno46qM2bkX6x0lNxZQ2/gQ3c1taad04OiN9ZFQXqe0vyFqK/R3IcITvYTg
UW2EdKBOOPQtxL8Nv0pmfwog9I25GSLlUTXIk1NkrTWB143b/T/ME73PkK/g09I83mzISL6VjaUS
8AXHCPlrKZ/4rfHisf2YaKZnuRlrtlDdEB8EVFEq/jh8uWIXrtDlrTa2tsMfPr0s2cgx8MsHNmB0
AwMwnXyqqdLnFYKVlzsZBqibjN0rv/jVXvn8aO6VDL03BAKnOLHesAnZ51NUBa7C0f1AwuenPdNB
8g8RDn41tH50qO2Bb9ESUbxiNqhjRMEkdmDlfUB5kmQJlB+nGh5yUOAU7+YwDk+bTgXdUrdNMHnI
XFs2d/j28MOqals8ETBjk9UCyvyCOcMQueGlURnW+OUxiD5Dsl+ZoXdyZi7s9EF22teCL0FT6TV9
xfesiPN/KGqjd0qKUqEOAqNlETIh+FmwJLLkwRVu0fccUKvq7MWpgfFV8JukkNIyekU8ahMblKCD
pbbObSpu6kl2/L6X5QzCzJvtqkehTlqiC4LQIAkq/HeiS1l2w+E2ja2bP2D8VTdxrTbvYUkeP7Jg
RVeQbBK6+TUGDi6W7oJXIaEKbRdyH5ub0HHaq6E00jH68hlRTtGfCYUjvLYmeKiql13uuzOLgd7Y
zYhf8gx2JHyXm+GhQV6WJLXnf8E5iOrYmuMxmIOULJTxYaAcXUtR985kZB7Yt6ojaXzXf/ioW/UP
lJ49GrFH2rDYjlUc9dz9WKH3TJcY0tiY2pRz4yII0imKwBN1j+3Fgz44sv3pQr3ZKq0b16xgdgg0
Ym4ljd+Ka/901gcyRENXKj06+IeMlwXVhgrm/Dk9ti4tUexx5S3AcVKGddi/bXINQZqylrqnLBC6
+ddzr8EQIpXmH3Cx5ytwznawaXA2leoOucgy4NdAH4CoM7A/q3rFElnJiSXlvQxlO/j8qw0F4bRb
w3ywVjOSbw1MCut6PUKfSpC1qscPYnfHka8Fp6gFsqF/IyDrviGdqNX3KjlkryFc2rbJjRMRburG
Xaqb/t+Hgccudq0ormzT621vTdSx5j4kBSAI/KWzLMBh8ITvDOWir5Q5p+C7bkngyLB+MezKEJue
lwk0+/Zt3ngyjYrRc6U5+GoDAqgcPdpKkELDjrb/FrevMdqOEtCg5heH5GkajqokK55As1OaFLHf
3pafupgaNdaHxbkO+6jCr8hb8H9PTJDGm4GSNYWQP6Gp/Vu4/zqRH8ZFXFIFpk7A0zRW7Q78hezd
8Rvb8N40vCqc0miVWVSVV/QhBA2qEpb+L4fSBle2DxtH3i09esz/Xodq2Tl8vd1uvOyMGE5XArMi
jPlL5jg8ymmDP9YP+0RgmX2QCkjRlWZoAf5YmHwi5w4hQMPWeP9IsICsMP0w2pLPt6ojNQDWrTTV
9ifyp9Ld/wHI42MsH9rYqoGXQQYi2h0zGuySjHi0t3diiNUQFIOtkphD7QD6LjDqPJPUMCmAF/bN
Su4H5Y7kwZzSS34lD/QCX3of9V/JnnDrekLrhvuMpfgKuqTv4PcE1A77DpNng7f4l1OODKl1JyTE
7SUQYKDwamfxzhvKZtWkSEBe3OPDijIBtEHWIppyY3UEFXrqoZEg/6djK4ygGRycGHuI7BMm/ZmM
ej5WOBa6cPOKP+m3rXjDaA+1Gbiyy7Y/Y0JIFTsEmWMk8NhSLbm7wDD/n3tu8Go8JjFO0itus4aT
j6ZF7feQyvCG7wJHR/OdPPbvInSmqMEgvPdTUSkIqYjvzj/W5WtpMZsNG3blBCSllkje7u2x/PlL
NvtHqnUPXlDL+JqcZjGslxwiW/450g3Z57OG+lzMFR8WIiR84vJo814qITHKcUctWyrZelClyaUb
q7+nu/+3PziJtyoBc0o62QQZEJWJNN0vVCCLpF/e6Dvtf25C3C2eIoA7zIuiBjScWm1c32GenaFF
mTwjnfkNk6uLMA8/ztcRSx4nk/9RvgvcIIMll3S6CFaAMxjSw9yKlqVTMlyRx/7rPMnpt4r6vpEa
5UcOVlBSu7ZOWGe+Yjxyxjg76nrGFXoepA71mOQNdmwS166RwXvcY52aDcW6+/dHC2dE6JYLIgXa
twHuSG2DN2aKSprZcpFWTB+7RZ59DhPXLGQN+pUUbonqEOLUx04ZgiawCwmk0OQVSgvuevKueLsB
mUh0bq/wER4uho0Y33sYE1RaRX34QRdscwwVX/g1so9LpzKOVx4pZKtDGc3qOSxUojBY/ksZDAaY
BOEozSXglOOs3vVpd/WCocjScexIENLurT96OsKSp3s47bNFaykrXsHDpb+3aGQhssWdfAr00HU9
1uQ3H72H1PE8nnRCk+uwGjXc6a2Xqr4cRN6uyaCVaFC7hoScZtOP6r9RUK1xfxQJ4ATfRttgi/3o
ktCgGb9CQ+ZfqbsbUW4tyZKcKwLV26hpkpgm1g48qw1CbbK2fQyf0PNyyzCw63foecshrG3E9bpU
HpqIeZdzlWK10IC8XifpifXDWreyQq7LHmML0jMOISCyO/UUubGkPmbuSAOFfBI6VCq6UsmKnaZd
qnm02kkj2FqbX6W6ERR3bNySjeFZIg0iRtn1su9oiG39a+FdJ3XSjpXFqSrNJBJNdrcugmm10zt1
xd5824kvJXFIrcthcy68769thNVGuavDyrinGlKI0ASjtm9f3N7ij+WJqfqsh92aMbe4bBpPVsP3
hg3sX674+7xag4eNKn3ll7KujWL34tH+AMFqxXedgHjkaW7KzNy2atZ4uaPQNPQs6B4JiKJ730yG
i7G5rQG4Y/b9+7+ddCM1YcFO9JlBUFBSK6mhf/qlppDdigBS1DK6/jIl9U5tNsXuqAIUPKC2bYAL
ORAFF5p7SIBEMKsLcsBqPVmCldDxkh/jbDQoDN9Hk7E+KO+5BprazoCEKeeO4NQcCcE52DosA3SJ
44pOQ9Ejwe0rUcwFh4j5YDcB3sxzI+YJ8EmeadbCrV+Q85gGCMDySHEwSK6Zwb0PbZbokWOT09pN
EAL/PBLevOJ5Nnhrj9eDPF+gjypawBth/+gB4/Mf5GDWQ+4XiiCHWiTWzjsFmta9eNrIHOhLT6SV
Op8qhOLim9pKlDInlAToezfUuRsF/ZMHRZ59p4vrVuDQ8Xi18hOr+eImtbfY0LR+vLa7mke1WCfs
xpZPt0l9OnkLKoZhfyUVryauXG/XJpA+i3k7xQf/ZagB0UTvi/tlG2ho+NRy4WPrYev5h1oRXxxs
OFPgWEMWNtQPnG+yG882Oi1z8BflAcfoKFIm45UBwiDkb3d0QtXBePKRLEckpDh6+zYapACbI5qF
6zc5bzYDJsPKLuabh6faJaCGgcHiezANOZhsnoCoFXvZgLMoRJeb9MkejBfjOK3800HMVnlcdJo5
xeBJN/bJ3IW5bLSElIQ6m3pqvBNHL/BAaiUXrsIJToyaW7Ug/6+jN4cVmxS4LlXgXpGX8pi+32Un
jr4Pq82jNi3zTIE7uybadVaujinXu9bY/LX8QN00Kbs+JikkjRRDsyTANxhvOZyR6GIMYe7RHVLJ
G0d4lNh8+sbJOshDaJ/wQvjiiS/qOm1tIhQ3RMNJ71LCm0DcTlio7PZ+L9kZzhQFxpZSQXWmpaST
gyPj4eTIR3CZBynSVpGoqT42sFq2VZRpBLXL40NXEwEgROxIyVPUyw+geJA/MqxVECRs2NsCNdnG
8qYuHm6K9vW7qxloqn4HFsidezForYlDGtUIaA/jhbcAzU269KXNxFU9/3Xri/G3JDrQ8OovnMKM
oOLJQoUfyG3YSQEGbhKDMrCYkJfZbOiP3ofT4upu6jBnDRT9NARYw7DEoNAgMeKPVle4/0zDl9TC
zXZdU7uYYx1IQ8NkBCVv4+UzlN4KJVIUwaRQKYKnojLZLnN+DtDvD7zHRy0fuF6a+uE/WofqLzpF
13dLGbavchTdQAQFZ4dDnNKz5apfnb16g+Cakk+rEk4/2oMTHTwlQCTsqY0kHGGTkQ53pJTXSG6w
mHA+ZHDr4VF1xHiIxXL8IBPTQeptxDclyyEr267MQljoI67Y5Lo3UvLgQguup8eaNfTjkvENlzN8
1q3LjQHFQClYzFdwRnI3BOWr5W1Ggb/gd86OXrW/IQxYqLGzaHScmcBt3NdjnGovDAgLZkhSsxX+
aFiHfkSuA+mEkK0SZur5hxX9R9R8ZIZgC7KhkwDtezqYIN7bVrnB6PbyhH9FFs3sU4NL4Ll8K8VM
LgtpxsEnYm9grM3zoZSuV7OzL6K/7+hsg4ZILes8bengpOEqFRLRtqsHZ4dbaLzIe9euBQO98p5W
wXn85eiG5SA/8TZ64BtzJMwN6rYzGFy+gay5kFPbQ9VGaKPPejgQY8lazTFOBQm2C5EmMnHgTOEO
1igs5V67dkvLryDdXL4Y6SXEZkHR5Nh+5mGIvTkFiOAEkgjk+DJNfSVaxEUA3mWobl2kBA5mNzr5
abMgLS+9WEIg2wzmTQ0ssW6xs/LRuHsrgSN1Eo0jXh5zWQB/cxBa9WGXB2s+W0I6doCS8ffmNWo9
1yLMpHymk5DhHC/ME66sKQdaAVGqB/RV+wnxeDxPW4sCp0TqIzfB5mrTrtNxX0v41Q0tMwcpbGfg
fHtsgIOUKaqmLU7+mmKx3v5ZXnNBXaEk3hD3hZmotcQlYnVSXUOGP2hA5ZjQPfkeFLJtaDp7+DGW
qohm3zc7pnoG9hbxoWDXHLm8ThyZHiRVFWoePM1oh/lLUV6pCYYgAogNGkhAOEJZQJ4tZfCyPEpC
bE8y06+/jCGrjWp26X+mcQOe6BuBbtSFuonoIojSNlAIWw/pmgwoS1YoO/tFIAM/SjFmBp594pTT
ZsJ47PZGFl5Q92tRePZ/CqgXsLupRrKwDrxByg1KcM0hSXgcpRZpKXpk+WZIh8HNfxWGJziz1xtI
hkGCawFjwlMQsxWHwKIhRGB6ZnGQABIoLnjBoKBnQRVbHkYwpQGt0CKFvVNt90MYUVssSFU93hMq
FgzrbM2AnZSWkhdZWNd1KHcYTN4CQcSr8rPVYTpY0Az11/4vSMXhqoJdhbqoQYJ/YazvelMByeTD
NhJ5fG+8iVYHiKvrF0005lKLhPFAfDAl0+NeReb+gx2vifgpXMEaXHs2tSAlfWB5I3/wkmxVWpu6
y4kthgBsK9TsGS9GjQowr7Igiqeh7XoOe4rap3TQeVP2Km0lqtz6Y7t0sa6PuXLotFegTHIVYqlj
pD7DIy2FKYy9EvxtrCC8kHsrgI+K0No3B7P6PFBi7xb08YS7uhng+foVdwRFjc1+vf632AfNUfyJ
qmzs7DYfPUn0SB9K+8Gap7oQd9FIBueYeCO3jpAxw1tcIG4dKuxhEBxsPOxcpmvtFbNtIOo94jIo
fCOep7qcB8trPN30BvKtBFoxW/trOUlsCsMRv7k94806ms0tfqlyJvmcy6xNHNvkq+/3eRW8NGEc
1qy4KAUPv+3vSNXotBPOiQ4hH+MF+RVRDDeAYvcjn3BZ9oh1X9Tu4yjKLrSvTjIEWhqLPw9nqIEn
+5mY+NbXghEh13jX66QYnL1h0qNRzD6lbJB6bbesReB8tSRI89U2RxxxKBvTm34uEIkMAWkTujew
F8Z3JX5f8WAUzZCtCeFLRHsyUC4iLHNFOiiiTOQypcY7/b6SI8Zv7vV+WADi82Lmss5TvuAHDp8d
vRS8De1gEDRnVq30je+gvepts21hXs+oaKnEkDGt04Rx0ammStVknbjZGOjAC8+zuj3zG+gaFVL1
ljGj3IkQdGYYpOhOZD+UA710v5JDFTFeh7SvzOJ0I30dBE0cM4KrJYY5bZplH345WZtE8DXsweav
ElY0WARetHRB8UvXz2NJQF1lovCQcuPhFm6a15x12Ofvnqvtlism/r1UpZXcfE5Sb43PBASRwrcX
5ubFDZb91M4mdQ1A2STtEgGXFc8+Au8dlWEjLY9YPokFcmG+AXRvXWh+iWy8JoS/VGhM9bmIceXe
07BnyslIYUN9FmyzCUoNOVjdDU1dUA/HV1Rfg7grhH3KUAvtdpL2CyJNy1Xe6oh7UG8OBztY0sJv
Xt56IS7VBoGP5zVCxk6gfUDs9U9aiLDRbHQ+2bN3clDfAa6HWxh/bR/ZK+5RQWnjNwWZFcor0zNf
ST4z1JNNK9HArS2FM8P5cntx21rG3XRQhk70x5Uzp4S433jee+YI0ktSXJoPOQnoCCBajWc6pxl1
yyxbsD9lZIUGHEuANK71l1JS62nNPeLrvFItncppYIiUYHUHhULU5mUSwEvYCR1FStgkujCt+G05
8OJCR3RJE8JrIAEZ/Z+/VT+FUKaoYbHCOYPsP+XiPhtjnPo8m6XxqHmKhLt+8h3lTvLkb5ljRglv
s2zpCa8hAC2q/ULc9WqgAi86g/hc5kB9iiq8UhTsNAwOo0XsgDdDny04o0OedHit516jzzZFW/YC
pA3Spw3DIvs90bx9LxQErWdFF0LGMTQ7ZQDhEtXj9f5Ex0MCR85wVkSJILTcT6jy++IPZsI+Rwmg
mGcRU/LmYTnb3Q+xDuHcP8YqV3TwwwIcEwUSZF8kKIaUJxb0+HSubibIsr4hvC+qeKmPrRej2ME+
pFWJfG0PWvzGE0b52JufxvSXxjRrwYOsi/H8beYTSqJx8Gliag9M5ZLY3KgdYT1ovDugFXv4o3cV
hxkT2UXZWeLLLp0FewSHtyrkH+MCQ2eV433QdyxEUwknOukmc5Udw2tbp4ueGxkzID1WyVyiNcFG
bgoaBhfS71qYQOxv7wpifbFlHIkuCN5OlqTE1OT2TgT/iUZ3Lsal7mXpy784xPheI/FfDl9DT+bA
St/ITBpqt1lPI/qnJpHfPkI9zzpCEhGmx7QOP8B3a02Jn5YJq1oAVymUH+oHONqdVlH16nAhfLMj
ibk+TBmeT46KvdMVQw3cCVoFbx18IivFgzkmm6w2Ed/xPkyY/98KFSkLhbZzXiAKbhg8hBWkL/LS
Y57Xcxo1bkDUliuQE8sZ/in3IqT3uUY9hDN+RQuo4dnwt3BRL9AJEJvguKzU2cDvvnX7Qgl2BrFL
wVkx1xntoTkdmSB9EN4Qy8zWmvo/b05jgNehX4zje73TtMKjVsL8Xdg3bfKi1znh8UVBKNuKgWlB
d0hQyPRehti0snM/jVr+0k/DNrLdKl4JaGgMiFzxiur84l2zeqsuD5B6JqhHStCVGnZ+FvpfEwU7
mR9LqIlWKbEoTLlhOWlQov5rNqbyq6MRDHAvl5/yYOR2wea4jaCq1HI+X1KiuR3Q3Pv885VLF+Dp
y0h4NmAsJtACmclsEeP4wn2UB/wA3RlG7BSjHW4LtDPGdm50yw+5iXxhphGUyRFtbq318QEN1nOk
Rso5/27pr1lK5031JhWTEQs+AZfU+//MfgqTqVMZ48Lisgy43mfEoCHR2+OwgTrC8AQT2IyAbRg1
W5n8XRcADy0twHl17Mf3QOt61MsS92tuSHTbyL6GMXS+Ppjb/dfGj/PPinDr4X8l5b0FOs9ORMEQ
h4gtpuPFLIAozz9y2LayqrZDN9xahOqntPTUsXj8MXj+ivkerHGEO3H1O9zJMj15wbU+rYTBS5MM
mtRkgsnWCvsdKlhKrb2R8/4rkf5z4jDGFitOG1cyr6lOHimsAAQ593kzCxS6gxLtD6Im3JW+YYd2
PCV/ryj6RKLwdY5p/Gyg+ZZwo84Nv+VF3CJiPnzCQkXkZwv8VoP0nWRKBZl97dpX4/AjbttPBKep
GCy2hBQYbQsOLPvgOW5OGdDAr6cXEH5gBNWQhifqPiv3Cl9aFcZ+mOF+89oFWMrnGxOL9A+/yJtS
Z2KNhESIG1RdVy/Z59BbchrEzr0H3MCMuag52c38qzyZObzcWeYURSmlz3Yboj7c/PyDj+JNj43W
FZ+SF+yayDtvc8IbJ80x2mkOhHs0AQIbEZqVldvnaPOXouDrQyqPR29R5C/wnWmL8bXHrqqSUAjf
ijHfzmzbCuWG2rTWGukqYgB7J4xmnMNWw6vOF582AgygId6gXlvKnX9zPTROqREJd4P+XStB79UZ
+g0Xk7+C0O/1yCFWRfWUQXrxGiiyHIqb8zsCba8meIAj//vcFuQkkiavzZwb7pHKjpr3dPBVoBUb
ti6nfVZ3mIUnVP04IFZYU3Ho5655UEKNI9CoKwGaEN+ZDTjCKNAjUfh5OrCE166Luzqou+foAk3l
VGaSVg+Q9oruJe2BzzKPLY6oylcEiuE3DKIgkuldbTqP5Z1Pj9cVlidMqvNuBVV03GhbxqAzbwrF
E6mWvEh8uVPJFI4ndCvohX/IHulhu+5vk+Vu02PoUjHxQAvSlyqowyMxZAxt9dmVGmQBMWsO15tK
QqUd90m1ayWRkIJbeCp42x76foMkU1My8pV910EJNdxc7tAJOKlcE51WAIzhbCN7obiUNAMdicGv
yIKPjrsdMIkwiEfKIbFe9UJb+XB971UZhvNptXcAmzWGONdKCH4MPDnpQ+QRVbqbfC3F9RZJgltP
XFniKIqDXkc+l57cCLMJ9cEJxdmJL3xPZ6smacGL6ZZJcrE7ewNwTNvrD7EPlK64fDt+9acr/0Ll
LmCpE9bH20SpwrzkP0+eZF+sCanqvMjx8p3QHy2XvtAOIno9bZeba9uz+I7cBJIsyuUeBNW3SeHg
gPjMEblHsXK7WkKMpecE05syBYjgPI4zNcid1KtFtrWqMJfHNxDIQUNwqOqydI0ds2xp/1HkrEtv
QGWKxS3ZOmoX6ltJbT8Z30ZB6jIrX65YDepzGFzFWIUX0zhh/CpldNosxjGYAtqsiHNb+iFIdVV0
qbrnIhZCGvKPrCzA2IN4NWraTNmDShy5kgjNmqohs9RV2AZSDrARUexEvadh61wHir7LFZJl7llo
XJIPCMLTZq6LU4AubcDgpaBUODpI2RKPBOigfLhQNiK/SKkBENsvI29HT8zVf7L8XhT9bVaeoHzh
H2+fW85zI8eE5qCL+HWAIvucs/tcYSEhs3eY58z2upFJzB1qyHPpVFGwa6dTjm9evTRS81P0lsO1
NPyVzTkSyvDCkkjoaRLaXLSQhkEfIh6CJt000+zbhIc0crEZlwpuayXaqvbbkJkfhmk00Vghx7Ca
6rX78EJ47xifhVPPL7rmtUcOekWOk81jAoOxFA7/8L5qgofb/TCGpDM6NbnssMAETV0sM40eqytk
avVlVG4x6FEgNHjRMOJTkDLg9/nrelrcLkV/OHdfbY5AoOXgGAZ0lmPC3Biye+iYtr2GF/n5tCPY
SJ+DUFUAxmJjSOQ0P8p9yzeutlGNRnXAfU7vgAewv+wOFJVF5lyiStN0aEDRBKoDdVFTNgpf1uyD
npJF9ss0lYxzm9C6BAspMtUWJXPM4RDJH29lANPIfSRvLrC/x+MfrGebAWrNmJRQfaIgGYjQYC+J
tZX160D+sTLMMhxiNtZ7EiymczQ5BBEb0kBMchNfXCMXoP21rYuE/GIe0CC1x9WnJQy6/Vw5gvAu
NxId+9rx6G2zIFGpGoaqqF1zkgfdjsow+6+eCaH/sQU6aAIGMdh7veaQryd1cTEW9eLfpujtQj+q
Wwha+AkJL5teadLvqWtHrcEULOaDnuKa+husAiAERWoW5+vnVRCkRN8WnO7fS2Y/xab0iaFI7mIL
2SPTymlJIwygLFBi3V2EApWeuZvuTqZSLsjGy5bNgyZEEaEHWjs59lxH7ZaPOBDl5E0OTrdPLJpk
qredVv4yeB47GcXAui/UJVacjzzRverPIbJ4MPZuJS8OS/h70nJ9hj4y2LBKxjKeopiwWwdYil+o
wnllu1/7MvUO6RfFcHYbnxpZ/pAoBl2Px4mU4yGRmVCghlq7uof38LddfUfxozzzwpZlOiJs3lns
PDixmL0ZT5ZZHPuVOyEoIv1kvfzn246Q62v9iWzeXLAk2Y5qcCnNJdMtZ5vO2gu2tkNhCX5pFIeX
7rkvVObANVAZNyKiXm+QlqEVi0C8T81CAAVQyMH4Wq0wbvyB7jUmQbU0W/nCW03U2I3/eN0cqTVA
flkgvhDneTuTJWxBLZfDGj5dT6ruGUojcTBVQoi5W8kcSFzJ8lTBH0+L2sL2Bjzcse0Ouk0ejnZi
dssjozawe35vj/iYbHoWdow1Y2e+1fZmq/CdVRm+kAo7/o7CEgSn0dDcDxcoo4PboLazYbWaTyj+
R5/dpBIbq9UtE77pLN+9Xqr5cgSMDmzTO6uPRHv3sPGUMA5XHfVTe2ImtXlJA3xy9/46fGrK3OvS
N3DnMUXrnTG7632oAJdsMXxq/twPZxUT/W/D8vPxceVICCYyuLugexNoBmhfkKy44Pb5/DIiZn3t
o5247+lcxLq32A5Jx8mGuW6VJY26/3RwkuX8xwRtannmD/CPR0HViWwKA5R0jsG6eXBdOfB/GN8P
ZHLxiZivGgvso+Mg74VeLfj07MYZrQcqF4+OfB6lXm9nT2EuDfh51eKW4UAEwICrCSPtkUi3423J
LSSsbVjVgSqxH0OPuVSgT46oY8AElp4XLdkJPprKJ/x1So8QHz/9bFJZiGXPi22cc+xRmhSLWkq7
JZTyPJsmEb15ryDPnHf7jZNT03SJme/76k8/R5N5fnGumavZo729a5q6USlqOqrYfbQlD2WxxM25
hCWo0Je2ajS2IH98d9OP4TQ5IzWl5kjprG9rOXz+DRilQJjm32ew7wQQ6TQQyI3hO+GAic70NySs
saJkRRldvSMCNej1l8fqTy3tHuUhgro1LQQOKS1OJw0gwy71nvmOro0KjNrGuxNw8TrkaSZTOiBV
UuIzyS9luoEjdirJ/voHAcBjrJ77jC4z3dy5J0hmb8j+aan9/LKJfN0ickkbT14L2F6t9LQNSyLz
+z6Wxq5ZE16oh7RJifNoAh7mZrC8HAcXyNL4EMvQiyGQZmPdFiw43MIWvRaHk4+LPrPcR3UldawA
X3vL8sKkNVbH5McJDb8TdGixtb+a1uMAJ9xG0Q8A0jlEfsIFAJRpAgItKFOy//JM8DzadgLhEwrR
cYqcwzJ5ROvdBrkvPe72wViPgEglXUshcjHplTqmHm3zbtAeVXp49AAehoy7WI0Bwo68Lq++5xzo
C4CsFc7xinvdF3Op/AE9o6591D9sM8bEv0NniTLLX+lfMQ8PwlvGCZ0bEBFtBgsyM9sMeY2H5wMX
NFWy7uHGCDUqzo1R7FD6WZqz9T9Pb+ojcXoijTIcLc5ZNYmgIPEauuncu73TUq6vFxLCJWwhpl6r
9hpVrNvwc/cOSb/Lvn8x/T4K3sQ6nGdujkbvyIlov1EdWgAIrlYWj2dhblw1gz2Utb7T7gpwP2n4
hPLBrMwrc8w+StZ7tE2ygu9KNlMg0yyr4I/OLFJbenRQWi1b7JPwn3LzvoO6uTNmtdUy9mXwKMD+
Ny35ImHw7LlAubVhDfFenn2uAt8krDqPOV42KnzL/n51+UXHClAk1IgrIjeGMRov4WvQiWIdD36C
FXwBv+Ri3v+1coLxm+tPloYP3mMsGVgjEUwne2+HYAppltpH1dvyjzwkEoXAaiZrOFPCy1aEwor3
3O+u6PWWifGlBkBYD7IbA8oprpg7PqNxCPiUbBDMEZffARFe2rZNPXJwkA/WLbtGe5spgol4IrKc
f77dPmp+FFz7gC1MKiH6YbQXQmIznwNX7P4tOgxVHoeM/FZJKTi/mjxSfW8+pfOHRNk0FniWRKZt
w/7ozUf7Wkar6dOAV46Jd1XePwDhQYa4ZOeepnM9BdNwI/RT7tmV9ydrYA2IhTFAkK5RkX1oblQZ
riPDQ/zdOt6FJdv3nbvQ5Rp7LCIQ5RDpPHBm899wYgHjAvTue7y00f+3VTJvTXgxq+B3T/0b3P84
FV5s84aCUkPssYDy/CJppHASyiC7enlJqvIqIEJGHK6ftuzCBWom74bS3yTUSrNcs5YLZ37OUkh1
zStbou92Bh8u6gEztUwhk8ibQPWAeufCp0dGtJTvoEbfVHdOwujQMizqx57YO8owFXZrP1/GLq2N
RdhKw4myU4/sgDygW32W9gkTL8UVGwfQNchJHfiOVAMRD7M4tBiygQzV/dVoe4Xs/r10OFWZL0my
FU2U9xvAqu+iA10QJ3VrA9BWPFO1R0fhBkt0K/1n4llrxfOHVnLKrZ9FpuTshy4ld4JvIZBQ9bAf
YFgZpqU3li505wbe2RpO4jtZmv6d2JUBYSVz8torWsN/CwdZOdmNgfbcI0bQQeFQwAhtDNnTMwfm
lerwzpfnw1dnaE1V6vTHhkGDemqlxMFepq9UnoJhN+EpRNmcwrWqePqqDFR6+u2o3pOlto5ESYr8
Jre+RWD2st7bV+5KZHVBiaT52rRKdc1HR6H2MH94nFXIjHABZBn2aYLtiWLfdQuf1YIceKskkY9S
ULH9pSbqNfy2hro7NGEVJz2oP/Uns78xdjNoSi/I9ApEXbvKlIUnJ+Kfz2I76QHKCKrW2GfQQ7av
/Ybb0ORu3alLyVQ6g+A480PVFD9j6CrDvhIUcc2u/EdTIc98Llp1mBso+yMlqQeD0/oKSy0A3dIS
5sXVarnFfXApTXOnuKr8TNyDfiya1EkN6e2vjFF/PjV2Yn4qMOrBmjY//SgQZ8DTuzP/GZPlhBGA
XNYblJ2T5sRXQJiOky38XTtkCZabncT2g7EopBmnh0+IJadzRmdPjoO2TKBJAKSK9gs1lq+LRLLf
+f3/HAmlHgNPuk0G8z3sVuvGm/rQB0HnEZk0jfLoZNNyrMJ/wx91vwJHkmUkfaXO38xwKSHMhkhb
Ip6+CcbNsn9WsaqmFGT6NToHO2LgYhJ4yjR/iHq3WN2RDE6+wmV/44wLPxFcA38RTOTRO6mF9/IZ
4nRKCqeTsoRSX1m+Of2IK0EUnw3ydytjy6FJF+eHU7aBcldAAejna2NBWdVLV3OyO2Pi1UgK/Z11
jbRrA6xpKPh5rUYiZj6pXKEQMilzPF+pdjzSqElfco9xv+dihgIJUlOPE5eXtGmtMC8a697xxQvi
qxHXZkKLRY5hq+s4VC0aBdnCyVJfBMuIMQRkMgRW2cO1wOLidW1SBBzYuvEXYY/T3d0Wv5etPIpD
CsVTJhDkN5Ymq12AYwfd7tLKhDsuTBsNTxqM9tGLXj2eXMm0Fo5zSG9od9+Wjpw714luO5YNjL5S
U6cWHaw9ZCGTg4XSSphm6nfi8cWzUO6RkLItYjotzJQPggdb1E4LQmcs+0l6e0AYHquibOSlVLkm
Dx20VH+qI0AbH/JBbuoARIargW7yx8lg1sZqtgz1+P3vqy26Qm96axM/JTYDV8vcyWb+VsVkfBfP
+TOdcDSCixVoClUxIyA0yDV4axCtCk5e8lPFktF/Q14V3npnUhJCG4ba3qrR0nmZ4ICdKm9fMAgb
wqrlb1fry2GFw37sNjQU17awV4qfWRX2p3ATI3tmanbiitWaLgMG8VqYwjMb6ctjIGy0pMDtN/uN
GrH9MQrO1Nlxfwrl8Zh5/sfxWUdXDFOT9It2kScj07058YLAgHnQ3/RndVCb8203HX/g8wMewuDX
zm6MuYlhFK8l9+OJPxlijLTrFrR60YGfbXZZ9ZlQTvNo5/2AoVOI9LFIvwUoJxoCjBX9+JLRAi7W
19vvSLqJNdOe/BK6ljJIFoHDKb1ORK+848Xknv72uqqfyL176SQDJjgdp9N4KWMXGCIqNXxjmdAM
AzyeMGzpvNtVCA6JOgt6mRaVh5C63kOKUUo3r0S7Cq1vrflW9sLtGjNWcxmHAqI0Pbk96kKC9N1W
WYfS6nZHyptpzlpQoX9iJYpNSyDSXMCcz2UbbcTuY7SI49aftnS1TPX1fcJSXCKg9UOanxCa22mb
3p2L0gj16SoytUGj3c0arrkIyCAigmTnYz/VRhmGqmDuGcclej8HRue/KOwWGssRNjPOfF2TDtdn
XkDhwleg68U6KRCxawFoFzeD7EiO3UL8q/Wg1HiJ99Sokm54x/E6RAjp2/HMyVUnPVNlD40GsmUp
au9TQfHztAH7hAhRTP/XbwYMrM88uw4cOr/43iJq/cQrPEAJhHDa8eJ6yRh1258QBcCOs9lYdu0f
aZnScVI1pu6o1UAbUpCavbf3bJS2NAwkbs7BFcJw0zVi81GVYDluDc4EQ9sQgmn+zWahqyg3IFWv
r0flKLQQnoJ6TDuMnZouqgGQKMMXl83kFjUP97bjdwrBjndj9EPDt4kKyqsdhiMNqKy8m4DhDsYb
MNH3PAzhUUmDRrc00XCFWd6s5OUjR3NYuqUP73goF3u0ykLKOmJAPfWPNuEUS5zOaBPWPR6HlLK3
R6JnIsVYVc903bx7lr40APzSwEoFKN4mRj7LWSXKRdOIdMCe/EE8s9H2r2SxPDkxuoE66AZvPHp5
zeWBDHPF6uoG0O7lk3nrdKySD7xQWq2G5wYBXKxv4AlXdQUPD3gcB7u6a9GFo2kNm+kkLAeed5cb
2y6Pz7hWSe4zW5o8kEqZOz3seffrdaikzt9DmoYbmcubjRre8HnJkGDKdmiVnOn77bws5WdzLAhQ
LQIIXUxI5UsYuPy6EldtJGpCXhwVM1410AEQ/VrEI4/QOxqifQkBOlLm3dlbmRRL8nvn5vNvSUjI
Ov7MJp46ehdSiHLP/r7qcGe+DyO7cjxXFGwboSh7Jd1in4Z6PtXjt+vtmqidJOK4aIAZvMRz/ZBb
DjBTbFunuG8EnnSzSAHk7giD+Y+JIlph8kIowtRjIZLHqdsTXWzUedISGZlk4EhUsOYnR0x1MjVc
RE0ZiNBeorDgOij74oXAylWa4bMKl68iDDN62O6z2QKgSmDksRwAqZSCEJAAd9rsTUKk2zOMzOTR
Ct289jYC2jb6dSUeBOZ8bul4gg9pqOp2zN5S5tVHzW5szavibAwP0VkxOLstLdIivkvEEOq+pZFC
J0OttgvybcLvUULnFaVEpMPv7EYR/7FnkfK+3GwJeINcrWs9pIVoj7gz+DDiwcw/poLHqVq9+HNt
5L4O7nciWQ1OLScrotWhaPbXLFHgCYWRnFZc+Mq0ioXxZF4fWVANVOq9Y0prxewWlDs9RVrDErv7
k8C5aXtX6grsv2lmciJ1clnJNdigOZmJq/9QZlXlRK6chYtyYYozLjyJwLHJDN2qyUSRGIX9HYQg
qNaB65kfS4mDe6UC44qwICr7cNSjGcWOBm7gfdYcLC4x3t3E3jn8ibmxpsrfWM55sz3lBQ9INTQp
fpzDTobaDmLbwBHXDY+E6uDHqeChgtRPOIap2Sk3S/kKV89CK3Vri/APEOkkiDGCaY+HT8hJySDP
b0/BoA1jcQdYOMEepQfjJJj6iBmWgz1oN5Bd+pJ+UjOTW6D9noUnKHl/jI6asB0WLSE1xiJ1CHd2
iQQ2t0Ed/F8DtxdILn3IZ27ZAPCVSDOCYnzMIOa/adjIzI/7AMMWAUGHev+JIfFLdnPXbz9JmNWV
Y6idczOVSt4R+wmOWQGaX3dpmjbsqAUtXSe+asTt0U/tFPSoLAWyIgA2qUitQzH+BKSQnL9PcyEm
isv08UrvAkPp7w7bL6I0r0ww3D5pDDwDHx3smFHb/mxObut7qz94tIJKq+LbecBAgu+pMYC+3vm6
I8Srw0I47EzpeTfnw8ue1Aql7f8E99d119ejGnRLeQQ63UfIsE2C6nBlA0ENeL7b9TKKgP6Mqg4B
rGP62VViVEwEwkKb5ZxVEcBMkQZo++/p1NgdlApYuEenyaIdaqV653Y9q6fMtyC1AxxaJj77jVWx
Vb/6JJ+vKqdjijNbXC9eqcmmw6UIMtEiV7LIbNAekrSsMlATmoCTcL85CG/74Wo+k/0JNaMxzezK
fOgjRiBBYl7CuwZhV304q19K/et5BExcH6ZPpg/6uCSnUiLFNLglag6yCrp6srYbz396MUYqKhXG
jQMk5HzF5p5KzmIT4TubgBflw4TcHJM3Qlc4N9EvoVag2oHO4IC/7bE/T1icco6O+KuNlkPON5Xr
PxeZjiCJM0cQWLLflTH1CukOIooA9kbwN65D7MgvTurkUVebp4wgVoADhNDouXCLpp1/ng9W57Tt
tQevY2vzZyg7Opfd65CxmyJe5RJjPus21vaJDhQhi/0bqCoAzzfWUQyC3I0F7X1/RqWR7kmHzHis
sCT+l6HMFYwDAcGQ4ly83fuU0xyPTsbpYbmfUQitVOVrAvrEVrlYs+n1XY8oMW+IMSmG/yL/AXLa
1rJBRW4YlNw9e0knuofS8ae8v+DLopVsILJLTgndjkCxf4bdzDre2vo7pNiQJBuUVADalaqk6Er2
iVeNghSSJgAKoD5Ryk0oXvxLSwH6POijuZ3ZEnOWPFOUkbJFdT3cR4+as0bnxiNMMXSVQ6HgbpIj
ed94VEMMAUGW3tTiCXEAXBTR7xeTIiNIHLItEQi/5hdabtxljmlANZKl0yOJcZobzA/ClG2qySlx
unacQQDIsveZfohzctrr1UMcOQELiIuwZsBrvP1Yv4nRv7Z6uxSmwXtjRUpjD6sRgy6k4MmfPg9A
ChMZa24m4FR72AYw/iZONJC0qyS3kYeibRMBq8elTLii4nI67sRBxGOe8gSt5y9W69qOMVY1peX0
Bbhne6/vlrAQ8JSYfRHPNYOeXV2P427KR6TAdHQ5+OUKVwjVVa+Pc3fw/QGSHY6rkUQeRknXv5gN
UGJCY8GMHrDb5RFddvlso90AhDS/wwtq/jDDPlOCv5mWM5MOXcj4KXJzbrjxlAM70DOghMTq49fa
DraXt182/juMMPmBM7IOhMqMcLC5vvrK6pnRysl40SBdVN5Gz/391VPmzEjKOnx+ln01B+cK3+MU
VloQiarY4ynkmREWhdpoJxrCGKc5Qde37EisBqJ8B0fS0VelM0EKryHuHgsyEUSedLty4OF6sMzO
nUyU7E0y5mw0KfBzdpYzasiTo5lKZQq06X2dM61ivQxeSKn7bc7AdaiSgrTa8H0TmtNKwZotph//
DEVikjfH4X55HJMTpEP9VfWCum2YzqZOZ7wvmMWhxaTt/vqB1kD9e56LY1rUqpo5moFMDnhPZ+7Z
0le1klJUXdv+WkoLdxeViCHFzBAV9fxsbhysRa1zumNLw+dz8JH5/M5WraG1LHAqRCMqTd5olu0g
zGmySmoE7pTTdEuWWnYjVuJvegHb72tVvhSi2Ya6xNi3dynh9JuLTIKy+eRVXhqgPHVGZHGpwZC6
LXzrc4g9wVa7bJttq3aUZyyAt1zuoXv9GrRucqNE/h779pl6nlt8DWhSEdk865IXTGe8w+4UaFYE
X4B4/8W9FPzZSFf0jmh32Bvr4lRkVaWvy1L6DuZI6NiR7ssck6pcDZgZwuHO2eRUWsSmV47AoAvb
Gv8Fbi7LiROHc9PHGYB4O6rfba/oN46NWbMEqsQCMV9BhLatj6P9lCIX/liOFNkh45CNfzOJ9MQ/
eT1aS9meUh1J0/gJGbcvIVLRlfMHXbSnNO9DJ/WYIXo5sccoDK9QGpbxhG5/Px6L0BAa2/rzUR9z
Zy7d+h4tPez9YDnRbvLyYIOKdxcZA00QvlsrkcJZw75dF4KmE6STjlxuuLJf+LmhjmVieDLmkQP1
btu2YE5Yi46rJ1vEJONQAV6pirg9ykzYGVW76zULRVLtuUl2L9YS32E9F7lFgEkjRPPpppOzZ+T+
JI0Wqn0ii9lpOGmAuTWoB7a6GgA//GsTRAI5k7EAQoObRRgriO882StxbDeF+UxnU8sPiHvJ/cqo
xLpC3cXhBQUQDHVxfYz5KbHkEwHXtDBZNCHl00ckRfzysmPTXXQhpsyIFxWTv2Z7B0nEp2CpcvPw
CUFUWKNBeYmEy5VV/qQ+Di3yLd2VXDHNGpV+U7JexyM6pR5m5ZgyU8pYHK03b5AIIv3E+QMRs45/
7MNklkWgk3ZP63PP21S/dvsqAlBMUaH32awR15TqX2TUBv7vXXmpdjjw5ZcC+2p2qpWLbe1aeOjR
O//zS0cSafxc22tD/gXV6mtSvTlIedEsJ+qaJD2qL203Nn/hd8UPWPyhB8mFzv6r6xk1JZR+r+6G
TPquKBmQx+oDwsnJZmPb+zh/trfBmU7qjcIuguEGAeoV7uYCsabri5EhpRUEQpSzXtB953eA3rah
ayrRpK78Up6lCrNozCwcOOaVaKglkJ53lvjWM35zN+GfA5ZBzDZ3VUG6fnyY7yrBmiFlSXcOjRX8
wDPT9lAHBBS1GHblSRkKOq8+tJ6wNg9nPUmUCfP7hncEYGusDsLqWR8hDn+adc3yacVgOzSiw6fX
Y39KmMV5PHhmd9QYS/QbUeoEpyEBrCjCmVz4NOOvArOQx5xn4SFzVxA1wNNRJ/YiwR7YES13a+15
DvCBl/B/QJbI6pgjmJJI2is75I3xHdBr8oCShrgUCo4q7P/DbUtfPKrds7YNGH5KDJAmoKZD8JIP
66SJGjUHZzn+ge1KP6xDmFKToWKYOcWUOVuzzf96joNsHmrJSNbWz0xO3cQL3FdeeR85tZ1HWiDU
9QonwerUU3ENLihMB1NGFrU47r8AFe6Kb1N/rzBKhtGRoxLbsLQ/Y6MA3AauW3jEOEO8XSpcgwwX
DmoPmByiqLN8J6P0jNibI2G9E6YKRrGzyj9bJBFBV2yBR1qr7t6O2UC5pI+GVzgCp/sitEEqyFMs
APTh56rzUSJUlbt39yRJtfnBleUDE0lXHv/mzByn3cfhAlBKYJhTuGQhu0FQtKUbCZmCbjtRGUmQ
6Qck0J7AJKBXkH8Uvvs2isjOZp+WjhdkuAKlXmnq1gPxgSNqrIk+DRXpJbs84rf89u0OJmPg1A+w
OLFMGEs4K7pZ7v2CUBQ0tUVke+gZWGO6/4B0qYavbx5J/g/57wre8Ae4SyzDBLvF++j0M7rMsu4F
lD8LVcekF+0hFe3STTwvx3U4tKvencNAKKiTUKOR/wnVcaCcdgaxhAH16uyDuS8clp63f13qaB/z
/Va5V/W0cwXCSc+rNX9rddc8iGfscaO6GEZhFyWe/laJwoTucNWW0y4Q708SqylpgKLQL3FMDwMQ
BlmEwU0cuRv39GGY5hgGCRj/9AcG7OPIpyzZHPGQk4IwPFbt07Q+W890oW1PgfosA92/hkwMDoZn
75J7B8jE+H9p5iA7jfJRtfnBq9JnOwsPGu0P6Ty7OoeB2OkDEnH8P8GTj3V0AkfamTqIYqlfVWYs
8oRiLTuU1odNTx8R0ePTRpaqdznSj/k88R6XPCgP/yFNuHadhTGm1ehz+v87KvE8RLVciIbOAsVI
rJpYNt5doxv33Y3kaWoZi1kl4fmC/wkFeQPQdYSBrLQOmg362VoYFVS9efIuohoKyAzG1Bsp9nIX
66k8qcabVEOs87S1RuV9n0O4q8ea79+IyRbUS7Pyfpfx3OzAnCUho2kR+arBTgV+yftWrFPUBFlZ
q5c33P36bXmH/JP9vsUsnPPtiiW5wyuYgq3ZeO6JkVsMxIuJxqz4q1mGsLfE4HCDScyZQgfi1vZ1
f0qb77IVgig+i3hnlSML0Z5RaSELcXlg1HMSFrM9OYmRz2gDrLEKNPGzhGmfxpaKja6aULuNkePY
meChiC7yby9bnQvgyxKyIr8PXrrDyoueZpYGpqN1H4+B11XMk2t4WkK6Cbmf2RdJT7XcHXqGSt+R
rRpEpN6Zx+1uJNCKmO72HmYZBl7I4nAwHZqrTJ8gRoXOWIwG4MiaOZGYB19LpF/wk7UV+ja0ptg5
Atwwwp0d8+NIZEg6hedMaH77CdhuvQJQI/ECTOp/EQtrcpkTPLcDEJ4LldJdH+ycoIVendtC36XK
J5meazq4hOKNA/dR/V6f5K/J/5Tp0uQtQjq+E79k+nNgEDRy7EHmMT4ney7Xj05e2OQXr24lV/5A
NjZqIPAzqabC6kx6wpvPIG5PlnGjjaaJRj5qZr1FdbrxE8wSEXJbFpioU7fTkOU/Mxq7CGZ5G7li
xupCpgW844r90y0+xckkiVLo9ntdwxUUgMZdjaTJVPSS1kFVw4yTCIlDdwV667XPzCUehzE1DOoE
zO9951LBD6rfdNFJxWU+XRorBL5CBGXGz5i59Eo/6TK6i2leMv/wBQjxlTiAGAm671wuZJpthu/B
a0XmEGXNn21X81vSd7OPEA9gF6X0CLLhAH69krsfJmM3lYw9FJXDCATI+IPwN6sRd7jieAj9z34j
arFySOrer7naCM63cXZI1xFKKGgQghd1jexlDlMZzyDADtHIa51aMhWVkTQqK6eyQUDGYmQb4mV9
sUFVlELKPFr50h2jZKA4V/aXdfes783Ob/MbVY8utbTUQSXHne/Ph9qK/vSHdpflU6Chu8TNxbcb
nLJE10eE9jSLardVujRXbip03/nt0KZgqACyCr1RUMaULZYjWyIJ7pFj5bT+Chbs+Lq+3MlKbLCy
M28V5INpsXz1lFCY01UGgROmcPG7JD5T04uJV7pET4rgomILH6TFbdijGqPLfCd0PJfs2ZM75DUb
CE7tBhQdDB4b/YLTow8riT4nd96NqWtFvj6vS3sgq59ygxezukrvxQBUYrV9LBZf3QgMqygLVvsL
RCWsB/CrhRRll1FPkwM1+aZqxyDBLidPNYyDlG5ZFIUj7Kbw2jqvxFuWoLuKMHb4LAzsh8gjJGlx
Pd0wCMLhuHefJi6I9AKRCc6kEzGS7z8VGbYJhYKiXBPB00kTgp5Kcj4meBcakuHKTwnQcfB180Y9
Nqimpp9zz+8ZynFGSpGl1Lecj1X+obDCblnp3PQ/QHmsjp0DoqGw7RWkaeqhIWrkeKgmoTPmQFSR
Nge29skua5EueOMdceh6h9P+bP7JoU2zgzaDqFCeWl601MYzrWjT2QK4sO+2yEFKqwniHwmYDm1k
Lpny4I/jRRQYuOjbu3+5kVnwZr7H/JLN4/AyHxa9879cO+8NZYvQobOJdJfvCUFJXjgmm1rFyQxQ
UrMIqpJannicb/apjgoWE/aQlkrhJR+1L/eX0JfYbtU2lCfHpiQqoyU9AADshT/NrYAdk4JL2dkV
P2cOJBo9yOGnGi1TtawuBcPw2hUlyFUznrQ4Dz81k1jgRpm+soh95r16R90C4GSn2mufiGnlyUmu
wkIB1woiU77LUB4WyAoOw3i/YWtxx+NUKj3CQeZvwTo6B7nva05cBb3UrM2RDOAUeyndMD+X4BaD
GvCTA+/wkMu9LmxpeSiPAYzlOAJpfLQtoxrqVixNAWTCV8K1u2e0TiQphAibfzyrFyTyiIDst/+y
3B2DfWqMPJxz+GDyp9nwM6gIq5HjyzRvNo2WuY7VuE1KyU+my2FeJviLkq6Wol8SLETyHy7/3IJ1
rMXHVzCj5n8M2nIx4O64MDXO9l7znbR4zKYaw7OOFjIgjUbgf7ZsRIfry0mxVxCqRYwH/5bkrHFp
85fobj6eKXqSSfVBBHKNqyRiJQZEj3wuRgw4BvmsUEQWQ6dlnHTkKlMmixaaCHbpcCHtPO2zDwic
pjXTa6qo4UG2GN8RVNahmux3ZmKYuO7MFm3wAMs47IqPnva6dfZxAPy99iY7tQsV/V5F83Yxc6Qt
BWGCflE9afpS7tzEUtHjnKnT9J1TMqrLIG4V6YZXnSBEcdr6M2TCX0eB92KpPZBd26leYijjOeOq
IVCX7RvIvpeal2HvHCcFm3aEDCOjOaAVUdQuiAAuWBZ/mFAJ9ZZVHenMJ6J5hthPAvJnjHRPhxCG
Upj4l8rnnCn6iHARoGmiGwhWk54/suZu0bCBFaUU/w+IWeWCBVonuQ4OdUof845HlhCT2/cI7fEL
FMfzcyowPdPuapiHMl40ADx9GfyIVQVsN0jiOoyA9SqlNS01yVlsOcPNFGhRW4F345VHNJN+iLlx
PfcXD3e2/+h/JaP9yKPvRduT2RkAUwiF7wu1T0xXduMK9GNbmkK9cRwPjcFZ2++ak4fHcDG0WsbA
SB3Lk9j5veTbdQPpeMS0eITj4j3s2Wp6Rr4KVi/J6iSYdd588X5mtxa/0ec53BbybZ4h9XAa/Vje
dC5gzDto+N5qf5p9Zi6eOHuYnn8L/e9ZN/p0TlJxwvvrKaQdVn+9ATxbUYl4UVixasOvJhm663Ze
kS/sHMCzegkFhciIUosS3HsbuTL3T2wo6MHbPQ7aqp/BfdOzfb3ocFch3vAbyLNlUPu/HkDSnG/7
LjFF1Ov+XzDVV0Dj9gLwoiiE53ua0gXVgzCMegdbRBgLmzoz/4L+oCqCuqxYe6imhXK7wn+Li5Sw
2kgvtjqQPn+xLp6mKdAwidCYy43GWkj0J4+vyJJTylGOUOKAPGje4FFNw3S6v65fJCvMWZ2ZE+VU
J/7uNbzYql4GgsgJ07uHAPwZEMt737xUE/vax/RldjUjfVsJ2nU/9lfJrq1YsgD7uEG2eLtagBDK
SJkZXNw3z7RM/Gkc+T9JpaSU7n+sJQzTCODJbB02RIB4UllJ/c19KBZ1NgSSB+Yx1qKzvLGUOBW/
3IzSy3FB2kHWhJXYOCVdcZeoeNU30Fsz/MGCHZs2aSCG+ZM0mivcOgay3X4ttKUY5gz2MS2YEHV0
Z6r+BnIJAzbwZqkGVujNC8thSxUfPmUSWTMf0IeLUn0jwhOAJksO+ZViXCx3bQhwoCB4iyM8BmGw
UcrfSW0BV6afAgVeZDE02ZZngHbcgkZ7rzfSaD26z7HzXkhAA1q5w5BiKIDaH4IH7/d/FlJBTsbq
XnXNb2mDdRV0pJJAQaQXpSCLLrQAOqldHCLT7jqewUtaJ7Ttj/DCpklN/SLW+yje+PxZRruK9kj3
2VjwXyUVpMjos+hLF6/qCa1EkUutu/2jk6nnjZ0fUgvyftIMuzq5T5+LL8UmJxcwOg6kKy9p2CTp
djHZ8PPgJLcWbxiYP+50lMfLELXMv6djRSezzmVzacTp8pJabrWvtI6YMu4RDuZRWeQFD5m4Pwob
By+6p9NbTXIGNPgUEU7vwlnB2Rf+VOI0muEqbgR2gV+UsrC/He1FqxJCJluCXEdLZHPAhgSDjHg/
qbVVi8lK63bYHCYsl6sM6Pfeby22KprUXd/t7wka4PTuqxE1watkShzMwZAhMCEuNXmip8Q15/Oz
bqiYeHA/rfrtLemdGWlOhnI1mvRtT+VVna7Uee/OWHvsmCfg9EWA7HR+xg8Y8Ly6dv1CiQ07jYsb
6ot2yaRBI7F1/Kn9nKGBaDnKwaeZo3NbpcEpTyzx8anEeDsClaL/u0QLUjZsNeFbdGIHXwWakMLr
HHTak0F69Z5AJ6VN3U6HIEO06usD3NMSuBsk2/YwSkfnJnbWmSO8DjQdShuA6BuNTNddwUAoA9Ll
278LJHcdqgHUk4iUuum52rPQk5rOcGp7LLyUThu0XtbBe+VnBRMge+jkEJg0lm0PL/SOhB/9PGaz
KVt75mF8iiLt6DWKlyjRezPt5Z5GldMH+sIuTsrQunhv+HHSQ7FyxB0IWtXGPEcbQyH1IxMwxmcD
fFpB1qOIBzpFkY9k/CbPSprL4EklMX35Gn1m21v72AaI22Z9PsZw1NIVoV2uO7xKnKYCzNPMhBtT
vDW68MyUS30ytjI9a87YeIiy0ZBk5JyqIeLxNMk39EYFiI8eMH+T9u5pA5NqhFM7dl10v6vGfmMd
I+qg7lFE1/4TfvyWgwaEywuQUuCfZHFbV3ZrFD1f9Y64dGO6X3E7TAe+bHvWVB0BfDJGPrn4dwwa
yQttTNGt2wq9ZJ/TB9qeek319kzY3zCznEYpayOhZ0G5vRx66bYGQDGhLPrIZbtc+ac3jMM8gm2a
HLVCBmVVoHtLIM7fgRAFbZxKMG4E/XmUD4cTWrH5jtb7GS9nvyHOndIxSLmm3dAJm8IABuBhXWIL
3R4eQu9GNpFLA22A6ky7TqGw9I+D+dFNa0Ea4lopHIu0lcIcViOEeSe/Pl9jzNy9wKTKjliYaiZt
uNHMDcNEFYhXnaDOvKy1wLkgUhftRQBm6rWrjBHx9gcTHhpyI6qAjzdLkUy+GfGW5n3r6Lb6L7/B
r7zVmHZ4fBURaqB0ai/h6nqZ5WjiUtFnntuA+FDWrHXexwsWWmpm1O/awlo0NRLug7bkIUKjqsl3
6M6oLS4PtlNNoDbPHZczD6O3RWTeJY0dDfyDYZRup9mwU1b5MbBPfN9tEid5XYNtddOQlZTmed8P
K6SjCDmaJfaEh4UpxyeDG5VX4gj91nIwTmIcUwWsQ4/fRDTwv0oy++cvUA/oNFef20iaD5L9Yi9R
0sH8fonOT4CTXw0SOUqC9DehnKuKQvXgprKtNxDQxjq58YHsaXV6dGG4kiPd9GFHbISsvQeClbpa
+r8T5N0xkCXp/VHwTj91slzGOm17crbcJkZqD+2B86ubwgrV6bg+bgv5KULHm6PgSRSW3zoPHOIx
sKtL59rLxxoN/gM30h0URdjFmFyF2MIVWzONOH9D6FIM5kJblcmb4Lfbt86cCVCm/ZR86JhGZTcU
acfMlBSyacnGtl89RxBdHlGbK703Rheyugur+8LLqCejerkWp8QIbJCxhWzvjcW8bcU76+/C2JSB
942/ymGZvaqUYsNuffDVeHEphDNbUK1ijqp6QlRU0BoLk29bdT+D9Cw/fUK6xE+ohwz4tgVhJuGZ
VWJIqhG+f+4nsdcsnFi7Z9vFDWARKxGuDLerxqaqn8ChSWyIo7wIdhqEtAkvY10peMXv3RTX8twQ
wwAJeMXTfETKhtFLwR+UJ9xsygVQZowLnfdok73NJdR17MVLYjZ1+Gi79RRN84h71fOWUe6jlLjM
gz2US0GML2+enxhNZihym4iGJSxCw+zHMhW7RwoyxpoIipGsHRP+EKIDsS2++9WdwxkKV+J1tXM+
eAVC1TKeMXYl9nv2NcNP+M3601Ou2DG2LpMkZkIrQpdmhyiMMY/tDwDCFfrW9/m/R21kCbderOwf
bgh1MKraRq3muFB8W9K9H3oN7Bl6J1I2mC38ITY77aC1uillRFfIcAoL+Vbmr4r6onPh7B0bY1CD
tRY4ZLcgya6ZopgPGNjVRS05vy3qBoszT8RjVAkZWCViY3ssmui72bWLDyRcU46ohUFXs+zKYI6V
n3gkaiegmPKH6TJd7RIZD0J1Ls32sbJMgKE0+xJhSmqUhA3RVl7UQbRzNE11DIqc7obc57ZkCYTu
bnG4e2/3XOd4LtPrBaDqqSgysSJItCdIb/pnDFuvDnjYRRpz4CK4ThcR7lqTcpX1aK5zkVo47fmN
jlfksAslWCoYMh1ZCr9do3XvOz0JF5+NjOFnT54N3qw7RC5ck635lDIdI4zug6xJYZ0TuMqJ7OkM
bD5fd+VuRkivXdAxZucHTP9yBJqEOiWSd0dxIJgz1s3TwuGLFPvbj25F8PraPoSTsBEwpcskWiiX
GM082qGY2jxklASYdizc/9peAuTpXpULdL7lQ/EKSfs7IOl5+5h3XuLHY0EkXW8GW7FzPqZL3fU2
0ut8rOVnLubC4nVydJ0+Mv5dgBPYuoTnoDxQdV5vgT4m3ZusaAbzQk70TGMrFVSoZVaCYY2xZVdx
gRxs5DnQB3GPR5x8BbDKO2DXzU+3tQdf2UT/42hB0zhLCRUPtIMOkmUy9243NoQXUQiXvJXdvkPW
VI+I7SxWU58QKPQdiJToCcUKI63cLsk8GV2qAX0Z0U622NZ/BaGMootBgHj6FDkpd4w0T4suzfWH
lfmIX12+BKMdkphlYVleKGxo7JIEQTr5w5AZ0qDENJZdnqdAJxPTnR6xcho42H0ydaY4VZIC/5+5
FqWu4/ZdlsC6OU+0BEXP/CJkO9nvkpeQ7jDoXkahrMPk57iclR5L95StzA7DSaGcLiEqPWJoB47/
EDCekY4RBFZ2rojTJF2TXid3hWFPhY8wcnolB1UL4/TQjw1gP61+dCqqpJ0xQ4I/XcJe7qT3MyFd
/uVDtvbYU2H9NhDweFDDiB4i9vka69cZAqe4xTvRMb5+QyUMJI7l/yrwZ74clMWH/4g0piPR9CUp
7rNg66kt9Bn9/5EGOqszz/VLjsYF6lpDYGgDw+YT4BBcwGJs1Cj6QUxzryFl7UknvBUAAPPAzZwg
bOjQZaLqnrd46WfHO0/1L9xF3afzKzCs2Ol/IZiTigOFN30bE54w/jx/BNCzPyvdX/GbTPrA9iFh
JcmCr+pqQTA/CrMS/4IeR5NPrq1hkcxBwHhSqFvYSGN8ieWcP2nEWrzskS3DzOUn9dDDZz7lhnFq
VPwIrns+ekB5cI/MDYwndDw77mzbCHXSbWMJDJx4B1F+LRShft4DmQ4z61D5JYcdrk1SS6TeDF26
xYrT2bZ5i/LsClcTrqjd7KMJiHIMfOkNuXhwW9WY7xbNXCyHWmZoXn6qYbBAEb6UMQwzmgeJL/jm
vhAfjZvxxd8Q8VF6gefj2kYz8uhDP7Ih3f7sA31SyaXKeF61C+MNTr0dNHwdgjQmVPjLfyMoivHg
LiOS+B6WFlqMaY9nEXsNq7QL0W4AaZrjhXAq5YzOGfytwQe4ki8v2GPb68ScOBdXsefTTW3W3ru2
BjUFkwpTlMakSqh3HD+K9wqqbBYppe/L/RR9QwWgCsHLUW6+8uToV9bMO0NM6116w5df5E7kwrTC
CtP0xErIPpRR4rjAuR7jyKj43My9GsNXsnba6gHuceQtddJy3gbSVYN8328Pbo2E2CragJXVw37W
bkTo9KT71EZgFQlKR39wKU4DaM3Z7BHiVc3d2JBqgTUsYR2iqce1r6VQMK+h0TTagUbo1CUjBy8O
Flfmfc3WqUxBj+COKcGfV6bZ879d1Ja+/btvrB48py8M+ATOjoYP6+VYKxx5lKE0EkLA15jv33uD
i55znHOtVExbZfH5zi8BW6G0IimxCmSMFvAHOeI88sKNu3h9xan/XBXK6ruIzqEA/txr0gE8ATeM
cm4wq9ZhU8tBH60eTT8llDVjiHLQV8i+bDbgvnffYX1ZYBA95nBZyV6KYmUeCbWZiWLX9oCYpDtM
Tr6qkyJlp4vkTLoRQhiYhs1Ns01H6f3KIcGcUltzLKpQKdtw8BrCtjzFQs/ajZ38aIjY+ld352Qe
Pi29DQ/Uvqtztf/xDshYhld1Xm+ocqw57JYnr10eYSVeDh0G9DV2WRTSK4lvtAbcXEwYISq8W6lg
Pj7o2g042w/Oey0+L+PkDfvDmC3uyOWhTkqhNwsGLFaB1MVodU4dymR6flf0O0GX5aI4wt3dKhe6
9vl1ejtN4iJbXWO9RjR35m72+yNkIaPu4p00q0p92x94Ki9Xfh1uOOnM8id2Oivj7GUzbj5+GbuR
F7hXXv6Oz5EE6BgxhilDiDbLFk5wkptLYkJcVyE4AXVbMi3hOENPEpIh7uJoot6PwdZwxWHj10ab
rFGHHRAdDmTJKqziTgPpOhxN6QjveQy5KbkmJuvku9r8RytIHuF/bGMbHj2/gVJXd7y9gzdXm1t5
Z79WcLZJyuxaiaIXlRVQb7uUyeJGURUE/gKuSCTIO0iS1jRwZ61n97r++mu0Y/XwVdqNCcKwQVgT
LKER8q8OFk4H/nZKr8YNkDBG0tQkvD/KkqTNrO9TWSPAfz+Y6SAZ06TlaTfQtESuYuKid+lM/mUm
23zy16zLZhWeQI54d+y9GiBinkScIU7DAt38ZAxYFLM8gJ0MN5o2UWQ8bVsi9jPqFa/lVCjeeW7s
zOvt7SURS874AeewolVy2XZ1wudV67KRC9PhhFgKBCsmWUtnejPEtdOdI9eDfGLLnA9WVJeLzhGK
J7haQT4/Js5GZqIzIJ4zPmZHwOj3NAvxLB2OLN1Ct0EgngeEVflFD+mXwSibA0iqitc0VPUrvWVn
eQYgjYrJVF8AzvHgFx1/wrem2AvtiP40p82+bqN3s1+lgjLJDPATLwS9t9R5SCbE8EBsT8bVL3VS
vvFLz1mXcT0W4OmG1vPPH2l6m43Ww8fo+51kCgOsZ+gyxKIO6FOk8d/M0eBQLizz2Oi+uvUO51t7
DuwdzIgtk75Rnbo5ZsBGMdTzA/Ilpg48weIdvMZMoLOeTh5BvQLIoFo4OSZCENpsA/Md6HLlumsJ
Z0jGLFap7DO7yzo6ay5l+0n/nBbhZ3TS959VrTfTwVWri0zZm18AWNy6FON1PHezac/PvjB9/Dhn
jzMGekxCDxBV3AcRBpCAmzdq/Fh4KATtnPMI63CBNZxN7jPqWC6jMWvHVcgwGkfwGhoQuhuWUMsK
8eoOnNZD3fgT0vxfzL2fraGP0ztQyRFQvjm6oSr51zHhdnak2jMBWQgRusxhrwN1AwpoII6mKhYB
VfxEw+Le6H/+Tk6goV+eGZmX6cQ1CXiaJrhX22AyYOkXJ7PN9/fUk6HqqgGK2KJ3zLMRtMuwswQC
F8MgNCtNiucyrBI1r0oFwFgIcGYkDwi6PS5MMK3RIVMdbPwml4Ty+30RXfeObin/wAvmXteaEhJt
Z601Qpl+M6TOBYAd6Ntu2Gt5T1ewec9eVhxhlLzoriE8BJ+2aEop6Uf9zDaNFRFOpJccBa42D6Vz
Cw5laSXGlpGouWhmUOwkNvkEPsejS+ZXIkMowWBsijBFGwCA368DOCErUU2ebCSyuJOykpS2WEO9
ru4jJPjnQgwuAfjfILQ7H7ej3x6qbOy40xbMqiun0AztaPAZ1xv1GqWhIZRe6hVc7pjKv9PDnpCA
h7rPHwU3fP6t0xe6DSl6qima85Cyhdq22wUVb2DdNE/c0qCUg6OqfH0SY89S5rCzKaljyfQFqadc
vo51iJguQ/Bt75c8Jq6iFmAvm4S5iGSTRLtlb7AcTHmTwL+7L4M90LsKwZY4zi5KYOPO6W4DJM22
NGP1BcitQolWf7Hd8mkr3h//V1NNdwPuPW+KgJ5VnFNa8LnTvTMeuI7UKqCTBt4/5Ohv5ZOareGn
I8D/dfEKtfb6MJ+QwcZUFHdhN2MsJ2Gn/k8/kQZ/aAZ2Ba2AX/urnYciY9BLVP3iTcxjcwJIoR9a
UEIlV6vlCWawYGsDLlKp7atwLy/9AdGHXq9eJV18pC5W9epUScHVf9O3cUPcUC6+63HkFPUSHFLs
69NlfEo6+zVabOdJcLthZORpl379TgU9VwtGdb3By+SsVpBznsnZ7sSV2Z/JfZSwCr2FD/DG6M6f
3ld8WKKk35XzY7VRZ1iBQ7hlyEoCODL7yT4U160YKrWwITmF+QXmzk98o5WbSl/vtv9rqft/i1cc
UEkqgmOIVTtjVZqj4jorQcoF2P7wbZRUytzDsuu+EVfQxJyalUdUaUSVMvoBXDHrfDXcbsygn8Vj
Ezl3/J8v4ZED4RW75XWfTHC3ENBPPFQLFNtCf3+XH7bdfAN7asE8gW0WiXK+QJVqS6WyTqwDp9aI
WPYjKLMogs/DCuUx0/4YMRdLqYn5ql41EvVhUqdgeiYnRUUAryU+UVoLQn/tl7V2x+h0hjqlhblp
rx/Knm8NtVlSuD5rcA97J4b1HlWljwdPXhLO0Rt/ek8mzh3kheouuog/3+G9QxpBEjtXnUzoEFJB
+CSv1D3glWOA2ue3+HHVupgwpEs+WtYaxpXiWY2BEjw+bYN7mRt9kme+RSSQsvnboXSMT1NuMKHu
bbg1JWMFBW93evMdt7sPrpWvI6UWcl2ZVj3N8vKAACvlqKqrHzr/aSdm3J8A8woRwIrz9za6c5ZA
ll4zWwVKFlZ6WTljfAchxFaCtlWNO4z1fZ8euu3+QrVseXyM3qh7ZFsfDP+oU1B6dvr1El6tfKf1
53flRZsu/5apa5LVi7pO92k5kuAYjyyso9rGQqAin5Mq/H5hZa4ke3DcUc7amWqELTux37CLpuNW
0KtudcX2LW45rq3E0/oSbsXDc4fEy7hJVgkiz59xt908f+3ozipGPnzS+q231/vfz9O8ayHh5Wb3
AcQB6gIdeAJYkt6qc2v97zKxJAtUHbmeojO+LF6wtUs+Lj9VYpEi5kbePSLMErGgkSYr8pebFawp
bRfAoWE2/MWMelOQj/4wG46qeIcMfEcNoaWU3JjaISPbbOxmZ6J5TpSHsLQ5mxJkJtq78QY998qi
C6pCQNef/z9eqIEt87RlEtfwV3Se6HRfcLbvtz66Ny6n2zmpJxufbBgcVl+LdAbUB1aqdm302Ml9
PsEV3SyUm5T14jyqDTHPnZvhK5UnoKlObpCMpTFKFDQBQQLx2B9Cb0LfvwFxqpzlXxpa5J5oqyZ3
QGYPMPULKqalM3n27teBASzM1Mjx8tF7gGHQkNYZJumdrh/2aZrXW6dM5kGklLfwhRpDIPv4He4D
t2sGs8evqwuS1++4j4+amuh4xfqqHWD/BgWCX+Va3sBBsiYRS48Q21aQr6jTDlEpy88WcWwW9uE7
Blhs6XvuKCVfMKVwjQAFSXnFDMX/gH/Jh8Eme8ReJcIbVj6sleYOEP9FBdkdtfRFMSPFBfsRgqJi
CZi9VOMKsPDd2z4y15apDtbA5M2vo/r3SWlO0OzvTCE1fYd1IUnm8S4n3Ce2uRsZzlLDkuaC311R
3mVCjsZXEKUyExbw1Hr4J9WcBMQs6+NNWfV4tANmKzICKDAFiUFRurxR1Z1NTEqMZfDNz73ZeiKh
d+GKaKE/zyDRb0dQnTettq5MZdRZNBV7zuWKCveMG58fcm85OJ2LtTBQbI+zxLkUxhU8lcp/XBAI
BHrqTLvnc+GF/y0BtWGj60wHRfZCNiwRw3FY84IHtkhumWnRzWCqSg2clYPpIFmiJzL/GtzYN+na
pVgIdZkPTEmZWMOe7Qg8HU24nLII9EebwxwNI5PwnwyJGTPUsZtVb8H4staiDozkYFYHyMgOoSJs
Gm2tbl2x+0MInMNgHSfweXCerfY2Kcmg32FyjCIrynLUjznAFXGJX7x3heeU75Iiiffy8H2WxosQ
EBSb4xu2FKR6xJ/HwYaJ0QL7gNVxxU7UZKua0UWQezPZGEGxHdYJryLozLH8BEBqePdU6ZatS0vo
sk+9SB12U05Xn57Uk9eGKrFH27AwJooZjQKQ/DdhIl+SG6H51rty5M5JGQ/OhkrQ9WpdKMbiXzon
cwsyqo5SXmQXQyKcxmKklSdVU9bC10Sx24btGOVskzkT4yOwaU0t+nHObvHTfXqOTErltisHn7s4
uOLZdgH39dqyST2AqBDt/36czj92a0R5aCbb6WZGxddc1cR2lnUjiRJrZBZ8ZWGCmuaKHhpLem0X
dUTn0Ss860yuOrJIYDYRXsHmbTXvcDrH4mbOr68F1czyDD9bLc82l80t4sqwg1+llB8bxQe2aB/h
lCcriMLcexZtBhJqQKT5t7b9ltyKR39TYDuSuX33oPflhFT3+BxNiBvP5+JElJzIV03OmYggI7v1
jpxt1h/k0K5bu/uZLLc7i6hi1bnY6SlloPH93nLQOx4hVDMsX8dddBoeveeUQGY9I3CeXEIXH1Kt
/9iMQRwP27FxeNFaQAkTSJChfol/o/Xw4u9sCqQeTNP+YLf8nSMGw0dH1fIqkpmI8xg4ICFDLcvL
ODcw7dK14mqOiSp09j3RJDDxUfNFk+9CPwJgF5mKTg1vzXLK61jVNysPbzGDJ/OuRF/+g/xtFMRF
JRzKl2ePotWYPp+CT/7W3ZswVQE+UKmJZ2NlLu+UNE1OFoEzH/aVQtT7tL1yu2ITdNeak2iH/IBU
/qfb33laaQUSkVkfGeF/kEZgNgltbEMJsOq4iE72NNIEbXHiiTjnsd0UzBkpSrpT/b4IAagNGowz
lkGvdfgaQeeIn+X+wTxzyHiTtKRU1CRPa7gwH15UVVC0XWn1+NuVheKeSQamt/mdIveumYHnktT8
KpVC/YYdjFph43lNgPAD0i8kmqW6f2gjfnrQciK2a1Ie/FfPyCMfaJ/LTqEzNQGnX5sKmL/CUySq
FufxaIaZRDznFkC9bD08TH6Hha7hluHQOMwyTENdxbDNQGy/MqCVao4fifuQawITVBsHyKE22y/q
VL9ThHKky2IFGca9kRPxt3V1eX3eENF03SZ3Bo75Fr9ufYYEFaDnJcay/3+bg3cZ1QO6LLT9o9om
s/2qPBO6c+P027roI+9ELPYmD4tDMSrWwkFSx6UnbvImqdypQwh0PldBxNhpli/HZMTga6taCHP3
60cBju5v1GauaqHq9hBYnyEBShK8CQZHBUSEGGhO86/ul2Wpb/UXfUb6nVpPRGjZS11cRT/wh22O
+9Q8gHf7ItA0yQoNqcaIjT22ygti/9hwUoBdSU20laRzGtOYZ8V06tF3s3olSF+rHwYNJ5Ag6XI5
0YM8r0NROCuBuaa/uBhyi4zMzBSspipStYPEh1p21nwOZfAMxoJ/fUT0jg3E1vpBepfGFyLnG/lf
WcMX+8Y6DBiIk6DIkNOCrPmLJR7+SgxkFzPJKjImx35r3/HO4rZa3MMKy1SrBxvlaTI0iRSFiAIj
FDy3vvAd2fyeasYFql9UKJ/wTAhs+40bWNzqNPO9pxCmZjmBCGhCEPdXDva18MIhpXxighT65Adm
UTVlc8UJfQvDtrIdtl6SZtq5CeK6VQ33wFE6STnEanMfhs4sHZlvYW0PSY8kURiAMGRoQAA26/jq
8ZSnPuPHQscBL72vVa+wVz0f2gPe3AS0TxFZ1gkBrQ4YySAR4bOy4sXdfx0JNKIRpmGDuw4zjY5N
FJTqSynJcONZX5BsWiExRl1MoApcjOMAGBkL6h/qm43aJVLTdFCbBsopdFWOcRdvdoQa6YXvQ895
ylCApJsBEaB0fMdwtlW85bCny8Xfv59zakX+z0shGDDaNo1eJ8srZSGSbxKcpBGRItzPv1yTqWjg
bhYQ6TRNh0qDMwQq7zG4T2RQuGFqwNPxhYJPcNyALDbed6f5OekgwKkAxQGi+IaazsguHhXBX/Np
KGf05EAlnqN32VZNi7RvQzYUP/oC46+g7IJ70C3zU1yf64qmGe/4SbvUipHz6S5jLu7pBaqtFokZ
EuVdOxkJlnKcn7eqtrXX9vLc+EzXYSBmm6HdDXWQi4fMfSez4a51CsuB0OCyHoIKboVzT93K2buG
eUbpjLjyGrHmd/nWnKc4cgaz/Tp+PhvxaI/xpNasZ+ljDks5M51f1bPPim94hdY7ELxhAD0GTvhy
9spNxZCtF7VPQcRGvgLTs0qD+MzCvz6GtyTlzbaVqsBnylbhLDtBRaKkNI9DuUTokhpSUb5bxBkk
4crfBr3OofW35MwcdCieM8ABG1mgluQM4qcL+3LMq0YiMYM+jTOju1O9rJxERkQCua3kl5T91UL5
1OV0B8U6ZExy1LDdrymEJkkZZAszUVvB4CzW0RVqC6YAS58HO/7Mj29ZCfHXRbaveE6Ujr7jFFY4
00A1ojpl1Frqc7q6URhzl2WcAH+1zs2waRxFYgpCNJAYWH27XSA+3P+sehl6yeeSSoXhm6+CbHAJ
SGdvOmy2uMQUuLLz8/luZ1G9lFyEqHjH3xkjNgCHJUOpnmWCk1dtjcM354EKdusJgEFXP5hKP3pd
00HWIElMfY579GnROdrezLz/LUAViJ5QLqtXrWLA2/TmJSMLK9oX778DoVbXWg96acxvCkwnS2IH
/VKJAght1y2f/XdWHAIVlI6O308ajBe7WEb9pb0lWIzFIx/K/wdHte1XfC8GCNao6p3Lr9Y5veVG
x2Zh1LjFQ1yES9Tan1jXd+ddXFSNNYVUTFROd1F1OYASso/E936erelORM0mF5fAKAUqfBn4z8AE
YnVWkqcpMFZ3Z1h72l1Z0z5p8oi4CreQ2z8kk7JJDwRdIeUSAzburLZrh83IkjgCHZaxEvazrvVP
ydH0Jthtl8fyraK3HDb8q0uFQV24Kk/Q+LHicpY2G0uTQv9IZ18AsbxoH3L4XxRjcy0w8y3b+N1d
4jE1eFuIRfun66ryulmeKGZsx09tg+2mtDh1neuM+H4EpXw0/dXPY6WIZJiPQ4MSTVAZkc7hdtAz
ssFOCFQkNbynY7i4cBfxTJNhSCH3izJfBet/idzQ77s6fTMszpyA9xWI5/DOdEh3SbMP7zi2fucd
cADyppWCKCn36kC4GZr6Ep5L4j8y2X8XHNewJYtUAx187YkU/4aLeQx2iAM2K1lnBtYQDgFr/ht/
A0hWIJ5dlM2i1jM8/jBt7ooB2l8BmDojj8D11ZhJUl17vMaiy2O+Ncz/bS+VQthsPzUfswWMSTaX
gf89MLsW0LlsbdBsaA1Rv0puPaavBSWtu0bgVv3n4ljG/B3kF5ipXTiBR1RWChadVThEUPWaZQDL
c5kJJy65oPwAioI8SwhjqqcL2fkriFAXmbGeK6L/r3s1wlT+jyb77e3F5H2jGd7/jeDn/V0ICwGT
zgY8P37DXNxDJpKMsRxq9RgP6+UO0MhQQ8pVtllQYr+4c4VXrS9CIGii27GIW7TX9ObF2GqDqOol
rwtKhcB+ThzNuuH9Rr1spGU8Aggaoehlh+4TL8XIMdUdne7PRi9hSKlBmXsgsvpne4webEZw8jEM
HjfUAwRvErdorVgRkK2k9rsYRzoJnGuwlXPjebF0gs5iM/qJpWiZIvr6NAeTyt73kTWMFxtr9QJY
at+XKj3dG0nM1z1SNZTAN9grQqxS65V/yiEJQl2gMdiwjPz5nIgihkkCWRX0ha2kz9y+l9pn+3ez
/K6XL2dEwglr307jYBR5nv+rE+4ORTFVZJ1ULd71NXk/zEdiYXggUF4l9HtDc4EHQgDW1WpVWCMq
B+IZk9KntPbh50mj3nmP0RR6nsX3Be3ZGQ65iG1zQnnCMCEdFJedQ3Enn850egVzHrN8WRaSm8Ue
iYklFlQwwntgsgI1bgQZ5R7/GAhgB6rN2wAyzST1eppxiLDA1UgfWkncdPMqPAvsB0m7Gw7R8arW
cjiR6f+iRR0HrJrhUQTGG/D4m1+fXlAPZZjvUnjKztztTXgGLUO1ecxXRB6ww1KImKH69p+9ad8R
lIMyzmQjuVQHfHkiwuSPZVjQtuMSO+DIUk4cNu+uUKHuFcE5rIgblahe7LCIojIhn0ZCYt3F9Yp0
RYxezOFYkJsph2KFpkWNYurs60aLg8f2CnmuxcQPV9slEbXEpEAMNGKeRIYiaCx1YKIF+abTAVIa
EvtYnIDgAyYFSpw5GeWiGGqQcmxxQpySW1BfG0RxdVAZAY1TiuFlcN2vXI+n9DvqZ8Oavr2Vbvf3
zwSigXX3v4ggKC9GB64jrMQCZpYP7qFw6kAtvfGBnPv8XH9BO+csRa4tbW0T03AwoINPvAth8lGI
q7aSHj4GT3cZyas0Wd46s+H7CtoqVIsMKfmQ7TjwXuhH6pFcJPkwra+gyjpbvSNZDbC1uHDNRzcu
nCbGQWTYg0UjZP4bd3nu6/WXboow8xsVRgS8g8meUaVTT4+e852iL9+x+A3vbukpxxMDyTcSmRSL
JXiEAk7vtXdxn1CQzDwHUEqwfur5uX3Iwxga5LzxUZ3DNBdfuCUwleOx3DLzLSxtOXn4ZcCAnLxw
hRK9Bl/48Et7jY70e3/3Qy5zF5HKTE//4/OJ0EQ25Lr6LGH1L2L0rJWGDkc8RUkQBhAR+SemSCd+
hkBZfWksJAvuJwfM235K74ck7vlNiY1WaJChY0S8TEXfpY2gRwFky4MUPnknNR1GgQ/NDO8dyCAZ
yI6zhVOQ8UXRAS//3itDWm4KzTzvynBaGrczX+4/zvTvKZKt90O/HjvrgZQ+pruEYDYSQ3l+kKL+
12glav1ARpDe4sK2WeA/F3blYAwOhULoBqn9xd3me56R8/lbdbcAT4OEL5k5kZPZe/3jgpXsrjeQ
mGzyaIDVsvebt6LqaJ7MVj1Iopu3xiIExJfePSLWcTZjZCtV7cnyDjz6DUf8tI5DwKtS4UztaGE1
fvO/cD/yyevGg1HgPVMHfiVMi2KIzxvDg1opS16B2s7DOMV1XSzgUuDosRACbsEIknXaPmNp90MW
hWCo9XSTiWzNMFcBTXbHdKXlygK+26WIu29K60Pu+v0z837KhJWT++hLcqusETxwb2zYBABPJkjm
xR/Cav2ppNfk/g5kvaphIb29tXtjd9keYkbm6ZRGXkHNcJMzdQp9CiRQSh5pdU9SgqMCkHwGquV4
zhZ0VaPGNm9gm2eg9PgIKlq8BfIHs9RhbxFjhz5f+1Q2joyQ+AOmbpGx1OeUAbBAPyLp1YCSnvIn
7zV2/RqHThz+YHesNU7h6fGuNJdqcreNSVW6BWhZk3JFDZWGW3QOxrwWSC/I8RQRycdO2nW+TOVb
Bk1zpshfgVqYgVkhTe34upJfYbo6IGYM5BhZmG0jwxWcYeYKM5vUMQxTCwJO0lDVqv78G7P5H31H
4WyAC9P8toa1lws/yOTy69+y4V03fJ4uUd2g59p4UNiD0UmupzuE1biPuYryAhtoeh4pFsjS21XM
yzkcAl7mVvxjmaD9y7lUMjDsUDGNntW4Vy6TuPVY6XgVjU+kGO9CzvWDhkQUhcovyPOpmx7iIJnT
feUBa7SW38v2ylayJzXTm4LGJmiEryzX7DABrKCJnkdQ7zbVu8zt8R6RWByfZotue43GdKyWGZQ/
PA1kdG+osxJ33XivEesTAB4F6K087H1U9aCrdExfYGnA/rpEVsjz7sWAbtIoJxYORltMnoQrZ77y
hrfxSuASXqyUIHzWDuzF9LIB9dD0gQNNmka9vsA8T2PfBNoSB12nKlZQ2GAhzo9MduT8WJz4KjPe
uVUjFU3iqiG9HU2YYBV/UYxZOCbIQIC3xKdGOs8n36LZeU6zZi9x3fvw26lENKesupGX7URHJ+VZ
gghKIQGNqSjGO5SMQQx8+djqXiwl+1JDOhLl0zQu7BfzIABu37pUU4dNEpz2u9XSZvs2i/Y4I3gM
1dYurdQ5jljw8/qQWb+D26dElO0844fxkP6KX6/SKHZOQx5TFA/TSGCftKU76mr0fD/zs89QaPzg
VNTR+W9h8TA4tElyN0O6kuCKdwH8FztJMxIGkoRoJRnj3pand652R3tR3f+ivO5H0AxGp5OR83/v
vc1sXzAvH8b4KgNmR9Tj+TyVgb/O8As7sn1ldhhBBT4bV6TmDnlwYhCEzUtu5ZEEEg8Oc+G1mZTJ
6suubwTEGvkVZE8CJSZ9cKMyyB8aPyFznmb+eWNcI84SIs6y7tGXQeGSQZtJpEysVGB4hx9iEsu5
O2doXh9f0aXFqxEzqfSnosiKK1IaciXPfwkGIANutryHiXgl4Snk7j4wJ5oEDM3TZ3OMVBvGZnQS
MVzHzEmmV30RS6u+9UQlfy8oiAlRkJg1BvBJ8mM7LfnqSHd7pRVidEYwKqgOURZJzofRQiD9tqA4
6IMunwaKuZTBsbdQ0zQU5g//rUhVaSzF8oEyaAxSpl2NN+w5z6IgpcB9TtQjLxL7y20J432ZOkLo
Q898tHDC/C9qlvX+ehX/eS9zmn4phbiWEHtkqlkqq/NHuqCJ2eSJLTdVKRvG+1tjuGvI/X8h7/Ly
167Z+JCGmLv8+D+MmEs32vYOayW4Ir6TkuowXH8iNWqxRi4ki5c/Bm0jMFncZLipsI6vdCZSU4eF
71LP5vlUFe9CpA9ZQRASt/zGB52jpw34WOUGos+YyroqTcGTXxHA+ogXjDlUkAbqylVMAB3RmsuA
sSHom9+zk5ngDkj73XJzLQnr+DjAIyYhBwvGg2aqPmCERP8gIQreMjNpJbtySq2RB0xioja+cegX
5Shf4JyvJkgd8h9tACC5KNeyol0qOKQ96Ivk35j8+MKPJU/+xejBhfhL26M9nI6xY8JbevfFghZ7
uq1kJKNF2zebtLPmGdmnAG94cS4rc60XzPU36In011pEBWHaDOOyJ6/Q4xdNTLvAin/yOpTjSigs
MNf3lv1fL6eYlI9eQsBqrXsdxpk8SoR3UoH2Tox83KxeM7wvkSwdOyCNNwDx5U2DcsQKnsDYwdfy
e5QPBX43/VsX8bB8T4ygFPd6dTguItNvOf/JMUey2EhJ3OH9S/kMuGqdtY2bG0ZM8B7SAgtFTvy8
vqwDBVxvllS0xMKk/v+om8ME7PTYqVTeqrEDw1Dv/nAAdetUQRZ1eiueQXwugts6OzPsilfcwfit
BalIs557Zeh4uOiyHQrZdbMdd9jSTbdS9L4nixm5jAYb6pmfhSev78yqG1+4E8DA3tgoG+/uUrzC
AZnYfRt+sEGcNTc0ROntG5O8XLUvMbJByMtijvBQ5vveG9Nv5oYh6/4DR5+WhU1lqhUh/vWWybDN
bbqJyJBVKk8/hLnXfYWLi52Gjd4t2ECuI08vd7la/h19ddL7ZbBDszugudzFPXI1m7z/ngc4V9m2
5o/prGQGCxPcFo4lxeEdsSEBjWahwaqWa8jc2UsZQhDSYvVnflbx2BZa3TFVhdyt2Qi6Vabd73K3
caYouvkTIJCWKB+AncO/xekDpRCdpdAESW0gF3uVI3op8Fd1uhjweIuEymmu8clNqQ3t6VMxv2Nu
Zec0d2e3tftT5ZgQ4qkDypwmhZ5YM/YVU8Q2Z9GsbqRfGNq5MRKdN3xb/TM3n89iRyN3A0kKr2+5
9oiAwee+pZ5b0vDxf6gqYXWmTPWnhkXylxAAo4FEJ/EsmRXKX710NururJ4qc7Xjl+MwUjwa7eCp
T4BOzxACMEsYQzOXcxRqhXxyVpXheHEz/fclMguWNryrCSIydvGuoHaUCFAMBNVX0CuZtPGMwtUp
5qRhU20+mdYWTUUya1fDb3gQKo9pUZhyKOYDcEy6psY7KFnkAKjszY0mM7XyO/NBGSNZ/nHyprkd
l42+n6hejRyJNMHOvf0iujFiaeQeiTFj0/crnsb5lmqObjj1+5Se+KpjiJotB0iJLxuerZdyzA6D
kdQdnHyEwUiZjuFS8Nl72qRazPDndeFQc8tqRSIjegG+xpBsWqeGz5FN8ObyG0FYXUHpW10d8zLv
IB9r5ihALZVcm5XcICrGKzrxSU+mOtLOndn2wtz3kYv1Hcem5wwV5cRj8kwkmwN4OKTAloyfyfsA
1cNl4jFwDwD8Bsu67GCfboQ0Gsr4GhlnE6NhwKi8m+V/xZ3rP6HQFNG6A3CQhrsgWQH6JHWOzrWJ
bPpfwaertENCx5Bte27E+NFrGTLhfnYz6dkFPzseuHfG7zazFIT1v2EZywEnOJBnFeAscrh9ndTb
pJMSk/GWBwdPHoVlNv6E9jWvbyGDXo5g7LZNfOcYvsoByIh9QkDxc+1tVFCPAaXwgYyFX6nK4s7m
pfDFKCpAqHBSbAsHvboSWTTcZHVJUzGs/x3l4Ry5VG2vYz5ZQq3PYwvkSJfSXzyGMoUVTduz5F/p
Dd10V32lgJUB4SSaYMPT2ZDYW11Dk0CmcwaVjjRZHnEsnXu6W2HcfQkPozbsLTs5N6bjYIBmZgC7
Z6zji8qfXPdv03C8bTbQBTpG20bO2cnmNMZGDoh4bDkK1pAkC+oJDt18RUO2sdvq7iD9R/EP7gZv
oab1ED/5wYHWo7MIKu6vizGTp1PzCfJ5eRd8QsULMmpYkoR32fPO+U8pdjnjiKMHkil0jqJhyH2q
LphTObIjSlMdPSASn3CT1clnOBXUJ/10eDWB7p6C24fCXCgyIXITKkzb+TD7Z6JlFF/0R9pG0z0w
9jSgimIXvOrfJCPgxDdesz0RAL/et1C36fc4+OyFAGd/8m5e9KkPia9kF2hZaIAfTUHv8jc+iPmC
aY9UX6mCqKhxQ3AvQjMfUha+YQUtRl+eIMsw+NMRBgjW6WCwXXZu6Cj+uj5BDE9XJOfuRqwX4Ip9
sgVfPKMMIEzljy9J8VvSZ0rfWb6HvbMJ1yZrm6wURS7xIodOwaThUBqS4kVnP6fG6xcvWSLchkMG
V2dzIhE3u+CGNMiiCstUciyIZTaD32VLvMuSg4D4xLcJoK5UG/rIims9l8swPa4PMkY32RyulxiQ
nGpD3sbCF0FkaJz7xctL552NFe19HxNVbiYGsTBPJJX25dldGJPO7tQytfIR9WSKzvrMfj6r5Urq
aaP6AZyZIfrGfNocbZKAEA/epymC+OIvmaoXAxtuE3fPEHQDV6eSm3qrItyBrsWaWHGddztfAx7B
1p9i4YCXuaGYTyAMrWaAQnM3o72g4ioMW+q6ZE16PSgWtb8mSm3sV8lj1Fso4YwaqE4SJ5N3FxJr
Fdppt3WYBUBh7wTlPKtocVaOGc2c9/bnhLYlFrXT6vLL5nkslDygEpjouoi9AzYdjUEYHkEOLxMu
zFrcNmt4zlo86hHnvG6eROZr+l4saIvH1KnFtMPt/h7Snk31j14hEgyYK8w+u/81cESyjukXPsQy
R4FGtuuMlBbOYa6ezH/sJCKlaFAOncQ3n8+3nI/efg2/8uQwm1xuI1T2EHGUEn5gMdNca+lmKqOs
lbKZ9f7Xi63Doga/fzmbeWx7a+1VyjH1tXghy5aLgxLhuXg4ufAxwdPzRbzQwg2049HTpguFLf4x
YvrJabfqtodn5LpvuT+xCvHVapvlIvXgT4P0+ZJl81M2dNWsRTI9tQWCEXAz7WDo3MpHxDqpMIeg
A/G3/y7nQn12VQ5AKyk/B6M227iibt/ScJ4HSi6i4CcTbPX/OhHDzZ6sHoInxc43f/Ugj4olWrWm
ovd/xJgpUoFfttlrFATPmsNaYmNnLIgzDdIQROgtjbSx3JebH2AjUiSq0IaqDt6GffQ/PCHC7O5s
lmerV0XkVuZTDXrgpTLfiQY0aBF3VFsgHWPFyVOlH/kku7kMu3E0JqlnHYaT8lEKQdMPFQw7xZha
w3BIMVfr7JnWrAxJ7/x1Af3WiscvFcmQF+sR6XBhr3gmnsb/EYEhVHW8fEP6FKA6A5uFiMZEXvWr
EpAj3odC33lm4FCuJas0eIt4pE/hFN2ZHHDDczOeRI85eHWOf5ADammT+nDTT9SR1l3cBm0KJ/c9
1R5EylVp6hl3jLUsxo3Oj0CiAIDvfGHthAvo2m7DjQcRzO3GVRsll4KbX11hIPvc8K+sslx/bHSG
16n/4yA+WeuLXrnmbzbTSODdW8U22JnWdqH/nnH9b9l7IAQxM9MIJYrghJ1R+15psLoGVoBDFBSV
Wz1jvZvmYS4ATsADvKiOW6yRQo4UfHMyaSfu1wzIVqamvB0MwhYbXpKn+RBWUZb02CSLa82eTn1P
Ss22iongUfCEHxb272TcQy0jaS/KHcVGJpWreWvVaNUYEz++35U/lSp2+2Pbj+IBkZQh5f9GuItf
rTvrfwpjSi+HvSazZIXQic9oCH1SUQKYAlYKgfwZ3cTGnCfxdcCEvefW4YeTjJsjibLsaZFKca5i
wpUsVF5ikhzaOK+ACpK6YRqQJyGRErZEw0xOe9dw5V9G7JaYt+ADh9fzZSo14mpx+E5WOgZjsNzb
ThHu1BayTy1pSjo8+naFFuvpIpUzkYHUp/LsykzS67Mzof9LZIdlNkx+cItWRdWZEkbbPC2XIVFB
bj3aAzce+PuBdsJXrF5gUDGJUg647RZC7LSzCXIaVWKCYTV2Fpr5O9zdWEQWg7WsGgaUhPejDnDZ
3yhucuO5y5LQKLCJGi8oPWYGgnCzL9F7FdMF3j/tkAtYD9PPiWNI3n0WRdKw1sXV/9ukA2h7yo+j
smlSf1pzKxtzsKlKdB9d79/p4gxVMCU3c0jyuL5r0mHabdLE2EEwRkir5CXjwu/cWUXfrzNPQNYX
tvyznYq06ljVxZXlPU/MD+r7fwsNBFsY9uh6DrDdoqjxlcoMFP3Yj+qAAuHqTsV0eBWHr83jqnSG
8qF2W3YojYJqDJppm47UH1vAoT3haHJu/0VVAXZKO5vCIZKXY/hePlEFM91mL40PNIhyI3FzbHo5
pWgVCoEg/C2yXP0AYK+RYeg3a4ENnsjhkpvOjmtE7q0R3cRsCDJY3Ye/o1o6Gs3JWhHZXw6YxWlx
CaYYF77TEq9g2V6kznlGmenN3M3H9xgsI0Gl2Ku17qQwNw+PlAZflBW5hiFYJpDehv9On+W+8DPx
rOdohgwa+n4I6XTqDKwUBifvNSH1vznZXo/SRfVYqvI8FSSYHyNV4gpW3FqEy8OHvBMcdeg6giN5
6ZW89jyH8SwKr9t70VotS3rJTOJdsk5StaXw6RZv7K4Wk148+ILLERGHwaDpTwG91n7MaEVUun8d
50DWOGEqLfCC9oeHXfxqu1SkDGowefHLNtKet2URKeq8VfnpUCruwjkO4Xs/8ukZdyrOO+/bX8/A
ThgSKBPscLZSOLCvKWbyAKXXDeXF+IbEaM5fc1Q5VmZVuU+aeNSZ15hgjL7KRAkXFhu9KdyNpZDN
yD/kJkhDK1uzySJTd6tsYe0tIRvBIh1AyuXqxexz9SxdGj1sCMAFflaTSAk3vfIr5S0XaDsxfsad
C3S9wLpDEec8tJeHXLyGVBpDSqi4cofPQzxXmPNMufTmuj3xf21lCXd29HKUk6lnDlsrYfX/oX+3
g9UuQLX6/rIKAJ2LAvw8YPGnh9ALDB4JKCJhJ63rnrkKJ60pdVKlyN0mGSiSpCKksZSFg+WbM/5I
8u97BlbNDN3uX53abee3hovI++4nFwuN3x7WP8pHADOwQqV8Na6KMJC1JVEIRrs6KdqQTCZghoAx
7Y6zaeUm4Xju4eQUKBZ65UINt9BAbA2Hm9hztAQ2Wrdmum8+edMIFhMtBZTKlTdhdcwWzSvuOuAY
JqMGp7n3b8eG6ssFKccVeO6PAc7Zp1nGiuxmXqarz3dFpFjdXqUlN6ADl+FxrpiQQWdCtu0rCvCw
pARn6m31YUkQwQElTx3EXOGv/CcksE8V9VbBBFaYwmn7P0zRjYPtZqzRZIupMZ28bGReTdIUVc0+
tHQCi5pEt7Txl+mzJDoYH15BCE8m6JyGNSvSzKmyILRcE2kDLaWyd2nTa7B9s4rdFgKm+rO1zydl
GHMY5afr6RRubqnhxQTNnc+LA/7DWw1J++OfqUEFAYYO9DLsg2icI0a6k30Xb/TDu3aq+rZyZFN5
l0sqtX3keh/40Wvwuo5B1xziABdALe86lhwpKdV3jUcRoPge8QBEsgi45XmJ1EmqQJyJTCu39qm/
nbeG00kQv5ECt0ZxNfyVkSNYRdT+5Cl3Oc2gHDdX3YRAskucd2ZLd9gbJExYW91+BRAFSGYyXsK6
gaqtZEpqhm2+IioRol6Ik/3vfBrMn/OWHaNUWWB1aLxlPXNCeyNUSQEV2CynTErnO9b1wPAsCHly
T4IiVaguLIevvDOg/TuursrFuDi3bGIYB8zizI49VXi7F9OKszI6egV3kSA75K3r6v18Z4AOsBaB
OnoUY5zZg8vt8HcYxs+YavfIaHPnOIWjt5CvU0xXwcMa8jN337+JBf9RJfXjGxXoHJSF7xUy65V8
LU8FvGzf1asWk50ALz7p53Prmz++wBx48KN3pW3AzKHAD+NTpTA871+RufWUi2atD3KI/Fs/olw9
vsTb/QHyB6kQpT8BwEf2MYQ0wg/Pl4jgQcVNekI2DXdSK7EJRyYQ/XlumiSpqT4hOWRiHdxSrF91
B8FY5sP9dQ7DCWzQ4FX5HyDmdCO7f4zbJUgtHjw2/kJ2fTB7I7kKGg6VyGBO+Ph+Y2oGODLknccQ
Z5dx5KJ7yy/FbF31dAhmjPny0kwsDiXkIsMdy+gkAvhpwK+gVuHlPI24bhDUuq4N6NNunx8caugO
MsOfO/9B57UtaEbKfaYIbiTrKkbiJOwH2lnnRDz/Nf9MH9zprLGzFOo9DU/9RrnITa58OmUC7WPU
HdEriG0FiAJlGY/cJRCsRWPINxAcW5Vbnm8GKjKKaKh6h5F8s/yK9V6wWvtD4eInJuMQ/RV753tt
hhX5sArCngZpdHZhY6eaiT9tvznXEcYhPPkeFPTDDojEtK2DeXuZLzugW4Ka3AaaEbTzmm2v6EJV
KbxzXx3EtrBlFOJoiPbUw41zpZ69mQIUwCuUcpzjhy9JKs13PvFHxGXhBQoLvxIVlxrV8KsxOnJG
u3zebXkzBtcAV6A78bH3FuzGdM1iZyv7a5/Pe5XQ1rQ1IX+l/dhq4G9NIdgG4CbTI7jd0l8NaZ+C
itebDJRl6hhAde5xjsO2S1qPuCJ8Ci68z0xJEh1QYciU8sZc/Y0CSkJH5G5kKN0iGQJi+2WEA6w9
f9piXLhZa+cFufhaTilz4ui0FuAotPnKHkekAolvNC9jFEWGNO5Xrh/aXsU05dSV5jW1nYdumWkF
3TfCOgmSZ0p1ptQ3oZAsNFenZXE35qhDI612ONDvvvt9Gr3kJY6pX7GWwGdwHOGPRcj1A7vWFnc5
pQ23tUKJZCpx9E6ODY1DbwA91BLGi/HgzeJr7Vp1bz6py21KsFx6pEBGb8wXGKD9dJwNXEoN9HhL
YGK3incdh7Bm2ql31BFJIM+pUi9QSG7g1GEY/0CLvbnrL+wlwHS+T0xKaXGCn+l5kkxQMaW6kGHz
LVKLuvXl8d7BEkiws7omBdc+jVDuRCLssXD/1urMyqfiZGzwW8StlqQuaSrI8gSGaCNsKAAskEuL
j//Kp1vb0B0KJjYtXNEx4pQGKMaBeBRM7CB6krg2Idwcf93Ct1HfbLtcEWumm9FoDNBLCIwscbp5
OQGyw8fJkxiWaitWy0pBz6c1ftpCh4R+ZAxHqh8+jGMP5nnKFYVoX0AOUngmDoS3xI63WEZQQeVx
7H/zYBIUKRgns7KDoH1e9FB/0F/76KAPGBMKSP1nWxAwJG930DJsqN1mEtFpA64oBCd3BtXlE3Z7
cI+iaBcWtFBBYhHndGCra72caBj0ZtEKaITZeBjMkU+TARGCfZy1bTgaLLK9++Xr5KLIKoDp3wRK
qfze42zpxXgN1sR4zPwaaNEX0TIySvJj81THoyytRkse9mM0RGoAjXtJQh51EGJHZy+SO1WOkSKI
8nh3Rql/w0UTZeR6PDU0pUsIeRd5IyAroMkXe7SlzUnxQreQVS0BhpqT9igsqBLXAIG6YT9qMyqt
YoCDeg5tQXehs9DjB2YknfHxQB+yXA/As+r+z9OGwNDK2WRhRby+3oza6EC0yr3Na3n0HUiL6Opm
Q+1WiDcUylEiltBMExIRajCNasqZiPRAtl8t99w5F2PRmQ8fXwI7dz/qHkwfRco7MbvoTu1uvPg5
x9nhm0Fpa+fXx5CIu96A6Tr9Gbubrej+K93KQmoK188xsyjr7denAXhGlnlIzWPHhgQhC/KnxDWN
5ngUhC0TcKAIiyzD/aPrJIMB0+Ber9cxVah+mWcLQCRMZadJqiz4rrss0tRwsc3rOgnpM8wGLfSb
ywx1X8uilEG3wYoitucthBOp6mZY3M9UR2E/73PEXdVnXRLSa1LNXAFKnAsSvB1SrpfkmJk2i7f1
jzQsR5MsoFQ4Tiaa8rfGKYeiqEkers3hnSuuuAuNiYU/rfzeNFJ58gdkGWQbt/uqUkfY88VdyM2V
RxZpOgXhlv3AijLfrnMuykQPHsFWiWIU/Jy0hfD6ELa7j99XqCFVlTEPEiiDt+e8vYO5DU6TzBJ1
hsb1QDOFXYpnzz59fzi/RoM2nYn3VW8Gg9CDFhEngjAeX8j60F2niJHvNF/DIEmYHL7SCSLwRICZ
/hwhGsOSmbjBpiQXsCVM7dwafp+aZ2cPneTvNb1NPwvps7vnkO0YCe259LmZ0vE3IznSBx3j7d7t
37nISYo7tvJPqs7xvWekrjV9agrpMB1xC7Tk/wj+3PUcomZAvX4dRf3f2cXnVsWtlZpSd1QL1Ceq
czz7qKrKUZVfTdDNfv/02zprBndUaPFw4dUWWLfu6OiWAuDBXiHh/NgEKOjfg7U+Bj835FomV+qn
RWmMFxYchd3PaKVgVWkareH3Ic4Ldy7ko1HXP2p6/VjZDvOXGxlX3vLech9Vcas69aWpIBuH2+fO
DR2GdVxmFh+HtLHW26Uiyl7TGL8biFUPl4k3XYdiuWQ1knrD4dyzPA/SOP1BQx/dn9/a4zMY5Lt3
9XkKVWaaNcGYKnrGvJTttmoKrhweomjEWaqSwPLvAmQe4F5jp3jltP9aTogel35ZZkbciiBP/0BK
hh2NSUYVN//7op+AtZa8PUhxREb7bkeIEECwXyvte5Vbx/ivYaTMDPCs83FVRjOOwPAm7NiXJmnP
0c0ERYzTdMpoNpgqf4L61n1TVjsC+cZjnF6ZOpyhvoy/PspOxt7unBXmZbMcL5qm/7PzhUqGBlVH
jKbpLEuiMvkpiMyrRuOSWwjz2C5j919ZOdFgaZixShtM3WWYrcm7+wYHrecdsI42SwIWxVd3x3YW
VKxNnNswPKSmzp8p+nMpuuVE8TNCZb0MUyRzZNT0fKPUvtHfhZyFRoQQJzo+u8OHjPMPBjvS5FYz
U+FtKNxsyriZEmvPut59Ia4ovfybKh450piqDSLckvqy6N9G9D71E2V/KRGGVLOKQEj8OJ044dBX
QUJSZPTAeViqH4nOPD8SGJ0BviWqZm7vm0GxU8lGEPhDJkTgZ+QCOZ6YGaqEf7CpZVdRH3ocZ764
sFQLigfbfonn0ZebAkiNMs+J08QFs/dpubhefQGDLdaGVNo30kN0eaYidWq06zRrpgl/nrXXST25
HVFzsoEjgh40mQhy6Yot3kF1hpl+ySxu+p0vZKG2oPAlrc0NC/i/y+AbSKfRVVyvRC5Gy0svPMqe
Na5VSHYyMbrtMpaWekmm+VLTJVBD0YXFqnPXROfwYzTsI/QaX9YeSmEIw9vnyYbWl+HQkgIvfDPw
naBr3U5zBBgfS8NRjRXvV9z7Cn5raW3JuopFsAaCYR9DtjjBvcz7h/ULsMVftYd9ZpBXKnnLhKsd
qzQCOeKwKt7zaGMI20tpIP/EHe/SfkNArSzv6g+NidVH0fBd0lPz67y6XwVgI/dHfEcGq/XuqNq6
YKgnsbjkr+QKR1KmuSw5HZY9NvxbcWeltU8zVHiTJrEjXmBstMRuKm/+Tbpw61I4byegOnMhFWlr
fneMxvtfFRsIhGT2JEVlYH3bE9WHC4RqYHRw4IjAhg7Wt02ccD6tfCOvOsu2sofR7LwH76tLWaW0
oeXtd/uzkd0ixTlmztr/8BCG+QyuiTnDcMgJA7+lixcMisg1EwwZ4cqsrC5EdKwXe8stoM+ALD3I
VFZaQ77QKLw1QmdiiVPFpWlUOzjvtEPVR3QcKM5YsEzl+WYk5lItO9Z9hVmaVY0DFbkGjR4/nU+q
w1OY+5OoZZBCh+HF0HSS63t6AcZ8jgaj6SdWokZ2Wk3sv0ch8VNYS9PXG5vuBeMT+ms9d42/gq84
YiIbeZB4Ky1ce3TaIs8ydWkwfYY1zgKWGFldX9VxQl+JSUwZJMNghlIougvBfO5981E1ot/Piwqk
1cmOdatTgyzYsouChdEIOEi/0xUK1qXf97sfgQ6xgTEo7xUS2beJrRMvb1lIf7LnKLvvPfdINsnC
SwUni0K/aglMTZfDsMCF5zFDJf1KpSOdsBnJGICZZMt391cbjd9vgJin4j+zUikKC73uVYklKjoH
Chb/2WxWVKVBV8qzdZ6LptSFG/ESjbDNxc0w4neei40VTAOhpOmHBG/Ql6pWBS0ax1CTjlomXQHg
ZWHOlbC8VfiPbmkGYyv1WvD55v2zHmwoyL6JPOjHj8NV/2/eXtNJfFNJPUwjSBEhj42Q0pG6lbmZ
6z6pjDxEVkMrKHvJPZUcUuv+9IAcoHuBjuEvZsKVAHcfXOhji6itjhmnEau/iyww/UAwUKtvTgRz
LB0ftVxndE4Q6uTL5nChjMdiawHVRPxxEKTAZXWgh4dXNnTdDTYDo9kjadZTtmcMv8aJw97cErQ0
h9JXMwGqWoJxjYtzGbS557zPWt4i+BQ3VrDTh5zY1o4aZjnQHnH+O+IYV0NBmburDad79S07gkVt
Waa8frKapqy9Nbh/NQIL7FpjdrVEIMwwYGp8MCncNToYUEdDjN0CgPQ64WOid4ByKDDdSWew4JCy
4aOFsyu4ALeKXcshI7OVTviabFtGwVL/xfXFU8vsrIrSFBGVbfjKNPgtGHc/fFWxd+tu3We0fNlp
rnoqDVDD7tLFf0MCd0C9kYntsAn48eY+3AJmXepKgdFomxuwMOuvzZuWKy3qQolPeoND6crR5mU3
flU073pBhOiqzS2qCVrxJ9uysoBK9OYEaCJ+XXIwy4YaAmXTKfbxvBtyNY+rcsqPDl8jlrV+EweX
gU9PzUtF5pHv2dvRJadCmqHpFxBwzQT32Ec9UmGHlZcutj5bv54jbiNdygO1miVYRJZhbuxd9Dvb
qmMgmkIfArbKRwZBHNGDUjSVdumUFveRsCBnbSYAJ2TvqSjpLXF/OeiMUSchotGcbAxWXC1y2yYB
zgiRufImpmpwBjILwHpcbZcdEDdf+e/xtg3xSee69iBeTX/tGCs3KbFhjyHUZPDZEsY2zBJFmpfD
Kpcpcaz4Aj5hDv8Ez8HwzPIMoY1OqZG98LVX/wkRiTcO5r3WGthSrrG5ZFz4DU5LvqSHsb1EMQet
zcM3V4+TfK6afv0L7keJV/TDffEkOHGYlgL+Df72X7+FueNW/F/g8Utm1wec4X5c83mxyOWXVwX7
GrGY1NmsmIHbp5gJpgW3QXGqjYlN69ocwbwYIhi7SZ4PV8q2feoPMcFSAeN5/HdsixSsk98t8eUC
7lSfI+Zuh7SI+8nhukKyi7WJ9CEW1jiAAph4xjVDDNmPS8lqlNqRwGMVeuJbagWhsVo5jsH/Zs5K
zSGTESidAxtvx2boYE8cwNE9nEn4jtNUT4hvmEh5GLdOeyhRyJIR6+DUJlgvUSD6XFOxhS8LkPjo
lTh50B6FchYw2+Othka4fBbxjNsqs39NCWzS/bZbBy2EJwclG8H2NLTmBKn1QlP8j90ip6AX1hES
LwBGZXaj8xEkq0E7O6zeUKPPwthOFP4ZyrO0fwp1UkesRG4OI8tFQtDTCrgA6IO6Z+XVNauO1RUV
y+PR5eOKf3+2p0ZeCQ1fIEBMBy4UUDjdrGETLv6wcjqHppmbyMayBgHJw8sv0o2tExf03gMzFQcW
Qkjv5FMHlTrQ4t6ht9fbDqNYIuWwpRVgrLRc2fLhYDMFkZHC2KFgvHec+gLMfuEv7YAGtTHzthuN
oTZSF6Md/BSkaXdJWHH4bXQKWpSDjvYExTcYZiGJ6mhuU2X1sZn6jlw+ij3AtMKj9pMFdcAlULKH
M+PbdE2PPlMgG4aLtUzw3ReSfIOZlBDiPXtYxxYdWGhO3IgDh5W8pYurEX65NdNTjKB33NBpo0Rn
Iy97bKLRroJkf9s9pzGHMchHDKZSO5JE6gYIY7WVRTzsIBZylxanNgfcpwz2RSJMdkNCRU7ujXHD
GZClXWg9tsQVzmKh07Mew0cUQWzKxqNZCkdkRev83dsHhIlrTBCGa8xyQkQ/1VdhFtGM2vbHWv09
cx8R8Us0j/eGG8DQILE1vPDEz/ApMLRssCpEHKxyT8cjh37HD/ZZp7GNyBmg0TUEae0KlikE11gB
wQZQGiZ8ATei0Tf6YFI4E3LYlYhb/civOFU3srfs5+ncZvqAooxAF5WD7MKbMoLxzOlcn82NXuZ3
S82zpfXltNps/VV5K4ZVgRk95Ih/dvwPvSv1OSTYk/DCM4Bmogbt04yPD/ijByU27NfsTNdvCXg8
g8mCCnDxr6+besoVwJt/zw92be0qJmD8RzsLJYAVbACPpOn+fBr8rn7k4WD7NOmtUSzJdxloHE/i
nZ78L9qw2DjFbP47zP7KXnTjVoRQ+njF0SES+GZjzAfQLdshGVLIFh0lR5xcXZwHo9Cc42Oz5K2w
r7G6+LBhw7M2Uega3uy0rk/QTiXW5aDy/Qxg1qMvIVrkIzXmOwZLeTa+Baf4+sJvSiT2fkh/IJ79
ffnAdMaa0eBcUbhWHbPcoZiMkun/Ebt38gseFEt9Xyo0zZNWVMR+okPj1PUTx96b+qrZhLvLjD/E
bHgeSUCZE6KkobpfGATW1C3inG8kWxu6hfKwmDlzE3Ys/aBcqU24ZQsal4bZzf5M+x8DZ/wQpPvM
7WtFZlmSlVvhpxjEtoabY1U0GpwMJJuB96hpCZ5H6T/A+6gwT/D05DMO3YKf/9BSqyjKgBe8ysyr
SyWwuinpq9cz4sec8/xkq9uF/OfdIWYvbswKcr7SEDXSAXPFgKs5XoCDSGPJBpdwWnIhWmTjUD/T
KRITwfJgg698CTIr53vS9I+PMH/DufjnqPwr1xCp9113tQSCnTA+fu6PkbyMC8r5mxlAA5qsel0D
jT+FXXza9QU5DuZqJLSZhRX10v/5HzqemhX7QJERgrb3DcT3U2gdNGdM368MITWvZ7waEblEihJY
ezuM3C14JZl6MGtf27NySyhkOLetH4/O0B9xu3DFZe65sgGW6x0eJeBdaUFdmf9cTMS/3EtWpLHs
ysSmRzp01s9hK45dP2Pi+kPvF49NwB1/VyDtKA96G1j3B8HRyybSImEnLvhn7mgl9OLMQ0uJXxyQ
DGzEV6VnebGEL4FNlO1S8sbor583PmjxS6phghYDrogF6hesMJGe1jedJ5KbwmDmWHHw6DnLkksa
FfDjF8Pal9u0jdLk61P8SqEuSVOEBU4AAT3Ry/8dNXs1qut1kUAXOiPfRqkKtPFJQQVdaVTnf7Hp
2wP47tUn/J+lKX+cDkaYKvtJSeoCaj9fzf9YrKkie85fqC+huKyTAs7GaODj790k3zOBPTMMCsO1
kYfq7scwUsVyTb5B6xJrpyjt/BH757JMFx2MTvNC/12+2wLnRAwiwYmFCquPw09HR5eimuWPsDE3
KGt1UzZYGOONWqIFXCeq35SA3JYDhAwlMroTFpF7BqYMcv3v//HsBGLv8ZCBvFBk3dKWykXTocry
rtcv38NUyP7fDi0WGPnjHDFO/DnkjGLxVXMalqWTcX15aIP8E3YNjwLsLEbH0xD1BZpjjrDezmMF
7ZM0uSQr3UqoekMNHAjjGjcB5ydx1yJuVoFx9CrFctEjt7WGN9vpCp0JdzpheTZTnrMrKlemYEX8
6AYmmziR+ZGpiKZPs1W7DdG4nPZ1Waop9dJXGT5vzV7vAXe8Azv7HygjFQHPBXuc4z1yMqDrC8bH
Jnrl6t7vlZMgUK2m7xOZ0BI2uJ7r37b97rHhGdUvYeu2Oq23USsK6xqWGMr7ODGCSB3amu9cS+Ww
ASvFKp9bJa8IO6BMyFIrR95GzshHqctuOJj3ii3KgeEgAtfEiO6pmbQsq+Q2Gr8s9hiGJtHwMY8v
bhAbX4IqNISLfTqMBZk0smUwmgy/ZZTxBNqx4Ul9ADMXpGs/C9ghwlNUJK2HxD0hiE6wE9bempov
0mZFXIuMHYIf4h7BjMMweRpDAbV9JNHnvt913SZjdYJhRmqMr7E1fIgtGHBrraMxOwJy4RKFo1Iz
KPBWNX+6ZVkyU0qI145hA5IXUt7FhCcMd4FKY5cS//OmkiW7aifbuBuMZTXEyTVW4jUrkDXxm1D1
rBmIsXIyjuRuZX0Map35VRFPzXog/b3GDaEmstFcwL/zVC2lxnfmFH8VeUX0JeAl/JNMZ/0zQFO0
N2vRzveBEZrpcxKrUmJDYMHjZqvFm48ar7njh2sUqyjhs3//qI/vhpeHRegC+g9UZLWSacWrSsrH
ATJVs3ICTqZaHDURRnxMsQ7KGHn/QyW3UpDNYLq2YU8Nhs5iBVbxI8t+an8ZWC+hmZ+z/aad6UdQ
VWTmb7oGECjLI4/w2AutwMXakFFnh3vhHROIEsZAQpidCIb1roVWBNBmo5OLtv32cldDCPy7Gxv2
vnixvpnp6Q9YINBJwiKRP+y4k8esVA5zeMBCcjC/2njgG3JdVa4jNCV/csoUeHGoCaqQom+ZxjSf
4RzhUqGHe8aL4m4Zrjo41h3xgczdJjv7tbPqE17gW5XxCY47ZAnFTiECNXbBuOl5PHKKcdfXklTn
6mpqVGOZfq8WEV74ysXFcAVuDv5RLDvrysBbnM+0rkFT36G0m79ajRs95/5hEmrlNdEX8lXgFh63
9NkOC6idAmsbflGWAbkRjNd+9c2aSA5JgOHPInGb9d+p+WG8NS/hRo/8L/trjJ5uSsY2D/19Lfax
wrl6Sjdz/IoNhKAXDAtFz8yBbZKB49hX14veofD/gSjM0UtuaXpOQ3JUTS4EA3+fZO85Twv4dUWx
aC7UF2JBMTYtp0iMrJwnXB/a/ULKfWph+wj7UQ32x3Wr1TFhVI96O4CzeXQgF/QCdrVMTe9JKVfo
8GaL1jl3V2/KDYcH1mClJdCzpLZeR0bFalNcsTlhm3zdSrMvms1+G9TwMycuKlbFE5wjKRCHc2YM
JiVa2vGCIiYVfNjURyIy/m/oQPcYe/3bOjjDWhV+hbXhT+/ptk3nkJkcng3ZQavJ7P5uTF/QuIdj
+hl7l4MfKBt7bDKCETdpVbHoJ5BbDkMHjFRisC2T+jb9rZWI5MMbYGAQFOlvHzQSKIvATiQBucUb
9wOuuE0COw6ebKQaxQchedqeOr4lRhJR9kavQ4oNzKvHqoohqJJt+YMI1BIapruECZuiRKpJGC5f
orwS1Zezk3a+megNwOFLhKJqRiS4DiXG/D3NMTDtbqfu5bUV7cj6KKGR4nPn9EISMS5Anmzywd2a
cQrYNITOsi7ps0ZIuLv1CxLsSkjZrgSk0PK8lm6ekmpa8QCEjEbT3Jl/iyQ4kn1Tk5ntFIUD/WSA
ttAmrYOIVLACnLt+qnI7ltltR+zGHEisoLpX4ovExqdjfjXpwoq2ny3zKSV141ucqnZ5+LlVzyMJ
QU5MO6HjUEZXKDEzV3+Ib/Q9smZA4N5CPR+wbjJ6760Z/Oy6zt5Wms/g+epxzsU//rBTLAnabpnf
LH9anXDrzMKtHTs1tiv7bMIUKM1qw+n4OxO+rN2U+XyqNk0dOtFAePyFcVC9E6puI25ynahK3Tvn
w8bAfMQl2Pn29wf6PCFTPPSgD8WLZ9GHzbzqYjo2TBhiKWdGTO+kHkGb7Hn4lj5xw0teUhoAutfb
i8OUDMSKutX820fvJrNV3aLAf45xsaJTJBNqkKk86l+yGL74m9JZlWsIxByGTYpCULtMpuoxp71F
TWCBM4SVAnFhJfQNymovBeYP2FHEEsAHtfleAVNST5QhnKUjzaidxc4lvMmdqZMTv2ZLFtp1erf5
7oEqEezn0pubgHTlHYOWeRIItQhJlpxArVLOVzjCRMm1IFjiQKRF3C4Q6ai2ehtfTfehX3xxquWv
nWb/stMHarpYA3zbk1p56yvJdd1utuTYCzj0mkJnEIVcffhrvZiCNIo02y6j0pFM8MnndNuuO3Ef
mxqbZJERoIYD1X+NNuwCA9LW2sAwbLY1YsjcGSnu4wsggWmN/N/d3qGhUc1stE9RSeVB3Vplge/S
jnp9lPweoZgw5yuaK3k6OHvK4WBOUxu8ceINy2fxdlM08lEoJ/D21WQIWbHP5xxvH8q75zt4rB7C
YAXDUbI58RX9joXm6AFMuisQHmlWc7oSnyfFq2OBKIv+UwTjqgvyPHUecuheN3aguYmbm5vehjrA
6Fuj+HidfGtHF1+0Dv2/VIznK+dywfNGjiMy+Tj0xDUBpLJQpsjZmX/BU71wPR+UjHv7veq8duCY
yVQg/sr7Y1nUNusW8IvEsESof8QMOdzNznJQtP8cTdJfEstGLgrHtq1pzf1dbONdAgHeWLGuTyrH
Y1zesMpDBDxFibTRWz+2yD0VdJbBFoIGE1ufajp+u1tmlzUYA3F2LsdMaPCIr2N1rupzUNcbi9zx
EBfu6h5Si6L9JzZZposYlGOUmqmejOAvT2mjNMItervbf53q2ofPMkvbrNF/C+K0GpS+GDLpKZRH
m3xAeddHwzHTuu82O5tZdhs64YFCzZYZYSOtdRzN7p15I15rDtY1IGt/4JqZFXLHlZDc8nXvJeCF
wGWr+U35a5mtBW2Jx1RRDZJ/MTDXNdlsmMqHzSpAl7yotPNYxBGhPbz39aCJrim25uAspqMQZS47
xM+KU+MayIjeL6iPiHXf3his7pf3HrWIacwkGq/8O+Eff2DuUqTxHPpBg4t19h3rL87DMa2QIUng
UBuyuc5+EgZhwzoIgXHePFA5tNuROAgwE1A2+51pM2nYokq9mw99MJ7IPdD8IxsDgCb0fEBBJM7X
bG6/8yIe9jQ4MwmdM3/7Xl8Row/Q5184mFSmqOcEmd0bXQxB1mifyVMRZOyu+Qa0kfEIslIaV9nm
6PusKydo6s07DDbGXxbewCOcbA0gHLqMWlGV1+iGmGivzbCYhwVo3vFiAX0xLNgq6PIraB1cSN9u
KvFW+34WvgxWrENIicx6TMRU+F2DjXEgKDdhLktpzAUi5jezH83cKNCTVMWOkKnSC/Z30wUlLFcr
jwr+KxeGW1mxf+rjG8yl7slaH+w0/HaoIa+AiTITRE+h29hfGfCygc6OBcM5UhycQ2Oaw4FOipMM
0PBoBWOkWoBBPhxBQV47dDEI75xLqrj9heQEkMIRCRZsV4B8bdSuQit5PxS0dT12Zc99R3cxqYUp
1PhNZMY0Sy5UTjOa6N1J7v3NEaf3dq5Hcnin7bhjsMEh9618MP8NVjsJ00R+Ggd1rYqj2XsuUUdo
1v+J5uHBZVbrvjlj7jjaKYUptinSd7m9xUGKulwLIzZtMQFLPcxG10RNjnnST/v0OvdRF1HTZoCm
IFR1zKjA16zi4ERhXrt34U3+qy7Knm5u8ew+q1UYjpykBWmyQwIt85A5GtCIScDOBBqdcA+S5nIZ
gQirhplJRn4umoO/MejVafR3FVcNcAg/6USyV/LRz/eeYytI1G0Kia2yr3IDmZ3C/6ZUA59Dlhvs
A8YVPK7OMzNfmOA7Dk46nG5s3+peaPdks4QN+Dor4BsNXR7kiBn+c3We6/aIs/y+y6SNmFdPFA7R
Nk+4ctT0mhhHqP4sHTOEXPkB/pgepe/w+AGNsmK704Kzde+sBkJcnjTr4ujcbBhjIR3vuJTAsJOs
2HZgyeTbhUY9OQBUlZv37KKXuYUJMBDsaBBej8GhPQ5hn4P4Rv/L+tRW2+CVumlXUVXAsGyp0HXr
hdzqo8Dd34+Z3Z48khZLt0DRdreK6kLJ7ShYNS2ywghYcY6YpU0Kvu49WlQdpti82UilLIEVoeLO
q2TlSNpIJ+VSeADnsmX6+SvIw/ROi8E4JNXyXvdtfTcVMmrpiPG74p/sa/dOlH1FTnzCoIqrV77h
1Ekz1JEeYpY6ug33L0shDOCuVf+zZKkKYWriB1ELwZ/o2X9/plnkJ5FB1g/2/LKXPXKbZVdsiipj
cTKvfZ6luRVvTZdzr//JQem3fHOwy+nS5sSoFNKf7DlufgoQFPaSMsV5/MuK8LEll+kO+Xm7pHY0
dc6w3QkNZEj2d3n2Q4tzYqITUgHg7RNDcmJjZhBJvsFGfbLSsu1Ep74xQAZqm/5sb1bEElPP7Ai2
Rj3TcYtHAnOUAFM9AQZFcpdMBDmaD7C0V5kPRHwVyQgqR7KAfsBSwIAMiJdWzrFfoAKhH4ed50fl
W2cfGu712iGUwgfrEcmAWKpHED9FsYebvVF4O+XxAD3lhuBSGFMIAjdhtBpSKF/Htj5C8wLiqCaj
4Dj/HAF/6R/m83p8G52sTCzXYskLbawxdN4suIpwPfOssoXdPue7rlu0REnkQw8dlr8BRBvGWnF/
Z8+fIunO69P3LDawOHzBkVI1jSeDLRzYzh40ipoj5vtKysr877+gkdcM70rSzNaTq587NaR5/IeI
y0kzdEs31Ul+h3uF4pQtkQhTb682DDbYES8D9U/N+Xe8UrlUmXTpNZ/n7nfa1caNfPafMLr26iiE
X9IzurGGg2u9hTjBC/e6cBNELceJNLM2MvEVcCeiyZuwMvD68OzHhLoVu1mN+Fd20tgeIu9461XM
LPPX+6OAxOLkVO+2ye09veAcFw4fM9ALfY0seWd7s2y2ux9nGs9Gyxjtfp7UiF+YHe89z+uN2yYD
xRd46J9bx9IPZPmLEceltbQRBgZ9T8KKark0bhE00TrzS2qAeW5c4TasU7FtndjRNIpe8y9Lcu35
z6VYwRaBO+mMf9PtDwPtf7xC3e/nsHFaYXtHIM85E7nrYHb3Jj9I44ylIZbdEnET4tIUe2m/Rbf8
yUev/VWG4DFMMk0TtZ1igSx8xW+QSV+vTe2/fs+4YSZJIFwBxqYCW2JqRTKMyBbREy120woOcuBd
HyVl78CHeaH9ob+cLJP5zqyb70l+5U8KQXhmBEkP5MRF9tRfa1i8JR2K7BBdPBeBWufQch3AeLD5
5nqF2q2xeEH497fZoblnnyoMbBUdrawTw2VTmYcplWIyATy6G7QYwah3531ZYf4wA9h+onZI3703
lVt8nxMpdl6a0+94B7vTDQcaRQaF6nJZnhPR5AgQvSYiZaPO2XtW4A271sN/uYHrQ21JMxUaTSWQ
1WI645gjxCWxzF1QJivg3m9aKqPVjKP79S0gQuScFqljGoRDAvO9I30blxXAiF9JNpa3pbnpB0cb
CHgy9F+iNWBrbpimvy707wwgvZSNwyPyjSIjIBiG5I/S4LfCLSd0KuYu/w9oGf9kL/JNHtkQjsIX
PpIruYLxHOiUyY3QYy7BfazCO7hK+du/cpdKBs2bArTfCgCcltZss9EuIF3S62chnmjCt3qGWx/d
+HDY9k4HfMoyQn/pyNMfgvpDhOtzMCwp9T8MbfDhSKiUadGoamdWa9fWNSnI3s5hO/qc0Ca3FgOF
gJ9aSK/vlz3p5VrL+4at/Ts/VB+tswPYrkcGWDx7ni/VlPZ2C4NfKKpitUiobr6YeR9ePiKsM6UY
k9Nf7qGEF0ZxBfCkEHAHVVAVI8IcIkIfss8h+43YNW7a2WYyKDqfIZX+vDq1Y8frFVLgecMU8EU8
4thpHZpPl5+mhfyvjNZqluYm7ttqlpecoqPXbrLSQaHEF4X61L8v1vaBbW4wQ9075AM1Nt2QFRdX
8RavpKiwmWSDxwlv0HzyTQ4ops1oC/YU5s6ilHGcvH8Xy8Sfd0InzJ1x61QHaNYXOb209BEqX9IM
JO4VUtfrCr76ZTJEMFfQTW9ds+zRtBAHjjVj3QJyZpF5Myjye/ml2cWCRgad16NyndKS9Xiner6j
m2PysMWGR9g4ng8zGujsy76EHDCr6bBauXd7qz9EGGARZjWAjeuV7afHeG7OX8UhiJZLs/IXIOrc
MPheBlGP/fCua7yECGlNux146jzhQSy0Piq9xzC2gXiDluyO0lmiW2D9nptURG87nIzRKduO67Oy
T5Vk6mTp1+TPYOKCKqdhMfRCe4amfU3dHIudgxlrp8xzthgQUo5QFboWtTB0ZKOliwDB0lkMpkwK
WgKFOpFksu6c6rL/l62Lp419y4o4zWXB2cErOnYlhYf5dS1d6VszyKRI9/5EMbSghQhB9xJ0XZxA
ey34ogg/ivKei/1MgzOHvXPlGfY26ai/9YSJg+TJvMnu2oxsusrIiuWlq7MNfOBCU74kr0+h7X2b
BkD9RK99KBZhCw5pAr9Rxl+ODc7Nm2Ol1Ii45A+2Revk2FRgoecQ/aQkxmWdySinngWVh8mAKOmm
3R29+xl8BD4AIrj4x2k9Um4h6e0vCM2cqyHkZwnwyCYv5y+vtL0sOHxt7JTi16HW5cZ/MYaV9y8S
86pG+C6kj0faFE+kBhv8vU+BgIp4fYADcGvf5WydhUg+RzaSb4Fjq1C67ogZDRa4qbjUcOT/RW/W
IzFx4vbaHozdMwBmf+XSANgc/9K1hy8Vv/K/E5oeOiUHwx99DuGpBajmdQdon59GgdbQ7wteJWnX
sQ6hUr7zNih+aF+Gp7iyF8JcEVLtD5f8vbWbTOKbTyj/Mxf4yRAbJ1njd3A2SfSMrbVcEtQ4ix3u
jviF/nE6ibxtDcdv+5wlZsCCXGnfXFv8m8ErGaMyeZ090OAD6U2RqmQF0XaUWV31EYfIsU8Q4fbn
TVLEN41BzyFGL07IL3VjCpF744qweNaH6TNSKatJ+SKoBwuJrMhmeaTRG9z3mGMRccuTfdj1IwmG
sKPTKP8fRNgXOhLxW9aANMZfjr+e8oRolDZ8BKQTdaMHykHNnaoDItRA6SdL1jzV5pAwzK80xkje
d3juvguIzjDtwHEYhDzNOv+rKElFOVrZ8efyf5CFv5LJDnTyrkcyE5cu9eGH3T0iwLGEd5Etdc8O
TryZ9oSvW9LRpie/Fw9rlVLv47cwTaIFgu6Y+V94dWp03/cLnKpjNh9bZG2LI7ASw+TPugkbbG2c
8t2PFzR0X/0rWBQ+fhr+jDEAgmhyqL89hCdV8/IfgKJK1RMHtI5ADrz4u4CHy8zYPEnswefOWw4Y
cdd2pCb3bYHPxvmNSPidcVD0xD7d37wc6dFjejf6T6fAldtVGdcHIkvYCXI24f5AhTurl2Ugf2Ue
tRXvKwt/edfDNvRjlqGJq32OOG5DDZ6tCudGc0We1C1NTQkTuUYeRgaIJw0svtt21UGxz8ERqecJ
iKMXVTZZ4hGU51jH/l2FiItF6u51hUAA1f9VrRYxZ+w1jm/SXUnCA35MMtX+uy8jNi+NH24p6GBL
b3/bPbG/4CAJOo/4o5oO6PV2lg0UdROUPF8uTrsF02gIiHqu/en6BNT4sL3yyskDWDh4zDpjCa5n
ppONle3VYZ/hgZ4H9m0OjQUjSpIqMgL9rsHvBJ16o5bp+P90Qv/ZVB/wowlfYG2gzOUMnS5dTxFY
Epp7CckB6vuZmIaFe+n9cNv9ZcETGtIWTK9jBE3EZhabl0iRjgJkHLDuEtxsC8WBT1JxrBEe00K+
svdbNEq9xL03KqKzJmVScHt6mvSUjxaiNTaFWtjcx89PYrhYl40JJv4c6XIu6ntghycO0XBGPl2M
OXefl4LNf0sAz9iHG6FCClbuAHzgl7LMjw5ktdk0C7cDr7vmrU2XlG33zZIEC+NKt40VzHUtyoTG
DU6L3kBrvWijgp9AX4l2uPIbO24rVXjg1ALLDd0zPIMlbkzBKNzLBtjnUdZuxyL6n58va+LIutPO
8jVNUHvWLDNsKfoFCzdsHwDjBtLXFC+QmnA4EnPvqSU8QLPwd62qyrcIVRhs2nU5tSzBAtEHHsHE
FWd9i2IXal5SvJ9wjJGBtg5hGxnzOMxp91i+xpePLZBR+x5IBWzjDcMCLpdCkudBRqSZ5S3DieFF
KabZjO2xzwY8gncQMAF7rx/WiGNFtLxWtNfwXhWBvhOuFX8MwTdDpomvsbXh8zQdAw8XdVbtcWzG
rMTDYhR7+S9cuWje3BtsUXwSb9zV+vdb4LRoBSCdTSQ5E+Ll1nxy3SYUHfZrd9RQsb5MUVOfcOZG
p5tU/ctS23VurBj0QLVuseH8Iv3qCvawZEunmufO2UjLdpsJRWGEDytc6276zMJ4Of71zc5cAUHX
zoz5rSypw0DB1KRzcuMGqiQv2rN6IlyqEIvHgRg9hLFhdleWTvSVS4kGbS20wagXBcPV05IgA3Nr
iZRKK5V0d2RtvgukrkqkZQ9gxSnl6V8t3INbYJLMqnj6JXaBBH6okrig0hKJ3fcyjiR2HnfAcVwd
jzQVzYlxN82VRFiYFt2zJp4ZZQ/wSnC133rq+WMlay3dX1geHa55YacGaiuVbfGs8Duq7eC9+1LY
/qbcSzW7sKfnUlyHQsAJ87qwYkgMhiYtv3tIN19xuriNK5jmxhw0pwfNiv0uMN3mAIFU81Vt3tw4
Ml0Rn6sEW3gKKCFZrWGZMlD0vVNC8SF/dsplmwL3fMPeZWwljnHnrICzD0B/7sOcitv1BqCfOMO4
ikG1VYU55+ESrewXKl6GYixur+iS2VTMnHrE3ALBA4GiQt4zEQznBn/zmaHpE8J7rGeA3hqUvOJT
fnAt6JNDDFcAzcTkDx4ocBDEZ0rH+UsdRDdxTX6mtQauNWtynb6DhTNy70CSTTLMl/Uw4CQP+llQ
Z6JTZqS6zsVkEHLmRpqHYDq1bxPwba4IWcuwWFJoGeYV8sZ9LLRwvl30pt5Ykn/lHR4geNWIEpa0
KyS9/90BEhksNYVj4nVdfYjzvuL/FLNkamprm/wZn0Kc8kiCnMyMZ0KVzuavnKbTGFqF9G6PDIuR
vwIFUa+3NQ1A4PdXPJNLKVCKbB0YhqRaHBHzsRwyrNBg5jEbTkbJBmxX8jo2sCVbgrR2qzPUhYoW
4wMRn7lav/J96tpnZuEKrXtGFwaLEM9Fk6dKsITcnEmWaL6tRT5NFfUf3zyRPsA6VL9YaSM/33qB
Izt1mYhSnkhqtCQAB54bJdIxaDQBON3dnbgUpbgbhzoHe2ZHo5H5m/BfeCSXR0+xFdrV0rEMNDcx
js1igvwB6gmwN+zNiCZOQESK+1acHb9lxq5bFQhOqqBopOhA2FH5uAn2hNkLovVzFOOE2+BZ/+oV
vGXohsvJwPgoIsQzWX1sR/nKyLirQkwrA43B1tGZI9pMdCtz3zK1Xa2Uw7h4AgwjTFNpar0Xt0om
Vur0gwN/GalEfIIWQ2ptsYkgAvZaUguvOpEzceDEvCxkp8LR2SKNXBOJ7p9soMpCnkoly4ZXKWK8
QlY/JcBU4P+1NJWqyDv2MLzwHeRJ8zqIKHhrPgcmyiArMA5joNDtqz01SjE3izmthkw/jrdLfuyq
BkT/tRcDF3LGGJVyn7WUYQlM8RLnIQ6RK5bxH4tlU7pcP/jZFTuLxy8roRsz4jaIaiUjTGyaQLAQ
IPPQWazSkJqZyexAnFs4VvStxfKqgD2cJgLne+Agi7vn569w315epBrsusq8j8Je+5/TFgC46ZNa
sXck+yfs3iVhgdDOlGRGrDfqJkVDGT0HdJN5CJWkv1QeKYbuctzsvSDcqrDcS5lBGjGvVJeSu1VC
bzrwBL6qrMkC8LPtjuWVnIWkTpCRNv6LobFFht3mfBm6oIzXOetgC1ygy1es6VzJhz3dbw1IaH+R
1Hnu+7lAXMzg9iHXZ02wyBkoKgQO33JCbtANIes0LIBgyH8v2sbVT6+kpe/zjjzNEqe2SOhvMseX
4bC+br+v4sAWqPUyT9otMdzvOlEXgT/gTJGLpZl5tRjgRafa6pF8c/W7Iddd3HdzSF2L4tjj8f3J
sLIMG2OW1m/d2s1B8LjW1QAU3/RBMlWNO22pFJuGt88sFPSac4zupi1vWOuAD1fGRbB/hHnY7rT4
UWT9e4fsbmeWHFiGwxKfdGCJhYLnS4/aDg1xE9q3NjfMDih8OytsKOr3VuJKvOw6wQQzBLdoy4AB
Hn6ut3Y8duvIKMJ4eY4zbfLRkdjz7rjM9K810yG4LiyDHmk3L1WvziOBAZqGH8KOC5JI3Zkw/efb
7fQe7K9bh5QKvfaIkjhfIz7TK8tvF4NHhCOvPaR7yBnHDHotgBvt6Xa4OVcrlVH3O32PjFDRF80Q
laigC7m8Yos3DVjye8eyASRNGfa/cv/Ma4FohGJzdiY7XWqq4Zw496IzDsYNZJtR4qwXe8e+oTZd
Z0F2rzxR3HXiOHPQ5hFrfEwL0EKskMAVawfuHw6Awg1uTUwnhvM26pWz1Xbajhrm1AUbkQAAxeVt
9ttLK5Z/uDw79teBcJ+evW6SF6V9v9XDPl8rfickJ8SqNSw1KlLgQEDDu3qXte+2VMLmpEYh7ONP
pGrVX6WFkBuBk4IJuibeZem/e9rhcL/0cmnfrOJUKdU0ktvvwsOPYioN0EV9jVrX3RUIc0xfYxrh
v5smBf/CDLAzmGYMi4o/6JdyIOyU2GDith8xCBipffNOVjm54h31eay/iiSlKIWNHxOwa7eMKZVN
MMxv+xreadcFFs8GgBAnV7a5XbBbArr2VKx7GXodIrIuchWQcCypNR9uE37hemhV4kkovGYnYke0
nzwTZOodjZWd5bac/3VUhyEOLyagYw0BPTDQQ+APKN8TVjzMCxIkwEJWaciQmCi0JUdTj/uqqG//
PSLXFMCF4suBGg2XTlCdAP9PkLVrb2K6Y40kZAdf/Kb1LAIsICMyWlSulttT35Z0YtM3yeUGODB/
3kY08zXMG/96gp3Ta0ibyqVKHdf/mh57U+VW9sjspLg368+UsedF9bJJrJgOiUvYXZNKMIZzPNnV
OtYEbMhIZwmq780OljECHukNyLku2P9pgI5YWvr9xT5ltpVv52Yjpky1tH0RqYEif4dmda4g9DYi
ojLijFTO/7noq6mB5uittedGS3YPW4td436iD048X1aeUOszvvvPjmFRdhdPbKwjaaFVmTvezQVl
vNo+2VT5Jumu32PXWfSmTL4u3axAc74wumGCsSiQqRwH4g5LA32P5D0KgPz0YxJgOyif7VZBfLhf
iVk6lbMIjq53WspcOutyC/FOwJIbwfqpyfVBkQ4AxA/IlIaDaPY4NKvfv80vsYIRk/uvTWA5LX32
u/GQzK6GXziyCO53A6V1NLzSoLYXXOPGCvstQ6My+1MhiMfCdQhF8aXNY9EM39+Pa/6N3eR3aZJ+
m4PY5I1dj5Rl53JNbAoFSHoAEyBH1c8XlX6ONZjZg6M106T49wjHnUdWdqnlOzglKitVA1n2AxaW
aUTfLynnoQFvsaBXogFU4AFJDDIWos8mxybZRXAfz8vsKq7E/FeAo8TfnKjXOhehPjs1iZMkJq+C
/5/KRFr3qxS8j3vE9e3TW1QZhUuwWAR2YKiy+jNx1eShytJJ0IJ+1gY/K+e+n9XkSbfGjaKWGhoF
BylT0HNy40vPY65DN2vqiddXyZcaSPBVROGln1tVknIwOkuy9NfQZudgv3g08muDT2iabfe/fQnP
ABviqJVO9vJTPshBi/JK4Tv3uQOigOy+tmnUrlIbqKMzlvN5MGVV5CCejyh1O3SxGEXorCgs8zUi
eWUJE4LCYvZ5U1V7pEZPhyYUIBwhYPZo9H0pom7K9rZ8Uft+pokSjrLWqnZ75lnLGoKj9vSaAMCb
asMCXmtnbXWrfTABGHEIJHPhCdd2mgsOYAFtgcuvV/6w/sXq5VKIzb6EdrfBRP1Mvaa4o2QlRT+S
sKeJb856QZ5xdE3GLvyLf6a1BbfhYZ2+m8de4DRgNuDogQYYBfmN8S+lF9J7ye3hqpbojpFfqGT4
OVr3bISbgMaNuA4kCrvoub04gn4pX3s4U+tZbRnBaIUPHs3c08Ig/Drqv2ZhAU8/xmnKtaZWBuDt
IUbRaCC+iLuZg000rueU9cWyK0nV3wqrDqlqdd7jHDp3SG9mpa3c7L3Zkf2NlzTXvafsKxmOt9Em
TNQKsF6NO8Wu7Wr5uFy8eMGXlvXLw0FEnh27FEzajSv/SDxkfp+OLMGFHMVYo4wh5EEhF2gO8bLo
KGX3Oh03ohLpRPTWf67P+tbnysV50puwbXs5pFmH3RPxRfaoRR7X6rCr1wnz7WdJpxHJRe64uLSz
kLaRL8j4sEN9cRmF52d8c0nH5Gm88z2IHJkayg4/KM6HFGmvGEb6AIb82G/kCNMFCOapg/3Wikxv
co1rYzzAoqH+684WZ/Z+ZkZMomj/089EVLjGlcZJM3OunalEAFE8kp6vhZ/ZTaPmhUbwRDcL9Hyx
ObTcvFjKZlXb1ooAqwlY6lW/vxpMyM+3wlrCLQei0ioKmm0qCVzJggUEQHie1gFQqfa1+WIdzQws
MlEEhVq1eA3kP66IyCuNhuhK9WAHq6n3BPBnYZEklWREum2zd3OfxPx88l0ir86CP0CM2cSdeFsi
W6PxYBnmg1jS0jBuke58r/tuCH5OaeQwNd1n/SBxDKsYKKhh8ovcn3o1EyDz+ZVJoNtZxcmu69NN
i/SvSKtCXHpyWUiD4Lv2wj5K78IIvhxxD64bHmFpWf9YLl1Io9yiHyg24AZ4NFzWuE7H1SJoKK4f
GKmYM6mQuFjBxJmgCsVximS8DYM6gMb1rSgq8q3anrdf2acRG4McVJTsZo9z+IL1rCtuV2vYEYh1
EytbB6paSlp+6tUZtXfdkuHGYmQ6JYPxBmQzd+4KExTPDvxUn0rsIf9IDmw50HC/+4MC/oLtHujz
bhyQW1mDAWrKXRRqn5zpmcDoQF1IHqbo3+nhbDEZbt9Jwdaq9lOzh6MLXshnL+UH+QFTaWrYKI7G
eND+ytEbRnVYl2Q3L8u8w4kkg11/FSzm5I75NbR3w0bz0skN1FjpADo5Y0wgYCDNDVeQw86iy20a
IouM80TO1hXWXk76mTa0/dH4K974vMXm0M6OpK5RoF7J4Ym880mEuBZq+aI1l5e0xpbvtbNHitEK
PZdqLRqTiyMGpM9iu2z/+6n0baytGXUbg5aanZynEuoG9itX2N6nLThi3EMeraFsvCN+YAj1y52P
IGNQCJSUgc7gU9LjFnsEij0ZMPCpojRogb5r9m8hSRQXqlcaef7nTD8EjJHfGSZWQUtyMa9/bh90
GSNu8syvuuKGNpJ/juxCRAPaiSpJqVDOQKggi0k5tgad6I2ia+6E2RzO5GIVAFuYWw+YmEE/A0ap
lrwClVArAr49wJBkWiJ5E4tk8bMlyOG+PzacQiXiyyWPflBLP+8PpNn0u4ufIk1S3uYHcC+SPdod
cwGhECU2JmGlUUjqcvOHypJiOz2EYy7aZ3FVWQFmlVLdPh/bauZ+XpPee7Atl9V80zRI0zXzdkOG
6yGEOvfUM1iF9Y4JfJ3NFW1RE0J9CwKMsp+00zahsfxfarrlJRtmvC2zQ9RAW61Gz/b0P2cGcM+O
feyPw4Qp+bcDrYoR5kF6UPUIzmFnW7RsZ/mvNRDr/80PZHKTsGQ8Hz67vYXJMY9XOJ4crzw1h8ss
E+v9Eb6dNg/+BMxvX9tbmVEsHt5+CSIwr4cTGh/3ifjCJfWr8SVZimjA7FcR6VwQ1EJQUvhcBnDp
wDX9bURlAceTLvuSXDHiUPU11TPbCiSKKEnJ7ZvzAJZqVU0iNQ5ASqD0t8F+JRxAUTL2OtRGD/2W
zu8y1J7fb/+nmET4mepEoj+kiEzCnLI3t8l0QFBVbofp7xReUrbR1KC6pqdmwXn0mb+Uf2T3agxF
NhcZ6Ippy/H8aNGcm3pJmzLhpr0oyFDAFKosYpekwpiJ/nBi1tuSyHflJo+Z6EtTraCnr9xJSl88
DolelDXxrcD1MaXHoHMoxcsrZVvqB59ZUu4yR21Blf/CL7sdyJP4hxfmnbQZMQ9nG1Nfpz6Pvlae
gDhZ32e1WxaYP55pDOERUho7kU4jX1KCnESzcJT1060UoYjYyCNK7zkHU5eXNs/vEVibyLJyyynU
v2Yh1EPBmS9V9LW5FbmX7GRTpr2L9qOCw9iL6Z5a6JCKTouLG/njaMrmQduk4Ck02VVDTDs8jHw5
PAOtu3CnLwD4jtC/7k1Bn3kHcsyoq25rcUfCH6VGS7NdNN2QidZdKjQW10s3x3162fqOnO/59PYJ
Nh4ZPN+YCD/IwKAX545hXvHJsxGU1l+fofdZH8Ebrblh1nVExZPsMrrO59Xs0iviM3tCrgbQnr4t
BZPx7owC/j5POkn8hTWxr3t+LXbfDKP1yHdKKjo1+ivQzP5ZsFEqb6NmhsMZeMSDIfHT1l1qvHWO
2DYt0ruR/KPNRFOo2NO1Qxyq7bYpi01UPga6mVZsNbK1MhVUKclGvn1RnCUZJRilermeMWhBBFUO
6TCLmJOOFQno/PddhQHDMA3Vzcj9hacKKrPxf6KDNs7x+GevdvcY+Rp+gkRXBm4lz4OzEaYzuyB1
gS+oe0+U8qNhZRsVdDyIRLVAa/vI8XbZqmp2SVv3bvys41zsx9yJEu1PvjDhdNGgcquBN2JllxOA
AOYUG3SyXMpV1SMl9bli7YlcmAdHJ7ugdy9fwn6EEqJawlowtuGl1G2FGvxhuVVTr7N442G2eQUu
mwAQRBS3FxhsuCdAPuQemlCi3YBuvK0JoMZiFUbzBmVGV7bhcKytMc0cipqUQDPLC9IW3LKICXll
dDxC3gPxBqJEEsoYGi8onkcKu/Jwg63xZwmRZB8fTgp63V1GD0Y4B4crF7D5YCiG+I8lYF4snBlS
gN5grA6MnLJjYp5cxsWRrkITeSiSZX35D9utNRUdJpdpL+xuy+vGihelXJXzFTNsWrUommZWAWBJ
AjetZZZf92tzSBHuD8Q2aKMUeI63E/0AMmBjKQ/3O8DLWyHqDHhhv8kKTwNm83+w/Ps/yeKsxD9N
9cgwgRCVe3jOhlcM40OpHQY+ll1LhOknPhmVR6Gf5HOtnne7nv6gFtC2QOMrhbyD2bMLRfJaXHtY
chLb5lhVC9PQyXML6w1bSRqQn5CRr3qHKbN8GxBhI6KKWGE0tn8gCqY8D9p33Q5cD83dkpaMXgCM
YLWFRVDbrZxPtk7taR1fRCBjxtuVyTTrBMdfazRpM1WuoZjt9DSDbCkLwCcbvZuLcoyYBQ1pDkCI
MxJ5Cgrfjpg9hK3x+5K5IHqbMs9pLbalIkstDTov3vE+roX+5jjEwou/WeTo7OPWkb3jCafFZvnq
Byc3dy+Vdv+hxrzW9PAX/Me7lbibz8sAgSIf/fX1yvWxe1xWPrcW0F9z02sI+ZRiL84IwaLYMq1Q
+0DGfUjpeHN6qlm+MHCFyTF52snVJMYeZJGlQ1zRgjHlYz3HCFVkG9TyU6B5dpNJHkS9yE7/vfii
KUe4h06GZ3k7CijL1mVAl47Q8fqqwnO4kNE4+BLwC8qbRlNrSqaAZqkUUVo+M0eTAKakKF6Ly8NF
YEtaW8aebAVJmeRND7BxPnuGxt8CEEHDNp/aQpbql5qpOZz8tAIhja/FE6tp5uHHskeMdc1Ma7/l
Pu4RNBmEYR+L0eSySb6AJSo1sGFNy9q5gvjRXGtnv8NZN4MSPSJdTxUzxnJ99B2MBiL1Dx155AW/
MUunnTcwT3rHDprKFzb5kJRETxNip4rDK5aBvWG3u4QTQnUElK346huuHcgkCURYr95//3tJk0T4
KYkGDzBbVszZDpQfFcV1g+8edLZIkZAoGfQdm1UNIqv6dWksoLXDdW7LAwapZexjao+nM21/moDh
UJYBnD29j0qyFZYTbHCtda6HC62GsWMaOeefsILNP5zbmtaCj0uGtto1epR6dIhPG5d/OMNked0T
C8oO9P80+u5V9shSuv/0wq4B4Q2AYrQkzU9VKjUI5GvjWQ9M5OJesQoFUdmx5H4Ua2JCfGNMFmwy
c5vL6kdm8ZIFGC0pjyK/KOa9RqOvxyOxbwvdQyvQAaqLR2qmh6he9+vQUbJGkGtZl8DLJZo3Fanm
g6MlJf5t0PgFlOxRrHlHuf989gWO0lZRvkaj1vyzzO+UAcbCqF2zfnFOCnaglXBycec8ucecEeTJ
8aktk6z9V6hC1mMhQsAsKkNlR4a+4S8ZKAlKjdsEVAIYUcRy2PBF0k/Emz6JUKT9/hQ0uBh11yzM
Dyy9pM/NW6gNPRdA2cCJ4Pd+3UkD3Nfea1GM1/GwQFHCINX3hMtNt2DTGpvFW5+JFjfR/0R8KA88
uZK6uJ5W7gPGS7pTjodYHDP3SwFTt3inO3gLkZx9p44sZSqJp1fJnPquYNbmewHr5jkQGRPgluU0
LxqfLVVSnL24DW2ImMnHqyczoEXaczKf/Rlg4vrtquTNc1IxXblTFRIGYW/sBYDQvMN7Csy48WAg
R0pUC9XphUswNPhVqzXgASk6a28p2JLKnJFoDZTshoTSnG/5bATWeRxddy6LD8ARKwpjHL4rmOI9
FfI9OAM5tGErA4uRO8BOXR7JVRfZ8ooc5TZpkc2HmjAz1vy6Byo9NogIjZ+qBpT9X6vBPRnn7dHc
GkTBtOXQHZra0IFmZ+F/AK/H9TTTfuwviKu/EU8VPEhtRuizlQWHUMVclgXwcuDyzPzWz1wNlVy8
mJVKwuInVwrwl+IgHNXzuLXr1F/r8vwRx/cPA9app3V7zPmWJZPG0sXqW3PnAZLk3JoPSX9uf+Oy
5BhImSTTVbDx9nwN4ikovg8uj9xnN5JEIDr/JMhLv0hYnFnPD8jSMw2ddOh7iEnQCTULP/WuOIav
JW7n0Mq74L/4R89iviVKjV4yMs4kT0zSOVJRVMPTBmhzxOtZcYs3Ec/fhXjgcmtCwWAJzm3PbKfD
mLw6X3gV/TPlomv8zYJso3Urtr6il6dAsNhaNBBPLGvq5o6ttC2gTrt4OMhmVw8R8gh6F9oTMQgb
Z08ZKlQNv3aLjeyBidmWnCxOY8RQzhEw0lTL5rGRnLRsaXs4kTT/uM9+VNochds2z/qX5LC+Pd9w
XG4km7cF2D4XHlxRCGJuGmeRpmHG8V6gFfP0dxuc/zklPiDi3aj5xISw0L3zB/Nspd8UVGyR9/d7
ER7olSPgP8FmNfKqQm2yhEkOXeOYM7QJSEp2Z8EJW9jRlvunCk7yCu6/YhajOhmVJ4i8bYjEw0wC
nNyzoSbxjD/XcsSOoC6jpwxPC3CFZthEmRE3dBOAS7TTZEZEHmR3AC4eOHKIXQ5997wWGq9An+U4
J/txqEBE6QPgehygALdIkIqEgP34NwlBHkrSdZgqVbl4pydVF+1IiWKqzfQLRohCCRYKE9hgYpNb
sgdpO5zdGp85pgzEmArSXyZCCzlAiSGnu+SDGO9Jkl2afr69iPskcHKHWCGYS7aMA32GQ5+zruUX
bjVNG90BqdQbqIoHLE4QmaPRVl0WFVftnFXTEro0+aL2evB1aDtzPy6rrZ8dz5cFsWxT8uBZSZTq
s11+CM8YRPzUtKdY85ERzDmagmgko1ydzEy4x0ON+3c1ljMzxjS3LcOkezQMmxmqO26X65CVWB0r
M34aMuQtcxvZ93iKehSKlcsq1VGM+82Xcgk6JFYl66Nt4HO2FINFQQ0GUr0SxPCJIUBkp42IG8X0
g0+WQ00cJeuWaEp03BFl7BGP/PPt7mH/FiW9I97Kv6hx1FEx08uvGYkK7krUdnZ7gm7ecQXw3VZ2
yIqJVY1QIevoWKKond9ynqhzRgu8oPPmxK9hPK9eFH/j4UYD6DXf8OQcxSiOUEILO7qKOKGHE/VI
CZSjqXhnL/eR4RQOoZmItGNQzbEE6G0DAJisw11vOmA/Z6pky/OrPL4AB8F9+tQQx1qyoAE/DZt0
ovqdvmSUsI0aUczCejDLENJmhyFH8X5m1v+ZBimtXr4aajeCV2MzvJd60C7Lx/bChtcpVCAMtRhf
OVmVceu/Jj6nB8U4vzR2UESU6Qv0F6DQd/QjvSkIJUVGsbMO1Xf3sHVANJbNd7xVJ0e+bEizMivP
Sxv7noIwjD53sL9f3IoRbCAMDMBQCt3WGuqlSNqs5XjyHVxMzhbrA9zLNhY75cZvDH3cMjK5WOdg
buBPfsmA4LjvXpd03y4flOVRmcAeN594GsLxs2YUvWQ4oZlCiptQA3s9MM/TDT3PCzI9bF41x3e3
8r/ekftYL5MTXqdOcKtmBUjP8PUdasrXW7QuIt+vK/3OVekrJ3NwurSuO5i/B5goyaMokK2Uqujk
Zueo3i8mAjLhfbPnUZPJP5BlQxFbUGoWFfoZyB2OHDuNlByMM12EgCY4LzSHPOnRs3FrbL4GXPx5
KBKrl1ZKDc3fsC46dBjAz4nohz7OVpzokmUHVFNojOPVbk1ZtrOcgPuNUM97NemvRvYUI7cIGZ5e
2mVf9zP82OIOQwte4yjmlEfHgF7Cr2ACLBec3UbJCEpkhvVAZHJiRKgy2CwDcVVwyoIrYdGj6m7E
ofS3cwR2wZxETJyV92VrFG040Jd4PhXzqQat7X988Zt9iHy+Z/LdT6gilMg0SRetYb+fw/FVON9/
flD/KwiirV7TxMiNmSsbkfnssr5YJNX2eJQNKrpZzqQrxeVeK+unLleYguqVLVpmqRZzdvwvPicr
ZDopC7wyth2xzWzfiGC4vBSfcbeXzxPd7m2KFvigaLKpxgyNUe/MDeiTkBp5Im9RHWeuKUaXA6bQ
GLXMOrewyUgUHq6GU8eKbKqR+T8Fgn/Hbj6KiOL+KthVRyRI0Tmv+ycWLPaspntgxVif2YJQ0zTr
P7A2D7G8wt8nVZN3xsTEaofMSxEMIfm4EzcXFe6JSoU0hoxGrK0S5Xeqya0p0bMnuez0i1cxKAj7
QMzm+9vC/CBgSA57hlRuVZgqP1fxeLuZJb4clc3iS5NDs1k+80UHDa4FfaRM+Ey+jJffD2Lba3aE
kVdZqFzJyQ3LOor/6OQWDw4CIbCuhrqlTqj0y/4pT4NJos8nbyTC75UZgGbz3aerl0rolzzdjC+h
KlUJSCfeQGQcdPvkJ2q6vvCD1YFhv978Fml9ZxKlh8/Y8K9g/n7MczT/Z3PCpuG5xGMQ1X9gEnm2
6hVwer9nUYuXbWKIlgmS402EXTTFDL+ECD/vnsBRWKwTIpQwP9TiLxTI2BuNyM/Z+G+rLulS9jZJ
EogzycdonpNT0gVz/YEmUG+247IFzVigNAmwK30VNvJ8XTKNc8DS86klXSh59VK07e4EyTNPAbdv
RNmNmhsqME/73awPAGn2uybUtmltMOVAHsAXcgtoX77BwTg9s4k2EOQLO9eayaegbq2UXtpENJPy
k0kqrZ/xqJ6RFSFJ6V/CME9lQWmVlBn/wRpi2DRX8g8b7MVi4fHBAqDSKlX23UmJTMQ8twdaJfmp
MUuCL4B5AeRMK4UJTyygClFk+sdiN6gDSXEuPUPS9oEZ+aRu+5nLJbnQTA3apz7j+Pfv0GmjuD9S
j8NwcsZ/RRHz9+TqwB1owa8PKN5NQI3LZCXBabXVriWcXHsh9Ao2HYjCDXJj+TYr84/lFi10t/7w
3LuPMch44APj3+tCyhEk2l0ILDPeVasbdw+UhbNHaZIGsHBT43teUe7hBH8rQkcSWRTXAj/0MKSI
rwCkV0dl9Meq4rwnDnIk2g79s++kmsejxqD1HPlzmB/WzhKlee34vEhkLhAe6Zsne2sH2gu5xvde
QOIzaZ/plGcXBHDqNooFdr+WGiE0Uqgu8V2FVCl/7vRM9d4F4As7SaRYaYbpLj5KQUCZxMgDUlsn
4nN4pzoit4D4CZgVtTN/XJd5CUjZFD87iS2l142Ffj2lL3FSWBKqp6q8B5Py2j2tOTExwm2a+uEn
QB8GgCwpm871Bq40mwwZPpYAH1+2lRJ3+k1wqhZ9B+JLtP5a+m4v3ykgV3i3Ps+UnQOyj6GcnJC+
x72RY4HkJSWh+Uw6dO4ENUplXuuZcJGxfCHaQn/8q2Qfkr0B0IK4LOUHRDdX38JhNdR65lX1yVup
8plxD6RyLiEmLqzWkc6z9oE4gjzbI6ZEGQKAuB8FpOiwxGdIkV4w20y0tG4udSFwQhVkSSEN3Akz
3+iajMk5uh2wO4FE3tyc6c5KE/AE5WgUR2i73i15R5uHGziouYX/wNkhCu4DAf4DHh5r3a8EokdR
GmvqFt+wFPf7we0lgqN50KZ4E9ksLIRuuXDm+wpEAQ1C/0XvDgIp6eSjad5lWtGB+lSmyYHzn4V3
XrhRJKJyYPilr1Ztuhlk/QkIjHYfUpRC1w5yD821lsnp8OPRpya/EvXf1qKbvksPsNgfedNwvGND
axY+EjyfzC4GOAfmdUE631/Drtak5AAmaGzBfB93g8GABiz3e3QbMyttrwSJ+FUs3DahYSqptCoA
jDIhV3XQcorlTAwYKNKf7r2L6G9C7WStbVTFgJwDdtpJqVqom+80MHCPauD+d2tCMd25dYxe07Fh
5FL1j617+V+DPTPu9P6SBoXgHQ6w4ToyKse2TQrDvv1hyNAwXAPY5+mWDX6aEwQZp8g5QmqzEZV9
2+fly2sJ66VxgWvw7gJCMWdkLucOFGRV+rireLJtwJLZ4UzBbRorfnVbbjQV7VqwhimbBBW9NTol
jYM29X1WZirQ+m59uFKB7s2QxMo9hsNfHJp/SiczFNsjTWMPgEfLNoHGaSzpGwXWpV2Ucy+nJRRd
BBN8Mp4IY94Zf4x0hgCE8PaFyTldbgBFfE3yxKez2FiepllpBit6cyt+5Ggdenz/RgRk06kyRsYO
lfSxDsZA6n11rKBB6KMJCUw9CgWpclnx9EuBuFRyBhQGPkFP8MtEX53zC+U0h59sG8xglw63d2eN
Q+U4N9/KeixhlsC0BUbaWeCsxoSBdZqSKAyCrbhQbtSPLQ4y0wpFXySE36mKOnL6pUaEQ0VgQE8X
NVox+TqdTYl4KHiMBUn4rR7nzLEARG1A0VTfEHggC26hIR8cMCwY6PR0SXlwI/V3Vr89QNy2P79C
SibnkZJ6lCquOIgQLE+IqS/Uv0SbUmR3vFPdjCyn4NM8b2M5gvUlrTrH2lvEv5g9GbmFfOiF7a9g
fz1ntIPGL+eW7BMNOFPKdnJ58IKAMhgubAnvbivS7Sbc/W99XEpZm04ZRuN7sC6tXvYmLSb6uUpk
Gqm3Oc/Zzwe7/QMe5qnjPQxoi16WuNyo8BoNjBB1IQ4RkYCnUJERHHTO1x1qbxjk6xhp9Ko2bscK
9NwCj4cCbB3Jw+jxXHzUPvSHWy7RgUjf9Ky1kj9iLugrdkDDBe2Ek/YbTZVMj24imLkuicNdHFrd
9HsPlFmmbZ84hVaFCYheGh+sBHJ9PKLl6/vz8JyeJxWurkoPSOElj5hbow1OIMLqSdQv3jrDX6Vo
ZpfUPmLkyBVpWl5gdtZ/TWpceM5LxTSieXm/M65LuQEZQJqh4crhvykta6O1KYzW/8rEt4XXTb4i
79hGrcfxRrAb24My70iLcdVa7SlErmCDo1YUZ6mz0eIPvGseXXRungB7ad0PG7y//B6Xbs8Op4Oo
+iJnMjJaqQlMGYvTtC00lGfWipKOghFxB5Pl27ibFtHUjueVOswRa7+E+CJ0HinCIXEqCIJ4ZZli
pn2KFUTwaYlrgaDULbusNLt513jumajRIsP5xhb8UnthNDin7ZFT6uyq+C9D40TR0vMA/PvJwMSn
VSky/jlJTQjHS4K2FzyW2ajiVwKFQrHi8Sc9RH+KjQyjHW3DJGPBBqZ3h5Cuv4jbtU7Pns48QNIV
kioptpdD1r1CEtXRqT2QdfNbuhTIJXhO89BYtm0hlmMS1BzGCNJDfw0UYE3iCgxixjfL87v662aa
yop02BEvo0dRT3taUy1x9AKkP3N61D3FNPv2D4I+0je1CHXDa0Cc59kDMSN74YY+4xfiXlJc/n/U
61sFMsekHw4gJpZFIdlzqtOovQbRKtErDh6fd+kEKCm4T/zCTBsUIG25bPHc6oUky4fuCF1o14FF
2WcAan7XTX/+gno5vpuHUszcr6ZcbmjbhOkEpIQcBFbLeoKXa+ndHlwZJpG/ghEWovS+9qCLeXj7
B9NJgymCCZnsKHjzIBMNUNHYuCVLyehlCcz2jh06Uq7Xq1oyK7RWKnXv422SeFhfjnMWySNjr/i1
/eHAhUg/gtb1vzxRiRarbNWu3GSmxMkXCeOlAq0Mus4Al5LR/3X6XwDoubYEg1YF7YzyALqgAUiO
HiqYd2agksa3wWHG2eE7TEUJ8Ks0Egx+rG87Lngd1IDLURkPTQrkNSfFkKaMT7OSYGt9gwSBJuqa
TZGovAMGFlFAf1j+FYakNarUS7pgpWErRHm91LwDUp1Y36P7hduTg02kM2pDtrvC08xesNYps68R
N9WD7d+OY3dgCpMTyDhrK7V3DW9QXvxjT6UDbHGZQJgb9mtx7S44W2LToBXeC3WIvxIpGIWpatfA
6SUvk0j6aGQbrt9SdULCIErNhghfLQhQ0UGJbh/pab7H1d4kIYZK/0mT7qgJgoeXeQelvX0x/exY
MH9h2m6Dn3x78U0O/kSw1D+ztIIWvd9VtGgJ9vwtS0MLUV+SDPCVXMk49xkoY//q55ENTKv5DTgF
0gRTW5E77/MH2JjFZKpSM5PncxzpzJei4hRNvhTm/1fulsFBH64SiKj26u0ObUK6YBnGWBT3AnjC
y1LuzADtH/+pbXda//Qags2w/8169/1ZSlxSKjHE+FMmvIyGhGbQlXPm7+z8sg8PqUjG5krw2PGm
0EZIrEZnfwHDwAm0ig2ag1OEgyxgZS+KMFS2wjKmEzpgJinUyO1Jh5sjC4P89RlSh+2vIIS3uYa5
CJP0P+hY9CUxDEega7rccyboQhfH7XlNeT5+RsLdv97VgeDBxz1226SnVHdliVj0gXfxVMdxYhaE
pWxczGvRna/XfHNpkJ+36t3uucf0PEKjCDQT+0Vz6YeV6sA1sBOl8n69j7LJmbkq9GWg35lhcVMA
pwEYBKNZMmBj1asaXsapPW/JfQ9dy2SiO+bGaKvM2QRQkF12O+PJRUF61EQMmeYoGuP/t9mylnXl
qXmJG1L/IvQSp4HgSp6c99oF3KAIb4ty9NMry9ffq4+ILk/uznoTklq+t6QM6c1wmFxSdwEy6A0R
K6z4804UPY+7yRNZicKlVx7VLB/wOv6U02HTJMr2TRtNIJJoiHax7XVJbJ3ze9W1yg/iF4aUUixu
qJxxHkjZUDn9cSR23I4rrn/dzA0iH5ZyYkAiNVx5+9NMUz5sg+LnACa/iV1/T5R1RX8T3nJ4G5uh
Sn8AbKvCKbxytHLKFYBLL7WTonwHi6KqyqLaHw2hI73pdmLr3H+cqbM3vBystqMWrbpU6Jd9wJoY
qNpeFQal4oJ6nkJiL8hph9jzX4NKAJaeb0YSREVPdtcy6YDz2vqF6P9vbRxz+eMsboPKOgYUo26X
SSq0G6YaTVjRDgUZsOK8JtK665I9wxz7QJQmgUwXjNaxPIGVgUmaDTI3Szc6EdNI/pbMcYJrbe5m
pNLHppCiZBNamlNudvybmQ+OQHdp05zLqqt8rDROUSPnUUeWc8mGLsvNZ4ncFn/roA0iOE+s+6qZ
3Ow+ZcPvFPo9JdIyuMTCXupIU2OEKDs54ZsEB8salitgujD0EbM90PK9cj/fE9Ib/P0n/n1RDxwZ
Ykf8dBE8u1cTh9UhWxfdN/QGCSXu9WgEUFy3xnYlA+gC+Sxsx+7yGWesdkUy1+6LpgTEPHk/U4TW
PrSvKFv7YFKXhOu9UhB/BF4TyFS9cmVug1Pldjs+vJlnSWjlUFWNKMTjGAkAs7fScaSS4OthIjf4
+05sktwptBIdwM4gi2IPjFfMzF641M84lEbDZzBojwCDD+6KmU/b81uVj2+0l6ycXrmns91io0Be
++en9wefJO1KdH6u+/m7YQAcxePR15PwDHlxLWRBIFKBttfsNJkossAo+lMuG1J3OwwjZBEXEdUS
t5EVg4imJuCXFR1hXDqqYzxENmhlWU5vPgD7nrdiuPLggBkjfX0v48M0ZEZS/8NXVLqQeH+taKz7
v9TNbZcodRZCCn51CdovGvPymIkj8CepiQtEgHk/NASF0W8B0DcPXztkQXVjMC71wtlr+X7rLcCq
X97NgNx00UPDGo7z0ffFcxMLmG1xCTNSOLf9OHTUYA+hd9MGelwq6kFYk8P86Tfp4UD3K0DxQhhj
WBdswXsKeAB2X15sCOQu8lbzXW3je7+M1DDLSQM8l5GcBo1njstscqHtGy4AhQPGQMsh/dC0q767
I4MyN/K3/vLvjIa9dLxtED3TFimGAbwSp5+lr69tPKGCwcDvl3E2bd+26RRUixy9ciVEnzLg2vyp
Cm7M/w5BcPP7i9yCot4RmiijDea9/uccPrYBDFe84vy1puTXg9DPxhfyE7aaV3r3yMG+2VVhjxYe
OvMDft4WJ065xG2Pq0Yo0pEilKoJPW9FEdQmraNMpc+k4/IfdkFuyf4FlLd/LVo7/tHFAUFnAZiQ
IwOQp+jp19QImq61d347G5YLDcZ6q2qTNtmJdfQfLq1pxe0A7k+7s3IYlt0x+gmeVQxZ3BABzhpf
CKbA1HOyVO6l75QP6Z/Eg1bQK44nyPATOZtYm5c43ZLYSdHM72crV68z02XJgWXhMZNxbjXMHWK2
GIuSiOBDMVKcoXW8xfMzKi3kHiMA1zEVD4QriQVXNTOKocaD+Euegin71k6BNtoJHykg7JhoPcy5
XUztjfms6uGlVDdPX42KEpwoyLTMnhzVxeobYD8102IQBYGdKbNsPNiZYWbmfb4CUkx9KL9XRR+j
phVV67an9HkklkoiPZzw+swvLxThCW4lEJEUldEawZ6J6j4lZjUCZJAk0WRLomshUeXnNtPMTLLO
HwC3gQRPK3fyhOUr1UC9Gpv76YlTbxcwFtBYEm7H1JF0FwFV4SZrITTcqPxrgmEj6mCw16RaUOPS
eYLABhxj/KWRUvGQOy6Aquj44DMLPDiGU6LVbcubQ8wLh3AijT2NX4pwVD3V2rxvZPkgNSDL214H
MqXTy68QSqaFFXQeEWnX0k0AdmDuvUDKrDsL+EICzIHCSwq57z6EsNaYykKReNH0wFoq+7hxw4E1
MCMWpcc3LuGOcbWTqlR/zMfEQVtmrDVwtscRuonkz58qQyOAi0fGRpnW+wDc47xjtkF/TwbL1hWV
KbHeBGdVV4a4YJ0S+HS34qHuFF280BOVuNJUFIX/R3KVJ6bSCHJJzPiIf0NQywW5GgTUCRbff40n
GyGEUOWaUZLvFM0w2PaTltsvbwxdW8DeGtw0OW8y01q+r6MTikjr74a/ZqN5MoDgtFy4vqATc7KO
uVrfWitnKB9uGo2eTxj2uxjiAeBoUi2okD4Ju/MoxdGxcOF1+fIbNKq/Ly+Dk+qWQNHWUWwmWJ+q
4HlXWAdGX1bw88c7oR9kCWOoM+Z+di27CLIDf9BeCCRVCex/RPnKay1gWMo/KHhKecSoO3v+fQmR
4h2SIL2AjbMGwb6dS8cOHgHN0LBbnCnwR5wvkEOktKefDRom99q5PQ1cW8Lmwy2a4CJZAk2ygnkM
PXcjTLTixBtKWts1LvHvJjLIs9lFhxIVF/6IA0/U2vMvUxEqoJpAjKq9Ot3f3iS7REqgMyhHW0AJ
6wiHp32tsnJG5HYqtqCEv89YaKM85ujl1zLBFfO7KOApYU+lbktphzQ2BwfKYkdUF6Jh1ILVKUPv
Y3+vw2o8TUrkMOs5TOxqxfUtsC8waBA3TR9OpXBsGbsJ0ovib923a/uuFClaP/sdgu5XZldcCujW
eJg5ukCxIvNDGPpj/j1ABKVN+/4OBfGWm2JOncyhY027m3VyvXudbFP9pCT4H0Va3KryPCK+JI8d
dOPhldHwd9gzVQ4fQ0Q7nhy0PDaEXzbBhj3gVAUa6mhE6gFLDO7MPlpNRGrJNtaAmE2EpgU3pC5f
YW7FDD3eywzuC9fpayki2OCb7M2c+8vzwavdz4alfIUF9YLalSG+DA4KMtc9qgoXYAFZRBmFJ9Sc
/uOg5XB6tKkN3TAJAQ2mWX2T+GM/jJZxxiFQfNV613TQWZqwFIILB9ibu7l4cegtGoR6cswusFlA
p+Emb3EyZIZ1MqlgmJjREgBmvXRRetV+YoaYPi79413SZQOOcv6AvzQbXnRZ3JNVvkjXhL/amX1z
PSYALLYzO0sjXiYd6ttmyDo5N0wn9DHoMAeq6l0dE1gpKJeACcKDq+GqMI+cNhO0h8C12t/xgKcp
K8hOrj91eZHPv051If89IqweORzD6EnLxWtC1cRDYn/m3z1SdY6wWzayjz3p2rnSAs9D+KdbYXfZ
P9htvC8373M/AbgCufTrFgJ3KPyCIu5n4ritAv5SL0Ttwf5Q3bS+sgbjKOJ/tMk2G5O6Appa0xyV
svTmtFmqcr25IqX5TxCDNXeo6+9wAmgDE7q4AIMjo2aP4bfxDB5FnvhkSPsL6P4yhSXgjIjw+mlH
TYNDlrPV+bu7HW6Oe0UEM39RJryojhkZx0ga0xIBoBCG8/Mp+06JMp42uAaxLtEhaPrBhIDhlSQ7
TYHfMv5QIkvbiCJLNY45NuVXy/J3VKb/smVotYvwvAa/nTFHM7T23TNvnZJPTd/+YJ2ZIVhju2ny
o9Phm/Okp9pq4huSLIKXKubQdF7hYmX/8KczdmaBbrtFLp+4nt/3DovcIU9fkgvF2TPXNGrd75Yr
9HAhF9IAO0++ujO89qw85T86u9AWGccCCu9OilM1HFXTmn/lKT6gOaPuqMOVJjWy9HARgogwuP17
twajO1cRYUFzX9jz38pu0n6ATuKHxP6Q1KPLDIUHy/9mkDeElKiMd4PhO1QqrTQnTB+vOa1g9iNR
9KfAzeJiDUlftN9WD1djVE+MV9oiDvtkaIoIUBRYGUwnecFE3rB57SdQs09aHBHf3DZ5nps1zsQX
JsrLKNpnDEwjHCWKiDhHdbgO4YhxYwuPH6LlMSedeO5QExneAGEuNC9PRmItj4y5CMih7p0PcJ5h
CH2l+KeaEFi+elRr23lAKTyp8iJSTZagMz/UEjolX0bT80QWqbX4LWOtwZ+d8hXgPv6SpGBqdrMZ
vSm1+ON8oAf+CXERKH5xFiT4oHblFFzIQwTa1EfVN9V8Nv87UqnSlAy17WHqXTFrkNIlYBGsvNVa
HTGQY769Si6p9eQfPB97jVH4ZvvTDiT15I3ECl70rgvepcoUI/QkqbkhysntnLwGLHWWxiixvPvR
izuK7QJHP2fCcuCZ8A3KXip5YvE4IxVI5O2mPFWlwksoZhHhKKNCoFmOwEfwfVCHHG1iYDKgt2xN
+5U8M0ME6VoMRBtz3zFwh9jrWhP24yPD+X++CSSBQZL7bpy8kZAZ6EyjNucvY2A9zIreN792OoZ8
t2cS6sVthUPpIKoHqYe6xXPm4GqQdEW5eJ1nraZ1OQsR9TsYxi0WWn9EIC+GUuVfng4dA3cicyKu
0syZ1WPcGoxWRClN9mVIgzK2N0guwGox2G5lM4hzffb1hUNVywUNr1PEEE/0ai/59/QrPiHxRlI3
2DQ6Z1xDlHFemvojJfr73AyqiRtnFrysHyjYWCiVxZbiNqsrSS+IYiFmGOSkwt5my9zCCL+Rb0Vx
h7illZf8cHQTQcevYvVAEfMVduWRv8VZ2aatcij5M3JHWvdyTV3CmPu+N4T9247ueSYu4HWBuNti
ZUiXpw9+bM69rCr6ZUxzY3gcm/6PDlcoGAsrEz6qq/OD5hK4HOnhqttTPhmfx9lqQVzal9qFyBPF
Fu8n4rF76gi3wlX86ogEbu+kgr5iBO4z2movKyHQMHUARLgflkNO5bDqNdAsNFc4/A+zKroQLr9J
31I6FmFl7wWXA0GIx9ZTtfd4u7TevHzXA2/PmIfVN74TCHXeoUT++2kiIW5s/Gqsxe/tZKoJnWP3
CsdqdVPUX04bt+vGoeOhyNMT3l2hr8J/9jHDFJgXBxuD55bxzukcJS+NF/rL8mX5nc5+1P9mj97U
XkMSEN+pWxm3gLgchG3szPSuzskxwcJf3ax/QBrlwUT2rAUZa3iEPNRQroaPSK8sxuzKSw3qO83+
1foZKL0ofSI4XyCv+6TWgwEnBxGna00Ntdzu68ur0mWfxx7rs/cxwvSqb6UtZBbu9UWwhj0oVEkF
lEF0YIGfQZ/eY0hNwQopnQhTbVCk5EgPRaNTf+CdMkoEdin1oWNWRRUoY+KZFHn11XDleQFYhSPX
NUWVlDHkfKxGwrWtAuZnUGH+LUEBlYzNvWgbgOrufWAWMU9pCRjqQGBGhKPdw/sqomgsLY1JbuHh
M0sIPais4eyYvI9/SJa5uCmW67T19jcxif/0G205wz9VeAUajnCKIsZiyd1VaelUgq96WrktvV5t
yhN9IRxo8yQPM1NE+4BVLwjh521jvirOZrQRMX2Pi/QGM7HT8g5yDPmsvQt4OjvBE0SNSu0X+Lc7
H1SH5xHf6CugjTZUwnaJwCRDcClXsiLIgNqY5sGFyjGc3ySd3W9Z1tIpXWnnZ8J6CKpK2bL/Ja/4
ve3H1YyBy7IQZgzSxUA21qTkIE209bPpWx6hlBjdgQyRb7kE3TMVQcIbSBtUAu5XuzJsZS7IcSZJ
TYbM1HdS8ZtE6qlzutHadt5KX7p1KDREZ9iq31ZF1/EJZ1Q55077e8aSp7K3YaW11CMBVWL71mak
oDfDNyndEeTfCJ1mLSl887FNl4AlyE7h/I4tYEpALEaffyVhTfeZNPJhNbQKy+bjmGOv/iP1UyXl
eggdRuH9/FxoP6hwEPycOPypUisgqIm43wlrYLLkHP7lWq/LPjDWxh3i0wxv/O659zwE3s6EraSs
L9iDGZ9WOJ5EKO4+dEmBb+O3geDqTPqSIpyR4BQs52p0K4ZKcw/ZVt0nw+IBCU9ahEeef4RGeizn
LPHnfduMASth3PlX4uKSwYcSU+NXSdoKMF1tBNkA3U+Wh+aLNT+shIke6gJMf5BvBs7X/BL01XuL
P+MHehoP2yTCB5ZczPaA7XVLGsm8te1tXMexq/9dCQUdD6+uTTQN6FvNok4R1rM0cQpdTdR9XE0D
g1ccIYuaZfRHdJSgO7+yGxbrGvumaNYz9De2of/9er6ztLv7G5TZhIkfkp1E+/R3KtIPn+AQ7MNH
sQG9hf+0qYREzFzl9ZhOAwExOY/piIxLmIh6poLmAh0Bl3xLT4wCHFB8Ye0lTz+yvwzPl5maqxcU
+oCmsLyNQyJ3aySLP1X9801wvy1PeYP7mheNeeGTVODOCDpHlVhIrnNdXOSEesX4ys8KYaQbYwzY
MteZMSGa5ZXyO/FFSnQ24ku2+yatkW5iP/hGgn+e7mTI8XKUOXrAV3NAv6zS1SiZggPmKo188D4k
5zRDqTERlH9TFEmZqKpo96UGpk1qNwA4wE0Fus/RNh4UGTMrqUnFD7Nmr+SPDUkwzhZ46A2/V2bh
Tu1TPwMjUyKEISzCPBSf1Fthp0mOvq2z1wu7mpF392aMSGJnHLUt+6hR5mbGBjw8LlkfIyjWtNBa
8TObfahpHlvrf0PIFAGRzQZY9cQedjidPAYKkbgrh9Hp2SaJ5IaoK7RteaGHoaM8DSkCgt2JIoI4
SmUgitdHXbITCFQ8n6aiWy0oLdwHY9lfanPKUbmhF+fPG+i1GoujnP54r7Yatfizkf/OpMcxwG4N
nODN5RYczGKGIqyeJJzTJtVkkTo7GarjTKCxVw52OFootOmCreBvAhH1L14xR589xNONotCBbCwV
uOVBDJDyE+iYuCcgUtg/dTh3AUT1smrPz4eMK01vEBTm2bSaIo9yaqcMC67U5yFG+TmmSfZrtbL3
C7yO1hXDsUBNRwGQlijdBmUWQk5Ap/r+4AUPtTkh7/60jnvkjm26CUp3oqyul4jDV87E8Lvw56TU
10vfwXmG5h6o0F1qKz+MA1GexOq4bzxBlUoUvTXx6CV8tlbfTwq+yM/Pqdn1L0TYkMIj50pi4OM/
U8MWyvLVI1q1EFUxz+cSM0Dem0caNI7bN5QFAVYvwaaGNq1Ymwp6nEq1IW9UCQMhPauuOC7ImuSg
UMv5X8uUMW8e8YICrqRRQ3lZJd75MyIwryUHJnQqgQypnI7GiQDmOhR8SaaUUwbYApkbsseMqTbX
hFvvQrK0VYWE3RwhXiE7GRh9NJfc0SKXhYX+gQNvrUgh1LXyqc+KhdxrUPjLyxOyc+0SkqbpgWuT
pZxoe2/iEa1BgisUhkeQHSdgRvxhf+FV6PzoCTGNFsZcpAI8bhdaoVuJJqtXMzs0LW+GFr5R4/tg
g3H7M10lj6FkkG3FYRoitMafTNp0EpAgWlfVyn3IjeMG3ifCH6RA8EmdWVjZNrkr5fx27PP0tQAH
UkqAUY0qii8HIcCDV+Q4Myw6dIBwYu5z8OXbzj0/UMW7+gobGSbDRfUGimdtnPZgqYL/FNPknmaz
Nv5CyMd8/R0N1umswaFsK7QB2KoMe6gh88VddbSChmmjqJO73+OVAcK/0pMOi7R4gCiqIzJmj9ku
ZifdhByGFCS3v3DZcC1DmpcnyEYQgRqLWcd2D6wpkOwH1GLYZ1YAvIKDatdel0fNSLTDJPUkggEq
IJAJcD3YigApWaYmrQ0lEa5lGrFXTXrlaLIJiWwy4J/wx6smQXAi93/PjZYg4mXyMoeYJXsjDq0n
RJ2+UjtEPWkqeGJUKauIqM+SgbsgmlADdE8ubfOt6m5Zg7iytn9NeRv63qKcCaEPhYzU9C4VxZNH
hjW40UC/cONLWNZQkzVDtmCJ7Ih+4EOwIm+SS2JzwDfKU/vvBMcBV2OJjEhwjkY6UiI+DlmqBXNW
aUve9j7Y4LVyAKGd+apu+2lTptiphKkDOHfQIrDPwEtKwUD6D+GGvk/hIHKn1PH9QzFx/Drv959s
HcyFopzDnZfXL6GolBOW//ywO0DL88cqRyzcPJ2EnYgqDsBCxDXk19kDh+rfn0ti4rJKA7mFyjbN
ef9NjAtqCiPmDbfvQbQfdPx3LWIoER8q5fMKVyQE9cZqetwtIAY01lkEAllOsPglZ97pyDADC5Eu
sI9Y8cVTL55AzS/FtbI5Dh60Gwjwl4JclFnHv0wHrxkRhabN3nPBLcRn13YrEG3E4MJVKlCDW/YL
Ya4uYZhjYgvIz1WR9dVkhyFbmPMDxhDz3Sgc+qp4CkgEGhTXCfUAV4LWC+K0Dr71STj65sSB2/bB
bF65MO3il+ofwblCoQCbLeyeYQbt+Yk55Pj2o2FGSRV0C7QY5kXMq/9FDM+gihqXa5eRV++nEzGw
myZH8ADOzNqWrmbicynafajPez1c6cGFFOcDBTqaU6mBCc54kKPUdN1xObsIjFRuV5oDHPhVIFZQ
iWkImyOarJkKwU+TbBjklN5ifaRPsiNY5ueqxXPgBH0+deBYImg16FSzEKMqYY8ZzyjS+qG1s5Vc
1wpjHXFcrYkLvlmyQkkfvz/j670JMVhVF9CErKhOVgy0vqZGbYyqEA8zxZaUIEM5hqEpDcKJ95dH
DxUA2N4L+WDY2WzqocZIbf6m84RnsqQpHlICqGCZ8foLlGXlbDqCr8PC8SCovet85SfTDR2/4JcQ
uiWjfguvMfU5O53YZxyvKexS3ZDKM0een87YbayE8EIbCXIa1samxVBQkVytn6CgzUHFSg7fxLsY
RLUPmkVSUOkQc48ZEiDD6eOR7r5Akug2VDFKCRirC5JJ1TCA1aUxSIA896g1jlWb0iTtWIGlQPJA
l23PWinDZU84vLXZLZlqxdT1kRUjI0rBlkypWcBKQMBRHogXP/JyAEyCMY3kSoDd0l5j1o8igwMl
v89PrgcOoi+FWCFeSiEJZSp0Idf6H331vvYgiAbOpiEMzgT5nSurRysFJL5Y6v5eS5DC0uS/3N1V
ItEu597HsgDDYq3lnSQTk0FthjBJxWP/ARwFvj7QVhNxTMUaZ+nxfNWv+gB/qZFQXvEKeHcZRH4A
XxYc4AK/ydiR1dw8KOLJa9X8dixfVpAB6UkArShO2aML4v4nMG+U9n5P7dGh64rkN2Tn8HUzCnok
F+J3tA8Lc20qjwS1UNL2BBJu8zgxyb1WllQvLKT1ON8GBc58WigOAPQK5Zusrbmv0gqymFN7JPFf
pUA1jqPelUqiQc07z6CybsLxfHSx0UHQ/FkAVNgaGdLsSrbMFNKK7gOpWVxY7T1iQ0y9fxHxIaix
cW1weJ1ZkTMsPG1Reqd+WfG7lJyriPS1FnKRCb+fR2CR//9KHBLhdVFPHI1CDXKqFuhsjvmwSFA4
lEhwjau7w0iHYtVFNh9Pvhyi7oSh5vyIJtKMV0pHbfoSdOdzXwKj0mSJreGB7BeW77kWhQykLZn6
6YW8RClWECnHBRla3EOkds261oKdeyd+Yr8wKLkbZhka63Xl+/rgIMZEHJG5ewqsyQbm3wfT+TxF
AFihGqzE/tSGAC2fJC13Zv4iraTeDhFU/LL2QHgHfWsRQ/9j75BbuzoYiUS61woX/pEZSPlYPAMb
pbHRG8dkraOtIlRgOpcj4KGbyI23lj8hATnn8QkiMCG8KjiObBmrrm2OoDxMOWJCy6ImpiPx8bH6
vz5z9V4EaNlTrZ9WL1fo+X5+FNhmdi34bwCYrQcDTNahViPQvYDBIrGD/S6m7VVnrko23fcd8pHK
jK4o44rikP/VNtgJ8JUNKla7TjD28HV7tUShLOjopDxVg55icxjB0A5llgj0lpkHXCekRqT20HCh
G7MMLnDeeq/wQzC6Ta9C2bLZvHMrWDyKtzVm7RToFWmME1Ko0YumFTsy8PPW5V0OL4F2yGBlRWPm
BARvA807U3cj9gB8vjhp9pKmuVTKuqGk1PGkFyhzq4x0CmyjddTMdAcltzG3AxZZ+6YF5gXjW+qL
bZKb3ohsibTuJVLNEwmQ48BxzQwjA1GQ6QugX1TzPdX90kB+ipZ5sZy2+oL50txeFkVRzdlyGlS/
FR7fn+i0StMRo+ccf+ViXOAv5xXNuRPCtjM34W/zFnuADDgI35yAnO7y1YT/80CY738Wy037F/E3
YG25ZKVyuqrLObKaoVwuKHuJ1xhPycxhKFFt4hX4ymoBeTPjiMmEx6wMhBkJOfcgL6SbMhWlu7Ay
9DRKFAI6/Zl8jhlXw1cVLNddkkUiQuz/a8FeNNcgDGVUuzUCwkwaB4atKJJGMOoQy81tHJCvDkUq
W3UEWi3hrp9Q4EVUzeFDwBJWXPJX6+0nUmBaZZYRB9U+RaebiYmI6loFjfBNIfYhW2WFW87bR2OV
yBFYjOtsRQn8N9E5T0tRFscnzPLNS88iKzopzOFEwucixPDJMrhlFYYaonR2K0b9oAwQM9Cyjvcu
ZcbSLrAFe0FUxxyDbahCdnStwkKThJXJSVOMOFd5+1diR2fGrzdxxn5GuIzEx11Hr0udBxrEFmMI
N3citcWHeaXR3QHNsP8JDXLu/l2ihzf5s0dL6XvyBTm8nlt49PNVja+pV1VtXyDU1vsUs0fMfTO2
m+dOoBEJtMjQmseJ+7uW0Txa27IXRbsrs5m5QNmN8X76Zi1r+zV9EQqzYTzOslQIKz1zm99CDD/g
c15OxjX4yZlOBg6VBagxf4fO91qiuGnOv8RaAwwyy+a5JtvP/VSWmnPUNt2aymvM2geTA7jjo+Cx
D0px2cpVDqRX8jei0CnBvTouvFK6EvcpDiLIu5cvd1CEo+Grt/jmHpB4+sWOMpmy/1jyC4941eIT
1DHJbwSP8xBrZhQa3vQaNn7cVks5ZjUjSoCoUzJV/l6bUYk0ZKqfhcB7uxyhFmuLu8/A5bic7TuU
DiWFeepzT2c+jAyL9sTCx3iK+rAUNjyoHQAkWa0ZbDiOEEe9XBf0/wX/nNDZU472zML/Sz8YXoMT
RAcGY67s1b4FodZurbdlLtheURDHZ7pu1Us2pZ5maaV2nv4Fek5dnWRd1B0BzZtoVNZgWfa/OuoQ
0s79ZtAL+KZBO279qEDq7k023MMm+cGZC8xIoRepvobRylIQz+tLmzMGw10IPwphZjutWH6O0XBr
3Qd1g+j+I8pbZR/Pxn+Hhn2JHHzm/3DdVXB68TT61uQE5pa2aDGCFx9G/6+XrqxDALSP1Dzxqdg6
nmqxIbVDFQ8opJp+9Fem7QVnNAFN5VUX86peSdcCAlmdfnBBtLFTSbZtCrcB5m8PVVFtMm4k39Fo
iCPD3jUA1P8PNdIEBe8XYafspY1jZbd6YtL1p+XXW/5idmOjNe+AuQBf5cmwMzU67bgXY/SG5Yqz
xgUSBwYhavIcD0R1voR6e3tHHV4MyAm1UqLMRHEOf5pEmfGSv03VkWaQNY6NVGIxFhqUT7dgFjTL
MvNtscHKSwgwBFGc6J8iLgCmXma7yYr8M/Z1RDTxtM3iuF6rVFXC/KN0Ilvaz56qrOGUwojl//Fj
C/nxGY0GelI/mG4p/PCKUVJeQerP1uO3dyOHsbPBzQKYiYAuV5+n5+ir/ZNqWvMwV/BNGUCUM+je
GKKxE5qbyAGQ24JZoLiVl1b+6gRUuPXhe6Y0o/NuAOruAqhEwExxKj+eBl88ZbJo97mBMpn2234K
LPLPH0lhKtUaTfL+XO2BZwYaT+jQwE+p1UzzAfAh+3UdDiMx4qNmj2XJCFYDNlJAFyPPjWwdAuzo
26GsIQZdCVNpjhjiwnFuhzRu4G+mXUEayreNY8QmtAqvHSf1cBQUC47L2YtWJmw+AoXYAynMPM4a
5ELIexvvFw052W5hOCK2wrR2IXBmEvNTPoOij2YEIvl8AYz+Xv86JfjOKMkdaDmr4jqEeRtYTTNT
05HfyVttaAIQVKbrW0+KD/09OyWpUUbc8+jdUrSlPzYLZR2oH8jb9FBpA+iyIRQSzXBsh1FXeyff
aQxMiLahVUw0CV1sZ4afEZpzmdZqHkRLsHt2BN8kJBB+X7TEc5EwnCe/EB4n2Z+HJvRUpWy35VyS
jJ/7uIJavWnzOQjq83kG1BxchhzLay8Ju13ldg++B0cylfO+Ew3O9IyTDkKt0PBBnmTBpJYqFb38
EguLRPq7d5c7rtnGbxKq2O3rrTSoSN4ZSNPXhxl1rQf8tN3/dTGZ5WOytSPZNavyg8I2ixJBxJaH
/tyWaIySb2VxZixuT/2yBwgG5ZATp+l13H5szm/V8uMRuge7TQdzmuZnn6TG5KIxNp5ltu4tMry3
fgLtpsNbXfY7GF2fkDUJnfq+jjxmzu0dgYTh46sBRyVnOjDp/ia1UpVr5QtDRGygn/BpW6MM+nsr
6nUstL53K2Bea2L0I5ibPyNWgj/M1qGBnrBXtzqJQlBvjFe7hLm3y5iUifziFRL6xtPwCydy9SNu
mqWBFH29xGN/QyB/Vv3lb35lQbZJEMJILbdw9gNvwUGxpmeKwLrfuhC0ZHqR/nJTrkglaMoGcz7p
X/KlUl9JUI9D3H3Nuq79Wom5moQb8xtSghTzg7Njg5PquV7+bc9vSew+yUW6t9Ow0jSfQ3L0bdYH
ss9eqbJKxRqKtSKV0UmcR2hs3t+VmShOtj5S04v2VoEUJQmrbHByxdJ+2q6iUQWyxCa1wu/B3i3c
h6w7/W4kcukv95saYYcJjsCdSTSENkdyQVxt3fnivbXIwINlmB6bOewTc/vyirAY9+lLrZ7vz1QI
BO+YuiYvWp6vu9wgWd4MWgOEJTlZ7HL0mt9m12fAE2vASfEuLvJlYj7qb80+INt3j8tQF33zq8Ct
acVp+YN3oriRWWwtPuGR3qWaEfMuxjrovsEOLlWyaIUnx52EwpNsitRNMJEJL9Xsya/grSXazZHS
arsdnQI0qUEkk5pRAWX2GnfK0uErZCs/Stb29X37x4Tp7NEj7hS4cWiSJK08wmR00do1xNjaehBY
Hp7iJ8eYNYI3gv5kN16dMp93/NZLh4G/d8fQ9AaPV57lFcOcnPuexi9d/ckf9a8OeLp5flFbmyy6
+z/HUQB78m3mrskLPqtA7r0IdKZ7ejsLzsx6ojTwXobJVDbjf1VvIPh7Gms2UfYo2rxdUAcviRRl
e4QkbTaRgGiy7mleoHnRa+Rzngb5vSDU22L+NkDDaGdpxAD0PoVRSv995PWadem2AGPjon+fyQuv
2+oSTSA8x0VcTocdqxiL6UwI4lHdGOgsDXgfIm+u+IrPxir2CByiF+mDFE5j16Bil/G8GZFVn8c8
O/gmk2ak8dLkxW4Hox4DQbU3hqW8yEzouMJvV/hGdUEXO/FVeq2qfI63eMLiKrYFkkqf3e14t9TY
E7p/xgCZwl5TJP+nGOe3eY8RtoTOwl0PLSR6jQOfz6+JKKu0nGjHzAu67chtFNPJIrr5Ud1+1NMP
RNjs4mnOg46X64RMuqa4w5UE98GlsQX2obxmIEVvHPDahX63woa8VI4kmQVRbT1Ojiwn9li+SmTg
LyTd+8GYhLfHQW8j/3aWM9Y96GtkxItzWDqgYXDaHawq8vLk3CEeznI+RonFU623r+5JeULB5z4c
3mz7n0amOuVQG/5K3iPpXfR76URiM2Urn7qOWjSv8DIxTIqxBA1wbtDTfMWq/Ssaf3bLG2Sia/nY
NEapJ5zaNz9tjyVvVZ6gHVL1SszQwnk/Q4LO5V5l0wWQAfoEgfVO1+EYigLXltQU/B3Yt5CxQ9XY
xOAKf1zifit04Y3lGxvQN0tOPBSdTpV38STK+rXlLUzboKN69wPDC8ApKNuvbIkC7MKPYScB+vvR
OL00AUgy29G2rdvR4K8/wJRi2JKkNFkd6gV0wjjcm3Jtdb5M/cagc5ZqtW1TozIwmddgZj9LQAX7
7b2b80Cg2MKatseSQ2Y9x7I6kGeN3y0dPdyr2MWnVeFuCBg663jd2gf/E090UGV/gcvNu/ZC3Dyt
AsEAkT3criZHzCgoHs6D5XKXKa/uwgaRAGPORp3tKH98Fqs7JuS3c0EDx3ZnPWcFibad9jxuFrDZ
aqUpWfKwTC3QhX3sRkYjOYfLwbsEQOzzk+7kK616H7wnEITP4mhIzj8S1seKov80QeT32rgN+U3j
iobIDFmYCJEBSWpylRHVkV03Kzlcjg8oboIBh8E5+jWjoRNKFhBfBJShEHfjj2VO7gK3zKkFVgml
p+1jgAOEW5xXyXFYggZVYCkKfz8czs1BbUT6f4PTxcaFJkWwlbE9fhU4Yt6aU2y5tpHJEe2OZ1ua
7v5HPxzVFz9oBkrDTOqhvbtNx0OvLc56nXermVUcQXDyKdd+W1dIR2SokyU45xxSo6xbLBGa1T1l
J1WFa3hWL5ryp2nLPJPRf5NicB4CDEPBBFmwAkcRMQZ/8rST36oz3m2yrHBjIWn1IHApPcygbIyx
hBK7jn/khMfvryC1zF3bsh9nW4Mv27MQXbCYQhVWS2MY0mUWOLJm/1DCA3ZJjfUVBgsDl2swYIV4
zcQzaagZj8d1eThD4vb0MJ+Pd7twCDChaUiU/yKuuDB0nyrUX0BfC93OkBMjAEhHTmxwaXn9L/Ht
4uugrXwCgzf6PJkEfYPkh+qcuYF1i5HRK/Q0WLG8gO7Mv6h8PIDHdpg+G4FJQHJcjMBT3Vq0mGZ+
wmUf7WzLtmmhOXjbjDIfsy6DqA1xqw7WWq8utoXIS9gyH6tFgFf41aF+Pnh3PT8AVs6H7PhBbR8W
KEc5MmwFOxnWokVJYJvSfr6/3gY+mXue/f0hsYOfHRVMZfuNHLACyQe5VnlcUYsexktpOEVsbUmI
xuGAkcM+NqJOMPdq0iBUGNtUQnA7zurUenkxnygqbOKzuwLa7ZpWS8/STHNFT+jOpWO45ZO8voln
fLRV4BhQIMGGoxNtP7UntB1bHLo4iQcoe8lo1q4/mruQKNZ7oL2O2hjmIpyavn7t2mGYG0wMQ2s6
JBo4F6fFt9kiNcs0WVF9681pWOn8qK9KIW0qWeOwkBOOOwuBKB+tSU4yfHLJoWnOA3XI8+Y8pAcv
D3FkAHqB4Yuq99zCSbhVUe/IAxnVxmTx8WWVbW1KVG6B0xYOSLC+8QDFa7bilFapWfNKmeH8+TNw
Vi4sY1YBjWlrltZdykLE67Jd+QyUEpfmoGSsR2oS2OSMfLBoEuM3Jd/L/AW5OQ4Br6Ix8zHyYbU4
YPIOuf/yAkQ7fX69wmp08ParGK1ZJxgkC2tr1L0LSztgKNwP8OFlgFIkCe0IuYU+uBJkIrqC51Ha
WZi8qxteQgA/Tyhy92rQf3HIj0nkkJcGl0CBF0DiHHBOqetJlPiH80EcKVc+mbYhRjJUaME6gSze
TI8LLyWRusj0sdAdpYC46iM441xIt9uS5idsjfkyZmM780O/gJTFAXZkxG0jKqK8sWQ957ayQ9+j
wgl19dpd6dFGbNnqh/LjjYFK4TYAxHZ6rd/cEVHD3LDJpAyLV9RgMAMDn7oveFPW4czXOzql7AsN
V4R6347vPH04/fdozut//+zKvTlwRahk3Tks1trzkQRhOhtkqsVKjkqZpB74ATsR8Ncuw0TtZxfC
goufC2wYuCHuL4cnrpc0LsJsCkp8ph7s6yl865O1JTlE5+afz94IJeyw53A8k5hAy8kgn9gfEV/8
iYTyr1MfPEu5M30OQmu8U6UvYa1G/jCveTVfwWrV7AUsyx5JNcGp1QVTWo4TWXQaW3+sVvv+Ybs3
R7LJ/0xsH4VdR9S+ntzRduWrg4cAknPzBnQNDP9yHmDR7mw9HxOz6xp7ku8a4jxDZJDTpDU8cAFA
qfBvQVARxS6685ontLme8miN/vX2ACrozS+bgN8qbdg6i2BR7Qde+S4hT1oeu1OheFTINQeB+bRQ
14DREmpvw9lnEoJDUQO4hYhzFYDOYdHdTiUdwSHrEA0AscsSc///rOGuetwO4cMnmsJaIwXxQRXm
ukTdn2nvQvgnLpEM9GbdaQX8wKbPr4dEnHFnavE1xCOPPdDq2SmMFX2rmLVMvT/A7U+eWtsQXjEp
bSexoFOK+Ubs8BlKBYkvsvXP+PJlIMw1UOT28VVEXYXUjOjz/RmoaztJQVFkzT+14utw7pNfSy2Y
ZJEujU0CIxL50Xby/gTq8tQ7PV+f/zSyt1kcwidmRe+PrzCoFnQhhecjsL/g9fDJqYGRSkrbWR4D
TG9Xacb3W4CM3bsM1HZuqtn+43Zk7PS7nRA4T6FhPKzI4C3Pl6qlQ9a4gr1y4jAuc0oeKsLTc4c4
K5d6g1zsdvP8/I+FZv06l+z6UzB0cConaz7hmRHriLqozgZHPrEUFS7goPe0G18uY8eUMtz9lgE1
rYmZ6hBfgiS8TATbLqwQo1imdmycdXCWfIm/vOEdGX88hq8Mt8+w1UwRjFvWDrcMbz5TkqvaIWkG
7BrD24PJNli6ICDgI6ePZz9I/r5WWjJCbkG3u1sjrvTFu8AvcvoZjlEqC7vOz2xuyy3WU8gTt8EH
GJkS4YeSLT6qlqdMu5p0EL3yn+S++L+f/rJakfzcVW07bQsR5MrpBkYzIsX61BxEmAtHQbi4lvUl
tuWq/UpTkwTZjpbWn9nEP5zsCFan1sV0bWUXwYaqeqSvGzy2rtv3XL8+PCDHq0ddmcxVM06n0WuX
xNAd9fU46bQcKiyJFDg0asL2xSW6OwcnxjMLG2xEj/KhCbmFtpF4XD2FV1b1X335h/o/W//R+MD1
Zf3u24dT+jSEZxEpY08pFr44wLi+Je01y3kpwNfG349LlxBgGnb9XcqfYzBdhg9w9jzXqUP/sN7m
bLSOjzsaVQk3EaC3k5dh9Yo2AsvrsA9DxrmMpJ2vjF+g+uD5wRHGeFX49keUHe+yzIZ23p4WL2Iw
qfsTb2XnkA0ER5+AsO8NTcUPilzR55yJZKr0XdyWKLCz/NDWrQHUl9OaFsxeVDincWA64MFM849x
wv4o24D1kGLGd+kGTBr7xQMkYchF61bb5u40XsHJZwun6L7AWdMxsSYdQw7gyTVJS8ad1Re7SyTA
sRYkOqkdoMmAuxesCJUah7IjRmSIUWCqdxMD0l3BHV4dOR5DYPfRGlT+Hy5Wexnh5zJQ3Osy3AfB
m1UODCNEt5lhNjrxeDzP3gecoNS7S1aG2NsNNb2pAtrLEm+bUpRXTZ+RMxepeL7EqL2TsArtONQu
EEAXm97EI0WtvkEbnA4+WmbGyXBRRFXENAgIYa92YCs2Y3tRchnHq93WyjfQLwsQfXJGfJNo8KKs
mOdqQrRVT3+2StiYfZqrkO8H4d5Hq68hOrRovrZQrPyHg3/2baKFxSi2q237nshAwyQzFSaKz6To
GYsnLrcg/dREOjfNAmJky0MykzwSYpaprvFpUyvv8dtAkMDsGrR+J16Jgcby8HjZiBgY6IU4oWN6
AE+Ytgsy+mz5gei22cOA1w8p8aeuWJLgAImtchl4P8cxlhnlJttVRYJGbSM/sL2NvWQHF6x7OUYd
RPYGpEexpmQSqy5gBd/h+JO6rZrTF5WjGNCsqrd0Nh4fcl7DAypksWDGObtBxOMv9lzvrD6fwc6M
8SZLtZU22ytZGmdrL/ZdWkhy56JPeZ7sTEW37W4L9xfKucw0ANOuh4A6IsoPlAEwiPHPmmjKwUSK
Tl3uMLL2gPA8Y8owFlEAoXRrON0Hv3x0qiWKxxDzmEvoLsiAIND+mS2VBPtPN9zyFNklE5yjwBG+
bDZwiJba7zifwA8etbY9oNgij1/hQagr5cY0q2BrrXmgy7cnNVg7ZBLJWQD+8MoqfAVnR8IOclRD
84ArnDKrUF5Efnkv1zIVe03IKW6427QNZMnYKu41CPJaJLifszCyUteO94kzkEWcoDJLBLk9DdKM
W27eCNGMEN2kQmFzSmDa6yQ8grpE5DvykvIifUVtm1F/uRUXP6LcFvlfLz49eG9Sv4pXP6swuruj
apTLfV8rJoVkpg9GFSmN/BUqAhVmcWoaW9xKhtPPkHkaBI6+fVTOVkZS4fQ25ybM2AE2uCYLLkUK
BEtk31bWzU9L0vyIfaoC4lGesv4JOXuxNl+XTLaPuXWS58mt72OvxK9n8kpyiIyk4Ie2gJ8xQK7y
RZAmdiztdlLiTbaFJTwKqWpklbiDVfhe3L/t7jwf7zKRvaoCubznTJmEinNd+tbC7Ralld6Q+lbV
XEc25BBVOim2IZsrV3nObZ7nX6Tc7hugpRikRTkx5YqIweq61kBBDVMxgeHbdcB572jcEv52htzs
OU25L5yCnqkyz/FvLNTi2mIsE2EMtzzBlRSlKoKHh7EeB3kXgFGwIISeldiE0J6tFmkUUL0Harhj
bScTrNxDJUFXgDatjhG6LAhlDK8+aOirlaa8UekCITJVtgOFadIRFm4/fnf4oY2GNIJ98litieqw
jDOgTu0J4A3oABOzY/MdqWAemsPjOxA940uqsrH4U/cbie/gaw+p8UJKlAqkMjMw6Y9wk+P5bn3F
0GXnNOJ3cM6FvZFmD/QY8aM3i78IueUCPzRGED++htoBgyL0iFJpH2/WXx/hI1rU85lnsiPIZsVL
wv+9sZdmORL5Pjdzp8tKAx+5rniFWtaQU/53vZORaeBfteFUAsVt1sz86giRFQX/lVzC83SDxRZH
/jnoxseilsbO40aXpQMRKbPrdnZdtdzZPmjAjqkTHlWUjMYWXVM7cthHvax2+663WQJ7O4D4xdpB
3i318n6op+gFZ7y46hjo7kunnwsB6IyRFA4JbVHUZL1+9dxCBsjPkeYCK2mqOocb997ZOsmyYnhi
HW6BnPoSvQ2LorU131LAgtYvr+6EZnYKSHy8KO/K8apB2gSOUtXtpq3Z1dJJdlBqrI3tO2LwDDNR
qG4+YQJYyJeQXew3rCn6Z9BGbo8AdhqvXCp6jzJZvyVAQeHdgrDhF1kH+zAg76VuKLTYmlCfW0eo
W6ITO/W2UWWc5IMEtQZ0GC00ZzRHuPR68ex4Djgsuk2E+mnrHSAZYIIjSoCHKWIJaPCPtdVtNUWn
KAA5QzvEfk/C+2DT+ClIhKL3Epc64cpiH7SZUBoEs5FCh8OoC7FfVJ0AmcRKYLNplRIgRQWsbdPU
f3VdkQm/2YySo3m5kqPCvZO496fknPRqMp3kFotEu23WZjaQYzjSdeSN/L97L1g2gAEM+6LqNOxl
FTl/3cNXPklhMWAcrAsqLtSeGVMmZrAEII1K8GwAcAqvtT1P0rdODc5VOYsH0yv7ADfwfHOV2sYj
rsTWloVRHV7aULJLKkiizUnLETRSvT6Fe5hv4rpbqUr2dMaUWLUDnyFdAc0EFwJ0Qv0nTyIW8YIi
p14Y1VtO5WrR3RS5U+VM2cXuLl9BAPaERIu1EulqR7fNxfc1PznCKjqZk8NRBpzlnJ/SIBUhYdeW
SfBjwNmbvYT+jzjkzK8CLzL4ysqvFcTE3AWE6jKhJ4TzToq96tBNFnj7Szvj41SG6enc5No+03y6
LaJLYcBoQH/FCMdqPL0Zn7b3aQ0uy4292zQagA/kzTSPStx/MBu2qSDk1xa1M6p6AtJg0nz0T6dz
GlijmHyigG0pvYnQpsJDllR4K4lXNbnuL3w6l2lkLpztf39EHAlUZB0u3filc+SvQDEAvZzFT6i0
tMHjz0m8VXq4Sy6irYlwvpO5E/3GRVnWtWNcpTP7fN4rvENSBOwTU0zxTtfUGeX/nu2EiazKc4Pr
VqRoelNXhi3byikArG5Wz0lhBnqS8tvsdPi45SXZy72IsD5dM83X1C8pJVQH2Aj0zY8L7lehxOO2
X3aIHivOKbgWrs4jMTZJsQ2l6mFidowaIUDzCP8jXKNB5MhJqUYHLybwbNyvrIyJ6ZOjcNNqHBfR
YO75O9FN8LJXZ1lqGqRtc4EaQZiyNoN8Ng48QSeuHj+lCxwaLqG/y9FVZ7viOdf8lDeLRgyHl5uy
qsw+Np66jXweLgeFRxgI581hF0CCbZ4BTtqxW5YBTuC4JKiBgoCCF6g3HuFPP2b4tZoHCaztxpzz
6DrJ9Zl3cIt6XhGF1zR/mrBPQybtIiImWdMlEGA00XYmGj2ygb5txckSAXhIl33TIrTiwTe6XjZQ
0PPHgpGH0u0GfbzpqIQBqUsdkM+0y9I8HvzT67fCwLaKYQfpISs3ivxHVHDBRoMIyFE5lmsmz8QX
rbAUb5VBpA2t10yE0bXlNmDUpMJJcwsKK5yNLsRAIlnyn/RdgPgI1ighEwhQvqb4N+bnEKnfBiA/
1OnOkZfxhSzjTHF1l1FjfjDPjLgTbErs/1hHiWFjBPm1uiOIubd1RvIvrI8PXvqIRimAv/3d7oU8
EErLr+D/Hy0y2q+7xwIzoxeTU+/ZjdbtBW2q2GzLq55Lwwr20ghvJQ2Zej53faz6sHH67OOz1P6+
NFQ3qvMga1me/q353MNAnxCHtalCktqnnJci9BolO7I4pzCqvTJYcjaOrIuto+zxQKkP2o1Pk1rM
+/65wQUu9/A1eMn4hz18SKWYS91vc9z+2p2L3LeQxfa79DZs4BBZqH9FvkWywiyMZW//Ch6/grR8
nmeKDZ9lqHQYU2pGn2IztaPY9qASLIvlcm8WaAxpCRTw+VL1MNNaeaAuftFRIS+QdZXNLRv4meAX
S6rX7Wv9dIlOVUXoMRbgnqJ7xtO00b63YXlyDQUlrH9KigG8+TVJHaHMn2UJL+i+X3sQTmf0ZIiZ
J/8OivpsqixqfMtJJY/mz9MjVGAMS9HbEyn1/sPvxI95jdta+m5GERDll4MmkFHRszB7zujX7ujO
G6qNyDZJHm/sBYgsrRdLyRSNO+FCBOneFZFMo8Kfind7hGwfL1OGnrrPM5D1Q7NGUUB2z1RwpvcG
19rK1lJhW8KjNI869U0fiCHPfwRgLQmB4EsiqFjDUi0WvtjWTtdeP4AawwM8qGg10Lmc+n/mYEFa
KbeXaBnxktbVZX5Ql/APINZtUgpczjhFXHggrsGcVGM9WUKzBsd7ozuGurc1m4q0ViJ4XNWWgs2P
Vi4ybpzYlPzsHWp01rJBa/rRjAwakY8VD/lS438nXdqQ+sPUXlrYInEOii4ie1l/AVQUcyoCrf21
dhpjvhDRegh2nUGjFaTgvCPPujruQtMOCjb9GyuNCyRLThcGY5uw0RPx1Rt/oMAr+1yt3puEBSpL
kKbUt7cUVLLrHIG3gTw/loDUCT5TWURWR+E4/gHodRVyKPiE5TjGm/Ct5a6JipNP/YI96J1ZaX9J
jkKOMPEfWy6jSLmIsglN7eocZbZm1x7C+D++EibQKnhvBynOGEgs5vy07dBqPNiQUeojDStomPKM
fAjHxXq+8yFQMNpBCG5028c/JJVJZ8V9C36mqwgOCU2ENHpUOt5amxsht9wdArzHr1aJPiW1c0iy
pMv4YZJPFha87dTREGKaCgij1eptUGSG/ob0Ff7s3v7MQxBzIHjYt+LKFs871n/o7SyRRIkfg7Hq
KGAoW5Z8lbtpOV+j5p9BUrLDVR/H/nCNKf9g7Ddeut+I7horUPpdKm9DGcy1T1tA3SWZTHOjQfQJ
ba/YmBfjn3ETQmDqMLdfwkwvk+AJAboUd9q7u+yJuZK5VuUSOrq9Xk7VJbSW7EUCyaQXYyhChNqC
ilC1fGe+iZCa40N2NxJS3Tw3jR7DlNf4xhJogvBi0wEtOBY9Sdy0Bn24r0+80w0SdGcJZfesYFXk
DelC6bdR/8YiikkceTYayJkhCEBlTaC9T23LupifgWpsWSJn0Vrm8fYf4oAWdXSsuRZCRV0KpE5i
YNV1bsBz9kkXnbnmCmqsXV4o63Am9qJ06YInajni85ISI6gxESh+b5gs4QVqSqR4TPFDqpTUb3lR
VLsuGkLF1B1SBOqD7koidOXLQwbRkyNDrU3fd5sJfSWwuV7W2VWgg204vtx5O/AxxR5aH/2f7wTe
jhDRs+hYV6SDfuw6NRRcPW5dcuYfqVG/wHjIJcXbFA0Q6jo0QFG0p91q5KHTEQDu8io3GE2Dfgsd
65s/hGx+cRrr5KO8hHPSn98jMmzmgz9Jciy8bO7Y89Kit6gVtv2CER5fHhgGF8rhWlelEX0mwW1a
B8wmpeFRILKoXP7TUhEeBgWG2eTfJJhaAZqPWF/b5lPeKDwfztRDb8A2FS5UdVEbqOeKxgnxvtFO
048trvFI9YBYbKlYtaa67VV3A65sXPN+GS//gFBZEu5jNLq8Nn8XlmNP9hdqnrEjMu4MFhsfDvgz
0v52Ip98LPZTojakDf27EJUi/bJGr58DkgNY1p+YSKvc/FdxjwYXijLc3XYlsJkQeFw4LTHhwAYq
OszoX8SzuwVxQACD6E8VtHNjumy+CUiOMiqmEL4WBGgpnskFj2bZdoD++Z75PXA5Ip08UOU5dL/e
HLqEMWaBat8mjFZ5/LC3CZVLXSFNNkUFrTOl5KBZyq22+r251B1/oSHGoQqTaGJozk5bbiPSwDJm
TAuyMFDV7ERtyWTdgQE9P5N+eyO6rwRD+GOo900FkkTGBHOSniq7h87wDbim65SambB4euy+PoPo
pfeIuARG/x1R2X8FQ7EHrM0NPyuwU2nGqoIz9LT2bRrdbhM2vCNg/S5GRJlhlGWCPr48rmGPFvGi
k0Tz4P7UTvr7XriySbJuUkNvBBmvXbzm4FV2IK83kVjyJmgYnCyW/1xOU/CG5aF4UCKEil7LBYL8
ROngUwbdPBbBTJ5/fPMnVjjPAhaaWeyfaSOSsjQrzzStf6rtYv3jG+fLA5rALbnCJz0aMc1j6R13
9+Rj6iU4vPsijA5p0D3wb4J5+NEdYcwS+I+fL8+o7N5ltu+kXz+Orq1eY77rvj7Vb/MR+f36br1y
qObgmql0VbD10Io6uvBSIbsfzcN9jVBRChsXhubGf5L4dBoqnR6lcgzWtI1MUpONT3juXpQvTEcP
YPGPvHFlM0K/hwV+SqcRj7ibZ1eujIhjyQ99eXTz6xdqyrZsFjA2ob78PiuqVUbUl37CoJPSAXLB
a03JS1t3gwnQyIgNSy1xhsvv2X5y9sjtow0aO7uSZWLiKo1Rtg7d85GRL9+cEquufYmsMEYEFG2/
ghIDOUmKuGTz7DCdcGDRskOdmPFSCYH5UUk9ggT4yljtYWg8LbGgTem/AI1BugAJF5Y9RnLfx4Hd
KsV0eQ6/Lgk9Bjz9O9Fqp3H+ulbkvoO9C5lxOd0qBNvLNHY0iHfNXrQhf8mLB24BZ/WRUUhDYa3P
3kg3OyIK2nr4hdlX8eEbPERFFztoqbyMdDxfpKxgAZl7eIOtPSggbFNHekxv3NJhen/kBOlhX5o5
jYzENO4kAMpFqbIxRjGIJt4n1sIBvZ1GRTMkz1lX9FMG5EVc1Qcf+CXYSRy3XCiSjZSKj/g6dauA
IupV6/P/tYLQdwKiG9IavkZ6OHbQbztwRf2IPIzl/jdx5wSbs2WNjLf79mzDk1FDPQkwp8avT2j6
klparOt+kYJrpB5ftaxgXMp5a4Ys2y66H0S8IogUSkQWBErqAp/HcoLpowvl+ZOwpyKMzwtyKIrv
M32nnUYcs7PY/tO7zI69RTwtMaKGoK9GnPB/aBKCj5IolmmTT6Kag8nXhSfiZ/y8NcZ0/d7UVeid
UCfBLxbA4gi3A5cFiYIM5CpPMDjFLXLcv9N/KPGgrQQ1EWD6ZlxTOo+h+OXT1wRXzMFXKT1nsCjI
HZv09oA3HdxDKa7TDhGW286CdKpTHREeq+q8Cgp4+Ajds9G0TwyLOcED93eVckbrthnt3HpaQYUJ
yrIaa+36U06Qrm1eMBpUbmd60x7GlTYKbyzNj7F9MErvR4JIaWapWbBGrE9AccUBdGSk3RtFqxhF
3i7p7Ye9cW44ZaMEU5edXq52AYfrR2hJFJn2T5+AjI88gD3dAVe/OqaXaMs1di4RIgiw3/27uCVJ
28pHXKiycOv3iOl8Dmt3HEumRyJHFjEuOVjkbej9A9LVKqlkDwJbLouW7/kLgmDxp9z9VOD14mXX
e5y0lncCg/c7RvJDQSHf6ECKC8GcO7LtBuWBbX/CkMTNoba4xhyECvwuT0Lue5PshhqvrRPxxukb
vzD1AEOfCBVd+Wcm6PVA40ohQHsu1GP6FOiZQH+dRlx6tKPjy1T2l/ocs9sqKHohl6shqnxfTgnx
UEt9KzB8Rn0swwVao4TpOtct0TlfACSU28lMcPe0h/+5ozbE2FmM6L2F9ZCTmPQehLnGs1CMxcZy
ibEeOeryJfmYm7hjBN5RGpUplNx1rWRAswYeiylJMk+bMStR+A0UsU2YC9WcMnuCbXCr4BW/v/8H
lqur68Ppsc++vmonF8X/ni7dlnI1HmCkpUL44NLxkU5aQp1S08dwl6o0Ns3uHsmLQvqei2oeTP/r
azSwEXjwUK6YpAPUtWaFCQyBEp9oENnyh0lYEb2s6eJMy0awOyfqdMSBwDQt8vc7lGsrvNIxl6Om
zGbvayrynIt4hLJzwI8nU3uv+SsG+Wgfm9wBBfm6cpnc2GcTHV9pOMPLR31X9d0gV9tHUoan8k7H
trE2LI8mBnpHDokdIPH3JgGujZnem1oh7UKpNBXSAow+5+44ObBzW5gpLwQhGdSEjnYH7iWI582M
dmD6fCj+i7m60Y87NTKsW0+6Iz6Vj815T6zQ6y8JLBjmpk+yA+4gD0e/aneaDnh5ZAObPqO9cH1g
WI2Z8GLN75iXQkuk9FmpwUIyABVcig21/vAbxDoJBbcGiBi6wyK3XkT9Xr/TKXI1S+GV1DRoTn5K
MLm2rSOw6sXKc//1GKk2RXutFTmAN8WbKnWYxc7MYr9KWnnrMPuPolni7llQi8oexOeu9nkFpucg
pTN32wY2TUynzbIRGZbouLJYjc8OB1NUcm63p2+xSX+7BACadES8tCpup0IAIIsqN0zBnKqRPPBJ
DqSZqaV/m9gbFcH1Yzkwk0KNTyRkV9REKTD/AolJZElj1bgFDcnfZ0HR/xnzQt+/2DcLVq4hpu2K
5olIcaOcUkWBSPiamx6soAjMlsrEsclA/e85zTy8Oxy64pg086+eWyClfzGfgg8XsEG9ToHvJlzN
mg/vnAwOf39+ZwWxrEuu7KAoYetVIJIoXBbCzloij27Cqa1zCHLRCZEfxzqh1qMjtWrtyTZ7ws43
7mCyOUrvJVdl2njHT2rzk3RMIO7JShGqhfnLM0QkVdDBU9+w6MWhx8XylJgzdaQXapNnfnhF4XyE
ypf4m02/dC0QedeO9p0y5cEefpILAzqm4gvnpHMfuXgqrdX/jRI0HtqG9J2wXZDhPzVcGPd+leyJ
ag601jw4yALIhFrqNiXcmxDmplXGo82WBLwfAVEhg3BnB9bagi3tlwLKG6jwQolT/6DYkPt9ArHz
KGWYzPFjmKcpphXUgpVG4v0nisTCG5mMm7TTxkH3ceRiaSP1VywhdicEBO8RVhhRkVNNo1QQdJqo
H2hYIu/4jr4NQ1dk20oGU62bkZ6Ta35R443ONjE8pixHlynxModZ2DtIQa0pZsor7zqe7g6/RaOL
OglE/Yq+AGpqo2K+/CN8YjWmpI0KdParJe9sDKkTqLf7q4DUE6JCQqqwQlZoOMcMXitsiRsWLOAG
rkq76PqVhyPjKGLmUnsXUKVLZJE/Uwaq63OXI/TGZw2KIEOvxGZMy3RCUMpAYpqohO5exXNOz5Y9
kmf0CTZZWcV6MMFpqywm1VRlVOjKDfXvjJ3Wk9dmmXVRR0u/X/8V9hPrlryKecAfJ3PG7jz83qE1
jw2btqmmiynFjwwMDcq2ZmTUv5fY5cP67SYZfRDH/rwYKCCgffN+GDa5/VoMn01pKxH3AHJXXoqv
stQi4Zwu1mWn2giLzIplukz1hsb4sWwqb7ANdXO/DVdG5orLBf6ArInujCA/e0zgGHetkYOe6pmH
ye0zKGTzZqtrq4ZKshoFDhOPsS4TJkRi8WrwcbN5zTeOf/bAbO42ddtQCGLLStKyR4mjMzv7N1pQ
6W1ZXL2ethzG9uMsoLr1EqnOhutOKjnHbAUtdp3F/G8d9tk0JaKmVXqpH3Wd6OdN+MMujRLfG34q
Yk5TUxVe9hHuKCY7HZSWrHiIXf88Nkx5GyMfJPdr29OJz5SvVYrhwxVziB4DJfXwJ3PlwV53jemc
cPlpez4RI73DF+ixIqLC0EYTrvwlks5856/TVneimYLwIuvOftb0VSsc+HMVseBJ46bmeNBVuooL
rHMvv9hgJz7sp1N+HO8FJQrOvgiwdOXwt4t0lIxm5NXuDAme4owZx96FCxORwyZWJsxp5j4+Ra9z
gPR61SqzqvprqM0hYpdAl0n5tyrfzLriG/ETW9tkSkZb5yksGczvuJNwjPH8Z3cE/2cb/xpQKFN7
ypMCUA0A6TlJYeDuQrd85iIq7+tBYWyo8UvErsHyLqpxKVMkzmnf5NgC5DaboIRHHaBf3YyEmPfz
9gjtqS+FruN5mBDNTEnr3gyyxM4gR3hYzY2vfmWmOrg+R+CqmG1v0jYZp/YSRdd0I8QssEeAdh5g
s0kkSLWCWt+GRfioDwclEiamVBtHD6mNdja8CpuyL7jYMGd7doihqGqiocv6ejFGR5B1uMz8GlMO
Hau8RWOnUuQyrz7JSNBvyQ7q8NSJLIOMjiUszOjiv6mF4i78Gp8LIPsxH7UTPcomFHgDKR1LFPMW
H6Vn31wprvipR0CCxcK8Y5fDWS+h/d/BLpmp2t7U3iyhdbZHvnFCtrbUUGrwh+Av3J/i5YABAsLK
bG/JC1GvjViOHpjoa6Pv+Qfr2EpAeRuAoqYIV8vuBvreFMBO8DTAfEhGJtXO9aX8w+6hSkmB6QYR
/OKOMnLp3vGN3XKo7oTfxiULwvqkc8h0Ajum8sh7A4y/KycwU4T4tUBLlwtZz8m2czXo7AeqI+zy
abxkqkb9qn/ji1SM22sbC3vfmvV8dVZXgcpH8jgPg0xOjACC6X1fgSD0/FZ/Jp0YxPoHEfvzqqwN
eerfiYhHXamx6Ps11AAUEkHDfr2cl1GDDM4noFddhN4da2lJ6gT6xBVdKJJcMFkRMFicW1KwOKWW
qLixPpd43l4KulEt2hCDrV7iSLz9zG9vp2caAl2F1/+s5jZL/+ES3RrT7o4w9cy96b7b0UCGf/Sf
BqD6ap8uOEJQTTrJXEu4sflQQljbfDx+j6yuWctNt3U3zrKGqLlh9F60Dq7X4SNQdagx5QZl5ll+
nu1kZEt3EYY4vtsjrj6k2fy+a7ZglKFHkO4qoVVHtr/2o6munJu5/4p1q6CFWGTttovROjS5bQ5B
YyaWXv6D9Wvqa4icp48NXPA6dpgF2eGdx8ibQ0o01mbnK/I9h3/Y4gPsjLT+4wXOdNM9Y/EBrKFZ
pQUcAjxB/tDLV36APC5Kq/KDNkhKkCpzchjPC3spJyzS6efsgkrvkhKv+9jA1jXNmODg4fSRZdtf
SJ2Nj1I97ddWgmusYF/ZRGGziEubNtXQ/TLq8KPD5OHcMRGL+PyS4/NcJBl46FHpnxHcjqvW9brv
Uwmmmb9DJybIjzjHdiqttHYfdhsJgBzb8UkwCmq0GbgkSQY0R65iGDmyTKCj0VrOElANeCadZ0zG
2I2ZhS//HuDxdaDyG5yKXwW7xYRHaIAzGt0tzJYAgEiDbOvRn2Ese0VOjlAoOseQ0hXS8VWPmNqT
mGES5CiY7Zjl8AXVdcrUPxZz/H5Nwqg5FwvCULNidJk4bhTC6hsPA1PBnhtwmjeoQCpy37Wba+94
RFUVlMlH/cL/5Cxt/voBwqxT+0Mno4KyzPR65KzorFJT4OY6SQh7ITymBpn0ArpiHJG0uxZcrf22
0pDjgXiew38Kk0uBGmGc2eX8xQUiFzMuYk2jDy9z9l0j+M0j6pi4fxjwcgUpRes7U2lJpex80K0V
f95odZA7M0cnfbQpOhP5kFBlQAwxEGLYqN6XX/W3vBWLv50zGkqtBKZuWDrlnBICz9e2rLyIsaD2
9mroGQAc4yD3qYs8hHGAWs4uIqsNoXpraVSDK4MuXsvys5U0b0wdMYafABsTOVok1zp0j43rI4PX
6cbPDWDLPxrySSmpx4oIOh7noc3fhNSnf1EPU+kfMm8DI7tn6RjEzW+3LhHmM9Oxjb1433qrjafS
YkPjJidtSSfjRujJ/qIs2S3B9lzVbF0R3zzyrN5yBNxF/KdeN5RZlFjhS+gENFA38JfbreMnneSs
Mp6SnGIbJnH9lA7b7SMX7I5qhcQKquPRv/IWcemE4iWw92ycqK7N635P9kGcqyAZgkqChwOnic3t
DnTkEtsjLhHzgPtIT1vpQrQ+ug99PS0Km4CKe2Uk9BF2Rxhn9G7whCT+2if3EB8NkX8zAfZ8JrYD
FdQGz6XGkg1zdwNGuvPcdxvnDp3TZ+vu1I6PFPLj4MtuJJKHavvNC/mVS9A/gPfiilWhF5gCghBp
9umFrkpnHavTpVkXXrG+RnTMp3d5kDysJRcjpjdYCSUSb3EDwbtkmDW1b9VMAmOLO202dJjEWTgf
nznUdcLOyg6J/xrMYthKkhakmDkhXpTd28Kze8S4yy4si20Mmc+noNdfzAKSJdWOMHm00hGZW+wQ
pWYdt7jKGdXEDVyV/PFa1FJi6m1PHT6gJ1NVKwRgdOVoYlZeTsgqOSF8if0GxJ5qQ56hza1o+yzu
5astsip+WCV/U1UDLbfcSAqwy45KrYbvqoicfq0+/vAW86k5fAlFvWtoZ0xj9SQTOHElL4ig++vn
dB/GHI2IQmeagwgrSFbFcKUpu1p3o/M2vlr0baeNG/vbTkNgiJa9Q+IZAslzlWmhofp1teVec9pc
bSqlDMRDTw2WkVd4AwtZ4QFnM7CR5Od+KiEgh4NjxeSb+O7bLmFd6zbNuanurT3pw9plLMquVUyu
SzW3K+KTvulLqpOp8fxOIyX5KhMVXuVff7H/YF7Rj/54cP+Etp+eeoh0QMVv3M9gbNoPYkFh31gd
JMfdZib/Tp9WtQefNQVasPAa1SkKhWqL5HfzZ6epCKs6Qa68ZZxIRuzDW53qcFJAsF4x6MQVbetC
p25gExPJOuDpyDY3A4P6zHSzmgHiVNj4dHDmTRHKo9VsGzc9NPQTZr/ivVBw7ztf19onfzqa+G3b
+TI+6BaVoPELQitFF9E4qBjk7UcpQS34gxqe2W9eQ3zqBdzL9PmCkuXRrx8BEcV363/LNUmVHpCC
SvPHj5NT5nnzotpVYprjGOli1czelRL4+BedRjks2BKC2LHHmp3HdvsbcPm1J7+vG3omrkWtoNis
NebHWyYqgy1TgcGu7KfqJxunYHOzUgjncktlisLpHRmdFXpRVjOC7XqQMWrtX1LDg8SUsGjpNIAb
wn2arsAW3cEOqDXaQV8hCDKUcbQEc16jd9byP7kM7JmjLhQ9ijJKhhNH+4yUoqb4r0psPUOb8ig4
DGztFMckI0No4tVPcGuiSxluJ0BxLFoQMCBgu/GNqBgIpZ5ibB0xNqON7LRICBSi2jzavFbNGz4e
0t7mcHDiDyVgGrVIIFA/p1dXrT5yARJVVfByU606uoENemVfqwLII/OcXPNkRuTYbh78bTmxNzxy
hCdHCQmeaUl+r7U/ngsZM+29jdLLHs5LUhv3QIsmJ9/LwDGXldZJdTyPqkluv5yCzaQPmHO0ppKg
HFTyNq/MSxI++8jfUTtwhrE5fvQQcneFmJyPH8XHP2IStOTg2qnay79lE0QDxgL18l6P3E0v/TvO
3VdvuWs77zolZCSsDH8Cn9uXdexI/NC6rjDMMnHbREdD8gP2kksGxiMXuK4MhbQ2HSHkJ8YF5CQ1
t4mZdLDdizPgv9xK83eav4Gwim6917zem2C1hWIn4ivFfQEx0zs2AVZqqH96ewADoWOhefTWIVin
UYQnTSxJD2UpNuv0mqWdE0saf0iODZsDF83JljTuX00M8FTA3QEj3onuWiWKJdVUAOzfmmWZrPI6
7Q92YDOWPos7AVQrWdDbUn6tXjUOiVgtC2OCllJ73eG1QCspSdNpksoHZClM74XVBi9drH3MKH8+
0BvlHaw3/i2YzsWqelcCFoFi8kM+F83gw5ZJH8OzC93mK0SdNC6GTMzIhiBaiah4IZtiNLUQQ1dR
OYbMlLBV7Bx1B65OXNFVSVF/FPBaBmThLwtdxKQLGl9c8ZlcTnxSaXsK+XZzI3kppt0uWYZ6RDHn
U0IvIfRqyTsS/M1SYHaqay9biehA26PYjQ9km5Poa5wa1Ca8B8yza08FX+g+Wf55ncwEby5ksHoj
EDiCiC0QxtLiEmx0mW6a+j/+/o9N5YYXl+psJC0vJSRbroDSpm70Bqf5eF2833XCGQ7bTty3Zlba
/nTnxOUgU6eO+rZLSUmV+FX6ok7CekBCS8fUm1K6IjOP8lQePuderon7UJYJhygllFpTJPALqWna
juVd+pVeSOPS+4IUep57HJslGqOknZ/6rXFUGDPICic+qomlJ75z12uVssL+0oWv3TLstxlhaO8D
ZQq8mErUKg43AKFcOlqtrORatgtIDOyhFIxQzV6Rp7aa5L77d471E8V5Hc0cg7IKIgcgm2ix/DXF
P3tmp1PZEv750A2QMEMLoDMN2WHTu03jzUl90ZoTxtIwfGbhGHdWHq8gO2xTCe2fB/0N8y8d9/km
YMxSjldzPFwomQ0gQaxpFnB+Oa1nXVCJ4Yj01hrhurSZ9jYN/rUCdz9yUzK2wNuvbON8mrBU7P/q
Ne8bBNr1YptZh0LlWgkccilHM3lpHOYDDOJvXEBQm3fN0QbWAyTFknwpFuI+sBZnl/03V1XrBKnY
Qm5SiBG+1m1seV1vIeRzIv6z2aOc/ZY6Oz7Ys2VjAU3FUrFt8NySkCQMnkwN82OhW59dYHOdj7ye
oBfzQ2N68Sumy4gA43yxNBnCCcUBgwT6OtIJ0dchU1A9Z0Nr+t++t5FQ5OYO5RiFe0rrtpJbL43M
lVyD5/7p6wuEe6+4JDY67Q+YSZAxq5eMUlwldfq25g20xvj1rPXH3yRwe7DQ8J7VYZagGjx4xp5r
15uju3xptgnTZLevZFlGMhjY8yTH8DFJ4OWBNt+JUbkxLiLlIEoWs3OgYT+aTVY/tewHLAocx6xA
bxmoGrTjD3PO1+137w3SO+3YzIe698WtbIrndDciGhxqa4Dk8861dyGy8ne755dauEkG6SZzU62e
suD7XY2mqoFDJZycqTb6kVx6b4+tHD/Y8FVUJMddn5R5tjFhqHYhADPaVtmF3AB8bwpkBTWc+iGv
F5kGvidB+ujceUhOt4LQXjxoYxDMTeOZ1c3xaR3bJ7ZGT+Do5azisw9AwOaeCK+ZhJXcTE7gJFL/
dUKeEPItu6+Y9IpreY+xxAQwkYHv7vW8Gn1y2a9baqfwnLqitVNuqLBGhmEVv66ybCIAEDsXj3uU
I9XIzDzQQl7j5SqcQa0cPHOmdmr6l0EwmD1knT2Ob49//+ZCJzcRt+z49xPcl2eUHYw/frqebpfR
o5YJjgGzgDaDeJfU2dWGaBmAjg798JE0PHk2DzZrRLbAJfypyRe46VJAj6oQnUsLgYvfW9h/pkjK
+PFrnHpEBYQG4FYjuChs10yPT+Nx67ZqOOLMzrRx8oPBCOXlhHSYqdQhX7aSKuRj3ScIC3uTOtxU
vhzyN2unzuSTvcEcoZXoEUoBZHRm3H9im4cJJg+duMmn5TexaHOQFXxjyhNHgrCVc8wjbowSB4Le
26LkqX0nVWyyEh5pycKMzEHTMOFVpu6GzeFidddWTDDGY+CNxKYjPKxkdbnksi4VbVlp0urFqdE9
cfghkm+IcdmFtxkDPD5bhqdDWr/rH5LvTWrypYdcF+r1JNTMPQwYEJZYCrEDncmJNXUahB+OjlhO
/ONayG/DrEVemoWEfsWtzd4OBXyAVJjXa/4+Zfbx/yDqV9aMDbemp4FkwRM19SJaLiXzcLK1GYg+
RMZlGCwPnoKZm5ExpFKFkyyOwgxHJFkns96kajbh4JU46Q5y9I0lJFJpDb29qdK6Rc+eTr819QzE
pwK6abw8/aQS9xglB8WAMbZlxO/NnWSkUpgNngYGlJDL0kCT1HH/xKTV/e4rKhHqn/P3fBLlcG/1
xxKPTj78CtmJvB5gMd6u/LEWc1oqqXurZlXiK12flHO3WqnCR+76ZkTWZZk5BbxQgt2iF2wJuxCF
bJWOLkDj0b81DAD8hek9UYVlZQARiJ4yJvqlDhuJvIipSl9PlsIieRoNHh6Kor3mbxgmItDj9uS5
/j8/iI21LArWCkrwy/0nxNkEdax/8UuBsoVIrpnDxRtRJd2lcEc/xX+bbbq00htBQLnlvQ4jRwpu
B3ZOkdTtsC0NVpNf06GAmmtUFQVGjdqb+dC/KUODoTT1kQuEiK60ULz5dClsSdGZ01xCADqDKXVL
+X5IVw2dFSzh0MV0Cg+JN1KN7SpLUhvCS803qoiDUzPOnSP9LRgeMA8s15raV8emg95iEHMSSsZH
e6YlCL6hWg/F+JryOIKUKjmVXbRusn/mJ6mCze2yDuWTslkc+MzuGJA5kwnzELTmM7HkICxRHI7F
W7A89zlLR/KXMMtj8FZx2wn/W/WJq/ZfuTpVSBxLLdwwtU6YHKRQceQWWQc7BRVkt9l40qd2nbQJ
YmEnsFpaTphuTmfyHwDAtKHb5C38uxxFfvlEsCK6b/BQ/8LRJeY/oSfEYUpOhWX2pXrgZc0rSCuW
eijZL1lJUijtqdKQXS6Xqy3XbtUkE06JqqR/X5ofkon8m82GHY7OP+qV+LSP/YwPdZaLhQO6wVgK
V1cTXl72L7XDWDYEjkRojETb93Ey+8hQsv5c6CxttVu+2zhYIFnzAchQknoXCM3JcwhBgjXxMyxZ
9hTL0VE3nqqhGtvrGKrskaxXcsObH2OBLfUMM+O6kw9bLRXaft2TxztsoCq/6krW15AJnurpvGtj
R+Knp76XSInuLi05u4FEogHXBtvpQCVxvjh2Dpd3wJOBqIRSgiyY0wNPaCqT5jY/+7r/StUmLnOZ
tAhEeRKEaUbU7T/gpDZDomyiV2oQMQ/mRO+WJSnwz5mLcHQQ6zwmciPmldIHKZQrUjNhYVHMGpMV
43VhiPt0ViSWU7khby6rlkdxN5LWXle+7CqJhyYLNTFhCytLfLFiv8tA137fXhOrd8gNXQXWtvzo
l3ZNFuk9MxCyd5vbE/0UubbEDDX7D8MRT4/ZT/c2jGyOFx4Zo9rXNMzR7Bfspbv2vxqZVZxg0m/o
I32GHRsLGVHIuaRnfmeIcirpcuEh0mmaGRRLrJo2YmIk8FLsgEsLNL/mMbJhwPPHeqGVpnXT7e3d
A7x3YEY6daVtSGNI34XU21xe+idZR/orBxxqul/k4Q4Ki8QZQGNtXhwK5kFzC/Qtefn/+DOxqSrk
BCoAK5/4gNaahSamyYki1M5M3ZddJRbc6p9QnhmzIL0dlTyJuCAiaGvAi+xIdWh5TKYo1e7xbr4A
IGCdwMzORkz9gAwys0t1lNpGZfbl6jYsWL7H75Nu/I6nTR9G00yneV6B+vxw0vl25J6tWmExDlS0
16j8MgtJsib3T0GI8mwWyvGwKn7toh2A6HK8uOdvtdIkaGoMYhRiv8zEAi84bE52kM6oCeIHaJmw
dS+Yh6a9AOp70bwAvZdWDeBM9xhetycdK/ddkCdMU/s9/mydCtWvgWQ4f/Ht1LBTaCA6IR6r9wi+
u+QuCmeCFNsO+DB6Q44EnI9EdngrXxXvjalEQ2aCZdyrOvwjvaaX1lWSPJZMVwz6S/eAEUJg8GPV
1W/rFI2XaGbnSBdDywDmobd3gA720PvC97uGFWRvE6QOxf0jlluUHbHdp0F0B1hmfMMqL9r7cUaB
ctinQOgz/uU2Vt1TiODRyCr9BkPmTgdP4EQnT8BPohHhX7S4OyLzkQmbqMLc7VgEJZQ81gJRzzan
y2I1oAZGE2DuFwFPVdtpkSSJV6HVwA12k9AEXMxNOXPRfgYv+6piRiwRCB1rnEonGG25ER3vubNe
bJttIEhZut+bYWDQH3XUxprlbY+YSsIaPOqIoPBpZuVci4Lyyg2FyRzoZ7CRCPk9ncTD49VmYWuG
d5BIUzaB8KoxsRBrpbmWpVTCS3hyb/fp4RsTZELHctGizw9FGFeH3D5GhmBD44KDtFLESoNkEG55
y78G3pAqVzqOoR5NW/2yYBKiLFXsd6iF2LzwBIPAwVHETJVDBnExeHjOH2idmekygXhdoPAe6Ysc
6fYeLkqF7GfHuAqoPWMsdILbFI+qPkt+4qcJrLHA0bi25qQOo1NOtZb4kh/dZeiWguIsnBMxjRQ0
w8tloGm25UDDMs3Ci7E9tftxtktCpwLMyhG39DmjhLaY0Qmhqlo1TI2bsWdZwP8KkQ1C8+HCW+Sr
ARw5++Lj80+EhaL7yAR2Zy9eyz+9u65QvhOMwe9G+tkeTwpxFjWHzlsBtBFMa6n7D0RH/G3SFX6z
u9SKCRJPHIvXMSZghckfNDzdERG3BbBEYLXlUoSER15JfmCpth7Z/bdq6lWwPPsbwOj4i9jrRaNs
KI9JDmjI30kiyHsIcAaobgHxyCrLmu7NldlTPIM0rNpDs5MhPr5FeVGUQXfWPigPxMswiH1AqDnS
WuWq3velS8UvJZ8k/achPkK0y4grszwE+xAsbp3fEk0LkevE0XLdJsv3pZdweyKGyesLe+/p0/EQ
CpkJfcFe74jlBkCtjM4n771MldVSRNf5KsJa+ba493keUPG/bjmKuZ8PezP+sdO7VE1urGkItz5V
PacFnHz0XnkkHBFLUOJn2egCutYDL1r2m8JYSrTihJjr6HUYCEMunlr5icbj8TszQ+zt2vnUmfz5
0factIw2KVXugFriQk40Oze/rSbB+L/ya3qKVb/51CUr2O9Shimh/S6qP+vHeBAEg2gRrl1pl1mX
mSQz6Vdo5kdwm9uTnQWVN+B5fLP4QnxRMooMFH9txTWzo8kSEShu7Dnvb81oBK+c9C/y7Yfa3hQh
yo0gX2HNYq9N0ntEsSltXxyRPi+yeDMHKikq6PjyQA9yjsaPCjjFI8bx0Z/qZOqZYx8rZTRhbUoO
clN5njKVbXu8knYfkqUiALUcQS2DsLMvy8/Etnc9NAkcDq8H4PpsIpl2xk9aB97jd/9Ld4BVZMW0
3Rbtnq6WlCj356ZYahl6M1pOEFJT0IMfIYhW4gIKp0ZE57J/eItxCTmlDFZ4g/n30ERB3D0f5GlZ
S6jiTQ44k1CdI/8wqOAKjbh2ZWwoOQB6rgbf0O4DjvZVkvZ7rmtOb9y3eZDsyiv1f1/otSgIDr4y
JWorsLiqY03PSS2hQD97Pumf58WmQ07TZH1/jz+kUBBQf6FpiOcVsNK39I5PCHRfS+6ho6N23xWi
mpfsKtHd+MyEh1uEhuSDQ/6Q9pZVXVdX1/vNy3OJjZB7CFQ+dFIgzsGxmrJwysrAuUHFuzj9Vz6R
nLD98RQdxsBb5KA7OwXY0xKCVm/pj1pcX2WBgnPfVVVFjXHhQhe8YvnmAu3zucVAoaxfppTAmf1i
4CFCWb/bfAW7fVGNiuWuzIQ0qzLfVCkMnCNLluWL6lbFlGJtM+enaGZxT6Lfm3pXwp20svPOVlW1
rxniaAruVmOze+x6ktvkdFsK40HtNWF8TzFg15j8vRGwwkhRJjn078D1gkz5R/+Bs7jAW4suiPiO
mJW6z0RyLPfeWHrMPDP+UmmZ3L1j9J7DQ3GzQtzkAFDrAxgiLU2Wya99mmDswf4YG9OuiKLLNvBX
NS0tDr2xOQ1U99KqnMBksQMBrsDY6NNWFlTc0nzj9Ufg5LR/X4hfftOdy2IVZFHS8DLKskpiXouP
2Mn5FxRWGgMJa1sUbdsdmH2JrPC5YotYlLo0FuA2zwqgsUG12AuEMJs3SYzd2ye0GS8TIevfJhuP
r+8v6C6Fa4AhgZvjAzIHbjZJQX/rMTBD+J+kFwPqKjhqy6igpKgbZoAZOUPn+9oMG5DzLQligDJh
AekG1YehnGBpzRgYsRqGeZJeMCNW9kcbeS7IjC4dLsUWOyDLEok8HI4IU30dAdRvZsqI1yGz71cv
gbZQDt+FFVP1rWU02Er08t1FTnsbXd/mkZsGfdRqlGYlYRbD2pAhdHZm1hnBniF4iyoSs66r4ZWQ
W0OBeWWpG3AR6huQCBfTYeEOTspO8PS/TNcfneJx3bHAKE9vlzjx7OIcG3+WfakzwvuURRVuHwh5
GX0FjP37oDd+QP6T9www4pjdU0H6COCD9nXPnxWxQlx+KPa6o8fTSf4QTCaXMOUw0BcOuOzOTg5i
eALCmthno9z14gM/+CfRuscdsL5BtF6oWtnvuOTJaRRbwvuqKfVc0aLpJNxZsqGUgIrLFjCFcvWb
HaWdO0iXt/yuTIBBNFSEY8gHXqubdn/XgKqRi++vfb4GrAAa+drJl2LUX+3c0915zfXLajYfr77k
o+7Kr5KZcxqMhE/SnBF3n21qbl7QAvd5v2f9dbIEW9FX3N6G3FHSgJmjs8GLPNPfHX95LCPh5ys1
p0jswfEr1adFPxT1GtgRR1gPFemzm5uE+MUY+8Q7+bBZS9q4W4eG8gFki5XvAM9Dbd09qR3hggK9
WP0tguzVHqJAk+9X4R2y+IApvqnrSWz1H0pWBEbngEOs40UhZPVPa/AxqsVrwdmdFGlOz+GeHyx9
fzbkf+9heBiSXp1FNXY5Pi8KDtibr6FQJKZmeouIr0tCMt0UkIdERiAQ1rM2YmzBFaSIraouFbxz
wwnrynkXn6IpJq+Ua1p3SSMajTliU2TPZdSVYiUB1NrnT3s0dkqehC8S1MnlttBFB4KpNZP1sDj5
QvfdEkb5lVR2bz3nxr4eO5D1+zj/bImEZbmZnKDZ7AlFeCSODhdjJ88GgniT8G8MoYrziQ3+WwjQ
9H5lSIDGV7dGREwF035PY1HK5WfQSdfzsEsGlkwZ6JXeFgkMs3gh+Eszb80+7c6tPZ3aI5R+pcW4
vY1BBYweXuIzR1wRjcMpPcA+H9gMfA435VpSUpcMtnGGn0X334ZAPM7DY8s8nWI7IVdJ68rMUhoR
jX65W6Tg9NcL3L2RHjNilWxkrsFykkdaH6gl/+KIRAJMfHSpf3/bROhXeoJs5uE7c+yXfyrQdw0p
AzjJ3TJDit2MK7A/w6bUE9PCsetnwhl/jf3JSACouhZ8CS+ypSCjMy20DxD6r/u9mzQ50e0PXAWX
ilxOrDXNacQDossVDF3Pf4YW9h9irbgTWEN/6pN7v+Ucx6gFkXxfz+kq2a+QWI+gTmDYY4GY+prI
0msQjt4LSHzOJwPAqV30i1QePkdPachsgtHxkUU7ZJ/QQa/6wZwom8Ux06v6pLAVEcammwcBzzjY
6rzib7YpUsfvK33xgDINnnrTOHidC2d85CPexW2ixQzUY+AmuJWbpBNesurAZEwruj0C5gPouN+a
pxD4uw2pbw/QJ+t/RoiNvEE31pVXpnSQcx889L2ndNzJvB8WUrJd5amRJz+kzDjvAAqbkL2rD2bo
3xTLBZbTcat6NP3FTfG1BGD4BdGZQmLjeO4gv2Dys7w5UqEt8rglswbhyjTGeQH43S+B14a6Zn4Q
Sqz32U481NetSZvki9IdxOZKfHYC/LF/Y9Bp1whnTTyalq8zqE0mfPFb/HE6bF4Vrf3tyJBng5cH
WLWQoYdCXAq/HxRMkpT99Eh73zk+RelHiZN2OTTkg8pIpYJZmS42MsE2Q3/XKMX2Frk7xUimQI0F
dfqzhz0lzE9q8BdSgXURwmBhZ8LjN5gzVeymb5gxYfmJICZRChcQp8qekL/lVyt2eMpXbVmqmfhw
EaDSHERnR2C0Bw72zTjzH7lPHqpYnYTND3IwMHzU5ocSr4S2YpiLxyEcg9X3YQSkZd/ygRTYZTe2
hComv4rEhGjTCEGhs9jmC6Vb7r2hk7GlynZ51khg//AiJjeJ0GH3iENORF60h1Ov5FzFsQJb67rR
3TxXhYlRiV5cbJaP2e3X7NhHPwkw1dFJpNayF3Eq4rUPBJ2j9fdLMv5Dw4dfKKi8tlJBtLsY0whJ
cGGcFkiNmjEVNmK9FHidpcNZ5981+LvMfskvCmChFDQob5qnDa585zHBozc/WMUtFkSswMg4Pkzi
meuxP0QQXoTabeHfBObrar3tltc0PzA34ZWRmQXsLdzl1A+k2jcp9pQYyTwfwRqfyl7JFxynG2KO
qPDPP9G1AaFRmiIRLK+rC9bVLhpKF4PYEKd0fI8PphBpCzCocs14J5tVZq51KDflieTseXHndGT6
YRqwZ7Y65GLpF6TwtO2kCc0XKPrkfBPKkLeHqdx1GaMpgLcfxLMIG8DWhLGFSoiJ3fyunEVM+YMq
Rw+yB4iJDVjaGC6mEp33dDNZxxTg8VnyOd0phc2+wvEUe0/d40smI1pYUbMdt65AG4QmLqLYlpIs
BeIC1c4sRjOPev8VUlb4D5aPaIoQ1Cyhf+kL753HngNGOsyRLf2lYlrnJqNtEecKFecNRiMb1ehC
TTEtcqrcw3YEB9O4E2O0vLHW9xApHmqV713sJx3XclQ4sb+A+61pgxd/ThP+szgFhA0BrrkeuuNI
0RTZ4kSAnarVYNUzKlnwp9jDZRosV6dH6j3r4iI6+U27ZLDyuFB0Y5alvDEYp6DISIlrywuOkOrh
ZOt6dG9oiJHJXaPWbDTlhJ48cUAqfFgitNJ1Rqp0nKz+gFa8NbDfl5GvEBwM/+qIPn8VFLFTIgdh
FhbgOVa88Lu0uFhX8IE4yuw6LG0Mn0+ppzwuNjn5fWEq0r1blT274c0XeVAe/q1353GZum/OxrN9
miX5UMnyV7Nq25e+kV/HUuUfFmVexQwIgAH6cJBC+tgYHKu/Sl6gRPL4lhn+rJyFXhzNi7Q5yJug
3e3nYC8ZgSyTylRF0eLodE2FsMk4bRXI06Q5MpbA1U7C35LOGJNHhvJ2/cxoeuc+FEZ49qWM8HsV
VEUy5AA3Pxyk+L6CZ5n9urWZskXXyL1vTZ2Xhw05g+DfHr1URnwHBA3wWbF3NrxRKcM6y7yVipXH
h3ahuuASIs0c+vuTs3b3FZeDc1/+QZOBsVoGzc2hro+pd58MnTr4LMHLmGNERDZvweQ6PoOrZ715
+Q23kdvg49ju0/YcvuAhlhwplGSrIDghaEjmTc0i4R7e5KAotK7k0jZdkTK4zLLOjv9Vu2P8PSHC
vYS87v1kfoYLcSGS+ZfEUKClvIyEbQ3eDEBNwP0Bc9Rh3ZTvs/Rfkxg9iaMiA8qpC3XOgLSNyP5p
BZh2Lwt0zGUP4nl5PXw0RK7njj0q9jnHspuQypgHwgOlvfS3Dmmiuf8Ugkfix6sU+Kq96lagnPsh
1STpKIlAykQfNVRRDFVtBlzfxmsZFqaO/1RlOoc1XFDgllrYmw4/zM06+LMZhPK7uB+v0Z+fFwz0
Syemysvr3WgtLXyCEY1oLPuRy73TBLq1djcJmNKVstx6i3KPwVbSgWWr1QArXjEcJnhmSxH3k5c0
2heedg8BxxVUrFuwx/R+zLTuh4KKvSYJ2chyCjwllsn2no4CqjmWC+0dqITxdgjRRARL4EEDAHUt
quM4d/UuifBciiZDNuhc2oQ58fGgpEHfI6KifhS6v4hlb69nqZqfDAaHSasi/odI+pfDUDBsopPq
MFiwRispCy20/0eRKm9Lev5BMiDyknkfN8i33E0Vlgtvqcl/Xqs39zkxWsZ35Nc3DOKpN/0ncCIN
rKoAh0aR+kehaJ46Yrm3SGGX5kn64z2lOtqlhiouA3UkEVc2UBy6NJV7Rovm3/3pqjFcp7xpSvp8
ghdvEIS+5MT60+epUbyB7GeJBxtEvZAFEmKD3/va6x3dQAkQLwKepn7Mi3v5Q0H0X8d/39CGkC/G
UCY+D0mG0+e0y+5Tx1/NwkL9yy6j49/6IjcyhPrILMFm7Yn8riYZTmgvg+sxNxtNCgr2IeOUhKmy
TiLzJP+0IrFR/l9pNw+H08rULcwhoJVMrwGdgT71IN5wbw/RbW0hxEELfgu7y0wyzIwJvFucW9Mq
/WRw2/q0P8v/nXAWY6Hfj5WZjGfd4usYUltGEGtuAf78bwcXwPN0EWH4W1q1n/Yl+iWR1YA2mnrn
Xqpb3IfnL4gniGOP+0xLO80RjlWGc+pL9e97yTLvNjAvdL8M6lErygJknQpPrkDnBUqGtOEemGkA
TYZVFlx3NJJj+KMWx7+fEhibQxIrea/y8OAX0Cf6lxF4rhZQE8ZWhr3TFMo4719FRaYnCJ9oLu+O
bcCXYAMyGZ4vywBIZR4UXkj3UzY9Zee4Osf8i5GyChiBWMGGJFia0Ad44+4maxrp/9ynI+/vAqhY
gCyQ+aLseSNRQBzN+lYW+yqvJULjBD/Bg/vKK56W4Ejb99rFj0yrYdMOTh/DiWk7UnWMUqtrdE6Q
XPTnecinnEwDNcfhny0C0VT2/DnbG7f8yupE4RXwRGGF0G+K02Db7c10fU7OkzDwNF1g2OYjrteP
OhHlI4a8X9ntWfcq3aq0R8foIOsZ7UOKvCTR3VGrnGdIVKtsst1ec9uqKJreyBbR9dbCmL1dgFq7
JZ8m+6oOXNluH/QuBOHj64GoAqRWPgKBDMZW3cAQguA/un06zQXoBH+wwiUT1+wv99z9kZU63sPg
ByDhutgSll/wnYgb9DcTu66uXYq/CSgSBJgVH4xDRZwX/zOpj1PUF6zhr9S3gifOQVFoYMZOHfXz
+kZa5PgQbhAlTR0+6cP5J797oLLh5PK9W9Mita48oVoNsksAOw0LHUqjbO9Pou2QNxxkxrbdthgW
oNfxmPjZBqrI6Vr08vZ2qXoiC5zT5Tf+x5VwmFLb/mitOw1zkviXg2EWW/yXYVvFhCJnCC2yveC6
Uz5I13g9b4k20qoEL/3zQu4uG/dhw//zFhTIgznGMQu9mNbVP6KymCt8X7IOkEkyP4lJisET31tT
7Dw9IJ8SDzFrJinjMC86gyqFBwnIvYniVJg7Ahi8dwoqh8QkAupMcb5nQIQPikDvDKbKD8SGQll3
shdZ8Ye3UY6EorvEQyqqgZJsgUKaxsk9bNKIcDwH4K3mWCUP4TC9WVYo76SawNfwulOMbvnIjUD+
8SGQXfe6os9hdkvpL3BCp3kzrPLdaKHnvQLlVRGiydHlvE4x/X9rjGI1hWxs4PklywnKZ28+qTjM
DV2zQXoBEYmUQz2ybxDX8y+QVT/oR8I1iTcj+2io5fUYJDieTaWywm8io2yD3GVeGzNOdyzqfaGD
Kcy14+TBXZ6SpDQ4crPxcspZbdeSp+bW+/Fb7pAPSuzq2OSeuxCUTWaykqOpOeR3zSsqM0IB82sU
QtFFS+A8qFPK0pZqlmE85iC+GRNmF8mhaJY6U3numIqIDppHv2uAI4ZV3j2x8kUWzsnRnYkfNJzs
xUaUprALrNlf/pQyEyd1Ouv69eszOmk6iESxNujHaucktBBOJcoPVQkCjfNwcGIybRzyaANMVrv7
efLEORQ+0bjnoKnemVIwTO578qtl5kXhXrlqgZuEktIPs0DaEzGvEdHILE+cojgcGaVqUBnwnERF
PC/Jj5BtNjcwWMZai2wtSK+aym0w4JL3cwHypPFqz8Njt5bifPVG8fMGwJvmQ9tdLveYn0gb9pZd
lX+uaiFOhRkKffCKCIa+Am1G4/uNcOLyNbaVXSDbcCFHAQvzqLrgX5Ej+JPZBu8Nd/i3DVWXGXju
OhgR+8XVBPHCKzzNcY4KZQ36pOPCMfb/SNxG9zkZMGcvwRxlqlJa+bERfM3R4X4M1SycrQRTA9fP
em7AlSUcIAJdvK9b8/2bJvsQvoMv2fnx+VmrPtziSpV1HJdgkVH2h4QCRvkPSEHnSCGZtfL9A8Ov
5KRng7Z8yK7TXgVFDN+oP7s5Aiqv9ExzIKr2pmG7xECrC02+IkXvfYLvvegFhuit5OdnzswoRjyb
e+hAL2noqrXqj5KEzk3e8ttZYzmgiUevw/0CjcnAas9BtEXLaJj3oIrtMUe9cLPIg2BxHUwifkEI
Sx2kkzb7N9ROFy0IdJvzrEQHwi/7QlhVe4oUVHbtcH9UsGQCwWA2co7zYGYU/7DseTlrf4rGkKQ8
kJspkhGV9IP9B6TLmzcmKsbO+S+UVFMWp8IAl1m5rhnloejbVO1u1+43S1OBIIJGYxgcCamNQZkh
Sou+L6VVW+2MlklN7zFEtLNPEvV9hVQm66KCtrbZEWdSboGZ4Zyv2eawOsvyPwOSj/NLhrndTrJX
z/p1A8v5j7lM/uCh26IZSQ2UuovRpAxcfZASUnOFR0S8bwYFV7RO7r0WZrvclhCbZszUkDtF3MFP
IOr01pwRGDhxb5+AAgXtC/zVp+XEqVTT/sL5FkAzXmq3ltV+e3h2g6bPzdOyF//i6HEZE+Jphcs2
LU1mseNrcJ3OCBvgl6QzyTQe9om8Y54YYF0eMmFZTqu8oymdPZq9vmoo65sdzNXoiPKC25lycYZO
t21YXQvId7/v4OWfjmLa37Sx2ahs5yGDx92bLSkN4HyaSDzjQGe0BxM7mGaU5UYymqg2ivrMKOlG
kvtZa47qeD5f9N0He11sh+tSue60ySnDMgh+wkXFTQhr2RilKzuoMHyfj5OlleaS05uARJzEJRa1
qTE/2ZuOIPHWgXPNdmRViwM+2Xi0gB82PkVR6ebt51pQlqxBdj7o2Xo3ma3E/rBqin9znbHDO7ys
KhDfROd1Ew3aMXl8xmc/cuVVQfsRQZWNU+L3y/YqSOnvbfjuuQusTCixIaox6wPNPVzEd3yKSz8W
XVTcZwOgyYnqUL4/HLWzKChfT3MhkuVf0Vq6XIJxDHDEHRR7P9o2GJoi4whskZmYqZnkx67eZ6un
ZQcdTxQYTs/UVLuWQ/jEu7xqpe0zPE06Zab8UflpH4A9nxmkQOtQvwVFCUjqmZ/l72NCSQ1OCzZ8
X58yHRf5j6Qo08RMvQEyRUXlX9Pqzc8GlvtuHNxIj8LafR/bylOaWsVDeSE475XyZDunZqNC7XBW
U8TCeKZN2glhRiHe8slxbQGaIkeP5W01YQU1bnKmBuN+Sr8Eg/xOgB7hTqCyulHI58SaxRauYjRo
WV5ShK9d+iYCjbvyih2VZolYTOp0XkGiTOqBhJNEGKEeSrdEM1IjOxkwM8Hwr7bugw/fHp6jaUpX
DlwyGdLK27BikWaxaH9ZbVK1e8EjH9lUXITcGisxAjtV6bUk+eyKv7cxvY4n/V+ElLE8BE+B9P0S
pLQMNWz+K3zCr9JrGkMjhxPwzqb6jSJs9smxcAS3ha87eoTBFo45VX15Bo8ILzwOLWLrXCQn4mwP
Ye/wQ1j/GRq61NGBtFiEgyzoy/j0J+UlghZtETTrhipimvHBkZYXimjfprREbem+2asApX4kzR3S
ZjZD/Ht8e7vn32U/8Y7jtYTbYKK4NyWc7TOmfZ+juq3qxoUvvQEqwUJLdDOr07jtar8+yqM3HxAQ
Bzj60PwB8P8W61QnZMM+9SpIgOks0d9oyfsJsUPmKUwL8btsGDDHsP9WCgCL5ZWq9tRwo+7Jym4B
JL74K54kjfhFkm73VBarxvnv0SB/y6C63G3veEfvqCMVvTG7GR/RUJDn+BCzmjRwg++V4vGHrpKZ
rNd8q1x2BdcZY91CL7KqFeIptCt4s8UIz//Rk/PVpVAUX/GVCjQeroCqmOSqfjrM+/052bgfny05
4mR72PjgUXzDAaDyK61z2yY4WkdTiqdTabmwpZ5ZOpooWbiEzHQbOc3ORTGdlmeRkb7JhwQhvgmJ
0ppzD4iXvW/yLJ2Rp6I2edpCng2CHN5fvUv8cD5051DpKAAw7stbDh+mpHxy74sMmPW8dqoV3ySe
j7YkqgK5usFb5xatj2H2MLsa+BP/tUgvHcspi250G62PRBSSjX6vm8vauIxMl4ZBlWlMCbDQbRpg
7g7WNXhFRsKHwkC2rpNNnLk9BMFyECH344XfGeoZOn0hBadfhpXML4bPG24K8lxzXJl11QEIs+lP
AuXhZzbe4FJvD99jcd0GSoUo9DbdOBybfUZ1P9v4R+51bXF9I1k3y9HxantGOruUKpxI5cmSFJoO
0ZFciGvyGHZCwBObCx3hxOmWX/LNWlThipa6x46EoEg02cRwMcAAg9+hD30kzppIQ/AoykFmV2nD
GvVXkvnMCdaIde9HXcIdvpxvHsNxmhjQlROkJ4qlYow/MF4XfBrbYvIhnvGWGA1T3lnKGkQHys2n
So4UGBTk0SwV+H5DoUDft79inCybzMCzCzMScl18zcvDQRsnYfEj9rXbtYOTsEx52qfR9W2YT2Oy
G855eCJyS2S+NAkSwpj5d9VowBohqBFj36QJkgBB60WHOwv6XSJzkhtZDpmpNgMnbLfZZoNr7zIf
BUF9AGDB4pBOBwQ2sybblO8xlG+pEWfvedjGx9geEUAr8yLooEIgPJh3JfG9gdycIg0INI/Q7eyN
7lTwBIoHqcsl1vVi1FI5oIOwVR+bH+Da2zIDu7pCow+uy1FP6IYJOmLVwyJr5x5jTQDLw21HKvtw
i3tSCgoVcMqfQCVIQj/Ag1Q6Q/MojZuCChJHIR1pN5zHRYDuG7+VWVXu/gfrgG9Jq3tmwXK8wBcm
DCFavSuNlCttzsEVTirZ7O9yZkFpUThj1wRX1jf6W9bGYKuzwBkcjHoDbY39Gh6Z6mQfxuqDMe8G
ZZpt6+jcmD2rRcC6vnIlKI8iGzG4+PADZKwLJyxO91cxvr/GlHal+Mu/3ex0D6/DNmXS9pnqcgEq
p5aqZbzIhhEhEtkyzFcz1+9FvN/MVY1aiECRu+mozbCS2TXEC7YdqBlrhyzf+OHjl5yJkoYWWxgs
wg9Oxof45YXslgjWl5HhJmsUxCQpmVz/q9qiqT9upLi40Jg0nip9RXqGYQOiYNm+jOfxn4ubvoO9
2ofB1fH528XvDsX8GgnIgffwwONbk3UKGgfVhMO7G4HKRUHRcoHDZOsA3HH0MbHZVD1s2lkS5hXL
wln70RNjlkYOAQE4rNV8je7f6N4lgeyXhxQ4M5yf2rG7To4G3TFm124aIKvqV8E1AdO2rKgP53xJ
k1ZFhl662OYUWMQ5iUIGMGgjZLDKOZdva7ZRW/9vG2vNvz92dK7fmF1DLZOH9bOK7nhq6aKTYhwM
qHBODKwOjyCSG2fzOACnsI2rFaKeh9BjvkV1U7HhL5eTK81HbYZrqUZ7sFfyHcccPzw8p0SdhtIU
6X/mok5b2yxduugcawF+Wa2GTdzNJJeyP724NARjOwdCGLXXGvXtuTT9UeNXGKUBAyLOJOI2SSDX
+B2QRIzuQc3+G27F8MsLTiU7dky9vyGFGanyRO27N1Lt+gnqQyspu7skhE6lmtCEJ58Ar9AWpbWa
GJfoNEDZE7+wNbYXKDEsJhd3CiJn/SkhgUMe+OKu3WUerDl6d5WePOUKHyXacjNmQu9X36qfCI30
vU9DnjFWQy2pc1hQ4iauw0qtZS62dn4ZEVHBqqenP+lmqk+MIukIsQibCsIkPD8CI/J0kb+nycW9
sgmTwnuIKRrHkFJPyVqdYPm9KDpfgnk3UHxU/6eLNGfkfYcAfUWxT6nZIJ3gCjB5oQtlyd0yA6OA
sVygVcQU2zGVtZvlvxJdo6Tr13dj8/u/JfZrMtVpBD9PYYaVq39Z71cC1gJWhZP8wUdUCmzlfWyE
qTkNTo6gcwSDcpvje+cBr+PEj84X5kyybFr442wOF7A5jokwmGiBxdwNHzhlxvBiFk/o9gizg9nw
cWtr6CI8rJ1MrFmoZlolQobbGUy5492L7k2JKKLkIwh/DNjva9OQ5EqVi/CYQN9CtgRmObKrlW42
LchzwU8uFvEBGTfLy8Z9C8cc+GHO5IbxwNFrOxvoXzZxcY29x695/BOLalklaUpE2PN4OaTuD8XI
ZqmzbHrD1TFSgw2G2qVBVIIkinVBe3oiY7aIZo4HO5ZDNYRx7bDLy8u4PycI4YvYNO8yAcxAqBTp
Y5OBnWVe69Gd76uwuhbkXHFSZE/N0QFz4orQ1/eL6pyNYiTkhdQcQN/apR2yVo8jW7p26FXbn2RC
/Rr6/rrhLiC3aOLQfjbaRWN9b+SJb1ZnJhzOY0sLmmyqcjT2iAC9uZgrzwCnahNu34n5BXUd5nRe
s8VjwoAe561bNMBCAN7L6kjSBjBf7ialt/1JRifOItWc6umEQmzpeh1Bx8D+89H9sMfytRnQr/5B
2rx3nfHD3jcl+8oVC9Voi4MG6sFg6XT/sl+TedX/UFu/Vh4eWlwjjpPAwhDxRMnGlZhEt/UvosJU
01WHMW/b5W7+QpA+emMF3azj7j3vcQH5cpn7SgPTchBwGvwIa9mAh2IpmC4OLIGM6OpgTCgLYclA
/WBBrMPCpxYuqVTgBxjL4JGhwhj3fYYs6U88EKJCtwAo9nCQJHq6jH6ubsFh1D3xAfyLO0FYfWYQ
K2SG+wK7gfgqqU/VoLfnKa+BaEL5vSO3eeY3XfTkIuwu/dl9Bo3sAxLn+sL/T+pP1x3b/r4YNJh2
uMh60+O+RdAJpq5W7lavWIYl5Y43tbh7n1TWJn48UXhV/yysdYB7tw/zRR5Gytrx4z5vhnI/Twns
z7shsHD++F6I2AJvP00c+/mTr9rDrGRQCifRpXMbtprjoBbljDfkvsIXf2cxak8Ci/SAaGcu9Uon
Y8w++BdKosebJtmI8EjrAk/CMOJxLhkZ34nIp1b+QpjItZyRg16l51p9+iSRrH5ThYP4NDV42oL5
tusaJOOW6lSbSWF3rvP5GoASN1kPpEEV1HVvubHXy551/m8UHGjxEQgekyjiLZtWSk3zVHIwyLUw
h5CCoHkWqJRYDwjzvdONiFA1XP+kkc/wIjBG3No1ls9pjMphAsEUGnJXWT8P4veK2FRNwGAiLuxl
IniaS9Z8jNEZaEZm+Rxll1hcwSVFXvaQgk0oQxoK/uwezWvO0B8Sjcz+joaV1TV/vRlaEVvD0CHu
Up9tDDe/WfRh4s2+OOf9z1RLTa2P2H6UOzaeDY1ck61ueoBZehIAXwhe1PzHGB0m5pZ8dPoMmOg9
HfelpgrL+lF7WOG/LwWrCcAAN7BGsGTNMGTmRZxe7GR32sCDemK1FsDJlPoSc+3t5C2fj3f/qacp
qD9H8TZ6hJ8cLOiXWcQ4MRjFWVBdtR+Z4eVt7VNT6lqcrW/mg9tGWAC+bz6tcDXJMENBGHBWy/cA
jRT0XZR7Z04yCXrJlVdOmiNQTruL3K1MYftAuOGRVfVin0zXR6fvlEnMkE+yjXSaFmUI6VPFeHBK
qU6EKEPfvM1BjLmydM33AqTBDCKR6fvEXGhU640TeX4dQkXnucoVfrESKXkAQTGgABaOpnfWomDg
TcUBkA6McZrkCKdjUzpKAcszC5ZbQJIjE9Y/2EczFHGnAoNP/viTheftmrdk4bUoqH2jUgujacEi
lcmdEWz+GXH9IjRX2HgOMqnQrM35uoGYFNwqAz2dhEQlvgLQq6CSFLxSZHWXUsc3sUmmw8hUkwBX
scDYBM7eF4NPpKly+LeGD8tIbicDbWEW+/Xx/mkmhVDWvVYBoEpBwkrqWZSHM7iP8DSvtJXHNlg1
/+KMatN1Vgv02JVRDLxxNHwUPJymuos6gCN2v7M6bOOKGE+l440NRt01C+rtFG5rmGLUtZ0JKaEm
VRPzr9XhCmQMutPJQQ6Gy4gP8KojZIsjntiuDNjcZe1rfI2NBP/QW8GQcSrwEWTZb8ENN11MBDtQ
8A4DndthxrYCPlRZhCfrtnGnU5VqPqnEnaFjvmKnT1yFSyQESsxFkSBp56YGnjbxZZoamIJEsSoC
/cVOeRpHMy5JKwlUCQ1ApdxpYxJMWJgxHlvGMnKr2AYJm7fNOk30NZ1SaLHXc85CZQ+kjfuo3clr
WrGjD/6FzcMmL0f7pKYBQDjfrTYhu4DWjGFwe17LubiG2gbPfcAA9xAORUpQ4vBhxf7GoH8Lcl2u
O3MtFHuBceW+p2EMUgyv+wS2h9WvUH9XZSHdU3JFXb1B79wKQ18bgtR+QcwpI/837QCxORw3TY9Q
a99xcAi6PL8pK30zq/RlfhlpD0uiMbUO4vt847fmSHlyxlhZNgOUD/QzxRXVFVoX1Ww+hotOyDIL
iEW2Px4LW2Z3tGQSdI8Hqepe8sO8qrHFv2z27tfe8N925K/2hFZgvNkBSOxS0DzIUFsvc5Dbsf9e
86Fz0kUiTVJ/pLNDxKY/1DTKl7VWUNirkW0ryPSYww3hf+qbGnyl7G8tqII6Grmz+mlGTAybq7zI
4YO4Ca7u19FfmuzKsG6AnFn57M5kKZ7wHcDJxE3MTLYkBqHaeTdkicdEoSNu47njKhKtQn+aEd7Z
UevUSdy/2USUtBnfQLOQfGZKqR3zIFXc/1iNDMqB6woCoUieYSiesD2US3w9C96OzLsfyAYQvpi6
5gPzBDRi8ZFYZ+bOQieuh8PIba0k1qfAUi3PqnpOmXcTeMpR1F+gCQW+c13zqDOlXsq6yHa72J2l
FSCmZuakXbHncKWG7WHjG8iawDuEuRZjteaD3mgX01mlOe7GDJ06+JltZUW0+fCLn1yugb4TJmz5
98IDHB4wbDPB/xiGQvfGNdRMSCHdvP4BUOsCDgMk0JFT39UBIKwfzdEc4qSfAqwsDat1cD+yPV+D
ElQkitrLiOORRr3sPmlkHM4oxCE/lVdNKun/X91KWedbCZx2f6zMxliNC/xuSevetBf98Zg/QDOl
6EGER/xvJsAkDlMEiXFo2qbZxwlGSt0vaw5lUUSXrw31aNmLhf/Yg2Vv5spKue2vBZlGTR97jlFc
gIYFwWhV3GAxOvi2A4x0RVRaytDPaOKc1Nh7GpzeMMHAhS8Hael6vkNHP4hNQvmjQ19kgdktwiya
zWtIeijslfZHdx5UZIgUqPo+rOZYiT1AsV67e8QKV/PKH3n7HuI12wPbNOtEV3I0IgsALA2EDnKD
4dt+loPq/UovIkEZt/QJTzOVTkqT87BP2MiVqHfRlNHYu/oFpEe63eVo34NCDMSK8m6zn3DzgQFn
cMajDw43hNE8fWq73FYRaI3v5lgYgr7Rz4SojuUkRTFkfpcXAwG9weDpL+XL1Pu6o7h1tqABArlk
HewyhE5FoBs1feI8ZwC3Q/H5OnM7MpPIi3t6g0DYHDi/BFEPZPSf+Vc9U/vN7ppPvv/4+jXiQez6
lTbgsxoS5mW/GQ9sA/ZvPLsCcTNyBIAMD9JdXLzcz0WiTqvO5dqxsVTndPhXgdoxTPqMRSJakLiq
qn2PSMw0BuCRG3b8D/OB81S8iwRCWabbU+zT/lr+mEej1WukKd9J39QDfO4achXilPerg19ylMOb
qoApwBLDLYNyEZxFS9d9ebxGEA8aEisJkvi8seuMpcqTPQljsuDYhujCh/AwWBC4i3i/MgBn8V87
KYpawdHiQh5k3L//FR0jZcUvIOKu94ZwViAGLsjtZSfM4DuWgatJENPv/FPoZ9BGRrEz3IpA11Uq
JyTO7T6rFJ8OenNOdfMWMYrM0MGNF0bBLTVnfeiwRw7dVUd2GuJqQtdoNnzwWuarH89Akym2q8M0
XS91ak97DQv3kfRM35f/pyKly/DyqfHZV9VkMo9ypdwhbgTQ5GQYJBI3uXCwxh0jKR5SN6y3/Uvf
WRwn3gCgrPTVmxipjOUPM6flkChGGgOSNQXpbJrxpfEMtOqGbTaN76+mQZZP8bvPrRqBK4lcP83J
ULIiBkIVrLVzVHlaD30wTg6zTb0ZyCURXibTHCi+nqaT5N4LlDBfPIiXTyKmiubk1vXCg9fozWNw
wg5u9lF4/8SDMFhKP8HSDt8YDCf1Op+sjaGD3EuhhcxkKPC4IY1fFWMgU22aa0dFO+KuZJxirB5m
nPHz+WRzATDluxThMZp5NI3a3rAIgp8rIJ8yo300GsmmYTzoDk/8ytHkkUo6Wh6Qkopgvord2547
lll3iRRIvEcBpryzuIsHOiZoHi/Mcc6VovAlPytYLnlowPrHPfGORZLxqkUke6pBn/aVKj+/VdAB
AjQAcNlgZlmHZpRlsaBSlOZ4YsMeilCjAXSPlvJFzqMSVPsixsKVoHr/ElOVSqvnie1mIksiFktP
hVWSPmrhrAt3VYUqJxKLC0NnUgL8Ap5y8KhfIjjNkakB0JUsWEraY8dU8lVRubhgghyI4KAGJpS4
KaD1HL+mIQSZH/+lsR5Gztzr0UasX+T9572hNvfI8aBsbyYukWqqwjvJ3uhqyLoQcR5VD68bgdPk
1VgR16w46dMw52EqTHLbsn0mmLcZLzUaaHnQrz2gmSSVLEkvuQrTJpVetuAoB9M5SLza97cMWyT8
8P/webNEH01cChuaB3IBdEVBKMn2FZJhNb6bl2w7hclpHHGF/yZYUCqCgbzgCs6qnKSgKcK+jk/x
pQSnPy7J2w2D7tykA7Fv96LVOh7wTiom3sJHCdnVH519XWf3KoYhlUKKSGoEVgLoie40I2nFMRD8
LqCcryqzpO1rM+j7EBC8/e5HSDNJl+qW/99949iCSATS97sDIglFHvyQPdD1Q7eT/SP/T9mLvqR6
GE8ZIkHzru/ZgvY0r9P76v8TZw+/eZBV0cCtf7u2diBoB6sXGST8ZXDN8WNT+euOPadHUrgm59Z+
d98v9NqqOu+pj7XvEy9epj0/zuTmIvdIN+2BkXABm4JiSdKdM5MWyictrIlAe81Gy1rPSqo6ELR5
pevf1S8q5SulG2+EmrXp5d9LSJmZYuCI2LN0vl61v1ADBSW07yUoid9j1f4aKdC6s6FnLKlppayA
7NqMt8pB04w76smALX8ICu6JF3cR5ZAj3k9dBgSNLqqFM+Eb2xJX1msnJeli32JtlbHq9hr5opmw
efLrtpqqtPlQmpcxB5DXYuwGFDUI5YjcblASp849/3o333MTUm453xWwvjCOvANTQZtqBKu6wumn
Gqah3XR3gOZhlfNPIijL2Xba4bTH2/sQ3dX/ocffFyAU7AZlvFro37j6wepRIJFDcEoXozLYCo4u
N6+N4w7ZExYVG2xQPbSxOJn1lfqzu1dJII8nScg8SX4UEeFXTvzVZ8s8g76/OV3J1YpwoPsH89nh
e2hQC7RhOkUI80jDqAhF8uIB8PezLg0X6YZUCUQitJO8H/HpAEvSWNwwrli0EaoIWnMj61k+Xwpu
KrmpyNc+8dW6JNvFfDGBJxMTPtoRKrCgm3QC2WcNJUsbMhlTLB0keMl7QQqtbEQyk5BztUhTkOf8
TGYXu+42/OLQmhLcWai+fWl/PVjPGiYzY3ByDbCxlL06JmWkcpZctzdYhJ271jnbzu0aUe4NtxIH
PQY02uy1HWCuscyze69T47vz4f86YnLragsJI+aDHk3HQU3MdyJ1sJFWkCPbjgk29itUdAL1AGff
A3VYvR+UmuWbSZxjZP1YT+5bFSG5V7LHMAp8yPrdPchQ4IJlmkyhf5VjJ7CudoAZLeIy6KwX1MPI
hD7VCykrAEf372+Xf6p8/hnMbwQQbEBNHlE2Nc2ZZIFIoPyP42lDVoSMtkliXnXf8R4fP/jSwvAx
eJvPQBz9ryU8DZZPUmVlG4BnGcYM1ZFTPTVpWP59ittsCMJHI4ypkCVK8Kckn5RH29G+hRo7zWdb
kns514DbZFhOtPXBFWIhQ1iAxNpqVlFdu5RTopCSjlGA7IEBzxmYxDIJOKCV3c39ZrkHD0zFlIpJ
ByhxZ0j8TMiBD4fKjpQmuTWvzARwE3MnwDCvA9WjDhh+oAcwtABqpmDu/sNHAgtEEbXWmA5jn3QI
2jGzYQsQdTzai8AyuQAMpSfMe9X+FHoJBBjDNmuTiZMi7gE2eu5dxx9TfdKYkrpylRukLLnpKSfE
1abjfKgYyZkXxIrisx71f/O+NLQm3CAkZQOqJ3WgJ3/qND+du0Y08XWzxZOVE4qw6n9c1Ipxxf/P
cw+nMf4H/isE6w06hhzlqdccd0KogUo7DBVNbqwAIQeAAsKhpa1OWd80qF9Kb6/VduNgcdI8Aol1
F1Vlaoj+9aiYEffZZODIdiV25x+PEaHI0ImG8OE5zAQnJ2LdSsI34j9Uk652ksXybTjpPRRRfMMo
BqDnAJo4nho9Mp/V30f+nmPUUqFqyS5nBSASreaMrvJmQVBXDsAe/FkjQ7O1mZgAfBK6+4rgQZAF
YCUSNJO3WX+5YSwuFSiGXZtHdkxLX/IGGy0LjAIwmncqRyNvPxwO5nMRaPl4IVdKgMYA81N6Bako
tGvlPVG5lKq7gknN4jZhyxsOtxHXeN2gZ4H8gHNtuRftlJeu6cW2uE24jEsQ5nv26oK1miyjMAW1
oDTcZq8sDgvRijCLzlFJW9uroxlL1wHx6ofJAvipGyElTblzYjP1miqh5lirRMKvhEMQWApKAF88
z9KwFwMOpEv6ujbYnFnuZnDScdbywMizXO8bSVrSOompAhlcRQyptE5GONycPqwq09Ke1B4PNJn8
nEWPpWs4IFNVnMIBv0oXzDKHXIK/WBJane91m3oiZhAPx5JqOHYLNz7nX1RUGMYDQbNaduuYIuis
3TsMBNvMZL9voZKliwsh28jvmwrKNPpwJ0LGgLAu19ZF7v79ZE1PtlKbEU9Ihr1zxZMMDly6q+kJ
xCRJb0vXYTN+VhQDViGotr2yQNgGKrh91bOLij1Y3dvT/AdPECr2KAF/+AAZbJP8Kmfak2uE5BdX
J2L3FfhK7mdxXEd2BOpvIr3YcyovqkhTVSBne7wpPNSsdTqOQINiT38/nFx2GGYeWw+K4NHahMc8
N3VNQwJPIeX9Rbc5xEOemKbl7VpYlwrUvkN08azhIyRk7Eet8vaorJr0q8SAW57EfynNwkLtBKNY
i+W4TDlAI4aypeQGLmaPhsAmpFheY78NExd4TIcEqgoHo5pnKVZw06ygsWJ9y7UAEi3kj/Hx1z+g
C4rj6lByQe98WpbguSNH/uSbg2aKvJOzk4TLaZIEsRr++ldlS7mUpEDSveqR6WLChOzXDhuAEhuN
hHly26Lzn+LsO38nppoaxx41+86pNf8muHjWr378aM2Lw97QMZbNfKV9wuRgngowXVh57V7KAqmy
fM27KiF38mPZ7X24olwxKq+ScQ3S11SX46Ccccl19u3olNIUzPK2E+/k4LSoz74dLde8Mj9k3dqx
VUuaVu9VzZkwsJNJe0puN6FKjR5uVTcuAWYEwE/3AYp0aoUGLl1Q6HnynTg0c3yx6MvsfsP1iITt
3T4joWMtq9I94BFTCRteuOfcD82r2QaZ5ufMl0pkjmVf1Y469RBded0hjifflSQmplAdD27pdLkN
Ej3rK9oK/GyC41vTKvZGq3maE46SF1ujzwSppDp7AMqkSYeBrK6O3ksY5eZtemhwSXoSOYTxos8q
SMN6O1D64wjbY0dY98hC0k9SYBUyHsezLTkdsxd/k+yfb18qTJBGD2eOgYYDgA0oZBZCEsJ+dhEM
PEc4GWxQ5t+da3TqF84zq3Wy+1xn3vMDmwvmyAVpD4mEEjXda/B+IM6KNevSW3YdF57VBHyG7+7J
iTLnTnt58iTK26XJu5sSEcEwSHr3BL6563s5sdQf02Iv20UUUNyvytYazcKv6M5QDm15yRyzx7Vd
3/U3YUZY/+UzRJaAYQzCP9Yw8b8BSjVedRtGmCc8n9xEGLwFe2hjaseb23DvYiN8OtM17zayH87y
udXwjxhF9CNmyVpZyTpASylMa302YQ7V5209Zl75UvBDgXjxPr04I9yCQUNnwYqKM27rNFEWzW5T
NQRBuguvImX/1THVCbnMiEuFiGYZh0+2JAWK/MblqOiaAUNOzLpSJYrwtSXHX38h6gSN8mwF23kg
933ULHy4355CcO8Cu6aVBzTIqn+w/fSbF7s8x0MkZjYkbTSyofrsdu3uTMYqUi6kWfgB2cEFiSCT
4kcQffnP1iE1WQbGySWTmlOLdEnMizfvokdWncdb3RbX00TdEE99R8/6aDmba+RScPqlVGIvarnG
mVEKhLo2b3cN16roupblgugnHU4xh8UxUXCUsBR34VlE4UPkirswb90cMjCU4xa/j1l9RTEGW54F
JOlWiquhbhPkTP5r+8U2vy3E5P/gJi3Ru1VNnrZzFK/8reh05XLU9aDqbeiVM6lEOsQglQt1qTE3
3WaltznkaxlVcVKs8/gwnj9fYMlfeQ0ocbZGVu9wHi0r62NNlSt6tOJqoVG4dTD9nZOsr2+tZks4
vPezRttohI+IEdvTrEHAfvT3T+jIxj03ExP/5F8DVFvzQM1+c1C3GQG4h9cs2V3qEAJZ0gAWYdsN
rvKBOs1oSU4gMXVEEl+nlxoH8/dCuVmOXSs/8HoIPvKes9aYDmAQNmsPUYq5puJh/GhDWq1+cq0k
4lPKy5RvdHheL//LzQfjJs80u7JDiu2xA8DXXDs1uLH2vJPt3HEWNmRLF8g2YrYq/ysltcmyeNL0
NiFP2X9AGJqE7nAxpMP39vXw3Ml/JW4WnBPk6p6FmMAUvNxSSlbXVOm3q0QQA0+pHb/BSTrycnyc
rk2wUeAxl6njTG0Ky46mYjulmO6mx79DiUssOyF7ZCSHqptB6afHyqFRwc0FY5Uxo6DTSM7Bfenl
q1HXMLCDGG0ruZHya7FV4Y6UcHZZaHZC/Sa5TjGjTjnCTA+VcjjP6EuOh1XfDDiCsJeHoQ/8i/G7
sfg3q4SxRXmJ7tSfsRNXFEMYSRKacsUehGDGy2apiNUJCs6uxVraybUjBcQkqn56An4TP72/y865
tg/Ii4jkDJlRHq9OB3QzIfwnOA/JfbKRmbuQDaFeLo44ev+YP1DrFhCLBUvFBZfYcXZXOkoKOQbU
9wLWAKh3hzQ+eiVccEOld1VEfGfsM6n6vQVbiKSKHJZz3k3ZDBK6sYt+JKeQgBQYWqObR9Ug2NsQ
jyt1vAmIjgimuAcXTW6pjrhW1QwQDCYwWQBVjP4V2aHVmYNijVRiTFjB2uS4aigICZ018/Kya2A3
2YrvjWiSXyD0eIyL6J7aYv5HVadwGaJwjK8iadrJcGzKFDsRTTgKsPFEhKh9SKp1VfEwAT/NCcsa
KrBznyrXDYLDn6yUYxASvwBAKI0spkSXT39IkuP7Ia6sRBTmD90zzo24ju0UznkIwEHO+h0aJS41
e0XTj34TJjBwHxnONXe8QQsXgNWviAsUzbrab/GqpJiXqWLhQ8gPoi5Y/qhXi0YmUgbhXst35tB1
GLiLRZYa8dwS56fzZe2PP2blYC/L7ZSTBidKZDOhI7VfJLBJYPhRMcfULM1E0sK0Yhuqg5ljmRIm
se1foMxWAFJVgunLvRDUjoHZQ0LD9vng4x3lpsPFP912maUBd6juYiRMUWUZ3bvyQMWwwu2nhpI5
uD0bWpYFozYiQRB4o1daanR49nwb5OH+RQQSmX/IKFVa239oQGfh1r5fwrsDV63If0g3roTztJ/h
Wmy7iL9Ksw+qsYcPlv6utGsUVrxkE/xorNq2C0/xBX+qIz8ahxReqfGJuZyIEaARRvCGGEJu/TDO
9Y4X57C3toa+lHO2UW+QA+ZVOPMwuNj/rcsBcH4ktOKxrCZHGWeK/nNAe0vUWEMujQzvY6a2HnFp
8cdGcdVQmYqJNsHUEugxbDr32kQRFhfLvUStOLn6GnfyXq/fCsmC6+yU39zD+BXbD3Kzi7TpwUe6
9HtnCFdAIZtO3+Uvj6Ep2+/ZoH8/pR1pyRPvWfVAstQeC1FJQNdRS64a+PwZ+d4DLeOokWgzbtzY
hP4N432lM0y+jZvAuZYpnvBH+R4YaSX8BQGACqdI9dQO6VsoOoHqpNwpqom0F4QLDmbkdNXZe1Cs
B9YoCnvioopFybj3nQ4gtc9k73kn8o3KTdWiCqK2QgyNXA11HUgiYZdMeTg2K5EHEd9eRV7s/aU4
SnoNMEY35MLDLJKEBqa5BCUr9zRA+KSXcD93pDE7me7yUn9kQPnWCizxWo62y/LCSzdeiblczeyf
Q6ulyKjLOZF3ypnasqj8UkqTOsWh5GFL01xIR1kJ3VT51YQstv83UMEkVlJ0kXgw/7gTzPLzySHN
VBdbj/HIu8jFN9yKnXwcC6951brRAJ3bt6UZE7Gqsa45GiAQGO5HbHHMxC6bgQs+Ge5WveH691jr
evkJBsxsM19yJZNvecPQJFFL4OVevg95Mu0Goa0e21PslFqsGazihOMJOSLLU3hIlZ+W3t+9sQyG
ED46ddaqG0GTC82tFTMphz8kdCMWFeAHx7MC9X0FmWx2UsNoUly+nE41gSi72KpJTteGQZjtnwau
ayVENz6XIb6sDSk+DGIxJbWmKCnK4WOsb38YYuMi79UBMQwoyv/UtHOMZDz+qkMWKtrf2ACDH7yS
bEZRWBXjl0ACQlXGy1gqKBA6z3zjlNVvUZHlLH0FOeWnm95U43pmnwh3ZGsyWFyrROF6f2ZALa2/
0Tipvi6v9FrtpoCQp8QrxycuW8sAQPtslfGCYLR8wwiCDyzlmu3UwJQJ2jIdMXnR1UVU7J/bvFfo
2DF4Gb4401IuI8TF4mlACD0G7ndp8Sza/kaNyYhi66hrc6jRKC7GVPUho4kddDRz20GD9km1KpKS
gdfakbzxJmLbFPZwCwxt36LLMz+hMaBZXdPysNpCmxfhiBhIRVL8ePr+zC3lUJ3wTXqUu34eCQXT
DINOjNKybj5oQ2UE+l5g++BbuZqaVO73Pe7E3y2fjmCVP3lOJ6YiGNPxAIKdFuqEDspiA5XA1K2O
JcqCyGbEIZ/gKynJCBvlZiC0ZJXOeXTl7IIXFP9WLT0YcyQoWt+Qtqpw+XUb9zLyEohANtcfM67F
HgeoeUxcr33wpnvVCAV88E1MzlQ/gqAdnQWOcwafqKJiIICYDYKoAItxcfowNQSG/X10eVQe3Ph8
SGCPD6gBfPxpWB7HcBIN/yrIZuF2qw89SrTPJQdM0FbfkPdt2q8UrEFDhtWd++LtsQQZy/YVrNvH
ZelFAXIwG6SK8ZThIkiXsaRsTUhehkr+59ZpzKzT52rEU/qzDC5ItzuiH2Gylx2eXUZyKf8mKpkM
GcZ/Mv6IsTQVCWLxqhHtdmmQ7zHsRUmoFmGakSzdlIOQgPlFCYTmVcJrNQsQys+U0/d8O5R+2Ky4
C0WTIzFxZZIq2TvcVJB2UGCo+J87p659aYvCGmm7QEVClxdAIuEL+eG1UEJC07YKBEAYeoV0hRpV
T4iHTIxP6kV/JDIMROLeLCQpwi8TaiTdrjxyRHP9xMzyERkPTO7WMF0xpzl1AL9e2msSHkiaaeU4
KD/iaoXuWEtFeb1LbWNqvv0kQTPlBCUWm38I9aJMRN9bei6WQaHPitpwFw5tdMEGdu+Rw46gBCe+
C+wN8oxgaleULHfhHmqQol2wElTjrevsTBF2pm8C8GgJ7rgDWC6BkKQhxLXBym5MYW5CTctacYDa
q1G6FmfpWawG6QFQNoBqBH8YsD5UhwxS2AkRZXY/pmG5fcBiuP/Y4RVcqfJBDZQBBvURkZCmFbEZ
4HEu1AHkpTcortCXOLmIUoVoEw8jGJ4BUen9HH3PoZLQqKp4D6oOaqhf62OJEJ19CIYZ2yXb51ST
d50ytLq5XV6piBmOIuvaOKAtjU0xYNOwMQM5et5a2tuSA+h89kgMDep7u2CtiYiSOHD4F7PvZ+87
IQkKy/0KW0sZ2LQu/6juYR0MupyFOJD+HJVtnAf9rmI/4jP9QpSu7UhzhOsccvD5FeSOCVERtxcX
fpfpZdWHfojcZ1B013iYQE7FHp1h/BMZIVqs+8RIKJJMlQU67LcQCeQhbZ18M4jB46/Tkcoob1bD
hLe+wXqTs/4DeZq3QlbEtpSdc/Wh1w+g6/GTKSIYB3RENetH0lDrbLa0w9sd9EY8XvIFWcJEsFi8
wrWlFz5EB0jFJ4W5D0ByplIX8YgNtBUZ4qVDq4kV9Vz3eDOgdKB7JXpAB6EMUS3dkgPe8DdhDuLm
oYJrqLCkf0jd6SVPAIBevBiRkOwpgh93uWEVddi5X8HCADvJ6SGJfRE0qrWI08uHU/J3J/W5Ceyv
dsA2iXe9SOx46zNrJAfTZgDgE0JLJ4D0qhSh7Yv2cV65/KaC4F+UntQkRfW5Tj7C3Bb9/YX/CWOP
DgV1EIx/8GrlUvtXcPT8r4GGlQJ0HCSVYSkC7AlX9ES0kSVlZovBnh7IUutbSK8Lx5TfhTwXvgaB
zYuZYWyq1r1Z84xUm+WxZK8mN7BSdH7mIaZiBpOnqKUABrEJqC/iieuR46C4SIBR8d+V4k/c3kPq
WuVZUcj2oT5RxT0yJJtrcC2LTesfWp6wHoZOIWfBjlKjw9/pYmMbbk0mDeKYBr1bhhHveWMhDHyo
5rZYvu6R31hpFy+ujsvpFnvWC8duwKeWFzaNR6E0qhbfOxBw5gyyZWxBWHIRZvIabHtIC+iEw471
vWwgKCv/jBwc6GgFzOilTO7y2ognzHImzLHRi18MgI5aW2DMNUphfSTvoZ0ISnwxD/ivmXYuknfJ
LrijPYYnAavCNL7mr2+oe51zrem259llIXCTz1UhNLcqbGSGnNErs5GC34rG/Hsr7RhN432dgRgH
JPpd1/O1Ke8GLwoM6y5TVS9tR1BLZnRsTTcREMtKx/MiQJw6LnorNTXkxYV0rCXDpdo0gyH9X9g3
a8Ocx+fZ3NWUv6vRbu2cpyV2ioXxYk7yI+sXjoZSmyS+Rczsqz9mTyyFLHDRk2HqkdfyoFUeD8IV
imv/GMjRChqzj73bCyx6L1zqTdkrSOhsBPw0NCfI6sNtFx0CFlpj0dvClXhz+i/KY7nUI7PZ4Sq/
pDOTbOKsj/Bp2uZWw3tp3HmgcIctLBaZsEycjShD5goB2wtDs6U4HLA+hRtQnjLxrD4Fkd9KXxMb
33Za3T6rbIUGa1P6j0VQdEEHbeaGW6lCC/Yqv0VF1RQF2buf2M83X0yjjKttLgQ1a9EfjuLzKMnj
ORRyu1lqB7aAhttSMDDG5QttFX9NWhF4mHhzxRZUEXtWyzMsa/v36KTcYA40yc8uMzhJOAJ/I4sB
2tRXSWAwe4Xs1gfvCddoXEv+Nb/zCCr3M3RMgoz1qLESBTjC0mYpoPLHBb2LlRkg0oj9f/xdrZCU
QcTCa9XPzXNzq3FoHcZiaCm9w8CfzB3swqF9VTERIEod9ff7OSu1LlqSiLV/7CBa/X75oVSXi2l/
+mruEUYkS6rvhEbsw9dWS5F83cA+pbglI+EPF+xv4ooHlKNSjrQaClqUse+eIPIao4vzW4PYL3lO
vI2eNkYpUMHTO8hFv0uRv7pgNbolf9nhjiggzKLviHFloiImkPLavHwCHDH47Krra91JzJYkcaSd
1Bzd47ItNe2ahyEcCSHr79meEnxdJaqbj9E6M6DaVUGmU25/DDIbEbTNeSJ6t+UwoDorpze53BAI
yrEDLJ9THPEaUquTJHmpZtD05JyOnoVgXNJgTRRVxo1Q+/5ijwhAsESgXBlw2hkzzdqUIf0LLLDp
MMd0LYHhY4lwjTUzAKTtUEOb0oKXwwtlp+Rk/63QIWbHo6+yg9x3Bs5ii2a6JGe2HwVMLHUFly5/
B3RgLLpFMrtHA6lBZggpP8jIqx4jOrTbV9TSWEwz42O0oGEA4zo+XdqhWm5QDDXdPsSm6ZZujSYA
zqGDiC73DTDQpTi59OJmGeE7jCLzgWftEMmWNIqJi8AeVeIsjHZ8yKrq43KJl3hY6M/ybS9k8j2h
TE60BxSxx7W/fqdTdLJF5DktvC6AZMK0aKAoiRI4H70D1JB4UYGoss3gXY+gMyPzSHCAJQL2qO3o
cvWhwWSuRK5mb9Zl1+TIKTm1BMmNRi7xPxm96mpkLxoEpm56/1N0AC2swyQZNvphHuNkp9JKTrIM
EwJqRmJIEogV09ZfLmPjn6Zx4ALbvKt3HPcoTozlhX+Yv3LVIMdSD1BRaHwfSK/GfJpxRNSmuDjY
OKdSmVVfvEq/Qf2h6iLWU0DHFEG89KI8AAI7dJlQ/B3f7Q/7G/Ier9/UMaWyKTFFzFl5hbTBxNXQ
Xq6iNY28hjZ/UoY9bCPb29MoctLhGrLnCBaBWN/SwlTS7AoQmOBq3pmc5zHDtmaM5wa/3w3Q0Dt2
ptSTHtJQ9K7SU8Sm3/jLXs9DoiIAyYiyp0YSpSKwCEVCFvINyvGLAmJAfSfBtvsiYDk=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity fpMult is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  data_a :  in std_logic_vector(31 downto 0);
  data_b :  in std_logic_vector(31 downto 0);
  result :  out std_logic_vector(31 downto 0));
end fpMult;
architecture beh of fpMult is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \(FP_Mult)/(fpMult)\
port(
  clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  rstn: in std_logic;
  data_a : in std_logic_vector(31 downto 0);
  data_b : in std_logic_vector(31 downto 0);
  result : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
FP_Mult_inst: \(FP_Mult)/(fpMult)\
port map(
  clk => clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  rstn => rstn,
  data_a(31 downto 0) => data_a(31 downto 0),
  data_b(31 downto 0) => data_b(31 downto 0),
  result(31 downto 0) => result(31 downto 0));
end beh;

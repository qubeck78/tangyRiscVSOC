--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Sun Feb 18 13:15:53 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_HS/data/fifo_hs.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_HS/data/fifo_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
cwjH8KICVYPfzkercoEQG+p4zkmHD+O7VWGKhKmt82XL5ID13lvVTkiTPzk+lrQiGUGt54aY7QSN
tiWlQgp4A44xG5uwj+UoIGfPE+5i/spp4aECPb8BatHXeWCTqjcSJHK1sDi4+X2tl7GSJxEC/n7u
mUBISeed0em12vmTOqk/J2EKNIkR+UCtxas9utRWRkjVA8Im4/ZODa2qHSEJxR/EnVDzS30MPaum
uLGKiEIHRT6ZGc3unscodVG/JxLxYL3YimX+WozIvYu7mSaFKWbyk5lu8Ssz4rjXOKWm02KRzex5
2drPwIGHH00B3AwR/umzNXRxCSiIz7mUaGW3lg==

`protect encoding=(enctype="base64", line_length=76, bytes=34816)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
qTKesSHGKICwapGL/m/zU6ApHLEjSf0nWd+8v3Q9pk+WVUHNOvOsx7cIEP9L0Cb8A9I9Y4OMkZlA
cMOyUxMJJntXCC9K2UuhcIoc0rzJv1wpmHYgz9+xszS7c/+xjC3vJEa3Qdxgcj7JH3lLJfLyBUS+
xQqdZ/qucaeTBQaisq9NQnPuJW8UuNyDnKolwUQPYegWiL6DPwmK41oZy+UTw0GDN8RdSYj//QFP
d0UEDBSmGYFm+GWtmkfxjSZwPVqs1ABo5XPQczVfcp64iKf0IVqQ8NjmgRl6H8Xf/fXaQ2jSXpwe
O7ZAxeuA+q0WMPsBF/s4deiTcIjsQFt/Z9btRoYPQj+ikozmiAKkqmN4pRMNKohRrFpNqhzirF5R
rFx/yKtnHM/egNrr0lNZvJIAEUutY1+VhKfeEH5JWdw/rtRUUOL8I5nzyG88wv1Z89QFkIacXLKz
jCOSk8OldwkI1zcP/dspgNxYo9Uhmy5r+Xo3P/RoNLtPdNSSDvu+ixRDR4/Xu6T0Ac3mfaYih/SS
9I08yXJFYwSJ7FG7wnH44caANKxWK9Vj9hyv5x9YslPNG2Tp0OFF+5l0m8wLLA4f+E2VDobSZpPs
mTxf8b1lCZAdnvlpPaSQn7l2hQVwIdqOL/kNeD1YXUNWtQfIsipk34ugy3wnNMQ0twTxbcXsFI4m
7LeHy8yYzKttWbmF4YjCDcuo4HjDbWNJA5jJnTWur0XSU4QSA3D7fjFsypQPl1ysm2YKd+sCmNxr
mF0AgI4phfMC3Lzxo8u5Hbx+Xrx2x9LbP9cuqJgmIMsokrRaWzVtHLw9yb7u+egcwYf5l6ichktr
FaQIit91s9iy4B+6tC0DaND23XARiXjB4STSRfzhZPmo72w8EoXVIQw/xndinvNmQRmi/1gy/6MO
ZG8C1tyjqIpTQcd+oVKxXdMfilT9lkbiaXABGft7MIyZSsvgyufajGE2EKATK4wdfXBBpF36fca7
UhVVR+D+JPbZr2okYckM5fC9o3TkKXlOv8l8nIGni0fooWhwBbRBVMUWIVOxwtEoXo7bIF4aYMtV
wUCR2KQyeiWrxC0vLlzsAMxJBac2BP81gTz6C3dYeo7lmV4FHShcMyp6DkPUEFTcxqSRQKJF/9Ku
tYDfiroEiXRffu1xCrBTtbA82F19fE1CTkHlXFcKLXCoJYC5+3bzttXdrl+IiO9yvz2mXpYQcto4
N/EjPvn4K7niWeW+OpTuFF3TAs9lgdoLMiDXc+yxwAB9b0pT10nqfZOeEoNFSRgzuPuiMTX0yIZW
5fXwWD31ou8M0luwpdwHTWYht9NPx9c1gE3eiH/Z54MY4YdS0gfDOvr+Y70Y8ziuViMrlFSZKCkw
MTiynzjOlgWTyTPSIn5muVT2uOuTZEk82TVekyeLyJ7CzYt8INt4NS7N65oFgVatbIeONhKC95lN
PBuIsg2JIbZ1tPVuoyKkIg00Rb44qgwakXDfPu4o1XjDaFb4tSRkOq03I9KMtq7R0fX/VZYatY3f
Bd+/9WfEQ/htd/dEHlAh08TYV1OZXxOCYqHFVsReS1FX2amnI1ECr5jLPA68fMSNYY9R1nqAJUEz
/NCirnhqTAAgLVsSOahSB46TYMHWHl270HF5oZPM7vAZv8ksAJ9rWTFAqHMootm4OkR65NjQKzKW
ZAibjhdSGTCW1VJoF34OfaWJ+4n0p9a9qPymgvQHOiUlD776hbF8UqnKscwXKdZVuEw+AYBcV+Hf
StSTcicyGvJPj+pWp72JQZVHxvC6yVClxaOixdTM/x/Vdi6zSdPlI8u4gft4yZkHkq315w88u9Tj
gZRgDdhDViL4rdUaIsf6H64sMvlHugxUQ9NA532Ljbek64e5mUTtFghwHZus2csomAsUI0IGj46C
UzwbSDun4DghtvKMjtKwYrQWFViQBsoq6P7w2USx6zv4gkNqtPX+icHxRQOGuqQ0BD6qKhE78wkW
PC8XfbIEvp/S4uy/va1tD/O8VgfgqmZEQJIw9rl3brB3R5ZhwsVGUImCrGGlRawhIniUdEb2kn08
+S50Zm+z+fYzfjWoLHlnW+wU1PxVvIooCdmvs199iEk93UnaqnSuJ4n8SbMA/buT9WDg6mzU3iAQ
pbzJPSLv0K2dkDoLEtodLE7v+BptWxHpAbNRTthK7C1UdN3yp0Cktp7mMG/OEGaKarBih87Q37in
V98gG0hlywpZ7tArRCTkOE+xT9+dKA08XUQ7HjgE8RfVki3OSN9c8Cz+/iAdnp7ArY5//aN5C6vp
Ha0DadYXYn7460pVEkwUL3EU4IuldczWEJsFQXdgIoMZGEnOvYNddTYr6LxDBMXc+EN738T22wUs
Q+vsPJ/pJH7yA3vS4GT0cvK4fKLuh8Kn2w8cQHSE9Z3Om+1s/mvy001DJUHI5qaZHWvpme3Dr4i7
+4q1Ap7myF+Rue6Xe7QawAsp94KZBre2I/1N8WUHRZaPR+d4dH86oVwMu8D1YChM9NVE/vAxoaeY
g7V8brOREaBo4i01vRgwV9i6nk2sO9Likrr+tKIg+eAbnLVGqnP9BeauSmgmXTmkDuE1rWtuA98p
XV4bzJ3UgiIMNaJtlAa21kZN4Qukh9HqFLwYNlQHMX+DZaRwIkaPCme6+xpqs85WT6hU3Ex3cilx
CVZxsXOGkkF8CYixUeuFkIOPEfY0FuR8dBSyPeDAYOQQJf/42yE9/JT1jLVyY3AKwu8RypZfxj7m
WhyUjpj0PQf6jcMyS9nyhakXJcPhvw9w8y9FctX+GJtDqaRB25fEBNarYbOSLLAtyG24jvANt9Dv
BuR2k5BEHZYD3mAOVWk9gbtKahIy9c+vz1UsP2kHYiqzt0rhyFD+j6hcZ6MURsneuOY+xfFa0q9J
E3Z6u9N8AG5OnksmXJX413CYfRzcRw/Yw4IxN0evLLXlyoaplGFkU1GJZGffJqlnvjFSyuw5j0GM
KfP5Os2OdzZec333e63Y/nUM61NkKDUSL+NYcqkORGU0u7iAkLUHSn5g0JLdNFeWMbnM3FFSWTOM
cz9a5MdwU4F8Zain3XJFba5olEkWGaSpgA4wBXV92sMLMg1La4Dcls5NgMwnASr0q6uqJABn0Z+6
drCtB9Fw1cOzcA5167k2BrEvhSyYZ3T5F8TT2Dv5InfLrjw3vzGVt3eofByiR8/mzuptW2NTtrSn
/nxOTLclA4FXcXizTn8csoFfYNtdZFLGi7MU8BTeNLqdNdkX00BwZPtTsW6l7YHR2UJiCbVI9HQ/
ZhnEdazQRiCU/BkHjyHnfAe7McsuWUiAgRThpx8PRI4udK/bJxocjfVR/HEVlQi9mXHV+fGTOd7O
cgfYxYtJRsOJMBb5h/vO068ihqLvVu04e/wVeFmWQmQAKLmr2R8PZ8ByaDVn12QK+IS61G7SNI2n
FR1o1czUCXrZWezuDQ0L8HnTFfvgefp6L6NSB+y5nomqJKlmpvQ7zTGHTBjegA61HKH8Rv2JnpUg
cNax08XTA6nAhm/pSSyXMp/B8+thw3L3+JUjcHVu0zXjKZERDNwB/Ham5JzshQO+r4xqHzkf73AB
uF6Vk2OIXfYkqVLuzXhgyW0nyLuoanbgUYlMoWlXb77qaOd+mc7zSyBvoKfFfSjn4dPHpReSOXIv
xxIu0L3JEoyuePD/GcFi5CLUKe5ehbYyEg99J1LZE5SYuq6ErHBLyuJ11BCKo3pnsMTb86scr3UG
Czy41ahJfX2UYB1yexg3aIBzF9s6nEiUTloXFLbNHP+sKdUaJvxJowILpDiWIxhtUG4pFTga5PO9
r1Qr4CoEMiMkP+5wgT1eWYn/CxczqA5ntf7LrId0DqkH679XjV1Lq/XuxznNxsSf2a2ot0PnSHgz
mqe/91NCGgB9nYj7tAxDRdZ/Lcao7thMN5kZcb/rlZqdb8/DdIIhCJ+/oB4vE6FmFg321Bwz6ePm
9nWUbVRQIgfNTHV0XOXUNZpLkUyor1piil40zs8i95tvmamSyfszNUlFB3OLxKnxAjIDvxTCnWva
Bq7irN/qwkQ5Jnfv+CMU7Ndz4oc+gJmQ36T57g6RzwMPHQqUgsP+JQDA+aCwkg0jGhYFLtoZOzNO
COq1xuhdvX4UpPDdk36nBXcmXhkoHkj8Wq4VZUD/s1MMI6t3Sfq7BjyMi3A2unFz+J0L44ZCpDQe
V7uuREJ4bZ6SS0ueFU1Alfg9RHU/Kpk1ecSJKCA0ac+eeIffWFlLOAqw9j3A1hsDLSMpvk/M9ttw
xv24FfE/aNgsCSNFq7uA7iNvfCkjtjpdbUZaUo9IGlndjBPeJyx26476v8lYqoJXbfQPHRdZ13mP
7fO0GXciim9HA8JnkC91N/R2d/rbiRXYu5lUu8QVgVi6VWLQVS7c2EiEkFclPiHmol7RrWRcr7sv
UQr6KHlbl8JG0ANDIA/moiiOJUiYRtNmfEU0h1I4XeyWCXXovecgFuwAGUXVHvNDvaGfWojjjt74
Y5fn+gE41YY4OHd9sZMVEtYP+H7Jc1HH8kVH5HnBe1wbHYbzoDoR/DCV6nXztdgO28mjoWkgupaZ
8PiSG1qoifKrGpmbZh0O1jP/X4MSLIohk9mY9Q/ubMmhmthHQjseXpmfZbplVkLYLxs2uCvN44cW
Tlix5wdPuVV97cuMKsLfyFn5L2kDcjYDLbGZU0EKqu1EfDfGfkrAZR9/FNO3NcBI5HidqqD46Ap6
IOWGu7A5P8QRUGLQhbnM+9GxooohOjwWY99Skf86jinzdeMAzpU1Iw4zML67731efm/g3HUwnEKF
EIjBCzGCTX2UDlzUjmbmKWv1GcZVlsGsiJ7bQQTg8LvVMFVvKE2G78UawW7jCkL0Srrcyx0E70zh
yZ19wa8EzQoa7fgm0j9+LwRK4D69cvHJGfrgsFJUbKD6pCqyDvNuL7WJksysze3/nUxteAUCs5x6
kIkODUNl7KfYl9Mh6jTctYyN0PlYBfrKD8JrCM+k5z6++xPndbPLndhud2fQuvKh52Svm2VQmVN1
txsvGoJhycErls65EybD4egvBCSmQDfWbrYVV7Ud2Rvanyid+G+7C3ua5+yp4ZGp70sT/7pxh62i
JOqJH0oJv+J+gCmpx28llSIE8k1RttzcWGdcVFQL2je3d54V3CGgRh0DfgfztBMueL6DguFPCb/A
7s65hKXHku+71+joIki2UGiwp8TEEec4+NFmAoUe3GX+BDwevSHydpBb9TwUaXyTilGEyvdGUzzQ
kfejliDHAFM02noi0+J2U34eJmktMuSjHbZ8SaYq55dFex2n3k/PNlUBmV9MTYv3TZLmuOsjGXWB
2QRBuuJL2sW6+PTYbiPtB3LzvbFPX8mo/pqYNQDe2vh/9n04GGJm36QobkbftNSe5BPxM0bh+u4J
lQs3lK2hndu92S1mGlzTNtHNwba+zplb6jmy6NStHh0s1ipQzcJXsO7a9lx0AEIVZEXBS0nZB/vS
9E+xcSt43x46I5b1y+0974SSesz3H3+KUY6WXJh4JNFKfOF4i5JsrWQf5EBzOLaJTAIw9f7gXXQE
C5U9gq6J7fsl/4n8GQ0vvV4cKDAznTzhglu35V9VdqBzQ6UrH/1STI2V2CQYKNeECmfN3Ydjouot
J3BK74IzUjQsqXujXbv2CB43/IbEBBz5GQtl/mCYgTawxNsvDDnipmyQ+FBtT/KC3oNzOz56zYeD
9P2YKKl1jhSCv2pJPY39sx9cNyHosj4DnR4cAdjBVjsJA8ZOPh9o+3AVXbHcKoJ2i76f/Y05ZAXb
4hv/wv7+ERc2qRHrzC9RlbLV2z0AD4BvTIt4WQeKhMA0nrBzQwYKnH+3h6oSxicpMcLHpmMRKY2u
NHhOdtyuKeyzvc8JEjyXpBTHPzMLPQ/GoODBS2uq5hsn/YTKJuGSTVE0YLEb3PEDeGQK+XX/o6tS
Ab3YSuI+mu7dvRHn8Fx9OhQsUaeCWLhSDHc6XinSmOer2xy4b1yUQOfyEqsrqn2hdVlSQ8xbQVCa
YiGmd9as4PPuvCaaIx599d7HPRlMM9QKAFHAw2UXI+thKDM8CFBF7TPD4v8srMZcPBk6cUsCSaC4
jx8qVNWRDIWLb/NLHJAsw/WPwns+cAksWuEsT/BtW5IW2FLjJwYKlZgVPe5Ow46YbdiQC+bIOMO8
EjSfs4nmfuBwWFbfS0tZP4IzYikL3xeByax1xY/Gw30ete9EeObL60x/6V/OtwZMcKnTuDsPGd8x
JvkKJzaB90kN5tnkIZrq5TKCypl0zoF/dQEn6H+tTcAdLRrMXk2LZTTo4wV6tlyrxlfNZHSFEkIq
tGEtRHEK4+hgcgyhfyRUNzlxc6fO+FyhnaulcYTaDxysYLxUmbmKqktlpZJbbEzEWGiIciIsArmu
u56NNwxv33kZ+khL1a+/EbzgJPch+zCABZGJvka4kzUbZOnsPjrXBOG25M+3C3mfol883TVOpQuz
ygcb/dNxkhSvE+nt6Oi8y7bMDJuCso8WKQr+Mj/WiuEwtXs2gy0i8hPB37N3+aAaUoVnMTFHNBi0
ekN2t6c+JPNAdRVE84kUWeTrSEYk0Sl9WH8vCPQffzqoG7tJl2QS1ZeZpek3HFzUFDAXJcIWJLBS
1keGlxRTtIb6c9cJzMANwttp5n97XLBwqpDUcpcUkgk8fy0q5xdKKbvpeEzja31fXJWPRep04jJO
ixvDXf86hBv4o2rrYzFwS+VApfrciEWauaYKunD6I0KBDcePWdSPoT1BDB/6QlEv8wbPZp3MY/Mi
I+dt6iTSOQYr1O87KAqzYO5w3q8uY4fxoDDEFiG/e2gXSz29296nuxFf7Xse3KKrGrLG1Fcsc3Y1
AhecHcU8GiIxgW4auM3hHYB24MIIlskNPSWx/LIlNq19z/m86UR6wovPsOeeZUuYIUPHXAYCAIEI
NdnpoTWQEdDKJPfGBr629gZPnIXJIFI04Izf7/V6/pKQrCC/1bkn2DMqFBrJrB/UEP6u7VlVwpjJ
9c4o4Sa6sJ2d+QHK2cTEACZX5ezq00kSj3oSMIOOSl9M4lB6Ja4CUk8DiPM2jO1M+U7C/GfTy2cF
Usa5gcIi7WW9UPuElo1OJOUFw2zIvN1UHraXyT53MFmmxIm9gyol8CsfigIajNxyOj2SelXUkMFW
7iVgmUv7Cr+Vbwc0IDCdaHEq+BF+ExZxJQULMYcCwSjgnnLbzcn1NsfYrH/3voggL6J4kdKG/ne/
/6lmLhh192U+dLgQ50dmhZqxS/aPI8R66R/eaOLwNvIUJ+cQF6GYCw3bi/NmeRijHI1K9LNGzA5C
NLwlJQUYjzin6JKaws8pfcF8MiFuKE4EcmYlJBhTwclQBlGL2cfnrxnzyF54FfYnBgak7s3ENxfk
msd/IwnPwtniqzyojNJryJwW4Lt1WcUz59MvLlm32lD6Mt6zgJ2a+jBii7g97OS00QwK4SUly/EL
Ie0x7/tvkTCUCa/IfcLyYodMsfggu5V5qMSSlndglOTt4DFBQSDIN9hfd8jqPHilb58lJ3qd+kpw
SC71XDZ/v/VCUp3rnzEQBjAOvNbqPbOz97awJFo4cWl+MnxwAUxOkmgiVnrLQYCgNXiRcEq8OKu0
773YiHDH8XdIPrgce1vCq6CpijcpcN9Qv5RYKXnMhps+5reW3IG7TSmNXtI5hVfO/bjWMpzLKERp
Z0t4vsjQftfiUIgdpD17HSuEWQayzqjZO/hZn8Y4KqGHzBVbSsRtv1G9z2MbeyIedvUn3ZpJ8d5+
KdE726IIYjYnCVNU7/vwml2yhrwF4zoG+XygIeNOfG5V99N+bPF67bh8qZS+QeEFs0caqRfRJ5Go
/a4ZZlXXTcFYosL0aNlPpLXFmSmtDjagt7gvG1bKwN/t5ZOJlzNAKlzsyhLYHXWTU5Iq2J3Lwhcu
IoCu1Ezbhr85jw4PejBcnBfc3T5SLsjzZiDmfjKZ9zf/Cr9mF6jSg0rNLvFyDlbSO+crb++3pEVK
Ti562KVwmNtYHyHWWP5AF0t69njf+FAEYkS7G1XoZzCgrFpcGQju/ShNVuhxmFM2HF+Phfi/byVN
50MNYkFPhq+A6ROM1X/O3+jL+3Gd8Ukbj0iOS64eQG5lu/Yd4pPi5YfvZSLPYdBppieKqTwNES1T
zynDciQyUl9gEYvdP3RQLLpjDZrfdBb/idbw6ATCIYNRDaJxB1PmxI35nzNoptueznTR6VvOgKcw
uKii6VdxEMrKj9S5YyZTHZbH/+xv0vmNIk7HBc6w5DFwxAGDk0i9jxhqWDuBnZGVHRdUj4lfAFwk
6WrTu05mKpLejFkMnshHM0gEes4igOT07jBqkCeSdGVUGi+TpsbZ296jt2Q46IE7PRwzxNlB+ld+
Ur1vAp5BETLtjpCZq2znY/QOQIHjGo/IFZDQihZQHEm26YwdGl9w4lILACJA06znb4jt4iZghG/o
dQAYuOqRzoKuuvvHUK4pFi42/SCTwMe8/TMAOPeOzD16cWWIkB99eDyrtpBC3ZMeCxViBcoKuxj1
ePrdiNIUqJFXFXl7g5q433pIOGQThn3d8IQcTJdvngz+lQTprXmgysPm+HiaY7r5sodf0JwDAExA
RbdvEglQpcGzyGkE17rCrMcjLIzYkYu0nS7VDlQ00S1JEbcW/pIiTzJdzRdQAGj9n20v+RXXQ7Qo
L6LcWiEUVFAOv49dmz3abkSQSjQxwg+yRALox0fODlINvOLq+zlvXV6GOKgO6Sis99DMhBKTwnns
oeihOfF20vmneE5HGaDGNdEW8Ee4Z6eGhnA3g9EklrkV9Mg6TRZsr6mIsY3Ir35eztSWyRhmmCWd
gNQMa5TJVb1OyH2MNb2gkcmssJrPJ50sva5FvyMOXfwpZ1aNqHpkQWgOl4lQF2mHUPMXxxLSVn77
HCNktUHXA+ajAfwPodYXxrYXl2Fv39DMvI8V6lDvh5xy1HbjYMOxGwpPAVRlqROBi9vZTEFmtO9/
Bjxg5ghUe1sLdjEDZ6k0+KK2LoFnQTU7Zs5OTeXAmoyLa6R46q99DDoSZKkFbgbpN3xC4M+VUzrW
NDfM1uErJS96cN/jNa2CB4F5t8VDcMXt2KQgLec2pCG+uq7WS2Wmyx0tIbzSn/RPFew7n0s/Xeav
t1dJUNqFYFSLBVwmli6NI4BfQ33AG6/dNbfbw72Jb1yXu2tdE5+Bg8mXTbNWv/RfzW2/+kF5AcLY
yK3zTIBWjQuPwlt230eVxN1jANNdgZEn01vdlWyHj1wJ3TqKNARklb9gifultzbDd7nRYR7L3MzB
FXTqZ08Myi/xiXtkYlBcfutKRatlGgCnQskLKdecosPc5JNc6cKLi5INavdWqhWLnJjX3sAV8y+n
7QC552KlSC0+gcpR595uyDPxWOcxiJ/U9wqgR19suh9ZzfW0jEATOVzUnmlLkS//v/S7UxQ++bbI
uqLEoMa/EEFIQT7facTuFOb0ySP90oZaQ1+JPDYwQ+MP1S4M/EIis1KoENmDL7WHwXRCuYbgS3Y8
S0tHTp1/VIule/lzOll/93P5JeqtX+s0FPj1u66tb6Erk9/U1KA3pPLMsUkva2PD6delXGdQCAJO
x+ox1CIB2WaYsJgGYJ/m7FEwpuBVO9TfdXyAVMyrqYOwq02KIg/uQvxmOIJhgjRUgl67jaiI7dSJ
m+jtJ9QQVyVUaooRyb5UqnOJjahrQg/Pabvrb3XuRXHnT01rEnCAlzQJ0edxzUjBXPkeLYqHUbg5
ANTczXsZqcM4CIzQyeXPxSabHQSLrtqnO5QvuTolgZ/fvBlRK074JtqCzEgi+cCL1xnkxzFug1Sf
gbVDe7a5jDF4QvvT5ik4AC9PCBVfQbXhA8h8fDBVbIcQoKvzGRyTJwt7pzjg8nNpTQHWuP8suU8f
CpfxONcNCmjOkJsU0QneQY8Lbt2YZPhI7scagwE2aq3KBt1hQASoYhwZZapaDiEHPM++hTnrkZ0c
TkuR1/wLZyiEdQRekpqbs+5XFUoykrMPqUMLb3TGPYS+9Sf0rhn+zuStsw3jdFRq5AAJN9/zY1KC
6fkoxd5RaKnpLd45kCVlAATG1DPBxamJIAJYJJsilShsJU/EjrD/2KJkLgNHhCk8SSMubl89CxLJ
dr53+g0uQBApSJ/UshdfXx4S0FttIT8gC7gMA1sLjeegaPado8rdY8s5xtyJR7WAFG43lq6zYhpi
lqqr9ZWQ2TfFXjFAndy9etYJSe0+yMKFiR9DpWpLk0qcoyw5wqyD1PvoVgGMbO73N+uGN9sFfOxq
1C2VhhJWd7DyWIQj/NFavKS+ePlk9jZKrLvSficg0j4ilihN1YlEAWnIDQ5ZSfApYHLzU454hTtx
hT9wpggU6HN0Dn+T/ALY4dxsYvC5839/17WkF5FdzA+wHgFBfFn8pTAtptLmU0cegUWKBmUjuIEl
grfWMkZmUdAXxZWmjo5S8rfM9olBOaiUzfJvbTILuDQb0si55XheNmXbrsxMBVfZscBOSI3sgM/C
+bMGOWNPE8E/F1qT9c0JaS+5hBaKowbK912JfFP9HnwLik5Kj6CxuU5CBaLhNI1aAyowyHBArdKp
N31YWD3LsgheQj0qSL+u7q2TGGWQWqeRj/A2uvnmKg50Z48XUTsczVEgsW6jG8pzxcy/iDh/AVOw
61kSlKqyDoB2TKR1JjJLqY9XTmvrwmc5NztcUtwO/Lgu5my5yezST9EgUZUEUi1J/Xxr/fpLhutW
G6aMq8lXYi+VA5exuyIcD9FrDW2MXn4NpBXsl53DH/PDNYQjleAm3g59ETpW/cu286Q0M2AyYOwx
zuHSpAlZdBGlbJmvUVxw17Y8i/lSiDvEG2DXWibQkBaPDprCjOYQgNquXfdcRG/1REE2FUKXRoBW
Zfk3wVy1WPP2we+2AYTzgE87uZMTauOUv5Do3Pog0DYF46w2730XYdxw8OBrngDMgb6dGc5kNZrb
GVAOXYQCXTVy+hG7h/UdamHA5CEJVkP3Q4e9app+JCWkDDn8cAl+ELL6yTs8vd6kloV7lS7zuPw6
R95wRktVXrF+vLO2XQOjBNoJLJGwAqMiRaaNuO+27U53WiyyLu/l1J2B+CBi0TFIueUnnF+CaUfB
4wf9sYq6AXp2EfwKbbtQS5S2KOf2Zk2ukwCH9mrjlTw2y6to8+4Qwrz268x1AdDIcuIULPV9lzxk
1y+TqI4NT634HQhluBTad80f+KoH5OF3HyiK3yKyM73dWdD32ph5MngAsfi5inz1artGuGQss23P
L6u7gq4yn5QqgMjXbhYbv3uXbuIZUUBb15lIHUaDs0aqC18bgHVejR2cBVDemtBCxiSlrLKscNDs
sK41R9uEQxc3DW9Mj1mHECJPaH7dFw5Cce6MNfgLhTypVvAT0UG5DzIrKt59gQkJe7wrPEfbyWHa
wFzX2olTi8eAr/RJ6SBp7nXH87TPIE7U3MsdzvWd+wH4aUoy1a1dZeexhY736EgaKcgU6ouMJLF5
Da0JwP2znzuNAGNANsHqNgbCRazBiJQ+x3emPl432b9SeBtoOfPkCpb8jWDIKWzy2AF/E+JfEKBn
jyPRAfC4SJwsRsh6Tb2C8vu12LyK9omfZB4+C5Jo+5VyuJbj+/v141zazIhKTQ5ZphY0yqyux+r6
aq5DNnCA01KYEK5+8JNYjCkoB/8yp8w2/pTAZdH0URXCVrFq7BHHTP0vsFL36DfZupN6DHWq4qHZ
SyTmIBVTxEstDrNnNqBNKqWQcpYiwPijazqhcQcye71r1p7WX4JjWdh1R3UgrNYpMK5UaOT4mP6f
AmqmwjQol2Rdu7Uv+WdQpL2b7h4kun/ppPkl/lBBHJpKV8AwlWRRAnZjgUSwKwvZCwbUBW7Je9Ge
fFindQHt7Y/XnTV41dF3yPDX/7KmTWduho/OtZjNxRtX8a2GP7nISn+21qnI+gUxwU9kVLP5pYhy
bIwcs+i4hxWl/ujBaWA63MLhTFNuhfrLeKn+b60tJCa5lwuVCTVrp/uEopO8C8L3R+xDjYJ3aADN
tHm+aSb3BesYgIobR+h2+WHK1OwPb6uX1J3Gkz0yyNSEeSAEzwQJo8+jRVsdA0NzlL+SoaeJVUIJ
XLlcVyuwaWYy4hvAjp7gmpcKmljk+UbZ7/moJ4Bvbhpbhyh3sxZADseVxjPLmZ8A68IblOEbYdcu
hhzEPFel0yQSg59UVySLLK4zQWAdZntSX0Kx7vO27E6FGtrECVPcmhtDdiIbsemeQdiS6gQmvZNH
G8kvWlNG0NwMxmgEajF9SA+waKatbdmwuOPDjui/X3REptqy8Ym11fQpxFmkeU4FxLwQ6DHFZvNA
45JXCMaRkIx8XVx1eUiUD0I9PscOYY1at+qC7TMuZoKSltZRrYJ6AQ5sPrtA84TEPeHKlJZLb9BB
fz1JHYGt4m2Ob7KDvHHrGKo//4a7r9/f/kQ3kMJfzVZ1hTs4myRH/axRJTEP2eqYw0aYzOPNOl80
VgamW9VAQcLdM1duhsJ++ILKFbFse4cy8wEjkb+VmbIB3Ms/4xkN8YgzYc8sAgcv8uiBIBCQZNqj
nTV71MDJLyaST7g9NEk2c/cK2Xx6Ch2rtxAVEOe6M0KFPWqA5LQRtWgz6Pmnd6dF4TJl2/vxeTkS
3dcTx1KZSnakDpAOVgl2fhavbBMpJCRD6UuL72r/k0N24Xm5a6PuX3Gvjnb7f0/HXqIoX39ABACS
Xsak9qZjzADUZABksqjeGc8g+JZgFLyxWEbh6XqZX2WkUi5a6CRVLXVjhBM6/L53IIr5bpeP5JgI
GXCYlHTXM4Ad4aql2gFXP0gSBc1OdAiLzMPsRs+qCNZVsbJX3y0jDG+IfnjaWmDOKXJgton7jASN
iQjZeCroG1MEmukAynmZ6fnkMDfPUnXZ3cs5prg/IKjqPNw0OBfYwrP8+91CuXTNrZL3FjZ/7qvO
GnGBp/K17g9cxWbms7OaQjNq/oXCmXUcyRJfvKjCNAdF+tMmFRHCwzfDmLzKqz+Xufpd6aOaQ4lH
XkXi6W0O6zp3gts1pRunoi3QGr0AmccyxKQzgbrqnxVNctPAfOIL+3rpGQD2mrvDe3bao6LsDwoJ
THuCz39zC3rn72Git4hvKwGo+GHDU/2LLqyCX1/sGByZZw56UiZmQSExlhcwIYdJgkr05OVH2hvN
5js57OhE5GyJlM71HL6ZE2OvKkp4loFGNQLejnSLgOJHC09W0g+a460HllSzk3/YOX4P3b5qXeUv
SlFEpoJFOtwWVWqpiy2gA9DdxtTmMF3qj4DTz87IEVdVQ9vcKvLmyLFDOpL+ZAqUvECsX5pDQv2b
sff8zy8+3sJwtNiBYpWXN5Ex6zlhyBewBGyNI+jljwveidm0co+1fybps1593N5UDsjn/1i9+2Y+
1kShCsOkiezkjdxIBBk0742OabUzDLzzwdOexFtQ7zSd2Ro/Rz0tnfJtpgUNwJwnu+iFUUv17+kW
Bb1tgzO4oRZemAHk/jJ2Q9PuhKhue23z3wd+a5FlaNhFC04j0yz2XZPLO2C4TGoEBn/CfvrUJStI
06sibZPdkT23PCAbEmrvPJ9Fg3qS97cNnBFmZucrLUsLj6ityl2RoMyFs9IIwihVn5sl4pZYgnl+
cPk9IRAD3+oFeiwC/Mml8k/5/NOImSDR0ImPgB/vMSRjOi7vx64TIVDkSsZ2vkFqOxd13pv49OzX
LVcDiVy5bd6D5gH1EEPDvkHQE+MI/VfLw8mHsunA4FRllZURxfEkE4SAj0y5e4yYmwSxeuqA0xN+
1NupEmzEJ8PatDQutmmXijfXvnBpmZro6KCke4RBdZYRMfY8AqX4UvzVR2/GSK0Kat+GSgkqsVsd
33Tjb4dDGTsP7668eeeE0zkIg3DCZa6nOH3lhnjxt1HCDEMwJNjUSIoGaViUIVdGUVm879cLupEz
M6wMlXfHsjuWDpmWtsF1TNZekSXsKE72uRwZ8YiTwDWZ2dt6LWDtAT/oleY/GUI2P651/6bUGNMF
j0GUKGsp63cf/Q8w0OuY0P5mWq3RPF2bH/JoJ9qUJh3MFNv5imtwjzxqjUVLOO6NLOR3smpxBnr6
Bg5CSVdYs70dHLzPsnbCFcQqBFKGkCHNzDvAb1CNIdpRwTIaSKydbab+KftBoH663PaFQjzr0Tzs
jDyZe3RTi19DJnYcuJiwUsVu6D1yTqj96k0n6cK2bcsWoxyUXOY1Ed6hednLWo42ATEBwJM/vmln
8SLvlnfiM3fc7fzjR5YGylxy4nVmOh026s1iK02RUUGwO1N3msJlqUIUZruIKLAmzZCJwqXshZLj
MrOQKrr8VDoK4y4afvs77Cuf5CPdMFYr+nd/vg7sYzSkKTgZjE0Tl0+32jSmD25RlOEMCP0TOqHR
CX9NmKcxKcup+lXHFurqH5px6BlKKLg/T3KWVRhXHB88eX4c25pWr/c80RrqQfTh/uJxK6RCbFCb
fjPREKYfDvy/B2vjOwjX/PVHseVng55TG0pw3RE4SCcgY0ig8HMaYUdiyDsYHx/UhVePEPFgw0fs
Fd29yWFqy9Yj1jDQXv13VYQlUJsY52k7CpelUK0UcTKX0l7zl3AgosA/hHxbSj8hPnnpry1zadW8
6tHAcN459IoJnYzpVLT2wUEIUk0D8vwig4AHhno9tuSf7c9dzDQOJ4r4/efUG5mRTf+uqDn55gO+
apqN6EC8oPOyRKt/QqsbfIVyra5s3uu9mFs6/E6kSJEzfFMXs/EWXqQ6R/GSvkHta1GIcR0GkZTc
C/8poRDh4/bSaqJybhKCT+QmtZEepXdM/bhFVxlmKur3ablZWif23rx8QUWjLeD8OJ+XEmzJPgAC
LojJVBIhDxHgRslA/lMpAVmpNcKj/huLCILYbDwY7QAH80MRH2kZYF1CpGXgmW38hJX4rJ42p+FH
vEA0JJPL73u2w8YYF3GYNfcqKe9sp2Aq+81+C+ZvK2dq8auNmJVThMLb1EUDUoP7yzbUPJ5XEvft
Rg8/3Geq8cauvuFVdKjZjFVj/a151D3cexL8Pw6bJoR1A9mLGyZ3j90ULiAOZTDyS3M633AqLRUH
puTGLr8dv1EkwcTloNiOegO9aMxnS1KH7aUgrk2CUY4X/u7eGcTkFn10i3JdUUipV0bnnV09Ildc
P8h3qUQRciZnZgeb1HHkk5tpBjO0Bqf7/lpwMvUVTzqtnZUXMledG86rskJPD+a93oRpHEZ95eK7
h6grEv92gVqNftqQECnc1vlimFSHM/ZvoHyjRXTF1oouKThpJ/MmkDmQXiyri4E/j01twGp5Unf8
x7Z6nqz0CGMpgg8YmxVsDfmH0PhItweDkuy7g497jnfotqv2QbIOanvlR1xDNAquohL7NQhFSc3o
x27LWp74Uynsh+0ocC9/FFERZziqLSugOcyvCBGgOE1/SZwVSD8PVW/XaOB+TyKBFFhSOvPuezFM
6+sq+b7h7oIHm/ylmt4ui2UOL0dMGFd03lIET2Uz3CqeW8MV7bmtbsZ+C3t6GdSmSrLrS0wcy1GD
AGWQXKuFmJozWBmQm3GkDROcN0av5aVtTpHXUUSi2YOFQ/OnseDosiET9LJ+5PpFMgOH2tvLEJGs
4+rNoGwh7vRcJyjEjG05VjpFwjLeUhL4HC1orY30+dD5b3y1m1PbVrrd6xBrn8CkyviXorkvyFY3
14qsyBOr02KQiQ9I5MFcFqeedm2SE8gaqr4nr8l6eChcIJQeFVA/qvlEJQwggurOrx/KTiA2nkAg
+Us2NQCBZYBOHn+VRaEcTogIP0UiIMGMEEZdGBQz5BUvcCkZX2O3ypHEXLmTxg+JWfytkBNGCmHd
snVHufg9rS1GK0k6LicsqCT5b3Vd8WZcSqthS0yvlmpOF0dnwzDM2vM5L+sC+aVkRDodc4pqjhMh
Ux+0jXfqi9x0ngUeIx0RTK8JKpL57leIXqRflU2D8m/YouDFvQyNiho5c7BVBgzIuKHZ8M9PmZwR
W/bpMGM7XCIZ95AdU4wZz7AMLKVFkDzasgkH0FYNdfHDQfQHCw3Fa4RdxpHW6qyguWbvLDQDl7gq
w+IP6nKV8Fk5alVSVM7HUhmmmG7ycKqCxs35zgxFmGxJcZ5aZoK5y47MKb0FO2YREstFX0Uqu+a4
6TfCNrDjJBkeKWjEfn2L8mp/9gEYyyKdQthxg1UNW48TSpPN9I6dRw4Kl2yUI7NfRB8l5nNSIjMd
UCvX0gyWJ1kQMyG2Mqfxr1qBhK3JReRGf9FECqOahYrEtTiCTE56tWkx9wcUd8lSaV7l7BXrxFKA
WL9HPYTXpn0jS+s6PBpHMLMKMWNs1DYhovHFKzjAoaPEKFk562XPcUVJkljZz6UpWxOjjWMJc9zR
/tDuNk9wJmttsHhZ+fQQsr4isH+cn/+FVcQt2V2Q9XKuInUeXDBKe0QeHlf1EkT1X9zXKJusHZoK
TKN9N65Pe0QZOZzmVE0Yw/zRjMcOVunkfvvI7JyTuU4gyNCUys4peWs19VVZ+cFYiQAF+8JVyH6L
ihd3NFWQDFTdVrJCgzWCvn3kEwrUKqYjiEq8xau6/LefUEcwA5yYrJSBWivO2dpqdg2AR4+rG2zV
SOmBepjGeW6FiRpCO0EUL3PSHNNg4muzfEacqce8IjihJ01UhUJQm9C/NynBoqGAZ3UUNGeaFX/L
yu/BRorzCIaZ1uJahrRpMoysmTvzo68eKW3WJ197le+ZuE+S7uyMIqmNU2l4PWqmQrH8i7RvO9fr
V5C3XQ0YHme7wYa6++cAfoP1kJdaQ6pmUM6MjDyTjBDRD0P6l3U8UrmUZcCUXQ7O3MT6Rj5c2Viw
gXyd79atu4xxNwvsHNoQb6i9ow0E6XHAJFCRFr7Rr8mVFGYBexPkOQeghFcD66KabSZ44UdIMF5W
aGoRvIyfRd4hibtvh/n/V/a4DO/5Qe8/vHedsROjwWxtfHhP1E5w8ENqSJwQALElV+OmMKsNhYSb
SjvemiJMOpti3XhO2I3YfZZcxjepsjNiYtXuvwK+nGoXQJKlMZ+DWBV3lxZ5tjwo5+yD8Ce0nIy5
83vxIhqr78WugZ3WlRsc9iiMybqKj7EocKxXF6TJf43fpVsOydWX44oOI8fT68uV+rrqd7FFxs8+
l8OJESGYtVo6zHnuPTdv2HZ1g5ljg8vnTUyRL88co84u2KMgUpNK15bQWHnMV5qpw9kOt3MSdpkJ
NykE8ZaN0gypurFcPoWvrfhUZNYPAfQllKDRetRfrBazmQYZeMYLMrCqY33KKD+YwTZeVDUNFbm0
EnuKlo7QwjLo4LmOOPU7I9K4jO4QwZ7KJ/mlnBy4bSBBVIiMGORCsVQtiXlAecfQm5SvfXT+vJpr
rGoVb/CyfxL0ne4cWuBYzgiqhwDXXvyrsou1gZisW0kDIcVdt2pM0j3+uVc7b9hoNJqc0Pb5l8wl
5w6Jt2e0Ky6jwzBg70I9yI2LFN4XQ+8MrkVu2/2kUeWbZIXc61oaLnf+YNIzyOrYRqHX43rNVcLy
knSsppRYg8H2IA71HYdhbQMC/mBZP0FR7EKpRJPJORFvIPOzA1hAEMZMPbi8Hm6rtaLgCmMGh32k
LkN91xOV5qpYUrTEY4wWF7F6yPGOOS2ndRuPOk3WIUFcP8xMj6Kbxe0shuqpglbHfc6Ku/KMDe4m
CE9JBWoghkyjw5LLLbgGq2uRqB9zpcHTzZT13+cPft7mXqWBuwgpOG24VUTr/WHTrAL+6x3qp4cZ
3a8NrpDeaxgcJNp4SxbTFZQgatKwGfMteNN40AMTLGApEUZqXQlipoA9srNkX7AuElum9C4ym07h
vwRkYQFitpeoJV+y5E1pyXwyYfDE4DObaiWBRXPyxE5467Nc+v8H6cf6kEX0ONFz9z1W6q17t4zp
V4esCqvc3sOhBBakxvF2casAdPpdlz3Qud1HDi3QcUPJFREcwKbJnHqCYud7xlnzl7vxFbNaNyBr
24nLbNtc2B/FEcDU7v3+OuZyOZn4dQFbxJRlra4bsGFtLVTBHsm2df0lhM3cCsGYa/KuTmlECqQl
UqrN24hcGzWITD9zeE/HpWVe5qwXwSTQ0Pt5Ztx6tZ1e61Rb3nOX/KmE/cgWPFhDaMysB83+4GnN
NCness3dGRhDb0+G+Z0xDUeQAAdn8CktgRNAguSUFKaGjyxyRW10KfeGs44Pn/gnYwlMEhFibGzz
tE8rIjDjqgYccDj9llECxs+OBlfJXn4z5SWr+v+MxiXxTHumfZ4dJU+mNIcLVN2Bb99sFqFD8wAN
zgYtdTrK08hhooY81SK7TiZCdzX8iQz5Mcwq0kONip6s1lDgqDjPeGenPEdD8PLZiMVuNhCLP/7o
++lVPVmB9RG6R1Bgi0e8nN56/w0BenuTj999bcBTdgB4EQe8tI4cI2PN6pHkK0UpVFkWiKgVPkEz
jq/fgNh7P3ZFJaSO7lXUyJIGkeM9gAkuQDoCoHtAE5Yy+WUhzjvY+Mm0zPX3/0n9ZOx6qXnKU6X9
nLvWY4xnt6ti/iYC0WF24dqJFdoMDHkysq1ZpHYSpAFG2kD3TzPzeeyWClHPWtYWlZ5EFKzlXGSC
A1X2V86RPmSrS4eEOT/zVrfMjjVzCC/sp05zoziv61YoyHuj6dTxuOcmItm/05X9fcp7JJg+nhca
ZJuJm7pkTl+QeMHpCNuQW5ZdC/LIZCuT8e3QGyiwG75TyvoE++Uq1MHpoDPCrza+qWrD9aQhq1yh
aF8baw4jWI/sWzd8MMo6Hdiz+ZbeYs6doTtW8ybBRHN9HVwwnZS9LSZEiYB6EVesSozH0S4GinFj
MzowrnOV8h6c1p+0ayRoW77/F69CsT7AF8VRqaFUa38y0kU7l0kF0g0e1Sxri7oETiFX2KhUxNK4
joAeJIqJXLfC0AuTr8yfJq43cUl34Yk5+KFSrz/u++/4YRv+hNUzVAQxmm1tdI3FQ2twIVBN/eEQ
HRj4Rn33N/FI20IVy5QQRtB8PVxes5Qt1++px/stAviQWRrje7QpEB2YDkDfvmYQIuzn08I/21d1
Y4tAUjemJOoy22ueuOYmme/Pgjwqg6LVXckuelPdQz4sO/nDWKNTqkH1e0fQ+w68/St8y/bck+qm
H7dw/SFDtkLWd6jRqNrNg1W2SuylZhL/4LehUI4vBPtFTDktocSyZx7WPqurdAnp3W9IUbWJnsxG
gRcUXN5B/rfdiXqjB8ZZpIeLSGUgf3S8G5F+9P0m+Hz0fFmWBcdtXdW7YP+fEBJLcY5sfoKDAdk0
a9wQYZv4h8TC34B1t1WDvTVSKp2kWTM+V8EMxpYapEUEbMKw+fO11swT52iT4g279ebtsgjqFGzd
eQemxfutHVeJNPIfxIbz/BWcyi4S/9I6pLJocRP+02yPEYHE7QXdQ9dgJdKHXBQ9JRHeBtRhMZNs
F/o3cGX0/nk5l5e4q6sjYQ/uOAMW3uw5mkNPhJjSHJKteAdehXgjWUo3aAapByN/rEWMET16bWWC
vc694P61ezJ9SnrFp3//9kAuMI7DhXOAt3eZzrudAIyIZ2gRt7BCj74Wo+VKu566heIxdiN58ZKQ
YGhU3CdAvdDAYSz6pTX+pbbqKsYA0fARBNhPlXiLu5lfPvb5s5qjAeidkbYCYWFdpdvCR0qZ+jAG
pnem2669yXSX9ay6DNS32TDUVb1IfpTnYBZGXvGnhSQy6gllsZqccP2cRLt2ppi7FG1aHWoF4gd4
eyUzxEo9B4hX58RgvzCZYcV1naXhWeZ7qex7y2u/rffRducgB8W/O23O7LOcsfJXpZkMG4JA9PP7
kDeJa/EEcZh0WqXfVyyti9Ro2IKyGa0hFEaTQLB72207TVSr/hYbT6a0Q6lTvedyxo6xJ5Wmm5sL
hekOh16RVTqfx5Kpc8p0QgJzVoOqI65/Rj82yRCjp3r3RIUOkECNvyGt1alCEyLp+QhI60oVxQbH
NEuPIaLkTiodeWWL7DZCshTuLY4nhg6LnlURZRITNWX8Dab0+fc7pR22F7AX+U5ZrjPlFwo6cQ7U
bE++oBT4ijfhjU4Jw/2dcT8He1oZ3qDvO3l2GewgbWpwCxFE3chajnku+ZoA2+hm568Dif14uNaa
j1kQBdNlw4sYsBSQ219J5UYHinTZievj75jIVhPP7SDRPtDlXt6I+k3tO0+/9OvuEWpl8ey3Ni+5
IEEtAiR+8ZFnvt6JTuGn7lxPTYd0WoodDa5wV7if0BXBgNPLYRpU8cwuoiMkGt9P98iXKWyn1uaJ
S0tpo96mRSISmjo9joSYbK0xUs9iPD4fT+okQKRx7YtWp5rnEqwuDBu4fUedXCNZKT8/oXWpy+l0
+f79fKAq8N4EF8UoNJrJBGtxIY4x9VGvliNbcjMGx6Wfc1VZDEfhEQ5axPi96Njk4SOtnFlTDELU
oi2Cy+dSm0qg65+uEXXVU6WLZoTfa3WGbMykUXhRidQYThZlUJiJX7WsJTKricM3grKwIBVdC7uP
QKr3Qv6nxfRBGOOt4LjK7r1zoy81zmeEbrdCtFWAJeRw3ncDJbsIR6Ba7lUJO05/BSNZngFeUwZN
c8IUY+JwOHB0wMhCJpJbOlqkgwI9YWlwDCZ0ZiNaQ544t5OVSDK16+7aK970jxy8V5WayRPEkRVD
xuCn4UXvsJpJhqAYBPcbwBJWYtxGLfmjT81KfS1OcqRMFgE82g2OHV5Ro7PU3y2NYddHwptjVwJd
EMWiawmylzghqwCHktVkL34K89BBJx5CkUiYi+eULzw8p6gawuGFvFpfyzRVDPv+nE9nttubK0bk
OS9h3Od0O8RPPnrzUNlrC0fd9jIKzTDwVz/poKR990oilrN8hjqDoSfpRDgiBLJY1Art/o/5AY+f
w10Yni8lxFBaLemIAMsA4J6lCUn8hq1IIkTLRsulGE87bMUoUP4pq/k1K9hRdtnT+J4LeSdDTfGc
AS1EZ+XSu67D5Ox5hoziVbE0zi+G6lp3BlztTtNTC0t5pZKPv8eAwNeWvh5TiBsVmZ/bl38u5JNS
ppcrWCcrEyyofj44/KfDNPzq7ha9nnQ7VQqSllmFLO+l8OgdDFqKHjfKKylfaMIxShf2q7ZGFz3+
UwTKUSyXUxD8Sjig0u02Ctxnzaat8Z14Q1g7XPsLuZriu7KjaZOE26OeVOirz3k3XjGo0ny5gIVG
jib2FG4mjng6ZMn0ZTnwUdEXo5AlTHHdN9PW772EWd/4KNFxYvgxMGq00JowlgZuBD5ytOP4ZBh/
1+oKl/6FZMEFh2m9k+9ywl0X2Uk4BdhFnHpzFmjr4OutXrowGlA5YKu6Jj4DIzNnCfbT5OG0r/Os
usWSskB2SgLafR93vADg9MClg4qs/jTojq/g6o2Cy1dRjVjB3kmcvbTka5O36DoNJ/b1WSwbEMbf
FodpuG/U1lnlSYgI33yOSJYzIfGEoLknofRPHf/evvLpIMypITyoUcck1d4cKQ+4RSFp70JJe+Ij
3oRqtbvzGikCQZgjfFwPXqJ2026wS9qychlhJ6em2jPhhUUvq4He2NPMr6bChKulSUujuN5YtuWW
wFIe8gDubsGZPqatkzv3slRChWoy3UChLuMMpoijxbcNH1A1+T1hyywfRDEGHAgS9M4R3nVmr0vq
aa5MpZFzuVfnDX1FkLBeRzRwi5c6wuTCGP51yIvXr7hUczxTiaiBESLXZv78DZ/r0bdKDzE60pTJ
kfJsGho4j04GtJvzInB4nJyC11a4k26ThxaCATT3G7LU3QoXEYoKuGfGpXdopIjlL9mhGao7BnYY
0r9ty+fROim5zwPxNm+C7ZXAOU4DZvQBngrmPCpg4rHfxlG378mfn3S0CbaWNEa35Cx6px3CkXFl
rXQV7NaoQ2zQNTSDV/lRk7T8IuTTgpIMXHDt0HODBbkJ/z93KRJAPwb8Df03RARsaRh3IZrh1XmK
fjWfr3Q3GtYbqN2m5/8cNpyACgo3rg5Y2d9P6Iez4LY3O8cikaptuoOMjuVeo8/bXijayIpmPt6W
QABsy8IlSoGoQZ4IW+AU4SaEav5XEU9KzPqBSjdhDODTj3mSBMsIGPs9KlxNVSr/HQUp4+7sKCVD
60q3IWnV8Ukx/Mm90Rr8cIEr41Rsh7AqvowPA6QyQGM2nPlKRNlQPnvHJlNcN+QFxTAoD1RwIEHD
wlY6DSHCZEfnRkcVGkQmz8DmRE/iIuXYjFyty8BK+i/4bfD8DlxBO9lT4LAMWwSboGJb/T3RUmw2
ncl+xPf9tkkLgHlzST3TcrwurOxB/9DNMQ5HF3DgWNT8oSnQM0DiwwDp+8b1YNbpiteydh/RH0IO
ygxItqcjFI91rb1f9ZS5b3QwuOKdprE5lk+3Af5TZigZf37DxGABwKMyWVOPW46ZP1F6K4Cx0r1l
oxekhDSes9j1M2PiV7uHJzSHbkvUzzT98qqaXeiibVi/GgPxMqViDjthGikVCFV3pgyHYFaMaH80
91SHC3H7V6NbZd0hSD/1FJXU0lb6E76+eQNc11tPQLzCEig8cC1i65uJDDPvZjXi/hTy3HtW7CRo
L/uZF9kd9vZ6agx4Cjc3iiVo93QBL65JJsrlw1RKTH0JVoTF++qtEfPpoTU7u4/GR6q+Xmr1sNfb
LKS62KA4SCkB5L/qs2vNodP5BvbP62c868HHhHlrkTrE44epyM3DrJfSxJJm/dVUvUt4HhziN+Fg
19el7aAH2PA+/4P3jLfmgt3TOD49wxp0RBhteRGe9fDl5+RZpm8JyPXOWyqN5hLoC+c3b/zjW8Sp
RTVAdMQrrzvM6HSGDVrjg/m3T2kfp6OFND3ZuCv8sNq30o1dQjIxU8Z0/cQlxD5paS7rLqHqxA8j
JrXt3Q4GvST5+ucwGgMT1qltpvvJ2andLV5sjD1CBP1ek7B7qi5QO2CNWxCCsf/lbQhEfpSqKrv4
6jXgkI9eDH6/DKL1mpFQf+JEPDz5DnRUBbYxhSpRlNZrgw8bHhGX5kP5Td8v1aXhfW2SZ2aQfSFS
Z78RwngGlCYhyAvGALIpxNl7OXZc/AssAuYboNio2g6EghmgUCFP6Q9HgRZv/leXZvf9yt/5KqXu
eQgV85LDDprLuxiFYHF+7TmGnH03mxVEDhx4gGoFDjwMrYXdpjyJNaHNYsVrEFZfXUCyUu2BNV8G
gRCKmZPH0ICzgPwc1me6owejnnzxIa4pZ59b58+UqE7vp0aICUlbXXU/iu6D3GUfWfzpkTI/MX3V
f45TlnEY7CakfypZm36BoN765UVJNP8YKC838AfODMZLm2C+gP2Q2bN9RW7CK0QGrXVq7INOYYSK
BM8moITrJqqA5+jWVn+1wJjRRxOOx+YHomUsYstjw8GYu867Ozkqaa/jZJM0E+HhaWWRmygn6Cl8
bCmgrRhc/uwn8ziI/ui05zWFaBCfTiri+cfU2n7y461NXIddtGugYe7TvjERBMQEomQMCN7XHbAX
rNcBUGmXrxmoMhR8PX/Q77yxKCD79GSdYMIYVC6qhm3n7WTyeDtZIwJGN0TDKDH3EQXbp4MMW8SL
hlkUcRzImXMwe7YQGtxBWQ/pNRFwZXxhmASRuXnzLxF0Q9cNroYxCMh0a2QhRy8zRBQDjk6+Hs2r
5VNH5hIUERzPmusmZaDjIOxTStfHIQVZxiwbDPXgqPaJQZidApN7JtpS3yZKHgzxKZyZgfSsxi/O
P9xzIzJa3kVn+Aimae+2yOzA5LeIhuLkweKlFVaTe1egUN6INCVGJ4NIQoYPjxFwzMVC7QANbSxR
gkdpzjVQzaFOZ6zZsGIXAA3jBzRLQmbvWfFcSuOYbFqqVawpuK6lsVm8IGLpqncXkf4wyu/LgxNP
TgPoHBg4HG3gQkmSNQZGbXMjQftjM65S+qYukA0SDMrbSG3D5/57744JOeYaYxUCnTjefRVE+Uk2
7aLdkMaLxa9oXtjpklQHXTp8F7FhvgPW11AA/L5pfVD0BPmA83wCy5N7tJmtJMvNiN7BcVS94xkE
sjZaidav6iSd1b7xA3OsaQSYd4CgeXBDrTwAvRb0GmJSjyO3i9lTw/G7PgTPY8id87W5JeFqESDX
zgkwT9KzuPkAUKEkeutkTTVpT2kr89xdxZOntEwBofbAWNsy+kV+aK3vz1LXhPRKpkJKda8/SZHL
BtSEJZ4jjT0eOn08otxViEbAkjXkk3NiD8azLcanGKXe0FTibut7IJKdyhPTb/4VPDIiL9vdzEwy
2y6N49Cl2MnpA2XqTw5JPXXIZaOT+PLxtiHBzI6fVxxMU5msJI/H1symjpU3vb6ssTNVEqxYQn6M
HpCg3XC0VmvUXBB7FFSJCSI9o20kP45kFJSRr237t6SxuE1RxJtTB1ZpJdte2YLphfEAC5HPulQR
kzmFyvOZkCOsjpN6S+UwEWhwOH7pLZ9e0dHGXIwjxgW4EAuObBm9PdlKGUGUg5Mc1Fh8rUyZU8C8
lOaZuklHOFUbYnJwnCMXVTFS6tMOiS1/PayN5ggy/G3hLuWYkToE7nor6cVaGs1fuXNbG40owY9P
6vsioH/G/lhia8xNifU0st7MHnkZZZKrFHnQyFvbTtaBbnWBDdsWAs8BLHKHBkmMadxSyz7QKX7d
s8B+odZL0PEViz1ceLoISBXQHeQ9f8Pr32v0mU7lKnIn29vZ5YlXpFJWi4AehH5qr54CX6mO5MJN
VuiqIqnLR+uZknY7wgxfMtHpOZ/ofqiq1n/rlIUTzmKvw+LKsHmNgpp/Lp9Y1w+4BcmvjrkcpmjB
SjxPBe9hrNmQ1tn4yTq9VwgJQm/sfSeQ+tOv+VIkmNN5IIQlbGWMfculrB8JXefAwLdHoJ87evh4
xWkDOzpoFxZUyBm7ApTgciGQn8s8aygD7OTT+TRkmOQN/D5s7j9wJfWrvanVwlKyxg79BnyAaxgI
L5hVoAbIjiaPzpOYQ30QhExmgqM6Wsbv9lDABx0QcigL3VkXb/YpZNm9NVFKSjPhjl8KgIj/duib
BAq13ADQq+bR8tkUxnZHF3Za+Dq0ZHDyTffipOfOffRUzK2OaE38zPuyEPMkEVhuPa8NsWLW2W1g
xRG3VbGaVN2vIGppb6K6k/xQlq03k1OIkgXLbHpX2hCcpL0AjXUEf5vs+wVS97OTONSaGwb9aOsS
rKQzU2FPjpd+JWFQKhhUwsGAbzgJ86UvZzoji5ZjEAybrWo3Wr3uSt5MZ9GgKK/CW7sjJYVZIk0S
PXgVAya5WEYyDaf3uK9McXNZQNj91vfJdooGQZdBJLXSAUNuu+WS7JMPQ2iY0IQDTWL+fDbaTeLh
kZqFhTGc4zN0wSU7B17iMlHrE9iGB9R+sbBa56OUiqe28saF/sql26fSCNohNAfEbwg7kBlKEfyQ
fl6Lnw9blWOVdmUI0oX8PEJTRyxtJgVkorIoCfdtjQPhjcJeGugypIL2NxK93AgemZ3cb3Yl8kcJ
WD9JGn7C3JkTh23HFMkTy7uz/npe9QCqEGbGBbQJ6whs/6JrUZGwftBtInZTDp/0yXZmQz+6hcV3
zzS3yfBzGaeQ0flnoPqZj0gSKfGZBWyQAsojWkWBVQdBPKn259SzIEmPbMpbOFH//aLvboHW77++
K+tnda6CV9J+QLs4qx6WqdgUL/k4m5bfRHxJnopXZHDeAc7ezQ/vBa6sqm5bXML2B94QSwubovti
waYilF1f5bQeTNg6SHIVynidaSFiqd9+RnBZ3MzkNaQJGVBUQehj1vfnWxCuPbg4cquSJIBU71Fu
5cs8wTABh6s76B3yNLqhUpaSr6XsD9GD7SNTdtH6zoA0TDhgGoLeR7C9Krxp0+CJx1OKPFR+spVq
tPAwZh2no0XZ7IAavMonRzwMVXyZcqDD8PPKXKfYWHFf8n/xBK66x4xs/gBtavGZzhlJ0icml/4V
lqszGm03uCQWmaLWmu6gqbymLBMph9i4v7wh9aL3NcKBYQNOAUG/5j/6gTgR1w+pOuydzFuXVnwE
iyWAmDXVa99wpDKGgf1EL5c4HbbOHQV92WxOVACxMPehkrvDYLXQ55lqfFXZXyqypTFM4cGo4MJo
JccRMdjgZVem70FOhgxFJCxJLWiYGmDwXsr1VNOqhYbecFAPQXRnIOj85WGJvzydPkDk0xLDkvAr
e98qeCtO2vhPxmRs5MYL2gsbSPXns8GWpOWeYgq83WJRyxkeJdLjtMze7XuwJRxqmBNVXcOuSLIo
cBTNJFHsj/hWjdbpEn1/6dJESnAIytZC4vKGTwyLqmvCAwrvZZG9+PIAxxGkPIT9mF8Q7cpcdExm
OacwhUORugCdtZTf08rRn3j585ZqbKT/edeFrDxZbkuZmdhn/batOQHiNgPrxeYXfrZVvoUlnhAr
15aMbQIEka27955Lc4qY2HZDrMtQkk5jm2gEfoHW8MTi71RA9jV3JDWR7lYsRN/tuJEobuIiLuIm
WOsfe9S7Pfh3E1OQmR2n36c14mAW8//WTB8t8/3cuPQUzrj51aYfdHAZozAN8dXxtFASzsTcPoVT
Tp5qlsBVelA42OTCqkvoP3kb0lt4OSLpfmPm60A+irAfI2evrHfIL+ssWX5DUis3YWUEOVASVxp+
y8tXvREYCkGZEi2dKKVCxYHij/V0VepGppUCJHJgTPt/Pd7eBOfUG3mgQBDJ0aWFQvm8JvVLvHpJ
IkK+OhueHPLMVREMAyKnBvH5hLPSnEDS6nbnPebJp7N4PeNa0tTzB68EKFs25Gp/ynQsYrnv4EEM
ewwAVX3TSZcK2wB41q+vyNsVXiR85l1lo5gVZ9qGJ+OPUsaWDwtRmJWJgvPJWaKBoq6vWhzm67uo
7OAQTCP1wqYj0YH16j+h8N/iVqFFPRH4b9wHZtVjlS5aX55IbJCwScfDl1eZQdiACaOZlymAhYah
7VYpFpKEaaWPL9EnzUSH1bPyFnkF2CbyEoD1cqGWUK9YYqo/xEKttJPPmUPb1cpCujllL0p1HUV2
RDt2hacEkhbjey+ckFKou/jp7xGQDJDg8IUBYu/e2VY4xPyFjbEKC6vUG887SLn/Gut7+IqJ+/Hc
S+E+tB2Fpx9FlCs+TSA4d40p+I6uzVnh0Uqmfm77teTyfhQaJyUxCO4f7TjRVPDECqIKJhlfWPdE
L8jVHSNECGdrmcodqiPbzQM8o8KTG4UFktq2Tmq+/DCkxRMUki2n9aYNOLICsNQ2NMV5HwCmhLp2
JRSEE+mz0aUMoDnNh1IT8A2w5aVtMNr/y2lDcJ22nfXmhHW/TUolnc8FbwWoyvWTHAje7t4bfeli
s9D+hbqgQfs82qvVvHBy6CPlekWfOLwTgWlu+KjGj55YUuVTrT6t++juBCquewDUqql+fys3kRlP
zreYkrk6LWqLo08F8X24cvT2kzvVKtk48AJbBGdwLEm/1t6AnvbYdZfErs/M/cYoJVyC2Eawvl7l
vT8Ypwg26fIU429mTQSiVCE7roXRjMIHpvRS/W09xnYeve5+78OORO9NdyCnX1To9Ix8Yb9kTLPv
yDKJhD8XG98eXyVlZ1v17ByT3XiN7Ovr0e+S38Zfjb4WZ9YhG1V2GhFGRDcuBbZThCGktB90TEhn
JfdpUDJ09jPewZ6uRU/3yeHWinKiuOS3xFZROiq0GCniqUwi6hZfXikzDW0mubg2S0ZcEwpQhxHM
efDMpqUeDSbjk6RP4kDaq9NK3WVLSkH+ZWwjibkDntJLqpXfnJEL4otjqaJ6Nrke86FqnyDLXhk5
vR3D+rKU8US3LoHhvYRkvr0isWARgJqUeAgPm6FB4ADgKbO+qPlkKYcTQtJMEc8zLKfEZ5dImotK
338SSF1we/cIjC7EJYUg368LL0kzoFb8vHNE3mfHO8IrQu+IjLNa9Dvn3HLWhHJXMB4ms7jJ9drT
nrm6bIlGv+5OP5E/EWYoD8XmouRn1xTM/1VvDW5rVkTq+c7JLMlIXv8A6KPzyykSxLrsqRyfGWqv
eaSDWNvHgcTBUwZCD0eaMf6T0p3ky0I6DcbC/ImvSI/bvAy8EERwztp43Pi2f+LPC0+moIoZH7/Z
EdjHdSrtgP7arYkfL/a6rKU3YDxTDf4IdLV8607dkAsPbL+qMMf4HxaYkfoqjjgJvAK18oYULwk6
3PTOXrND64DxpBsc92rSKFu/nTBdNuv1LRWq3jYQsZ1Ot/7tcdmOi99mY6Flv9TcAk6jOE8toq4Z
EYMCuva/ZVaBxMfjT9wAR/X/WmRUfy4UEKfrUmqUa8uO+pnNEJt6NJe89vfQ8NJSO21LFDPOvtnG
TgPwsro3tjMecLKngel54nYywYi2dRKNZ4c3nv3G1tNW7DcKOIGS2jJCvSxkapePCP/rYwneWd8u
yL35CCdPC4KwFWcHqKCH0+O3SHsTx/UpNiRKSdgBFOAWiqOeD7vVps9PQaS+L8nx64mfPzYXP9RO
UcQ9NyN1cd3Osgbo2FMLl/4MDPna8JO0UgKiBEZUyqBa0A0ejfoTVsF7PdVzemDlwcf5bU5bWZow
eqQljfJOYywx3lEmYRyDfxzxwJ+K/Ouna5mfZ4WCG/AYBA96xKsyPA7qCxo2grT7vc48d3fsL25c
46/dgxjzc3sJOvColt54DSmVPAFu9cWFd/JdJy6e3iQhGeU8hr5aZP4obr4s3tynORHrSFZ6ZnB4
G0oPbqVq1eH6Wu9+qZIdeBm7kMNSh9WdmcT8aXkPfOXmsrmQhnBSaRyiz7xOQhatCTIeb8JN7Byf
zT+F9ovBLt2/p/+KiL11G+W/mpYL4l3BmmnGuNZHDRls2auyjlcw0MF35sQ8s2gX8PvmPAYsz/t3
WgMNVTEQZMffk4i0hCq/KAlBYLSQ1wyx3B8Nz8Q6LwnGKIUPMVRrCWyFDidU0sc4aV9ZftxQ9bjH
nkatTvf6WvIBlR8fWepH6TLCzDZYIcFDg03VQteQ3JKuyVaDP+IVPC2ET5aBAvt1QG2i9+y0xeNI
xv4qoPLSeRj1JvkK519HLl9qGQGDyZwvATNbBKpb+0bn0rqPrWp0WG7Z+tPGYwV4ZVCoGoWn9z2s
iZvfvLV6BVRn8ilyh2csv2oaRm262+0LOdvP9OarGXOVRS5UbP9XNF+9BEThzXQqtspE95BOYT9x
MKEWAxyK3aMmlIiwS13BhjpjsVGce5uyi27zNs91Ftk/bHTeFODgVgXOdLVXuaovCIbDGnmZUp0Y
Wlt+J4tBwDh+VeCi8QcfLq3uQCxuTQEb3GuW6HU8RrUVtvTomJmHWc0LcuWeXHq0fX9KZTrB+2+O
DvD9sK6dPJ4suukAW387GCD+BdePSaKqdWBYnKPAmuGxrbsGjA84nY36TfXT0JyFzmrmfES6L1HU
R/C8KHXkv81xrbsuws6jAlWoGs9CFIXBzgAL6h6UrT967iChkDNYWXwcaf0vyu11ngdAkmnpRz5O
sP3Chv16MmCOgpE/wtOMGoHOo9upshpiXB9R5IGqgpEiY7cNPzzWVbcEPDpuu7mwI9MBGMmDs5zg
Er2w5KWfIguVDZ6S3BRmUmJR1bwtx7ctZbyaTY5q3s+1iwuUu2X2pKSEKMzYsofC08ZFzy294J61
e08XxoDcZQeuYFQV/piCOnFj48tj/uVR5amrmMHVFUAN+eWbUyg7efw1Q5cky2VtywKYNHKsADxx
l1ONLUDWl2hydk1WHa8Ru3BVxl5P8Hk14zJQw5VlSLue+nupUP3CzryMYA9/a/J+nS+TTMdPOU8Z
LRjgq0lP617zjt4NdfwDbO/fs9JpUn0qGz5KIFAVEW7wQEWg51JdAq3pL9EsYqqw8vziRenumoGy
DoxPTlMJGCQQ7HFmalrmjrYbnFTEwTZovGfYBY5R/SY3//4OL2nm51ReEZ+yfxVH7VLOeoQhExpw
qK6VNLBML9zSTslwqtYJwrdaGzyxbPkThvQkOeX5Q4uUMlFb0CudAELaFJMC6vxklv7Dl4aIeYCy
yeBHMFMn+FFEeNMqKVcJXv+/9Hf9IH/eoa7fIYhhgsTC7aFxxmPrNVfzafx9aIrTIJuz5lM/sEuY
JjO/r+5SyU50o2h+32U4byRlyrVMPabUKkPaQIWSDvvGklwv1ZVS93ri/7x9mMtSgIL1V8cIlgTL
B9NxiEY09wiAaRZ1j4gwD/XVfnNPr1crYXbJt7Z1Rkrlz204WoTQ1Fg33iq5jyJhLjcSbDHUAMZb
GC7EvSqEtfaHZmNi6mYWmc97xqoNH9paKJ/8ZWg0fqHlDyAb8jJxirGLiwn5A/I2N7vzgCN2vHtU
WBYMrzyGDiyEXvAkZ9+UtzVHmKJZPUzbxvx2OM58DcuUtk7hjiA3NGBsURX28HdOcTrAFq6hcfx1
c3j6+uo6sU2TimXY//svCe8IoQ76SAi4ZcyhPKyaFDT6w3+QE4Y7k6fah3WhXmkPZ24yDkEMUPdm
nlw4u7HnlY1g2nhMMKPHZCqBrI/lk965cAJ10g79QH+OiZn08B3nTB81h5uF9GY94zlhVaQwq6kM
zn/A9KXIQwZHgra9fzu0CLVWIZgkOui49WaBPq3cufdybSeaeRlHUgx7Drv/BO3X7TqipribGBIH
lzoR7e1wXd1sAHhtv6bMWlxp3xZpsyU4FQxyBKW9BcMer7SIiYUUS/cjx+l1BgAZo5KeEsmTeBoa
GN/6zsYVQVSO4Fm29F68JvU1cVJBWoER8i4Myr4xHfXGSj1kCGc/S6sdmEqCT348tHgzkuO8X2iF
MxvoOJWnQn0ZNQniZmur7FXhvdc5TJ6J65fuc2E8t3ojF1mI8VwNXaSFHL5D6yj1kjIYsUPeg3/i
IMArB12RSh3kIfOueQKwYQEA8fHNnJulgJhlyJGxFXMHWHw9Z3hkjMOI1Xx1WRWyULoPoctQ8RKz
Qi0obf1DQ9DRPvIRSliKArRdQhR50XnW5tYAWicYH/PTMdnDLZJ3zkwyTzc2ATVOXfZpl/4tXEYB
DyCAgAcqyTpMLHB8w9ID1Ay6Y7iBN0UCxX39LXD27Fp2Q1F05JzzsRLmKgd9CLWnqfr9U7sSFhXK
Q7hQN5elfL4ixzTB2j5FJX59L7rDU1csAZJkk6Ll1MPHDqvo0mrf4Rs82ju/0dzUqOxOG7hoMq8U
ABdxynyu/+S5vuEaPH3GF5zniDQw3RNI2ZNhCay6ndqf92wnh/ISNEFhk9oTTr20OYTtlCMfcH36
PQB/9w8lB+/og4oX6IsYOTk/uqMIFEogfFwdl+ggwM8J6O/fzMu2+VPfdXIu8A2z1OiIJfgjVM7B
KD8e8swPzGqKINRxh60qC0xdUR/HxDYgp87UD6/FZbzyVqSVwmn7dfFQS5Fvac+e6E47VCYXQ4V0
upu4yE/QNmNQ+GPU3iOct07u2WQ6puBv+FuyryCiGLLIq1fjtnRYTSq1/wB7kL9l6IyXlk7i/7HC
w16hsfmuvnpVopeQ3XNdcZ5UzhtjRA1K1QzOYfeg4xXiflTjpsBfrb1Qju9gO3hK7Q/gfKmQK2Ss
QdhPIui7bl2mTO7mzx4jkxc199cGnizrlgQH63zjZZBgbuh3L5ER+8nikS5VLibxQ5BklQf8fh3u
GMopmyKJx91Bwb8tgOKCYy6rLgCzv2vQ+IZZxRMvzQaK1rd5XQtNWfa0XYahMrrxX+JF37FeK0EN
IHLa9LJ0orEbVI9VUHHemir8FgjuvYgODFBPSX3pFJIsDyDk0yknzWGW7iEUPa4gGFWsJi3YBsn6
pGAb9CHk4VZoAi5Pz8Gu2sTgS+XkLSg94OUvS6KsFhru9EIj0znBpuj1q2+cPy8NC+573M62eqqR
oPIqwhq7gr0CG7aTGWs7elsBtFeky0Xat+dZM9EGxpcsDW2X5XAtGs3mZMtMJ7nEuuK0mrbxjUqD
itdL+OA6u6xL4kfJ9CPyX7unQNA9tqhcykwwhHq1TYUVhNEIU11Dlf7I/gE8KSQQiIEAr7rvoRpK
/9WTGWxukHYxaviJdDhO8PqIc2F0hBTAPEDkWE2pwSCPDFw0pkZW1SeIb68pIb7n8dn09wsFsSe5
kUL2bHnFFEGUgasC6pLE1qPoOeF0FeRuEZ391PD4BV4fAD78JPb4wINqKIbvEW6RypkK04hNjBda
Cb/nkjIeZM96xdHS8NXg8YT/jY0GdQ9APMPtRKahQ5be+5Jn/+jIXGwNbPt6mk9QNALtp3vNrTgz
5raFXHa1BulqJRZveX1GUB5ratxq0GpoGoZcopzCjOCSCZ9ci9hy1DfYGIzMVRQe0PwOi0P9wgIX
d+ZkPxbeRkwNU5N88T918H+SH6mOFb3gQax7UWu4aCRV6SKNQB288L1TDjRBAipp2ATlZsGjuJzw
mhae2PkWam9llaY5QZVODImVlqCPhSmEUzXTSoR6fgog11xrQVlQuMJI4gEDA0CcDmxPI2EeHy/O
L3c9n6XcYBUoCX3AikjHCTTWtS7gfNDp6uQB/JDt/fC9nZ1cfpG3nLlDnAn2b+1WHq//GO7P0PfN
rQWE1DkC+ZUYqY7JWjbnrWO9U0FmUZTbjCiLy10k1Ql+AEWZkPcce4tIPQdkQwZ3zE2OhaH9w7g0
/HjFT4ZLMBTSbdrBjh3BAY0bzvqpztF/Z1dp5tuGnOzuVRafWzxdvnAKP+eHmekDUZCsPy8ajw0a
4jXCp2+t3kusg0uZUqS9DF1rcWT3VOYlHjQ8zP03PmMB0IF9sF3UJKJWqCaO1huHCsIKcogcG1A3
HEkjJHDPg7aenqJcHccnLHQ8uEWx7EMyrD5wqiWeuRuohOA6M4C461VBDuMOE0wlAWvx4Ls7t7MP
NZSumkReCH03Tu0zbggfWefO7xmLGbtCubkh88lS1QV7aamSrJSGN4VNU9padR1zWcSWo9yzYXsU
26mrnJri4xzxLoK60TdR9hf+d09+5o7KwxOpiQrWWznv2YON2r8trQh5eGjC1/O1kUBEsetpgoLT
LWmD7my7UxEqgPJyZwkhydHwN1QsbIRbFyMjiC23OocVaVfWvkRSe5XFyz9UW1SIsCBTSdnoYRL9
R6vk7uKQaGW3qiAINDd3yTLxnmdtyN3+50C6iawexLIpwf1AsuVxd3V306rdxcPlM8wCyMavHTmK
rHycp1hrvfWX3TnnJFnZBK7AK0UouxpTCWGoW5buL3/1LGxI1velx27RLhfNXbXZwK9Rads7scd8
A22oWRPb0qGWCrL80mpJSAnVfu8zzwYpU0FMLXms+OLmzPvMn00i7QZlKhXY1PS3OiHfjg1MXrnM
qNA4HCW8djhLrpW2b5uWCmI48kYdPo03kvN4Cb9cmXm5ro0oumj/zHFOh+aIwHKPrFd93dgtRdvB
Qxb00vGrl0vXDTmUTRQsHIjODxQ7O16ZJiM8RuF9FwezxP4QorLzxSyofm7PGcljA79kBzSPph8+
aT/0XcCDWs4x91IkR0MpbX3bidTozzs2koYuyT4IGPiarpgp7ofirzPtYIjy97VTuWLpUUAc4OlD
r8rn7e8MjY/TKc9rsWkwjYZGuuS5v81ylFdkyv20e0NaCuG/x0Z31f+FqfSjZNNU+Jw0iRlEQ0R4
l7GGGA5ENrJRe9tMd53vpJ/XtBBFxyhILcU6AJyAOP0pzosHOltbsYuM3+/I08bIBC/GD5gBQ2eh
cnA/cBzN2lLScIrU/CF+MspqnknCDFrNqbH+upsOtXrlG6AlVaa/KNqfuK9HIgbVtW0lfO4Huc+n
5Ae80rFE+Q5ZdjpD3LqJXNZ9pr9KcU0Eu/bJFFIn7BngTlUGFWp5u62I1FaFy5WWlcUtqgV9I3hH
uRLRRcRZpEosMGUOA7OfzaueVgLASnMfgD4bAcZtsMpRXMO9LH7uQB2/BorUk6tdsZMcDtcmQtpC
yFZpVsn43gDd5fAaOr5LXdBmIe78TWCcfSls0vUzi1XMZWiGcmdD08MdyLEbqB+EQvyrv2DFfdLQ
hoSzOktFwRt8L3JkvzGGML1WQbJOv6OnTgB5atdF40TRVc/fSzNoSR0DdpB4zmD2I//Bkd7onD+J
8m3qC43JSz0I3mOAoqoWVwtAYf6AhamyqD71uGm/0jeYF1B5JLaMaYdUWaFrfZ+hVJzckVJZVtkz
dhlyzqCG7Ui0TmEhigVuz+vSBGOXmwkl2UyQ0qhipaSXznppvYEhsd2a+z/1GPC+Ke5NNnhZJLp4
JO/tCUYl+Gth8JnBY/HWmLxCZPKo/mc9yPomCFh14bWNrIYIBSSuoeS8D8OldAHymmRPOYKQXtgR
pZUMKUiD1J1ddHGJTdVgnosOHO5Tv9oEJ8v2uyzaOESMC/AibXkK33HN0enr6GBN/r/Po5UMiIEO
Xj3Bmvul+tsmI8EZRRvCfSpDDYW7RfMfN1eIao/keEEpZU3VJO7K5KdAyyUm6j1W6vglsxnHEukw
QKFS52+1mJmanChykyeiknl57xVeZSmyP+lC2AEpuGDhENt7cMV+iILENtLSz5e27Kk7PhFblCzM
SaRKjVeAQsZntDMi9kx2vXkiHcAXCIxlKlz+c4KX4VPdsb6cwi0OmjYtXcgKEX3nYmB3aZg3LkFk
wic0Xl1H6tfm+kcKIjcnL0vyZzXTW5q471sXAAm9QScIXuIrOt89YbBWR1AHLMtlUeAsWHtPlRwT
KJP+0hOf6ySLJPfabH+S/4IW3nSm08wAIcEdnIpVuySgCJpkZEWRWnTAntTje3a/6ZM205tu+6ON
IR8+PnSjjAOndLKVKQejUuvAca+c73fAK/W39ra5ZIcvot+MnrtfabpRNmM2KrD3chFLSHmTwe/f
ORIxhrhLAYa927pcX9Q3xpDJs609QYl0+mANVtoh9L0iQ1B/Yd21zjSKg+kwnwdXd0/uY5Hi2voU
8qt9+GXImshva5/bU7WD6b6ZXJJ/gsQcUNeQWDfjaDBq6uvSmnbcjSq8u4QrTsg59KVgOrz6DrXL
rcT0oqsAyz5wWNvXo/wiqsLMGa2jRIMDDrsipt2/atH+WZbIYDLlVKgiZh8BpdCqlawWOYV27u7B
zaDFX3FZnYNkXScO1aykNusoaLxcXZrXlccm00Zi1s9efg4t8doJdw402QKU7Jpy5QoJQxLFlLLm
0VgGfl8IHltWh0u1yeVSTJNnXQlUIro8MH6WjhpK+5rZ/FICbdw7HTkRdffjDu3XjTDJo32XUS/+
7eYjS3SbjBeafTf6UqikfKpS98B5+TzJoCg6nv7L8ttBO0giZX8aFtdPX96Z4G93HOl7GBU8MGIR
8MkMI1C2FCRsDj6lCYTrpGgabpmqAkFTU5ZmcMgvrueuJppVRNg0y+owxL/Yw9WDl/wyVx89FHOg
kWU8vj32RoGte7KL0z/1q+zw4a7hiyM6lAyHbwmQqBajKiqjJGIE+qLmuSAPaZn+XThRoXGCYLFn
EFZhj4KFofC6LItNV8a/SWr/X2pFUN46EQKze7Jj63U6B40drVkAaZASGtPxf7U8m0hGJ089ZX0v
TDxxh58FWkiNNge/hUA+0RgZMI4S8v94C7Yl+hhhd47MoCs4CjrATQz9HqvZtQ0OxXhLkZxk3sUy
uzrvJtaZKvo8jTVcMCt+ZVWmvkXDPSQwlDAxtjvABWgtX2TO9do2MKO2f1RqNK9qiqUYFA4WCata
XdQNr9Vxe1ppkWqpll9QVpWjgb/w4o7VyQIpdQz5pZR5rhDxkvYC0gS6SYumWHQkXN9QYZpdABUv
Wi4yPlAjz/hYdzO41OasF4g0pxScjOS74QgrTmXabjXasSuPygNxZPmqTihGRMKBc1sIHBAoFOCK
Ayce6yvI16nqDDw+PG24hjoFNFRii8PqSk3lfexnXBhCvsZQcFoQ1tjz86v6g84kSGrHks2htCit
4BUQSu4jo52FwQHzymcp0BtBhkPbiGywJLsuhemJ1E9pf9ZQba7BE+g7QCYCr7qpf1GxKs+UMlED
BHxDe0fSTW7nXVUEN6UAEMlU1+vWrhylIqfWq+cJK8hkrXXx5QQyDpFeFvlpkmvasI/3UY3GOnC+
3XVwQHC9Fu2q9jn7oWr5QLolJGpd1JSyF3VkoXZ4cvVwFep+7LxhSnoa0W8GJC7QY7EFEJ5TGVeL
Hmwqtb2T73QQG4SC9FFnGD/CdO2XKDfEQmMc8NEO4uQbcyTt+9cEWjLbb/Rc2KLHxsQswK94GsQB
1KDo9E075RF+n4v0Ifs19L8YCf6/0KQ97nYeYfFVUDsQfXPecqKKadGZAJiN/Nvj4fJAHmMxCc+S
LJ7Fxm1LSv9uPTCrmv+ZYKjk2vXcMJ6Lu13CCAdAdE+uia8sCA6IRJswMySvl9Swqf43LZrAlVde
m6h6qL01MokJslTKQR5j/LPbkDq1B32Ow87GMC+S72SKjFD+VerOhHPaBnk4npjy8I3bFF75NdFl
4+iEXc4Anic1n2OzVngwqQE87dMMcHQr/wFWd2QOPvSxGnyMRF0aD4rW/ErPiXfwsYFcpqr9EVHK
xjzKsEVqJBjo/xCev+5FLSGJh9NJel9uDW/h2NW7rGhg9g9CVOkFOcZAO+x9FZbyV0es2zmGgN7+
LJiMK0bX9Mm8ceUR5AY8fTDlijZE0N8M8zSFYET1ww0a2TbnHSXbikBd3AAoWRmsib7Ul0I9QgvI
Ybuku/5L6lcDRR4sfrhzsAEq0I0VERPOZPkDgHt9A+0iBW+eZdrTRXhgAeXmEyLuQeVmA3DNZFLK
vUHkwbQbKDgwrDE+f4MlRGcoezEaMlffg3lefWRnytuaFaAw6JVl1V/i7D5Npf6ikGmBrxcZuIyW
+bvzIQEGYEbZmWGyzsD+POH3QqlWuskp7RMA9Hj8xtC9hj27FCVigsrtij2POsNDNVzHPNhU3oMa
UynHw3PBDwtsNs+6mUWzE/ulIY+LvZ2zg6evmPHnyyY6IfvhgI2WfmFcZUNB2bJ5pZfLps30M+MC
fArW4fFgQHAM9RDofc3hAXEe/DqCqOsDU7m4a+IbHNMS1D8v34XBhSo1bWrkxEUbLMlvA9OSdH1n
SzxkWDEPbEFvCTlt522Q4KWJ3wblm7fwBSGKTMro6U1rNY/g3ej0TLeNy3aPPq+Svai7I80ud0DH
8Ti4Tg/eC1YkxgfAwaeVMyjTSfRJal2bPfAlUz7cd7yHcq5Unproi2ItPYLU5HsFf08aUIc58QdT
AMQiD/lLIqXymC6B+NX1unc+P5HGdK6ld0r+ndHGOX74wqeEX5tWdG9MuJI1GTs1c5R1QiaeILtJ
e9oEXT02NMSq6JP5jzckMDP0+0oMhdirSuAoCgAkA1DpnSQFppDYKFo/6kv+zAkO0hTzY4H3XM88
pagDRJw2COC9NwSiVk4KZst34LikUFfEAIed0fArPWICWtk9KkXct/N8veNo28jJqzpJ3f38XZs6
EzNgD4cXWNNYLzYclZQXPliL9RfIY6MUfRvz8eMwDg2pTcc3Ywmg41TbUoxBCWw8q+hd+3oF2aVq
q6XOBrYP4spXmDZ6I4JiHt4y3tZb2Aum/V+0yvoHtOgSLUFCacIA2dngrkH1yX+JSNahb0IddzZn
hYGneqPQl+E/iju75NDv05+qbG6qBuc/+60GVksWloHszFeaV8Km45CXJrHEMX30liMQPRphH86w
lXokbRdUnj8wHVUQO7wrH5wqeE5ZGi7G8HYcIxedyXt4wzrbnqNCtrx1FH0golmYhGqu8rycOXFc
/gsRXR31lNlgoYKFa2LvJW4uXRCRx9739QA1oNmNPczolQBFU5WHggfpuVIWX/QBwb6UrRFxOU/+
iMuszF6uWUt8SwyjwxxqRLQaLk+1rJ/2/e7AvRrAyGR2l2NL0Qoxezi3NcrkBtYvrlLD173tColp
fGU2EgFf6sM3941vuhQUYrRWSARiAPa6vNBPcmTJlND+S+7iCTocmz+WnK0AmvIXH563/T6+ArxJ
3B2ap7/V7har+/GYzhYkxUtQJje3p9CGzOLQYkXvFlfxlrl9XJGn6t6vgZ6McwQSX/dvZiJ77P/v
yEKyR/t33FA76+qK7uLGsXjtCrT/NvwPn+Z52WJrxNTUJ+o52W7N32OdSBtXVxdLVa3pH9Ek7xje
Ig62E2mCimWroUBBQi3zi7CunYGtaA9BdSfL7yl1AJtoKNY6TzVzzJA30mhcPmBKDJkGCf4kly7q
2bKXKtSktxCRGJ7rWkcf9Iu8GlWAkiETf8aVT+nYfTuBBR9RfakgpBqHkMCfvNB+T8l0CVpYV6H7
HlZfoM1ceDL2QRF1Addz5T8dwgj8wtxDu3Sn0Ju+6o2/eP8A8VdLvJ0fxMjlxEAFl21VEKSE7nGl
GJ/VV+MD/k6WEJ0QMZBQ+eJG8iz20n9qNYSdYRveTvNeIsA2OilnuhtnDGxa+E6ZkFK+7R1bUy0S
SqT1V3rURH8v+ToahHHx6k7Vnodb/U5CV+40c6bZZvm9aEpN76pyzf2g+LdfFtXJgjU2kGkcfyED
eNBa/nWZslfY1P5sJZGWi8iFMchq062+W2UYwHBUbHXiAe0da+ZAXD42NoQxR3dv1P61XqxeYFCS
qL2twrX3eyl5dQ/YXVp9W0p8W2MkNKDS8SaeWK5Ats4X+Smr9eVWCPI7pB7CLog4MtNrjCOJCucb
a5c+XktL6ZAv87CoyMwmiZ4WA14/39rmNc+wuLiiDWeApCT1Sj2KzbmTWYb/0HqrUAkeoS6+rJS0
LZXg0mA/tCOjbYZtRLW2P0AC2NzFVD66AwN2dHwKd09ebgRjnGSWoC4UgdRVH6nVu9D3BtPrF3eq
HnlBXAge2YOc84QB/41rEiFNnUIMNpxsyJbbgO3WFl/ZdODpT+ewXZKkmwT0PD2+L24A6onofpCj
RpsnJaqjmFGlBRp2dqo2omYHRZ4EZXZSM+ZxhKigJLuSFyrAmXOMcbLaW4VaCrvKV5XOahugcq+M
XkL7cbGIz8Zld5gOf99I4ub/Q+q09bz5zn7uYT3v1QEePngF9/cmiZjzr7piatq2aO6OJ5k95uCV
9cMcX9az39yKfJGkZwsXeUcboKeiHI2s3O8FHIWNwkjk/wfeiZk8KfiVjuqk+8y9WWCI8ySvGaHz
XtlbHj0vSUq5vD6oo0f7T85p4lLec9sTvJGTzfjSloWPW9LFfBXaqu0RNdr3pLLmSTgx5phYd4PS
ZtLSz8RiCPsWIkt+G1/ImgpKMO/1pnGq7UF+vNRxvhUSD9t8edGok+vhUuEJl5yDZIpjua5OtvTS
aECorTzFzlTEegGVhB+p6iYdTd0zOmegPzPZFWsqIrEiBfoke9v+h3pU/xCPxdzCxSBY5ZabsSyk
laNsJSQxwh+UXgMoTqGTqB96TvjsyMNOH/xZ0Q7joLae3aEWg5InPL48inDSi1L0wEQhPFQyLT1e
tPYyerCby21G8dKjhfd4o+maSAQem5Jp2E5/Cf86olJ/gDuBiv1lZmiCBSEmXenBakwmrA/FRi2d
g/gxaLxVjyXIBc8mUPO54YUmr/yXie3YMsVY0otcBKZ8ZSNkJDFAZo88ks95zjZQgar21R0++OZH
YJ+gwShAG34M0I3jjN+VJ1p5+ML9L2TTrHHQLjv10tsKoqHSU54q30lMOVJr64GawAYdbjXQR13i
BiTiKAP0+rm9kM2/1bZXh6tJiQf+gFgNXEiZ+6qeyhHuLGnTNI7GSPkE5joEGEbYautLeyhFo4KC
FEtG892MUN2/7g7NVxXrtB86FklBbhZT3xGgv5rWa1QyyFq1Cdj9RzUCIY6cEKFJLe1ehaza2AXE
XH4rUqKIE14fP7KOGnDhgTu6X7wx/ts23LGBboj8DHd2s/t9ZElMCii5UMyzH7cQeE7qjr9P7Zt1
nBGj+Vs3VF1HrfQm7AupvpcRWOxjaZKUUR3QsNUzKviakMdOeFR8mxrZgEJYp/8xDxsVUIyuTWSv
g9oDQIuvLqdVe3JLWw+UBnAPFdCG9+u6kV9B0eY/CDVWIAunek469+FGWGZ/HQaeYdfJfM3Fzjyb
b4NHWC519ITrfW8EW3oKY4DaoHbeHXlKZjqbSFbjzsChks+AlFp/rSaZwi61WDk6o3k/9PHcVgs/
9YdQJSKZxyWX+HPKntb5hmdio+PYFLB23uq/0z5EQSXrWddfAtekvuO/2BI/7te4mmjAjuLzwyur
HMgrIcBupDryniVfJQyzDAlCgfDjwxGZWzv0lVtjhx34sYD/Wcx2ir7cMsnyJ/EUuhGOy1sNwXBq
yKIl1CkYsGkO388kOshbngzt399ESOm7QmwA/VNAlXgbKyPQMCAKqpadmR5a8ow1yv20fVm47RqT
isj6vlP7YWMQ8UDPT4rrSEz4wUQL5hM8oLJPx6P/f+Lf4yX232i0KD6f5VprJ6cnVrQyOgsDi4qX
SmZ4A6ge2VQ5vjH9iftFMgxNG0HiEB5uy+7Fi7fS0tLXKp3ILX61FxuL198vfF02TxmQ5zIlfzbO
TuLglH2QCXKac9uFVdn53mC34ahpWBLrHWlyvIcCj5vcDFGhdnA4TC73I/fU7LxR7R6kSWAK5RMV
8M2JyBRk8GnuDXY36AOZOPzt4EhW8l95s9i66RTD6rDM1gOVfaMt+rWbOVr9x76CEzAdPpQYKbTJ
1WHH0w6RWd3R9gM24oLuLC++LXlHPr74SIQeE8bFf46k9HUACGYXBMN8oa2WaH1Tu3Qx3088C0l+
ltP7uV2EbGgWMFmGACT8/dEjyIf7BQdKO7nEvHeXQfFjvT52VkWAdptifwyjt0eTFKm8dRFpTA5N
+cHvu2ewztZCydKtEcwfoYJ7U+8R1fKkWqdJs5dezqEXNSrYDIOxqEcvVuaHey0zVyNS0ItOU+L9
F+jpYJhe5cYMns6v3Bnued9g3FN3/ruhBgoZL3YhfFF2CrtmQQU7zxk4RGPt022TnNRwW8BzbJb/
NrPRX5kVjxcCdgOHaWgaB7UgpOjuNzRcSpkY/bGxqwycYDoUggHNEsTmEIUCSccs3gYX2tfadsW9
qEJUNqEoX0MFmh9VHEgIEyL3rq368HjbpC00M7Ld5ZaxQ7J7uFz5a1cW18HY5+j27oMAibvcYHSg
QAXVTy9IRxAO5pnz8Sf9yqh7HdO6Oeh0bc38P1kknkqW/BC/0G7x/tLynUI86mWAUHI55lbG2N4a
Zi6+SUQQIxD8vTOBrj0tOcwzyl1j8JTwgE2sKTru0qqFi6hqu/HI1t4Z1wVxQnuQqSrtxv+bBK7n
7VNrrfVf+wMqBO0JH5lxoTKs7kEwaBYXaf5dQpC+XPq+BEHBgGkCNZxdX4KsEHD8CgFgZkPmyI4b
SZ+d2hhVidFtudSr8Olm5VCtvrsukFIZkXlNS99qpGfoY6QE+3/I6gql9qGAX+PXnsHdweYDh7ne
hLUM9aIl0hO0rjfZ/IDOy/q8FtP+6858m/rux6kZCRwgtDgES0drP44rKUPtRftaJNgWqe5qyg51
hbMmXPItZFyUiAGRWn5zXMbD/Vow+hi4rqje72Dqr2EBoT0JIhLvtfak+9t+dcJ61zJLgwnRqwyI
HZNW7/qvUL3PRytxHvbN1FxdC2lZcvy5NPKjerQG1BD7WbyJ1L+4yvwtdus+uaq3ULnhkY5aItys
OhpDnsEsdLIqo+nhoL+7eswSIw96eEQGRwX9+AfKyxBfHppLr3hcI3qF+bgzZVi/hh+n8y6Lq+4/
gMSqNiu2gOFVnGWb2uvyO0Sj9+OU3QbPwStBJZWzP7YdztkiXYBfeBYzL6pMyNewIm4m4pssRytc
GDT3V3eOWfcr2RPyoUev9NH5+A0FKfDQFYYLR3C6C7X8iTFiCelgO5Rsa4Msvd5MEPNIYU2TBkaj
+x7PQBU6ffXBYweT9D721UAU8uNbzxj6/IaDXPDUJSETQ3/GKoLvjszgUIVHtOfIut+2Frh+lfOD
X/fobxkdUIcjd04t9jGSpeX9ko/Pm/Il4rvqHL6mtEGMZI8hR8ZJZKR9nqvRa9PYc/ccXZAq+TjU
nNuFgpkmnCHNRMbQ/Hg02TuFuS5leB9TUPUeKXB2qSGDLxlqKkS5reUfQdluYgS+IXqtSJta38jR
/WkauhgHJwBM87EGLOmbySBffrc4uBxmb17ZriA8nsniicVJ67ODHx8lEeLJlQMwHAEmBr/93OtI
8LqIlLssNHooJhPFaUnxl+AGS9Y/LZmr9OARtyuCePetLnI8P/JzrzedAgYYGyFvm3OHMpJq9Aog
jzFW7YtYXXCrnJ3SnI7wEW73p/Ayw9P20WJ8eggr+voEAZh0G3PerAgN0iJz3TlhFZXBIbvyO8Ot
v4vqSqVbRU1iTE1lV6yr5X78rmNU88kzJUuQC2IRyqTcLuy2H0BmKj8j5i3W25Kt81FzRcZXZOU/
U33VlYIRDjt/KtW8nK3FcmKNuhzE+XhEKJonNe2QHmiqQIb0pJ/bJfMcS5yCaR29IVG8ZiMVrDha
DXjFWhd+Nuh6aX6gBKfs7+omGlOThfh6GS3vdslSOP0o+3+OESnDGZ1Xm+wGku/HINYNPvmAzgDU
A0NyeIrNM3QYbAlpZ2k91rLMJxJcrfnO0t0gNFQ7ptMne6JkWZwjDhb44bA8rkoD5xWgKEkiQvKP
mih7EbB2zpHKXsuR5Y9bOH2HDBHKJ6sAUSVL35OepbqRmJucvInXrw2vPBe9BcqD3c/PWJhjyoNA
nl84Y1MGajmZiOGJyzw3xiEFS8tcImcVbE/WCuQMjOH9FZs9sjQ5hUn0pVCl8bE/PeT64Asmiv9h
tQCV2VLtPCW9IpsD/Lav9UqDDtpQM80C5GFgc0fnQSoxqPkoSFzOKnSmNSPvYaYIQeM5eYewRhhj
EA0QniMTD/XQcOvxCvBYNarArHJpwnx4mjPt/r8tYUyB1RX8n9PbQCTWjnP8a64OZTddxptqqBbK
RPZxEDSz3x+gzvymnDTUHQO4FhqS19N5Wpw3OiL3MBNkW7hBd8VDfUhx0FN+STTk5vwvcKd8dk++
ePlCo82TEtZ+gQ34NyGvZhKEQFhbmAxrQopVvX48pLj4wIr0O8UDOkgCmw6YbEdkKkbxrY2uJUE+
tMYDM4z17zYLX5Sq0jwzt97pbneQ0GkPXPU/YO9wAuANZFNy5pC1Q7py8PZn0XHlnWQgxmqmgJjQ
7SdrgJzovD5cv/dpB35jkr/geM+Pe4ZuT11FX7vOQJOJjgcR4we+FSERBaHRP18ANhOaBjZ5fT+2
Ac6/6ld8pooc0g5HGcdTeursg9LmTKOCcZPhJpDX4UNE2kLOGK1Y5EPhYZPTfvFomI5Yow0Q/f20
bb9N07N6fKBzc0BXuLw9gvp/frEhGInyJu4sQEhZkaanYdvGyoPqJ+n2nQeNoz3JS5QEEno40g00
1H9X1we9kDSiQp0l3kak3pYEo66PUw9R1c1yAHd0bwb2zchX9wu6iAUKNSjqeR4+7zcHpACfbQSD
LaLNDYjNCD5pXZ/dt/QL3ETQwzi4i4Ng+gtH2EqYDacY+jOquPGb0vo413uZZZQs+1o/vuB0evJd
LDfr1WqZdVZJDMdKPUwl7G8vNsm9JdSkeei/1GN9oKqUHmK2gV1qzgwMMRR686a1BFWrBX5tIGKh
NYbXPmmr/tCtXCKiqVHAnjo7G+W53QDQLurE3O3x/69I3fIGk21byHrS8jDB4kSQb9aQ7UxfVHVq
TXyndkP97Ivx33G30s4+gSe1rvS00knWnhcg22CsMPMpm1a7hXs2TS1zcQKAvofhlHXQhBro/AJb
Qg5acPZJBQXwbZM7/R4CVCTbgiFSxkS1dL67Yjh2w7dV8qZtMIUsGoJ/UFCeJUgHpcogbsTPrPJe
UwTj9rlhzlFZes4FQ0fVeByTlk2L/TwC73VyVZjHd0GBUMf8SAPegDOwhJW2vc8wRjj+14rluq0X
uiDqOaFKG1UGCYmnRdM3Yr/7zyo9rln+qNn2MzTu+nr3kuo3zA7xUD+fN1H70G/QX1Plh2DPQ80q
Aqnjp1nE8C+uIt845BeWTm5u69Kogew3WifmJIBIYx4Kpl/CcX3XoTREibvrzR/fHRHahPnu758N
Blox5y/JGTAZPGElIFoDW9IY8JsPq71FrH9ZRa/EKiSzGLu2TPF2NGGhku6IPtthFAjDFkUivomD
Pzhh7WhjqptzCE7DyknaikktlWDrt/CDU8N1ZZYlBDPkkOJfXNMvJTmBNnGK3cHepew6Lh8LAj5T
hxhk9cDRC0JSopVB06OxC0mF6eePaRfhjn3kYgerK9qU4wVSI87+VYIvTEakaa14X7fyKRTc4bcZ
D3pOfABjdl9CKXeJox9j8uNUEInQ6tDwKZ39upJlJkBCmIXM9UH7FbVfdnj1VWGEbcqSV7X2TO0o
WTwU9eAO9kBKN5UrkXJ/fRlC+1ZxHwqyVbWmtDnHYvCvG5Y9UBrBRVeVZgjSz4GbUYsXK9AFGxy5
ysahLWkCkgW74P2hUbSAsAkCYbEtko35NH1vgfjr0XeF4YHTx4dWjyOo4ac7bCp0EycTptKw3sA6
JI7TVYqmTDrarSy54WFuTCCzaxtBkv/YG3EZVCUZB8HqjwfX6KCST+U55onkAB6dmmaGyFAsHVRC
J+dohyURyFOLQ9JgCIM2et6zhTQ8YgbyhGrxOBowHmOqTsTNXZVSyBsoF4x9yivPqTn2/aPUr/Mx
j+5hO/to1RicVKeJOmVwuesQG91aGeYLDk2a7VWjPeCLPlcSg2bYndiIuhOQ4coxiq2akNvzQUPp
PPbu7mEKlCmK52j97ZBr2KGssQYTKp3iKMISy38gPz+fRtpU4EI2n5r4e0f0eSTRQcDXR3hhIbuu
0VMM1nNA5R5ukQ3G4IJ272A9QMA7llAp++pLeCkbYo2gx46K0zUTLguVASgcicwfgiWbAbWWUqY0
Dw1QxmFlDq/ILBITCY7IsiOv6Nix33ArftzfS2m5hHemHO/SuD6CqXvX2+1yp8YGN26IqYZxXqNb
V8C1PTp0orrVH+ZDZZl5RH/YLZWHWWFKyk8xso+cxqL+OUFsLNSz/Y3kd63bHb63GpmP8Rl98rGs
NeEVYrSRGkSMY1S2DgFizHDv4a+tDnHg7ca08rcpnTERDRznYqNqeNgqB8gdumwxEPZmyPf3KihI
q/wrsLXVODaDWttGkz0DKsFjHzY1y8IKc1PfAhcFAXyNiM3RLCoHM5JZOz1qWzPxdJsWr3xkwdQY
pBr8tQj7XQcaxW7UFDlcsjIJG+6kjsC6HYrdwpqCJKDksZgyCqjtPu8WSPixjyO/vpypcGIobsHG
9bSjNyTKZg74z3XPjsKRup+YVeLEWkxQeJ9XEhEVsNAqk1PqlZuAZ2zAd7cFXYmStw8GxZ9P2B+C
cY1li93XAiuU6xqyID9xzql5WQaPVKf+XbGQhc5aUWIrmfy7i92+4BDd9WsPuivX7BXoQXpLJqfg
l3GlGpwVxXAQIp9hN5p0IwZe+WlQSnOEcEGhjqPMuzk9CNECShDVzK8refX1ysxL2ZoYBLOuktzA
hZgwK7cmn4Tgyx6+RgPlURRbFyYIyvUCFRrBjJ5UpIN3VdZvln1Cwpvdg0UK6vanLhoYLTdSL8Wh
NuW7zpD3ClxDtMI31gEvKF6X05kdjqZIqaCw+F9Gc/Yg3O0tt8tuFMPFzKdaC5wCMM/m3bprAfY0
tbRQ/dEjoKAB8YSDs8HAve0ysSNf/uhw5ME5oNB0vQ6MdvVYoDIrthXYt0mTuAuWB+zma612BsXi
GAFpGCWzAgXbEUm5LcU7okoyS5AWhG3LM0AUsQfQhmwyeW/musjoD6lSn/H5bp5ttaAuiaz0BYZK
dgk/9T2kvcsYEvjaya3YpFIxsXtNpoSs5+rd3+cz9Xzj3TAs6aqLbNe9ZH4Ev4duMbtToZbtCn35
fCKgPzJjgf9ZHsuyFnDzPojv7XpQns5dtfX6tncKzjDpsDc9nREKZR7SB3F8IP3K0UNHPi2InGuB
HQXp9mTmbLEmkjFNGubQC3a/yFJTyxoo+T0KF7plg9jyAUYbzM94DvVfd+E1oZJ5pbTjjrJFX878
cnpaq8BDEdXqauPbokQ4Tmq6Kzqw6IVMIoHxy7EDedSro8p5WQJ2CYNbLfOIO/9TQ2aDpQ1vlxBc
Bcgt/35F0ORAFkp7e/UhzQ6GVJ4Q6qiG57OUZDFqTUb8EchWxd1vHsbNM7dKzYbjm4nY2hxWsIfw
ecttWyNH5dkOeSB+rTl8t7VJ+vi8Z9JVv6sKNz7DeO7l7TukBXlKWUkPyOs1oGtrLB1NISCQBPW+
E3Snhw3u2wCvryLQEGjVLo+tbhbdQZ960a181HpYKUL9s0h63nrwms6nBE6HyJV4lAInIcI7Vjgj
o+L8DNRApdiWFAVrJu6gvFL2dP2tc4ZS8DBsO71DRSK8VDfhe8F9muC1ugye/QtpwTsOOawl4huG
rY6lHXjLosMGMK1UELG+KZmQmWJMkuh0HjHVGXSeQAxTD5ZWpey92aPOYXOAqBdp8tMJyko4FRlp
a9kTxgtp57oj1GwnpQ4vReytR6xQ9YIDG+t2sQr7PMYcTjtaNWD4GSc1G7M0H75a8msxQaIOInVW
WfuuOtSHxDeDuK2BOxKEo1ZuAd6MAoWsjNZI6uwV5F9QnLtW0oLfDCd2EuI0KQ==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity i2sControllerFifo is
port(
  Data :  in std_logic_vector(31 downto 0);
  WrClk :  in std_logic;
  RdClk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Almost_Empty :  out std_logic;
  Q :  out std_logic_vector(31 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end i2sControllerFifo;
architecture beh of i2sControllerFifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo.i2sControllerFifo\
port(
  RdClk: in std_logic;
  WrClk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(31 downto 0);
  Empty: out std_logic;
  Almost_Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_inst: \~fifo.i2sControllerFifo\
port map(
  RdClk => RdClk,
  WrClk => WrClk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(31 downto 0) => Data(31 downto 0),
  Empty => NN,
  Almost_Empty => Almost_Empty,
  Full => NN_0,
  Q(31 downto 0) => Q(31 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;

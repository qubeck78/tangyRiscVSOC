--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Mon Feb  5 12:34:05 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/DVI_TX/data/rgb2dvi.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
Zcwvws4ZL0Si+OTncFjagR7U6q7eZ6sJsM+Z9bWy+HlEtOrQ6f4YPne88GWFn2YLS6yVlm2h3jLl
21a5Vwv92vW/h5H6hryoLT9pqhOwwPcf9yKmVfpWmH9vhYddI6I3a5CwORtBwDWx8fiUYu5UQZ8a
c0ogw11EkupFiphTzVPDwa9j1YCiMQG6lfmibo+U2b/O0jzxkS7ETozJZ7PZBHcysxvEGsUSjWHb
siVgXAuDVoxBjHtvAmW9iLe8ZkjNQ+QsWP9AQL4E9BEMI3Ho+ZqIsi8FBfI9p6CRimNxYlkq/jjF
QSG+hLQ2qR6TtZKdNjQsBKiZNHQk5bX6IM8sfQ==

`protect encoding=(enctype="base64", line_length=76, bytes=65584)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
8GBFZkfGFTdScuxdHolyrFHKb7VMaEqaQ6BhCWDTd5/2/mcyhdsjXdNc68J5MXyXcvb0SVYM4GJu
mkfbB46KpRorNRGvMra+Ln1rNqt+g84OsYoWGLFaQXvLL+IZlq4e6E/IhimqIhtqXJgdXN8jiG9+
/PpWVoFTCmFJ8jYV54FtKNgHAf4l38VqOQNgSsF34M8dl6cKIngRCUvktfPTfV0wF9vXvYSmY+sz
hTA+P+gGbbwYzH4K3D3L+RwDC9HpYaSoFOG6zN0oVFwJOJfxmw34ovnPqdPuZ2JLXhsEUP/ayEzu
+dwuwqUS/Bk2Th3J9sM5AgcP/LK01eWTkLyBxc8rTTxf1PLqX99VyL5pmbttR+GftmkTOtE5ADPr
6K120MWJuHr5Cl1+Gpw612QL5W+kH3YWXNT1+GezyawqUbPIPpV9lthbpp1lTfTJ4lSnZccmvlWb
CM9iy8CeiUZtDhZpuTEhrhyGHCISxGrAwGh7fcwObfAyJY6dy88L/UQg1SRwfzYnvOgz45/NznaF
3TxMD+QyQGRCZhqq1YtBkDg276vwtETmJXtSTP+XDCExIV7uGhndxat15mtbMY6AiBuq//NKMEZE
oJKIeebMgv4v+vTQVu8AsBwGNegR/3fL6FKXDOKsoqPuVUS2KhZ0aYjAzdwZne7TO7B7nfUg/oBH
d2/KdVOkG2ub6GuLnr6YUTV8sMjSjUwrUiTIReC0GZ4pdHB83yr/sSt55leGbQX86PZYwWoqOfB/
NxtUjh6p1/KE9xwm+yHVWH1khigSTEX3Tm38tpv6nXE69rn0OU4e8OA0LGvZhT0J5qgKLUMgtbpw
H+/ruTpqoofsg8IZEIVuGInkpO58/Fy1HjNTwcjv0HjEFwzM34/HwIr7OdJIxejdXI1c4IXG6x+R
DEoJZNEQlArc7/IYjony9P/oW/pvBbc+ZuMEjbkVgg7P47W4Q71HkATwy/g6ACn1GvoKc/qzQKvz
H3A/jES+xv+mbVF3vIG1SSw3q5hIBqiuVKdX2e5NippKhfBTbOd9OFGRBhjL1Z1DI3Lsafc5iaOX
8k46AnPKHi9mhYmg5hPoXgkiFxBNkG7vp1W+lo911E1bByd95HAu3tnaHfd+UE5B9ECMhaof6BbV
PVEYy9c2MY7Xu+UJ7xd+Mg+A0kNArE/wZjU5ATb3paOcVLDztQ5OpoMuiFWyjCSeBLikang/UmLv
43jILyUw10M+nR360m7t4FlWkqn5jN8AXza/RVdpAdEx+uwyXGue9DraGMQTGVMXjOrEcBhj7cqE
4cbCMChKcB7TsEoD/d12eU5CEFZtbgZgE5HAKKZSu/Dgbzr9kAls8BGNfJlWC9vLoZ+u7Q6MGCb/
6EdOf0ckFaoly/e68OaxvwOMcjbgS7QmDo5tCJc/ylvR7J2L5B663yGKLGXuC5oeIY1Wtqb/1Dij
mqjkNTXc3Ff9afEBnhln6ekAFv50vcZhjngNPmmM9QIlpgNHp0HCQkPm7OKlzpyAA1jbr7FTHk8y
9HBPmESjJPpkiMVvEnD6mOoP477k76qYGs48okWOcL2fvQ7r+JQ3qi1WVFdFxWYhut5lUukez5g5
R8j/LXM0mwRZ8wdiDCLLbZFWop3Q4G/e+W+GbygojoaYTxXRnrp67JToF15qUydmS9CFujqiRY/r
xjx/vBXMsWXUxWJaxYzNezre/gkbFp9ANPJqTIHQPBMvx8DeQt88PBVYkPXQknL7TwD9up4DJQNt
mjDQ81UeivLN0lrXDpeXClXP+i208D2750h3lvV7+9GTMnuz++MpCZr4mFn0mxokjS3kW+F8OUIJ
uRhlyk8j2XlBxV6JY20zWJ54UfBoHzvPcVfU1cDDZgcI3TvCZ1AjU0/Q8llAF2isjcH8Y3StZMde
sfFUZ9AAuUQppxH0zu3eut9oLRYizfcJ9pw/07Tl+eXOE4c2oDHG1SVyferNLNZjnUVsQZxoWhmg
D/UMPF6TKsBIHDhY9HKuurQigiuKz+9E7fNsNtu4k3iTGEuzBXZn97Go3LbcjZZ7vV0gppM0wRQg
PpNBbd6ReAbAyEI/CLUoa6qupB44wvyPcZ33849JGfcp6NJCTfJW0H7YelUAxhlDcHdEeGhEM0Sm
rqcG1L3tS9Vn/v5dRhxgHxlAn6ifvcKO8oIWIz2ypkR7/0nYtEmCfaAIQ3Wo/EnlbhoRg7uP9/HQ
a69j2gbE3DQQbgJhrZMR7xyKFvQvGRRDjmpC8MijzjEDqW6FJGlznVwRWtfsiZwmFuX+HLIZxe4G
nvxkzJxShYpeiAPqcZj/PVq3S0bCTzipmnoIFbHyxjPhF3mAaxpbBMFA+4XkPE1glhpGrqGlbE7e
zosHRWhzJqH/Tp6C+xbn0LDp4ndNM2Kg8vQ3zpJIA09CE8vLsQ2CFGB47YBJ/1PjgqPgQ9fSb7Ap
h2xf1G1b1VpBD9hVlo1t5TG/BIb5YizUGzOjwa2JBrQZaDPMfYgJn0sYV73tAbTIa8XKgJX7JHX8
V3fuDo/LGzJwWiFcL8C3uD9o0HRsVC1bgQaIpn9nhkGcaaphLRupbn1qUuRh5H+poQk9tezjXCDQ
dSC1E0bVXWE9GXjnrcc0ShRKAf8imDN7WBr9lx5V3nJhJcv6YHkOc54aDKxBXGuDE6YjARq8Lwdk
KF9K/zTY11T5icLtWAK+N0T+buNFhJeOkgt3BecZjUzCFZGtVM674H2l838IsOR8qCDtR8wgIaBY
UmNFiNW5U4vxzy/fgku84c14HwfsSn5IAfRInJE5/Cd5B/vMuAYakJytof23yoIcXED3iROb0M/m
dBPmRhayg1Yy/adO2cKJOf6qpZ7JtUJVfLuYI+HysUbdZffqpcCPQf2wTQyWLTHPooVqHd+FmoTH
P+IlV7cSB59Od6KcV8fSGB1nqQYarENsOyWgCshCQEOeKyi5+ugRRqabzP3xwMKirVLGWOmGgTQi
YsdKUPsl+RRsqZPu+E2RvjCag93lXDyZUaf1huIR9k5bjXDkxV8xrVhV1SbvuaHlcZbQx1YSpSVZ
CvVOiBykwu2mkRYLX9oAiNyS/Ko/HmJMEI8w4DgxxR+BqUwxpP8K/hSLqE1t2SNfQjpGBrQZzdBE
Razt6ItteoZR1AumvJuHS8zQc9ZmjYy+w4VHTJiP1ueDhf7XyeYLQrnp0QC6zJEM4jvXUmP2xtdb
9u+42SVnsBLwCqgWj0YEP/dByaX4fzgLdoseZUZK9AdV03qJeAeexIFCdGuv5T+ezFreyIeoQ6nf
pRAr/sP8hGLhQ+LwzuO3WUNv3M05Z/xvbMQ3ZbZ3ODE0f9KfsU5gr8R3VnFUuAQUJPFvGszkxFOb
4CViNO58zuJEtYC4UF2bnzZCeRGS/dFWbvJdP5DDAkVC4l9vISW599y5FrIHJkFMuf9j1qwhhLEx
dYV+z7ONaotevFh82NBQuAeLmBUpJ4yTP7OrvNxQ/P4h2KRmOFzSBYZQpTQ4g1QVLVH22VmiIkKh
J9dJlb5ubi9DNiNDYL3e3pDo5BusKzPkpWcSWb31reibBFTalXJpzxBoCteGcqsoMMhTi5YO8mcE
KSvA5asdOQeUKFQOhzOSKRa6cbvtyVNIt4f9cz1FahqLTKWy+kgRf6zjxFVJkCYwypQoYFCrCjHu
Tw4F/DUOLmdD4eCUGjO3MKSF6JwW8StNaUZDEWT5A0DZqI+WVPfzu4GB9XzoALGnaHWYaiDOjdFX
+jNLU53w9BzZIoe98lQQLCGhPZr17XyOhAAjbBtYJ1JkKdLQb6Qp5kcPP5CMdicaqMwoHJn07Ao3
xI7rB5jAqEfoZ2CWrYfS/0BOLY/fZGpY/laT3OW5HzplmLBBpw6WAmZUKKAcIbOkSFS2v7pm/Mew
XDXWQ0AmMRMEtY4RuT8QJ172uZBxxZG10Hy+pfVGOTMcaHwq8aEtm1E62/j7yBdJiCL2xbiCOEK7
CWkvdM2otTPZHrBiEBXh196/fdJzqpKeP7Z+7WFP/ETEzHiwNInbyNUJLQ39UArEVQc7sRFB5H0Z
PFfmx+nX0N4VXPIA0uJ61Q8g3OMBFqTz2khQbpuR2ErQRHfLWPCDSi793Y0rRawO/V4WjJWMJLwe
lP/09WhUcsmuICAoUOGMc0FEfgOh9y5x3S/7VDQJCqLlyfJ8pB1d9KR62szYjxDGBm/vJFID1Iji
7jr5OUD71vymFnKho9sEwGUkHI8yufsIZfU/xU58choZo1n3QNBekGJxVKdHr8gho4oYnVRVEX1O
bjEbUAlfmU4U2+XbxpvMGlFuMLVtXRjR+LNUR34Xm5F5xLPENHU36ENftapBe+0FuPt7CxN4b9PJ
Lz1S5fYFUCvgQkNpbpK/N00tN2lccrHK2g65eJgqnrmRWxWe/kZTPXsHv5+Daq3jGVLYfQxjNh7N
IJC4ILkp27E1QfCpoxq+GuKaNiK80tu3nIOCsDQgQ8tLMIRkAgnrtQY7gL74lT4vTbcAGwP1w5e+
UhiBGo6JNZPrc0IxjRq5pQHgBAp46xjqPcscSKXgJqGEB413LR9NMNnjhkwfu+hz+DLPN9Ip8ctO
uFWYGvvGg42Rt1h+lPpOSOqjIHr3mFl/4THyavjZG025PzHxD5wEkUyhi/v+wIx+ayCN+xyDcP6R
Wfa7T74vv+b8tdfgsR70bzrHp43BV7doEIne0ZdF40HjbEYq8jK6JPpN9/jxaTya51t/a5txyRVM
TCXdZLmW+9rxQDqPvnsR2Ll70BkABFyqmyAKqNN07RhG3q0nnXt8ExCztvku9qbi9RaqB1rZ++QF
V7zWHM2YhLzSNwz1K0Uu4v5VgOP8yoRpXMTEIwEBW5suRQUuu5WkVfkOiu4ws7/l3n/YwRtNP/gA
DKNUvBda/lbM4nT610uYIVLtbs2hKiCVzsxTvKk+/vFQf4BDIZBpR4Ix+Sgs9uBYbnanKIV4cQQ8
7ZXEwd04C1GKDKt6ucPsbp+r1QoElG4bcaovoHRXY2KG3lDnE+2DOB9tUszK44mzpuP8v48z1dWR
IP0V1rbbN5csTsthNUb4bskJuOVopCqnfD0es6ux1sr01JEPJ7Fz+viNus4sqP5IvuG4sS6LUScZ
cVVN7cPAGE5Wt9nhlyUwDKbtROtg5s16stCFhDHoU/1rnAoc4auiGHKeZ1i33Kj4Rhd0H5vahVpU
/c9jUGcAos6GIE7FAZ/lymkoPqIv9aahj/DI3uY6HciZUfdoaX71CF45p/uoPQGxPp1T+O45U/Mc
iuISwu4IeoB9ve7csAN0/67ZLZDJNxu3IvOJm34680h0nuPyfytW+e9b8rQi5AMyfHab8e+JQsXS
jHrb3leJIC8RsqnafC+kqhMe26OSWvxENYm7Z8kIYcTR39aGgJVwfYRQW5xIaUa4GYLTpDq1rSsb
K0hGRxPNjdnsle4ZF8W2fsPVEAxxt4tbZOGVcQt/c7t8YExEiZXJQtxRFkbGEvgC4tVE7N9PGq2R
x4WKTmmiT5GF/5/A4oC1DSb7F8GkHX2Wm11gK7n4R5nAXn8S+oh2TMKb4SLwtWA4XL648c2feTdo
TfYcCViylJZtBEta8M0KNW9V7qjSdYM+1aAGMpa4kcOzR0xAv6Yj6dinBqxdF5N2St9Z4GDHPiaf
HsMhkirEztoCNDTeKrdNX/UUdBrYT5qnwpbi409dXlRidy7mhD3zMA/kWQLDF0y7sOsTSGw9cDPy
umkSwIAbrC3ODD2DkxWnyCkmnPMRho2whpVpmJZJK+anE94svuudmSVnEzrMu+qppDaO0MqmLmIM
Yio7WjOO7P0k2i8z3hcNr3nIBTMoBx/vuTeEh6I61QrxKiFe+OsTXTNPZNGkE3fNkt5PMDPxMc3b
pN6QxMHcPBWjmiJyP6P6LiSVQcAOpkkjxeFkxFbd06eaJaGiO1fcFWThVhrw3IwndI0mIa7ltJWM
RamO7uiXvnHSYa7yRe57eLIDEc6bzi0adxPBrgA46kYT2qBw4Onwo/8ht1p9gtu4XEaxGuaD+ZFC
yFLY4FFINUkgJ3GtmRLhCxF533KZShFBB/V99fmPsfGs5Irk8M8V2oXZziRFyxAsIeHn7QSMFidi
U0JL19FWZ+HhiMRZG3hKxCPIVm004Ur6ct28KD71tX3h+Yjg5aokqoXIduf3hbvkLbqLROPKLgyT
+5vUt6yCvA1OOZy3YxinJ/zih6J2aflvPOg6H5GlALyTyJVTAzkJE8K5zVRHUv/kuUxwKzEnSBsR
e+wLLqv6kwduhaML71GVm3Vf/boPdnFYRrAPQRLxXbo8F5rkHpCZXcGIIGtQeYMQ0MeFIzuEUpwj
jAkbYSi9Ssd8ikMRaHylGmQ2MO3/HlFhq5coKyWKrfhntPSfqLC35T+4TUvSBORP3ZE/iEnEbTF1
dnIIVJQ6Z22EhhKg+Jdu6OXDUmMw1Vw/afVdMT+SZZ5K4sxWT/sEZFT8LLdx9fnedYsnGuPO6Hmk
/Cis3roiACVfEVCLWCnFHTdTdmgoP+rADrRcbRCgC2VHFYsYyRlrb/NwPLDq/EQu0X1nF3oauvMi
K+NV8e76XtWx45QjiEv303oEEEfcnJi/vj5Bv1PzXj3SH5tpP4Dlp2luCfqOmALVnpOChrvg1nbr
u8JtxEp5wsF5SeIKtaouHZn0xEcPjO1UxOtmEq9C0Pk1O8zUjEv1NBa6+8MCoL8rwUx+yBVj+rch
mEGhpcUKMSpXkXTMFF+ypuHTIGSLHVqQQ2VI9LLxrCB+Fgz7//7KsQ3XJ8MWjT6PIGc/1P6rDRYm
6OjrMnWVPqw3vGHmC5VNB4Yc2garv9a94aAGcY5aSX4Xygm9R8kAgpnRntgLxcXSf8k0hdUqIiTO
vV/sTEoybmYHmPN1OMwFWN6E5guXDmTCm9byEbKXG/XdwfUhh3d0LMMuNjvvYAWG3JHCI6ISaTTY
Ix0nExDx4Jyho0zWtN12LczZTyo9HuvrEzkQAkxa/hXJvojLpzqONPXdbsdLS88jl7t9/9EpbrVN
XguWUdNf9voalCe8nknUrVJNEMD+aV41p4ZV62iSKxjQO062YDdf71c5Z+O6PlokFEhnOXwoTAdX
te2L2m3zzkvyz0IvnUjb9iZxpmlsTjf9ssySvFoCyycA1eMAWE0+9e519XC4jI7YV4DtwZmYVpLJ
pL1XaJs7QIKUHhjc2uFXGcZikIPcWWAIG35Pdt8R76Yn1MMWRwWFVoYuT2f74RK+5tJHrNjqWNbA
/hiGPtMwRSaBFOASRIHFNAlUQKLpvw9zOHYW5MlI5UMuA5YZqI+653HN039x8rjoQiy7RM04YpNL
Cnum2EAhKmGUtVwSzNLr93FJo60iQ7gNwr9PBq8vhA+Ic0u76DNukvS4xfcXbmzL3EBguV1iLDKA
1Vimu7buDCFWgMseAJ69q7ghq4InnAB/Ow8yn3cEydQiWNNTvAUDmYyXgaHW9Ba1jvpw5tm+1puS
IwOlyUwgIYPbxnc3TrsLkJmKRMOIMbC0RTp0Tfn+T8dUveVJg6RC93LQPZ0h6fg3TFmoSzL01TK9
Mi6BlAk9/L4y9ZVuzuH7QCk7OpBIvSNRIhc9maPi5CkI1bWjFICTr3H1F5p9UuYVEAmPbTjECsIq
hVFV0KTltoZKrdHqxlA/rOmlp6mBG1EfCxt+uOtlYsk2TABLSvDZ5HUM+ilMKgnLyd/XUWtTGqoB
IA38E2G0aSJ6qb5USsBpI0U/X7TRr7xZJ0AQkZZgBTlAln/yb4TH4Cf1nAKr2guKhIOsmPBkE1d1
Y1I5RrSXsz4qp96d6oHg+c+ipAV+GvogxstrTwtKJTG/C4KFSYVtroLc+vpzaqlBZFP4qB1dmOI3
nR6OhI1WDTgSD+mf7RW3HJphtFayODuI6D6Sp3r+33DfRzX3fMy/1a1Og5gkNVoo8flY5WXZo+Xj
pOhr26pq1Y8wk0dNkQ4MlXxfoAg+VZIBf31SiEulpoU2FAQA2D9mjAwlL8t2QEQ2kw9VTviGx/Xk
36/DKF2iS+sE7O87ZI1HdCvaoXk+1DDfvamb7/UYXM6zyMKvKlD8NEj3Y41HKMGj4DtLrLOD3FPS
BBGY7dVPOAfDwpf+fVno7ViHbXGDkwTYAhmhTHVyMcwkBReeV+L6RKM9QP/kV99Iu7lixDHUwMod
dmJYMqHqxKv9NriSR3ChLiC9oW9ZOd4tTww5RfJOMxTDlLPrYpKLbgkNdjW2JPmeAzsHaekDd8rb
mYQF8JLZCEcD1WDNkyDMXjXayr+s8fnpkSIWyH+8t0aFP7T40UivRSTmB+pWxdzdKX4R7IHtBDCC
drBTN8lbrVS2vjbuY5KlQv4Cs1aZsRdm98YqrQZd05iu6eNTMgL2Fbyuv/adorlqmTKoL21d0qIl
xN6ddrUCs0jPuQnmSbYCNqLboRhAuV+gZ77gnUSJz2c32h+WeIISYJ5v04woA0Y7AtrN1chIHpYE
2Y0IM6TngUoOpLBykV5gdI35EUwnPtTosxIyPwlhBiOHrUzl050+RRtqp54eOKusC4FZcS1C5/rP
URwjkx1gvU7EbypuDhEWVJRWa/k66Px7hM+jU+gbZYnWC48xt0H6P9kE5e61JVRd4vr+tyRVboCa
UBwJwPhoND6Vvb2E/LTycefUU4yFP1jeqBQW5rJAdA6l79GYP+Ld9+rYfBxRFE9qVGpQA2GVis26
Sm23NkZfj58Mrxetbcpwbuh8WxSDygqi4+4fDcYkDe/mYEr6azlWG+ouKuNWPIHmJCmYQ/dUHMn3
obpLQnRdr3HMpruYpQbTrEFuHc/ezx6wrDrjaRNQvPbvXUAqd/Em+ab1PfZRE6K1e11oZyjAGSSu
qDgP1CiWklcu/hKRHkMVdkAu5kZgLqkM8c4LSmfvkdRGeK1Rfz8r8Hd48R2OForWwK7tzqLivbN1
w7AY+GouVCOp1M6AnMXqLaGLza9sbRx1Br/aK/UVUHhPZyftp0MEBwFlrvvZJwj1gnzsxYYK1HgI
6itFWbQ5Xv7+a3VME/3jvpLkP2DOwT9INyq0ezKDeaInos1fJTUkHX77cH66ygBA2FEpZOLutfji
Zsu69+bw8+N/oZ8OYGOOsxv+lOrBraDoEeuCFBd5HQoKmvAc1e4P5NmoN0sBHRDu2K4wgwqQdJaw
alujaKNbyyrbjX0KhxeRNUzQNY9e3s0VVmVNPzDP9oZjEd9JgnnwCszZ938gGb5kyxeGLtCbdHfo
+kbunBD6rEtHQAMusC8fba56vC/kdrvDlV4/Gkb/1pdO0Y+ELcOLKqYHSSSg8CS8bPoIv4N3cnlj
oXGrwgg9gzSr7/kqbP8WBethlPDDLrFPLSCwA8fTkJTOYat+ZxGZBrQqxqT3CBGCERCPpCHouYra
d26DLL1A4bc/LQee+xdCvGm3Kfe2saXSnLyGpO+c24iv92LqAGH1I/J5lO8eHLtSnp5j+QkatWgy
R4iAJ4tnb3ii/D8ct79AbY3LQFuskBqZtNmFpVAgQTeEs0A5g4wQU+KJk6OoNQfTTOXIxezO1wmc
ADoKedBb9YPACIg51pD2x9wshwSlVt/lz1sSXz8ejk4Dn1DKixNnt4CPVTtlgX0B88R4ms8yQH7g
ALrW7rIObZqCCO7fZVLfae4520h43aD0AsPba0lUCAXvF2AbRiHwxKMq2jSRI3QKaizsOHj4LuYL
Hb8+I9FFLR9gzEM3OEVhKMKXPs9mDuoyIT81eBJaM/Fgw8BwJtBFEvnJ9LmSmyJK+8pMuHdZeheB
R74WARRY//CgUrjxE3bRRijBPdEDlinw4Rm4mfRaJ6llhAZiK1oOTy0r74JgUR7llGQu0dYU33zt
mzTwQmdHtP4L7mCni42ekc5RuQUiD76ghsFtxmCz8O7pt/FSoGTw2mKTlJPmOX4umiqfBcHP+fxF
LG0ehW8EoxT6RNiPYUfCbDb2c/+6FkmJgTMl7usdPfx3geaVoLJNbXc3c+myd0ne7nrDP1wEtnTP
GNlzRVuWtzL5uNvRBUEXfmq9OSit0gzvl26t9UawrzBsyBhqZapfP3/uucnPzaJDHZYujnDh/lvL
UGO6OTLd11/Q1WVvGz2CdkMEKm6/VP1D2vzYs+RzLzpBS4b5ep1Sh+cB0pgls1MWlPflhY1g4XOt
m+wv5pxHLiTEJudwCOCybpNDkAYU9C2I6oOSjZMrRGk0HqZBmstbLTAsxR7c+u8rFsxwnnEGaFBw
mPwxh7uGo2YSIonyg9f2OOv73b+JFMfTPWIOjNK3IwSVZ+2LjQFGQCbLlOJSGU9rrxH2gCCqy+1p
W29rImgid3sgXPZEr5dKckHA0yMBUU2HszoGj/hCQvTL1drEvfgCCT+yUqDbba9WpwFRU7QBzJTd
OvGRKPJWTbrNJNpLjmrLzXnnLnjFVQSTtqJ8UEFYSuDtyLDRHt4jnItS4DYMA3tQBrZIrdxLrhWl
r0WMyqtEthWJqPyDPOaLmvh5jUWAhrIeupq01UvGQXaim/Nvr7NJyJgWk3PcSxL31tsX3KPHBWwg
FuiWq4aRVES9bJYafptmKGSDyMAqbrgo2U+akd96loZqnKMA9MPv81l/EefI8g8eBst8Cbp86UE3
GxeSJQoOBa40bmj4mpx2klmf4GiqOhNAv9tPGBSSuLQYLurqUZBpKUAreYJU183Js7CNHb8pLNMC
Fr9HVV1LBtb8BWMvt1pTi7HQtmtb+L7jsT7uh9XW/Ds2NxEFX5ZGxGQDYiABg07slBMy4M9iawFg
DZKzWZmqhczlsutYVNI69hMFi9/r0iGxQLyd9w14+0lzeYN+Dt6Po9rdxXcBZnIrTobmVatF5cYg
wV9/7sL6TpnHII8Va6DZpZDaqZhx2jS52GlqSBgDJOeS4akw0r7uTeUjamaxsWdJJiQFGQG3+jLR
u3DwIbf2Aa9jvWDkIuaUKpFIi05Q1E7lGkrpjYm89/IQ1MtWZabrf2/nqOv7LcY/yRQEFDKHGiQf
rNUKR6ZDQTxHMkP3qOFnZS+01WvieLVq/bxkJa+3K81rVwNtA5iiZxs7re8PAGmpytl6HUFOv2uT
M5mA/r4IcFccsDDshCgz8V7f165iKfx8XrkLKt9LEbhSSZ0+kNYT9kJa3DuTXOvz1jkSYglLcHjP
VCBwSe6yRcwSEIxF2hhBGh2iqXvcFelx8y0HrQLiipsSEWwJt0SM+/fYiHnyyDj1sWjIvjsD2Kds
YyYN9kxZpoMaLzh+TNskF4vS0PirFaqcQks4mdmkerizNnGRP9Bk3t+UhCKzDKsS4cUMPauPJ+FT
s1rAJZlf1MVXUND4UJnHpXETjx679523LDrxbH57Sl4pUhCYHQtIeIBkMaeXaGo1ZAJUoknSsSuD
fbnXiMP/Y1/hBTN5oP+VaReRIM5u/XxwtdvP/SMb287lBJFneIiW/L5JsPEP2JerkDh/hf0v2hvw
2lOh9/kejmuYESsa8nRb94mnmPRlFlvOdsXuvg9FRAZJtU/ZsvTgKr/CRHVfP/OMgmO/Xp0kZqII
X7kd++4ECigVcwqWlQNm2g/qioSLS7YjXawO5yA/7Fhk5HmR3INm5pZlh1zSC/6ClfzM+f4Q5GKz
nalxmvUW/Tr0m2Zn4b4JUHuFemqqpchbdUzkltrMo4JRj1+ch8BwU0t+gMeLGeoC/4ctTRdSJBTN
lY9pT54HqjJPf3E0L0Kcv0W8k6kQDqOuYQ2mQQdVhs1xhlK7bgD33IBM3Jh/WpPlCNJSO0yKZEHa
zUrIoweMOUUgtM53kqIRNcjFCEYlsE+4gpKOBPycuUKxbNBnrbIxE4+MOnztjGHj4a/wRoZC8TfN
+SadYclhRUPf6qA3EA+JfFCPFor7rj3ZmbTn528ugx9R3pb5v4fLMBulre+TcLrtex0QTKZbuBZF
N2rd9TeA5S88P8SiKoIPwmim9za90uEVjNQXh759w6jfcFuV82i3lATa0CmyEC0LZ8LHK2FoXi4H
9399M4E30z3lkO1mh+Voob8gYD/bY7XQq/6xb1wRbL+A1MId39ne2Q5GstSVbuRVtOWtpAXwJVbK
u6qvQHJPYQJiuZstf2uJ2RQFgGoxECOeAqQU2nllMzhKVlUMgBGR9Jc12efDs2vGjPB4ziwCGWUz
TuweZnmkecnEw/y3LgQY41RC9dOXc9hyVULtf3/Ge/eytBkPb4AO1TmA8w8pw0gILT9HkWm7v5aH
CKhV6LAzOlezkC9FOB7G1lvnxmT2PxNgSO80jmkdJtBgodpvS/mtk54bbww0Fd6iScTzbm4dg56e
H138fBlSYu335VTMU318OtTk/j8h3H6NAMFivicSyX9hT76n4tBVnea/YgmXTSkoc4j5iqW+KyVb
wKqGDTzoq7Jv9+qKFHz+Y+e2iHxiIAxUZggpRPzd5u9wZ9ppP5EHDrmGQrRheNoRIJG76gW4sUSD
rhYfvmrn2KrpUI6EQVVtMYFEflHBTk8kYW4vyx635zDqf3dca7taEkOwKfhknqDxXq6wI6eYzW6b
pLCSd7f2MpoUQ/pPmtwJxedUOVJfIbn27HG8bRDZAgwhSEd+rl2ITON4ETbiWYT44Mz102QQ4vIH
AOo6bvoZ/oL6FK6la/iAXujzyGwKZZfmgeglKmvoASN0arTW7qNhZ1xnF8MMsPa8xZtKZYn4bhT4
2H3HSduYkcnebuILYCNveGf2ICPJ1lV+Iy3n4bX30fAHwelocUFLjVU9AT7sSSMXE9L/0KbdB+Oc
OU+yF6RWExIuQ2Y12qW6p5XRPXJMmMcgjae1AIcmomBfiGjLFjq+TyY5raD1fV2IdoLg4pYIml0n
lr5kHZPDpJbW/UCJb2ofdcByGFjm9+BYM2gVHMOX0m4voJylYH5jHT6eGYjy9QjkADB0U7KnRvwP
AQrblKQ6aaVPvcfiuqPlpe68oW5ujZ9RNHwJ0FgJzQ2ViC6tR/Fmy/8j+/elxXwxngBlq54b7mu2
YU3VLoccU1MQu6Z/rGL/NZDyDCEavgEFSyrqw2ZegAH8ENXAIRTM6bisrpANSmDIP2uuLlXTqBc8
+55D9nRTB26pLxxboW0e6MFrjt7yTfHBisulvK6IiEybBjdYUtf2XRGct72ifevQbAPek69GBmKj
N4mRFecdz/jRjn1fuyh1aapsgu2ntfAgfzXQNs0YlaCFEn28x4t0ntw7c37EVaXOUf1GlXilGb6m
+giaonBoZUG4zRQk0KjwHaz32E/aLbB3e87r2O+LqomuW788TIdSfgQWdj8oZgJvprWxxWcbMY+w
Q+A1phz92tpumzSAsNROSBCstuOIt/vLnNkZhEP21X0Sk5QgcnHbF+jc2nUybjLSIKzb8AhE5Tvv
AlLIof9SSat1mWHo8uiNBID5Yh7fKQY9LhrcK6S56UcLKOnhoFYwwXB1T48WxTilWHG6CI+XmwFZ
xfgiQ2XP7rqBYkP/A8w54H2pYLrRFTR6Kgf9tkb6ASJe3RYyVdjK7cIEtomduEwAuZUmvAsDhdIC
bWrkm7mxGQkZLy6HUhCpNrVx4y+QnPSwCoB3ElDvI597nF+/igPtkuMkN7574I6iDZ6RooZZcvq4
V1VKgEWrh8Kf7XBWKrjd8CBM/n8TTSRA3BfmwX3ayGc6eKQTxT2BF4url6LGS+jqinAV9R51F47J
PyVqwDsT52qTYRdsQF3MMp3/zfSeijR6hxWb1nptjBChKy8o+UfFDFMqaoM+MPyq/q8jfNYXx985
ExddJbY8uWnsxX5eYsP+ZKqcaSsgv5izDAgHG6/t/a6puezgNJre7KWq2gpHvojHcxVzspEpiJaP
KGAxZ27WoGWBvF8Z9tTED84xvapeSZAhxOAucUoSHityHZQbPFD3o6RxM9We86FL0p8FHtqoQIY7
BN73u5YsCpMQ47i+xgQ+iMs60m/4D0gdufYoR4TuoFRPdpnAtAs5dTv9kQbA+c3MVYaO0GYx4/lF
srRaEWhrwp0m+VGcj0mFV7PBi6QFW/EQ+JzMyKpbWq76C6SkLGA4bhuBL8SuaMR1itbsLvX4OsxE
wzxHozEjSjd7Dmkmnccb/ieZfer8fPoAwU04wERcvU53QVFvXS0ui8rryDCZzRIJLp+Xm7qd9DHN
Xc/zvvo8J1KWxbDTFSYuNdd8Fat6WIwJZrfkkQCWa7CmUMky7zKksKC1en+d2I+2SMJUmcyBwHw3
qhvvEDQU54bv39a3kMgxJDN6ANl66qMMhZhTHpN1dH6HNiiCBTaWaNnMN0+vp6ZMTipV/iIjqLTj
1BtPgQ6QS8PpsvTMq/Q/r1eWwPOYxkyPuJhlYKxS9GHPd5M6w98al6vgQLqw2sDP5Pc02tmPwuJB
pYv6WM3CSfj5gtw5/n8aLRvAiepLBaqXC56sxAPQCGv+eld32Cet3ORrIHkNj0RkzFILc4Ev/3gm
Hs6L6GUDOg60/K3LWIZakLU8XA3MwBLmpbqMVmf3cP3qBTxAT4fR5XozynkVJtfjNH0bpmObei66
5zLeDOvRJk6HaX+exq8ttRkFTnxE/wtwv7l/7i5IsWq7HjphOVAUpmwOsNUrkD3ISx+rw1ip1XRN
gcrcHhmodXT93kBBkOdyUslgh8l4LyXTkPjIw3pq6dCtUrMrgUUfVAhj+n/EJ6lsCdcgN45wg5cZ
ea0+VLi5UqNKsgXObPWa7BGZvpjY14jtDW/JOO0PSFarRmFAD4hI7HkRn5OnGt1DZvImtfo2Qoqv
0pMLskG70SSnPZP1fR526fPhfrmgHs2KhkbV/RXi97lkZ9/v98SbTsVjSzkWS4d8Agh43Jk988fa
d/2WXYgioyA5k4X+aTiMzVsweREYkxfMAFg4XW0PsS5Oc7IlJ4z4thJ4hf6xVP3l5tDbBYXB5w4X
H73Iq02rKf9yJfpzWBN/aagWJVNL/EnSb/vPNJqFjqm/BIN3nJTa0MopnKFRYI69PobEtinLFR0i
elqME39CZMQc7Cq7CRnhL34KaqhRK5qEmxjTQEXcsn7aHcK5QHpCucbA6pwK4J0TXclz21th9N2I
aBH/NyifAHXsDLPevjpeHhyM8T/k+XQRzEelbjR8YyG6gCUmdhvlYMWT+B9tC0TmK11us7HIMJ9q
yYgym0k3JyqqTBwRjqzR41qeYSVHeZ3RcrIq0QAb3FDAZYbGDYu3/0QHOySwYTGnOChYST9eshqP
WlKoAFXKL+hW7kWBOST474F7H02bliz/GW/IbmT2UqUDpmFTZk45iGKKI9+VJaKvNFJXEGZe/A/I
FeWQHusYcn6SnT/aBuRi+7KJ+SnpuqIdI2gkaFSWiqxi0g/o5mis3owkG/eYY3AEP8WeqAT9lkoe
aSlKpfkzhWBv/PKrnzBrD+4LAljuvclwFyAtwyV+IXRldTkroocPS4LOngNhhwT85U7L+FD5VYPf
UMA1aopViVlZFY32WSvJEkuCkngYKHXWyxEasRDorL2cHai6gPwadQaz4srimf/Raw1TjaGTVuiK
UR+cEavHsDn/S8pPGfCPC2GCGVWmPwICU9tp2jDuF6Yz3VJ2mTx1nL24SeFdfzIhjdAvfvqd5hQH
I2OUHXC66UMti5Jg+iIKyrMUkxNTdjvarJo8zMGWESw2Hmwrv8HYIntJyXstKMi8l4SQ/KMsQzwz
R+0cAuFmFGUv683CtwREhI6dMPL/alGkMgylhbO9lsL9eWsVg+m6dBMyJF8FR+pQautOlde1TBPZ
X01UblPuw1uJJ1WvZi3gaZK+nZT7mekMwpsNIlkxK37b1ShkRCag2bdEkqqqFHOkb3o6sKMdMvms
I01b91IqNWpqlTLQtxp0pBl8ViIiq6xKgmLi2ZdXmg5HW3BSblUt9M0Z+htoWxPAhD98yR+Y11Mk
idVdH6jlu3np4tiIQcTsIGB8R6fN1TEhy6Bxt6WLA5Ce4yQIyIETC2IdK/C00Wve0RTrwHMekG9L
r+QqxNjdSmO3bq2XHNC/YUF6rswh4Ssd2vsrYZ4LsM9OnmA5IM5ILwG7VzwJgpyN/AXt5NUhJGFk
O0iVIxUjBzXqQ2M9Kos22tiXKvK9a3MejxhpDLwLvKbIa1E0tWGnBOqPCQQzIbiiBk4Kpg7iAtG9
lEq1654Z+S750unep8AxbnnVUuGt5IVioZDTQ3r4px7keyaOzQkL/0DTarBO6r3F+1QmKr4OZYg4
SDJpUGL0WK2AwtDTo70ZYAaQK8/uqqQBwoAxD+YD7aI8IAkrs3pfqwbGhiIAf09/th3zq0kjraEe
ENQyArKdO3a4Qbc22FJqJsvo2aSsKZwBBmcg+f3c81d6M4OPx8cHngtQhEBnpLnI/UPv6GfJ+cwV
k3NBSdJ3E1oZR2ZhQjzq9fCWeHmCDk2tGQ1bGLNoFiBU+ijtFbc2JF8jWjWUVQsTkFHICDlWkjSP
M6Mutt76nPcl+a8bYjrXyECucEOT7e0j/zGiGoKUYZz6XLwWL1gSk8fBChmW8AfoIaLoXO8I8jiF
LwBat4yrut3lF7+qXwL+KBljfupxxXdNB7kDDtMhv4smGVZ+9owddiAP4vR+5diYwesNrZsPbKeO
2crg1V9n0rR0EdtZejw5cR2SCcrp2MwELg2tdAt4T4fLECeNYEsvIqMd1n8hyxbWmGH1O2JZYw/9
vNhOvXhavvrwGyUa5cm7gnmVnD83pKr1BBkFR5Et6ahyk7WJYNTztfug7r8D4iBPVuE376a4UGPy
X1p1K4YV7Bvx2TfrPV5E9uuXMWED0T4SypS0Kxuy/r5ZNgoCFv/t2G7of4Qu6fJb1W8c1I8TBogE
h/E7V1cBIPhQWOrfBtw1Ze+7hfFK9fvOrcwu395diGaJeCsOHji4WYomodqEguEq0rMp5VDWpq6Q
/BpqWRYfvvPabfGGDHW6oFrZBqSBmFgopHgSUIKuSOXamVr+AbpX/lPEtOnktZ88/QUTPRWojiVW
p8MzJN5ZqEqv8crYfIlE0E1/vJSGeOF0mns+E9/XtpMJeOzCHURDL25AySf6P32EL63d7jSwjQDZ
DPoTSLnK+lS4BEGUK+l8bvAR3tvQH12skJhLmkqoL3ogLg1n7O+0h1eD17mHbXUMk8ervVqyrmKU
GypUo8dRpWbfChgjCju6tjERSl3sAQ0GBJiZILR6ZldXqVFJ8rFeOIS2CyINwHLjkkPWI8tAgTgz
obOD8UpbyvzmKIfWSsKfwG/kSAz6kBAGaJWf2kd9TC6WAQOtAyOLaxFp7ICOdAESSz3b2i4Iiaoi
booF3hzjGhDbYOylHAwXRkpG3jyla4g46G+Ez/vODbPZm/anA6lxWMR4ZXG5B6F7XIeO4DDCGHBN
W1efjqvpBSGZ5Eg9bPwZR8E1RIY5e0quBEpbbC1f9eAg2+aVN8NltDXG04fCBztU9dHwEIQM5i1f
481Ar5Mk8p5aS6o3iU7XsZaM/t/84/0znBCoJ2GFiKAW4WdSAncoioPtzFZmo0tIEGHykUcGgMBj
j51vW5VghG7AXfHCm47x6Gp1oEgMXxqExxGWs2jmhrRom+bpDH7y2AzC4qMhlhOrlfLPszJUxM7s
d8SnbeB3gEHkveWa99ca4i4VN1Mj32ZApi7lGMyW49LdbpMnloH7Em31i/Fj0+Z5Stjd7aiJio+g
L6xx04WL3fFbWCHlVVppfaGnQpTuFPWoAamULTKQxSl/fzZXmCXI4aoogmeJDBh+0kYMSlgDDNvf
1XAwo0iC1zqoWhhBXmUQCjAnZi8MuOT0mew+QBwugRPr9SoRS5HtVlTwCZExjHX5fMXHRNZeWOyu
ghOCa2wZ4LY/4ATE/x5BeqQjCcSM3LLOYOYG9F2OneqWMMqmlxots4JLyyXmaF3SdPLDh1ZsTVH+
2E7kURPxxX358bX1ZiIp4BCsSA+/mETYLtMqQO1D2vHc2wLIUd8IeS2Nr7Cr1BmtMpG2KFTirvp8
QYD3lJKGc8SRL3K0n1x521a+FOrJv5PDzDcWdKLk2pbQ1Vc4pmiLexeRDX3tqocQDiVZpFtPuPZK
BsS0zffwD4lwzewvFP6Im8r8HW7YW7aIwJpJkEscBOg+0HFnwXB0ReyV8TSAbDJuDbOr+Z+5Wj3u
DmJdb4kaegkP5KS4ozSkOAnc9V1losopfAIVc2e9/fLaJLt2KgJm+dD5dlXYJN0d9G9rKFiycBMA
6bYL1/Npda0Ec0orFfSclwMP1781TPJk8PNR8MaQcByDTqsemkXKZeBLBZNPH3d2e1q+mWmelWfI
RiVcaHi4BYdsmaqcdkY+tNspL+hscEfJn7vxgkHJpd39IRWyypnK96dcCNGhvmGuLTZL/63+vSb6
t54ksmpqKLgLnLB2ggaFwJk2w7toesiap+13tEiURWj3N0sOFcmF+/GHfmKwS1N1ulYjTUlLzhq7
ozS8dOWT2PahFo1JcqgvfiAHMv+5kEoTjX52+gE65GNFVpd8bfBX8SlRYmeXkthxY2yD/q2AveNe
0LMzIorCdQ7WRW1ojWo5V+ppSl11ml0lpMfaqEyrn8r8eNwUguFaKChblQN+rhVPwzzSsh12jHFz
xw2Je8lIMCy2duwRILZeDSI8Rk3QVQmbXpde49W9Rzv9o6wkNMXH74k5ViqlPgllMze8gB4sejZq
cSVTC4D+hqFGEC+sJp7D9maeqQcJmoQ7mE2YbsCnia3atmPo3xRBZa/aH2dZQWAKwKsZ3YMxKQ3D
anIMgNPwtNws6G6PvEsmjEjkglhe0E4ySdjdf3yMawxUUNUYuh0I/hMMWX4YT5Cr76EOHL6nwujV
rGWnof8W6xE9c9K8l+dwnE/Pu7wrV1E15OYbx+aw+Q1kr091kGEs/k1+8SMAtUcven7vnFoWr3Kw
SLxGv0kkFYGVUbLCAWzt0wGnpQ0KTgjlkBnQwqTF0CVWhGayFfaaSllPOC0mrq9SiRUzWSvrWYjU
QJW3guPvf+ZLeH0XO4z3GuVMt2ZKdKF02t6Hex/fgAGcFSMSLX76NAsocMHKcU+HMX/rrXE3cMXz
qEzTocr351pl+LYehFCuQ0j0kcbP19fiJURzuE2g0wobcwTB69ZAk6t0yCw58rwuurk+JFIDFzRb
G0kfmkwvaX9e7QCA7apNfaHlihZwLKadisypu8iApKO2drfLB4YhMXOx352GW2f4kzmTI9H0tIjY
l8nw7A/ZN72PPmHUqFTGlTZKIWK+FeuV/pl2o5gxzs8f5qZaVKdxdknJEhRtT7LNKtzl31b/DcfJ
0p0wK24ZuQx+4wSelchqukAVSTtWF6etoOBMgSEMeGh6dJYJgGBVpxNIg4UmdyLHKZndryx9D/kz
YYyvv2/NaYdkVd17cyWgtr3FdR/XdTHUD5d7/J41QQAkB2L143RZTbChFcnE9T6g6wWtFW1kYlYz
3K4f/tIezWoHpanQ0U/+mb8skXVIpE9P1SAt41a7uxD4LTg0nV6qbGgpppPkXNdYzTiXYCZodnf9
ghiilvQvFOZhYo7qTj0mfphqvoxGN3NQpblZuHBsFyLEx1bDh1G+a4hZU9pEPs0uq6JSNG/Jt95A
P8shmSb15uvPLle1c+moj6HqJNGRK+zkdOtUfp7+UZNqrfpnqMfHqL7UmhtVlWLJImENIMmgMog5
Au7fFUUeRQLM9h1F/Oq1GiBCA5W+6kb5BMQroIpuFjMBii5tmZYXWQBIrw9ND2sGO331d8DxIQp0
fPo2DI4s2VZVQxhqay12iKI4P2vdQ8/4XL3TrKpj95ph55Xzf6B/M4YKaqQzwDR2YF3WcVXoPNtB
Y7JoP7FTiXvdnGTUQRL07klMRrhcV84DkM4jzmqHVza+4sEre761w/I54EXc3zh+q87M9SHbXPqL
joHBLV03cSQevNIS/rGauJBBpJnzdkEH8UqT+MERdzKpznazxdptxvlYP8RNNMELRfnbJJZJEapd
lo5wH4uklsOp3cCLZlfUJOYZ5EQOqAvho8XCqzbaC5VPYWZDrV3f/vwIt4zdpN5ms9EhyRVXwXQg
VN3YXjlLrgWwmufvsGXJ7VxHFIp5dNUw4IC1DT37VpVpEuMsHeVknWpGU3tQ81qgJRYRwaKGLDR+
Frj0UQuFeeCX1iEAWosxkSEbO3n7rI4nlblZJZFTjodCRQ0DJ2mue9BTkBflmcnoO3WonlqfXeNh
/H9fpUB6uMgnhyE5FWam16zpGvTQ8aQ/EgdL9/2ErH24Vycd1Ae+acsssSnKRlIVunlJS2abet9B
ItgCTWPxVRdxJXM8pq3AfBeZoGGE71u4tFtC+BF4YtQ/jC4b490Fxx9pdkCSDzqapHA7AGxXTnK9
zrr6nb1b8hZ6lnz9bNxkXO8GN4vXuHeHc8oLm3nIuz+T0ZomyAtV5bhSz4Lauv2L5oIteLLPeV9q
luO/7ZN2mOBUzH2vhxZi2H4/9kogxKYjHP4K8wnzNw7syzNu5GIfDBMg776IX+87txKb/WA5yuYf
gN8EFakDkTgF/So7DdRVixltv6q3GsuM+nzM/h7ZtNEYcT9TQJaDmoDw8s/X2xq1L80J9zyd3z4Y
Q1CHoL5QefMeVYXLxIyiI/nfExAc8VJOXgCoYyQFCzc2R91+dMjdEwNQhqg93MpRknfbGFEq4wpQ
SCFjR+FCob1FoYBL5RL6DMX5xwCS5VEDE3h3/Y2DTqwJOSv31xjmCNMZTsQa/PIG/Zv/hy4SFCKT
VULUdSzcPjdOcnPHMLUMLnu9T8mkn9Vc/JBOpo5wDqQdY5n5g2BuVzT0u34S5q3GeRAuAP+KI+FM
c7YEcf0bvcJqa4MxZEffh+1c/RF+Dy13XeAmpmdug8OjNAdfMQgdmC/mGQl4NqKJSXS08L+t0sxd
JtujuwQXgD7HX9dzYyQzKxLnPqa1CJkjrl/h5Ze+hBk8wc1EDH1p4DG9BUHxzDfxAZ/hPzJwf8wp
OMvLKv6FpUZnjNVTKyb0TNf/gLMCIfBN6davYeScxY30nBCPnC+hID4PJYeKYJwthPjn0430X46d
KoMkdRlyPoTRqS8wKR+aHzgc/F1qjiGBzEM1HidfVPiHquaHcnaXDjCEzMZSaHNlfnl5oxYUQj9R
0h4dGz9Ag1HK93RexaAHv6GZ+SHFolFiQwIfJo1Qz6uv8NdVbc5K4Xw5Xafp77DLkBbJ5XdMTikK
VgXKWukxt7HzmgjRd65Bk7GBB6oUWTHpjKWb60v587EOCK+dpbaslsfhz2sQ2BYNXd+f1kAmgT47
IcKF5fDVfEQawBpQPt3NOcwwdbzdWwTBZpLoyHdIWMw1MgC9SPUkzHtN7y6QJQoQNxcf2nMCMEc1
r+rt/01ZyYcgGd1DmZ1bum/MvqbjGM6OJqCmKW7YUs7EkABD6k1KeU7JKFZTieg3U3Abx3qyG3qd
Tqvip0fNXNO2xmtp8h8Oq0W6jDpQqwkzR5ioi60sB90MsdAwksyVPqAiSr69aXylSVZyLv1czt4N
JG/j9/oT8sxM8HDE/K/cuZ8zwBT9u2YB1aNE9NN5Yd4PyJogcn9zI2zyfVZJnheH7zmFjGkq9GeQ
shFvICV0yWnDnoDQROl5YB9EA/8JDpD7cjHPI4Bu5knK1xtvTtExWLzFYUFkpz6BxI5AjZ6L5pr5
1XBlKmNf8FmBoxX13R0uR9/B+pFUISdv0S3uVSvvhwTBpB/H4mhDyCWelK3cQBDvZbVWwuGkd5UG
3sLh+JjD9iT7+oIRHp+KbsVaK2zKr2KP1BvaoYs1b8pXKOs4P4m0NEbgFpBMDsiw6plheP9mmEnc
6EtoCnqrFvIOjjuLuIrmZudl/fQbKmvQnStJG+Ut1++arywEfcCJ6c1dxYQi4qu6ys3LBLIwaVRr
qvIP+IJmpDrBrk+aH3uRaqT6+eAaWpriGTkzuDOdtKV8KlxC2K/mT3S3a/SyGBQhccw4PUsGmQ37
0Pt7UX56XHacdBQXQkzr/27T9TiMwfqxE6IGAZxnmRkKdEotzOTGB7FdTJS+UR2XhBZN81Q8aUI6
neeVbExkTpd6KIq25WKhIL+JSCAe6Q6j4S7PS94ZuiAiKCQGPk4SvTOPFeMknG8+dlyexuFph9UC
Q/fct16lejJBUv/4ODYn7n/AAMckJYpkJHlS4LYZatqNcCGCAJzWMo2WRQR5mAEv7JHpgKuVX/V0
71ZPUFCdnnSjZ6+lduBpN1j3j0HA2agr1VpkX6v8hC91XGaZEv9B4XYEvSlSzlKttLCrC6rTgG5O
8ou4DDGgqk+Rvd8QDba7JLvFwVt3klq8yUD1gfB9m5dbw8tJ8//kfHWrZ2tNU/ZeJG3O/Yvi2Ivm
TiGtXu+EefZ3cfkyGzxemnFRhmpiFtuhtgx5Su6BXHGF0YA37q9sRwyJzUF+O0hvJu4w0kxnCijn
XUczNX9xSx1YzfSqeaxU4WMR8c5s0xZrJfjQkN3HYjvEIPLmKUKXk/aPuvA6MHlA3Apb1c0Kf4JH
4+dGLQL+qU9YdaDAo/bBZVhNsJTgjiADEC8J6Ec/uLo5te4EzPpKiyXB6kFdNjEEZMEnOyq9UySy
M+PHTzRKKsruKtXsgL9FuxgsPhxcMQYPumPh8Enz/BhudWugvwba8uEaVfLq7SBt0OYxQVLrvLW+
LP7EXzObpu3IUM+Mwmb6s+Wbxj4YB+u8ktlgKPD6Y9+2e6Gs51Cl/5m80Qq0DQouqLv7/W3gw4H3
TZq3T4z8plK2dvLXYHhfJFsu0PrihcM8sUDdPGL9I8rAHnJp8qVHAK3zZYw/cz/eZdmIdCf17m/0
ZAv83LQvBTbn6xIrcmDVuNI3xKIYyxu87uBVEBhksoRLIbfEANX0f87Bfo7qcrlGkuH4srbeNY2k
/ItvN/lZAVHoAIRi5WVHXTWVFlYGD9MBaiJKkdHVqDq3eCuQLAF8xhIG8266TE7WaDZgkWItHS+j
fADLmbJ2jF9i7sLyqD7lZxSuK5JY//WqkrOcefP4vhV7nUrvkkex+iYgtHRg4TjhtPyWaMpOJ8o4
0P3VVWNzB9iplkzzLlIv8oyZMoHFVDcN9/sOltPXDQaxklgE31a+LTpxZZkKA74RFamBmX94cwYB
ZGt/SIbsWtSR7r1+Hv3jsaz1p1VCnrx7w0zl9Cr1g0+f1gPjuSkfcwi4Xz2Tt9j49TYFxKcxW0j3
yvc4JUfRxaqCT4ZMSJ15SpP7R22YBH0dc68jvJ7mwaT7TGTmJe1GYQGQfQGCQqwQo5a6QgGs49ko
ZqgGy0cY110bVbyw8e8D42/4X4rxIfD7PAxnHoH3j4GL+eDcCd22ehmy5/UD51H+yMXdS+j4+a7J
lmqPQxqg0SF4195ej9badirhlzQ1ilIKwOkSmIPFuN/cSiZymGz8pvaJ3Z8/WTt4HRbCeh7ZPRdB
UMckmN1qOYavtpmomUtrTlqb/mnPYQu/5DUMoPABJsfQg+pTftx/1RJUNtZv/4v5PztVVUlZBZEf
vUxjVeClPxD4fZ7FRUd5CwHnfeGA4lYuaP7IjDEJ0clsXhPxAdrnwXxO/EAlds1WonZgBi/jlf4d
Pg3uiB0rgfnxhftMbqmYCu+WjnbPbZXoaMyU8R45L4kB2gyrAmKEL7gI2kv2SqTbJ/8fzc2smGWb
76gqph1EKNUVvvHy13Np4OQq9LV6+V3VFbrtq2hB0kzoQi4PCGZ7m/0brD6oQb3nw6fOKUtQNruq
9D6qw5e9PZKBYLyEapcxeI0pG1dLOTSA4j1kW3+QLmVElwfQFG9FojnPFeF0NH8aCwutXth/xnUV
GYUgw3Uhqnv45R8N2Xh8yQhN0iG0gDgzbk5Suy5fVLvZ9OH/5T6bXUwcrVube2FySPjJkLnynH2H
/v7xE47CTGNDIYbUpdfT/KMqUraYUAY9S+eZgxMSElEG3NCY3CPvidSWNxK6m+PKS1mDRPN0piAo
gZyR0DrsDNP2Nf0WRi8dTrnb6fEAswLhA+yJ5bc9lH8/KxCUfmWv2HRkXrHTbNp8Vxw5tQxvS7pI
Cc/5kcmcbNu25/6/ByC3HKwmtbao0At6OoE9UEL9ZvuzHIhfbe9JgUTYGzSJpJfEN9iyOjX8KRZB
xatocwwPfqPaejhvw8WY5jo1HiPTfzemihfqtFLTEFEw4HcPRFKa3smSJ6ufTN0LvHQPL/r6QVqo
jzxb4A8M+QrZVPFUA5KzVChOFJqyW9GdnzSoX2S8T9t0UQi9LXZbZXsaRZREYTrNBjObld3qAROr
BaeOxHcRMZwsm0t0JuGhAupoPn0PLnru5Hi5WiwmAWKC7wBUzMljSRREYO4F6m1rNptJjE/kSG1I
UZi5j26fT0qbWeEnFVqnXS7K2XZObYoiRwHW/SAjqhy+Er8/dbtCYoMd0cGuvgMVCp3+gWgNH1QP
4FN+qlnmaaOq2yvMrsC59dYhic9YlaHYZ3PwDDL3D7eWUn9vqvSdDsZ3Xx/2Pg6O3AwGgl8t+Iz+
cIIY2oGK+oL2Ex8pBWrHXonWIBNdeInho0vewREYsOzYK0X27Q8fNcE44aUKgl8re/+sUbRPhXIX
C7VM0+VUW3Lrd9HcF84mTUT/DYhmAhhkEdmNFMrGOzZJvaHoW2cGinC3vF1k4DSXgGlPkV72Pb7O
X3o/ceTafxwh5YG2Byw9aGBA9LUJAAPa6Mi//hN5LwYhvx5S1o/mTSaRss1ltFVBCg5sazSX1lhe
C6EaIpA4AWBbmpfk0MaNqZAarwvxGFb22htu1h4an/ndUGc59t10UeBDVD5+HMuqLl5ZxsUqVGkV
C80Y1N+l1Ey1GWG7vFElOcnItLb4CRvUaP842K6800hPJKqAKKjOqOBRpPK8Q74v1Muv80VPWtLF
s3fFtmrdR0Tgc9yP7u0lYwgxBS2tQT8NYkQKC28zl57Us3aq1TXFfXxqx+Dp4Qsdw8huc6TRxdwb
tB+YTtOE0v5VFBIJvVaASv6R8unmqcXWrf22SDEPt6TWDzFUOcHBKhdMzqD8CwvlmqAZCCMb2uxk
DdE7Wk4nE1JCajh68OaID7fWboEEYnGZPQUQgODT982uS5jyYPBHa2LdJs+1+V7AfJFczqgPs+Z9
moK34bzVuxy6Anc8MvfWP/N4lvD7F1SwQhW9iWk92P8wC39MJ+qJL2c3g2GmnlNkHlBa3nHYLfMH
lgGKOyszZLM0ytRZydVDE3SiEY15ANJuptr8+tMJ0FyDi4SNL5S6dZX0QiKw7qvJI8pYjpDc1J+l
EqggchPH/R3Ki9nkDFJvcvVOudBzWEvIzUJHR70L8gXyAolPN4AOivWOQEFjx4jdm5hVwhAOJiJN
evnrnSc15EIgtRjpRHJEJmQLcQVXq2kQbsStnOrOZ8lJecURZPmjrbDtsPyFEG6uDNtJCfb1hKjr
q599hSUpGTE8Yug7zKMfr+/LdPOm/ftzt2QJncto4/BxpVQdz+PxoSRTwiopol/S3d6hQLwn+aWc
Zr5ahJZmZPnwFz6/6om5pxvYfqEFb9s6LcVrRYYs2RTkHMmW73pzGtFyjB4Tz9OVtRZsB7zHgC7G
kOQm5JloERfAa1Y/GvvcG6pAX3wg/HMT1wFiccAhWWRopWwb1cYlp6BEUFSJxk4cQ7blJcY5U04z
oT40jHkhgSWEms0qFlZQ/KNJkylO0phsXfbPmL0FOQRo9bj2Zgq1/D6AIRnous9Bi2nR/KiedldL
hN1BHXLSwahV9b2qMjMT04SJWAkmM6WHiwiR/H6v7ap4GS1e0DxnkqqUl0HNBXEaVhkqRQlpJlHV
aP1+bgmeuhBXdIKKNipvq2KfwY2KGO7l4h0UeV6kCyW/z+86DJSvH5XUh2P0ZLCbhXDuj54A5rqq
bmgGXPZFTlHhgotZAdrT6T/zS6sbFyeKBy2TsduZatA1kaxc+KJyg7v/Dr+RlO4V1rnHGPPhD140
sAl71/vckJ32Ys6jEBtqikUrZMS1uQcikdUXdapOUqPsmsBQryAuAJKdaROk7Om2QZH2l4v7oILc
Gf8kFkW8z0uxouAPYtU/7n8Q+NHzL4oCvNgJMV2n8LmtShD7E1BjomrzgxuEkKmRbZlMv30nEaYx
79D5aACo3V6v3XBV+2W3mg3QBtyRfy6gu7zKcflqtCfImjoKzoecZX2BqZLa6rZ03+Aa0qyBnuHB
Nf7BDrA5biMQo2Xi7fXxCXrHKlF4PpnwA4FKRShT7UjtTG5yWSEInzYoAiMfQUeFQd5YyK3wl6N5
MWx5Rr0RGnwVg7DPc6WRyVWiP1SzMcp0WLCJhJaWWJKqSNAYV5C2DgUK9WUektaeL9dkZ6bCMB7Y
SJekVcsO3Yk3FLP6Cl5oDe3c1CLKVWcB/fMHKrRctWn+2tKP8pmF9gKX501ooLaGB3EkySbbfoyT
YHHrL2NaYpD+Tg3Gui/v1RA/ujnqknZ0rJMbTHMCHqqc0kVyMDe3PyzS44HJ0TSJZ850eXaqlJsn
fj0WO6HwVRL2HVHSrY4WIseDujPA3V1OpzxZAJnUxnhPjOpJGZILt4T5lLlrYjd4HjSB0AmHvwCZ
wRWwkjejR2Xl5d3DT/hEsAsCJBSGOzOQDvk28HEPODFQjIobJB+xY1QsjwhYQ4u0ryx9L6xPsdW3
g2j8BmX/A5lGTKckQyaRpFD4NnhS+fkfn/c80bETXhdAA7Wn8KYnS33C2NbjIPdL6dwiyowOuIw/
l8sMw5D8nETCeI6ff80OUiMNsO+bswaq69YG4Tmg9C69sKmyEZQD1E72oWRxnv7thuuGVXyovZQ2
U1s0Fom+gy90mODqt4E6Sm2TSOHURu5F/h3d+Q5hZBvnzfqYMqrij9EnmrnHMg5yjTivV1KBsvaz
VfrCVvBjI1GKItzMZOW8luY4R4XWFx3KfRT5Z51wK6x0YKs065CS1WiEmqD+pPaes20yQM52W2hu
I0xTnLSXtSjYycK5P6N25KBzgEEKHaZmAH9f0s4PdAgY/CZEuAyqzak5bOzkuQcbBhwwWjRW785P
+ijc3q4rMk7XGPO1zH9nB3BE7KyzHP+vZHR2sDlA/2NmjD8RWejMxQ8hOQz2Z3S79efM+In5K77w
IN2hnk3ZODUIYQ84KW938EL7Z44pX0nLPEnfVFKks+S2qkuzvvGI21HitU0DwPg98+eBeqtm5XPD
QXcbN0HbM1Xs21XE9ll4fZOVdnsu1h3vgkziOY12Mbs1bBjHDl1FK+sJwquhprud71Po2GhU5vrn
eKKW1OmUZV9U36CPKr+/c+253SLtFXFZJXaCsB2+rDN9tatl+GsMoB7NWMKF4bcLbv+naDJ95HGp
RLVskxnFBhxV3baMaJidplvUycsDjIB3u53dMX1jgXknyJXP6BSwx02oeVrdJuKS3gK3c5qQ/TXi
juJSbTDP16K1QFdGPLG+xs40w8KVBLX5UMoRIvyYKeEQR+O1gPSR39MHcxmlk24/dCfZIYlo+LYM
wZfGYBOIQLuYa/JWdMhsZcpc/VO6A0uHjbNvIAciyIUFaIqfULJqsTgowiiY6JNHuKRCnPug5PVe
oZa9Hu7wB+7uhtCHHGFPijPfV1KxTrINLY0p6SgdfFQZE1kvaYh/2sB6Q+BvcsVtgNSq4z1KB5z2
tS8NFJaq4kQ0WDlGf6LKdHABi/xvFtAEl5QlXtKAm87yD0cdweOij4NGO+fcuy6bfaghcfJ3bWgz
WkcOAcG20xTYdfSMCzV8yF/+YUWW3L+fCpJq9nQ5Ek/2dQ70wfIaDi/BH9Dkg0ijcObgRxiiXsOr
x5C6lwyVlmtsB6FHmsrYzMVi/XV9udG1R9g+Xzi6UM71AGhbeKUurBlFOzH2l84sk64INwCw57+D
6evZKXtAPnOfIK4ns8xOgDwA5aauinahTUFHanu9/ODJV0sb/sAR8aIJKnqGUa8TK4eg8CSutF8I
tZFYd9pFlpaolYY6h8nrUAf5Dn+B/wXaqsvD4f0pMspmdSMnriIXHXZ/anjUy/4gVNQ+BNCaGnNQ
z9m/UJgSIz2Lpf2dNsqL5J+HHoraN8Q/B30BHCDxjfayOINKGZOwljch13+ZQnetfTsWbsJ0IABQ
SrTOoEMpepnsbOkxWaGHQ6DYyFgWoI7TqgoS5bdFNG+PGkaZCBnJwFgyb9CL6jbG4gf+AtLmpAoV
5egveZ/E5vSlS+81EkE1B4iCUJOS11/DMbi/q4jzWnNITEcLwd7I0U0Dxhorrvo+V0nINZByUvAv
8Uxg/JbXXP9drm8AWuPDUjeOvH22jJ0+QxEadY5uSwMfmdPO/7Ryer/14rM6GwUpIz3Uw36Wann6
tUjKM03xizwcDTDo8KW87qVmfvxBmviQOEh7TS/pFJOuRqvGBZWURWBSB19ev8JTdtIvl78uU6tG
VR201YfvRfx819ZcsD2lvqguIAyEpHHHYhnX0Le4+27lQK5Dr0WYjX6v1ZNFWUvUD7afFTFR6chL
54o3qvokR3/kFylLPdW7OPK9gHxOeLWMbKmsM1CWrHwQYwgjIZ1IIyyocmCwjtmDx4IRpPuQh/+4
zoWTm2dmqn1DmOvXD1aP37KVMqaDacIJJfvDMkVeupQMJ/jRSpbEmZwtqtZzAwsuLrLEmrqH9dVI
6gtf5hpUF0Uf/zLxRBZkKTqF2vDKWZ6wWn5hxeaDNfJVr/+uphN9vEr05xExRu8xFM+BabVwdrln
ZmxhMH3XtueMqpkGWA2pFY02SdR24mHacheZZv9aKK5vHTI8jQvAZhkPW0oza6dP4DvvbXf9D961
bviWWC4vybx+vFP50VzhC9A9uWxMxFHpdS8hhjJiRQjJvMWCMAcmjRgVqYL5vznpb+xUcnAD/Gjd
JXG76MV+GDaI67KCo4+KQTyoVuKmPM1ir5V6HaWnlPEeCn2lhCSS1azmMvri/8gjK6xrN8+Wr9TK
deIMJVeOJCkXd2jQzh9a6skYVtSu+b+6QaPUUIkMPN0W5QYogezGlg0zKKYrLaOUmFf4WK+22rLV
70qz/gVDaYmG0plTEPhk2kYWVrgUqOaTJGvpe4YJUun70KVH5kqsIov4DTM6BT4hidhbdiqGuH1p
RJX+aj3ZgK//Nn/l0lOm5SetB3yx118umPn9uurk9aL7JAbuOiLrpoHhkeI/pueir/7vsyUu8Bla
5Ih5wyOOUy2yxSz5UzVsFdlE7xhjqojPgiwCsI50PpCWpmAiIjxwkHEWg9g/yvR6Cvnn884K70ys
NXcX64bFrnnHg7F2dEKzdPKiizgvhQu+qpJp2SheEQWKDlOeS2sD/EPpgN1MZ33s+8DR8jf3u2PJ
KTdImvxypAwWhSHUxnuK/pox385lQIpPxmzcpXGRhqOeyuGJc02ZxaJwZ/PTvE8jqt7Rs7m63I5D
Ya+2ZDpisR97GgpXDJlsfcGXOrYg212gSQSj0LzBOxEhRDxQ9C7F6rlLKFGU/V+nsd7D5fo8aPQW
mrhs0Ny7ILpZ4sRFjcbx9OLj/KBN4r/ZIfP6nSmN/s5jXiXKhnqbE5t8GAevXcmVb9RJjcbOCImH
GjweL3dfiUo8UKDjGUr4hpIB1dGMHvOgk/xTkElJgxw+EiqdiBggk/4S8qeCe5jk8JVV3uFsJ0PL
aqs9Xc6XDbwrZZKlWq5dLUMUl5lvo4u9jxe60mvYUom7Rkg8Yoc659FXJUcTYrDb62UT7rYJ6Xy+
aT1VqpD3c5O9ttiFYV9dPtBEZDlDbm0cxeme7M9z/WrTgw5pGROawxSsQzUIjvTdUR58dXp2qW04
kesujkxCtg0XhRmaNBxogv7hUKVysuhhf85kNCKwKW6J5gtA1W1NAeg2gCtaFIIn3UlabP5kREY1
vB06CieLVuB/IfJQ2lkRJDQqaQlMXvZz1FjYS8SVzQimimfMbiXsZL86Gql5rgxhfpd3ZiRXw393
efhs5CD+Nx1nW03Y9dgAZ/OCQ8Xg/RTNxZmTqihjfG8h9izASqiUSEWkK/xMzjj7A7ZTwsjsxm/9
9z/gcqIGnmm41NN8uK3a/3CIxuvAE9b1q2WaDxGHrx82KAJPtDIVE1Cxx5ejm9V0yH5WokuHYPwN
xAG2OSyAk7pp7vnvFXCztQlEM/O3efTVV01k0M1CUForZeWoe6NXnIQk/YckdIZPa/NK969YQ9QM
muHZI/SfkhV2sxto4DkJN0a81TpKd58qigI1wvY+XkOwV2j9vUNZOFWEuRz3BCUpmh1H5wYhlsY2
ypVTrBMH5QvWKkfYMvVHMeKuf8OgG91WcG54vENVm4OFrty0dk7QB+9d81RwMpshZ5qJzLZQ3uPO
TRfh5e680GubCC0ocT8cmAkXd8zo2Q8trDLLBKQiuqXgOpLUKjBErNnoFNwZl1xaTRF1Uc/dg7bv
KCML7rmDhLz3Ry1Rhhe+b3o9VLHwtXW2lTK4LdHhVyOarOawe1w8Y0kwMTNQQoSdzlYaUNtklvsR
Hc+ozk1Kgw/BzrY2fj4UMq4yxUQ/n+lXJywNZSnb8vzXW8565D/jI2WIPk5o+GY3NXAblofE5VK9
VHFCZ4oH7B8RPQxW4HkP7vmtm/lxfTrYQz3B4phZvNzBaYJh/ZxLlescY0N9i5uqO2bYz8/f9ElV
22Luw+tRWTyI1aascr1KTO5u0G50YDtODvTMUuRr2hTH3ZhpPaIEWif1IzGjOHF7TTiqH3T1xfKl
ckLkgZh5dermQsEYf7BLuklzR/VEj0C5SaqfyQIAOBL0jD9x6NZZlBx7cSUy4D+/pre2ADWvj/WG
6rpIyPo2ODe6NN30fBMz+vQJRa5Yh3RBD1QJliA+xfVBgkeK98e7Dbgl/0C3abZpFutYjEkHLfjP
JfE8Owu0hCWblfGfwOjCBXNw9IBYHJYSygz03igqBYwG5W32LumkazHwDqEjd5+r7ykF7iW6zkVU
3IhbvaQx+YxUpDb/q5gaSdlVYdOgkM4EEvg5SprgpSplD6x7xx+1J01ym40KtxoqGvk2tNTNhyez
9rB5K54O6XF7mAMtpa5I3YijvMJdi9PKZKoFhKgdn+5iUIc0LEi3Mm5wPa/wIyiXMAbD8ffL0QIx
gN6ZbU7n0dyjgWWWOSjUIG/+4ZXEtWygdnn9o1WHXM7etDuvPH+rF+lafCPq72XiuBOLVJfjuSls
WloV2tT6J5zHzaWkucSCM7fexQetxJKIw0RS/wpj4sAK38yPhs7bkoALm3K1RujdV9FRImOzXJnT
R969QHoBa4aGjG7itXbqB1ZPZU15x8RUjFhKHvbYJsT2MSVIrDU6Zy4bPEmEQ37Zg3puWWvZ1Dfi
SMkx/TOyYF+OhbHYXdqrVjXmSPpO44sflI2GkY/4Vba6Y0Je2r+5kWkIBiBGbNfS7s00vDhVNNHc
TCeh87VVR0YfdVF+HsI+l5zG99JyFjxZQ/nknxiOJCZPpwNvgfXA1GIcgeis/72eHBWJw1fICrBT
wGZBYX/4jQyVzYPLT9/mBl7VPZT+BQrPQzyhx7kNs8IANrzyhU1iNhyH40t4Pj/k5tn/NF6cXLbG
a+2k3YsKoFbVshQe9VFTqjNsAZu+v/UfKj9AIaRUSXgCOi9ueyoRlAHgDne1JCU5yyio7LxgbRrS
sqqgcU/s/ezxBBDw/0ntAgYti40L991TpCOIruYZUcYDTvNKtiuBx86hvce8NcVGMXAeNX81UaJX
S5NeFFDA/+6xaxQmfV8UWJ3b3TOMFsaEfTntAw+GboUzdfUW+4IpqGOp7/HLHmYDi/PRI+lzb2UW
C72zZZsgG3eHBvcvY22wOjfkBgoQDUuLHoIEJczv+JOIncS0OYQa7jFNHTj2owRsiEmYmYExxFK7
NfFqCnNqeBETvliBFhCuUOvM+n6zuVD/NK87KV0vx0MgYrsAMLhCcitD5B4D8OVslBohoVl/Wbfm
x3AyzP2lgKPE9ch60syfYmBamAhYA3nlAnDQOHpL+9/b8sXI41end5YCgVWvkAz/E6hKAz21Z8fR
CZNSGXfomAqhFCX59SOTp7+ElmMCnTCvv4vVQ7lN8PnCWlBPWUgY3c8hyuew5WnwmJ+4UCMfKq15
feAO8qM9y1kp9HRLe7tH+aD8J+lVl06Je7acsk6VtpcSaAXHfbxwWXlUWPDEIKyXXWDP0L4DYP2z
Z/At1I8HoL6BWqRG/OehDdAMZNBMW8yn2EtZ1GDi6wtS89rcM0jbOPs9v1s1IgsMFR+NkiDY8uv0
vsWeD5v1wyiYV+9Lz7t3JGhcLsi0v8oNoRujTJtNsVRrmoWh6p1wSWe2imsM2p6OGfOyVmzNjufZ
s3KaUC+r0/Ed+/xdreMDstKD/p1qYqd3VuTsQl5voepMJm1MDSTN0jxtansnw0+gFbD4PqU0EgUX
qUqxd6Pp1dRKE59ol9Rwlx3aofYm874IErBG3NAqJPzciLpBHUjtjOa/jO9jDjWE32lA5jBqHQGv
c9Ub1OvaiBvhPgeGDckEm3mcgm133hcDd221zxYqGgx3yrWed1+EQmFxwyptffNkcoIq5i6c2sKK
SterJag9yBPugtednS1KRIHvYUFVrdybyvROxiBxd93BGfpdjy1rbTcF/hFCOkRLYbYKHm3FG0PO
jYRa2ibyiLFgmMKomzwtx7dbZSEglYEKI3EEZ2v0jTUbgKRuUYCHV+bjH1NQvqR3AsSq+Q2p/0lW
cPaNZepeaAJgi808qa9FMyuF11jxOkuuBfBAht4hXPgzMCrAmnCQd2/HgeRsmoPz0q/4t5FdrQ9H
P5kao58EW2ByRYetO7vqadoR10bDDYUlc+zxiSZdTcDTpYOcrbDspCL6lio+bvj4q+AgK2laIFnT
8o2VWXrwFsCtsnNRsuF92TS7EuwihHBeXil+LtGNe8xOSwg9Z/oBdoRrhG4tJGKYgVdy4nap4ZkJ
s9KENYEOS/hEzxoQiG/XpMzswscPzMOvwgngbgtoA9KlLxZNvdSflFxjU4EOx//uy0oyMszv2izx
0rJUpW35O66s9kxZdQJIHXMId6nZR7r+Wrh+XPQsvwaGjZKD9WhIVVv5es1Q1Dav4DEp7roYVZW4
HCujJNlxG5KSU6lYg9Fds4t278yFmMJ3mjpOYqVIlEHs9WQmfY5HBo67TUyT09YuhVdCbxI6C0Ep
Mq5VZmwwR5z6THQ+zHJck0eEQ2kdJKT9I/rVsdj38DIsCyi5XZ8lpOMyrNJtYgx8V8nyfepVrI6G
AvMKxsWXAQbUwaKjAxHYThack50EJMeq703Wsp4DDDM4nwQiDG42G1FYZt858FmC0FRTY059mYqu
U+0AfDYvABHsSHPnxO88ZIfe3GBuFZ4zNUbC7ITy5pbYw+V4fwpgw8/K7cT9npRV79NxrWdJeQHG
Oz/8GpbgnlBsKQvCWxtZG4DSZ5fOpgSsyyELf8Hri8jn5ucIy1Rhvzt85wwMGioBGqpig3xZ5lcc
4xVoyJfGLVDxNZhMwPYZG2mXAlJVXgFarbzVb0mpG3YAmSnS2mhTw2aUOcDNE3dRI02aXHWSPywu
4z9hWt4FRZ5OLZ4UxF1WKEJdDbXNJi5GDEMtHYex7qozd2r4GbYo2ETmQqDImeal6Rd5sWHOuiLw
lO6xfohEXGWBDB5O88a8F+Lf2jn//kqX+t4k3A5T0rmbDH1VfiXQznpS0R89NOZiPP/A68xseXv5
e9b49IlctoxxNWfXng9cMLzXMUivQ3LH2g+yKqmW3a/g0sN8MAmD+WtQ17PfSIOm2ucPbH7PaTE4
E6iWx2BLPMcMtyJCNx+mKKCmwu2JsHQr/V9ZjCIMxVO0h6KbPr35UD3HUBDxdo6fCRoGkJKI7lhD
iXqJu/sdgpaRhRXtyXiSWHmA4FZa7agddrT74l/X+Qx87jnXqSjGpALmWyM14kSywQP2Sak8VQG4
g9V/8NT6zen53pbNV8L0+sdn6XnAxcJKDD1I6ogMJFAK+4POxqatk/Gt79TpapsWl9YNVTsbt4iG
R/xt8J+Lngax0Dplbgkax+InRflflPApi9hYxFVhhId/dVlPj36/1b5FVlG4EluIESecUa2x0952
i5HQBkUfVIntZqqeqjCIiB06mOCUqy3b6lo0AMIlGhZVwRZnmM8lLpLub6oH2yZHx/sF+sWkEACC
BDQO13A8kcDSlP/wOTqIhvICKkak5h2mgfDabX5WmvkWiKGUhEYsnChOJ8F495BRiYamAgWfBbzQ
OgdkIchrDgrYIupvBE1xab7K1srlK7wBp9Pg0YmK/+kgmSswUORpjvt2H4q92F/j/tYapNpXRsYo
mAwHZ+T4nz1DJL2U3BRgN1wIj8RaARIflsS0JvR65XXFPok7F+zgbeypj0x26Hj6EuKEsVw4I0Jj
/LS7AwMZqOP6sKZHgBv3AZ3bZZylOx+pCiYzRE9zwku+hKwsh76r8l76PPIfyOtnZzUq1NuI9kOb
RU64MbyvDbkgXdYVXn1yepGVGtxpz/jlmf3/IQdaXKZqNDzG/QzDaRQQu5tAKUOFwJGaB1QshbhQ
cDoRfxZhfIOcHzg1Qrk60ZxsQ0X1MFdyx0BmLR9tYRT8iK3piJO9dmo2PCJp03DZ5RrbHLxNbcN1
RtP+SApKThVZxq38OPFApdZLCb+68I0Ll7Z8JxnrQsm7Q/An+c3OjPnLsujvxu/BPOp/ORRhohd8
2vrfraWD+r7uoBqBKSs/SHaLZXXQZv3n2v2pxarZu4+mSTTQ9RYacZAb/HxoC36ZRtMFMcPirnaX
LksK54nvj4I7y/C3C8TkeOrOSS8WXIRhflq+GrQUz3KIXx+vNQw3VtokYHM0RHT4VNg8GjaTYIyG
KPq5yVcYkmnRGr4ztgzxEIA4fLYlLo6A0rEx7JLor8ryxk/ClgCXMLwREEOsMtgm6oChzOb5ZgyS
IZb9sJi8QbuDOd8gpjUQbnPVMoMNmTn/OkH/9zWPFxuAebviLNr78WtSr5ty9cAaWcAFynn4UUZf
/O61X+b5jo8o7XOlPNlV1tLcgXYQQsQujXitEyKl08qeUF/b/lKeqvfVQ65vfgxXSu2EqPe2B+ue
ioTVszD1UPJj7QiFNiX+G6vPFa4AJCKSCYJRMQ8ZO8oiH1O9e2r7jQo2q7VHptJRSBjb74Ql9/vL
Y7X9Hgbv7j8bxhVr1TsfyLc6OA3rQUynkKUh8S1j4VC5CXP7sDHcLJT8rnN/iDjjx5KcARv3cNBe
kSjEC5s0ojMQgWKhyIw+7jcT8b8j9UFQB/IRt6ZsKnM2zeUD4RAReTHOzd2isLsAEaC+LyHAn5/x
IVuTYblsGRQwN2v7lGljSMOIxgXETythyH23Wsxwk75/UgGhyIfd7E4VbIpDSPY0Hkv/bPs36k9D
JrpIZNMvhzFH1SerIj0BN+MKHg0yZu8PeYyjHvZN3nCtUdlv18FD/GORl7NGS36k5uRoN8R4q2Y8
4O07qpaOzdKkkbf0VKoBzYQYtlgKVO8/JT+Kvt5sAiQLH6sl0m3bsZXDFxB01P9Wbq2vhR1XD7jU
oj+KVGyeafr/D4DzODtUjlUfKYug9x5XTe9RHd+CWgVHTw7trUyS6s3CBnQdX8GNbrivnCyRP5ZK
fq4gc8uwVkC8mkYD2GTrBZvheVJYTH/64pjPAXq+mIv2TEyf9qpl/2HhTyaYr+weGydoTKue+/oT
bT8X5BuG9Yr4mQ5qKRu1mQdFLCirH0qPPE4PrZYoXfTUDxA/Uj/wteJ1YA4F+6SciTNHsoak8tnM
8Laeeh2V6uhYFwoRX59YKIJNOR0nAxGgMVfqgfsp1CzP0/UfMYxh/Stw2w5i4VhV34O5ff4YowKd
uK4/3e1J9KmN/TA0VI0ZtfXusiiWAxFiCmDy8m4GMCg+yv+3Xi1x0CBPQBSkfrV8Pmm6xJ72md88
8U0I/Xx3zmlqi5dyB6ZmOL8mLmKVSELHRWXK9p6CuHNPLPhhoSLhW3rEocdCqhHncgvBEbvuYSIX
n6IENONgsf9aFKccmtaGuIQQhXNVl07Ol9gYiU5IT0a16IF+q+Z4sIDkxLv1mwP4dMldPnS4XBk5
wqbi7JDkoxpVq4IvO88/XWBbBtVTsnMMkInNNpcotEgXHCAMkUrA5xysoTvFHMN9aXOKyQmdB627
ybIDEzAA7K2FMIro1uFSOwWGsh5IUv5bbccKzdXKnrpDC597vjYIOhRR1BkEWLnCW1WzqmsGOWvl
O1ajyl9kvq2P6oNRZRowwP02s48seHUwOwVKjSkB5xdAPYxvGhJZPLbDOtCbXcMCjTr9zd5D1nCi
N6DaowPtRKJ4UXXhGCfByS8C5MMC21DeKQXIdhUC62sMwiojUTWAW40i7CaO08990uCk91x3HRLb
M70FwUO0HQMIUkpLLN73muhk7aAiDWj9CEVLhvYF8BllzuPlq/nDzw8y+acdL9wj2nmR+oSIHqOU
imaixUeeiLnz0Za4ilXx0yfNBB+f4FG4+5f71NWYpl+O3ec5mIqlwhzelM0ku/At2vRP/4kq0d1F
5RzewmyLrsMRTK+7pCSW+jVCfC64v9odQQ4ZCIlZ8tOCIGnjjZdb++wCeCgnQETI2TNtTFSpBdMG
gIHfJWl3Mqrh7iNgQFuS3EVOQ+7l0iWv6SToNl/yi7tPh+uh6nVTftCpAJQyPoxMe9zO3cSwncOg
rkFswrY8ai+L15ZcptvV9AwBIhlp8smagmnLop2ZuxDwTp6oFyg1qcJJBNSeOpJTfINjhJRoqiDV
k6m3HqLG6OM0aCdleveS8XJuE6hK8/QrPA1ah7OOFx526oeF24wkc2lhd+lOIp4/4s+Nz0LMRQXe
7wZDfyBU6CHdXxKqgWE79Qp/VJgMjJfaAbYEZFyVuRKvHOktUYRJoSIlvktEH2tzfuK7+4S+t6F/
z8j/0S7Pmbr8R0XN0QKjaimiur8Ppaz6dV1wMNepKX1cP6rsWdEIzgQP/kn94NL6uTF5WQSoiSFO
2zx59Ru2sfa7SlOQd+OzDozJ7KDItu8XTalyWzNOFcKp5fsLUcku4kh1XfbaldJ9FEE+5rQHPlT3
wJICo7PnOoiApMXSlvj4QtElQyDVJ6UmRNj9sA7nrOTWsNN28u5DXGj/MsBCXLgXrGhPL6YGhwgD
Rj9218UHbfXB/sMrY1RyUOfK5drvEJR73juZBIp3yPSRQgya0FrjiEsxH5r0fHfZZLeuCV8yqZlD
wqoxxMQPyF7GIU8S5C1gME5mvsZvbaUnVGfsJvBk6D5RXyGmRlQ8jwTg0Hpg8PvWEC7JQrtSUkLD
Z17nuzPutilejcP1cfEebqcBEPeDIxe7Nqbi1e0pua6QoJ1MTulRs0bXyzAD/AkW2Ngd/+31neK8
dD/cSqmiDpVrOV8AXx/UZAzsRYJMMe6Sk1CvWuCl+zx7toXy8hkzXhmcsOSZiR759B+BjJ+yffFe
1fjxXMxobqsx1cD+E4iBe6noEbPfgFv4j1un8ZlnY06ZTqzMbg06b+ftLL/4BZS++JTeri/LvOZD
P3/xMEjkgHSk/oBMy9BsnbpbATyWPgEHo4BZP0IZviECdTBWkttM22UJu9wJXKocNPV8CLxH4fJw
kqxkpGlRtoGkisnJpWjPrL9IUk6KpGGLHYr8KJMg/KwNcBJupdcEBvYu6n0hg0QA2rpY620+Bioc
wKuWVf1rtVr9tOdGPgjR5KpHHMDIElvagyVDkgroUZtlu8GydYLQC1mXqyXKyhNM7Jo7GB9gz5If
tTkOU6D0vBWPr2v5K6KaWS0Hnysf++pf+QpWv3XzKaFwwpDUI3SDy+b4QaDhNXTSsLUYzazqIwNP
pga3AFfu1lrnnHjwgPGatT63q3D6V/26D18uwGUmi+stcsCGC8nXjMs8pReuSCenDKpFutF9k7er
ihKcRtT68hGA4UcuFsqA9+2q0Z9VmaZSzOwm2PwfJvqx11kCn1ZJ4VpZ1FOc/4W7x9SVm3lnAsK1
prpClb9lbken7gJqUbzXWQoNsGucGx6EWXzkOU1xo83BSd5JxDrMfXq1ybj2FmBUE6sXc078Yh2U
soEWsqr2VLdb3W5uFKxaUy35T1fH0szt8M4ka2dZDghWC0tT8Pu+6awWkMKegP8qLt5CXJN901Zp
QabFNmwPI+U/+W9Et5kRPAut1QdXynwQzl4NsW8kDlJUJ/6gjUgwf3B5WB4elNi1XwpMBPdqx+n2
cOSacoduDmenHMPCtP/x9lYlNwrRQw5RJLGTjYfs7aUkYbR3DbGvZrLbmosV9iafxfd/ZxdsCUa3
ACRA+3Sp1vBA4QoqYvZlzELNsslWSv3GPZHQs4puUz7qT3CHXQ+M9gYH5MQs08c3X8XzRQFzJHmV
XoI44SYIOjBAf9taE9I01QpUN9avp2r9dK1aNTzPlJScQPmvAxbNvWIWLPgg6wVRUyzPpLSRYrZ/
/t2pE8MXxp8Oxuweh7EKBtV5cF536FG3w0mxA43rCw3NRJc64nFFddzMexmKp2b57u4Y/h3HbR2k
qwHazZL0SwwtwthAK3I7JYVcJO0MOA73anUL4AvyvhJdRr81D8LraE7o45H0Y/umBVChYu4iTCn8
eOakk5rESk3a2Z6CcH70IpVHGI5WrD+gOf22vtn/KhualgMHv9AGvLPyUvHwnoR98Nd+ThRUfl8/
tnxVzpvO+YNNjE1nDZeruIzZc2pCWiu9XVOfKcXwbMeD+i8dxbqPM7dRWmIBKSr0vGgT/sQKcI8f
zLValSwv4ZsYAgy+ZuKeY389F7F9BINmiWybv083YrrbGavZJ1FgLXYHmAp94u/FT8RcVCTuYezd
W7rCckxcWzc9dv2XfPNC364BFf6lgJsOaNVYl3jUVQMRuit1zt638pJCnCWxGhSCj5Aw2kSpTSO+
1j/LNam38hlu15rgHk+KEyzLQlgYbY8zNvsAPk0IN2RN7anyyhZFuPG4z9fnlZfwIH48cGJd+CUw
gywNNjji23c3dZkHuKDMX9JQJ4teE9o6Oamvgr1oNqLdTVO7bOmjudEkTTwhU3IKwQrXdzYd2ShJ
jrbV6wAkOJRxnRlaV4SXgW4XIUtQf/bMj6E1ZoEveMDg3YTOI48jYnOCKzMEAAJYRI5d4L85cGWE
AJzSAGrWa4m7yI/DFsiOLHuZOk87KWQxx8DgGvp5iH7m8Wc4hcofYMwJ9bL2Tfs92YNz8dO7jndL
iZ68IZnZD0R5W4BrLYW7G97YD307tTvzGk6L7OXUMw4Lp3LgmVymURUZ4/wutzhQOEbC9dThwKsN
LjZntlw5j2KzK5hRDN0PjzqmCPbHAF0Gz71waZG9MBtg2MmDwsa+XvNxd19cpRzpH2v6PK/ZazZO
zi4nsjFcsMsKF73EvA9SWct0fxM4I/XOmEopUh2pTRf69bjuwoIYGVGiuCrGJ/8UgnrtVr5VzcYM
zO0LKMcNgj0XiY44lidrAV43zifLgdevtTl7j6DciRrK8vQELzyBuSLUaXfzxHQug86PvKGENQ+0
feRTXXyEbz8HSP3enVZR79Q/GhoaYjhK4XVqmYZR71XEwQjoKwRcnihBQtNf5INK/52jfpLz+ibT
5mRWM8E6RrX1jM3QlMHPuGEykwCtzDrb3T+F2HImI0gJdZ3pVxPuYY3l+GgEnNd2iALqXWAmTsow
2wC8dkzOWaA8h4vJh9yzVZH6HA0AUbwXJLHH1O8dFRSla7fFnmjh1aEfM+ToYxmuWprQNkTCaA58
xBPyGgJjVYvlISKeF/XVQLxvQGHQkxX7hmE2UE74KDOytv/7DuSfCSDzUjI9S6Wwminb7UrSK67n
+4XCmT7ePd41i1mzcTBgDFRX4q2gY/5dGEESbyzCXxmBajutw3Uc8Ve8AFrodP9J9E6dhf7axe1M
JACOjMS3iol4IpXXRfrwX3f+N1aqIS1v7y9Ag1p5USX1F7A0Uug10/ZGuFgkf2A/fPt8ht8pnyEq
QD8KhktUXPuemnVbldqzMrZeTexuc34sNoMFA4T8EDRd5qjqDaBtfGvq/mZPdm/+TmLC18R0F3s4
IY+XcuklWJQ2NKPRybm5WYbxKKmc2sBC1lkQoTy8Lb3tXiqErggktm7cOdJy+zgqYoZl38QZba1y
s2eRXHweVhVslrj2oqP0Ni84yEyCA5pV1HNmcUNvtq5HMuiGNALtj3PWLfdLV0eXqauJtDfnOAYQ
QAyAscTCzlFcy23H80qSZoiPspjWKs8uo64poCKvwUdsDCZ1PI9MqgkLKYLZWDIJ0kCv7dAaQz/J
l1XqZKBcM/grl0F2bhEx0LOHi4Kj1aoOJtwZ5UkgaWoUhl3UnExzQ8m+JBHrthEjSXOf6+wX3ptT
xOZ+0XKYk34TPVeNkRywKUmqHgpsZDnyvEgWzjBP6OJ7QOuxvjBQFZ/ubCF/O4Wjs/6GAgh4X+Zm
XWayzOs13piAhz9dEJIIzQSUH0nG8HAgiQl/ysn3M1wFvyXLKNaI7GeyigWPTallUti8VnqGKCY0
yapU4K+uXIqjFz/pcXZ28TeQ9VuAhRvV8elmpKNBpoy59nDGmTRKh3OKDlQgRGbH9PHrfbMjEAW1
JMKiDHQ7Myj82x6XE5aL1T0moo9ldXPxAGVgcyvc0iw6ZF7R11flM7ESoHqfAScI5Dc5tH77xxF+
gcCPtLUh+Uo+AdfxVccXzJ2fNfBf0gBCecEgledtXS109xBVVSUhb8bzNw4CuwiWrLTTXETiWx2a
GzRudZU7Qw0gnI8H49kQNy5RcB1zWTLP2CZyUKlrTDb1JHfe65iYjpRAE9WpuvFD81d+/4Q0BjJz
FxT6MUTT3vZNt7UjzKotvSszHT+4yZD2lVPl6o+pe+hf0DLe5xy5EGXJcZOL7hxhs4o3CxOTEw7y
Yk7BR7d0IvfHZJe2iOQZeLNb6042wXdDn+vdBg31YIOk9QPLNUMsmUvSGPH7sutvu2IzbPiZvPQ6
KzEFU4NephDScuVrGaD29nwAnOGSUHqnWP70OBGnros8XE2f0Rc66TcM9dgGfl88svcSAUB7SNof
YH7oDWuwL/jyTK72rAXw5s9Rlg/Mp0kM21q7y5XBqmMR0TyS19ceAA4byJz8QjGnFlEfsEVKsf1D
P0tjhihdur24lPHg9ZT5ndQbwFmBGqtL8DDvH93JDkXSTR9vX3VTT05KehgoW0+nWCeBvdMhOMUm
CKhMKhdHmrRIJFUeUUioL3urhd8NsOalLijF3D9rMIKOLQmv06VhFzfGHzm7zLmjBNvVikJp8qOa
YDtQQ/pzyY7h3MbATglRtbGCDuqB+QJptO2aqjBVCkJVmYaW64FR9ebFvCd4d3Cp0vCEM/x5r/rv
OUTY+AQ0XrZMmiwnbiKJX7uid7PclbUFxmfILAI3ys7GkQi4hPjvw1cx+S7iC9Pa94ddJkwm6rks
4+J8A5/WObn5xYpHKscEOTcfHNqgkl7sDBnwtBP4BJ+JiAvOlFY7cDvPRjt5h77RU79XLiQMNytv
V6i7kgjjKo0aANyYSBa6f4qm+/aVfQuHe5BVvOT5IA+L8XW3oPSB4/YuWUk18JNz3gOCdIomFRys
YktDBAG2uUcop4L/6em6dN0cQa0Fg2Sy0cSKgcdExvgjYDUKzZCaaoLC0i9CmJPwhaVi3KhniDR6
RgMQd9AryQy1H6LXh1o1y3Y5xah4S4C1vybyq/7lMizeDzJalpqO3LC/rY1ooYUq5+RFIFxylVMY
ST0I04TqG0dTR/+qYtS2tgqMSPw3uCD4K67DC5G6yXk4ymfy78bs2hy6ozgdfdlpT+b5A7/LhlPD
oMGrhEpTIbOj1wPfonnbSI16EGJdEZKqvRja2Bj8Vzgr7E/ACRTmDbNW2K+7SchOm+U54/HcOe1J
ASGQsg60qvC4ngtZPk+DLjSVjMCmMrImOePxzmDeO6oWfa608LlSZO61nViSyKS19/P8E6thzQpA
5UfGX4jvZ3j8AMS9MawNka683MHXZxOTR6BrGk5mPIk21TwwNQsmIDiVrCJsdHw6C8/uz8RE7L6i
/619+jtGFp7Mf34KF0MWGcVskxfm3Xv7jz01R2G5bSL34g1T/M8d6eeHErm9SLtPCmJg7mXCwoS/
0eyUHIZBthm5RC9eO2vSTJLmWLJ729qqKIEuaLxMplh80O1NbWifwdaXnck8bkj6DKsLwzYC6Bo9
I0qfI9mmbJZtiW52qquCGJ7KedWtOAuFKvSbF+GSb41BZ5/SUAiSLxUBEBjrg/fQVrZhyRoCtuLk
6kPbhEIgeL/cOnvGEYoQYTDOWld3xSXdt60EzdLNfLwSV3F0Wdci1zn96bUTAlYRE0ZnyH9MM8sQ
ZG/VivKkTQ7dXA2AbElX8kgtqWjJKtsHXr9WOl3RjVQgH3LLANi4tDff0FjtGCJfycv8/8rbg0Ql
7GTsLfvCONocaGEhaGJbXtJ6ua5fVqRm4AHx8W7v7M89b0z8rKRMbd+Rqq8oZRm8z+ybfeXP9KfX
NxmoGQg0/zTiu0BuDrCKE4ZmR14RW2Rg/lO37DdQffRRcxrUYb+qqi3So46K3lkJJTv0+AP4EDdI
tulheMFplCN+x/NOS/vM+JmhERIWyngWYtgkV05NMQfmLoWOTU5H3e1ZTPK858caGiOjXB3pmysE
X8T5a/JC/+ti51NeAAoR46ttNg9F/x18nvIa27n36zS9GWls1K277RsgD1ACVAUUcLzFKH6oK5ed
5yRXoM11GSfYdzy9dbS2iJKYE3JFZQDjwDlbM/BwHVUPUE0NvaxPUxRpTGFVDO6nwPq0CULUEEDx
1j1cmVVRdJn6izMjw+48EaUkuBOOmQZvUhVlLxLeJN3TT2cB9ghmjHSFot+GkIQkZdEDgKFmE7MD
yVFRoCnrx/1lCIAKpxA5p7r4XJxH6pxIhX3AH8ncYMTCbe08glPXZBw+ARxuwUEcPsN1eQCild65
TZDtRl1FNjDW2HbHJ4p8Q+/JzdwKDem8+GJh9bWD4oskVzvEAU2ak9Fm+azZWo2no1PjBju/9oRS
nftbaBhpvJFbx/jP9jXmb9HYB3mhyNLIliy4HcJPujckPDk1g4ExxterP/B3Kty9x3+jkLpMyQrZ
tYYOseYyQhXRboGMfqjLqxUE760+R0yiBZBb/WaH+7R5WORQyDhkaOFJz/ToETsMYhBqm+SZCF3+
C74iT2f8uba6jzXIeF8+Z8b5AJZttZ+n+7OjAKHRs1Y8BnGiSHVDL9rgcsMvLGrRdI+psnrqLnn7
sFFifrVqaA16U6v9TlJqDa3/ENvwQMmabIMY1I0Jjb8I2/eABFZeUTYLw7JKJZQAERTKHK/ETgVb
LdOqiQSl1klc8txQVA+RkiNhKBg9p6y+l1Ftoafa7kVL9C4H29J5Hkd4gTDWcH4z88CjcATQ8WSx
adDMW+5sB3RWMiyk21JGRNUh0uqOQ+XLhDxyYDrWMQr8+uIgMqCBrTJez/2CDO7XCHqTrN7E6QZ0
uFxOuaNU+ochAjVR4oB+MQhNTnlPFil+mA5KT+md4/H12E97j2gLgDw7irHUDA2apO84hujneT43
OWcbjefTNir1FvSPY9tCcw/usSCp8JlgAD1b7SahDcwZ6WIqvIyrSIo1WPTDtsNby/hIk0OvYMmC
YQYVzn9T+0u71XBRAErvjrlXWENfQRZpSlKUXEb0yPWcOEQf1ratpqPmc9YGpRM+SHPN/+kAN7j+
C+N8jIqZ7rpI3sgGvIst1j/8gf28zd+eld5fNEivwefr9J2kBp5zS9TS03xIohe/Tl0MkgdfiEPl
Fd8EK9bys0lJqA8rOvh+oKl2aR1KxP7+SfeT66uaqiPgIgiroOutMZw1JcEQ+bkZEzZ0/7zUk3XV
enhFiusaP4iRUKnmf//Oj64X52SCNmkCtJTm5pIagf7pK/NkIztrJQT5B/Ym5eSYBF/AmhXhbIqr
8+7XuNMB90AfoyiVnlbn75iZpsar9oIcX7vS72RETe0Ksh1gOa4PcAFzk/xVwwEXDK/GVGI5wVnf
0md7Fb0MZUudxmJXIZgScndCJJClxnbKjgYNANVS/4q4jwaQAeIqGwkWnQDIqtgYa2yxE3PT9Osf
vKDCmGIaLV2ZqA082IWlRjdJn1MQHfPTSNDoCfWBMo4iyr0BvO2mnX8a6FgpVE6q46vd2/CIWbw8
0tNzufQWD4lXAoQ0RMd+rAU3pA+jDn1SmkZw5dq0ie0tvrZwNT2Pdo5ihEIW5aU365RDQZvjfkd4
KIoN5cEy8ugh7d5Co0cWhVMHfVALuooAfZxoli5t9DDyOq075j4puzptSjASkVk5rt/5Aal8FVP9
kG9P4cg08T/l8bp2G2ec4zyTgzTDZDya1mRtAPapBKfPYIzyPSVYG5kXWMs3vyDffRKwEB5mTqcx
QGRW6oaF8/M9JSd8VHszNy+W5BBNHBDwAqTyCz7WIq/LAddMtm5q4TWVhXitj1n1O6ZLpVakPHpS
nE3rlrw1EBMHIKoBUuQC8SFuMWndjBfkRS2DJbaGajqdZwN/YnHYd85//genl0g5SEW/xxfYWHDs
2zhvbT+zPf/1YmtZRo+h2FTkfnFmtlLWEfRaT4Dja0OP5u4fohJcLxehyRTEsy17/CzLslVwPkya
kcO6/9lWDr17wOAfN8vabBjQRwpx8/nGUegBvGv1DSpdzU3TWj6pOvl2O6PCB60HHrSsGvwbvxJ+
J/jof/vApzDGZtp+wgAe+gqFeKZHna1sjEmvf0aIDE3QmCfd6WGgLnvclIGLTYiONSGGxfWqdkX5
zgJ/ZghKnYzbbKoYPYqP+G47lQWuH/OdMyTkCh4HvLkHObJpLLywEzHolx9eTir8ZVCqI246Q6UO
b6nx4yKJdEimxXHpGb1Ezdrn5FuSGlZ1V+lB4kJyz9gfwFEooxfR9LSU8+2HQ6bFemrAZtzSP4rr
F+mXxFrvWdd+uYTbITXzGm5uWyCimRXrZIwycClW3hXe+oDLNlgJ/5gwhSfgKficA0hXQVOFDg+K
bBnNPIZrsG7NKVh/jWK5w4MhJgCLYihEmztQ5X/g+EGbhmrb7vhcdFtbrxLyziEUjxfGPMjqBBFo
ln8FsHorn80EvMuHVde1AtA6g6fp4KFgsb3XX/Lyh5qJE9294rg7GfRJpAuB7hR8THVCaEwjCk2y
vnkWEJrqI97AwcslHp1PcxLSeNylsLYOcKQ+gxrOHT4r8N9nIXvvHwGnR+LwfVglrgA9mQl9p2U5
V2XJW44CsNmYbAtWjKdT8KRaImWgkJwetwQhgOMEv6jO0+b07oAjmbzKJiYQtdtqF8rQ3Ey85rj+
O2bb4N/OOOx2whwvdNgEVEsSDLdqpEJwq4h3ihJ99jZof0noOBLG8w1QGqv7uT/u64kbZmq72o/Q
KeRbVG18UyoZjhabn3Wrzy3CdjGnBu8w1AXcKpQCiGFMLRIfz1plLNH/uD1FsX0zeXvLD3S86o2q
PEoqWyxkWEuZsKJsh+nI80Jgh++YSPvCcCnqvClEJiUU/+41EGgD8Cd5mHyo6e+EvT8Jiv+l+rBw
G6BwKVB8zoG6Yc2CbcLq9AqCHiKpOsCsJCaWC5EB0x+isWC4Mez8K1bEo5XMRlpBFoz+Y+3Ko3rK
WGGTpKQBTLS7+dCvOnmdBjFPfsXBZCxVkZgFQmot7ww4kU4XlXBrg2/v5C4BTSlO+9TSc7OjpNOF
iHS+9CeYRiGsDr0ZKcmH86HdBAP3jv+0CdjWOvjtWHbAFS7iQMwf7TaQVfB15yfI4G/Q45fo9QW6
WD14zapiXGbtF2MnmLB7QDvpSsrpbDJR1Jc+ZpMeVm4Bsddi35LtGwvcM6CD9pQY9NNeUJ+uf8Al
eMnxBOEPNQ95M9VTc0H7k/1Xf6Tc+CZa7dY0U0wczo+BINNt+B30PRD2snIU4M273a+HRf1XYSwn
M/9r5tEVdFEogPm2VRovySF1nVuZ7LSJKJQTD2CIjugKfLTpJrn3I/lMRbVZsPkoesLUsEFW6CDJ
GN0h+JB6Qc2inqk4x03TKZV3/npL85vVhHi2/0/sw7/Am12PGgP6I01rW5GXZjIMzO7PnIQLKp0e
ZlrelgDYxx1ElqCLXYrIQb8o5cvEmV2+y+DQ7PV1Raxbg6m0LKzBPxL22SLLceCCB1NOLWLZWc44
66o8MRzg24lS5uibtGs3MfOKXSZqaB9UuzrX7tETwhywaIh07hV7TnRrq4fjgZ7oHJ3Z7d65rwBQ
9aPd49BD0SWaRJMmOIJ0BXrQb3wZRN6/fuvMVsGicu4wCn/L6FSvO3OkD5/62aPbHTEBkcckHk9k
g57VCwnBA4jZUx3JZ/7fiaDaMJEkhfWafdxzgpIt5WWfcMzMjYYhaA5Bh5k7SnWZDAOnLmUX+ZVf
aNQfEix3NP47EpnV55wq6KAEdK/U0rZiVKkl+64Y4TghHOKz5GlFnuQu8nxwrtzPqDkqP1B5hECY
YHVDKE4x3K9yKTb26Hy0DjapKkuZmE67PvewuuBwUN3s+Y39GIkW338SXIjUeUZWpL5Cd+qrxuzL
1oLuikZwJejVuKzd36fctyLBX+B5jM1fKYKxaVFhWCaZrmVBLV7BBz9kLcE2yP5hppfvUAKhBvsJ
eTf4JwdiyxN9QAPoDeHpvoi1VwuICRdBUOiRBpJnwQ1mhruBzlVkU7bNoTjqF3r2iEieTe4AHogh
HqbsyFpERZHfFjdUwBzZ4rG0qKUhBpSq2NeclcVL5maprLy/tfsNOOpeI0zYdRc/ER7Fp5G227Yc
7PwDOLrkqwgVtfrQMm4bOoQMGVxnfI3F9d0yJ6w/qo5KSGxoFvqAW0d9Uz3GykRvtsZ0IFVcKUMH
iFpSZb4RnNzm1PRS3wol6nmMjb3zc1Z+l9d8NA1p2I+k8NG/wTjNRNtbuBXqGs+Uz1u2YA+ent3R
slxd7pm4rZM1z/9mFFrsvOy2VU5HFhklhjTRXBX8esQ9USFoOLbUeFo5+GCVIun+uE1wo/dpLxAV
4y0UOk2M5YqMCmZr6ETmz8aZ4/Sqvodok7jo+KkJu4rl2NwMNzNbZwzNaE2MwT3EOp44i5UKF7di
uJw6bImviA9KJTUW0QxjsZxH57RHROnfD4pQYdSCL6JMMaXSzOoYxhbsUEGlGzr//65aySosU0ut
b1DjCmS8//ErKh8ob6pIIrL4DmNFAA4D+Bd29eHjda3TmADnpCeeSyFQDEk2rwxzeicFuCrLjh+m
qcPGOd8kwGhcKW7i7jB0Ej1G0fP2OIj87cfWjX6MeI9kzUuXQQkM+JA8FMJtx02SiINavhpgHmNz
Zsk5wscHlqeeV/dIi2Zd6cWUVE1gjFfDTG0Qbdn/eWEzoBeoC0P3XmvcJYFp5TRkPmlpEOO+dkWL
Quk/TwcFWLflt2fAwWgXUP+wBsvu5r9Ve4wxdpu1DkhlQt8CbbElh9/XTmUAcJCwiqM2vNo0XLSx
JHcLQtoI0caiH74IkmaNY7RnRUp3J2Xih8r57oGAfT+AMt3hRIWLpE7yefGxVqeODvZfCEeFqVO3
LtfZEihvovIQWz3gnbYNaoE3CpisIZNMK6osXrYpOqD7pGemllnak+FdGK65osYLDU6gaP8d8Mcn
HEtmCyT0uw21pAf9k6LrB0kF08vZBydMiHkhzxQGZY4JmstKszivrs0pqqEIXGQoBjdCIgVN3dMA
eoSZFvbJsfxA2OtIFkCS+caug+gD96hS4i/VKJJ5Yj/W2he7OADQhCscBaNBaJu89O0fgNyRa6g0
m7iv9LVtW9gvCLg/GjqIkgqNJHcKrN2SLf/Mb53utp9uYqNBH6T9/N6g8a1iBTlY7/B2FZ6UZbnO
M0WbYSPhhY+VkaqlqIiA7s3BUyIg9/LuIOlghzw8rVdDWGzSMcNRGMMDXtnyVtIOyhfaNN0hOCRl
h0082HLVX4kLOT/zZvUKmvA9HOhS3yFew19FogeeFxnvANF7hvaCSPigttAXXdcswVJLOr+VqJBX
+YWPT22aUkxTq68Lz0r2MBTDfUYPeJhsaJE2tguLJcdAPahk/rOb+Gd5WyCwVnG/TQDFrx2/4NwU
A1XxLe9+Yn+MEYsi3rZ8SHGo558CHQ8bZuI09fImsBQyc0rA0Oz0WhlyzLKq5w3WBFa30V37tQmH
wZzHro0FWnMeSE7HmCMOsF4bQ95TAGfs84wCq35GvvDZuoSHB5r8LAMvJ2s6+IpndMxFizRmdZHN
5y5wC+Sfbxy9cOn3Ax4ZnnFFOaWqxBKpGAQ1RBJgyAkrhRg8xkYEKcW3EQtDmxrcNvPB0dRXZiwN
wquJufEzNZw52pOKXIriGEYyPRBNc+zz23co5Y8X76Uf+1nDHlgZHxuB6nm3I49yF9oj/h9OeJxM
Zryomg07KGDwIpf4aANrUURrsZrwvm3aBtsKyI8V8o2XE4fkuHW8crku2iSWQ/Or3bA1e2aAqZqF
CFmfV1RzvtU7Xdt5LbLstOhqC9BPPkmQZ0UOC2rfXHgTVrsIBdgvZWuzR+ppZcUd+03q4yVu4B4f
A1wtgKZRJ56rETq47nRXH6eZVhvZ4nHpRoWorMqAcZYBM1xR9EMPsIOjA1GF1g/QIhjDTgXYCWK1
Rn4r91mU69osGB79tjJdG1uzCUmIOea4b21OfdXvPr1rnrFOQfoIQUZpNDHYGXUg/kg6+6I80EAP
XNbiOOTqRKoMv8n9DNxlk/nSeLkfTjcTpFMe4n3onOfeEDn5tA5CrMC0FlFSSlX5lAwmNSovMXCD
Q4fCcvRz2uOMnfJwujR525/vK/MRhhVgqSzc4Mz4K6jjLFDU8mTZHHtgN+pGwd00ntKJrj+d4q2O
8fQx3ePzhYgQ9zkTMFlekeR9/VXXFy1Jh2yzMfS9zWrwvKRAgKtHIgnfyBaPOHsY6bkt3EHPf+qN
frJpb3VNQcj8JREwH7YPvpNBjOP4XmPurIkc/nW60ygnKWF8kSA9o2GviHwfNZgTKvhoqgVti4Zk
AgSlhSrUg00ttiF/7iU6f5+PBFlugt3PrissEWCVpG0dH1cCE10J1OxV/fitKfBtPbt3PzKPYOvn
6FjkJ7UYeMNih/DIHJsND7lkbr4XuKMKEN0fTJH5MUjYeoDRxSflYtXmsYrVH36WPNIq8eF23dxw
FtVLS1F23+/UWBjk2i6bSECGJMZXkHvp6LqkRCx8j4T3HLt5sesc1hK2h5vPBaxdZXvc4KyHeuDB
CjUM3YGxZB8GfqNykmvnmxq8fhwSpkj23+CtA31IdOGdJSz2LeQDvhiuBvm1qH0NZRmrLl1K1S85
TP9sWg+ac0Y5t3eniGVPt2hFhB2CkZP/6f08AHbfvGx69H2paNchcsuNcQWe6QDYif3803BA8f/1
P/ofBpNcoRArQTH1yHCYo2Qo74T28yMcsJlpQOKewQEzcE1EyQVv2jFYgaprtU6/3w2/QQGgVW0p
ddQ84/5nJcwPVYhd3CHLEykGTRPpSr20oqy9bkX7N2twZiYX2kZOSeYpxzjSuBE8Zuk/dxfHlJiQ
jzXN/WvN9Q/Qk/TCrmDM29jzpLB/aUblsrwWNqD5uDTfLSDkkW9nrN+9Ui2HOVSjsRyysNxQiL8T
LnZiQxKMdPAQhvc/bQ+HrcoyF9d2nyMGkWEKH76bk/h8dioKEz1SWaLdsce8qr64g7eGEgdn6OAI
rvItLi9THZ+LOXdOf/c7I/C4e6bkEKIvVy6DTflpypPQ/qBY8B4Q2OCt3l2g4nA4s+VeA+hhv5Yt
mjURhedgJE5og0Hc0MSWYFS6Evwtzx8cbelSwRJF71QJlbOIEFuzqVUVvDcl8iQXj3ghG1IPn6T7
g4emPod0QG2jb+uTb/9mVMYrpxN+unPtFrcz6tiXJVkxD/azSDx3itspp31/hOJ5gtnLy4VTWRLc
Tk3IyC3ti9GW2XKjye081THp6NDlIwUov6UmutlV/2XLcc+hAz1CVRR/nb2kWS62QWFvCprRU0ed
0Kh4kgz55KGDgI3vgB8bzoyTlqHvh8mALLVtbAkSi2lwJiUafCmh11VlXQVPGS33h5flkN7aNQSu
wpiwaTXgVrwqGJycmjzPdZzDKLzvVNx25pyq9Aq51enTlHAG0jw9Z1xInbgyNzrhMIjIS2f6jJ/v
NNaMJtXhIoTz0tXG5OBKs3jtbpMrsRNPY6lmHaFHd8PrfwyFXctyF0auiCZFAQLKUd20tsVR1Qcq
VmrI5yBHuKIWVttiBqhH279i5n8oAxxtWd1s6hQlMZWhIaQgNwOzMT8Lw744BPS62PBmKmVbSe/j
ddRQ6eyLoTkxkPpDkhS6/M/fafavvm5cO1tYeWzpp15GtZbKBWyA7p73vh5I46L9anOF00ISMtc0
nElWpqnsWvE48pGeaJ4A+dxZ00SVfatAmoh/67Y9J2Y0Lz1nxCm655VQcQKIYQrioRG9joNF4wro
jXxXL3/CKu2FemxG+hYUmJgbYkuF+7brVuf2aw6XyhB598uerYxWOUDBJBCCaVbAqsvsJ5nff1KN
k/Ct9UaC05QaC3PNNKVlOXpP5sXXfSADJMAO9JXuaXOZEW9rM57M39xf628y7BsfDeYHrRu2sx1d
hz4x10w+7dgF4BV+BZSwHbO8a0M0pywO5H4Ghg76/v+wixcGf59D0j4snBnYgDFtT0CfpwN2BJx9
TbWqQjmnLEWaQ3o/lGpaKGAeyhbOZcnyqrNGxdt1jTEYd6nB0HR78DfXOP8AMtCkCtsueFumuxXU
tD5s2E5BfzfSW+zjoAPRLt2J/k1NqMtoo2CGxlXQOKB6jy5Grhff1R2+DAT4cviikZYj0GcpUhrx
+Bb6GD7+uYC96SnhLaThXNs+/x2ZHjogG4V7WBsVKNuPz5rsksjXR4sBKD8Ksi5rzyNTT+ysk/E5
vRm1ORQgA18PQsZ8x/n0t5HtG4gg/O6Q5rYacgoxlFoam1CoDsAI6xgJJUQ5SQ8mVaDVvMqHr8te
VOsgqo8xDxvQ0zDatxn1hazhmUS9sId8cAoUjwk/mnsk6yfasnrjeDXtj8uqkzPPJdMOeOuG3DLF
JTmbmmM6BSEI3AYzXxA8eBB5Flo8xJdFc3SjYA78BRWtRSDAzJZdkKsnzauuc8qklZljSECHpfxW
79l1RiQVTipuI5NuSw/K3LAoWfv1EozPab3341XlzCDtEuQMtn7u+/bhemHvYfP4rABeM9rPTTpR
SoDST9nRTupKRzXGb0ZJrqgHUTlL4YwN7qCt0f1HJLCm5HMMo2RuPXJkT/5skwYm21yARP5HymAk
AXLrXLyA7Khshh6ZUbk41n0sAH8gWCSfHx4LgCJsTjnN/EXefP7ariO1gSCBgv2OsypWjeTNvZkI
pX/ZyC1NdHxbie6qlOkd04uYD8dx847C/f0LuIilOr5agVv39vEaOlwmyeCveaupQH6b8P9qFRyW
wOmG9bCuKyfFyCP2+Z0JESKMxhlNh3AjgY8/km7/44giSCHJlsW27gJbaTnZvQphqIKuCTLD663e
za25sCuc6ODOzfZA4maKWpG09+5sWqBmFUjEPczhctDDJFJWITE/6tvBX9siGtUU+Hez658bgC4f
J3IjpgeU9x3XlTe4ACOl8wWg460d/xazg3nLvtWY9aUwzB1gSZnssMB+e1b4IlROyyviGr85scKy
hy8ZU48/+aYzI7l1U/wOak57TwcnF6OiRlfmbENl4G9BvnU4J+YiZVKMD7UdLg5LxLhV2avMO+sz
ZcKV2iCABleDDYhdxsx5T9ks/LPHCcDNWsQB0YLG1tq7rbdFsVXzUFWJjL0edtFQ9XAEzvesd7KA
Bv5Tj67DLxs/6EEghJErlF815+uumN91XJjSyIA5BD4ckqzx/ng+A8P0pAhRSybJNkKsuKRMKFjR
xJbQvdqIVl+OKtMq1b1uEzh9tZ++vgEnzyO/Dh2rqHSAoXw+lkdMS8UODj0DKS0JgGgtQyg9UCS/
QKqVpmBybwYOr61OroVGmvmg4zvGm4wIY+ywj4fIHKxD2DM37UwihPS7yMuc7X5UfJtjH/6qPd+8
Wdhe4HtPlwUwVAXnGnen0ro5CnDbgSieaJaHsf/2DKcW6spmH0Rd5KtVlfVF7LdVYi3p2vz+feVh
MhQvTh3XDfJ31ZS13rLJecTJprKq9SRcuJM5VXvusfYYVOTsJnwYPNFD7NyUIVaw8Qn/e+O/eH1o
66q4yNm9XAecdx/9RtMIyOptE2rimITUWK6ABMO4Mks1MKreJ7dDChVcyxm/x8XbE4/vbd41fB5d
b7KstcufpAtbeb30Ayc4NSGqSwQ51KfX2/Sef+cMrvH0+gygq2mzSEiY7eshytGV18/gXTIiPVjw
BBU6cIUfDJ4ooGhfFHhKMRpDrivfASe/kuXaPwuBWobLndf2mA/Du2uYtkcW6d4u1N6+9u0V93Wi
9camBqNbGJ2ZBeUqrZ1FoI6B4UXRqjyyisNfcvb1O0Zx/9h3NfXPTl9OTzCBJ/AaHcrmPJ+kBBH8
D1mK+XodUNYCsu6kN7UDnEo3nHlhIdzp8IxoRvI+5fnZNxrj/O20QDphnJjNpNbtojEBA6JKioSx
oL8IXI4k8PRm7ixDGqExJ9i8js9Axe6QsOuNsxx2BaEmWPF060q/J/WSAJzlrsYrfdepAFV/n6K+
nNkyvNU4V6a13TWNzGA3I1oUj0wgUQdQE0c+qp+iJSxea87laaw/rUhHfPN7zLApJ60HoPr6MSl3
dM03OfJosLFUpR0XYLaIVsHMGLx7s3SqzKsOii0M94NFwsGHjIiB2jvzYkN5HdnRAbUI8PJ2LXkk
OrP+mNoLinKD/NF36t2zui8IDaWw9KVR/ycaVLgZRcM6ofTQh5OkA6YC6Aqg2rP8TBqcxKkDPirE
A1m5oDsxqgm5qn3IrRH2N2iQgy4pn65r+2S3GPnYAshji1EEITmNzqnIsaIqJux+LVmKnYurZqdC
3LJGB4TnjFnwegZmqb3qw2TT+rULpQ+TIQb5KWqNSpbJ0/E04Dj97x5yc4mK6xSuqvJCE2thHPOY
HQdXGY/GRn+f++/MxZKEVNpBImbC8Oew/yUDs0SgCMoNbxY2QsH5QRgf53rdQMUckLRkxQVvP6l7
pNPUAa8cb3hSuuNaEACdauDqZCC+uDBqDMbsjmlFtcH1/7+jXaauqDBUVu/H2ydGg4ECuIXpD13v
vIQSZ1s5V4sAluspuMDsQHxDp/bgbNZWOE5y8XOOw83DAQa5HzbrY3j+YUTGxzlvKCivwcLWf4cA
J0SLh3/wkjttA0eOLAEoeKIC+sqo5o6ILwQhDkUXEwx0Qs8/mjmUjhf+ZHzXHEDeoB7zcAi2qbLx
jpTiCdTApxz40j1q9X9lON50Tu6AxwPQpySR8tSD+wltGG+3iqQQKSlJ+DLhDfLX+RclmLJJqvSU
FMf9t/gRCcH2Z3LtqyNdMTX+n+blsllltwsUuQOPeSto9XNjvf6gIfde2rb9PGU9ABBXYyQi4WJ+
nstECJTTNrzfPRHkmvCxCYXfhD7X60DHnhn0UhYasAEZ0wMwys8kIo+TwZixBdfKieK77jqMyDb9
1+mn6eHf7Sko0btvQedGgFgGF8zQBrVFH0TlgQR7yWbcETTbcX7HxEY4chCXZ0/dg0sGSjONH8T9
klqclJ9D93kHd3+urizXC1GxA/NyO3fEiqomASA2tOMqnb4Xa5mGHUwNtiV2gJ56Exd3vMhMfdep
DBc3wiM3EK7OKksGuyfWeP06/OsUuz/LzXiUj+BwvFKASPpAUhZQPvkAY7eiIunPorHiB5aSvZKU
9iOjmESD7tfWVLT5ktzqwm5C+E3JyZiXp+U7cVqE/BsPmcdfEuW0YK2gpbdBAVyh4kZW/mhR9DOH
Rn7G4w06C4cTznipB5ZN1YVEGZVTYRGvEXuuMDVRy/7JJ9DFVUSXWBasUEzHn35DnUTOjlnF7h5Z
3yEhsm7ED+FQfRXWNVO/bFWmo2Qsqll2xAyHFnAXsWAWPHu7fkInWltTRXDNV/yBQ2uS8A9CXg4t
Hiz5Wmgcqy4puFcw5sLgkfLd0QwGo0O3I+hejnxIq+LmpJYhf7Fj5gyNDslnkJvLDfltuhFUA9qu
wbaP7aG+FmSqbSVX4qd7/17Dm50lFf6BroTfLQqMWjNPoHWCi3Px9BnsUGuMGGxdFENqwgnKMG6k
9/AL7wcdplgsy7DcX5X52sphjYH5TQ0mPeNcOFkYQEHX3sjKPE2iOzjOi93cbC4kQ+qsx2+vpTSi
DwZZa1nmbrUlR8sWVf8TMW86JfdGXCutnQCYXHZz0s8nRnn8ZtNrcpn2gqgbvjZ30ZpgZKAAqNar
OHmedisH0tz1bOYbDZ9EK5kH82KjbDymPHrWsNlNQwE9TYYlzKlKniMRlBwUXsBbyNZ+snIyR4sf
icaOI6z1slXFsj9RYOSeQMTRkzlHvcOfIYNAr6NY9TvU2khWwwQhfcupczOgDzTZKx6c6H+07hQb
+IjplOTXx9BtU67Dh7E7OV/SBgSb/qoGd3rW1C2e0OxYDVyEab7beICmcySDLZx9J0JIxB83GXq1
SALlUJbbXsPSXaUOFiDKM65V9zJGjkKsbBfr0dLy+4AhANm+08h2W/bEzhk04cSRLKKokKDwJPYq
qr92+WPCaLVq8zouxCeLf7gr2IS7BpBHDByAnFczFgi5qSRPKe4zOkNGASfXteBUZHeEm4Q4lYgx
jbiK4Nu0CRPSLsJSdXqwPYXyQevxfL3h1MvI1JTM5sODK9ueb1v7BOeKRRAx8VaCM2wbu47Qpkne
pqSR0GYZR/9KAYUbVQ5R9J+nXNHUyLWixXItzDTjvkerB3MKOZZS9NhPnzVbcmoaJJiltTKmfLqa
kTfW33WAhOvlgNr/YfIMsuobtgMY6+2AU3Drm3VIwDy+04s7Gq99pa2WxtOWAmuy2E1CME/ZVHk7
dB1FybEdhRB7XtS3GZzT9/kdT0MDACrY6/ckimhb7ajEp+7+UwpcLuMordKBUiyrp76HbY+R//D/
tTyjOZhi06N3/1jDjYKZVhxhHeFud/Jghe/VgP337lZhdjgHEDDBpRwDXlN5Hxv2j8+bC4b1HTL/
MkXi2FDQnpdU5nFrt+0gUNRNSWhdhLB07/e5sw13Rb/XGaciygW55TA1sZOb8BbXejKBC76ox0e2
olK0qR01snDSzJ5HfGQNNS+B0gZKy9xlwdUzD2+KVdf2xQ+rPO8xFabLa+vNM82qCE4Ld1S8fut8
Pi63R+Nxr0RzCMx2aUvIh+tTJWv9vfWKFV8yPTbUjlKdYb8goxX6UfjZm+ByaJlYA2oXql+RKW3D
9IXqJIC9OAf9ApTWRctL98+VSnN4dmaoL0/ysjGC9xLlNkiVdfx1wsfsCDdcH+bP8aSVFE5ilUdQ
EjdmmuFh7w2HGvmjQX36I2yW+TNDq84djClml4CJnRdu05F3YHWPUDJY4Yla7VLSebJdc2G5c3oj
ZXIxz7PS7vpO7BMO8RZSAU8T6R3BpRc6Q8YW2SH1VUjrQHIB+sjy8tBOGoZ6ekMmy+sjMuzeku2q
WuRt2D4ZNlD8HMKbAj8+6umVk8koG5y9wraBoo4+UBH/uzXO8y+2OauZSskPqtkqIvb3unH7KjY0
vUt4Z2YWvfIRSjtqZ/GbSc+/DqEq/AufIeurvj216vWqnb513wEl09OPmlBxkgN+QbvtnhjmcytZ
P/t21YNS2wiAS4AREqic125DxM7DlROl+TuFLhUsjMdiJkmIU58u+g4a6xIc/Jo8oz8+Uci+NGeh
pHPBtvBBbWN7ULaCulRUxwJu9+5lLIz3/wYwltPXBqEJ649+Sn3PFAI0r0g4FOTWigy6l2ptVpuL
ebmZrnS43lLlaCc+S1dXpVnEZ2ADKBrhA0MnqHAdm1QnZGc5/SCSx/hvuNmskVRLqr8JLippD11t
fjFCgMRgEfpJ4CYTwhL5n1xiysDbN7XkCE/QwHgtbGPeXVfP0Iyn60MKWS/ea16ky/6syQsYkJxD
PQfNct0oN6Oa4ifl3ZUliTMzFaqLqDv4tUhoWJgOI+LYGl2PX8xnjHQmSJV5Y4G5vryMolNqh9bX
nHjd6+czYwSG8JASyJXsVsgTs9CIVYDGhbds4Tp58E3Az0OMOi3usdabX6DZjXu/vQJqgyoN1Tlk
IH92akPVzLa86mVuTo2RCrhUl/MQrraYpvLax8jTg8/cyYyRjmXPQHpyFLYzoXn0RxeaRb9P6K0K
N6tCZQCqK9SozC74y/SjsNp0ZuzZ5WelpArxHDe3fbLXgXlyPxAu/PxVFSFtKvymQvmsIUkkXCfl
rgL08LkQXCyoKqqr8gAiKqtkGXR9SXPnP6Kj2UR56fOnkW9vSID7WCkkHy5TW4yULbGmqCf9IDAK
9UhoSh3x2MhPO3rCh/FAP6Eywn5G/v4zl3tttUo5AnLSfbS5QjOO597bB83hr2Q5wb8czpPNdko8
qcO/ojLXfkibBzIuzBwaTKSgumfSKH/tcByDbDu40CBGRNX9q0+YNn6XTVCs/IiNpnDFiIwehXCq
Y+YAP8a4ObsBF7t5VPGSxSQIHThPt0Lr5ExlhTJR7PwM2PH4qM9rLmEjGgtxDs9sD+RzfnM1ALZr
JhvTuxmqqOJJy7eAse70fnpharcwRPENwBLaxcZDnRsApNoB37MF4T1q1LFT2VbXMt0S+PK2AODw
Mpw0kLlPJqkMc9tA08cP55fwNUaY4d6me/yX9zWVpdq4YPzTWJ/tjCcZV3z5YHQ9eVMeYCVZoLIO
hS9OIj0b9SSJIu5mEwoNJgx6vpQ/ZLb8mt1DeIDS+lvC9zVZqaPHtThGmcufUtnCPKz/RS208QAt
4Qu7zIaEt+PESzcOzC6U8VBpTL5Vyj4Wln8TfH02bK0/pL3AAPkRcQwcsaW/4eLmgh4FeBwb9rGH
Fvbkj2rk8BWgmtHrhSggobUvh9bLHBVajvCJHf2kyi3ouAvpiZUGaER7F/wVyTK58FOHeC0ygLRg
+KrQnXiiLnEP2WCNRoZXBvkfQhAN594DVNer3a5nz3mtNdCgStFYe1vVZ0ZOOUkAVB67zpeSNXze
ff5m2J0Mrh1RjLg6GPauHlvhjXp4d/dcmR2bxptMJoDd4bbQg/9YRjn2ossnfpC1XsTmPLNbtTAx
4NsZ7b88+RiugBx9ex1x1n60C4HueTthIio8CZ7cSP8vcDi9O4GR4wPPhH6Qc+0T1G68J6u9tUYn
fpVl49ljQDwliQmFnfphzke18IU/JlG+NQWbrmw/BJU4slrHhDlEWOHtoV0q9B781iQK9btPGaww
wOqZ2Xw/pucfw7nNDhb9DhD12v+R02Y1PR8E1H3rc+4vO6ziGA6BB19Xhv9xFRzi0Yy6HdVHN0Mx
MFu/FzC7TkMwZtJWsmggtuzpSaOMx2gQRrQO8YGB1B05ix8C0gAZuSu+qZRj+LQ7EMh4fkuFMFhk
Dp3h/tzI9kBWk9WU8tK+cdLleaYc4g62Ei0s5iOfZA1gkPIsBX4JEx9egk23WcBiEpB0IGeACsUh
NRrW+IyDXsBxtFGQRnBIvjTDNl2Eukg3q4zpWqM8vjfdmY8WunHMVz/9jkpqxbudQ7eNshKiyBQ1
rKYdL9gbqBLacVmTPpjHtMvUVLHRynNQpDiURgNp6P/8VtlHNsD9NfCjWximbSU2tpXT42w4wYaf
I8iUIJ8VJIZS/3pRwCgyhxDf+n+OxMycWmN+CfiNub8k3Cb72P+AbeP2zIfk+4qs7GZrb4Uolv6e
/0Nk62+JoAvlAybp73Y7II39UhSk2bXzzVans2pwzy6vAaFv3GpfbVkBm/Bxi1/oQK1dko6fuVmc
qXxFlUnQKlWTcZpaGPRE3/Ue1RYpu8i715coiLUJvODaddORoFTOnrBswgdW43BftctReFF57G+O
WkllvIWOi/XwHoITHWBfjAKr5+h4xfNBwEkWKpeAbxxvKHVhLujJXojCCC2LnnH0jnHJZh1VY4di
fEBu9mtbebEULuRuOh8ahzpkbF5QeSORk3eOLNIHWEZRknuTlSz1mcBFECl9jYBVHEQaSwl05n/3
HrXtyH2uY/LENByvZNMYB/v9e4HTbrFKIx1J+mvTmcv+AICF6g8Is/XCpIwxgnp/uHgdJlk6dAKf
MioUluimkxc6OOEGyyaxuuxrZn9tsQRtwjIYy1gI5xQ0FOVGCCcgmYel2HyW0CKWroTnXVxnkpaW
Hh/uNV1w3+V+BP/2D5fOVyW4l2M7y5/tBTYvBuImbttvQypE1py95J8gE4DMhzAhCn+VPmpAwsR8
77HLetH7vEBjS1vGkLSZbDcPV7DINZ/c2+eBrqkM1ni9MfZM/TyNtqgSuqXSljEZGuiZqxXWT7Il
4XHx0Drxrggit8BEcG2Nz/FeGs5vtC9DaC8bP7X2B48jc+Y2rXXOmJOWpc9JFelda2JrUxXJc98U
XgilQS00CErrkKnhEVFgYS3IJgnG+qd8Y2DfscjpoAHkvxW5vH8Udvyv8VmR3UfdeU+5zKEHQmuc
TLKbrmOphBh+Prh5+u/h1EgsMGhld6fGoNK38AgEyBglwjoJxhd/bUWbVYKWWLq2eRTVHBOgz7oC
geapIacDVY+5Pq94Y/TP2kGO6f9p5XKkxNjhsu/NHzRDjOthv2ftZOU+Z3I+HkX30lsj9OaTyoGs
dkX3L8aTX/QTv//s7lhBQlI2o04TkzghnH8LQa46KUVKg42CQBkpXJoA/p857GVLirm9oRG0xT3F
B7o2agVn0Bu6Yc3XqMwHKVbAiGELUyBmnyDVxz8OUNzl+tDct0MEvMwEzglJkwTb8BZIVn0hhx5b
K12mxtAc2XRQ/Baq/XnSTG4YXzyy67oOlks22SLC4HwWcs1gsZuVgcwmxZi6u22R4d8N2VVmnK0F
xvMN2oHNymmlpIKFrZkmJ3fzv54nzgzAzqXe+ZdZoJWp9A4LA9dWWH9KDH6A2Qx08pPGklDV8TD6
/u1pz+vbeY5Y/IGOlOzSjGo93XY3qKD6Cj6uzwE2iIC9KN8wpVKO5IPmkAXUUuNIWcmyj46W50jN
d8s58ZnS2cVI89WNukNJ3CP+nqtxB4Y6p3cs/ngzjB0TSQ6IIkjYchZsHrpGxcEIcGKOrjCBVCf1
HU4GH8AQJD36WoEDBhj68yjfa+GMx/wEItLJU/5/7ro8Bkb0rnQfvZieIwAhzBMaKStygNZPr2Jf
SHYLmpQpE+shQahu4tcgMu6gMaslMRxIrqBFzC92+KerVP17Q/7yAIFoSqhzKy+6vV/CHluCaNxW
NKBC+jZshtNFar/sRrjHWkH+prO7BOVCPL9Gl8cffGUYTcuJOqN6OWX50HIkUp2ic5+7SsKhC7pe
UJfXP1HXXkx6smkpF7AhVgTe1v5kG8SG8NBZruu1f+SoEOyMW4uZRcGZzPuVPx6SrtiRZTz3dVoa
F1ed+C+xFoT2iW2GvuTYiCJsNnQQmDOWSqdGP8+fMfb/YoyiiShijdN2nXtWjytXyPeLofJyCNow
763KM3awPAntE4hxErEXJTbcRczVUAsO+KSVSUhVGd7Anv/Ej40/+AuZUl7eT4bERkxf57BYBGdr
/8YD/Jtms0L3gt2Zd2c9pj66JrGgYm8dvgpq0xRoviNDSHDwJ5NdbyuyPpl1Hc+A9OF5uacXUUxi
qkD+zgm2O8G8omAtSbl+oWqsp8+8lHkv7BHX058DpCc93b335Xs7b6V0W1C2h1dvpaQpPiUBKZq2
rZ+HUXXGC3u2LOba5MC5nuR2nyBgQdx+HZL+wWOSbDX+jLfUvCSIAMTPHrRJ8XyyclSz1MQ5AEsG
5kF2LpH1Twl0MKQyIS6vkFaUrVuLAUNk+8Tvt2EpllqI9VMhYlDl81hVL3yjRSsHVTotQ5+uyJEY
wEPQm0t9MJdJzf0SlI6YOOMxE6GQABpFZdw9mYSf/2AHXp6gQbEVwzyeD5nhz5tMcRH72MOiGmgY
shV/Za0tXhwYTQPKaOXt4NnJVqY+e8NJh90OKvy+cOP7ZkWfHaDirV19TVVvps4MLSVTQPmV/IH+
VRqSVBfeRvByv4ef9Ib1qFGuoWlxvczNt0lg7t0UwYpMa67DZYXkPt9rDxEf51Fw+tVG/jawEF7c
jJIpe7yJpcyLQa/RuuKYJW2UYhV5QlRvYYd4LJvtij+q6BukTwA8a4GPSXbsljk2g0AB1pb0Pgiz
wrEhvqXakqHELzA8JfVq8uh2bfENMQLxccYH87ZDbU1MVFhaEzRMJiQxVBg5F7Nz9GhLsBaV+LK9
V866f2PIQJKhFyUHuFROroz+6xzPRmI8lHqymJYrhqCdBbhNNphVTDBZl/geESFKU44frZ/ED35z
lGkMbjYnvF8L3Y/wLQ4b/8mKaDbrtw4MV+zfUCW70HtI0tNB0tFSdPagKLCKEGVq1PynTdyLqM7d
R+0Ik9dZwo+5gYZSDVIGNNUC4XNNavqAw6hav01OLW7qhXMdjxkM08+fuW526N4Qn3sMESGNm5un
GCvIBo/TiABCYvo2x1IKnVeSJVs1iOBXiXynLulp4S8S0Vcm7liQoJ6pH2I9iJQRHJx8UPR3OLSq
gAwTjT3EPhcz/nCok6G4i8zErEs17qXtL3/4EueKJqQOOSds2qbtbl6fLNiwbkEuwdGh81/xMDSf
nunkdlvXuPHHSZkd5YGSEvkGVpveMrfNYKPFQqG2Qy+tspiZXzmfABzc+1rGlccW39yRwTb0B+FN
R4yUOjAKXgI3vsnw329P/Euc5CtxYr4Fc9SM4P9vSSpX725g0a9k5Ir4/TPEWCD6ZICLRMoFTo5e
RdVxU8vf0IYDz+l1w0LNnAxAUEphWnqP+NxLo+NDosakUkSPH6RetqEhTfKVyJiP2NY1p57dSemN
r3rLGZenWPFKF9gpWXoQN/47PeBeRIA2R+S61dTim7md1L5c+xTuQ1y18JBRY+mu59KrE+eWGdAH
ojzDkkXUO4y0t+UYp9hKCGgjm8lrDiEs3N56Bg9G33va78Om/o3DLjQIQsNWbZ2z2Lx3eZaznXwA
UYaccbNybjCyfP+/nWkcYIrZIEg8Z7z7P34gz9H0n3WLPQ1MfJMWxK1x/Z54sOoS2u6ozQwHYlCM
uZehaxSkoOzy8Z3JbZROegFK5hMM1JnRJ5eTWuKysXHr62fNfL618Fd8rpnJCUs9xhYZALmi1eeu
wF0hxYmx+vTVtJcJ+se8TLAwUtgkWTCyUcIUDbznh2wL2XxKO7c/GQbUJtzhLaR0cCPOKEoUKrsO
twsOzEU4MRBFVzougie2hR7D8Tc7+lUDozACx8C0CwW6IXLi++7BJRGkJDSdlJ+Mpil4CI30mRB3
ADGsryq1DH5oO6ygn9/BCQGLAtrXhBf5bOXl9hH5eO4PoEaN6duhH11Sxrb96o7E4YA064rgckpE
QK3//6mQj//yfCa3jwksLgzJ6UVJBCDA2lLgk3c0korApUCTxsWSHruuTf4AxPqNycCEHvlfpKcl
zPnzP2gnuZm+kLRbXC2YrjCKpKb4Ckf5XDITn9zG3+xGW9Ly60gM+U3W5UJgRrxuXdg1eZvxID7u
37p2Dwfx7WajmsLi5PAjUWCs1hMWfKtlmYaAaaPTQ+o2Uru2wZeUu/uEbwqplMcmpGD9uzt9+BPo
EI6nypt/0ZRZonx+bIMNc4K7GFfNDrxqvBxVeWaHkrtN56lCkF1+FCCGymta7d6EP9z28VYOseIL
mJjeb0Ej7fN1M/+1z0ITzk7omII5tX1CbAgWQD/y2eUAz52HbMUTYi1h9ttr+wvj5AWUqjzeuKr5
kUy11sqiD/mhKWCjs60eaiSf48wMuFE9pXyuqHTrpJB9NihXiKvg5989scAgqz7UWwAOAVZ97Q+g
jSkDRsPuAVMPf728s6YAhnek1dqfSS0B2bx+Crkr0B2FeU1ZAriLFpwb+HaEFhlGAXM/gKV7FAEh
CSOIMVFCRSnj5AiABr91hk+rHZG2K/J8sYkOwYcdKwiY8zkOUnFv+YKMGl1yxk01hFHyCzonSq9h
EjjSXfFHB2keQV29uJ3A2Ah16vDcjHsk3XdmhqQy2m8ifhWOQ6OUf4SAIjNqzpN0ChM2blqPy5PQ
pUy3lwWuZpJymP526ABxrZRJXtLd6tbIsQNgqsN8l/bBJXG+nIjZIk+fdKkv2MvHIoiwk1igvjpT
CcQyK/OiVKyCMduQmK1G/WTlOPYmo/ybxxaDkJjMIXJViyKpvfbZpRbjFZ2bQwpoq7i5/FJ3NOLd
rTXhVwobU5LoeE6AqsQfwBu3slvEEude6gPwGBPTxrMjk+e39cQkkAz/xtwUOt754gXKGGjSQHSH
rkWcdqfb1g822LzoPaZRyq2gpnIrZqfBAbfJ0qWbX7BD+35QthzTzIYfwePguMsEv45dISDB2ORY
/vxyMolgjinq0zaFEi0Bp2wIsDKvxzg9EiPJfOCcn9MY9Xa6AtKJOjvascRHZc6X2t5alGo1gSC0
eDaEktYcVgt1j1GAPLeUVasfRAw4L4AaJu9MPE5tiDhz9rcVYaatLiyP0hEaLJAgRVLg6fjZACzd
ITISpVlSumiZOzpQ6ApD9F/LCDytpA30+7Ml6XBgIkqVBihQJrEH9RymKqhX7v/pHSh5wPSSIHar
OPX+tggA8un8f4S+HgHRKH3UYmWdhCQ3OI8i6bOK0Cpj2p3m+Yw5wRgDf50AhXeXoqY37UEHuIQ8
KZs2hTxOc4RaF410Al7B/DtaMDiu+2OmlZWxeK15NBjCvRCqgzgZ5eVa9J91qxQCL99xhXSG8gRX
fdnQqeEoIgHAEC6RFr7fEMhMQgF5KV1JnZx9Km54v+f9BFtD8m89NdV8Vg5c4dJpCa4FitggeKxf
hw3PopJWtauPQEcJq9QvPghhspm4iy3I4Pp9PKrfdq0mZ4Qe+tmabEqd8KVcEcl91goqfeYKrim4
pFca4PMWMKPGD4nonY9SCn4Ytk6HyRORB5+/oUx93xd1w62XWYemfAMYaZekB30uDG0M4+fq2J9E
O5NxZ+JHDL4bYPj1pMd7MPsKMCTAxNz/r4iYL0U/aJGMIkDSq0KKNhiIyk9msuKhJPl+IsGbyjtc
5ntpMiXZ+KYRYIO1s01FUP1tnaXX0WE6NOoowyAIno7Cjd5S5Z8Eq/z4mSrspfXJA6ItRzB2QkLP
TM/KMnddb3eM3RMmFaEOfdBDbRny87wLCLkFs+sQ8G0qsiSH8nUrmVRCoVm8uPUBd+bsCno6zvRa
oVBaUB0i11BF9jqf2cLtlfFCeLrXhXQneEwA0NScbUnkzeqaNIblN2Pl/mpPjvlD254MxVyYDxyj
6MIL7dobQ8iZ/kppBQyOZviLDKrwfFNh7PxdqA3D4Jiy/7EfvJNGTOpq8ZLdIWx6subAlApoJriZ
pVWTuBIh7WCrRQXyvh/hAYI0ae7D/e6vFujJXgo7Y7DDhf19MKj4bZhsZkfZO0O4RR157OsEcR0w
zXPr32+VdJi1u2o/KT5TkLy01zJjJX6uSbjehQXrpT4XrLfJh4WUECo+7qkZVfQLgKpNKPBt6dbl
0LduQiLwwvLIvB4UgF8blvAuvRM8SXjX/DHxhAggkL+fWZUpEajy4y6kebuLd6G7B8ijciyT2KpT
QE/FUCloacytLrf0RCBYkNlBhUpuv1Wle1YduRBTRYYuChvKKIe6elDRelomP0uJdQuha5Ifibk1
79G7L0SCub3Zf6eIOp+2CfXEnM5tk21e2n1y2WAdC+EwVhgJl2Jey85GBmVlXymfGlP6KRm9gR55
d9gnL6S/s6LN9OWvyDCOrlRbH+vPRTsCaufxB1YDFom6vZ00+Brtb6rXqMay8tZu3Uk4JzeNiseU
dq50OodK5LUe7g9AXCz8yXCxn/ts1ydqEgDU31hG/Qkpbwh4g5UVaxVVjWADRxWZ9yr99drpucXd
8LgimrJAZDJDdCtmYkl78PMwLRjYr2dO2+Gcfm+4bBPvpe92xmOos3yck6zz9S9HYPK1etoLTCnQ
2zPEj940JyGuRHt/Qd8K3Ch5NmFRrL24qDTrYq7i58gVzhmfouiTiKvke9E7mggqXuRV/vuOerMJ
zwod6YnhnAFcMIFC3qfxQcjtKXHZJkzVBgQO25i2g9RYNc02qoPhf3RpoGL6dQGYA88gXDhkGrAC
swos2qIIU75vd/3lvvfSU0GzYluYTEYwA8A444Uhs6V30qjiBrRq3U4xPELdw+5lGcCJ9wqK+0F4
XBUNxDPtKHSCb32BiM0UzT9bqEAczCuzG0rIa7aiQz1X7wAatUHJSwgiSMc91OrmByZZx+Iu3o5W
XQlZVYpxYd0s1vQOZOglTR0RC+QTMHRqtbaiPUlGJ5IrM3SysXbgEpxj9PJjCJi8VRI//otk86pv
nkpTM1lrkenkkEnrMlj3wc6F2QD2T9arzyfnzlZrNvx6KwmSuBKa1cygmNA6CKyFyGpPWzh4Kyi3
lkEUtMh3hPbosRUFjZb2wHooKe+Pq4QyA3PvdfNhAvHt32Xm0R29fQP8mecENqc3eQblhQpboqrX
nrKkmNv0I/yX+MsHi9OysuQwtzEH/cCbtwLOKnBog6H/LA4nyOWlYhckBafFUPp+KcnOE8KaCL3F
7Smkg3FAYkK7aQttdYEIm1ttythL2EuqvP7L3e15AVWUaEHdu4azZ+n5O3YwY+Kg5D/mlDoFrwf0
0YhHXAtodOob/4A7UV9Q1nNozTqMxO1cIq3ILUz95HkS0J1KcL/v04zXpivqtzR3zkRN9uYy//au
o1qtd+Pc+PFUvAMLL1wSH0IQpHo1hFGVz4JX1ZkiWPJYkL93mKGGSlUbRTLs43io5KG4NhpFA2ZJ
yMnYhgFzYrLaBtc8fKI2VZfrm6t6DdsvxH+RQYwX2XyWQBYdbxNoRQCwWFWmT1DkHsNfzYIQ2Qyt
DwcB08B6scK0xdNNbkKy6v46T5WaDQNxkGaApv/jkXMUlkKOWTRTIiBlYkrZYf86KelbrQU9jHVK
8sQRVx4k+MWawxSuiS6sWkhZaOcYRZqNfkEf1SfnLvMU76njdQWhQJAGYjcNMkWsmEQdqjoxGxAc
aUyWJWimOe+egKvn9D75vFeiKvxeBnipDczglc3BXo4phV3YANouheePvXfrDcjiqlxgnUeX5GUb
GjnSzyvYK8jieORsE/RHf+JQSUXd90ZH1wRuwkPKhPwyYh+bnFPequPqtOa2dDTZdwfHURWMlJay
x1TDvq0JU3Ip/UV2pN2Y2TqPGh4Tul2lLDaHYT+u/EpsoquBYMK6cOv44TQdz55xCnwcI+g/GunG
HyTF2KNr7WGqLrF+5vw5d/mcdKmpu9HPPYXxmb4+HmCgeRTz2vtqTyQ/zbFxra1sAs9N79xzSuB5
9caun64l2qDkYPajrMi3eLjqK0dhrJ+fWQURIq+fR6ORA7o2Z93wCp6n7RwrGMC4hs7k2dCC1t0A
BMuY+0ATeUPxylLNT1fznffS8vFInm4hulVFLPPn4V951OGj1/IncX4022H0jPshr1nhoEG1Dup1
v6qgwVdqB7Z7rJIhppAy9S9iBlMzWd7bxfADwncEXzq1U8Qd3MMtsZltWoRGoKEj1lIf42heAUKb
FxkkAWQOR4LeONnhK6euUdPn3BLlsBPoLs2oThi5gco1xHBUviprrOxqXtMnHGZeMlnVfFr2fcXZ
ZL3rRN4cXXEnimAlVT8nj96tyKTqwKNkkqEiijmoTOLdYg/PbATwK8nV90x+JR6MHvbm89Ug32n5
x2hi3YuYhmDHcp8jGl/vVacTzvkYeiOn1nVtTUfYT6nVQqRggvdQjuXEYLSOcD9Z3XoqLEqrgfhj
191hLT9agZQ75Hc6+/MWpYR2pR/FSva2BGa0+bUYWWAIte7w3E9wLW3j5DsyE4L5oeui1/SRSNGv
85E7OjoBO0t6Xo8H50SuIE2WNFkWo2qFUSj6Md5XWAsomVojYIxtVBI6b1t9CfjaFt5KOhJqFllw
ZUDOwxwY0EtuwzL97kY/dYguqcaE+50+xnKz7XrJhusRp2ovABToiijqqTYIeJLypJydqr/AeU8h
/F/XorQ67LgBMF1WZIAIG2aJWaa8aC+GnLJxZk0AroK8AW6N6QyBtOPTjP6TFfO55HqXR7AQihQ8
Zq9CobuH0nh+sUmYbMuug+0MI5QaTsEGkKMLaNY6CxF99IfiiJUHVq/pfof0kYbZg5WiBWD9GQAS
FG9o3H122TQa0etscd/2rMUPjp6lHL5+d16KAK7WMlroM8OoUmuQaFKmF2/4ww6n5UrW+TBnHxWH
lvYggJ34M1Ojz+5/73H16hCYiGHNzDOWQMB+6VFqjOuHfw9DkHinj3e2TT8AKSQcWCfXrUF1ypIS
qr2iZV2UDZski297iKk56jaK3UhqRlT72gRPl6IVVnPDmapzjkF7OjKjLtAIqFZcV3MVaMCRmtfS
KzjC6ZrfYvcVM6EuBZBvQ2x8ZQ3ZU679cHrgOXVv6ZLGvW8L5BxtA8m0Q+47CCXzeok/K8EtEcsu
T6VnwxJnR7uAzGeQOt9KumfJG2jvOUS+44Hg0SPHieKXSJje6jKCPh9jS24KpMfDs7ylJpz4b656
ftr10yf2/L9ey5RfNk5s4kUlcRt/9yrkxsgtyFjcIlnpku9zgwAVqjELvKOo+Vi4nWk7/lCKaMBF
F68vpj6CH7Lbcs3nJwlK53DYu8U1Nac8YeH7DwErI5dGslNaum1GkK5QFjY6eD4TtJw0eh4jrzPb
Sho3KoMHJ0nXmVqhcOc33a3FYSrB6uV3g48OwptAaFP5mry9ZAv8QP8LfpKNjZfxbPvlMmhP4cYY
wAuEQ5uMHVykaj1PIq+Atp1UqgBVooh+MDMk24gGQ6UCKPoBctfKWiIRcoQpgIgQs+QM+vcDHYJq
BJQ6dy3+bD05AUWAUnf1l3evsh7F8WoaXxsVVqCZZhE4weY8qWxJuq2Io3vGFI/IqSoInjQ28uvj
pcEfAcGBe/k2xB+34/O3NHv19vA8qlIhUICLZqZe1x6UhaDj+uiEOmqjbIeR6xasgnzlRe1hodDr
4TIt9AQYBpt8+1xA9S4ZDIGovc5ndBLYKwog4mI+WrG3AgZPmnI2hRo5rzSWjrRkSEW4AyyIFgXM
44//8FxUvuJvzMl7UQLbsMAru1itkMIdm+xMn9RCS0VkfKomQ8BeEnzc4DOX1+cob784S2QLsn1p
wWekaaQBULUqCSmvB+fd5bYp93s+PFC7QvUheuHxeUHo6QY5avrlYPN1RQI+EbIg0OVMNftf9SFm
Tej5TQN7E0B85fBF1Yx2SibI01rxugatJza9LbfUZ/NdHV0PFLMoCrLvZjAZxfh8/rxflE3S92bl
CVkEyJSrtaupq1HTgBv5UBOuEhb5iJr9ilRSpP+16DWnuOcku1wlnhx2jJeX6ohkyGmGDhFySag9
FKMt2mLdMRwocLu7uE4muK+UBl2JaCAbNOCmbg5ueSJWejK1Ii+SNva0oTQMgd+xpksLELvjmPM4
Ja2BD03OpqIbLE42GFDOIjqPRV23Ue+bE7A12EiiAmdWnqF6ifSZkRY5vPzfDeNhCQXGcZOedZWK
kJSgp58pvgs0fJiDu0AC4j9kqBSUG99BcT5kR+/+OcBWGLYuRNhnkrDE04LB0+N64T3FM3WHl8ik
NDBL8FLi7iLPYmMYwxeHIoWTjAKKNFJeGaBmKm+GgtNqckoJp/PvbkLMldvC4xk8eBM9BETmcly9
QMGKXIU3+BRSx6JVS2UappEUtK/1VyLh9cXOK6+7zpLJfc7vI0WS9+k29Qt2tEUeSq+h/EwGRZSt
6/fRvkjXQYOv1/zu0bXPXy+mjGODJ0pJdetWUJoo7x+pLOpOcam8MFzA4EaFDVB7znkB9+9n01+r
WfGXN08nm+lIiiBKXuEZUzGTD/6ypRNFoxhTN60fe16uARrPehtn6cqD2cREppqximeU4QCkNLD5
gA6L+axgK7nIoPUJibd9xmAuQRzWN45ozW3dBk9qnjCWl4b8XLmRm4wnWE3KC+UBMV+3Tjty+sjq
wA7q/XCZaevPzlAfktnNfRrj+zW1yC15Hw2lG99oVa3jjVPoIeXplq+fYJ04UZkmh/dMONKF/cWc
NHG3gblJkjzoqBvU8gRZJ7ECMPNohqhGoZaT6SoltrvmuEwaELEybtm58vnVoAlBnq0xpAGlPjDg
qDRQs+Otau2uB3TkN2CMw4K/u584wL0PLsoQ6rXGEBFzJim77n+XfNo1xcFeauS8MaU+x5Ezumko
XAyBxAHkkULeeWA760aRf7nGXQbvIYIudj0emHrIQICHmzD9i2VBqwnoCJamNyOtDv3+lJXErl3K
L/ZhMvIaYKmrdBd2a5nvzV7ZULg72GckMapnTHIp9wYN1U3rGZcOfDmfpnNjYoaF99UYXw9FT0Fo
e1mhw+XXCYBHZulGws/mPGQ+Nx8reLaif5/ijZn4S62rPoDb+YqUMzl+hb7tslglxL/cCO9On3v+
OnvKkD5VZMA1EKxr995Of9yYaFvQVaGV9c+LJwsMp1LSNCXwdZbEk5XQ0dDDJFDq3iU5nFy3iiDy
ZFQ5Zls5A57Hq8G1dbzWQToUv8OGA16Cqzhj23f0Fb/lzyJTAUpfq/nO/DuQFglRFwQPlBpPaoKf
Yq1FuxOI/ORGbnWD+Uj7yj/h1gNo+Exu69nCbJTWXHAkgxOKYRpsWXNbY/6JPzX5u/V7f23VxTM5
SsLkMUCWsOTZbr1dZ/srIopcY6KWTmoqmDtyMVdm3qUfswHTeuGFLP74Ldpfqjz1KY/GxpVFyN65
a23h8wYgtIY6H+Ao43bwWFkHIeieyBghscaR9Aj2MT0C0x8baGvkmdyIglKZykrMu7que0G58nVN
4Nt2b79PeJXg4ZTcpoPLmFZSKXe14aC7Ixf1Dm6a9nwJ1yY2+Fnqs1Ye4TWB3HJtLl8HCFDLRHRx
Uk+6Tff09/Re4IEFgEicUsRhncfDhOvl/+6j82694SLtagK9UNb9DUH46pLBPDkABCobAjX0M8F+
d3LDDKjfzoegI0eXPUBUox5CyWsy7Vljk7SeZ4s581nV5c7RVPwCfyEjUY4N9K/ZzM7mrOid87JC
fNutFiNGCm5yWULhvyGBTm/VlggEgcXWAwE/2b7javp1bQlYplN0F0JUOEsttIvxaYuqaksuHi+C
gpOLDW7jzMD4EZ+Xg7o1Bgh8jR8wRsdxZRxwXw2Z53VYlybo+MqXOcddqXm7dCJP5J9M9G/XNceC
doNv0jURZu3wiE/OYKSmT+mRbt9nhJIUbVyn0eJsBhQCtQwUFrto9gNb3fx0T/TQ3syrr9PY9S0k
lwzysM8WCz63Waaf99/cs68mZyWmNUzVFDO/KRnPtNwsfHQ1CIBhQg0AF+AByMtHYKaxiUQL6YMt
IvowRAZEpP4bRiItzrmzmHqwuh5WqDNO7mpnXPxkAmBG0xoqCKAdTw85xXXtMAWEHGUWmrZXBOKa
sovEQsmypJdaS9HHaID42iTVJxG2FahdOPOjDYhkIAO1hfvQzPDK+morT3dpmm9LvUW2AtuCToh4
q8biC0P8ViID84eKcABgelT3ObISWiZ+w9dMTmIz212J0npdN0tdi/eb9FaFlz5MOiN1XUwEEeve
FxiYIQfAWEYiYdgVE00ygUGEhditoq47sTWcUUMDsfnr8WDTNuDQ+dj/VDdA1vL2UkSo+OZGsy3o
M9U8vrOAqi+wrcXNzqQU2CKfEkpRDEfSW00WKlrQzGXZJkUZvd3ePTaEFQbb3rDwoHrtC3qx522l
2SSlxqyOAdTB1iGTBZ2GmvFjqVEPWppwd8VEgs98IZ3hWVWbWe13/pOotli8yvNK9FMSMb8L+r4F
JoyPz3cTaQd0rkZL9PQLbAwh32DCm0vi2j0kWg+N9P9PQMmNN0W4mOJOFpdkHjwjFafRQM9ycIho
LgwwCSqaOnEx/OAx4XFVUXOwIKlL7TQPxhAVdjkPIwOTwpbvgKvk+Dl8+Sc02e1nYaFIliaLMHFV
aRTOaOaeTzZrqUemCBuzNbRKqBU3sqVTxWeoPQu6e9/1Ftx4MVWMqfETniNezjYnNLkmUOE3KP3k
qLzjQdZC1JLfBboXsUdFsLWdD1j+Y7RPw2VVyyme+1MweImHADK6eKpJYcqU2QbNkq4OEt40+Yzz
y3J3z/D+8lO+2Le7O6epntiYFYjY11rotJKAomC4NHen3kk2hWQfRvWnhASNBMvnpO8gyaQX1Uom
tpymaL8kSBtCGfrgvYCbcLaZSq0Hoj1eBuoRkOFVaG9ZTYnCq/NJOjv15NS5pgJH9TfX9Zr5Fze4
+NywGYGFmbMgLv0+vyGYGAzGYBMyAlarmDrUg9+gWi7OrnP/PUOgCEUxtUcGMaCRf6cmDVvkyGhg
PbvKfHM7Y3EcDhr7z1h8VY5SeGA11JY4SIcTr7gQwPuT+Hwzt2H1lobEr3prznZrb6dXRQ3vZUYB
FZ5U7oRDlLRTQjpLUFb8z0jzcJlWwnW4O2BA6oR35NRsGSoxcHge+NRrKwB34GgaFRka6iHuZ85u
V496CqBeQv4e976uskc9QRhBA4L/uLOQ3O+mZ54X2wz9F+e+vskMRP4cV33bx4e763KU/Vg00Km2
Fn8ftp3hZiOd8ajpV6Mynlz0O1DQhxiMJqEn7YHHrZI+/j9jcv3C+ZbuJTXM7FQVhZtqK3S1Etgi
9hdLTVc4iXjHcQnmJT4CAA5tB/tbDFBnWxOxCfRFk2a5rVUi6rjkjM4Sz7Nf43WMJGbHzwfHRNpw
iGWwqzjMTlfS44y9VUVV1s0DZ2SWVvNKTkW/PEbor4OOfkNVKgbHM3TiYTKUSlOh5w3dENvGW39I
fOOh7w3oBM4eOkvo9sutAJr2CQZDSFAoXvgdctbMINhPQSb+bfcTWHYIAjb0OaOb/QaMYq9zfTCM
b07kvgiqJi18NkRpvg2yHRW+URoXcQsZG5WuqOYZMwkrvMwguJa/p+HeUQ2/Av4RYsTN93p+dxa5
+Af2CdH8bYRuTaJt830alYPJ7Tctrc8b6/y//AHFJjlYvYHeJN/BL4aFZ7IZfJHjSMWl+m655XZW
XzUhqtrMYWhpHAZC6AwI+sieS2jT1cMiGzIbyEBDcG6Mc0Rfk+rLQxTsMpR6Ir/PK1xH2+/ujxYY
EeN0LZulWaCPGmSbmU3vWXCOzH3GfIjmzHvr2wk/5WzRsDaifZeoehc3ylOHwMrtHstBUs/Zq0ny
U09CZTJo6zDckJom61t6k1wg7QVWwpPuIZLY/F3pUI3R4O3E3h+bNh2i0P7bNDYJClXOR8di4V1X
SUI1GdF9wCjP4bh0MjIt1V5w4bFwM/9DpObSdc8wgl7ffeQXXjKuxDmz9nc+xXDkPLtfFfgQpcwq
35m0UZpj62I1Dhd/fOUk0wOvQDkf7VcAyMIc8d2QW8IRf9Ck2r3gps7lxlJnb59qTsWf+VpNrVlH
EceoTARh70o4jDOCjzNFSj84FOm3C3sxxqv93DlUNeCrZYUQdk1ISHno6DsqbgwWIu2NeFvtYx37
drAD0DRiOqbbo69INgKxskZVu1l+CXS5KUsIfI4Ji6i3SB2ka2969aps0YPs1RrH2+m58SZnYcr0
xN+1qDAaRgQNEQ+jHDbxwBED/iDmjVIOVthX8LUVYHHt9mVSw+ko80lqTKkfLpdekpR6f2c1mF0R
ZWZMHLKvD/3NPg05YU6ycHdeXEYK3y+7L8hFVYZmXPMvJvX7AgUtC8Ou1jYapHS0jF/yd4cjVY72
fAW2NAjCyPlJ/N4GBFyr5Eyx6r1RvNyETLWy+cFA/3OkFw7hLYoBTzWipGNMhOJmUIt60gEYnkPc
BOtKnF68UfNVSGEnx2Z/8ZjwDr9MCe8Dl68JjndgLaigUOUVkFbPKF9Ddz3tlxu6dFwW5u4kBLBZ
nnaUtg3rIBTw+kicGF8NJQu82dIekIZfn5+vFSLHlvAxeO6fN5BoWcD4H44mIWVaXRWX3AYK04Ad
EraM3ECNcUV/yxII13VJB5BbDn9ZUsrW2NmVPXTkRpJNqkyHn31SKU5uvxTBq2jjCaosTwSGZB4f
gOPq7zrlY5hNR0Md3VYinJW8571qTGb7nt2wOIIFNgW4mZMh6YHZBAq/SYAtQNdOgHDYPk+klirF
D/fXZljZ0rDpdYbOfKTlIkpqA0LEkFfidNKPVvrmgEN1FE034bHHWBahh9ICwW3ncIwqKiGsqlxR
NwkCNyWZgUExr0yPCBKQswjDIrNLduuU3fP4fNyJGwuox5QrcUiz23JKyf1D3UEz+dhl0zZA4kst
XGadGkHMzK6qodtAuschR61NqflYm/gUvdANMWITGB1TI7NKDNt7DeIA4nuKvNXRsZ74QtO9TqpQ
Ucm92Jl1EBWloS7K7iyfMAm7sGMtTdPUKenr3sd7DbwJaHiygG6bkjNMRB5BaqYmgXJMcAPYx58B
L80c/ySzzJPZWHzzO18FHphtXrCNCKki5tyKWGrEXnNPHWodao5YmKxKYZsMsWwl9a121G1QkWqW
yyplWKkmQeO/krXYzU5gRA/ihmVfayNrb3NlqxUaULNRH+v8gs2CpmWGiPkmazKkrAzXZQ0fr3wg
Y9Ve4M6Rv4eqLvAoYBrczZF1GCZvu4HoTLdLIwJru+cSZyyQ1sEGXAhagiHVfRUZ5M3tWcerDLvL
0V0DDCKonALnRZnL3f9ZA6ufb7WoQiJ/1YQvBkoyso7eyLremoVDeIcyMWr47W/NKWidsalvlIy9
qOmhXUEqMIY7mYrWQcrvsF+PMPWFIuaZQWneeOFt0Tnb2zv4DOtp+hs+xQNtE51SSKYNWCz6VnCw
rg+nzP/h5rLgxqDlm47jhqifgDFLMEiEH/b10eVR8wP50hsOI02IU5xXdMBO0beolQycmwJzCm66
t81qCNwva/fywnHBbM7qRqg2XNOHfC9ba1rxG/isaTw7djWUJmFJDDgIIbWFVjHsrWdOsBdglXeg
4LAdsv9DQHIVAgDF3zmDIbV9zmMVHwGu/+0vvy6y7bKi2AjsL0T/hWMX1YY+SpPW9ZodhSEQogCt
80EgSIomcfdH4ZO+oR4MY2Ajnk/UnF+DzK3ZbiJOvtFZwHAzzn2wBVoVJeNQKjtV6xmlA7hItMMs
5vAa1A9wwe6dYgxWMngptwzvtkHk7TWW2dXPIw2Y0f45Ant7oGHVhHIm32ZuBCVpM1wSIgBYvnKC
BNBd+JKsTUi1+kzoU+ZXaNOcfvO3p/zPPrmUZ4LghQXhvLHra59adGjujEvD97jtIkNR5/r6Ku2F
QYgQ7Td8ob2IAtJhv0Ifmp48pIvjm8YjaFcJk2dS5DxqWo25H5fveCMX1zezIwwYk7H/uCwhHpZi
NujQlid6ZSOgRo2jPJoWcSEFNCssovvIi5TdhNtpe2I3chSxWEwzFgKYlZjWSvsXLoO9mj4msqdC
8pKhELI784A9/J57gCCbzUM9dd8QIEuhZWEtnSrVIwzK9wDq6keODAwLN2VdjosDQtBqQ7sIXkZM
iOZ/KzlgkTCl3RqhNolUo+4AnNfWPSuDgAqcD2dPvtvZqCdJT61ay6J7n0ZwReoncbOYpZ9KUcUY
dOUe8C8ZZDkgSzO0e51GGEa3xBauPWKX6VhojyL3ouU9FyAomGwJNt0PqbrH7l/7ZxJ/Hf+TfJWq
Lc67em+gGTmgQr92ESNni4KnDMAz+mOxSPjEa73VOoXUHxlCthjf4eXdmKFwl72OnRhLq6+JX+4w
0ETE7qCpJScVGB3HlHF9vD0m5ZaCan9ZFHyxv2UUrcs9RpzOcxmr1FdHzm9+rqJGgpyrTvR2484p
yULC1qK+1BMCSTy/I3eWmicY2CTawvIi+rAyIL95F7yXpKWWyMobYr/vToS1zZCon7+1hdoiipSG
OZBS2gK7l7UiuOpN2jmtGTCAjpjYnB3u9A6bBhjuEvK4/AQTNp++w6Xu7mUKqZDuA08ofMxMk4yn
m4pQWyje15VBPgzTe2l1y790QBhTVw09dstlMc+vywzKnILvnGP3dA2feCEJKG5dKmEhSGvwqjHE
oOIAbWeFO2yfwukfAzn4BeXLKftlkmsBCd1AJqw6sZEC274/et3n4e3BywLL7sX05UDytxYeaQNf
wmKxzUOjaYstMMDdc0wKiTuX9js+wbuJu8QcdYD7spYlnGUr4+XO5QuW6iDqcKH9o4/xW7FiqzU0
fK4uKffxQvMz8LWfUnhH09NBb1v+qAI/5F3oI/gcLS24LHpauhXBmJC1bgcdHz5h8aZKo4T/CFL0
2QOghYmAKxkQtEHiHPjks59Nx+RLzZvGSiVtkIxup/4Sohj4ESHKDH5ERozUMZHIz3Zfb3jN03z3
5h2DJKmL9cjwLjDmX3se05xbdW4PToSK8gITZtJ1we5onuL0r4jtQpFJbGruvn521zIa2lYV54CB
O5UfPaMF6MjF5GfTVXLH6WeBxdqzESNXBBdST3ixIIkBwuR96NaNLR0wOzEQEfa6PES6HNCSJorE
gTWzGb0Ex7kDJLUV8juUmkEHuEax17mG/wWCO5TlRVrSfvTdYV42Ufl7rDOdTP48BZqzFIviAhGI
8ntPORZ7vfKs8GyxdzUxOaSJ78FvM1ZD46sLJFz9HCOPQgTL8sDJwS/y2FfNJ+tduEq9Xc8HBUXz
nkS/5/ofDxI/FViKGRgTQwnq3D8t7i/9vmETgaZVDwjDLME8fg5o0biPbCVp8IcFR27GW+nXzjoo
N4upO5zfaSb0ygv7WH3y4aAe7YNSEjV0dZMy7YnGV/yw34QLHLfr5osz09JESBVjlKkscfn98UVi
tmYKmrJQYoTODbN+JdCPcKktrZCZBf//tQl2Ug7jC+T3RocOR+f99k4n6ru74SAVdqQL3tUJ57jH
of8pZMLPasQd5djfNJrvruhoAQJD+JE5HAsZmfIkqwBgra/mAdoncORX3KWdaxdlnrFXp/Y1zkcu
ZyvLUSJ+06P6VdG/cgpxOORkAlnEV+uJjoWrFIgL1TYxoyBkFBRsoLEVMpjZZE1K5WElC2WSng2g
MDrbHFurKs0hGpHVDHTmPxzu8HTglgTVT2h0/WXyMnqfcdgos4aQiptmQc3jldsTyf5VZucJ2LS/
WcoIW9HQthJSwBQhldH7zIhl4nlgYFff6J5Uxvx8ldRVY2504zymZG9J6BlgQMD93C6EF3kXWYY9
jnlwmbuNJYpWbul6wCYT1qXbTih6K3N6k4iXHCzuS8m/FBEInYrsgU9+yVMItbujaR8sszsfPW0J
xedBJ5gW7DzrmSklZmM8tQIO2c03BvkOdyj001l6bj8cDoDcVX40lpZYSOe0vDPVsZyOU+Fg0n/h
lRsBafGQox7rmz51uJk/vbJlP3zmWrEsZAmNJMBa93Nl8pnnyDdUz77PU8Pjdnpt6ytQu4ny1hSW
JM3rPlTIWuqQHog8jPdRRO4uc//1Zanbgnk+hnVceea2tbe7l6s6aC00YuxqjluuQsE7s4+5HukI
twhwlRznRP60G7+zvmdYoBlFfv4u74amVBUesqiVPmfpR0IwPWfiHvdqHL2OrULMuXocOT3oo7yj
G28Pn2+h1HLPNM7WZU7zqA5JBgDDd7ZAHL/RlQLB7xrPWvmCIHGTZ3sJ3vRxVfbhAmR08SKPXHV9
N6Err0WnQhlvyOXXvK5ZOnYrVLbxQLpxNpFJMb4/nCTuW75Q5u56opjga1UUut1Z2aU0V+a0fLEA
ExxgD5/P8lCj4GNwxd5WSk97BgQg/X9iZgOqpceAzyzmsZsq3E1AW0aza9sW6A/FcJGEIaEDhIdP
nq0ddtORHynezKn5RK0HPPHPpun+gCnOc0XftxIHFh6EtbRWnkDOe66NZupbf0xWnnbEMPRC91WR
ATJq1UCXwaL4hREypXOAxhFzHRWPFaTUe0rR6Bo2JtMgHBs/sbsxIUPfBViI4PHJPK3xl27m/BOe
Y7jRjYFdWH4ic9hhIAZyVRBkOFkKuxdItGod36308pUQ/CI5j0Zqm3s8Y0IsT49PnFF3mHoh6Nzq
Juiu1RtKbKw8IRrPEVk1vFBscRS51t2W9OfqNz0tvHdVeD+MSwFlxZfKgiHvjJCcLhKixe6NiC8q
7iLloSNNAV5qe7VJkr4BYbYAb0eYJqcAt4jRwEBR8h0uA1ixfJgyBGg25Mmeqgw2sVHZHx8fA478
dfc3TP+gcAzTC/AgAof+hml9dGycuCfBAhaAxUzqRk1zPpm0MHJvu20Ds0/XRKq3RzKKZZwcEAj6
sYqBCg4mcxrCAtqBg4Jas/tS6ExsbQ14XyZBON9mOsoX01Yf0pYCamocAnp2/1Uj51z8S+IYYcPn
L48AADyZNGoNd+G+RAbamXVCNg2inHh38PXltk5Xd9qasei7r8UTvtiBSvgT/hoOA11V56X8i8yU
vqIFjZYwfdgDDQvju4GZUsoROusmRbnHndkaRupGPS2oEETY+sMOfdWuiJHbTkUOCUWKgg4CKgn+
wOsDBAex8vMfvsVKzqQR42hLNvyHpbp2GYxGy3MilGcm2YDVVuT+2HMet0Q1hQ/E1OCHkeV+Iz3Z
1lB7BByLBQ0vu17zRH6XrsGIzF53vD5C+UNkQBkYs2u1ek1dOwRrXmi21K51N7BYcfzzltZK9hTi
uKGqkQ52W+Bd4dPLFg3AruBEwtVJoy5GIqgWW/ICfVhNM3+9P3wJkTiGgAnrQiB435OkMBapNQ2M
Co1yx+xCNyTJ8ZGCfhJIPZOzltDJrtnJppPY36kmEOVIvBrSEUQViWmOogclp7ANIR0og213zar3
XajZlBRLA2ANCaQqlq06Fl3f5GM4LgNBVxI8NxzFc/me+xdDSV/L8JTVCcMQDMPqxOp0n88xahf3
f+1Nno76lDtBbDXtjph8EWWnyUY2TxxyZeohLvOEqQZINfHKZDmUQHub1k07vNkwgzpbIq/wK246
zTiVRVYKMVOqdtgy9FaiZxTUTTKx2mfV3jyj+KMiCbszA9384U//3s66cSMMyhgQdPBcDGQT+M/J
M4Nqp1vrCEnq96tDDvBhx2Txdd1DmJg9GQ5IHvuusTbwfbkfS5Y9h7KQMdI0yKRdx34MWiVwg8EB
8lHPhwU0sxKoJap6emyXfSeCd9nPY/srqJVAJHesmFggoPr38M5vzTjB/6XMgRxD5eblOcO6EdT9
UM5nKDErY1BsfqmnrC2Gv541dlPw7PCMEnzKI4Bogurk4cyAlfxfKPsS0IT93Z4A+mUsbj2bi2O1
WjsLvp+kcLoebk7tgHDGgnj/gyhHA+oK7/3XXXLnjykFWzzTbuvsdy1zKGANZsnB9WrXyFmXxXYA
xVkOFLOpDNk4GKu43ZjZygUF6SzH7OepK9lNYebLYfiBfaVXyRgnKkhHl3uM6Pm9NA9ASsiI6ObL
dOTeWixrKemY1+//cBVOewaIx3ozve703hLPOp+JRllt51ipdKNc3Z5lfC96+hHPkoK+nIoQLqo1
IYmpN7Say3QDw7gN5Rsdra7r55YDIb6944IR1qiUq2MvnD91Qzeo2IMbZlZqFJiX6WYtUiAJFgjE
tVWyveqdYFqyB4IEeXi8GKNsgyXIdcjbgsqZq3whXfDNV7YVXDwiMmSzgDGjepa0u5OcX0Ciw+zc
DGGpIINPcQHmLDddIVbyQoLrkNIFQMGtTSeJMLdsaEMQ5G4tY4j7F1A51oa4hvWMvJl6O6eZVZXA
aJihfcMcyh+nnuAvqrEty8GjPQCjDtykDwtgq/r/fCzGkjdezshjruz1Glg5c/12OeltknxiXRPT
hl0zfFTla/ZdMGl+Ylsg5XUvdQ2Ecw1FnwClsOupPXICtDfeXVekW2NsYoqdL6DZc9dD0ot2hcef
SlT4SW1F+wNAqnE1ix74UrxBd8ZEoJOHjM1wyinmfsqu3voKE/lJX66GcI6HVZb/91Q+xjXfw9nU
EkxgC8YhIYbQ8nzCQZTJ4kOdbK7OesY/9dDd8vFhZDu0Au1jQFcFfE1bc9QS5k641wgICk5gkxP1
zKh5bHOq5TnhXcH3UyIa8RpPaglk10IDR0x8yygxRgAMyQvGLXsrJfCGm2QotknNFgFH+28cq2jO
c2HdWddha29NvIX7gLWU7PRpjGxEyoKesDigNXnNVMuPn/eD7OLZhijxjLQiyp+d31iryM/V5Mor
AVHdyJmLHT9J8sVPND+Q+iGq+B25YHUGJK+Fpp3szk7Wf/rromNshRGTXdU59JVkVZ9wsHKHHkBT
WeEFXCuZ3BYvldIo/2bptFAcus7cjvM03GHy8deETyvB8UwI9pGsl7YupSgmSR5uJZXHnlWbZqc3
t04onzmVYLzNnrNFHnd6MaY7gfcmA6AaphMh1No5bdFr/1CQnlQnVnUfhWtKuFUoTzdKyi/bxWx3
V3fYwQTE3RMv5FTX0JApXYoEUR3B6SCU/Rmq7Xflg8FEljVu9DmGKOp2ROB85t2ajTvw9qRei7nE
HgAXAPuAK4TXzlXzKfBf7RN1QIOS8Sd55+nYNzIpnBgXrwiwlwskoildCfTcuAYi8FLHlB4wyZhZ
S8yicLdabnvHssEZpr+eNpkvIJ+VYvf5/aJTZ7wQUgAP5RwZGp3cdM1BKO9vjDJYZp+RY9HL5LBg
YwX9or3vQVKWrgjXIeYgNmpvTFNZ0JGCflGfssOG4PGnabIPirD+TT3jNScNnY4zW+IQrZOZlQXv
If1UYLB/2wrDurpT3M51vvqDvapIT2AQ//dHukzCwQhYcYgkzfoyWD4KIVYuDYPKljY2xcjcxKOr
zd6M5BxVWOW0RBatC69aqCa0AwkHWcIWLl1yU7nxM6VxBOwhsw86cn8sCVazDWkUEYSCVxi+tGYj
jrZkBOXQ5Z9AonQA7QCiqFQJbJpNyBZYyCLoV/IIo8sGTJidK7o955l5JuSuX3nQUpB5Z0T076c0
DFW5G8RLh5Ki6J9xQQcLOAcugQG6kEw9KLYL6gFldpe0c//FnTDcYhjD/FHW2nKEmAZNlgsas4hZ
+u/OcyRpOtFtlYZcDE10yxZ+/OG5xLz6yW/4ocWyukz9BDFB61jpqiCYp/5WBvz9bW0a6WoEQwd0
Mj6SHtbTdeyfATLQNid7ts/5Lf7xizn0wqMABfYZ6CPeP/yeJXaFb/GGAKGlQq69miUK5HdxdhgQ
nu1Wrn3F1yQHUkclZdGFn0wmY6lw/4rnZpboEJgOjt43YhqJGEao5ydvqnnRy+LhXxF21eoZJjSC
MgmJDZPM9KjQRQ8mCEhUjGQ/5dUCTgdp6+8WFvYyULiIQf9VAj7WziS5kW9/QUUy+36c6y1xiBJD
5/8e9l+DKLB680/UID/InU9f+8gDv9LqT0TDKoIi4Qi1r0KH7uAI2o5mVvKTjkzTRtVJIBv6tVCj
3AbXxnUnUD+ycMvVu3fUf8IaGXLZEi58CQ/5T3rReg7OFi4KbhxMjDMgUihXq6xzOZim1pUBw51a
2nX6lY6gVfxSfzEh+65ILMcq8sqOMwYRwMlIU+Tiu9A5ygbswvMrQQ0HL32Bwx37jgXkSvd8RSLC
trUp1YQiXOIO1Wigf219PYoDWnQPKPXnDttcl481gZ0lfW+VKZ/TZmkacN1e1i/kS4MtS63jlkzH
m6jOLpxOm3y4ptbDQmy4eX3PmChNDrShCZVo2je+KGumd3iUFxs/sEXNp/qDy4huYMh6QRkeSSCq
q5t1rRUXl9j0hs6yN2njiBZ9QQIgdYoNIB5huGlNn814Zfpu2pAm/hW3L8+5+hAcrxlWI9jAO7HM
69a6taesGrBD+5N5yXdJPBYdXdbC4+GZPf7O7MmxzMZmU9c0dIkiMhFRJhv3Mzx/NO2dOZb18clr
JEg6mw+tPlcepsx8Ag0iUcMo0NdcdBWEDZygogGvG5aYIh8NcDAYD9TKgMahNOwK/9V7FZop3XAv
iE7T8Mc9+HKqbBcRYvAwhtIJ0b+xDhQC97b0vYwYnnz6VYUJOz30oB+PczWmu1SmoPetG1TdUsq9
Toub/AFt+sKDlqFl+zCV5Gc6NFH4UWThIOL0g8d0E++MmBK/T9Y1AlKpBeQ/w7jj7FjYL+SzA+PC
z7nCXAm4sfxISHzfmwsnPODn3ytIpxuw5iFijHFUFAMTGBPK/q0KxsM4Rh5THPbiS1dVNNSpcBf2
6TYk0w9MKC9kRGGutnVUls9K4Jyv/nI0dRPWHI0tSs9hGpmN4kbQ1Qq/2MqRVD06vBWL8LSczR//
tdoZTdQrbPhuuCo9rpTLYIkhksVXEgcZ05NFEOIx/jAbafRRROykHByHG9lOb4P6nDj9pkJh122Y
CbZh/IyNrAFEzM4ZDBhz1OomDLZaz4XkO0mjp6j4hEj7rtJW7az0pyYCqk4Nk2ZtUkKceldzrSQX
UwHullUOcVpMARjy86zkjwtGQybj7timR1i1AZbFis33ZMZIY9VCfxaclX89dsm0nt7h8uCmZd7j
hyYxKZBIep0hcr9DSyYYlmBM/xkHVYNLIrz9UJE/yokJpXpFPoY8xp89HPLWQrha4kUJijoCTmqk
WEsfVXIMh5unqmIjbaIPE+qhPdYJ4H2HKfZxIxT8tdfdwHlLlibZKXx8f402flS8w4KWoRLbRN3/
nqDtaIbIXtL+8Zc9oXXjq67JSlCc3VyZY1q/5Xijv0/sqD+ojd4RAo1coCPz/tD0+id1V7WTFfdU
0qnS5u81q2HxEqlLirSP6+SK1suxvjuR4hXPqz68NIikAONhmHGZPYsuZkkcXTIo8+YFrLk7fVwK
R3N1JtvBf2bSj5HXVvgUT0eGcmfzemwFUywlFxQ343gnXvP9UhZXJKuJ2LEgmkqTcJlg8SBTmd/k
1HiKqC/r4bK3Okp2dkI3iLU9ChETTZZeaCral3aaqR887lU+D61w5vQu6eYADfwjtxJ0MYRsfJYZ
mWXsJz4nFW3hKb0Sqh0usoIn+xBCxi9WjpDUR1YSASAp4WVrlUCuheaqTIixoM1Ayci2e1eEuTWG
jRrOmMXw7RfdL/HwD9tLhd6hCYBW7YNAZ5uAtq9nb140Ig0TWSxA20UwEy7Jbei80xT/2y2yXf9H
4/L+wntXGENQqpfzQJM80qOIGMQF3tT3QVL1xX7LDXgz6rjpu8bUNZJhBubBranXNDpDVybEsIRe
6Mp0RuKagk+yMQY71KPFVbWzC9v8zdA1ZwqATYl3mp5deuw2eTzul3VglcWBXGQ67bre5r4fzN/z
tRBgK8vAjGjoif9O+0W6OCQSaRLM0jtgYe1pkQsm37U4zbOGK10xVv/Ct2kmXBL9AF6Wf+/qrNFR
RB82qqBd8FyYhzxD0wDEY5U5vdIy9q1aSHSfpy+6tR0BPNhCFXIhoRK+S+4j+DoD7XQkNIzLdAr5
gEyHfaqDVGHgp0A9nFGcxjxUdHOZF3hDQKUTurpGtn8KxybC4k8QU08D2F5A52sb/qUJt5KFr7fa
iQzIIq28f48U6fHcp5UenDVg5fJYqJT62xME8SUxvI0tpFwca+krvJExIaXg3fKsp9xkuhrOvwv9
eK/Ab3gSasNsbdP0Pri3J0wPL+ABkIw4PZ40Oh8tdewD4hB0ss7NRRd/EvYlFkOL1RwG8Ss7ad7L
dFmeBJyHkcykZ9k+yXysiU3qhv0a6f/1rNSljiPoGeF2NzwzFOI/UEsMBKCypmibStNGRDmcKxAE
Z2fqGT/RfRs9HxQ/c0e98oGbAWQcsDu0uVGY7M2qSAgcnglGGvHNuXQ8fqf0CJeMXzC/p4qYsMiw
rVJ5/KQgi57uMCZ/XPmHyS6vxyeX1SjbbSfQUe+CA+7NZNLvZugHFsFqJr+r4vYpwJoB8oSf7y0X
P/HFhkbtrcoYuQq22z/sEZNTs7znRp9Uxcv9Jxy88zPpH6yz5eY7Fuw2/klD0xYaUsoMbqb12c6G
BzzFyhnqJrMm7yVQkIuhfks1LbjODIN+tRtmeknIE63xX12VhMaJgWULmpW7zhi0dzJS7q9cfKLS
v/+XYIeX/Ae+Oeu1Qv079BZfZ0i3HON1MZXhyZL+3BO6swfqfOZMMb8UI+U/HcnpStRP5zXa7J7N
8/zJbLohyyyxgywnhEKqqYgpW8V9Uk3aO7pnz+Q/eFgBM3ldXdxTkGr/SgeTEJ2+ihJ7nRRPCSxB
aZcZKn0wacovmdxO5At+mV+FBcdKIn8xxCtJu0btVOxLEHzFNa2W5ClQKHb58F2Op1pvEj8G1U/f
CV5xnQ57WX1kLBU0AX2TjYwGsDgsyW4GwEGCJTQ256UrrdT+wZNxqwNhyKZ/h4+9df5eLlW5XO9r
gikK7swOfmj5AuxGaLVFi34qINlc2mIesB3wzaPT1z6APsyairWGl95qJO9dwIzjYBYaDK7GsXe7
262+ZCRiYucLbbA5f45t1qbwJyyTmgORj6OnfGJlG3mtwa8GlLwDJlvsrIqz0gfECZHJ0Fv39OQx
6goZqOPRxZk8Tlr5QmuDn9veEG4CxvFlbHDmOxlv25vKzXgBK2nBy2FF/KOXw7DAC/qHtSVviISn
vMhQjgTveM5UsnnT1r+IrLi6Y3FPpxuCduYjREGO5Gonjl1cnhgSz3MT3D+AjMeJ++jN3is8XLE+
vWxsjyuxkUNFFtNzr1Ejkiy+wwhaFUPzoPGNoIH0+SyGYLnvgcMeRBCIJQSqHdGfMVM/gF8uvgdL
cHavK48xk00hz0OO/QEvjEG2x0/3qIa3DSn9/OuR3S4J8iQzmtNwy2lqNGUMX/oiKtrHquHOGUvO
yej52r+fWYxlhPPXrJYW3Iq/OM/3rShiifq6Qm9UsXs2y0e5aMgLZxnGPD7tM8bRQou6Cm3zLjqP
G9Ig3Tw7/QZgJqy0/ikxp31ibqmwyIS7Rr2QcIKXppRkr68/3WpbL3jMa5LS5yeUb/ZdQ5Ca2MdU
a8eO59xM7I7Ane533UwXK07taX06k5cQ90I2it36RY1w0O+H1jXk1+Io1gjrYzXZPGmtEMSShMSZ
8A4uneb1P7peC39r7Xkf6NsMb2LLCpT6CW6oXlNExy5rUgHZvTBhRrZhz7hVxLvrmVh5jRMzJHLY
j6qRD/iAFhBOg2Em+G7QJemvwUHXTkgWQZjGqf1czQ1dw54Lei+hExmVMmAh9CMCWwm0Izyfl4Se
dDrQApKSxtZk+tYRBYbvxEYK0w9pZH92iFwvddK6BRIeN/urpdtLsgyYxFllb4tG5Ia0WMeFBh1W
16rmc2ZrM8Q6AMQn+eRmYx8zY3Nfjsaty53nm2m1Js5VPIvSsW+GT6uFc48eMua5rtlJ2Fe3GWps
SEkkoyvXNFuPnebDYgBgagVvEvYmLBk33WAUzmgAnCQoUCK6U0no3FqJRevrsIJkAxjPGWCBQMx3
G871zWJy6bIZBaAsHET2C5igsU7ao6HZXdCQAxf267OwFGfrthWB0ozY1nTkezWl1/QHfY3/VIVn
uW+wc5MmDR3d9Jdxc8xj0v5dTaGlA5e3D7rP0Rh5ggg3o4zM+z+DjiwbdDoOxu2/Qt1VtSdQq9Jp
OOKrvOvwH0c54RzAsDGHjRdrx8RPcCKRfCpLJ/E3WdB9EIM5dIXyT2OZbPoQ1v3ZfcRoElCTj1N0
dW5cFNWrjmyR1twmeO7dvGtJCMpFgSrQndCZYd2YF342p3FgsZpMQGEUmRMJ0m0toG7yr+tGbjbH
2zFS/3Eo2CEDEjcto2VrQni+7KQuOUjkcwA+TXh6/ggA9+uymvKlKEcYOvdHM90mYVS2hErGeY7W
V/3sngcl+pwgCLo+lWoDv33ANpQHcTaCLiWyfWp31Icvj4Z8TbRWYgz1UF1xmKGga7vbGyFr8Xel
KfSKkDkxnMSYoRE0rz/vQbMqJqOrSTg8wQ7+VKPYrKkWMIogh6PKhAlamU9FAO33mMnQME9DUDhh
fesHYIzqMtxfner9+cIDbJS0tp+jMKjxZuj7stG9NngM0otRON/Sj3r/iT+3xuWsIVK5n9lRjpV6
yoK6DWs4bDwvyL5OPWOhEjvhz13s+eSihE59QPervubLiuSckM0zAK6BS9WNVGvUwwpoICJ7HOcQ
ElodDlJ5Ss4c0r0Xg1YDqvCHrxvUN6lJABWc03BY7lU7dbP0Ae9nj+1boo9WcOQxgF7cj06jNeHo
NLOPCci8sgS1oD+O2mj3GeCN4Ynl4UzCCE3KN0Rp5tGv1NxaZiGflmOZT0AWIKz4ozmK5MY8v8FR
JCt5j4OoABUv/cjI2N+5w3tAqGNBSXRtGr5DWh7UkPe5EPM0BmWCewdAEe/PoHZxlLIzQLGRAWgT
t1dazqyEEq4XDy8rDgrpgpzatD7GArU1aoY+qzN1T0EVraX3UOWMCMR1fZx5yILT9WZpKbqfXQBR
5AvmxUO2ielnTyllu0BRjGl8cZbJ5U1BUlqu8JceS238xMEBzsMbp0nhOjgiC2u+jjl8JvDxkmnW
kqyFxka9HES6lwxSgFGCERCWockjWfdL00priYCiXa7x1o/gEb4o/LTJp7jEmSnWmItfKLE9hWw3
yf3dqu5iDLRr4Y+nr5anHEh1gy5QuPG5LAGZjEcuBYySn8ciBxiX0cxhiqZi6Pw8KDgA+PUmqGTn
nO3mo1bmooCWEZrfRW+lO5auwNIqzzi8kaBesIs1c5qFkoHY4qA72Uzo5f69mkPjBdWELmr3A3XE
Wts2gXDMjvR1uDAT4nB1LVgE8tVHY3na07QU4B7vCbqB3ewSSQ2MGB/elVbKtWwfNktQuMKcCbwV
7ARCFg7MDfaYvlj5BwJNAvkUZPurf4DBTU0I0AHXzCYaBhlEicGIv04sNUgNBrsMFeTAMO64EK24
jjLF2RouErwubQepr7gjU1dx9c4/2R4zfdfZi8oQMDXDIYeWrBj9VnB5YohnZppmCQJY1rF+0vaV
L/NdTUuduBaZy1jZTcUjHxeDnQy5Vk+f2eRGCCAt4PhnnTq3ytxlGsaXYGgZllNm3JOZsWGSavlb
eNtlk6T0wGB+Payi72bxx7YrMCu9T1D3nqXUsSRtdhRn0efDxB1gqviJ9WWeM4hrlgEUNdJdwTLU
LWi4sbAzsQfmWW/dYs7mqtXxYeiBF56Z4QenGfXh45De4oob1uCqJ4vyhE5EhLra7KRh0603EOAt
GcQ+aG+nzDJYDNJka95/plJWyr8Sdt6YQp0KTO8kVMRaYmhAFPvpNcZiRx7cUDVMMrpz7MH2Bp3j
wRij1rwHEz67W9Mup5CSSR0w28Y2i5rGpCIqrxlf+ccc3nUZp9/KwFAPAddKqlIdD194N7bUmCN/
vGmWK1OfaJ4E8AgQQJP4fHlmrD2T0Xq5862OsEf1h4TRRxao3b4Vsl4+2qCbvDVR+jjDDCzAOljb
c4o155UVHOuGeUHA9kxfKIK9flg9XcRj2S8WKgF240fzhcNQQnJRPw2zjsSJ3wbKPCmQLr+d4stK
zVd19zBZJzpu/r80TsUTnhrCw1NQpFRhQWy+6bTfPKdd0tqPhQ2WKkhsbfR/skQO/L39y9HaLH4C
E45QVyJIEzduqAUSuOse4OS7VvlGV3XcByvCraGaeYsdidJxdctBZavlFZddrHjEBkrU9sygsWwH
//Meu/zBaoxRw2qzzCvI042U5rAFV0CPm21ngWq97gYE71U4r8Ks4eWOL1GCVx+zvh8JL07PWMal
BZsvEC5I7NItD2I92a0GTOYT11xP81tjx7TRMUcc6iIJ9ZJu+OkWLiV0br502rgeGn8x4ABV0lcI
FpkDkBCGLIxZ8LaH3MxARerm9K4FmbwYaM4/gCUNSKBy0fLwjwG/plKnZ+Z0nRdTjXqapbAiU1j/
4iUFI5/87cx1SnTEwcCt9s8kmJzYNCUYW64hFI+1MzS/qE3ChieJ6Mg5kAPCMhGNA999+1ZH5bbs
Msu2RdnQ981HdBOR/CU1PLX04Vd5GWrbRHA195LYjzwBG0jEydOTrj0x8kbYCfsMrsX8IbLNsmKJ
EgJDMFrK9NcO6Uaag3d0HmAIyBlrMO38Ej7iJmEZFDx7jA1AHZdRMEphh0SR3V4r0qPYnxm4+e4V
/JE9c7SoKRks/1GWoHMjN4bllBqVvmuTZGW3DE3ztgj1h0qr+nSjT+HfSACs4fqiMfFnztoPSA+/
l4XO8yUVgYxm5Q+kOWzFq9J5EnAC+1OTrQiLvryIkP48K5rQeAt93UrhaCCZw+V4/fQ13yjNPgyP
N6S3V0/zLEcOIeAUXNrrvVCpv5t2Bq9mPIbHwitGsnmn4yUlSwqMipqbBogwQdisac4xIPaXsABL
N/ci3+t+E6yhiSZ/bHN3daXfOOD8tSDQZrJjhl0qO+QF8vW/izAKZOxC35arJBCO5PmXnrxHAUxG
NuUMb1/02E54oogDCwzrL+cNColnD7qYGnomSM0Zn8RXGvUD06akGZBwp1/wCxgeNhUXPL6+KKxd
rNAYeGbObnXpHupKefhPIHAPQBPulSwCTD0ZW09vYR90ijmN1IfLeDIZCOY4uOp1JmVE1OgMR8Ou
YUaOSMyajzB6CkOrGZhCXeUadygjmKiZ32+tkxWL9VVi0/faoFWqZHPTOG9Ujw9ATT5hI5d19GBb
jPQbAxNkoBg7FSyqKRMogXNuSCDAVe8Y6p0gvKW454UmE4cld5C5PFahr2hkyywMVPl8wT0ZX2uR
nVZVy0k+9V4wmwJpspEF0LopOqbAYya818WCScZHlleXqlgvPv1f83tawPUz5p3Qlp9RMRuLThP/
dvfeN8mnFrRAvp70gA8AB6Ghj8O6Sn4rH9NoYyg3SBsnI160X1o/nl7T4v2RtYfGXKrVGohF3BtV
W5+tlZyQjDW6z2VtSL93oTyWcflW20UiWOgowQBzaikpKq/7G6e1QLPJlz8neJoQGK1GVuV2CD2V
nAP6UFiMGeoAWvEtd1j1dWteNfiSjaRm2/pDhxQfQSndBf41sngIDCl1bs8Oe//JCZTjbT45OEW6
NRx48HkPCXpiqoqLJkLoO6Yllv4n59X7Gy9JLVXbYTRmr6z8EjM+oa2rsbjU8xlDNkhMqnhU+RMp
GuJELN2n+99xbVY2M10BopUocqXDAXRJs0OPAhTPB+o1epYQj4ZMdAnB9mfdxGOxtl2Y+6ugpvKv
evPJEsGvPqsbvC+w2iWYqmn33it6xn2j0gFBq64b9xH2Dup15FtK9jI3982JYxUeW+btoLKk098S
tAionm9PlknvZKRjv0AQbjaB6FSo16MPiFXhoaVauPT8TBIVoIfJIYHfB0A2soXB1TEUaG3+nonD
jfpiOPACel/nbDgC2Kqp+UxCBZLWv1p7HxDLW/KCiwWKFA7uGfC15+7ZbrY2wHpqwlWTt9YLCBL5
DGjit4aYMgv+FMeU16l9ULMXhOxuCCB/w6/T/nqOGi22ruDYlIvwhxHi4F8fFhuvvymsP6Gf7GaL
F8aK+cqzXXyZr82gb79l4D7672BzLWEJM8FDGMsc2HtLpooFpsTJKR1sxZ9ABGIZ3BJe97HAyH21
QLtHvQZNOc6rpA5i1wKJPvzE859J42HgxkIo2GYWEU+Zij/ZYz1BuDlqZkpM+gDJH8YieYVKu4+B
oJ/re8acWMCGnuA3onz1vlR6+79Py/1xX6cAITnKisJBaBfZc538PqULMwdOvz9PG/UamSFZT6wN
6snaYx/S5/FBhyDt6GwvTMQvUf6uEIqPjVNTW9YxOodYeAIs7E6PdU94+MlPyItBxNwcuObhXnpV
Qi3gjQPBqCKuq2wmTT68JdwOfmS4kn9+yIdcVNmUFOUcVVCJl8FCyv/RNOxDs0do9qx2aSipCwzq
bWqiOag2h+oTxuJ2kQpqP5fau98Kn3jQHvGs/+YOLWFh+EuZvCsM5XM0eY1wUELJEfnKrJENhwqh
qVlpgV88x5BAZwpqIP6MJr5TZiHGdJPpjiPJUULKtQ1nCg==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity DVI_TX_Top is
port(
  I_rst_n :  in std_logic;
  I_serial_clk :  in std_logic;
  I_rgb_clk :  in std_logic;
  I_rgb_vs :  in std_logic;
  I_rgb_hs :  in std_logic;
  I_rgb_de :  in std_logic;
  I_rgb_r :  in std_logic_vector(7 downto 0);
  I_rgb_g :  in std_logic_vector(7 downto 0);
  I_rgb_b :  in std_logic_vector(7 downto 0);
  O_tmds_clk_p :  out std_logic;
  O_tmds_clk_n :  out std_logic;
  O_tmds_data_p :  out std_logic_vector(2 downto 0);
  O_tmds_data_n :  out std_logic_vector(2 downto 0));
end DVI_TX_Top;
architecture beh of DVI_TX_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~rgb2dvi.DVI_TX_Top\
port(
  I_rgb_clk: in std_logic;
  I_serial_clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  I_rst_n: in std_logic;
  I_rgb_de: in std_logic;
  I_rgb_vs: in std_logic;
  I_rgb_hs: in std_logic;
  I_rgb_r : in std_logic_vector(7 downto 0);
  I_rgb_g : in std_logic_vector(7 downto 0);
  I_rgb_b : in std_logic_vector(7 downto 0);
  O_tmds_clk_p: out std_logic;
  O_tmds_clk_n: out std_logic;
  O_tmds_data_p : out std_logic_vector(2 downto 0);
  O_tmds_data_n : out std_logic_vector(2 downto 0));
end component;
begin
GND_s3: GND
port map (
  G => GND_0);
VCC_s3: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
rgb2dvi_inst: \~rgb2dvi.DVI_TX_Top\
port map(
  I_rgb_clk => I_rgb_clk,
  I_serial_clk => I_serial_clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  I_rst_n => I_rst_n,
  I_rgb_de => I_rgb_de,
  I_rgb_vs => I_rgb_vs,
  I_rgb_hs => I_rgb_hs,
  I_rgb_r(7 downto 0) => I_rgb_r(7 downto 0),
  I_rgb_g(7 downto 0) => I_rgb_g(7 downto 0),
  I_rgb_b(7 downto 0) => I_rgb_b(7 downto 0),
  O_tmds_clk_p => O_tmds_clk_p,
  O_tmds_clk_n => O_tmds_clk_n,
  O_tmds_data_p(2 downto 0) => O_tmds_data_p(2 downto 0),
  O_tmds_data_n(2 downto 0) => O_tmds_data_n(2 downto 0));
end beh;

--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.9 (64-bit)
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Sun Mar  3 15:15:44 2024

library IEEE;
use IEEE.std_logic_1164.all;

entity systemRam is
    port (
        douta: out std_logic_vector(31 downto 0);
        doutb: out std_logic_vector(31 downto 0);
        clka: in std_logic;
        ocea: in std_logic;
        cea: in std_logic;
        reseta: in std_logic;
        wrea: in std_logic;
        clkb: in std_logic;
        oceb: in std_logic;
        ceb: in std_logic;
        resetb: in std_logic;
        wreb: in std_logic;
        ada: in std_logic_vector(12 downto 0);
        dina: in std_logic_vector(31 downto 0);
        adb: in std_logic_vector(12 downto 0);
        dinb: in std_logic_vector(31 downto 0)
    );
end systemRam;

architecture Behavioral of systemRam is

    signal dpb_inst_0_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_0_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_1_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_1_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_2_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_2_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_3_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_3_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_4_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_4_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_5_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_5_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_6_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_6_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_7_douta: std_logic_vector(15 downto 0);
    signal dpb_inst_7_doutb: std_logic_vector(15 downto 0);
    signal dpb_inst_8_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_8_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_9_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_9_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_10_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_10_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_11_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_11_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_12_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_12_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_13_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_13_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_14_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_14_doutb: std_logic_vector(31 downto 16);
    signal dpb_inst_15_douta: std_logic_vector(31 downto 16);
    signal dpb_inst_15_doutb: std_logic_vector(31 downto 16);
    signal dff_q_0: std_logic;
    signal dff_q_1: std_logic;
    signal dff_q_2: std_logic;
    signal dff_q_3: std_logic;
    signal dff_q_4: std_logic;
    signal dff_q_5: std_logic;
    signal mux_o_0: std_logic;
    signal mux_o_1: std_logic;
    signal mux_o_2: std_logic;
    signal mux_o_3: std_logic;
    signal mux_o_4: std_logic;
    signal mux_o_5: std_logic;
    signal mux_o_7: std_logic;
    signal mux_o_8: std_logic;
    signal mux_o_9: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_11: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_14: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_17: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_19: std_logic;
    signal mux_o_21: std_logic;
    signal mux_o_22: std_logic;
    signal mux_o_23: std_logic;
    signal mux_o_24: std_logic;
    signal mux_o_25: std_logic;
    signal mux_o_26: std_logic;
    signal mux_o_28: std_logic;
    signal mux_o_29: std_logic;
    signal mux_o_30: std_logic;
    signal mux_o_31: std_logic;
    signal mux_o_32: std_logic;
    signal mux_o_33: std_logic;
    signal mux_o_35: std_logic;
    signal mux_o_36: std_logic;
    signal mux_o_37: std_logic;
    signal mux_o_38: std_logic;
    signal mux_o_39: std_logic;
    signal mux_o_40: std_logic;
    signal mux_o_42: std_logic;
    signal mux_o_43: std_logic;
    signal mux_o_44: std_logic;
    signal mux_o_45: std_logic;
    signal mux_o_46: std_logic;
    signal mux_o_47: std_logic;
    signal mux_o_49: std_logic;
    signal mux_o_50: std_logic;
    signal mux_o_51: std_logic;
    signal mux_o_52: std_logic;
    signal mux_o_53: std_logic;
    signal mux_o_54: std_logic;
    signal mux_o_56: std_logic;
    signal mux_o_57: std_logic;
    signal mux_o_58: std_logic;
    signal mux_o_59: std_logic;
    signal mux_o_60: std_logic;
    signal mux_o_61: std_logic;
    signal mux_o_63: std_logic;
    signal mux_o_64: std_logic;
    signal mux_o_65: std_logic;
    signal mux_o_66: std_logic;
    signal mux_o_67: std_logic;
    signal mux_o_68: std_logic;
    signal mux_o_70: std_logic;
    signal mux_o_71: std_logic;
    signal mux_o_72: std_logic;
    signal mux_o_73: std_logic;
    signal mux_o_74: std_logic;
    signal mux_o_75: std_logic;
    signal mux_o_77: std_logic;
    signal mux_o_78: std_logic;
    signal mux_o_79: std_logic;
    signal mux_o_80: std_logic;
    signal mux_o_81: std_logic;
    signal mux_o_82: std_logic;
    signal mux_o_84: std_logic;
    signal mux_o_85: std_logic;
    signal mux_o_86: std_logic;
    signal mux_o_87: std_logic;
    signal mux_o_88: std_logic;
    signal mux_o_89: std_logic;
    signal mux_o_91: std_logic;
    signal mux_o_92: std_logic;
    signal mux_o_93: std_logic;
    signal mux_o_94: std_logic;
    signal mux_o_95: std_logic;
    signal mux_o_96: std_logic;
    signal mux_o_98: std_logic;
    signal mux_o_99: std_logic;
    signal mux_o_100: std_logic;
    signal mux_o_101: std_logic;
    signal mux_o_102: std_logic;
    signal mux_o_103: std_logic;
    signal mux_o_105: std_logic;
    signal mux_o_106: std_logic;
    signal mux_o_107: std_logic;
    signal mux_o_108: std_logic;
    signal mux_o_109: std_logic;
    signal mux_o_110: std_logic;
    signal mux_o_112: std_logic;
    signal mux_o_113: std_logic;
    signal mux_o_114: std_logic;
    signal mux_o_115: std_logic;
    signal mux_o_116: std_logic;
    signal mux_o_117: std_logic;
    signal mux_o_119: std_logic;
    signal mux_o_120: std_logic;
    signal mux_o_121: std_logic;
    signal mux_o_122: std_logic;
    signal mux_o_123: std_logic;
    signal mux_o_124: std_logic;
    signal mux_o_126: std_logic;
    signal mux_o_127: std_logic;
    signal mux_o_128: std_logic;
    signal mux_o_129: std_logic;
    signal mux_o_130: std_logic;
    signal mux_o_131: std_logic;
    signal mux_o_133: std_logic;
    signal mux_o_134: std_logic;
    signal mux_o_135: std_logic;
    signal mux_o_136: std_logic;
    signal mux_o_137: std_logic;
    signal mux_o_138: std_logic;
    signal mux_o_140: std_logic;
    signal mux_o_141: std_logic;
    signal mux_o_142: std_logic;
    signal mux_o_143: std_logic;
    signal mux_o_144: std_logic;
    signal mux_o_145: std_logic;
    signal mux_o_147: std_logic;
    signal mux_o_148: std_logic;
    signal mux_o_149: std_logic;
    signal mux_o_150: std_logic;
    signal mux_o_151: std_logic;
    signal mux_o_152: std_logic;
    signal mux_o_154: std_logic;
    signal mux_o_155: std_logic;
    signal mux_o_156: std_logic;
    signal mux_o_157: std_logic;
    signal mux_o_158: std_logic;
    signal mux_o_159: std_logic;
    signal mux_o_161: std_logic;
    signal mux_o_162: std_logic;
    signal mux_o_163: std_logic;
    signal mux_o_164: std_logic;
    signal mux_o_165: std_logic;
    signal mux_o_166: std_logic;
    signal mux_o_168: std_logic;
    signal mux_o_169: std_logic;
    signal mux_o_170: std_logic;
    signal mux_o_171: std_logic;
    signal mux_o_172: std_logic;
    signal mux_o_173: std_logic;
    signal mux_o_175: std_logic;
    signal mux_o_176: std_logic;
    signal mux_o_177: std_logic;
    signal mux_o_178: std_logic;
    signal mux_o_179: std_logic;
    signal mux_o_180: std_logic;
    signal mux_o_182: std_logic;
    signal mux_o_183: std_logic;
    signal mux_o_184: std_logic;
    signal mux_o_185: std_logic;
    signal mux_o_186: std_logic;
    signal mux_o_187: std_logic;
    signal mux_o_189: std_logic;
    signal mux_o_190: std_logic;
    signal mux_o_191: std_logic;
    signal mux_o_192: std_logic;
    signal mux_o_193: std_logic;
    signal mux_o_194: std_logic;
    signal mux_o_196: std_logic;
    signal mux_o_197: std_logic;
    signal mux_o_198: std_logic;
    signal mux_o_199: std_logic;
    signal mux_o_200: std_logic;
    signal mux_o_201: std_logic;
    signal mux_o_203: std_logic;
    signal mux_o_204: std_logic;
    signal mux_o_205: std_logic;
    signal mux_o_206: std_logic;
    signal mux_o_207: std_logic;
    signal mux_o_208: std_logic;
    signal mux_o_210: std_logic;
    signal mux_o_211: std_logic;
    signal mux_o_212: std_logic;
    signal mux_o_213: std_logic;
    signal mux_o_214: std_logic;
    signal mux_o_215: std_logic;
    signal mux_o_217: std_logic;
    signal mux_o_218: std_logic;
    signal mux_o_219: std_logic;
    signal mux_o_220: std_logic;
    signal mux_o_221: std_logic;
    signal mux_o_222: std_logic;
    signal mux_o_224: std_logic;
    signal mux_o_225: std_logic;
    signal mux_o_226: std_logic;
    signal mux_o_227: std_logic;
    signal mux_o_228: std_logic;
    signal mux_o_229: std_logic;
    signal mux_o_231: std_logic;
    signal mux_o_232: std_logic;
    signal mux_o_233: std_logic;
    signal mux_o_234: std_logic;
    signal mux_o_235: std_logic;
    signal mux_o_236: std_logic;
    signal mux_o_238: std_logic;
    signal mux_o_239: std_logic;
    signal mux_o_240: std_logic;
    signal mux_o_241: std_logic;
    signal mux_o_242: std_logic;
    signal mux_o_243: std_logic;
    signal mux_o_245: std_logic;
    signal mux_o_246: std_logic;
    signal mux_o_247: std_logic;
    signal mux_o_248: std_logic;
    signal mux_o_249: std_logic;
    signal mux_o_250: std_logic;
    signal mux_o_252: std_logic;
    signal mux_o_253: std_logic;
    signal mux_o_254: std_logic;
    signal mux_o_255: std_logic;
    signal mux_o_256: std_logic;
    signal mux_o_257: std_logic;
    signal mux_o_259: std_logic;
    signal mux_o_260: std_logic;
    signal mux_o_261: std_logic;
    signal mux_o_262: std_logic;
    signal mux_o_263: std_logic;
    signal mux_o_264: std_logic;
    signal mux_o_266: std_logic;
    signal mux_o_267: std_logic;
    signal mux_o_268: std_logic;
    signal mux_o_269: std_logic;
    signal mux_o_270: std_logic;
    signal mux_o_271: std_logic;
    signal mux_o_273: std_logic;
    signal mux_o_274: std_logic;
    signal mux_o_275: std_logic;
    signal mux_o_276: std_logic;
    signal mux_o_277: std_logic;
    signal mux_o_278: std_logic;
    signal mux_o_280: std_logic;
    signal mux_o_281: std_logic;
    signal mux_o_282: std_logic;
    signal mux_o_283: std_logic;
    signal mux_o_284: std_logic;
    signal mux_o_285: std_logic;
    signal mux_o_287: std_logic;
    signal mux_o_288: std_logic;
    signal mux_o_289: std_logic;
    signal mux_o_290: std_logic;
    signal mux_o_291: std_logic;
    signal mux_o_292: std_logic;
    signal mux_o_294: std_logic;
    signal mux_o_295: std_logic;
    signal mux_o_296: std_logic;
    signal mux_o_297: std_logic;
    signal mux_o_298: std_logic;
    signal mux_o_299: std_logic;
    signal mux_o_301: std_logic;
    signal mux_o_302: std_logic;
    signal mux_o_303: std_logic;
    signal mux_o_304: std_logic;
    signal mux_o_305: std_logic;
    signal mux_o_306: std_logic;
    signal mux_o_308: std_logic;
    signal mux_o_309: std_logic;
    signal mux_o_310: std_logic;
    signal mux_o_311: std_logic;
    signal mux_o_312: std_logic;
    signal mux_o_313: std_logic;
    signal mux_o_315: std_logic;
    signal mux_o_316: std_logic;
    signal mux_o_317: std_logic;
    signal mux_o_318: std_logic;
    signal mux_o_319: std_logic;
    signal mux_o_320: std_logic;
    signal mux_o_322: std_logic;
    signal mux_o_323: std_logic;
    signal mux_o_324: std_logic;
    signal mux_o_325: std_logic;
    signal mux_o_326: std_logic;
    signal mux_o_327: std_logic;
    signal mux_o_329: std_logic;
    signal mux_o_330: std_logic;
    signal mux_o_331: std_logic;
    signal mux_o_332: std_logic;
    signal mux_o_333: std_logic;
    signal mux_o_334: std_logic;
    signal mux_o_336: std_logic;
    signal mux_o_337: std_logic;
    signal mux_o_338: std_logic;
    signal mux_o_339: std_logic;
    signal mux_o_340: std_logic;
    signal mux_o_341: std_logic;
    signal mux_o_343: std_logic;
    signal mux_o_344: std_logic;
    signal mux_o_345: std_logic;
    signal mux_o_346: std_logic;
    signal mux_o_347: std_logic;
    signal mux_o_348: std_logic;
    signal mux_o_350: std_logic;
    signal mux_o_351: std_logic;
    signal mux_o_352: std_logic;
    signal mux_o_353: std_logic;
    signal mux_o_354: std_logic;
    signal mux_o_355: std_logic;
    signal mux_o_357: std_logic;
    signal mux_o_358: std_logic;
    signal mux_o_359: std_logic;
    signal mux_o_360: std_logic;
    signal mux_o_361: std_logic;
    signal mux_o_362: std_logic;
    signal mux_o_364: std_logic;
    signal mux_o_365: std_logic;
    signal mux_o_366: std_logic;
    signal mux_o_367: std_logic;
    signal mux_o_368: std_logic;
    signal mux_o_369: std_logic;
    signal mux_o_371: std_logic;
    signal mux_o_372: std_logic;
    signal mux_o_373: std_logic;
    signal mux_o_374: std_logic;
    signal mux_o_375: std_logic;
    signal mux_o_376: std_logic;
    signal mux_o_378: std_logic;
    signal mux_o_379: std_logic;
    signal mux_o_380: std_logic;
    signal mux_o_381: std_logic;
    signal mux_o_382: std_logic;
    signal mux_o_383: std_logic;
    signal mux_o_385: std_logic;
    signal mux_o_386: std_logic;
    signal mux_o_387: std_logic;
    signal mux_o_388: std_logic;
    signal mux_o_389: std_logic;
    signal mux_o_390: std_logic;
    signal mux_o_392: std_logic;
    signal mux_o_393: std_logic;
    signal mux_o_394: std_logic;
    signal mux_o_395: std_logic;
    signal mux_o_396: std_logic;
    signal mux_o_397: std_logic;
    signal mux_o_399: std_logic;
    signal mux_o_400: std_logic;
    signal mux_o_401: std_logic;
    signal mux_o_402: std_logic;
    signal mux_o_403: std_logic;
    signal mux_o_404: std_logic;
    signal mux_o_406: std_logic;
    signal mux_o_407: std_logic;
    signal mux_o_408: std_logic;
    signal mux_o_409: std_logic;
    signal mux_o_410: std_logic;
    signal mux_o_411: std_logic;
    signal mux_o_413: std_logic;
    signal mux_o_414: std_logic;
    signal mux_o_415: std_logic;
    signal mux_o_416: std_logic;
    signal mux_o_417: std_logic;
    signal mux_o_418: std_logic;
    signal mux_o_420: std_logic;
    signal mux_o_421: std_logic;
    signal mux_o_422: std_logic;
    signal mux_o_423: std_logic;
    signal mux_o_424: std_logic;
    signal mux_o_425: std_logic;
    signal mux_o_427: std_logic;
    signal mux_o_428: std_logic;
    signal mux_o_429: std_logic;
    signal mux_o_430: std_logic;
    signal mux_o_431: std_logic;
    signal mux_o_432: std_logic;
    signal mux_o_434: std_logic;
    signal mux_o_435: std_logic;
    signal mux_o_436: std_logic;
    signal mux_o_437: std_logic;
    signal mux_o_438: std_logic;
    signal mux_o_439: std_logic;
    signal mux_o_441: std_logic;
    signal mux_o_442: std_logic;
    signal mux_o_443: std_logic;
    signal mux_o_444: std_logic;
    signal mux_o_445: std_logic;
    signal mux_o_446: std_logic;
    signal cea_w: std_logic;
    signal ceb_w: std_logic;
    signal gw_vcc: std_logic;
    signal gw_gnd: std_logic;
    signal dpb_inst_0_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_0_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_0_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_0_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_1_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_1_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_1_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_1_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_2_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_2_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_2_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_2_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_3_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_3_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_3_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_3_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_4_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_4_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_4_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_4_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_5_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_5_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_5_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_5_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_6_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_6_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_6_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_6_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_7_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_7_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_7_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_7_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_8_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_8_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_8_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_8_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_9_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_9_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_9_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_9_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_10_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_10_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_10_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_10_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_11_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_11_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_11_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_11_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_12_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_12_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_12_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_12_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_13_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_13_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_13_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_13_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_14_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_14_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_14_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_14_ADB_i: std_logic_vector(13 downto 0);
    signal dpb_inst_15_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpb_inst_15_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpb_inst_15_ADA_i: std_logic_vector(13 downto 0);
    signal dpb_inst_15_ADB_i: std_logic_vector(13 downto 0);

    --component declaration
    component DPB
        generic (
            READ_MODE0: in bit := '0';
            READ_MODE1: in bit := '0';
            WRITE_MODE0: in bit_vector := "00";
            WRITE_MODE1: in bit_vector := "00";
            BIT_WIDTH_0: in integer :=16;
            BIT_WIDTH_1: in integer :=16;
            BLK_SEL_0: in bit_vector := "000";
            BLK_SEL_1: in bit_vector := "000";
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DOA: out std_logic_vector(15 downto 0);
            DOB: out std_logic_vector(15 downto 0);
            CLKA: in std_logic;
            OCEA: in std_logic;
            CEA: in std_logic;
            RESETA: in std_logic;
            WREA: in std_logic;
            CLKB: in std_logic;
            OCEB: in std_logic;
            CEB: in std_logic;
            RESETB: in std_logic;
            WREB: in std_logic;
            BLKSELA: in std_logic_vector(2 downto 0);
            BLKSELB: in std_logic_vector(2 downto 0);
            ADA: in std_logic_vector(13 downto 0);
            DIA: in std_logic_vector(15 downto 0);
            ADB: in std_logic_vector(13 downto 0);
            DIB: in std_logic_vector(15 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_vcc <= '1';
    gw_gnd <= '0';

    cea_w <= not wrea and cea;
    ceb_w <= not wreb and ceb;
    dpb_inst_0_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_0_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_0_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_0_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_1_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_1_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_1_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_1_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_2_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_2_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_2_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_2_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_3_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_3_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_3_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_3_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_4_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_4_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_4_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_4_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_5_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_5_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_5_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_5_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_6_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_6_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_6_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_6_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_7_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_7_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_7_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_7_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_8_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_8_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_8_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_8_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_9_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_9_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_9_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_9_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_10_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_10_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_10_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_10_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_11_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_11_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_11_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_11_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_12_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_12_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_12_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_12_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_13_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_13_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_13_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_13_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_14_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_14_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_14_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_14_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_15_BLKSELA_i <= ada(12) & ada(11) & ada(10);
    dpb_inst_15_BLKSELB_i <= adb(12) & adb(11) & adb(10);
    dpb_inst_15_ADA_i <= ada(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_15_ADB_i <= adb(9 downto 0) & gw_gnd & gw_gnd & gw_vcc & gw_vcc;
    dpb_inst_0: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"2E230413262301130000006F00EF26232423222320230113001300130013006F",
            INIT_RAM_01 => X"04E3079347038463F79337B3478305A3C78387B3278387132623871327832623",
            INIT_RAM_02 => X"17B78713A78317B7AC2317B70733F7B30793A68317B7A70317B71E6307934703",
            INIT_RAM_03 => X"959367B3879347B7571397134783F06FAC2317B7F8E3879317B7A70317B7AC23",
            INIT_RAM_04 => X"85130793F06F90235713971307B39793AC2316B78613A78317B7A70317B7D593",
            INIT_RAM_05 => X"A783A78317B78A63F79337B3F793A783A78317B704132E230113806701132403",
            INIT_RAM_06 => X"B793F793A783A78317B707A3079304132E23011380670113240385130793006F",
            INIT_RAM_07 => X"041324232623011380670113240385130793A0234703A78317B7F06F8463F793",
            INIT_RAM_08 => X"0793470308630793470303A32783F06F1463079327032423F0EF26232C232E23",
            INIT_RAM_09 => X"07B3270327838023470387B3278387132623871327835A632703879327830263",
            INIT_RAM_0A => X"2C232E23041326230113806701132403208385130793F06F0463079347038023",
            INIT_RAM_0B => X"07934703006F87934783E86307934703FE630793470307A3C78307B327032783",
            INIT_RAM_0C => X"006F87934783E86307934703FE6307934703006F87934783E86307934703FE63",
            INIT_RAM_0D => X"250385932C23871327832C232E23041324232623011380670113240385130793",
            INIT_RAM_0E => X"006F07931663079327032423F0EF25032583006F07931663079327032623F0EF",
            INIT_RAM_0F => X"25030593262304132C232E2301138067011324032083851367B3278397132783",
            INIT_RAM_10 => X"859387939793278350632703879327832623006F07931663079327032423F0EF",
            INIT_RAM_11 => X"2783F0EF851307930EA30E23F7932783006F07931663079327032223F0EF2503",
            INIT_RAM_12 => X"2E232423262304132C232E230113806701132403208385130793F06F26238793",
            INIT_RAM_13 => X"0C6307932703086307932703006F07931663079327032C230793F0EF25030593",
            INIT_RAM_14 => X"079320230793006F2423079320230793006F2423079320230793106307932703",
            INIT_RAM_15 => X"079327032A23F0EF250385939793879327837463278327032623222300132423",
            INIT_RAM_16 => X"F06F2623879327832223E7B327838713F7932783222397932783006F07931663",
            INIT_RAM_17 => X"07B327839713278374632703879307B3278327032623006F0793766327B72703",
            INIT_RAM_18 => X"7713270307B3270307B327832703006F07931663079327032A23F0EF25038593",
            INIT_RAM_19 => X"2E230413242326230113806701132403208385130793F06F2623879327838023",
            INIT_RAM_1A => X"006F22230793006F222307931463079327030463079327030463079327032C23",
            INIT_RAM_1B => X"F0EF2503859397938793278374632783270324232623006F0793006F22230793",
            INIT_RAM_1C => X"27832623E7B327838713F7932783262397932783006F07931663079327032023",
            INIT_RAM_1D => X"240320838513079380E7A78317B7A02317B72703F0EF851317B7F06F24238793",
            INIT_RAM_1E => X"87932783F0EF851317B770632783270326232E23041324232623011380670113",
            INIT_RAM_1F => X"F793A783A78317B707A3079304132E23011380670113240320830013F06F2623",
            INIT_RAM_20 => X"F06F8463F793B793F793A783A78317B7A0234703A78317B7F06F8463F793B793",
            INIT_RAM_21 => X"2A232C232E23041322232423262301138067011324038513F793A783A78317B7",
            INIT_RAM_22 => X"D7932783F0EF8513F793D7932783F0EF0513A6237713A78317B7A703A78317B7",
            INIT_RAM_23 => X"F0EF051304B3278327037863278327032623F0EF8513F7932783F0EF8513F793",
            INIT_RAM_24 => X"208385130793A6236713A78317B7A703A78317B7F06F26238793278380230793",
            INIT_RAM_25 => X"07B7F0EF053705B70637F0EF851317B704132C232E2301138067011324832403",
            INIT_RAM_26 => X"006F80E7A78317B7A023073717B7F0EF851317B71663879307B7A70327832623",
            INIT_RAM_27 => X"17B7A823A78317B704132C232E2301138067011324032083006FF0EF851317B7",
            INIT_RAM_28 => X"E7B32703A783A78317B78063F793B793F793A783A78317B72023A0230713A783",
            INIT_RAM_29 => X"2783A70317B7CA63879317B727032623AC2317B7AE230713773717B7F06F2023",
            INIT_RAM_2A => X"851317B7F0EF0513F0EF851317B7F06F26238793278390230713473707B39793",
            INIT_RAM_2B => X"F0EF851317B7F0EF0513F0EF851317B7F0EF0513F0EF851317B7F0EF0513F0EF",
            INIT_RAM_2C => X"0513F0EF851317B7F0EF0513F0EF851317B7F0EF0513F0EF851317B7F0EF0513",
            INIT_RAM_2D => X"F0EF0513F0EF851317B7F0EF0513F0EF851317B7F0EF0513F0EF851317B7F0EF",
            INIT_RAM_2E => X"17B7571397132783C263079327032623F0EF851317B7F0EF0513F0EF851317B7",
            INIT_RAM_2F => X"17B7222307932423F06F262387932783902357131713171387B397932783A683",
            INIT_RAM_30 => X"006FF0EF851317B7CA6327832703C86307932703CC63079327032623AC230713",
            INIT_RAM_31 => X"2783F0EF851317B7006FF0EF851317B75A63270387932783006FF0EF851317B7",
            INIT_RAM_32 => X"F79327B3879387B7270320232423D46307932703242387932783F06F26238793",
            INIT_RAM_33 => X"B793F793A783A78317B70013F06F2023879327830A63079327032223F0EF8663",
            INIT_RAM_34 => X"2023E7B32703A783A78317B78063F793B793F793A783A78317B720238A63F793",
            INIT_RAM_35 => X"851317B70593F0EF851317B7F06F046307932703F0EF8463F79337B32783F06F",
            INIT_RAM_36 => X"F0EF0513006FF0EF851317B7F0EF05138E63F793B7930793F0EF851317B7F0EF",
            INIT_RAM_37 => X"C783879317B7242312E30793C70317B7F0EF851317B70593006FF0EF851317B7",
            INIT_RAM_38 => X"0593006F2423F0EF851317B705938067A78307B3879317B79713606307138793",
            INIT_RAM_39 => X"851317B70593006F2423006F2423F0EF851317B70593006F2423F0EF851317B7",
            INIT_RAM_3A => X"0793F0EF851317B70593006F24230793F0EF851317B70593006F24230793F0EF",
            INIT_RAM_3B => X"851317B7006FF0EF0513006F0A63079327038A632783006F24230793006F2423",
            INIT_RAM_3C => X"64610A0A00200A54420AF06F006FF0EF0513F0EF851317B7006FF0EF0513F0EF",
            INIT_RAM_3D => X"6E6F73206F6C2065656C2C6574616973696C6E49000A4F42656773206F632067",
            INIT_RAM_3E => X"000A0A303030302020796D656E6F617269666320504674206461746F20657473",
            INIT_RAM_3F => X"202020200A2029202020204F207C20202020000A7E2820202F5F2E7C20202020"
        )
        port map (
            DOA => dpb_inst_0_douta(15 downto 0),
            DOB => dpb_inst_0_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_0_BLKSELA_i,
            BLKSELB => dpb_inst_0_BLKSELB_i,
            ADA => dpb_inst_0_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_0_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_1: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "001",
            BLK_SEL_1 => "001",
            INIT_RAM_00 => X"20202020202020200A202D2D2D2D202D2D282D2D20200A202028205F2020207C",
            INIT_RAM_01 => X"2020333034324220202020200A2065646C7462205379617420200A2020202020",
            INIT_RAM_02 => X"20200A2020446D6F20746220202020200A2020206B2061206572202020200A20",
            INIT_RAM_03 => X"6165202D4F520A2700276E6965630A0A00B000B10A202D2D2D2D2D2D2D2D2D2D",
            INIT_RAM_04 => X"0E240E6C000065732065656C2D207272656C72656365550A00720A2774657220",
            INIT_RAM_05 => X"EEB4001800200D1B7C017A01000000100EAC0E900E740E6C0E6C0E6C0E540E3C",
            INIT_RAM_06 => X"005C002044C8080C88444400004CEFAC003C001C020D0108080C88444400011C",
            INIT_RAM_07 => X"C844020044028148440000BCF00C008000240002C844080C884444000058EFD8",
            INIT_RAM_08 => X"814844000090F12400CC00240002C894080C8844440000A8F0A000A800200002",
            INIT_RAM_09 => X"011C00240002C844020044028148440000C0F18C00F400240002C84402004402",
            INIT_RAM_0A => X"0300440281484400011CF3C401440024020D44C1030044028148440001C8F224",
            INIT_RAM_0B => X"44000084F4E80190002044C878004402814844000054F4B8016C0020020D44C1",
            INIT_RAM_0C => X"00240002C944C1CC080C8902814C440000F0F54801B400280002C870080C8844",
            INIT_RAM_0D => X"440281484400054CF6740208001C0002C84402004402814844000090F60C01E0",
            INIT_RAM_0E => X"00000000000000000000000000000000000000FF000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_1_douta(15 downto 0),
            DOB => dpb_inst_1_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_1_BLKSELA_i,
            BLKSELB => dpb_inst_1_BLKSELB_i,
            ADA => dpb_inst_1_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_1_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_2: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "010",
            BLK_SEL_1 => "010",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_2_douta(15 downto 0),
            DOB => dpb_inst_2_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_2_BLKSELA_i,
            BLKSELB => dpb_inst_2_BLKSELB_i,
            ADA => dpb_inst_2_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_2_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_3: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "011",
            BLK_SEL_1 => "011",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_3_douta(15 downto 0),
            DOB => dpb_inst_3_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_3_BLKSELA_i,
            BLKSELB => dpb_inst_3_BLKSELB_i,
            ADA => dpb_inst_3_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_3_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_4: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "100",
            BLK_SEL_1 => "100",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_4_douta(15 downto 0),
            DOB => dpb_inst_4_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_4_BLKSELA_i,
            BLKSELB => dpb_inst_4_BLKSELB_i,
            ADA => dpb_inst_4_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_4_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_5: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "101",
            BLK_SEL_1 => "101",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_5_douta(15 downto 0),
            DOB => dpb_inst_5_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_5_BLKSELA_i,
            BLKSELB => dpb_inst_5_BLKSELB_i,
            ADA => dpb_inst_5_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_5_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_6: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "110",
            BLK_SEL_1 => "110",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_6_douta(15 downto 0),
            DOB => dpb_inst_6_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_6_BLKSELA_i,
            BLKSELB => dpb_inst_6_BLKSELB_i,
            ADA => dpb_inst_6_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_6_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_7: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "111",
            BLK_SEL_1 => "111",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_7_douta(15 downto 0),
            DOB => dpb_inst_7_doutb(15 downto 0),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_7_BLKSELA_i,
            BLKSELB => dpb_inst_7_BLKSELB_i,
            ADA => dpb_inst_7_ADA_i,
            DIA => dina(15 downto 0),
            ADB => dpb_inst_7_ADB_i,
            DIB => dinb(15 downto 0)
        );

    dpb_inst_8: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"FCA403010281FD01000000001BD00001000100010001FF010000000000000100",
            INIT_RAM_01 => X"FCF700D0FEB40C070FF700F0FEB4FEF4000700E7FDC40007FEE40017FEC4FE04",
            INIT_RAM_02 => X"000005074187000040E7000040F702F60500418700004187000004F700A0FEB4",
            INIT_RAM_03 => X"010700F7F007000041070107FEB4F65F40070000F6E795F700004187000040E7",
            INIT_RAM_04 => X"00070000F11F00E70107010500F7001740C6000000174187000041C700004105",
            INIT_RAM_05 => X"000738C7000000070FF700F00017004738C7000002010081FE010000030102C1",
            INIT_RAM_06 => X"00170027004738C70000FEF4000502010081FE010000020101C10007FFF00080",
            INIT_RAM_07 => X"030102810211FD010000020101C10007000000E7FEF438C70000FE5F00070FF7",
            INIT_RAM_08 => X"00A0FE7404F700D0FE74FEF4FE84FEDF00F7FFF0FE84FEA4F41FFE04FCB4FCA4",
            INIT_RAM_09 => X"00F7FDC4FEC400E7FE7400E7FDC40007FEE40017FEC402F7FEC4FFF7FD8404F7",
            INIT_RAM_0A => X"FCB4FCA403010281FD0100000301028102C100070000F7DF00F700A0FE740007",
            INIT_RAM_0B => X"0600FEF40500FD07FEF400E70390FEF400E702F0FEF4FEF4000700F7FDC4FD84",
            INIT_RAM_0C => X"0080FC97FEF400E70460FEF400E70400FEF402C0FA97FEF400E70660FEF400E7",
            INIT_RAM_0D => X"FDC40007FCE40017FD84FCB4FCA4030102810211FD010000030102C10007FFF0",
            INIT_RAM_0E => X"0140FFF000F7FFF0FE84FEA4F09FFDC4FD840380FFF000F7FFF0FEC4FEA4F2DF",
            INIT_RAM_0F => X"FCC40010FCA4040102810211FC0100000301028102C1000700F7FE840047FEC4",
            INIT_RAM_10 => X"000700770017FEC406F7FEC4FFD7FE84FE040780001000F7FFF0FE84FEA4F55F",
            INIT_RAM_11 => X"FEC4BB9F0007FDC4FC04FCF40FF7FE440340001000F7FFF0FE44FEA4F11FFCC4",
            INIT_RAM_12 => X"FC04FCB4FCA4040102810211FC0100000401038103C100070000F99FFEF40017",
            INIT_RAM_13 => X"02F70030FC8402F70020FC841740001000F7FFF0FD84FCF40005E8DFFCC40020",
            INIT_RAM_14 => X"00C0FEF400400180FEF400A0FEF4003002C0FEF40080FEF4002004F70010FC84",
            INIT_RAM_15 => X"FFF0FD44FCA4DE5FFCC4000700170027FEC406F7FE04FEC4FE04FE040000FEF4",
            INIT_RAM_16 => X"F95FFEF40017FEC4FEF400E7FE4400070FF7FD44FEF40087FE440D00001000F7",
            INIT_RAM_17 => X"00F7FE840017FEC406F7FEC4FFF740F7FE04FD84FE040880002000F70000FE44",
            INIT_RAM_18 => X"0FF7FD4400F7FDC400F7FEC4FE440380001000F7FFF0FD44FCA4D4DFFCC40007",
            INIT_RAM_19 => X"FCA4030102810211FD0100000401038103C100070000F89FFEF40017FEC400E7",
            INIT_RAM_1A => X"0180FEF400300240FEF4004002F70070FD8402F70090FD8402F70080FD84FCB4",
            INIT_RAM_1B => X"C59FFDC4000700170027FE8406F7FE44FE84FE04FE040A40001000C0FEF40020",
            INIT_RAM_1C => X"FE84FEF400E7FEC400070FF7FE04FEF40087FEC40600001000F7FFF0FE04FEA4",
            INIT_RAM_1D => X"028102C10007000000074207000042E70000FEC48DDFF2C70000F95FFEF40017",
            INIT_RAM_1E => X"0017FEC487DFF347000002F7FDC4FEC4FE04FCA4030102810211FD0100000301",
            INIT_RAM_1F => X"0017004739470000FEF4000502010081FE0100000301028102C10000FDDFFEF4",
            INIT_RAM_20 => X"FE5F00070FF70017001700473947000000E7FEF439470000FE5F00070FF70017",
            INIT_RAM_21 => X"FCC4FCB4FCA40301029102810211FD010000020101C100070FF7000739470000",
            INIT_RAM_22 => X"0087FDC4F29F00070FF70107FDC4F3DF003000E7EFF73847000000C738470000",
            INIT_RAM_23 => X"EE1F0FF000F7FEC4FD4402F7FD84FEC4FE04F05F00070FF7FDC4F15F00070FF7",
            INIT_RAM_24 => X"02C10007000000E710073847000000C738470000FCDFFEF40017FEC400F40005",
            INIT_RAM_25 => X"2000EE9F007000022000EC8FF3870000020100810011FE010000030102410281",
            INIT_RAM_26 => X"014000074207000042E720000000E90FF507000002F706F701000007FEC4FEF4",
            INIT_RAM_27 => X"0000000739070000020100810011FE0100000201018101C10000E68FF5870000",
            INIT_RAM_28 => X"00E7FE0400473887000002070FF700170017000738870000FE0400E700403847",
            INIT_RAM_29 => X"FEC441C7000002E795F70000FEC4FE044007000040E7D40700000000FCDFFEF4",
            INIT_RAM_2A => X"FC070000CD5F01B0D84FFBC70000FC5FFEF40017FEC400E7F007000000F70017",
            INIT_RAM_2B => X"D34F01470000C99F01B0D48FFF870000CADF01B0D5CFFDC70000CC1F01B0D70F",
            INIT_RAM_2C => X"01B0CF8F06870000C5DF01B0D0CF04C70000C71F01B0D20F03070000C85F01B0",
            INIT_RAM_2D => X"C0DF01B0CBCF0A070000C21F01B0CD0F08470000C35F01B0CE4F03070000C49F",
            INIT_RAM_2E => X"000001070107FEC404E700F0FEC4FE04C94F0BC70000BF9F01B0CA8F03070000",
            INIT_RAM_2F => X"0000FEF4FFF0FE04FB9FFEF40017FEC400E70107010700C700F60017FEC441C7",
            INIT_RAM_30 => X"0400BF8F0D87000000E7FE84FEC402E703B0FE8406E703B0FEC4FE0440E74BA0",
            INIT_RAM_31 => X"FEC4BB8F0D8700000100BC8F0DC7000000F7FEC4FC57FE840300BE8F0DC70000",
            INIT_RAM_32 => X"0FF700F76A070001FE04FE04FE0400E70770FE84FEF40017FE84F85FFEF40017",
            INIT_RAM_33 => X"001700170007388700000000FC9FFEF40017FE0400F70530FE44FEA4C88F0207",
            INIT_RAM_34 => X"FEF400E7FE0400473887000002070FF700170017000738870000FE0404070FF7",
            INIT_RAM_35 => X"398700000800AC0F0E070000E99F00F70530FE44BFDF00070FF700F0FE04FCDF",
            INIT_RAM_36 => X"BDCF021001C0A80F10870000BF4F02A000070FF700170005E58F39870000C70F",
            INIT_RAM_37 => X"001739870000FE04FEF7053039870000C14F3987000008000000A68F0F070000",
            INIT_RAM_38 => X"002009C0FEA4E74F3987000000100007000700F71387000000270CF70090FD07",
            INIT_RAM_39 => X"3987000000700640FE0406C0FEA4E44F3987000000300840FEA4E5CF39870000",
            INIT_RAM_3A => X"0005FB4F39870000009002C0FEF40005FD0F3987000000800480FEF40005FECF",
            INIT_RAM_3B => X"10C700000340AA8F02A0028000F70010FE840007FE840000FEF400200100FEF4",
            INIT_RAM_3C => X"6E696F4C000000004F4FEA9F0000A78F0210918F1107000001C0A90F0720930F",
            INIT_RAM_3D => X"20646365646170757361702072756E67206461760000544F000A6174646E6573",
            INIT_RAM_3E => X"00000000303037787461726F6D20697475676E6F4147206F72656F6C6F626761",
            INIT_RAM_3F => X"2E5F20200000292020207C20204F202020200000205C20207C2E5F5C20202020"
        )
        port map (
            DOA => dpb_inst_8_douta(31 downto 16),
            DOB => dpb_inst_8_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_8_BLKSELA_i,
            BLKSELB => dpb_inst_8_BLKSELB_i,
            ADA => dpb_inst_8_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_8_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_9: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "001",
            BLK_SEL_1 => "001",
            INIT_RAM_00 => X"2020202020207C2000002E2D2D2D28282D2D28202E200000202820207C205420",
            INIT_RAM_01 => X"7C2020203330303220207C2000007C72616F6F6F434F676E7C2000007C202020",
            INIT_RAM_02 => X"602000007C20532072666F6F6F747C2000007C207965796E737350207C200000",
            INIT_RAM_03 => X"65736C702052524500003A677669655200000000000A602D2D2D2D2D2D2D2D2D",
            INIT_RAM_04 => X"0000000000000A74657273617020726F65206261766F726E00000000000A7365",
            INIT_RAM_05 => X"FFFF000000000002010100520000000000000000000000000000000000000000",
            INIT_RAM_06 => X"00000000020D78004401200E0000FFFF00000000000044C803004401300E0000",
            INIT_RAM_07 => X"0D44C1A0080C8801300E0000FFFF0000000000000D4402004401200E0000FFFF",
            INIT_RAM_08 => X"8801300E0000FFFF0000000000000D4402004401300E0000FFFF000000000000",
            INIT_RAM_09 => X"0000000000000D44C1A4080C8801400E0000FFFF0000000000000D44C174080C",
            INIT_RAM_0A => X"0100080C8801300E0000FFFF00000000000044C801AC080C8801400E0000FFFF",
            INIT_RAM_0B => X"200E0000FFFF00000000020D44C1080C8801300E0000FFFF00000000000044C8",
            INIT_RAM_0C => X"000000000D44C844020044038801300E0000FFFF0000000000000D4402004401",
            INIT_RAM_0D => X"080C8801200E0000FFFF0000000000000D44C174080C8801200E0000FFFF0000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000F070F060F040F030F0000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_9_douta(31 downto 16),
            DOB => dpb_inst_9_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_9_BLKSELA_i,
            BLKSELB => dpb_inst_9_BLKSELB_i,
            ADA => dpb_inst_9_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_9_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_10: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "010",
            BLK_SEL_1 => "010",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_10_douta(31 downto 16),
            DOB => dpb_inst_10_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_10_BLKSELA_i,
            BLKSELB => dpb_inst_10_BLKSELB_i,
            ADA => dpb_inst_10_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_10_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_11: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "011",
            BLK_SEL_1 => "011",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_11_douta(31 downto 16),
            DOB => dpb_inst_11_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_11_BLKSELA_i,
            BLKSELB => dpb_inst_11_BLKSELB_i,
            ADA => dpb_inst_11_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_11_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_12: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "100",
            BLK_SEL_1 => "100",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_12_douta(31 downto 16),
            DOB => dpb_inst_12_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_12_BLKSELA_i,
            BLKSELB => dpb_inst_12_BLKSELB_i,
            ADA => dpb_inst_12_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_12_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_13: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "101",
            BLK_SEL_1 => "101",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_13_douta(31 downto 16),
            DOB => dpb_inst_13_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_13_BLKSELA_i,
            BLKSELB => dpb_inst_13_BLKSELB_i,
            ADA => dpb_inst_13_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_13_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_14: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "110",
            BLK_SEL_1 => "110",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_14_douta(31 downto 16),
            DOB => dpb_inst_14_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_14_BLKSELA_i,
            BLKSELB => dpb_inst_14_BLKSELB_i,
            ADA => dpb_inst_14_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_14_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dpb_inst_15: DPB
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 16,
            BIT_WIDTH_1 => 16,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "111",
            BLK_SEL_1 => "111",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DOA => dpb_inst_15_douta(31 downto 16),
            DOB => dpb_inst_15_doutb(31 downto 16),
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpb_inst_15_BLKSELA_i,
            BLKSELB => dpb_inst_15_BLKSELB_i,
            ADA => dpb_inst_15_ADA_i,
            DIA => dina(31 downto 16),
            ADB => dpb_inst_15_ADB_i,
            DIB => dinb(31 downto 16)
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ada(12),
            CLK => clka,
            CE => cea_w
        );

    dff_inst_1: DFFE
        port map (
            Q => dff_q_1,
            D => ada(11),
            CLK => clka,
            CE => cea_w
        );

    dff_inst_2: DFFE
        port map (
            Q => dff_q_2,
            D => ada(10),
            CLK => clka,
            CE => cea_w
        );

    dff_inst_3: DFFE
        port map (
            Q => dff_q_3,
            D => adb(12),
            CLK => clkb,
            CE => ceb_w
        );

    dff_inst_4: DFFE
        port map (
            Q => dff_q_4,
            D => adb(11),
            CLK => clkb,
            CE => ceb_w
        );

    dff_inst_5: DFFE
        port map (
            Q => dff_q_5,
            D => adb(10),
            CLK => clkb,
            CE => ceb_w
        );

    mux_inst_0: MUX2
        port map (
            O => mux_o_0,
            I0 => dpb_inst_0_douta(0),
            I1 => dpb_inst_1_douta(0),
            S0 => dff_q_2
        );

    mux_inst_1: MUX2
        port map (
            O => mux_o_1,
            I0 => dpb_inst_2_douta(0),
            I1 => dpb_inst_3_douta(0),
            S0 => dff_q_2
        );

    mux_inst_2: MUX2
        port map (
            O => mux_o_2,
            I0 => dpb_inst_4_douta(0),
            I1 => dpb_inst_5_douta(0),
            S0 => dff_q_2
        );

    mux_inst_3: MUX2
        port map (
            O => mux_o_3,
            I0 => dpb_inst_6_douta(0),
            I1 => dpb_inst_7_douta(0),
            S0 => dff_q_2
        );

    mux_inst_4: MUX2
        port map (
            O => mux_o_4,
            I0 => mux_o_0,
            I1 => mux_o_1,
            S0 => dff_q_1
        );

    mux_inst_5: MUX2
        port map (
            O => mux_o_5,
            I0 => mux_o_2,
            I1 => mux_o_3,
            S0 => dff_q_1
        );

    mux_inst_6: MUX2
        port map (
            O => douta(0),
            I0 => mux_o_4,
            I1 => mux_o_5,
            S0 => dff_q_0
        );

    mux_inst_7: MUX2
        port map (
            O => mux_o_7,
            I0 => dpb_inst_0_douta(1),
            I1 => dpb_inst_1_douta(1),
            S0 => dff_q_2
        );

    mux_inst_8: MUX2
        port map (
            O => mux_o_8,
            I0 => dpb_inst_2_douta(1),
            I1 => dpb_inst_3_douta(1),
            S0 => dff_q_2
        );

    mux_inst_9: MUX2
        port map (
            O => mux_o_9,
            I0 => dpb_inst_4_douta(1),
            I1 => dpb_inst_5_douta(1),
            S0 => dff_q_2
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => dpb_inst_6_douta(1),
            I1 => dpb_inst_7_douta(1),
            S0 => dff_q_2
        );

    mux_inst_11: MUX2
        port map (
            O => mux_o_11,
            I0 => mux_o_7,
            I1 => mux_o_8,
            S0 => dff_q_1
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => mux_o_9,
            I1 => mux_o_10,
            S0 => dff_q_1
        );

    mux_inst_13: MUX2
        port map (
            O => douta(1),
            I0 => mux_o_11,
            I1 => mux_o_12,
            S0 => dff_q_0
        );

    mux_inst_14: MUX2
        port map (
            O => mux_o_14,
            I0 => dpb_inst_0_douta(2),
            I1 => dpb_inst_1_douta(2),
            S0 => dff_q_2
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => dpb_inst_2_douta(2),
            I1 => dpb_inst_3_douta(2),
            S0 => dff_q_2
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => dpb_inst_4_douta(2),
            I1 => dpb_inst_5_douta(2),
            S0 => dff_q_2
        );

    mux_inst_17: MUX2
        port map (
            O => mux_o_17,
            I0 => dpb_inst_6_douta(2),
            I1 => dpb_inst_7_douta(2),
            S0 => dff_q_2
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => mux_o_14,
            I1 => mux_o_15,
            S0 => dff_q_1
        );

    mux_inst_19: MUX2
        port map (
            O => mux_o_19,
            I0 => mux_o_16,
            I1 => mux_o_17,
            S0 => dff_q_1
        );

    mux_inst_20: MUX2
        port map (
            O => douta(2),
            I0 => mux_o_18,
            I1 => mux_o_19,
            S0 => dff_q_0
        );

    mux_inst_21: MUX2
        port map (
            O => mux_o_21,
            I0 => dpb_inst_0_douta(3),
            I1 => dpb_inst_1_douta(3),
            S0 => dff_q_2
        );

    mux_inst_22: MUX2
        port map (
            O => mux_o_22,
            I0 => dpb_inst_2_douta(3),
            I1 => dpb_inst_3_douta(3),
            S0 => dff_q_2
        );

    mux_inst_23: MUX2
        port map (
            O => mux_o_23,
            I0 => dpb_inst_4_douta(3),
            I1 => dpb_inst_5_douta(3),
            S0 => dff_q_2
        );

    mux_inst_24: MUX2
        port map (
            O => mux_o_24,
            I0 => dpb_inst_6_douta(3),
            I1 => dpb_inst_7_douta(3),
            S0 => dff_q_2
        );

    mux_inst_25: MUX2
        port map (
            O => mux_o_25,
            I0 => mux_o_21,
            I1 => mux_o_22,
            S0 => dff_q_1
        );

    mux_inst_26: MUX2
        port map (
            O => mux_o_26,
            I0 => mux_o_23,
            I1 => mux_o_24,
            S0 => dff_q_1
        );

    mux_inst_27: MUX2
        port map (
            O => douta(3),
            I0 => mux_o_25,
            I1 => mux_o_26,
            S0 => dff_q_0
        );

    mux_inst_28: MUX2
        port map (
            O => mux_o_28,
            I0 => dpb_inst_0_douta(4),
            I1 => dpb_inst_1_douta(4),
            S0 => dff_q_2
        );

    mux_inst_29: MUX2
        port map (
            O => mux_o_29,
            I0 => dpb_inst_2_douta(4),
            I1 => dpb_inst_3_douta(4),
            S0 => dff_q_2
        );

    mux_inst_30: MUX2
        port map (
            O => mux_o_30,
            I0 => dpb_inst_4_douta(4),
            I1 => dpb_inst_5_douta(4),
            S0 => dff_q_2
        );

    mux_inst_31: MUX2
        port map (
            O => mux_o_31,
            I0 => dpb_inst_6_douta(4),
            I1 => dpb_inst_7_douta(4),
            S0 => dff_q_2
        );

    mux_inst_32: MUX2
        port map (
            O => mux_o_32,
            I0 => mux_o_28,
            I1 => mux_o_29,
            S0 => dff_q_1
        );

    mux_inst_33: MUX2
        port map (
            O => mux_o_33,
            I0 => mux_o_30,
            I1 => mux_o_31,
            S0 => dff_q_1
        );

    mux_inst_34: MUX2
        port map (
            O => douta(4),
            I0 => mux_o_32,
            I1 => mux_o_33,
            S0 => dff_q_0
        );

    mux_inst_35: MUX2
        port map (
            O => mux_o_35,
            I0 => dpb_inst_0_douta(5),
            I1 => dpb_inst_1_douta(5),
            S0 => dff_q_2
        );

    mux_inst_36: MUX2
        port map (
            O => mux_o_36,
            I0 => dpb_inst_2_douta(5),
            I1 => dpb_inst_3_douta(5),
            S0 => dff_q_2
        );

    mux_inst_37: MUX2
        port map (
            O => mux_o_37,
            I0 => dpb_inst_4_douta(5),
            I1 => dpb_inst_5_douta(5),
            S0 => dff_q_2
        );

    mux_inst_38: MUX2
        port map (
            O => mux_o_38,
            I0 => dpb_inst_6_douta(5),
            I1 => dpb_inst_7_douta(5),
            S0 => dff_q_2
        );

    mux_inst_39: MUX2
        port map (
            O => mux_o_39,
            I0 => mux_o_35,
            I1 => mux_o_36,
            S0 => dff_q_1
        );

    mux_inst_40: MUX2
        port map (
            O => mux_o_40,
            I0 => mux_o_37,
            I1 => mux_o_38,
            S0 => dff_q_1
        );

    mux_inst_41: MUX2
        port map (
            O => douta(5),
            I0 => mux_o_39,
            I1 => mux_o_40,
            S0 => dff_q_0
        );

    mux_inst_42: MUX2
        port map (
            O => mux_o_42,
            I0 => dpb_inst_0_douta(6),
            I1 => dpb_inst_1_douta(6),
            S0 => dff_q_2
        );

    mux_inst_43: MUX2
        port map (
            O => mux_o_43,
            I0 => dpb_inst_2_douta(6),
            I1 => dpb_inst_3_douta(6),
            S0 => dff_q_2
        );

    mux_inst_44: MUX2
        port map (
            O => mux_o_44,
            I0 => dpb_inst_4_douta(6),
            I1 => dpb_inst_5_douta(6),
            S0 => dff_q_2
        );

    mux_inst_45: MUX2
        port map (
            O => mux_o_45,
            I0 => dpb_inst_6_douta(6),
            I1 => dpb_inst_7_douta(6),
            S0 => dff_q_2
        );

    mux_inst_46: MUX2
        port map (
            O => mux_o_46,
            I0 => mux_o_42,
            I1 => mux_o_43,
            S0 => dff_q_1
        );

    mux_inst_47: MUX2
        port map (
            O => mux_o_47,
            I0 => mux_o_44,
            I1 => mux_o_45,
            S0 => dff_q_1
        );

    mux_inst_48: MUX2
        port map (
            O => douta(6),
            I0 => mux_o_46,
            I1 => mux_o_47,
            S0 => dff_q_0
        );

    mux_inst_49: MUX2
        port map (
            O => mux_o_49,
            I0 => dpb_inst_0_douta(7),
            I1 => dpb_inst_1_douta(7),
            S0 => dff_q_2
        );

    mux_inst_50: MUX2
        port map (
            O => mux_o_50,
            I0 => dpb_inst_2_douta(7),
            I1 => dpb_inst_3_douta(7),
            S0 => dff_q_2
        );

    mux_inst_51: MUX2
        port map (
            O => mux_o_51,
            I0 => dpb_inst_4_douta(7),
            I1 => dpb_inst_5_douta(7),
            S0 => dff_q_2
        );

    mux_inst_52: MUX2
        port map (
            O => mux_o_52,
            I0 => dpb_inst_6_douta(7),
            I1 => dpb_inst_7_douta(7),
            S0 => dff_q_2
        );

    mux_inst_53: MUX2
        port map (
            O => mux_o_53,
            I0 => mux_o_49,
            I1 => mux_o_50,
            S0 => dff_q_1
        );

    mux_inst_54: MUX2
        port map (
            O => mux_o_54,
            I0 => mux_o_51,
            I1 => mux_o_52,
            S0 => dff_q_1
        );

    mux_inst_55: MUX2
        port map (
            O => douta(7),
            I0 => mux_o_53,
            I1 => mux_o_54,
            S0 => dff_q_0
        );

    mux_inst_56: MUX2
        port map (
            O => mux_o_56,
            I0 => dpb_inst_0_douta(8),
            I1 => dpb_inst_1_douta(8),
            S0 => dff_q_2
        );

    mux_inst_57: MUX2
        port map (
            O => mux_o_57,
            I0 => dpb_inst_2_douta(8),
            I1 => dpb_inst_3_douta(8),
            S0 => dff_q_2
        );

    mux_inst_58: MUX2
        port map (
            O => mux_o_58,
            I0 => dpb_inst_4_douta(8),
            I1 => dpb_inst_5_douta(8),
            S0 => dff_q_2
        );

    mux_inst_59: MUX2
        port map (
            O => mux_o_59,
            I0 => dpb_inst_6_douta(8),
            I1 => dpb_inst_7_douta(8),
            S0 => dff_q_2
        );

    mux_inst_60: MUX2
        port map (
            O => mux_o_60,
            I0 => mux_o_56,
            I1 => mux_o_57,
            S0 => dff_q_1
        );

    mux_inst_61: MUX2
        port map (
            O => mux_o_61,
            I0 => mux_o_58,
            I1 => mux_o_59,
            S0 => dff_q_1
        );

    mux_inst_62: MUX2
        port map (
            O => douta(8),
            I0 => mux_o_60,
            I1 => mux_o_61,
            S0 => dff_q_0
        );

    mux_inst_63: MUX2
        port map (
            O => mux_o_63,
            I0 => dpb_inst_0_douta(9),
            I1 => dpb_inst_1_douta(9),
            S0 => dff_q_2
        );

    mux_inst_64: MUX2
        port map (
            O => mux_o_64,
            I0 => dpb_inst_2_douta(9),
            I1 => dpb_inst_3_douta(9),
            S0 => dff_q_2
        );

    mux_inst_65: MUX2
        port map (
            O => mux_o_65,
            I0 => dpb_inst_4_douta(9),
            I1 => dpb_inst_5_douta(9),
            S0 => dff_q_2
        );

    mux_inst_66: MUX2
        port map (
            O => mux_o_66,
            I0 => dpb_inst_6_douta(9),
            I1 => dpb_inst_7_douta(9),
            S0 => dff_q_2
        );

    mux_inst_67: MUX2
        port map (
            O => mux_o_67,
            I0 => mux_o_63,
            I1 => mux_o_64,
            S0 => dff_q_1
        );

    mux_inst_68: MUX2
        port map (
            O => mux_o_68,
            I0 => mux_o_65,
            I1 => mux_o_66,
            S0 => dff_q_1
        );

    mux_inst_69: MUX2
        port map (
            O => douta(9),
            I0 => mux_o_67,
            I1 => mux_o_68,
            S0 => dff_q_0
        );

    mux_inst_70: MUX2
        port map (
            O => mux_o_70,
            I0 => dpb_inst_0_douta(10),
            I1 => dpb_inst_1_douta(10),
            S0 => dff_q_2
        );

    mux_inst_71: MUX2
        port map (
            O => mux_o_71,
            I0 => dpb_inst_2_douta(10),
            I1 => dpb_inst_3_douta(10),
            S0 => dff_q_2
        );

    mux_inst_72: MUX2
        port map (
            O => mux_o_72,
            I0 => dpb_inst_4_douta(10),
            I1 => dpb_inst_5_douta(10),
            S0 => dff_q_2
        );

    mux_inst_73: MUX2
        port map (
            O => mux_o_73,
            I0 => dpb_inst_6_douta(10),
            I1 => dpb_inst_7_douta(10),
            S0 => dff_q_2
        );

    mux_inst_74: MUX2
        port map (
            O => mux_o_74,
            I0 => mux_o_70,
            I1 => mux_o_71,
            S0 => dff_q_1
        );

    mux_inst_75: MUX2
        port map (
            O => mux_o_75,
            I0 => mux_o_72,
            I1 => mux_o_73,
            S0 => dff_q_1
        );

    mux_inst_76: MUX2
        port map (
            O => douta(10),
            I0 => mux_o_74,
            I1 => mux_o_75,
            S0 => dff_q_0
        );

    mux_inst_77: MUX2
        port map (
            O => mux_o_77,
            I0 => dpb_inst_0_douta(11),
            I1 => dpb_inst_1_douta(11),
            S0 => dff_q_2
        );

    mux_inst_78: MUX2
        port map (
            O => mux_o_78,
            I0 => dpb_inst_2_douta(11),
            I1 => dpb_inst_3_douta(11),
            S0 => dff_q_2
        );

    mux_inst_79: MUX2
        port map (
            O => mux_o_79,
            I0 => dpb_inst_4_douta(11),
            I1 => dpb_inst_5_douta(11),
            S0 => dff_q_2
        );

    mux_inst_80: MUX2
        port map (
            O => mux_o_80,
            I0 => dpb_inst_6_douta(11),
            I1 => dpb_inst_7_douta(11),
            S0 => dff_q_2
        );

    mux_inst_81: MUX2
        port map (
            O => mux_o_81,
            I0 => mux_o_77,
            I1 => mux_o_78,
            S0 => dff_q_1
        );

    mux_inst_82: MUX2
        port map (
            O => mux_o_82,
            I0 => mux_o_79,
            I1 => mux_o_80,
            S0 => dff_q_1
        );

    mux_inst_83: MUX2
        port map (
            O => douta(11),
            I0 => mux_o_81,
            I1 => mux_o_82,
            S0 => dff_q_0
        );

    mux_inst_84: MUX2
        port map (
            O => mux_o_84,
            I0 => dpb_inst_0_douta(12),
            I1 => dpb_inst_1_douta(12),
            S0 => dff_q_2
        );

    mux_inst_85: MUX2
        port map (
            O => mux_o_85,
            I0 => dpb_inst_2_douta(12),
            I1 => dpb_inst_3_douta(12),
            S0 => dff_q_2
        );

    mux_inst_86: MUX2
        port map (
            O => mux_o_86,
            I0 => dpb_inst_4_douta(12),
            I1 => dpb_inst_5_douta(12),
            S0 => dff_q_2
        );

    mux_inst_87: MUX2
        port map (
            O => mux_o_87,
            I0 => dpb_inst_6_douta(12),
            I1 => dpb_inst_7_douta(12),
            S0 => dff_q_2
        );

    mux_inst_88: MUX2
        port map (
            O => mux_o_88,
            I0 => mux_o_84,
            I1 => mux_o_85,
            S0 => dff_q_1
        );

    mux_inst_89: MUX2
        port map (
            O => mux_o_89,
            I0 => mux_o_86,
            I1 => mux_o_87,
            S0 => dff_q_1
        );

    mux_inst_90: MUX2
        port map (
            O => douta(12),
            I0 => mux_o_88,
            I1 => mux_o_89,
            S0 => dff_q_0
        );

    mux_inst_91: MUX2
        port map (
            O => mux_o_91,
            I0 => dpb_inst_0_douta(13),
            I1 => dpb_inst_1_douta(13),
            S0 => dff_q_2
        );

    mux_inst_92: MUX2
        port map (
            O => mux_o_92,
            I0 => dpb_inst_2_douta(13),
            I1 => dpb_inst_3_douta(13),
            S0 => dff_q_2
        );

    mux_inst_93: MUX2
        port map (
            O => mux_o_93,
            I0 => dpb_inst_4_douta(13),
            I1 => dpb_inst_5_douta(13),
            S0 => dff_q_2
        );

    mux_inst_94: MUX2
        port map (
            O => mux_o_94,
            I0 => dpb_inst_6_douta(13),
            I1 => dpb_inst_7_douta(13),
            S0 => dff_q_2
        );

    mux_inst_95: MUX2
        port map (
            O => mux_o_95,
            I0 => mux_o_91,
            I1 => mux_o_92,
            S0 => dff_q_1
        );

    mux_inst_96: MUX2
        port map (
            O => mux_o_96,
            I0 => mux_o_93,
            I1 => mux_o_94,
            S0 => dff_q_1
        );

    mux_inst_97: MUX2
        port map (
            O => douta(13),
            I0 => mux_o_95,
            I1 => mux_o_96,
            S0 => dff_q_0
        );

    mux_inst_98: MUX2
        port map (
            O => mux_o_98,
            I0 => dpb_inst_0_douta(14),
            I1 => dpb_inst_1_douta(14),
            S0 => dff_q_2
        );

    mux_inst_99: MUX2
        port map (
            O => mux_o_99,
            I0 => dpb_inst_2_douta(14),
            I1 => dpb_inst_3_douta(14),
            S0 => dff_q_2
        );

    mux_inst_100: MUX2
        port map (
            O => mux_o_100,
            I0 => dpb_inst_4_douta(14),
            I1 => dpb_inst_5_douta(14),
            S0 => dff_q_2
        );

    mux_inst_101: MUX2
        port map (
            O => mux_o_101,
            I0 => dpb_inst_6_douta(14),
            I1 => dpb_inst_7_douta(14),
            S0 => dff_q_2
        );

    mux_inst_102: MUX2
        port map (
            O => mux_o_102,
            I0 => mux_o_98,
            I1 => mux_o_99,
            S0 => dff_q_1
        );

    mux_inst_103: MUX2
        port map (
            O => mux_o_103,
            I0 => mux_o_100,
            I1 => mux_o_101,
            S0 => dff_q_1
        );

    mux_inst_104: MUX2
        port map (
            O => douta(14),
            I0 => mux_o_102,
            I1 => mux_o_103,
            S0 => dff_q_0
        );

    mux_inst_105: MUX2
        port map (
            O => mux_o_105,
            I0 => dpb_inst_0_douta(15),
            I1 => dpb_inst_1_douta(15),
            S0 => dff_q_2
        );

    mux_inst_106: MUX2
        port map (
            O => mux_o_106,
            I0 => dpb_inst_2_douta(15),
            I1 => dpb_inst_3_douta(15),
            S0 => dff_q_2
        );

    mux_inst_107: MUX2
        port map (
            O => mux_o_107,
            I0 => dpb_inst_4_douta(15),
            I1 => dpb_inst_5_douta(15),
            S0 => dff_q_2
        );

    mux_inst_108: MUX2
        port map (
            O => mux_o_108,
            I0 => dpb_inst_6_douta(15),
            I1 => dpb_inst_7_douta(15),
            S0 => dff_q_2
        );

    mux_inst_109: MUX2
        port map (
            O => mux_o_109,
            I0 => mux_o_105,
            I1 => mux_o_106,
            S0 => dff_q_1
        );

    mux_inst_110: MUX2
        port map (
            O => mux_o_110,
            I0 => mux_o_107,
            I1 => mux_o_108,
            S0 => dff_q_1
        );

    mux_inst_111: MUX2
        port map (
            O => douta(15),
            I0 => mux_o_109,
            I1 => mux_o_110,
            S0 => dff_q_0
        );

    mux_inst_112: MUX2
        port map (
            O => mux_o_112,
            I0 => dpb_inst_8_douta(16),
            I1 => dpb_inst_9_douta(16),
            S0 => dff_q_2
        );

    mux_inst_113: MUX2
        port map (
            O => mux_o_113,
            I0 => dpb_inst_10_douta(16),
            I1 => dpb_inst_11_douta(16),
            S0 => dff_q_2
        );

    mux_inst_114: MUX2
        port map (
            O => mux_o_114,
            I0 => dpb_inst_12_douta(16),
            I1 => dpb_inst_13_douta(16),
            S0 => dff_q_2
        );

    mux_inst_115: MUX2
        port map (
            O => mux_o_115,
            I0 => dpb_inst_14_douta(16),
            I1 => dpb_inst_15_douta(16),
            S0 => dff_q_2
        );

    mux_inst_116: MUX2
        port map (
            O => mux_o_116,
            I0 => mux_o_112,
            I1 => mux_o_113,
            S0 => dff_q_1
        );

    mux_inst_117: MUX2
        port map (
            O => mux_o_117,
            I0 => mux_o_114,
            I1 => mux_o_115,
            S0 => dff_q_1
        );

    mux_inst_118: MUX2
        port map (
            O => douta(16),
            I0 => mux_o_116,
            I1 => mux_o_117,
            S0 => dff_q_0
        );

    mux_inst_119: MUX2
        port map (
            O => mux_o_119,
            I0 => dpb_inst_8_douta(17),
            I1 => dpb_inst_9_douta(17),
            S0 => dff_q_2
        );

    mux_inst_120: MUX2
        port map (
            O => mux_o_120,
            I0 => dpb_inst_10_douta(17),
            I1 => dpb_inst_11_douta(17),
            S0 => dff_q_2
        );

    mux_inst_121: MUX2
        port map (
            O => mux_o_121,
            I0 => dpb_inst_12_douta(17),
            I1 => dpb_inst_13_douta(17),
            S0 => dff_q_2
        );

    mux_inst_122: MUX2
        port map (
            O => mux_o_122,
            I0 => dpb_inst_14_douta(17),
            I1 => dpb_inst_15_douta(17),
            S0 => dff_q_2
        );

    mux_inst_123: MUX2
        port map (
            O => mux_o_123,
            I0 => mux_o_119,
            I1 => mux_o_120,
            S0 => dff_q_1
        );

    mux_inst_124: MUX2
        port map (
            O => mux_o_124,
            I0 => mux_o_121,
            I1 => mux_o_122,
            S0 => dff_q_1
        );

    mux_inst_125: MUX2
        port map (
            O => douta(17),
            I0 => mux_o_123,
            I1 => mux_o_124,
            S0 => dff_q_0
        );

    mux_inst_126: MUX2
        port map (
            O => mux_o_126,
            I0 => dpb_inst_8_douta(18),
            I1 => dpb_inst_9_douta(18),
            S0 => dff_q_2
        );

    mux_inst_127: MUX2
        port map (
            O => mux_o_127,
            I0 => dpb_inst_10_douta(18),
            I1 => dpb_inst_11_douta(18),
            S0 => dff_q_2
        );

    mux_inst_128: MUX2
        port map (
            O => mux_o_128,
            I0 => dpb_inst_12_douta(18),
            I1 => dpb_inst_13_douta(18),
            S0 => dff_q_2
        );

    mux_inst_129: MUX2
        port map (
            O => mux_o_129,
            I0 => dpb_inst_14_douta(18),
            I1 => dpb_inst_15_douta(18),
            S0 => dff_q_2
        );

    mux_inst_130: MUX2
        port map (
            O => mux_o_130,
            I0 => mux_o_126,
            I1 => mux_o_127,
            S0 => dff_q_1
        );

    mux_inst_131: MUX2
        port map (
            O => mux_o_131,
            I0 => mux_o_128,
            I1 => mux_o_129,
            S0 => dff_q_1
        );

    mux_inst_132: MUX2
        port map (
            O => douta(18),
            I0 => mux_o_130,
            I1 => mux_o_131,
            S0 => dff_q_0
        );

    mux_inst_133: MUX2
        port map (
            O => mux_o_133,
            I0 => dpb_inst_8_douta(19),
            I1 => dpb_inst_9_douta(19),
            S0 => dff_q_2
        );

    mux_inst_134: MUX2
        port map (
            O => mux_o_134,
            I0 => dpb_inst_10_douta(19),
            I1 => dpb_inst_11_douta(19),
            S0 => dff_q_2
        );

    mux_inst_135: MUX2
        port map (
            O => mux_o_135,
            I0 => dpb_inst_12_douta(19),
            I1 => dpb_inst_13_douta(19),
            S0 => dff_q_2
        );

    mux_inst_136: MUX2
        port map (
            O => mux_o_136,
            I0 => dpb_inst_14_douta(19),
            I1 => dpb_inst_15_douta(19),
            S0 => dff_q_2
        );

    mux_inst_137: MUX2
        port map (
            O => mux_o_137,
            I0 => mux_o_133,
            I1 => mux_o_134,
            S0 => dff_q_1
        );

    mux_inst_138: MUX2
        port map (
            O => mux_o_138,
            I0 => mux_o_135,
            I1 => mux_o_136,
            S0 => dff_q_1
        );

    mux_inst_139: MUX2
        port map (
            O => douta(19),
            I0 => mux_o_137,
            I1 => mux_o_138,
            S0 => dff_q_0
        );

    mux_inst_140: MUX2
        port map (
            O => mux_o_140,
            I0 => dpb_inst_8_douta(20),
            I1 => dpb_inst_9_douta(20),
            S0 => dff_q_2
        );

    mux_inst_141: MUX2
        port map (
            O => mux_o_141,
            I0 => dpb_inst_10_douta(20),
            I1 => dpb_inst_11_douta(20),
            S0 => dff_q_2
        );

    mux_inst_142: MUX2
        port map (
            O => mux_o_142,
            I0 => dpb_inst_12_douta(20),
            I1 => dpb_inst_13_douta(20),
            S0 => dff_q_2
        );

    mux_inst_143: MUX2
        port map (
            O => mux_o_143,
            I0 => dpb_inst_14_douta(20),
            I1 => dpb_inst_15_douta(20),
            S0 => dff_q_2
        );

    mux_inst_144: MUX2
        port map (
            O => mux_o_144,
            I0 => mux_o_140,
            I1 => mux_o_141,
            S0 => dff_q_1
        );

    mux_inst_145: MUX2
        port map (
            O => mux_o_145,
            I0 => mux_o_142,
            I1 => mux_o_143,
            S0 => dff_q_1
        );

    mux_inst_146: MUX2
        port map (
            O => douta(20),
            I0 => mux_o_144,
            I1 => mux_o_145,
            S0 => dff_q_0
        );

    mux_inst_147: MUX2
        port map (
            O => mux_o_147,
            I0 => dpb_inst_8_douta(21),
            I1 => dpb_inst_9_douta(21),
            S0 => dff_q_2
        );

    mux_inst_148: MUX2
        port map (
            O => mux_o_148,
            I0 => dpb_inst_10_douta(21),
            I1 => dpb_inst_11_douta(21),
            S0 => dff_q_2
        );

    mux_inst_149: MUX2
        port map (
            O => mux_o_149,
            I0 => dpb_inst_12_douta(21),
            I1 => dpb_inst_13_douta(21),
            S0 => dff_q_2
        );

    mux_inst_150: MUX2
        port map (
            O => mux_o_150,
            I0 => dpb_inst_14_douta(21),
            I1 => dpb_inst_15_douta(21),
            S0 => dff_q_2
        );

    mux_inst_151: MUX2
        port map (
            O => mux_o_151,
            I0 => mux_o_147,
            I1 => mux_o_148,
            S0 => dff_q_1
        );

    mux_inst_152: MUX2
        port map (
            O => mux_o_152,
            I0 => mux_o_149,
            I1 => mux_o_150,
            S0 => dff_q_1
        );

    mux_inst_153: MUX2
        port map (
            O => douta(21),
            I0 => mux_o_151,
            I1 => mux_o_152,
            S0 => dff_q_0
        );

    mux_inst_154: MUX2
        port map (
            O => mux_o_154,
            I0 => dpb_inst_8_douta(22),
            I1 => dpb_inst_9_douta(22),
            S0 => dff_q_2
        );

    mux_inst_155: MUX2
        port map (
            O => mux_o_155,
            I0 => dpb_inst_10_douta(22),
            I1 => dpb_inst_11_douta(22),
            S0 => dff_q_2
        );

    mux_inst_156: MUX2
        port map (
            O => mux_o_156,
            I0 => dpb_inst_12_douta(22),
            I1 => dpb_inst_13_douta(22),
            S0 => dff_q_2
        );

    mux_inst_157: MUX2
        port map (
            O => mux_o_157,
            I0 => dpb_inst_14_douta(22),
            I1 => dpb_inst_15_douta(22),
            S0 => dff_q_2
        );

    mux_inst_158: MUX2
        port map (
            O => mux_o_158,
            I0 => mux_o_154,
            I1 => mux_o_155,
            S0 => dff_q_1
        );

    mux_inst_159: MUX2
        port map (
            O => mux_o_159,
            I0 => mux_o_156,
            I1 => mux_o_157,
            S0 => dff_q_1
        );

    mux_inst_160: MUX2
        port map (
            O => douta(22),
            I0 => mux_o_158,
            I1 => mux_o_159,
            S0 => dff_q_0
        );

    mux_inst_161: MUX2
        port map (
            O => mux_o_161,
            I0 => dpb_inst_8_douta(23),
            I1 => dpb_inst_9_douta(23),
            S0 => dff_q_2
        );

    mux_inst_162: MUX2
        port map (
            O => mux_o_162,
            I0 => dpb_inst_10_douta(23),
            I1 => dpb_inst_11_douta(23),
            S0 => dff_q_2
        );

    mux_inst_163: MUX2
        port map (
            O => mux_o_163,
            I0 => dpb_inst_12_douta(23),
            I1 => dpb_inst_13_douta(23),
            S0 => dff_q_2
        );

    mux_inst_164: MUX2
        port map (
            O => mux_o_164,
            I0 => dpb_inst_14_douta(23),
            I1 => dpb_inst_15_douta(23),
            S0 => dff_q_2
        );

    mux_inst_165: MUX2
        port map (
            O => mux_o_165,
            I0 => mux_o_161,
            I1 => mux_o_162,
            S0 => dff_q_1
        );

    mux_inst_166: MUX2
        port map (
            O => mux_o_166,
            I0 => mux_o_163,
            I1 => mux_o_164,
            S0 => dff_q_1
        );

    mux_inst_167: MUX2
        port map (
            O => douta(23),
            I0 => mux_o_165,
            I1 => mux_o_166,
            S0 => dff_q_0
        );

    mux_inst_168: MUX2
        port map (
            O => mux_o_168,
            I0 => dpb_inst_8_douta(24),
            I1 => dpb_inst_9_douta(24),
            S0 => dff_q_2
        );

    mux_inst_169: MUX2
        port map (
            O => mux_o_169,
            I0 => dpb_inst_10_douta(24),
            I1 => dpb_inst_11_douta(24),
            S0 => dff_q_2
        );

    mux_inst_170: MUX2
        port map (
            O => mux_o_170,
            I0 => dpb_inst_12_douta(24),
            I1 => dpb_inst_13_douta(24),
            S0 => dff_q_2
        );

    mux_inst_171: MUX2
        port map (
            O => mux_o_171,
            I0 => dpb_inst_14_douta(24),
            I1 => dpb_inst_15_douta(24),
            S0 => dff_q_2
        );

    mux_inst_172: MUX2
        port map (
            O => mux_o_172,
            I0 => mux_o_168,
            I1 => mux_o_169,
            S0 => dff_q_1
        );

    mux_inst_173: MUX2
        port map (
            O => mux_o_173,
            I0 => mux_o_170,
            I1 => mux_o_171,
            S0 => dff_q_1
        );

    mux_inst_174: MUX2
        port map (
            O => douta(24),
            I0 => mux_o_172,
            I1 => mux_o_173,
            S0 => dff_q_0
        );

    mux_inst_175: MUX2
        port map (
            O => mux_o_175,
            I0 => dpb_inst_8_douta(25),
            I1 => dpb_inst_9_douta(25),
            S0 => dff_q_2
        );

    mux_inst_176: MUX2
        port map (
            O => mux_o_176,
            I0 => dpb_inst_10_douta(25),
            I1 => dpb_inst_11_douta(25),
            S0 => dff_q_2
        );

    mux_inst_177: MUX2
        port map (
            O => mux_o_177,
            I0 => dpb_inst_12_douta(25),
            I1 => dpb_inst_13_douta(25),
            S0 => dff_q_2
        );

    mux_inst_178: MUX2
        port map (
            O => mux_o_178,
            I0 => dpb_inst_14_douta(25),
            I1 => dpb_inst_15_douta(25),
            S0 => dff_q_2
        );

    mux_inst_179: MUX2
        port map (
            O => mux_o_179,
            I0 => mux_o_175,
            I1 => mux_o_176,
            S0 => dff_q_1
        );

    mux_inst_180: MUX2
        port map (
            O => mux_o_180,
            I0 => mux_o_177,
            I1 => mux_o_178,
            S0 => dff_q_1
        );

    mux_inst_181: MUX2
        port map (
            O => douta(25),
            I0 => mux_o_179,
            I1 => mux_o_180,
            S0 => dff_q_0
        );

    mux_inst_182: MUX2
        port map (
            O => mux_o_182,
            I0 => dpb_inst_8_douta(26),
            I1 => dpb_inst_9_douta(26),
            S0 => dff_q_2
        );

    mux_inst_183: MUX2
        port map (
            O => mux_o_183,
            I0 => dpb_inst_10_douta(26),
            I1 => dpb_inst_11_douta(26),
            S0 => dff_q_2
        );

    mux_inst_184: MUX2
        port map (
            O => mux_o_184,
            I0 => dpb_inst_12_douta(26),
            I1 => dpb_inst_13_douta(26),
            S0 => dff_q_2
        );

    mux_inst_185: MUX2
        port map (
            O => mux_o_185,
            I0 => dpb_inst_14_douta(26),
            I1 => dpb_inst_15_douta(26),
            S0 => dff_q_2
        );

    mux_inst_186: MUX2
        port map (
            O => mux_o_186,
            I0 => mux_o_182,
            I1 => mux_o_183,
            S0 => dff_q_1
        );

    mux_inst_187: MUX2
        port map (
            O => mux_o_187,
            I0 => mux_o_184,
            I1 => mux_o_185,
            S0 => dff_q_1
        );

    mux_inst_188: MUX2
        port map (
            O => douta(26),
            I0 => mux_o_186,
            I1 => mux_o_187,
            S0 => dff_q_0
        );

    mux_inst_189: MUX2
        port map (
            O => mux_o_189,
            I0 => dpb_inst_8_douta(27),
            I1 => dpb_inst_9_douta(27),
            S0 => dff_q_2
        );

    mux_inst_190: MUX2
        port map (
            O => mux_o_190,
            I0 => dpb_inst_10_douta(27),
            I1 => dpb_inst_11_douta(27),
            S0 => dff_q_2
        );

    mux_inst_191: MUX2
        port map (
            O => mux_o_191,
            I0 => dpb_inst_12_douta(27),
            I1 => dpb_inst_13_douta(27),
            S0 => dff_q_2
        );

    mux_inst_192: MUX2
        port map (
            O => mux_o_192,
            I0 => dpb_inst_14_douta(27),
            I1 => dpb_inst_15_douta(27),
            S0 => dff_q_2
        );

    mux_inst_193: MUX2
        port map (
            O => mux_o_193,
            I0 => mux_o_189,
            I1 => mux_o_190,
            S0 => dff_q_1
        );

    mux_inst_194: MUX2
        port map (
            O => mux_o_194,
            I0 => mux_o_191,
            I1 => mux_o_192,
            S0 => dff_q_1
        );

    mux_inst_195: MUX2
        port map (
            O => douta(27),
            I0 => mux_o_193,
            I1 => mux_o_194,
            S0 => dff_q_0
        );

    mux_inst_196: MUX2
        port map (
            O => mux_o_196,
            I0 => dpb_inst_8_douta(28),
            I1 => dpb_inst_9_douta(28),
            S0 => dff_q_2
        );

    mux_inst_197: MUX2
        port map (
            O => mux_o_197,
            I0 => dpb_inst_10_douta(28),
            I1 => dpb_inst_11_douta(28),
            S0 => dff_q_2
        );

    mux_inst_198: MUX2
        port map (
            O => mux_o_198,
            I0 => dpb_inst_12_douta(28),
            I1 => dpb_inst_13_douta(28),
            S0 => dff_q_2
        );

    mux_inst_199: MUX2
        port map (
            O => mux_o_199,
            I0 => dpb_inst_14_douta(28),
            I1 => dpb_inst_15_douta(28),
            S0 => dff_q_2
        );

    mux_inst_200: MUX2
        port map (
            O => mux_o_200,
            I0 => mux_o_196,
            I1 => mux_o_197,
            S0 => dff_q_1
        );

    mux_inst_201: MUX2
        port map (
            O => mux_o_201,
            I0 => mux_o_198,
            I1 => mux_o_199,
            S0 => dff_q_1
        );

    mux_inst_202: MUX2
        port map (
            O => douta(28),
            I0 => mux_o_200,
            I1 => mux_o_201,
            S0 => dff_q_0
        );

    mux_inst_203: MUX2
        port map (
            O => mux_o_203,
            I0 => dpb_inst_8_douta(29),
            I1 => dpb_inst_9_douta(29),
            S0 => dff_q_2
        );

    mux_inst_204: MUX2
        port map (
            O => mux_o_204,
            I0 => dpb_inst_10_douta(29),
            I1 => dpb_inst_11_douta(29),
            S0 => dff_q_2
        );

    mux_inst_205: MUX2
        port map (
            O => mux_o_205,
            I0 => dpb_inst_12_douta(29),
            I1 => dpb_inst_13_douta(29),
            S0 => dff_q_2
        );

    mux_inst_206: MUX2
        port map (
            O => mux_o_206,
            I0 => dpb_inst_14_douta(29),
            I1 => dpb_inst_15_douta(29),
            S0 => dff_q_2
        );

    mux_inst_207: MUX2
        port map (
            O => mux_o_207,
            I0 => mux_o_203,
            I1 => mux_o_204,
            S0 => dff_q_1
        );

    mux_inst_208: MUX2
        port map (
            O => mux_o_208,
            I0 => mux_o_205,
            I1 => mux_o_206,
            S0 => dff_q_1
        );

    mux_inst_209: MUX2
        port map (
            O => douta(29),
            I0 => mux_o_207,
            I1 => mux_o_208,
            S0 => dff_q_0
        );

    mux_inst_210: MUX2
        port map (
            O => mux_o_210,
            I0 => dpb_inst_8_douta(30),
            I1 => dpb_inst_9_douta(30),
            S0 => dff_q_2
        );

    mux_inst_211: MUX2
        port map (
            O => mux_o_211,
            I0 => dpb_inst_10_douta(30),
            I1 => dpb_inst_11_douta(30),
            S0 => dff_q_2
        );

    mux_inst_212: MUX2
        port map (
            O => mux_o_212,
            I0 => dpb_inst_12_douta(30),
            I1 => dpb_inst_13_douta(30),
            S0 => dff_q_2
        );

    mux_inst_213: MUX2
        port map (
            O => mux_o_213,
            I0 => dpb_inst_14_douta(30),
            I1 => dpb_inst_15_douta(30),
            S0 => dff_q_2
        );

    mux_inst_214: MUX2
        port map (
            O => mux_o_214,
            I0 => mux_o_210,
            I1 => mux_o_211,
            S0 => dff_q_1
        );

    mux_inst_215: MUX2
        port map (
            O => mux_o_215,
            I0 => mux_o_212,
            I1 => mux_o_213,
            S0 => dff_q_1
        );

    mux_inst_216: MUX2
        port map (
            O => douta(30),
            I0 => mux_o_214,
            I1 => mux_o_215,
            S0 => dff_q_0
        );

    mux_inst_217: MUX2
        port map (
            O => mux_o_217,
            I0 => dpb_inst_8_douta(31),
            I1 => dpb_inst_9_douta(31),
            S0 => dff_q_2
        );

    mux_inst_218: MUX2
        port map (
            O => mux_o_218,
            I0 => dpb_inst_10_douta(31),
            I1 => dpb_inst_11_douta(31),
            S0 => dff_q_2
        );

    mux_inst_219: MUX2
        port map (
            O => mux_o_219,
            I0 => dpb_inst_12_douta(31),
            I1 => dpb_inst_13_douta(31),
            S0 => dff_q_2
        );

    mux_inst_220: MUX2
        port map (
            O => mux_o_220,
            I0 => dpb_inst_14_douta(31),
            I1 => dpb_inst_15_douta(31),
            S0 => dff_q_2
        );

    mux_inst_221: MUX2
        port map (
            O => mux_o_221,
            I0 => mux_o_217,
            I1 => mux_o_218,
            S0 => dff_q_1
        );

    mux_inst_222: MUX2
        port map (
            O => mux_o_222,
            I0 => mux_o_219,
            I1 => mux_o_220,
            S0 => dff_q_1
        );

    mux_inst_223: MUX2
        port map (
            O => douta(31),
            I0 => mux_o_221,
            I1 => mux_o_222,
            S0 => dff_q_0
        );

    mux_inst_224: MUX2
        port map (
            O => mux_o_224,
            I0 => dpb_inst_0_doutb(0),
            I1 => dpb_inst_1_doutb(0),
            S0 => dff_q_5
        );

    mux_inst_225: MUX2
        port map (
            O => mux_o_225,
            I0 => dpb_inst_2_doutb(0),
            I1 => dpb_inst_3_doutb(0),
            S0 => dff_q_5
        );

    mux_inst_226: MUX2
        port map (
            O => mux_o_226,
            I0 => dpb_inst_4_doutb(0),
            I1 => dpb_inst_5_doutb(0),
            S0 => dff_q_5
        );

    mux_inst_227: MUX2
        port map (
            O => mux_o_227,
            I0 => dpb_inst_6_doutb(0),
            I1 => dpb_inst_7_doutb(0),
            S0 => dff_q_5
        );

    mux_inst_228: MUX2
        port map (
            O => mux_o_228,
            I0 => mux_o_224,
            I1 => mux_o_225,
            S0 => dff_q_4
        );

    mux_inst_229: MUX2
        port map (
            O => mux_o_229,
            I0 => mux_o_226,
            I1 => mux_o_227,
            S0 => dff_q_4
        );

    mux_inst_230: MUX2
        port map (
            O => doutb(0),
            I0 => mux_o_228,
            I1 => mux_o_229,
            S0 => dff_q_3
        );

    mux_inst_231: MUX2
        port map (
            O => mux_o_231,
            I0 => dpb_inst_0_doutb(1),
            I1 => dpb_inst_1_doutb(1),
            S0 => dff_q_5
        );

    mux_inst_232: MUX2
        port map (
            O => mux_o_232,
            I0 => dpb_inst_2_doutb(1),
            I1 => dpb_inst_3_doutb(1),
            S0 => dff_q_5
        );

    mux_inst_233: MUX2
        port map (
            O => mux_o_233,
            I0 => dpb_inst_4_doutb(1),
            I1 => dpb_inst_5_doutb(1),
            S0 => dff_q_5
        );

    mux_inst_234: MUX2
        port map (
            O => mux_o_234,
            I0 => dpb_inst_6_doutb(1),
            I1 => dpb_inst_7_doutb(1),
            S0 => dff_q_5
        );

    mux_inst_235: MUX2
        port map (
            O => mux_o_235,
            I0 => mux_o_231,
            I1 => mux_o_232,
            S0 => dff_q_4
        );

    mux_inst_236: MUX2
        port map (
            O => mux_o_236,
            I0 => mux_o_233,
            I1 => mux_o_234,
            S0 => dff_q_4
        );

    mux_inst_237: MUX2
        port map (
            O => doutb(1),
            I0 => mux_o_235,
            I1 => mux_o_236,
            S0 => dff_q_3
        );

    mux_inst_238: MUX2
        port map (
            O => mux_o_238,
            I0 => dpb_inst_0_doutb(2),
            I1 => dpb_inst_1_doutb(2),
            S0 => dff_q_5
        );

    mux_inst_239: MUX2
        port map (
            O => mux_o_239,
            I0 => dpb_inst_2_doutb(2),
            I1 => dpb_inst_3_doutb(2),
            S0 => dff_q_5
        );

    mux_inst_240: MUX2
        port map (
            O => mux_o_240,
            I0 => dpb_inst_4_doutb(2),
            I1 => dpb_inst_5_doutb(2),
            S0 => dff_q_5
        );

    mux_inst_241: MUX2
        port map (
            O => mux_o_241,
            I0 => dpb_inst_6_doutb(2),
            I1 => dpb_inst_7_doutb(2),
            S0 => dff_q_5
        );

    mux_inst_242: MUX2
        port map (
            O => mux_o_242,
            I0 => mux_o_238,
            I1 => mux_o_239,
            S0 => dff_q_4
        );

    mux_inst_243: MUX2
        port map (
            O => mux_o_243,
            I0 => mux_o_240,
            I1 => mux_o_241,
            S0 => dff_q_4
        );

    mux_inst_244: MUX2
        port map (
            O => doutb(2),
            I0 => mux_o_242,
            I1 => mux_o_243,
            S0 => dff_q_3
        );

    mux_inst_245: MUX2
        port map (
            O => mux_o_245,
            I0 => dpb_inst_0_doutb(3),
            I1 => dpb_inst_1_doutb(3),
            S0 => dff_q_5
        );

    mux_inst_246: MUX2
        port map (
            O => mux_o_246,
            I0 => dpb_inst_2_doutb(3),
            I1 => dpb_inst_3_doutb(3),
            S0 => dff_q_5
        );

    mux_inst_247: MUX2
        port map (
            O => mux_o_247,
            I0 => dpb_inst_4_doutb(3),
            I1 => dpb_inst_5_doutb(3),
            S0 => dff_q_5
        );

    mux_inst_248: MUX2
        port map (
            O => mux_o_248,
            I0 => dpb_inst_6_doutb(3),
            I1 => dpb_inst_7_doutb(3),
            S0 => dff_q_5
        );

    mux_inst_249: MUX2
        port map (
            O => mux_o_249,
            I0 => mux_o_245,
            I1 => mux_o_246,
            S0 => dff_q_4
        );

    mux_inst_250: MUX2
        port map (
            O => mux_o_250,
            I0 => mux_o_247,
            I1 => mux_o_248,
            S0 => dff_q_4
        );

    mux_inst_251: MUX2
        port map (
            O => doutb(3),
            I0 => mux_o_249,
            I1 => mux_o_250,
            S0 => dff_q_3
        );

    mux_inst_252: MUX2
        port map (
            O => mux_o_252,
            I0 => dpb_inst_0_doutb(4),
            I1 => dpb_inst_1_doutb(4),
            S0 => dff_q_5
        );

    mux_inst_253: MUX2
        port map (
            O => mux_o_253,
            I0 => dpb_inst_2_doutb(4),
            I1 => dpb_inst_3_doutb(4),
            S0 => dff_q_5
        );

    mux_inst_254: MUX2
        port map (
            O => mux_o_254,
            I0 => dpb_inst_4_doutb(4),
            I1 => dpb_inst_5_doutb(4),
            S0 => dff_q_5
        );

    mux_inst_255: MUX2
        port map (
            O => mux_o_255,
            I0 => dpb_inst_6_doutb(4),
            I1 => dpb_inst_7_doutb(4),
            S0 => dff_q_5
        );

    mux_inst_256: MUX2
        port map (
            O => mux_o_256,
            I0 => mux_o_252,
            I1 => mux_o_253,
            S0 => dff_q_4
        );

    mux_inst_257: MUX2
        port map (
            O => mux_o_257,
            I0 => mux_o_254,
            I1 => mux_o_255,
            S0 => dff_q_4
        );

    mux_inst_258: MUX2
        port map (
            O => doutb(4),
            I0 => mux_o_256,
            I1 => mux_o_257,
            S0 => dff_q_3
        );

    mux_inst_259: MUX2
        port map (
            O => mux_o_259,
            I0 => dpb_inst_0_doutb(5),
            I1 => dpb_inst_1_doutb(5),
            S0 => dff_q_5
        );

    mux_inst_260: MUX2
        port map (
            O => mux_o_260,
            I0 => dpb_inst_2_doutb(5),
            I1 => dpb_inst_3_doutb(5),
            S0 => dff_q_5
        );

    mux_inst_261: MUX2
        port map (
            O => mux_o_261,
            I0 => dpb_inst_4_doutb(5),
            I1 => dpb_inst_5_doutb(5),
            S0 => dff_q_5
        );

    mux_inst_262: MUX2
        port map (
            O => mux_o_262,
            I0 => dpb_inst_6_doutb(5),
            I1 => dpb_inst_7_doutb(5),
            S0 => dff_q_5
        );

    mux_inst_263: MUX2
        port map (
            O => mux_o_263,
            I0 => mux_o_259,
            I1 => mux_o_260,
            S0 => dff_q_4
        );

    mux_inst_264: MUX2
        port map (
            O => mux_o_264,
            I0 => mux_o_261,
            I1 => mux_o_262,
            S0 => dff_q_4
        );

    mux_inst_265: MUX2
        port map (
            O => doutb(5),
            I0 => mux_o_263,
            I1 => mux_o_264,
            S0 => dff_q_3
        );

    mux_inst_266: MUX2
        port map (
            O => mux_o_266,
            I0 => dpb_inst_0_doutb(6),
            I1 => dpb_inst_1_doutb(6),
            S0 => dff_q_5
        );

    mux_inst_267: MUX2
        port map (
            O => mux_o_267,
            I0 => dpb_inst_2_doutb(6),
            I1 => dpb_inst_3_doutb(6),
            S0 => dff_q_5
        );

    mux_inst_268: MUX2
        port map (
            O => mux_o_268,
            I0 => dpb_inst_4_doutb(6),
            I1 => dpb_inst_5_doutb(6),
            S0 => dff_q_5
        );

    mux_inst_269: MUX2
        port map (
            O => mux_o_269,
            I0 => dpb_inst_6_doutb(6),
            I1 => dpb_inst_7_doutb(6),
            S0 => dff_q_5
        );

    mux_inst_270: MUX2
        port map (
            O => mux_o_270,
            I0 => mux_o_266,
            I1 => mux_o_267,
            S0 => dff_q_4
        );

    mux_inst_271: MUX2
        port map (
            O => mux_o_271,
            I0 => mux_o_268,
            I1 => mux_o_269,
            S0 => dff_q_4
        );

    mux_inst_272: MUX2
        port map (
            O => doutb(6),
            I0 => mux_o_270,
            I1 => mux_o_271,
            S0 => dff_q_3
        );

    mux_inst_273: MUX2
        port map (
            O => mux_o_273,
            I0 => dpb_inst_0_doutb(7),
            I1 => dpb_inst_1_doutb(7),
            S0 => dff_q_5
        );

    mux_inst_274: MUX2
        port map (
            O => mux_o_274,
            I0 => dpb_inst_2_doutb(7),
            I1 => dpb_inst_3_doutb(7),
            S0 => dff_q_5
        );

    mux_inst_275: MUX2
        port map (
            O => mux_o_275,
            I0 => dpb_inst_4_doutb(7),
            I1 => dpb_inst_5_doutb(7),
            S0 => dff_q_5
        );

    mux_inst_276: MUX2
        port map (
            O => mux_o_276,
            I0 => dpb_inst_6_doutb(7),
            I1 => dpb_inst_7_doutb(7),
            S0 => dff_q_5
        );

    mux_inst_277: MUX2
        port map (
            O => mux_o_277,
            I0 => mux_o_273,
            I1 => mux_o_274,
            S0 => dff_q_4
        );

    mux_inst_278: MUX2
        port map (
            O => mux_o_278,
            I0 => mux_o_275,
            I1 => mux_o_276,
            S0 => dff_q_4
        );

    mux_inst_279: MUX2
        port map (
            O => doutb(7),
            I0 => mux_o_277,
            I1 => mux_o_278,
            S0 => dff_q_3
        );

    mux_inst_280: MUX2
        port map (
            O => mux_o_280,
            I0 => dpb_inst_0_doutb(8),
            I1 => dpb_inst_1_doutb(8),
            S0 => dff_q_5
        );

    mux_inst_281: MUX2
        port map (
            O => mux_o_281,
            I0 => dpb_inst_2_doutb(8),
            I1 => dpb_inst_3_doutb(8),
            S0 => dff_q_5
        );

    mux_inst_282: MUX2
        port map (
            O => mux_o_282,
            I0 => dpb_inst_4_doutb(8),
            I1 => dpb_inst_5_doutb(8),
            S0 => dff_q_5
        );

    mux_inst_283: MUX2
        port map (
            O => mux_o_283,
            I0 => dpb_inst_6_doutb(8),
            I1 => dpb_inst_7_doutb(8),
            S0 => dff_q_5
        );

    mux_inst_284: MUX2
        port map (
            O => mux_o_284,
            I0 => mux_o_280,
            I1 => mux_o_281,
            S0 => dff_q_4
        );

    mux_inst_285: MUX2
        port map (
            O => mux_o_285,
            I0 => mux_o_282,
            I1 => mux_o_283,
            S0 => dff_q_4
        );

    mux_inst_286: MUX2
        port map (
            O => doutb(8),
            I0 => mux_o_284,
            I1 => mux_o_285,
            S0 => dff_q_3
        );

    mux_inst_287: MUX2
        port map (
            O => mux_o_287,
            I0 => dpb_inst_0_doutb(9),
            I1 => dpb_inst_1_doutb(9),
            S0 => dff_q_5
        );

    mux_inst_288: MUX2
        port map (
            O => mux_o_288,
            I0 => dpb_inst_2_doutb(9),
            I1 => dpb_inst_3_doutb(9),
            S0 => dff_q_5
        );

    mux_inst_289: MUX2
        port map (
            O => mux_o_289,
            I0 => dpb_inst_4_doutb(9),
            I1 => dpb_inst_5_doutb(9),
            S0 => dff_q_5
        );

    mux_inst_290: MUX2
        port map (
            O => mux_o_290,
            I0 => dpb_inst_6_doutb(9),
            I1 => dpb_inst_7_doutb(9),
            S0 => dff_q_5
        );

    mux_inst_291: MUX2
        port map (
            O => mux_o_291,
            I0 => mux_o_287,
            I1 => mux_o_288,
            S0 => dff_q_4
        );

    mux_inst_292: MUX2
        port map (
            O => mux_o_292,
            I0 => mux_o_289,
            I1 => mux_o_290,
            S0 => dff_q_4
        );

    mux_inst_293: MUX2
        port map (
            O => doutb(9),
            I0 => mux_o_291,
            I1 => mux_o_292,
            S0 => dff_q_3
        );

    mux_inst_294: MUX2
        port map (
            O => mux_o_294,
            I0 => dpb_inst_0_doutb(10),
            I1 => dpb_inst_1_doutb(10),
            S0 => dff_q_5
        );

    mux_inst_295: MUX2
        port map (
            O => mux_o_295,
            I0 => dpb_inst_2_doutb(10),
            I1 => dpb_inst_3_doutb(10),
            S0 => dff_q_5
        );

    mux_inst_296: MUX2
        port map (
            O => mux_o_296,
            I0 => dpb_inst_4_doutb(10),
            I1 => dpb_inst_5_doutb(10),
            S0 => dff_q_5
        );

    mux_inst_297: MUX2
        port map (
            O => mux_o_297,
            I0 => dpb_inst_6_doutb(10),
            I1 => dpb_inst_7_doutb(10),
            S0 => dff_q_5
        );

    mux_inst_298: MUX2
        port map (
            O => mux_o_298,
            I0 => mux_o_294,
            I1 => mux_o_295,
            S0 => dff_q_4
        );

    mux_inst_299: MUX2
        port map (
            O => mux_o_299,
            I0 => mux_o_296,
            I1 => mux_o_297,
            S0 => dff_q_4
        );

    mux_inst_300: MUX2
        port map (
            O => doutb(10),
            I0 => mux_o_298,
            I1 => mux_o_299,
            S0 => dff_q_3
        );

    mux_inst_301: MUX2
        port map (
            O => mux_o_301,
            I0 => dpb_inst_0_doutb(11),
            I1 => dpb_inst_1_doutb(11),
            S0 => dff_q_5
        );

    mux_inst_302: MUX2
        port map (
            O => mux_o_302,
            I0 => dpb_inst_2_doutb(11),
            I1 => dpb_inst_3_doutb(11),
            S0 => dff_q_5
        );

    mux_inst_303: MUX2
        port map (
            O => mux_o_303,
            I0 => dpb_inst_4_doutb(11),
            I1 => dpb_inst_5_doutb(11),
            S0 => dff_q_5
        );

    mux_inst_304: MUX2
        port map (
            O => mux_o_304,
            I0 => dpb_inst_6_doutb(11),
            I1 => dpb_inst_7_doutb(11),
            S0 => dff_q_5
        );

    mux_inst_305: MUX2
        port map (
            O => mux_o_305,
            I0 => mux_o_301,
            I1 => mux_o_302,
            S0 => dff_q_4
        );

    mux_inst_306: MUX2
        port map (
            O => mux_o_306,
            I0 => mux_o_303,
            I1 => mux_o_304,
            S0 => dff_q_4
        );

    mux_inst_307: MUX2
        port map (
            O => doutb(11),
            I0 => mux_o_305,
            I1 => mux_o_306,
            S0 => dff_q_3
        );

    mux_inst_308: MUX2
        port map (
            O => mux_o_308,
            I0 => dpb_inst_0_doutb(12),
            I1 => dpb_inst_1_doutb(12),
            S0 => dff_q_5
        );

    mux_inst_309: MUX2
        port map (
            O => mux_o_309,
            I0 => dpb_inst_2_doutb(12),
            I1 => dpb_inst_3_doutb(12),
            S0 => dff_q_5
        );

    mux_inst_310: MUX2
        port map (
            O => mux_o_310,
            I0 => dpb_inst_4_doutb(12),
            I1 => dpb_inst_5_doutb(12),
            S0 => dff_q_5
        );

    mux_inst_311: MUX2
        port map (
            O => mux_o_311,
            I0 => dpb_inst_6_doutb(12),
            I1 => dpb_inst_7_doutb(12),
            S0 => dff_q_5
        );

    mux_inst_312: MUX2
        port map (
            O => mux_o_312,
            I0 => mux_o_308,
            I1 => mux_o_309,
            S0 => dff_q_4
        );

    mux_inst_313: MUX2
        port map (
            O => mux_o_313,
            I0 => mux_o_310,
            I1 => mux_o_311,
            S0 => dff_q_4
        );

    mux_inst_314: MUX2
        port map (
            O => doutb(12),
            I0 => mux_o_312,
            I1 => mux_o_313,
            S0 => dff_q_3
        );

    mux_inst_315: MUX2
        port map (
            O => mux_o_315,
            I0 => dpb_inst_0_doutb(13),
            I1 => dpb_inst_1_doutb(13),
            S0 => dff_q_5
        );

    mux_inst_316: MUX2
        port map (
            O => mux_o_316,
            I0 => dpb_inst_2_doutb(13),
            I1 => dpb_inst_3_doutb(13),
            S0 => dff_q_5
        );

    mux_inst_317: MUX2
        port map (
            O => mux_o_317,
            I0 => dpb_inst_4_doutb(13),
            I1 => dpb_inst_5_doutb(13),
            S0 => dff_q_5
        );

    mux_inst_318: MUX2
        port map (
            O => mux_o_318,
            I0 => dpb_inst_6_doutb(13),
            I1 => dpb_inst_7_doutb(13),
            S0 => dff_q_5
        );

    mux_inst_319: MUX2
        port map (
            O => mux_o_319,
            I0 => mux_o_315,
            I1 => mux_o_316,
            S0 => dff_q_4
        );

    mux_inst_320: MUX2
        port map (
            O => mux_o_320,
            I0 => mux_o_317,
            I1 => mux_o_318,
            S0 => dff_q_4
        );

    mux_inst_321: MUX2
        port map (
            O => doutb(13),
            I0 => mux_o_319,
            I1 => mux_o_320,
            S0 => dff_q_3
        );

    mux_inst_322: MUX2
        port map (
            O => mux_o_322,
            I0 => dpb_inst_0_doutb(14),
            I1 => dpb_inst_1_doutb(14),
            S0 => dff_q_5
        );

    mux_inst_323: MUX2
        port map (
            O => mux_o_323,
            I0 => dpb_inst_2_doutb(14),
            I1 => dpb_inst_3_doutb(14),
            S0 => dff_q_5
        );

    mux_inst_324: MUX2
        port map (
            O => mux_o_324,
            I0 => dpb_inst_4_doutb(14),
            I1 => dpb_inst_5_doutb(14),
            S0 => dff_q_5
        );

    mux_inst_325: MUX2
        port map (
            O => mux_o_325,
            I0 => dpb_inst_6_doutb(14),
            I1 => dpb_inst_7_doutb(14),
            S0 => dff_q_5
        );

    mux_inst_326: MUX2
        port map (
            O => mux_o_326,
            I0 => mux_o_322,
            I1 => mux_o_323,
            S0 => dff_q_4
        );

    mux_inst_327: MUX2
        port map (
            O => mux_o_327,
            I0 => mux_o_324,
            I1 => mux_o_325,
            S0 => dff_q_4
        );

    mux_inst_328: MUX2
        port map (
            O => doutb(14),
            I0 => mux_o_326,
            I1 => mux_o_327,
            S0 => dff_q_3
        );

    mux_inst_329: MUX2
        port map (
            O => mux_o_329,
            I0 => dpb_inst_0_doutb(15),
            I1 => dpb_inst_1_doutb(15),
            S0 => dff_q_5
        );

    mux_inst_330: MUX2
        port map (
            O => mux_o_330,
            I0 => dpb_inst_2_doutb(15),
            I1 => dpb_inst_3_doutb(15),
            S0 => dff_q_5
        );

    mux_inst_331: MUX2
        port map (
            O => mux_o_331,
            I0 => dpb_inst_4_doutb(15),
            I1 => dpb_inst_5_doutb(15),
            S0 => dff_q_5
        );

    mux_inst_332: MUX2
        port map (
            O => mux_o_332,
            I0 => dpb_inst_6_doutb(15),
            I1 => dpb_inst_7_doutb(15),
            S0 => dff_q_5
        );

    mux_inst_333: MUX2
        port map (
            O => mux_o_333,
            I0 => mux_o_329,
            I1 => mux_o_330,
            S0 => dff_q_4
        );

    mux_inst_334: MUX2
        port map (
            O => mux_o_334,
            I0 => mux_o_331,
            I1 => mux_o_332,
            S0 => dff_q_4
        );

    mux_inst_335: MUX2
        port map (
            O => doutb(15),
            I0 => mux_o_333,
            I1 => mux_o_334,
            S0 => dff_q_3
        );

    mux_inst_336: MUX2
        port map (
            O => mux_o_336,
            I0 => dpb_inst_8_doutb(16),
            I1 => dpb_inst_9_doutb(16),
            S0 => dff_q_5
        );

    mux_inst_337: MUX2
        port map (
            O => mux_o_337,
            I0 => dpb_inst_10_doutb(16),
            I1 => dpb_inst_11_doutb(16),
            S0 => dff_q_5
        );

    mux_inst_338: MUX2
        port map (
            O => mux_o_338,
            I0 => dpb_inst_12_doutb(16),
            I1 => dpb_inst_13_doutb(16),
            S0 => dff_q_5
        );

    mux_inst_339: MUX2
        port map (
            O => mux_o_339,
            I0 => dpb_inst_14_doutb(16),
            I1 => dpb_inst_15_doutb(16),
            S0 => dff_q_5
        );

    mux_inst_340: MUX2
        port map (
            O => mux_o_340,
            I0 => mux_o_336,
            I1 => mux_o_337,
            S0 => dff_q_4
        );

    mux_inst_341: MUX2
        port map (
            O => mux_o_341,
            I0 => mux_o_338,
            I1 => mux_o_339,
            S0 => dff_q_4
        );

    mux_inst_342: MUX2
        port map (
            O => doutb(16),
            I0 => mux_o_340,
            I1 => mux_o_341,
            S0 => dff_q_3
        );

    mux_inst_343: MUX2
        port map (
            O => mux_o_343,
            I0 => dpb_inst_8_doutb(17),
            I1 => dpb_inst_9_doutb(17),
            S0 => dff_q_5
        );

    mux_inst_344: MUX2
        port map (
            O => mux_o_344,
            I0 => dpb_inst_10_doutb(17),
            I1 => dpb_inst_11_doutb(17),
            S0 => dff_q_5
        );

    mux_inst_345: MUX2
        port map (
            O => mux_o_345,
            I0 => dpb_inst_12_doutb(17),
            I1 => dpb_inst_13_doutb(17),
            S0 => dff_q_5
        );

    mux_inst_346: MUX2
        port map (
            O => mux_o_346,
            I0 => dpb_inst_14_doutb(17),
            I1 => dpb_inst_15_doutb(17),
            S0 => dff_q_5
        );

    mux_inst_347: MUX2
        port map (
            O => mux_o_347,
            I0 => mux_o_343,
            I1 => mux_o_344,
            S0 => dff_q_4
        );

    mux_inst_348: MUX2
        port map (
            O => mux_o_348,
            I0 => mux_o_345,
            I1 => mux_o_346,
            S0 => dff_q_4
        );

    mux_inst_349: MUX2
        port map (
            O => doutb(17),
            I0 => mux_o_347,
            I1 => mux_o_348,
            S0 => dff_q_3
        );

    mux_inst_350: MUX2
        port map (
            O => mux_o_350,
            I0 => dpb_inst_8_doutb(18),
            I1 => dpb_inst_9_doutb(18),
            S0 => dff_q_5
        );

    mux_inst_351: MUX2
        port map (
            O => mux_o_351,
            I0 => dpb_inst_10_doutb(18),
            I1 => dpb_inst_11_doutb(18),
            S0 => dff_q_5
        );

    mux_inst_352: MUX2
        port map (
            O => mux_o_352,
            I0 => dpb_inst_12_doutb(18),
            I1 => dpb_inst_13_doutb(18),
            S0 => dff_q_5
        );

    mux_inst_353: MUX2
        port map (
            O => mux_o_353,
            I0 => dpb_inst_14_doutb(18),
            I1 => dpb_inst_15_doutb(18),
            S0 => dff_q_5
        );

    mux_inst_354: MUX2
        port map (
            O => mux_o_354,
            I0 => mux_o_350,
            I1 => mux_o_351,
            S0 => dff_q_4
        );

    mux_inst_355: MUX2
        port map (
            O => mux_o_355,
            I0 => mux_o_352,
            I1 => mux_o_353,
            S0 => dff_q_4
        );

    mux_inst_356: MUX2
        port map (
            O => doutb(18),
            I0 => mux_o_354,
            I1 => mux_o_355,
            S0 => dff_q_3
        );

    mux_inst_357: MUX2
        port map (
            O => mux_o_357,
            I0 => dpb_inst_8_doutb(19),
            I1 => dpb_inst_9_doutb(19),
            S0 => dff_q_5
        );

    mux_inst_358: MUX2
        port map (
            O => mux_o_358,
            I0 => dpb_inst_10_doutb(19),
            I1 => dpb_inst_11_doutb(19),
            S0 => dff_q_5
        );

    mux_inst_359: MUX2
        port map (
            O => mux_o_359,
            I0 => dpb_inst_12_doutb(19),
            I1 => dpb_inst_13_doutb(19),
            S0 => dff_q_5
        );

    mux_inst_360: MUX2
        port map (
            O => mux_o_360,
            I0 => dpb_inst_14_doutb(19),
            I1 => dpb_inst_15_doutb(19),
            S0 => dff_q_5
        );

    mux_inst_361: MUX2
        port map (
            O => mux_o_361,
            I0 => mux_o_357,
            I1 => mux_o_358,
            S0 => dff_q_4
        );

    mux_inst_362: MUX2
        port map (
            O => mux_o_362,
            I0 => mux_o_359,
            I1 => mux_o_360,
            S0 => dff_q_4
        );

    mux_inst_363: MUX2
        port map (
            O => doutb(19),
            I0 => mux_o_361,
            I1 => mux_o_362,
            S0 => dff_q_3
        );

    mux_inst_364: MUX2
        port map (
            O => mux_o_364,
            I0 => dpb_inst_8_doutb(20),
            I1 => dpb_inst_9_doutb(20),
            S0 => dff_q_5
        );

    mux_inst_365: MUX2
        port map (
            O => mux_o_365,
            I0 => dpb_inst_10_doutb(20),
            I1 => dpb_inst_11_doutb(20),
            S0 => dff_q_5
        );

    mux_inst_366: MUX2
        port map (
            O => mux_o_366,
            I0 => dpb_inst_12_doutb(20),
            I1 => dpb_inst_13_doutb(20),
            S0 => dff_q_5
        );

    mux_inst_367: MUX2
        port map (
            O => mux_o_367,
            I0 => dpb_inst_14_doutb(20),
            I1 => dpb_inst_15_doutb(20),
            S0 => dff_q_5
        );

    mux_inst_368: MUX2
        port map (
            O => mux_o_368,
            I0 => mux_o_364,
            I1 => mux_o_365,
            S0 => dff_q_4
        );

    mux_inst_369: MUX2
        port map (
            O => mux_o_369,
            I0 => mux_o_366,
            I1 => mux_o_367,
            S0 => dff_q_4
        );

    mux_inst_370: MUX2
        port map (
            O => doutb(20),
            I0 => mux_o_368,
            I1 => mux_o_369,
            S0 => dff_q_3
        );

    mux_inst_371: MUX2
        port map (
            O => mux_o_371,
            I0 => dpb_inst_8_doutb(21),
            I1 => dpb_inst_9_doutb(21),
            S0 => dff_q_5
        );

    mux_inst_372: MUX2
        port map (
            O => mux_o_372,
            I0 => dpb_inst_10_doutb(21),
            I1 => dpb_inst_11_doutb(21),
            S0 => dff_q_5
        );

    mux_inst_373: MUX2
        port map (
            O => mux_o_373,
            I0 => dpb_inst_12_doutb(21),
            I1 => dpb_inst_13_doutb(21),
            S0 => dff_q_5
        );

    mux_inst_374: MUX2
        port map (
            O => mux_o_374,
            I0 => dpb_inst_14_doutb(21),
            I1 => dpb_inst_15_doutb(21),
            S0 => dff_q_5
        );

    mux_inst_375: MUX2
        port map (
            O => mux_o_375,
            I0 => mux_o_371,
            I1 => mux_o_372,
            S0 => dff_q_4
        );

    mux_inst_376: MUX2
        port map (
            O => mux_o_376,
            I0 => mux_o_373,
            I1 => mux_o_374,
            S0 => dff_q_4
        );

    mux_inst_377: MUX2
        port map (
            O => doutb(21),
            I0 => mux_o_375,
            I1 => mux_o_376,
            S0 => dff_q_3
        );

    mux_inst_378: MUX2
        port map (
            O => mux_o_378,
            I0 => dpb_inst_8_doutb(22),
            I1 => dpb_inst_9_doutb(22),
            S0 => dff_q_5
        );

    mux_inst_379: MUX2
        port map (
            O => mux_o_379,
            I0 => dpb_inst_10_doutb(22),
            I1 => dpb_inst_11_doutb(22),
            S0 => dff_q_5
        );

    mux_inst_380: MUX2
        port map (
            O => mux_o_380,
            I0 => dpb_inst_12_doutb(22),
            I1 => dpb_inst_13_doutb(22),
            S0 => dff_q_5
        );

    mux_inst_381: MUX2
        port map (
            O => mux_o_381,
            I0 => dpb_inst_14_doutb(22),
            I1 => dpb_inst_15_doutb(22),
            S0 => dff_q_5
        );

    mux_inst_382: MUX2
        port map (
            O => mux_o_382,
            I0 => mux_o_378,
            I1 => mux_o_379,
            S0 => dff_q_4
        );

    mux_inst_383: MUX2
        port map (
            O => mux_o_383,
            I0 => mux_o_380,
            I1 => mux_o_381,
            S0 => dff_q_4
        );

    mux_inst_384: MUX2
        port map (
            O => doutb(22),
            I0 => mux_o_382,
            I1 => mux_o_383,
            S0 => dff_q_3
        );

    mux_inst_385: MUX2
        port map (
            O => mux_o_385,
            I0 => dpb_inst_8_doutb(23),
            I1 => dpb_inst_9_doutb(23),
            S0 => dff_q_5
        );

    mux_inst_386: MUX2
        port map (
            O => mux_o_386,
            I0 => dpb_inst_10_doutb(23),
            I1 => dpb_inst_11_doutb(23),
            S0 => dff_q_5
        );

    mux_inst_387: MUX2
        port map (
            O => mux_o_387,
            I0 => dpb_inst_12_doutb(23),
            I1 => dpb_inst_13_doutb(23),
            S0 => dff_q_5
        );

    mux_inst_388: MUX2
        port map (
            O => mux_o_388,
            I0 => dpb_inst_14_doutb(23),
            I1 => dpb_inst_15_doutb(23),
            S0 => dff_q_5
        );

    mux_inst_389: MUX2
        port map (
            O => mux_o_389,
            I0 => mux_o_385,
            I1 => mux_o_386,
            S0 => dff_q_4
        );

    mux_inst_390: MUX2
        port map (
            O => mux_o_390,
            I0 => mux_o_387,
            I1 => mux_o_388,
            S0 => dff_q_4
        );

    mux_inst_391: MUX2
        port map (
            O => doutb(23),
            I0 => mux_o_389,
            I1 => mux_o_390,
            S0 => dff_q_3
        );

    mux_inst_392: MUX2
        port map (
            O => mux_o_392,
            I0 => dpb_inst_8_doutb(24),
            I1 => dpb_inst_9_doutb(24),
            S0 => dff_q_5
        );

    mux_inst_393: MUX2
        port map (
            O => mux_o_393,
            I0 => dpb_inst_10_doutb(24),
            I1 => dpb_inst_11_doutb(24),
            S0 => dff_q_5
        );

    mux_inst_394: MUX2
        port map (
            O => mux_o_394,
            I0 => dpb_inst_12_doutb(24),
            I1 => dpb_inst_13_doutb(24),
            S0 => dff_q_5
        );

    mux_inst_395: MUX2
        port map (
            O => mux_o_395,
            I0 => dpb_inst_14_doutb(24),
            I1 => dpb_inst_15_doutb(24),
            S0 => dff_q_5
        );

    mux_inst_396: MUX2
        port map (
            O => mux_o_396,
            I0 => mux_o_392,
            I1 => mux_o_393,
            S0 => dff_q_4
        );

    mux_inst_397: MUX2
        port map (
            O => mux_o_397,
            I0 => mux_o_394,
            I1 => mux_o_395,
            S0 => dff_q_4
        );

    mux_inst_398: MUX2
        port map (
            O => doutb(24),
            I0 => mux_o_396,
            I1 => mux_o_397,
            S0 => dff_q_3
        );

    mux_inst_399: MUX2
        port map (
            O => mux_o_399,
            I0 => dpb_inst_8_doutb(25),
            I1 => dpb_inst_9_doutb(25),
            S0 => dff_q_5
        );

    mux_inst_400: MUX2
        port map (
            O => mux_o_400,
            I0 => dpb_inst_10_doutb(25),
            I1 => dpb_inst_11_doutb(25),
            S0 => dff_q_5
        );

    mux_inst_401: MUX2
        port map (
            O => mux_o_401,
            I0 => dpb_inst_12_doutb(25),
            I1 => dpb_inst_13_doutb(25),
            S0 => dff_q_5
        );

    mux_inst_402: MUX2
        port map (
            O => mux_o_402,
            I0 => dpb_inst_14_doutb(25),
            I1 => dpb_inst_15_doutb(25),
            S0 => dff_q_5
        );

    mux_inst_403: MUX2
        port map (
            O => mux_o_403,
            I0 => mux_o_399,
            I1 => mux_o_400,
            S0 => dff_q_4
        );

    mux_inst_404: MUX2
        port map (
            O => mux_o_404,
            I0 => mux_o_401,
            I1 => mux_o_402,
            S0 => dff_q_4
        );

    mux_inst_405: MUX2
        port map (
            O => doutb(25),
            I0 => mux_o_403,
            I1 => mux_o_404,
            S0 => dff_q_3
        );

    mux_inst_406: MUX2
        port map (
            O => mux_o_406,
            I0 => dpb_inst_8_doutb(26),
            I1 => dpb_inst_9_doutb(26),
            S0 => dff_q_5
        );

    mux_inst_407: MUX2
        port map (
            O => mux_o_407,
            I0 => dpb_inst_10_doutb(26),
            I1 => dpb_inst_11_doutb(26),
            S0 => dff_q_5
        );

    mux_inst_408: MUX2
        port map (
            O => mux_o_408,
            I0 => dpb_inst_12_doutb(26),
            I1 => dpb_inst_13_doutb(26),
            S0 => dff_q_5
        );

    mux_inst_409: MUX2
        port map (
            O => mux_o_409,
            I0 => dpb_inst_14_doutb(26),
            I1 => dpb_inst_15_doutb(26),
            S0 => dff_q_5
        );

    mux_inst_410: MUX2
        port map (
            O => mux_o_410,
            I0 => mux_o_406,
            I1 => mux_o_407,
            S0 => dff_q_4
        );

    mux_inst_411: MUX2
        port map (
            O => mux_o_411,
            I0 => mux_o_408,
            I1 => mux_o_409,
            S0 => dff_q_4
        );

    mux_inst_412: MUX2
        port map (
            O => doutb(26),
            I0 => mux_o_410,
            I1 => mux_o_411,
            S0 => dff_q_3
        );

    mux_inst_413: MUX2
        port map (
            O => mux_o_413,
            I0 => dpb_inst_8_doutb(27),
            I1 => dpb_inst_9_doutb(27),
            S0 => dff_q_5
        );

    mux_inst_414: MUX2
        port map (
            O => mux_o_414,
            I0 => dpb_inst_10_doutb(27),
            I1 => dpb_inst_11_doutb(27),
            S0 => dff_q_5
        );

    mux_inst_415: MUX2
        port map (
            O => mux_o_415,
            I0 => dpb_inst_12_doutb(27),
            I1 => dpb_inst_13_doutb(27),
            S0 => dff_q_5
        );

    mux_inst_416: MUX2
        port map (
            O => mux_o_416,
            I0 => dpb_inst_14_doutb(27),
            I1 => dpb_inst_15_doutb(27),
            S0 => dff_q_5
        );

    mux_inst_417: MUX2
        port map (
            O => mux_o_417,
            I0 => mux_o_413,
            I1 => mux_o_414,
            S0 => dff_q_4
        );

    mux_inst_418: MUX2
        port map (
            O => mux_o_418,
            I0 => mux_o_415,
            I1 => mux_o_416,
            S0 => dff_q_4
        );

    mux_inst_419: MUX2
        port map (
            O => doutb(27),
            I0 => mux_o_417,
            I1 => mux_o_418,
            S0 => dff_q_3
        );

    mux_inst_420: MUX2
        port map (
            O => mux_o_420,
            I0 => dpb_inst_8_doutb(28),
            I1 => dpb_inst_9_doutb(28),
            S0 => dff_q_5
        );

    mux_inst_421: MUX2
        port map (
            O => mux_o_421,
            I0 => dpb_inst_10_doutb(28),
            I1 => dpb_inst_11_doutb(28),
            S0 => dff_q_5
        );

    mux_inst_422: MUX2
        port map (
            O => mux_o_422,
            I0 => dpb_inst_12_doutb(28),
            I1 => dpb_inst_13_doutb(28),
            S0 => dff_q_5
        );

    mux_inst_423: MUX2
        port map (
            O => mux_o_423,
            I0 => dpb_inst_14_doutb(28),
            I1 => dpb_inst_15_doutb(28),
            S0 => dff_q_5
        );

    mux_inst_424: MUX2
        port map (
            O => mux_o_424,
            I0 => mux_o_420,
            I1 => mux_o_421,
            S0 => dff_q_4
        );

    mux_inst_425: MUX2
        port map (
            O => mux_o_425,
            I0 => mux_o_422,
            I1 => mux_o_423,
            S0 => dff_q_4
        );

    mux_inst_426: MUX2
        port map (
            O => doutb(28),
            I0 => mux_o_424,
            I1 => mux_o_425,
            S0 => dff_q_3
        );

    mux_inst_427: MUX2
        port map (
            O => mux_o_427,
            I0 => dpb_inst_8_doutb(29),
            I1 => dpb_inst_9_doutb(29),
            S0 => dff_q_5
        );

    mux_inst_428: MUX2
        port map (
            O => mux_o_428,
            I0 => dpb_inst_10_doutb(29),
            I1 => dpb_inst_11_doutb(29),
            S0 => dff_q_5
        );

    mux_inst_429: MUX2
        port map (
            O => mux_o_429,
            I0 => dpb_inst_12_doutb(29),
            I1 => dpb_inst_13_doutb(29),
            S0 => dff_q_5
        );

    mux_inst_430: MUX2
        port map (
            O => mux_o_430,
            I0 => dpb_inst_14_doutb(29),
            I1 => dpb_inst_15_doutb(29),
            S0 => dff_q_5
        );

    mux_inst_431: MUX2
        port map (
            O => mux_o_431,
            I0 => mux_o_427,
            I1 => mux_o_428,
            S0 => dff_q_4
        );

    mux_inst_432: MUX2
        port map (
            O => mux_o_432,
            I0 => mux_o_429,
            I1 => mux_o_430,
            S0 => dff_q_4
        );

    mux_inst_433: MUX2
        port map (
            O => doutb(29),
            I0 => mux_o_431,
            I1 => mux_o_432,
            S0 => dff_q_3
        );

    mux_inst_434: MUX2
        port map (
            O => mux_o_434,
            I0 => dpb_inst_8_doutb(30),
            I1 => dpb_inst_9_doutb(30),
            S0 => dff_q_5
        );

    mux_inst_435: MUX2
        port map (
            O => mux_o_435,
            I0 => dpb_inst_10_doutb(30),
            I1 => dpb_inst_11_doutb(30),
            S0 => dff_q_5
        );

    mux_inst_436: MUX2
        port map (
            O => mux_o_436,
            I0 => dpb_inst_12_doutb(30),
            I1 => dpb_inst_13_doutb(30),
            S0 => dff_q_5
        );

    mux_inst_437: MUX2
        port map (
            O => mux_o_437,
            I0 => dpb_inst_14_doutb(30),
            I1 => dpb_inst_15_doutb(30),
            S0 => dff_q_5
        );

    mux_inst_438: MUX2
        port map (
            O => mux_o_438,
            I0 => mux_o_434,
            I1 => mux_o_435,
            S0 => dff_q_4
        );

    mux_inst_439: MUX2
        port map (
            O => mux_o_439,
            I0 => mux_o_436,
            I1 => mux_o_437,
            S0 => dff_q_4
        );

    mux_inst_440: MUX2
        port map (
            O => doutb(30),
            I0 => mux_o_438,
            I1 => mux_o_439,
            S0 => dff_q_3
        );

    mux_inst_441: MUX2
        port map (
            O => mux_o_441,
            I0 => dpb_inst_8_doutb(31),
            I1 => dpb_inst_9_doutb(31),
            S0 => dff_q_5
        );

    mux_inst_442: MUX2
        port map (
            O => mux_o_442,
            I0 => dpb_inst_10_doutb(31),
            I1 => dpb_inst_11_doutb(31),
            S0 => dff_q_5
        );

    mux_inst_443: MUX2
        port map (
            O => mux_o_443,
            I0 => dpb_inst_12_doutb(31),
            I1 => dpb_inst_13_doutb(31),
            S0 => dff_q_5
        );

    mux_inst_444: MUX2
        port map (
            O => mux_o_444,
            I0 => dpb_inst_14_doutb(31),
            I1 => dpb_inst_15_doutb(31),
            S0 => dff_q_5
        );

    mux_inst_445: MUX2
        port map (
            O => mux_o_445,
            I0 => mux_o_441,
            I1 => mux_o_442,
            S0 => dff_q_4
        );

    mux_inst_446: MUX2
        port map (
            O => mux_o_446,
            I0 => mux_o_443,
            I1 => mux_o_444,
            S0 => dff_q_4
        );

    mux_inst_447: MUX2
        port map (
            O => doutb(31),
            I0 => mux_o_445,
            I1 => mux_o_446,
            S0 => dff_q_3
        );

end Behavioral; --systemRam

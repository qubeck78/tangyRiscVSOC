--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Thu Feb  8 12:48:04 2024

--Source file index table:
--file0 "\C:/Users/qubec/Documents/Development/ProjektyVHDL/TangNano20K/tangyRiscVSOC/tangyRiscVSOC/src/uartFiFo/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/Users/qubec/Documents/Development/ProjektyVHDL/TangNano20K/tangyRiscVSOC/tangyRiscVSOC/src/uartFiFo/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
cTb2kbtzurGWBtalgAEGL8KnfEJyqsTFeVBgUGUpa47Om/voE7x9R9GRyUrYP53C5Ra5N9e/jGLz
eVXN1oK7Aq8ZZslYFygFPE01GFBONuKtu2dkDFc7P6+bC60+cMVXVVDKpJQ4+146Smrb21lQbyYr
EnecTDhh7QEsmeMkK4tiiF2lhXfafXQwGcoJOPfyWOe6FslcI/z2/tSdEsInipDKe9m/cS5KGvWJ
+14XxrYZ60U3mToIl/xS1oQjgHGBEv6JJzrQ6t+2lNb9MjzDpbcEUzkoH8mQF6knDhG16ygRMZoF
wLSQiCtHMjCFFHXDEihy8cGBNXjWq7xIFjh04g==

`protect encoding=(enctype="base64", line_length=76, bytes=53808)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
ChHoT0gDTLSkiS7zdaxAh7rcVWfYYkH31otPn/eKzi18GeF1RcWI6ubsO4jovOVMrugsRHqKF0oH
W3D6MFtU1FDpp4nuiErTA/heHRYwh1lOhM8tHxZf+u8bPXjfrhuFzBzNsiLgEmeQH7/5/8zLrw1e
juxJqVM+Zxwdx7Ta+jgAYpkbwSJqfBt+RBeOe0pSiTH3R//iuQC7LqJ2RAgD6QTP9nw548ijIUj1
s0bn7FKD3cUPOVDl8SB20h1icUnXuEObtVQaWAZUh0EZqZtKtOopdofcVr1GH8Gx6gN9C8zDz4pQ
ZuxnwOczRjuZC12TGlTufj7JEmpGlg5wnoO4WJP8wc9arAi8Aja3iwY4w8jsddRL6j15Zc2WNHYa
7LM0vxYqTnuMgpwh2fOyQpuOwZB6sML4wPDo5zJcVC9IG8NuW5neyCrcD3u/VU2Dn6sYya4KDHs3
floa2AHRkqMBzE1EQyq9eDEfizAsgkCo6bsgK8YFtfkLEeolJOoEChahcbzhnbkZ5u6iDEZaSKm0
MASGO5d7nM7KU8CuuEdKxPi4yVDaZr5V420SwFByx5fnFnfKxC6LumOOg5fIxEwxWfy0Yhtw5jmG
RLPbsYx0j7xk3qseXuFlEwYtpxAi977FnqihB+pSn/B3U6ZKToQOqa+Dpe/uH3Jd7AZpdF7xzOlu
J18vL7t+HmC5MLyrE4EW4GUL6y5EtmIOw1r455MndMa7c2PLyRpa4R7NAosjZCqQyWeNhQBtq4jr
8hw19ntGXP1VQ3m9bycp5jbCNH2sQ3ANlKd0PXqyq+A3uKhWux+SamsBHOiMLj7eKxYTPnTqDBQ5
vHWyYTx6IbZex6hqw0z6z4GJen49Bv/6/abOQqXl2riF7RAXFfllj2myLr9MPoCSfjIIA5q9XuYr
1Ezjprureh6RQoteBRLqRNDy7ka+tij+VcfjmmIK7wVISX8hoJxTcDRvNsUz5J6WLPSAqNmJPFXV
BbpSKL4OXdeHzRfJwsR/vPZiebJRTPDqAYbz8GgopJH6Fk3MjWcOz9LdFen8qkAYCeMjGFo7ECaS
avJ2mtPi+rpzRQOoTdfpV29fm/nb+OQSraR8RFexUmuiAfuECJVaUYWIxA90lsb41ZyFtFTCyOG4
mUC3FU9Vd4wk+/sZQtUmyBDE6DohA/BgJuHqdfUgNub1Ny3anR6E9EitqmW+Z9bz95YHBuCbPNAI
v8H3JI/Nd+efDizLMZWO4RJ/riEsKXnhIrSxtinb2IoFv8VPLb8yOkuZrFvifT/vPRgHzgKLv4XR
23fm+b2lA0WgQY4aAW8Cj6+jyu4WWnMs3VI2io/vGaKhchog2PKCCLAIAqM+s3yiAJNXT8hS/rPR
J+fGF2CD9Mpe4a8WqHwRlEiLlHFVj8udsMVwJXYF4j3Kl243UZo7po4ZVqd72g73WDpSfXPimU0Z
pEaBFIH85WGrSCX99l1RkMHN4FEknQACqQH0s+VB6usTI+QfGF5SkKf1KqUu45cEjBIRifdo2Dh6
u3qLfeORiH8H7IBOhUsObnEwmslmFvcJYGl/wQXEX9KjhEJEet/W2539GkCaHtpS4dSreMaXxF88
wUyRgiSsqX0U55Foi0iqewLSAGgczhfLX0Tt9f1y2P0/kex9VCcWJD6IOGUTTal2XKUx7rsMkIab
jldqCmM83DTmyaYro6g9C/y9S9f46iHv0CoctMoQGbaLfaXOad57HkUucofHgzXPLw1p43S/k/9L
z30DngtsH9pxPa+aPTWUcVtFt+acIGA6pugd3+uty5eaYaB0LXCdECc3n3bkZC/oNNwfgazRGO80
i+MTNDV9EWOSVPz4FIBRGoHlttHuCoKPwDzFB21raiYRVCXy7Av9wn4+wevg8pi82Yc4q+dJpfbQ
tj+IWAnKP0tsYhOWRGGyfNb4RbxIcuohFv/mG1kvInyfUPmVI/9V3dS85Rbq+FEknXh9SvqevXwp
VEKAO5ckkY6UJYBNuP8n4gA8UG2FbwZT83y036M4JvGaz5drYv8JwfshekY9P71fuzkUhC4K0weQ
3Fw1wQQ1VxTDbWmgAJhi6SH6uDrkbbYuc89MdFma8qUU0lgy23DY1pPcPLkdzjeMvyblY7D/BzR6
gZWXj9I/Fk8NxvXcTldAKZZosJFcWFRSjp8ZSwn9MZpgFAdGB6RED3PnFfpaIdKvI3ua1WEsBWET
b6v0V3noFzTHuzfpKs69YXqNvEpp1yG1qcie+tUvpiop8hFlucwQgNxFGTQPEeFHCIErFg+P+6ke
HiRgplQTrR0VpME9W84HMpzur1QQ6JfgPbvhtfIwI7A+AIpNzI2gxrReMiOoouawWl7+HKI5tokh
zs3doTIB8IOXR4XzIN/OscbhlLFgtZskHzijXdteVWuioF34RqKVXRC2oU/x/lsn6pSqoTLBaw8Q
7V4ea556w04b78KVl1/RjHZujTM+WQwg/LAxAvT1l7iMlXal8duqeC1By8OJxtCfucSuKZXd/ug1
64t5C6E47AneYDuxCjvFE5FOiYlndYXkJUme75FgQtKGQxSNeeeVYPqMTOkpOgqYrn4++vr73xX/
vYLgQJ+v5XCQhQxms3bXrSmPrvcIfTn0uW0xHeszNvgtd9OzP63HpLwHwv50XJobLcJbD0Z4D1Q3
gBne8ijkhbu63i6ullSNSg0Qg1eldBMWO8mEAPHlhS8ssp1iGBKxNE/iyZjy2kAkZmBRvTBMOh9F
PxF5Yro4z6NrXkAceFUg1L535v6z+mkW3oLAeeQNQb3Moz06a0JAE/2Xm/fYL4Y5iyQa5b4he5i0
jSO7FqwlBILR87QGdmRGCLj5F24rIKozJSB2GG75Dr6lQrmTfhdwCsBNTrzgZ9Kq/X+C9/B/wxo+
In/VZg2XBeYEEiLBKmdkR+ZzNjOZ+am+giIeaKgm9lf9yLDFqr/3yI9xT2hAxIBxex0LehJOQuJ3
HdQwSqlJbUx7kdAk/opzZHzniDtiD+Yf3jvSaPIscWz8dzuN9JF44BXr9idQm73i87N65yzI82zh
ZaWte9Qi1+07EzYzUFHZJMCawwZqIKvMAf+ckOzIKSw/Fs8/Rhj4DSEW2yDEGEZgkXIHXL3NBCAN
2Ak60TaRfwqP1Nozej+lxapNX6jF9gAKwilo2aH+zyDgj6nIyO6YRelX/3FVc7mZA+NbHEjJz0QU
UHbwaN5s6zrcGB22AmJmLq0zjue2H1AYGV2V928gZqV3ICu7KmxsgsAbg274YQyJvQCc99VMpM+n
vy+03bgl1JJRVmmifHLgLWax94cZTErJzkjNeLbAZERzSOiVsaASIPaENhkPVLdAz6geTwlqeO1P
cRAJDZSISVN/3nCCphOBGZHCA0utlJjZ9F637R3QCfORDG7FvGmTGTouDZ8bzDzqWvT4X1VlxRyV
IxS82AHOJe7X3d7wAUfIvJkZKsa+/s0h/PC9ojQMBvMRiczYGPc9WTgNv7uIqviklL0yxtUQzTv2
tCxA8r2/GkORcuKXI5nmgQT6O7b6infabr6+ido7qIB0RJ7rXtCCCQviQ2BvnchzAsaky79JhD1y
tdGoqqNvyynG6xgE8E8xy3jez+Vkx5lctR+RXxkNCth+E0GX2kng4+x/+KHGv5miqx74wiBdoazD
z2pB4H8Y4zQxKR7yIN6ruotDANbk/bYEI5W/abA9ivKuO/eWia7Av3flkSYbgBFs4R5A5eKJkk4S
rVoPVBwYAwYDZQ9xgreW4JKPbpMEEA7cpD5/XdETaokDpuDHhz0x2l9O1BTgwWeI/ojVGJ1BmZ1i
LDO1AXPu7A0UvEQSdSMz//9DYUMw6Qz2/sFSBiRMYeaH3rKLymqBALZrCwphMmnRji9JtuFemUih
p9ZmsVIllub0o4JlZufTGxm/9HzywerpNfiwZTa/p0Z1WrAcNObgKkOPTmzN2d/8f2WCXmdsSsjb
VsYIrpN8T8Eajv18frJIX01/BDjoH/bDOdktpgg8p1FL/imSy9tSuhS2NUl6Qf9eRr5vy5//IWsW
3ttEImczc4q+T1J95dWL2zG1e+3sIxItW/vVkGyDLwK6g0nk4FUm735gUaJmhGeJIuiGg5vKh+1S
GYjOy/SejTVioSjvddlnkorY9KedRy+FUJqemotE10iLtS4K3CPhFeAWPAIg30bFkGAICQKWYaeO
16mH03YdXWonWTcj2Np+pPQPcJaUZysxT6wl/cOIdwlFoWsSXLypwlj6BZTGeQaSdUCntCBSm1/+
lzyhNN0ay8UFhnvKARChRa6BGNRAr1hk13DrkB6XemHXY4kUdGOvgnv4otcjF6y49Ir8KBcjx99j
RIKLdDHVL0bq3CUFq94T41yhSYBNVfHdvwDKRHTuvR8ay8xeh72d1tlzsXVsi1Vki9ZRwQ/2BsK8
6U7fyZWhvflwN29Pp5UXk6P6Vee0yi8vHWvVB3sXonyf6imxLWK0/Z6YX2Nc9c65KgH1zWMQowTI
IV1TuyTxNCOFeAl1GmF47VRXj9ZKkwTZYl1GQTQU3zQ4ihybuRF3p2FSPF25okXy8fqBd3SPHOgF
TotaIt2I3aJAULVdlcFaWVDl1fw5+pom9TEAZaTkfNYqmBigIQ4xUvVAYegen1DcXpaphuTr5KR8
9tBkuYSkbDcAetbbbGCjLV6GQcFv+m8Iz1UN1tLc7iMGRrrXm7CneYxL+I3+HepysWtXZhcfUYZF
z0zx4X9+lh3XsnuKn5HKLDa8EokBOsCVwAxykjBUJgh12VXknjSdQCRlZPnQJEOkv+9Ym7PqapyQ
RIMglPUQJY93VPcOlUUq8Sqg4uA2Q2yYLnDSKJ7ubWx+m2iyYSxO00Y5ojq9InITyrMJdEaLbppx
hEDbmFarMiuam8ZTUlwCllbMxIOrViTbJDeDJvnICuixYIFZQmi6aZk+lSJqHPOvv3/cnY+NJDJl
axv8cl8Gkwuh8G8RrOrkKDdGlsXRYn9mTzXkxI0sxfdbrMwVNWK5e4fU6rBBzbgdkqd2fM0fuks+
PTb0WDwWjHr0bOMwRKtLD9k3FOjT1nVLzK1/BOHOla4GDnGXil8d+ndK/Rir351gf6EgB53FJf/x
Vq9BQDmhugeE/XK0IhJ+06bbLznDifDQvHePUwZg6qREjMUMi8JGQ13JFPUGpUzroc8JSIrkHJ5/
bbIhUOz6SZhFERYXBYQUaTHgNTPgLKxj9CRqiCyhhG8nqmy/ftY3n/KHW8gUYdfL0ybmlI2QP5J0
dwhR5ExHNgpVkjra4kziCK7z1C46WYTmRHEgUluhNSS42Vst0rEtKlWQXbqLDSsy0OuJLlvJZ1t3
0rDKymNFO4uML//QSsS7g/IVPFRlv88Ezuh8xt84CS+4M6T1TH7d0nNpw4XFDRbh6C32mhvgAEQI
/SacG3zG5Fax0NL09AuVVdHod7g/Arb524u7zDroUTXVh0muEZFEcLDijiln0BbBIu5mMt2Zbsq7
+JcUEg9Z0gJYdZqsp7rJ+nIu4F8zNTLcBUTVOEwlbfZ4TZH+KqnJ6VN99e2rrB1lRZcYPJYNbhRN
GlL7f5mq64dg+q9XsO/dwHOJ3JevIvVSMD+D5pB58Jdb4mypuGiUpkj2SdO1uR7LfdUSBkjVdbUe
kEAnpXNCTZubKotOyYxzb4jtykFRefsWjvqYesjzt4vw80aKdVDzXpjMUMajbKEeI+eln16sK72Q
k/mD+a4J6UeMwqyGKIxqtOY6GIj/RU6i5dh/5iqDEz3uNkujP45AsFjs1ebUcvK82bQAdeFveQo3
OYfZILo6//KDh8F7xc1kdLlwla3SJuOxv+VOfwoGml7ahW1CLugHMZ/9bbry29gOnJaTpmEDCJmd
gBM1ThSm5KWCMDO7R2PcnH9dGYo6bhhQvgo4Bad02jmiX+KHR/y/40VRWYWtY25lNhfaTq/PmXpt
yupUDSi5gMMfye8NBKLpimI4MTuz3xPp3hSTwX7zci0vOe+8wZP4o0eMeYaWGUWcBhXhn/IrwvBG
TAQkK6CjI6A26XXQ2WfnajR1rsk3gtoMHBj1XIqSngW0u1kyL8ATVUuyxoMD1Ye8L5IoIepEwLeF
aYwBfGkYDOLMHvZeNcCAImeGxK1vYARmrhhqpyDnQV33tOvQ6EZS6wxutJf5VSX7UvbJqTmTa/zj
XV5hCS6F/YEhOIEWXG5B659GjwkpuqqOzkn5CpNFCBYGtreyL+6+Q4lmEtmxwqS/2ZvjsJEKgEzs
aWXLomFmEoVeG/4GaW5yp2e28uurmX1lfUEp8kwqlhWNE5VWqtkXfCaT5OJzMjmcCggityJrXm93
Y35Q0ZiXBnx2JyxumYhVe8Z03JeUzwi4JXcu7k2sxSSy4qrHL5HL9ffpty+zWWqvpdHZubFm7XkG
9tyyLaaGA76citSsvZQoO3NOUcCglX6umYW+sIugoY9V1ouFsrSdwX2I2Pe541LfhtwhopdWGE9n
wUHZl/WuYxPPhYZm78/YlX6qF6D7adk0N+SE8HbK/dRUO/OBK1cyp2N3NvACMVWIxDSIF9C5JJTL
6E79SBd8vd2/lK75EhOxcoewDaobQes0SWQDEhkxeE+DvsTfkUTouiPv9omIR9EMgTiw5XuPuDz+
bZDuptOWGmWDzg/kHbblEG2zjQl8QCHZ2Rf0J3QhkRVf34XIv4YkzhGZuzG/5TDfAxZXfv6Uhdhr
RDQmZ1zvSkAi54jXZAOPmD2X3ulSDz4B7stjnNV+C0+4gPTyWkqAjdCer9NSpRg4GCkbmKnoWjzb
VhwWlFXRvTLM2eh7+jj7/IOCUxVsbO3c5or4WFf6fV6x5mzhpTJ+fOAvml1rV2JE/g+KEwGaOLwF
dL6XKl8gzEILC/eg9R+if2aDtY/YZlXq74BRYI3DGVJZi97OX3G2QY+hRiuea3FW8839NWHDxouh
Eflr9pLas9ebUkwh+7nwoIbLwqQdLP+AXEUp+6ghKlUdXHZ4xDRPEyO5G/w10rrVrF5nHvZCuUNi
8UWH+B7zFUnc0x84DltZQsUDrWrbWpQ2lHZI01/WL2NwbGfqjuDJxVuhrhXKXodtYZVP128iJAgh
VvATJ8k+GoBGHFhsahnd3Icubken9pG4p3THExdQpSqca/d8emwKv9XRfFj+bChY9EijjAcreHd/
eLoL4vPRXqDecWbRowduQWJ6peaIsTr5UzBR5q6aoFM8+PqhMJVhOKrYkm4SHkqyfFUKg7WxrXcG
+kdgnsux10bbH3gAw6A1Rr0ivQn5hxitO8DRtKbj6MXndrrG70Fhr9hkkm1daqwXE7eBae2D9mTs
avjKlNASRUeZAA2Cq5D23geE77Xe87eaChlhmFZI08Iv9onXl0xcbfd3LiN5QuwswnaxZ/ITprBh
/y4b8Im8rM2uLRtxQuP8gp0htJWUUd6+DzI1czAKHLGhSKGeCG4r3xBjoYg/Nhu0TjWIlz/Tx0rU
faa1tNUyRH4ubWcPsTiTqgdSBXcXTusrBU4XObAIGCjLQ8PsBImcfM9Z4HuGJBGr5jQM39AQwVPH
sjkWgGl2ByB50lXlWYnU9Ik4zef4RNpAiLksA+rDFPhbQvUKNgLNHI2CaWKMwEvOL3KLevgvqILS
Uxv1F65z088eDU5OnrnPFsm64Z3AOIW/TE+uasRbpNdODsxs+gCnw3m51UB/3i7TuOwiCLQzwnRU
zQ8u69J/6qAju1GRvua/j0C4oGe71ZBtumr7wFSfqjqBm/I1baHQGFLCf44hSRqXQPK17Cys4Spj
C9CqT0XfH+LIGt0cU0v8A2OIyyedLw5Pnn45FFvE/jQqW86z5zqaTvLnyvZx+BAo3ggwYl4/uHsO
Ob44wjnIquc7g5YLxnExMQrn4oLPo9HDRuxGzMno7bO39/8VyNGSNychwgpYnUyP2PJmccIrjZoc
jsrQ6viy8rUQn/SojCEmuQ2/4d41cFNXv/k9Cj9oZSGIZNLUoXeYfAqe020vtReHicDBZYgk3RCX
PrmBK7dI8HnsTyAFCJMQqHrvUjT8NgNvqVZ+XfEfEyjgHKSfuZd5Dyey/J393WdMstQOWUBnBuEO
7Fha6Ge1wMTgNkFAnYQ1/uqq3KpIVBvhxORk28NJORSqHcTTckE3F0S8uX/g05uRxzYjOAYONDYq
bvCf1EHrXEsCjhv8UVX3zqe+7gIJ6PkS1IPOo+5+uYAfbThTL6kcUga29nVROi5fgy+1yRECIWl/
IrKKRfxyC5k+9IskmeMGoGiS6UXpyXIj8RArLAlqlNs/1WDbG0VtE+wc5YwkdAws60b2rruT4+Dj
P6QtM2j5Xtsf8pC1Fxntm1Fx/QgIOL7C6vOHwwnQD6NQpCip+b0gpdY+/I7HZB/t1sBArOLH8E/U
S5S6kkcrNHjX6z0GwQgLzvN3y7f/mENyBA8mjJMxIpJtkJpwdUCg+7gG4VNs9urSeG2vBM1thcmw
zv+JfrGV7o8oIdGDJZTJa7t2tNKMmgXukKTmwpeG78WbBcUt/cyImYa1VpeuRGIgiJw3yWLgMoc1
g6XhqczGRHlK4SMZtbrbnfpaLZfCH/zyChicheXH7MHmTKB/dBSGo5kpINVi1Ov/wRn4caKCwB7O
siuoXzSfZ2G7FslyQzbZpdMpBKFjjMheipnzD4FrST+anaBC1pKtqatYazuOjAPvbVBI2WsPsAPS
y8z1iLiGdyXAPUHN3NlZS+maWXclr/LxGTkNt6/Ezm5cJ9uiwfTGuChZLDMpJ0uA0TyAUkyCauin
NXWcEQykBhGL5/Xujj/8Tb9o5Qpz9hgz2ic6EtrYanp/c/Nx7ntRHx7FgyuDQts9nrXPOr53FWTn
4leOztNGtAfMIz5UT86DzuFz29OvsqbIl++Qii4QOLZCiJdiKoHnhDlUg9YAFAklzxw9nYd/44QL
8zr3exERXbPgrCJ5xdlcwe2dsl7NBvzLY941e8NTLRgYREXqpWjuPLnaUkCUFFYo1qf3tG4mSXlz
8aBeCV8lhiioVa+pUcm6QluXBKZJFkPv8sr3pYLol0ysqfYf8DI0PsoRDQWFKKlzx7FLLKc2d9GW
STI8EG0is4UMAUdFq4sEi8HVnQyefMYbV4QXr2xzkR+ag/I658Jd4it3ErqLj5idAqCBS3w1dnkQ
8J1OB2RZNGvzYmvX6J41aoHsnSjoi5aAom+E7K461ssFDJ4oAbsYrdDI5tuheIcW86dk/Ouo0dPK
3ssLojwD7KE0Yp2ahcnGEJOYcBIHajVjZ+6yQFfkEhLcXoujOR0F5wzTMdr7uV+MG9zRBhFMPxpX
S9oAmqgt1CPrvCPiUa/5AmgCouMn2Cbuiqy1ppbDaiNPhdCxVgGTfi5TTWAz3c2x4F7qCnWrK550
7+MRscMtV9s8TvXnXwNMZrCnPv0+bpGR5GMTPiADxg55uKHyI5zwNmdYFqc60pAuF563c8MryQlc
MPX8tsNSdVFttWbyZTK3CJfyS1WR09bcYSjv2wIcECwOZ724KeBL+jHjC7uockS1tcJfYqCcxVdE
L6rHNEVrIVSzXTnrLsX1gRUC0BjisM1b1SsUgXVcl6xDOlrl9UdGSurgYKStpc1b/aVifr4PnqF0
7Gv4AKezbt54BhkfiugOyUEnIJisciFJHFxXMcTjRw3TW9CeXSbMhzrWmz/umNhBJxXJ+2v3tigJ
SBrljxNGNk03W8U0OZUQhRJLFud3ZYTsLuWm8zubxpgi1Zn45uVRwinV/KOAcrRjEFDP8uBWjX5t
r944rSqq7z7AHtEq3EizbycxcKz5lMqeS0xhAv3ZKV2MwEStezs8DUvWsPGyB5hZ9qzq1KafUTTh
5peBgazoqhwLtjNxsyQylcL7ZtM0yKefK9CT0GySq3j17YCkYt8CvP3LGCjpx11u79xDQ+cPOOwp
GpbkTd8+m6Mh52FgF413eUvR9WfC5m3AMoNseQwpRGu2SIFk7evek5OguS0JO++zTJzfWTIa2l3j
5Xor9SZQESf5lFf66mrkpq9CCasR9lWKFKkVazZ0dRjNIT7U92+75VpPK/eK6+YThpIWWakiH0jc
N8BypIsYrMD8xV3E3W8BYzHYHvePn/lhk4rsMEiKplT3GiYZ3thF+hXlmz07PKlXyJb7XoaC1mVX
9qAiNgdu4p6rCofWNObvvvrnvr07lHtIH+aCDJU6InrCh3mmUWcBmvTNA4dwtOJ+vFfV0wuq7ivE
esNHlJ9hFaARFh7cJx7VUKK7Pz2E0t1xyCf6qVwJ/Cv+6rOm/LjFvckuhyK07g/a1WHeyagTZhF9
fO3N7yu91uGYb79rasPdPD2aDFOpIqdsuolIddZd7M5p/UjOb+GbJWcckpqOcfb13LiQDu7O/y6P
PrJPnDAYhQWxeay/XR5CyX1IbNoyl/hZF72dJsRQuKZcVgcXvaiLxjFLPxIPkfajGYsYxIR6/KOA
qicTH2ZegatbQE/K1TRPDQ+Q4FXn+LSBdMPVN2erUIfdHLj0ltpSg5DKs3i0x2pEVqeDSgN2/5zK
gebr3hY+TpUx4zCPfTQImo+GKdWD/e45rBKddni8q7dWjeR3OXm62SP473isMGupV2pxVtLR/kQc
Eoe/4PZVJEsL5uVosh9wTXxB1QMO95h4CE9DcVDHDroeA8glB8aVyfieiocUy2fU9fAj93Ejy2z6
RiqlKE5rj8wAnb8jbTIx2qiJrFgP2Zdr14oCCLRV6Y83yMz+aOlkUBm/W+KufsQB7yBBnvX0vwmp
rcGOrtap4ibdfMVr1JffBNfOwsJiNtQrcBD7dC8vHLNtvWggxICcBD5ijX5yCuWQDyXjsYXReFTj
XsxtijPsc5yFB5qsqM9WoJznEE6XuBRZ3VsCsjumlK3I3/0CTUsRqE8UCcFsgsHscVqsyn+cEMRD
nwCxFzhmzkQ6hZ/NAEUT+EG17PuypQT4fiAi0DZxBmmbab0yfhdtWo3oMfedKv8qvAXaGhmp+CUs
RiaDOCn1iAHVBD1aInn1GWZXyT60Xjst5n9VIUITEyaZzKzdmTnAqgIvsNjb8p7Xcx8LpCH3PvOf
L6FXdQ3Xv/hiJ9GOTcJbeuoqPMjNQb9gfu1kvTYK49XIiPyrvBnyuqWIKUhLzca0sb+4HvcinRVp
6uU5xQsLbETL5rugNTue2CvRG7ZDnM1l8PI6HBjrNNizoc/K0SLSYZG2tOaRWEcmGG8qrJbOy+GM
F+GkvsA4M+a76shsgPP9542YHSa22SUiAJljgscBVu1hyHegTK0pXLzD2UBd9IgUtVydey2dIT8+
1iFOwiQZfNnJPhVWqBb6y3CCJLNiuJZ+JMyQZTdI2O5gXaxitsSSx6CoGzN8XqxHFsU9fK4d8L/j
rpR6hc0GQmBpzPgQ/e4O0ng+u981DiujhTIQxAMk+UmQrt7UMiGBL1ykrPJsrYMJnDdYaAcD3iMB
Gj/idUTcPiD1Rb+fWqvVqRjNwfaPkQFgj7o2PUMNjXNro4iNhHMycXTL2zGBRQXibzf1UXLgjOdG
I5crkcHTfhr7inKsxeu8cd3wQtT2qOdV0j6FobQ5CtZXYMf7316fOh7ntCsogd+VhKw7N7YFjZGm
+XXarIJfkrbhcLYofcSSC2HvPLXtRpDOYIiajug2icXi+YhstD77d0ZjwtixQHTOcvyNGRs4QqFN
svm25vJnu8z/yLEssooj7RAExp/e5LepJyA8OTjc/oDnuFah6l+DsJbOGSh1QVGWzAPt4MRRA9T/
1aArzq6Ad07Z/p0jlk4E1w7SHSRsOkpuwT3Qv+0R012DgUoiyrTgbOLV7abacpd569iaTauNeEfO
nhnFR5UIBysX20BKo9nLNn9WuUx6hxO8b1YcKjpvE4SGz88/i0P76Y52OmUw73gGIGfSb1MtMtKR
MJvMCP7uW6ute/+RDfw6nHSh9LQn8utJdduXIXXvAMf4rjDaxaTkLV2DvSGzLy1XlwJA9ssTGD0Q
KZxEnEQYVxPlmymi72XDtP13/CWJp4IYnrdj84bs2Y3GsTlS5ePDvFDCU77J3fp7mAgaQou/cq+8
6y7eVXHhnL+ML+WW9Ngq83OimP6ZOD8NzKKNQ0mBR71fs7pH1OJoBnq6JkVaz7c8sRtukcpeluaT
eTeqjPse+kp7HmJx3UgNk15KhOAm+8mbuUFDhKmepWD9OTtAyNb3mGaat0sjZ2Tp8Dz+DRzQ/geU
lXYHDvNwLlR+qc+5/F/MPNL0RvlRuTNnox5bKRR2aJvQoCZX/dpet7G7hnM/NG6cFxfsqEMZUnuM
XMXbQjBgBdB7yFukc/bmERbs6MblvMQ773eEqqx+Ha9g9A8BwdgXpc9TwP+GplAMgvpcf30gSOjn
SwHXYGg7j+hDIlno8nFx+Rup+taCXvdZpB74Xn2EyGFY1pRjwrvTVnzhZUEui8WRg8YyP1uNMbSV
vR0HMlPtd75YEGp/TnmU3ELAtp13+2kQ3jQ0+FAM5ez5367vXj9fUd5R1dwMZVZM/gxQEUZkP2XO
pEYNZyC+BHQuoLPWS24eoEInM9UIlXL+LENByiejDTyCuTG8lSVS6XGYU9dpl+rjl0Dr92koIw31
NeMOAR3ZAuDZ68xymQmftEseY545LUEWqUaSBb0r+tF7YmOvGCBLjVrNrrvkPetNBfFEMHrNm+Km
H9nWkX8T7YdiWTZPXMyHB4wFQAxIPst+CzF0r6aBgJez9NfxNc4sviQjhSzVHst8PEe92Sba3PgP
qEnkLsd1gVL47n8RepwTNGeEIGto+tilfW9Q4XePQdQRZ75Ac2/8sz/XAJvnCdBd9RCR7sVyIwNK
8x/UPDgjKUYFbvlvirTltZfvhiQPGHZ/uQZYkVrXZ0vcmqetXiQAB8LoauTkM3xz+ZQWkJtfDRNX
plB1Vp8HagaWWQlGEo688RzxMaogQF7d2IsFiVhyNzw+sMwtNKI6h8be/zuENc+Q5waDuJgG5cDO
l+mIxAYOdffACAdwTpV8qqK6lKaRlSE0FCk1wu89pI335FS4Sc57NCPUoyKaPcgdWWu0bv1TtQB0
ZP+OV9myqRAriMOTGgjCySf3YHNgf86KytkM8NP144IboHINLFPbVorh+q89vP5YqyQMt1ZyIeiE
00T5TFoDanhCC/SaUrhU3VB5F3RWnn5T9sz8de5jiXBqEiPLMRoBTGcVa9yzcjIZtCyuUKsIEZx+
OV7gUnv5EEp1UCcXVj0WnVmslcHOBEwS157L2aQ0e8OPgOtJL3ca+IoWI98pAPQMF51aMK/H2ecL
MEnuC+ei/lwibx/KxEY/WE+Nvl9j1UYcqKcO+SWkoPCje8kU+l7VDfLzAaqtAQ2+kbvwgkCaNX8N
iXlnH9asp6lHgPSXu9/palZPOzvnGsXKsPOS8+tfOBUpUbJ5XAkEoB9j2NU9iHfP6zvR1rTbSbDI
LNgmbncvmrdIL6gWC+goRwxRuuNco+m6DDhYdbhgrmlDuzamS5ldrOWVOhFexEvidDHZM+shGTh7
54IkiRNEKY+XShFFypu0aCpmOgHP+JPkWZgeDZnn0rjkstHUQixl1v5hCvUS6MsWYE9bbSTAyyAE
tdq3n9UiYOUlclGBjEqKHCE4xia/aP++3Myg7iSTCDqDBm7m8r5/HhOqrEvgKhBMJRjevAtn+4/r
hvhF6NORxR7uX1zYVFKr7Hc3goJwRZ6RYZL3NfWpVUWTMAMdewZ/dTe5AtqYtGmH0iHzPTcq/jy8
0Dy47qUH2wQw2QjYsjqPqtFHS+T3QxyZsUct7/V1ftrYuMYuBr3oHzF/2qa7SAbe3vd3xr0tj7fW
oChpI+cbBW3VElVSgdGWNxrytFF6bshV9p87+2JhaWotK0fsXi8ISfn5nBlqMfxEsfxZAFk9fhzT
OeOtXZYP3ObYZsMuhlRpSX7XtohGym+7/7PJ5xK24BT2yQx04zr2dQH+YIa6BHaxw5UudXFBHkcv
T+x3Jvm5YtXqvvCHuJDBdPMu1hAp7uKv/hUwFxOFvxBmj0LTHHDkJaI9q8Ou/hlXSPRLqa2Nlsle
GkuZuj9K9aWurbMCa/VGtBQfBiXY28xDwXoIgGAPWfcvzZeWQ5fe2qoiFlWuJvsYNcHPCSvz/s0q
m/6ud4PHSc4K1CJv5NHFGYIbLH0QFhCODTQQQsi55aGxcVfAcw/cx7c1hX82HkO7XECZwzef8ANn
0fhUWcO45SvtkihywpH4LvgQnPJm4zuuYwWS6srE4qlkzrsz20QhLWOxiDb5O2fzt+FsESutfftT
UntQiPnmxCZr9YiaLha+aTVO9XER14mGhJwsLi7kFfKzbgSwxSPETaaA4uFZ5GQT9vEcDaLA52ZA
Pc8BcJKV1oGHjb3A3nvvDZMKSbirVy9s+ICMzb+Xi5S9yVWyFiNQH26jsy8XLhtbUobnfHIKI6Zs
ZgAv6RDXsyTQ8JUH1at2nMqTjLiwodu5eVHQrg1NVxVPGdHZTZI3E64uDlbn37ZgXmE4FXnajs1Q
QDWQawD4wF3/6v/m6JcZmlzHdLwMlFDi/4suCig0FwnrJfJpa8FJIHoIYbHARvQvAJsPEAcLFBQh
IeUS7fUhd4IZwLvH5fDB91pG3dD752wrpqhQTQGp/mGvp8HTFAJIJyISaWamf8FLS5pXjSYJOyNR
k6CPA8fAn4DxlxPH3TuWF+B57o28jtsziVb5R0O1N8zEdeUmypKAKBgbI+9pGTWTgF54SVI9aPjf
VRbVMBKBDnEBqQPzXjDXHJ+p2aCmATLFMkjTJA5etGSPjbGFj5LO20IiK2o82WHnYFdJoqx33Nmv
9K2Ck2oiiv/78Ax1htSVfBgE/5wNNKjOuwW+uPnKZMAm9BssmpSH3hxGaMS2poaysiphAxA1IzX1
lY0xFL8redx2n73h8BPKGzYoMjd4y+R7flJ/MVEdTh7qtwtLJVAnqhBNNJznx3Uy5qj0z6ygjveL
pEqfXiH6mS+6NWZY2n3SbUAPbm5X366gIW1yo5C4nW3+QxwSKaH9sQPRoxXZ5OfOPXBdJD8653Mu
4HXfHtTOxddSRsBUy3y7HNW+jrmDy+lGE1Vri292AZbb2jifbePp9eEuE2bMMbARzzOagHW/4udc
XdAiWvCupZo5qGCxpB10n2vZcv8BeYwiKr4wbkLGbUyZtyO29oHFZD4ESQl4+lKBjgtXmkuZ3hAb
28Dltq6a/OMBKTwjbr8YXjyUtb/vcmJBos/g14cz6vnfsm/VrIP276fiv/dzbGYlXLXY5SFnX7w3
BQfm2uYvBBiCCbOucbgQB2xpCFsdKoDOsV8YJk4CV6gi7i2lcDGphpEzJdkhI9NX/OwtyxMDE0Tx
OhUYN7G5uJUnDDGcW23+cOix5N+vOcAgmsvD0txgLrLFntwR+6PcYK8MA+iZsdvuMi/DsumvIyJp
qu02pqO55DRE+50E+oRvpAXdvgCkiT//nS7GCP8+ev7857FyM+B7DMwSsiUvuagNITc8BmAwFy5O
FqwkCkt1WTfiXGjDpjWBHORnZiWtYDQh65h5UO3NcbHPvEEaqiGHf/reBGbHF0rZxrSiq1zGsmSJ
6Ll0fNYTa+L89KErWiPfaGIHmtxHOeL2WZ+2s9I+kVqu9xsPq38v7MWutYtlVmNDC1+zMJ03s4Mj
hbAwiP1BdyNJKiudznlMoDq6H0M3suPOT+Lc3XQQZRJKZpC7JMMNmNRHN8JYleCVYs3B9hNjINFF
5N+vL0oLVVOw/yb2lRpEYijZB0AC4gg6BLnGcxIsbyckKyz1fJXrFAKu8MP+vV+bIdX9puVE6LSw
eqIGzcxSGm1enbMVN7kD93/4frgMCU8diozx8VF18AASbTY2Izk/RdpeZ1qnzk4SOCv8VcmEg3ss
vI7UWf3onErVEW+UrrCBZKjcAWCW7y6YUqnWKqV1zB6gXFVv5tvba5P7i3baPSMTw4GgpKNIDUp3
cXguQRWqgdnB0oV5cgmHVH/YHE1wOah49iDqykVQPibP/ErgachFouTc67RYNFKBIPXsH7ryRPtH
exNZaxttLRPqANefI8CumCK5aWMU3ZIIJYxLwviEMlX0063NkZMUUb/C7iM5SsxmZzqFRjVnvroo
xUEBTV6bpacgyRXAPgu9jjwqXQTCUnENG/867X7Wn51Byoeha6H17lpAhQ079nDF4gRS1Vrrr6MA
YsvI5wu9zmqVLWBjKDHgdos7x+ZkCNs/3/P3hwnKb4gPrAiO0k3WFft7unYkXQERQ/Ji0qmlvrgz
x0zfoLe8ftXM+D7SkpeQwBloawIQgy/JJmkU9EHKPYwbB7COkKBR5YeMEBDu/Wlkz4AFdEQeKR6m
qiu30cA+vQi9BfKbN8tC5jL37eGEBK4DhH80ZfrprOudkRbnOJQx/wZTCbc/H9M8gPVDki3lAsyW
w8DJYx3CsElA7FaZKd9nEg2l5eNas1ZBr2IZClRwX2Ug1XfCEQ7mgZdAYLoehameoEjEG4K3QsIT
5nMVd2NiXcmV/cAhkvTzG9VoakJS7AcLvMkKKRzMNIJC4yDdnoCEPaSJWjP6jBb1SL3ELJ21jVKM
5aCqrDm65ryANGxEiG9hTcc1bmxvS6UB8BKXL2NSoPhbJtSWiEoAn+fOIiaprzyyCELmxXPRr15D
J/kU3crcQ0W5H0Vr3QVI1Ydb/u/kgxgnHittKo+QF4Xl0Dq/Lvn0A55rbLJCaRyhghaYCqeM64VX
K+a8TECJLsNzkCh46c5/mJ+FEZYvre+iaPMIWV32bx7wY86UxhEJDhDurCHlm36bmbK0mS/+Qiuu
HOk5Rfa1HdrxAN90/UCpK7dS8CDV9OZfSLuuwC/xn9TCYMYHXol96aw8fPnAPAcxwXblX9I/HxK1
SnHxj+aFvLtNCGuy6RT0BvieGzlPzWmSj+aNUuygDw8FlFJIRlx5Zm5a50a9MKkLIrytcJ4GHNZf
Wcjs1y738sOSNYfwr/+Aw4/pjb5OAK2k/Twzke97DDQzhFhzqU6/dkg60sSy+MF3i3Qk6uhurOHl
NiJxL7lruse2fek5be+XtP54OydZfEZPVddTlwpLjowE39NwfL6cG4pCwegTRP7+xZ0rviP36al/
ln8W5Hvy4bPoxqxMLwHCk7w9qiGUfZ4Nh/dGvwyWewbyJHh0ryLBhXaQD+U3C1Zna73f6MNf41WB
P7j6KnRimpn7vROM7Hia/Q1lwe8dYICR7bv0YmoinEBKtJgHdLr5jJMTmX4rcDS9Rkz8p/myCD5C
iAVQfQtgOZ16Y88IOf0wBD7C/14YYVHAug7hndLEuhD3MWLhdC1bwfdNW4d1l4PCh21fh9NEbOcs
9NDGw9SYr7uUccE1T372/fnDa+E1J9qSmJhfrvWwFXfXFA5k1FkI5sXEC8QkpmV6iTMAulcT6GsM
fVaEdrSXhjsW9gMKNf+6nEUaBoZEfFFKNtmLN8zzDbR9fQ70syQEoXJFfBYqGi3SJ6OORBOQ4DxS
xsGEOZA7HWGqULL5shUIIylSIrBN8JoZ9z8wbDQaOwurdpIAnQiPVd2lYFgiYuc79Hb9WffiCavG
n6U+UP5K0CC2zWh35gQ3CpkPNeXqMXsqr9ksgP7rAS8qrGOO/vIDPpbJE77KBUTVCuCnWq3DMAIx
BFjG5VtKY14ShlAjtzT7HEutIHtOewheRZp3U+XQseFdhzBW82sonzqbf4gS2a0asR1oSeRVqWGE
FltUYfjrmWeQoY6WnmmvA1CiCAcqBgUCuDDf+TuwRExMipsbTtOL0ASxxF1xHTnGtI1VrPqD3AkG
xWZSHOgx2hwYAw5bZVM7dHj5E/q/Pb2h4eap5cCT1bppwOlYFIsWFkSQrrnaibw4krC+MIY9a6Wu
xrCJ+eN+lIXc1vI8mEV+aLzXlY4A+EBjJWi6nhwhAb2TgSVkZ4MSUBfW78fzT6BbnILdElbHGHW+
qcDX8t+RYDJLmgurg8FkUmBo4zf5nGcq0q6Mf0YluN4vaQVlgx6kr6H2BxPDenRgsSyPJKBHBAjA
YWrq3WORWSZbYH72S+pKv910ttq2odRSfmoLpBaK7nep1ZkAWlVC6x4aGy69utEdNt4312R9YHbA
y20Y+md/Ufb4agj2OlaXsyHLR2sXVjap/gH3k4PHOMST8D8PC/+1PyYhvXMGuR15vVXOWW7BbliJ
JepuzTHxGHXhcZrK1ItTRk+Iq/YmuYV52A5263VrciEERMBa2hhBtGGtI/8AswZBslOq0lUjKaLo
JO9T0JAhljUcwhGhWl0HBHCQO8sjt9nonvpyQ1jiaqWTFYjy2Zrf56fO9nReqQFV9APDmAbg19WK
nO3quUPC1yfBqNpqirKjKAikp1jXc7rpUXa3gjHS3P1iRgTvIu0sTdhZDncPFTiZbzBLs+z4sZ3u
K9BWmvoPD3/MS3/uzM2yPmCWcqslEN9PbRkkjE4CvZUkmY0tlAlIf6pB3GTbVbvRenhxVfD0D6CH
K6UfNUB/7VSOPELICrizrkX+vj8Hds7hOxqYZAWY6P35QvwiuSgptra/5HB0bTtyWapN36t+iQqy
w9KG+Fe0n7T6G3w9J591NyyWKYMgro+rbiqMSUd+YIdXJMdmIzV+x3F3i+AwZu3b04IukKwLufuJ
tgt/vuj9kBuuWdHVAXpBztsYPB8XaOxoDhBDQWjI/gyCPrcNCBEBRNEXjs5JbCIiwXxBMYdjBEfs
NThvDeotZfkx5DghDRXmXaOmcdBguz9hOLOWfK4fFQXNR5VSZfpEbarkzO1L/3WjvGqJOkvGtjz9
yF3kc8/6Zw1LLL7rIypwr2/NTDxffB9ALpB6q0Q0GSR6aaxAzNVNv4oDEcUDjE8dvOetIj63I4ho
M/m6QuQGGh1GuSB5UOKxEylnEjmbNaGR9Ct61qhZe8lN0Q8h9J7ky09+qVPJuxPIVk9zwGu6IuFe
RmHOgihu85LxTkKeXDHiUUqBdUqYYbnFVQNHWB7gd2hMov+aAU+jMP1LOYTOXRBrmwgg80NZUwAd
S+pUwlNfTWRFxWtiWyageTUC8GVL9O2nIvA80t8sRttSQX4LreRMguX3jPfSkudS7v9ZMohkcFkk
XD38Aqxg5OdacO8JXjIUHfoDDX9ObSPGBQxdMO4eg1cmtFhPuSkqUhJzUsCshmeCEzbQ1USlNgin
8ExMkSSqNzEe7+wpEul3ASVHpIaAVfTySuU1n+59OoNlkI5kV49aHYlofekC/HswAC8+67uyeqkC
DTF16pXxtMZSp4la8oZP5lfF+gxoJBZedlO5poRQ4XF+Nb4h5q/qlEnap6gsImpdGTD0R/B3w8xZ
sb3GnhLLc11ylT+ZYkkZZpEPPxjNooFwDkutYw5W93Esl4exaWg/pxqZj69qOyi9NdZqpisIq8tp
xgLR8vG0WXRFKMIvbw05W3A+ArJxWQELEqa8rRpDQJk3O+URO2d4QwqocV55JomOcu4sR/Vd/Ypw
qcBx3o0PEx2qIpoX8PUT2mLkQgx+b7RInXqRdWg4vyMLQuwI6atkokeJiJfRANOnfAmtGaCNm9tt
AWUcKDmTkifkGp0XoARLXTGsZxgalIfFaHKt+NPM3SLIzPotAjb0JZaurr21hyXbdcaFVkh3mKZH
1nB7gh+q7HHBlSWqRsUjgOSRSvXT31gi29d7SH13EzoNmb7Qw+SKmrJ8ipzfWApH3zwi4jYw/fMU
8ZTbeZhxDjXWhsAPirHWM4IU4+n1Nl6iG9lSPhEfTBczSK1fdVQbUUGzqAQytYN81t4bRIj2A3pP
owGFV/vgMCU4vPsNTNnHiFstxPgbg4sesM9ufDEOIykMjjX7Sd737JKul2rGiErHaNy1AU5GSRQb
nKVxC1LL6T1w5Kp5JhP/qs/nkdwOJxV0i5Yb8MSPVWkY/c4i3FSU+R7J6ts/SVy+X6pT+gehQPIi
k7VJc8JTnfxRHpbXYKOQqvAJOB4qqGSmKnTQ6dadL6LoiS3SnXInXdNNRXXYyfGP0Oix/rkGOzHr
dxXg6wD5k16IHfBVgOPaJhua45Icl6Z7Bh+imVyn0O+V+cdtk+trAmI6OQEUUhXWvrEA0nylOfyV
k3o8Fg87XkBMNkDZJJ/mSRfcGZDsyUscHWlMmEJCiY5QQ9Jm252ymRdFuHaYLKuTXg2bXe2ufmvJ
jvT7qehECQ7NOAB8j5IDI9m2uHErYD9Vlqgc7RmmATqz9znmUhu5/5vRRDIJYeGUVtIhgYoX9KmU
V6+7JNPlm2U3uEvQyvTF78Xy93VPCmE2i0dEZfhLnFjkMD+psTiZXZMjPBGD/G97f4Ytd/FtD7mg
PxuaLc5ef7zXipeAqlDqbVzQUOhYykdM9rqX5Jy4TETINU/Lxs6tpChm/kZu64kTJR2vaYW1Vz9Z
9/WbfrrpaaVKD/KoSzBBIGQXudA5YTV5Qqf7vf4XJV3CHFrddjM1fpoiy5DcxQY7nF72+JMPTD+m
2vE8iTu4eBz8j42ll1VlWydoLCbJmV+V9BaVvh4p8Ssot6c3Mnmr5czMPHfKk3xWwi2aOccmflq2
ouD1mnXdilOOZ9EijoeB9lWBUontanI6ZWpi447F9X9hH/1EhowRqkBAv+PLyN+9FPoWF17ziJKd
YOWdV53/SAyqJCIw1hY44jks1wVmObhEQvsL/BFQoGj9zQAfP7xNWT/LqMfNDAuZHI9YpSAT3KBT
mLk7jopSX5I83/n/foKvx1A+i2sYZsEyIluJri9s3SZoEt8//xTroZWpPYQXhv6jX5gJWOrQq0f4
KYJZ7kkXoCW9VY7Pe/pC2oRw/Xs5+fKr6mFg1XELuqHrwH0HPVctCGIwvPLQ5ux3xilHlQ/srDo/
FIl/DhSrbNxpoiZg4yHpsImxv8ve3hkV3iclwYfKNhTQDRN/vBg0raWueCn/sF1HYKCvFaZg6Sav
QGLJSU0N5srBzTBoWlXtkr9ogKNMPDFb9QbbHTyiPG4JNawwivJIYUHPDfZ/aBD9eLFlryQoQnB3
qTQ8jSFulQalL3vxf0GABvwd+uT8yC4BSZ7jMDgFP/ExSftEOfvxxkPFsmhqfJhV38uQt/l+fYmQ
cwpoUn6CzNeQVDD1hnhnpQkVamIS62Pc8t/Vg5NHiVVySbbGSUZk7r5RVVu1v2o8+/exbzxg1QaL
7Ytzb9IYkzOkhWWi54K8C83qalQUek9Ch7YzY9LvoCDmME8syB09eXDRuuo6o8Iv87q8Vumk6Ukz
U86QNW4kYQI4XKP3+99kMLuxfxflUhhwExpaJh2D4MQPrFwvXqORgsyENKOzN/vNXQ/YANXcQ0ug
5VkRBTKrczYBy5X7Bbx5k/C2uESsbT8AQnteZY1h2R9caNIa2jTx9CsvK8GPXeb9pu/AjtV5souV
T3f8FIEQRklyQYQ4EEXuVU+xYKG5sNy78OoNILanGEoypfE4DRDZImjYoIksHg7bu6l7b1StITGp
adluHi3otT9Z1VaYzRBU3+0EGrNZkXvWc6MSKB5xbwSDWAuL0mcnKA4PqAFtV1862/QarA3TnVmV
H6a5gkO17e58ANr7antHmHINI7D2RoDoeprGpwd2KcgrrYQibkqW2vyyZaOQs2bNoMZhbOrLXDL6
3ohawtnN/l/Y1UrKXrxSLVnOTSTH2FTA9SfWV5JLZLrPpuI6/v4QJBqbzgaHcxNj2OpHqP2XISrS
FolXSRK6ye0CZhv4fgIyGFXUhtGei//4UrQJycQdhj3NWReiM6cqSVOwGzGv59/WcuLajKfpxLbY
02BhvT0Uuogu+RZyPgAGHZQXx8pjBuJMrzUhzwl3jU2d1WIR5FS2DxyzpAwps31Glz+ZP05xeCzK
rajZmsGCHtGoaoPNf4euJE/UrbUOGBF1IBlkXVPr5pFiR+5sygYZTrPV8k4z+Yzb1EOZW3xhTqST
2WNDS8dSHhkrItdQJAPCpgj2tLHyurZkfJGfrdJOA9QV3TKX4XVSWFK2g0viTsubbIc15KhGW9GU
PnjqQvpEkcUibDom8LqGT/4tYKTomxS05K19rv3BUOCw8aQVwxWXYbWTEGdYY4wXdcnnMsTdlk2a
vPHnCDzp23lLCudL2PaQf5N3y61ezLFaqVjBAShO9JaZyHnsLo4F/tXCHc0zDtE8b1eK25u0NVxo
oe8obct11nKM+3hWUdRRQuvqDQ6Xtu5l9+2bF7QCuuZhgKVNuEg+QVM4ABAY6WArWfRSlN0DzR4/
rg8+avLZKpBQkajf3M0g+UZLxNRm9vfBubGOsqhDPR+fIPvokGVLU3ugI3M12nXMDyVEpnOLPKsI
qn6sxv8RpeG37TATdTbYqyQs1IGlM8S6TGz/rIweskryITndTkDYeWzeHrAGzBZVnjQ5n6v7PqEp
3sfWmtA9SOpNzvL37+fHSOGglrGE30Vrxce510zIbyIa/1L6LOkYi8AvH8mPJZyKJq4YIrQ4TK1O
B2mAzQBMNxT4IFAloTF5FmcnTOXUSyQeltk1qmFxDQ5D/Zodw1zR+sdgB1ZOV2T4vwITXLHyQUjt
27pufNudTqvbZS3KXEO3Wx2vpsSDemIAd1S0jvODafOLWYJIxc6X+EfoYo68wwmBz3vE5ef5Uw+5
Gw9a5BgoQvIINycvwkvHxTqZJmMVxggsAlgra4yJ8Q4f/t2+dUCn/r0WwpveO/SOuJKQmieFJC+/
ONc24sfQsxFqjqvuLaikXrlsAbRRFAWG/s1KMicXYG+jAl3Ht7KEv53OjwGrOCyT928TJAz0Klb4
imQIRSBI3mUexCFLqo0N5wVRytdWdY43TVgXZ2dSIbpgP6dc+PHdQ/OeS+fhFspzzepoy/LGFgtI
8J8ow2i0gFciz8byqDZN34reWVDQrpt0OvaeVmPgdTMzSog72uNtiaYLHrEE01eQw5JTmMltAuz8
k6GP35SnyN7U6z4FRtc5GZKcp/xRZ47Qiw+6W8PY7yTSk4c5fzkyZjMgP4RK4+GLtQr24pAT7zxZ
FSIzSNRRrqT9QCkyRhta5a6/3zJuQo3GAPKJ+18FB/JsFXeAHZvoi/ASRAU9vhh7S9IZaiD9HTCn
b+13BUawcup0iq3sRcjsQh/uNsroBVgZ9q5Tb1C/Q6M+YeC276HEr1th+EdWasCMEjqhmIob0zhw
pAqLlWPNz1dIUusRkRoCIPdnqFBgDyT72i8Mu1OR49PqEcOjnj2SnWAb17cELQVU8vLnIlvdeQo6
09ii5NLpzMkAAu8mHCGV81qs9a5jnlML17+RqqQRivWphr4uuL1ndMmsJ02QnS5BySidKf698yoN
2gCJ92mS/jBEGFL2Xv/m+WMxhUQMoq6ze/SZah/pah0drj7pb55P7B+nqSKT00/Alyg908ZkVFiL
hHbYmIqB1a/CVfCL8JXTuMyecnhk5DYLOxITiFgmzgR7fnrkhfwFrbS1m35sswVl+fdv9C7kRbZI
SK3WDdX+Z4CzvImBQLIGAcGsD/wiURXSWM9wKPvCKYp/XT7YFLGLq7HLWQE6jUU0rLzfqTz0Guie
dkrLpWALgA81866TG3SBXOmnblO1HSLFic+Db80oDYsX3Be71byreJQU/KHRHJgt/IZ5lw5/LFcV
qFhv8z1+2SS65lc0XHQ3VYXZ5zQA8O9dIMs9mwrfo2dhmCbISUaOorCzz+RzN/zDnQPwMkTI3uh7
r63MgA0hdHDXsan21EMrCs+Dj3J4TW5kkP92bpyh2lUwckjPJV3W0Y38mh4Saei85oapGw9z7VWS
AuIPOZLygynfGfTC5sW1v+lFSYRWyMCVsZvo2itEqWvSiaOMhoTYo7x0qc5svzV+UuRp9o41MS7u
4ANoRkGQpc1kS0gzD1mPq3Mxh34kAatVrxNf9dplxeAyhyk/CxlfhNnVCQRVCnYfUSGO6GRMqu+z
kzNCG6Xf8Ipz9Hjv+qkTe7QpwbZqimMSgSRiC//nkAEGnpgL+U1/hYskDCOUC1/rRR5gmQQD8ZXm
paWAI4EsdJu5Qn0ntWkrqjYirPz7z5kdP2m1WS3Bf1AEcoGQH6ok6PYuRqvRYhANzTdQRlnATyQL
CiAxz7pj2JM2m3DpE4uREeIApcCYSKM4o//HFrH1SfsP9fMoDKHmsL0eOvFCNDumYsgBu2wQvqFR
Ev5TLtMjoTj8pG2SDh8yrygGoNVMYBGsdiAzyUbvFyuFb8i6yj6rCVf9VJJ2PSsgOKu1TP1yCH7V
9oi34XZBerKwmnQvetRVLCkxhPG6rEHhzKx55pQMqhAKty+mo4s+sNnmt2pQahHOyil8YY7c9Prb
hl+GD0jsdynsqq/njZbXbqUxmw9W4jcSPnjm5HIFea8/YV/OodruoQNdo6Qac5CSUnBiltkHdvbv
LWZ0Ch3Ti0zgJ7/aNsQBNmFgijF4braJmd313lgMptslZiUEhkEdX74pbfq7tefjIqVSSnC7QBqX
L71MvWvKX26YTcFrpci7bZRG36SepDjAcDz0UDGPEWynSU+m+1Wk0fB46kw9HK+hShGCi8YUqUPP
L3gjXSC0e2EgxI+Qp6slhOEguVHehtW4mqp+eZ+3oK8tsa8uN6ZSXq5/9xfxMKkZ+9uPWTVbzRqD
2czYtkukC9Y5CK1XF5KiTSmNHXNEKN//Sb9KWvi6+KIshSh5fkp9yyq6suWzgMXdUJp83Jpc07SQ
zl9wdW6/DWeL0pPqE/Apt3QMTpV8IwGbw+hZAOKHQR5wFfR7G6yTrkoBjSSJ92BivnF6+7B7LI5u
AvcqmJuxOF7qZs+yTjvRnaK6A7gotb7KeexnJ1ADCyL11X7ObT6jT8ksBXo8azKF0O++fRgzRgmn
8b1ZiPuNMZSWHXuhATR527tRXTvrwTU8N+5V4K0XH3ZGEUha+y8h0fiQxfqbYrXW6SX2ahIAPpvO
3VE8v+XB8aoGZsC97IwEGo9fDXbJt3ZcGx0JXxQdKOeK3zmk/phBj9KMf71WcS1feq9/8LUyh7Fu
FoBuaHxzPO4NSpFIzPqwAUNbyxkiujcHwRzHzPpyQiutsRDhLgEPdU3SLTykUfl2GFmJS4qplkIl
aoWDHIuStOPwGZS+EOEkL6lVLOxPiXkV5CuJESLVAaQjk7OuT50TO2Q+++yhmgZAJka8DIb9MVyV
priCEq2ftTZ8VIiisLGXp92/Dg5HG+v1KgOSaRtGx6anbjt6YpTv9uPR8D/ZYjv/z8DdM3VrYLb0
NwPcovRRqdDmENQjrA7iP9x9dbtWIpqg/mshsZ1fmZn1x0m/6PaKSYHccKbwkTAieIXIx2ZM9jCD
YJtEH8IM5bnhSZ84vLiOX6HAgHXl3rMasZoSWYtwiMxEHZZhHHTakHyTIYUJWKhsnkm0PF1O4q3e
BHfOqQlH4q6LEHj4hc7bW+KBI+kBQlebjWknZR8A6JvMduGFs+fyjo/0gT3fD8St/RHZ0aycQ1DO
8UQ3IJY/hMGGmnutJS/W5fC5FodjaJp55CDa1g2dFbsNVCwrUIhuVZE3qBk243ZbcVR8qwe/jyVV
zFkScPYKNT3zvhmAAzhc7tHo0e3I0qUE3++pOPnalDwRmUwZGOdMA2yXKF3vA9GlbD0qFxZb23q6
6vGfC6AUzFftkRKp48aH1WlfngBWJ7aZqFcxhUzdrf6xVUVv1jetW9iYr3Pv/ai4n9vRMqMamYyN
SttSs8LQCoM05KGMtmubcczLHAUhfshc4xuC/tvo42DjZWdPiUrSyZxxWaVxbkTOwTQlBBtg+kk2
UNvBG+sOtzTMQ+KTNrZTEPyZkSJ6/qrlEZDY/HaWKunRtuMa/4+S8cF2EwnP9iZu9Y6NA2BOgGIv
uyOuC3QSsKstNiSsGeM5rDhPuI946XqaNXf0CTQh5VIV+JKwmZzKY5otV4VGTs4dH7cJ9xpWlyWg
LRicJWudQ5nUlZr1e6Po/McC8Gvs8WsvQ82iaCnOYRgtcJ7Fa0lL5pC6ZW+L/H9ddxVhNpRT9xst
YoP8GMa3FPBjg5fxIhplvgODYFLPOawjUBovMmDOxMBsWxNf6A6SYMFBLqCqpw3bFe5z5JlZ2nqO
8RDJAzzyqvhRjqYa3TVscOCIW6kGGOVt3sfUiY8esKWDmOt70APddZGEiAit8HoMEkey7yzya7OU
pG9RS7a/SSYqCFESb6uJVC1uF/9hKG8uxE8nXz/Z551/hd8nb6NsMNxKV92OFnWD+MHwmG2ODy2d
0qrwLkjfb/7J96FuCHEgKRKu8mS+9J8tSsJviK3e4M7uXHUnpOhOSVnbSjh0/IN9p5BeyHoLuFgz
6U9P2tMgeby1aNY5/5bu7SuYoBuskhOUk4C2GJJQy7wBpKRNFcrGaahM40DKqOjd1jrNwRaKrfeR
ttmTrhRMbUnFbCM45Wy9Tk9s+xwZ2anGfFFOapCUGtiw1cHHTjxVLtvmcsY3Zb0250KCE/2CCGXg
57lwYsFXLMh/ShVXT/trHoFuJRC3coFrzyN7M4/WmaoYnX1jF4f1T+9pVXTrnbCRiU8kxLjc3hX6
1rMUvERHHC9LJQcFbueiwLi9PVUUczR8Pn7C7sXVkco6g2sYHUu4EN+voNmvLRfrhYKqIQxzHSQF
ruSGNGgj65kyQvHfaDICWGCwfmRadzlRceOmSH0qOja2GuTQQb7Dix7vyAmUUUKap7GWmUSXHeIx
AzzCYKfanZftBouX0xphoN2qUbWfKwbATv//zawJpoZHaehzl5b5pDfarZM4jvaQr+M2xodkD+ai
Xnsnlt6e3Ee3ir899Ynj8ZzO9NXjpKm1XnnSMxE1clohdyAR7B3ylnfPqem2eJ/I2GzhfR3ZI/6e
o+dkMkfR/tnXeLyYi8/9IwMni+LEv97sLJ8YkohPJUVJLKIAQBSP2qN3mXrH/p/9p0Ut7eFUwjxc
zgchnU218RDK8Iu3E+VMpMUq7VX5dESqe9HzAaRPDyLPMPC7Dvi/MLBuDBnwqWekFGvis5cFi+9Y
WbEipiI1mbI0ab3O7PPid87xw3cwnNxUycfLERtUKV8armX2MyO/9ZeDM4uJyOBjG1grbxHldOc1
VK6L0V0RikN6IwdWNwxFSfOg3/Nebfxpdy+x61a5cZH4Wz25XTlzqPyJgahHIGmUE2HhFYYSsE5A
GZx+UXVSLkwoJw/XPBk7oJGD3iICO81kp7N6j7spu23MiEx5ovwRry9uksIpaO1xYvVr4Dqp7w+A
l/DgbMM9tXlwS2AYxU0PbagfGmsW4fZrkQQtObzlvORfPnWBlyz1pM8OLoUg3y5m/DDYCG7JkBsT
EB+jAgWs3M1wxgoVowQ2CJ0FopnPH11i1aOGrMfS2qOHOBekcT2rTyIDlaHLWUPW/lpk/xhFQYn8
CYUpM7N1s9GbzML+0vVuZdW2MiJAIduIO54YG5Q7S0d8v3dNYkUIfF6LcTOUfnXSirCBjgU4g1G6
3J0cU44YbKpai9RRx/P9MVrncSgYjpGOpC2Dd7qunodkC9nR5hXvUxIUYdOKx9xYJsIhuSGudPpH
FEWLsJjyLP3kwc04VeO0rlCE5T/bpIhQjk6A4qbgs6l1M0AlXdrw9yrWyrzVWVhorHmEGjTJ605O
cv4fjSPZI9dSclml0f9t0ufyiZv9KePZAJ7EmIwMrSrwEXASMgQwDnqTNVVeGnM1k7fRzNI2+T+D
tdv4Q/ozDjIlDj0JdSEBNcFj09CGKpOcLxh2SW2V5S7d8dm7ctSonUdsFG+PmyIYkqPJT/Wl0+Hf
5hBj58FNEE2y798v2bbiwtVyW6rm3aiwWS8RJu5+8SKkFL5QA2l3wW6g/P+WVTgrWTNjtkBPS0Cu
DBmbaOvdnZy7GWgiCECMLnzdSVYs9Iq0qr8QGQPdafsYxw9oXZgdMVoIZ2yUNMyd999kVDo9GBzg
ndMeLRU11HXBIA6XbP0Mb9AR6WRuMHooegRLpfHTeJA7pjNcpZaw1ycKU2seoT6N3gEg34m6yC5c
cB7RVxyWQ0vTT7l8Sg3Ug/3p2tuC0f73N3QPPSn/Jcurh116uRc5KUG6hDC7h1vu7HL2jv/sZlkQ
SMoM+Nt1BRqsq6l3ooLPGYEGogIn1+o79jBUyhdK9GqBnmnezzKHO1L2qVubJ92brjuCJPaO+1CF
mGCgKU5rKd5ZBzIln/80VIhplM4NL0r8POfAqNX7LhHawX/vxoutnfJbhwdQYWNHeTPNAebCaKjg
TwnpUuFwx2i9S3lS6exoi+Z8NoLGRuQH2BzyVgLpvBWeyEHAXgtJYb2LGj76Z7yMssFiyrxCpYzJ
0yFm4w5YhFok50txDFUhbyr+MTY3opkQXIC5Oxepgqu6AmiabAVUUk4QLH4MyMIxAHpmDgBf12Mc
tQl6SHA4OLxpycyMZ4gGBMvXBaR3xxDg2rdndKzBk8RX/4EPqHU7An8kniTI2mCXC8lvqhhGevNm
kWA4ROn9cUhC78KwVwJszaat9kJYvLCf/prUVKuV6R+140fDNlqffoF0PQhNh/lMNSxVjsxSV105
Aug9sUHF4pXYUiqljFqHLyukqiMQzVy8ibUrPa3CnwNNZQl075emzDyNEd6c5GgJj/KcKHmTGA3/
3PzdB3Ehpy/hIDf5+H9ppRHMjL4HfdqgziXwn7uU0o1vPtuwOeJ5SM/VIU9PsItYXwSofUYnESy5
gmfjB+3VTeuIkeWuqz+Fy1ImYFxS0m7oR1q2eEWwoxapLpiXAgwri5ybuj2hGcz7gM95/umE3PEw
AzHaZ4/TzcQRZkxdb8no16d/suoCFz2N0k4H+J6UnE/lOqSsdafrFBsS4SOCCIy3U2ACnBqSlnF6
jHmcP8YCe13q/BVxCK3JDAydpHvQ0mJLQJ0I2qrKQCBsdcUm+e07w0fClqDVyHgBH41GuEqFSpg7
RQaYsY8bW3rq7BVJatQATEIQ/HPNBOqEpnoePV4mByb3gK5/Zhfvxmz463twnDb9Ev9WynbdcjCy
9gOkTwdp2qBsYMiKHSSprNJCYax22K+QKbOvsscErrYNzIhxNUwqZneEXIVDZZAwUd5y24Mja3ir
vwL0725F6aLgbi+IrhSu9/Q7chfRZjcCGuRNvqoxhf7AIAKTOQHxhsiGa0P4hTbERrmEiBzvQWBT
/hbnUBsza5tDot2+KiOhloCSaxGMB7DXFgD9eAv9wqgj/cowc1hLt7a9YczXLtOT4pQp74fjaqq0
zNJljcBemJ+8Mmfvi+gpE3sJ9qoIdEOXbP26saNn5X8olfkM53B7hUkfWOI3kWUmBkthF6FWnCj5
d1BmTmmwYwHIPTMNsCIcUuM0xcKVedJlZ7G3kPRr1Xs/nuo9zlzfpd1wf305lryTtbnRCOVPN2Hn
yyc/aPpgVaF/MdbVEPf+7vh6/mPSiivJEcLM+XZ15n45lX36mxd3lxORmKF8m4o1hSuzp6EYsg4T
pNottiGvL+9PLM84F7lPWfPGI2ocT0gUglyAebhKltQStY6vhr8j+qmTwwEMbMw4P8KjlcQZnCsX
OFuW0rqphFG3boyDXhw7B+uFzI/3WmudaMBkKuGBhqjoSRoYpS/FJ4S95Ln0qVH3ky/Eun0jOda1
A+1VJkcCHaqtfpszBXqXcUYj7toEpH4HWegHCxhUTiC5HVwHbxxidHpkCut8nqPI5q6jLJBOnabe
VVwB3lTDFSOb5+AJ3U8LqIHLQYmoIu8rO8B4dFA9LfZ+uLOkAVBKsiR8QWoCYSzN2ZekawjOul1f
fBs7PxROSaf36C5H4QH8eIWT2GyZsIYu52yF69vqd9ZzesXlWHHvaWuKXRIPhN7Joy8bpVGkQmls
yNm9FvQpOJeEBmrMVWvKNlo6EkQQ9nlseXAk5OOmw+xBAV0qH415uaLKwdL2E3Gchyx0Jr814KAW
CDFtOXXkzWeVFLZE+jMKSCsVRoKFx7V+4FtZ7XZu3HzKsEs+x2WPSfT4GF9S74JfQqZXT8203cSG
PcjmU1nG8AWiJeAw+D3h9dr/1V/e7qfdnTuC7Xqzyk9fdIXZ07uI4hIp6wDPmwjf4oxA7u6umUb/
EMHMhV5X8uhurIDnp6s9AdGh3qCu2LYdBbP4KA3/HsopvHeSUHsJS7Ah1b0zSyj0SbnbQYGeG9wj
2BkRUEMbHJnauOJIve0YPOX35uDEwsZ4351rhdHagRqYntx7Yuy2mastgZUi9iAiYaIcXOkUZg8O
3VSdb0bJ2jNQhs1f5bV9+VMFGJ6UitMjpKiR8c0bo1wK9ZbSDCgaqApx2QIpRr3gpmewZrU8g1q+
AGPqC7YjJeuSd02AiLnUNxGR+MY8ixQxC5LSHTOuA4lMJTYQSlnHYPG1okIVh1br0TyPMLTPsXo/
PAJgBx39CjZ7Cgkk9BZVhWj95RMTUHz/IlNhJrPWQIyK9vtFwTIX+ZQTNw9XZfGBu+vffsMURhzB
/FpIQVLz2I+5iyhYXI0sR3NHBfe1djLj80tQ29DVdeHb89Q7U9uWKZ562XJVYIE3Gh+cYXTDkjEZ
/s/uF1diaTJdRpZb6fzO1x8JGoB7yAm58GmAJM0Mj1cc8mzycZvy9aBV5PtqEwJT9l3YRUtf7oxE
7nSCHu2RKhgB6jnAxzCJrhh09okvFMyA8moL4SYIA/a1NO7bsG/oAJctAJgB2hKVvS3yPI6lrrqq
X/gSbuDInF+aklugoNyaUbH9eIiFpavAVHNOC834XIhzqse+L8RsKneVw57GEtxcbsRrZxbbqyQI
Xw9SA3NV/7BpWTtZhimJdoteDI0gRB7BqugnSIMltZks2a6I5T3ZOBCxpTYxnEYv8q95b/bwV3hP
MI0uSGnV96M3E0hE06jtCG/XDkcyOT6gF0LFjuinc4rtMsWjaYw5/tqjOdKDbcrgzpAPgk7eKwel
cCI2yZViJOewITrXomWmkFEjhM5MyoL603dq1uywR6yihDd9Bb62M+00U2yZS/6HZFUy0UanVe+z
c48GV/ssReIMrrNsVmtlACCBs6t4QfVyCaElBnhLhgbjfBIEixewawVd9q3eUt2MW8QsZmrzsWTt
PMexl5hW7MQJwdz0mb1NcAKN7z3aYcSDLtACHneo8/uypT4Z1fp0F8SWHSBDlbENfqcvk6f+qbD1
Y1ZLrzi8xOSqNQz/6w/ppBMpVbVqD7SXAdI5RSAOHHDItJx5igi9Wkr3HXlR8juy0Grknhh0SxvX
JGzrc7nld+IN/kmHO3BSMaGKXtFgzoAMfC7uVb8KESzPTT8ULh8mpPRbxA/Txkx/uqwOjf27EssT
8m0we3cU8GgwFcjWhtF+qMlcRfrJFhxemhCGwXv2wxLAKNPt4QP+oyvtYDT8OYtRqsQi907FIYhg
EwtYFpnT7DMVHTIxiQcMKZYhc3P4oyMaF20kD2k0BjsqYPrc7Pb56jI72Aes4uJKDepbilFxRmrQ
0OgdwnJXckFp+twmTJ+E0cb7NjZW9gVJY+T3CpqOZ4P3Jk0rgD2cHq55asKBA7yJVOyJRQelcazH
5+241KC7LlLuxfUPY0eqo4MuqRo1a6RLgtx8TomEnMke0J9BGG38QfDBizxgBHyz4d95EQVDXbKb
ROTP+8YJz3Orira6ADC+nEVDvupBr/cE9ACftMKp1Wymc3S3L9e7vW+DEyY2PqOjM2fi4rV/EK8M
Dy095Ij14NGqM+K9a9txUvZFvOWdWO22HAHFPQe23HJcfcgpmcm+Y04OjLt5YG/BGaOfwAQPY9cT
NoWRziA7XQhaBBbwBubclt7wKkFcTQaLaO+yLKEZS546VtSv3bQmVYA5KX09wU/pGZ625QGv0ruo
xBoxCaky52gAXQqTMObvImvY/K1F8MNVH8xpljFqeieNca+zLp9OESGYqqKQ53zUi3Rb4jxTvYom
wYly+xOHxngnNXv7yB++bv9vTnhAtukFPmQhB/kqq0/WncgOv6OuE03VdMik+jFM+3IGYgRKL2IL
BQKJFgKF0Atb2ABVLiHjAqf4juKuaPE2KbPp06pj0gsqHGBYnKZ2IVKaeiZVymUoNVkVOm8kvXde
U/z2gECL4xwhGPKWQaKdins5v8uXD5Fj7/2atOmQCOYO6n0u7q6tleoVxhKYfLSEqQoH+ErmVNWG
apehnx3A9e4fVKfb1eCBClOhBiypD9LHUv1QOymTZqfe9RHPv48ZF2Dw+tmwt/NTSl2H7Npso/c4
BL6nEV5ij2CCvvDVxFYsACy28t49YHRcSWzzsJ9fcyXwh0LjMtm3hbSxZ1o0XuSzQuwO/+VXWZPK
3JRl/ctfxjO8htp3D0RESvmX2HAHX9BsnMyvZwn624LfTcSYhx585EKybQkC32GN/pS+btodb7h2
TGi2MatfmDWJO1raFXtv7INPFRvw++VUZWL3pRZxiaMFdFRwikm/TAtPaVEaBZXAcxVWeSf6DrPo
afT0Pk3iVxwsbKJUflCQwYiFtGhksvpx6Zk4g1SPAkoTcjlPZ6UFCVPM2i3Dzxbwd/dfV12tR2Xp
CyPd1H0IMMNYpfQOLSo04PAD+/D8N2/A+pncskDFhcPqDnc5Qfo2kkX4PXH499/9S1f4YTZSn3fa
+il2tMTkleSq4VewHpVw6E8bHYSxaddOHekp9tE2N/8fZoXx48EdHJ0N8B3dMmsEN6nMISRw+twX
aZjC7aQQmLQKld9VGpXrpMNTCdwJoIC5MQYO3nMcWJPURZrI352NAvjm38F+VG+dbNc2TUZTYFJq
wvZvVvuftJ3k+EFJAwYFgfl8DOqStY629mIO6L7G+q8fBPM9mQKmbFr2ec1v0T+2ESXh5JRXx9X/
LPxgnduKLMgonhPlUtb/lKIWlhjt0nCtlJ4J/WG9gFbDS3DwyOVkiGGvlZu+rkGRl0iQTn9m5bhx
xPLT7KUW+n7IDZKcCNjjsPSisSJCtXgFF3ZVmnfhGvAYM6PhpGoejTWcPCCMPqAsotZRykCfsOBm
K5Zg4ht+zkzXZi0tUhVLEcO5DvByAPq+CpKO/9oSE6KUMmv7d6sr+5kKxbo6/tTEJoefRDzp7f7S
ltYHku3acIIYRV9zBHIGFRmf0J32k3f0ngm3HJD5OCg9Ah91X4bxpqCfXQbN//EQqcqIpSlx00uw
sVEwOzFS+hyh5NCtk8mKLsCRC9hPtumFamvTpnexfcVSObzdpw6eaHudeTQvdnUprS4cv2Q83oOS
qY3pY00iOuIfzsqDiSQMOhZkQk2NENpvkq/j6sxMwG2so02gZdd04BBJcRjrf8xQJ9xeXWOa3G9Z
Zj08iGpI20grQWhSBmemPAFCIRvMP9lq6Afu/1p+iuBy0A4T9yBqHFS9tHwEPYzXdcoZElAPVALh
uBMfS4Jbx70FlvXAfSXbc8uHWSoUn6eXBtYopOXvG/mNAXN4vzAVzL8XpjgOVe7XaSSdwOgo8cb0
H1a0BeQmtww3siuMoljx4fwyFwYPyvUUvOOW/KjjZEx0ZMXK2mCcZkXId9N/2LpMBrXeHEAbSQaD
GPZMFOOzWYu4F3ifnsMT09pId40fRanLfo3/mRmN+1f8EaasUUmjVDUTDa+3pfaD0Y1zvfG/+JHH
1tcCpsTxPvLVL5TxwLSvutuczB8hjXDR6x12w6WMcldKsHsVjWZWbSZkRLrWB1v/aAixGU1mmUOv
vR0eLW27bOhmfa1vexIdL9Va80O2gbJW1EuNjxQDIwcrOzqzokYD+GAF3mFze1/mIQelun4wMuow
1tgV+5otK49RbbQRzL54JQM6hUKpjJEUb7yMadnvMEBnAa4AV+pg0iUTexZ9q5pUU55FApX9EfrX
q1qNIx29SexqAMgjPH1sCHGd+2sDxBTnyc47j+99dq3Q2SHP07dI1DMQqgm7dhsotcWbLDi30GVb
CIbZNlwHgvZRfNxI/hwQY76Bv0WKNaf4RzT3+beA9E9vqPctf+hOcjhMyJX6cbx9pQtiN4ZEVeoJ
MbHo4Mio2MQyIMmtMOWyJTozRmcCDAmN4ARJhVmmPNb+54KIoJfdXMUY2FoaUidinl0UfF1iPu4W
OvLaYlWlekpHmcrY1NWn6ablvg7JlTtNOm04H0Ag2ef2flrOEMO0D0zvaaD4cuZbnodp+lOfQ3sw
KbQM37btdbge3NH1UoyfJe1pzGjULUkvHBUAcI0iYKIVbcr2VDe9jt5CyPXb0bCguwUFgT+QfJXy
eBVpPo7oxiOTz5PjQoIO1yOHijqiLq5hzto/KHTHyINh3RFSNcZVlZpoHHmx/CJasDV7bRkwZUx+
Lpla2Zm022w2XJ2VpLa24dX0nUFjHCxxJY/oQD5g959TNp9clAN2bltI7jJBMgT8wrOHcXz3t2tz
3v+W0FtNWdGlSk5D4w02ocKGln/OUNJqSfP7R8cpZQHG2jfzqtYv+ntehhNsMa89usV7N9Zb40FD
UIbmmeJ2R/eQxZiAm3HgcLJvl0SWhkyA1NgWEXriOkU81zOC1XB9MjJYLGZKdVs4PQEYjLVyNf4Y
QZtJbl3BxziKNiqAlNu09MtKipFY7p41NCs27Qr/6naqSPI1Upj6CX26W1bfyLYzgbNdcc5X1VGV
1FL9PDit3RCkRGsghXtubU1n/OGJDwe6qG1ayTVQO/NNFc8kNjJG1e38bLLkTkCly9yMQnQsDd5H
zMMKnrC+wpAznSD5DDN93WqsmdPN4LyOFgQuTClNSIIFMwpxSo2AVvSYKB2YI0RhUKrRek/PQUJf
+1n+T8di4Ex0/jnpF6gApNtCvvmven7ePbrwzJSITO+YCKnmf6U8IgMV1KvTQLCX9eb5NDpAqFT7
7ZmX4fkq8VYoaJMlkdWFfQIt+jKhLBKQ/1sjkkbL33GpEYmoHsMZnQmK/ePzLmm5H8YBfITpqLCk
LElyUIzd1uE1v4A6g4pPt8M7sMBxs3wCsF73Bb9s6+lnT16qb0a5nO3pyTNuQUDcV7iZeyNVH2JI
MFk88OtMmRSvvuGdSjUM21lYSrKH5o4LGESPI+UiRJ0KWXUnNpfuDkDXMMrGCnRHsqH3kEVh9LWV
xTmh88PNNhe0aZ9fqjolBdcw1tyK+Kb3ELoVOOOqWPLSzqj0dS1v3CWVazJiq5QX9m0E6cBVGjgQ
CnKh2SEtxFlD6wjt9vFjdWRtOB2sNcM6HRZ0PeRlmr5WYykU4F0Gr63dOPoHBV1HAYmiJae6A72N
Vy1tlSnKfvUhXUAAOwQC9g0zigw7ZQSLsetZrsEQuNQb/8fLvNpCXQJdh4i+HpKDVamSf6XdXYqO
KuOfncUgmEXwMd2u3Q8vor4BHDe49j4ueUa/kwH0nSTa7oviEXyH9Y31XxBKSvso+6oYYnBzWi63
xrP0vkSavFZjA7n20boa6PamXkV7vndw17CMzI90dMZ1P4mWrBKEYJt1MnaCLtyut/QR0Gr+2V+a
U+3tMJ6GS8DIujmJ2drGBhGDkE8TAYzl4w0AcjfE7HJa4SdJEP/1JhBxnN4P+tdj+x465S5dnZMg
FiXXLfYWyuDr+NffQBukP0r0O7vUCuJgpQSGPe4vrFtV+1pnPrlG526emOjGSpvkpUeh8dSbHsHk
NCTLkg9nqusHp4sHcBurxOsNs4N+41BRA7ehAiZ5RBDVFu9MEhdlE7elXBYQWr7gxWC3OGuFLwJP
7mTzqPwAeWFVjmRPPb2LDiMwbRYCfG6BcpgBnLSbHuT8trDZCsvaOTY47qRzG78o2pKX4n57xMBy
OrRzcMBg3qOnJXm0uRnTJjAec3YkwODw2kWzokZsR3IhB6wQ+dkIsxWrpNN6p8ryMti1FDy+tCNJ
WERhQ6ibFbVnfIvlVqyIZ5Ij5x6RvjlZoWhpy34AvNGB6xedDoawnfazfQY5YfygXqYJ6bMqo/u6
2TAkmOZzr7IFG45xMwKnQw6aipGsm2LAxuZG0nsE1S68hJLCdC4B6012asWTZvUX0XBqS5W0uoE9
YbzgAXJ11oEa9X6CcGqJSJ1D7xVKNbsWPhknWTFU8fOUb2hs+LCadfKOQ8VphKB5EnGWm96yWbK8
Th1hYqocu8gDgUjdsd3/LmihYrXRFvm5oDVOwvNKJ1bJzITIVPwHwxkohU0UkxFVGFxdrumTlUzy
mXb7N1mzalvmqv2Xu2t/WzEIRJM05iSkxDrF0Q0HEOpFr4VHIy4dy483UzZvC9CdReCRzrh2jhcG
KpleiKC+G7NHp5vLKRySc5I3g6Qs0mQchWpYTiCwezx03HzQ+rhkYlETAYTNoCSer7TCK1blh902
LHTPwAJrkJNRKH+FOJhVogYYhO/uocktGi67+ovIq5aP7+mbK9TGljJwRgznyjjdJmnL7Ddl9laY
304gv2QLnzRxqImZSxKDDldeDyoHtqYWNE09DP/VK5J2D1wUNOyrrWa/NA8ZKkCvdXFlUUBI1/tG
8RQpjJffcFBiU9QQv2fFboKqWAPm/KIZ31sVeGJsCUWJZwF3LU2k5iHMgnUda6G3pZrlYXGFPE/1
aE5a3AD2BTaK41TuDmXbJfrPFedW7FkbClDW494Llwem8K0DbSO2+CiPcasD9bCZNGOlZTOt67YS
GJl5ytlkK00Xhk4e52aKEmxf6WPxsAYxDk3pjxIHj04BXehjsHL2GAFbn8CP3Ef2HMpsOs4Fg4W8
dWaCP3D4ErBqtwmtO/hwgdYGMiiqsRd5vLXASN2uA7r5Q12DbuF0l0OpJiaHVGefIR3BYo/dmSdq
MDWyi8EmSjbIMHHgD9OouRUSxSL+2W5oRDD2vM0s2SBh8rorLJC+k9gOUB7y9rFzHZiXXH+/c0JM
YE4dBEwPs7OwIkvKgnoAHBPyAqgDfYXcEAFoaD9tHlp21/Emot3+IbsteRkffPScN28ZapRFvKem
3g4VIMLehNQxaiaavaZDCnEHYL+K2iKHVwGc26RlbNdErWISJ66bLigLALwCc76PxD6o6lE+zOIO
4ZwWPYaNR4NhFkFt1qee9e7N1duFhUZHhvEzEilqNYAOSJsG+SmDTPpM7TU7kKaQozONNsF4h9yM
3Q43EULRPwY5Eby5KhoUC3fDMtimens5NkLUvK6oY+lzvsDYiWP4UDwIAtthVOwaPpBV8YsvNvoi
zmt6X6IQsoKznf7UU5ZP9HR5YyR1XesOuHWW/ujxGHeruJTY2/lEuLUR40oyv6u+0u/fmJctOBUB
D6RQT0bGAaKIASOBxkoAejAbQX6OZujoLiYx97e7fXRWnvl1U+DZ5xrENazDxgHzC9xbGhjdLV10
tyCLe1jEWq6i7ZyqzrHILFLfH2ilDhTpoaGgRtvCoWucYTHB4o4D6oCmqfHT3m2ydEkZTE5xqC93
GHFvyehkn0DJ/M1sirQFFw4ZhEamRL+JgsTf0CA1q5PNkKyIKq8kNORef7SEk2L9hTUZwGdFNikN
tigNCHKupTqkrpOxUPSf7BGx+RTrRznnDZwKefAp4UkWS4rKjBm17aV0p5iQeoheVFVnLc8kBFNN
MCKQgzIY4z2qb6YHrLFGASWcznxNFFAFyTPGGiJM+G9eb+T6Pk15847aDhRTMIt9+zBW/JsNlLsv
8Sy+8/MXsRmGVd6VuQuI4PyrCIMsxjuhPQuou3Cxv/Qq8sgM/TghLiT4g3v0pcV+X1YkLyvf8kgh
LJnCYs4QtiipX60og9tCiQoMOC0uUW4y7bjhDh7looXFYdU8L98GDk/KNq+6+7gXHZENvRkwKTng
xekAQCSk+rjZplz1IZKnrAqVn4g5cXinKcB8ogOovYJWzrq+YMxyxPN+RvaAv1vuPRf7QZoa0DxU
AltpxBkPkOT2ii4sVU24C0KbNeftsvc603EnWdDt/oYdaTNtLZxCnqkoYnKSj6wB27dl6QjyUaJX
hnnJ1cMaEXC4RQ4qttFOQNOb1LWctbBrRCcVCqi9byK5ZnfeX1zmSEPqC9X1cRjw0imudM8kTpLj
xwZ2vCwg2yKomGnl1f9bBWCpdSgXdJIETtMWOV6FGhFcyCWyCNmTHXqPzU8lhVIM+nq4vpegZzvv
ot9ZL9psvg5m5vccjP3ze9OSdiRZsyrwALsDB2JAdSmML977ZUTOgiOIfrBCUA2RBJEafZ8HShM1
4GPk3FJI4TE9yKiKUnecI0S/YI4Hb82tdxp+OO6ZrOm5FdAPOj0Yd9X8YW337hY/Ld5TCpo8FsST
g3bINAWQxN6tuNv4s1+eAFdBt5sGZta2KUxuJFOdsPIWdsLXqU4n+TyFSvBG4OXXtFxEwVfDHIjg
DInpkH10xdhWmrkNeR5fiV6q0+xTUhE/SFpegc95E8bTeaHYNhISULxb5laZf19kWvOd2cDst1+C
YEjAL0ERL9fM8M+bKg0O40TI73G6XqEqx756ozjlFuYnIPdybEfDfVC1+keF/lumVb6+AALNg5DW
q45SehOCnr1AStLK+JGy7uf9vZEGzYdmOKsgrWMpjepsV70OpIzuXdGF2ZiiktggXCrtuVRm/jdu
0kGg+g9n/P4T9JUVtQsUttPRrlGrxza/7SnMUlvPURLEGetbec+cYpqHBfwZkRIjKZ4Q7Dk6an8s
hj8wrDsx6wZDzncjK6uzSrwsBgTfwYZ9nKJUk8qpnGxBgQzIU2Dl6xCAD2vSSRAnthZJNisPEIO0
bKdechFpWw0tw6TAouN0diLfsCVo6V2shG3Cap9WAzi13jcNox9i4379/+65SwuZbSc2mfrB7JYp
PpIeM16UgbuyeUpYewqITTmQTQ/MJrFmKeQgRcU10G3XBwzqgH2szygb9C+lq3D8AMDHNgHGmChf
AFZeXv2eFKCCaVwfhlNPnmy1vHRlCnEfMLhUSrQK8dkzc9RiXe5jhGjqzLjDuH5O/F25Yb6NcNRE
jSsNyvVvXUbF5LhMJ8BGpV9rMN4M6q/AjRLMG5W+Y+FSM1ijiPSUJjxbtXkEWEhNOTj/Ffd6l97c
70k+iQLmvWp57If9jk7kKbWd2+4DB6qD0kCmCXmo3U+YAJe8/Dmb2ReIBVnq6OaQj2ZpD7pQG0N9
sExmnsH/TJZMEkQNVORT6HU0Cm9k3yHWwdThFHcy4t+2ixMaTl3Y2ZI19BUHxNO6vqurCYX2g/aN
mapVwwfmaztIs3UUSfahU8MuxQGay1veWHUUhN5dBwsCSKXDodzXkBlZvy/kCBr+adQDtZvfmF8I
xNEZ1nkJYsGRsp2qazI4wUepss9WlMH074WGZvV2z944EwCt94cFw/0dSj99yupgABAXULgxHuud
94H0aMlk9pKdtoyW8qSGIyfx+5SLJsn87m3yfXe/iSPq5eXLjkmLIhEyOs+TLVqzD2WULmZtUXfa
qhxv4olwxNpd5jX9EX/pux+k6gjLvtZl6n6/7XkuB2Bm1NdXGtX0kpwiEpKj+JVd7TTDzeQ7C2Tl
iiun1ZSvCf8oloYvuVweyzpu3zg7z0O7shdnjQE6/sZqkKq28DN/6qrJa/EKKdC9shIv/VYvcFUu
UyXMKfN42omRC3SRZDpnc3GUms55JR+vqLEsae7fEyl8nQz7ZNRryPBzvCNpr9qqwRpFeJriQF6O
zejdqcMWB1StfoLowtulacO+j0xyrtVEVkjh0Tw3MrFXhcFK1A7EaixfhN1/Q5kLlnU2KyqUqRZ4
9FvUfV+YMbNqCdxxEOUrzu0mE/yDYER9sNgFhAFPCFG0xtlOy3EeHFnjonFTq5kkAJDVzk/C4gUN
g+Aqo2CSSue0/ylFgficQfcMKM872J1RRYHZHf4IKkDUcZHxsPdIzzPzZYsDizWVUBBKZjI8Dun2
fX0716OfVCQU5rvi6qspliGSJoUEAhBy/1Fcsz5UIJlXEPaA69Zg17EeaKckVLsfnCosp63crXrp
6z7+txQcJJpwYV2J/nOg4oVDj1hgxp4ViQIQ0P0W6SYL4VsBP2sjBKtmuaNozMfk1d/p04Ij90F8
/Xmlr7fZjc0bjv7wHiCcTTcKPBqTdJ/HRbSC000Qy2Gu+Pjytj4BrtA29TbiVhhrEPXH+CdqphEV
tRSG4+37qF6Xy4Ohm+5wHVrPHpYXOk1MrMDgzWiwr/JazECYlpnqFXe6g550OmIvsM5BD1HwfJyH
rMkNSELan6IpSj5qd12xXZm8eS27iSmXAKPTVKB4ZPauABsZOxI69wMsJ+zPWy7AOyjboKDnK7xa
dqBRLIsdXeZwE0i8okjfOMIGlRqvghfr9Jq0mpWlLUyul2GdDwyDpZuKZoxPOiMBSRNZyMHM6cEC
ewXwJWwv8XNXw7IBRndZgsDj1U+JzM4BLG3WaiH1fruBg3GuoYih63UUcLQNthpPor6sAv9lrwya
Igz4kaaFlF6AIeHlhH+wix291uuuKyHnajrF61MbUb+friQEl/Curk/W9sCaCZ17YOwT0bMR1v9z
uBWbDe3k1nMBZf2NdQmLOxhlRphA3HCEP9/X4NFsMlf9eRwMCox5bd+BabXDQeYhCygUL5jarRiS
lvLll5wrj4akAQOIRf5IsisWV86wCByL0dNJ5Kv5vZbMQuJO7pnuuLLQjt/KHaO1eW7Ln3BhO26j
FC+KsAsMl7L/hZ9uSgzwGlxUUqjuiA4ld7trqgiQ9dSAJQjDC1heF28hO+vDaFMEjG1goV/Tx77V
FE0U5TggGd3i5Bi99NEKZCEMwEE45U/L69NV3JD+rEPu4mdY7lMTGibFyG8pW+PMwhzviTy/1tqa
wv0dlgoH7yhCbVYO4aV5YDS6eB7H7D6OcI/bwhNjiHMoScag0k5OcxrgS/+D1EXKgnmbOJ6g4Ewg
Y0NW6swd4uCmbN8RhM01pKZxfNXSfUNqiXOKxHTgr/e0py1KphwjPgF3gTSQBxZleax71JB+lwRw
0d/M61nQY3IVFP4Lk5YxoBOen5MEHKk4Izu+hUHvu2drm0cH7C19b3u5zvbksR3JaoYwyK2Le3WB
+3MnoOLviUtdNEfb4Pu9dQS/Y8X1K9KDKzDN6M8R3k+jsA6MNgUEP0nu2OVuLHsJWwxBuZXgsoti
ridEQhm0Kil31lYLQGDn0J3MzWH/JXdGx3hW50/0TC62qE3QFqdN4dugRR9/BL6EJ7SxiUAZDMa/
u311iRYwCLbOctjAEppXUOuhVycAQKZZf3h650Fu6z9iXnrBDnx+V0nv/q6Z9j+6QTCgvCGaYibN
mMNSln5ZkN0gV2UV/rU5Y9lzys4+JeLMUqAi75l6jqZotllYvyUeGMTrw8b5KcuRfMi+XnaMPJfo
JTf73IRmWxMOJGhmzT/Gv55lAFYgjjoWKasRVjn9q2Suw46BZe6sX7NDn42xBjMcF7fCN3OXtlIK
R5jrBemo6NjHRUaem/xqp0gSyCQWQeJRmIX1YBi4q20SPQMb6XK9eIzuiTofx1/IzZVIO8AGMwtq
JmhJtq8eQvSIC4lZp1xhtA20RyLEz1E2ZwgpYLqr966LPsCtrNrUYgkx/rXPhKXBNDagUD7F7+oL
8WlmZ3zmZC8Kkgzska+2E9k5iaJAwm0yljFhprHBWo7UMPpBGic3OGWeXHBV415YkWzjmA4bC2zg
HrfiM2mNFMBb4eDrvayRW66ljxo1rJ2XXqad7M9SXSztp0joRJDLCM+uONLdpbJxrpLvhQjotO6Q
Vc7WzoMPh2hdWuS7a0cZo7F8JzUL07OIuyI78UNvv+LTItfl/smAQ3xaxjqHuw6S8A2tP797IpfG
YtWFJDdSLNNTI/38YKFBySvRN2OG84MIBa06+1dPjyBhCoLOnFSzyt1GATLS5tKvhti9vniLpO7B
0wGnXSi91tMErj6wSXO2WBTYpVF7rosgnslEjauec67YQduIZZJuA6XJQ9ii4h82kRdzy03nRPS+
e68810J0L85kCiI1erJDXGzNFAfhat4XA9cWn7p1gcwRTCd8bm/+nXSUgq2gwQGHe9PTRZrmC6ki
nWBmvEDBvvdFU+QqkT0xr4nbrPokVsaB9Lp2/MsO6+CbZCndyYz84N35KznijH7urg6F9O1HQysJ
QoIheliZ8lYNsx2P6GkRpFKfA6glnjS/oz2RauzVjjpN3sZvFnpkbchYPc0lwwo4sIUgfRE50dhZ
6b7WPJvCNvJWWoQZ94dx2f6DLDfzRjBa8z0CnSYHT1CT+BhgeaMoPSE1NnuT+If82HY1c53SOq2h
a5MXmClBAxdDVJ2yxVDsfdZDOLpqhwe4OXVmC3Dxwb3cQWRemnAnaR39drMqTY/6IpY7jayerrfZ
ytb0QrKsKWwzI2siZV4OXY/RRopJBAMUGsbw+2Nj55rdNAo6fZxRxlobrUx06mcFeoayBWrelhA3
WnKbYqafncIeN39znrayBpsMmVZsIpQYL+VdnXqa0U/yFhh62+ykgSye3ETiOQ6SsM6fLOvSxfgh
F4LGAANzusTjeamDLzCJcUOjTyZaaeJ5Q0RejCCaaxWKhEMSJftRe2grPFXif4IqZ39Wvej5Ycpt
y/xIELgdAl6q5I/FtRH9ugVdlxhGKBHvctdSf3rqLPAcrP3HzxuoPPcKro6mhpJXacGzNdY80fL/
4Dv1WBqmK4VMquDh+gVa/nThnhhrq3JDFqPpZdvdEXQgjDUvpfXG0AqWTmAqXObASwNsv6h2wxyb
+GDg0a3UUOvX3mlwxUF1SZZ9tyLWPs1mJuLmS7YYxSqWckZ2+pKdO4BTanreR+Y3YiMWG5NVtR8E
PVffPZlSfU+v8ga1a2xTgV8GOSn8gRuQSwDXCYrNbsTeFZ6lyiRcYGFbCXh4W8OhO2jqVtwtlAzD
3Bi/Gk37v5D+zjKisWsJlQlZqOrOiyixlqKbMd7DNAv7x+LQCz3px4DMctW/OD9avuOV+oHCLIvp
jFC4Ilslu8oYl/ZdjKY0NOhxlEQTPiZ2NUIZL5wD1rwha582hGSzm3leXSJAR//pabiMPb1APeJs
s/xKG3aXf8SbDUO2ATHAgJBsNvU0uNzFCNomV+Qse0T5fIjadei3jWn8T57PwFK4G27Jea6/g8r/
tYX9xefCW7M91I8/KZZMRZEIpH+l21HjtsR2KLrxAgKzHtjvaE2GL28/WoCMOSqJfU1Fc93Xxfv9
OxY58NL/H0brqi0icOHAv0wgYfQwoBsT7XIk5guWYybKbNHtxyTgfnDmmEngVOAIXme6etEZ6z7C
SGXDUI8FAT2KCF6uhiBydUT6jBV6evttnAt5x1DBIso0oizPGwvSNKluvi/9/fv1XB/KjPAm7qXz
SWRPvu5nK6Zwml8ta7iQL3TR2QUIrvDxiNeegeUT30012uXFTfbOCAHK50MT8TBhDtdJN++ugO3g
WJA/rgSG+SZqNW7VDX2pSFkcFKQoyz/t9DpbTZY8sYi6kE+Cad/Ky3aQvMF0rKrktvf0Uk/sKTdG
r6Rc2U2AQNsPWodUtm3utEleLQt4DmRNyGlAMteY6vMOkfYc9piJbubcbPSXI52MsHtbXdgtOIpx
tXPhKQdZXKDslWJ5cJEVTh9bPjRR73HWBLxwYaOyBOwuvH7tM73tNCgmxK/YxfAHvrgzGbMuEzXB
aOS7nGKnHmJZxiSLprQFTJyvYDnaODKhp3007WTm5lS8C9gqFztkqUjEXrvOj7FigPq7JR0vm1RX
84eYVt9d4hAtzFSeYTEnQzcTp6aecGZsHMrTzu57gzt33r0c7MF1UXvPpLNUbIx2wzwCVN/HY3Jo
/14ChXhZung6MOdDI9ZDnWSzMjxuVcRuAzzEQUwV7ZSKMUZdKpNRzmt5k8qUrJw9eVQXFtiXV5lr
mlFroqEwkg1maajPcJtYBubMC87hW0cvKtrTHtdu5TPm6e+UCzGyk4qkccIkt3lOWSUHtl+3JtlH
1O+yr2BMG4VzasCCLigXkUpMY32347vI1nVO6xAaeM9GQOSPqAhSm3YG5+EqZ0oPE0crOlRwdA1o
P4WNYBYMnbbcp1KNBK6jkQ8GxKEtwx6Fy21JJctccPEd8GEdhm2Sc9TRfRDxJtzfYeC8V8gcJS/1
ayghTKl2bhWlWlqsyCe8B/FosRRL1gmMWtaq6bYkRkYJ9Gb5q6EY+0IPnAam/GfGp6ExQhpObN9l
cBHJcR2e8xMgRItMphd+Gr9ZBguYWEsrHYw1VGjTnh3nH4xzmA9S2spPE5Ns18jFmdqBoQ6sxX9/
s1kz+wEseaOVTR0IT0PYUrYhyzgjnESRH8QyTxeoexBJS3Of9DIXuwBmt5urGQH+j1GJUFaqaWYJ
436InzzBneAgNnZFhPg3HNd2dmP+LfnvG/R5jELmT37ISZz4QsyuJMXGOrRaVWwW90ObslpLOBJJ
2+0K02IsjvBcsiS+irZvCHWVlArFG5+zXkWBJnbszpBTRbOcp33dYr/4FD4hXXDz8E7VDQHvp3ld
z0Phapqf9CgaxTz7a/IHNPpSie/qiuRbm1NlOEx+7gKHjUWjNN5LJv+wSr1MqdVcO5MSAIMamL8e
rsmKspwZi5tryVs3tIGezfaJpg90YS6e+xm1oIKMs4Ii+QkmpjneEa0ESFVboSf5Gl/iPgR/PrPZ
62VUAWYEHm/lKryy4dceGFVCIXIQpY5CQYIHSW/YOUVgDxNjWORTmxMoZSjKqNBVEKrrIe5s6ruN
ZIWHy+D9SjhwiSxySixFKc1prJyUdyVnzLsETB/8Qo1mBqmr5b3NeFPZ26FkStNa4auKMTERn8f9
r6V4whNWPf8Bcm+4e9mH/fFvcLrMLhak1I8FAM/0Eqx9R2qb+bQgG7B7x+tblWx21Ig4kSjtIz4q
LtX2CCudWxVHSBzpcQusjQhTZjwUTxMKrbT2NSuYqvvm9MWscyvzaCWn1oDFHQ9dZVk7Gzw/VkQ2
ykGppHYarkEfkfl/W1/+JpLmjn55H4SPF75WdZxXNtAaLbXSv6qiNpfYZYR9HaApcD2dtpZkJg3O
zkUccVtjeye5cbbmCEjDgrb2IB53n3bsF859ysFsbHCMye9TwUZA0OLs8Kx/eGjDf4jf4IfaNlQt
G2dIEf2xGLwz27aMfYygtoonlfCaJn9NmCR9iCEeatwoqt0+INXKISF7+Dx2WhAS3uSbjjxoBWUg
kZiXtCt8W/HFgJCIFhfou/AvYfXD3YanGCp/EOV4Np3kJpLAunHbM9A8cYjWt0SKq4IGl4jGk8j9
1x42HSmPsBwAOhlfUwvaz0rIlVDFs6jxOsKSHzwqco9A40oz8bcvJQ2UM4XTnJ6f61XqsuNQZq9R
aP/vPUUjndDHphklixhkANyq9vExUa5dUXp49D/w0QG0OWiQtlvNoAaLzoBn/UlhhyQQrTlbVvTg
uh9uROv05aFNScmy4fisZH0C9bWR66KPb91TxmHXcjQJ1WP2Gqdjt4xxLkngx3LdNQoLporxdquJ
dVc32SvaUACbU09Y68Mj8MSxQy0RshbriFsMMJtfzcIhKZWOWJaBkSwW5/3D9yu81IGNkrIogFQJ
IKwM0sWTcOyl9Ic6OvTbRysmNqcZjrx6nJJTbQDwLDDXbVe1eATHQKaasDiFVUY7PsFTRTw3Fo8S
vwp8xkrTgvV/l9PuIQfcmXuLX1e/oza0WxMj6dpwVh7VNvPBKiFink7Za9PUbWjxMjQowneRqnJo
IkLKiPSlQ6e5MjsB2EBkibMZOqPZ6YM7ObgS6wu1vHNvIttRV8JmiEjCyyf06nPN8zzFtasggBJ+
EDpaHyx1HOubbBl0ZT2DvdYJdMYsA/Bbi6Ee+YiknCz+xDiaXRjCwpV8gsao1BdOOgGOOJMYnN2K
injx5Ibmj8MUsDwMf1cKlX+l3lYlBfYGNQCqxpcJUQiA3v2urGgHdvU4oidesrwFI6cjt3sHyawD
HQEYiysHnQn9yZUsLBDGUGD9hepXtmXbl+YSPukii/rh8ei8y0kTQL2aCROkzKXOiyTvEse1Utro
iE7aEfhy7TIJwH7UbU9JavnIfdKK+QVi+F3qVreDA86rf9NQaty5nn2e0a7YwGvPBG7+yN7mZ9at
eXXc3Rtuci582NHJgIvpDjk4H9Jp5jKhGuEuTJZH24If1qtCYDvBWo8SoNJSjWtslyvM6JPykV5N
gs78BWlk+ZAm7xWTu/uF5Bf6qms1uX+cidfjo6s6HxrnQ0e/qE23w2mJlUlq6vShxNGvbH6O3jr9
ndnMqUYuAvjeatueWfeD0lxOe63J9k/ZDLEpI5U2Gy4Vy/mNwlsgVjFFf+PbXQlSVhu359iyLkGU
cpeJ5xoBp0g45xLJNBF3jOqSFlsmBiM1qfIAi0CpBUV+mahgCxjNS/Ssu/MYH1JAUddzPjL5s0c7
6w2vVjCB3MYd+O7goot0m10qzqaoWEpBsUJbFKJfgQWitI0sehmSLyloMmKPzw6x7nPgr2vV/pIr
/WOFgUPKLEgRgjOvROxyeAdoMko+KtvMlLMRdP01or9nqiR90MyQQG8Ta2OFEMWOyEo1tRz5JEK5
EpDpaU7S3jpz53Xab3dzpHfpDOzYu10UC9XvzLpd4JxxBgTPn7wT5fLWFwtOZtCWpgzkJg7U/04Z
EQfrWDqknxwpUTzFocH5tqmHFMSbxE/RMQ8YeC5LBkwomYCSvtkvYEjufqAWgh8wP6mpUVSmTiKV
ZDE8KqHVGBQBbuay+v1Nd+Xcr4YmFYTcahAzrhJbeYoZxS3HDJp8DeHf5H5yHnNndC3+AWQWlHDa
+/HjszsxU+NP+NrRsw5DOZbmb3Q+API1Db+e7S9ntxrs6RD8VEGQhIxlPAuZzSR4MUGiVFU6nJYF
NIwIRRU1XJQxz6ferC3MsVl+AiW8zZmk8sEcImQchrbLxiaFVc8OMYOePhJCxMN3Kx17f4u6a8m5
Lx2jjI+Y2i3sjnGtf+be8Nt3UiEdEQoSzsIntF+PzUXt/XO4gOJpjU4+ofdz+jzN9DQAbdn1B9t3
9o5cKetzcGur3rIE1ib57HafQDC9eQrW0RLAPC4aykWb/GjO6xcrbsduh4ISAQ+kYwL/13cfEtHr
DlKAjHJQer1C8EgrknAf72sqyhqYrm1IpGtCUrLnZcdH0hX9rzerzrF5dQ4kiml9P+N+VCRW9hz3
KMJtzSZ7J3oGJ4H/lq5u+RuHUbkCAG7WfgMqYutUIb4fFhspQbVILVOfivHCYIF9rKjZy1qE51CB
yV8CeDgR+FoOBEPdni6BJpTBrYWn1T4efvy44qb6G+fMGUCMAFwD5UOSABXBXpyJn36IU3zdHheE
5IjHIsMrKveQgckC9vp+ezk66VZerF+0XSQ/9lqeflCBQC4NFKn3bA2xoWaSxkP46brMrKNdUKym
G4BOE9OLpP9HKx0yxqf4c/bU9gcj7LfMTfSk2WomcHM2DoR/o8fp7VIJ9eUYAnwcbDUQShLwqy2t
R2jvphFvWUmrU67qInPoKBJwU6JwWYk4knqhNs0c6jZ9WYYzqSDKhWxDSxXQ4JQ8opLxwo/dH48E
X41H3ZEjTS9EdWvbM87w8hBcdLEA991ErhxkWZTrhv2mhGoY90acUFPKUdj65u3nAbeETAnYETWs
mfa/gpm9tE/29Q4I1mwuTjlvOmxW9RcFHI7ktrdcwmKeyiCnXCTY2zvIaiWhI+V0TeyCjs0iuk6d
4xqryx2p2EVu+NWbhNq/dAkyO/3ILOzkilgEKFTK/VYlrsG0ln1U5F5/pFyT7e6toQQ5q4Mglpe8
PaSstzRZyP182BfC2VeboE9Ehyv8CWRookLnN6B8rCqwzhgQ7xHfjmBhHvW8m5AIbTX/3m16z4yw
XZfag4cALrpF5t3WkLZZhnvRYs1aJJ1a2isBEPjnm1Lq4pU3LiGXexp7tz1WYuaZD0grpnZXTDJS
yVT9o6AfX+Ubo97j4CCX5Y/9Ayq+RSQKsLYNaie9gKiYJGs1WfGWHyeyD2Jwlm0WffxVO9+QdcKk
xexz81X093EqWvvNR0mGiNHCRkyVZjs0pCqyiAZbYLGRmAUz2WFos6bmube1Twu7kxbg62NE5rdh
HcV7dz7S2iP+B6ZX00VVD7AduT1mIvzuZUllYgTkcb46P0zbfvqHfBOUPhXHhldadnSkgE0+YWdK
J7r6o7H/xLnWeZvlOY+ij79UiL6/O71ZiBrGaAAb0LXr74cSPClyxdByBzAKXbtZ8o1179X7jO82
EvaSQR2bi7cS9gKDK5MALQxqKNfo9U9eJ9cAHVZfU9Gz2SsZ8WUf/Izuz9QoPAp3gU9s7sHiC/Ye
ZU4ORW7ZC36iBAXY0diqcRscCIItSPN0qdLrjXSE56kwhEoxH5+uFEbgD1XDCWTccq6J94x+F9LQ
PYQsaermp+rmV5g7wV0HCYJEkUPd0qllLgCOJRKj2pygiVp2ZY7ivKZ8o0R+G7BG7zq6wEa/B64q
9ATvBAsLyH46jYB2HSe6vYCA2rb/KdkSLc9DbiCcmJQ4dRjlM6TkGiD2JmvDz3mYlpwCzYMqKipb
xKliLiwh7QSeUgjVrvcugfNMWIlsEB7tBgp+gj6AXPD8GRHC+QaAp77FZfN6WQl4zFMPknJlDWNi
F745lsyy1iEAodxiSbZYUv7C2PnEV06ezt6x9CClMkyUjr2vS4vuIf270GPOj3yrRYwhHWSHDKrp
xKvoF9FURWfR7/s17yeRX8cb80JDUF1zKZkiXDjGAKw154Xx+/wksZXW8VBw3O274GKyNLrAZnLr
wKUxmAGADSv0NAMvfWckEIuMonvMtYIcSZ45agD7kOtG6hHeHXxgeNUNgGcLtOStuLR0VCVkJRm8
1kiD2gT2AwOA0xLoFR1EneJUNGUkrcUkpiULWfb3ztUF6B3Lvt7NK8LTr5mlDkAbF/Wt1szoWuOG
bs+JigmWcp55DHxxu9gi/WS7fEAGR9coSJrZoyPFR5EqiDJfMTG6Af8Jyvk68fbqmbPQ8S2A7omy
Y2QuGkD92sYCLUgLkknKKC4tz0xQ+GQvUiYqE1vqwS6ZIaKwSxJmgMSFzzP7tvBoCXatu6KuSqOe
+s8k2B4ojdL2OHMB4+i54fFnAdjx9o3Rc3XBxkr5GOa7WL3hq0EMwfgT4WvjVKiClYW+qTKQNF66
rZRJnCshCw6E3wAICE3kqXm7TWdo62o4ouVhUaNA95cglxBk0d3m8PbzVpdjFAC/IOl6CBTvWJtv
Ju4Hkftx8T8k2Lo/GCprp5LrshqCaFpYB7GeAjEjrlnZC7PTmOO+ztTtj4XIGm/nKXZCykjyOQPI
0V2KjVi6MGW6SO0ZtWJovUchBfHVSI3XFpnIluWqYBI2v/klrNEmVn+4GZBbAN8clb3YNnNT0+Ff
YmJQ7kPDE/5VyffEt2uG5PszrE6m2/Lovlr2OUDfrobuGhjFLxv1chzL9E8FcVwbopmlFq/Uxb06
FqhyHGA4QV7UindSxbnF5LW0rEM+bgDKHTgjIl4M+J9cIgj357p3vhI43ZHcF6lLLjGDX4akmn9g
hUper1mkGlGp92GTVbAoRBcDr29588LpU2U58WwqfDQ0lQJLuFDQRHd0L5AR2ZkCir3qq42LUJEw
tde1dkmqtrJVA0STkxaZ17aFHFDTOxV0Ym+gPd/urUuvNxcx70AzIdMQzn46eNqXC0piV6PGx6Pz
4PkfM8rL0gNk+46//DcUB8kzVOFT2XvlY+C97s7fbAaeyrSpK5MI2xvfdSA8XDqCmLR4v8QUhBeR
KA/vXEHzNg3bB4wmBkv6iGDjRs0P9BQDH6EuYTUG6wZVbuUlReaskQ9XPtFyIZesn23/zWehAHq6
5nsjHeZW3EIsO8vp98y8xSO6pwBxeBTtGRQgDWDVZgidUfXzkEjF/u9simZN2EIoZSQqZczOmM6n
C7aMTrlh9y/A1iyXwLYD7JKOgvHbbJpKB2I99zTE1GqLjFstrLf5xNlH2wxe2ybSnZHZQ3yRgkR+
+Nd1QkwWMlgQrTp/wT70ZqhYxKv29EeLiG5FFo2zqpBym6Hl2n9KQQIo5wCml3ymEP+APezpsesW
aSZ9fPvR0uUPnsU0DwNWm75MMda8xKMHY3hlhw71sbfFba2IFjO0GxVHdeHG+HJEQ1tM8ldD9gBd
GbqKDhKYZzwsm6yl87E9UGRGWxkaTj1f6b1TtPSBwtohh/WFENRxQveEwkUGWg9A54l3VdPAc4p8
lg0cQzRkT4x+T0CyhtOm+X2uWPuXaPetZv3dddp7fS1oDfLiayQDaX5prcoJr27ugyNWPboOKNMP
nGsUzw97IQWTptxEVCvLKYf2kTwWENXr990ihxs0AltCLSYV8Vb+CbgbfIZX0Y0zJs7RYauLBUG5
peaofKEsJwLoL3K5nBg3ZR9tIYEHnfunxRJ3NetL+rg1EDVE+DaNl0zNvnsLqtWRDvEkgQS6utns
JD5mxJ1FuSopaeNygAWTsDspjRVktekiMZTdmQ6TFNhfO1CXL01DsuXmcU4Jyx0AG18Ebl//RYjS
2sxQZjE7GG1Tz9kYai2aHdCQEm21puZNkRqH1tO50jUuwmTBKXH9SYFGO1JBT5tfeI6IpyhBNYjY
TAJFMN9f1e3aGTBnOyzDiMQ+g2sQVCG4STwvf3d4L50m33eS9MbBB7jWLeMnKNR3MJCzO8w5Z8wH
FPtujCbeGLIVNi0lg5/AcELCMzWzHp7zxPEgjimatuQa+kiElOOb8BEp+ViAQo1SiLMFSTayzNQN
feP2eQ2OC8/22khtbPW8oXKcq2sTBjIPL03YdBq6q8j+Go5sUOYHUH3mOxPnbHab2g/4nT1tyXGJ
skOesNgH3l/+9fhOSeCn8BfUg823bt0zZvldLjgGWwWlEiT5gg0KS9RVtqVvEMDQJUt4+Kn9d/U0
ftufUw9rdJt2mbBJJ7lqnrVHAmjymMInZz+sHvrN4cu4kNf36Xw0+q0b9HGu7kTlmv958UN9mclq
ELI9vDFpHXU1hk3cTiU7JyfxfbzVjJL9MWt+incnDaiTttUmBPcxybAVbkW6LWez648OeV0+ZLH1
MeokOrhjfo3Qca/JB+s4vKQCuqLHjzFoElj2VZhlHXdEALlP3IfhpGp3B1y1ly0/rpIG/EfVtUle
Ji1nZQbLwVm0ipIdH6L7rP+qHp9N0tDg4E4CG16EWpYvmICUzR6k+6kyHS/Trn+jBun3SV6IBzqX
tB2GsM4g1BeCXW2bqdoCLK187IrLOY5d4qSNjCq679P6d8Abi077x50v6xkEEZI5Q6dIV5JGWG3h
5itc+QV2zMQIClxjlljmjIEW/U/7h9g3xe6q7ztntyQTgSXOWxc/kwp33Le8Lav3sZH8e61wIWLb
XTgxWjaiq5fnfW6z0g6UjtdNpyJaySQ6rqFA31yYBleBQtB7MJrU7TjaLZIRjswJ8m4rmeng5Xzj
Hm+PecOZkJGcLw6b2/zoWBeEW6btRRM5fIR9zvfTNMYS0Yu0fcUdDVoq9vap2e9Z33VCgMweKjVk
IRBZ6uN9Kd8WwzYNmpZ3iB+zA9bA8OJUCJhLbkqXuszEpePqZbtMEbX++xK9MeLQiSUsXVevjlmu
T1OYnyyanoOR+pnhoe3JJ+OccJW3rzs6zzoVNkLSiAi8kcoFIJ5mxLnhZw7QtGOILlxNYUr4SlB2
Hmm+7VkK0QARnlscVydMKzOapGo3+GO/19Rgexh5ghFomI9hTK04pix6fkTV2ygOHh0dbefqrjBi
jUB2XVRA27KsGd3UdLD37pVD/FClOXJx7Vrpi1mDDmocwL6x5NtP2VxHSEnS01tAn7K8L23X0as2
GZn5RCjsdxIbtaOVbYqyYT4dcTtmtTgQh5meRsO6cYp0M/dskZ/3A1KNXr90o8049xUwgIVRD5yk
K5reqzwWCTDNqQQ5v5LOi1AmPTMyU+gkoYLt2UI5UAsMdjOXnDUptoiWahYFY8f24QPX6XltmM3U
9VyX453ZJTMRDO5GmfN7k8urNZ7Ib6KU7JF+qxghFLm58Oy5UZzFmgr0cDM5YlnNRaKkB7SK9r9x
a+AMozyyRvsTkSVpjO3dGGfJkd6t6gdMMrZWTGtpf+L12N+q+c5Qi7Jm+oNxT8zRZZ9F8kd2jtwK
ApqZOWJpv9O3fpJgD8L/TgkNeFbnRIDwBJA+dYHipgiVkqnolKqrWTTDeRt9C+D/vHf0ohhuWANk
B/P2MVR0X2hGxbUIwuB+SL49B6KwwB7+J81TDQxEz0HGbEVmIUJVJIHZ3457T+hwJ5o8VO0cj8xq
EmHfOyJRvzdqNRlFW7cfOUvZmt8VVCKsA2f5rkNkKxxpgmm+JLPUNzP39hMls3JOFVKKdvf6zDMh
PVPZ3phoQVf3amdWe222MTFN3OMNyllawxgtfNdeXoO0upwfE+EaKn/Ab+vCgpYf1Vl7HPZTbjbh
C3J9fpOI2a7x2qwDAZmAH7p4cjCDjfHD/i8xRKzqF3G6k4HI4CNnmDjW2hAKVef17Pvk1f0gay0I
yX29afPGTXHxNaCo1SffBhFEBlxMbbx7X7Duz1qqn/vMm7vtX6fsYVt9cwxshJXPqBfvbNOg8JwJ
Z7H7jznDovo3nv8atDDY1Bh4/xX2cC3BsLQf0InLJo46pHih6yQOlt7NugU5b4pd50uHZ2NPORvv
K0z5anj/1LAZDdkdnME66lt9SXzBsQCrJL4Irfx6r6OWGsZg8IvZ1l6VhtSvYS65k6P1m1xGTj2F
IA3ZrrPGTZtP4POwC1n/Z2dk5HI0kLgnf0ZonNU20BBq9+kCT0kil1h2tw7GFoCqAo74GYAAOAl3
p0Vua3D/9Z1d93gc04GcZiUE7HtrbjdpWY33bbCscfyCOUeOWUzuaamDl+ovkei198mEyfhBjz8T
ZIFTpEazctzNmMSDmSX6LcJXlZequORrR0hL8uyZQ4qD8wEoDnYYZlab44fmFiDMWalT1bKTfHyd
lWrO/a7PBgpgmNEy9bda514rzOmsN32DdHBw2jq4v/URywPPxiKCEZGVlUklmj4BkAIbZmzydWWq
hK6aE4qhO8Tz5tBT6g7621/lgpxb0lvHxwvWgtIxlsmkovOW2c5PmKJUjh5q5tg5S5xfZApOYwgL
xS/3f0S3ytLH379mezs/YblWktt9WRZAx3duESMdrdAseTm9/Lqk2zRFFJSJoWRDQxuHZE5gIB9G
K6dzY2U/l5TM5U2IzscuE30tNgLVrNk898I8C7AAS2Rbwf9xVc0hroNDtISBdGJ+LzRx0eeQBtgf
JKRwaxSthUstTbN29qfiAd4QSC/Xec10GIRerI+JMPZ/sRmkiDrY3COs9hfoHPneKIo6xEE0wYk6
vg2TUBL1RTlDY14323BTfHQ/cyFR9L9OVp2bAa/RmV196bmXFBVWzQRv+PAWjGtlO2VwVGiN2tq4
ZfpzbVFcsPXb1tDSxlLgLjlZlO9zk2fWhgWDr7vEsRsUlWes0ykyapII6aZNNa8xa5XSt9KZ5Luq
YkppiDy1pZod0YhVwAzo2qg0qYkofn0a/dZG5YjJtdC1pTilzg7YGbfq0gFZ/XTBk9IxceVhSt0E
Qk06l+/KHQkr4COBG2fbXpVNNJDiPFSKGbqNxURH2fWqq90y1WRM1SeiLhXDMoTK3g+ziPiE9yA8
TWBCeuGHBz/+wTHyLkNzu/HWq0NgvsDg+ypY6Bphs5IF6Zg1+ImnJp5+O1zdncN4oK11qleLjYT7
28uh+31CgjdH/5dDWNDA4Gz0pbVcfjDuif0SZvmTMI6lEyWTDfie7N2w0bdKLeX2xeCxOX8onX8p
QOncNPJPtA/rj/SLiRPc7lGyc41anutah2YivOjYAfCLFOxnNZFnImnor3K9lDJx2g+rHT7kOlqj
DMmfZZ3fU0S5NxhXhLULyS0k20BATrYGWs0QRxF5CDRvKrMpnQngwG7ZtfcEc//EV6PRyrjy4fyd
WJVl3ZaABvh25Gyi5Rfqbq39ptsZRMhfubXs/UbksZ+F470HAJ06z4yagBm17JY0JLdmKIaQqN7W
UneveR4zytrKsBjfoDFFoFUIhcKltuhHX2MUwV4x8A4+mNTAEb37CcC1JtX8EZpTlUTP47GSN+i3
rIlYy4V3xdqIz5yTgxcQDfYfJlM5Eadkd09bpZnO/aL075ETe50IzYmBpPa/HOo1CIwg7fszlR6m
fvzRGSnYRHY/XQau4j9dx5SnuuFrUiKHZTl0CZwkbw2zTIlgEagW9MUnEcJDv1C5ZNZgQHyWSh2f
R+uY3N38Z2EmSfeetuRYHpHun7IfG+NQMv0BKMzhni1R3c83qy1aARnvKD4vqnv84OUPs7IxjqkD
FXkOHzvtQke7XtXXyK0KrSL7XA6jIZGY4gZ3/Ia77jU48fJErvBqFX3JVppelKpOuIIreEEydIyN
ZXJa4Rl+5MYlSVZU6BeYWJ4hJfm1TyqHHWT0TCjzBZdqCK3/wQEJuF6te7XpohpxGynpZASz2xmN
TtOWclQLH+9ojqmLU6hYRcJC5fQvJy74zkfUzRCtE9fNVcXcRRwtO4BxjqWYrjkNp5hh8EuhMG29
10yDqNu8QMpfxHnU9Fs29Unkw0Ue+1tx/ptsnxmH+x/+9BUfcSdi6JPaNPK7NJWnYv9jUSb80lDt
kanqpz4MSD7CuGAvmYn79Zb6bMRCbkTjbdfbTXHYUI4D0ZwVgnthz2lHaUwmt6Jta/eh175x9zQz
fV8Eu4WZzLv0G2j6P7+6I+hLwucEPCCto1bk3J+DuoMaTvGEYAI7qCj3dYzpB/Hnz3aujg1nvejo
d4KdzgD9tlk8uueJbrqKkisCSRdshODC4oLo6O9rrbeOV/lpdAfAXhWiuX6T/u7t0eHTuN+ZT6cm
1Udm62TnYimYvs1yuv4+VsXhum1V19uFV7pk2mjMrl7+9FQGPK3LH5Ew8CbkMBmK3R/P9GeUEIYs
+lVUPUvBRvL6rvUsXsncQ4Nodmd4hPvRo+dJjFmF1y3drG9q2l6tKRhjfrhAgbAVf1Ou6gIbcH9j
FGiyx2EE4d1JIMLYdtOPq5Sh3hpypv7HM/VnOeFn8B8LFilRuPwOZhBtDM3r+t0ldVx6ySagEsk2
xWjRwy1/badebmQ3Dg4NISEyIW/PzLZ9brACSgtDNGxtp5Gzk6d4jqeVXfGdscbaeDmRQAga4t4O
zBfJYTFgFfDqek1pWBC3FqW4aMzb15qsWJ7lVsy2GtJzit3iZR8YG1DYHrGXT717d6Fb3luWMfZg
XZL8Q1bgGbS9q/QcjKQ8A1jeTi0uUWCdSvRScWC9geP+qiQ7xpEKFcIIOnMwjcVy0WuwbJehMQGa
RTljTaGtdtM5KkNnoPEEFdhw5RPKBluODsqtyd33BaR906sIbvxJkwEnpya8Qn1/0gHtk5/E0xNr
niFDzFCL38HvWSJjc+NnPZ2HX0Wci3hUHFqhEtOPNjB/pQslDbUSe+CdS3N9hgVgWSjo5lv7ef52
cQuqE9xtIfR1w3VrtfO7JmTlQ/C5dFBT/OVAImX+ZwEwcvw9ChcM5bvKj5PS3VimhsuS5RBKDa+z
zEwQRjSioQ8HgDEu9elN7djpGxvML6+sdJG5BsqieMSRJAeqcBm5V2b1ScByFMSA+BiSI/ku35QZ
RYPjJ08d70Q4xNolnxacwN7L9sjcvuQX0lsCgemvc4Krn7ve9Ib905ECroDz2v532f1j65q/Yov0
QNVE+Jy4Rlv6RGqv4NhLfchOMKaeGqzZ2B3Os2tIera6qmPM8M896h3YoBnCsSVwdJGr/x2gO3VE
2aVhheQKOifLzGxIoiK2BKGHTWRAJvOuOppDh7x+uCwS1VJQF3mN6yrFMLQoSoSdLrGikdAmmmhm
4cNw/Q0IR45IOLyANi4zlajuuc3MfUUihnRUffYL1UIXOdrCNe6feLLguZzcRE1odboWLkvLmg+0
Jb7JfhohHMOd7SNwPw4t+4XoLv14uduv89nDBOM4du8kJLdUZZAM675UlIKcKc9+mQVDRMzKfdeH
CPuTVHNKRus4z1wOjkAmpSbiMao7EtnqSPLVyQsoYNvwkgsnTuBGBjvtEWNo/0uYu44DaLdx+wb4
HXetAxBdjfLvAwB9nT87bk4h9vBxuprJ+WEzv1qZeG6ZfhJbbEV1FrM9dIUwuniVlztEaAEb1kvY
C+iKR4vcuaUUp8RNU/Sb8H4SaPj+SZqojsIqzwMqWSq+Op5ny2/Wg9Bc0fMyTzcQQ/gI95+y8jWZ
GeK4ueP/7WStrK1aqXVPpXj7I//YPu0s7OxrUCYa5n7uewI8b+oqlM9TtNVZbca5nNjUZrOCBV3N
CKJC2qDTtMu3V0ocm8YPFiXnL+GwePhK2KNKTlXp8U8AZkSAfIEwCyCO0sZHOr+56VioWr5hyntZ
1kSUjEIBjwubTG/Scn9MARvTVU7EuIzVAXGTXw8uRWeeyNUsE3nh3oCylods6Nli4AZM5zLlzjm/
BuuuoOwZsJVKJ+Nh9n3kiU60UnShAhbSrYJ0gX2sScVSNFO8r4cRsH7/u6U7EZzpeY1yRy6GLP39
SZxSXUYxFMSo95VjSQftpDQPNmriiPvzSz7V9anveinOnjdVaKXbqoGYsJO+pbMaqaGxKuojnFRA
S2ZCjQ4U86TYN0rmny3canglEuO4DlZHJD4AkGhUhSbGAvHFccLSEQ6/tzHgecbqd5IZSArnVm5E
p+DYBn5KMzMarkZdDPm6Ca45jeDtbJAYI/xVeu9U0PHu1j7/ixf19JO2bv/QQVYRDpnkAspBWnyx
TY0g7kt8dyvOPt2+78vQeCffJaBIk70VYiFSwpQiJWKZDme4Z9+oNQTSOJ8cQc4oIi0KT/L/NXsv
k1cjcj83uUuFqdadB1iff7q3kzCoSPF7Gdz5OA6fXa4T6d+ptFlwpgexmZntnEtFohQNziuIg7Qh
368u1GR80hxYyuAZAahAwU8WEw8F2fV4Q0rHRq2tAZaS0KOLBmxK1mjAGHTZSZXs7TlsDdtabPIS
XxGJNt/5j1YGvucbhEuw1Z6jRE34wFbE5+G6mxtWjk3JIe7YeVU29n1B2VJrhyjnRP9r0eqRzgOB
Nb+lhFqoftb81VuSwpw+9G0LqFR3g6WziMNmrwJmA89c40mCfhJ+O/uE/GjxpYeJHIMCxvfPp8Zd
QS/rfETpRkSAkmuevhx+J5/OEiCV0J7KDCrwma+wVRF4y/kzNLNH4ef3btLYsuW2oyofUhTwrzgH
TaZ7plPXVg5CZcQTjsbIBxn+GM3OhzoI5nCS8kOM0UP3MhlvsCLiX2uV3rAH++/mzvzPlJGxy39q
zLrE+MlpHi+VnIRWoe2gpXnV59qMkN0bEStnulrnH93xtIQST+CHM68MfY4Xw2XLchQLX7T683Zo
tA6EirNWkQ0jKejvna5eafMxpORHz4wxeO20WzFM/7qk4uuC+/Shp7xObBkIIuo8WGM51TfwhnTT
pGTDk010BqpDksKwb9S3tttoPjLd4evJElmCBH56TgRlMex73lxJ1zFfH6T+KOVotK3qHFfsKgof
3bMrbUNNDZoTyziKOK1JLO+RxLqpMXnXDFgF9pI3Z+UnbNwweSpVCBuP9N8dXHzBIOfN8VLGYbef
jfEiRpSpJmnsC6wsfHw6PcL87pjBjcP6kaUGzz7Jxz7MVn2JmykCIgEqNP7zqBhQnTcKp04xHbSH
EJIP9nkfINZRkEdDqcWMzLjkic5kCVGX2TglSfRA2Xk2nkYV8C963I98QZgPzcwEIDF04gAoFddv
gF5jwRsHgHzOQTTm4N4Q/x0u/hV9tDfaGv+03BIB5F3EBwGJ/ccS8+KGKGg9TCJgSw0rfhPu62L6
KOzwmoNywiK55FFOIGqiIfBZQ2yRXe1py0q3ZK631yJbid/V037SHPX99InZtUNn9PWNe/H5r4MX
SHYs4SgFhEG/rnE38Fv0He48L0H4oTMQJ9U5ylOCOt3kD/lfbCnw3o4QI9nAXhvyBSNl2mB0dBSB
4O7fBfAK2RwnuOm81fT04WEFq5KQ2Uq6wCRSgiFwyD1lP97owi3EP1FItMB2ccIDpWchkoV8VT1p
KB0MW2V3ZW0sLxN+PVjTZp2N+SLc5nh2MHt4fijDHK3uLdIzAF71mveYTArte3Hp2NaM8LuTtBhA
y/4o+Rg2AsFVZhCUxI8MFALX+e7CpznROCXhI4KpBAsYEuQAKxjH/SwEc1CQPVgXv/GP8POHXm6Z
tnulGhZEYhZIMzFIyJzrf3OXSigjx0UAg8iAohm3W76wucQVgS0c48s1o+9qV6dHXO4u5b5R+Cm0
bohmP0QqhD04MAicn/EJVdVfXL5m0e7QENcwNWsDY7Xr7k2ayhkhkRhnTOIw7/L0o6NG+ajCSvNI
aaPbE5lajWVePOgCGsgXpYBz04kcTkVk1r17ulwvV6hKmsAbFTRW5K7sihqKea9MVjWn9yOzdqgN
SwvhBV94HLM0CMBW4QyGraaZZV4P2AW2oWFbvaKltVq/aUfrJPoau2dFp+t9SahEmraJv/2ARgKR
l7g+JKPf5EbzMVFvZRQqTNdHjUfeOh2hVaupuBRu9heSRZyjs4zawbW4WC2Fzi/6t0Yb6gjVHt04
dp1UzNQmv22R6BK+5SUPE/lZzZecZn8cfS03VnoDx17o3tuTYt+ci973UIRrSgR3djMtQvx+EtY6
laGij7miVYiDsPdlIMrEIzXMBQy0AURPsUcjiGtuLF1PPx88y+AcKLq1eXJ80K0+mCmmyXlOHIJO
LNKbLzo8lZDM/tOz0ida2sGj+ilAu+03VQrgTLaGmeqOHHy+Dw/vjildwMXn5ImIFVA2DsVWU9ic
dJR5/a2AD4pzubThA1IplBq/pAiSiYrYl7VNgAO/ePgKu9h0LMNnn2uNGzwmhXaXL3GwjrqBjv8I
dhryCcCstA3ZzvnN/d9rW+2D/Xf8t2E9Vnhf5/wMdaJ4RN3w/wPTTueWNPobL2QZyb1LGQPOqyk9
V6/D5pYteU6rZwnujm7o+M61kb+BRzbxYEc96iSFRHmxANqNXN0Ri4tapaDhw/45HkA4zyt3d2OO
jACDWnzX1y2hXfS6bRTwcMc5G8ihPP6o6/zZDJii8H4xP27evCOizuVg2gMiv5tp6dA+90LivDJy
vtBQ7slISpl8yD/kUOyzL9S3mPjc41KuRPpVKa+Zh4K6gcSb24doDROrte9cByryMk/c897BwZZ7
SgzxMjtBTSzRW+GCEdZl8fcgHxXdkv/e8aqGazZ4vSPQSLXTXI0vWVHAQEtajqIAgnfc3AUV1qAO
bu5EnJhjv2C4V5jdysAPaE9Pw08lkKChZUhi0g+6bK8cgfH5hrtZNWpnmoePIBGxkOsgI+j1zJI8
21bgr5w/ZNM21//MPHVevdghXYq2OU/tDaUEJ0IfwJdxWewW8GrJf8I61WI82KvfbmEzm4JasGyz
BX39GLY9ES4WV4Rk2e94lnEY51i0EBef/lR5BdO2Wj0gIq1+96JlZjimZDztk1eInvPnI08x2jUi
N3ouAkgCefm+14Amu1DSMDrQIxqZ9HFQhL6dkwd6NQmCeGTghEPkKmbimK9UMiG0JjHDV5dLo7I6
s8mjzd3aOyrj1VtBXUlD2xz5FpUAaFhjvijQ22ucBeZxE9lsk80ccQpYj5L/TTER9HFswqooq8kF
p1GhnA2llBdb63dkLhhYwaqww23QJcI9k+J2vt+2xAPoBxk9U2cNVMD9r1cyWhOUvCUVP/zbNdj7
tvi2Qxoltwi2451nXHJPmgG3rYQLDThXDRQS++wwmxsXkKnCbkckFLTtrsT0j8IG0b9wvGVHw9zE
v5ACl4wKSxJRaOyEQ49L3TFqj8m0a7K1pZPVc5hBw1WUEBrH+pqnu3+0qBOp0K5tKvzsH3gsFKc0
CYF/r75Qaxsg8yGf/MQ1fEllBZxcFx5vI7ScGOMtf7AFjFhx3uCr8pMcb0CZT2lP+cSpP+rkBPF8
MpVmezIbMNsm6LdNFAAUi9b8PsG1W+RIYSDB+NzynswLaetbA/niJTECcK/8LjQx26RRGSAvDDHt
4KEjQdl3a+vyJQzs9sGfKpP5Fr6XMfUySSxH3PFbLPjz6Ak9nyKRuwJhHIffqj/EFs8dBpjDDQuV
mh1hR0XMq4P+uXbd3UFlNIpFnaG6iMypAT9h32gn9ARqQa/6ZyeIz/x4OWRR5Phiy7BHxDqHl2dl
ngzFRUWxoEC3ShcFNVDXVWQGv7ZBiN8csQXBewppRt36hugCX4yb6jMASx87lZmBgnWTMj5PPM/B
XWdfeI42dPr/kHDuF7qkKLoGV8J7HT/sY0tTidfGCHkxWzXDt8dbWG57VgD1XD20AbftC2hadDzO
Nf9IxdqCHuzH2FvQA0YImFsEyk/qpUu7lDJJ5EnXBU9A9iIBwztgUfc3C0VTIGR+Z+edgoGOgHuV
CF0vrBRz7qjPXknNHIhiZSurqLj0GJZFdHiVthke0knOr2AgNoRc4n+2fw8vNcgV139h2Za79WwJ
D6TSevMj3WDv7k5Z8s79dX5mhISf6X85u1FdtPaANNkDTgMT3Yr0tu8Mv018dBXxMSafoi9mcCDU
MJlDyvQwOH8V7q5k6nrfgy1XQIqgFGmZWPfW0leGINRM9+VnbtjIIE9/1UHxWcULJ2uNEGkE+w/g
vps0OL5PCxYfefQXPehJYCRtSIChdhsSACJGR1MR02aU3UhvZnQjPUU5fXeFpUoHusrAaG6URB2G
ssyxypLutcoxrvmWfnfnfKN6t2/0DB64atUmklWWJIJFdHnwaHHz0N5HA7tUuCv4X4QsnZbEk9vX
/zK3dJx4Ddu8mFjCUExVgN18YVgojiqFoYK3IYpLusFojIHb/7EI24WVR8H6VVIn8h0k1NWn70cn
sKeOj9lpXb3YFCghRWDLl8Kltb+mV8HQAB4bxs4g/jPqjsThrIG8oVjDUK15f45nVKW3Cl44z/1K
ohhl7EQ3sPYcXFNb8sYvangZFt3+kxOgucjqvlpNpcT2RoG+I5q659itWrb5GKF47jBabqG5sujr
ceP74z1d9JrPil2xbTezxmeR6usGGki53sUfIYpffoI8e5OrzoRI8imtdCi05HBtywRfSq89W3je
CsDkIrw/46DEpY5r8wddpKp3WHD47e5Y9S4endCyD8uwoPX3m2UW+w1kCxCedm5WzW9zYXfdz2di
cdItNLYrB1H1c/cesVTclhXJsbtBgnNkUAqXbSRKOuAILMmgyPhOv1GAxoOT1ShhZ9ChiNAbPUCw
XpQ4c1rsgElkHgSLNLELmA0AhN1SaZJqNUohKoaoffT4FH8MG5YJIiUpznItgS5WPDIX95IaTOfx
IoDPzuKtll4Mu3eN+s3vO/8WQtC3lMOQ8C/ax44aAweqJ7dT0/ZM4fAmkaUpIaDTapJpaPP90QPl
r4uo2Aiyu4jKea2BeZtUg1xqQa0B3OrUXcrV3jgxTnpAaT+bvKuJ7zCjMnI02g3u/Ml6QpJM5vG9
xZ7/gldfedggPwBApDPvckU+Dv8vmIf09dxcut0UrdXizVyZ0RUFbIg4Ck3R2YpTIZZ6iDH2JEaA
j1qoW5eqNEsH1i/DjR65wLhvlulOJdXjQy7rYV5RIaUuCr5ddIJwrTtf7Duvt09NBDerQ+/rHbBs
dNpr3mStyl14HmcPtRGJGh7D0/bqxzeBYsoVXtXpTsKGB9FNKWFsHzupkFp8AqvfdBPyu8OR4rbi
BCEi1ST3/n7JgxTAWidb91No1wGb8uZ6HKN0EJM/p+Qyutoy7an584LImmVVXLM5PzRrz/K4lacm
R7mhDgK72vWSiRY9fm9U9OxeHxLv8w8/Hyc8x7Ds3SY9O2BmThaXHYu7q/LrwzCwMc2nH/wxjbe7
QgvUC0X5CfbNMxRZHdhi8+U8Dm80MfjmkCjVZgcDHO2tBN2CNpB7ztMDdcXdnlUgY7qof6sgPnip
R35qE42C9wOnAnj5Er/RF+9xoKeWfdfJffFbycrqLBfYSJtN4Rc+Un6FYjwIBvk2EeELeeXQFXAu
Bfz+R6Q+gVhm7J2VFniNwiauP2LEMmJngTJoSDRfqyzs204Jg6KTuXP+4htYokLDjg360b5Xs1e8
y00OE813u2F6EjFwxSKFUFrwhwSc7jaSNqDBY8Ic/VqaWoxBKex9ERNLJmrgrLqXigB4y5iRv5PL
S3bXuh9m+7mJLJt3TajZ1YMxMCV6w3sfn3BWuF2jfKW41oaOQb7R4Gdzqll7rc8r2qL8f5HTFHRH
kdbvB/ZViw/2BRNmLt0l1SsiUE0e3NM5A/RSVyZ/oEhqAP1VoRbtXG6U42BwV9SIxLI6UJL2uR6a
/20GHnkabCpUGiaenTh7SwmC6pInZF8eKr0OAYC19gBBjShl54HaEC6ipnab3e2vvjJQl3a7Vp7i
D7zXOyhPDUQPdqYpUw2mzAxQ5JuE4OJ2Zkps7XM62+pMwN4GzNDcn2F72lEAFu78GbcaKX9/Ilrk
NuldsUtidQHTxk/7U21HDTuXcShmvE74Ha30dKT+N2cMOltGrM56Gja5ALQOg76bKaf8dn7YWkOq
RvMYcqBIIpYoPFoiPC8b/hElDZ0juH4VzTY109M6bI5eQnjQ5laOVCS8Vc/3z5ZJLj+kCpmI1k84
Fpdil1hqifXAfv7DqwcNy6WS/gT9PmSrejUjawB5g3NcMI7Y+OM3YX9d/U2kDGlMOfwZ4eRVm5Ha
LXA8Yj5ywPm4N8Ge/CfUICG/FzbTAAR4FMofk3Tt9wYSP7FvT74ZR/CGhQVehjiRN5EznNfsXC8f
QBvtviPpgIJKVnrgrRjQu5JTud7NvbD0S9fBijq6N+NDqeovKN2fXt8Hr6x+rDRC63xVA3TLh9lH
T4NBbkxvYkIqy8j3rridXOCW9OmcOFGqJtBCPx7TPa6CTgy182QEwkQ8zsjsjd1K0Kj7PipGkfg+
1ETki5Q/23DjEj2k3OzIdEigPBSjBqi30bT8iiHEn7JFuisriHqZoJsQusJ/l6fb0iisdIJ2rT8u
7nkFs8Jp2EQUH5+2Gck8KAAGGFy5oKf0hPPEIoV4EdH89eJowIEef1ApuOhy5NBxZ6eyZaExSSQS
p5yYO8h+BfV8W83DSoZ5dS/WnKETsjSAsELJtRvkz9ld/D4YHW8NeV4dCk6rxt+jNRLawgszu4CP
Rt8B1oLr9eo1JNpaPZq90RUPLkGCraCszPv/ZhhRtaLKf1wLWlifOnvMUKfHOBzvkJ6lZwzfQhUq
RSnQErdeqxQAEnkZYhaPqnPY8QyOUUqjsSQf3LGjZHc3LJ1Q+CqvWsimQ6G91R6/ggxaxbudIziF
8Wjvy8hWveBsFb6V33uyEVKukh4SEjZpKoGfHc30gaMa7vnS9HVTcVES9cfiLqhxScla2FisuhbN
3GWq5bwqqJh+kvrQfcJjoj8q97LjzAbd24yPEhkXJkATvZUPY02mBE6ozx4na0GGNQRY45it6acx
bkA4uAhWCQfkQegeGqj+z9Mid0OicnFpeo7fMcP1bdHRAeS5oPgS4nYYpImYEz/sylEUx3k5Ilaw
b88smnn77V8NUuA0oYga3NUFTqo77v/jp3/1D3LOif9vj7ihZnFZHr9SJgetRUJzXJFA68gUX/RF
5q9/P6LQbQaSUiWxppaGK5YILS1inYjr8IuRq9IQXqjN33baBOH1XELyhL0ZXu2znfK5McyY/iQU
cfqjXHTESTrTTErnbN2af8x/PbagKAKH/7YM4VKpuhdVENW25ACeFuvmhwhPbpLCl65OIicWB9+1
xk0PaBsXB+kcCws2pzH8JFD1Zs9etQdN4Q/DNbZwCLRYJk0ozMCRH3Q1pD6n+DWJWUdEUyWknS0N
I0ndoVe/G1WUTczAKm5Bup+VuHSq9EWwdXcbahfbbTN7AELtFhUnOuZLTJ5XbYOR4p9m6OE3K7qB
ZthGtg+TV6qnKyFVTOCEyuCcddiVUF6uP3RvzzfukVza3FctEWQAhWopAR5Dezg0ysnB63+OOrjI
QjlY3tC9CV2utVdBec6zELJ0UiCbpnfnK+z7KUI6vhsIsAFi2/KDWoqMe6fbNpY+PeNRyGwtKfuk
AKIIvvlMyPj1J/JGgAHF3qXKQtk5ZNcR/mFLhpim2YyJ5BNKhats6kvxlIE4VikOx3h0mhjteii9
aGlE5XGJMJUPHWbXRkScABgUY5ba9y+ZaeAeRSpwz4NN3ntb3Oqz9ISuzrxRtpAd6y7+eDruPa7q
bmteWZtvBFKJpQyWAVHsR4GRIJbEFDlhG25kcN4JUXtzvGgZjTFfwEAZlt1/7bX765dcP2aywuQv
Da8KnMOuIitq7MUZ5OBi4xgOEHgE3sTbDdoUIzXleTcqtPFoE6Ffb0StTgoqMASAwBr9Lk/67eR9
NwtZNUW8dmohjYZakrO15e120jjLBdzPVQBAx2usYvP/fgQCiXMp6VIl3NRsbOWvr74YoitezFqD
Ke4p/PRyj4Gvj3uuZPIDF+dYCzIpcC+KipvogGQzHY3FCSyA3uabY2e1KDFz4oaN71R5aD2gQ8pF
FADSWckQJQ+YxM+GV68WnSqArz9OOdN9MSjqrRd3bm1vDCYGuTlu1xIVi5G3MYdI+hrp1sM4B04F
YlNsL30hTsB7QdeVNvK5cmD6BG/UtmT15BQUDc5K8lCfVof1vqDHT/6RINBeD3ankltm6nlYtc47
9f/GK5gTZ5Ty+CsWVly4U1d6ocxLoeRcezG6wAbGefMSOaMQU/RfcagZ3QBQMKOck43qLSqNZNdr
Hhq6mVtPfd/cEbER42USv4+fvozwruK7i/z9m9ejHr9W9QxOP4YiV2WkMR6cyO6/Z75cYQarokOA
vQe+XmjEBhSnKRVNX7ZMdY9vTn6fgFeLH3WWFlSFwX11hPaePjXyPrA7UfGzMiXxUN46lM8Qq5DV
PZ/cS6t+q9bxPr4HJ4JN4bAhT1XQgu9eddCJPARsFIm2W5KepJFdYNiyB/XD2GCS+ua10bQeQaPl
AIDZMmE7H5xTUaWk1MxmSjqs51BhsKcvMQCIGh5xUAQwV3BKl55vAxgJOlAvKqqMdhY2oxrv2yeu
udd3P46L5I9FoehkWFx21oCjT3Dw1MbvLsAeF33okeXQXkL+Dw0ulmKAqHPfPUFlnBM+Px7FnTFf
6xCzILU+sgqqO2U38tq/JAxSC3YJ4ll3S+CJRhmgzFVc9FkIAmDCyDwaZLQFosLspT2eDrlhEniN
hFZh3BKPU7AFU11Dp7XyvrI7CyBaMCTcMYzabj42iKSh6XoAs3JtEcf9vKnLpC4Pc5C9nu0iRnTS
Fnefh3eEBTIpwz9ceVma6ikqoZhzvbM0XQxUd03YpKrdlGCafY1bxln89HCPSyO6C+vqX8m8Uwm+
wG9eC2UxfiivVugI5RK38XJqal1w3GTkxSm2H2mcPBlAiT7MPnqoq7I3m3xaymwGq6YeV9zf3m5R
bCJW6nRcgdK0qkXza+t5xdUIpjKZFggpxRh3cN1Lv52cnlwJh1jGKOSnBwP7tbXLsZmS7JjVW+F6
HRpOZbqe+tJ0JcrshFwNtXD3Ar3PjbmyVY8ZFrY27aZOTToxxcZA4ZeYmS6Ipuh9eMWKioP5SmAP
NTFk/buz0B95HwQnPFgSEIJEJ0kqk0u8Y22STgTAvRhcLA9orRogoT4E4CwQuYMI6FAbGPRXJJtT
NeJz59v/OoieHI88Reflc3i+Ak2oprlQcpRvRmTV7EEMzwEXvndFmLTXdh2je6BjxxxeeqQd4By8
iYP1Hp+XxICYL/xq/RUb9ip+WJS/Z34U37TaPzQSJVOz9tGH25XRUglGmfsKAyAwOaueHBKuV101
9TSGmvnZg9GR8dBci6FPY+QrdXA4uX8peDb2Vwi+zoWyQSWDOHIJLc70P9rFbZUyzasq+q1G7Ouq
6vRpA32VrZOozz2uW0Pi1UudFxUJW3yxZREFMGLu5ggTTMrMKODyefXiZRroTfjY37cbJn30tsoq
R2a0Hl9iS3Tv9EPpDDWcAFDK0W1AVb9GqU2Knl6nszhwt6taF+GC77ZJdqsdp3X0I835j/ZxJCbh
Lvdt+BHE5ieepQpGdQ4UZyaxiGBa6oQe+LZVVpHIS1PwK557yRuLUq7qRsZHUycTYL4PkW52EGRw
RAgev/fcCfHFoQbVwf7kOJDfHSo3kgtEJgIw0YPlyeOUnPaVxDWOLVt83ZAN/LQaYqhxcr3q6AyI
ntkzQ7ODJAo0WG39p0M8yAvz7XZOf3bsIK4CwQ6d8t9a/xMpDq0+UcMnskh6D3J+8MFSImFnd2DS
Z0XWuLUClze7vuKXYVlBfwUeaT9i+R3ql1cgnY0dW3cDcgnVjH1ZiKSeqUFGmHxPIV30Cy3MvUy9
UrRAgVBCEaY+PJAGRNr8Ya1JT+eB6M4BpqC+YsxGTVDjoFdy+Eu8KHV4U87ULnHfDISNMpqk9EfK
7/RAiIuhVCGCn15f4g0Kl83Ca4YgqW0XGE+l560+XyTsxVAV6YYVdAa9MqB8HVxbaG5v7UKxr9IW
xtbR6r+9X2eNugeMivgRhr5M8PEKnywgP8fw0lXRVU6osI2SEuTEMT+Qx27mPDaewnxkPYk17cgk
/WG1ojKginmsE+bf9xuRjApOarJa0F2hM4F8vAId/E6Chz8IeR+ZCIMNYdC/FX9MS6sljnM6j9LF
L96UFxzwGG4UKHW/CmHClTamw4TucaFn9vUyXxwlIdK16+DDmBTcAzRzpmFvNdQqCF+CPC4pCYjm
vMTsKqrNCZMEYEOlEplINlqHMxl7QA467B86rzRuVCQeokcSkL/3sU7rri3xRVz4k79sULC40K1e
XvXtcHnIxJnOF0h3QuxN6uvTcN1fR3dPjwxArn/ZRzmmZFldWyCc3rmSCxVM2veorvFUJtvT39oV
C60o3V0a6nL+jTfI9tl9POppM2wUNuyNa5lQ+IhueY2HE5p0KUVpuj5597/1nxO8T4mmB7Yg4aOs
4C1Qwk8eTmm7XZVxO2nNDmCelWL9FcwqBZsqv88fDw/GRW0VLoB2BSarVOt/bzLAXT4gTwh8RlTw
FoQ2SBDcA6jnEgFaVf9CcG3lfUJvLrvDKzSgedZzdjbA7uBye0SGYnymJTFrov/QAClJPk5qRoOr
//tuvdL6N3r/b3V5eIwJLz3xo/AsgwnpNtYeiIRN+MsvzR+zQ9v6hdNWPS0L64DMm2J+60GuH4lw
VXRSFQsIoOjr8SFlPHIf3iP/5C1h6nmEXL6So4DeZfi9ovZMOwP0BlsSjWrwU3JmqGaOW7SZPekB
OSe22+D+XIspd/tmW3nocKEZrPZjZGwaXLXrhnrj+PAbDSbEjLwTRXnGbXhgf8xjlWjfoLH0yY4W
0WGR55wT24XRER5IaLjH4hjGIvPBeBqi3xxJYyT/uoTMo2LHBhlaqgoXNOhsnXxlwinF4UvdFv8k
FMdN4stipIjpe8uXH5KXf1BX/TX2Dw1ocXkizPqBqP78XgFh3Fw2bdJyZc6bP5dwkKg37TW0oDf4
Spmt/Nd7RmKmXAByWDHwhDUp8Wa22g4o91lNZb+Eh8A00zGmS8JGqaR06K8C0vuoRyVIJw2te1LR
aFi7p07e5UnNOdi8erQHeZOrksSkxH2RfaZQWe6f5cxSFJAitQg2Yo8hN8VZFpYSpGT60qPfI/UC
+llwe/TCHq2VMGFioMGQ9PhLUjI1J7a4Fpzv45LYdN8JreF0s72KXUdKXnLp24Ps1/Q80I6ufE82
OpIebHVblFMaS9XF59r3ncxcQ4IogRJbmhdTyONImPYWu/LtZqxzT9eeawRcksetYRpFD8OUp2Ci
u1gXbcpw7jHpLudcDMsm+9a6zYmCiNZxkBe3sHyeUz3VVbaT9rILJ+SqWby/3wNDg7nlvctkGvM6
KEBJQTHbMwj7uXW8u1FkeDMpCuW/ACqRGN93+duRWy5tZ7h2q3g4dEZItl0+2MzqdQi5Br5WnCYX
7Y9mQXR0EMdZh2XP9OPRTLL69CcpoEiToQBuYl/n8/NhZr0MGL7TxCqEH6XQekvq8+74kt6IWgyG
ZOKCVR1nHhp9tB6ZsBmBO2cIZ3T4eItRBXO12ykNDAqYu6v5IOXhkh1cKlx3FhLL9nRRseGaC1a+
Okc1kwAec0YO7WnqZ3HGEa8wPF7YddCSYcQ6qyMxWdmtZ1SKIAPr8wdrQ/KCPdovz1AJ8cou0JUW
FP9xVM5l9mcQq5ZqPwRRb8Ky13BQTpM1w2cSKihH54Z5hDuyDWBQ+HFT+LPCHS7XHqmqckCFxwxY
nWYNnx7bFnmAlzx5CT1BcUDO5ofb7xYof9PMVCAER0h10TXs0DjOI3grKyBnkR0Tm4pLCeFUGveU
pWV4wy8m88+tRDlfC14vo7s9kolYXoGS4khDYtf9r7dOgDyI5jQkqn7XdGvKighm3IbsZFAawF4n
BdbzxQjyu6GeUkhJdUF7g5w6nrixXcfgLBXMWopmDVp/FnfukUg2tBAjF3dU9W7xd2wCOlXreRJQ
WBcXWmdbZoccM2Jm+UOh5numqGfWRfaIN/oVeYFilx69VJx9BI+/oxEZZ0poKGL5PgwGG6owpZUX
vhGWCSAU5SyJgcpmBSNDbVGudW508HDGF13zyYQAV2Usic0yJO7x7UIvqHB4qxvyjp2STNrE9F9O
otS3pjWE/dnHKK+piBpWASpvYmdGGLyU4BzeL8Lk0hbn8TxUWTMwH1UJe8OgXpatcu1jbLwp8UrB
z16TDatZhCu6MLzPQjJzBoLczI6c74uqrgWmlairMcJ6wBsIOT0YbpqHot/lk+Melj98n/gbgrb9
gTOt6YbeOqMCXHnWnxOOPzDtDc541FfYJUSnjYtCRJxmTQ4o24q79+Wr81Lx2yKakxxVjJICFSzY
slWgKgNNpYliFyHYLMJpgg/UbPYhLrldDW6DEZcBf4U+6bhCNtkdp2eQvCNVSNysMFv5ZvpGPYS4
soTdz+XNM0Y7gdeDeQubSjtONy82Lu+yw+dFBhY6+X0MpWvrdoy/8KCGWiq3bO7nf8JgFob5d/O+
qDEwLJYzPKeUh9gsjhxzx7f6AClmxWXaXXASbf+p2zy9QskGBfzB9G7UGcVnjZhz5ZYpkEq0x72b
XnLSgD+qgohGCuGoocvLIzX2XJNMAknOsB81Q5FQejkqVk0vNT0Pc8Vlu3X6PIkWzWo6nedf6IEO
QheW3KiG/EnB0N02bDxFQvvVDRk6GRqaTNWeHJbVSeXSKChXTQZFNN6FHyP0DwNJ5GVqnqspZbN4
LZH21LuWe6y+MtL48Ocy/69V8uLhrYHReFinNTc79p5Groarf6eWOXMgfKjt6/DH6kNTND0BOuab
rWTME+LQJk687DfNcMXWzAVBvo7M1Hgtk9CaVROwU0qFpk1lLe8iKxNdii1LFg5TSmBCTkr6ggLy
8RsBtXjiJWYmtEqoWNm3b++q+eyYfuWPDJh3r9qakOCXm6qBXCKQqXe0Cf7/AH78tbuBQT3/x32p
iQh9mPjto/o4JsWx2C1Lxv3J6WnoYdD1uSWsUmq10YMcGH/RqCJQ4tFABBPOQnP+doBprXO0vvgJ
MaOgAO+0rVgZU7IqBQaPzAq0FvYYG+RyISMvZP3FDjBSNtuDdHgVDO4sR4pFrA8U8S3+w5vmBNEO
z4bNLq/W9c6ySll0G6Vb7C6OXdG9Q05vUC7vp0/H1FGcjTM4SKGkwQZGe8G1CB+Gj/q5yCuogS/z
hC5SWSk7OchwCohSCWLTTsjghpxaw48rfsrhEfHLQDTTABTc+eoCBU5lmzM1XupmLhi2KRV7VBVm
kOOeVkDRV9kEZkAe2kTLv+A/Uq0lgAY3YJH9+ImaPdrYmoLcTmyHK33RD+BGSuqkCQHkmlcddNJk
mfc7lj8XOlU9Va5FJrxqcXoFDTGDC8OiuSnoj2eB/+f8InHIYfzkkZGXHYQpKlkAu6klvkP6oPY7
ghT+QvwDe/VCepIMfiqPF3QcWmsqPIBJFLBhX88q+ebs9i1SchFRSlFonGvze3QAo6hqicX6vlOr
qDagNNipZctt1OaHGG3/NZCavl1lfOyEEHTTXqWuQJAUs0dvfQaGVIZ4kvI57MWM8ijfHpyaqZ2E
mG3SwNhWHXbuAcYk2hKTOKqnZKYOpeGJtPT2dqjp0437IazCQedgR8EnTk45xZAt5Lh4NGhwxVhv
V4h8ujBSjlZrPTLZ3QUjhXp55DTqSYnn+JDWHO+LCySF4w45U8rcqZxVJy2FFPKaUyaX7K1oEsBW
zdZepPXrPcvQYdRmoZtd+0Ki+gama83k4Z3KVX8ReucPXYkIgYOslOeiGSrfxk0jzXEJmO7PERz0
u2uzJL80i7asBaHFJnq2e22M6cmDqbPwCaOluhZG30+ltKrU6oHMsWM+o8qNqTjqa3PzIns/iHGx
5SCovlDMPU0CLYOX66+Trii2YRb90cyd4tCWore1LpNN3kqWzLSz/w9n/Ln//9KtMMOX24JDCIv2
emqlxbUjWEbhlygfXgGfE5Or7ZDwbm6k6kUHSJxA5ZR1WPyWnw4h0SOvrHZLSFdggmbxIlHw8Gei
Ezy31xJIQFr8qIEZ3TYaomzaIPdpF/KzFGSKrgf/KlyGq1VSif89AM2DRGWmZGzJVbfd8LIGMfc1
Vv6YwBwXuTFIiqqYg8PvASSoGEU9j4rc3siAai5pNTNp5hHQPUK3TwiEJuovlwwQiTWB3V2K8Vf6
zbYOA0qgzRK0HyQ8rvuI66RxSEW8MkwNP2VlkIVH6ZssM89e8/+Wwx1rXNQsA88kW5dvl3MmVjUE
GTOzZOeNccqmOJDM40A7iyhIF+ZhJ3DVoBrcZ9VUmlAqunJo/i6ZsU+zd6IfhpdjlE+dfF3Om9pz
GDgX9S4klovcdnRSt/1dg6Uqn5sxf4FZsidq5KGsJCqjyBqHh1sX8bc2pi+46M4cZO0fi1UW2uZQ
HOyxadN2FoRVlWY0m8lHgGw+PxzKVvl/KxjcEHugL4tRkLCInLhLDRgNYXOf7/JWloh0u757RRdu
HTbzBZWRsOu+qAA8I1ZErjjkZRlnTrZBdi+bf5euQ5eEDdqgzBccpWfjcikS5RfySCFy0o/BJa5P
Z6UaE82s1uazMJdRHTEgzxju/xq6EJA9Zwh3Tl/fIHNEd0toHxhUEYeImw8U+qY4U03qFQSwRYZB
n+t3j7Jb4pLG8Ip5uJJp255N5mP39ewEjMWNBzYrH5W7GT66pSLVVtbYW7qSxEIybVfdIfB59yMt
t9GQOhDUrfler7CK3NxeTdVWc9wWmJN2JY1oiGvyodh7Ee/ff1VlD2vYPEJAturyFjOvjXiLjex0
qLanqYns8u32Bk7dsaf7MLB3jJUlIQMmC2IC+7ARh9NaW4Wm9V60GzqZRAa1NFasIelIOCd908Jv
2Z9kt3G0Erp3pQ2pdkRNaRrAcO4oFbDRtU2hQ58vqMV1KJAfI+tD9iN7cCKZ8bZ36M2BIixhWy/q
oOJC0S5odNwTtbB95IhEWb2iWd/oVymP0NWZWkNr7HT4VC/RY/a2ShGQ0MaSXW3AuBKguKtON1gb
hsJmFfDgBABlpwFyXDYJebwusliy1aSN1/udNPdA7e6zUv77A/2K4DaqEu27m5mTJGXwaHFgM/XU
XJOex+itLLeQAoJ0McZAWg1Y1dO48zjWbM4OeUiRiXXNikns+xfRXBl5SesRRR0UNGfocVE/whoP
dY9y3/LtQqOTaMbpijKaPUB6B+ou5LNk2o71e+TTu1c4WTsQvyJGh9vPzHXC2fo6XzF8kIu2ditv
SXk5vCFuIi7OhiMKH74zXEqqEZMfgi55YLv66wcVxfdwgzfvshiZSC+ZdB4AsG0ZC7d9HVbcwK+V
P87M6SxVn5cdkNwRtVFtuObIxKR3fklPCI/w2AYqLChdB1lCn1pi0HRh6e8PFV59o6UsFiReI/aG
AvbBlMio2C54cRxlFPhsO/l7PURY0/uHs4AM0fxSU7EtAt9bseSr8rsZAoeSwyJTxPDG14QHjMqv
WqOyCtxjlkHZv1rP6AuH0W05BxLZxz7AlzpZd52ipBFQ+NZ0gcYTu5Qk6Q06mtYhg6qnqliLBAPD
vJHQktiq38a7bsAt33G6k9v8QT4+pf/duVxkLi0W7c4VH0FBjGOR34s6Keiv7zKZ5nYIOy7D5q3T
m+TftSAzIjDHkMjvt7Jy4ZBzBMSmxvr7hLTzgR01Eyne1JKf5Q/oU/t8T0I4Hl3ziNPZNtrXz/xu
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity uartFiFo is
port(
  Data :  in std_logic_vector(7 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(7 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end uartFiFo;
architecture beh of uartFiFo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~fifo_sc_hs.uartFiFo\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(7 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(7 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.uartFiFo\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(7 downto 0) => Data(7 downto 0),
  Empty => NN,
  Full => Full,
  Q(7 downto 0) => Q(7 downto 0));
  Empty <= NN;
end beh;

--
--Written by GowinSynthesis
--Tool Version "V1.9.9"
--Mon Feb 12 13:36:18 2024

--Source file index table:
--file0 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_HS/data/fifo_hs.v"
--file1 "\F:/Gowin/Gowin_V1.9.9_x64/IDE/ipcore/FIFO_HS/data/fifo_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
UMlZN96vbvedkvzqbMh0cOLvum5Z/GkNrhK8a7XASrzq23Mj4NWutdHv43PgvqmN4yxJ+j5r+VmL
nT1sMnScZmwot/V7hDx5xnwKz9duwk/WCjSftb82DyLcY/JtunJ/3tYk0iLQYTON0De5qqKs2N1P
mPL/tr4DOMfSasPrBMC2DQBQx6ei8Kt5mYue0sECgSbaWlTHK4NNIQLUlniIeV93bHJhHU9eo6Ky
Evm3KyjRZ0OpIiNmScend/Hn3WnouVlpFnTBi5BCKV7CLIGN6cR+TDcLGT/qP4RIOwtWALGuTfM6
F0zwkFPcznCUsrzRKhzMDIBwnPpZNsCRybwUUQ==

`protect encoding=(enctype="base64", line_length=76, bytes=30768)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
fRFCGMnMcK7lHNDbtej+26JtHJvE7aaJmZ534O2ILzAwww5ql0mXbpY9pQFcrqimKgQDn1DlgV3t
D+nNTg4hfDLTu5CvKw4kK9/1B20vsW9SU6LGQWXiQCoDWikE6hgNLivsgcf0Fh+g+6M9LTzvTn9v
cqQAj9qh9AYGJWMpHu4XtHoBog2A2qE0ALPxta9xsEGtQk46BbRR+fHNqcdMdzWisZv06ynclG93
3VK3LN/0a6nvWoxqBkgVcqHQhDT3FoKExV/YWpoEKxJii8jrDDHZBMkxLaiBwfU75a5p1A1KN6MF
4vcQV+Ly/KgqLNKsmQk8pZ/Q+VxKiRJruj0Wsyd4fx7cB6SiyO3k33bQTFBRjaX9XZw5xwR0ryVh
GH3HD0G7omR6tC920ehlliy82EDYd8GDQL9YrViS0mzlIOL02CxCT4CBuTs95+P9piEblixF59Fm
Z31aj3FRWkukZ5g+WB7XevgrHulXtZYtJX50ARRESe5USQ/DfnZUR/RKgD1Ajt9ic/SxCce/9u1e
EJcQhf5rDvFnD73+WCdHgbpHFGwASMoHLV0DSKgDS3FSS7GWhJoOmEuq/C2tD0IujbWoE1BSR5Tv
kafSo5MTF83k3hPAdq/JtQH2KjhDXfLMP7R7CN+LUID+64VA6aYeWt5fK/z9cUmT+eDJ59v+53Bz
RqXOM6lfxoXNf496UrNb+bdJDPGtrtOBTj1CgMsHEGnMrPbKvpf4goTxvMH+fZM4KKv1Vzv13JNw
5HeVSRZku1mheyqOHq82LpFn4RvjOw342+zvtQMgV8lVDIsRvoeFehGo0iD5SJk1ZTXFjIiP+5PC
cLlUdXfx4cUt1ngB8rhPZRyP0fFP1nuw0EL/VqfnW4WKtl6dTyIYPUiD4+KKf9Qby4DkoZwcfA/T
ILTWu0yBQ1u9M6figbl5k8qWeLxCQyTTwhDAPXFl/WBWM2ap898MpRXceP/8BKv2XAyeDcmfNF8Z
0d7IF6yJd41JF5sdCPaMSbCBGo9/8VonjFYCOG5ttbo2/hn6pKNMuxUtyDda7IA+9/E9oAM0V6Ca
HzLoG3ulYoo8JeMnDMyrD89mePupxW/VDJnd4iwA8bUjVlOvsXFKWLXY0fY13YFVZkZlnPMeFVzb
1emP+5lod7LPqxzOTSZwwW60vm2/cFe00NJE39l7E2g6RjmFOsAIrvNQcPQvgbIH9GtLaKizdtfg
Ev5bzFlQxYUtEW+Rla35rcSaEtDVdJ2lWypqWYu0juk//hTcr/rjiS4JKZqsQmefGqhNnIOCAbU+
tTc40A8/ogLofILJHjjuMNfQuWWsWWQgcDNwZeZXsM+aX/yFFIqEm4Ca5gprmUAftBcFWV9Zk9mg
tvT7LbEckNd9ZTFYgxOEpAwAF/lAIu9+/bAGFRY6xggQIpi0hPWiJD+23zM/pJDajRV80MEl9StH
Fb7z8X/d825S+JqrEZZEA23AOyX1t0/GgNazku7qM6jUYgG4j6fWbEVA3rL3bxTgFpVmwwk5VcAf
cVNQPVbOuFv7KzYOy2GZGUdTsjUS2lsXrcBo7C5qwLMSEV0eQEIwdfrwsjxSX2qwR+vHWwNRlCmn
0+t8tNxciGgFC5PP4IXKXsNVSHFFRhEHT/gZQtMA+J0rJc6qvtdCsnE4A1XeDaGK++WVvYiBywEn
WIPRa2w5cNoRRTFreJhowCL9FN32bOayBwi7lFw95iGZSl5aMcnkLqStT1V0nvWn1t+i7rQcYDIg
9+vjYpOfMrnCnQ8wZXkrsIYGYniDKgZgC/xZ2HKDLdc5BRRoY4TT8Ma7Lur5uwLAW6Z+W685tpcF
9D8bV3KGWXgszD485gTrWxynffvphGB9zK5trFV8H9if9+dgC9AS1nOss7BjOrlZdGSDDBEQ4w08
3lvKNNA5gVQgVob1DKZBfVRn4FRJQUODFJaAFt6mQD2Q7VR61XVXDAdjLDTzpziXebcm57iK0P1T
ThNPWzWrCO39oS119vUQyPYRPk+ZQdGfUb9DWNzbfp3XPZYMHFW+XMcSeMVmN8bZzN15d3zC40wy
caUeyUv5m1agLolJhWjHN2OtmgfgTUlwaxeZ0b1/a3nAMV0NfFhPb5yAYiKxUK737ik1qtM8DalO
X7a/jcPbbeHOCEBc/T0QoUW4q8zLaOVWinF/9JspEE0GDT79MZavyt+xQayfWTN0T0R3Ln6zsGzY
RCqjpL5251r3vzJIzuOtqgGVTOy/pj/Qz16UmVeAOMiUTkI0STNYFtjz7aCN1zn1rgFFsvnnFWbC
QdfU3mKo/MgBXuUF6ZB9gMYDKE4+KZOMt1b01uzuwf7wXcd/5jjSsVCC62uZoopLJIqZTcmUKdgW
Isq2ZLqpICWKhBKccxqFZ/FYmcx3lDqDuBqeH9OjwfEOJJd2YxrXAPT8uzjmCCfOul3sCF+4ben3
dXjC0Ozi66G5aLOeCuKxU/qjzy0pM1L0c9GPXQQbQPrg7uqoPyF3+FUmg7LcOKq0yYT73FYjQCda
efb2duCqpREZi7D9XWlsGasLaMv3I0scBECTcSPFeuPhwVhzDIzQxXkjx+ra+O1yOoL+tbbvUvTS
Sjqer1jXq3r0hchNvaEv2w43VIYMnC47jqeZ1Ks18uscVoWrZAgq2rTWgfJBvdSpY0eRxeZGV7Ta
V2E1JkiqWmh4YctMqE/tojMaPAlGONgI/lppoKul+ZWY2GdxeL8o78eeWXu5nOPiKSKj//ToHSQt
xsPHaJiViBBqD0FhaGQjJDdDdmMZdF7gWTtT1cLrMVr3JsK8AAfWG3cJLFrzjJ/BqgAcl7d3aTy7
/u+sS8B61DtYcz60pz37hTGnx47Sfm6v5S876tMcPzFyv34qXaQAubvBEOIR4r72sUm4dkG5bmnt
l8PwEZVPBueTLMiZgiABx9G9M4P22rlhUKBL3JIUZimGOiBJSPE+N2KhV1HzTfkfg44gRMgXOicD
03OKLtmWhN7bDF9WkZXBUjHw5VfPjzE/oErGOonGQGhq3eYoYTf/ZJPEz3Z2oJL7AqIUer2t8PyK
s7+i2dfvpc3TjpC5AMOn9af7qGezm2Nq4fGDANIhwJ9b9nsonaFJz0o6zqjebTb2kYjtHrL5zyqU
SM3bXkK6hiynuuxj8uc/4YafioIfEFhwGwHXzAhCxoF0FC9Asy9TboCFCl37Mmc7SPsqpZgQFwg4
bbqxwPPqg8o7lGWU5fcMX0xRns7kTUyjbg7QwauZwYipF/AdI9HMOAe5pnvtUjglg/byTNGlErcO
+V+JK9mELl9PTB9Ra6mmurb/JgIM1LkLGgzxikcNkeT1uI0YI2kAoT+rNfkiP3vOS7rYtcodl7/9
P251DCAAqgrGmItrV2G+YbvKpYiOd0Yllurs/yXIE2Wg9jInJL3Jfkp+gT72hLoMzfr3yf4LctAP
5Wu5CtmJfVAqKNQpKSik7Pqeev0weFYY8qks5fQlo9g7Sg7NglyAyEqfcL97r1j+t1GwXdHq5fha
6ibZ9sA6K+JGr+U2i8DBssgYGxSCxGqHAFwXipFfHrKxsvGuPt0ze2b0IVghrOY6D5v+TzedlxR8
Ts+frA0rOKWAU1Nh24vK/KmIOPZ5+awSg1vJ52oZ9jW/6mlYVGndhCwXwI4v0t0m/jKA4a7DOq3Y
wkECksVIm7BSYMqwFU7pNq3IjpnVtATqGT2nkMbtad2ijWHTAREdY2LZ9ou3etTo4Wqr1XH00Zff
TfzJucxFPNXAeqtpyjLj60Q4tU4I8ZwSG+It/nkYtaXGrVwv986FQ1lyGJxFKpGOdNRUe1HDHEYE
C7Va9gl3Zm3mUbNhM2KnJ9eQSrWGM3vHXj9S4OOQUxd5xEgpsPx15V5LUlpE/e8oJXoS3OOaQM3l
rVPrsmFjb/XgsQf/CvW8GlNQ8Jv5q91CMcFKE9P2bWrvAg7vV8of3/3m3Q0O5mhvz50PJt/N5Qow
BrNrPzJFNz60EcYFGYOqF5sUAm2YMPE5+CeojUzv1KxXBjPFEOID42dT3k93oN24EXG+Z6CwUi5E
yCrt+Wl4WuCoIhZIE4sEe2CtcaiHlHUek6MpxqpC76KnD0zDKhNtMYeDpPymyz7hQpbDpHz40Yo6
7044PUAGiOnOndU7hM2vE1D2kM/F8BZUWAEAYvl1POYwNVd9UOhcTdToQPVwzX7/k98re9L+XCVr
d16lREA3y4IV21W/DcKbC5K+88ZeoVunF/zhC5uqmmzmmyITXuV3bk5EbojlXeu6FA16YNLFjLHI
LACjZ3L2roEQWSOTe3sKCM4wSYGPpztMeJoZsAB3SeWR4iWp5lJskRcNev0G45F1hhAu8EgqGJOT
3sP3oF7woGSpAIWVO5R/BLT4cwuqUzQBukxYh+P5Bg1Aw/aTRzcc8O0knZSHhHTaKAVx/Ua09Eoc
w+796QY5fTNA2YqWhHmHUvWvYAI55tBlRrBQzZzPT1OClZ8Iqylpdno856vRiHFdw3D0DHeE2P5V
X9ILYMytv3SDDEl4d8BhIYVXgmAuBM3X9h4emOLse6+FYGTQmfDnwuGkC0Vmgr+lLudjegy/58/Z
cO8QioRctBgSSHawAGqknx05Wxyg5jrfwrloiONNd3/lIYYP+KhrB3N+2bOmXctBnI1IkKhCg3qn
dC0lC/O6a0iyvReDRp81fNijhBR4nL8QzYkcuuK2Lfb3wZOhUm06K+navN438xzn0AYHbRzJU++x
LzNX4R5wMqFQ9fw46Wlc7i6QcFyOC4FhtJFJULJ09E18yEID4JrmKhBAtMMNhhXP2WzHJBuq/5BV
+cx/NuyLZGiEexPZNLj83NT4cV+JP1gSEYeGP0GhomtVDFnau9izLn3+4KiTUIaZqoj8Y+wkGSSJ
NPgrcawGkmkFndzSpkcRiqmpgfLuO64z1HSoWQ14NE8K2JJRb7Kgmch+CAYWlLsA0PxgDaU5iQHX
NncY+LTofgej6ldqOpgfRXsvPAoysAPLXjETe3BONHE5J6uVn7bYwQua9kLi+2Wt6YcFWainS7ID
0A8hI+4AMq6qYCkDabxbmIub2WBTXNLUERskg5O7DpeGPj6aHbHQGGHYrU4yKOJ1CZPM+hwlJsjW
QfsXVybb4/UqCLWfFD54dOl6xgzDJT2cYvy48qMMsEEl4NbkxhwscQ1bTBCm4mLgADsGjY1s89hK
ETBDU3hyev4Tkyrw8/KZKXXq3JAaPyZf8NaAUVa98sAQnNP00TshBm+AvwECAp2HdiASFigJlGnc
EhjuyqiBnfset+oR5+A9AsX5Zx906czdrtkReqKLBjlCWgOdUargj/BXxYKvOegVkGxQh4CqBSkP
aeVfBaxdLUAsFYtzFLk/1gKRnJ4XjgeBlJMkzAKpTmoaMq4tKwf8ueSmiiAS3bjWR0Hufq35FY0H
y+LJ92d9cvgrFH6i5hYZTX3xkks16ah3pREQzoJNF7FMPrQ718rAmu+/nqCZOWJRsxEGhGkqZxv2
iww+9uBbEz+WxxFdfuwnw3iYeYSibYMlBRSu64H1i2JFNg4plXr3sy3Lj7gPAIO5MmmcFiPHmG3F
nuJWdqkV9aA+o812EYPCnMTjsna/pJxoETrn2FYhFIsfBO6SjhNRBQ26amKPBPgdZfmGUQx2yKKQ
pXZRwFy0XSWaqsY7UmU3AvZI2lEVEWxEquTdjjhRiYeeAo/sBq91EhSoHWxX+O0BSpHhcIvzrfH7
y2Oid0Dk5xUUBApSWtRTkkt3RWhRopiNTegwOBYPvehkKQoOOlimr88x2exZnmnzjb1YpRIfZFKk
0JhN+KM9twul1M3m6BJa4NKB2Ag3cnykiXECajFqUrNJDm4mobglSzoSTYsXIGyi+zNdudo8yfGX
Qn+MRK8jzXUKAmJJ3ZZSVfT/TLX91znWxqRm3WwhvyDkOVHu4ELrejoB4y0KeejLZFNB8CH/3XQU
VKGb2KhomQmUr93oJi04SawJQWpgnKAA0ZSDkivQ/TTfZPxJyOum73qYWTRpqzXiKPWAKZyvjxlL
FYkrCBtBzb1HFv2N5wpDBFm5zLfbFj+kham96OSYRkmmHYiS3uKibwPKVJCOVNRa27+fGdWEKpy0
EdrqSuoStVF5lOo81uyUcaZu2rM4AClx9br1z5tMz87qe+Y8A5dfoSYIvoIg05dSBP5QZOtX08XE
d33D78+CffvsTV3K9Him97ZfVOFtJgrR6Sc2y96TkfMyI79DFb4a3PK67kXfRFbNHXCCW7uHdsa2
cEeMhMnSKQvHwKM57ABEW2yDCOAu2EEJEDfBDt9OC7L0XD685GWpiK93y8wwNqa4f7YSMG6sGS0C
vNCTCfElFC4lLii6ngWEiWi5BKtKwfSMuNn8/672VMfb/f3+WZ+X7I8qFIjyGZh123hoKPTC4CQm
0cA1xZXpca16/djhri2d4nN4+KXSBu2+uGASQbUJpWUleP7/Wf2BySbZretoYzPoVqrieS9b0EX6
wp+z+VNYrljIbwegZoEyFr5f54/+RkhANkoZJ8tTG8zmZ7d4ObrAfU07Hlk6ef3H+vOTD2KE24bA
pxC4m5D9GGK1YaQEa3jL8T6PIKzMJfgNnmdXI+XYtC1umg5OLlTavn9Eh7zzm2Bym49EB9tJ0D7A
ZGfTXLcuE4xiWZyXDLGoxx4FWLzaZuK4H596AW1VifR5eRC1jsv+Ok9zS0ZeRKd0NAM+VnqRIWlk
AN2//hSMSgAu3t+ACyHiJ51uQ+BVpcjXbyPOl5lh+u60++5L9+Kp7XuuLlvFC6EJ64mjoxAyjn4/
TXHUvK1JX57drRsvK1ny/vC/wCHWlmeQaYUAMRWWxf5IzTnNWH8PpH+Lu9+tX0rOI5ovb6kST991
M7z8wXcQLvwVMsS44NHjxSqtQSpV99IvupbD+DXUzysN+Ed5QEqUGiS0RbAkxrWtbBbHe6vBirMd
uE4J/8o9oGDWfsrGc7j89zOx9uCejHEzKk4vcdLzuE6iCRZxn9z3SBSNC7rZIyoucnWj3Ay/7oOZ
WJLvFqtZX852GJPNnJUfabAloCgFW2oHGOqTvKwDPqmBlvQdvzo2MajUsjve9VqxQRoSje9Smzsa
JClnL53j28uyp4lc3RHsUeHoO1sGeF4ACBG/+8h2gVLmA/7p4DVEXnrnxOso1LD+fB6ajwl5Bu7n
mQJAfXypLwxUkg3ldLmiGv4IPHt/VEnPkbQdAjRJC1Ts2hKLQbTjbmpHBQMgxhHWfpq7zYcIAZnx
mJahFvM0ik84qnHD9CVQYDzyG6i1/Kao5LkHpQZLPLZvl3n3+huHaLHKgAQ9wzxcJYAN0vMlsDP1
rSnVXjyQildz5BecEYmgTof2eB8OiIHC0j1mMCHOy4/nd7zr6tD9NJgVxB3fZlp69w8jQqPvI1l/
5vTwYLiXpCHaCDrDfXweE5oIJWp1RCyr6+Dq+PTM2khmwAfd1H5yzbBcAFR1EVNbMsw3cs0EhDNr
iRk5sbiztUWfE+7/eOW6se3AXx3TuiW42QEOgiAiwwvadNbYcpJay3ACaQHGeKt0V0NJAVTMnTQO
ss99ng6aHcAVtL8SslDFEfrcr/PCmwYn9HMTEUiPac41lKxicuYjEHkVgRClNrb4GXJE+wQau+wk
DxUMx/Tgzn7+9oQnl4MEvGeRcb37iVyxZlwuFX/4DcPqc8XnyWDeJCHpl3m4Z8plwWh5OuKO3YzL
A0cpXyphWvgE4EKhKqMH57EFNP4mEwKk0gAD9c6LxRTIecjzWUElwfoZGIkIS8NfvCyIrZu6uMOi
rWTocU91yzkYSf8p8KlUCxPfhmrW09Mx7ms21uENjLcOU8BJX4Co8MEGvECbg4iE6KWdI36h9A0b
nj9uGe9e5EPs2GvRgou9fE5XHp7FwXYWHaGS54schg4+HiX99qNRJJD0IjKle07RYCdjweh0UB7o
QM8D3SiWU2Sucnei/QaU1xfT5tgN2kqwUvof/ldfTma8+8PmIytPTgBncEVzaE+jsYbQbtBEf2oo
VF+7E1dOEmnAoFWIyLN+tlD2ZLiOtnc55vPpIRnwYcLRvpfCYFhWceis6rYoiolIJemYSBWn0Pq1
QsmWugLRL10I1yiwy1F5HU54vjpckqcAaL3XSJCk6/6pYNjGzI6RiKrQRZQZcyUiUYPpDQvLBnRI
5WPH5wWFdXdE5rnEB7W5/3prdOVJDmaDz8Tofv/6T3tlf8hsCT9gBFms1fBJp+lazVcfh9UWOZJR
zlddE3M2diXrx4xh9dg1XPecgfJVakz4lTn+LIu94XFRsLXM5BBqY8rEsmO1yFA/GwMpoyYFUsdQ
xz3uWq/kEK1esgSx2ZtFYQYy2bMLJV3We15Org47u6oT6iuRgfuPxpkUvwJ4M2e9vMVuBADUdnSg
+xBNGsonSIymnWfzmeOxkUAm1NmStLp0io9OWNj8gZInTPs8OaKnAVmPSf69Dn42YbcwujLJ8pLl
QjZKRKZkqP3xxfz+CMZNWlS9p6fU1Gq3J8HPJEyj9KOMV+NVVVygnY7xu6zkYo9fjtJxkOOhaUZt
MK/K3EIKjF1wPE1jpTaJjxUX3bbe9JiCsZ+OaaDLIaqrQALwtqVfUPjrOKJ/vRv4sCNghq1FzxA2
9MHzxiwjUJU6bighBkhyW6H5RvCi5trkdeG9nItuvXugtJ/1qT8YIBqjGgm4E07bNeetyDdJO8Pc
DuNm6NErFyeAXgZi+gJNAGe52P956bSNT07kExBaf6Iv28CEsk7R3SLumwXS8+pxkaOrwXKjDcSB
6fZ+HXOYRdANNN51MQYe9DydruNHMIm6cZ/hYDPrFIUUeP/3+Cg5aeGoSUXCk9dFwi25UflYDRHD
fuUs5d1aaU9IOrUtIZsmKT+qb7wmqsQoHemKWxAeRdXpxujoYFnTtllxaVUeCZ5Kzhueo//4fzPb
39Vh14WVAcjViapZ+HBOCUkR+HS+Do4y37maz7oJtNZQ4F8i15eJerm8oHhV+puYGU37w5SWOIb7
GkMLsmTTWAAyGgIYvz7qM8S1gqMB3boCOShi4P6YuqzZf3RTJaYs0pRHygxHtLyKE2+lz/mmP0bR
kBFvDKoFVq8cjTbdtBz0+JFT7PIGLkAs6g2u2AYRl0JSEbH+q2F79IWlAdw6EjubaciG9n6ozVDH
k9BzwAPZ43NyUBUNPXjfwSLLd60ilAJ4nGG+5GKIMfyBgjXPgt4w5+9uogFlWxvJveKWoeJJ4Hk7
+D63pZL3z0gvOkLfV/5ZQ0lwYi1VR7sU6obqs+1T4b7e4CP9VyFtTHT5otx3AM4f4A81IXUZfRJa
kg1+w5JqMysk32JQsgjFKku0MLOeyr7P/sxHZJydDvXwt05/xgUzFS0kzAMKgxGOPZDWOHhHJ7Zt
53S/OjZvdD/dzTwm5m5r1kmly5mrAmhAer1TiteWpzwOyDzfHT5nxLtc6yn7drVGxbuT/Cniz6AO
WkB50tv9dccAvFt+uMT+eE37xyI4KzUpLlx6Z1S4vGAhfD/DLxOY1em3o+WNAcqXBSpQ5lmXb4vu
jQ7tfBMTGmGUyOKOeo0T9f2dSL/FOXeTyOeTPaiokOGgot8QONRQG1uWNeeYrd+0m18jfhavVLWP
BEbVu8GgOx6fb9kRssH3yySFH8LX/y/IvvA1ekHiiA5GhPc6Ln6/3b1a7+KIsx//dhk0ewjnSl5s
IafXW0q48NJuXzngcdpjgNwVq2XWdO+5CsJADjfgzQKypooAmBDViQOoDLNlBkTZYQSdjzHKbBIl
8n+A2ScmHyjprmry3kq9RGGZdZ38Q7kwJB8tbQWNsAOIiyFKRPY+cKQ5clDJWyPAz91YPeUmZWxe
3zx9ivaNJpSj0D+Pq+LKNjELwlbs6u9jNrckTxV+6oqhKrqrj0fhflgVE5i0COOhBvyvufbbDmi9
m61PVOkoC7TDJ24BC4pZRmDVj5LwOWkOGJJGsDT8gskGceOcVoEIuEo3ijAOQfUTyVjy8u5J+mRY
8BqVPZYDQdQvS789uTy1SelSMwdUq2GHZO3ddeTKy4tG3F8CkrMrUZun7bNIbrbiDlUUfLVgsgmL
42iTBvuX7GorL0eLeKuF27Q8XbeFcaAGpOKraJvHrMwGdnXkX5bONszkVLTlp3beEPlp6v1PGo3b
uBNxX06uscRBhe5zwd7wEnUSg3kCP2BKmuNN/iV3SXkOsiDf5lY6o1cWVO2XNa9oVu8+iwPTsIgI
34LD9CF380JqAKhIayJ1yCSh+UaqOfSCRrV+BmfCytb1T5uGvqAzf2ziI1ndot8YvHQ93tTyQAcQ
cllYx48dhl6PK4zp9BmzWZRBbzGcUWqEg34507uTnDxIxGwa3RuFVfF3rVijvgQhTtViy/gHHZQq
R863Ql1V6tbEJpsnumqLm7YU7raNVZ5MXkdc4qYFf59BFR2/dKsAnEMvWlbj76ZNnHrSOTbNRAWa
jT/TITcwp1Gfs6EcSXJN0HGL9ppQKFs/6nY4N36gbmiHlh255FuDdzkXN25KTgwE6vVwzBtEzpwd
QRvjeyY6Vn7ze8VoHK6awouGCUDNzy7BtDqQGafV3PKCB8lUbpLglXS69Hv12Lk9AwJTesuiG5mo
B5JDf7bjmtL4CqyRbLZJaZVv9WtaHLHRXI6EqYlRvUg0TA86ieg0gF5wQBgPLGc5agBMjfYDJ8r/
xLJx4igmlazswb4BSStS+H4IfNPzYQwdiOXFzB8mhZKfTdMC3FiLDwGga3qkhiu5D6fzRfyNM4CU
lk5QC35qS6BJjf5fizHCE5B0ZgrWdpJYWE87qXwPl/bv/LUhLHTCK9m43Wi8S7AswWQc2lDMQ0KX
wGVSphvE1yu4NNiD64LT/iOwykkU78lPeRYGlJtWUnYUo7wOcftQjqS4kgQfAVwXNaEMdMR3Vegu
5FXxsQkGkpNP/J+Igk3wA/pBW4v3kzNslicujxD+C7FD7XxzTFTjVKspjRc+PdCrnqgOado1rehZ
mHWDOVZLLezgk/4grGbAlpWPcz1pY1D9zrhG7fs0FF5QGqvv/qGc6nASunYPoX7m5u/YZD0NfTej
E/IXBzfptU9CFsfHeZB6dxImZgUCaxD49kBaRe9MEJjySTZKqXVXE32pP7q6OtPhs1u/4dQIfjKc
KrFwX2+B8Y6ZcOxYv3P+NY0A4VmSHydewduPafR7wd2OgMScGqT3f1okXbK8UHpPLIk9IdqJblI5
eOC7CU35df54UH2NIw/Tb0SA2JojqVNCtQNN7sHipnHoMcsdiaTQSkDlcdddS/pzNcXLQoElEh+j
E/HRQCMvTKF+RxgJIMRy7bRDRbMRysQlO25HMcXxE+JeHGIWaP4Xo090a40XECXfli83yenNXmej
oTpRmkpiHg+Jr9MRrEkDlZi65M23epqn2OVY7Y3NBiEr9UlVUGdF7JUKxAt/KTVJ07TeV2Ryb8mX
fWkImMIGnudDPyNKVTWtLgYIhamCHDuwRGFENUrjWr3V6x5m28pe1A21cS7iG73h8pzwqFUDQHUK
Wpb4rrUtfugzCVRIqZNbJkL+5MaRp61f/EOacV65S+qctVcOmqTCsDHmyrIcMN88S4sBa5s/WeXV
vV2RygtvF9BD7kqHOWw5rNuhio9x/wvpaDur1+Cn9FbF63F7Tenc/tE5DgrkBPKLVI0OxliURRQE
kMEJxIPFmMGERIDcHF4WnIjt2fbmyvXGUhim01NO/rJ4HKxCGz8TtQen8mF1b1Gexeecq/UE38XQ
50uoBsW/ibGv+KP8gAhq8bARaduoI75hY3ArjJdw6i1gtZc+LiHVTt7HC0Yetg1CH/fSIaqJzjII
N87DLB2SlFzo0J8mp8rg5LAtTNPg4Nm38P4eFEvHRMySzFtx5KxagerK9pROkF0Fxu13ZKwbhRzf
KUAykCXV8lVg9/YdrhxU6eoe40iyOtWxUAJ6m9hW9L3vqp1Q40+WzSgzl8UvZF7DcfyQdi9mIia4
fXBQk+v37BbcQOxUbo2uXentDc1Z4YTKLyq4YsOoXu/+rVRBlnPwiOBqemGAOM61eKjAJCSmZLZU
PY1098RCHE8/Q6vwGCL0emC1J7ZcaZS0y+Gjcf/5+CDLii4dxaVpTaDC8vn0FiXKEe3te1xWKhu1
L/y3KW2blEI2QNiKoIzFVsB3Iny5DsK24YM9q1DisCCNXuKsvLWGNlLSwvVBZNGhPg5bM5+FQTFk
9N54uH1lgZc7X2U3jpXJCEdB4pYXc7Kl34Fyu/FlwnpdLYpeBRKvWfrz0Mtadaj9+D8y0eJNermG
RtlCqCnsLQ6JCeHy4lYBXb+xeB2bf6XDPzZbJjL40Nj59W7Dhr3tE4ABtCke+2EoGk/+My2nacSr
MCmFeu0WDU8s2/MDz8ywbZ36Sr7EJ2guGIcdeCDp2Nk2X5+C9ZGw9YMPnun1uRWy28LigAp5xntO
YQ0NI1k5GGBjWhhS5MOTR+p1eMGOplKLkB0vTnGiXedAMFiXrcNmwwoC0DOFiDURRG8QYivrBpY/
qZUZgDrOAULlqsIUnP7mpq4hL0hLdEFNGdyYGxFBmkx+BQaCwn26LpYpPiETrvqTqVdpQJDwm1g8
3AlyPR1qG3ohIzG5xtvW6jDmJGk1m4INy3SW4SZRKDcUX7wGYRHQpwMqHw5vHu9DJOLcErgPQZdH
8IyMw1RHYToTRttWsux6VHrP0VW0CnoXGXZGVGsWGmK403wtHzuYJKkVM67CtD4EOgdPx8KbwZZY
5IJYBRvAcehwhHNWlMQ5NsmSBHYf3ZiIA98e8LcVhCrlVjhTsuOjRRsshkg5nUNVZdFQQpEaceLw
3/wUwKOTj+PSLqoYDj64o+U7rExuKTrGuerYdxxzrK5XO6968pfNlx8tzc5iEdPPRK+DxCf57nKV
Zr9eTwbum1U8WLtJ9xWW3savcSsWBJDfz7Ti/Nt944THck092hnroqSPS/nhKptnJfEUVe0IEjPq
Y6f8Gm3yqG63iFZYp5c3I6hG37qD9u3mix4UvCKrrvCk3xhAqu3kGglb6SRmqywVDp13CzqgQGD6
0hizb/RVUi0Wq9+3fGxNlPr72WQug6KAJ4XU3OZTCgV6VZ2enR49AAN/HsyRCy2+lTwwp2clvSwZ
5nvCBWDd0rs9wcrbW2/Hk6IXDpPy4PV9kCg7db2qZzsdJ4FQTegn/Q5hFuxHF2Pgj1QajBpWbuYv
bcYMALNirRl+8tB/VrGqx6/pSWjdVrAP44JR6sqvmjJbDlpLlcnAfxHb6brY4zo6IY9QEqlh570H
89cHxTT8wKlG5t26dZKV/ZYrUaEFtfUJ5hKB9/AGAw+8X6HePngvM1iCFd9lXqj0BSnzBmvLwFmE
52NERMWy/J6W/1AJ2QGXpWBr9c2zqYtEdfvFCRtMEfK0fFpWkt1HM5HeDoSS9eqpP0HU5I+8RviQ
p1XxnSAh+tYDFgEK9F3ykIJycrYiW5y/YkYxPghXhGL/XIByJHng3+Iow4FtBWfPbuOCeOmgUFTL
kE3rP6OQlEvFMWrxIkcrHljgk2pGxU+K3Xfug8l+T3WKTcr4mkoQqInoljlyemkSHdGgo+GxpJuV
iptR9tB6wVxCQOP9qEwWTzAPss/qi/lX4yjkowqfaLzZZas1K5NVMSgCyLOLYU0reXCG3VnHpjwD
sAU7JKelIy5/bu5nBCqFHwdWV51bP+HtC6XEzQjhR5bDw6wQV669ueaJTk3n8Xom6zJp3EEUbS5k
1qVLyoljp8qouBZFjbVN/k0zOeaER+9CKyeOHseHLor5PcKDVU9xV3jSbLiABNevdvyr40N3whXa
optI1cFuFDPV2eEl5TDrW5VMJhIVp/N9voxjUmiM2+wGhWHSEorVOI1aMVummaO1Mu3pfFfWPhOh
f/zaJQAopAMEJ38mW2SrVTQAhFln5JyFac/Pq9fr5WPn/PA3N034lJHp7pDpoNt4k4860s52ZkFy
MUHRoYhYVhdAclWxQ6bD7Pp2hIzZhiXY/GLo0UxJAQN7vpWkVV2nf3cWv6aUcMKbbQEGhjqPpAMB
l85tcPpE5zq5tEpXpq+Vgnrug7/+DBK43wE17tmrnzY7+N+7ZVXjVLuVD4Af08/pM3KMWw898mUe
KKKhEwp4DAKiYGM5HoViyqMo6WCTVT7ktLcTwBJtUsQhvED8GYjAk/d+XarkvmdYFyv8+VruY7NU
m+oIhQFwy56MYhTFATRIMWaEPxqQzQecTIbyodluQSrtOfrvO+Y4662JxI4/Xa6E9JYcDF+ciqNX
zTaUYdxuLGb6CrkAAiwswu9lXKm+Gcj17Iii8Y0XUqpt7FEfvKuw1vIMsGJd1PulWBDprl5QibEP
Pku8hE1AfuSeEelfdZuLnfo4j26Cg6gzkmomD3U1vrTaB0IS4069XRGjTs2+VdJJujnLpZwiaT5A
MZNDNavvYxbFkuH0IKsbeqKk2l82Hsd9CEloS9BP8nvUlopS/k5KK5HWK72UOX5PMsgtj3cv3iQZ
+Coq3zd0EvcSd6EMfdgloYnLpByfTt0id+Rb2NC5nLN0bxf715gY6+UCjVUDC1LKr6zhokxBYT0P
V9l6iXNrk6wehRuhDlH6T6OulXZiTa3Jo9jTbWyZ3ZcAcKj04C271r5ugqL7VQvWlC/emRDgKuXo
m6k7MGVWo2ansAWve3ZziujVclkx/syu8jvG5yxWDWo1ETMkDCH3eBn0bw4c+RFbguGfbzfmIshK
69SW6ZsDx051LaPHkkUlgpdezoeL43akUcc31ydsHrXTgNWZKLZ4JmmJqAHPhFVZfnpsxOQXiJBX
niac4VGodn3x980N/J3p9k/TbeYH1ZFzZH4W5BrtcspWEa7wCIoomavhcHfkcNEmc65FJfGD34gs
9kbz78d3fO51p+ItZfQbrDBC70hjt+KxLXAQym9dGD3r04UBq0Gdbo/8O2coTY+ZlTW3PVefTXEl
PTRGmikYh3CKlXU6HfOj4FLNoavht2jACjpaSo/86XvaDyQv/YeAeJObCduEjbWlZbCM68Zz4U2r
VbVcAO5g/ooZbV1Al4FAARktpwcML5QvZLg/6bhPplLlqM5+CxwF+V9yJfiUpdPsY+4zzc696XLb
VPEqfe1sUfw+w6aF2LZmTdYvHW1d6UUU9RCR087cT7sjTT3cpTojxdF2YV4LATSF8n7lr5y43/mc
rQI2uypgtdUEBeIQjK1W5TZXzXM3kK3JbLzJ2NGaQec0Ba1U1mNSbOu0iHRnn8aA3QSHuLWHdfmh
4ILnCl1+K0zHjEmDcqz6cb/KOh3YDz1ahCpzuVb7j19Si1OcZc0APmnvEf2YDDwec+RiXghy40pi
2UfgrjX5jXVYVM6VTWf96vAwiF6ToyWHSEOoSY52CRiQQbM1hfwMq9E/hu+48BQbp5U93fQ9PpWw
/W52H11xmPeNM967m9m6HCpZ9+bdeekWUxhz8T87ur9FCe7ASRgiCgbz0VMeDqJe7bF9M3dLhVSd
l+5J+yHGba6citCIkKw8C1kVBekOuyw7m/hyLH11/28khEUZLHAMHw34vVPJMPwYHNQ4W13CvhhR
S/5Th9bM0qbnlgX3XjB6k70NX/YqyPdHweKeoaCtllAVC5d7Kdn2Jc3KnZQIv4e1Y2SRRkpfbmUz
K4UC5nntcgW9wWhI5r8jGItHpe1LXLL17VaaGap/8BdSChxfoLD+04uIpNl/aYBZw/vVVi+gT/0i
y3pTVWEzJE2gTgCpYeE8nf+p0SeWPDblG/jBBAs4JEFCrGuGLZ97OPzf7yilPkMPQKcdVXagJ1Lx
hTSf+f5HGeKPrdbCjvBBstrC6PaWtMDByabd7DNSBoDwKufvRTvmeG9kk4d/k70q9RwyeGqInBPj
SXf0K73y2mc/gQpjDbcAHdtkYYfR7yL2nr07JNAvt+suPgot2dFvqt9PxwHyXfzEUM4c50VLUj9k
xEoFaGlvWE2ryK5axmplzB1Kyc8mSTjne1sPEMrXZfiln9q/D2BNCL9hgRst3EdF/BEnbqI7WKHG
/nxXo4K6/5OmCqpKHcqJg+7IQ8i/cxfo0DX2b/LO7dP0vzKs01cPqExtkAcG2hXek9+UdbaJZyq7
Y37P8jUmDRTsbmxWgpsH9s/WBoFLO8KMUvdUcP66FxUq7rkmp2xDn6bzeJeFNB5y/MtLkz9ffREW
TsVi41LyFW71HwoioZIpz/FYCiIEkSaLdc0A2oJ3IV4QTRJ1cE8XoHHyx6LdZocp9o2QEC/yIc1u
sdOt/VETe52JFrZBsI35hJDhgmp2NJr+MqGZRY9+h4PGwlZIr+QoHGiHb5qfguoEEhDxSMpmt/6F
pZ3d0gwhUyOy7AboNMxPHwsUezkQmtDjUshzJIimzfkQCsHulojAqK8kXdUTHaEq+GAjVm62TTjh
Oxczyb2BrSEJRSKbnfUA6qvdXaO/reNFvSwipyizbrh84qI5VT9rjp+EKdlSgEPfyiEdUDCIVjAy
8Ge07N9bqUdvrEhmGEMEp6XtLeUy+4m6+HLo/gy4X0WU7kuvI+AIu7lc6pw0OpjxtBEcnM4JxEUQ
qlvP3da980syYRKI3PFvD6dw6qlmbFZrhO6FVpEyx9JSNDjbUshmtapAPQ0TK2IvBMAH112XYiqK
uCHDYdAeZ8oeIjNDS5AJoRtt65VxTagn1qSCbVp/fb9Ib55OKIWaXx41pUvjT4nGWnrQgOfj7/C7
mc2n6Admr6dokgQD9jOqJue5ccn+pXDCYxoqfZwKvaY1uPdlPXf0swcf3wAIz9pLqA9H00vTpOpQ
1uYX3j7mw5N6utCmXlH3bPHh7cUd5ViVcgvq+XqjQ65sR2ONXDKek4q3IktM6N6rGgc+mqHJ5feB
wSECb1756lUW6JpL7FyHm/Is2DUBvX79RlwHAMYNbszae5fAPfhS8U713fSDneDTSZiIYrt2r0xF
j7G9VqpZIJ54t1UoBvZHBvYUxqa/A5XfXdkdnVw8YAewKZ+pU5qCDx7EvLj0+OwoRO2FcDQ9NHiD
MM05UHLo8zMwoy4OhbqnVDqeXuNrjbODo2ai6aM+Rnx9c6yyuWHwHMO1Od4DWqCq4KusVwTAc7+p
FUqphS7bfUTFOaPRlKpjCUqWe7wcRXsSLyfu8yHeDGs2q6ClKv8K3rl9BmxjNaa1n7O1PuJnJimJ
MRnrdidGcMl2nfA6M1UEnEcJMdP6jwXmQ3oWsscyQOSWMNDVsTQ47AlcEtXZiqe28vH6HmBjYIaP
anx4TA80YfQQctJCLWK7yWwd8NMsQOr9ZxWDs2uqezEm7YQl+8Ms7JoMWXI2vecPvHPRiJUf9KBC
9scymJLEl5fm3PHEoDcgBOJpsOElwcYGwOVnAOM2/Z0J9RIgoJkjYTaRvxKxxGuhcZ+HPaPcTtfH
49k2gCkNehl9x421k7jg6zXKwPisbdcZitH1GLYZORjdBjwmuvPIlLioFK5TN7DVNjwoM18AgkJ1
rdN8kx3zk9FFJis5VLqER8NHK0MG9+KVJHcPWjEcK7qSf3PmKvIFjaeFZDY9GgzLWT36O9e1KpMM
lurvos3wkIUvxGofsEtjF33Cy56TUmdMIwlk5DOx1OutQQ1MFJ+K7f/Eeu82oMbXRsmXwmAmgTJf
z1dJZF6zTDD4gHTdDeF40GdN+lzeS6gyquJxXt8NzFjyCmCU7szHWULdSRP/cyNmynGqY04mt82a
+NrUdmK0qc8PQlhMt5BeMkUnKqjNR7UZUGnoFHKs+2SwONRjMpqujA3Tkby3asIEoCpzAbPvjyZ+
3V/2lL8i/FV3n0J3MnnAR50EbNdPCQU34TiAvnLIVO3H16QcjaE+b28uWrofHBXp9TrGyoEjxAwt
t0gytuWtiVy50+EQVWZgKDmGWqgpAJ9Kao4QLGPPP4b6TXBD0B1zYIiVHeNyP4peGcyH5HcMwf4c
RI7EixE0J5KXxN3XkvYLgNs137AHrGtZNJoJzaCNQKTyPht4kAVXuCt/W4lFCd313Pp3py+7oqaH
/YHuABQy52/kOx5SVlCoIvC+N1sB2JA+HESq07tI5J0J0FvX6FL/7eTU8pK2R/31Zbb9qM3LBPaC
fhT4Psa+mZP0YTZLhOZc46nURWdl8oWjDAFoE//yWXURWtTY7JYMzfKCwzbX6ar3IOHmxerDTSbz
TQfqRBoYIhSnWbTYheOqDm/P2mSx2xp6LQdt1oMHN+VkRno28uhJZ2+XQfqwZBKavFlSi2tH1and
y/dsukrCrhY/iYuejmBodYwoxOVx0KlQWOq+AfO9GufMp/DgLTBf2G0UYYAg8pLO6YrgULkRCtkE
oTcpAMIkuou1sWTfYNAUfsJY2dAt6BcU8xT57QeqSbtGaCtZy0tH/fyrb4taIdMN1ND7DvYyAUcp
iSozrj9wkCFWDMtjroDRsMdDoVJ8O2xAUv3AG+ZikZ0ZIT1VSueeARSOrNkPBUJXVfYh2V/zn1wE
1gpDk7yF+lGpoletlFnwXiMRIwtC5EHewE63Xg2C8ZdPLAcSDV665oHgUQa2VWVBJQn/ToObKaBa
tnTfrmBSqWB0+CBS6ZcpSUeqyPdP6KwqymTWkRGagPXnl9Qt3Aj42qIUDM69sS7HX0uM0T2Sdkwd
7pqn7todRdkDhVx4cfuQ0tQbUaVEnrUroUnfs0Q8WlUtHYRPP8MJ+dzNijXWQqJjXk8TCmL67KdB
NRpSpB4FqLrDtmi34i8nBLb3R7AWgW/vWKF620kqFI5X9dX+12ch6vlk1zRB4SpGa4K7SF77S+GT
2hwAFAkfU/Jcko19U4/Azy6gvUHk72F/wJKICd5JhS8jvBVla3ZccP7QdnGU/Xda6DWDjLLYo8e2
TwG9IbYbr0cNGnmHXi+gJ7DhGfu5yPwL6KqOhb+RwYi/AnWzSTQGwOL9qbEA9+pmg7vqN2ntPYCC
lLe8XSrEc7wkvBEbkI9DkaAYRFAVk7A++2gBLRYlPdzTxvHHFYR+4SIQkEDsdUFeGJPpLALz9AmI
jLOqeobZvOfNNUeSoQGrnPa6VYuZD/EJLNLdLWeseiu1t9Z4pO3+0RhnEi2L0RpT8x9KRtORFS+8
Myu5oyWkoL7Grw7WWua1U7hkH10r8H+B9kh7f0t1vcBjPH1XDCsZdXzGLDqjGFK74MSeJRUARpnt
+BD5qtjFmMjP3FLDUJBAH4dMA9XVuuJgXL/jBUCnSF7CYUZO7OSNo3I/RPyADrGR1/YdZRDtbZuJ
FgXah+x9yOkFqtPHp5pQHbCe9Z6UZCnUyjaQ2IhJkNiBQSu0k3ZEmyXGar8TbcUYsUZa8hUNF+LM
a0P2DyORRf+4cXj+Bpg2nQl+r7IVJL2538hGgtKQPP8H+1gfoEV61DiqZsozVsnZHCReAfedtGGo
lIawdu6aKlrPmnWwl7zeJqldywdPBjo4yldw4ssW7PyvDRqFl90u+363MBTpmG++jl/FsMTtA4GC
/kvkUyVP3P1lHqC8yLCU2sey9nZOuWoHbZ/sbCP/KFjCB+Jq23f2sj1MuahhAOmGemwHtPvsbRDH
rnV3QbedzBc6foAyg/Zg+vIHJ0/UKQxsmje5+Jfp/c62JC8PieXH/sC4EBkh7PBOTlCLsSf6iaq7
MVXFFaDSHpxBeYP7Yqkob5bS2PQna9fRQgPnxEgzG+W8j8dqSuYvLQnIZadq0uMpfHwp2DMy7Ez0
GL29i5qAnbiDzr5OQH6IHEa6fohH2jngB+ViQKf0+WVqwL1XlLwI/SNdWTA3YyLqABgMzS5mpGQL
jnWCOolCYTL0a1r/ffNzZtdvh6VBAR8koJbe+ZYBRXlKr83swAUrz8hGzCZpgEbKNDBODHKzpBZj
mRCiRhKTHc8MeurA4XvIJuo5w6r22ozOWOREvE1RKoK161/HXth/njinOlNB1X39vEmCIS1Jh1Iv
g5Rah4N5ISudV9RxKIaH5MEsaP+GSEToVu1F4EcK8vrqE3zpdF7cd56MCtJpP3gUmliaKLDgJESF
D4EDakUg3JVN/Htv8Fp4K2jbAf2omhTXTGXRz7rtGx+ype6lXSvGcA/dFOTKH1IuSO8Ii0IGvyM1
9VCAL7+aDEcTIgru8l1xvRNlw5Q7F/33FTfbizLHwyrlI6Tbk7aikFyxMjrG2+DdS3tc6/+Lzo5H
fTTheaNUMW7iomBK694d806PI4DXR2xRCt+HiSqmtFWda4O4Go+xnExn+cmDazOb80bJXmBpuLxX
ZiLRW4tjXKznRavDMCcnk8o6AHbmTRM9VXzD9pOeRK/hbMzqCfOif2u9ki7SYyI3eOqeJ/UJIPxy
cUQcZQnEAHJhI6bBmcT2gq+NptH+1IGVyKHdafk17tYqgpxGtg6mkWnsWSqPIsqoUJQdLa+HmaYw
953u0ArKT3hCjesuF9PjxkZyzKqaz+6MI1i0CYaRXrgQzLphIMevl9IBRzw9D4T0Vt4dXh7SAIOH
1JUzh1moChAEoMP8wW+WqYjAC3DTkl/7fZD0nl6W25SDnnwGWOGFaesxgmvlantobk6IVv68jGC7
6u4puHtydqb7C37G3KenhUDyVTrWadIuxkD39/heNuS4AuGWMvGjeynmoTAVd7JWydmToj3OtCxX
qBPn1vWsJHiNpnVJS8U5hMeEMMIfy+9N8vIqh3qAVmoLAnqwgfqeQ2feHSbtFK5bX9EFVlFH5TqE
1K7WsqqjaLCpKa3X3FYw4pURDRbTxEFYXfnnOEbAOr0YbwdPEMNvqqpTJ5uKep7ZxhsNbeDD4bGv
hCPV5mlPxVS2oxFP/RfIbCpjM0diwo7S1i/HVHLrSulPaa2mSfXmTcgAWbFhfmtKprmRpOH+XJBC
a0Ruh2VOybn2nXgvsXUG+ZJa4aFOhFBZp1l88kUSJzJG27f5g+Oi6GKa5lt5fB7yjigHdK4E21aq
f9PZ6D1q593Q/cEOnG6JkBP4flnIbzuoKrPoyDX7Z/u7vJuP/Vyd+RBA/9qw2x1bwj1FxE76FGr2
qD+PWqZ14832S8lqU/Dwgf3jHlE8sR6G6jnPttBP3XijL7KswWGS6+Z6V/JtLdVNAta71xA9N+O9
ag8kVVFRFUsqj8opx2pw28ietbtWzWtmebC7w1/C7GfP8bKFrp+dSo9AnEX5umsulki3ThWNMNsg
o1aqJKDm2Mirc1qZxNd7FSKKgtbEuiRd2zW/gsQ/ec8YDRmepn+TpXibV0GViRP4k5a4mepSa/a8
FVhD4berdMXbpXa5PAN7DuF1n2xYL3hYUaUH6z6GRaHnQ5/eDi+lT2x11H1B2yEdVmzs9R+PwMYe
sUxhHtemHRU/zA3KlnOYYzrX6jnKymr2E30nLDzjXeo13e8e2gXdXAqDmV6H+iDI6gZBqk7QwMMP
u2Mm+RrQtSbAUACB4ozoBX1CPDjF9Zfa6kHz5YlQsvg31WMNabIS5RszLFQAAsc4u32POLacOaO3
d8JgbKL1gcMzT94ANPBUvfsleGAapMKuO9/UrKO+QzIgEYLC18wSz0fln49qoXLHP3XBJLGafqrg
HuR+s0JBVOncX0Qg0e8A8wQwB+vA605lGOxd2CsBD4D4LEIQE4iJyzTZAxMgpVr3HjRLRtKlp3gH
a+RTE3btq1inx8fdTTZCA74IltgHvq51uxf+E11qAsb6mDiaK0QiIC0R/eycFo8pIqk6oHbv3CZR
xJV9bv8fee+A1JJEAiABCzbRhyq0TRKCg1yFaMqhfn0xbK8Ic8oUBkUILPTyxqUXGfLK/GZBdTpC
LwYBoQbRADS9vj762RK3hbXxzYMtMAmk182zqp9vbmVvsdVyrWHrDGiSR1pqwjXBycq9mclHyPfE
ou2wHZXrC6KbNAdzgEctxOvWSa1q2bpWb8MMT7vNB17yD0jZxzXx+JeNKpkPYdgYZzZTgJgS9dt8
bZ7kJwh2w3bUuxAAmoM3cIs4R8Ys5GG+oxMJMkB4vlY9rT+BoXtLDX2T2+osXE73udnfj9U6gyfQ
wefSA8HfbTLMsxnHlDUVq9Q1LxPbW/+77KYaF72Frx5KOuCmmhawA9ULcV1byqHJwcyIY7paI4wf
5DvkbTHjHL+mUbZLx/4Il9gSPXnBycLpBNrV4/5Lo9+PdODCnafj5K83whgI1vrrCNWaTam6pjDX
SYWRma4Aqr0avBIBl3dTnYX8VumcjI+ZPcZKAJZFgQLUDdKPoWRZwLtJ7cVc+JlZn7J1ZOGQgUTq
H7apPEJnk78/qBSU7WE0BII6SncB+0EkFKk66Bn87f7lYq2397g4C2OyZiYx+GggJedeXMDFiCoH
Atr5mPuJ9XHBPPiHwNzUmYsy6eW+33w+b42jxFQOUQ3a/cxNECrVetwphRwu9gkxc4rlR2y9wQ2z
lFS1UfKBzCB3FlT9CfxkokBVDdOXYTfbMXQJdOLx5kT3OHzGQJmrbgz1lJFfI9A8Ubgtg6ScOLLj
RmgpX2IVYV2iW6BdM1JRp72Cq53ZYomBy7m0A90bsjTbjtcLV5qYHJRsp3K7NUzLsE0aPVxY1Xo4
D5w9+1eRwhOQ5U3n/bXDO94uzv0Q2X33fc/2yo4fJu8rBBY0Anlbgxn1QYFvRsGNLpaB528ngLJ9
6eoSH8Ipw13qlHPELHeARFXmpkf99TnS9OLvR3Tkg7RnW0/jNZhk2w+bLU63NEXTGNnLEtzVrbVI
fQRUQbdTM5Wx3Nj7PggUTKrGyMekjH5nx9/euTp6kMEv84krVL792X7YiwrvdRy4eV7w1OlnaW6M
Oz7Zh8PdIb0CPWn0chyYyKDtscBwHFvN0mdlGEM548ORqBpPGJUsiqWVh2eW1pRjMxJOHSgCPv0C
VcVpEaB3ilhj10SK3ZXQA+nbj7TGBvDqkd4kA+8Q7UYmt0tmBtxL2NuE3NH/0gHU5RQsYy1at/3Y
e/97JkrioMjXCyM/3NKQzUOZ/ETD6YaJXHQEWakMoXmrrNpMOEe/Q/bd6hGAGedQ+lznFkUpAkaK
ZMjDEc21FkLU3nmiL70VwUZbvi4Jh+o6IfsY+CMlcN0SQXW0YJ5ryigiWGA0geIqgtyKJL7ZoWP7
Fy749AInyJ+wLQS+W2BajpRNwgct03JzaJ/+Pdmv2y5JRrjbOwRFqjtJDMa5iVEuE0mvQrbnADhj
173IHpu4bL8gEqG6MOe8sKlZPQJWqeuYkv9+S70KHKoMHjpaqRhEwguS308Rxu1E/I3oyudVR4Yr
99OSBpw8FXLPlmyW0YEmsgSngHd1xN7lCvdVIQuT1rEcatDfvZXqH+2Y+wK+BODah0Kizd68gWbl
fc/YJc+1E7Liz1bCpcVFtZooWu1ilqSrm9ryALESmZJlMWacSHAqJudgVPylyHMGmCTFbcwT7gzI
pn/K4qdl53Qp/eXRDkiCnoPlB5j3cmcXhUC3e1cMtaWtupAiZ/Hc6Nb7G86lmai3V5JRbrCA3wrA
2IIOdFsxFJUlNRXwvlE2zsG0LmeaSmapZ8Fb7CTK5oHtNT0wTl8q/bkcJzCxU84T94I+2T3neemd
ABKDSRrFqLU/3O/zwwTwuOjvE/7JKSqiL7tIRn/Z6cEJzZyrB4jHmhcs/gHfu7jpsOAA6z1JqUEp
BdxlAtk3m6GJWev+50U6EFk8JDrLXiuUioC7sh+CqB8pX/Syk6gub9RDFQBsWonguiTQhNWG9BDK
yF/wgc34WBrADIEWzx2zQl2fEXZvrujU88RY6K+mOw+K0jDHJhAe10xws/bK6I6CHbhwlTxBz58M
REqDZt+PQ3SPEoImUEkK05UWLtNNoJpVA9w/uknGrliAuSVMernvMwARCOMGr0/4usVpiLmRFd1l
1J+ICHstTpDR98UkHqr4qFNpN83iLTVoBYr1aclKJ5/qdEeMZ1SjJBzkRCbuMSMm96sF3YWuTTgj
ug5zKCw2fjVCfcuClt3LpG8SELdTdvvJCvnYEC/nzbVJf5Z8/20kSACBQ/X8+h9kwyC5kVNJ75xt
/JEPHbIy2HBbHOzn6iEciX1iOM7uf5l20vnWFi+EGXyURseY6tBwSOEseCXENsSjaUbjcq5rSIJj
BQDAJsYcLQyBGf+gMfxZgMauPlKkjVbKfnpli//lYHVkdOrqAKe8tnK8s0tX7UZ5Ng7FHSCZoh3t
7+d4pGfwSCbLuoGgDE0xw6mPy0HxKG01GZoRlx/OcA2snoNEFenP5XNBAeFhmr249+u2L4MvGqV9
i4WpnAA9dafHas9Y3r+WC0rALxSV5e9Rfq1NKeOK1ulUSVFSq8Mtvs4YAiKvdPDGGB1J7L8CAozF
8nyutu6yrVqiVrE5azVdO2mhCD9KjCl4HT6W/EqE6pQYfYKemyuspLR8eQxpY73ESYDdK4qtcQhj
ltZWXS3alOow6m2yov1gW16iaZCNC7TnrDTnFHx6lVHs2D7MzuRKyFuiOJvsXhGFpw6oU3cfH0Li
MbOhMd7WKxJ8erS4+zoDCO+VKy6oApwjZ451YT+/CHMu9Q+bzYwJFHnZ8wzei7K3xx04lmBojXSo
eNYapJ9Lkco1I2g4FbaDv0Cv2Bg20R23SWD5S5kNfqzfAQWpwZl1VpbjAs1RBUuI93y7+QsWKTbk
aIbqBJ3G+s2p3LVui11+Sv7bdYr/yJ8fOt0Ffg5ZfLY23WgpUnLaWb5eB25iUfTTFjhKi8d7waV+
BH7qKOAQ+oh7EDyl/WIzEzhHo2Ej72DrU+iR9p04xIsjQifBAIuVACdu5zhuMpaM+3A8yUwmnO+l
ePdiaNWFqF8d7XyjjOvjHWb98ix2S5pfK5J9Jtaj4DVhWQCyXRoo/EdtAKo9XHrbZMhbG2PbQ4xq
2V4BUcnIacgDlJkoCaai/iX0KjvmVIsK/t86FgocNbd+G3t9nvt1VLsJGIEXdMtBwd/sFqaZ92oh
AkARvjHgPI1yolwqipmlr3X/OWoxEFtlRVFGSY6p8Sed4MtEjLs9sKjNT+ZYIIj6J4J/dl1wvbXL
n0JAOrr6fBEW84PcLIymBBuOz/6EH+FQTtz987Kh1RopEnp9up6xIuCmaZuHpWdpqPctO9yJ/0rK
Uk3fY0ruvZdkU51K5QLiN7i1pA4uX+J1C34qMMsK2uYvFf92qFM9oIxU232e5AhQM9LRYeh0WxqT
A73oWl1YQctbYHFtyXxHG1atp5xvWf9OGNvTpX3scy/Gc0pYwnqeqQypXKfwL4BWhQj75i1vVai9
UlqUrHFMaIsUQwvbmnwiZ9a4ruBYrF4ojnPl1wIBXpFJzxXnf+KB3vngmRkgti+eGSEQEwfUK3PL
S5jxmaDAKoYbjp2lvKaisJMxLFjKEwWPagAkq2CS3gni48noiZC+dad2LKZ3+Mzp5PsbfGZLIjf7
Q/rWqM0y1H9H9RHNprneknSnnAH1M2dnRYTvbdCEZ7AlbaiCRvWTGLItg/NSV4X/A/8F+6XyF8cd
M+6sEB8RLpm3ql43XhT8Eav1ErVVBTfjymYQjxZ0XNK0wbFKc2cXDkmaxzHnMpT+x1r7KEXaKJSt
fqYU4+46bRKIk6tpPjOJqEAILVLZhjOshSSIgfscaKsvYtuGs/L3QdOD8HoDYJMWEySTw4kE8Mc5
P7a1COX8QlVipLcD4d+ktpR/XGUMWfVAhHf92dx2sYNeyxCQPbh79tPxoSyYjT19NS1snqkXXSKe
de+j2FQ9neOO4XHG4c+dot3Ry092Q54V6N1cTEJKwCXk+y9gu5js+vU6aSiWyxT9POvLTbIjJLcI
FF/jhBwR310CUE1Wazf8O9yedRuo9tvxapIsnQi+AWScEue2UbT35Lst4u8WiNKuExP02ANeEOhI
pT8WvLc50/EsLXRDqtpUCIbMqoDGzNAZftvMlFkeO7aBWOmPTq2+nbsDPd/XpwefTqChcai/Q1AS
HGjmHCLPHZ02fRC7mg9RQYMoVTfJ4Y+t9+2VIBA19h5Es+gGSqbUgNDmWYSAc9o2uk+t1JIA/536
jPTg1xngKG1Xe3S9DSkstLBsaLYO6qw+ImfVqZqgJQYnHnupOer5tm2gRmHaPuCPa2GG1qsGn+zP
qUYj3fLHl1i1tMCD9Pv6cfgTLyLBGlo/bqXpQdRgn1NqseGjPX9R9ucI4pabmMzMzkaA3vMSugA5
2tY9chU1VcOydUGr0DU06IkoGuKkwbIxkN33xeAWo9eYOC5akkDoFfVA5BwPRSk8vNpxoDyTLJWO
HPvom7YGl7nkitLIFqwqA3mtcTSMqvnv+S8EDgAfA3L2MSKGgM4zgF39DuRB2UA0mJYeHmR5vjTE
C2QJUhvjsPhRcYCUbZfKqRBpKDEdAW4zFFCB5pNsKvSv7JTSjDh3ixKCr2Vs6ladyPL/7CaFVDUu
sJzBRv7oqcZshztZBwDxrYAsBqnS98KZdSkXzzLxY8Ce4JH0LYsq5l+pdNDd5mlFPO3c5LiTVPr/
+L8YuOuB+uEsdFGXp2mGHCCYd0uoS+XxFuDwvag3heOMJwt08T4V2DW/XOanD1F+2XexFEEsHpzN
h1ObWG0Cgv+HtzM2bSMIL3PkLFlv4mp02R5g68MqFfTNc8vmJATw2jAhlT+Z7v+5MxS5pz1YpObS
SFunyv0SYDIrHIjV13LzWQhu1r2BlXMxEAHbzwO+TlVUfNpz8okDZkVzBedNLX1Z61nyHtJ9WtQK
mHg46bBszPLkaVUBc+qKOTVWX9DhZZ4UN2u4FbNnXWmKxLecg9mTIBGj2wCzi9Wbc2b14+pvsAFp
pQMiLHAl7e6kcMNq/8k7taF7jhyuJIs5Ka4YziR/lWRQ2HncZ4YrNV9sjA/iBsM+IUKO/fcRFlJa
s4QDOk/dmc9b4oXz0HdQICDe5bwu9Hn6Qr8C34g/rd9LOYcJC0OSKmsixf61j0SQZ6yDDt29oJtq
0NK7Pwb1+gejJPnqDzWfpv1XSxJ/lyPoMypG61CEbrFKrQ0f2YyYrFr+/TYdGCPd6bqOU43tw6CY
Xqv8gI8C5E/S+PKKDmNuiTqizH2J+Glo04DTAautqZt0QoobKvp9T0qBri+ckBB9St+VN7+1QbEY
twMdRgV95a21G+d00tjV6bQmuZuJeAa2u5YH5poZLl8hYvxbYeMBVijYYI0A05B+Es3YSPfamk3g
oOofEflBxVOpCcelyi9wjPsSDkqZ2Ct3xaB7er4EtUL/nyzbXZsa1t5CKTGe5sQNdkjzP406oS0x
2uQX5IwacoyL8X+GP5HoumgrKYdb8KOJYnM1J+egbST4GiGFsZrs8LJxe5TOmpPmPIkCMOKN+dlG
EMmAA2zO48kPMRfA/coagJR6+v8Pm30IxQe5BfNW9DU/ay83bGK1QFcmTvqI1w3HfF5UpEaP7iFa
86z2Cd9X/J7VTkDcgHOCo2ptUB7vJnSgLZUrSfCzEOZutwUPf66BFTpoKL/k3oZe1OHKKng9rMxG
YSRDHZXtajxw9GYh7m80AoICXkZBKm5KNAYq17QdgjW57iPzzX271TB2GvfkgonGkbEaJ7QtS1Ya
FDzRTlwjcuvQ9LkP53iLH6qhQmBLkOaWebKfUxL/Ma1/mAwTzekuu/DXOsUsKIxxaI+7WORDsxbR
rSxr2NQiHeO+viYJ8/B57CXAO2gWrWiZmjRCDEDpxep2L3I0CGrO0nX4dekY6tkGjTIAUo/toAUv
a8m4HcYd4VRSqUrEWkBmeQrpPIUb+zBoRQYtUIcMBDpgeqaiZgHVOtmSgUMm/tPy7bu2TxeQBJYT
ctTak+rSejslS1BEjhIsNHMWFN2ZpeGAwoCN8J66Obl83i+JcCRqfoDLTdcnsZW3UUNdD00SgiUV
2zZ9SzQo7HNmq6jAajpHFPouGKtYvP3edDTalTiklF3MoOS1lco3n5w+6Js/xhF5lRQs+4hppjeC
p+D0itjQNsTYvcsBFOyQ3YQX3+jdoxQ71XONkubrvvqNH66T+pJQj4hexSPr+nbIW1U2ilut2SAZ
+PISDj8YqB6bsh8DbfN7uRROs9oDhmhW5pRtpU5xJgA3fJ4sA0ChIJB0juttlv7ilwKZOFRS0Zf+
KNjby3VFkEtr1BZo7Nkt9VjQrF2oL0RP6t926P5gmj7p7MQ+7rl2MPoGJW/BSNSO1+O9+/Yidcxl
nALyNBjbzrP7uTxqhBkVpf5JsuLJeoTPfsLQ4g+DJGtmsmzeVLMUoH3o44Bh9G3cN4ISFwvGaf16
fjwu6vr48X9YCxUH7igdFeuy9SZaMPZjHvepfB6B1vUc90MO5xjH7P0cvtKXMzKOotRVjxezcoAe
puxR2EK03vbt3LV0fZUJDXsUh8raunJ1mpRlpnYkIc5xymP2GsB3iSGuAitzqeyFVOsA0+YMf46/
vu29+Nbc+Bnwum0jNI3AehmdiKSptJrJWS+OxD47ey+suQt2m6TV7+8E0H1dhlWy/TDy9WehKWuB
Rp26AhS06T+Wv3Zvm0g9gztC8F/wnX7S9wae0RJIh6c1eKj3tK58/54Aam0GR1tUTMlAoXxTjkza
p4NhCfbIOrmPnNZgyMcbMfGdZ+yZ7yExYvVPUJXPJkCGDjO/wt9zMNYVPVTK9wctITOKwJBx0AeH
R/DPwjyVEmIaikPm7i8Nu6hgdrdsJAmCz8OJyKP8ckbrxvjHZjJCb7hLsITpsAIjuZDOP8Y195yi
/CqDHc/UnVdxnA39bE6kAbebxeMVu81HiXM43OHO98hLCfiec9wGfYrOm5J4C4wPfZn6QYx7YAFS
x+yQOAfRSKBoqhQKO6HJoGCqlVsrUB2CxH9ArP1zwRP1L39jjVHzgVS8HsEN1zcPFvQATogGS4Sz
c3sYKMvjLID6ITtnEybpgqUcgZ44OTA+/DuNcnEgAStcFQTZ214IsRRjh8ER1vtDJfGflldcaxpl
Bz/h/Y1k5nbaW3QwtsWj42JDM7Ybpp5IAa0K+33Tz7aUvE74iNO4qtrJGqrOc2y9f5pKuoSZXaoU
fvAOb2aob64xKr7mD9H1HPb8nvHKKr5/Aq6rE/4nN353UQrcdl8czksa3VpdICn0MkBpgDA4p2ly
Zv9USPlyXPi1zk+hoTkNOPIOPBG5cv0V8S0JmHI9qJnL/+OYtQtbKMy0XRoh8uqfDYs2TCVWJDwc
8eJhZe25bxqAbWJoF9JK/kxM7VEQQ8R8TdUv/ZVoUJf1JgNxc+N4X0zHAcg/ps9f0QfgwP9lVeff
wmajgw0VhscknSnwS+7SxP/3S4SH+WIosNhqacgdKQi40rC0esejsV9WWuzlB8ZG3ARdo6FrDdR+
BJHmdeYEgK5cPOKf8xSxOa8rvzDBr0JCdb3Y7a1rRBqBKl8jFxzMj39bAdY28TEZqiPSSbN8aT5g
0QMMvsvIftaRNBK/toZE7P6BIeDoQQwiIadpvzPFBHtQ5eu0/Aqp30cqawzOGaRQH9DKD/WKPuCV
8L7AxnxAwDJRzzRqpmhN/FGDnynQ0frIG4iF7cX/GiPCXmVULp0j1WdbNbv8cKnLlTGmcZL8pXFY
JjcPTHk+E65bqbQFXBubfxaqD3G5woUepx6B7RPSkr8OTR5SZKCQ1/gaQUSCbNLCryjibZJuBoX6
IdQJyB823NkSRnLHPJHQrVc/0K/cFngrc/lZ33O+WvrEmca5m0lrOrbgmgLHIf0ghE2JQleK/qCr
xlLhDHI4p+NRzHUQ/f7/P4NL0UoWFoc9Dpx08eeqm8ajhspGK52nNXsN6Q4xnLrWlmArpVhdzlO4
foqxOENotu6LMu2jCQVPWVVQu9UjMVwMZqjmYPHAKu9nrT4s0QqVwDojfcEBxJZNNJ5919SmPeFc
jZrUZOkQavewah0TXPS3X9XQDcHVzpA0VH8NpmQ3NtkebHpDZCVS9ne1vqReg6xbLFL4m0wtimWh
EqZY4DwIeYIFZ6iP8EzSVQJIGagUPZRpzpGwR2UiwohhClO8NNaXXMZ5rqNRmO9K9EEhSyXaBg4F
ypgAXCiRiotooSbnVARjiH6MDjx495dOLivUfH0VZ1aQVSS1XUmRQCUsrZjCy3Jo2Oc+FjIjwTxv
bWpsH/FSNnh4R4M9VjdAWV+Xx7H+1rvorZBr5dkLbj6NiThdMbcxE8VlaZBsS4FwwfJQDzKOmacl
ww95sWOXgRPHNNLMdYjMeVaz/4+m96QkTXb9wUaRmr8uaXPU6nnCC8Qqm6Dv8CV8M8sqNX8xwE8t
k5Lhj4AwFAnN4DXd0qYvM9OtTTgbG7pdOIK2u6osswg7R5yf7GXKapYfFGkFry43GWGfs74/awmm
q/x3KjsxkoMmIf9T6KjO9WQ7Fob4xJ010ZutW02ojWOfeWhxC3Yc5xRXG6Zi0SUf/CzlzbBXUF0k
HCy1BEbQrdotStHhnzxiXfa2mwnenwzFgbCna5jj8nRCvhXk6s+HXKcXzIZ5m5JUYg5KphP/9P5Y
aVXDl79rm9n3jqIVUbkEGNVaYVlTdMPLKZozOw5NXVVRmeEOKMa9+F9NQepk7UZ/Fl04fo15SPT8
I/MHaCCQ0M0n0vygCEevp2zriFwMbaA5ZsjkbOUBoJcY2ZSaQvfNj7w/ltdaz/eDx35Sjbdoksg8
tQCMiSIvDH7NOpvQdFgY4YTzVGZqStfVngXk+02j3Hq0gke5/s7XgEPHvAKQgfm/bJRUsHoKu0nU
zbEtP0IBZyxPAaND+EilpNUJxxY2wVAxZGDHu1l1en0pNrjGgPb+0tUvqXUh7mN6CRWXanYOghCi
gbTqrITGKwTzI22xKKTd/3IoXvany6oFOrQXbuvBXnzFrYR1vc5RVVG2hf/+KRpmMRO0Zs2vhUOP
40engePiJHvCBBEKocLG3URVgguxSe/VpH5eLK6W2T2hvxQVMcLTt4csZnngREpiqisE+1oduCck
N25B0Hz6IxWZ6xIwoonhsWa6oabOoUYUKjZdI6l1RFG7pKlEnTs7+hvag8UrfmjtvhP7FNzBDPau
TFAGARmvH9mfYdECA8GUYlg2L+wOYwejq0asKXeCEo9vgakp97EcaPNLMx9o4o6s689ByIeZpf3I
KSNKjHaSLu+pOpx6zq0lLhlmP4/NoQBmk2TDbN0v3sCd4K7qGCAl0DJh4b45YcahldmfRzmxf7y2
KRGK+rKoPwDAbCk6sROUULMZh2aPWO9gal6Jqpk7+4H1a7lYsuHF+NNC+I91N7NsOkuthfsnzX/R
QLes5XSPKiLBFUQCFlt0O+e6Mydj5nTQ+64bxroKBye2EGlmibTjffuuSDdIwszj90P6MaAATn//
jeu1NPoG6sc7W6g0KfAO7MiSnVRjJZ1UY6nxzEtaJEwL82YSJPXPq61m4fmSAfPBYUPuA7XVQzj3
QglyNfl54TLGAXQGeJP8z/gT/zyF7bNqpxG7RjVpUyMVNrcxPgpDtQE529d0S/SHP5/kgT4B/OE4
zDv5Wxx/+QIeT4b0kQI0dWIeJLIurYTFyi2OtJ80AQIIUlp6Xltdk9BI233uQaQ+GUwgmjfOPfSa
MAq2sFR/lS5U8HXvKkjxgTuCmcMQ4Kdlu6H0TkbyVe40RCTKfFCcVqaVC6ADXsXG+qEbYdUuCsNB
0kkLueRdlPU8R7VsqM2Gazl/kHRXl9PEKvUCmVuaXxGPOKlwh1yFEmogTY5NaSMxjpycbsU9Uy3F
5ZZJY0ygb09vTHCHhtvgV1J44qMTJgzpJjWOikJ41ep7C2g/E6Z+LzAU6NcOc+4HV3WdvFpZCW4Y
qW5RuA7U/1B4S3/OQe0jPtzjfndVPwWHIjsqukg8NDKz0pG9P1q6mFC4dKKM2DkpCR97DLxDNP+c
1rg2bzolUX36MOAhA9upp1GGTCLjgRy5rKvxUVd8BR0ssRNMGLN+DdYg1g5m7W3J/vmMaORnR/Us
CmP/jmxPbg8RTmFRJcJMjiypfpRwoFvNdg6Qw9v0k27+CVGTZpQuW2CIFpqr8hLw5LGcHEGhyIQh
+HtL05p0eqye+WGZOiVnuA+tNGcIlre7eWE78BcNZbvlxCSb711EhA2dPUTfNGJcgG4tYnjhNiyX
G8nk3EdM8YgH42/6M0BBODVRmtbbDO8LSap/54hx+JekCtK5RNcHeDrc5xNG8d7bEzudGl4M7W2n
LeeWflB13WoF4Fg11pZEmv8I3BREkfkXXlOyAaF6V27psgi4C0NJXD5VZK+GDnDMnnkaS28UdYJA
XwWCjKkgG3RkOinT7TMSyyaURPmm8Ron6gyJSQPGsGF60uhk5x6OaA4u0qXThh3ZMpU0n+3fHZbD
anY5Vg2Gl0MhtSbxUnUkJAvl2gFwnGj17Bow/06eOApURO0Z8YnWj8VQs2mDnJekhLQfYJF5d2zC
87YD+11QxTVDsPBo/EhrQhkWpjj+Lsj5eSsFnsb4L/xsBvLIf4930cQHd7OLo2vymcY3stQ7ecA1
K5cZHuyE4oZ0Mv4R9fsVzmpgDzWLfnvlEdVZi8rxlalHIS0WWc8uGwOkR/2fc5Gp5KBDNIOKyDpz
38zu4i68GvfJkn9PPFO8KDpCaGj/8oqALCdiRkQWSyPovBg8fvp/Go2hecsdaDM6/Fr7aLDykdCe
l14y+fYwP2GAIb+WkRDhIqVBKlcoHlaiuDz3ymMTlzQOdrDxkrmaLSg/zPR4amMl9xm1lZ1rzb8Y
PwfB4SiXdoQdIXtsi03yqDsm1vqpQ0kI9KSVsL4UqYIKI1swhIEvjIW/f+xQAZSWzeyemiQ+6DlO
91sdpmvAaichiqJVN3i63Vj6OoX9Q6ymRWi5N9zvCdGxchzkdPHABc+Nr7uc9bC5mP+9Y/Bcy2BH
k0pFvXHjDQx2yc8GGKMLd97YSS5KVNW16eWKbv/elNZqECUOHfCsb+AqDzKItAkG7eJ5YbTHvU74
8FnEewbvZlj1Wve/mtLsKM2WBP5yAEb7aGrJHTNlGWJY55XNbuoydTXJ88sxp9fQVZTJadQE5nCM
6WfmBTjuUdX8T8d4phvvXswCnUJIyNBEZfQvC/YKOE/1Bmgh7XlF4imQuUvSdFCAgKowGh7Aw6zI
0xPIXT4eFDhGkBBqjtticGGs//4GT0/hSr9EDcpy2Ln+QgagGs0TycjoHD6GbtBhi0HC0lgQjNDW
GgNCW3LRqnSi1BQs7KYudq/2HbO/Q3kU1xAYTB/tSqkQ9Qb0T5/WDzjoJQK9pNfv9mODszf/KVaa
UHt7/o3MTtn8QQj0y6SIYJhmBh7Z8kWXBAK0vWa0MoeIGBL3FtCzLI2/RIzJTs3OdiUaHLgG7iLp
65PWiG+4ZkK/DuIkQpe2q665HsRMw435emRTF2LnaeW6JvtauHv6K7cmGUWS3a0u+Vg7X71bducA
kYqFhqDfS/SbVQizwnstBP1MH1lOs6wVRjNul2Xciae0Ke3z/6W28AI8gaRNhLdreszXuZgj6xDV
CAqKr0zFlEF13xaY8eFtkd/n1hRRKNgpp+LMOd2lOYxP+Ic9xjO1r1a4uRiHZZf7EBH4Qowuy9p5
ppUAigLDNvFavQXvvFI4h+bzNN0Q0WeHZE9diCzyqgWZQrCcrShEox5/9T8LrT2e2BXnS3HZoUC3
vZ0+3C7CqvKJCG+EwcUQ/22fcMsVOWRnV667h8iiHTcnQ3mpl6OvNMGMdNAUrdoBFt5uNv+42pu6
tpY2xTAYKtJgD+ooVqMHvVvjpt5qBsu8OO0LO7SsDcZxdyGUdQbtaMChopPElD/7Q0Vsq/4CbQvz
KNaoy5ncQCQsTzQQThU0xnXnR67Hyxu8twCoaksLp6tvcuYDWrukwuoAYt52JC+02UnQCZRgAm9n
8uWytDHe8CTq/+uKKRwDoRPYQdkj+XU/z+uQJ+8XKc63B1506x19Po2pBYRz40/IG1PmJ98WGa60
C1SEK9qPC+7oHTJ4xeaNeCfOKgJ6ay6/sxbTruvCMn9D5zSZYQrbnNiPI+6w9S1Dh7If/pEF6tjm
kg+iZgpsGBiVwHYB71eF4MY7YkssYrHWjUUmvja16VJUFSYcC+pA+J+JCUPNWiXjxVxDbekmouzM
dYHHS8GyUo321B1OywQUwZz0MT9880hVtaVcKcNFIUNMBn5PadiqX4blftC3WqAIU8G8Zj1I6E9E
ZYC9FpRpli31cnYdvjpqUKLIkKtTrUWfIQC395MQTDynXdshle7+hcg0onISWqhqq4L+gqTRgb1F
RsSOjIhAj1ElN3oNgtiqIXfE3Ha86ohwgf62vfp9sOFFixSc9sSzbcRyRNF86+aOprebiyEWVWrz
ENg9K46qRVbMbKzfm1vyIxKqCcE5BWpo1xTC9hYeiW5vLWBGc+GRV5+KIvabb5jSLF5KQwC2DfsY
xxdxvPPcYGnhxj9VapzSL71mAbKyF/jotTDPxwiuLuwQtGYpF0WHBBmFb+ZRYRhPdhoNklJxmKDB
ko6CQA7p+xvMEmwpUIxoxF7nqWsEYprdB7kQSxyyCp17Sr7s6BI62hvZuKZ4iqt26WNiZrm8XU9e
vjaGUxyEN6ykawscIPFnR8g4DufBVZLlNm3bNhCiQfbRc+V1UhnHuc5E5KRpQqatnr4vlW1QNsrp
tggCGfH/Tn4L+9ySNuBOAO6b33LVrciJzYaJe84U9s0okAUILpi8EzAm8L5vRa/snDoME6u+UJ/U
xVUc36vVAAX2gtkAH7YBhg6YrNoaPIr8NK2fWWEA7LR0hpDxpMfXaO/I4pF0/9DYVCcj2RissXUV
yc6xYH/Mnm5EpvHq4nZ55Y4ZuSpu52wpS5mpVzjHVWbOGgzcdVEOlZMRO1tRjRkrAFv16y8z4WDp
UHMpKRRPJ6JzMMg9Nk1SIbFHQ971btTnHre3VQ8vThdk9ol+1d/FpFCOaeQHspBbiJJ1uokwGgjX
ejqN/6AYVEvNdMEt8ekGd8VDsnCZ9BU8F0IOdKfCn6ecUNnJXXbuq4JzyERzunQ0DKA9vYyG3XeM
vx+nu29QEDnAig7fc5pd+wgjk7DSiAWZ8fihu/n8VmVDUB8VkmtoxHdsOciISA33pSfXBV5QkZcz
ohwDYcjfTrXNQ0FSCgatOaco1sK60RsKNfv8tepfn0rbiKmMHFdkgpMj/0JgQ1Zlm6LEdGxcw17y
c+GhU84gqFdeH6N2GmYmNBJ+rAuu3JJFix5kJxfebdFULOqN9relHtsynb3bUNe+nr9KpjwcFpYE
VOk/MTrsWOPgduiRkwswPlzEjxucmWt3s/J386cGhHIXcPuG+2zwbbH9yxANkptzFjcrYTV7KLYi
HKGtzbo2tA1h1VyTWOJUY5hjvigUvLiLjYxH6GZSC8WPoF4xZOIKRMqqDiEBkCu9BhO6Pqk+YXVC
zC5K20f2/vLwOaGx4i5E/mu6XMJXwtYyFshWHISsFsjSl070fF4DseSfgKBHMqJWEJ7ODQvDq2jy
whcd0M0kwaWMt32DC/n/htJSru5yP+m2QquI9scQI3odmVZQtogmAU3pM7rGMUKkj546SNWsqmQ8
d86S3j/4hb2G/Di0z7pmHSvaY869g0NRN98sVZTqo+LDC5oxEWwdz8R++d4eQ0ObXEiNBPkaocPf
SxQhWHx7U062dZmix1d+zgkv/xzo9z2oeRFlIxq6f5gzj2Drjoi35/Dfgj5fEo4vbORStnHSPk8S
+y/AQ0B81tFzv2G66zN235In0u7LN2Hu0HpJ9pe6lYVE0Bcqj4g/TOJ8qkrA2M502ZHdRNALqABC
2uEEq7eaKYA3DfpHrmxBhQt9b1XhihxlTjHZJ5GxU9t7iCyB2MWRmjsjJLVjDbtXrlBMOX/8LVZy
5xMX5JnM8kskUX5y75b7cJA2sO/C+1JzuFOLbJ3pajf4/YClnpeSRC5z+pd87W8pBDjwfJwISbb6
GjT5DVt9Bz3oAL2mp1I3ezUx44GKoqhuUhzaTypHPZsxEru4oau1HnORlLMyrhBn4u8o6Z9e6BCr
HtrhefFXmefFexKYhP2RL53PS7qH5TxngrlDgfN7f4LsDvaHs1Fu5Pj+2ow8GkZ9QkBUDheL1tgL
fMuO2TlQ0NDduVN0seLp7Qkgm7LSdhqgX2//wJC4gJ8YH62fT/PnJK78E+WoagXLEnStY8BdokZD
jaR3mau+aIEmOK780zhgrJEqEKG4khoC0HXoA8MmGaLibirx+xwcHs6AyMML6hFRkERkGDxOqvUU
HwU+uGMo9HKVC24Y0awwzLzxIlgPgcHqRxj8EOx6Rs3qYj+5pPzIYMxdyvE4FPT0eBFA03IpYSN6
Vu+uAdevsR+WW4O+uszIMt6jiHpsoYdhPk0niuvEcXKT04BfNSgstphe89I19wQSSSdi2vgmQcMA
1XcHmoTe9iCA+0MHqwUPbzxXgQogsohOaD2/aLi1r6asHRYOwjsa4sjxyysSKA72gezuybluUoki
DNgNbsKfw+/P/lKqyDL1YkiMiPyWSTrcow6FHIwQiUR8u/lNsg7O31PkWaPO0+r+6Azf3ZZH4XRc
J+ZOEx4Z16xbJnvbvekOrJAvVb0xOJJCJU+XDUjnCihchsTqlcS+f5FHoi5L/RN5eMr75NNV2r3e
XrbQhnPSp84aYVLnV8QKPj3xQw5IJk+apLxUtNFCj/c5627N09TyyJh7pFyaLYnwO8E9Y+DnTZV5
nVTzPJDaSNg5QPX2dsnilBdH+MkHIU5vw/NzcrUPlSQ4czVVD/Z3RgK1dlrGA/OT2gKqNtu6SKao
Eo+Rsqs5Q5tFQjCAUPE/vTukn+8fjmw9mHPl2VQga9vW0fEOVxoYJmD1waAdx0hvbsSetIa3+usX
KJz+FeFn0W9jdlcf5gPrSyk7GSSi8/vjNDfh1DWgOCdEwWu7pt4fK0uRTTgdgw8COQtVs4Ya5On9
b6qPONZi2F1rl9KaIqbXnMYLHdF0oH+0d/DOgxiJBqdkFWyVfearMk7a8EYV9ik4DX7OK6eP8rKI
uEe5zUKiDKe/mUobvnlxkO4KJG0ktwkA3vynCb17vdko2nUxb4hpTy0Z+RXxAb+QgCmCEmt7feOV
DbOyooj7LFs8oMk6a5pYiAecSW3cPliBf72hhtXpZoY7IWT51vu/iBgZknQTCjsFoGWkSCukw2sj
BETtJLftqyB9yF88OM+nk9AOFLK7nWHX7ZLWkMyoXlpfZl0bNLcig9jNf4akA/L1EVUxHRVCzj0i
FMs2FSUsEmnZYmLeVdRwuv/cx0oV65ciPNyLqJPeUsrkWkN0X2GToU/yuatzF14AOF5iw8B+C6r+
OaBqN4n9ZS94jpCULZTCSJDAncLhvhxxslfqJdngqN1KsLZGqnOUiloiZgFA8IC7nx6vniaHRnsR
Cza+sRh+7EYgq9ly6q7+eqw/U4djRW+NCGvjdyv8jzshiLUWStr19SO1yEy2Y5ncv3Xvj4BKeQ6D
t5gU0br+zW/FYGdI5J8nNnZzZ4GJvwG+J1EpzXCUdmm+jk+SsvvktQzTrrAeEe4pwe+VQdvDBYP7
zADLT0sQBQDvECFzNbZyrdrs4EiZEwASUrNhv3tBWz0el0Od42SEqh4L4x/7CuEXNdXzQ+4FN5lh
hy/fIMytEBOImkUDVQtZDGPUalUaTcBJJtbLK19mVGXpipeR6WuNGPo/eGk1uexkXnpJe/uKdVFD
7SaOvizyO2dXGzskTesT4NRJZQveLFV/m2bRj7bXCCsVRxn7+U6zwGW9dwFW9npM6GCt4GNEKN6Z
H1w39Ha5xCQETume2t59h8HcfcfW4FkLvzSgSIYoRglGWFoa/GfBSlMTJGz65oA5j9Sp6wfaEOVz
UhpnV4KMCJf0HXJjvtX4UPj6YWHi3osJu87r/lP97zESH3YtoIdiXH6T1W5dWr/+guakJmHol3Ym
UvPgtniybx2P8GAnyiu+0BUXc6ryLFUiKlpoBt+0TRvze3Sefp0orbxiYQwL/oweBcC/fYreyCjH
kc06/C4W/q6Aizqo90XHZoTS6HqOBi3boDynYZcfwrD5EOMQ/uoA5KcLZOvzUdFdEUrv+BLtw14C
3LtxBI1gGu3WTlI4muS9XyyZEABa6hb7pFr7SqgCs+cGfFzsM8WaVrOijVdnIo5HlrLFc1IHTzbT
blQeQ8etSKxHDMWOsdpIEvELlEDAb6l5+vcEVkutbM03gb9Nugr4BBLX71FISO9pPpsIA0XHt0Bw
PPizRcQJF3HF+0vqjru5RjmTe6z7lW5W+5ZKgr6s2s40VQvhk3MvgRucDkJLj2nqqDknsvYvzd31
ibwwo6DqDNZ1au+t9LR6esnMiU9gt5gM1RVO+k1YIpbk4ClrN2fNZaczC2rKwtr6+p3cmozPYKXY
JP8vOBi0nRneheArQMamqwjkKZDM6cXiTfmQyP+7SI7SMfXrH6jDYwvJNl5U3abUVduCdLyVTERp
pPWwLxRa10EiWzUKwWQzl5Ebb+EcDZB3c43yZFJzDecKlzGjVQAjje0Q3zjzol6oNIhP+QwBioQW
p8wG8R4wPD0WQgE/qiuqOJpw3re2WwgVde07hsGxktEXsNzmm5wNidQuDKrznTs1KsYAW7a6sOk+
VLBi+1gBw5GRs9yizQbVRQ1sB6SFPXInNoIE05OUsJ/SfoU5ez74xYfo8KCVHTOtSEFeXAnqqWX6
q+kN517SNJJvP1e942HQgZ9o4BLqU6cWO1jeaPBo0D+ouvJYH54cf4Rq5EVA5WgCTz+VbZVAigA6
L7jS2Zwwn1cUx08EoNH16PVQww0Xpm7X2y5SqYUs8FSb4rluP8g/r84Y20DlGc4eOqtTKmIufCyK
gCI+bKXFApq+Jwh/WrIuvr4I7VBvXVkiAfKMSJvfSY3mDoVzOdZwzkKqmeh/Yi+v3V/n559eHnRl
Yy3goTljMsSJ0u0yqmfLaRDjxjSxB3Klu6v/tBGJqH4paKK+KkeRXibkol5WHnAGjQ+8lmz2iCKk
EH9jwCqT1y/jN61L/ZIDH0ajz16UAC4geQGYSUrtQsZC/VanokF3wtvnQSbZhLFsV0RQQRlGi5lO
E3cTLRKSgs5iCw86dkcbLL+P+O9Eg22gNR+w6VVq2ef1I0x/1cjHPxhVEPrW5NSCyyv1zc4rYqCq
j572T4Njvf7qkREZEQ6LdnwS/Y4BmxhfM3JI37lBF0uZbGnu6E9kZ4k1gxJLoPbIsegkrZZZtAUJ
GkalMaS5xt+i0giFgSW5iC4M9H7sa+wR37Z5eS9bcYyYIyGyNxWxCA+ZFzbuWaXhviq+Z8mUgzEW
biDdOjSWS9qdnn7nYW0ngXsHq36DiKIq/DRlg7DH9ioC9igCvgzpNmd++2sx/Espm3SMczwhCY4C
CmByjVG9jVhpB+hAwv/DQezFUu1NFDSJeBroCwB4NySACTfd76XZCB6P72+7ff+ClZOS5t2XaMZX
oSd7a4PTI6KRmvkktVvX4k5zE/pwHBZ5aJfCHNSDYLS7BR2JByotzNsxqleeRlWILqZU84W4Nhq8
wnhYkj6ZJYbdBmG5TAJ04BDaEpO4hFlZ867bPoSTAqdKAIWZumS5GrG+XfJZ3nTbX4YRX8m7Wudf
HhdBk98dbb4oSbDHj2vyoaI4yQtlDFlFpAEaL9VcwB4TFqGEkocOw1FlaqiTzoaLsMoSGYKyQnDT
wGc0ihgVVaZTiPKDBMacc2wDZIsIsnSpNyvVfHgQRnhbB46j5TFdHaZt9fzGc1W/swqmwHRcRRoi
4ponrOVR4jT+xJS6mcnT39Qch482lGilhrzwhvnaiTMoEYK+f8/aI2Sze83+3I4gd+2aJ+RR92xT
W0Jhp6p8Ah0m/A/E+xWp95FOVwly2iZYF8cbggOPRzTt7Dp20GQVtLywJ31b0fGJMwp0lvmZ8cZ1
Sv3AQiHURtcf51F4V46TA8zVikV0oTIUATOu2GElAPZWzsWjA91q4V4aM5uYjvzyqhs9/t/0bqHq
i748siAcI3oj/cSWMdG2BqftXJfz+fqS6c3e9q/o+cWwbBzFVJHuDyuZbMj2m3Iwn/vTMP8tEQ07
oZdzm0oI7iWObzSvwNyEPZ7KwYHGVfFeXAyvteEaj8g6gyKXke8crhbd8f+aixK79s0DRgP0ZzuQ
toW54Sy+2wNO2mdoa2uxPxNcDWrBCXYuWZFpKf9As5UcMbkrTU/FtpUjLryk1MT7xhDPV5OPSkhs
3c/MEvVEKU7J53wwZKgN56PLLTvmRLOK1Jgvm7CQInbtDg2gdCPlQEnhf5MXy6V+waWCW6E54KsZ
I1ReGv83to2mZklOwQmBtjJpE3abQFDqtFlEguZL+3AUPydFwm4kUoG5AzbwuLyKma/MtXfLF/IE
f2Lma0IX+uLAjKu+uM3P4perqZYVvdiO89z1FhswQlHKNpBmLb8diZG1euqF7UtsTxtEqf1l5KGt
kYzva6U+gl8PGXfw/6e+HK/TaPZuy15n2SdO+/W+DQTxJane32QRcuZLUL8dAX/fXfQwnDc464SH
WU6h7BxyXb9TMM0Yu02dJgEbP25NEn6o1vtNbewE/DtP6a1fGLRx4B6TBnYC3zmcQ4SCycSCGAtg
xEr1Sfz09NosWtAuCp9HFjuX7k08ImZPxNtNIqci5cIbl9fOGgKBVqwWW0quVWvRO0dw+DiHKbm6
jcz3YYeqEhGuaYroa8WfYAlPD6l0AKbMo/xJaD4OZkyKrrxtSSDLYkG8LPz3of0249d4m03NmpnX
7kPgMlOZnBhAayagAJQaU94GjRD7PkRevpidkK7Q91UL90i7/+UWsZwC8F1/Xal1K07jAKUNL5Xo
N/naVvnA9yblHaR1mLC0D7ie8p1zgNI7z+2+z2aXkBTdZi7ymrClKuFth4lIXk+sjd19GuBbm5EY
DK73jyjZClrk0yqzYx9pQvmPeYFWfbfVEQ3xzv1f7yFBf1i5a9qPRpNPLg/ZCQDI71qXh1Pb3G4F
cOt7kcT+dmbK+833S2rzCcMhH+PBvFVa5VPS0vv58WVGhZ/0NjBRc7+SdtP3wktNc+OsyDRQvk4Z
LF+lg0embL6ROjVqj1H2HT4qJTnmqimixRnLpJp16vWkNeUgwBF+c1ruGrJYXhWOfPgt6i4+C6WJ
YtZc2uvpVBtICGh4qf42iis3zs3kGTFfPMIsbT1hcmMK/wrjgwBGX2l1TIKh7e+e80wkTDvqfpxC
z4uj49nCUKtwYUspI0ssF/K9rurityggoJr1ECjIMBF/WRNipLjqBV6Hs5H560yLMgMZ/0Noki48
R4skP5v1NpdfqFS0jp/Eug/ezCpgrLDQwgjwtHcr65U80mQSjfNXp2VBGtiy
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity keyboardFifo is
port(
  Data :  in std_logic_vector(31 downto 0);
  WrClk :  in std_logic;
  RdClk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Q :  out std_logic_vector(31 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end keyboardFifo;
architecture beh of keyboardFifo is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo.keyboardFifo\
port(
  RdClk: in std_logic;
  WrClk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  RdEn: in std_logic;
  WrEn: in std_logic;
  Data : in std_logic_vector(31 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_inst: \~fifo.keyboardFifo\
port map(
  RdClk => RdClk,
  WrClk => WrClk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  RdEn => RdEn,
  WrEn => WrEn,
  Data(31 downto 0) => Data(31 downto 0),
  Empty => NN,
  Full => NN_0,
  Q(31 downto 0) => Q(31 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
